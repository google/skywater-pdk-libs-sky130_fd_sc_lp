* File: sky130_fd_sc_lp__sdfrtp_4.pxi.spice
* Created: Fri Aug 28 11:28:36 2020
* 
x_PM_SKY130_FD_SC_LP__SDFRTP_4%A_27_74# N_A_27_74#_M1000_s N_A_27_74#_M1002_s
+ N_A_27_74#_M1021_g N_A_27_74#_M1020_g N_A_27_74#_c_323_p N_A_27_74#_c_309_n
+ N_A_27_74#_c_310_n N_A_27_74#_c_311_n N_A_27_74#_c_316_n N_A_27_74#_c_317_n
+ N_A_27_74#_c_318_n N_A_27_74#_c_319_n N_A_27_74#_c_312_n N_A_27_74#_c_320_n
+ N_A_27_74#_c_321_n N_A_27_74#_c_322_n N_A_27_74#_c_313_n
+ PM_SKY130_FD_SC_LP__SDFRTP_4%A_27_74#
x_PM_SKY130_FD_SC_LP__SDFRTP_4%SCE N_SCE_M1000_g N_SCE_c_396_n N_SCE_c_397_n
+ N_SCE_c_398_n N_SCE_c_399_n N_SCE_M1002_g N_SCE_c_400_n N_SCE_c_401_n
+ N_SCE_M1035_g N_SCE_M1029_g N_SCE_c_402_n N_SCE_c_416_n N_SCE_c_393_n SCE SCE
+ SCE SCE N_SCE_c_395_n PM_SKY130_FD_SC_LP__SDFRTP_4%SCE
x_PM_SKY130_FD_SC_LP__SDFRTP_4%D N_D_M1023_g N_D_c_476_n N_D_M1038_g D D D
+ N_D_c_475_n PM_SKY130_FD_SC_LP__SDFRTP_4%D
x_PM_SKY130_FD_SC_LP__SDFRTP_4%SCD N_SCD_M1032_g N_SCD_c_518_n N_SCD_c_519_n
+ N_SCD_M1012_g N_SCD_c_523_n SCD SCD N_SCD_c_520_n N_SCD_c_521_n
+ PM_SKY130_FD_SC_LP__SDFRTP_4%SCD
x_PM_SKY130_FD_SC_LP__SDFRTP_4%A_851_242# N_A_851_242#_M1031_s
+ N_A_851_242#_M1004_s N_A_851_242#_M1017_g N_A_851_242#_M1024_g
+ N_A_851_242#_c_565_n N_A_851_242#_M1019_g N_A_851_242#_c_566_n
+ N_A_851_242#_c_567_n N_A_851_242#_M1013_g N_A_851_242#_c_586_n
+ N_A_851_242#_c_568_n N_A_851_242#_c_569_n N_A_851_242#_c_588_n
+ N_A_851_242#_c_589_n N_A_851_242#_c_570_n N_A_851_242#_c_571_n
+ N_A_851_242#_c_572_n N_A_851_242#_c_573_n N_A_851_242#_c_574_n
+ N_A_851_242#_c_575_n N_A_851_242#_c_576_n N_A_851_242#_c_577_n
+ N_A_851_242#_c_578_n N_A_851_242#_c_579_n N_A_851_242#_c_580_n
+ N_A_851_242#_c_581_n N_A_851_242#_c_598_p N_A_851_242#_c_582_n
+ N_A_851_242#_c_583_n PM_SKY130_FD_SC_LP__SDFRTP_4%A_851_242#
x_PM_SKY130_FD_SC_LP__SDFRTP_4%A_1047_369# N_A_1047_369#_M1015_d
+ N_A_1047_369#_M1022_d N_A_1047_369#_M1003_g N_A_1047_369#_c_785_n
+ N_A_1047_369#_c_786_n N_A_1047_369#_M1045_g N_A_1047_369#_c_780_n
+ N_A_1047_369#_c_781_n N_A_1047_369#_c_789_n N_A_1047_369#_c_790_n
+ N_A_1047_369#_c_782_n N_A_1047_369#_c_783_n N_A_1047_369#_c_812_n
+ PM_SKY130_FD_SC_LP__SDFRTP_4%A_1047_369#
x_PM_SKY130_FD_SC_LP__SDFRTP_4%RESET_B N_RESET_B_M1001_g N_RESET_B_c_882_n
+ N_RESET_B_c_883_n N_RESET_B_M1033_g N_RESET_B_c_885_n N_RESET_B_c_890_n
+ N_RESET_B_M1009_g N_RESET_B_c_891_n N_RESET_B_c_892_n N_RESET_B_M1036_g
+ N_RESET_B_M1026_g N_RESET_B_M1018_g N_RESET_B_c_888_n N_RESET_B_c_896_n
+ N_RESET_B_c_897_n N_RESET_B_c_898_n N_RESET_B_c_937_n N_RESET_B_c_899_n
+ N_RESET_B_c_900_n N_RESET_B_c_901_n N_RESET_B_c_902_n N_RESET_B_c_903_n
+ N_RESET_B_c_904_n RESET_B N_RESET_B_c_905_n N_RESET_B_c_906_n
+ PM_SKY130_FD_SC_LP__SDFRTP_4%RESET_B
x_PM_SKY130_FD_SC_LP__SDFRTP_4%A_881_463# N_A_881_463#_M1030_d
+ N_A_881_463#_M1017_d N_A_881_463#_M1009_d N_A_881_463#_M1015_g
+ N_A_881_463#_M1022_g N_A_881_463#_c_1068_n N_A_881_463#_c_1077_n
+ N_A_881_463#_c_1069_n N_A_881_463#_c_1095_n N_A_881_463#_c_1161_n
+ N_A_881_463#_c_1070_n N_A_881_463#_c_1071_n N_A_881_463#_c_1072_n
+ N_A_881_463#_c_1078_n N_A_881_463#_c_1073_n N_A_881_463#_c_1074_n
+ PM_SKY130_FD_SC_LP__SDFRTP_4%A_881_463#
x_PM_SKY130_FD_SC_LP__SDFRTP_4%A_975_255# N_A_975_255#_M1011_d
+ N_A_975_255#_M1037_d N_A_975_255#_M1007_g N_A_975_255#_M1030_g
+ N_A_975_255#_c_1223_n N_A_975_255#_c_1224_n N_A_975_255#_M1010_g
+ N_A_975_255#_c_1209_n N_A_975_255#_M1006_g N_A_975_255#_M1031_g
+ N_A_975_255#_M1004_g N_A_975_255#_c_1212_n N_A_975_255#_c_1213_n
+ N_A_975_255#_c_1229_n N_A_975_255#_c_1230_n N_A_975_255#_c_1231_n
+ N_A_975_255#_c_1214_n N_A_975_255#_c_1232_n N_A_975_255#_c_1215_n
+ N_A_975_255#_c_1216_n N_A_975_255#_c_1217_n N_A_975_255#_c_1218_n
+ N_A_975_255#_c_1219_n N_A_975_255#_c_1220_n N_A_975_255#_c_1221_n
+ N_A_975_255#_c_1366_p N_A_975_255#_c_1237_n N_A_975_255#_c_1238_n
+ PM_SKY130_FD_SC_LP__SDFRTP_4%A_975_255#
x_PM_SKY130_FD_SC_LP__SDFRTP_4%A_1524_69# N_A_1524_69#_M1019_d
+ N_A_1524_69#_M1010_d N_A_1524_69#_M1016_g N_A_1524_69#_M1042_g
+ N_A_1524_69#_M1041_g N_A_1524_69#_M1044_g N_A_1524_69#_c_1412_n
+ N_A_1524_69#_c_1413_n N_A_1524_69#_c_1447_n N_A_1524_69#_c_1414_n
+ N_A_1524_69#_c_1432_n N_A_1524_69#_c_1415_n N_A_1524_69#_c_1416_n
+ N_A_1524_69#_c_1417_n N_A_1524_69#_c_1418_n N_A_1524_69#_c_1419_n
+ N_A_1524_69#_c_1420_n N_A_1524_69#_c_1421_n N_A_1524_69#_c_1422_n
+ N_A_1524_69#_c_1423_n N_A_1524_69#_c_1424_n N_A_1524_69#_c_1425_n
+ N_A_1524_69#_c_1426_n N_A_1524_69#_c_1427_n N_A_1524_69#_c_1428_n
+ PM_SKY130_FD_SC_LP__SDFRTP_4%A_1524_69#
x_PM_SKY130_FD_SC_LP__SDFRTP_4%A_1747_21# N_A_1747_21#_M1016_d
+ N_A_1747_21#_M1018_d N_A_1747_21#_M1039_g N_A_1747_21#_M1028_g
+ N_A_1747_21#_c_1596_n N_A_1747_21#_c_1597_n N_A_1747_21#_c_1598_n
+ N_A_1747_21#_c_1599_n N_A_1747_21#_c_1606_n N_A_1747_21#_c_1632_n
+ N_A_1747_21#_c_1600_n N_A_1747_21#_c_1607_n N_A_1747_21#_c_1601_n
+ N_A_1747_21#_c_1602_n N_A_1747_21#_c_1608_n N_A_1747_21#_c_1609_n
+ N_A_1747_21#_c_1603_n PM_SKY130_FD_SC_LP__SDFRTP_4%A_1747_21#
x_PM_SKY130_FD_SC_LP__SDFRTP_4%CLK N_CLK_M1011_g N_CLK_M1037_g N_CLK_c_1708_n
+ N_CLK_c_1709_n CLK CLK CLK N_CLK_c_1710_n N_CLK_c_1711_n
+ PM_SKY130_FD_SC_LP__SDFRTP_4%CLK
x_PM_SKY130_FD_SC_LP__SDFRTP_4%A_2555_47# N_A_2555_47#_M1041_s
+ N_A_2555_47#_M1044_s N_A_2555_47#_M1014_g N_A_2555_47#_M1005_g
+ N_A_2555_47#_M1027_g N_A_2555_47#_M1008_g N_A_2555_47#_M1040_g
+ N_A_2555_47#_M1025_g N_A_2555_47#_M1043_g N_A_2555_47#_M1034_g
+ N_A_2555_47#_c_1766_n N_A_2555_47#_c_1776_n N_A_2555_47#_c_1785_n
+ N_A_2555_47#_c_1767_n N_A_2555_47#_c_1777_n N_A_2555_47#_c_1778_n
+ N_A_2555_47#_c_1768_n N_A_2555_47#_c_1769_n N_A_2555_47#_c_1809_p
+ N_A_2555_47#_c_1770_n N_A_2555_47#_c_1771_n
+ PM_SKY130_FD_SC_LP__SDFRTP_4%A_2555_47#
x_PM_SKY130_FD_SC_LP__SDFRTP_4%VPWR N_VPWR_M1002_d N_VPWR_M1012_d N_VPWR_M1003_d
+ N_VPWR_M1022_s N_VPWR_M1028_d N_VPWR_M1042_d N_VPWR_M1004_d N_VPWR_M1044_d
+ N_VPWR_M1008_s N_VPWR_M1034_s N_VPWR_c_1877_n N_VPWR_c_1878_n N_VPWR_c_1879_n
+ N_VPWR_c_1880_n N_VPWR_c_1881_n N_VPWR_c_1882_n N_VPWR_c_1976_n
+ N_VPWR_c_1883_n N_VPWR_c_1979_n N_VPWR_c_1884_n N_VPWR_c_1885_n
+ N_VPWR_c_1886_n N_VPWR_c_1887_n N_VPWR_c_1888_n N_VPWR_c_1889_n VPWR
+ N_VPWR_c_1890_n N_VPWR_c_1891_n N_VPWR_c_1892_n N_VPWR_c_1893_n
+ N_VPWR_c_1894_n N_VPWR_c_1895_n N_VPWR_c_1896_n N_VPWR_c_1897_n
+ N_VPWR_c_1898_n N_VPWR_c_1899_n N_VPWR_c_1900_n N_VPWR_c_1901_n
+ N_VPWR_c_1902_n N_VPWR_c_1903_n N_VPWR_c_1904_n N_VPWR_c_1905_n
+ N_VPWR_c_1906_n N_VPWR_c_1876_n PM_SKY130_FD_SC_LP__SDFRTP_4%VPWR
x_PM_SKY130_FD_SC_LP__SDFRTP_4%A_372_50# N_A_372_50#_M1023_d N_A_372_50#_M1030_s
+ N_A_372_50#_M1038_d N_A_372_50#_M1033_d N_A_372_50#_c_2064_n
+ N_A_372_50#_c_2057_n N_A_372_50#_c_2058_n N_A_372_50#_c_2059_n
+ N_A_372_50#_c_2060_n N_A_372_50#_c_2066_n N_A_372_50#_c_2061_n
+ N_A_372_50#_c_2062_n N_A_372_50#_c_2063_n N_A_372_50#_c_2067_n
+ PM_SKY130_FD_SC_LP__SDFRTP_4%A_372_50#
x_PM_SKY130_FD_SC_LP__SDFRTP_4%Q N_Q_M1014_s N_Q_M1040_s N_Q_M1005_d N_Q_M1025_d
+ N_Q_c_2203_p N_Q_c_2157_n N_Q_c_2191_n N_Q_c_2152_n N_Q_c_2153_n N_Q_c_2158_n
+ N_Q_c_2195_n N_Q_c_2159_n N_Q_c_2154_n N_Q_c_2155_n N_Q_c_2156_n N_Q_c_2161_n
+ Q N_Q_c_2204_p PM_SKY130_FD_SC_LP__SDFRTP_4%Q
x_PM_SKY130_FD_SC_LP__SDFRTP_4%VGND N_VGND_M1000_d N_VGND_M1001_d N_VGND_M1036_d
+ N_VGND_M1039_d N_VGND_M1031_d N_VGND_M1041_d N_VGND_M1027_d N_VGND_M1043_d
+ N_VGND_c_2209_n N_VGND_c_2210_n N_VGND_c_2211_n N_VGND_c_2212_n
+ N_VGND_c_2213_n N_VGND_c_2214_n N_VGND_c_2215_n N_VGND_c_2216_n
+ N_VGND_c_2217_n N_VGND_c_2218_n N_VGND_c_2219_n N_VGND_c_2220_n VGND
+ N_VGND_c_2221_n N_VGND_c_2222_n N_VGND_c_2223_n N_VGND_c_2224_n
+ N_VGND_c_2225_n N_VGND_c_2226_n N_VGND_c_2227_n N_VGND_c_2228_n
+ N_VGND_c_2229_n N_VGND_c_2230_n N_VGND_c_2231_n N_VGND_c_2232_n
+ N_VGND_c_2233_n PM_SKY130_FD_SC_LP__SDFRTP_4%VGND
x_PM_SKY130_FD_SC_LP__SDFRTP_4%noxref_24 N_noxref_24_M1021_s N_noxref_24_M1032_d
+ N_noxref_24_c_2367_n N_noxref_24_c_2368_n N_noxref_24_c_2369_n
+ PM_SKY130_FD_SC_LP__SDFRTP_4%noxref_24
cc_1 VNB N_A_27_74#_c_309_n 0.0303728f $X=-0.19 $Y=-0.245 $X2=0.267 $Y2=1.93
cc_2 VNB N_A_27_74#_c_310_n 0.0170886f $X=-0.19 $Y=-0.245 $X2=1.335 $Y2=0.945
cc_3 VNB N_A_27_74#_c_311_n 0.0360573f $X=-0.19 $Y=-0.245 $X2=1.335 $Y2=0.945
cc_4 VNB N_A_27_74#_c_312_n 0.010626f $X=-0.19 $Y=-0.245 $X2=0.267 $Y2=0.912
cc_5 VNB N_A_27_74#_c_313_n 0.0216212f $X=-0.19 $Y=-0.245 $X2=1.335 $Y2=0.78
cc_6 VNB N_SCE_M1000_g 0.0397638f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_SCE_M1029_g 0.0261891f $X=-0.19 $Y=-0.245 $X2=0.267 $Y2=1.93
cc_8 VNB N_SCE_c_393_n 0.0671492f $X=-0.19 $Y=-0.245 $X2=1.3 $Y2=2.275
cc_9 VNB SCE 0.0326712f $X=-0.19 $Y=-0.245 $X2=2.605 $Y2=2.027
cc_10 VNB N_SCE_c_395_n 0.0394595f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_D_M1023_g 0.0666232f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB D 0.0120694f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_D_c_475_n 0.0197933f $X=-0.19 $Y=-0.245 $X2=0.267 $Y2=1.03
cc_14 VNB N_SCD_M1032_g 0.0376276f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_SCD_c_518_n 0.0352528f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_SCD_c_519_n 0.00747201f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_SCD_c_520_n 0.0174565f $X=-0.19 $Y=-0.245 $X2=0.267 $Y2=1.93
cc_18 VNB N_SCD_c_521_n 0.012027f $X=-0.19 $Y=-0.245 $X2=0.38 $Y2=0.912
cc_19 VNB N_A_851_242#_c_565_n 0.0236663f $X=-0.19 $Y=-0.245 $X2=0.255 $Y2=0.795
cc_20 VNB N_A_851_242#_c_566_n 0.012171f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_851_242#_c_567_n 0.00969086f $X=-0.19 $Y=-0.245 $X2=0.267 $Y2=1.03
cc_22 VNB N_A_851_242#_c_568_n 0.00509852f $X=-0.19 $Y=-0.245 $X2=0.38 $Y2=2.102
cc_23 VNB N_A_851_242#_c_569_n 0.00435388f $X=-0.19 $Y=-0.245 $X2=1.3 $Y2=2.275
cc_24 VNB N_A_851_242#_c_570_n 0.00213752f $X=-0.19 $Y=-0.245 $X2=2.77 $Y2=1.935
cc_25 VNB N_A_851_242#_c_571_n 0.0070315f $X=-0.19 $Y=-0.245 $X2=2.73 $Y2=2.027
cc_26 VNB N_A_851_242#_c_572_n 0.00262319f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_851_242#_c_573_n 0.014382f $X=-0.19 $Y=-0.245 $X2=1.335 $Y2=0.945
cc_28 VNB N_A_851_242#_c_574_n 0.001144f $X=-0.19 $Y=-0.245 $X2=1.335 $Y2=0.78
cc_29 VNB N_A_851_242#_c_575_n 0.0142281f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_851_242#_c_576_n 7.38858e-19 $X=-0.19 $Y=-0.245 $X2=2.77 $Y2=1.935
cc_31 VNB N_A_851_242#_c_577_n 0.00330352f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_851_242#_c_578_n 0.00545072f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_851_242#_c_579_n 0.011552f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_851_242#_c_580_n 0.0474813f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_851_242#_c_581_n 0.0303231f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_851_242#_c_582_n 0.0158251f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_851_242#_c_583_n 0.0339641f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_1047_369#_M1045_g 0.0429192f $X=-0.19 $Y=-0.245 $X2=0.255 $Y2=0.58
cc_39 VNB N_A_1047_369#_c_780_n 0.0064922f $X=-0.19 $Y=-0.245 $X2=1.335
+ $Y2=0.945
cc_40 VNB N_A_1047_369#_c_781_n 0.0122587f $X=-0.19 $Y=-0.245 $X2=0.38 $Y2=2.102
cc_41 VNB N_A_1047_369#_c_782_n 2.67424e-19 $X=-0.19 $Y=-0.245 $X2=2.605
+ $Y2=2.027
cc_42 VNB N_A_1047_369#_c_783_n 8.6638e-19 $X=-0.19 $Y=-0.245 $X2=1.45 $Y2=2.027
cc_43 VNB N_RESET_B_M1001_g 0.0170581f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_RESET_B_c_882_n 0.0263412f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_RESET_B_c_883_n 0.012806f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_RESET_B_M1033_g 0.0997745f $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=0.46
cc_47 VNB N_RESET_B_c_885_n 0.183923f $X=-0.19 $Y=-0.245 $X2=2.75 $Y2=2.635
cc_48 VNB N_RESET_B_M1036_g 0.055192f $X=-0.19 $Y=-0.245 $X2=1.335 $Y2=0.912
cc_49 VNB N_RESET_B_M1026_g 0.0396359f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_RESET_B_c_888_n 0.00749069f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_881_463#_M1015_g 0.0227069f $X=-0.19 $Y=-0.245 $X2=2.75 $Y2=2.635
cc_52 VNB N_A_881_463#_M1022_g 0.0141749f $X=-0.19 $Y=-0.245 $X2=0.26 $Y2=0.58
cc_53 VNB N_A_881_463#_c_1068_n 0.00173856f $X=-0.19 $Y=-0.245 $X2=0.267
+ $Y2=1.93
cc_54 VNB N_A_881_463#_c_1069_n 0.00161563f $X=-0.19 $Y=-0.245 $X2=1.335
+ $Y2=0.945
cc_55 VNB N_A_881_463#_c_1070_n 0.00117261f $X=-0.19 $Y=-0.245 $X2=1.315
+ $Y2=2.46
cc_56 VNB N_A_881_463#_c_1071_n 0.0014127f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_881_463#_c_1072_n 0.0149461f $X=-0.19 $Y=-0.245 $X2=1.45 $Y2=2.027
cc_58 VNB N_A_881_463#_c_1073_n 0.0088511f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_881_463#_c_1074_n 0.0582437f $X=-0.19 $Y=-0.245 $X2=2.77 $Y2=2.1
cc_60 VNB N_A_975_255#_M1007_g 0.0159424f $X=-0.19 $Y=-0.245 $X2=2.75 $Y2=2.1
cc_61 VNB N_A_975_255#_M1030_g 0.0287825f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_A_975_255#_c_1209_n 0.00362284f $X=-0.19 $Y=-0.245 $X2=1.335
+ $Y2=0.945
cc_63 VNB N_A_975_255#_M1006_g 0.0411279f $X=-0.19 $Y=-0.245 $X2=1.15 $Y2=2.102
cc_64 VNB N_A_975_255#_M1031_g 0.0236269f $X=-0.19 $Y=-0.245 $X2=1.315 $Y2=2.46
cc_65 VNB N_A_975_255#_c_1212_n 0.013701f $X=-0.19 $Y=-0.245 $X2=2.77 $Y2=1.935
cc_66 VNB N_A_975_255#_c_1213_n 0.00991328f $X=-0.19 $Y=-0.245 $X2=2.73
+ $Y2=2.027
cc_67 VNB N_A_975_255#_c_1214_n 0.00219262f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_A_975_255#_c_1215_n 0.00501326f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_975_255#_c_1216_n 0.00185708f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_A_975_255#_c_1217_n 0.019482f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_A_975_255#_c_1218_n 7.18436e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_A_975_255#_c_1219_n 0.0305903f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_A_975_255#_c_1220_n 0.00231989f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_A_975_255#_c_1221_n 0.00468421f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_A_1524_69#_M1042_g 0.0130706f $X=-0.19 $Y=-0.245 $X2=2.75 $Y2=2.635
cc_76 VNB N_A_1524_69#_M1044_g 0.00836612f $X=-0.19 $Y=-0.245 $X2=0.267 $Y2=1.93
cc_77 VNB N_A_1524_69#_c_1412_n 0.00877012f $X=-0.19 $Y=-0.245 $X2=1.335
+ $Y2=0.945
cc_78 VNB N_A_1524_69#_c_1413_n 0.0107016f $X=-0.19 $Y=-0.245 $X2=1.335
+ $Y2=0.945
cc_79 VNB N_A_1524_69#_c_1414_n 0.00366019f $X=-0.19 $Y=-0.245 $X2=1.315
+ $Y2=2.46
cc_80 VNB N_A_1524_69#_c_1415_n 0.00267182f $X=-0.19 $Y=-0.245 $X2=1.3 $Y2=2.102
cc_81 VNB N_A_1524_69#_c_1416_n 0.00166888f $X=-0.19 $Y=-0.245 $X2=2.77
+ $Y2=1.935
cc_82 VNB N_A_1524_69#_c_1417_n 0.00910172f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_A_1524_69#_c_1418_n 0.0171805f $X=-0.19 $Y=-0.245 $X2=2.73 $Y2=2.027
cc_84 VNB N_A_1524_69#_c_1419_n 0.00311855f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_A_1524_69#_c_1420_n 0.0103873f $X=-0.19 $Y=-0.245 $X2=1.335 $Y2=0.78
cc_86 VNB N_A_1524_69#_c_1421_n 0.0229622f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_A_1524_69#_c_1422_n 0.00353514f $X=-0.19 $Y=-0.245 $X2=2.77
+ $Y2=1.935
cc_88 VNB N_A_1524_69#_c_1423_n 0.034375f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_A_1524_69#_c_1424_n 0.0151314f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_A_1524_69#_c_1425_n 0.016831f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_A_1524_69#_c_1426_n 0.0394704f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_A_1524_69#_c_1427_n 0.0161629f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_93 VNB N_A_1524_69#_c_1428_n 0.0201381f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_94 VNB N_A_1747_21#_M1039_g 0.0242554f $X=-0.19 $Y=-0.245 $X2=2.75 $Y2=2.1
cc_95 VNB N_A_1747_21#_c_1596_n 0.100912f $X=-0.19 $Y=-0.245 $X2=0.255 $Y2=0.58
cc_96 VNB N_A_1747_21#_c_1597_n 0.012806f $X=-0.19 $Y=-0.245 $X2=0.26 $Y2=0.58
cc_97 VNB N_A_1747_21#_c_1598_n 0.0177048f $X=-0.19 $Y=-0.245 $X2=0.267 $Y2=1.03
cc_98 VNB N_A_1747_21#_c_1599_n 0.0249664f $X=-0.19 $Y=-0.245 $X2=1.335
+ $Y2=0.912
cc_99 VNB N_A_1747_21#_c_1600_n 0.0081825f $X=-0.19 $Y=-0.245 $X2=2.605
+ $Y2=2.027
cc_100 VNB N_A_1747_21#_c_1601_n 0.00349984f $X=-0.19 $Y=-0.245 $X2=2.73
+ $Y2=1.935
cc_101 VNB N_A_1747_21#_c_1602_n 0.0063686f $X=-0.19 $Y=-0.245 $X2=2.77
+ $Y2=1.935
cc_102 VNB N_A_1747_21#_c_1603_n 0.0506059f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_103 VNB N_CLK_M1011_g 0.034515f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_104 VNB N_CLK_M1037_g 0.00217083f $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=0.78
cc_105 VNB N_CLK_c_1708_n 0.0470028f $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=0.46
cc_106 VNB N_CLK_c_1709_n 0.00464418f $X=-0.19 $Y=-0.245 $X2=2.75 $Y2=2.635
cc_107 VNB N_CLK_c_1710_n 0.00350064f $X=-0.19 $Y=-0.245 $X2=0.38 $Y2=0.912
cc_108 VNB N_CLK_c_1711_n 3.00037e-19 $X=-0.19 $Y=-0.245 $X2=1.335 $Y2=0.912
cc_109 VNB N_A_2555_47#_M1014_g 0.0215698f $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=0.46
cc_110 VNB N_A_2555_47#_M1005_g 4.20731e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_111 VNB N_A_2555_47#_M1027_g 0.0213234f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_112 VNB N_A_2555_47#_M1008_g 4.71631e-19 $X=-0.19 $Y=-0.245 $X2=1.335
+ $Y2=0.912
cc_113 VNB N_A_2555_47#_M1040_g 0.021894f $X=-0.19 $Y=-0.245 $X2=1.15 $Y2=2.102
cc_114 VNB N_A_2555_47#_M1025_g 4.7181e-19 $X=-0.19 $Y=-0.245 $X2=1.315 $Y2=2.46
cc_115 VNB N_A_2555_47#_M1043_g 0.0273556f $X=-0.19 $Y=-0.245 $X2=0.267
+ $Y2=0.912
cc_116 VNB N_A_2555_47#_M1034_g 4.91762e-19 $X=-0.19 $Y=-0.245 $X2=2.77
+ $Y2=1.935
cc_117 VNB N_A_2555_47#_c_1766_n 0.0167915f $X=-0.19 $Y=-0.245 $X2=1.335
+ $Y2=0.945
cc_118 VNB N_A_2555_47#_c_1767_n 0.00262554f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_119 VNB N_A_2555_47#_c_1768_n 0.00224475f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_120 VNB N_A_2555_47#_c_1769_n 8.26908e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_121 VNB N_A_2555_47#_c_1770_n 0.00127147f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_122 VNB N_A_2555_47#_c_1771_n 0.080415f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_123 VNB N_VPWR_c_1876_n 0.641339f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_124 VNB N_A_372_50#_c_2057_n 0.0198151f $X=-0.19 $Y=-0.245 $X2=0.267 $Y2=1.93
cc_125 VNB N_A_372_50#_c_2058_n 0.0094698f $X=-0.19 $Y=-0.245 $X2=1.335
+ $Y2=0.945
cc_126 VNB N_A_372_50#_c_2059_n 0.012502f $X=-0.19 $Y=-0.245 $X2=1.3 $Y2=2.275
cc_127 VNB N_A_372_50#_c_2060_n 0.00710098f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_128 VNB N_A_372_50#_c_2061_n 0.00330174f $X=-0.19 $Y=-0.245 $X2=2.77
+ $Y2=1.935
cc_129 VNB N_A_372_50#_c_2062_n 0.00320714f $X=-0.19 $Y=-0.245 $X2=2.77
+ $Y2=1.935
cc_130 VNB N_A_372_50#_c_2063_n 0.0102239f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_131 VNB N_Q_c_2152_n 0.0030484f $X=-0.19 $Y=-0.245 $X2=1.335 $Y2=0.912
cc_132 VNB N_Q_c_2153_n 0.00263859f $X=-0.19 $Y=-0.245 $X2=1.335 $Y2=0.945
cc_133 VNB N_Q_c_2154_n 0.00899605f $X=-0.19 $Y=-0.245 $X2=2.605 $Y2=2.027
cc_134 VNB N_Q_c_2155_n 0.0217882f $X=-0.19 $Y=-0.245 $X2=1.3 $Y2=2.102
cc_135 VNB N_Q_c_2156_n 0.00200864f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_136 VNB N_VGND_c_2209_n 0.00888741f $X=-0.19 $Y=-0.245 $X2=1.3 $Y2=2.275
cc_137 VNB N_VGND_c_2210_n 0.0063073f $X=-0.19 $Y=-0.245 $X2=2.605 $Y2=2.027
cc_138 VNB N_VGND_c_2211_n 0.0798227f $X=-0.19 $Y=-0.245 $X2=0.267 $Y2=0.912
cc_139 VNB N_VGND_c_2212_n 0.0122954f $X=-0.19 $Y=-0.245 $X2=2.77 $Y2=1.935
cc_140 VNB N_VGND_c_2213_n 0.0115225f $X=-0.19 $Y=-0.245 $X2=1.335 $Y2=0.945
cc_141 VNB N_VGND_c_2214_n 0.00801233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_142 VNB N_VGND_c_2215_n 3.99129e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_143 VNB N_VGND_c_2216_n 3.21684e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_144 VNB N_VGND_c_2217_n 0.0112246f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_145 VNB N_VGND_c_2218_n 0.0297893f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_146 VNB N_VGND_c_2219_n 0.0581579f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_147 VNB N_VGND_c_2220_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_148 VNB N_VGND_c_2221_n 0.0173303f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_149 VNB N_VGND_c_2222_n 0.0580217f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_150 VNB N_VGND_c_2223_n 0.0492511f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_151 VNB N_VGND_c_2224_n 0.0449164f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_152 VNB N_VGND_c_2225_n 0.0129398f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_153 VNB N_VGND_c_2226_n 0.0156677f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_154 VNB N_VGND_c_2227_n 0.00613348f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_155 VNB N_VGND_c_2228_n 0.0034624f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_156 VNB N_VGND_c_2229_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_157 VNB N_VGND_c_2230_n 0.00631381f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_158 VNB N_VGND_c_2231_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_159 VNB N_VGND_c_2232_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_160 VNB N_VGND_c_2233_n 0.762644f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_161 VNB N_noxref_24_c_2367_n 0.00427584f $X=-0.19 $Y=-0.245 $X2=1.425
+ $Y2=0.78
cc_162 VNB N_noxref_24_c_2368_n 0.00393461f $X=-0.19 $Y=-0.245 $X2=1.425
+ $Y2=0.46
cc_163 VNB N_noxref_24_c_2369_n 0.00224633f $X=-0.19 $Y=-0.245 $X2=0.255
+ $Y2=0.795
cc_164 VPB N_A_27_74#_M1020_g 0.0235814f $X=-0.19 $Y=1.655 $X2=2.75 $Y2=2.635
cc_165 VPB N_A_27_74#_c_309_n 0.013109f $X=-0.19 $Y=1.655 $X2=0.267 $Y2=1.93
cc_166 VPB N_A_27_74#_c_316_n 0.0349461f $X=-0.19 $Y=1.655 $X2=1.15 $Y2=2.102
cc_167 VPB N_A_27_74#_c_317_n 0.0239626f $X=-0.19 $Y=1.655 $X2=0.38 $Y2=2.102
cc_168 VPB N_A_27_74#_c_318_n 0.029772f $X=-0.19 $Y=1.655 $X2=1.315 $Y2=2.46
cc_169 VPB N_A_27_74#_c_319_n 0.0168578f $X=-0.19 $Y=1.655 $X2=2.605 $Y2=2.027
cc_170 VPB N_A_27_74#_c_320_n 0.00356547f $X=-0.19 $Y=1.655 $X2=1.3 $Y2=2.102
cc_171 VPB N_A_27_74#_c_321_n 0.00393449f $X=-0.19 $Y=1.655 $X2=2.77 $Y2=1.935
cc_172 VPB N_A_27_74#_c_322_n 0.0333894f $X=-0.19 $Y=1.655 $X2=2.77 $Y2=1.935
cc_173 VPB N_SCE_c_396_n 0.013503f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_174 VPB N_SCE_c_397_n 0.0603914f $X=-0.19 $Y=1.655 $X2=1.425 $Y2=0.78
cc_175 VPB N_SCE_c_398_n 0.0109496f $X=-0.19 $Y=1.655 $X2=1.425 $Y2=0.46
cc_176 VPB N_SCE_c_399_n 0.0209409f $X=-0.19 $Y=1.655 $X2=1.425 $Y2=0.46
cc_177 VPB N_SCE_c_400_n 0.015707f $X=-0.19 $Y=1.655 $X2=2.75 $Y2=2.635
cc_178 VPB N_SCE_c_401_n 0.0161611f $X=-0.19 $Y=1.655 $X2=0.255 $Y2=0.795
cc_179 VPB N_SCE_c_402_n 0.00534401f $X=-0.19 $Y=1.655 $X2=1.335 $Y2=0.912
cc_180 VPB N_SCE_c_393_n 0.0205886f $X=-0.19 $Y=1.655 $X2=1.3 $Y2=2.275
cc_181 VPB N_D_c_476_n 0.0306218f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_182 VPB N_D_M1038_g 0.0386408f $X=-0.19 $Y=1.655 $X2=1.425 $Y2=0.46
cc_183 VPB D 0.00585641f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_184 VPB N_D_c_475_n 0.0179228f $X=-0.19 $Y=1.655 $X2=0.267 $Y2=1.03
cc_185 VPB N_SCD_M1012_g 0.0316639f $X=-0.19 $Y=1.655 $X2=1.425 $Y2=0.46
cc_186 VPB N_SCD_c_523_n 0.0156176f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_187 VPB N_SCD_c_520_n 0.0109701f $X=-0.19 $Y=1.655 $X2=0.267 $Y2=1.93
cc_188 VPB N_SCD_c_521_n 0.00861177f $X=-0.19 $Y=1.655 $X2=0.38 $Y2=0.912
cc_189 VPB N_A_851_242#_M1017_g 0.0389006f $X=-0.19 $Y=1.655 $X2=1.425 $Y2=0.46
cc_190 VPB N_A_851_242#_M1013_g 0.0295214f $X=-0.19 $Y=1.655 $X2=1.335 $Y2=0.912
cc_191 VPB N_A_851_242#_c_586_n 0.0243424f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_192 VPB N_A_851_242#_c_568_n 0.00535688f $X=-0.19 $Y=1.655 $X2=0.38 $Y2=2.102
cc_193 VPB N_A_851_242#_c_588_n 0.00188342f $X=-0.19 $Y=1.655 $X2=2.605
+ $Y2=2.027
cc_194 VPB N_A_851_242#_c_589_n 0.0366336f $X=-0.19 $Y=1.655 $X2=1.45 $Y2=2.027
cc_195 VPB N_A_851_242#_c_577_n 0.00259642f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_196 VPB N_A_851_242#_c_579_n 0.00776905f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_197 VPB N_A_851_242#_c_580_n 0.00155643f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_198 VPB N_A_1047_369#_M1003_g 0.0264748f $X=-0.19 $Y=1.655 $X2=1.425 $Y2=0.46
cc_199 VPB N_A_1047_369#_c_785_n 0.0240078f $X=-0.19 $Y=1.655 $X2=2.75 $Y2=2.635
cc_200 VPB N_A_1047_369#_c_786_n 0.0338754f $X=-0.19 $Y=1.655 $X2=2.75 $Y2=2.635
cc_201 VPB N_A_1047_369#_M1045_g 6.58841e-19 $X=-0.19 $Y=1.655 $X2=0.255
+ $Y2=0.58
cc_202 VPB N_A_1047_369#_c_780_n 0.012146f $X=-0.19 $Y=1.655 $X2=1.335 $Y2=0.945
cc_203 VPB N_A_1047_369#_c_789_n 0.00139803f $X=-0.19 $Y=1.655 $X2=1.315
+ $Y2=2.46
cc_204 VPB N_A_1047_369#_c_790_n 0.00375498f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_205 VPB N_A_1047_369#_c_782_n 0.00337392f $X=-0.19 $Y=1.655 $X2=2.605
+ $Y2=2.027
cc_206 VPB N_A_1047_369#_c_783_n 5.19703e-19 $X=-0.19 $Y=1.655 $X2=1.45
+ $Y2=2.027
cc_207 VPB N_RESET_B_M1033_g 0.0519307f $X=-0.19 $Y=1.655 $X2=1.425 $Y2=0.46
cc_208 VPB N_RESET_B_c_890_n 0.0208497f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_209 VPB N_RESET_B_c_891_n 0.0143356f $X=-0.19 $Y=1.655 $X2=0.26 $Y2=0.58
cc_210 VPB N_RESET_B_c_892_n 0.0085377f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_211 VPB N_RESET_B_M1036_g 0.0117926f $X=-0.19 $Y=1.655 $X2=1.335 $Y2=0.912
cc_212 VPB N_RESET_B_M1026_g 0.0257931f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_213 VPB N_RESET_B_M1018_g 0.0201233f $X=-0.19 $Y=1.655 $X2=1.3 $Y2=2.46
cc_214 VPB N_RESET_B_c_896_n 0.00282931f $X=-0.19 $Y=1.655 $X2=1.45 $Y2=2.027
cc_215 VPB N_RESET_B_c_897_n 0.00401655f $X=-0.19 $Y=1.655 $X2=0.267 $Y2=0.912
cc_216 VPB N_RESET_B_c_898_n 0.00439565f $X=-0.19 $Y=1.655 $X2=1.3 $Y2=2.102
cc_217 VPB N_RESET_B_c_899_n 0.00240857f $X=-0.19 $Y=1.655 $X2=2.77 $Y2=1.935
cc_218 VPB N_RESET_B_c_900_n 0.00134753f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_219 VPB N_RESET_B_c_901_n 0.0194582f $X=-0.19 $Y=1.655 $X2=2.73 $Y2=2.027
cc_220 VPB N_RESET_B_c_902_n 7.70891e-19 $X=-0.19 $Y=1.655 $X2=1.335 $Y2=0.945
cc_221 VPB N_RESET_B_c_903_n 0.00336323f $X=-0.19 $Y=1.655 $X2=2.77 $Y2=2.1
cc_222 VPB N_RESET_B_c_904_n 0.0330111f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_223 VPB N_RESET_B_c_905_n 0.0440374f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_224 VPB N_RESET_B_c_906_n 0.00636775f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_225 VPB N_A_881_463#_M1022_g 0.0243381f $X=-0.19 $Y=1.655 $X2=0.26 $Y2=0.58
cc_226 VPB N_A_881_463#_c_1068_n 0.00409007f $X=-0.19 $Y=1.655 $X2=0.267
+ $Y2=1.93
cc_227 VPB N_A_881_463#_c_1077_n 0.0267189f $X=-0.19 $Y=1.655 $X2=0.38 $Y2=0.912
cc_228 VPB N_A_881_463#_c_1078_n 0.0180522f $X=-0.19 $Y=1.655 $X2=2.73 $Y2=1.935
cc_229 VPB N_A_975_255#_M1007_g 0.0567717f $X=-0.19 $Y=1.655 $X2=2.75 $Y2=2.1
cc_230 VPB N_A_975_255#_c_1223_n 0.199996f $X=-0.19 $Y=1.655 $X2=0.255 $Y2=0.58
cc_231 VPB N_A_975_255#_c_1224_n 0.012806f $X=-0.19 $Y=1.655 $X2=0.26 $Y2=0.58
cc_232 VPB N_A_975_255#_M1010_g 0.0252119f $X=-0.19 $Y=1.655 $X2=0.38 $Y2=0.912
cc_233 VPB N_A_975_255#_c_1209_n 0.00541981f $X=-0.19 $Y=1.655 $X2=1.335
+ $Y2=0.945
cc_234 VPB N_A_975_255#_M1004_g 0.023388f $X=-0.19 $Y=1.655 $X2=0.267 $Y2=0.912
cc_235 VPB N_A_975_255#_c_1213_n 0.0138956f $X=-0.19 $Y=1.655 $X2=2.73 $Y2=2.027
cc_236 VPB N_A_975_255#_c_1229_n 0.0140714f $X=-0.19 $Y=1.655 $X2=1.335 $Y2=0.78
cc_237 VPB N_A_975_255#_c_1230_n 0.0168353f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_238 VPB N_A_975_255#_c_1231_n 0.00364405f $X=-0.19 $Y=1.655 $X2=2.77
+ $Y2=1.935
cc_239 VPB N_A_975_255#_c_1232_n 0.00147063f $X=-0.19 $Y=1.655 $X2=2.77 $Y2=2.1
cc_240 VPB N_A_975_255#_c_1215_n 0.00790569f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_241 VPB N_A_975_255#_c_1217_n 0.0198368f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_242 VPB N_A_975_255#_c_1218_n 9.26678e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_243 VPB N_A_975_255#_c_1219_n 0.00962316f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_244 VPB N_A_975_255#_c_1237_n 9.98093e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_245 VPB N_A_975_255#_c_1238_n 0.0437039f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_246 VPB N_A_1524_69#_M1042_g 0.0720716f $X=-0.19 $Y=1.655 $X2=2.75 $Y2=2.635
cc_247 VPB N_A_1524_69#_M1044_g 0.022984f $X=-0.19 $Y=1.655 $X2=0.267 $Y2=1.93
cc_248 VPB N_A_1524_69#_c_1414_n 0.00101163f $X=-0.19 $Y=1.655 $X2=1.315
+ $Y2=2.46
cc_249 VPB N_A_1524_69#_c_1432_n 0.00137446f $X=-0.19 $Y=1.655 $X2=2.605
+ $Y2=2.027
cc_250 VPB N_A_1747_21#_M1028_g 0.0293761f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_251 VPB N_A_1747_21#_c_1598_n 0.0181846f $X=-0.19 $Y=1.655 $X2=0.267 $Y2=1.03
cc_252 VPB N_A_1747_21#_c_1606_n 0.0150029f $X=-0.19 $Y=1.655 $X2=1.335
+ $Y2=0.945
cc_253 VPB N_A_1747_21#_c_1607_n 0.00442836f $X=-0.19 $Y=1.655 $X2=1.3 $Y2=2.102
cc_254 VPB N_A_1747_21#_c_1608_n 0.00685116f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_255 VPB N_A_1747_21#_c_1609_n 0.036204f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_256 VPB N_CLK_M1037_g 0.0252155f $X=-0.19 $Y=1.655 $X2=1.425 $Y2=0.78
cc_257 VPB N_CLK_c_1710_n 0.0468803f $X=-0.19 $Y=1.655 $X2=0.38 $Y2=0.912
cc_258 VPB N_CLK_c_1711_n 0.0200972f $X=-0.19 $Y=1.655 $X2=1.335 $Y2=0.912
cc_259 VPB N_A_2555_47#_M1005_g 0.0188277f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_260 VPB N_A_2555_47#_M1008_g 0.0192305f $X=-0.19 $Y=1.655 $X2=1.335 $Y2=0.912
cc_261 VPB N_A_2555_47#_M1025_g 0.0192147f $X=-0.19 $Y=1.655 $X2=1.315 $Y2=2.46
cc_262 VPB N_A_2555_47#_M1034_g 0.0225169f $X=-0.19 $Y=1.655 $X2=2.77 $Y2=1.935
cc_263 VPB N_A_2555_47#_c_1776_n 0.0263273f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_264 VPB N_A_2555_47#_c_1777_n 0.00422168f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_265 VPB N_A_2555_47#_c_1778_n 0.00401432f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_266 VPB N_A_2555_47#_c_1769_n 9.19819e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_267 VPB N_VPWR_c_1877_n 0.00807184f $X=-0.19 $Y=1.655 $X2=0.267 $Y2=0.912
cc_268 VPB N_VPWR_c_1878_n 0.0101057f $X=-0.19 $Y=1.655 $X2=2.77 $Y2=1.935
cc_269 VPB N_VPWR_c_1879_n 0.0129392f $X=-0.19 $Y=1.655 $X2=1.335 $Y2=0.945
cc_270 VPB N_VPWR_c_1880_n 0.0203059f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_271 VPB N_VPWR_c_1881_n 0.00602232f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_272 VPB N_VPWR_c_1882_n 0.00733303f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_273 VPB N_VPWR_c_1883_n 0.00386019f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_274 VPB N_VPWR_c_1884_n 4.02668e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_275 VPB N_VPWR_c_1885_n 3.16188e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_276 VPB N_VPWR_c_1886_n 0.0105563f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_277 VPB N_VPWR_c_1887_n 0.0392694f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_278 VPB N_VPWR_c_1888_n 0.0517434f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_279 VPB N_VPWR_c_1889_n 0.00631679f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_280 VPB N_VPWR_c_1890_n 0.0513897f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_281 VPB N_VPWR_c_1891_n 0.0432568f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_282 VPB N_VPWR_c_1892_n 0.0474515f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_283 VPB N_VPWR_c_1893_n 0.0277157f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_284 VPB N_VPWR_c_1894_n 0.0227641f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_285 VPB N_VPWR_c_1895_n 0.0206876f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_286 VPB N_VPWR_c_1896_n 0.0439372f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_287 VPB N_VPWR_c_1897_n 0.0133881f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_288 VPB N_VPWR_c_1898_n 0.0134822f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_289 VPB N_VPWR_c_1899_n 0.00540054f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_290 VPB N_VPWR_c_1900_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_291 VPB N_VPWR_c_1901_n 0.00450185f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_292 VPB N_VPWR_c_1902_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_293 VPB N_VPWR_c_1903_n 0.00382106f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_294 VPB N_VPWR_c_1904_n 0.00866685f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_295 VPB N_VPWR_c_1905_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_296 VPB N_VPWR_c_1906_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_297 VPB N_VPWR_c_1876_n 0.146251f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_298 VPB N_A_372_50#_c_2064_n 0.0152959f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_299 VPB N_A_372_50#_c_2058_n 0.00857798f $X=-0.19 $Y=1.655 $X2=1.335
+ $Y2=0.945
cc_300 VPB N_A_372_50#_c_2066_n 0.00482227f $X=-0.19 $Y=1.655 $X2=2.73 $Y2=1.935
cc_301 VPB N_A_372_50#_c_2067_n 0.00342651f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_302 VPB N_Q_c_2157_n 0.00241216f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_303 VPB N_Q_c_2158_n 0.00293074f $X=-0.19 $Y=1.655 $X2=1.335 $Y2=0.945
cc_304 VPB N_Q_c_2159_n 0.0126062f $X=-0.19 $Y=1.655 $X2=1.315 $Y2=2.46
cc_305 VPB N_Q_c_2155_n 0.00399136f $X=-0.19 $Y=1.655 $X2=1.3 $Y2=2.102
cc_306 VPB N_Q_c_2161_n 0.00153535f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_307 N_A_27_74#_c_323_p N_SCE_M1000_g 4.49244e-19 $X=0.26 $Y=0.58 $X2=0 $Y2=0
cc_308 N_A_27_74#_c_309_n N_SCE_M1000_g 0.0319394f $X=0.267 $Y=1.93 $X2=0 $Y2=0
cc_309 N_A_27_74#_c_310_n N_SCE_M1000_g 0.022439f $X=1.335 $Y=0.945 $X2=0 $Y2=0
cc_310 N_A_27_74#_c_311_n N_SCE_M1000_g 0.00547964f $X=1.335 $Y=0.945 $X2=0
+ $Y2=0
cc_311 N_A_27_74#_c_316_n N_SCE_c_396_n 0.0121199f $X=1.15 $Y=2.102 $X2=0 $Y2=0
cc_312 N_A_27_74#_c_316_n N_SCE_c_397_n 0.0242535f $X=1.15 $Y=2.102 $X2=0 $Y2=0
cc_313 N_A_27_74#_c_320_n N_SCE_c_397_n 0.020464f $X=1.3 $Y=2.102 $X2=0 $Y2=0
cc_314 N_A_27_74#_c_316_n N_SCE_c_398_n 0.00732621f $X=1.15 $Y=2.102 $X2=0 $Y2=0
cc_315 N_A_27_74#_c_318_n N_SCE_c_399_n 0.00179838f $X=1.315 $Y=2.46 $X2=0 $Y2=0
cc_316 N_A_27_74#_c_320_n N_SCE_c_399_n 0.00342718f $X=1.3 $Y=2.102 $X2=0 $Y2=0
cc_317 N_A_27_74#_c_319_n N_SCE_c_400_n 0.015353f $X=2.605 $Y=2.027 $X2=0 $Y2=0
cc_318 N_A_27_74#_c_319_n N_SCE_c_402_n 0.00937969f $X=2.605 $Y=2.027 $X2=0
+ $Y2=0
cc_319 N_A_27_74#_c_309_n N_SCE_c_416_n 0.0435057f $X=0.267 $Y=1.93 $X2=0 $Y2=0
cc_320 N_A_27_74#_c_310_n N_SCE_c_416_n 0.0259988f $X=1.335 $Y=0.945 $X2=0 $Y2=0
cc_321 N_A_27_74#_c_316_n N_SCE_c_416_n 0.0271947f $X=1.15 $Y=2.102 $X2=0 $Y2=0
cc_322 N_A_27_74#_c_310_n N_SCE_c_393_n 0.00938374f $X=1.335 $Y=0.945 $X2=0
+ $Y2=0
cc_323 N_A_27_74#_c_316_n N_SCE_c_393_n 0.00249879f $X=1.15 $Y=2.102 $X2=0 $Y2=0
cc_324 N_A_27_74#_c_310_n SCE 0.0460279f $X=1.335 $Y=0.945 $X2=0 $Y2=0
cc_325 N_A_27_74#_c_311_n SCE 0.00877681f $X=1.335 $Y=0.945 $X2=0 $Y2=0
cc_326 N_A_27_74#_c_316_n SCE 0.00619643f $X=1.15 $Y=2.102 $X2=0 $Y2=0
cc_327 N_A_27_74#_c_319_n SCE 0.00877048f $X=2.605 $Y=2.027 $X2=0 $Y2=0
cc_328 N_A_27_74#_c_321_n SCE 0.00823536f $X=2.77 $Y=1.935 $X2=0 $Y2=0
cc_329 N_A_27_74#_c_322_n SCE 8.36472e-19 $X=2.77 $Y=1.935 $X2=0 $Y2=0
cc_330 N_A_27_74#_c_319_n N_SCE_c_395_n 0.0028594f $X=2.605 $Y=2.027 $X2=0 $Y2=0
cc_331 N_A_27_74#_c_310_n N_D_M1023_g 9.71503e-19 $X=1.335 $Y=0.945 $X2=0 $Y2=0
cc_332 N_A_27_74#_c_313_n N_D_M1023_g 0.0626452f $X=1.335 $Y=0.78 $X2=0 $Y2=0
cc_333 N_A_27_74#_c_321_n N_D_c_476_n 0.00113723f $X=2.77 $Y=1.935 $X2=0 $Y2=0
cc_334 N_A_27_74#_c_322_n N_D_c_476_n 0.0216649f $X=2.77 $Y=1.935 $X2=0 $Y2=0
cc_335 N_A_27_74#_M1020_g N_D_M1038_g 0.0171312f $X=2.75 $Y=2.635 $X2=0 $Y2=0
cc_336 N_A_27_74#_c_319_n N_D_M1038_g 0.0163173f $X=2.605 $Y=2.027 $X2=0 $Y2=0
cc_337 N_A_27_74#_c_316_n D 0.00797832f $X=1.15 $Y=2.102 $X2=0 $Y2=0
cc_338 N_A_27_74#_c_319_n D 0.0636786f $X=2.605 $Y=2.027 $X2=0 $Y2=0
cc_339 N_A_27_74#_c_320_n D 0.0255298f $X=1.3 $Y=2.102 $X2=0 $Y2=0
cc_340 N_A_27_74#_c_319_n N_D_c_475_n 0.00758203f $X=2.605 $Y=2.027 $X2=0 $Y2=0
cc_341 N_A_27_74#_c_321_n N_SCD_c_519_n 7.17435e-19 $X=2.77 $Y=1.935 $X2=0 $Y2=0
cc_342 N_A_27_74#_c_322_n N_SCD_c_519_n 0.00862957f $X=2.77 $Y=1.935 $X2=0 $Y2=0
cc_343 N_A_27_74#_M1020_g N_SCD_M1012_g 0.0382697f $X=2.75 $Y=2.635 $X2=0 $Y2=0
cc_344 N_A_27_74#_c_321_n N_SCD_c_520_n 2.89551e-19 $X=2.77 $Y=1.935 $X2=0 $Y2=0
cc_345 N_A_27_74#_c_322_n N_SCD_c_520_n 0.0203253f $X=2.77 $Y=1.935 $X2=0 $Y2=0
cc_346 N_A_27_74#_c_321_n N_SCD_c_521_n 0.0283447f $X=2.77 $Y=1.935 $X2=0 $Y2=0
cc_347 N_A_27_74#_c_322_n N_SCD_c_521_n 0.00226005f $X=2.77 $Y=1.935 $X2=0 $Y2=0
cc_348 N_A_27_74#_c_318_n N_VPWR_c_1877_n 0.00310866f $X=1.315 $Y=2.46 $X2=0
+ $Y2=0
cc_349 N_A_27_74#_c_319_n N_VPWR_c_1877_n 0.0233053f $X=2.605 $Y=2.027 $X2=0
+ $Y2=0
cc_350 N_A_27_74#_c_318_n N_VPWR_c_1890_n 0.0130355f $X=1.315 $Y=2.46 $X2=0
+ $Y2=0
cc_351 N_A_27_74#_M1020_g N_VPWR_c_1891_n 0.00430542f $X=2.75 $Y=2.635 $X2=0
+ $Y2=0
cc_352 N_A_27_74#_M1020_g N_VPWR_c_1876_n 0.00544287f $X=2.75 $Y=2.635 $X2=0
+ $Y2=0
cc_353 N_A_27_74#_c_318_n N_VPWR_c_1876_n 0.010973f $X=1.315 $Y=2.46 $X2=0 $Y2=0
cc_354 N_A_27_74#_M1020_g N_A_372_50#_c_2064_n 0.00901268f $X=2.75 $Y=2.635
+ $X2=0 $Y2=0
cc_355 N_A_27_74#_c_321_n N_A_372_50#_c_2064_n 0.0113619f $X=2.77 $Y=1.935 $X2=0
+ $Y2=0
cc_356 N_A_27_74#_c_322_n N_A_372_50#_c_2064_n 0.00317122f $X=2.77 $Y=1.935
+ $X2=0 $Y2=0
cc_357 N_A_27_74#_c_310_n N_A_372_50#_c_2060_n 0.00759774f $X=1.335 $Y=0.945
+ $X2=0 $Y2=0
cc_358 N_A_27_74#_M1020_g N_A_372_50#_c_2066_n 0.0110893f $X=2.75 $Y=2.635 $X2=0
+ $Y2=0
cc_359 N_A_27_74#_c_319_n N_A_372_50#_c_2066_n 0.0198266f $X=2.605 $Y=2.027
+ $X2=0 $Y2=0
cc_360 N_A_27_74#_c_321_n N_A_372_50#_c_2066_n 0.00817964f $X=2.77 $Y=1.935
+ $X2=0 $Y2=0
cc_361 N_A_27_74#_c_322_n N_A_372_50#_c_2066_n 5.06953e-19 $X=2.77 $Y=1.935
+ $X2=0 $Y2=0
cc_362 N_A_27_74#_c_310_n N_VGND_c_2209_n 0.0243845f $X=1.335 $Y=0.945 $X2=0
+ $Y2=0
cc_363 N_A_27_74#_c_313_n N_VGND_c_2209_n 0.00285585f $X=1.335 $Y=0.78 $X2=0
+ $Y2=0
cc_364 N_A_27_74#_c_323_p N_VGND_c_2221_n 0.00660406f $X=0.26 $Y=0.58 $X2=0
+ $Y2=0
cc_365 N_A_27_74#_c_313_n N_VGND_c_2222_n 0.00349398f $X=1.335 $Y=0.78 $X2=0
+ $Y2=0
cc_366 N_A_27_74#_c_323_p N_VGND_c_2233_n 0.00701926f $X=0.26 $Y=0.58 $X2=0
+ $Y2=0
cc_367 N_A_27_74#_c_310_n N_VGND_c_2233_n 0.0135299f $X=1.335 $Y=0.945 $X2=0
+ $Y2=0
cc_368 N_A_27_74#_c_312_n N_VGND_c_2233_n 0.00102567f $X=0.267 $Y=0.912 $X2=0
+ $Y2=0
cc_369 N_A_27_74#_c_313_n N_VGND_c_2233_n 0.00634764f $X=1.335 $Y=0.78 $X2=0
+ $Y2=0
cc_370 N_A_27_74#_c_310_n N_noxref_24_c_2367_n 0.004008f $X=1.335 $Y=0.945 $X2=0
+ $Y2=0
cc_371 N_A_27_74#_c_313_n N_noxref_24_c_2367_n 0.00766371f $X=1.335 $Y=0.78
+ $X2=0 $Y2=0
cc_372 N_A_27_74#_c_310_n N_noxref_24_c_2368_n 0.02259f $X=1.335 $Y=0.945 $X2=0
+ $Y2=0
cc_373 N_A_27_74#_c_311_n N_noxref_24_c_2368_n 0.00403618f $X=1.335 $Y=0.945
+ $X2=0 $Y2=0
cc_374 N_A_27_74#_c_313_n N_noxref_24_c_2368_n 0.00508143f $X=1.335 $Y=0.78
+ $X2=0 $Y2=0
cc_375 N_SCE_M1029_g N_D_M1023_g 0.0178978f $X=2.445 $Y=0.615 $X2=0 $Y2=0
cc_376 SCE N_D_M1023_g 0.0180919f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_377 N_SCE_c_395_n N_D_M1023_g 0.0192623f $X=2.445 $Y=1.295 $X2=0 $Y2=0
cc_378 N_SCE_c_400_n N_D_c_476_n 0.0143003f $X=1.885 $Y=2.13 $X2=0 $Y2=0
cc_379 SCE N_D_c_476_n 0.00181258f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_380 N_SCE_c_395_n N_D_c_476_n 0.0177311f $X=2.445 $Y=1.295 $X2=0 $Y2=0
cc_381 N_SCE_c_400_n N_D_M1038_g 0.0616745f $X=1.885 $Y=2.13 $X2=0 $Y2=0
cc_382 N_SCE_c_397_n D 0.00253516f $X=1.455 $Y=2.13 $X2=0 $Y2=0
cc_383 N_SCE_c_402_n D 4.48282e-19 $X=1.53 $Y=2.13 $X2=0 $Y2=0
cc_384 N_SCE_c_416_n D 0.0158547f $X=0.715 $Y=1.295 $X2=0 $Y2=0
cc_385 N_SCE_c_393_n D 0.00223362f $X=0.715 $Y=1.295 $X2=0 $Y2=0
cc_386 SCE D 0.0951316f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_387 N_SCE_c_395_n D 0.00138741f $X=2.445 $Y=1.295 $X2=0 $Y2=0
cc_388 N_SCE_c_402_n N_D_c_475_n 0.0143003f $X=1.53 $Y=2.13 $X2=0 $Y2=0
cc_389 N_SCE_c_416_n N_D_c_475_n 5.10582e-19 $X=0.715 $Y=1.295 $X2=0 $Y2=0
cc_390 N_SCE_c_393_n N_D_c_475_n 0.00488854f $X=0.715 $Y=1.295 $X2=0 $Y2=0
cc_391 SCE N_D_c_475_n 0.00439839f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_392 N_SCE_M1029_g N_SCD_M1032_g 0.0374024f $X=2.445 $Y=0.615 $X2=0 $Y2=0
cc_393 SCE N_SCD_M1032_g 0.00617333f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_394 SCE N_SCD_c_519_n 0.00433856f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_395 N_SCE_c_395_n N_SCD_c_519_n 0.0374024f $X=2.445 $Y=1.295 $X2=0 $Y2=0
cc_396 N_SCE_c_395_n N_SCD_c_520_n 2.7498e-19 $X=2.445 $Y=1.295 $X2=0 $Y2=0
cc_397 SCE N_SCD_c_521_n 0.0072346f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_398 N_SCE_c_395_n N_SCD_c_521_n 6.21144e-19 $X=2.445 $Y=1.295 $X2=0 $Y2=0
cc_399 N_SCE_c_399_n N_VPWR_c_1877_n 0.00337203f $X=1.53 $Y=2.205 $X2=0 $Y2=0
cc_400 N_SCE_c_400_n N_VPWR_c_1877_n 0.00220396f $X=1.885 $Y=2.13 $X2=0 $Y2=0
cc_401 N_SCE_c_401_n N_VPWR_c_1877_n 0.0149865f $X=1.96 $Y=2.205 $X2=0 $Y2=0
cc_402 N_SCE_c_399_n N_VPWR_c_1890_n 0.00457417f $X=1.53 $Y=2.205 $X2=0 $Y2=0
cc_403 N_SCE_c_401_n N_VPWR_c_1891_n 0.00379792f $X=1.96 $Y=2.205 $X2=0 $Y2=0
cc_404 N_SCE_c_399_n N_VPWR_c_1876_n 0.00544287f $X=1.53 $Y=2.205 $X2=0 $Y2=0
cc_405 N_SCE_c_401_n N_VPWR_c_1876_n 0.00457201f $X=1.96 $Y=2.205 $X2=0 $Y2=0
cc_406 N_SCE_M1029_g N_A_372_50#_c_2060_n 0.00605239f $X=2.445 $Y=0.615 $X2=0
+ $Y2=0
cc_407 SCE N_A_372_50#_c_2060_n 0.0215923f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_408 N_SCE_c_395_n N_A_372_50#_c_2060_n 0.00435587f $X=2.445 $Y=1.295 $X2=0
+ $Y2=0
cc_409 N_SCE_c_401_n N_A_372_50#_c_2066_n 0.00184782f $X=1.96 $Y=2.205 $X2=0
+ $Y2=0
cc_410 N_SCE_M1029_g N_A_372_50#_c_2061_n 0.0111226f $X=2.445 $Y=0.615 $X2=0
+ $Y2=0
cc_411 SCE N_A_372_50#_c_2061_n 0.0312464f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_412 N_SCE_c_395_n N_A_372_50#_c_2061_n 0.0021331f $X=2.445 $Y=1.295 $X2=0
+ $Y2=0
cc_413 N_SCE_M1000_g N_VGND_c_2209_n 0.0131547f $X=0.475 $Y=0.58 $X2=0 $Y2=0
cc_414 N_SCE_M1000_g N_VGND_c_2221_n 0.00383152f $X=0.475 $Y=0.58 $X2=0 $Y2=0
cc_415 N_SCE_M1029_g N_VGND_c_2222_n 9.15902e-19 $X=2.445 $Y=0.615 $X2=0 $Y2=0
cc_416 N_SCE_M1000_g N_VGND_c_2233_n 0.00378113f $X=0.475 $Y=0.58 $X2=0 $Y2=0
cc_417 N_SCE_M1029_g N_noxref_24_c_2367_n 0.0114573f $X=2.445 $Y=0.615 $X2=0
+ $Y2=0
cc_418 N_SCE_M1000_g N_noxref_24_c_2368_n 8.45104e-19 $X=0.475 $Y=0.58 $X2=0
+ $Y2=0
cc_419 N_SCE_M1029_g N_noxref_24_c_2369_n 0.00106586f $X=2.445 $Y=0.615 $X2=0
+ $Y2=0
cc_420 N_D_c_476_n N_SCD_c_521_n 0.00256385f $X=2.245 $Y=1.755 $X2=0 $Y2=0
cc_421 N_D_M1038_g N_VPWR_c_1877_n 0.00240528f $X=2.32 $Y=2.635 $X2=0 $Y2=0
cc_422 N_D_M1038_g N_VPWR_c_1891_n 0.00430542f $X=2.32 $Y=2.635 $X2=0 $Y2=0
cc_423 N_D_M1038_g N_VPWR_c_1876_n 0.00544287f $X=2.32 $Y=2.635 $X2=0 $Y2=0
cc_424 N_D_M1023_g N_A_372_50#_c_2060_n 0.00789148f $X=1.785 $Y=0.46 $X2=0 $Y2=0
cc_425 N_D_M1038_g N_A_372_50#_c_2066_n 0.0118526f $X=2.32 $Y=2.635 $X2=0 $Y2=0
cc_426 N_D_M1023_g N_VGND_c_2222_n 0.00347949f $X=1.785 $Y=0.46 $X2=0 $Y2=0
cc_427 N_D_M1023_g N_VGND_c_2233_n 0.00635675f $X=1.785 $Y=0.46 $X2=0 $Y2=0
cc_428 N_D_M1023_g N_noxref_24_c_2367_n 0.0148566f $X=1.785 $Y=0.46 $X2=0 $Y2=0
cc_429 N_D_M1023_g N_noxref_24_c_2368_n 0.00101608f $X=1.785 $Y=0.46 $X2=0 $Y2=0
cc_430 N_SCD_M1032_g N_RESET_B_M1001_g 0.016346f $X=2.805 $Y=0.615 $X2=0 $Y2=0
cc_431 N_SCD_c_518_n N_RESET_B_M1001_g 0.00542897f $X=3.145 $Y=1.365 $X2=0 $Y2=0
cc_432 N_SCD_c_518_n N_RESET_B_M1033_g 0.0311684f $X=3.145 $Y=1.365 $X2=0 $Y2=0
cc_433 N_SCD_M1012_g N_RESET_B_M1033_g 0.0257005f $X=3.22 $Y=2.635 $X2=0 $Y2=0
cc_434 N_SCD_c_521_n N_RESET_B_M1033_g 0.00359082f $X=3.31 $Y=1.455 $X2=0 $Y2=0
cc_435 N_SCD_M1012_g N_VPWR_c_1878_n 0.0084767f $X=3.22 $Y=2.635 $X2=0 $Y2=0
cc_436 N_SCD_M1012_g N_VPWR_c_1891_n 0.00457417f $X=3.22 $Y=2.635 $X2=0 $Y2=0
cc_437 N_SCD_M1012_g N_VPWR_c_1876_n 0.00544287f $X=3.22 $Y=2.635 $X2=0 $Y2=0
cc_438 N_SCD_M1012_g N_A_372_50#_c_2064_n 0.013294f $X=3.22 $Y=2.635 $X2=0 $Y2=0
cc_439 N_SCD_c_523_n N_A_372_50#_c_2064_n 8.39989e-19 $X=3.31 $Y=1.96 $X2=0
+ $Y2=0
cc_440 N_SCD_c_521_n N_A_372_50#_c_2064_n 0.0367383f $X=3.31 $Y=1.455 $X2=0
+ $Y2=0
cc_441 N_SCD_c_518_n N_A_372_50#_c_2058_n 0.0024106f $X=3.145 $Y=1.365 $X2=0
+ $Y2=0
cc_442 N_SCD_M1012_g N_A_372_50#_c_2058_n 0.00102196f $X=3.22 $Y=2.635 $X2=0
+ $Y2=0
cc_443 N_SCD_c_521_n N_A_372_50#_c_2058_n 0.0418807f $X=3.31 $Y=1.455 $X2=0
+ $Y2=0
cc_444 N_SCD_M1012_g N_A_372_50#_c_2066_n 0.00184071f $X=3.22 $Y=2.635 $X2=0
+ $Y2=0
cc_445 N_SCD_M1032_g N_A_372_50#_c_2061_n 0.0131819f $X=2.805 $Y=0.615 $X2=0
+ $Y2=0
cc_446 N_SCD_c_518_n N_A_372_50#_c_2061_n 7.1136e-19 $X=3.145 $Y=1.365 $X2=0
+ $Y2=0
cc_447 N_SCD_M1032_g N_A_372_50#_c_2062_n 0.00380547f $X=2.805 $Y=0.615 $X2=0
+ $Y2=0
cc_448 N_SCD_c_518_n N_A_372_50#_c_2062_n 0.00658393f $X=3.145 $Y=1.365 $X2=0
+ $Y2=0
cc_449 N_SCD_c_521_n N_A_372_50#_c_2062_n 0.0289934f $X=3.31 $Y=1.455 $X2=0
+ $Y2=0
cc_450 N_SCD_M1012_g N_A_372_50#_c_2067_n 8.16079e-19 $X=3.22 $Y=2.635 $X2=0
+ $Y2=0
cc_451 N_SCD_M1032_g N_VGND_c_2222_n 9.09582e-19 $X=2.805 $Y=0.615 $X2=0 $Y2=0
cc_452 N_SCD_M1032_g N_noxref_24_c_2367_n 0.00800592f $X=2.805 $Y=0.615 $X2=0
+ $Y2=0
cc_453 N_SCD_M1032_g N_noxref_24_c_2369_n 0.00679692f $X=2.805 $Y=0.615 $X2=0
+ $Y2=0
cc_454 N_A_851_242#_c_573_n N_A_1047_369#_c_785_n 0.00234508f $X=7.775 $Y=1.295
+ $X2=0 $Y2=0
cc_455 N_A_851_242#_c_574_n N_A_1047_369#_c_785_n 4.36016e-19 $X=5.665 $Y=1.295
+ $X2=0 $Y2=0
cc_456 N_A_851_242#_c_571_n N_A_1047_369#_c_786_n 0.00230901f $X=5.375 $Y=1.295
+ $X2=0 $Y2=0
cc_457 N_A_851_242#_c_574_n N_A_1047_369#_c_786_n 2.06305e-19 $X=5.665 $Y=1.295
+ $X2=0 $Y2=0
cc_458 N_A_851_242#_c_581_n N_A_1047_369#_c_786_n 0.0213082f $X=5.48 $Y=1.29
+ $X2=0 $Y2=0
cc_459 N_A_851_242#_c_598_p N_A_1047_369#_c_786_n 7.89316e-19 $X=5.48 $Y=1.29
+ $X2=0 $Y2=0
cc_460 N_A_851_242#_c_574_n N_A_1047_369#_M1045_g 3.63802e-19 $X=5.665 $Y=1.295
+ $X2=0 $Y2=0
cc_461 N_A_851_242#_c_581_n N_A_1047_369#_M1045_g 0.021747f $X=5.48 $Y=1.29
+ $X2=0 $Y2=0
cc_462 N_A_851_242#_c_598_p N_A_1047_369#_M1045_g 9.13873e-19 $X=5.48 $Y=1.29
+ $X2=0 $Y2=0
cc_463 N_A_851_242#_c_582_n N_A_1047_369#_M1045_g 0.0256607f $X=5.48 $Y=1.125
+ $X2=0 $Y2=0
cc_464 N_A_851_242#_c_573_n N_A_1047_369#_c_780_n 0.00691981f $X=7.775 $Y=1.295
+ $X2=0 $Y2=0
cc_465 N_A_851_242#_c_565_n N_A_1047_369#_c_781_n 0.00841785f $X=7.545 $Y=1.095
+ $X2=0 $Y2=0
cc_466 N_A_851_242#_c_573_n N_A_1047_369#_c_781_n 0.0213301f $X=7.775 $Y=1.295
+ $X2=0 $Y2=0
cc_467 N_A_851_242#_c_571_n N_A_1047_369#_c_790_n 0.004005f $X=5.375 $Y=1.295
+ $X2=0 $Y2=0
cc_468 N_A_851_242#_c_573_n N_A_1047_369#_c_790_n 0.00516485f $X=7.775 $Y=1.295
+ $X2=0 $Y2=0
cc_469 N_A_851_242#_c_574_n N_A_1047_369#_c_790_n 0.00387828f $X=5.665 $Y=1.295
+ $X2=0 $Y2=0
cc_470 N_A_851_242#_c_581_n N_A_1047_369#_c_790_n 0.00159855f $X=5.48 $Y=1.29
+ $X2=0 $Y2=0
cc_471 N_A_851_242#_c_598_p N_A_1047_369#_c_790_n 0.0128597f $X=5.48 $Y=1.29
+ $X2=0 $Y2=0
cc_472 N_A_851_242#_c_573_n N_A_1047_369#_c_782_n 0.00781254f $X=7.775 $Y=1.295
+ $X2=0 $Y2=0
cc_473 N_A_851_242#_c_567_n N_A_1047_369#_c_812_n 2.55326e-19 $X=7.62 $Y=1.17
+ $X2=0 $Y2=0
cc_474 N_A_851_242#_c_573_n N_A_1047_369#_c_812_n 0.00602878f $X=7.775 $Y=1.295
+ $X2=0 $Y2=0
cc_475 N_A_851_242#_c_577_n N_RESET_B_M1033_g 6.76405e-19 $X=4.56 $Y=1.295 $X2=0
+ $Y2=0
cc_476 N_A_851_242#_c_580_n N_RESET_B_M1033_g 0.0366865f $X=4.5 $Y=1.375 $X2=0
+ $Y2=0
cc_477 N_A_851_242#_c_582_n N_RESET_B_c_885_n 0.00979198f $X=5.48 $Y=1.125 $X2=0
+ $Y2=0
cc_478 N_A_851_242#_c_575_n N_RESET_B_M1026_g 0.00196567f $X=10.655 $Y=1.295
+ $X2=0 $Y2=0
cc_479 N_A_851_242#_M1013_g N_RESET_B_c_899_n 0.00560569f $X=8.235 $Y=2.875
+ $X2=0 $Y2=0
cc_480 N_A_851_242#_M1013_g N_RESET_B_c_901_n 5.18957e-19 $X=8.235 $Y=2.875
+ $X2=0 $Y2=0
cc_481 N_A_851_242#_c_588_n N_RESET_B_c_901_n 0.0132847f $X=8.375 $Y=2.22 $X2=0
+ $Y2=0
cc_482 N_A_851_242#_c_589_n N_RESET_B_c_901_n 0.00438376f $X=8.375 $Y=2.22 $X2=0
+ $Y2=0
cc_483 N_A_851_242#_M1013_g N_RESET_B_c_902_n 0.0149829f $X=8.235 $Y=2.875 $X2=0
+ $Y2=0
cc_484 N_A_851_242#_c_588_n N_RESET_B_c_902_n 0.0128651f $X=8.375 $Y=2.22 $X2=0
+ $Y2=0
cc_485 N_A_851_242#_c_589_n N_RESET_B_c_902_n 0.00122199f $X=8.375 $Y=2.22 $X2=0
+ $Y2=0
cc_486 N_A_851_242#_c_565_n N_A_881_463#_M1015_g 0.00914384f $X=7.545 $Y=1.095
+ $X2=0 $Y2=0
cc_487 N_A_851_242#_M1017_g N_A_881_463#_c_1068_n 0.00193416f $X=4.33 $Y=2.525
+ $X2=0 $Y2=0
cc_488 N_A_851_242#_c_571_n N_A_881_463#_c_1068_n 0.00387234f $X=5.375 $Y=1.295
+ $X2=0 $Y2=0
cc_489 N_A_851_242#_c_572_n N_A_881_463#_c_1068_n 9.19145e-19 $X=4.705 $Y=1.295
+ $X2=0 $Y2=0
cc_490 N_A_851_242#_c_574_n N_A_881_463#_c_1068_n 6.19539e-19 $X=5.665 $Y=1.295
+ $X2=0 $Y2=0
cc_491 N_A_851_242#_c_577_n N_A_881_463#_c_1068_n 0.036478f $X=4.56 $Y=1.295
+ $X2=0 $Y2=0
cc_492 N_A_851_242#_c_580_n N_A_881_463#_c_1068_n 0.00280941f $X=4.5 $Y=1.375
+ $X2=0 $Y2=0
cc_493 N_A_851_242#_c_581_n N_A_881_463#_c_1068_n 2.57155e-19 $X=5.48 $Y=1.29
+ $X2=0 $Y2=0
cc_494 N_A_851_242#_c_598_p N_A_881_463#_c_1068_n 0.0022421f $X=5.48 $Y=1.29
+ $X2=0 $Y2=0
cc_495 N_A_851_242#_c_571_n N_A_881_463#_c_1069_n 0.00365481f $X=5.375 $Y=1.295
+ $X2=0 $Y2=0
cc_496 N_A_851_242#_c_572_n N_A_881_463#_c_1069_n 7.66037e-19 $X=4.705 $Y=1.295
+ $X2=0 $Y2=0
cc_497 N_A_851_242#_c_574_n N_A_881_463#_c_1069_n 7.51009e-19 $X=5.665 $Y=1.295
+ $X2=0 $Y2=0
cc_498 N_A_851_242#_c_577_n N_A_881_463#_c_1069_n 0.0023084f $X=4.56 $Y=1.295
+ $X2=0 $Y2=0
cc_499 N_A_851_242#_c_581_n N_A_881_463#_c_1069_n 5.1983e-19 $X=5.48 $Y=1.29
+ $X2=0 $Y2=0
cc_500 N_A_851_242#_c_598_p N_A_881_463#_c_1069_n 0.00586848f $X=5.48 $Y=1.29
+ $X2=0 $Y2=0
cc_501 N_A_851_242#_c_582_n N_A_881_463#_c_1069_n 0.00147577f $X=5.48 $Y=1.125
+ $X2=0 $Y2=0
cc_502 N_A_851_242#_c_571_n N_A_881_463#_c_1095_n 0.00675359f $X=5.375 $Y=1.295
+ $X2=0 $Y2=0
cc_503 N_A_851_242#_c_573_n N_A_881_463#_c_1095_n 0.00521395f $X=7.775 $Y=1.295
+ $X2=0 $Y2=0
cc_504 N_A_851_242#_c_574_n N_A_881_463#_c_1095_n 0.00421778f $X=5.665 $Y=1.295
+ $X2=0 $Y2=0
cc_505 N_A_851_242#_c_581_n N_A_881_463#_c_1095_n 0.00455827f $X=5.48 $Y=1.29
+ $X2=0 $Y2=0
cc_506 N_A_851_242#_c_598_p N_A_881_463#_c_1095_n 0.0140128f $X=5.48 $Y=1.29
+ $X2=0 $Y2=0
cc_507 N_A_851_242#_c_582_n N_A_881_463#_c_1095_n 0.0128552f $X=5.48 $Y=1.125
+ $X2=0 $Y2=0
cc_508 N_A_851_242#_c_581_n N_A_881_463#_c_1070_n 2.25477e-19 $X=5.48 $Y=1.29
+ $X2=0 $Y2=0
cc_509 N_A_851_242#_c_598_p N_A_881_463#_c_1070_n 0.00282898f $X=5.48 $Y=1.29
+ $X2=0 $Y2=0
cc_510 N_A_851_242#_c_582_n N_A_881_463#_c_1070_n 0.00146301f $X=5.48 $Y=1.125
+ $X2=0 $Y2=0
cc_511 N_A_851_242#_c_573_n N_A_881_463#_c_1071_n 0.0151543f $X=7.775 $Y=1.295
+ $X2=0 $Y2=0
cc_512 N_A_851_242#_c_574_n N_A_881_463#_c_1071_n 0.00203161f $X=5.665 $Y=1.295
+ $X2=0 $Y2=0
cc_513 N_A_851_242#_c_581_n N_A_881_463#_c_1071_n 0.00112005f $X=5.48 $Y=1.29
+ $X2=0 $Y2=0
cc_514 N_A_851_242#_c_598_p N_A_881_463#_c_1071_n 0.0156447f $X=5.48 $Y=1.29
+ $X2=0 $Y2=0
cc_515 N_A_851_242#_c_573_n N_A_881_463#_c_1072_n 0.059136f $X=7.775 $Y=1.295
+ $X2=0 $Y2=0
cc_516 N_A_851_242#_M1017_g N_A_881_463#_c_1078_n 0.0072156f $X=4.33 $Y=2.525
+ $X2=0 $Y2=0
cc_517 N_A_851_242#_c_586_n N_A_881_463#_c_1078_n 0.00266134f $X=4.46 $Y=1.88
+ $X2=0 $Y2=0
cc_518 N_A_851_242#_c_577_n N_A_881_463#_c_1078_n 0.015564f $X=4.56 $Y=1.295
+ $X2=0 $Y2=0
cc_519 N_A_851_242#_c_571_n N_A_881_463#_c_1073_n 0.0296395f $X=5.375 $Y=1.295
+ $X2=0 $Y2=0
cc_520 N_A_851_242#_c_572_n N_A_881_463#_c_1073_n 8.74157e-19 $X=4.705 $Y=1.295
+ $X2=0 $Y2=0
cc_521 N_A_851_242#_c_574_n N_A_881_463#_c_1073_n 7.16574e-19 $X=5.665 $Y=1.295
+ $X2=0 $Y2=0
cc_522 N_A_851_242#_c_577_n N_A_881_463#_c_1073_n 0.0115618f $X=4.56 $Y=1.295
+ $X2=0 $Y2=0
cc_523 N_A_851_242#_c_580_n N_A_881_463#_c_1073_n 8.25632e-19 $X=4.5 $Y=1.375
+ $X2=0 $Y2=0
cc_524 N_A_851_242#_c_581_n N_A_881_463#_c_1073_n 8.89831e-19 $X=5.48 $Y=1.29
+ $X2=0 $Y2=0
cc_525 N_A_851_242#_c_598_p N_A_881_463#_c_1073_n 0.0116531f $X=5.48 $Y=1.29
+ $X2=0 $Y2=0
cc_526 N_A_851_242#_c_567_n N_A_881_463#_c_1074_n 0.00914384f $X=7.62 $Y=1.17
+ $X2=0 $Y2=0
cc_527 N_A_851_242#_c_573_n N_A_881_463#_c_1074_n 0.00571686f $X=7.775 $Y=1.295
+ $X2=0 $Y2=0
cc_528 N_A_851_242#_c_583_n N_A_881_463#_c_1074_n 0.00187899f $X=8 $Y=1.17 $X2=0
+ $Y2=0
cc_529 N_A_851_242#_M1017_g N_A_975_255#_M1007_g 0.0200304f $X=4.33 $Y=2.525
+ $X2=0 $Y2=0
cc_530 N_A_851_242#_c_586_n N_A_975_255#_M1007_g 0.0193825f $X=4.46 $Y=1.88
+ $X2=0 $Y2=0
cc_531 N_A_851_242#_c_581_n N_A_975_255#_M1007_g 0.00117768f $X=5.48 $Y=1.29
+ $X2=0 $Y2=0
cc_532 N_A_851_242#_c_572_n N_A_975_255#_M1030_g 6.96361e-19 $X=4.705 $Y=1.295
+ $X2=0 $Y2=0
cc_533 N_A_851_242#_c_577_n N_A_975_255#_M1030_g 0.00134707f $X=4.56 $Y=1.295
+ $X2=0 $Y2=0
cc_534 N_A_851_242#_c_580_n N_A_975_255#_M1030_g 0.00300113f $X=4.5 $Y=1.375
+ $X2=0 $Y2=0
cc_535 N_A_851_242#_c_581_n N_A_975_255#_M1030_g 0.0193132f $X=5.48 $Y=1.29
+ $X2=0 $Y2=0
cc_536 N_A_851_242#_c_598_p N_A_975_255#_M1030_g 3.20873e-19 $X=5.48 $Y=1.29
+ $X2=0 $Y2=0
cc_537 N_A_851_242#_c_582_n N_A_975_255#_M1030_g 0.012421f $X=5.48 $Y=1.125
+ $X2=0 $Y2=0
cc_538 N_A_851_242#_M1013_g N_A_975_255#_c_1223_n 0.0131732f $X=8.235 $Y=2.875
+ $X2=0 $Y2=0
cc_539 N_A_851_242#_c_589_n N_A_975_255#_M1010_g 0.0131732f $X=8.375 $Y=2.22
+ $X2=0 $Y2=0
cc_540 N_A_851_242#_c_567_n N_A_975_255#_c_1209_n 0.00445223f $X=7.62 $Y=1.17
+ $X2=0 $Y2=0
cc_541 N_A_851_242#_c_568_n N_A_975_255#_M1006_g 0.00818034f $X=8.275 $Y=2.055
+ $X2=0 $Y2=0
cc_542 N_A_851_242#_c_569_n N_A_975_255#_M1006_g 0.00277117f $X=8.19 $Y=1.277
+ $X2=0 $Y2=0
cc_543 N_A_851_242#_c_575_n N_A_975_255#_M1006_g 0.0096129f $X=10.655 $Y=1.295
+ $X2=0 $Y2=0
cc_544 N_A_851_242#_c_583_n N_A_975_255#_M1006_g 0.0212212f $X=8 $Y=1.17 $X2=0
+ $Y2=0
cc_545 N_A_851_242#_c_570_n N_A_975_255#_M1031_g 0.00580232f $X=10.83 $Y=1.06
+ $X2=0 $Y2=0
cc_546 N_A_851_242#_c_578_n N_A_975_255#_M1031_g 0.00679501f $X=10.8 $Y=1.295
+ $X2=0 $Y2=0
cc_547 N_A_851_242#_c_579_n N_A_975_255#_M1031_g 0.0182722f $X=10.8 $Y=1.295
+ $X2=0 $Y2=0
cc_548 N_A_851_242#_c_577_n N_A_975_255#_c_1212_n 7.23768e-19 $X=4.56 $Y=1.295
+ $X2=0 $Y2=0
cc_549 N_A_851_242#_c_580_n N_A_975_255#_c_1212_n 0.0193825f $X=4.5 $Y=1.375
+ $X2=0 $Y2=0
cc_550 N_A_851_242#_c_575_n N_A_975_255#_c_1213_n 0.0278818f $X=10.655 $Y=1.295
+ $X2=0 $Y2=0
cc_551 N_A_851_242#_c_579_n N_A_975_255#_c_1213_n 0.0105538f $X=10.8 $Y=1.295
+ $X2=0 $Y2=0
cc_552 N_A_851_242#_c_579_n N_A_975_255#_c_1229_n 0.0233337f $X=10.8 $Y=1.295
+ $X2=0 $Y2=0
cc_553 N_A_851_242#_M1004_s N_A_975_255#_c_1230_n 0.00742021f $X=10.7 $Y=1.835
+ $X2=0 $Y2=0
cc_554 N_A_851_242#_c_579_n N_A_975_255#_c_1230_n 0.0193617f $X=10.8 $Y=1.295
+ $X2=0 $Y2=0
cc_555 N_A_851_242#_c_578_n N_A_975_255#_c_1214_n 0.00203673f $X=10.8 $Y=1.295
+ $X2=0 $Y2=0
cc_556 N_A_851_242#_c_579_n N_A_975_255#_c_1214_n 0.0263461f $X=10.8 $Y=1.295
+ $X2=0 $Y2=0
cc_557 N_A_851_242#_c_579_n N_A_975_255#_c_1232_n 0.0222565f $X=10.8 $Y=1.295
+ $X2=0 $Y2=0
cc_558 N_A_851_242#_c_575_n N_A_975_255#_c_1217_n 0.00595381f $X=10.655 $Y=1.295
+ $X2=0 $Y2=0
cc_559 N_A_851_242#_c_568_n N_A_975_255#_c_1218_n 0.0247471f $X=8.275 $Y=2.055
+ $X2=0 $Y2=0
cc_560 N_A_851_242#_c_588_n N_A_975_255#_c_1218_n 5.59489e-19 $X=8.375 $Y=2.22
+ $X2=0 $Y2=0
cc_561 N_A_851_242#_c_575_n N_A_975_255#_c_1218_n 0.00701373f $X=10.655 $Y=1.295
+ $X2=0 $Y2=0
cc_562 N_A_851_242#_c_566_n N_A_975_255#_c_1238_n 0.00411426f $X=7.835 $Y=1.17
+ $X2=0 $Y2=0
cc_563 N_A_851_242#_c_568_n N_A_975_255#_c_1238_n 0.0118652f $X=8.275 $Y=2.055
+ $X2=0 $Y2=0
cc_564 N_A_851_242#_c_569_n N_A_975_255#_c_1238_n 0.002059f $X=8.19 $Y=1.277
+ $X2=0 $Y2=0
cc_565 N_A_851_242#_c_588_n N_A_975_255#_c_1238_n 0.00142254f $X=8.375 $Y=2.22
+ $X2=0 $Y2=0
cc_566 N_A_851_242#_c_589_n N_A_975_255#_c_1238_n 0.0221794f $X=8.375 $Y=2.22
+ $X2=0 $Y2=0
cc_567 N_A_851_242#_c_575_n N_A_975_255#_c_1238_n 3.04264e-19 $X=10.655 $Y=1.295
+ $X2=0 $Y2=0
cc_568 N_A_851_242#_c_576_n N_A_975_255#_c_1238_n 2.30471e-19 $X=8.065 $Y=1.295
+ $X2=0 $Y2=0
cc_569 N_A_851_242#_c_583_n N_A_975_255#_c_1238_n 0.0178191f $X=8 $Y=1.17 $X2=0
+ $Y2=0
cc_570 N_A_851_242#_c_579_n N_A_1524_69#_M1042_g 0.00132813f $X=10.8 $Y=1.295
+ $X2=0 $Y2=0
cc_571 N_A_851_242#_c_565_n N_A_1524_69#_c_1412_n 0.0041865f $X=7.545 $Y=1.095
+ $X2=0 $Y2=0
cc_572 N_A_851_242#_c_566_n N_A_1524_69#_c_1412_n 0.00583069f $X=7.835 $Y=1.17
+ $X2=0 $Y2=0
cc_573 N_A_851_242#_c_567_n N_A_1524_69#_c_1412_n 0.00470044f $X=7.62 $Y=1.17
+ $X2=0 $Y2=0
cc_574 N_A_851_242#_c_568_n N_A_1524_69#_c_1412_n 0.00549364f $X=8.275 $Y=2.055
+ $X2=0 $Y2=0
cc_575 N_A_851_242#_c_569_n N_A_1524_69#_c_1412_n 0.0126033f $X=8.19 $Y=1.277
+ $X2=0 $Y2=0
cc_576 N_A_851_242#_c_573_n N_A_1524_69#_c_1412_n 0.0164225f $X=7.775 $Y=1.295
+ $X2=0 $Y2=0
cc_577 N_A_851_242#_c_576_n N_A_1524_69#_c_1412_n 0.0027192f $X=8.065 $Y=1.295
+ $X2=0 $Y2=0
cc_578 N_A_851_242#_c_583_n N_A_1524_69#_c_1412_n 0.00120361f $X=8 $Y=1.17 $X2=0
+ $Y2=0
cc_579 N_A_851_242#_c_566_n N_A_1524_69#_c_1413_n 0.0126432f $X=7.835 $Y=1.17
+ $X2=0 $Y2=0
cc_580 N_A_851_242#_c_569_n N_A_1524_69#_c_1413_n 0.0287683f $X=8.19 $Y=1.277
+ $X2=0 $Y2=0
cc_581 N_A_851_242#_c_573_n N_A_1524_69#_c_1413_n 0.00305261f $X=7.775 $Y=1.295
+ $X2=0 $Y2=0
cc_582 N_A_851_242#_c_575_n N_A_1524_69#_c_1413_n 0.00911232f $X=10.655 $Y=1.295
+ $X2=0 $Y2=0
cc_583 N_A_851_242#_c_576_n N_A_1524_69#_c_1413_n 0.00360237f $X=8.065 $Y=1.295
+ $X2=0 $Y2=0
cc_584 N_A_851_242#_c_565_n N_A_1524_69#_c_1447_n 0.0113517f $X=7.545 $Y=1.095
+ $X2=0 $Y2=0
cc_585 N_A_851_242#_c_566_n N_A_1524_69#_c_1414_n 0.0014071f $X=7.835 $Y=1.17
+ $X2=0 $Y2=0
cc_586 N_A_851_242#_c_567_n N_A_1524_69#_c_1414_n 2.61905e-19 $X=7.62 $Y=1.17
+ $X2=0 $Y2=0
cc_587 N_A_851_242#_c_568_n N_A_1524_69#_c_1414_n 0.0133902f $X=8.275 $Y=2.055
+ $X2=0 $Y2=0
cc_588 N_A_851_242#_c_569_n N_A_1524_69#_c_1414_n 0.0108913f $X=8.19 $Y=1.277
+ $X2=0 $Y2=0
cc_589 N_A_851_242#_c_573_n N_A_1524_69#_c_1414_n 0.00441098f $X=7.775 $Y=1.295
+ $X2=0 $Y2=0
cc_590 N_A_851_242#_c_576_n N_A_1524_69#_c_1414_n 0.00657677f $X=8.065 $Y=1.295
+ $X2=0 $Y2=0
cc_591 N_A_851_242#_c_583_n N_A_1524_69#_c_1414_n 0.00114893f $X=8 $Y=1.17 $X2=0
+ $Y2=0
cc_592 N_A_851_242#_c_568_n N_A_1524_69#_c_1432_n 0.0245708f $X=8.275 $Y=2.055
+ $X2=0 $Y2=0
cc_593 N_A_851_242#_c_588_n N_A_1524_69#_c_1432_n 0.0199905f $X=8.375 $Y=2.22
+ $X2=0 $Y2=0
cc_594 N_A_851_242#_c_589_n N_A_1524_69#_c_1432_n 0.00743506f $X=8.375 $Y=2.22
+ $X2=0 $Y2=0
cc_595 N_A_851_242#_c_569_n N_A_1524_69#_c_1416_n 0.00984189f $X=8.19 $Y=1.277
+ $X2=0 $Y2=0
cc_596 N_A_851_242#_c_575_n N_A_1524_69#_c_1416_n 0.0120793f $X=10.655 $Y=1.295
+ $X2=0 $Y2=0
cc_597 N_A_851_242#_c_576_n N_A_1524_69#_c_1416_n 2.06729e-19 $X=8.065 $Y=1.295
+ $X2=0 $Y2=0
cc_598 N_A_851_242#_c_570_n N_A_1524_69#_c_1417_n 0.0129462f $X=10.83 $Y=1.06
+ $X2=0 $Y2=0
cc_599 N_A_851_242#_c_575_n N_A_1524_69#_c_1417_n 0.00124934f $X=10.655 $Y=1.295
+ $X2=0 $Y2=0
cc_600 N_A_851_242#_M1031_s N_A_1524_69#_c_1418_n 0.00719648f $X=10.685 $Y=0.345
+ $X2=0 $Y2=0
cc_601 N_A_851_242#_c_570_n N_A_1524_69#_c_1418_n 0.0208359f $X=10.83 $Y=1.06
+ $X2=0 $Y2=0
cc_602 N_A_851_242#_c_575_n N_A_1524_69#_c_1418_n 0.00596748f $X=10.655 $Y=1.295
+ $X2=0 $Y2=0
cc_603 N_A_851_242#_c_578_n N_A_1524_69#_c_1418_n 0.00160399f $X=10.8 $Y=1.295
+ $X2=0 $Y2=0
cc_604 N_A_851_242#_c_570_n N_A_1524_69#_c_1423_n 6.56351e-19 $X=10.83 $Y=1.06
+ $X2=0 $Y2=0
cc_605 N_A_851_242#_c_575_n N_A_1524_69#_c_1423_n 2.97663e-19 $X=10.655 $Y=1.295
+ $X2=0 $Y2=0
cc_606 N_A_851_242#_c_578_n N_A_1524_69#_c_1423_n 7.47514e-19 $X=10.8 $Y=1.295
+ $X2=0 $Y2=0
cc_607 N_A_851_242#_c_579_n N_A_1524_69#_c_1423_n 0.00407641f $X=10.8 $Y=1.295
+ $X2=0 $Y2=0
cc_608 N_A_851_242#_c_575_n N_A_1524_69#_c_1424_n 0.0480455f $X=10.655 $Y=1.295
+ $X2=0 $Y2=0
cc_609 N_A_851_242#_c_570_n N_A_1524_69#_c_1425_n 0.0170792f $X=10.83 $Y=1.06
+ $X2=0 $Y2=0
cc_610 N_A_851_242#_c_575_n N_A_1524_69#_c_1425_n 0.0447149f $X=10.655 $Y=1.295
+ $X2=0 $Y2=0
cc_611 N_A_851_242#_c_578_n N_A_1524_69#_c_1425_n 0.0016068f $X=10.8 $Y=1.295
+ $X2=0 $Y2=0
cc_612 N_A_851_242#_M1013_g N_A_1747_21#_M1028_g 0.022286f $X=8.235 $Y=2.875
+ $X2=0 $Y2=0
cc_613 N_A_851_242#_c_568_n N_A_1747_21#_c_1598_n 0.00222819f $X=8.275 $Y=2.055
+ $X2=0 $Y2=0
cc_614 N_A_851_242#_c_575_n N_A_1747_21#_c_1598_n 0.00194947f $X=10.655 $Y=1.295
+ $X2=0 $Y2=0
cc_615 N_A_851_242#_c_575_n N_A_1747_21#_c_1600_n 0.00205781f $X=10.655 $Y=1.295
+ $X2=0 $Y2=0
cc_616 N_A_851_242#_c_568_n N_A_1747_21#_c_1608_n 0.00513121f $X=8.275 $Y=2.055
+ $X2=0 $Y2=0
cc_617 N_A_851_242#_c_588_n N_A_1747_21#_c_1608_n 0.0131957f $X=8.375 $Y=2.22
+ $X2=0 $Y2=0
cc_618 N_A_851_242#_c_589_n N_A_1747_21#_c_1608_n 2.92986e-19 $X=8.375 $Y=2.22
+ $X2=0 $Y2=0
cc_619 N_A_851_242#_c_588_n N_A_1747_21#_c_1609_n 9.80769e-19 $X=8.375 $Y=2.22
+ $X2=0 $Y2=0
cc_620 N_A_851_242#_c_589_n N_A_1747_21#_c_1609_n 0.0219598f $X=8.375 $Y=2.22
+ $X2=0 $Y2=0
cc_621 N_A_851_242#_c_570_n N_CLK_M1011_g 8.50689e-19 $X=10.83 $Y=1.06 $X2=0
+ $Y2=0
cc_622 N_A_851_242#_M1013_g N_VPWR_c_1888_n 0.00386228f $X=8.235 $Y=2.875 $X2=0
+ $Y2=0
cc_623 N_A_851_242#_M1017_g N_VPWR_c_1892_n 0.00431487f $X=4.33 $Y=2.525 $X2=0
+ $Y2=0
cc_624 N_A_851_242#_M1004_s N_VPWR_c_1876_n 0.00397221f $X=10.7 $Y=1.835 $X2=0
+ $Y2=0
cc_625 N_A_851_242#_M1017_g N_VPWR_c_1876_n 0.00477801f $X=4.33 $Y=2.525 $X2=0
+ $Y2=0
cc_626 N_A_851_242#_M1013_g N_VPWR_c_1876_n 0.00625424f $X=8.235 $Y=2.875 $X2=0
+ $Y2=0
cc_627 N_A_851_242#_c_572_n N_A_372_50#_c_2058_n 0.00179861f $X=4.705 $Y=1.295
+ $X2=0 $Y2=0
cc_628 N_A_851_242#_c_577_n N_A_372_50#_c_2058_n 0.0571411f $X=4.56 $Y=1.295
+ $X2=0 $Y2=0
cc_629 N_A_851_242#_c_580_n N_A_372_50#_c_2058_n 0.0131254f $X=4.5 $Y=1.375
+ $X2=0 $Y2=0
cc_630 N_A_851_242#_c_571_n N_A_372_50#_c_2059_n 0.0053532f $X=5.375 $Y=1.295
+ $X2=0 $Y2=0
cc_631 N_A_851_242#_c_572_n N_A_372_50#_c_2059_n 0.00463079f $X=4.705 $Y=1.295
+ $X2=0 $Y2=0
cc_632 N_A_851_242#_c_577_n N_A_372_50#_c_2059_n 0.0194052f $X=4.56 $Y=1.295
+ $X2=0 $Y2=0
cc_633 N_A_851_242#_c_580_n N_A_372_50#_c_2059_n 0.0083561f $X=4.5 $Y=1.375
+ $X2=0 $Y2=0
cc_634 N_A_851_242#_M1017_g N_A_372_50#_c_2067_n 0.0057489f $X=4.33 $Y=2.525
+ $X2=0 $Y2=0
cc_635 N_A_851_242#_c_573_n N_VGND_c_2212_n 0.00244285f $X=7.775 $Y=1.295 $X2=0
+ $Y2=0
cc_636 N_A_851_242#_c_575_n N_VGND_c_2213_n 0.00227525f $X=10.655 $Y=1.295 $X2=0
+ $Y2=0
cc_637 N_A_851_242#_c_565_n N_VGND_c_2219_n 0.00329011f $X=7.545 $Y=1.095 $X2=0
+ $Y2=0
cc_638 N_A_851_242#_c_565_n N_VGND_c_2233_n 0.00504432f $X=7.545 $Y=1.095 $X2=0
+ $Y2=0
cc_639 N_A_851_242#_c_582_n N_VGND_c_2233_n 9.39239e-19 $X=5.48 $Y=1.125 $X2=0
+ $Y2=0
cc_640 N_A_1047_369#_M1045_g N_RESET_B_c_885_n 0.00999911f $X=5.93 $Y=0.805
+ $X2=0 $Y2=0
cc_641 N_A_1047_369#_c_780_n N_RESET_B_c_891_n 0.00331099f $X=7.105 $Y=1.64
+ $X2=0 $Y2=0
cc_642 N_A_1047_369#_c_782_n N_RESET_B_c_891_n 0.00103837f $X=6.04 $Y=1.76 $X2=0
+ $Y2=0
cc_643 N_A_1047_369#_M1003_g N_RESET_B_c_892_n 0.0156215f $X=5.31 $Y=2.525 $X2=0
+ $Y2=0
cc_644 N_A_1047_369#_c_785_n N_RESET_B_c_892_n 0.00924683f $X=5.855 $Y=1.74
+ $X2=0 $Y2=0
cc_645 N_A_1047_369#_c_790_n N_RESET_B_c_892_n 0.00103837f $X=5.87 $Y=1.76 $X2=0
+ $Y2=0
cc_646 N_A_1047_369#_c_786_n N_RESET_B_M1036_g 0.00186845f $X=5.595 $Y=1.74
+ $X2=0 $Y2=0
cc_647 N_A_1047_369#_M1045_g N_RESET_B_M1036_g 0.0828343f $X=5.93 $Y=0.805 $X2=0
+ $Y2=0
cc_648 N_A_1047_369#_c_780_n N_RESET_B_M1036_g 0.0119585f $X=7.105 $Y=1.64 $X2=0
+ $Y2=0
cc_649 N_A_1047_369#_c_782_n N_RESET_B_M1036_g 0.00495466f $X=6.04 $Y=1.76 $X2=0
+ $Y2=0
cc_650 N_A_1047_369#_M1022_d N_RESET_B_c_897_n 0.00262473f $X=7.26 $Y=1.895
+ $X2=0 $Y2=0
cc_651 N_A_1047_369#_c_780_n N_RESET_B_c_897_n 0.0158813f $X=7.105 $Y=1.64 $X2=0
+ $Y2=0
cc_652 N_A_1047_369#_c_783_n N_RESET_B_c_897_n 2.44208e-19 $X=7.21 $Y=1.64 $X2=0
+ $Y2=0
cc_653 N_A_1047_369#_c_812_n N_RESET_B_c_897_n 0.0147455f $X=7.4 $Y=2.02 $X2=0
+ $Y2=0
cc_654 N_A_1047_369#_M1022_d N_RESET_B_c_937_n 0.00309755f $X=7.26 $Y=1.895
+ $X2=0 $Y2=0
cc_655 N_A_1047_369#_M1022_d N_RESET_B_c_899_n 0.00224935f $X=7.26 $Y=1.895
+ $X2=0 $Y2=0
cc_656 N_A_1047_369#_c_812_n N_RESET_B_c_899_n 0.00378432f $X=7.4 $Y=2.02 $X2=0
+ $Y2=0
cc_657 N_A_1047_369#_c_780_n N_RESET_B_c_905_n 0.00463759f $X=7.105 $Y=1.64
+ $X2=0 $Y2=0
cc_658 N_A_1047_369#_c_789_n N_RESET_B_c_905_n 4.06718e-19 $X=7.215 $Y=1.9 $X2=0
+ $Y2=0
cc_659 N_A_1047_369#_c_782_n N_RESET_B_c_905_n 3.29608e-19 $X=6.04 $Y=1.76 $X2=0
+ $Y2=0
cc_660 N_A_1047_369#_c_812_n N_RESET_B_c_905_n 2.30182e-19 $X=7.4 $Y=2.02 $X2=0
+ $Y2=0
cc_661 N_A_1047_369#_c_786_n N_RESET_B_c_906_n 9.16824e-19 $X=5.595 $Y=1.74
+ $X2=0 $Y2=0
cc_662 N_A_1047_369#_c_780_n N_RESET_B_c_906_n 0.0258344f $X=7.105 $Y=1.64 $X2=0
+ $Y2=0
cc_663 N_A_1047_369#_c_782_n N_RESET_B_c_906_n 0.00609156f $X=6.04 $Y=1.76 $X2=0
+ $Y2=0
cc_664 N_A_1047_369#_c_812_n N_RESET_B_c_906_n 0.0073767f $X=7.4 $Y=2.02 $X2=0
+ $Y2=0
cc_665 N_A_1047_369#_c_781_n N_A_881_463#_M1015_g 0.0131981f $X=7.22 $Y=0.5
+ $X2=0 $Y2=0
cc_666 N_A_1047_369#_c_781_n N_A_881_463#_M1022_g 0.00422199f $X=7.22 $Y=0.5
+ $X2=0 $Y2=0
cc_667 N_A_1047_369#_c_789_n N_A_881_463#_M1022_g 0.00845198f $X=7.215 $Y=1.9
+ $X2=0 $Y2=0
cc_668 N_A_1047_369#_c_783_n N_A_881_463#_M1022_g 0.00825996f $X=7.21 $Y=1.64
+ $X2=0 $Y2=0
cc_669 N_A_1047_369#_c_812_n N_A_881_463#_M1022_g 0.00807902f $X=7.4 $Y=2.02
+ $X2=0 $Y2=0
cc_670 N_A_1047_369#_c_786_n N_A_881_463#_c_1068_n 0.00170818f $X=5.595 $Y=1.74
+ $X2=0 $Y2=0
cc_671 N_A_1047_369#_c_790_n N_A_881_463#_c_1068_n 0.0157193f $X=5.87 $Y=1.76
+ $X2=0 $Y2=0
cc_672 N_A_1047_369#_M1003_g N_A_881_463#_c_1077_n 0.0157734f $X=5.31 $Y=2.525
+ $X2=0 $Y2=0
cc_673 N_A_1047_369#_c_785_n N_A_881_463#_c_1077_n 0.00121672f $X=5.855 $Y=1.74
+ $X2=0 $Y2=0
cc_674 N_A_1047_369#_c_786_n N_A_881_463#_c_1077_n 0.00487723f $X=5.595 $Y=1.74
+ $X2=0 $Y2=0
cc_675 N_A_1047_369#_c_780_n N_A_881_463#_c_1077_n 0.00501688f $X=7.105 $Y=1.64
+ $X2=0 $Y2=0
cc_676 N_A_1047_369#_c_790_n N_A_881_463#_c_1077_n 0.0456033f $X=5.87 $Y=1.76
+ $X2=0 $Y2=0
cc_677 N_A_1047_369#_c_782_n N_A_881_463#_c_1077_n 0.0142423f $X=6.04 $Y=1.76
+ $X2=0 $Y2=0
cc_678 N_A_1047_369#_M1045_g N_A_881_463#_c_1095_n 0.0124188f $X=5.93 $Y=0.805
+ $X2=0 $Y2=0
cc_679 N_A_1047_369#_M1045_g N_A_881_463#_c_1070_n 0.00572527f $X=5.93 $Y=0.805
+ $X2=0 $Y2=0
cc_680 N_A_1047_369#_c_785_n N_A_881_463#_c_1071_n 0.00131004f $X=5.855 $Y=1.74
+ $X2=0 $Y2=0
cc_681 N_A_1047_369#_M1045_g N_A_881_463#_c_1071_n 0.0043062f $X=5.93 $Y=0.805
+ $X2=0 $Y2=0
cc_682 N_A_1047_369#_c_790_n N_A_881_463#_c_1071_n 0.00418019f $X=5.87 $Y=1.76
+ $X2=0 $Y2=0
cc_683 N_A_1047_369#_c_782_n N_A_881_463#_c_1071_n 0.00629751f $X=6.04 $Y=1.76
+ $X2=0 $Y2=0
cc_684 N_A_1047_369#_M1045_g N_A_881_463#_c_1072_n 0.00585292f $X=5.93 $Y=0.805
+ $X2=0 $Y2=0
cc_685 N_A_1047_369#_c_781_n N_A_881_463#_c_1072_n 0.0157023f $X=7.22 $Y=0.5
+ $X2=0 $Y2=0
cc_686 N_A_1047_369#_c_782_n N_A_881_463#_c_1072_n 0.066169f $X=6.04 $Y=1.76
+ $X2=0 $Y2=0
cc_687 N_A_1047_369#_c_780_n N_A_881_463#_c_1074_n 0.0151158f $X=7.105 $Y=1.64
+ $X2=0 $Y2=0
cc_688 N_A_1047_369#_c_781_n N_A_881_463#_c_1074_n 0.0113402f $X=7.22 $Y=0.5
+ $X2=0 $Y2=0
cc_689 N_A_1047_369#_c_786_n N_A_975_255#_M1007_g 0.0707164f $X=5.595 $Y=1.74
+ $X2=0 $Y2=0
cc_690 N_A_1047_369#_c_790_n N_A_975_255#_M1007_g 9.31864e-19 $X=5.87 $Y=1.76
+ $X2=0 $Y2=0
cc_691 N_A_1047_369#_M1003_g N_A_975_255#_c_1223_n 0.0103107f $X=5.31 $Y=2.525
+ $X2=0 $Y2=0
cc_692 N_A_1047_369#_c_812_n N_A_975_255#_M1010_g 0.00324311f $X=7.4 $Y=2.02
+ $X2=0 $Y2=0
cc_693 N_A_1047_369#_c_789_n N_A_975_255#_c_1209_n 0.00137554f $X=7.215 $Y=1.9
+ $X2=0 $Y2=0
cc_694 N_A_1047_369#_c_783_n N_A_975_255#_c_1209_n 3.14285e-19 $X=7.21 $Y=1.64
+ $X2=0 $Y2=0
cc_695 N_A_1047_369#_c_781_n N_A_1524_69#_c_1412_n 0.044314f $X=7.22 $Y=0.5
+ $X2=0 $Y2=0
cc_696 N_A_1047_369#_c_783_n N_A_1524_69#_c_1412_n 4.22248e-19 $X=7.21 $Y=1.64
+ $X2=0 $Y2=0
cc_697 N_A_1047_369#_c_781_n N_A_1524_69#_c_1447_n 0.0438751f $X=7.22 $Y=0.5
+ $X2=0 $Y2=0
cc_698 N_A_1047_369#_c_783_n N_A_1524_69#_c_1414_n 0.015091f $X=7.21 $Y=1.64
+ $X2=0 $Y2=0
cc_699 N_A_1047_369#_c_812_n N_A_1524_69#_c_1414_n 0.00370879f $X=7.4 $Y=2.02
+ $X2=0 $Y2=0
cc_700 N_A_1047_369#_c_789_n N_A_1524_69#_c_1432_n 0.00658961f $X=7.215 $Y=1.9
+ $X2=0 $Y2=0
cc_701 N_A_1047_369#_M1003_g N_VPWR_c_1879_n 0.00907365f $X=5.31 $Y=2.525 $X2=0
+ $Y2=0
cc_702 N_A_1047_369#_M1003_g N_VPWR_c_1876_n 7.88961e-19 $X=5.31 $Y=2.525 $X2=0
+ $Y2=0
cc_703 N_A_1047_369#_c_781_n N_VGND_c_2212_n 0.0307994f $X=7.22 $Y=0.5 $X2=0
+ $Y2=0
cc_704 N_A_1047_369#_c_781_n N_VGND_c_2219_n 0.00987454f $X=7.22 $Y=0.5 $X2=0
+ $Y2=0
cc_705 N_A_1047_369#_M1045_g N_VGND_c_2233_n 9.39239e-19 $X=5.93 $Y=0.805 $X2=0
+ $Y2=0
cc_706 N_A_1047_369#_c_781_n N_VGND_c_2233_n 0.00775071f $X=7.22 $Y=0.5 $X2=0
+ $Y2=0
cc_707 N_RESET_B_c_885_n N_A_881_463#_M1015_g 0.017097f $X=6.215 $Y=0.18 $X2=0
+ $Y2=0
cc_708 N_RESET_B_c_896_n N_A_881_463#_M1022_g 0.00300243f $X=6.495 $Y=2.285
+ $X2=0 $Y2=0
cc_709 N_RESET_B_c_897_n N_A_881_463#_M1022_g 0.011299f $X=7.2 $Y=2.37 $X2=0
+ $Y2=0
cc_710 N_RESET_B_c_937_n N_A_881_463#_M1022_g 0.0103295f $X=7.285 $Y=2.725 $X2=0
+ $Y2=0
cc_711 N_RESET_B_c_900_n N_A_881_463#_M1022_g 0.00363939f $X=7.37 $Y=2.81 $X2=0
+ $Y2=0
cc_712 N_RESET_B_c_905_n N_A_881_463#_M1022_g 0.00657128f $X=6.385 $Y=1.99 $X2=0
+ $Y2=0
cc_713 N_RESET_B_c_906_n N_A_881_463#_M1022_g 0.00185104f $X=6.495 $Y=2.012
+ $X2=0 $Y2=0
cc_714 N_RESET_B_c_890_n N_A_881_463#_c_1077_n 0.0162587f $X=5.91 $Y=2.205 $X2=0
+ $Y2=0
cc_715 N_RESET_B_c_891_n N_A_881_463#_c_1077_n 0.00858899f $X=6.215 $Y=2.13
+ $X2=0 $Y2=0
cc_716 N_RESET_B_c_892_n N_A_881_463#_c_1077_n 0.00313482f $X=5.985 $Y=2.13
+ $X2=0 $Y2=0
cc_717 N_RESET_B_c_896_n N_A_881_463#_c_1077_n 0.00676296f $X=6.495 $Y=2.285
+ $X2=0 $Y2=0
cc_718 N_RESET_B_c_898_n N_A_881_463#_c_1077_n 0.0111496f $X=6.58 $Y=2.37 $X2=0
+ $Y2=0
cc_719 N_RESET_B_c_906_n N_A_881_463#_c_1077_n 0.00178039f $X=6.495 $Y=2.012
+ $X2=0 $Y2=0
cc_720 N_RESET_B_c_885_n N_A_881_463#_c_1095_n 0.00877968f $X=6.215 $Y=0.18
+ $X2=0 $Y2=0
cc_721 N_RESET_B_M1036_g N_A_881_463#_c_1095_n 0.00102243f $X=6.29 $Y=0.805
+ $X2=0 $Y2=0
cc_722 N_RESET_B_c_885_n N_A_881_463#_c_1161_n 0.00192855f $X=6.215 $Y=0.18
+ $X2=0 $Y2=0
cc_723 N_RESET_B_M1036_g N_A_881_463#_c_1070_n 0.00114026f $X=6.29 $Y=0.805
+ $X2=0 $Y2=0
cc_724 N_RESET_B_M1036_g N_A_881_463#_c_1072_n 0.0161629f $X=6.29 $Y=0.805 $X2=0
+ $Y2=0
cc_725 N_RESET_B_M1033_g N_A_881_463#_c_1078_n 2.12412e-19 $X=3.805 $Y=2.635
+ $X2=0 $Y2=0
cc_726 N_RESET_B_M1036_g N_A_881_463#_c_1074_n 0.0190872f $X=6.29 $Y=0.805 $X2=0
+ $Y2=0
cc_727 N_RESET_B_c_885_n N_A_975_255#_M1030_g 0.010166f $X=6.215 $Y=0.18 $X2=0
+ $Y2=0
cc_728 N_RESET_B_c_890_n N_A_975_255#_c_1223_n 0.00993652f $X=5.91 $Y=2.205
+ $X2=0 $Y2=0
cc_729 N_RESET_B_c_897_n N_A_975_255#_c_1223_n 0.00492349f $X=7.2 $Y=2.37 $X2=0
+ $Y2=0
cc_730 N_RESET_B_c_898_n N_A_975_255#_c_1223_n 0.00396108f $X=6.58 $Y=2.37 $X2=0
+ $Y2=0
cc_731 N_RESET_B_c_899_n N_A_975_255#_c_1223_n 0.0016622f $X=8.19 $Y=2.81 $X2=0
+ $Y2=0
cc_732 N_RESET_B_c_900_n N_A_975_255#_c_1223_n 0.0029302f $X=7.37 $Y=2.81 $X2=0
+ $Y2=0
cc_733 N_RESET_B_c_897_n N_A_975_255#_M1010_g 0.00159845f $X=7.2 $Y=2.37 $X2=0
+ $Y2=0
cc_734 N_RESET_B_c_937_n N_A_975_255#_M1010_g 0.00439243f $X=7.285 $Y=2.725
+ $X2=0 $Y2=0
cc_735 N_RESET_B_c_899_n N_A_975_255#_M1010_g 0.0160783f $X=8.19 $Y=2.81 $X2=0
+ $Y2=0
cc_736 N_RESET_B_c_902_n N_A_975_255#_M1010_g 0.00105611f $X=8.275 $Y=2.57 $X2=0
+ $Y2=0
cc_737 N_RESET_B_M1026_g N_A_975_255#_c_1213_n 0.01091f $X=9.435 $Y=0.805 $X2=0
+ $Y2=0
cc_738 N_RESET_B_c_901_n N_A_975_255#_c_1217_n 0.003266f $X=9.36 $Y=2.57 $X2=0
+ $Y2=0
cc_739 N_RESET_B_c_901_n N_A_975_255#_c_1218_n 0.00644019f $X=9.36 $Y=2.57 $X2=0
+ $Y2=0
cc_740 N_RESET_B_c_899_n N_A_1524_69#_M1010_d 0.0111852f $X=8.19 $Y=2.81 $X2=0
+ $Y2=0
cc_741 N_RESET_B_M1026_g N_A_1524_69#_M1042_g 0.0229853f $X=9.435 $Y=0.805 $X2=0
+ $Y2=0
cc_742 N_RESET_B_M1018_g N_A_1524_69#_M1042_g 0.0169837f $X=9.545 $Y=2.875 $X2=0
+ $Y2=0
cc_743 N_RESET_B_c_903_n N_A_1524_69#_M1042_g 8.09313e-19 $X=9.525 $Y=2.34 $X2=0
+ $Y2=0
cc_744 N_RESET_B_c_904_n N_A_1524_69#_M1042_g 0.0205745f $X=9.525 $Y=2.34 $X2=0
+ $Y2=0
cc_745 N_RESET_B_c_899_n N_A_1524_69#_c_1432_n 0.0203787f $X=8.19 $Y=2.81 $X2=0
+ $Y2=0
cc_746 N_RESET_B_c_902_n N_A_1524_69#_c_1432_n 0.00438751f $X=8.275 $Y=2.57
+ $X2=0 $Y2=0
cc_747 N_RESET_B_M1026_g N_A_1524_69#_c_1424_n 0.0134562f $X=9.435 $Y=0.805
+ $X2=0 $Y2=0
cc_748 N_RESET_B_M1026_g N_A_1524_69#_c_1425_n 7.53791e-19 $X=9.435 $Y=0.805
+ $X2=0 $Y2=0
cc_749 N_RESET_B_M1026_g N_A_1524_69#_c_1427_n 0.0612574f $X=9.435 $Y=0.805
+ $X2=0 $Y2=0
cc_750 N_RESET_B_M1026_g N_A_1747_21#_M1039_g 0.00890808f $X=9.435 $Y=0.805
+ $X2=0 $Y2=0
cc_751 N_RESET_B_M1018_g N_A_1747_21#_M1028_g 0.0125287f $X=9.545 $Y=2.875 $X2=0
+ $Y2=0
cc_752 N_RESET_B_c_901_n N_A_1747_21#_M1028_g 0.014655f $X=9.36 $Y=2.57 $X2=0
+ $Y2=0
cc_753 N_RESET_B_c_902_n N_A_1747_21#_M1028_g 0.00105702f $X=8.275 $Y=2.57 $X2=0
+ $Y2=0
cc_754 N_RESET_B_c_903_n N_A_1747_21#_M1028_g 6.75833e-19 $X=9.525 $Y=2.34 $X2=0
+ $Y2=0
cc_755 N_RESET_B_c_904_n N_A_1747_21#_M1028_g 0.00330484f $X=9.525 $Y=2.34 $X2=0
+ $Y2=0
cc_756 N_RESET_B_M1026_g N_A_1747_21#_c_1596_n 0.0104164f $X=9.435 $Y=0.805
+ $X2=0 $Y2=0
cc_757 N_RESET_B_c_904_n N_A_1747_21#_c_1598_n 0.0416982f $X=9.525 $Y=2.34 $X2=0
+ $Y2=0
cc_758 N_RESET_B_M1026_g N_A_1747_21#_c_1599_n 0.0416982f $X=9.435 $Y=0.805
+ $X2=0 $Y2=0
cc_759 N_RESET_B_M1026_g N_A_1747_21#_c_1606_n 0.0105429f $X=9.435 $Y=0.805
+ $X2=0 $Y2=0
cc_760 N_RESET_B_c_901_n N_A_1747_21#_c_1606_n 0.00858789f $X=9.36 $Y=2.57 $X2=0
+ $Y2=0
cc_761 N_RESET_B_c_903_n N_A_1747_21#_c_1606_n 0.02463f $X=9.525 $Y=2.34 $X2=0
+ $Y2=0
cc_762 N_RESET_B_c_904_n N_A_1747_21#_c_1606_n 0.00486514f $X=9.525 $Y=2.34
+ $X2=0 $Y2=0
cc_763 N_RESET_B_M1018_g N_A_1747_21#_c_1632_n 0.00334005f $X=9.545 $Y=2.875
+ $X2=0 $Y2=0
cc_764 N_RESET_B_c_903_n N_A_1747_21#_c_1632_n 0.0049086f $X=9.525 $Y=2.34 $X2=0
+ $Y2=0
cc_765 N_RESET_B_c_904_n N_A_1747_21#_c_1632_n 2.44495e-19 $X=9.525 $Y=2.34
+ $X2=0 $Y2=0
cc_766 N_RESET_B_M1026_g N_A_1747_21#_c_1600_n 0.00143721f $X=9.435 $Y=0.805
+ $X2=0 $Y2=0
cc_767 N_RESET_B_M1026_g N_A_1747_21#_c_1607_n 0.00171438f $X=9.435 $Y=0.805
+ $X2=0 $Y2=0
cc_768 N_RESET_B_M1018_g N_A_1747_21#_c_1607_n 8.05544e-19 $X=9.545 $Y=2.875
+ $X2=0 $Y2=0
cc_769 N_RESET_B_c_903_n N_A_1747_21#_c_1607_n 0.0301364f $X=9.525 $Y=2.34 $X2=0
+ $Y2=0
cc_770 N_RESET_B_c_904_n N_A_1747_21#_c_1607_n 0.0027865f $X=9.525 $Y=2.34 $X2=0
+ $Y2=0
cc_771 N_RESET_B_M1026_g N_A_1747_21#_c_1608_n 0.00141084f $X=9.435 $Y=0.805
+ $X2=0 $Y2=0
cc_772 N_RESET_B_c_901_n N_A_1747_21#_c_1608_n 0.0246233f $X=9.36 $Y=2.57 $X2=0
+ $Y2=0
cc_773 N_RESET_B_c_903_n N_A_1747_21#_c_1608_n 0.00445513f $X=9.525 $Y=2.34
+ $X2=0 $Y2=0
cc_774 N_RESET_B_c_901_n N_A_1747_21#_c_1609_n 0.00672284f $X=9.36 $Y=2.57 $X2=0
+ $Y2=0
cc_775 N_RESET_B_c_903_n N_A_1747_21#_c_1609_n 5.96631e-19 $X=9.525 $Y=2.34
+ $X2=0 $Y2=0
cc_776 N_RESET_B_c_897_n N_VPWR_M1022_s 0.0121162f $X=7.2 $Y=2.37 $X2=0 $Y2=0
cc_777 N_RESET_B_M1033_g N_VPWR_c_1878_n 0.00573692f $X=3.805 $Y=2.635 $X2=0
+ $Y2=0
cc_778 N_RESET_B_c_890_n N_VPWR_c_1879_n 0.00638698f $X=5.91 $Y=2.205 $X2=0
+ $Y2=0
cc_779 N_RESET_B_c_897_n N_VPWR_c_1880_n 0.0267445f $X=7.2 $Y=2.37 $X2=0 $Y2=0
cc_780 N_RESET_B_c_937_n N_VPWR_c_1880_n 0.00704815f $X=7.285 $Y=2.725 $X2=0
+ $Y2=0
cc_781 N_RESET_B_c_900_n N_VPWR_c_1880_n 0.0137815f $X=7.37 $Y=2.81 $X2=0 $Y2=0
cc_782 N_RESET_B_M1018_g N_VPWR_c_1881_n 0.00619053f $X=9.545 $Y=2.875 $X2=0
+ $Y2=0
cc_783 N_RESET_B_c_901_n N_VPWR_c_1881_n 0.0257073f $X=9.36 $Y=2.57 $X2=0 $Y2=0
cc_784 N_RESET_B_c_899_n N_VPWR_c_1888_n 0.0232601f $X=8.19 $Y=2.81 $X2=0 $Y2=0
cc_785 N_RESET_B_c_900_n N_VPWR_c_1888_n 0.00559239f $X=7.37 $Y=2.81 $X2=0 $Y2=0
cc_786 N_RESET_B_c_901_n N_VPWR_c_1888_n 0.010534f $X=9.36 $Y=2.57 $X2=0 $Y2=0
cc_787 N_RESET_B_c_902_n N_VPWR_c_1888_n 0.00435918f $X=8.275 $Y=2.57 $X2=0
+ $Y2=0
cc_788 N_RESET_B_M1033_g N_VPWR_c_1892_n 0.00431995f $X=3.805 $Y=2.635 $X2=0
+ $Y2=0
cc_789 N_RESET_B_M1018_g N_VPWR_c_1894_n 0.00411452f $X=9.545 $Y=2.875 $X2=0
+ $Y2=0
cc_790 N_RESET_B_c_901_n N_VPWR_c_1894_n 4.10716e-19 $X=9.36 $Y=2.57 $X2=0 $Y2=0
cc_791 N_RESET_B_c_903_n N_VPWR_c_1894_n 0.00393618f $X=9.525 $Y=2.34 $X2=0
+ $Y2=0
cc_792 N_RESET_B_M1033_g N_VPWR_c_1876_n 0.00544287f $X=3.805 $Y=2.635 $X2=0
+ $Y2=0
cc_793 N_RESET_B_c_890_n N_VPWR_c_1876_n 9.39239e-19 $X=5.91 $Y=2.205 $X2=0
+ $Y2=0
cc_794 N_RESET_B_M1018_g N_VPWR_c_1876_n 0.00648382f $X=9.545 $Y=2.875 $X2=0
+ $Y2=0
cc_795 N_RESET_B_c_899_n N_VPWR_c_1876_n 0.0256962f $X=8.19 $Y=2.81 $X2=0 $Y2=0
cc_796 N_RESET_B_c_900_n N_VPWR_c_1876_n 0.00524087f $X=7.37 $Y=2.81 $X2=0 $Y2=0
cc_797 N_RESET_B_c_901_n N_VPWR_c_1876_n 0.0192559f $X=9.36 $Y=2.57 $X2=0 $Y2=0
cc_798 N_RESET_B_c_902_n N_VPWR_c_1876_n 0.00517715f $X=8.275 $Y=2.57 $X2=0
+ $Y2=0
cc_799 N_RESET_B_c_903_n N_VPWR_c_1876_n 0.00629104f $X=9.525 $Y=2.34 $X2=0
+ $Y2=0
cc_800 N_RESET_B_M1033_g N_A_372_50#_c_2064_n 0.00703491f $X=3.805 $Y=2.635
+ $X2=0 $Y2=0
cc_801 N_RESET_B_M1001_g N_A_372_50#_c_2057_n 0.00958959f $X=3.235 $Y=0.615
+ $X2=0 $Y2=0
cc_802 N_RESET_B_c_882_n N_A_372_50#_c_2057_n 0.00114357f $X=3.73 $Y=0.18 $X2=0
+ $Y2=0
cc_803 N_RESET_B_M1033_g N_A_372_50#_c_2057_n 0.00869271f $X=3.805 $Y=2.635
+ $X2=0 $Y2=0
cc_804 N_RESET_B_M1033_g N_A_372_50#_c_2058_n 0.0485487f $X=3.805 $Y=2.635 $X2=0
+ $Y2=0
cc_805 N_RESET_B_c_885_n N_A_372_50#_c_2059_n 0.0117311f $X=6.215 $Y=0.18 $X2=0
+ $Y2=0
cc_806 N_RESET_B_M1001_g N_A_372_50#_c_2062_n 0.0024097f $X=3.235 $Y=0.615 $X2=0
+ $Y2=0
cc_807 N_RESET_B_M1001_g N_A_372_50#_c_2063_n 8.03796e-19 $X=3.235 $Y=0.615
+ $X2=0 $Y2=0
cc_808 N_RESET_B_M1033_g N_A_372_50#_c_2063_n 0.0198806f $X=3.805 $Y=2.635 $X2=0
+ $Y2=0
cc_809 N_RESET_B_c_885_n N_A_372_50#_c_2063_n 0.00511773f $X=6.215 $Y=0.18 $X2=0
+ $Y2=0
cc_810 N_RESET_B_M1033_g N_A_372_50#_c_2067_n 0.0105004f $X=3.805 $Y=2.635 $X2=0
+ $Y2=0
cc_811 N_RESET_B_M1001_g N_VGND_c_2210_n 0.00137133f $X=3.235 $Y=0.615 $X2=0
+ $Y2=0
cc_812 N_RESET_B_c_882_n N_VGND_c_2210_n 0.0201786f $X=3.73 $Y=0.18 $X2=0 $Y2=0
cc_813 N_RESET_B_M1033_g N_VGND_c_2210_n 0.0105224f $X=3.805 $Y=2.635 $X2=0
+ $Y2=0
cc_814 N_RESET_B_c_882_n N_VGND_c_2211_n 0.0778328f $X=3.73 $Y=0.18 $X2=0 $Y2=0
cc_815 N_RESET_B_c_885_n N_VGND_c_2212_n 0.0214596f $X=6.215 $Y=0.18 $X2=0 $Y2=0
cc_816 N_RESET_B_M1026_g N_VGND_c_2213_n 0.00748219f $X=9.435 $Y=0.805 $X2=0
+ $Y2=0
cc_817 N_RESET_B_c_883_n N_VGND_c_2222_n 0.00720663f $X=3.31 $Y=0.18 $X2=0 $Y2=0
cc_818 N_RESET_B_c_882_n N_VGND_c_2233_n 0.00927548f $X=3.73 $Y=0.18 $X2=0 $Y2=0
cc_819 N_RESET_B_c_883_n N_VGND_c_2233_n 0.010567f $X=3.31 $Y=0.18 $X2=0 $Y2=0
cc_820 N_RESET_B_c_885_n N_VGND_c_2233_n 0.0834297f $X=6.215 $Y=0.18 $X2=0 $Y2=0
cc_821 N_RESET_B_M1026_g N_VGND_c_2233_n 9.39239e-19 $X=9.435 $Y=0.805 $X2=0
+ $Y2=0
cc_822 N_RESET_B_c_888_n N_VGND_c_2233_n 0.00613456f $X=3.805 $Y=0.18 $X2=0
+ $Y2=0
cc_823 N_RESET_B_M1001_g N_noxref_24_c_2369_n 0.00630151f $X=3.235 $Y=0.615
+ $X2=0 $Y2=0
cc_824 N_RESET_B_c_883_n N_noxref_24_c_2369_n 2.05582e-19 $X=3.31 $Y=0.18 $X2=0
+ $Y2=0
cc_825 N_A_881_463#_c_1068_n N_A_975_255#_M1007_g 0.0239716f $X=4.905 $Y=2.135
+ $X2=0 $Y2=0
cc_826 N_A_881_463#_c_1077_n N_A_975_255#_M1007_g 0.00452892f $X=5.87 $Y=2.22
+ $X2=0 $Y2=0
cc_827 N_A_881_463#_c_1078_n N_A_975_255#_M1007_g 0.0146647f $X=4.7 $Y=2.22
+ $X2=0 $Y2=0
cc_828 N_A_881_463#_c_1069_n N_A_975_255#_M1030_g 0.0104021f $X=5.13 $Y=1.21
+ $X2=0 $Y2=0
cc_829 N_A_881_463#_c_1161_n N_A_975_255#_M1030_g 0.0050139f $X=5.215 $Y=0.797
+ $X2=0 $Y2=0
cc_830 N_A_881_463#_c_1073_n N_A_975_255#_M1030_g 0.00585847f $X=5.13 $Y=1.295
+ $X2=0 $Y2=0
cc_831 N_A_881_463#_M1022_g N_A_975_255#_c_1223_n 0.00961975f $X=7.185 $Y=2.315
+ $X2=0 $Y2=0
cc_832 N_A_881_463#_c_1077_n N_A_975_255#_c_1223_n 0.00469715f $X=5.87 $Y=2.22
+ $X2=0 $Y2=0
cc_833 N_A_881_463#_M1022_g N_A_975_255#_c_1209_n 0.0388643f $X=7.185 $Y=2.315
+ $X2=0 $Y2=0
cc_834 N_A_881_463#_c_1068_n N_A_975_255#_c_1212_n 0.0015413f $X=4.905 $Y=2.135
+ $X2=0 $Y2=0
cc_835 N_A_881_463#_c_1073_n N_A_975_255#_c_1212_n 0.00900183f $X=5.13 $Y=1.295
+ $X2=0 $Y2=0
cc_836 N_A_881_463#_c_1074_n N_A_1524_69#_c_1412_n 0.00121091f $X=6.91 $Y=1.29
+ $X2=0 $Y2=0
cc_837 N_A_881_463#_M1022_g N_A_1524_69#_c_1414_n 8.89602e-19 $X=7.185 $Y=2.315
+ $X2=0 $Y2=0
cc_838 N_A_881_463#_c_1077_n N_VPWR_c_1879_n 0.0421468f $X=5.87 $Y=2.22 $X2=0
+ $Y2=0
cc_839 N_A_881_463#_c_1078_n N_VPWR_c_1879_n 0.00517766f $X=4.7 $Y=2.22 $X2=0
+ $Y2=0
cc_840 N_A_881_463#_M1022_g N_VPWR_c_1880_n 0.00518229f $X=7.185 $Y=2.315 $X2=0
+ $Y2=0
cc_841 N_A_881_463#_c_1077_n N_VPWR_c_1880_n 0.00267942f $X=5.87 $Y=2.22 $X2=0
+ $Y2=0
cc_842 N_A_881_463#_c_1078_n N_VPWR_c_1892_n 0.0100972f $X=4.7 $Y=2.22 $X2=0
+ $Y2=0
cc_843 N_A_881_463#_c_1077_n N_VPWR_c_1893_n 0.00613787f $X=5.87 $Y=2.22 $X2=0
+ $Y2=0
cc_844 N_A_881_463#_M1022_g N_VPWR_c_1876_n 5.63543e-19 $X=7.185 $Y=2.315 $X2=0
+ $Y2=0
cc_845 N_A_881_463#_c_1077_n N_VPWR_c_1876_n 0.00932806f $X=5.87 $Y=2.22 $X2=0
+ $Y2=0
cc_846 N_A_881_463#_c_1078_n N_VPWR_c_1876_n 0.0134762f $X=4.7 $Y=2.22 $X2=0
+ $Y2=0
cc_847 N_A_881_463#_c_1068_n N_A_372_50#_c_2058_n 0.00878037f $X=4.905 $Y=2.135
+ $X2=0 $Y2=0
cc_848 N_A_881_463#_c_1078_n N_A_372_50#_c_2058_n 0.0137131f $X=4.7 $Y=2.22
+ $X2=0 $Y2=0
cc_849 N_A_881_463#_c_1069_n N_A_372_50#_c_2059_n 0.00107097f $X=5.13 $Y=1.21
+ $X2=0 $Y2=0
cc_850 N_A_881_463#_c_1161_n N_A_372_50#_c_2059_n 0.0274446f $X=5.215 $Y=0.797
+ $X2=0 $Y2=0
cc_851 N_A_881_463#_c_1073_n N_A_372_50#_c_2059_n 0.00314501f $X=5.13 $Y=1.295
+ $X2=0 $Y2=0
cc_852 N_A_881_463#_c_1078_n N_A_372_50#_c_2067_n 0.0214076f $X=4.7 $Y=2.22
+ $X2=0 $Y2=0
cc_853 N_A_881_463#_c_1095_n N_VGND_c_2211_n 0.0116733f $X=5.785 $Y=0.797 $X2=0
+ $Y2=0
cc_854 N_A_881_463#_c_1161_n N_VGND_c_2211_n 0.0025919f $X=5.215 $Y=0.797 $X2=0
+ $Y2=0
cc_855 N_A_881_463#_M1015_g N_VGND_c_2212_n 0.011301f $X=6.91 $Y=0.665 $X2=0
+ $Y2=0
cc_856 N_A_881_463#_c_1095_n N_VGND_c_2212_n 0.0115333f $X=5.785 $Y=0.797 $X2=0
+ $Y2=0
cc_857 N_A_881_463#_c_1070_n N_VGND_c_2212_n 0.00130941f $X=5.87 $Y=1.165 $X2=0
+ $Y2=0
cc_858 N_A_881_463#_c_1072_n N_VGND_c_2212_n 0.0246366f $X=6.77 $Y=1.29 $X2=0
+ $Y2=0
cc_859 N_A_881_463#_c_1074_n N_VGND_c_2212_n 0.00388739f $X=6.91 $Y=1.29 $X2=0
+ $Y2=0
cc_860 N_A_881_463#_M1015_g N_VGND_c_2219_n 0.00482246f $X=6.91 $Y=0.665 $X2=0
+ $Y2=0
cc_861 N_A_881_463#_M1015_g N_VGND_c_2233_n 0.00970391f $X=6.91 $Y=0.665 $X2=0
+ $Y2=0
cc_862 N_A_881_463#_c_1095_n N_VGND_c_2233_n 0.0185493f $X=5.785 $Y=0.797 $X2=0
+ $Y2=0
cc_863 N_A_881_463#_c_1161_n N_VGND_c_2233_n 0.00434512f $X=5.215 $Y=0.797 $X2=0
+ $Y2=0
cc_864 N_A_881_463#_c_1095_n A_1107_119# 0.00537784f $X=5.785 $Y=0.797 $X2=-0.19
+ $Y2=-0.245
cc_865 N_A_881_463#_c_1070_n A_1107_119# 7.92695e-19 $X=5.87 $Y=1.165 $X2=-0.19
+ $Y2=-0.245
cc_866 N_A_975_255#_c_1213_n N_A_1524_69#_M1042_g 0.0128268f $X=10.22 $Y=1.64
+ $X2=0 $Y2=0
cc_867 N_A_975_255#_c_1229_n N_A_1524_69#_M1042_g 0.014209f $X=10.305 $Y=2.325
+ $X2=0 $Y2=0
cc_868 N_A_975_255#_c_1231_n N_A_1524_69#_M1042_g 0.0034218f $X=10.39 $Y=2.41
+ $X2=0 $Y2=0
cc_869 N_A_975_255#_c_1209_n N_A_1524_69#_c_1412_n 2.46211e-19 $X=7.69 $Y=1.74
+ $X2=0 $Y2=0
cc_870 N_A_975_255#_M1006_g N_A_1524_69#_c_1413_n 0.0189f $X=8.45 $Y=0.775 $X2=0
+ $Y2=0
cc_871 N_A_975_255#_c_1209_n N_A_1524_69#_c_1414_n 0.00927858f $X=7.69 $Y=1.74
+ $X2=0 $Y2=0
cc_872 N_A_975_255#_c_1238_n N_A_1524_69#_c_1414_n 0.0077589f $X=8.375 $Y=1.65
+ $X2=0 $Y2=0
cc_873 N_A_975_255#_M1010_g N_A_1524_69#_c_1432_n 0.00844683f $X=7.615 $Y=2.315
+ $X2=0 $Y2=0
cc_874 N_A_975_255#_c_1238_n N_A_1524_69#_c_1432_n 0.0123806f $X=8.375 $Y=1.65
+ $X2=0 $Y2=0
cc_875 N_A_975_255#_M1006_g N_A_1524_69#_c_1415_n 0.0037133f $X=8.45 $Y=0.775
+ $X2=0 $Y2=0
cc_876 N_A_975_255#_M1006_g N_A_1524_69#_c_1416_n 0.00307622f $X=8.45 $Y=0.775
+ $X2=0 $Y2=0
cc_877 N_A_975_255#_c_1217_n N_A_1524_69#_c_1416_n 0.00376461f $X=8.625 $Y=1.65
+ $X2=0 $Y2=0
cc_878 N_A_975_255#_c_1218_n N_A_1524_69#_c_1416_n 0.0107039f $X=8.79 $Y=1.65
+ $X2=0 $Y2=0
cc_879 N_A_975_255#_M1031_g N_A_1524_69#_c_1417_n 0.00295477f $X=11.045 $Y=0.765
+ $X2=0 $Y2=0
cc_880 N_A_975_255#_M1011_d N_A_1524_69#_c_1418_n 0.00719769f $X=11.815 $Y=0.345
+ $X2=0 $Y2=0
cc_881 N_A_975_255#_M1031_g N_A_1524_69#_c_1418_n 0.0180061f $X=11.045 $Y=0.765
+ $X2=0 $Y2=0
cc_882 N_A_975_255#_c_1214_n N_A_1524_69#_c_1418_n 0.004371f $X=11.175 $Y=1.675
+ $X2=0 $Y2=0
cc_883 N_A_975_255#_c_1215_n N_A_1524_69#_c_1418_n 0.0157927f $X=11.79 $Y=1.51
+ $X2=0 $Y2=0
cc_884 N_A_975_255#_c_1219_n N_A_1524_69#_c_1418_n 0.00189695f $X=11.175 $Y=1.51
+ $X2=0 $Y2=0
cc_885 N_A_975_255#_c_1220_n N_A_1524_69#_c_1418_n 0.0190634f $X=11.955 $Y=1.06
+ $X2=0 $Y2=0
cc_886 N_A_975_255#_c_1216_n N_A_1524_69#_c_1420_n 9.37757e-19 $X=11.887
+ $Y=1.345 $X2=0 $Y2=0
cc_887 N_A_975_255#_c_1220_n N_A_1524_69#_c_1420_n 0.0143801f $X=11.955 $Y=1.06
+ $X2=0 $Y2=0
cc_888 N_A_975_255#_c_1216_n N_A_1524_69#_c_1422_n 0.008716f $X=11.887 $Y=1.345
+ $X2=0 $Y2=0
cc_889 N_A_975_255#_c_1221_n N_A_1524_69#_c_1422_n 6.00847e-19 $X=11.887 $Y=1.51
+ $X2=0 $Y2=0
cc_890 N_A_975_255#_c_1213_n N_A_1524_69#_c_1423_n 0.00504594f $X=10.22 $Y=1.64
+ $X2=0 $Y2=0
cc_891 N_A_975_255#_c_1213_n N_A_1524_69#_c_1424_n 0.0391112f $X=10.22 $Y=1.64
+ $X2=0 $Y2=0
cc_892 N_A_975_255#_c_1217_n N_A_1524_69#_c_1424_n 8.27848e-19 $X=8.625 $Y=1.65
+ $X2=0 $Y2=0
cc_893 N_A_975_255#_c_1218_n N_A_1524_69#_c_1424_n 0.00485425f $X=8.79 $Y=1.65
+ $X2=0 $Y2=0
cc_894 N_A_975_255#_c_1213_n N_A_1524_69#_c_1425_n 0.04434f $X=10.22 $Y=1.64
+ $X2=0 $Y2=0
cc_895 N_A_975_255#_M1006_g N_A_1747_21#_M1039_g 0.0468539f $X=8.45 $Y=0.775
+ $X2=0 $Y2=0
cc_896 N_A_975_255#_M1006_g N_A_1747_21#_c_1598_n 0.00400663f $X=8.45 $Y=0.775
+ $X2=0 $Y2=0
cc_897 N_A_975_255#_c_1213_n N_A_1747_21#_c_1598_n 0.00989616f $X=10.22 $Y=1.64
+ $X2=0 $Y2=0
cc_898 N_A_975_255#_c_1217_n N_A_1747_21#_c_1598_n 0.0205761f $X=8.625 $Y=1.65
+ $X2=0 $Y2=0
cc_899 N_A_975_255#_c_1218_n N_A_1747_21#_c_1598_n 0.00106005f $X=8.79 $Y=1.65
+ $X2=0 $Y2=0
cc_900 N_A_975_255#_c_1213_n N_A_1747_21#_c_1599_n 0.00119711f $X=10.22 $Y=1.64
+ $X2=0 $Y2=0
cc_901 N_A_975_255#_c_1217_n N_A_1747_21#_c_1599_n 0.00291507f $X=8.625 $Y=1.65
+ $X2=0 $Y2=0
cc_902 N_A_975_255#_c_1213_n N_A_1747_21#_c_1606_n 0.0611806f $X=10.22 $Y=1.64
+ $X2=0 $Y2=0
cc_903 N_A_975_255#_c_1229_n N_A_1747_21#_c_1606_n 0.0130074f $X=10.305 $Y=2.325
+ $X2=0 $Y2=0
cc_904 N_A_975_255#_c_1229_n N_A_1747_21#_c_1607_n 0.017061f $X=10.305 $Y=2.325
+ $X2=0 $Y2=0
cc_905 N_A_975_255#_c_1231_n N_A_1747_21#_c_1607_n 0.01314f $X=10.39 $Y=2.41
+ $X2=0 $Y2=0
cc_906 N_A_975_255#_M1031_g N_A_1747_21#_c_1602_n 7.66892e-19 $X=11.045 $Y=0.765
+ $X2=0 $Y2=0
cc_907 N_A_975_255#_c_1213_n N_A_1747_21#_c_1608_n 0.0187946f $X=10.22 $Y=1.64
+ $X2=0 $Y2=0
cc_908 N_A_975_255#_c_1213_n N_A_1747_21#_c_1609_n 0.00210664f $X=10.22 $Y=1.64
+ $X2=0 $Y2=0
cc_909 N_A_975_255#_c_1217_n N_A_1747_21#_c_1609_n 0.00237283f $X=8.625 $Y=1.65
+ $X2=0 $Y2=0
cc_910 N_A_975_255#_c_1218_n N_A_1747_21#_c_1609_n 2.06729e-19 $X=8.79 $Y=1.65
+ $X2=0 $Y2=0
cc_911 N_A_975_255#_M1031_g N_A_1747_21#_c_1603_n 0.00914148f $X=11.045 $Y=0.765
+ $X2=0 $Y2=0
cc_912 N_A_975_255#_M1031_g N_CLK_M1011_g 0.0234152f $X=11.045 $Y=0.765 $X2=0
+ $Y2=0
cc_913 N_A_975_255#_c_1215_n N_CLK_M1011_g 0.0061399f $X=11.79 $Y=1.51 $X2=0
+ $Y2=0
cc_914 N_A_975_255#_c_1216_n N_CLK_M1011_g 0.00666082f $X=11.887 $Y=1.345 $X2=0
+ $Y2=0
cc_915 N_A_975_255#_c_1219_n N_CLK_M1011_g 0.0123287f $X=11.175 $Y=1.51 $X2=0
+ $Y2=0
cc_916 N_A_975_255#_c_1220_n N_CLK_M1011_g 0.00461023f $X=11.955 $Y=1.06 $X2=0
+ $Y2=0
cc_917 N_A_975_255#_c_1221_n N_CLK_M1011_g 0.00229563f $X=11.887 $Y=1.51 $X2=0
+ $Y2=0
cc_918 N_A_975_255#_M1004_g N_CLK_M1037_g 0.0161209f $X=11.045 $Y=2.465 $X2=0
+ $Y2=0
cc_919 N_A_975_255#_c_1232_n N_CLK_M1037_g 0.00357225f $X=11.175 $Y=2.325 $X2=0
+ $Y2=0
cc_920 N_A_975_255#_c_1215_n N_CLK_M1037_g 0.00748648f $X=11.79 $Y=1.51 $X2=0
+ $Y2=0
cc_921 N_A_975_255#_c_1221_n N_CLK_M1037_g 0.00154674f $X=11.887 $Y=1.51 $X2=0
+ $Y2=0
cc_922 N_A_975_255#_c_1366_p N_CLK_M1037_g 0.00340337f $X=11.955 $Y=2.835 $X2=0
+ $Y2=0
cc_923 N_A_975_255#_c_1237_n N_CLK_M1037_g 0.0272919f $X=11.932 $Y=2.67 $X2=0
+ $Y2=0
cc_924 N_A_975_255#_c_1220_n N_CLK_c_1708_n 0.00469362f $X=11.955 $Y=1.06 $X2=0
+ $Y2=0
cc_925 N_A_975_255#_c_1221_n N_CLK_c_1708_n 0.0121281f $X=11.887 $Y=1.51 $X2=0
+ $Y2=0
cc_926 N_A_975_255#_c_1215_n N_CLK_c_1709_n 0.00377579f $X=11.79 $Y=1.51 $X2=0
+ $Y2=0
cc_927 N_A_975_255#_c_1221_n N_CLK_c_1709_n 3.53117e-19 $X=11.887 $Y=1.51 $X2=0
+ $Y2=0
cc_928 N_A_975_255#_c_1221_n N_CLK_c_1710_n 2.3236e-19 $X=11.887 $Y=1.51 $X2=0
+ $Y2=0
cc_929 N_A_975_255#_c_1237_n N_CLK_c_1710_n 0.00131264f $X=11.932 $Y=2.67 $X2=0
+ $Y2=0
cc_930 N_A_975_255#_c_1221_n N_CLK_c_1711_n 0.0127443f $X=11.887 $Y=1.51 $X2=0
+ $Y2=0
cc_931 N_A_975_255#_c_1237_n N_CLK_c_1711_n 0.0679451f $X=11.932 $Y=2.67 $X2=0
+ $Y2=0
cc_932 N_A_975_255#_c_1230_n N_VPWR_M1004_d 0.00251651f $X=11.09 $Y=2.41 $X2=0
+ $Y2=0
cc_933 N_A_975_255#_c_1232_n N_VPWR_M1004_d 0.00582566f $X=11.175 $Y=2.325 $X2=0
+ $Y2=0
cc_934 N_A_975_255#_M1007_g N_VPWR_c_1879_n 0.00784611f $X=4.95 $Y=2.525 $X2=0
+ $Y2=0
cc_935 N_A_975_255#_c_1223_n N_VPWR_c_1879_n 0.0259247f $X=7.54 $Y=3.15 $X2=0
+ $Y2=0
cc_936 N_A_975_255#_c_1223_n N_VPWR_c_1880_n 0.0254156f $X=7.54 $Y=3.15 $X2=0
+ $Y2=0
cc_937 N_A_975_255#_M1010_g N_VPWR_c_1880_n 0.00478407f $X=7.615 $Y=2.315 $X2=0
+ $Y2=0
cc_938 N_A_975_255#_M1004_g N_VPWR_c_1882_n 0.0116897f $X=11.045 $Y=2.465 $X2=0
+ $Y2=0
cc_939 N_A_975_255#_c_1230_n N_VPWR_c_1882_n 0.0014994f $X=11.09 $Y=2.41 $X2=0
+ $Y2=0
cc_940 N_A_975_255#_c_1231_n N_VPWR_c_1882_n 0.0152368f $X=10.39 $Y=2.41 $X2=0
+ $Y2=0
cc_941 N_A_975_255#_M1004_g N_VPWR_c_1976_n 0.0136341f $X=11.045 $Y=2.465 $X2=0
+ $Y2=0
cc_942 N_A_975_255#_c_1230_n N_VPWR_c_1976_n 0.00923846f $X=11.09 $Y=2.41 $X2=0
+ $Y2=0
cc_943 N_A_975_255#_M1004_g N_VPWR_c_1883_n 0.013088f $X=11.045 $Y=2.465 $X2=0
+ $Y2=0
cc_944 N_A_975_255#_M1004_g N_VPWR_c_1979_n 0.00441239f $X=11.045 $Y=2.465 $X2=0
+ $Y2=0
cc_945 N_A_975_255#_c_1230_n N_VPWR_c_1979_n 0.0138843f $X=11.09 $Y=2.41 $X2=0
+ $Y2=0
cc_946 N_A_975_255#_c_1232_n N_VPWR_c_1979_n 0.0160117f $X=11.175 $Y=2.325 $X2=0
+ $Y2=0
cc_947 N_A_975_255#_c_1215_n N_VPWR_c_1979_n 0.00790796f $X=11.79 $Y=1.51 $X2=0
+ $Y2=0
cc_948 N_A_975_255#_c_1223_n N_VPWR_c_1888_n 0.0182077f $X=7.54 $Y=3.15 $X2=0
+ $Y2=0
cc_949 N_A_975_255#_c_1224_n N_VPWR_c_1892_n 0.0179753f $X=5.025 $Y=3.15 $X2=0
+ $Y2=0
cc_950 N_A_975_255#_c_1223_n N_VPWR_c_1893_n 0.0309709f $X=7.54 $Y=3.15 $X2=0
+ $Y2=0
cc_951 N_A_975_255#_M1004_g N_VPWR_c_1895_n 0.00486043f $X=11.045 $Y=2.465 $X2=0
+ $Y2=0
cc_952 N_A_975_255#_c_1366_p N_VPWR_c_1896_n 0.0104694f $X=11.955 $Y=2.835 $X2=0
+ $Y2=0
cc_953 N_A_975_255#_M1037_d N_VPWR_c_1876_n 0.00294353f $X=11.815 $Y=1.835 $X2=0
+ $Y2=0
cc_954 N_A_975_255#_c_1223_n N_VPWR_c_1876_n 0.0796734f $X=7.54 $Y=3.15 $X2=0
+ $Y2=0
cc_955 N_A_975_255#_c_1224_n N_VPWR_c_1876_n 0.0116041f $X=5.025 $Y=3.15 $X2=0
+ $Y2=0
cc_956 N_A_975_255#_M1004_g N_VPWR_c_1876_n 0.00600843f $X=11.045 $Y=2.465 $X2=0
+ $Y2=0
cc_957 N_A_975_255#_c_1230_n N_VPWR_c_1876_n 0.0236052f $X=11.09 $Y=2.41 $X2=0
+ $Y2=0
cc_958 N_A_975_255#_c_1231_n N_VPWR_c_1876_n 6.23327e-19 $X=10.39 $Y=2.41 $X2=0
+ $Y2=0
cc_959 N_A_975_255#_c_1366_p N_VPWR_c_1876_n 0.00933894f $X=11.955 $Y=2.835
+ $X2=0 $Y2=0
cc_960 N_A_975_255#_M1007_g N_A_372_50#_c_2067_n 0.0011385f $X=4.95 $Y=2.525
+ $X2=0 $Y2=0
cc_961 N_A_975_255#_M1031_g N_VGND_c_2214_n 0.00335808f $X=11.045 $Y=0.765 $X2=0
+ $Y2=0
cc_962 N_A_975_255#_M1006_g N_VGND_c_2219_n 7.27384e-19 $X=8.45 $Y=0.775 $X2=0
+ $Y2=0
cc_963 N_A_975_255#_M1031_g N_VGND_c_2223_n 0.00341315f $X=11.045 $Y=0.765 $X2=0
+ $Y2=0
cc_964 N_A_975_255#_M1030_g N_VGND_c_2233_n 9.39239e-19 $X=5.03 $Y=0.805 $X2=0
+ $Y2=0
cc_965 N_A_975_255#_M1031_g N_VGND_c_2233_n 0.00469358f $X=11.045 $Y=0.765 $X2=0
+ $Y2=0
cc_966 N_A_1524_69#_c_1413_n N_A_1747_21#_M1039_g 0.00353208f $X=8.54 $Y=0.67
+ $X2=0 $Y2=0
cc_967 N_A_1524_69#_c_1415_n N_A_1747_21#_M1039_g 0.00383104f $X=8.625 $Y=1.135
+ $X2=0 $Y2=0
cc_968 N_A_1524_69#_c_1427_n N_A_1747_21#_c_1596_n 0.0103062f $X=9.885 $Y=1.125
+ $X2=0 $Y2=0
cc_969 N_A_1524_69#_c_1424_n N_A_1747_21#_c_1598_n 0.00299173f $X=9.72 $Y=1.255
+ $X2=0 $Y2=0
cc_970 N_A_1524_69#_c_1424_n N_A_1747_21#_c_1599_n 0.0198322f $X=9.72 $Y=1.255
+ $X2=0 $Y2=0
cc_971 N_A_1524_69#_M1042_g N_A_1747_21#_c_1606_n 0.00778096f $X=9.975 $Y=2.875
+ $X2=0 $Y2=0
cc_972 N_A_1524_69#_M1042_g N_A_1747_21#_c_1632_n 0.00532878f $X=9.975 $Y=2.875
+ $X2=0 $Y2=0
cc_973 N_A_1524_69#_c_1417_n N_A_1747_21#_c_1600_n 0.0133393f $X=10.4 $Y=1.135
+ $X2=0 $Y2=0
cc_974 N_A_1524_69#_c_1419_n N_A_1747_21#_c_1600_n 0.0149364f $X=10.485 $Y=0.71
+ $X2=0 $Y2=0
cc_975 N_A_1524_69#_c_1423_n N_A_1747_21#_c_1600_n 0.00466358f $X=9.885 $Y=1.29
+ $X2=0 $Y2=0
cc_976 N_A_1524_69#_c_1425_n N_A_1747_21#_c_1600_n 0.0202205f $X=10.4 $Y=1.255
+ $X2=0 $Y2=0
cc_977 N_A_1524_69#_c_1427_n N_A_1747_21#_c_1600_n 0.0117062f $X=9.885 $Y=1.125
+ $X2=0 $Y2=0
cc_978 N_A_1524_69#_M1042_g N_A_1747_21#_c_1607_n 0.0212868f $X=9.975 $Y=2.875
+ $X2=0 $Y2=0
cc_979 N_A_1524_69#_c_1418_n N_A_1747_21#_c_1602_n 0.00611739f $X=12.3 $Y=0.71
+ $X2=0 $Y2=0
cc_980 N_A_1524_69#_c_1419_n N_A_1747_21#_c_1602_n 0.012724f $X=10.485 $Y=0.71
+ $X2=0 $Y2=0
cc_981 N_A_1524_69#_c_1418_n N_A_1747_21#_c_1603_n 0.00226205f $X=12.3 $Y=0.71
+ $X2=0 $Y2=0
cc_982 N_A_1524_69#_c_1419_n N_A_1747_21#_c_1603_n 0.00440176f $X=10.485 $Y=0.71
+ $X2=0 $Y2=0
cc_983 N_A_1524_69#_c_1425_n N_A_1747_21#_c_1603_n 0.00178258f $X=10.4 $Y=1.255
+ $X2=0 $Y2=0
cc_984 N_A_1524_69#_c_1427_n N_A_1747_21#_c_1603_n 0.00140604f $X=9.885 $Y=1.125
+ $X2=0 $Y2=0
cc_985 N_A_1524_69#_c_1418_n N_CLK_M1011_g 0.0162481f $X=12.3 $Y=0.71 $X2=0
+ $Y2=0
cc_986 N_A_1524_69#_c_1420_n N_CLK_M1011_g 0.00309178f $X=12.385 $Y=1.185 $X2=0
+ $Y2=0
cc_987 N_A_1524_69#_c_1422_n N_CLK_M1011_g 8.99584e-19 $X=12.47 $Y=1.27 $X2=0
+ $Y2=0
cc_988 N_A_1524_69#_M1044_g N_CLK_c_1708_n 0.0113192f $X=13.115 $Y=2.465 $X2=0
+ $Y2=0
cc_989 N_A_1524_69#_c_1418_n N_CLK_c_1708_n 0.00444405f $X=12.3 $Y=0.71 $X2=0
+ $Y2=0
cc_990 N_A_1524_69#_c_1421_n N_CLK_c_1708_n 0.00322163f $X=12.86 $Y=1.27 $X2=0
+ $Y2=0
cc_991 N_A_1524_69#_c_1422_n N_CLK_c_1708_n 0.00492964f $X=12.47 $Y=1.27 $X2=0
+ $Y2=0
cc_992 N_A_1524_69#_c_1426_n N_CLK_c_1708_n 0.00279431f $X=13.025 $Y=1.35 $X2=0
+ $Y2=0
cc_993 N_A_1524_69#_M1044_g N_CLK_c_1711_n 0.00134326f $X=13.115 $Y=2.465 $X2=0
+ $Y2=0
cc_994 N_A_1524_69#_c_1421_n N_CLK_c_1711_n 0.00787326f $X=12.86 $Y=1.27 $X2=0
+ $Y2=0
cc_995 N_A_1524_69#_c_1422_n N_CLK_c_1711_n 0.0151549f $X=12.47 $Y=1.27 $X2=0
+ $Y2=0
cc_996 N_A_1524_69#_c_1421_n N_A_2555_47#_M1014_g 2.94605e-19 $X=12.86 $Y=1.27
+ $X2=0 $Y2=0
cc_997 N_A_1524_69#_c_1428_n N_A_2555_47#_M1014_g 0.0232866f $X=13.025 $Y=1.185
+ $X2=0 $Y2=0
cc_998 N_A_1524_69#_M1044_g N_A_2555_47#_M1005_g 0.0232866f $X=13.115 $Y=2.465
+ $X2=0 $Y2=0
cc_999 N_A_1524_69#_c_1418_n N_A_2555_47#_c_1766_n 0.0108416f $X=12.3 $Y=0.71
+ $X2=0 $Y2=0
cc_1000 N_A_1524_69#_c_1420_n N_A_2555_47#_c_1766_n 0.00222847f $X=12.385
+ $Y=1.185 $X2=0 $Y2=0
cc_1001 N_A_1524_69#_c_1421_n N_A_2555_47#_c_1785_n 0.00843997f $X=12.86 $Y=1.27
+ $X2=0 $Y2=0
cc_1002 N_A_1524_69#_c_1428_n N_A_2555_47#_c_1785_n 0.011682f $X=13.025 $Y=1.185
+ $X2=0 $Y2=0
cc_1003 N_A_1524_69#_c_1420_n N_A_2555_47#_c_1767_n 0.0111469f $X=12.385
+ $Y=1.185 $X2=0 $Y2=0
cc_1004 N_A_1524_69#_c_1421_n N_A_2555_47#_c_1767_n 0.0209874f $X=12.86 $Y=1.27
+ $X2=0 $Y2=0
cc_1005 N_A_1524_69#_c_1426_n N_A_2555_47#_c_1767_n 0.00102421f $X=13.025
+ $Y=1.35 $X2=0 $Y2=0
cc_1006 N_A_1524_69#_M1044_g N_A_2555_47#_c_1777_n 0.0152979f $X=13.115 $Y=2.465
+ $X2=0 $Y2=0
cc_1007 N_A_1524_69#_c_1421_n N_A_2555_47#_c_1777_n 0.00770832f $X=12.86 $Y=1.27
+ $X2=0 $Y2=0
cc_1008 N_A_1524_69#_c_1426_n N_A_2555_47#_c_1777_n 2.92379e-19 $X=13.025
+ $Y=1.35 $X2=0 $Y2=0
cc_1009 N_A_1524_69#_c_1421_n N_A_2555_47#_c_1778_n 0.0143644f $X=12.86 $Y=1.27
+ $X2=0 $Y2=0
cc_1010 N_A_1524_69#_c_1426_n N_A_2555_47#_c_1778_n 0.00101687f $X=13.025
+ $Y=1.35 $X2=0 $Y2=0
cc_1011 N_A_1524_69#_c_1421_n N_A_2555_47#_c_1768_n 0.0155271f $X=12.86 $Y=1.27
+ $X2=0 $Y2=0
cc_1012 N_A_1524_69#_c_1428_n N_A_2555_47#_c_1768_n 0.00518864f $X=13.025
+ $Y=1.185 $X2=0 $Y2=0
cc_1013 N_A_1524_69#_M1044_g N_A_2555_47#_c_1769_n 0.00416796f $X=13.115
+ $Y=2.465 $X2=0 $Y2=0
cc_1014 N_A_1524_69#_c_1421_n N_A_2555_47#_c_1770_n 0.00999458f $X=12.86 $Y=1.27
+ $X2=0 $Y2=0
cc_1015 N_A_1524_69#_c_1426_n N_A_2555_47#_c_1770_n 0.00241163f $X=13.025
+ $Y=1.35 $X2=0 $Y2=0
cc_1016 N_A_1524_69#_c_1426_n N_A_2555_47#_c_1771_n 0.0232866f $X=13.025 $Y=1.35
+ $X2=0 $Y2=0
cc_1017 N_A_1524_69#_M1042_g N_VPWR_c_1882_n 0.0124046f $X=9.975 $Y=2.875 $X2=0
+ $Y2=0
cc_1018 N_A_1524_69#_M1044_g N_VPWR_c_1884_n 0.0162124f $X=13.115 $Y=2.465 $X2=0
+ $Y2=0
cc_1019 N_A_1524_69#_M1042_g N_VPWR_c_1894_n 0.00371605f $X=9.975 $Y=2.875 $X2=0
+ $Y2=0
cc_1020 N_A_1524_69#_M1044_g N_VPWR_c_1896_n 0.00486043f $X=13.115 $Y=2.465
+ $X2=0 $Y2=0
cc_1021 N_A_1524_69#_M1010_d N_VPWR_c_1876_n 0.00327078f $X=7.69 $Y=1.895 $X2=0
+ $Y2=0
cc_1022 N_A_1524_69#_M1042_g N_VPWR_c_1876_n 0.00700579f $X=9.975 $Y=2.875 $X2=0
+ $Y2=0
cc_1023 N_A_1524_69#_M1044_g N_VPWR_c_1876_n 0.00954696f $X=13.115 $Y=2.465
+ $X2=0 $Y2=0
cc_1024 N_A_1524_69#_c_1418_n N_VGND_M1031_d 0.0145629f $X=12.3 $Y=0.71 $X2=0
+ $Y2=0
cc_1025 N_A_1524_69#_c_1413_n N_VGND_c_2213_n 0.0232571f $X=8.54 $Y=0.67 $X2=0
+ $Y2=0
cc_1026 N_A_1524_69#_c_1424_n N_VGND_c_2213_n 0.0241534f $X=9.72 $Y=1.255 $X2=0
+ $Y2=0
cc_1027 N_A_1524_69#_c_1418_n N_VGND_c_2214_n 0.0248493f $X=12.3 $Y=0.71 $X2=0
+ $Y2=0
cc_1028 N_A_1524_69#_c_1428_n N_VGND_c_2215_n 0.011338f $X=13.025 $Y=1.185 $X2=0
+ $Y2=0
cc_1029 N_A_1524_69#_c_1413_n N_VGND_c_2219_n 0.038593f $X=8.54 $Y=0.67 $X2=0
+ $Y2=0
cc_1030 N_A_1524_69#_c_1447_n N_VGND_c_2219_n 0.00539113f $X=7.655 $Y=0.67 $X2=0
+ $Y2=0
cc_1031 N_A_1524_69#_c_1418_n N_VGND_c_2223_n 0.00974322f $X=12.3 $Y=0.71 $X2=0
+ $Y2=0
cc_1032 N_A_1524_69#_c_1418_n N_VGND_c_2224_n 0.016786f $X=12.3 $Y=0.71 $X2=0
+ $Y2=0
cc_1033 N_A_1524_69#_c_1428_n N_VGND_c_2224_n 0.00486043f $X=13.025 $Y=1.185
+ $X2=0 $Y2=0
cc_1034 N_A_1524_69#_c_1413_n N_VGND_c_2233_n 0.0376065f $X=8.54 $Y=0.67 $X2=0
+ $Y2=0
cc_1035 N_A_1524_69#_c_1447_n N_VGND_c_2233_n 0.00542958f $X=7.655 $Y=0.67 $X2=0
+ $Y2=0
cc_1036 N_A_1524_69#_c_1418_n N_VGND_c_2233_n 0.0456177f $X=12.3 $Y=0.71 $X2=0
+ $Y2=0
cc_1037 N_A_1524_69#_c_1427_n N_VGND_c_2233_n 7.85159e-19 $X=9.885 $Y=1.125
+ $X2=0 $Y2=0
cc_1038 N_A_1524_69#_c_1428_n N_VGND_c_2233_n 0.00583049f $X=13.025 $Y=1.185
+ $X2=0 $Y2=0
cc_1039 N_A_1747_21#_M1028_g N_VPWR_c_1881_n 0.00945383f $X=8.825 $Y=2.875 $X2=0
+ $Y2=0
cc_1040 N_A_1747_21#_c_1632_n N_VPWR_c_1881_n 0.012531f $X=9.87 $Y=2.935 $X2=0
+ $Y2=0
cc_1041 N_A_1747_21#_c_1632_n N_VPWR_c_1882_n 0.0169159f $X=9.87 $Y=2.935 $X2=0
+ $Y2=0
cc_1042 N_A_1747_21#_c_1607_n N_VPWR_c_1882_n 0.0113423f $X=9.955 $Y=2.825 $X2=0
+ $Y2=0
cc_1043 N_A_1747_21#_M1028_g N_VPWR_c_1888_n 0.00422429f $X=8.825 $Y=2.875 $X2=0
+ $Y2=0
cc_1044 N_A_1747_21#_c_1632_n N_VPWR_c_1894_n 0.0216426f $X=9.87 $Y=2.935 $X2=0
+ $Y2=0
cc_1045 N_A_1747_21#_M1018_d N_VPWR_c_1876_n 0.00224111f $X=9.62 $Y=2.665 $X2=0
+ $Y2=0
cc_1046 N_A_1747_21#_M1028_g N_VPWR_c_1876_n 0.00694756f $X=8.825 $Y=2.875 $X2=0
+ $Y2=0
cc_1047 N_A_1747_21#_c_1632_n N_VPWR_c_1876_n 0.0158055f $X=9.87 $Y=2.935 $X2=0
+ $Y2=0
cc_1048 N_A_1747_21#_M1039_g N_VGND_c_2213_n 0.00905916f $X=8.81 $Y=0.775 $X2=0
+ $Y2=0
cc_1049 N_A_1747_21#_c_1596_n N_VGND_c_2213_n 0.0251144f $X=10.245 $Y=0.18 $X2=0
+ $Y2=0
cc_1050 N_A_1747_21#_c_1599_n N_VGND_c_2213_n 0.00520779f $X=9.075 $Y=1.17 $X2=0
+ $Y2=0
cc_1051 N_A_1747_21#_c_1600_n N_VGND_c_2213_n 0.0156774f $X=10.01 $Y=0.8 $X2=0
+ $Y2=0
cc_1052 N_A_1747_21#_c_1601_n N_VGND_c_2213_n 0.00771614f $X=10.145 $Y=0.355
+ $X2=0 $Y2=0
cc_1053 N_A_1747_21#_c_1602_n N_VGND_c_2214_n 0.0044287f $X=10.41 $Y=0.35 $X2=0
+ $Y2=0
cc_1054 N_A_1747_21#_c_1603_n N_VGND_c_2214_n 0.00168329f $X=10.41 $Y=0.18 $X2=0
+ $Y2=0
cc_1055 N_A_1747_21#_c_1597_n N_VGND_c_2219_n 0.00854661f $X=8.885 $Y=0.18 $X2=0
+ $Y2=0
cc_1056 N_A_1747_21#_c_1596_n N_VGND_c_2223_n 0.0355164f $X=10.245 $Y=0.18 $X2=0
+ $Y2=0
cc_1057 N_A_1747_21#_c_1601_n N_VGND_c_2223_n 0.0205159f $X=10.145 $Y=0.355
+ $X2=0 $Y2=0
cc_1058 N_A_1747_21#_c_1602_n N_VGND_c_2223_n 0.0270013f $X=10.41 $Y=0.35 $X2=0
+ $Y2=0
cc_1059 N_A_1747_21#_c_1596_n N_VGND_c_2233_n 0.0378679f $X=10.245 $Y=0.18 $X2=0
+ $Y2=0
cc_1060 N_A_1747_21#_c_1597_n N_VGND_c_2233_n 0.0115248f $X=8.885 $Y=0.18 $X2=0
+ $Y2=0
cc_1061 N_A_1747_21#_c_1601_n N_VGND_c_2233_n 0.0103038f $X=10.145 $Y=0.355
+ $X2=0 $Y2=0
cc_1062 N_A_1747_21#_c_1602_n N_VGND_c_2233_n 0.0142879f $X=10.41 $Y=0.35 $X2=0
+ $Y2=0
cc_1063 N_A_1747_21#_c_1603_n N_VGND_c_2233_n 0.00986114f $X=10.41 $Y=0.18 $X2=0
+ $Y2=0
cc_1064 N_CLK_c_1710_n N_A_2555_47#_c_1776_n 0.00177271f $X=12.405 $Y=1.625
+ $X2=0 $Y2=0
cc_1065 N_CLK_c_1711_n N_A_2555_47#_c_1776_n 0.0489729f $X=12.405 $Y=1.625 $X2=0
+ $Y2=0
cc_1066 N_CLK_c_1710_n N_A_2555_47#_c_1778_n 0.00158259f $X=12.405 $Y=1.625
+ $X2=0 $Y2=0
cc_1067 N_CLK_c_1711_n N_A_2555_47#_c_1778_n 0.0145654f $X=12.405 $Y=1.625 $X2=0
+ $Y2=0
cc_1068 N_CLK_M1037_g N_VPWR_c_1883_n 0.00551575f $X=11.74 $Y=2.465 $X2=0 $Y2=0
cc_1069 N_CLK_M1037_g N_VPWR_c_1896_n 0.00572634f $X=11.74 $Y=2.465 $X2=0 $Y2=0
cc_1070 N_CLK_M1037_g N_VPWR_c_1876_n 0.0125062f $X=11.74 $Y=2.465 $X2=0 $Y2=0
cc_1071 N_CLK_c_1711_n N_VPWR_c_1876_n 0.0167943f $X=12.405 $Y=1.625 $X2=0 $Y2=0
cc_1072 N_CLK_M1011_g N_VGND_c_2214_n 0.00614479f $X=11.74 $Y=0.765 $X2=0 $Y2=0
cc_1073 N_CLK_M1011_g N_VGND_c_2224_n 0.00341315f $X=11.74 $Y=0.765 $X2=0 $Y2=0
cc_1074 N_CLK_M1011_g N_VGND_c_2233_n 0.00498864f $X=11.74 $Y=0.765 $X2=0 $Y2=0
cc_1075 N_A_2555_47#_c_1777_n N_VPWR_M1044_d 0.00180108f $X=13.305 $Y=1.84 $X2=0
+ $Y2=0
cc_1076 N_A_2555_47#_M1005_g N_VPWR_c_1884_n 0.0144719f $X=13.545 $Y=2.465 $X2=0
+ $Y2=0
cc_1077 N_A_2555_47#_M1008_g N_VPWR_c_1884_n 7.35335e-19 $X=13.975 $Y=2.465
+ $X2=0 $Y2=0
cc_1078 N_A_2555_47#_c_1777_n N_VPWR_c_1884_n 0.0165445f $X=13.305 $Y=1.84 $X2=0
+ $Y2=0
cc_1079 N_A_2555_47#_c_1809_p N_VPWR_c_1884_n 5.55389e-19 $X=14.655 $Y=1.48
+ $X2=0 $Y2=0
cc_1080 N_A_2555_47#_M1005_g N_VPWR_c_1885_n 6.82734e-19 $X=13.545 $Y=2.465
+ $X2=0 $Y2=0
cc_1081 N_A_2555_47#_M1008_g N_VPWR_c_1885_n 0.0115861f $X=13.975 $Y=2.465 $X2=0
+ $Y2=0
cc_1082 N_A_2555_47#_M1025_g N_VPWR_c_1885_n 0.0115861f $X=14.445 $Y=2.465 $X2=0
+ $Y2=0
cc_1083 N_A_2555_47#_M1034_g N_VPWR_c_1885_n 6.82734e-19 $X=14.875 $Y=2.465
+ $X2=0 $Y2=0
cc_1084 N_A_2555_47#_M1025_g N_VPWR_c_1887_n 7.3263e-19 $X=14.445 $Y=2.465 $X2=0
+ $Y2=0
cc_1085 N_A_2555_47#_M1034_g N_VPWR_c_1887_n 0.0149339f $X=14.875 $Y=2.465 $X2=0
+ $Y2=0
cc_1086 N_A_2555_47#_c_1776_n N_VPWR_c_1896_n 0.0174527f $X=12.9 $Y=1.98 $X2=0
+ $Y2=0
cc_1087 N_A_2555_47#_M1005_g N_VPWR_c_1897_n 0.00486043f $X=13.545 $Y=2.465
+ $X2=0 $Y2=0
cc_1088 N_A_2555_47#_M1008_g N_VPWR_c_1897_n 0.00564095f $X=13.975 $Y=2.465
+ $X2=0 $Y2=0
cc_1089 N_A_2555_47#_M1025_g N_VPWR_c_1898_n 0.00564095f $X=14.445 $Y=2.465
+ $X2=0 $Y2=0
cc_1090 N_A_2555_47#_M1034_g N_VPWR_c_1898_n 0.00486043f $X=14.875 $Y=2.465
+ $X2=0 $Y2=0
cc_1091 N_A_2555_47#_M1044_s N_VPWR_c_1876_n 0.00371702f $X=12.775 $Y=1.835
+ $X2=0 $Y2=0
cc_1092 N_A_2555_47#_M1005_g N_VPWR_c_1876_n 0.00824727f $X=13.545 $Y=2.465
+ $X2=0 $Y2=0
cc_1093 N_A_2555_47#_M1008_g N_VPWR_c_1876_n 0.00948291f $X=13.975 $Y=2.465
+ $X2=0 $Y2=0
cc_1094 N_A_2555_47#_M1025_g N_VPWR_c_1876_n 0.00948291f $X=14.445 $Y=2.465
+ $X2=0 $Y2=0
cc_1095 N_A_2555_47#_M1034_g N_VPWR_c_1876_n 0.00824727f $X=14.875 $Y=2.465
+ $X2=0 $Y2=0
cc_1096 N_A_2555_47#_c_1776_n N_VPWR_c_1876_n 0.00983606f $X=12.9 $Y=1.98 $X2=0
+ $Y2=0
cc_1097 N_A_2555_47#_M1005_g N_Q_c_2157_n 8.61148e-19 $X=13.545 $Y=2.465 $X2=0
+ $Y2=0
cc_1098 N_A_2555_47#_c_1777_n N_Q_c_2157_n 0.00999132f $X=13.305 $Y=1.84 $X2=0
+ $Y2=0
cc_1099 N_A_2555_47#_c_1769_n N_Q_c_2157_n 0.00145317f $X=13.39 $Y=1.755 $X2=0
+ $Y2=0
cc_1100 N_A_2555_47#_c_1809_p N_Q_c_2157_n 0.0169449f $X=14.655 $Y=1.48 $X2=0
+ $Y2=0
cc_1101 N_A_2555_47#_c_1771_n N_Q_c_2157_n 0.00256759f $X=14.875 $Y=1.48 $X2=0
+ $Y2=0
cc_1102 N_A_2555_47#_M1027_g N_Q_c_2152_n 0.0139613f $X=13.975 $Y=0.655 $X2=0
+ $Y2=0
cc_1103 N_A_2555_47#_M1040_g N_Q_c_2152_n 0.0145139f $X=14.405 $Y=0.655 $X2=0
+ $Y2=0
cc_1104 N_A_2555_47#_c_1809_p N_Q_c_2152_n 0.0469373f $X=14.655 $Y=1.48 $X2=0
+ $Y2=0
cc_1105 N_A_2555_47#_c_1771_n N_Q_c_2152_n 0.00246815f $X=14.875 $Y=1.48 $X2=0
+ $Y2=0
cc_1106 N_A_2555_47#_M1014_g N_Q_c_2153_n 0.00129639f $X=13.545 $Y=0.655 $X2=0
+ $Y2=0
cc_1107 N_A_2555_47#_c_1768_n N_Q_c_2153_n 0.0120231f $X=13.39 $Y=1.395 $X2=0
+ $Y2=0
cc_1108 N_A_2555_47#_c_1809_p N_Q_c_2153_n 0.0153308f $X=14.655 $Y=1.48 $X2=0
+ $Y2=0
cc_1109 N_A_2555_47#_c_1771_n N_Q_c_2153_n 0.00256759f $X=14.875 $Y=1.48 $X2=0
+ $Y2=0
cc_1110 N_A_2555_47#_M1008_g N_Q_c_2158_n 0.0164983f $X=13.975 $Y=2.465 $X2=0
+ $Y2=0
cc_1111 N_A_2555_47#_M1025_g N_Q_c_2158_n 0.0166791f $X=14.445 $Y=2.465 $X2=0
+ $Y2=0
cc_1112 N_A_2555_47#_c_1809_p N_Q_c_2158_n 0.0481817f $X=14.655 $Y=1.48 $X2=0
+ $Y2=0
cc_1113 N_A_2555_47#_c_1771_n N_Q_c_2158_n 0.00365612f $X=14.875 $Y=1.48 $X2=0
+ $Y2=0
cc_1114 N_A_2555_47#_M1034_g N_Q_c_2159_n 0.019233f $X=14.875 $Y=2.465 $X2=0
+ $Y2=0
cc_1115 N_A_2555_47#_c_1809_p N_Q_c_2159_n 0.00541669f $X=14.655 $Y=1.48 $X2=0
+ $Y2=0
cc_1116 N_A_2555_47#_M1043_g N_Q_c_2154_n 0.0177674f $X=14.875 $Y=0.655 $X2=0
+ $Y2=0
cc_1117 N_A_2555_47#_c_1809_p N_Q_c_2154_n 0.00203336f $X=14.655 $Y=1.48 $X2=0
+ $Y2=0
cc_1118 N_A_2555_47#_M1043_g N_Q_c_2155_n 0.0204755f $X=14.875 $Y=0.655 $X2=0
+ $Y2=0
cc_1119 N_A_2555_47#_c_1809_p N_Q_c_2155_n 0.0132586f $X=14.655 $Y=1.48 $X2=0
+ $Y2=0
cc_1120 N_A_2555_47#_c_1809_p N_Q_c_2156_n 0.0213824f $X=14.655 $Y=1.48 $X2=0
+ $Y2=0
cc_1121 N_A_2555_47#_c_1771_n N_Q_c_2156_n 0.00376674f $X=14.875 $Y=1.48 $X2=0
+ $Y2=0
cc_1122 N_A_2555_47#_c_1809_p N_Q_c_2161_n 0.0161378f $X=14.655 $Y=1.48 $X2=0
+ $Y2=0
cc_1123 N_A_2555_47#_c_1771_n N_Q_c_2161_n 0.00256759f $X=14.875 $Y=1.48 $X2=0
+ $Y2=0
cc_1124 N_A_2555_47#_c_1785_n N_VGND_M1041_d 0.00396699f $X=13.305 $Y=0.925
+ $X2=0 $Y2=0
cc_1125 N_A_2555_47#_c_1768_n N_VGND_M1041_d 6.6282e-19 $X=13.39 $Y=1.395 $X2=0
+ $Y2=0
cc_1126 N_A_2555_47#_M1014_g N_VGND_c_2215_n 0.010323f $X=13.545 $Y=0.655 $X2=0
+ $Y2=0
cc_1127 N_A_2555_47#_M1027_g N_VGND_c_2215_n 5.65914e-19 $X=13.975 $Y=0.655
+ $X2=0 $Y2=0
cc_1128 N_A_2555_47#_c_1785_n N_VGND_c_2215_n 0.0162168f $X=13.305 $Y=0.925
+ $X2=0 $Y2=0
cc_1129 N_A_2555_47#_M1014_g N_VGND_c_2216_n 6.25324e-19 $X=13.545 $Y=0.655
+ $X2=0 $Y2=0
cc_1130 N_A_2555_47#_M1027_g N_VGND_c_2216_n 0.0109423f $X=13.975 $Y=0.655 $X2=0
+ $Y2=0
cc_1131 N_A_2555_47#_M1040_g N_VGND_c_2216_n 0.0111552f $X=14.405 $Y=0.655 $X2=0
+ $Y2=0
cc_1132 N_A_2555_47#_M1043_g N_VGND_c_2216_n 6.15114e-19 $X=14.875 $Y=0.655
+ $X2=0 $Y2=0
cc_1133 N_A_2555_47#_M1043_g N_VGND_c_2218_n 0.00344465f $X=14.875 $Y=0.655
+ $X2=0 $Y2=0
cc_1134 N_A_2555_47#_c_1766_n N_VGND_c_2224_n 0.0178111f $X=12.9 $Y=0.42 $X2=0
+ $Y2=0
cc_1135 N_A_2555_47#_M1014_g N_VGND_c_2225_n 0.00486043f $X=13.545 $Y=0.655
+ $X2=0 $Y2=0
cc_1136 N_A_2555_47#_M1027_g N_VGND_c_2225_n 0.00486043f $X=13.975 $Y=0.655
+ $X2=0 $Y2=0
cc_1137 N_A_2555_47#_M1040_g N_VGND_c_2226_n 0.00486043f $X=14.405 $Y=0.655
+ $X2=0 $Y2=0
cc_1138 N_A_2555_47#_M1043_g N_VGND_c_2226_n 0.00585385f $X=14.875 $Y=0.655
+ $X2=0 $Y2=0
cc_1139 N_A_2555_47#_M1041_s N_VGND_c_2233_n 0.0024321f $X=12.775 $Y=0.235 $X2=0
+ $Y2=0
cc_1140 N_A_2555_47#_M1014_g N_VGND_c_2233_n 0.00824727f $X=13.545 $Y=0.655
+ $X2=0 $Y2=0
cc_1141 N_A_2555_47#_M1027_g N_VGND_c_2233_n 0.00824727f $X=13.975 $Y=0.655
+ $X2=0 $Y2=0
cc_1142 N_A_2555_47#_M1040_g N_VGND_c_2233_n 0.00834786f $X=14.405 $Y=0.655
+ $X2=0 $Y2=0
cc_1143 N_A_2555_47#_M1043_g N_VGND_c_2233_n 0.0115649f $X=14.875 $Y=0.655 $X2=0
+ $Y2=0
cc_1144 N_A_2555_47#_c_1766_n N_VGND_c_2233_n 0.0100304f $X=12.9 $Y=0.42 $X2=0
+ $Y2=0
cc_1145 N_A_2555_47#_c_1785_n N_VGND_c_2233_n 0.00604388f $X=13.305 $Y=0.925
+ $X2=0 $Y2=0
cc_1146 N_VPWR_M1012_d N_A_372_50#_c_2064_n 0.00399362f $X=3.295 $Y=2.315 $X2=0
+ $Y2=0
cc_1147 N_VPWR_c_1878_n N_A_372_50#_c_2064_n 0.0253521f $X=3.52 $Y=2.77 $X2=0
+ $Y2=0
cc_1148 N_VPWR_c_1876_n N_A_372_50#_c_2064_n 0.024461f $X=15.12 $Y=3.33 $X2=0
+ $Y2=0
cc_1149 N_VPWR_c_1877_n N_A_372_50#_c_2066_n 0.0228765f $X=1.745 $Y=2.46 $X2=0
+ $Y2=0
cc_1150 N_VPWR_c_1878_n N_A_372_50#_c_2066_n 0.00879107f $X=3.52 $Y=2.77 $X2=0
+ $Y2=0
cc_1151 N_VPWR_c_1891_n N_A_372_50#_c_2066_n 0.0142054f $X=3.355 $Y=3.33 $X2=0
+ $Y2=0
cc_1152 N_VPWR_c_1876_n N_A_372_50#_c_2066_n 0.0118456f $X=15.12 $Y=3.33 $X2=0
+ $Y2=0
cc_1153 N_VPWR_c_1892_n N_A_372_50#_c_2067_n 0.0116964f $X=5.36 $Y=3.33 $X2=0
+ $Y2=0
cc_1154 N_VPWR_c_1876_n N_A_372_50#_c_2067_n 0.0155229f $X=15.12 $Y=3.33 $X2=0
+ $Y2=0
cc_1155 N_VPWR_c_1876_n A_1662_533# 0.00520703f $X=15.12 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_1156 N_VPWR_c_1876_n N_Q_M1005_d 0.00467071f $X=15.12 $Y=3.33 $X2=0 $Y2=0
cc_1157 N_VPWR_c_1876_n N_Q_M1025_d 0.00501859f $X=15.12 $Y=3.33 $X2=0 $Y2=0
cc_1158 N_VPWR_c_1897_n N_Q_c_2191_n 0.0131621f $X=14.045 $Y=3.33 $X2=0 $Y2=0
cc_1159 N_VPWR_c_1876_n N_Q_c_2191_n 0.00808656f $X=15.12 $Y=3.33 $X2=0 $Y2=0
cc_1160 N_VPWR_M1008_s N_Q_c_2158_n 0.002216f $X=14.05 $Y=1.835 $X2=0 $Y2=0
cc_1161 N_VPWR_c_1885_n N_Q_c_2158_n 0.0177485f $X=14.21 $Y=2.24 $X2=0 $Y2=0
cc_1162 N_VPWR_c_1898_n N_Q_c_2195_n 0.0128073f $X=14.925 $Y=3.33 $X2=0 $Y2=0
cc_1163 N_VPWR_c_1876_n N_Q_c_2195_n 0.0076925f $X=15.12 $Y=3.33 $X2=0 $Y2=0
cc_1164 N_VPWR_M1034_s N_Q_c_2159_n 0.00300749f $X=14.95 $Y=1.835 $X2=0 $Y2=0
cc_1165 N_VPWR_c_1887_n N_Q_c_2159_n 0.0242438f $X=15.09 $Y=2.24 $X2=0 $Y2=0
cc_1166 N_A_372_50#_c_2064_n A_565_463# 0.00422339f $X=3.78 $Y=2.385 $X2=-0.19
+ $Y2=-0.245
cc_1167 N_A_372_50#_c_2057_n N_VGND_c_2210_n 0.0209093f $X=3.78 $Y=0.98 $X2=0
+ $Y2=0
cc_1168 N_A_372_50#_c_2063_n N_VGND_c_2210_n 0.00700638f $X=3.78 $Y=0.895 $X2=0
+ $Y2=0
cc_1169 N_A_372_50#_c_2059_n N_VGND_c_2211_n 0.0119009f $X=4.78 $Y=0.805 $X2=0
+ $Y2=0
cc_1170 N_A_372_50#_c_2063_n N_VGND_c_2211_n 0.0087902f $X=3.78 $Y=0.895 $X2=0
+ $Y2=0
cc_1171 N_A_372_50#_c_2059_n N_VGND_c_2233_n 0.0161927f $X=4.78 $Y=0.805 $X2=0
+ $Y2=0
cc_1172 N_A_372_50#_c_2061_n N_VGND_c_2233_n 0.00197315f $X=2.905 $Y=0.94 $X2=0
+ $Y2=0
cc_1173 N_A_372_50#_c_2063_n N_VGND_c_2233_n 0.0117026f $X=3.78 $Y=0.895 $X2=0
+ $Y2=0
cc_1174 N_A_372_50#_c_2062_n N_noxref_24_M1032_d 0.00157942f $X=3.075 $Y=0.94
+ $X2=0 $Y2=0
cc_1175 N_A_372_50#_M1023_d N_noxref_24_c_2367_n 0.00992221f $X=1.86 $Y=0.25
+ $X2=0 $Y2=0
cc_1176 N_A_372_50#_c_2060_n N_noxref_24_c_2367_n 0.0239361f $X=2.115 $Y=0.7
+ $X2=0 $Y2=0
cc_1177 N_A_372_50#_c_2061_n N_noxref_24_c_2367_n 0.0125954f $X=2.905 $Y=0.94
+ $X2=0 $Y2=0
cc_1178 N_A_372_50#_c_2060_n N_noxref_24_c_2368_n 8.93443e-19 $X=2.115 $Y=0.7
+ $X2=0 $Y2=0
cc_1179 N_A_372_50#_c_2057_n N_noxref_24_c_2369_n 0.00454663f $X=3.78 $Y=0.98
+ $X2=0 $Y2=0
cc_1180 N_A_372_50#_c_2060_n N_noxref_24_c_2369_n 0.00148907f $X=2.115 $Y=0.7
+ $X2=0 $Y2=0
cc_1181 N_A_372_50#_c_2061_n N_noxref_24_c_2369_n 0.0124136f $X=2.905 $Y=0.94
+ $X2=0 $Y2=0
cc_1182 N_A_372_50#_c_2061_n noxref_26 0.00147531f $X=2.905 $Y=0.94 $X2=-0.19
+ $Y2=-0.245
cc_1183 N_Q_c_2152_n N_VGND_M1027_d 0.00176773f $X=14.525 $Y=1.135 $X2=0 $Y2=0
cc_1184 N_Q_c_2154_n N_VGND_M1043_d 0.00239587f $X=15 $Y=1.14 $X2=0 $Y2=0
cc_1185 N_Q_c_2152_n N_VGND_c_2216_n 0.0171443f $X=14.525 $Y=1.135 $X2=0 $Y2=0
cc_1186 N_Q_c_2154_n N_VGND_c_2218_n 0.0224079f $X=15 $Y=1.14 $X2=0 $Y2=0
cc_1187 N_Q_c_2203_p N_VGND_c_2225_n 0.0124525f $X=13.76 $Y=0.42 $X2=0 $Y2=0
cc_1188 N_Q_c_2204_p N_VGND_c_2226_n 0.0165068f $X=14.62 $Y=0.42 $X2=0 $Y2=0
cc_1189 N_Q_M1014_s N_VGND_c_2233_n 0.00536646f $X=13.62 $Y=0.235 $X2=0 $Y2=0
cc_1190 N_Q_M1040_s N_VGND_c_2233_n 0.00447057f $X=14.48 $Y=0.235 $X2=0 $Y2=0
cc_1191 N_Q_c_2203_p N_VGND_c_2233_n 0.00730901f $X=13.76 $Y=0.42 $X2=0 $Y2=0
cc_1192 N_Q_c_2204_p N_VGND_c_2233_n 0.0102248f $X=14.62 $Y=0.42 $X2=0 $Y2=0
cc_1193 N_VGND_c_2222_n N_noxref_24_c_2367_n 0.0891012f $X=3.355 $Y=0 $X2=0
+ $Y2=0
cc_1194 N_VGND_c_2233_n N_noxref_24_c_2367_n 0.0543934f $X=15.12 $Y=0 $X2=0
+ $Y2=0
cc_1195 N_VGND_c_2209_n N_noxref_24_c_2368_n 0.0284909f $X=0.69 $Y=0.525 $X2=0
+ $Y2=0
cc_1196 N_VGND_c_2222_n N_noxref_24_c_2368_n 0.0202612f $X=3.355 $Y=0 $X2=0
+ $Y2=0
cc_1197 N_VGND_c_2233_n N_noxref_24_c_2368_n 0.0124489f $X=15.12 $Y=0 $X2=0
+ $Y2=0
cc_1198 N_VGND_c_2210_n N_noxref_24_c_2369_n 0.0205756f $X=3.45 $Y=0.56 $X2=0
+ $Y2=0
cc_1199 N_VGND_c_2222_n N_noxref_24_c_2369_n 0.0224826f $X=3.355 $Y=0 $X2=0
+ $Y2=0
cc_1200 N_VGND_c_2233_n N_noxref_24_c_2369_n 0.0124647f $X=15.12 $Y=0 $X2=0
+ $Y2=0
cc_1201 N_noxref_24_c_2367_n noxref_25 0.00456442f $X=2.855 $Y=0.34 $X2=-0.19
+ $Y2=-0.245
cc_1202 N_noxref_24_c_2367_n noxref_26 0.00151984f $X=2.855 $Y=0.34 $X2=-0.19
+ $Y2=-0.245
