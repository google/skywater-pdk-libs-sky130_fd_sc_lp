* File: sky130_fd_sc_lp__or2_0.pex.spice
* Created: Fri Aug 28 11:21:02 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__OR2_0%B 5 9 11 12 13 14 15 16 22
r34 22 24 46.1517 $w=4.2e-07 $l=1.65e-07 $layer=POLY_cond $X=0.545 $Y=1.005
+ $X2=0.545 $Y2=0.84
r35 22 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.5
+ $Y=1.005 $X2=0.5 $Y2=1.005
r36 15 16 8.85098 $w=4.98e-07 $l=3.7e-07 $layer=LI1_cond $X=0.335 $Y=1.665
+ $X2=0.335 $Y2=2.035
r37 14 15 8.85098 $w=4.98e-07 $l=3.7e-07 $layer=LI1_cond $X=0.335 $Y=1.295
+ $X2=0.335 $Y2=1.665
r38 14 23 6.93725 $w=4.98e-07 $l=2.9e-07 $layer=LI1_cond $X=0.335 $Y=1.295
+ $X2=0.335 $Y2=1.005
r39 13 23 1.91373 $w=4.98e-07 $l=8e-08 $layer=LI1_cond $X=0.335 $Y=0.925
+ $X2=0.335 $Y2=1.005
r40 11 12 44.1654 $w=4.2e-07 $l=1.5e-07 $layer=POLY_cond $X=0.565 $Y=1.36
+ $X2=0.565 $Y2=1.51
r41 9 12 546.096 $w=1.5e-07 $l=1.065e-06 $layer=POLY_cond $X=0.72 $Y=2.575
+ $X2=0.72 $Y2=1.51
r42 5 24 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.68 $Y=0.445
+ $X2=0.68 $Y2=0.84
r43 1 22 5.95879 $w=4.2e-07 $l=4.5e-08 $layer=POLY_cond $X=0.545 $Y=1.05
+ $X2=0.545 $Y2=1.005
r44 1 11 41.0494 $w=4.2e-07 $l=3.1e-07 $layer=POLY_cond $X=0.545 $Y=1.05
+ $X2=0.545 $Y2=1.36
.ends

.subckt PM_SKY130_FD_SC_LP__OR2_0%A 3 7 11 12 13 14 15 20
c41 11 0 1.4009e-19 $X=1.2 $Y=1.66
r42 14 15 16.4002 $w=2.58e-07 $l=3.7e-07 $layer=LI1_cond $X=1.235 $Y=1.295
+ $X2=1.235 $Y2=1.665
r43 14 20 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.2 $Y=1.32
+ $X2=1.2 $Y2=1.32
r44 13 14 16.4002 $w=2.58e-07 $l=3.7e-07 $layer=LI1_cond $X=1.235 $Y=0.925
+ $X2=1.235 $Y2=1.295
r45 11 20 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.2 $Y=1.66 $X2=1.2
+ $Y2=1.32
r46 11 12 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.2 $Y=1.66 $X2=1.2
+ $Y2=1.825
r47 10 20 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.2 $Y=1.155
+ $X2=1.2 $Y2=1.32
r48 7 12 384.574 $w=1.5e-07 $l=7.5e-07 $layer=POLY_cond $X=1.11 $Y=2.575
+ $X2=1.11 $Y2=1.825
r49 3 10 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=1.11 $Y=0.445
+ $X2=1.11 $Y2=1.155
.ends

.subckt PM_SKY130_FD_SC_LP__OR2_0%A_76_473# 1 2 7 9 13 16 20 22 23 28 30 31 35
+ 36 39 42 44
c70 20 0 3.06547e-19 $X=1.68 $Y=0.84
r71 39 41 8.69362 $w=2.58e-07 $l=1.65e-07 $layer=LI1_cond $X=0.895 $Y=0.445
+ $X2=0.895 $Y2=0.61
r72 36 44 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=1.792 $Y=1.67
+ $X2=1.792 $Y2=1.505
r73 35 36 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.77
+ $Y=1.67 $X2=1.77 $Y2=1.67
r74 33 35 13.7882 $w=2.78e-07 $l=3.35e-07 $layer=LI1_cond $X=1.745 $Y=2.005
+ $X2=1.745 $Y2=1.67
r75 32 42 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.935 $Y=2.09
+ $X2=0.85 $Y2=2.09
r76 31 33 7.36005 $w=1.7e-07 $l=1.77482e-07 $layer=LI1_cond $X=1.605 $Y=2.09
+ $X2=1.745 $Y2=2.005
r77 31 32 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.605 $Y=2.09
+ $X2=0.935 $Y2=2.09
r78 29 42 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.85 $Y=2.175
+ $X2=0.85 $Y2=2.09
r79 29 30 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=0.85 $Y=2.175
+ $X2=0.85 $Y2=2.41
r80 28 42 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.85 $Y=2.005
+ $X2=0.85 $Y2=2.09
r81 28 41 91.0107 $w=1.68e-07 $l=1.395e-06 $layer=LI1_cond $X=0.85 $Y=2.005
+ $X2=0.85 $Y2=0.61
r82 23 30 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.765 $Y=2.575
+ $X2=0.85 $Y2=2.41
r83 23 25 9.07985 $w=3.28e-07 $l=2.6e-07 $layer=LI1_cond $X=0.765 $Y=2.575
+ $X2=0.505 $Y2=2.575
r84 18 20 71.7872 $w=1.5e-07 $l=1.4e-07 $layer=POLY_cond $X=1.54 $Y=0.84
+ $X2=1.68 $Y2=0.84
r85 16 22 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=1.88 $Y=2.685
+ $X2=1.88 $Y2=2.175
r86 13 22 44.7816 $w=3.75e-07 $l=1.87e-07 $layer=POLY_cond $X=1.792 $Y=1.988
+ $X2=1.792 $Y2=2.175
r87 12 36 3.26277 $w=3.75e-07 $l=2.2e-08 $layer=POLY_cond $X=1.792 $Y=1.692
+ $X2=1.792 $Y2=1.67
r88 12 13 43.8991 $w=3.75e-07 $l=2.96e-07 $layer=POLY_cond $X=1.792 $Y=1.692
+ $X2=1.792 $Y2=1.988
r89 10 20 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.68 $Y=0.915
+ $X2=1.68 $Y2=0.84
r90 10 44 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=1.68 $Y=0.915
+ $X2=1.68 $Y2=1.505
r91 7 18 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.54 $Y=0.765
+ $X2=1.54 $Y2=0.84
r92 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.54 $Y=0.765 $X2=1.54
+ $Y2=0.445
r93 2 25 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=0.38
+ $Y=2.365 $X2=0.505 $Y2=2.575
r94 1 39 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.755
+ $Y=0.235 $X2=0.895 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__OR2_0%VPWR 1 6 9 11 18 19 22
r24 22 23 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r25 19 23 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r26 18 19 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r27 16 22 12.8484 $w=1.7e-07 $l=3.13e-07 $layer=LI1_cond $X=1.785 $Y=3.33
+ $X2=1.472 $Y2=3.33
r28 16 18 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.785 $Y=3.33
+ $X2=2.16 $Y2=3.33
r29 13 14 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r30 11 22 12.8484 $w=1.7e-07 $l=3.12e-07 $layer=LI1_cond $X=1.16 $Y=3.33
+ $X2=1.472 $Y2=3.33
r31 11 13 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=1.16 $Y=3.33
+ $X2=0.24 $Y2=3.33
r32 9 23 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33 $X2=1.68
+ $Y2=3.33
r33 9 14 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33 $X2=0.24
+ $Y2=3.33
r34 9 22 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r35 4 22 2.61429 $w=6.25e-07 $l=8.5e-08 $layer=LI1_cond $X=1.472 $Y=3.245
+ $X2=1.472 $Y2=3.33
r36 4 6 14.0659 $w=6.23e-07 $l=7.35e-07 $layer=LI1_cond $X=1.472 $Y=3.245
+ $X2=1.472 $Y2=2.51
r37 1 6 400 $w=1.7e-07 $l=5.47723e-07 $layer=licon1_PDIFF $count=1 $X=1.185
+ $Y=2.365 $X2=1.665 $Y2=2.51
r38 1 6 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.185
+ $Y=2.365 $X2=1.325 $Y2=2.51
.ends

.subckt PM_SKY130_FD_SC_LP__OR2_0%X 1 2 7 11 12 13 14 15 16 17 26 44
r24 44 45 2.8292 $w=3.58e-07 $l=6e-08 $layer=LI1_cond $X=2.135 $Y=2.405
+ $X2=2.135 $Y2=2.345
r25 37 48 0.480185 $w=3.58e-07 $l=1.5e-08 $layer=LI1_cond $X=2.135 $Y=2.525
+ $X2=2.135 $Y2=2.51
r26 17 37 8.00308 $w=3.58e-07 $l=2.5e-07 $layer=LI1_cond $X=2.135 $Y=2.775
+ $X2=2.135 $Y2=2.525
r27 16 48 2.97714 $w=3.58e-07 $l=9.3e-08 $layer=LI1_cond $X=2.135 $Y=2.417
+ $X2=2.135 $Y2=2.51
r28 16 44 0.384148 $w=3.58e-07 $l=1.2e-08 $layer=LI1_cond $X=2.135 $Y=2.417
+ $X2=2.135 $Y2=2.405
r29 16 45 0.576222 $w=2.58e-07 $l=1.3e-08 $layer=LI1_cond $X=2.185 $Y=2.332
+ $X2=2.185 $Y2=2.345
r30 15 16 13.1644 $w=2.58e-07 $l=2.97e-07 $layer=LI1_cond $X=2.185 $Y=2.035
+ $X2=2.185 $Y2=2.332
r31 14 15 16.4002 $w=2.58e-07 $l=3.7e-07 $layer=LI1_cond $X=2.185 $Y=1.665
+ $X2=2.185 $Y2=2.035
r32 13 14 16.4002 $w=2.58e-07 $l=3.7e-07 $layer=LI1_cond $X=2.185 $Y=1.295
+ $X2=2.185 $Y2=1.665
r33 12 13 16.4002 $w=2.58e-07 $l=3.7e-07 $layer=LI1_cond $X=2.185 $Y=0.925
+ $X2=2.185 $Y2=1.295
r34 12 26 11.0812 $w=2.58e-07 $l=2.5e-07 $layer=LI1_cond $X=2.185 $Y=0.925
+ $X2=2.185 $Y2=0.675
r35 11 26 4.34634 $w=2.6e-07 $l=1.98e-07 $layer=LI1_cond $X=2.185 $Y=0.477
+ $X2=2.185 $Y2=0.675
r36 7 11 2.85366 $w=3.95e-07 $l=1.3e-07 $layer=LI1_cond $X=2.055 $Y=0.477
+ $X2=2.185 $Y2=0.477
r37 7 9 8.75273 $w=3.93e-07 $l=3e-07 $layer=LI1_cond $X=2.055 $Y=0.477 $X2=1.755
+ $Y2=0.477
r38 2 48 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=1.955
+ $Y=2.365 $X2=2.095 $Y2=2.51
r39 1 9 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.615
+ $Y=0.235 $X2=1.755 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__OR2_0%VGND 1 2 9 11 15 17 18 19 26 27 30
c32 27 0 1.33616e-19 $X=2.16 $Y=0
c33 26 0 1.72931e-19 $X=2.16 $Y=0
r34 26 27 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r35 24 30 7.13466 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=1.45 $Y=0 $X2=1.322
+ $Y2=0
r36 24 26 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=1.45 $Y=0 $X2=2.16
+ $Y2=0
r37 22 23 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r38 19 27 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r39 19 23 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.24
+ $Y2=0
r40 19 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r41 17 22 4.30588 $w=1.7e-07 $l=6e-08 $layer=LI1_cond $X=0.3 $Y=0 $X2=0.24 $Y2=0
r42 17 18 7.94884 $w=1.7e-07 $l=1.47e-07 $layer=LI1_cond $X=0.3 $Y=0 $X2=0.447
+ $Y2=0
r43 13 30 0.067832 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=1.322 $Y=0.085
+ $X2=1.322 $Y2=0
r44 13 15 16.2698 $w=2.53e-07 $l=3.6e-07 $layer=LI1_cond $X=1.322 $Y=0.085
+ $X2=1.322 $Y2=0.445
r45 12 18 7.94884 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=0.595 $Y=0 $X2=0.447
+ $Y2=0
r46 11 30 7.13466 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=1.195 $Y=0 $X2=1.322
+ $Y2=0
r47 11 12 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=1.195 $Y=0 $X2=0.595
+ $Y2=0
r48 7 18 0.543863 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=0.447 $Y=0.085
+ $X2=0.447 $Y2=0
r49 7 9 14.0637 $w=2.93e-07 $l=3.6e-07 $layer=LI1_cond $X=0.447 $Y=0.085
+ $X2=0.447 $Y2=0.445
r50 2 15 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.185
+ $Y=0.235 $X2=1.325 $Y2=0.445
r51 1 9 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.34
+ $Y=0.235 $X2=0.465 $Y2=0.445
.ends

