* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__a32oi_lp A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
X0 a_56_409# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X1 VPWR A2 a_56_409# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X2 a_56_409# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X3 a_465_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 Y B1 a_56_409# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X5 VGND B2 a_140_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 Y A1 a_357_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 a_56_409# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X8 a_357_47# A2 a_465_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 a_140_47# B1 Y VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
