* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__dfbbp_1 CLK D RESET_B SET_B VGND VNB VPB VPWR Q Q_N
X0 a_755_463# a_767_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X1 a_1823_430# a_1091_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X2 a_531_47# a_225_47# a_617_47# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X3 a_1499_98# a_1545_332# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 VGND D a_531_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 a_1091_21# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X6 VGND a_2317_367# Q VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X7 a_1545_332# a_1307_428# a_1823_430# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X8 a_225_47# a_114_57# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 a_1307_428# a_225_47# a_1419_512# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X10 a_1545_332# a_1091_21# a_1705_54# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X11 a_767_21# a_1091_21# a_917_47# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X12 a_617_47# a_114_57# a_755_463# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X13 a_767_21# a_617_47# a_1046_379# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X14 a_2317_367# a_1545_332# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X15 a_1307_428# a_114_57# a_1499_98# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X16 VPWR a_1545_332# Q_N VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X17 a_1319_54# a_225_47# a_1307_428# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X18 a_2317_367# a_1545_332# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X19 a_1046_379# a_1091_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X20 VPWR SET_B a_1545_332# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X21 a_1212_379# a_114_57# a_1307_428# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X22 a_719_47# a_767_21# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X23 a_225_47# a_114_57# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X24 a_1419_512# a_1545_332# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X25 a_1091_21# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X26 VPWR SET_B a_767_21# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X27 VPWR a_2317_367# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X28 VGND CLK a_114_57# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X29 VPWR D a_531_47# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X30 VPWR a_767_21# a_1212_379# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X31 a_531_47# a_114_57# a_617_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X32 VGND a_767_21# a_1319_54# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X33 VGND a_1545_332# Q_N VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X34 VGND SET_B a_917_47# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X35 VGND SET_B a_1705_54# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X36 a_917_47# a_617_47# a_767_21# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X37 VPWR CLK a_114_57# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X38 a_617_47# a_225_47# a_719_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X39 a_1705_54# a_1307_428# a_1545_332# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
.ends
