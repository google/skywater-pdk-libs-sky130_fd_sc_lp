* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__o2111a_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
X0 a_289_65# B1 a_389_65# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X1 a_32_367# D1 a_32_65# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X2 a_389_65# B1 a_289_65# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X3 X a_32_367# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X4 VPWR B1 a_32_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X5 a_289_65# C1 a_32_65# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X6 VPWR a_32_367# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X7 a_741_367# A2 a_32_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X8 VPWR A1 a_741_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X9 X a_32_367# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X10 VGND a_32_367# X VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X11 a_32_367# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X12 a_32_65# C1 a_289_65# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X13 VPWR a_32_367# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X14 X a_32_367# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X15 a_32_367# A2 a_741_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X16 a_389_65# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X17 VPWR C1 a_32_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X18 X a_32_367# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X19 VGND A2 a_389_65# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X20 a_32_367# D1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X21 a_389_65# A1 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X22 a_32_65# D1 a_32_367# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X23 VGND A1 a_389_65# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X24 a_32_367# C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X25 VPWR D1 a_32_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X26 a_741_367# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X27 VGND a_32_367# X VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
.ends
