# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_sc_lp__ebufn_lp2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_lp__ebufn_lp2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.840000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.376000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.545000 0.440000 0.875000 1.435000 ;
    END
  END A
  PIN TE_B
    ANTENNAGATEAREA  0.626000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.525000 1.605000 3.235000 2.150000 ;
    END
  END TE_B
  PIN Z
    ANTENNADIFFAREA  0.404700 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.670000 1.075000 2.000000 1.605000 ;
        RECT 1.670000 1.605000 2.275000 1.775000 ;
        RECT 1.820000 2.075000 2.275000 3.065000 ;
        RECT 2.045000 1.775000 2.275000 2.075000 ;
    END
  END Z
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.840000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.000000 0.000000 3.840000 0.245000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.655000 1.350000 1.915000 ;
        RECT -0.190000 1.915000 4.030000 3.520000 ;
        RECT  2.715000 1.655000 4.030000 1.915000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.840000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.840000 0.085000 ;
      RECT 0.000000  3.245000 3.840000 3.415000 ;
      RECT 0.115000  0.265000 0.365000 1.675000 ;
      RECT 0.115000  1.675000 1.490000 1.845000 ;
      RECT 0.115000  1.845000 0.445000 3.065000 ;
      RECT 0.645000  2.025000 0.975000 3.245000 ;
      RECT 1.055000  0.085000 1.385000 0.545000 ;
      RECT 1.160000  0.725000 2.350000 0.895000 ;
      RECT 1.160000  0.895000 1.490000 1.485000 ;
      RECT 1.160000  1.845000 1.490000 2.395000 ;
      RECT 2.180000  0.895000 2.350000 1.255000 ;
      RECT 2.180000  1.255000 3.725000 1.425000 ;
      RECT 2.575000  0.085000 2.905000 1.075000 ;
      RECT 2.840000  2.330000 3.170000 3.245000 ;
      RECT 3.370000  2.330000 3.725000 3.065000 ;
      RECT 3.395000  0.745000 3.725000 1.255000 ;
      RECT 3.555000  1.425000 3.725000 2.330000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
  END
END sky130_fd_sc_lp__ebufn_lp2
END LIBRARY
