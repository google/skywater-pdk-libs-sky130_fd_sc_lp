* File: sky130_fd_sc_lp__a2111o_2.pex.spice
* Created: Wed Sep  2 09:16:19 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A2111O_2%A_86_275# 1 2 3 12 14 16 19 21 23 27 29 30
+ 31 32 33 35 39 41 45 49 53
r94 52 53 12.2413 $w=3.15e-07 $l=8e-08 $layer=POLY_cond $X=0.935 $Y=1.36
+ $X2=1.015 $Y2=1.36
r95 51 52 53.5556 $w=3.15e-07 $l=3.5e-07 $layer=POLY_cond $X=0.585 $Y=1.36
+ $X2=0.935 $Y2=1.36
r96 43 45 27.5175 $w=2.43e-07 $l=5.85e-07 $layer=LI1_cond $X=3.212 $Y=1.005
+ $X2=3.212 $Y2=0.42
r97 42 49 6.81202 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=2.42 $Y=1.09 $X2=2.3
+ $Y2=1.09
r98 41 43 7.11011 $w=1.7e-07 $l=1.58915e-07 $layer=LI1_cond $X=3.09 $Y=1.09
+ $X2=3.212 $Y2=1.005
r99 41 42 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.09 $Y=1.09
+ $X2=2.42 $Y2=1.09
r100 37 49 0.135687 $w=2.4e-07 $l=8.5e-08 $layer=LI1_cond $X=2.3 $Y=1.005
+ $X2=2.3 $Y2=1.09
r101 37 39 28.0908 $w=2.38e-07 $l=5.85e-07 $layer=LI1_cond $X=2.3 $Y=1.005
+ $X2=2.3 $Y2=0.42
r102 33 48 2.68691 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=1.845 $Y=2.1 $X2=1.845
+ $Y2=2.01
r103 33 35 29.6841 $w=3.28e-07 $l=8.5e-07 $layer=LI1_cond $X=1.845 $Y=2.1
+ $X2=1.845 $Y2=2.95
r104 31 48 4.92601 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=1.68 $Y=2.01
+ $X2=1.845 $Y2=2.01
r105 31 32 16.3283 $w=1.78e-07 $l=2.65e-07 $layer=LI1_cond $X=1.68 $Y=2.01
+ $X2=1.415 $Y2=2.01
r106 29 49 6.81202 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=2.18 $Y=1.09 $X2=2.3
+ $Y2=1.09
r107 29 30 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=2.18 $Y=1.09
+ $X2=1.415 $Y2=1.09
r108 28 53 35.9587 $w=3.15e-07 $l=2.35e-07 $layer=POLY_cond $X=1.25 $Y=1.36
+ $X2=1.015 $Y2=1.36
r109 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.25
+ $Y=1.36 $X2=1.25 $Y2=1.36
r110 25 32 7.77087 $w=1.8e-07 $l=2.15349e-07 $layer=LI1_cond $X=1.24 $Y=1.92
+ $X2=1.415 $Y2=2.01
r111 25 27 18.4391 $w=3.48e-07 $l=5.6e-07 $layer=LI1_cond $X=1.24 $Y=1.92
+ $X2=1.24 $Y2=1.36
r112 24 30 7.93686 $w=1.7e-07 $l=2.13307e-07 $layer=LI1_cond $X=1.24 $Y=1.175
+ $X2=1.415 $Y2=1.09
r113 24 27 6.09148 $w=3.48e-07 $l=1.85e-07 $layer=LI1_cond $X=1.24 $Y=1.175
+ $X2=1.24 $Y2=1.36
r114 21 53 20.1192 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.015 $Y=1.195
+ $X2=1.015 $Y2=1.36
r115 21 23 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.015 $Y=1.195
+ $X2=1.015 $Y2=0.665
r116 17 52 20.1192 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.935 $Y=1.525
+ $X2=0.935 $Y2=1.36
r117 17 19 482 $w=1.5e-07 $l=9.4e-07 $layer=POLY_cond $X=0.935 $Y=1.525
+ $X2=0.935 $Y2=2.465
r118 14 51 20.1192 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.585 $Y=1.195
+ $X2=0.585 $Y2=1.36
r119 14 16 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.585 $Y=1.195
+ $X2=0.585 $Y2=0.665
r120 10 51 12.2413 $w=3.15e-07 $l=2.0106e-07 $layer=POLY_cond $X=0.505 $Y=1.525
+ $X2=0.585 $Y2=1.36
r121 10 12 482 $w=1.5e-07 $l=9.4e-07 $layer=POLY_cond $X=0.505 $Y=1.525
+ $X2=0.505 $Y2=2.465
r122 3 48 400 $w=1.7e-07 $l=2.23942e-07 $layer=licon1_PDIFF $count=1 $X=1.72
+ $Y=1.835 $X2=1.845 $Y2=2.005
r123 3 35 400 $w=1.7e-07 $l=1.17584e-06 $layer=licon1_PDIFF $count=1 $X=1.72
+ $Y=1.835 $X2=1.845 $Y2=2.95
r124 2 45 91 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=2 $X=3.09
+ $Y=0.245 $X2=3.23 $Y2=0.42
r125 1 39 91 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=2 $X=2.135
+ $Y=0.245 $X2=2.275 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__A2111O_2%D1 3 7 9 10 14
r35 14 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.97 $Y=1.51
+ $X2=1.97 $Y2=1.675
r36 14 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.97 $Y=1.51
+ $X2=1.97 $Y2=1.345
r37 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.97
+ $Y=1.51 $X2=1.97 $Y2=1.51
r38 10 15 5.40652 $w=4.03e-07 $l=1.9e-07 $layer=LI1_cond $X=2.16 $Y=1.547
+ $X2=1.97 $Y2=1.547
r39 9 15 8.25206 $w=4.03e-07 $l=2.9e-07 $layer=LI1_cond $X=1.68 $Y=1.547
+ $X2=1.97 $Y2=1.547
r40 7 17 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.06 $Y=2.465
+ $X2=2.06 $Y2=1.675
r41 3 16 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=2.06 $Y=0.665
+ $X2=2.06 $Y2=1.345
.ends

.subckt PM_SKY130_FD_SC_LP__A2111O_2%C1 3 7 9 10 11 12 18 19
c38 3 0 5.59569e-20 $X=2.42 $Y=2.465
r39 18 21 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.51 $Y=1.51
+ $X2=2.51 $Y2=1.675
r40 18 20 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.51 $Y=1.51
+ $X2=2.51 $Y2=1.345
r41 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.51
+ $Y=1.51 $X2=2.51 $Y2=1.51
r42 11 12 11.5244 $w=3.68e-07 $l=3.7e-07 $layer=LI1_cond $X=2.61 $Y=2.405
+ $X2=2.61 $Y2=2.775
r43 10 11 11.5244 $w=3.68e-07 $l=3.7e-07 $layer=LI1_cond $X=2.61 $Y=2.035
+ $X2=2.61 $Y2=2.405
r44 9 10 11.5244 $w=3.68e-07 $l=3.7e-07 $layer=LI1_cond $X=2.61 $Y=1.665
+ $X2=2.61 $Y2=2.035
r45 9 19 4.8278 $w=3.68e-07 $l=1.55e-07 $layer=LI1_cond $X=2.61 $Y=1.665
+ $X2=2.61 $Y2=1.51
r46 7 20 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=2.49 $Y=0.665
+ $X2=2.49 $Y2=1.345
r47 3 21 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.42 $Y=2.465
+ $X2=2.42 $Y2=1.675
.ends

.subckt PM_SKY130_FD_SC_LP__A2111O_2%B1 3 7 9 12 13
c30 13 0 5.59569e-20 $X=3.05 $Y=1.51
c31 3 0 5.87692e-20 $X=2.96 $Y=2.465
r32 12 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.05 $Y=1.51
+ $X2=3.05 $Y2=1.675
r33 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.05 $Y=1.51
+ $X2=3.05 $Y2=1.345
r34 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.05
+ $Y=1.51 $X2=3.05 $Y2=1.51
r35 9 13 5.17764 $w=3.43e-07 $l=1.55e-07 $layer=LI1_cond $X=3.137 $Y=1.665
+ $X2=3.137 $Y2=1.51
r36 7 14 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=3.015 $Y=0.665
+ $X2=3.015 $Y2=1.345
r37 3 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.96 $Y=2.465
+ $X2=2.96 $Y2=1.675
.ends

.subckt PM_SKY130_FD_SC_LP__A2111O_2%A1 3 6 8 9 10 11 17 19
c39 8 0 5.87692e-20 $X=3.6 $Y=0.555
r40 17 20 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.59 $Y=1.36
+ $X2=3.59 $Y2=1.525
r41 17 19 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.59 $Y=1.36
+ $X2=3.59 $Y2=1.195
r42 10 11 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=3.64 $Y=1.295
+ $X2=3.64 $Y2=1.665
r43 10 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.59
+ $Y=1.36 $X2=3.59 $Y2=1.36
r44 9 10 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=3.64 $Y=0.925
+ $X2=3.64 $Y2=1.295
r45 8 9 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=3.64 $Y=0.555 $X2=3.64
+ $Y2=0.925
r46 6 20 482 $w=1.5e-07 $l=9.4e-07 $layer=POLY_cond $X=3.5 $Y=2.465 $X2=3.5
+ $Y2=1.525
r47 3 19 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=3.5 $Y=0.665 $X2=3.5
+ $Y2=1.195
.ends

.subckt PM_SKY130_FD_SC_LP__A2111O_2%A2 3 6 8 10 17 19
r28 17 20 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.13 $Y=1.375
+ $X2=4.13 $Y2=1.54
r29 17 19 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.13 $Y=1.375
+ $X2=4.13 $Y2=1.21
r30 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.13
+ $Y=1.375 $X2=4.13 $Y2=1.375
r31 10 18 9.52433 $w=5.38e-07 $l=4.3e-07 $layer=LI1_cond $X=4.56 $Y=1.48
+ $X2=4.13 $Y2=1.48
r32 8 18 1.10748 $w=5.38e-07 $l=5e-08 $layer=LI1_cond $X=4.08 $Y=1.48 $X2=4.13
+ $Y2=1.48
r33 6 20 474.309 $w=1.5e-07 $l=9.25e-07 $layer=POLY_cond $X=4.04 $Y=2.465
+ $X2=4.04 $Y2=1.54
r34 3 19 175.127 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=4.04 $Y=0.665
+ $X2=4.04 $Y2=1.21
.ends

.subckt PM_SKY130_FD_SC_LP__A2111O_2%VPWR 1 2 3 10 12 18 22 25 26 27 29 42 43 49
r55 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r56 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r57 42 43 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r58 40 43 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.56 $Y2=3.33
r59 39 40 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r60 37 50 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r61 36 39 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=1.68 $Y=3.33
+ $X2=3.6 $Y2=3.33
r62 36 37 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r63 34 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.315 $Y=3.33
+ $X2=1.15 $Y2=3.33
r64 34 36 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=1.315 $Y=3.33
+ $X2=1.68 $Y2=3.33
r65 33 50 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r66 33 47 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r67 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r68 30 46 4.70928 $w=1.7e-07 $l=2.28e-07 $layer=LI1_cond $X=0.455 $Y=3.33
+ $X2=0.227 $Y2=3.33
r69 30 32 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.455 $Y=3.33
+ $X2=0.72 $Y2=3.33
r70 29 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.985 $Y=3.33
+ $X2=1.15 $Y2=3.33
r71 29 32 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.985 $Y=3.33
+ $X2=0.72 $Y2=3.33
r72 27 40 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=2.4 $Y=3.33 $X2=3.6
+ $Y2=3.33
r73 27 37 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.4 $Y=3.33
+ $X2=1.68 $Y2=3.33
r74 25 39 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=3.605 $Y=3.33 $X2=3.6
+ $Y2=3.33
r75 25 26 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.605 $Y=3.33
+ $X2=3.77 $Y2=3.33
r76 24 42 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=3.935 $Y=3.33
+ $X2=4.56 $Y2=3.33
r77 24 26 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.935 $Y=3.33
+ $X2=3.77 $Y2=3.33
r78 20 26 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.77 $Y=3.245
+ $X2=3.77 $Y2=3.33
r79 20 22 29.8588 $w=3.28e-07 $l=8.55e-07 $layer=LI1_cond $X=3.77 $Y=3.245
+ $X2=3.77 $Y2=2.39
r80 16 49 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.15 $Y=3.245
+ $X2=1.15 $Y2=3.33
r81 16 18 29.8588 $w=3.28e-07 $l=8.55e-07 $layer=LI1_cond $X=1.15 $Y=3.245
+ $X2=1.15 $Y2=2.39
r82 12 15 33.8748 $w=3.28e-07 $l=9.7e-07 $layer=LI1_cond $X=0.29 $Y=1.98
+ $X2=0.29 $Y2=2.95
r83 10 46 3.0569 $w=3.3e-07 $l=1.12161e-07 $layer=LI1_cond $X=0.29 $Y=3.245
+ $X2=0.227 $Y2=3.33
r84 10 15 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.29 $Y=3.245
+ $X2=0.29 $Y2=2.95
r85 3 22 300 $w=1.7e-07 $l=6.45174e-07 $layer=licon1_PDIFF $count=2 $X=3.575
+ $Y=1.835 $X2=3.77 $Y2=2.39
r86 2 18 300 $w=1.7e-07 $l=6.21068e-07 $layer=licon1_PDIFF $count=2 $X=1.01
+ $Y=1.835 $X2=1.15 $Y2=2.39
r87 1 15 400 $w=1.7e-07 $l=1.17584e-06 $layer=licon1_PDIFF $count=1 $X=0.165
+ $Y=1.835 $X2=0.29 $Y2=2.95
r88 1 12 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.165
+ $Y=1.835 $X2=0.29 $Y2=1.98
.ends

.subckt PM_SKY130_FD_SC_LP__A2111O_2%X 1 2 7 8 9 10 11 12 13 25 47
r18 47 48 3.80025 $w=2.68e-07 $l=6.5e-08 $layer=LI1_cond $X=0.76 $Y=2.035
+ $X2=0.76 $Y2=2.1
r19 12 13 26.5598 $w=1.88e-07 $l=4.55e-07 $layer=LI1_cond $X=0.72 $Y=2.32
+ $X2=0.72 $Y2=2.775
r20 11 47 2.34757 $w=2.68e-07 $l=5.5e-08 $layer=LI1_cond $X=0.76 $Y=1.98
+ $X2=0.76 $Y2=2.035
r21 11 23 0.640246 $w=2.68e-07 $l=1.5e-08 $layer=LI1_cond $X=0.76 $Y=1.98
+ $X2=0.76 $Y2=1.965
r22 11 12 12.2584 $w=1.88e-07 $l=2.1e-07 $layer=LI1_cond $X=0.72 $Y=2.11
+ $X2=0.72 $Y2=2.32
r23 11 48 0.583732 $w=1.88e-07 $l=1e-08 $layer=LI1_cond $X=0.72 $Y=2.11 $X2=0.72
+ $Y2=2.1
r24 11 23 0.341465 $w=2.68e-07 $l=8e-09 $layer=LI1_cond $X=0.76 $Y=1.957
+ $X2=0.76 $Y2=1.965
r25 10 11 12.4635 $w=2.68e-07 $l=2.92e-07 $layer=LI1_cond $X=0.76 $Y=1.665
+ $X2=0.76 $Y2=1.957
r26 9 10 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.76 $Y=1.295
+ $X2=0.76 $Y2=1.665
r27 8 9 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.76 $Y=0.925 $X2=0.76
+ $Y2=1.295
r28 7 8 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.76 $Y=0.555 $X2=0.76
+ $Y2=0.925
r29 7 25 5.76222 $w=2.68e-07 $l=1.35e-07 $layer=LI1_cond $X=0.76 $Y=0.555
+ $X2=0.76 $Y2=0.42
r30 2 11 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.58
+ $Y=1.835 $X2=0.72 $Y2=1.98
r31 2 12 300 $w=1.7e-07 $l=5.50568e-07 $layer=licon1_PDIFF $count=2 $X=0.58
+ $Y=1.835 $X2=0.72 $Y2=2.32
r32 1 25 91 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=2 $X=0.66
+ $Y=0.245 $X2=0.8 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__A2111O_2%A_607_367# 1 2 7 9 11 13 15
r22 13 20 2.68365 $w=3.15e-07 $l=8.5e-08 $layer=LI1_cond $X=4.262 $Y=2.1
+ $X2=4.262 $Y2=2.015
r23 13 15 29.6342 $w=3.13e-07 $l=8.1e-07 $layer=LI1_cond $X=4.262 $Y=2.1
+ $X2=4.262 $Y2=2.91
r24 12 18 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.4 $Y=2.015
+ $X2=3.235 $Y2=2.015
r25 11 20 4.95685 $w=1.7e-07 $l=1.57e-07 $layer=LI1_cond $X=4.105 $Y=2.015
+ $X2=4.262 $Y2=2.015
r26 11 12 45.9947 $w=1.68e-07 $l=7.05e-07 $layer=LI1_cond $X=4.105 $Y=2.015
+ $X2=3.4 $Y2=2.015
r27 7 18 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.235 $Y=2.1 $X2=3.235
+ $Y2=2.015
r28 7 9 13.0959 $w=3.28e-07 $l=3.75e-07 $layer=LI1_cond $X=3.235 $Y=2.1
+ $X2=3.235 $Y2=2.475
r29 2 20 400 $w=1.7e-07 $l=2.4e-07 $layer=licon1_PDIFF $count=1 $X=4.115
+ $Y=1.835 $X2=4.255 $Y2=2.015
r30 2 15 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=4.115
+ $Y=1.835 $X2=4.255 $Y2=2.91
r31 1 18 600 $w=1.7e-07 $l=2.75681e-07 $layer=licon1_PDIFF $count=1 $X=3.035
+ $Y=1.835 $X2=3.235 $Y2=2.015
r32 1 9 300 $w=1.7e-07 $l=7.33212e-07 $layer=licon1_PDIFF $count=2 $X=3.035
+ $Y=1.835 $X2=3.235 $Y2=2.475
.ends

.subckt PM_SKY130_FD_SC_LP__A2111O_2%VGND 1 2 3 4 13 15 17 21 25 28 29 30 45 46
+ 54 60 62
r59 62 63 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r60 59 60 12.3913 $w=9.18e-07 $l=1.65e-07 $layer=LI1_cond $X=1.845 $Y=0.375
+ $X2=2.01 $Y2=0.375
r61 56 59 2.18804 $w=9.18e-07 $l=1.65e-07 $layer=LI1_cond $X=1.68 $Y=0.375
+ $X2=1.845 $Y2=0.375
r62 56 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r63 53 57 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r64 52 56 6.36522 $w=9.18e-07 $l=4.8e-07 $layer=LI1_cond $X=1.2 $Y=0.375
+ $X2=1.68 $Y2=0.375
r65 52 54 11.9934 $w=9.18e-07 $l=1.35e-07 $layer=LI1_cond $X=1.2 $Y=0.375
+ $X2=1.065 $Y2=0.375
r66 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r67 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r68 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r69 43 46 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=4.56
+ $Y2=0
r70 42 43 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r71 40 43 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=4.08
+ $Y2=0
r72 40 63 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.64
+ $Y2=0
r73 39 42 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=3.12 $Y=0 $X2=4.08
+ $Y2=0
r74 39 40 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r75 37 62 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.92 $Y=0 $X2=2.755
+ $Y2=0
r76 37 39 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=2.92 $Y=0 $X2=3.12
+ $Y2=0
r77 36 53 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r78 36 50 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r79 35 54 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.72 $Y=0 $X2=1.065
+ $Y2=0
r80 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r81 33 49 3.915 $w=1.7e-07 $l=2.28e-07 $layer=LI1_cond $X=0.455 $Y=0 $X2=0.227
+ $Y2=0
r82 33 35 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.455 $Y=0 $X2=0.72
+ $Y2=0
r83 30 63 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.4 $Y=0 $X2=2.64
+ $Y2=0
r84 30 57 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.4 $Y=0 $X2=1.68
+ $Y2=0
r85 28 42 0.652406 $w=1.68e-07 $l=1e-08 $layer=LI1_cond $X=4.09 $Y=0 $X2=4.08
+ $Y2=0
r86 28 29 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.09 $Y=0 $X2=4.255
+ $Y2=0
r87 27 45 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=4.42 $Y=0 $X2=4.56
+ $Y2=0
r88 27 29 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.42 $Y=0 $X2=4.255
+ $Y2=0
r89 23 29 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.255 $Y=0.085
+ $X2=4.255 $Y2=0
r90 23 25 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=4.255 $Y=0.085
+ $X2=4.255 $Y2=0.39
r91 19 62 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.755 $Y=0.085
+ $X2=2.755 $Y2=0
r92 19 21 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=2.755 $Y=0.085
+ $X2=2.755 $Y2=0.37
r93 17 62 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.59 $Y=0 $X2=2.755
+ $Y2=0
r94 17 60 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=2.59 $Y=0 $X2=2.01
+ $Y2=0
r95 13 49 3.22816 $w=2.5e-07 $l=1.39155e-07 $layer=LI1_cond $X=0.33 $Y=0.085
+ $X2=0.227 $Y2=0
r96 13 15 14.0598 $w=2.48e-07 $l=3.05e-07 $layer=LI1_cond $X=0.33 $Y=0.085
+ $X2=0.33 $Y2=0.39
r97 4 25 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.115
+ $Y=0.245 $X2=4.255 $Y2=0.39
r98 3 21 91 $w=1.7e-07 $l=2.44643e-07 $layer=licon1_NDIFF $count=2 $X=2.565
+ $Y=0.245 $X2=2.755 $Y2=0.37
r99 2 59 45.5 $w=1.7e-07 $l=8.15107e-07 $layer=licon1_NDIFF $count=4 $X=1.09
+ $Y=0.245 $X2=1.845 $Y2=0.37
r100 1 15 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.245
+ $Y=0.245 $X2=0.37 $Y2=0.39
.ends

