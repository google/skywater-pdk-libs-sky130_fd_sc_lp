* File: sky130_fd_sc_lp__decapkapwr_3.pex.spice
* Created: Wed Sep  2 09:42:27 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__DECAPKAPWR_3%VGND 1 7 9 10 13 14 16 19 23 26 36
r31 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r32 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r33 27 32 4.62272 $w=1.7e-07 $l=2.5e-07 $layer=LI1_cond $X=0.5 $Y=0 $X2=0.25
+ $Y2=0
r34 27 29 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=0.5 $Y=0 $X2=0.72
+ $Y2=0
r35 26 35 4.64076 $w=1.7e-07 $l=2.45e-07 $layer=LI1_cond $X=0.95 $Y=0 $X2=1.195
+ $Y2=0
r36 26 29 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=0.95 $Y=0 $X2=0.72
+ $Y2=0
r37 23 36 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r38 23 33 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r39 23 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r40 19 21 5.30815 $w=4.88e-07 $l=1.65e-07 $layer=LI1_cond $X=0.415 $Y=1.77
+ $X2=0.415 $Y2=1.605
r41 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.575
+ $Y=1.77 $X2=0.575 $Y2=1.77
r42 14 35 3.12541 $w=3.3e-07 $l=1.18427e-07 $layer=LI1_cond $X=1.115 $Y=0.085
+ $X2=1.195 $Y2=0
r43 14 16 13.0959 $w=3.28e-07 $l=3.75e-07 $layer=LI1_cond $X=1.115 $Y=0.085
+ $X2=1.115 $Y2=0.46
r44 13 21 39.2878 $w=3.28e-07 $l=1.125e-06 $layer=LI1_cond $X=0.335 $Y=0.48
+ $X2=0.335 $Y2=1.605
r45 10 32 3.14345 $w=3.3e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.335 $Y=0.085
+ $X2=0.25 $Y2=0
r46 10 13 13.7944 $w=3.28e-07 $l=3.95e-07 $layer=LI1_cond $X=0.335 $Y=0.085
+ $X2=0.335 $Y2=0.48
r47 7 20 36.8902 $w=5e-07 $l=3.65e-07 $layer=POLY_cond $X=0.66 $Y=2.135 $X2=0.66
+ $Y2=1.77
r48 7 9 44.344 $w=5e-07 $l=4.6e-07 $layer=POLY_cond $X=0.66 $Y=2.135 $X2=0.66
+ $Y2=2.595
r49 1 16 182 $w=1.7e-07 $l=2.86575e-07 $layer=licon1_NDIFF $count=1 $X=0.975
+ $Y=0.235 $X2=1.115 $Y2=0.46
r50 1 13 182 $w=1.7e-07 $l=3.01081e-07 $layer=licon1_NDIFF $count=1 $X=0.975
+ $Y=0.235 $X2=0.335 $Y2=0.48
.ends

.subckt PM_SKY130_FD_SC_LP__DECAPKAPWR_3%KAPWR 1 7 9 10 12 14 17 19 24 26 35
r36 34 35 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.13 $Y=2.81
+ $X2=1.13 $Y2=2.81
r37 30 31 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.215 $Y=2.81
+ $X2=0.215 $Y2=2.81
r38 26 35 0.224086 $w=2.7e-07 $l=4.1e-07 $layer=MET1_cond $X=0.72 $Y=2.81
+ $X2=1.13 $Y2=2.81
r39 26 31 0.276009 $w=2.7e-07 $l=5.05e-07 $layer=MET1_cond $X=0.72 $Y=2.81
+ $X2=0.215 $Y2=2.81
r40 21 24 9.31427 $w=3.63e-07 $l=2.95e-07 $layer=LI1_cond $X=0.755 $Y=1.042
+ $X2=1.05 $Y2=1.042
r41 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.755
+ $Y=1.06 $X2=0.755 $Y2=1.06
r42 17 34 3.21187 $w=3.3e-07 $l=2e-07 $layer=LI1_cond $X=1.05 $Y=2.675 $X2=1.05
+ $Y2=2.875
r43 17 19 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=1.05 $Y=2.675
+ $X2=1.05 $Y2=2.29
r44 16 24 1.32393 $w=3.3e-07 $l=1.83e-07 $layer=LI1_cond $X=1.05 $Y=1.225
+ $X2=1.05 $Y2=1.042
r45 16 19 37.1925 $w=3.28e-07 $l=1.065e-06 $layer=LI1_cond $X=1.05 $Y=1.225
+ $X2=1.05 $Y2=2.29
r46 15 30 3.69365 $w=2.7e-07 $l=1.94808e-07 $layer=LI1_cond $X=0.425 $Y=2.81
+ $X2=0.26 $Y2=2.875
r47 14 34 3.69365 $w=2.7e-07 $l=1.94808e-07 $layer=LI1_cond $X=0.885 $Y=2.81
+ $X2=1.05 $Y2=2.875
r48 14 15 19.6342 $w=2.68e-07 $l=4.6e-07 $layer=LI1_cond $X=0.885 $Y=2.81
+ $X2=0.425 $Y2=2.81
r49 10 30 3.21187 $w=3.3e-07 $l=2e-07 $layer=LI1_cond $X=0.26 $Y=2.675 $X2=0.26
+ $Y2=2.875
r50 10 12 14.1436 $w=3.28e-07 $l=4.05e-07 $layer=LI1_cond $X=0.26 $Y=2.675
+ $X2=0.26 $Y2=2.27
r51 7 22 39.9593 $w=5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.725 $Y=0.665
+ $X2=0.725 $Y2=1.06
r52 7 9 14.942 $w=5e-07 $l=1.55e-07 $layer=POLY_cond $X=0.725 $Y=0.665 $X2=0.725
+ $Y2=0.51
r53 1 34 400 $w=1.7e-07 $l=9.42404e-07 $layer=licon1_PDIFF $count=1 $X=0.91
+ $Y=2.095 $X2=1.05 $Y2=2.97
r54 1 30 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.91
+ $Y=2.095 $X2=0.26 $Y2=2.95
r55 1 19 400 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_PDIFF $count=1 $X=0.91
+ $Y=2.095 $X2=1.05 $Y2=2.29
r56 1 12 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.91
+ $Y=2.095 $X2=0.26 $Y2=2.27
.ends

.subckt PM_SKY130_FD_SC_LP__DECAPKAPWR_3%VPWR 1 8 14
r14 5 14 0.0108064 $w=1.44e-06 $l=1.22e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.208
r15 5 8 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r16 4 8 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.24 $Y=3.33 $X2=1.2
+ $Y2=3.33
r17 4 5 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33 $X2=0.24
+ $Y2=3.33
r18 1 14 8.85771e-05 $w=1.44e-06 $l=1e-09 $layer=MET1_cond $X=0.72 $Y=3.207
+ $X2=0.72 $Y2=3.208
.ends

