* File: sky130_fd_sc_lp__nand2b_m.spice
* Created: Fri Aug 28 10:48:39 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__nand2b_m.pex.spice"
.subckt sky130_fd_sc_lp__nand2b_m  VNB VPB A_N B VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B	B
* A_N	A_N
* VPB	VPB
* VNB	VNB
MM1004 N_VGND_M1004_d N_A_N_M1004_g N_A_46_54#_M1004_s VNB NSHORT L=0.15 W=0.42
+ AD=0.12915 AS=0.1113 PD=1.035 PS=1.37 NRD=87.132 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.3 A=0.063 P=1.14 MULT=1
MM1001 A_282_54# N_B_M1001_g N_VGND_M1004_d VNB NSHORT L=0.15 W=0.42 AD=0.0441
+ AS=0.12915 PD=0.63 PS=1.035 NRD=14.28 NRS=8.568 M=1 R=2.8 SA=75001 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1002 N_Y_M1002_d N_A_46_54#_M1002_g A_282_54# VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.0441 PD=1.37 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.3
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1005 N_VPWR_M1005_d N_A_N_M1005_g N_A_46_54#_M1005_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75001.1
+ A=0.063 P=1.14 MULT=1
MM1003 N_Y_M1003_d N_B_M1003_g N_VPWR_M1005_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1000 N_VPWR_M1000_d N_A_46_54#_M1000_g N_Y_M1003_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.1 SB=75000.2
+ A=0.063 P=1.14 MULT=1
DX6_noxref VNB VPB NWDIODE A=5.1847 P=9.29
c_52 VPB 0 1.69314e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_lp__nand2b_m.pxi.spice"
*
.ends
*
*
