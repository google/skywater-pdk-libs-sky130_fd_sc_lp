* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
X0 VPWR D_N a_196_535# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X1 a_27_535# C_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X2 VGND B a_332_391# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 a_487_391# B a_595_391# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X4 a_595_391# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X5 a_332_391# a_196_535# a_415_391# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X6 a_415_391# a_27_535# a_487_391# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X7 VGND a_196_535# a_332_391# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 a_332_391# A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 a_27_535# C_N VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 VGND a_332_391# X VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X11 a_332_391# a_27_535# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 VPWR a_332_391# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X13 VGND D_N a_196_535# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
