* File: sky130_fd_sc_lp__nor2_1.pxi.spice
* Created: Fri Aug 28 10:53:14 2020
* 
x_PM_SKY130_FD_SC_LP__NOR2_1%A N_A_M1003_g N_A_M1000_g A A N_A_c_30_n N_A_c_31_n
+ PM_SKY130_FD_SC_LP__NOR2_1%A
x_PM_SKY130_FD_SC_LP__NOR2_1%B N_B_M1001_g N_B_c_51_n N_B_M1002_g B B N_B_c_53_n
+ PM_SKY130_FD_SC_LP__NOR2_1%B
x_PM_SKY130_FD_SC_LP__NOR2_1%VPWR N_VPWR_M1000_s N_VPWR_c_76_n N_VPWR_c_77_n
+ VPWR N_VPWR_c_78_n N_VPWR_c_75_n PM_SKY130_FD_SC_LP__NOR2_1%VPWR
x_PM_SKY130_FD_SC_LP__NOR2_1%Y N_Y_M1003_d N_Y_M1001_d Y Y Y Y Y Y Y N_Y_c_98_n
+ PM_SKY130_FD_SC_LP__NOR2_1%Y
x_PM_SKY130_FD_SC_LP__NOR2_1%VGND N_VGND_M1003_s N_VGND_M1002_d N_VGND_c_116_n
+ N_VGND_c_117_n N_VGND_c_118_n N_VGND_c_119_n VGND N_VGND_c_120_n
+ N_VGND_c_121_n PM_SKY130_FD_SC_LP__NOR2_1%VGND
cc_1 VNB N_A_M1000_g 0.00179493f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.465
cc_2 VNB A 0.0211263f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_3 VNB N_A_c_30_n 0.043153f $X=-0.19 $Y=-0.245 $X2=0.35 $Y2=1.46
cc_4 VNB N_A_c_31_n 0.0203861f $X=-0.19 $Y=-0.245 $X2=0.382 $Y2=1.295
cc_5 VNB N_B_M1001_g 0.0015777f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=0.765
cc_6 VNB N_B_c_51_n 0.0203861f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.465
cc_7 VNB B 0.0214155f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_8 VNB N_B_c_53_n 0.046066f $X=-0.19 $Y=-0.245 $X2=0.382 $Y2=1.625
cc_9 VNB N_VPWR_c_75_n 0.0641695f $X=-0.19 $Y=-0.245 $X2=0.382 $Y2=1.295
cc_10 VNB Y 0.0106863f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_VGND_c_116_n 0.0121567f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_VGND_c_117_n 0.0352805f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_13 VNB N_VGND_c_118_n 0.0121567f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_VGND_c_119_n 0.0352805f $X=-0.19 $Y=-0.245 $X2=0.35 $Y2=1.46
cc_15 VNB N_VGND_c_120_n 0.0146145f $X=-0.19 $Y=-0.245 $X2=0.26 $Y2=1.295
cc_16 VNB N_VGND_c_121_n 0.114861f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VPB N_A_M1000_g 0.0249895f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=2.465
cc_18 VPB A 0.007988f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_19 VPB N_B_M1001_g 0.0251437f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=0.765
cc_20 VPB B 0.0100018f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_21 VPB N_VPWR_c_76_n 0.0112967f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=1.625
cc_22 VPB N_VPWR_c_77_n 0.0484529f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=2.465
cc_23 VPB N_VPWR_c_78_n 0.0261756f $X=-0.19 $Y=1.655 $X2=0.35 $Y2=1.46
cc_24 VPB N_VPWR_c_75_n 0.0479422f $X=-0.19 $Y=1.655 $X2=0.382 $Y2=1.295
cc_25 VPB Y 0.0032435f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_26 VPB Y 0.0350453f $X=-0.19 $Y=1.655 $X2=0.382 $Y2=1.46
cc_27 VPB N_Y_c_98_n 0.0139933f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_28 N_A_M1000_g N_B_M1001_g 0.0473735f $X=0.505 $Y=2.465 $X2=0 $Y2=0
cc_29 N_A_c_31_n N_B_c_51_n 0.0130856f $X=0.382 $Y=1.295 $X2=0 $Y2=0
cc_30 N_A_c_30_n N_B_c_53_n 0.0473735f $X=0.35 $Y=1.46 $X2=0 $Y2=0
cc_31 N_A_M1000_g N_VPWR_c_77_n 0.0222058f $X=0.505 $Y=2.465 $X2=0 $Y2=0
cc_32 A N_VPWR_c_77_n 0.0252511f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_33 N_A_c_30_n N_VPWR_c_77_n 0.00129037f $X=0.35 $Y=1.46 $X2=0 $Y2=0
cc_34 N_A_M1000_g N_VPWR_c_78_n 0.00486043f $X=0.505 $Y=2.465 $X2=0 $Y2=0
cc_35 N_A_M1000_g N_VPWR_c_75_n 0.00827383f $X=0.505 $Y=2.465 $X2=0 $Y2=0
cc_36 A Y 0.0377377f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_37 N_A_c_31_n Y 0.0119963f $X=0.382 $Y=1.295 $X2=0 $Y2=0
cc_38 A N_VGND_c_117_n 0.0252511f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_39 N_A_c_30_n N_VGND_c_117_n 0.00141307f $X=0.35 $Y=1.46 $X2=0 $Y2=0
cc_40 N_A_c_31_n N_VGND_c_117_n 0.0146695f $X=0.382 $Y=1.295 $X2=0 $Y2=0
cc_41 N_A_c_31_n N_VGND_c_119_n 5.35643e-19 $X=0.382 $Y=1.295 $X2=0 $Y2=0
cc_42 N_A_c_31_n N_VGND_c_120_n 0.00400407f $X=0.382 $Y=1.295 $X2=0 $Y2=0
cc_43 N_A_c_31_n N_VGND_c_121_n 0.00775088f $X=0.382 $Y=1.295 $X2=0 $Y2=0
cc_44 N_B_M1001_g N_VPWR_c_77_n 0.00206182f $X=0.895 $Y=2.465 $X2=0 $Y2=0
cc_45 N_B_M1001_g N_VPWR_c_78_n 0.00357668f $X=0.895 $Y=2.465 $X2=0 $Y2=0
cc_46 N_B_M1001_g N_VPWR_c_75_n 0.00626226f $X=0.895 $Y=2.465 $X2=0 $Y2=0
cc_47 N_B_c_51_n Y 0.0018192f $X=0.935 $Y=1.295 $X2=0 $Y2=0
cc_48 B Y 0.0417627f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_49 N_B_c_53_n Y 0.00613187f $X=1.07 $Y=1.46 $X2=0 $Y2=0
cc_50 N_B_M1001_g Y 0.0206888f $X=0.895 $Y=2.465 $X2=0 $Y2=0
cc_51 N_B_M1001_g N_Y_c_98_n 0.0155419f $X=0.895 $Y=2.465 $X2=0 $Y2=0
cc_52 B N_Y_c_98_n 0.0242366f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_53 N_B_c_53_n N_Y_c_98_n 0.00135012f $X=1.07 $Y=1.46 $X2=0 $Y2=0
cc_54 N_B_c_51_n N_VGND_c_117_n 5.35643e-19 $X=0.935 $Y=1.295 $X2=0 $Y2=0
cc_55 N_B_c_51_n N_VGND_c_119_n 0.0139636f $X=0.935 $Y=1.295 $X2=0 $Y2=0
cc_56 B N_VGND_c_119_n 0.0269149f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_57 N_B_c_53_n N_VGND_c_119_n 0.00128577f $X=1.07 $Y=1.46 $X2=0 $Y2=0
cc_58 N_B_c_51_n N_VGND_c_120_n 0.00400407f $X=0.935 $Y=1.295 $X2=0 $Y2=0
cc_59 N_B_c_51_n N_VGND_c_121_n 0.00775088f $X=0.935 $Y=1.295 $X2=0 $Y2=0
cc_60 N_VPWR_c_75_n A_116_367# 0.00353023f $X=1.2 $Y=3.33 $X2=-0.19 $Y2=-0.245
cc_61 N_VPWR_c_75_n N_Y_M1001_d 0.00215158f $X=1.2 $Y=3.33 $X2=0 $Y2=0
cc_62 N_VPWR_c_78_n Y 0.0409085f $X=1.2 $Y=3.33 $X2=0 $Y2=0
cc_63 N_VPWR_c_75_n Y 0.0244227f $X=1.2 $Y=3.33 $X2=0 $Y2=0
cc_64 A_116_367# Y 0.00136968f $X=0.58 $Y=1.835 $X2=0.455 $Y2=3.33
cc_65 Y N_VGND_c_117_n 0.0275555f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_66 Y N_VGND_c_119_n 0.0275555f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_67 Y N_VGND_c_120_n 0.00932149f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_68 Y N_VGND_c_121_n 0.00704609f $X=0.635 $Y=0.47 $X2=0 $Y2=0
