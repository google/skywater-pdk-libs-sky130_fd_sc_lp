* File: sky130_fd_sc_lp__o21ai_1.pxi.spice
* Created: Wed Sep  2 10:15:58 2020
* 
x_PM_SKY130_FD_SC_LP__O21AI_1%A1 N_A1_M1003_g N_A1_M1002_g A1 A1 N_A1_c_41_n
+ PM_SKY130_FD_SC_LP__O21AI_1%A1
x_PM_SKY130_FD_SC_LP__O21AI_1%A2 N_A2_M1001_g N_A2_M1000_g A2 N_A2_c_65_n
+ N_A2_c_66_n PM_SKY130_FD_SC_LP__O21AI_1%A2
x_PM_SKY130_FD_SC_LP__O21AI_1%B1 N_B1_M1005_g N_B1_M1004_g B1 N_B1_c_99_n
+ N_B1_c_100_n PM_SKY130_FD_SC_LP__O21AI_1%B1
x_PM_SKY130_FD_SC_LP__O21AI_1%VPWR N_VPWR_M1002_s N_VPWR_M1004_d N_VPWR_c_121_n
+ N_VPWR_c_122_n N_VPWR_c_123_n N_VPWR_c_124_n VPWR N_VPWR_c_125_n
+ N_VPWR_c_120_n PM_SKY130_FD_SC_LP__O21AI_1%VPWR
x_PM_SKY130_FD_SC_LP__O21AI_1%Y N_Y_M1005_d N_Y_M1001_d N_Y_c_145_n N_Y_c_146_n
+ N_Y_c_147_n Y Y Y N_Y_c_148_n PM_SKY130_FD_SC_LP__O21AI_1%Y
x_PM_SKY130_FD_SC_LP__O21AI_1%A_29_47# N_A_29_47#_M1003_s N_A_29_47#_M1000_d
+ N_A_29_47#_c_171_n N_A_29_47#_c_172_n N_A_29_47#_c_175_n N_A_29_47#_c_177_n
+ PM_SKY130_FD_SC_LP__O21AI_1%A_29_47#
x_PM_SKY130_FD_SC_LP__O21AI_1%VGND N_VGND_M1003_d N_VGND_c_198_n VGND
+ N_VGND_c_199_n N_VGND_c_200_n N_VGND_c_201_n N_VGND_c_202_n
+ PM_SKY130_FD_SC_LP__O21AI_1%VGND
cc_1 VNB N_A1_M1003_g 0.0253206f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=0.655
cc_2 VNB N_A1_M1002_g 0.00692134f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=2.465
cc_3 VNB A1 0.0201848f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_4 VNB N_A1_c_41_n 0.0468897f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=1.375
cc_5 VNB N_A2_M1000_g 0.0267018f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=2.465
cc_6 VNB N_A2_c_65_n 0.0250035f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_A2_c_66_n 0.00397097f $X=-0.19 $Y=-0.245 $X2=0.295 $Y2=1.375
cc_8 VNB N_B1_M1005_g 0.0295549f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=0.655
cc_9 VNB N_B1_M1004_g 4.99662e-19 $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=2.465
cc_10 VNB N_B1_c_99_n 0.0494453f $X=-0.19 $Y=-0.245 $X2=0.295 $Y2=1.375
cc_11 VNB N_B1_c_100_n 0.013048f $X=-0.19 $Y=-0.245 $X2=0.295 $Y2=1.375
cc_12 VNB N_VPWR_c_120_n 0.0840719f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_Y_c_145_n 0.00951404f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_14 VNB N_Y_c_146_n 7.58946e-19 $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_15 VNB N_Y_c_147_n 0.0273454f $X=-0.19 $Y=-0.245 $X2=0.295 $Y2=1.375
cc_16 VNB N_Y_c_148_n 0.00896706f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_29_47#_c_171_n 0.0174052f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=2.465
cc_18 VNB N_A_29_47#_c_172_n 0.0142392f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_19 VNB N_VGND_c_198_n 0.00557173f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=2.465
cc_20 VNB N_VGND_c_199_n 0.0167643f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_21 VNB N_VGND_c_200_n 0.0282571f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=1.375
cc_22 VNB N_VGND_c_201_n 0.128948f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_VGND_c_202_n 0.0063111f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VPB N_A1_M1002_g 0.0246212f $X=-0.19 $Y=1.655 $X2=0.485 $Y2=2.465
cc_25 VPB A1 0.00733017f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_26 VPB N_A2_M1001_g 0.0193062f $X=-0.19 $Y=1.655 $X2=0.485 $Y2=0.655
cc_27 VPB N_A2_c_65_n 0.00628254f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_28 VPB N_A2_c_66_n 0.00965369f $X=-0.19 $Y=1.655 $X2=0.295 $Y2=1.375
cc_29 VPB N_B1_M1004_g 0.0272128f $X=-0.19 $Y=1.655 $X2=0.485 $Y2=2.465
cc_30 VPB N_B1_c_100_n 0.00716433f $X=-0.19 $Y=1.655 $X2=0.295 $Y2=1.375
cc_31 VPB N_VPWR_c_121_n 0.0106587f $X=-0.19 $Y=1.655 $X2=0.485 $Y2=2.465
cc_32 VPB N_VPWR_c_122_n 0.0484153f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_33 VPB N_VPWR_c_123_n 0.0108797f $X=-0.19 $Y=1.655 $X2=0.295 $Y2=1.375
cc_34 VPB N_VPWR_c_124_n 0.0503601f $X=-0.19 $Y=1.655 $X2=0.295 $Y2=1.375
cc_35 VPB N_VPWR_c_125_n 0.0298023f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_36 VPB N_VPWR_c_120_n 0.0437806f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_37 VPB N_Y_c_148_n 0.00378797f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_38 N_A1_M1002_g N_A2_M1001_g 0.0557605f $X=0.485 $Y=2.465 $X2=0 $Y2=0
cc_39 N_A1_M1003_g N_A2_M1000_g 0.0327537f $X=0.485 $Y=0.655 $X2=0 $Y2=0
cc_40 A1 N_A2_M1000_g 6.05496e-19 $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_41 A1 N_A2_c_65_n 2.88282e-19 $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_42 N_A1_c_41_n N_A2_c_65_n 0.0557605f $X=0.485 $Y=1.375 $X2=0 $Y2=0
cc_43 A1 N_A2_c_66_n 0.0327225f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_44 N_A1_c_41_n N_A2_c_66_n 0.00305778f $X=0.485 $Y=1.375 $X2=0 $Y2=0
cc_45 N_A1_M1002_g N_VPWR_c_122_n 0.0298791f $X=0.485 $Y=2.465 $X2=0 $Y2=0
cc_46 A1 N_VPWR_c_122_n 0.0252511f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_47 N_A1_c_41_n N_VPWR_c_122_n 0.00125434f $X=0.485 $Y=1.375 $X2=0 $Y2=0
cc_48 N_A1_M1002_g N_VPWR_c_125_n 0.00486043f $X=0.485 $Y=2.465 $X2=0 $Y2=0
cc_49 N_A1_M1002_g N_VPWR_c_120_n 0.00818711f $X=0.485 $Y=2.465 $X2=0 $Y2=0
cc_50 A1 N_A_29_47#_c_171_n 0.0223937f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_51 N_A1_c_41_n N_A_29_47#_c_171_n 0.00187244f $X=0.485 $Y=1.375 $X2=0 $Y2=0
cc_52 N_A1_M1003_g N_A_29_47#_c_175_n 0.0241841f $X=0.485 $Y=0.655 $X2=0 $Y2=0
cc_53 A1 N_A_29_47#_c_175_n 0.00170291f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_54 N_A1_M1003_g N_A_29_47#_c_177_n 5.71696e-19 $X=0.485 $Y=0.655 $X2=0 $Y2=0
cc_55 N_A1_M1003_g N_VGND_c_198_n 0.00336601f $X=0.485 $Y=0.655 $X2=0 $Y2=0
cc_56 N_A1_M1003_g N_VGND_c_199_n 0.00425094f $X=0.485 $Y=0.655 $X2=0 $Y2=0
cc_57 N_A1_M1003_g N_VGND_c_201_n 0.00680801f $X=0.485 $Y=0.655 $X2=0 $Y2=0
cc_58 N_A2_M1000_g N_B1_M1005_g 0.0237406f $X=1.015 $Y=0.655 $X2=0 $Y2=0
cc_59 N_A2_M1001_g N_B1_M1004_g 0.0284192f $X=0.845 $Y=2.465 $X2=0 $Y2=0
cc_60 N_A2_c_65_n N_B1_c_99_n 0.0139038f $X=0.935 $Y=1.51 $X2=0 $Y2=0
cc_61 N_A2_M1001_g N_VPWR_c_122_n 0.00445507f $X=0.845 $Y=2.465 $X2=0 $Y2=0
cc_62 N_A2_M1001_g N_VPWR_c_125_n 0.00585385f $X=0.845 $Y=2.465 $X2=0 $Y2=0
cc_63 N_A2_M1001_g N_VPWR_c_120_n 0.0112227f $X=0.845 $Y=2.465 $X2=0 $Y2=0
cc_64 N_A2_M1000_g N_Y_c_146_n 0.00353813f $X=1.015 $Y=0.655 $X2=0 $Y2=0
cc_65 N_A2_c_65_n Y 0.00395012f $X=0.935 $Y=1.51 $X2=0 $Y2=0
cc_66 N_A2_c_66_n Y 0.00533665f $X=0.935 $Y=1.51 $X2=0 $Y2=0
cc_67 N_A2_M1001_g N_Y_c_148_n 0.00357145f $X=0.845 $Y=2.465 $X2=0 $Y2=0
cc_68 N_A2_M1000_g N_Y_c_148_n 0.00448715f $X=1.015 $Y=0.655 $X2=0 $Y2=0
cc_69 N_A2_c_65_n N_Y_c_148_n 0.00236193f $X=0.935 $Y=1.51 $X2=0 $Y2=0
cc_70 N_A2_c_66_n N_Y_c_148_n 0.0314039f $X=0.935 $Y=1.51 $X2=0 $Y2=0
cc_71 N_A2_M1000_g N_A_29_47#_c_175_n 0.0204918f $X=1.015 $Y=0.655 $X2=0 $Y2=0
cc_72 N_A2_c_65_n N_A_29_47#_c_175_n 0.00388545f $X=0.935 $Y=1.51 $X2=0 $Y2=0
cc_73 N_A2_c_66_n N_A_29_47#_c_175_n 0.0204582f $X=0.935 $Y=1.51 $X2=0 $Y2=0
cc_74 N_A2_M1000_g N_A_29_47#_c_177_n 0.00568997f $X=1.015 $Y=0.655 $X2=0 $Y2=0
cc_75 N_A2_M1000_g N_VGND_c_198_n 0.00439036f $X=1.015 $Y=0.655 $X2=0 $Y2=0
cc_76 N_A2_M1000_g N_VGND_c_200_n 0.00415251f $X=1.015 $Y=0.655 $X2=0 $Y2=0
cc_77 N_A2_M1000_g N_VGND_c_201_n 0.00598651f $X=1.015 $Y=0.655 $X2=0 $Y2=0
cc_78 N_B1_M1004_g N_VPWR_c_124_n 0.00663507f $X=1.445 $Y=2.465 $X2=0 $Y2=0
cc_79 N_B1_c_99_n N_VPWR_c_124_n 0.00161206f $X=1.65 $Y=1.48 $X2=0 $Y2=0
cc_80 N_B1_c_100_n N_VPWR_c_124_n 0.0240385f $X=1.65 $Y=1.48 $X2=0 $Y2=0
cc_81 N_B1_M1004_g N_VPWR_c_125_n 0.00585385f $X=1.445 $Y=2.465 $X2=0 $Y2=0
cc_82 N_B1_M1004_g N_VPWR_c_120_n 0.0119726f $X=1.445 $Y=2.465 $X2=0 $Y2=0
cc_83 N_B1_M1005_g N_Y_c_145_n 0.0175628f $X=1.445 $Y=0.655 $X2=0 $Y2=0
cc_84 N_B1_c_99_n N_Y_c_145_n 0.00724399f $X=1.65 $Y=1.48 $X2=0 $Y2=0
cc_85 N_B1_c_100_n N_Y_c_145_n 0.0250843f $X=1.65 $Y=1.48 $X2=0 $Y2=0
cc_86 N_B1_M1005_g N_Y_c_148_n 0.0190519f $X=1.445 $Y=0.655 $X2=0 $Y2=0
cc_87 N_B1_c_100_n N_Y_c_148_n 0.0329163f $X=1.65 $Y=1.48 $X2=0 $Y2=0
cc_88 N_B1_M1005_g N_A_29_47#_c_175_n 0.00255208f $X=1.445 $Y=0.655 $X2=0 $Y2=0
cc_89 N_B1_M1005_g N_A_29_47#_c_177_n 0.00423437f $X=1.445 $Y=0.655 $X2=0 $Y2=0
cc_90 N_B1_M1005_g N_VGND_c_200_n 0.0054895f $X=1.445 $Y=0.655 $X2=0 $Y2=0
cc_91 N_B1_M1005_g N_VGND_c_201_n 0.0108708f $X=1.445 $Y=0.655 $X2=0 $Y2=0
cc_92 N_VPWR_c_120_n A_112_367# 0.00899413f $X=1.68 $Y=3.33 $X2=-0.19 $Y2=-0.245
cc_93 N_VPWR_c_120_n N_Y_M1001_d 0.00476222f $X=1.68 $Y=3.33 $X2=0 $Y2=0
cc_94 N_VPWR_c_125_n Y 0.0265345f $X=1.53 $Y=3.33 $X2=0 $Y2=0
cc_95 N_VPWR_c_120_n Y 0.0162509f $X=1.68 $Y=3.33 $X2=0 $Y2=0
cc_96 N_Y_c_146_n N_A_29_47#_M1000_d 0.00236306f $X=1.36 $Y=1.06 $X2=0 $Y2=0
cc_97 N_Y_c_145_n N_A_29_47#_c_175_n 0.00183148f $X=1.565 $Y=1.06 $X2=0 $Y2=0
cc_98 N_Y_c_146_n N_A_29_47#_c_175_n 0.0165697f $X=1.36 $Y=1.06 $X2=0 $Y2=0
cc_99 N_Y_c_147_n N_VGND_c_200_n 0.0178111f $X=1.66 $Y=0.42 $X2=0 $Y2=0
cc_100 N_Y_M1005_d N_VGND_c_201_n 0.00371702f $X=1.52 $Y=0.235 $X2=0 $Y2=0
cc_101 N_Y_c_147_n N_VGND_c_201_n 0.0100304f $X=1.66 $Y=0.42 $X2=0 $Y2=0
cc_102 N_A_29_47#_c_175_n N_VGND_M1003_d 0.00671177f $X=0.818 $Y=0.837 $X2=-0.19
+ $Y2=-0.245
cc_103 N_A_29_47#_c_175_n N_VGND_c_198_n 0.0214761f $X=0.818 $Y=0.837 $X2=0
+ $Y2=0
cc_104 N_A_29_47#_c_172_n N_VGND_c_199_n 0.0170745f $X=0.27 $Y=0.43 $X2=0 $Y2=0
cc_105 N_A_29_47#_c_175_n N_VGND_c_199_n 0.00297106f $X=0.818 $Y=0.837 $X2=0
+ $Y2=0
cc_106 N_A_29_47#_c_175_n N_VGND_c_200_n 0.00255347f $X=0.818 $Y=0.837 $X2=0
+ $Y2=0
cc_107 N_A_29_47#_c_177_n N_VGND_c_200_n 0.0186967f $X=1.23 $Y=0.36 $X2=0 $Y2=0
cc_108 N_A_29_47#_M1003_s N_VGND_c_201_n 0.00226765f $X=0.145 $Y=0.235 $X2=0
+ $Y2=0
cc_109 N_A_29_47#_M1000_d N_VGND_c_201_n 0.00223559f $X=1.09 $Y=0.235 $X2=0
+ $Y2=0
cc_110 N_A_29_47#_c_172_n N_VGND_c_201_n 0.0103698f $X=0.27 $Y=0.43 $X2=0 $Y2=0
cc_111 N_A_29_47#_c_175_n N_VGND_c_201_n 0.0107147f $X=0.818 $Y=0.837 $X2=0
+ $Y2=0
cc_112 N_A_29_47#_c_177_n N_VGND_c_201_n 0.0123168f $X=1.23 $Y=0.36 $X2=0 $Y2=0
