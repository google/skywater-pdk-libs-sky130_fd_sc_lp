* File: sky130_fd_sc_lp__or4b_2.pex.spice
* Created: Wed Sep  2 10:32:34 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__OR4B_2%D_N 3 7 9 13 15
c23 3 0 1.36172e-19 $X=0.495 $Y=0.865
r24 12 15 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=0.315 $Y=1.46
+ $X2=0.495 $Y2=1.46
r25 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.315
+ $Y=1.46 $X2=0.315 $Y2=1.46
r26 9 13 5.98103 $w=3.93e-07 $l=2.05e-07 $layer=LI1_cond $X=0.282 $Y=1.665
+ $X2=0.282 $Y2=1.46
r27 5 15 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=1.625
+ $X2=0.495 $Y2=1.46
r28 5 7 215.362 $w=1.5e-07 $l=4.2e-07 $layer=POLY_cond $X=0.495 $Y=1.625
+ $X2=0.495 $Y2=2.045
r29 1 15 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=1.295
+ $X2=0.495 $Y2=1.46
r30 1 3 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=0.495 $Y=1.295
+ $X2=0.495 $Y2=0.865
.ends

.subckt PM_SKY130_FD_SC_LP__OR4B_2%A_189_21# 1 2 3 12 16 20 24 29 30 31 32 33 36
+ 40 42 43 45 47 58
c130 58 0 1.66734e-19 $X=1.45 $Y=1.5
c131 45 0 6.20762e-20 $X=1.445 $Y=1.5
c132 43 0 6.34071e-20 $X=3.58 $Y=2.005
c133 33 0 2.92444e-20 $X=1.67 $Y=2.095
c134 31 0 3.08793e-20 $X=1.67 $Y=1.09
c135 29 0 2.36599e-20 $X=1.585 $Y=2.005
r136 46 58 0.874306 $w=3.3e-07 $l=5e-09 $layer=POLY_cond $X=1.445 $Y=1.5
+ $X2=1.45 $Y2=1.5
r137 46 55 74.316 $w=3.3e-07 $l=4.25e-07 $layer=POLY_cond $X=1.445 $Y=1.5
+ $X2=1.02 $Y2=1.5
r138 45 48 8.46025 $w=3.18e-07 $l=1.65e-07 $layer=LI1_cond $X=1.51 $Y=1.5
+ $X2=1.51 $Y2=1.665
r139 45 47 8.46025 $w=3.18e-07 $l=1.65e-07 $layer=LI1_cond $X=1.51 $Y=1.5
+ $X2=1.51 $Y2=1.335
r140 45 46 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.445
+ $Y=1.5 $X2=1.445 $Y2=1.5
r141 43 54 2.68691 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=3.58 $Y=2.005 $X2=3.58
+ $Y2=2.095
r142 42 43 38.764 $w=3.28e-07 $l=1.11e-06 $layer=LI1_cond $X=3.58 $Y=0.895
+ $X2=3.58 $Y2=2.005
r143 38 42 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=3.15 $Y=0.81
+ $X2=3.58 $Y2=0.81
r144 38 40 9.7783 $w=3.28e-07 $l=2.8e-07 $layer=LI1_cond $X=3.15 $Y=0.725
+ $X2=3.15 $Y2=0.445
r145 34 36 30.0171 $w=2.13e-07 $l=5.6e-07 $layer=LI1_cond $X=2.167 $Y=1.005
+ $X2=2.167 $Y2=0.445
r146 32 54 4.92601 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=3.415 $Y=2.095
+ $X2=3.58 $Y2=2.095
r147 32 33 107.52 $w=1.78e-07 $l=1.745e-06 $layer=LI1_cond $X=3.415 $Y=2.095
+ $X2=1.67 $Y2=2.095
r148 30 34 6.93832 $w=1.7e-07 $l=1.43332e-07 $layer=LI1_cond $X=2.06 $Y=1.09
+ $X2=2.167 $Y2=1.005
r149 30 31 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=2.06 $Y=1.09
+ $X2=1.67 $Y2=1.09
r150 29 33 6.82373 $w=1.8e-07 $l=1.25499e-07 $layer=LI1_cond $X=1.585 $Y=2.005
+ $X2=1.67 $Y2=2.095
r151 29 48 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=1.585 $Y=2.005
+ $X2=1.585 $Y2=1.665
r152 26 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.585 $Y=1.175
+ $X2=1.67 $Y2=1.09
r153 26 47 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=1.585 $Y=1.175
+ $X2=1.585 $Y2=1.335
r154 22 58 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.45 $Y=1.665
+ $X2=1.45 $Y2=1.5
r155 22 24 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=1.45 $Y=1.665
+ $X2=1.45 $Y2=2.465
r156 18 58 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.45 $Y=1.335
+ $X2=1.45 $Y2=1.5
r157 18 20 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=1.45 $Y=1.335
+ $X2=1.45 $Y2=0.655
r158 14 55 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.02 $Y=1.665
+ $X2=1.02 $Y2=1.5
r159 14 16 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=1.02 $Y=1.665
+ $X2=1.02 $Y2=2.465
r160 10 55 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.02 $Y=1.335
+ $X2=1.02 $Y2=1.5
r161 10 12 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=1.02 $Y=1.335
+ $X2=1.02 $Y2=0.655
r162 3 54 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=3.44
+ $Y=1.925 $X2=3.58 $Y2=2.07
r163 2 40 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=3.01
+ $Y=0.235 $X2=3.15 $Y2=0.445
r164 1 36 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.05
+ $Y=0.235 $X2=2.19 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__OR4B_2%A 3 7 9 12 13
r37 12 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.015 $Y=1.51
+ $X2=2.015 $Y2=1.675
r38 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.015 $Y=1.51
+ $X2=2.015 $Y2=1.345
r39 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.015
+ $Y=1.51 $X2=2.015 $Y2=1.51
r40 9 13 4.20303 $w=4.23e-07 $l=1.55e-07 $layer=LI1_cond $X=2.062 $Y=1.665
+ $X2=2.062 $Y2=1.51
r41 7 15 235.872 $w=1.5e-07 $l=4.6e-07 $layer=POLY_cond $X=2.105 $Y=2.135
+ $X2=2.105 $Y2=1.675
r42 3 14 461.489 $w=1.5e-07 $l=9e-07 $layer=POLY_cond $X=1.975 $Y=0.445
+ $X2=1.975 $Y2=1.345
.ends

.subckt PM_SKY130_FD_SC_LP__OR4B_2%B 3 5 7 9 10 11
r42 10 11 13.3251 $w=3.18e-07 $l=3.7e-07 $layer=LI1_cond $X=2.605 $Y=1.295
+ $X2=2.605 $Y2=1.665
r43 10 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.555
+ $Y=1.32 $X2=2.555 $Y2=1.32
r44 9 10 13.3251 $w=3.18e-07 $l=3.7e-07 $layer=LI1_cond $X=2.605 $Y=0.925
+ $X2=2.605 $Y2=1.295
r45 5 16 38.7444 $w=2.79e-07 $l=1.92678e-07 $layer=POLY_cond $X=2.465 $Y=1.485
+ $X2=2.525 $Y2=1.32
r46 5 7 333.298 $w=1.5e-07 $l=6.5e-07 $layer=POLY_cond $X=2.465 $Y=1.485
+ $X2=2.465 $Y2=2.135
r47 1 16 73.2963 $w=2.79e-07 $l=4.20743e-07 $layer=POLY_cond $X=2.405 $Y=0.955
+ $X2=2.525 $Y2=1.32
r48 1 3 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=2.405 $Y=0.955
+ $X2=2.405 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__OR4B_2%C 3 8 10 11 12 13 17 19
c43 11 0 6.34071e-20 $X=2.97 $Y=0.915
r44 17 20 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.095 $Y=1.29
+ $X2=3.095 $Y2=1.455
r45 17 19 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.095 $Y=1.29
+ $X2=3.095 $Y2=1.125
r46 12 13 13.9408 $w=3.08e-07 $l=3.75e-07 $layer=LI1_cond $X=3.09 $Y=1.29
+ $X2=3.09 $Y2=1.665
r47 12 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.095
+ $Y=1.29 $X2=3.095 $Y2=1.29
r48 11 19 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=3.005 $Y=0.915
+ $X2=3.005 $Y2=1.125
r49 10 11 43.7534 $w=2.2e-07 $l=1.5e-07 $layer=POLY_cond $X=2.97 $Y=0.765
+ $X2=2.97 $Y2=0.915
r50 8 20 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=3.005 $Y=2.135
+ $X2=3.005 $Y2=1.455
r51 3 10 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.935 $Y=0.445
+ $X2=2.935 $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_LP__OR4B_2%A_31_131# 1 2 7 9 13 15 18 22 24 28 31 32 36
+ 40 48
c80 48 0 6.68483e-20 $X=3.365 $Y=2.88
c81 32 0 1.66734e-19 $X=3.1 $Y=2.44
c82 31 0 2.36599e-20 $X=0.74 $Y=1.92
c83 28 0 3.08793e-20 $X=0.65 $Y=1.07
c84 24 0 2.92444e-20 $X=0.65 $Y=2.09
c85 18 0 1.48027e-19 $X=3.575 $Y=0.84
r86 40 42 7.15912 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=0.28 $Y=0.865
+ $X2=0.28 $Y2=1.07
r87 37 48 17.4861 $w=3.3e-07 $l=1e-07 $layer=POLY_cond $X=3.265 $Y=2.88
+ $X2=3.365 $Y2=2.88
r88 36 37 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.265
+ $Y=2.88 $X2=3.265 $Y2=2.88
r89 34 36 12.0329 $w=3.38e-07 $l=3.55e-07 $layer=LI1_cond $X=3.27 $Y=2.525
+ $X2=3.27 $Y2=2.88
r90 33 45 0.89264 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=0.83 $Y=2.44 $X2=0.74
+ $Y2=2.44
r91 32 34 7.85115 $w=1.7e-07 $l=2.08207e-07 $layer=LI1_cond $X=3.1 $Y=2.44
+ $X2=3.27 $Y2=2.525
r92 32 33 148.096 $w=1.68e-07 $l=2.27e-06 $layer=LI1_cond $X=3.1 $Y=2.44
+ $X2=0.83 $Y2=2.44
r93 30 31 47.1364 $w=1.78e-07 $l=7.65e-07 $layer=LI1_cond $X=0.74 $Y=1.155
+ $X2=0.74 $Y2=1.92
r94 29 42 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.445 $Y=1.07
+ $X2=0.28 $Y2=1.07
r95 28 30 6.82373 $w=1.7e-07 $l=1.25499e-07 $layer=LI1_cond $X=0.65 $Y=1.07
+ $X2=0.74 $Y2=1.155
r96 28 29 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=0.65 $Y=1.07
+ $X2=0.445 $Y2=1.07
r97 24 45 24.4 $w=1.75e-07 $l=3.5e-07 $layer=LI1_cond $X=0.74 $Y=2.09 $X2=0.74
+ $Y2=2.44
r98 24 31 11.5222 $w=1.8e-07 $l=1.7e-07 $layer=LI1_cond $X=0.74 $Y=2.09 $X2=0.74
+ $Y2=1.92
r99 24 26 12.5413 $w=3.38e-07 $l=3.7e-07 $layer=LI1_cond $X=0.65 $Y=2.09
+ $X2=0.28 $Y2=2.09
r100 20 22 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=3.365 $Y=1.74
+ $X2=3.575 $Y2=1.74
r101 16 18 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=3.365 $Y=0.84
+ $X2=3.575 $Y2=0.84
r102 15 22 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.575 $Y=1.665
+ $X2=3.575 $Y2=1.74
r103 14 18 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.575 $Y=0.915
+ $X2=3.575 $Y2=0.84
r104 14 15 384.574 $w=1.5e-07 $l=7.5e-07 $layer=POLY_cond $X=3.575 $Y=0.915
+ $X2=3.575 $Y2=1.665
r105 11 48 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.365 $Y=2.715
+ $X2=3.365 $Y2=2.88
r106 11 13 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=3.365 $Y=2.715
+ $X2=3.365 $Y2=2.135
r107 10 20 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.365 $Y=1.815
+ $X2=3.365 $Y2=1.74
r108 10 13 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=3.365 $Y=1.815
+ $X2=3.365 $Y2=2.135
r109 7 16 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.365 $Y=0.765
+ $X2=3.365 $Y2=0.84
r110 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=3.365 $Y=0.765
+ $X2=3.365 $Y2=0.445
r111 2 26 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=0.155
+ $Y=1.835 $X2=0.28 $Y2=2.045
r112 1 40 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.155
+ $Y=0.655 $X2=0.28 $Y2=0.865
.ends

.subckt PM_SKY130_FD_SC_LP__OR4B_2%VPWR 1 2 11 15 17 19 29 30 33 36
c32 30 0 6.68483e-20 $X=3.6 $Y=3.33
r33 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r34 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r35 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r36 27 30 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.6 $Y2=3.33
r37 26 29 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=2.16 $Y=3.33
+ $X2=3.6 $Y2=3.33
r38 26 27 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r39 24 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.83 $Y=3.33
+ $X2=1.665 $Y2=3.33
r40 24 26 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=1.83 $Y=3.33
+ $X2=2.16 $Y2=3.33
r41 23 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r42 23 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r43 22 23 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r44 20 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.97 $Y=3.33
+ $X2=0.805 $Y2=3.33
r45 20 22 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=0.97 $Y=3.33 $X2=1.2
+ $Y2=3.33
r46 19 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.5 $Y=3.33
+ $X2=1.665 $Y2=3.33
r47 19 22 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=1.5 $Y=3.33 $X2=1.2
+ $Y2=3.33
r48 17 27 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=2.16 $Y2=3.33
r49 17 37 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=1.68 $Y2=3.33
r50 13 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.665 $Y=3.245
+ $X2=1.665 $Y2=3.33
r51 13 15 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=1.665 $Y=3.245
+ $X2=1.665 $Y2=2.8
r52 9 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.805 $Y=3.245
+ $X2=0.805 $Y2=3.33
r53 9 11 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=0.805 $Y=3.245
+ $X2=0.805 $Y2=2.8
r54 2 15 600 $w=1.7e-07 $l=1.03263e-06 $layer=licon1_PDIFF $count=1 $X=1.525
+ $Y=1.835 $X2=1.665 $Y2=2.8
r55 1 11 600 $w=1.7e-07 $l=1.0761e-06 $layer=licon1_PDIFF $count=1 $X=0.57
+ $Y=1.835 $X2=0.805 $Y2=2.8
.ends

.subckt PM_SKY130_FD_SC_LP__OR4B_2%X 1 2 8 11 15 17
c29 15 0 1.36172e-19 $X=1.235 $Y=1.07
r30 17 19 3.55902 $w=3.38e-07 $l=1.05e-07 $layer=LI1_cond $X=1.2 $Y=2.015
+ $X2=1.095 $Y2=2.015
r31 13 15 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=1.095 $Y=1.07
+ $X2=1.235 $Y2=1.07
r32 9 15 0.0262452 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.235 $Y=0.985
+ $X2=1.235 $Y2=1.07
r33 9 11 32.9809 $w=1.88e-07 $l=5.65e-07 $layer=LI1_cond $X=1.235 $Y=0.985
+ $X2=1.235 $Y2=0.42
r34 8 19 4.80115 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=1.095 $Y=1.845
+ $X2=1.095 $Y2=2.015
r35 7 13 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.095 $Y=1.155
+ $X2=1.095 $Y2=1.07
r36 7 8 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.095 $Y=1.155
+ $X2=1.095 $Y2=1.845
r37 2 17 600 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_PDIFF $count=1 $X=1.095
+ $Y=1.835 $X2=1.235 $Y2=2.01
r38 1 11 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=1.095
+ $Y=0.235 $X2=1.235 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__OR4B_2%VGND 1 2 3 4 17 21 25 27 29 31 33 38 43 49 52
+ 55 59
c63 43 0 1.48027e-19 $X=3.485 $Y=0
r64 58 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r65 55 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r66 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r67 49 50 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r68 47 59 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r69 47 56 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.64
+ $Y2=0
r70 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r71 44 55 9.14399 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=2.815 $Y=0 $X2=2.635
+ $Y2=0
r72 44 46 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.815 $Y=0 $X2=3.12
+ $Y2=0
r73 43 58 4.13127 $w=1.7e-07 $l=1.77e-07 $layer=LI1_cond $X=3.485 $Y=0 $X2=3.662
+ $Y2=0
r74 43 46 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=3.485 $Y=0 $X2=3.12
+ $Y2=0
r75 42 56 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r76 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r77 39 52 9.6488 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=1.89 $Y=0 $X2=1.695
+ $Y2=0
r78 39 41 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=1.89 $Y=0 $X2=2.16
+ $Y2=0
r79 38 55 9.14399 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=2.455 $Y=0 $X2=2.635
+ $Y2=0
r80 38 41 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=2.455 $Y=0 $X2=2.16
+ $Y2=0
r81 37 53 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r82 37 50 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r83 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r84 34 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.97 $Y=0 $X2=0.805
+ $Y2=0
r85 34 36 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=0.97 $Y=0 $X2=1.2
+ $Y2=0
r86 33 52 9.6488 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=1.5 $Y=0 $X2=1.695
+ $Y2=0
r87 33 36 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=1.5 $Y=0 $X2=1.2 $Y2=0
r88 31 42 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=2.16
+ $Y2=0
r89 31 53 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=1.68
+ $Y2=0
r90 27 58 3.08095 $w=2.6e-07 $l=1.05924e-07 $layer=LI1_cond $X=3.615 $Y=0.085
+ $X2=3.662 $Y2=0
r91 27 29 13.519 $w=2.58e-07 $l=3.05e-07 $layer=LI1_cond $X=3.615 $Y=0.085
+ $X2=3.615 $Y2=0.39
r92 23 55 1.16013 $w=3.6e-07 $l=8.5e-08 $layer=LI1_cond $X=2.635 $Y=0.085
+ $X2=2.635 $Y2=0
r93 23 25 11.5244 $w=3.58e-07 $l=3.6e-07 $layer=LI1_cond $X=2.635 $Y=0.085
+ $X2=2.635 $Y2=0.445
r94 19 52 1.39532 $w=3.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.695 $Y=0.085
+ $X2=1.695 $Y2=0
r95 19 21 8.7172 $w=3.88e-07 $l=2.95e-07 $layer=LI1_cond $X=1.695 $Y=0.085
+ $X2=1.695 $Y2=0.38
r96 15 49 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.805 $Y=0.085
+ $X2=0.805 $Y2=0
r97 15 17 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.805 $Y=0.085
+ $X2=0.805 $Y2=0.38
r98 4 29 182 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=1 $X=3.44
+ $Y=0.235 $X2=3.58 $Y2=0.39
r99 3 25 182 $w=1.7e-07 $l=2.82489e-07 $layer=licon1_NDIFF $count=1 $X=2.48
+ $Y=0.235 $X2=2.65 $Y2=0.445
r100 2 21 91 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_NDIFF $count=2 $X=1.525
+ $Y=0.235 $X2=1.76 $Y2=0.38
r101 1 17 91 $w=1.7e-07 $l=3.745e-07 $layer=licon1_NDIFF $count=2 $X=0.57
+ $Y=0.655 $X2=0.805 $Y2=0.38
.ends

