* File: sky130_fd_sc_lp__or4_2.pex.spice
* Created: Wed Sep  2 10:31:56 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__OR4_2%D 1 2 3 4 7 11 15 16 17 22
r36 16 17 15.2287 $w=2.78e-07 $l=3.7e-07 $layer=LI1_cond $X=0.225 $Y=1.295
+ $X2=0.225 $Y2=1.665
r37 15 16 15.2287 $w=2.78e-07 $l=3.7e-07 $layer=LI1_cond $X=0.225 $Y=0.925
+ $X2=0.225 $Y2=1.295
r38 15 22 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.27
+ $Y=1.005 $X2=0.27 $Y2=1.005
r39 14 22 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=0.27 $Y=1.36
+ $X2=0.27 $Y2=1.005
r40 13 22 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=0.27 $Y=0.99
+ $X2=0.27 $Y2=1.005
r41 9 11 274.33 $w=1.5e-07 $l=5.35e-07 $layer=POLY_cond $X=0.7 $Y=1.51 $X2=0.7
+ $Y2=2.045
r42 5 7 197.415 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=0.7 $Y=0.84 $X2=0.7
+ $Y2=0.455
r43 4 14 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=0.435 $Y=1.435
+ $X2=0.27 $Y2=1.36
r44 3 9 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.625 $Y=1.435
+ $X2=0.7 $Y2=1.51
r45 3 4 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=0.625 $Y=1.435
+ $X2=0.435 $Y2=1.435
r46 2 13 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=0.435 $Y=0.915
+ $X2=0.27 $Y2=0.99
r47 1 5 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.625 $Y=0.915
+ $X2=0.7 $Y2=0.84
r48 1 2 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=0.625 $Y=0.915
+ $X2=0.435 $Y2=0.915
.ends

.subckt PM_SKY130_FD_SC_LP__OR4_2%C 3 7 11 12 13 14 15 16 17 24 25
r43 24 25 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.15
+ $Y=1.17 $X2=1.15 $Y2=1.17
r44 16 17 11.6823 $w=3.63e-07 $l=3.7e-07 $layer=LI1_cond $X=1.167 $Y=2.405
+ $X2=1.167 $Y2=2.775
r45 15 16 11.6823 $w=3.63e-07 $l=3.7e-07 $layer=LI1_cond $X=1.167 $Y=2.035
+ $X2=1.167 $Y2=2.405
r46 14 15 11.6823 $w=3.63e-07 $l=3.7e-07 $layer=LI1_cond $X=1.167 $Y=1.665
+ $X2=1.167 $Y2=2.035
r47 13 14 11.6823 $w=3.63e-07 $l=3.7e-07 $layer=LI1_cond $X=1.167 $Y=1.295
+ $X2=1.167 $Y2=1.665
r48 13 25 3.94672 $w=3.63e-07 $l=1.25e-07 $layer=LI1_cond $X=1.167 $Y=1.295
+ $X2=1.167 $Y2=1.17
r49 11 24 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.15 $Y=1.51
+ $X2=1.15 $Y2=1.17
r50 11 12 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.15 $Y=1.51
+ $X2=1.15 $Y2=1.675
r51 10 24 38.6168 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.15 $Y=1.005
+ $X2=1.15 $Y2=1.17
r52 7 10 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=1.13 $Y=0.455
+ $X2=1.13 $Y2=1.005
r53 3 12 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=1.06 $Y=2.045
+ $X2=1.06 $Y2=1.675
.ends

.subckt PM_SKY130_FD_SC_LP__OR4_2%B 3 7 11 12 13 14 15 16 17 24 25
c46 24 0 5.50976e-20 $X=1.69 $Y=1.17
r47 24 25 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.69
+ $Y=1.17 $X2=1.69 $Y2=1.17
r48 16 17 13.5366 $w=3.13e-07 $l=3.7e-07 $layer=LI1_cond $X=1.677 $Y=2.405
+ $X2=1.677 $Y2=2.775
r49 15 16 13.5366 $w=3.13e-07 $l=3.7e-07 $layer=LI1_cond $X=1.677 $Y=2.035
+ $X2=1.677 $Y2=2.405
r50 14 15 13.5366 $w=3.13e-07 $l=3.7e-07 $layer=LI1_cond $X=1.677 $Y=1.665
+ $X2=1.677 $Y2=2.035
r51 13 14 13.5366 $w=3.13e-07 $l=3.7e-07 $layer=LI1_cond $X=1.677 $Y=1.295
+ $X2=1.677 $Y2=1.665
r52 13 25 4.57319 $w=3.13e-07 $l=1.25e-07 $layer=LI1_cond $X=1.677 $Y=1.295
+ $X2=1.677 $Y2=1.17
r53 11 24 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.69 $Y=1.51
+ $X2=1.69 $Y2=1.17
r54 11 12 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.69 $Y=1.51
+ $X2=1.69 $Y2=1.675
r55 10 24 38.6168 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.69 $Y=1.005
+ $X2=1.69 $Y2=1.17
r56 7 10 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=1.71 $Y=0.455
+ $X2=1.71 $Y2=1.005
r57 3 12 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=1.6 $Y=2.045 $X2=1.6
+ $Y2=1.675
.ends

.subckt PM_SKY130_FD_SC_LP__OR4_2%A 3 7 9 10 11 12 20 21 41
r50 41 42 3.12273 $w=3.48e-07 $l=6e-08 $layer=LI1_cond $X=2.18 $Y=2.405 $X2=2.18
+ $Y2=2.345
r51 24 34 2.424 $w=2.4e-07 $l=1.6e-07 $layer=LI1_cond $X=2.125 $Y=1.675
+ $X2=2.125 $Y2=1.515
r52 20 23 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.23 $Y=1.51
+ $X2=2.23 $Y2=1.675
r53 20 22 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.23 $Y=1.51
+ $X2=2.23 $Y2=1.345
r54 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.23
+ $Y=1.51 $X2=2.23 $Y2=1.51
r55 12 30 8.39637 $w=3.48e-07 $l=2.55e-07 $layer=LI1_cond $X=2.18 $Y=2.775
+ $X2=2.18 $Y2=2.52
r56 11 30 3.39148 $w=3.48e-07 $l=1.03e-07 $layer=LI1_cond $X=2.18 $Y=2.417
+ $X2=2.18 $Y2=2.52
r57 11 41 0.395123 $w=3.48e-07 $l=1.2e-08 $layer=LI1_cond $X=2.18 $Y=2.417
+ $X2=2.18 $Y2=2.405
r58 11 42 0.62424 $w=2.38e-07 $l=1.3e-08 $layer=LI1_cond $X=2.125 $Y=2.332
+ $X2=2.125 $Y2=2.345
r59 10 11 14.2615 $w=2.38e-07 $l=2.97e-07 $layer=LI1_cond $X=2.125 $Y=2.035
+ $X2=2.125 $Y2=2.332
r60 9 21 2.52097 $w=3.18e-07 $l=7e-08 $layer=LI1_cond $X=2.16 $Y=1.515 $X2=2.23
+ $Y2=1.515
r61 9 34 1.26048 $w=3.18e-07 $l=3.5e-08 $layer=LI1_cond $X=2.16 $Y=1.515
+ $X2=2.125 $Y2=1.515
r62 9 10 15.51 $w=2.38e-07 $l=3.23e-07 $layer=LI1_cond $X=2.125 $Y=1.712
+ $X2=2.125 $Y2=2.035
r63 9 24 1.77668 $w=2.38e-07 $l=3.7e-08 $layer=LI1_cond $X=2.125 $Y=1.712
+ $X2=2.125 $Y2=1.675
r64 7 23 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=2.14 $Y=2.045
+ $X2=2.14 $Y2=1.675
r65 3 22 456.362 $w=1.5e-07 $l=8.9e-07 $layer=POLY_cond $X=2.14 $Y=0.455
+ $X2=2.14 $Y2=1.345
.ends

.subckt PM_SKY130_FD_SC_LP__OR4_2%A_72_367# 1 2 3 10 12 16 18 22 26 28 30 33 35
+ 36 39 41 42 43 44 48 55
c126 42 0 5.50976e-20 $X=2.145 $Y=1.015
r127 58 59 11.5066 $w=3.77e-07 $l=9e-08 $layer=POLY_cond $X=2.795 $Y=1.45
+ $X2=2.795 $Y2=1.36
r128 57 58 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.77
+ $Y=1.45 $X2=2.77 $Y2=1.45
r129 55 57 18.5652 $w=2.3e-07 $l=3.5e-07 $layer=LI1_cond $X=2.715 $Y=1.1
+ $X2=2.715 $Y2=1.45
r130 46 48 5.36482 $w=2.88e-07 $l=1.35e-07 $layer=LI1_cond $X=0.485 $Y=2.065
+ $X2=0.62 $Y2=2.065
r131 43 55 2.50919 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=2.575 $Y=1.1
+ $X2=2.715 $Y2=1.1
r132 43 44 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=2.575 $Y=1.1
+ $X2=2.285 $Y2=1.1
r133 42 44 7.36005 $w=1.7e-07 $l=1.77482e-07 $layer=LI1_cond $X=2.145 $Y=1.015
+ $X2=2.285 $Y2=1.1
r134 41 42 7.82015 $w=2.78e-07 $l=1.9e-07 $layer=LI1_cond $X=2.145 $Y=0.825
+ $X2=2.145 $Y2=1.015
r135 37 41 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=1.89 $Y=0.74
+ $X2=2.145 $Y2=0.74
r136 37 39 10.4163 $w=2.58e-07 $l=2.35e-07 $layer=LI1_cond $X=1.89 $Y=0.655
+ $X2=1.89 $Y2=0.42
r137 35 37 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=1.76 $Y=0.74
+ $X2=1.89 $Y2=0.74
r138 35 36 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.76 $Y=0.74
+ $X2=1.09 $Y2=0.74
r139 31 36 9.30461 $w=1.95e-07 $l=1.63783e-07 $layer=LI1_cond $X=0.945 $Y=0.78
+ $X2=1.09 $Y2=0.74
r140 31 50 20.3333 $w=1.95e-07 $l=3.25e-07 $layer=LI1_cond $X=0.945 $Y=0.78
+ $X2=0.62 $Y2=0.78
r141 31 33 9.33876 $w=2.88e-07 $l=2.35e-07 $layer=LI1_cond $X=0.945 $Y=0.655
+ $X2=0.945 $Y2=0.42
r142 30 48 3.86198 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=0.62 $Y=1.92
+ $X2=0.62 $Y2=2.065
r143 29 50 1.54022 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.62 $Y=0.905
+ $X2=0.62 $Y2=0.78
r144 29 30 66.2193 $w=1.68e-07 $l=1.015e-06 $layer=LI1_cond $X=0.62 $Y=0.905
+ $X2=0.62 $Y2=1.92
r145 24 28 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.34 $Y=1.435
+ $X2=3.34 $Y2=1.36
r146 24 26 528.149 $w=1.5e-07 $l=1.03e-06 $layer=POLY_cond $X=3.34 $Y=1.435
+ $X2=3.34 $Y2=2.465
r147 20 28 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.34 $Y=1.285
+ $X2=3.34 $Y2=1.36
r148 20 22 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=3.34 $Y=1.285
+ $X2=3.34 $Y2=0.665
r149 19 59 24.4204 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=2.985 $Y=1.36
+ $X2=2.795 $Y2=1.36
r150 18 28 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.265 $Y=1.36
+ $X2=3.34 $Y2=1.36
r151 18 19 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=3.265 $Y=1.36
+ $X2=2.985 $Y2=1.36
r152 14 59 27.6612 $w=3.77e-07 $l=1.47817e-07 $layer=POLY_cond $X=2.91 $Y=1.285
+ $X2=2.795 $Y2=1.36
r153 14 16 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=2.91 $Y=1.285
+ $X2=2.91 $Y2=0.665
r154 10 58 39.1678 $w=3.77e-07 $l=2.13014e-07 $layer=POLY_cond $X=2.905 $Y=1.615
+ $X2=2.795 $Y2=1.45
r155 10 12 435.851 $w=1.5e-07 $l=8.5e-07 $layer=POLY_cond $X=2.905 $Y=1.615
+ $X2=2.905 $Y2=2.465
r156 3 46 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=0.36
+ $Y=1.835 $X2=0.485 $Y2=2.045
r157 2 39 182 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=1 $X=1.785
+ $Y=0.245 $X2=1.925 $Y2=0.42
r158 1 33 182 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=1 $X=0.775
+ $Y=0.245 $X2=0.915 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__OR4_2%VPWR 1 2 10 11 13 18 21 23 31 37 41
r33 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r34 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r35 35 41 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r36 35 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.64 $Y2=3.33
r37 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r38 32 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.855 $Y=3.33
+ $X2=2.69 $Y2=3.33
r39 32 34 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=2.855 $Y=3.33
+ $X2=3.12 $Y2=3.33
r40 31 40 4.35645 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=3.43 $Y=3.33
+ $X2=3.635 $Y2=3.33
r41 31 34 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=3.43 $Y=3.33
+ $X2=3.12 $Y2=3.33
r42 30 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r43 29 30 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r44 25 29 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=0.24 $Y=3.33
+ $X2=2.16 $Y2=3.33
r45 25 26 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r46 23 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.525 $Y=3.33
+ $X2=2.69 $Y2=3.33
r47 23 29 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=2.525 $Y=3.33
+ $X2=2.16 $Y2=3.33
r48 21 30 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=2.16 $Y2=3.33
r49 21 26 0.468274 $w=4.9e-07 $l=1.68e-06 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=0.24 $Y2=3.33
r50 18 20 5.06779 $w=4.38e-07 $l=1.65e-07 $layer=LI1_cond $X=2.635 $Y=2.01
+ $X2=2.635 $Y2=2.175
r51 13 16 38.5472 $w=2.88e-07 $l=9.7e-07 $layer=LI1_cond $X=3.575 $Y=1.98
+ $X2=3.575 $Y2=2.95
r52 11 40 3.08139 $w=2.9e-07 $l=1.11018e-07 $layer=LI1_cond $X=3.575 $Y=3.245
+ $X2=3.635 $Y2=3.33
r53 11 16 11.7231 $w=2.88e-07 $l=2.95e-07 $layer=LI1_cond $X=3.575 $Y=3.245
+ $X2=3.575 $Y2=2.95
r54 10 20 9.7783 $w=3.28e-07 $l=2.8e-07 $layer=LI1_cond $X=2.69 $Y=2.455
+ $X2=2.69 $Y2=2.175
r55 8 37 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.69 $Y=3.245 $X2=2.69
+ $Y2=3.33
r56 8 10 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=2.69 $Y=3.245
+ $X2=2.69 $Y2=2.455
r57 2 16 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=3.415
+ $Y=1.835 $X2=3.555 $Y2=2.95
r58 2 13 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=3.415
+ $Y=1.835 $X2=3.555 $Y2=1.98
r59 1 18 600 $w=1.7e-07 $l=3.62077e-07 $layer=licon1_PDIFF $count=1 $X=2.215
+ $Y=1.835 $X2=2.5 $Y2=2.01
r60 1 10 300 $w=1.7e-07 $l=8.23954e-07 $layer=licon1_PDIFF $count=2 $X=2.215
+ $Y=1.835 $X2=2.69 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_LP__OR4_2%X 1 2 7 8 9 10 11 12 13 24 32
r22 30 32 3.57993 $w=2.33e-07 $l=7.3e-08 $layer=LI1_cond $X=3.142 $Y=1.222
+ $X2=3.142 $Y2=1.295
r23 13 44 6.62042 $w=2.33e-07 $l=1.35e-07 $layer=LI1_cond $X=3.142 $Y=2.775
+ $X2=3.142 $Y2=2.91
r24 12 13 18.1448 $w=2.33e-07 $l=3.7e-07 $layer=LI1_cond $X=3.142 $Y=2.405
+ $X2=3.142 $Y2=2.775
r25 11 12 20.8421 $w=2.33e-07 $l=4.25e-07 $layer=LI1_cond $X=3.142 $Y=1.98
+ $X2=3.142 $Y2=2.405
r26 10 11 15.4476 $w=2.33e-07 $l=3.15e-07 $layer=LI1_cond $X=3.142 $Y=1.665
+ $X2=3.142 $Y2=1.98
r27 9 30 0.294241 $w=2.33e-07 $l=6e-09 $layer=LI1_cond $X=3.142 $Y=1.216
+ $X2=3.142 $Y2=1.222
r28 9 47 5.44345 $w=2.33e-07 $l=1.11e-07 $layer=LI1_cond $X=3.142 $Y=1.216
+ $X2=3.142 $Y2=1.105
r29 9 10 17.8506 $w=2.33e-07 $l=3.64e-07 $layer=LI1_cond $X=3.142 $Y=1.301
+ $X2=3.142 $Y2=1.665
r30 9 32 0.294241 $w=2.33e-07 $l=6e-09 $layer=LI1_cond $X=3.142 $Y=1.301
+ $X2=3.142 $Y2=1.295
r31 8 47 9.01912 $w=2.28e-07 $l=1.8e-07 $layer=LI1_cond $X=3.145 $Y=0.925
+ $X2=3.145 $Y2=1.105
r32 7 8 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=3.145 $Y=0.555
+ $X2=3.145 $Y2=0.925
r33 7 24 6.76434 $w=2.28e-07 $l=1.35e-07 $layer=LI1_cond $X=3.145 $Y=0.555
+ $X2=3.145 $Y2=0.42
r34 2 44 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=2.98
+ $Y=1.835 $X2=3.12 $Y2=2.91
r35 2 11 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.98
+ $Y=1.835 $X2=3.12 $Y2=1.98
r36 1 24 91 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=2 $X=2.985
+ $Y=0.245 $X2=3.125 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__OR4_2%VGND 1 2 3 4 15 19 21 23 26 27 29 30 31 39 43
+ 49 55
r65 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r66 49 52 8.39153 $w=5.67e-07 $l=3.9e-07 $layer=LI1_cond $X=2.525 $Y=0 $X2=2.525
+ $Y2=0.39
r67 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r68 47 55 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r69 47 50 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.64
+ $Y2=0
r70 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r71 44 49 7.95352 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=2.86 $Y=0 $X2=2.525
+ $Y2=0
r72 44 46 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=2.86 $Y=0 $X2=3.12
+ $Y2=0
r73 43 54 4.35645 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=3.43 $Y=0 $X2=3.635
+ $Y2=0
r74 43 46 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=3.43 $Y=0 $X2=3.12
+ $Y2=0
r75 42 50 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r76 41 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r77 39 49 7.95352 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=2.19 $Y=0 $X2=2.525
+ $Y2=0
r78 39 41 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=2.19 $Y=0 $X2=2.16
+ $Y2=0
r79 37 38 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r80 35 38 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r81 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r82 31 42 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=2.16
+ $Y2=0
r83 31 38 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=1.2
+ $Y2=0
r84 29 37 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=1.26 $Y=0 $X2=1.2
+ $Y2=0
r85 29 30 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.26 $Y=0 $X2=1.425
+ $Y2=0
r86 28 41 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=1.59 $Y=0 $X2=2.16
+ $Y2=0
r87 28 30 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.59 $Y=0 $X2=1.425
+ $Y2=0
r88 26 34 4.30588 $w=1.7e-07 $l=6e-08 $layer=LI1_cond $X=0.3 $Y=0 $X2=0.24 $Y2=0
r89 26 27 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.3 $Y=0 $X2=0.465
+ $Y2=0
r90 25 37 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=0.63 $Y=0 $X2=1.2
+ $Y2=0
r91 25 27 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.63 $Y=0 $X2=0.465
+ $Y2=0
r92 21 54 3.08139 $w=2.9e-07 $l=1.11018e-07 $layer=LI1_cond $X=3.575 $Y=0.085
+ $X2=3.635 $Y2=0
r93 21 23 12.1205 $w=2.88e-07 $l=3.05e-07 $layer=LI1_cond $X=3.575 $Y=0.085
+ $X2=3.575 $Y2=0.39
r94 17 30 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.425 $Y=0.085
+ $X2=1.425 $Y2=0
r95 17 19 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=1.425 $Y=0.085
+ $X2=1.425 $Y2=0.37
r96 13 27 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.465 $Y=0.085
+ $X2=0.465 $Y2=0
r97 13 15 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=0.465 $Y=0.085
+ $X2=0.465 $Y2=0.44
r98 4 23 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.415
+ $Y=0.245 $X2=3.555 $Y2=0.39
r99 3 52 60.6667 $w=1.7e-07 $l=5.47723e-07 $layer=licon1_NDIFF $count=3 $X=2.215
+ $Y=0.245 $X2=2.695 $Y2=0.39
r100 2 19 182 $w=1.7e-07 $l=2.755e-07 $layer=licon1_NDIFF $count=1 $X=1.205
+ $Y=0.245 $X2=1.425 $Y2=0.37
r101 1 15 182 $w=1.7e-07 $l=2.498e-07 $layer=licon1_NDIFF $count=1 $X=0.34
+ $Y=0.245 $X2=0.465 $Y2=0.44
.ends

