* File: sky130_fd_sc_lp__ha_2.pex.spice
* Created: Wed Sep  2 09:54:30 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__HA_2%A_270_95# 1 2 7 9 10 12 16 19 21 23 25 28 32 35
+ 39 41 43 48 53 54
c111 41 0 7.01745e-20 $X=2.695 $Y=1.35
c112 28 0 2.76446e-20 $X=3.76 $Y=2.465
r113 53 54 31.8081 $w=3.75e-07 $l=7.5e-08 $layer=POLY_cond $X=3.217 $Y=1.26
+ $X2=3.217 $Y2=1.185
r114 49 50 15.5114 $w=3.5e-07 $l=4.45e-07 $layer=LI1_cond $X=2.155 $Y=1.332
+ $X2=2.6 $Y2=1.332
r115 47 49 7.66857 $w=3.5e-07 $l=2.2e-07 $layer=LI1_cond $X=1.935 $Y=1.332
+ $X2=2.155 $Y2=1.332
r116 47 48 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.935
+ $Y=1.35 $X2=1.935 $Y2=1.35
r117 44 56 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=3.217 $Y=1.35
+ $X2=3.217 $Y2=1.515
r118 44 53 13.3477 $w=3.75e-07 $l=9e-08 $layer=POLY_cond $X=3.217 $Y=1.35
+ $X2=3.217 $Y2=1.26
r119 43 44 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.195
+ $Y=1.35 $X2=3.195 $Y2=1.35
r120 41 50 3.36558 $w=3.5e-07 $l=1.0361e-07 $layer=LI1_cond $X=2.695 $Y=1.35
+ $X2=2.6 $Y2=1.332
r121 41 43 17.4613 $w=3.28e-07 $l=5e-07 $layer=LI1_cond $X=2.695 $Y=1.35
+ $X2=3.195 $Y2=1.35
r122 37 50 4.31381 $w=1.9e-07 $l=1.83e-07 $layer=LI1_cond $X=2.6 $Y=1.515
+ $X2=2.6 $Y2=1.332
r123 37 39 36.4833 $w=1.88e-07 $l=6.25e-07 $layer=LI1_cond $X=2.6 $Y=1.515
+ $X2=2.6 $Y2=2.14
r124 33 49 0.543965 $w=3.6e-07 $l=1.82e-07 $layer=LI1_cond $X=2.155 $Y=1.15
+ $X2=2.155 $Y2=1.332
r125 33 35 9.12351 $w=3.58e-07 $l=2.85e-07 $layer=LI1_cond $X=2.155 $Y=1.15
+ $X2=2.155 $Y2=0.865
r126 31 48 44.5896 $w=3.3e-07 $l=2.55e-07 $layer=POLY_cond $X=1.68 $Y=1.35
+ $X2=1.935 $Y2=1.35
r127 26 32 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.76 $Y=1.335
+ $X2=3.76 $Y2=1.26
r128 26 28 579.426 $w=1.5e-07 $l=1.13e-06 $layer=POLY_cond $X=3.76 $Y=1.335
+ $X2=3.76 $Y2=2.465
r129 23 32 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.76 $Y=1.185
+ $X2=3.76 $Y2=1.26
r130 23 25 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=3.76 $Y=1.185
+ $X2=3.76 $Y2=0.655
r131 22 53 24.2915 $w=1.5e-07 $l=1.88e-07 $layer=POLY_cond $X=3.405 $Y=1.26
+ $X2=3.217 $Y2=1.26
r132 21 32 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.685 $Y=1.26
+ $X2=3.76 $Y2=1.26
r133 21 22 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=3.685 $Y=1.26
+ $X2=3.405 $Y2=1.26
r134 19 56 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=3.33 $Y=2.465
+ $X2=3.33 $Y2=1.515
r135 16 54 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=3.33 $Y=0.655
+ $X2=3.33 $Y2=1.185
r136 10 31 40.7811 $w=2.24e-07 $l=1.98997e-07 $layer=POLY_cond $X=1.6 $Y=1.515
+ $X2=1.525 $Y2=1.35
r137 10 12 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.6 $Y=1.515
+ $X2=1.6 $Y2=2.305
r138 7 31 51.5401 $w=2.24e-07 $l=2.6024e-07 $layer=POLY_cond $X=1.425 $Y=1.135
+ $X2=1.525 $Y2=1.35
r139 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.425 $Y=1.135
+ $X2=1.425 $Y2=0.815
r140 2 39 600 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_PDIFF $count=1 $X=2.45
+ $Y=1.985 $X2=2.59 $Y2=2.14
r141 1 35 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=2.045
+ $Y=0.655 $X2=2.17 $Y2=0.865
.ends

.subckt PM_SKY130_FD_SC_LP__HA_2%B 4 9 11 12 15 19 21 23 24 27 29
c76 23 0 7.01745e-20 $X=2.38 $Y=1.875
c77 4 0 1.61446e-19 $X=0.995 $Y=0.815
r78 27 30 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.15 $Y=1.66
+ $X2=1.15 $Y2=1.825
r79 27 29 45.1865 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.15 $Y=1.66
+ $X2=1.15 $Y2=1.495
r80 24 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.15
+ $Y=1.66 $X2=1.15 $Y2=1.66
r81 22 23 69.5192 $w=1.6e-07 $l=1.5e-07 $layer=POLY_cond $X=2.38 $Y=1.725
+ $X2=2.38 $Y2=1.875
r82 21 29 100.466 $w=1.55e-07 $l=2.1e-07 $layer=POLY_cond $X=1.062 $Y=1.285
+ $X2=1.062 $Y2=1.495
r83 20 21 71.7618 $w=1.55e-07 $l=1.5e-07 $layer=POLY_cond $X=1.03 $Y=1.135
+ $X2=1.03 $Y2=1.285
r84 19 22 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=2.385 $Y=0.865
+ $X2=2.385 $Y2=1.725
r85 16 19 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=2.385 $Y=0.265
+ $X2=2.385 $Y2=0.865
r86 15 23 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=2.375 $Y=2.305
+ $X2=2.375 $Y2=1.875
r87 11 16 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.31 $Y=0.19
+ $X2=2.385 $Y2=0.265
r88 11 12 635.83 $w=1.5e-07 $l=1.24e-06 $layer=POLY_cond $X=2.31 $Y=0.19
+ $X2=1.07 $Y2=0.19
r89 9 30 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.06 $Y=2.305
+ $X2=1.06 $Y2=1.825
r90 4 20 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.995 $Y=0.815
+ $X2=0.995 $Y2=1.135
r91 1 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.995 $Y=0.265
+ $X2=1.07 $Y2=0.19
r92 1 4 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=0.995 $Y=0.265
+ $X2=0.995 $Y2=0.815
.ends

.subckt PM_SKY130_FD_SC_LP__HA_2%A 3 8 9 10 13 18 20 21 22 28
c67 20 0 6.34558e-20 $X=2.775 $Y=1.875
c68 13 0 3.48876e-19 $X=2.745 $Y=0.865
r69 26 28 8.3391 $w=2.89e-07 $l=5e-08 $layer=POLY_cond $X=0.515 $Y=1.66
+ $X2=0.565 $Y2=1.66
r70 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.515
+ $Y=1.66 $X2=0.515 $Y2=1.66
r71 22 27 7.62099 $w=3.08e-07 $l=2.05e-07 $layer=LI1_cond $X=0.72 $Y=1.65
+ $X2=0.515 $Y2=1.65
r72 21 27 10.2233 $w=3.08e-07 $l=2.75e-07 $layer=LI1_cond $X=0.24 $Y=1.65
+ $X2=0.515 $Y2=1.65
r73 19 20 47.3682 $w=2.1e-07 $l=1.5e-07 $layer=POLY_cond $X=2.775 $Y=1.725
+ $X2=2.775 $Y2=1.875
r74 18 20 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=2.805 $Y=2.305
+ $X2=2.805 $Y2=1.875
r75 16 18 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.805 $Y=2.995
+ $X2=2.805 $Y2=2.305
r76 13 19 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=2.745 $Y=0.865
+ $X2=2.745 $Y2=1.725
r77 9 16 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.73 $Y=3.07
+ $X2=2.805 $Y2=2.995
r78 9 10 1002.46 $w=1.5e-07 $l=1.955e-06 $layer=POLY_cond $X=2.73 $Y=3.07
+ $X2=0.775 $Y2=3.07
r79 6 10 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.7 $Y=2.995
+ $X2=0.775 $Y2=3.07
r80 6 8 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=0.7 $Y=2.995 $X2=0.7
+ $Y2=2.305
r81 5 28 22.5156 $w=2.89e-07 $l=2.22486e-07 $layer=POLY_cond $X=0.7 $Y=1.825
+ $X2=0.565 $Y2=1.66
r82 5 8 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.7 $Y=1.825 $X2=0.7
+ $Y2=2.305
r83 1 28 18.0918 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.565 $Y=1.495
+ $X2=0.565 $Y2=1.66
r84 1 3 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=0.565 $Y=1.495
+ $X2=0.565 $Y2=0.815
.ends

.subckt PM_SKY130_FD_SC_LP__HA_2%A_227_397# 1 2 9 11 13 16 20 25 26 27 29 30 31
+ 33 35 38 44 50
c131 38 0 1.1966e-19 $X=1.64 $Y=0.815
c132 30 0 4.83823e-20 $X=3.97 $Y=2.56
c133 29 0 1.50736e-20 $X=2.25 $Y=2.475
c134 26 0 1.2842e-19 $X=2.165 $Y=1.77
c135 25 0 2.15799e-19 $X=1.572 $Y=1.685
r136 49 50 56.8884 $w=2.33e-07 $l=2.75e-07 $layer=POLY_cond $X=4.345 $Y=1.365
+ $X2=4.62 $Y2=1.365
r137 45 49 27.927 $w=2.33e-07 $l=1.35e-07 $layer=POLY_cond $X=4.21 $Y=1.365
+ $X2=4.345 $Y2=1.365
r138 45 47 4.13734 $w=2.33e-07 $l=2e-08 $layer=POLY_cond $X=4.21 $Y=1.365
+ $X2=4.19 $Y2=1.365
r139 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.21
+ $Y=1.35 $X2=4.21 $Y2=1.35
r140 41 44 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=4.055 $Y=1.35
+ $X2=4.21 $Y2=1.35
r141 38 40 8.29153 $w=3.18e-07 $l=1.65e-07 $layer=LI1_cond $X=1.645 $Y=0.815
+ $X2=1.645 $Y2=0.98
r142 35 36 15.3453 $w=2.56e-07 $l=3.22e-07 $layer=LI1_cond $X=1.25 $Y=1.965
+ $X2=1.572 $Y2=1.965
r143 32 41 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.055 $Y=1.515
+ $X2=4.055 $Y2=1.35
r144 32 33 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=4.055 $Y=1.515
+ $X2=4.055 $Y2=2.475
r145 30 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.97 $Y=2.56
+ $X2=4.055 $Y2=2.475
r146 30 31 106.668 $w=1.68e-07 $l=1.635e-06 $layer=LI1_cond $X=3.97 $Y=2.56
+ $X2=2.335 $Y2=2.56
r147 29 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.25 $Y=2.475
+ $X2=2.335 $Y2=2.56
r148 28 29 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=2.25 $Y=1.855
+ $X2=2.25 $Y2=2.475
r149 27 36 5.57291 $w=2.56e-07 $l=2.34915e-07 $layer=LI1_cond $X=1.66 $Y=1.77
+ $X2=1.572 $Y2=1.965
r150 26 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.165 $Y=1.77
+ $X2=2.25 $Y2=1.855
r151 26 27 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=2.165 $Y=1.77
+ $X2=1.66 $Y2=1.77
r152 25 36 2.98828 $w=1.75e-07 $l=2.8e-07 $layer=LI1_cond $X=1.572 $Y=1.685
+ $X2=1.572 $Y2=1.965
r153 25 40 44.6805 $w=1.73e-07 $l=7.05e-07 $layer=LI1_cond $X=1.572 $Y=1.685
+ $X2=1.572 $Y2=0.98
r154 18 50 32.0644 $w=2.33e-07 $l=1.55e-07 $layer=POLY_cond $X=4.775 $Y=1.365
+ $X2=4.62 $Y2=1.365
r155 18 20 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=4.775 $Y=1.365
+ $X2=4.775 $Y2=0.655
r156 14 50 13.0941 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=4.62 $Y=1.515
+ $X2=4.62 $Y2=1.365
r157 14 16 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=4.62 $Y=1.515
+ $X2=4.62 $Y2=2.465
r158 11 49 13.0941 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=4.345 $Y=1.185
+ $X2=4.345 $Y2=1.365
r159 11 13 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=4.345 $Y=1.185
+ $X2=4.345 $Y2=0.655
r160 7 47 13.0941 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=4.19 $Y=1.515
+ $X2=4.19 $Y2=1.365
r161 7 9 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=4.19 $Y=1.515
+ $X2=4.19 $Y2=2.465
r162 2 35 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=1.135
+ $Y=1.985 $X2=1.275 $Y2=2.13
r163 1 38 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.5
+ $Y=0.605 $X2=1.64 $Y2=0.815
.ends

.subckt PM_SKY130_FD_SC_LP__HA_2%VPWR 1 2 3 4 5 18 22 26 30 32 34 39 40 42 43 45
+ 46 47 59 67 72 76
r74 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r75 72 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r76 70 76 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.04 $Y2=3.33
r77 69 70 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r78 67 75 3.55231 $w=1.7e-07 $l=2.32e-07 $layer=LI1_cond $X=4.815 $Y=3.33
+ $X2=5.047 $Y2=3.33
r79 67 69 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=4.815 $Y=3.33
+ $X2=4.56 $Y2=3.33
r80 66 70 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.56 $Y2=3.33
r81 66 73 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=3.12 $Y2=3.33
r82 65 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r83 63 72 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.28 $Y=3.33
+ $X2=3.115 $Y2=3.33
r84 63 65 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=3.28 $Y=3.33 $X2=3.6
+ $Y2=3.33
r85 59 72 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.95 $Y=3.33
+ $X2=3.115 $Y2=3.33
r86 59 61 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=2.95 $Y=3.33
+ $X2=2.64 $Y2=3.33
r87 57 58 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r88 55 58 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r89 54 57 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.72 $Y=3.33 $X2=1.68
+ $Y2=3.33
r90 54 55 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r91 51 55 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r92 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r93 47 73 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r94 47 58 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=1.68 $Y2=3.33
r95 47 61 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r96 45 65 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=3.81 $Y=3.33 $X2=3.6
+ $Y2=3.33
r97 45 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.81 $Y=3.33
+ $X2=3.975 $Y2=3.33
r98 44 69 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=4.14 $Y=3.33
+ $X2=4.56 $Y2=3.33
r99 44 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.14 $Y=3.33
+ $X2=3.975 $Y2=3.33
r100 42 57 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=1.78 $Y=3.33 $X2=1.68
+ $Y2=3.33
r101 42 43 6.25164 $w=1.7e-07 $l=1.07e-07 $layer=LI1_cond $X=1.78 $Y=3.33
+ $X2=1.887 $Y2=3.33
r102 41 61 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=1.995 $Y=3.33
+ $X2=2.64 $Y2=3.33
r103 41 43 6.25164 $w=1.7e-07 $l=1.08e-07 $layer=LI1_cond $X=1.995 $Y=3.33
+ $X2=1.887 $Y2=3.33
r104 39 50 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=0.32 $Y=3.33 $X2=0.24
+ $Y2=3.33
r105 39 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.32 $Y=3.33
+ $X2=0.485 $Y2=3.33
r106 38 54 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=0.65 $Y=3.33 $X2=0.72
+ $Y2=3.33
r107 38 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.65 $Y=3.33
+ $X2=0.485 $Y2=3.33
r108 34 37 53.7909 $w=1.98e-07 $l=9.7e-07 $layer=LI1_cond $X=4.915 $Y=1.98
+ $X2=4.915 $Y2=2.95
r109 32 75 3.32263 $w=2e-07 $l=1.69245e-07 $layer=LI1_cond $X=4.915 $Y=3.245
+ $X2=5.047 $Y2=3.33
r110 32 37 16.3591 $w=1.98e-07 $l=2.95e-07 $layer=LI1_cond $X=4.915 $Y=3.245
+ $X2=4.915 $Y2=2.95
r111 28 46 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.975 $Y=3.245
+ $X2=3.975 $Y2=3.33
r112 28 30 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=3.975 $Y=3.245
+ $X2=3.975 $Y2=2.92
r113 24 72 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.115 $Y=3.245
+ $X2=3.115 $Y2=3.33
r114 24 26 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=3.115 $Y=3.245
+ $X2=3.115 $Y2=2.92
r115 20 43 0.512231 $w=2.15e-07 $l=8.5e-08 $layer=LI1_cond $X=1.887 $Y=3.245
+ $X2=1.887 $Y2=3.33
r116 20 22 44.2216 $w=2.13e-07 $l=8.25e-07 $layer=LI1_cond $X=1.887 $Y=3.245
+ $X2=1.887 $Y2=2.42
r117 16 40 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.485 $Y=3.245
+ $X2=0.485 $Y2=3.33
r118 16 18 38.5894 $w=3.28e-07 $l=1.105e-06 $layer=LI1_cond $X=0.485 $Y=3.245
+ $X2=0.485 $Y2=2.14
r119 5 37 400 $w=1.7e-07 $l=1.21318e-06 $layer=licon1_PDIFF $count=1 $X=4.695
+ $Y=1.835 $X2=4.9 $Y2=2.95
r120 5 34 400 $w=1.7e-07 $l=2.67862e-07 $layer=licon1_PDIFF $count=1 $X=4.695
+ $Y=1.835 $X2=4.9 $Y2=1.98
r121 4 30 600 $w=1.7e-07 $l=1.15288e-06 $layer=licon1_PDIFF $count=1 $X=3.835
+ $Y=1.835 $X2=3.975 $Y2=2.92
r122 3 26 600 $w=1.7e-07 $l=1.04592e-06 $layer=licon1_PDIFF $count=1 $X=2.88
+ $Y=1.985 $X2=3.115 $Y2=2.92
r123 2 22 600 $w=1.7e-07 $l=5.31742e-07 $layer=licon1_PDIFF $count=1 $X=1.675
+ $Y=1.985 $X2=1.89 $Y2=2.42
r124 1 18 300 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_PDIFF $count=2 $X=0.36
+ $Y=1.985 $X2=0.485 $Y2=2.14
.ends

.subckt PM_SKY130_FD_SC_LP__HA_2%COUT 1 2 7 8 9 10 11 20 36
c25 20 0 1.65987e-19 $X=3.545 $Y=0.42
c26 9 0 5.44689e-20 $X=3.6 $Y=1.295
r27 18 36 2.6489 $w=3.33e-07 $l=7.7e-08 $layer=LI1_cond $X=3.557 $Y=0.848
+ $X2=3.557 $Y2=0.925
r28 11 33 4.40024 $w=2.73e-07 $l=1.05e-07 $layer=LI1_cond $X=3.587 $Y=2.035
+ $X2=3.587 $Y2=2.14
r29 10 11 15.5056 $w=2.73e-07 $l=3.7e-07 $layer=LI1_cond $X=3.587 $Y=1.665
+ $X2=3.587 $Y2=2.035
r30 9 10 15.5056 $w=2.73e-07 $l=3.7e-07 $layer=LI1_cond $X=3.587 $Y=1.295
+ $X2=3.587 $Y2=1.665
r31 9 38 11.734 $w=2.73e-07 $l=2.8e-07 $layer=LI1_cond $X=3.587 $Y=1.295
+ $X2=3.587 $Y2=1.015
r32 8 38 3.36228 $w=3.33e-07 $l=8.6e-08 $layer=LI1_cond $X=3.557 $Y=0.929
+ $X2=3.557 $Y2=1.015
r33 8 36 0.137605 $w=3.33e-07 $l=4e-09 $layer=LI1_cond $X=3.557 $Y=0.929
+ $X2=3.557 $Y2=0.925
r34 8 18 0.137605 $w=3.33e-07 $l=4e-09 $layer=LI1_cond $X=3.557 $Y=0.844
+ $X2=3.557 $Y2=0.848
r35 7 8 9.94197 $w=3.33e-07 $l=2.89e-07 $layer=LI1_cond $X=3.557 $Y=0.555
+ $X2=3.557 $Y2=0.844
r36 7 20 4.64417 $w=3.33e-07 $l=1.35e-07 $layer=LI1_cond $X=3.557 $Y=0.555
+ $X2=3.557 $Y2=0.42
r37 2 33 600 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_PDIFF $count=1 $X=3.405
+ $Y=1.835 $X2=3.545 $Y2=2.14
r38 1 20 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=3.405
+ $Y=0.235 $X2=3.545 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__HA_2%SUM 1 2 7 8 9 10 11 12 13 24 34 37
c23 24 0 2.76446e-20 $X=4.56 $Y=0.42
r24 35 37 4.05935 $w=3.33e-07 $l=1.18e-07 $layer=LI1_cond $X=4.477 $Y=1.862
+ $X2=4.477 $Y2=1.98
r25 34 48 1.84848 $w=1.78e-07 $l=3e-08 $layer=LI1_cond $X=4.555 $Y=1.665
+ $X2=4.555 $Y2=1.695
r26 13 45 4.64417 $w=3.33e-07 $l=1.35e-07 $layer=LI1_cond $X=4.477 $Y=2.775
+ $X2=4.477 $Y2=2.91
r27 12 13 12.7285 $w=3.33e-07 $l=3.7e-07 $layer=LI1_cond $X=4.477 $Y=2.405
+ $X2=4.477 $Y2=2.775
r28 11 12 12.7285 $w=3.33e-07 $l=3.7e-07 $layer=LI1_cond $X=4.477 $Y=2.035
+ $X2=4.477 $Y2=2.405
r29 11 37 1.89207 $w=3.33e-07 $l=5.5e-08 $layer=LI1_cond $X=4.477 $Y=2.035
+ $X2=4.477 $Y2=1.98
r30 10 35 4.81618 $w=3.33e-07 $l=1.4e-07 $layer=LI1_cond $X=4.477 $Y=1.722
+ $X2=4.477 $Y2=1.862
r31 10 48 3.38042 $w=3.33e-07 $l=2.7e-08 $layer=LI1_cond $X=4.477 $Y=1.722
+ $X2=4.477 $Y2=1.695
r32 10 34 1.72525 $w=1.78e-07 $l=2.8e-08 $layer=LI1_cond $X=4.555 $Y=1.637
+ $X2=4.555 $Y2=1.665
r33 9 10 21.0727 $w=1.78e-07 $l=3.42e-07 $layer=LI1_cond $X=4.555 $Y=1.295
+ $X2=4.555 $Y2=1.637
r34 8 9 22.798 $w=1.78e-07 $l=3.7e-07 $layer=LI1_cond $X=4.555 $Y=0.925
+ $X2=4.555 $Y2=1.295
r35 7 8 22.798 $w=1.78e-07 $l=3.7e-07 $layer=LI1_cond $X=4.555 $Y=0.555
+ $X2=4.555 $Y2=0.925
r36 7 24 8.31818 $w=1.78e-07 $l=1.35e-07 $layer=LI1_cond $X=4.555 $Y=0.555
+ $X2=4.555 $Y2=0.42
r37 2 45 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=4.265
+ $Y=1.835 $X2=4.405 $Y2=2.91
r38 2 37 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=4.265
+ $Y=1.835 $X2=4.405 $Y2=1.98
r39 1 24 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=4.42
+ $Y=0.235 $X2=4.56 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__HA_2%A_45_121# 1 2 9 11 12 15
r27 13 15 13.7316 $w=2.08e-07 $l=2.6e-07 $layer=LI1_cond $X=1.21 $Y=1.075
+ $X2=1.21 $Y2=0.815
r28 11 13 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=1.105 $Y=1.16
+ $X2=1.21 $Y2=1.075
r29 11 12 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=1.105 $Y=1.16
+ $X2=0.515 $Y2=1.16
r30 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.35 $Y=1.075
+ $X2=0.515 $Y2=1.16
r31 7 9 9.07985 $w=3.28e-07 $l=2.6e-07 $layer=LI1_cond $X=0.35 $Y=1.075 $X2=0.35
+ $Y2=0.815
r32 2 15 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.07
+ $Y=0.605 $X2=1.21 $Y2=0.815
r33 1 9 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.225
+ $Y=0.605 $X2=0.35 $Y2=0.815
.ends

.subckt PM_SKY130_FD_SC_LP__HA_2%VGND 1 2 3 4 17 21 27 29 31 33 35 43 48 54 57
+ 60 64
r62 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r63 60 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r64 57 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r65 54 55 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r66 52 64 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.04
+ $Y2=0
r67 52 61 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=4.08
+ $Y2=0
r68 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r69 49 60 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.225 $Y=0 $X2=4.06
+ $Y2=0
r70 49 51 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=4.225 $Y=0 $X2=4.56
+ $Y2=0
r71 48 63 4.71369 $w=1.7e-07 $l=2.27e-07 $layer=LI1_cond $X=4.825 $Y=0 $X2=5.052
+ $Y2=0
r72 48 51 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=4.825 $Y=0 $X2=4.56
+ $Y2=0
r73 47 61 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r74 47 58 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=3.12
+ $Y2=0
r75 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r76 44 57 10.2049 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=3.22 $Y=0 $X2=3.007
+ $Y2=0
r77 44 46 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=3.22 $Y=0 $X2=3.6
+ $Y2=0
r78 43 60 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.895 $Y=0 $X2=4.06
+ $Y2=0
r79 43 46 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=3.895 $Y=0 $X2=3.6
+ $Y2=0
r80 39 55 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r81 38 41 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.64
+ $Y2=0
r82 38 39 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r83 36 54 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.935 $Y=0 $X2=0.81
+ $Y2=0
r84 36 38 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.935 $Y=0 $X2=1.2
+ $Y2=0
r85 35 57 10.2049 $w=1.7e-07 $l=2.12e-07 $layer=LI1_cond $X=2.795 $Y=0 $X2=3.007
+ $Y2=0
r86 35 41 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=2.795 $Y=0 $X2=2.64
+ $Y2=0
r87 33 58 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r88 33 39 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=2.64 $Y=0 $X2=1.2
+ $Y2=0
r89 33 41 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r90 29 63 3.05248 $w=3.3e-07 $l=1.11781e-07 $layer=LI1_cond $X=4.99 $Y=0.085
+ $X2=5.052 $Y2=0
r91 29 31 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=4.99 $Y=0.085
+ $X2=4.99 $Y2=0.38
r92 25 60 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.06 $Y=0.085
+ $X2=4.06 $Y2=0
r93 25 27 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=4.06 $Y=0.085
+ $X2=4.06 $Y2=0.38
r94 21 23 13.1514 $w=4.23e-07 $l=4.85e-07 $layer=LI1_cond $X=3.007 $Y=0.4
+ $X2=3.007 $Y2=0.885
r95 19 57 1.63918 $w=4.25e-07 $l=8.5e-08 $layer=LI1_cond $X=3.007 $Y=0.085
+ $X2=3.007 $Y2=0
r96 19 21 8.54164 $w=4.23e-07 $l=3.15e-07 $layer=LI1_cond $X=3.007 $Y=0.085
+ $X2=3.007 $Y2=0.4
r97 15 54 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.81 $Y=0.085
+ $X2=0.81 $Y2=0
r98 15 17 30.194 $w=2.48e-07 $l=6.55e-07 $layer=LI1_cond $X=0.81 $Y=0.085
+ $X2=0.81 $Y2=0.74
r99 4 31 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.85
+ $Y=0.235 $X2=4.99 $Y2=0.38
r100 3 27 91 $w=1.7e-07 $l=2.88531e-07 $layer=licon1_NDIFF $count=2 $X=3.835
+ $Y=0.235 $X2=4.06 $Y2=0.38
r101 2 23 182 $w=1.7e-07 $l=2.91719e-07 $layer=licon1_NDIFF $count=1 $X=2.82
+ $Y=0.655 $X2=2.96 $Y2=0.885
r102 2 21 182 $w=1.7e-07 $l=4.02803e-07 $layer=licon1_NDIFF $count=1 $X=2.82
+ $Y=0.655 $X2=3.115 $Y2=0.4
r103 1 17 182 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_NDIFF $count=1 $X=0.64
+ $Y=0.605 $X2=0.78 $Y2=0.74
.ends

