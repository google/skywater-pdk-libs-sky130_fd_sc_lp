* File: sky130_fd_sc_lp__or2_1.pex.spice
* Created: Fri Aug 28 11:21:14 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__OR2_1%B 1 3 5 7 8 10 11 15
c31 1 0 9.68154e-20 $X=0.645 $Y=1.26
r32 13 15 16.6846 $w=2.6e-07 $l=9e-08 $layer=POLY_cond $X=0.27 $Y=1.26 $X2=0.27
+ $Y2=1.35
r33 11 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=1.35 $X2=0.27 $Y2=1.35
r34 8 10 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.72 $Y=1.725
+ $X2=0.72 $Y2=2.045
r35 5 7 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.72 $Y=1.185 $X2=0.72
+ $Y2=0.865
r36 4 15 55.6154 $w=2.6e-07 $l=3.73497e-07 $layer=POLY_cond $X=0.435 $Y=1.65
+ $X2=0.27 $Y2=1.35
r37 3 8 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.645 $Y=1.65
+ $X2=0.72 $Y2=1.725
r38 3 4 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=0.645 $Y=1.65
+ $X2=0.435 $Y2=1.65
r39 2 13 15.628 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.435 $Y=1.26
+ $X2=0.27 $Y2=1.26
r40 1 5 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.645 $Y=1.26
+ $X2=0.72 $Y2=1.185
r41 1 2 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=0.645 $Y=1.26
+ $X2=0.435 $Y2=1.26
.ends

.subckt PM_SKY130_FD_SC_LP__OR2_1%A 3 7 8 9 13 15
c40 9 0 8.30388e-21 $X=1.2 $Y=1.295
r41 13 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.2 $Y=1.35 $X2=1.2
+ $Y2=1.515
r42 13 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.2 $Y=1.35 $X2=1.2
+ $Y2=1.185
r43 9 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.2 $Y=1.35
+ $X2=1.2 $Y2=1.35
r44 8 9 17.561 $w=3.13e-07 $l=4.8e-07 $layer=LI1_cond $X=0.72 $Y=1.357 $X2=1.2
+ $Y2=1.357
r45 7 15 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.15 $Y=0.865
+ $X2=1.15 $Y2=1.185
r46 3 16 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.11 $Y=2.045
+ $X2=1.11 $Y2=1.515
.ends

.subckt PM_SKY130_FD_SC_LP__OR2_1%A_76_367# 1 2 9 13 17 19 20 21 26 28 29 31 35
c64 19 0 9.68154e-20 $X=1.545 $Y=1.77
c65 9 0 8.30388e-21 $X=1.785 $Y=0.655
r66 31 33 3.54598 $w=2.58e-07 $l=8e-08 $layer=LI1_cond $X=0.97 $Y=0.865 $X2=0.97
+ $Y2=0.945
r67 29 38 45.5639 $w=3.95e-07 $l=1.65e-07 $layer=POLY_cond $X=1.802 $Y=1.375
+ $X2=1.802 $Y2=1.54
r68 29 37 45.5639 $w=3.95e-07 $l=1.65e-07 $layer=POLY_cond $X=1.802 $Y=1.375
+ $X2=1.802 $Y2=1.21
r69 28 35 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=1.71 $Y=1.375
+ $X2=1.71 $Y2=1.21
r70 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.77
+ $Y=1.375 $X2=1.77 $Y2=1.375
r71 26 28 10.826 $w=3.28e-07 $l=3.1e-07 $layer=LI1_cond $X=1.71 $Y=1.685
+ $X2=1.71 $Y2=1.375
r72 23 35 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=1.63 $Y=1.03
+ $X2=1.63 $Y2=1.21
r73 22 33 3.22376 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.1 $Y=0.945 $X2=0.97
+ $Y2=0.945
r74 21 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.545 $Y=0.945
+ $X2=1.63 $Y2=1.03
r75 21 22 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=1.545 $Y=0.945
+ $X2=1.1 $Y2=0.945
r76 19 26 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.545 $Y=1.77
+ $X2=1.71 $Y2=1.685
r77 19 20 57.0856 $w=1.68e-07 $l=8.75e-07 $layer=LI1_cond $X=1.545 $Y=1.77
+ $X2=0.67 $Y2=1.77
r78 15 20 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.505 $Y=1.855
+ $X2=0.67 $Y2=1.77
r79 15 17 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=0.505 $Y=1.855
+ $X2=0.505 $Y2=2.045
r80 13 38 474.309 $w=1.5e-07 $l=9.25e-07 $layer=POLY_cond $X=1.925 $Y=2.465
+ $X2=1.925 $Y2=1.54
r81 9 37 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=1.785 $Y=0.655
+ $X2=1.785 $Y2=1.21
r82 2 17 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=0.38
+ $Y=1.835 $X2=0.505 $Y2=2.045
r83 1 31 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.795
+ $Y=0.655 $X2=0.935 $Y2=0.865
.ends

.subckt PM_SKY130_FD_SC_LP__OR2_1%VPWR 1 6 11 13 20 21 24
r18 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r19 21 25 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r20 20 21 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r21 18 24 13.8148 $w=1.7e-07 $l=3.58e-07 $layer=LI1_cond $X=1.875 $Y=3.33
+ $X2=1.517 $Y2=3.33
r22 18 20 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.875 $Y=3.33
+ $X2=2.16 $Y2=3.33
r23 15 16 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r24 13 24 13.8148 $w=1.7e-07 $l=3.57e-07 $layer=LI1_cond $X=1.16 $Y=3.33
+ $X2=1.517 $Y2=3.33
r25 13 15 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=1.16 $Y=3.33
+ $X2=0.24 $Y2=3.33
r26 11 25 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r27 11 16 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.24 $Y2=3.33
r28 11 24 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r29 6 10 7.10956 $w=7.13e-07 $l=4.25e-07 $layer=LI1_cond $X=1.517 $Y=2.11
+ $X2=1.517 $Y2=2.535
r30 4 24 2.90666 $w=7.15e-07 $l=8.5e-08 $layer=LI1_cond $X=1.517 $Y=3.245
+ $X2=1.517 $Y2=3.33
r31 4 10 11.8771 $w=7.13e-07 $l=7.1e-07 $layer=LI1_cond $X=1.517 $Y=3.245
+ $X2=1.517 $Y2=2.535
r32 1 10 300 $w=1.7e-07 $l=9.26013e-07 $layer=licon1_PDIFF $count=2 $X=1.185
+ $Y=1.835 $X2=1.71 $Y2=2.535
r33 1 6 600 $w=1.7e-07 $l=6.48074e-07 $layer=licon1_PDIFF $count=1 $X=1.185
+ $Y=1.835 $X2=1.71 $Y2=2.11
r34 1 6 600 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=1 $X=1.185
+ $Y=1.835 $X2=1.325 $Y2=2.11
.ends

.subckt PM_SKY130_FD_SC_LP__OR2_1%X 1 2 7 8 9 10 11 12 13 23
r16 13 40 5.76222 $w=2.68e-07 $l=1.35e-07 $layer=LI1_cond $X=2.18 $Y=2.775
+ $X2=2.18 $Y2=2.91
r17 12 13 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=2.18 $Y=2.405
+ $X2=2.18 $Y2=2.775
r18 11 12 18.1403 $w=2.68e-07 $l=4.25e-07 $layer=LI1_cond $X=2.18 $Y=1.98
+ $X2=2.18 $Y2=2.405
r19 10 11 13.4452 $w=2.68e-07 $l=3.15e-07 $layer=LI1_cond $X=2.18 $Y=1.665
+ $X2=2.18 $Y2=1.98
r20 9 10 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=2.18 $Y=1.295
+ $X2=2.18 $Y2=1.665
r21 9 44 10.8842 $w=2.68e-07 $l=2.55e-07 $layer=LI1_cond $X=2.18 $Y=1.295
+ $X2=2.18 $Y2=1.04
r22 8 44 4.57673 $w=4.08e-07 $l=1.15e-07 $layer=LI1_cond $X=2.11 $Y=0.925
+ $X2=2.11 $Y2=1.04
r23 8 21 2.52975 $w=4.08e-07 $l=9e-08 $layer=LI1_cond $X=2.11 $Y=0.925 $X2=2.11
+ $Y2=0.835
r24 7 21 7.87034 $w=4.08e-07 $l=2.8e-07 $layer=LI1_cond $X=2.11 $Y=0.555
+ $X2=2.11 $Y2=0.835
r25 7 23 3.79463 $w=4.08e-07 $l=1.35e-07 $layer=LI1_cond $X=2.11 $Y=0.555
+ $X2=2.11 $Y2=0.42
r26 2 40 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=2
+ $Y=1.835 $X2=2.14 $Y2=2.91
r27 2 11 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2
+ $Y=1.835 $X2=2.14 $Y2=1.98
r28 1 23 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=1.86
+ $Y=0.235 $X2=2 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__OR2_1%VGND 1 2 9 13 16 17 19 20 21 31 32
r32 31 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r33 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r34 21 32 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r35 21 25 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.24
+ $Y2=0
r36 21 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r37 19 28 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=1.405 $Y=0 $X2=1.2
+ $Y2=0
r38 19 20 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.405 $Y=0 $X2=1.57
+ $Y2=0
r39 18 31 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=1.735 $Y=0 $X2=2.16
+ $Y2=0
r40 18 20 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.735 $Y=0 $X2=1.57
+ $Y2=0
r41 16 24 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=0.34 $Y=0 $X2=0.24
+ $Y2=0
r42 16 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.34 $Y=0 $X2=0.505
+ $Y2=0
r43 15 28 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=0.67 $Y=0 $X2=1.2
+ $Y2=0
r44 15 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.67 $Y=0 $X2=0.505
+ $Y2=0
r45 11 20 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.57 $Y=0.085
+ $X2=1.57 $Y2=0
r46 11 13 15.3659 $w=3.28e-07 $l=4.4e-07 $layer=LI1_cond $X=1.57 $Y=0.085
+ $X2=1.57 $Y2=0.525
r47 7 17 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.505 $Y=0.085
+ $X2=0.505 $Y2=0
r48 7 9 27.2396 $w=3.28e-07 $l=7.8e-07 $layer=LI1_cond $X=0.505 $Y=0.085
+ $X2=0.505 $Y2=0.865
r49 2 13 182 $w=1.7e-07 $l=4.04815e-07 $layer=licon1_NDIFF $count=1 $X=1.225
+ $Y=0.655 $X2=1.57 $Y2=0.525
r50 1 9 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.38
+ $Y=0.655 $X2=0.505 $Y2=0.865
.ends

