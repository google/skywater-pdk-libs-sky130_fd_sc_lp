* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__mux4_4 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
X0 VGND a_114_119# X VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X1 X a_114_119# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X2 VPWR a_114_119# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X3 a_1525_119# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 a_27_119# S1 a_114_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 VGND S0 a_1041_333# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 a_27_119# a_1041_333# a_1525_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 X a_114_119# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X8 VPWR a_114_119# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X9 a_84_277# S1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X10 a_200_119# S0 a_1157_431# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X11 VPWR A1 a_999_431# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X12 a_999_431# a_1041_333# a_200_119# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X13 VPWR S0 a_1041_333# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X14 a_84_277# S1 VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X15 a_1367_119# S0 a_27_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X16 a_1589_431# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X17 VGND A1 a_952_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X18 a_1110_119# A0 VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X19 X a_114_119# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X20 a_114_119# a_84_277# a_200_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X21 a_27_119# a_84_277# a_114_119# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X22 VGND a_114_119# X VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X23 VGND A3 a_1367_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X24 VPWR A3 a_1403_419# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X25 a_1403_419# a_1041_333# a_27_119# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X26 X a_114_119# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X27 a_27_119# S0 a_1589_431# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X28 a_200_119# a_1041_333# a_1110_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X29 a_114_119# S1 a_200_119# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X30 a_1157_431# A0 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X31 a_952_119# S0 a_200_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
