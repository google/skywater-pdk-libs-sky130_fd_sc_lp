* File: sky130_fd_sc_lp__a41o_m.spice
* Created: Fri Aug 28 10:03:09 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__a41o_m.pex.spice"
.subckt sky130_fd_sc_lp__a41o_m  VNB VPB B1 A1 A2 A3 A4 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* A4	A4
* A3	A3
* A2	A2
* A1	A1
* B1	B1
* VPB	VPB
* VNB	VNB
MM1010 N_VGND_M1010_d N_A_80_153#_M1010_g N_X_M1010_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75002.5
+ A=0.063 P=1.14 MULT=1
MM1004 N_A_80_153#_M1004_d N_B1_M1004_g N_VGND_M1010_d VNB NSHORT L=0.15 W=0.42
+ AD=0.07035 AS=0.0588 PD=0.755 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75002.1 A=0.063 P=1.14 MULT=1
MM1001 A_335_47# N_A1_M1001_g N_A_80_153#_M1004_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0819 AS=0.07035 PD=0.81 PS=0.755 NRD=39.996 NRS=15.708 M=1 R=2.8
+ SA=75001.1 SB=75001.6 A=0.063 P=1.14 MULT=1
MM1006 A_443_47# N_A2_M1006_g A_335_47# VNB NSHORT L=0.15 W=0.42 AD=0.0819
+ AS=0.0819 PD=0.81 PS=0.81 NRD=39.996 NRS=39.996 M=1 R=2.8 SA=75001.6
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1008 A_551_47# N_A3_M1008_g A_443_47# VNB NSHORT L=0.15 W=0.42 AD=0.0441
+ AS=0.0819 PD=0.63 PS=0.81 NRD=14.28 NRS=39.996 M=1 R=2.8 SA=75002.2 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1005 N_VGND_M1005_d N_A4_M1005_g A_551_47# VNB NSHORT L=0.15 W=0.42 AD=0.1113
+ AS=0.0441 PD=1.37 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75002.5 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1009 N_VPWR_M1009_d N_A_80_153#_M1009_g N_X_M1009_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.1113 AS=0.1113 PD=1.37 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1002 N_A_300_508#_M1002_d N_B1_M1002_g N_A_80_153#_M1002_s VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.9 A=0.063 P=1.14 MULT=1
MM1000 N_VPWR_M1000_d N_A1_M1000_g N_A_300_508#_M1002_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75001.5 A=0.063 P=1.14 MULT=1
MM1007 N_A_300_508#_M1007_d N_A2_M1007_g N_VPWR_M1000_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.1
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1003 N_VPWR_M1003_d N_A3_M1003_g N_A_300_508#_M1007_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.5
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1011 N_A_300_508#_M1011_d N_A4_M1011_g N_VPWR_M1003_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.9
+ SB=75000.2 A=0.063 P=1.14 MULT=1
DX12_noxref VNB VPB NWDIODE A=7.8703 P=12.17
*
.include "sky130_fd_sc_lp__a41o_m.pxi.spice"
*
.ends
*
*
