* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__sdfstp_1 CLK D SCD SCE SET_B VGND VNB VPB VPWR Q
X0 VGND SCE a_324_102# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 a_124_128# SCE a_196_128# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 a_1810_463# a_871_47# a_1912_463# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X3 a_196_128# a_324_102# a_27_408# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X4 VPWR a_2598_153# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X5 VPWR a_1912_463# a_2158_231# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X6 VGND SCD a_124_128# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 a_1810_463# a_2158_231# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X8 a_1502_125# SET_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 VPWR SCE a_196_408# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X10 a_196_408# D a_196_128# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X11 a_282_128# a_324_102# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 a_1135_57# a_702_47# a_1221_463# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X13 VGND a_1135_57# a_1847_125# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X14 a_1221_463# a_1263_31# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X15 VPWR a_1135_57# a_1703_379# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X16 a_196_128# a_702_47# a_1135_57# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X17 a_1912_463# a_702_47# a_2116_125# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X18 a_27_408# SCD VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X19 a_1263_31# SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X20 a_702_47# CLK VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X21 VGND a_702_47# a_871_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X22 a_1912_463# a_702_47# a_1703_379# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X23 a_1263_31# a_1135_57# a_1502_125# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X24 VPWR SCE a_324_102# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X25 a_196_128# D a_282_128# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X26 a_2224_125# SET_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X27 a_1221_57# a_1263_31# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X28 a_196_128# a_871_47# a_1135_57# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X29 VPWR SET_B a_1912_463# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X30 a_2598_153# a_1912_463# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X31 a_1847_125# a_871_47# a_1912_463# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X32 a_2116_125# a_2158_231# a_2224_125# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X33 VGND a_1912_463# a_2158_231# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X34 a_2598_153# a_1912_463# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X35 a_1135_57# a_871_47# a_1221_57# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X36 VPWR a_702_47# a_871_47# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X37 a_702_47# CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X38 VGND a_2598_153# Q VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X39 VPWR a_1135_57# a_1263_31# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
.ends
