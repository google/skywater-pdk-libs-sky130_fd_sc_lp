* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__nor2b_2 A B_N VGND VNB VPB VPWR Y
X0 VGND a_40_131# Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X1 a_283_367# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X2 Y A VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X3 a_283_367# a_40_131# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X4 VPWR A a_283_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X5 VGND A Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X6 Y a_40_131# a_283_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X7 a_40_131# B_N VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 a_40_131# B_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X9 Y a_40_131# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
.ends
