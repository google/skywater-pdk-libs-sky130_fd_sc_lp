* File: sky130_fd_sc_lp__o21bai_0.pxi.spice
* Created: Fri Aug 28 11:06:27 2020
* 
x_PM_SKY130_FD_SC_LP__O21BAI_0%B1_N N_B1_N_c_72_n N_B1_N_c_79_n N_B1_N_c_80_n
+ N_B1_N_c_73_n N_B1_N_M1007_g N_B1_N_M1002_g N_B1_N_c_74_n N_B1_N_c_75_n B1_N
+ B1_N B1_N N_B1_N_c_76_n N_B1_N_c_77_n PM_SKY130_FD_SC_LP__O21BAI_0%B1_N
x_PM_SKY130_FD_SC_LP__O21BAI_0%A_39_51# N_A_39_51#_M1007_s N_A_39_51#_M1002_s
+ N_A_39_51#_c_114_n N_A_39_51#_c_115_n N_A_39_51#_c_116_n N_A_39_51#_c_117_n
+ N_A_39_51#_c_118_n N_A_39_51#_M1005_g N_A_39_51#_M1006_g N_A_39_51#_c_119_n
+ N_A_39_51#_c_120_n N_A_39_51#_c_128_n N_A_39_51#_c_121_n N_A_39_51#_c_122_n
+ N_A_39_51#_c_123_n N_A_39_51#_c_124_n N_A_39_51#_c_125_n N_A_39_51#_c_131_n
+ PM_SKY130_FD_SC_LP__O21BAI_0%A_39_51#
x_PM_SKY130_FD_SC_LP__O21BAI_0%A2 N_A2_M1001_g N_A2_M1004_g N_A2_c_202_n
+ N_A2_c_206_n A2 A2 N_A2_c_204_n PM_SKY130_FD_SC_LP__O21BAI_0%A2
x_PM_SKY130_FD_SC_LP__O21BAI_0%A1 N_A1_M1000_g N_A1_M1003_g N_A1_c_246_n
+ N_A1_c_251_n A1 A1 A1 N_A1_c_248_n PM_SKY130_FD_SC_LP__O21BAI_0%A1
x_PM_SKY130_FD_SC_LP__O21BAI_0%VPWR N_VPWR_M1002_d N_VPWR_M1000_d N_VPWR_c_278_n
+ N_VPWR_c_279_n N_VPWR_c_280_n VPWR N_VPWR_c_281_n N_VPWR_c_282_n
+ N_VPWR_c_283_n N_VPWR_c_277_n PM_SKY130_FD_SC_LP__O21BAI_0%VPWR
x_PM_SKY130_FD_SC_LP__O21BAI_0%Y N_Y_M1005_s N_Y_M1006_d N_Y_c_310_n N_Y_c_311_n
+ Y Y Y Y Y N_Y_c_313_n N_Y_c_309_n Y PM_SKY130_FD_SC_LP__O21BAI_0%Y
x_PM_SKY130_FD_SC_LP__O21BAI_0%VGND N_VGND_M1007_d N_VGND_M1001_d N_VGND_c_357_n
+ N_VGND_c_358_n VGND N_VGND_c_359_n N_VGND_c_360_n N_VGND_c_361_n
+ N_VGND_c_362_n N_VGND_c_363_n N_VGND_c_364_n PM_SKY130_FD_SC_LP__O21BAI_0%VGND
x_PM_SKY130_FD_SC_LP__O21BAI_0%A_320_47# N_A_320_47#_M1005_d N_A_320_47#_M1003_d
+ N_A_320_47#_c_396_n N_A_320_47#_c_397_n N_A_320_47#_c_398_n
+ N_A_320_47#_c_399_n PM_SKY130_FD_SC_LP__O21BAI_0%A_320_47#
cc_1 VNB N_B1_N_c_72_n 0.00179832f $X=-0.19 $Y=-0.245 $X2=0.36 $Y2=2.085
cc_2 VNB N_B1_N_c_73_n 0.022919f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=0.785
cc_3 VNB N_B1_N_c_74_n 0.0279338f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.46
cc_4 VNB N_B1_N_c_75_n 0.0185785f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.625
cc_5 VNB N_B1_N_c_76_n 0.0536042f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.12
cc_6 VNB N_B1_N_c_77_n 0.0240474f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.12
cc_7 VNB N_A_39_51#_c_114_n 0.0193853f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=0.465
cc_8 VNB N_A_39_51#_c_115_n 0.0195134f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=2.235
cc_9 VNB N_A_39_51#_c_116_n 0.0174462f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=2.575
cc_10 VNB N_A_39_51#_c_117_n 0.0156525f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.12
cc_11 VNB N_A_39_51#_c_118_n 0.0194732f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_39_51#_c_119_n 0.0213458f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.12
cc_13 VNB N_A_39_51#_c_120_n 0.00510976f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.12
cc_14 VNB N_A_39_51#_c_121_n 0.0151788f $X=-0.19 $Y=-0.245 $X2=0.26 $Y2=2.035
cc_15 VNB N_A_39_51#_c_122_n 0.00759449f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_39_51#_c_123_n 0.00768913f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_39_51#_c_124_n 0.00543769f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_39_51#_c_125_n 0.0233587f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A2_M1001_g 0.0367985f $X=-0.19 $Y=-0.245 $X2=0.92 $Y2=2.16
cc_20 VNB N_A2_c_202_n 0.0215034f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB A2 0.00741604f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A2_c_204_n 0.0158701f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_23 VNB N_A1_M1003_g 0.0500264f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=0.465
cc_24 VNB N_A1_c_246_n 0.022727f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB A1 0.0246633f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A1_c_248_n 0.0185469f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_VPWR_c_277_n 0.123877f $X=-0.19 $Y=-0.245 $X2=0.26 $Y2=2.035
cc_28 VNB Y 0.00800137f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_Y_c_309_n 0.0046936f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_357_n 0.00635798f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=2.575
cc_31 VNB N_VGND_c_358_n 0.00524934f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_359_n 0.0169422f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_33 VNB N_VGND_c_360_n 0.0303161f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_361_n 0.0178095f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_362_n 0.181844f $X=-0.19 $Y=-0.245 $X2=0.26 $Y2=1.665
cc_36 VNB N_VGND_c_363_n 0.0052564f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_364_n 0.00507191f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_320_47#_c_396_n 0.00206415f $X=-0.19 $Y=-0.245 $X2=0.995 $Y2=2.575
cc_39 VNB N_A_320_47#_c_397_n 0.0218029f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_320_47#_c_398_n 0.00323573f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.12
cc_41 VNB N_A_320_47#_c_399_n 0.0207109f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.46
cc_42 VPB N_B1_N_c_72_n 0.0280032f $X=-0.19 $Y=1.655 $X2=0.36 $Y2=2.085
cc_43 VPB N_B1_N_c_79_n 0.048833f $X=-0.19 $Y=1.655 $X2=0.92 $Y2=2.16
cc_44 VPB N_B1_N_c_80_n 0.0152268f $X=-0.19 $Y=1.655 $X2=0.435 $Y2=2.16
cc_45 VPB N_B1_N_M1002_g 0.0240814f $X=-0.19 $Y=1.655 $X2=0.995 $Y2=2.575
cc_46 VPB N_B1_N_c_77_n 0.0297966f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.12
cc_47 VPB N_A_39_51#_c_117_n 0.0238244f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.12
cc_48 VPB N_A_39_51#_M1006_g 0.0213131f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_49 VPB N_A_39_51#_c_128_n 0.0170764f $X=-0.19 $Y=1.655 $X2=0.26 $Y2=1.295
cc_50 VPB N_A_39_51#_c_124_n 0.00799139f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_51 VPB N_A_39_51#_c_125_n 0.0178478f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_52 VPB N_A_39_51#_c_131_n 0.0135602f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_53 VPB N_A2_M1004_g 0.0386062f $X=-0.19 $Y=1.655 $X2=0.535 $Y2=0.465
cc_54 VPB N_A2_c_206_n 0.0157837f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.12
cc_55 VPB A2 0.00397468f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_56 VPB N_A1_M1000_g 0.0456174f $X=-0.19 $Y=1.655 $X2=0.92 $Y2=2.16
cc_57 VPB N_A1_c_246_n 0.00480606f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_58 VPB N_A1_c_251_n 0.0184709f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.12
cc_59 VPB A1 0.0279655f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_60 VPB N_VPWR_c_278_n 0.0192873f $X=-0.19 $Y=1.655 $X2=0.995 $Y2=2.575
cc_61 VPB N_VPWR_c_279_n 0.0123127f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_62 VPB N_VPWR_c_280_n 0.0375394f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_63 VPB N_VPWR_c_281_n 0.0354573f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_64 VPB N_VPWR_c_282_n 0.0297359f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_283_n 0.0066101f $X=-0.19 $Y=1.655 $X2=0.26 $Y2=1.295
cc_66 VPB N_VPWR_c_277_n 0.0883773f $X=-0.19 $Y=1.655 $X2=0.26 $Y2=2.035
cc_67 VPB N_Y_c_310_n 0.00604478f $X=-0.19 $Y=1.655 $X2=0.535 $Y2=0.465
cc_68 VPB N_Y_c_311_n 0.00408715f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_69 VPB Y 0.00268694f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_70 VPB N_Y_c_313_n 0.00332759f $X=-0.19 $Y=1.655 $X2=0.26 $Y2=1.12
cc_71 N_B1_N_c_74_n N_A_39_51#_c_115_n 0.0172275f $X=0.27 $Y=1.46 $X2=0 $Y2=0
cc_72 N_B1_N_c_77_n N_A_39_51#_c_115_n 0.0025504f $X=0.27 $Y=1.12 $X2=0 $Y2=0
cc_73 N_B1_N_c_76_n N_A_39_51#_c_116_n 8.09487e-19 $X=0.27 $Y=1.12 $X2=0 $Y2=0
cc_74 N_B1_N_c_79_n N_A_39_51#_M1006_g 0.00984439f $X=0.92 $Y=2.16 $X2=0 $Y2=0
cc_75 N_B1_N_c_73_n N_A_39_51#_c_119_n 8.09487e-19 $X=0.535 $Y=0.785 $X2=0 $Y2=0
cc_76 N_B1_N_c_79_n N_A_39_51#_c_128_n 0.00733077f $X=0.92 $Y=2.16 $X2=0 $Y2=0
cc_77 N_B1_N_c_73_n N_A_39_51#_c_121_n 0.00107237f $X=0.535 $Y=0.785 $X2=0 $Y2=0
cc_78 N_B1_N_c_73_n N_A_39_51#_c_122_n 0.00812617f $X=0.535 $Y=0.785 $X2=0 $Y2=0
cc_79 N_B1_N_c_76_n N_A_39_51#_c_122_n 0.0102899f $X=0.27 $Y=1.12 $X2=0 $Y2=0
cc_80 N_B1_N_c_77_n N_A_39_51#_c_122_n 0.00141328f $X=0.27 $Y=1.12 $X2=0 $Y2=0
cc_81 N_B1_N_c_76_n N_A_39_51#_c_123_n 0.0108848f $X=0.27 $Y=1.12 $X2=0 $Y2=0
cc_82 N_B1_N_c_77_n N_A_39_51#_c_123_n 0.0222758f $X=0.27 $Y=1.12 $X2=0 $Y2=0
cc_83 N_B1_N_c_72_n N_A_39_51#_c_124_n 0.0044343f $X=0.36 $Y=2.085 $X2=0 $Y2=0
cc_84 N_B1_N_c_79_n N_A_39_51#_c_124_n 0.0159302f $X=0.92 $Y=2.16 $X2=0 $Y2=0
cc_85 N_B1_N_M1002_g N_A_39_51#_c_124_n 0.00527689f $X=0.995 $Y=2.575 $X2=0
+ $Y2=0
cc_86 N_B1_N_c_74_n N_A_39_51#_c_124_n 0.00235336f $X=0.27 $Y=1.46 $X2=0 $Y2=0
cc_87 N_B1_N_c_76_n N_A_39_51#_c_124_n 0.00877317f $X=0.27 $Y=1.12 $X2=0 $Y2=0
cc_88 N_B1_N_c_77_n N_A_39_51#_c_124_n 0.0680934f $X=0.27 $Y=1.12 $X2=0 $Y2=0
cc_89 N_B1_N_c_79_n N_A_39_51#_c_125_n 0.0196413f $X=0.92 $Y=2.16 $X2=0 $Y2=0
cc_90 N_B1_N_c_75_n N_A_39_51#_c_125_n 0.0172275f $X=0.27 $Y=1.625 $X2=0 $Y2=0
cc_91 N_B1_N_c_79_n N_A_39_51#_c_131_n 0.00218086f $X=0.92 $Y=2.16 $X2=0 $Y2=0
cc_92 N_B1_N_M1002_g N_A_39_51#_c_131_n 0.00293115f $X=0.995 $Y=2.575 $X2=0
+ $Y2=0
cc_93 N_B1_N_M1002_g N_VPWR_c_278_n 0.00448979f $X=0.995 $Y=2.575 $X2=0 $Y2=0
cc_94 N_B1_N_M1002_g N_VPWR_c_281_n 0.00457151f $X=0.995 $Y=2.575 $X2=0 $Y2=0
cc_95 N_B1_N_M1002_g N_VPWR_c_277_n 0.00492109f $X=0.995 $Y=2.575 $X2=0 $Y2=0
cc_96 N_B1_N_c_73_n Y 4.75045e-19 $X=0.535 $Y=0.785 $X2=0 $Y2=0
cc_97 N_B1_N_c_79_n N_Y_c_313_n 8.74624e-19 $X=0.92 $Y=2.16 $X2=0 $Y2=0
cc_98 N_B1_N_c_73_n N_Y_c_309_n 0.00349463f $X=0.535 $Y=0.785 $X2=0 $Y2=0
cc_99 N_B1_N_c_73_n N_VGND_c_357_n 0.0107489f $X=0.535 $Y=0.785 $X2=0 $Y2=0
cc_100 N_B1_N_c_73_n N_VGND_c_359_n 0.00346638f $X=0.535 $Y=0.785 $X2=0 $Y2=0
cc_101 N_B1_N_c_73_n N_VGND_c_362_n 0.00512229f $X=0.535 $Y=0.785 $X2=0 $Y2=0
cc_102 N_A_39_51#_c_116_n N_A2_M1001_g 0.00668904f $X=1.385 $Y=1.175 $X2=0 $Y2=0
cc_103 N_A_39_51#_c_118_n N_A2_M1001_g 0.017798f $X=1.525 $Y=0.765 $X2=0 $Y2=0
cc_104 N_A_39_51#_c_117_n N_A2_M1004_g 0.00680097f $X=1.385 $Y=2.065 $X2=0 $Y2=0
cc_105 N_A_39_51#_c_128_n N_A2_M1004_g 0.0186867f $X=1.525 $Y=2.14 $X2=0 $Y2=0
cc_106 N_A_39_51#_c_120_n N_A2_c_202_n 0.0112845f $X=1.385 $Y=1.25 $X2=0 $Y2=0
cc_107 N_A_39_51#_c_117_n N_A2_c_206_n 0.0112845f $X=1.385 $Y=2.065 $X2=0 $Y2=0
cc_108 N_A_39_51#_c_116_n A2 0.00494825f $X=1.385 $Y=1.175 $X2=0 $Y2=0
cc_109 N_A_39_51#_c_119_n A2 0.00202342f $X=1.525 $Y=0.84 $X2=0 $Y2=0
cc_110 N_A_39_51#_c_128_n A2 2.93821e-19 $X=1.525 $Y=2.14 $X2=0 $Y2=0
cc_111 N_A_39_51#_c_116_n N_A2_c_204_n 0.0112845f $X=1.385 $Y=1.175 $X2=0 $Y2=0
cc_112 N_A_39_51#_M1006_g N_VPWR_c_278_n 0.00700688f $X=1.525 $Y=2.685 $X2=0
+ $Y2=0
cc_113 N_A_39_51#_c_128_n N_VPWR_c_278_n 0.00368392f $X=1.525 $Y=2.14 $X2=0
+ $Y2=0
cc_114 N_A_39_51#_c_124_n N_VPWR_c_278_n 0.0153616f $X=0.84 $Y=1.34 $X2=0 $Y2=0
cc_115 N_A_39_51#_c_131_n N_VPWR_c_281_n 0.0059371f $X=0.78 $Y=2.575 $X2=0 $Y2=0
cc_116 N_A_39_51#_M1006_g N_VPWR_c_282_n 0.00499542f $X=1.525 $Y=2.685 $X2=0
+ $Y2=0
cc_117 N_A_39_51#_M1006_g N_VPWR_c_277_n 0.0102159f $X=1.525 $Y=2.685 $X2=0
+ $Y2=0
cc_118 N_A_39_51#_c_131_n N_VPWR_c_277_n 0.00958487f $X=0.78 $Y=2.575 $X2=0
+ $Y2=0
cc_119 N_A_39_51#_c_117_n N_Y_c_310_n 0.00459372f $X=1.385 $Y=2.065 $X2=0 $Y2=0
cc_120 N_A_39_51#_c_128_n N_Y_c_310_n 0.012979f $X=1.525 $Y=2.14 $X2=0 $Y2=0
cc_121 N_A_39_51#_c_128_n N_Y_c_311_n 0.00509219f $X=1.525 $Y=2.14 $X2=0 $Y2=0
cc_122 N_A_39_51#_c_114_n Y 0.0132673f $X=1.31 $Y=1.25 $X2=0 $Y2=0
cc_123 N_A_39_51#_c_116_n Y 0.0101687f $X=1.385 $Y=1.175 $X2=0 $Y2=0
cc_124 N_A_39_51#_c_117_n Y 0.0187624f $X=1.385 $Y=2.065 $X2=0 $Y2=0
cc_125 N_A_39_51#_c_118_n Y 0.00302019f $X=1.525 $Y=0.765 $X2=0 $Y2=0
cc_126 N_A_39_51#_c_119_n Y 0.00678522f $X=1.525 $Y=0.84 $X2=0 $Y2=0
cc_127 N_A_39_51#_c_120_n Y 0.00202444f $X=1.385 $Y=1.25 $X2=0 $Y2=0
cc_128 N_A_39_51#_c_122_n Y 0.0149004f $X=0.675 $Y=0.78 $X2=0 $Y2=0
cc_129 N_A_39_51#_c_124_n Y 0.0886628f $X=0.84 $Y=1.34 $X2=0 $Y2=0
cc_130 N_A_39_51#_c_125_n Y 0.00414202f $X=0.84 $Y=1.34 $X2=0 $Y2=0
cc_131 N_A_39_51#_c_117_n N_Y_c_313_n 0.00151821f $X=1.385 $Y=2.065 $X2=0 $Y2=0
cc_132 N_A_39_51#_c_128_n N_Y_c_313_n 0.00231004f $X=1.525 $Y=2.14 $X2=0 $Y2=0
cc_133 N_A_39_51#_c_124_n N_Y_c_313_n 0.0143864f $X=0.84 $Y=1.34 $X2=0 $Y2=0
cc_134 N_A_39_51#_c_118_n N_Y_c_309_n 0.00385488f $X=1.525 $Y=0.765 $X2=0 $Y2=0
cc_135 N_A_39_51#_c_119_n N_Y_c_309_n 0.0017629f $X=1.525 $Y=0.84 $X2=0 $Y2=0
cc_136 N_A_39_51#_c_115_n N_VGND_c_357_n 7.11221e-19 $X=1.005 $Y=1.25 $X2=0
+ $Y2=0
cc_137 N_A_39_51#_c_118_n N_VGND_c_357_n 0.00262091f $X=1.525 $Y=0.765 $X2=0
+ $Y2=0
cc_138 N_A_39_51#_c_122_n N_VGND_c_357_n 0.0252169f $X=0.675 $Y=0.78 $X2=0 $Y2=0
cc_139 N_A_39_51#_c_121_n N_VGND_c_359_n 0.0136331f $X=0.32 $Y=0.465 $X2=0 $Y2=0
cc_140 N_A_39_51#_c_122_n N_VGND_c_359_n 0.00249195f $X=0.675 $Y=0.78 $X2=0
+ $Y2=0
cc_141 N_A_39_51#_c_118_n N_VGND_c_360_n 0.00564615f $X=1.525 $Y=0.765 $X2=0
+ $Y2=0
cc_142 N_A_39_51#_c_119_n N_VGND_c_360_n 2.13818e-19 $X=1.525 $Y=0.84 $X2=0
+ $Y2=0
cc_143 N_A_39_51#_c_118_n N_VGND_c_362_n 0.0118895f $X=1.525 $Y=0.765 $X2=0
+ $Y2=0
cc_144 N_A_39_51#_c_121_n N_VGND_c_362_n 0.00975073f $X=0.32 $Y=0.465 $X2=0
+ $Y2=0
cc_145 N_A_39_51#_c_122_n N_VGND_c_362_n 0.00581473f $X=0.675 $Y=0.78 $X2=0
+ $Y2=0
cc_146 N_A_39_51#_c_118_n N_A_320_47#_c_396_n 0.00116416f $X=1.525 $Y=0.765
+ $X2=0 $Y2=0
cc_147 N_A_39_51#_c_116_n N_A_320_47#_c_398_n 3.10725e-19 $X=1.385 $Y=1.175
+ $X2=0 $Y2=0
cc_148 N_A_39_51#_c_119_n N_A_320_47#_c_398_n 0.00146055f $X=1.525 $Y=0.84 $X2=0
+ $Y2=0
cc_149 N_A2_M1004_g N_A1_M1000_g 0.0246803f $X=1.955 $Y=2.685 $X2=0 $Y2=0
cc_150 N_A2_M1001_g N_A1_M1003_g 0.032956f $X=1.955 $Y=0.445 $X2=0 $Y2=0
cc_151 A2 N_A1_M1003_g 2.7091e-19 $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_152 N_A2_c_202_n N_A1_c_246_n 0.0246803f $X=1.865 $Y=1.66 $X2=0 $Y2=0
cc_153 N_A2_c_206_n N_A1_c_251_n 0.0246803f $X=1.865 $Y=1.825 $X2=0 $Y2=0
cc_154 N_A2_M1001_g A1 0.00372822f $X=1.955 $Y=0.445 $X2=0 $Y2=0
cc_155 A2 A1 0.0333779f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_156 A2 N_A1_c_248_n 0.00240552f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_157 N_A2_c_204_n N_A1_c_248_n 0.0246803f $X=1.865 $Y=1.32 $X2=0 $Y2=0
cc_158 N_A2_M1004_g N_VPWR_c_282_n 0.0046928f $X=1.955 $Y=2.685 $X2=0 $Y2=0
cc_159 N_A2_M1004_g N_VPWR_c_277_n 0.00899983f $X=1.955 $Y=2.685 $X2=0 $Y2=0
cc_160 N_A2_M1004_g N_Y_c_310_n 0.00530149f $X=1.955 $Y=2.685 $X2=0 $Y2=0
cc_161 N_A2_c_206_n N_Y_c_310_n 0.00136982f $X=1.865 $Y=1.825 $X2=0 $Y2=0
cc_162 A2 N_Y_c_310_n 0.0320222f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_163 N_A2_M1004_g N_Y_c_311_n 0.0171742f $X=1.955 $Y=2.685 $X2=0 $Y2=0
cc_164 N_A2_M1001_g Y 0.00104254f $X=1.955 $Y=0.445 $X2=0 $Y2=0
cc_165 N_A2_M1004_g Y 8.49723e-19 $X=1.955 $Y=2.685 $X2=0 $Y2=0
cc_166 A2 Y 0.0568556f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_167 N_A2_c_204_n Y 5.79218e-19 $X=1.865 $Y=1.32 $X2=0 $Y2=0
cc_168 N_A2_M1001_g N_VGND_c_358_n 0.00316751f $X=1.955 $Y=0.445 $X2=0 $Y2=0
cc_169 N_A2_M1001_g N_VGND_c_360_n 0.00585385f $X=1.955 $Y=0.445 $X2=0 $Y2=0
cc_170 N_A2_M1001_g N_VGND_c_362_n 0.00619488f $X=1.955 $Y=0.445 $X2=0 $Y2=0
cc_171 N_A2_M1001_g N_A_320_47#_c_396_n 0.00183058f $X=1.955 $Y=0.445 $X2=0
+ $Y2=0
cc_172 N_A2_M1001_g N_A_320_47#_c_397_n 0.0114368f $X=1.955 $Y=0.445 $X2=0 $Y2=0
cc_173 A2 N_A_320_47#_c_397_n 0.0116487f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_174 A2 N_A_320_47#_c_398_n 0.0211702f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_175 N_A2_c_204_n N_A_320_47#_c_398_n 0.0012279f $X=1.865 $Y=1.32 $X2=0 $Y2=0
cc_176 N_A1_M1000_g N_VPWR_c_280_n 0.00540376f $X=2.345 $Y=2.685 $X2=0 $Y2=0
cc_177 N_A1_c_251_n N_VPWR_c_280_n 5.95696e-19 $X=2.435 $Y=1.88 $X2=0 $Y2=0
cc_178 A1 N_VPWR_c_280_n 0.0251108f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_179 N_A1_M1000_g N_VPWR_c_282_n 0.00499542f $X=2.345 $Y=2.685 $X2=0 $Y2=0
cc_180 N_A1_M1000_g N_VPWR_c_277_n 0.0101119f $X=2.345 $Y=2.685 $X2=0 $Y2=0
cc_181 N_A1_M1000_g N_Y_c_310_n 4.68513e-19 $X=2.345 $Y=2.685 $X2=0 $Y2=0
cc_182 A1 N_Y_c_310_n 0.00634384f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_183 N_A1_M1000_g N_Y_c_311_n 0.00282382f $X=2.345 $Y=2.685 $X2=0 $Y2=0
cc_184 N_A1_M1003_g N_VGND_c_358_n 0.00319852f $X=2.385 $Y=0.445 $X2=0 $Y2=0
cc_185 N_A1_M1003_g N_VGND_c_361_n 0.00585385f $X=2.385 $Y=0.445 $X2=0 $Y2=0
cc_186 N_A1_M1003_g N_VGND_c_362_n 0.00717808f $X=2.385 $Y=0.445 $X2=0 $Y2=0
cc_187 N_A1_M1003_g N_A_320_47#_c_397_n 0.0143967f $X=2.385 $Y=0.445 $X2=0 $Y2=0
cc_188 A1 N_A_320_47#_c_397_n 0.0351651f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_189 N_A1_c_248_n N_A_320_47#_c_397_n 0.00238f $X=2.435 $Y=1.375 $X2=0 $Y2=0
cc_190 N_A1_M1003_g N_A_320_47#_c_399_n 0.00403231f $X=2.385 $Y=0.445 $X2=0
+ $Y2=0
cc_191 N_VPWR_c_278_n N_Y_c_310_n 0.00432261f $X=1.21 $Y=2.51 $X2=0 $Y2=0
cc_192 N_VPWR_c_278_n N_Y_c_311_n 0.00314598f $X=1.21 $Y=2.51 $X2=0 $Y2=0
cc_193 N_VPWR_c_280_n N_Y_c_311_n 0.0102293f $X=2.56 $Y=2.51 $X2=0 $Y2=0
cc_194 N_VPWR_c_282_n N_Y_c_311_n 0.0158621f $X=2.455 $Y=3.33 $X2=0 $Y2=0
cc_195 N_VPWR_c_277_n N_Y_c_311_n 0.0109918f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_196 N_VPWR_c_278_n N_Y_c_313_n 0.0267375f $X=1.21 $Y=2.51 $X2=0 $Y2=0
cc_197 N_Y_c_309_n N_VGND_c_357_n 0.0197662f $X=1.31 $Y=0.445 $X2=0 $Y2=0
cc_198 N_Y_c_309_n N_VGND_c_360_n 0.0205969f $X=1.31 $Y=0.445 $X2=0 $Y2=0
cc_199 N_Y_M1005_s N_VGND_c_362_n 0.00216892f $X=1.185 $Y=0.235 $X2=0 $Y2=0
cc_200 N_Y_c_309_n N_VGND_c_362_n 0.0140002f $X=1.31 $Y=0.445 $X2=0 $Y2=0
cc_201 Y N_A_320_47#_c_396_n 0.00884662f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_202 Y N_A_320_47#_c_398_n 0.0106271f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_203 N_VGND_c_362_n N_A_320_47#_M1005_d 0.00356149f $X=2.64 $Y=0 $X2=-0.19
+ $Y2=-0.245
cc_204 N_VGND_c_362_n N_A_320_47#_M1003_d 0.00224632f $X=2.64 $Y=0 $X2=0 $Y2=0
cc_205 N_VGND_c_360_n N_A_320_47#_c_396_n 0.0121144f $X=2.04 $Y=0 $X2=0 $Y2=0
cc_206 N_VGND_c_362_n N_A_320_47#_c_396_n 0.00894468f $X=2.64 $Y=0 $X2=0 $Y2=0
cc_207 N_VGND_c_358_n N_A_320_47#_c_397_n 0.0168087f $X=2.17 $Y=0.445 $X2=0
+ $Y2=0
cc_208 N_VGND_c_362_n N_A_320_47#_c_397_n 0.0110909f $X=2.64 $Y=0 $X2=0 $Y2=0
cc_209 N_VGND_c_361_n N_A_320_47#_c_399_n 0.0162611f $X=2.64 $Y=0 $X2=0 $Y2=0
cc_210 N_VGND_c_362_n N_A_320_47#_c_399_n 0.0110561f $X=2.64 $Y=0 $X2=0 $Y2=0
