* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__sdfrtp_4 CLK D RESET_B SCD SCE VGND VNB VPB VPWR Q
X0 VPWR RESET_B a_372_50# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X1 a_27_74# SCE VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 a_217_50# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 VGND a_2555_47# Q VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X4 a_300_50# D a_372_50# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 a_1107_119# a_1047_369# a_1201_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 VPWR RESET_B a_1747_21# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X7 VPWR RESET_B a_881_463# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X8 a_1902_119# a_1524_69# a_1747_21# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 a_2555_47# a_1524_69# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X10 VPWR CLK a_975_255# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X11 a_372_50# SCE a_504_81# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 a_1705_113# a_1747_21# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X13 a_565_463# SCD VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X14 a_1747_21# a_1524_69# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X15 VGND RESET_B a_1902_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X16 a_1005_463# a_1047_369# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X17 a_217_50# a_27_74# a_300_50# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X18 a_27_74# SCE VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X19 VPWR SCE a_407_463# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X20 a_407_463# D a_372_50# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X21 a_372_50# a_975_255# a_881_463# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X22 Q a_2555_47# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X23 a_851_242# a_975_255# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X24 a_1524_69# a_975_255# a_1705_113# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X25 VPWR a_2555_47# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X26 VGND CLK a_975_255# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X27 VGND a_881_463# a_1047_369# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X28 a_1047_369# a_851_242# a_1524_69# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X29 a_1662_533# a_1747_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X30 VPWR a_2555_47# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X31 a_372_50# a_27_74# a_565_463# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X32 a_881_463# a_975_255# a_1005_463# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X33 VGND a_2555_47# Q VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X34 a_372_50# a_851_242# a_881_463# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X35 a_881_463# a_851_242# a_1107_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X36 Q a_2555_47# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X37 Q a_2555_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X38 a_851_242# a_975_255# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X39 a_1047_369# a_975_255# a_1524_69# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X40 VPWR a_881_463# a_1047_369# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X41 a_2555_47# a_1524_69# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X42 Q a_2555_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X43 a_1201_119# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X44 a_504_81# SCD a_217_50# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X45 a_1524_69# a_851_242# a_1662_533# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
.ends
