* File: sky130_fd_sc_lp__buflp_8.pex.spice
* Created: Fri Aug 28 10:12:46 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__BUFLP_8%A 1 3 6 8 10 13 17 19 21 24 26 28 31 33 35
+ 38 40 42 43 44 45 46 74 76 87
c120 1 0 2.10106e-20 $X=0.495 $Y=1.185
r121 76 87 2.62209 $w=3.35e-07 $l=7.2e-08 $layer=LI1_cond $X=2.088 $Y=1.347
+ $X2=2.16 $Y2=1.347
r122 73 74 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=2.645 $Y=1.35
+ $X2=2.715 $Y2=1.35
r123 71 73 42.841 $w=3.3e-07 $l=2.45e-07 $layer=POLY_cond $X=2.4 $Y=1.35
+ $X2=2.645 $Y2=1.35
r124 71 72 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.4
+ $Y=1.35 $X2=2.4 $Y2=1.35
r125 69 71 20.109 $w=3.3e-07 $l=1.15e-07 $layer=POLY_cond $X=2.285 $Y=1.35
+ $X2=2.4 $Y2=1.35
r126 68 69 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=2.215 $Y=1.35
+ $X2=2.285 $Y2=1.35
r127 67 68 62.9501 $w=3.3e-07 $l=3.6e-07 $layer=POLY_cond $X=1.855 $Y=1.35
+ $X2=2.215 $Y2=1.35
r128 66 67 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=1.785 $Y=1.35
+ $X2=1.855 $Y2=1.35
r129 64 66 11.366 $w=3.3e-07 $l=6.5e-08 $layer=POLY_cond $X=1.72 $Y=1.35
+ $X2=1.785 $Y2=1.35
r130 62 64 51.5841 $w=3.3e-07 $l=2.95e-07 $layer=POLY_cond $X=1.425 $Y=1.35
+ $X2=1.72 $Y2=1.35
r131 60 62 7.86876 $w=3.3e-07 $l=4.5e-08 $layer=POLY_cond $X=1.38 $Y=1.35
+ $X2=1.425 $Y2=1.35
r132 60 61 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.38
+ $Y=1.35 $X2=1.38 $Y2=1.35
r133 58 60 4.37153 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=1.355 $Y=1.35
+ $X2=1.38 $Y2=1.35
r134 57 58 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=0.925 $Y=1.35
+ $X2=1.355 $Y2=1.35
r135 55 57 39.3438 $w=3.3e-07 $l=2.25e-07 $layer=POLY_cond $X=0.7 $Y=1.35
+ $X2=0.925 $Y2=1.35
r136 52 55 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=0.495 $Y=1.35
+ $X2=0.7 $Y2=1.35
r137 46 72 8.62477 $w=3.31e-07 $l=2.34e-07 $layer=LI1_cond $X=2.166 $Y=1.347
+ $X2=2.4 $Y2=1.347
r138 46 87 0.221148 $w=3.31e-07 $l=6e-09 $layer=LI1_cond $X=2.166 $Y=1.347
+ $X2=2.16 $Y2=1.347
r139 46 76 0.240809 $w=3.33e-07 $l=7e-09 $layer=LI1_cond $X=2.081 $Y=1.347
+ $X2=2.088 $Y2=1.347
r140 45 46 13.7949 $w=3.33e-07 $l=4.01e-07 $layer=LI1_cond $X=1.68 $Y=1.347
+ $X2=2.081 $Y2=1.347
r141 45 61 10.3204 $w=3.33e-07 $l=3e-07 $layer=LI1_cond $X=1.68 $Y=1.347
+ $X2=1.38 $Y2=1.347
r142 45 64 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.72
+ $Y=1.35 $X2=1.72 $Y2=1.35
r143 44 61 6.19223 $w=3.33e-07 $l=1.8e-07 $layer=LI1_cond $X=1.2 $Y=1.347
+ $X2=1.38 $Y2=1.347
r144 43 44 17.2006 $w=3.33e-07 $l=5e-07 $layer=LI1_cond $X=0.7 $Y=1.347 $X2=1.2
+ $Y2=1.347
r145 43 55 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.7
+ $Y=1.35 $X2=0.7 $Y2=1.35
r146 40 74 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.715 $Y=1.185
+ $X2=2.715 $Y2=1.35
r147 40 42 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.715 $Y=1.185
+ $X2=2.715 $Y2=0.655
r148 36 73 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.645 $Y=1.515
+ $X2=2.645 $Y2=1.35
r149 36 38 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=2.645 $Y=1.515
+ $X2=2.645 $Y2=2.465
r150 33 69 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.285 $Y=1.185
+ $X2=2.285 $Y2=1.35
r151 33 35 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.285 $Y=1.185
+ $X2=2.285 $Y2=0.655
r152 29 68 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.215 $Y=1.515
+ $X2=2.215 $Y2=1.35
r153 29 31 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=2.215 $Y=1.515
+ $X2=2.215 $Y2=2.465
r154 26 67 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.855 $Y=1.185
+ $X2=1.855 $Y2=1.35
r155 26 28 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.855 $Y=1.185
+ $X2=1.855 $Y2=0.655
r156 22 66 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.785 $Y=1.515
+ $X2=1.785 $Y2=1.35
r157 22 24 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=1.785 $Y=1.515
+ $X2=1.785 $Y2=2.465
r158 19 62 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.425 $Y=1.185
+ $X2=1.425 $Y2=1.35
r159 19 21 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.425 $Y=1.185
+ $X2=1.425 $Y2=0.655
r160 15 58 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.355 $Y=1.515
+ $X2=1.355 $Y2=1.35
r161 15 17 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=1.355 $Y=1.515
+ $X2=1.355 $Y2=2.465
r162 11 57 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.925 $Y=1.515
+ $X2=0.925 $Y2=1.35
r163 11 13 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=0.925 $Y=1.515
+ $X2=0.925 $Y2=2.465
r164 8 57 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.925 $Y=1.185
+ $X2=0.925 $Y2=1.35
r165 8 10 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.925 $Y=1.185
+ $X2=0.925 $Y2=0.655
r166 4 52 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=1.515
+ $X2=0.495 $Y2=1.35
r167 4 6 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=0.495 $Y=1.515
+ $X2=0.495 $Y2=2.465
r168 1 52 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=1.185
+ $X2=0.495 $Y2=1.35
r169 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.495 $Y=1.185
+ $X2=0.495 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__BUFLP_8%A_27_47# 1 2 3 4 15 19 23 27 31 35 39 43 47
+ 51 55 59 63 67 71 75 79 83 87 91 95 99 103 107 111 115 119 123 127 131 135 139
+ 143 147 152 153 155 159 161 163 168 172 173 175 179 217
c393 127 0 4.02565e-20 $X=9.565 $Y=0.655
c394 111 0 6.98894e-20 $X=8.565 $Y=0.655
c395 91 0 3.31432e-20 $X=7.135 $Y=0.655
c396 83 0 1.06511e-19 $X=6.705 $Y=0.655
c397 79 0 7.1545e-20 $X=6.615 $Y=2.465
c398 59 0 6.55541e-20 $X=5.415 $Y=0.655
r399 214 215 8.74306 $w=3.3e-07 $l=5e-08 $layer=POLY_cond $X=9.565 $Y=1.43
+ $X2=9.615 $Y2=1.43
r400 213 214 78.6876 $w=3.3e-07 $l=4.5e-07 $layer=POLY_cond $X=9.115 $Y=1.43
+ $X2=9.565 $Y2=1.43
r401 212 213 8.74306 $w=3.3e-07 $l=5e-08 $layer=POLY_cond $X=9.065 $Y=1.43
+ $X2=9.115 $Y2=1.43
r402 211 212 78.6876 $w=3.3e-07 $l=4.5e-07 $layer=POLY_cond $X=8.615 $Y=1.43
+ $X2=9.065 $Y2=1.43
r403 210 211 8.74306 $w=3.3e-07 $l=5e-08 $layer=POLY_cond $X=8.565 $Y=1.43
+ $X2=8.615 $Y2=1.43
r404 209 210 78.6876 $w=3.3e-07 $l=4.5e-07 $layer=POLY_cond $X=8.115 $Y=1.43
+ $X2=8.565 $Y2=1.43
r405 208 209 8.74306 $w=3.3e-07 $l=5e-08 $layer=POLY_cond $X=8.065 $Y=1.43
+ $X2=8.115 $Y2=1.43
r406 207 208 78.6876 $w=3.3e-07 $l=4.5e-07 $layer=POLY_cond $X=7.615 $Y=1.43
+ $X2=8.065 $Y2=1.43
r407 206 207 8.74306 $w=3.3e-07 $l=5e-08 $layer=POLY_cond $X=7.565 $Y=1.43
+ $X2=7.615 $Y2=1.43
r408 205 206 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=7.135 $Y=1.43
+ $X2=7.565 $Y2=1.43
r409 204 205 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=7.115 $Y=1.43
+ $X2=7.135 $Y2=1.43
r410 203 204 71.6931 $w=3.3e-07 $l=4.1e-07 $layer=POLY_cond $X=6.705 $Y=1.43
+ $X2=7.115 $Y2=1.43
r411 202 203 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=6.615 $Y=1.43
+ $X2=6.705 $Y2=1.43
r412 201 202 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=6.275 $Y=1.43
+ $X2=6.615 $Y2=1.43
r413 200 201 27.9778 $w=3.3e-07 $l=1.6e-07 $layer=POLY_cond $X=6.115 $Y=1.43
+ $X2=6.275 $Y2=1.43
r414 199 200 47.2125 $w=3.3e-07 $l=2.7e-07 $layer=POLY_cond $X=5.845 $Y=1.43
+ $X2=6.115 $Y2=1.43
r415 198 199 27.9778 $w=3.3e-07 $l=1.6e-07 $layer=POLY_cond $X=5.685 $Y=1.43
+ $X2=5.845 $Y2=1.43
r416 197 198 47.2125 $w=3.3e-07 $l=2.7e-07 $layer=POLY_cond $X=5.415 $Y=1.43
+ $X2=5.685 $Y2=1.43
r417 196 197 27.9778 $w=3.3e-07 $l=1.6e-07 $layer=POLY_cond $X=5.255 $Y=1.43
+ $X2=5.415 $Y2=1.43
r418 195 196 47.2125 $w=3.3e-07 $l=2.7e-07 $layer=POLY_cond $X=4.985 $Y=1.43
+ $X2=5.255 $Y2=1.43
r419 194 195 27.9778 $w=3.3e-07 $l=1.6e-07 $layer=POLY_cond $X=4.825 $Y=1.43
+ $X2=4.985 $Y2=1.43
r420 193 194 68.1959 $w=3.3e-07 $l=3.9e-07 $layer=POLY_cond $X=4.435 $Y=1.43
+ $X2=4.825 $Y2=1.43
r421 192 193 6.99445 $w=3.3e-07 $l=4e-08 $layer=POLY_cond $X=4.395 $Y=1.43
+ $X2=4.435 $Y2=1.43
r422 191 192 68.1959 $w=3.3e-07 $l=3.9e-07 $layer=POLY_cond $X=4.005 $Y=1.43
+ $X2=4.395 $Y2=1.43
r423 190 191 6.99445 $w=3.3e-07 $l=4e-08 $layer=POLY_cond $X=3.965 $Y=1.43
+ $X2=4.005 $Y2=1.43
r424 189 190 68.1959 $w=3.3e-07 $l=3.9e-07 $layer=POLY_cond $X=3.575 $Y=1.43
+ $X2=3.965 $Y2=1.43
r425 188 189 6.99445 $w=3.3e-07 $l=4e-08 $layer=POLY_cond $X=3.535 $Y=1.43
+ $X2=3.575 $Y2=1.43
r426 184 186 6.99445 $w=3.3e-07 $l=4e-08 $layer=POLY_cond $X=3.105 $Y=1.43
+ $X2=3.145 $Y2=1.43
r427 175 177 5.5876 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=1.21 $Y=0.765
+ $X2=1.21 $Y2=0.925
r428 169 217 68.1959 $w=3.3e-07 $l=3.9e-07 $layer=POLY_cond $X=9.655 $Y=1.43
+ $X2=10.045 $Y2=1.43
r429 169 215 6.99445 $w=3.3e-07 $l=4e-08 $layer=POLY_cond $X=9.655 $Y=1.43
+ $X2=9.615 $Y2=1.43
r430 168 169 14.528 $w=1.7e-07 $l=1.7e-06 $layer=licon1_POLY $count=10 $X=9.655
+ $Y=1.43 $X2=9.655 $Y2=1.43
r431 166 188 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=3.195 $Y=1.43
+ $X2=3.535 $Y2=1.43
r432 166 186 8.74306 $w=3.3e-07 $l=5e-08 $layer=POLY_cond $X=3.195 $Y=1.43
+ $X2=3.145 $Y2=1.43
r433 165 168 225.599 $w=3.28e-07 $l=6.46e-06 $layer=LI1_cond $X=3.195 $Y=1.43
+ $X2=9.655 $Y2=1.43
r434 165 166 14.528 $w=1.7e-07 $l=1.7e-06 $layer=licon1_POLY $count=10 $X=3.195
+ $Y=1.43 $X2=3.195 $Y2=1.43
r435 163 182 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=2.9 $Y=1.43
+ $X2=2.9 $Y2=1.77
r436 163 165 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=2.985 $Y=1.43
+ $X2=3.195 $Y2=1.43
r437 162 179 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.225 $Y=1.77
+ $X2=1.14 $Y2=1.77
r438 161 182 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.815 $Y=1.77
+ $X2=2.9 $Y2=1.77
r439 161 162 103.733 $w=1.68e-07 $l=1.59e-06 $layer=LI1_cond $X=2.815 $Y=1.77
+ $X2=1.225 $Y2=1.77
r440 157 179 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.14 $Y=1.855
+ $X2=1.14 $Y2=1.77
r441 157 159 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=1.14 $Y=1.855
+ $X2=1.14 $Y2=1.98
r442 156 173 2.11342 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.365 $Y=1.77
+ $X2=0.24 $Y2=1.77
r443 155 179 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.055 $Y=1.77
+ $X2=1.14 $Y2=1.77
r444 155 156 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.055 $Y=1.77
+ $X2=0.365 $Y2=1.77
r445 154 172 2.11342 $w=1.7e-07 $l=1.44482e-07 $layer=LI1_cond $X=0.365 $Y=0.925
+ $X2=0.24 $Y2=0.967
r446 153 177 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.045 $Y=0.925
+ $X2=1.21 $Y2=0.925
r447 153 154 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.045 $Y=0.925
+ $X2=0.365 $Y2=0.925
r448 152 173 4.3182 $w=2.1e-07 $l=1.03078e-07 $layer=LI1_cond $X=0.28 $Y=1.685
+ $X2=0.24 $Y2=1.77
r449 151 172 4.3182 $w=2.1e-07 $l=1.46642e-07 $layer=LI1_cond $X=0.28 $Y=1.095
+ $X2=0.24 $Y2=0.967
r450 151 152 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=0.28 $Y=1.095
+ $X2=0.28 $Y2=1.685
r451 147 149 42.8709 $w=2.48e-07 $l=9.3e-07 $layer=LI1_cond $X=0.24 $Y=1.98
+ $X2=0.24 $Y2=2.91
r452 145 173 4.3182 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=0.24 $Y=1.855
+ $X2=0.24 $Y2=1.77
r453 145 147 5.76222 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=0.24 $Y=1.855
+ $X2=0.24 $Y2=1.98
r454 141 172 4.3182 $w=2.1e-07 $l=1.27e-07 $layer=LI1_cond $X=0.24 $Y=0.84
+ $X2=0.24 $Y2=0.967
r455 141 143 19.361 $w=2.48e-07 $l=4.2e-07 $layer=LI1_cond $X=0.24 $Y=0.84
+ $X2=0.24 $Y2=0.42
r456 137 217 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.045 $Y=1.595
+ $X2=10.045 $Y2=1.43
r457 137 139 446.106 $w=1.5e-07 $l=8.7e-07 $layer=POLY_cond $X=10.045 $Y=1.595
+ $X2=10.045 $Y2=2.465
r458 133 217 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.045 $Y=1.265
+ $X2=10.045 $Y2=1.43
r459 133 135 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=10.045 $Y=1.265
+ $X2=10.045 $Y2=0.655
r460 129 215 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.615 $Y=1.595
+ $X2=9.615 $Y2=1.43
r461 129 131 446.106 $w=1.5e-07 $l=8.7e-07 $layer=POLY_cond $X=9.615 $Y=1.595
+ $X2=9.615 $Y2=2.465
r462 125 214 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.565 $Y=1.265
+ $X2=9.565 $Y2=1.43
r463 125 127 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=9.565 $Y=1.265
+ $X2=9.565 $Y2=0.655
r464 121 213 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.115 $Y=1.595
+ $X2=9.115 $Y2=1.43
r465 121 123 446.106 $w=1.5e-07 $l=8.7e-07 $layer=POLY_cond $X=9.115 $Y=1.595
+ $X2=9.115 $Y2=2.465
r466 117 212 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.065 $Y=1.265
+ $X2=9.065 $Y2=1.43
r467 117 119 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=9.065 $Y=1.265
+ $X2=9.065 $Y2=0.655
r468 113 211 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.615 $Y=1.595
+ $X2=8.615 $Y2=1.43
r469 113 115 446.106 $w=1.5e-07 $l=8.7e-07 $layer=POLY_cond $X=8.615 $Y=1.595
+ $X2=8.615 $Y2=2.465
r470 109 210 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.565 $Y=1.265
+ $X2=8.565 $Y2=1.43
r471 109 111 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=8.565 $Y=1.265
+ $X2=8.565 $Y2=0.655
r472 105 209 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.115 $Y=1.595
+ $X2=8.115 $Y2=1.43
r473 105 107 446.106 $w=1.5e-07 $l=8.7e-07 $layer=POLY_cond $X=8.115 $Y=1.595
+ $X2=8.115 $Y2=2.465
r474 101 208 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.065 $Y=1.265
+ $X2=8.065 $Y2=1.43
r475 101 103 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=8.065 $Y=1.265
+ $X2=8.065 $Y2=0.655
r476 97 207 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.615 $Y=1.595
+ $X2=7.615 $Y2=1.43
r477 97 99 446.106 $w=1.5e-07 $l=8.7e-07 $layer=POLY_cond $X=7.615 $Y=1.595
+ $X2=7.615 $Y2=2.465
r478 93 206 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.565 $Y=1.265
+ $X2=7.565 $Y2=1.43
r479 93 95 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=7.565 $Y=1.265
+ $X2=7.565 $Y2=0.655
r480 89 205 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.135 $Y=1.265
+ $X2=7.135 $Y2=1.43
r481 89 91 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=7.135 $Y=1.265
+ $X2=7.135 $Y2=0.655
r482 85 204 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.115 $Y=1.595
+ $X2=7.115 $Y2=1.43
r483 85 87 446.106 $w=1.5e-07 $l=8.7e-07 $layer=POLY_cond $X=7.115 $Y=1.595
+ $X2=7.115 $Y2=2.465
r484 81 203 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.705 $Y=1.265
+ $X2=6.705 $Y2=1.43
r485 81 83 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=6.705 $Y=1.265
+ $X2=6.705 $Y2=0.655
r486 77 202 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.615 $Y=1.595
+ $X2=6.615 $Y2=1.43
r487 77 79 446.106 $w=1.5e-07 $l=8.7e-07 $layer=POLY_cond $X=6.615 $Y=1.595
+ $X2=6.615 $Y2=2.465
r488 73 201 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.275 $Y=1.265
+ $X2=6.275 $Y2=1.43
r489 73 75 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=6.275 $Y=1.265
+ $X2=6.275 $Y2=0.655
r490 69 200 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.115 $Y=1.595
+ $X2=6.115 $Y2=1.43
r491 69 71 446.106 $w=1.5e-07 $l=8.7e-07 $layer=POLY_cond $X=6.115 $Y=1.595
+ $X2=6.115 $Y2=2.465
r492 65 199 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.845 $Y=1.265
+ $X2=5.845 $Y2=1.43
r493 65 67 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=5.845 $Y=1.265
+ $X2=5.845 $Y2=0.655
r494 61 198 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.685 $Y=1.595
+ $X2=5.685 $Y2=1.43
r495 61 63 446.106 $w=1.5e-07 $l=8.7e-07 $layer=POLY_cond $X=5.685 $Y=1.595
+ $X2=5.685 $Y2=2.465
r496 57 197 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.415 $Y=1.265
+ $X2=5.415 $Y2=1.43
r497 57 59 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=5.415 $Y=1.265
+ $X2=5.415 $Y2=0.655
r498 53 196 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.255 $Y=1.595
+ $X2=5.255 $Y2=1.43
r499 53 55 446.106 $w=1.5e-07 $l=8.7e-07 $layer=POLY_cond $X=5.255 $Y=1.595
+ $X2=5.255 $Y2=2.465
r500 49 195 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.985 $Y=1.265
+ $X2=4.985 $Y2=1.43
r501 49 51 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.985 $Y=1.265
+ $X2=4.985 $Y2=0.655
r502 45 194 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.825 $Y=1.595
+ $X2=4.825 $Y2=1.43
r503 45 47 446.106 $w=1.5e-07 $l=8.7e-07 $layer=POLY_cond $X=4.825 $Y=1.595
+ $X2=4.825 $Y2=2.465
r504 41 193 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.435 $Y=1.265
+ $X2=4.435 $Y2=1.43
r505 41 43 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.435 $Y=1.265
+ $X2=4.435 $Y2=0.655
r506 37 192 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.395 $Y=1.595
+ $X2=4.395 $Y2=1.43
r507 37 39 446.106 $w=1.5e-07 $l=8.7e-07 $layer=POLY_cond $X=4.395 $Y=1.595
+ $X2=4.395 $Y2=2.465
r508 33 191 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.005 $Y=1.265
+ $X2=4.005 $Y2=1.43
r509 33 35 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.005 $Y=1.265
+ $X2=4.005 $Y2=0.655
r510 29 190 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.965 $Y=1.595
+ $X2=3.965 $Y2=1.43
r511 29 31 446.106 $w=1.5e-07 $l=8.7e-07 $layer=POLY_cond $X=3.965 $Y=1.595
+ $X2=3.965 $Y2=2.465
r512 25 189 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.575 $Y=1.265
+ $X2=3.575 $Y2=1.43
r513 25 27 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.575 $Y=1.265
+ $X2=3.575 $Y2=0.655
r514 21 188 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.535 $Y=1.595
+ $X2=3.535 $Y2=1.43
r515 21 23 446.106 $w=1.5e-07 $l=8.7e-07 $layer=POLY_cond $X=3.535 $Y=1.595
+ $X2=3.535 $Y2=2.465
r516 17 186 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.145 $Y=1.265
+ $X2=3.145 $Y2=1.43
r517 17 19 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.145 $Y=1.265
+ $X2=3.145 $Y2=0.655
r518 13 184 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.105 $Y=1.595
+ $X2=3.105 $Y2=1.43
r519 13 15 446.106 $w=1.5e-07 $l=8.7e-07 $layer=POLY_cond $X=3.105 $Y=1.595
+ $X2=3.105 $Y2=2.465
r520 4 159 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=1
+ $Y=1.835 $X2=1.14 $Y2=1.98
r521 3 149 400 $w=1.7e-07 $l=1.14521e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.835 $X2=0.28 $Y2=2.91
r522 3 147 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.835 $X2=0.28 $Y2=1.98
r523 2 175 182 $w=1.7e-07 $l=6.26259e-07 $layer=licon1_NDIFF $count=1 $X=1
+ $Y=0.235 $X2=1.21 $Y2=0.765
r524 1 172 182 $w=1.7e-07 $l=7.64068e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.28 $Y2=0.93
r525 1 143 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.28 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__BUFLP_8%A_114_367# 1 2 3 10 12 14 16 17 18 20 22
r42 20 31 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.43 $Y=2.195 $X2=2.43
+ $Y2=2.11
r43 20 22 24.9696 $w=3.28e-07 $l=7.15e-07 $layer=LI1_cond $X=2.43 $Y=2.195
+ $X2=2.43 $Y2=2.91
r44 19 27 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.735 $Y=2.11
+ $X2=1.57 $Y2=2.11
r45 18 31 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.265 $Y=2.11
+ $X2=2.43 $Y2=2.11
r46 18 19 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=2.265 $Y=2.11
+ $X2=1.735 $Y2=2.11
r47 17 29 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.57 $Y=2.905 $X2=1.57
+ $Y2=2.99
r48 16 27 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.57 $Y=2.195 $X2=1.57
+ $Y2=2.11
r49 16 17 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=1.57 $Y=2.195
+ $X2=1.57 $Y2=2.905
r50 15 25 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.875 $Y=2.99
+ $X2=0.71 $Y2=2.99
r51 14 29 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.405 $Y=2.99
+ $X2=1.57 $Y2=2.99
r52 14 15 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=1.405 $Y=2.99
+ $X2=0.875 $Y2=2.99
r53 10 25 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.71 $Y=2.905 $X2=0.71
+ $Y2=2.99
r54 10 12 27.7634 $w=3.28e-07 $l=7.95e-07 $layer=LI1_cond $X=0.71 $Y=2.905
+ $X2=0.71 $Y2=2.11
r55 3 31 400 $w=1.7e-07 $l=4.19196e-07 $layer=licon1_PDIFF $count=1 $X=2.29
+ $Y=1.835 $X2=2.43 $Y2=2.19
r56 3 22 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=2.29
+ $Y=1.835 $X2=2.43 $Y2=2.91
r57 2 29 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=1.43
+ $Y=1.835 $X2=1.57 $Y2=2.91
r58 2 27 400 $w=1.7e-07 $l=4.19196e-07 $layer=licon1_PDIFF $count=1 $X=1.43
+ $Y=1.835 $X2=1.57 $Y2=2.19
r59 1 25 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=0.57
+ $Y=1.835 $X2=0.71 $Y2=2.91
r60 1 12 400 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=1 $X=0.57
+ $Y=1.835 $X2=0.71 $Y2=2.11
.ends

.subckt PM_SKY130_FD_SC_LP__BUFLP_8%VPWR 1 2 3 4 5 6 21 25 31 35 39 45 49 51 56
+ 57 59 60 61 62 63 78 83 89 92 96
r141 95 96 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.32 $Y=3.33
+ $X2=10.32 $Y2=3.33
r142 92 93 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r143 89 90 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r144 87 96 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.84 $Y=3.33
+ $X2=10.32 $Y2=3.33
r145 87 93 1.20413 $w=4.9e-07 $l=4.32e-06 $layer=MET1_cond $X=9.84 $Y=3.33
+ $X2=5.52 $Y2=3.33
r146 86 87 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r147 84 92 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.555 $Y=3.33
+ $X2=5.47 $Y2=3.33
r148 84 86 279.556 $w=1.68e-07 $l=4.285e-06 $layer=LI1_cond $X=5.555 $Y=3.33
+ $X2=9.84 $Y2=3.33
r149 83 95 4.69206 $w=1.7e-07 $l=2.32e-07 $layer=LI1_cond $X=10.095 $Y=3.33
+ $X2=10.327 $Y2=3.33
r150 83 86 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=10.095 $Y=3.33
+ $X2=9.84 $Y2=3.33
r151 82 90 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=4.56 $Y2=3.33
r152 81 82 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r153 79 89 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.695 $Y=3.33
+ $X2=4.61 $Y2=3.33
r154 79 81 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=4.695 $Y=3.33
+ $X2=5.04 $Y2=3.33
r155 78 92 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.385 $Y=3.33
+ $X2=5.47 $Y2=3.33
r156 78 81 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=5.385 $Y=3.33
+ $X2=5.04 $Y2=3.33
r157 77 90 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.56 $Y2=3.33
r158 76 77 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r159 74 77 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r160 73 74 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r161 71 74 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r162 70 71 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r163 67 71 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.68 $Y2=3.33
r164 66 70 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=0.24 $Y=3.33
+ $X2=1.68 $Y2=3.33
r165 66 67 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r166 63 93 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=5.28 $Y=3.33
+ $X2=5.52 $Y2=3.33
r167 63 82 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=5.28 $Y=3.33
+ $X2=5.04 $Y2=3.33
r168 61 76 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=3.665 $Y=3.33
+ $X2=3.6 $Y2=3.33
r169 61 62 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.665 $Y=3.33
+ $X2=3.75 $Y2=3.33
r170 59 73 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=2.775 $Y=3.33
+ $X2=2.64 $Y2=3.33
r171 59 60 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.775 $Y=3.33
+ $X2=2.86 $Y2=3.33
r172 58 76 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=2.945 $Y=3.33
+ $X2=3.6 $Y2=3.33
r173 58 60 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.945 $Y=3.33
+ $X2=2.86 $Y2=3.33
r174 56 70 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=1.915 $Y=3.33
+ $X2=1.68 $Y2=3.33
r175 56 57 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.915 $Y=3.33 $X2=2
+ $Y2=3.33
r176 55 73 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=2.085 $Y=3.33
+ $X2=2.64 $Y2=3.33
r177 55 57 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.085 $Y=3.33 $X2=2
+ $Y2=3.33
r178 51 54 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=10.26 $Y=2.27
+ $X2=10.26 $Y2=2.95
r179 49 95 3.07411 $w=3.3e-07 $l=1.13666e-07 $layer=LI1_cond $X=10.26 $Y=3.245
+ $X2=10.327 $Y2=3.33
r180 49 54 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=10.26 $Y=3.245
+ $X2=10.26 $Y2=2.95
r181 45 48 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=5.47 $Y=2.27
+ $X2=5.47 $Y2=2.95
r182 43 92 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.47 $Y=3.245
+ $X2=5.47 $Y2=3.33
r183 43 48 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=5.47 $Y=3.245
+ $X2=5.47 $Y2=2.95
r184 39 42 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=4.61 $Y=2.27
+ $X2=4.61 $Y2=2.95
r185 37 89 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.61 $Y=3.245
+ $X2=4.61 $Y2=3.33
r186 37 42 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=4.61 $Y=3.245
+ $X2=4.61 $Y2=2.95
r187 36 62 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.835 $Y=3.33
+ $X2=3.75 $Y2=3.33
r188 35 89 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.525 $Y=3.33
+ $X2=4.61 $Y2=3.33
r189 35 36 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=4.525 $Y=3.33
+ $X2=3.835 $Y2=3.33
r190 31 34 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=3.75 $Y=2.27
+ $X2=3.75 $Y2=2.95
r191 29 62 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.75 $Y=3.245
+ $X2=3.75 $Y2=3.33
r192 29 34 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=3.75 $Y=3.245
+ $X2=3.75 $Y2=2.95
r193 25 28 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=2.86 $Y=2.19
+ $X2=2.86 $Y2=2.95
r194 23 60 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.86 $Y=3.245
+ $X2=2.86 $Y2=3.33
r195 23 28 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=2.86 $Y=3.245
+ $X2=2.86 $Y2=2.95
r196 19 57 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2 $Y=3.245 $X2=2
+ $Y2=3.33
r197 19 21 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=2 $Y=3.245 $X2=2
+ $Y2=2.53
r198 6 54 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=10.12
+ $Y=1.835 $X2=10.26 $Y2=2.95
r199 6 51 400 $w=1.7e-07 $l=5.00125e-07 $layer=licon1_PDIFF $count=1 $X=10.12
+ $Y=1.835 $X2=10.26 $Y2=2.27
r200 5 48 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=5.33
+ $Y=1.835 $X2=5.47 $Y2=2.95
r201 5 45 400 $w=1.7e-07 $l=5.00125e-07 $layer=licon1_PDIFF $count=1 $X=5.33
+ $Y=1.835 $X2=5.47 $Y2=2.27
r202 4 42 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=4.47
+ $Y=1.835 $X2=4.61 $Y2=2.95
r203 4 39 400 $w=1.7e-07 $l=5.00125e-07 $layer=licon1_PDIFF $count=1 $X=4.47
+ $Y=1.835 $X2=4.61 $Y2=2.27
r204 3 34 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=3.61
+ $Y=1.835 $X2=3.75 $Y2=2.95
r205 3 31 400 $w=1.7e-07 $l=5.00125e-07 $layer=licon1_PDIFF $count=1 $X=3.61
+ $Y=1.835 $X2=3.75 $Y2=2.27
r206 2 28 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=2.72
+ $Y=1.835 $X2=2.86 $Y2=2.95
r207 2 25 400 $w=1.7e-07 $l=4.19196e-07 $layer=licon1_PDIFF $count=1 $X=2.72
+ $Y=1.835 $X2=2.86 $Y2=2.19
r208 1 21 300 $w=1.7e-07 $l=7.61791e-07 $layer=licon1_PDIFF $count=2 $X=1.86
+ $Y=1.835 $X2=2 $Y2=2.53
.ends

.subckt PM_SKY130_FD_SC_LP__BUFLP_8%A_636_367# 1 2 3 4 5 6 7 8 27 31 32 35 39 43
+ 47 50 52 53 57 59 63 65 69 71 75 77 78 81 82 83
c122 47 0 7.1545e-20 $X=5.735 $Y=1.85
r123 73 75 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=9.83 $Y=2.905
+ $X2=9.83 $Y2=2.27
r124 72 83 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.065 $Y=2.99
+ $X2=8.9 $Y2=2.99
r125 71 73 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.745 $Y=2.99
+ $X2=9.83 $Y2=2.905
r126 71 72 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=9.745 $Y=2.99
+ $X2=9.065 $Y2=2.99
r127 67 83 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.9 $Y=2.905 $X2=8.9
+ $Y2=2.99
r128 67 69 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=8.9 $Y=2.905
+ $X2=8.9 $Y2=2.27
r129 66 82 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.065 $Y=2.99
+ $X2=7.9 $Y2=2.99
r130 65 83 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.735 $Y=2.99
+ $X2=8.9 $Y2=2.99
r131 65 66 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=8.735 $Y=2.99
+ $X2=8.065 $Y2=2.99
r132 61 82 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.9 $Y=2.905 $X2=7.9
+ $Y2=2.99
r133 61 63 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=7.9 $Y=2.905
+ $X2=7.9 $Y2=2.27
r134 60 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.065 $Y=2.99
+ $X2=6.9 $Y2=2.99
r135 59 82 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.735 $Y=2.99
+ $X2=7.9 $Y2=2.99
r136 59 60 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=7.735 $Y=2.99
+ $X2=7.065 $Y2=2.99
r137 55 81 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.9 $Y=2.905 $X2=6.9
+ $Y2=2.99
r138 55 57 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=6.9 $Y=2.905
+ $X2=6.9 $Y2=2.27
r139 54 80 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.065 $Y=2.99
+ $X2=5.9 $Y2=2.99
r140 53 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.735 $Y=2.99
+ $X2=6.9 $Y2=2.99
r141 53 54 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=6.735 $Y=2.99
+ $X2=6.065 $Y2=2.99
r142 50 80 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.9 $Y=2.905 $X2=5.9
+ $Y2=2.99
r143 50 52 32.3033 $w=3.28e-07 $l=9.25e-07 $layer=LI1_cond $X=5.9 $Y=2.905
+ $X2=5.9 $Y2=1.98
r144 49 52 1.57151 $w=3.28e-07 $l=4.5e-08 $layer=LI1_cond $X=5.9 $Y=1.935
+ $X2=5.9 $Y2=1.98
r145 48 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.205 $Y=1.85
+ $X2=5.04 $Y2=1.85
r146 47 49 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.735 $Y=1.85
+ $X2=5.9 $Y2=1.935
r147 47 48 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=5.735 $Y=1.85
+ $X2=5.205 $Y2=1.85
r148 43 45 32.4779 $w=3.28e-07 $l=9.3e-07 $layer=LI1_cond $X=5.04 $Y=1.98
+ $X2=5.04 $Y2=2.91
r149 41 78 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.04 $Y=1.935
+ $X2=5.04 $Y2=1.85
r150 41 43 1.57151 $w=3.28e-07 $l=4.5e-08 $layer=LI1_cond $X=5.04 $Y=1.935
+ $X2=5.04 $Y2=1.98
r151 40 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.345 $Y=1.85
+ $X2=4.18 $Y2=1.85
r152 39 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.875 $Y=1.85
+ $X2=5.04 $Y2=1.85
r153 39 40 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=4.875 $Y=1.85
+ $X2=4.345 $Y2=1.85
r154 35 37 32.4779 $w=3.28e-07 $l=9.3e-07 $layer=LI1_cond $X=4.18 $Y=1.98
+ $X2=4.18 $Y2=2.91
r155 33 77 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.18 $Y=1.935
+ $X2=4.18 $Y2=1.85
r156 33 35 1.57151 $w=3.28e-07 $l=4.5e-08 $layer=LI1_cond $X=4.18 $Y=1.935
+ $X2=4.18 $Y2=1.98
r157 31 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.015 $Y=1.85
+ $X2=4.18 $Y2=1.85
r158 31 32 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=4.015 $Y=1.85
+ $X2=3.485 $Y2=1.85
r159 27 29 32.4779 $w=3.28e-07 $l=9.3e-07 $layer=LI1_cond $X=3.32 $Y=1.98
+ $X2=3.32 $Y2=2.91
r160 25 32 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.32 $Y=1.935
+ $X2=3.485 $Y2=1.85
r161 25 27 1.57151 $w=3.28e-07 $l=4.5e-08 $layer=LI1_cond $X=3.32 $Y=1.935
+ $X2=3.32 $Y2=1.98
r162 8 75 300 $w=1.7e-07 $l=5.00125e-07 $layer=licon1_PDIFF $count=2 $X=9.69
+ $Y=1.835 $X2=9.83 $Y2=2.27
r163 7 69 300 $w=1.7e-07 $l=5.29693e-07 $layer=licon1_PDIFF $count=2 $X=8.69
+ $Y=1.835 $X2=8.9 $Y2=2.27
r164 6 63 300 $w=1.7e-07 $l=5.29693e-07 $layer=licon1_PDIFF $count=2 $X=7.69
+ $Y=1.835 $X2=7.9 $Y2=2.27
r165 5 57 300 $w=1.7e-07 $l=5.29693e-07 $layer=licon1_PDIFF $count=2 $X=6.69
+ $Y=1.835 $X2=6.9 $Y2=2.27
r166 4 80 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=5.76
+ $Y=1.835 $X2=5.9 $Y2=2.91
r167 4 52 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=5.76
+ $Y=1.835 $X2=5.9 $Y2=1.98
r168 3 45 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=4.9
+ $Y=1.835 $X2=5.04 $Y2=2.91
r169 3 43 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=4.9
+ $Y=1.835 $X2=5.04 $Y2=1.98
r170 2 37 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=4.04
+ $Y=1.835 $X2=4.18 $Y2=2.91
r171 2 35 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=4.04
+ $Y=1.835 $X2=4.18 $Y2=1.98
r172 1 29 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=3.18
+ $Y=1.835 $X2=3.32 $Y2=2.91
r173 1 27 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=3.18
+ $Y=1.835 $X2=3.32 $Y2=1.98
.ends

.subckt PM_SKY130_FD_SC_LP__BUFLP_8%X 1 2 3 4 5 6 7 8 27 31 33 34 35 36 39 43 45
+ 47 51 53 55 59 61 63 65 66 68 72 74 78 81 82
c148 53 0 4.02565e-20 $X=9.185 $Y=1.01
c149 45 0 6.98894e-20 $X=8.185 $Y=1.01
r150 81 82 9.691 $w=4.38e-07 $l=3.7e-07 $layer=LI1_cond $X=10.215 $Y=1.295
+ $X2=10.215 $Y2=1.665
r151 80 82 2.61919 $w=4.38e-07 $l=1e-07 $layer=LI1_cond $X=10.215 $Y=1.765
+ $X2=10.215 $Y2=1.665
r152 79 81 5.23838 $w=4.38e-07 $l=2e-07 $layer=LI1_cond $X=10.215 $Y=1.095
+ $X2=10.215 $Y2=1.295
r153 74 76 5.76222 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=9.35 $Y=0.845
+ $X2=9.35 $Y2=1.01
r154 68 70 7.15912 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=8.35 $Y=0.805
+ $X2=8.35 $Y2=1.01
r155 64 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.565 $Y=1.85
+ $X2=9.4 $Y2=1.85
r156 63 80 8.71846 $w=1.7e-07 $l=2.59037e-07 $layer=LI1_cond $X=9.995 $Y=1.85
+ $X2=10.215 $Y2=1.765
r157 63 64 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=9.995 $Y=1.85
+ $X2=9.565 $Y2=1.85
r158 62 76 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.515 $Y=1.01
+ $X2=9.35 $Y2=1.01
r159 61 79 8.71846 $w=1.7e-07 $l=2.59037e-07 $layer=LI1_cond $X=9.995 $Y=1.01
+ $X2=10.215 $Y2=1.095
r160 61 62 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=9.995 $Y=1.01
+ $X2=9.515 $Y2=1.01
r161 57 78 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.4 $Y=1.935 $X2=9.4
+ $Y2=1.85
r162 57 59 1.57151 $w=3.28e-07 $l=4.5e-08 $layer=LI1_cond $X=9.4 $Y=1.935
+ $X2=9.4 $Y2=1.98
r163 56 72 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.565 $Y=1.85
+ $X2=8.4 $Y2=1.85
r164 55 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.235 $Y=1.85
+ $X2=9.4 $Y2=1.85
r165 55 56 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=9.235 $Y=1.85
+ $X2=8.565 $Y2=1.85
r166 54 70 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.515 $Y=1.01
+ $X2=8.35 $Y2=1.01
r167 53 76 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.185 $Y=1.01
+ $X2=9.35 $Y2=1.01
r168 53 54 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=9.185 $Y=1.01
+ $X2=8.515 $Y2=1.01
r169 49 72 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.4 $Y=1.935 $X2=8.4
+ $Y2=1.85
r170 49 51 1.57151 $w=3.28e-07 $l=4.5e-08 $layer=LI1_cond $X=8.4 $Y=1.935
+ $X2=8.4 $Y2=1.98
r171 48 65 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.565 $Y=1.85
+ $X2=7.4 $Y2=1.85
r172 47 72 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.235 $Y=1.85
+ $X2=8.4 $Y2=1.85
r173 47 48 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=8.235 $Y=1.85
+ $X2=7.565 $Y2=1.85
r174 46 66 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.515 $Y=1.01
+ $X2=7.39 $Y2=1.01
r175 45 70 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.185 $Y=1.01
+ $X2=8.35 $Y2=1.01
r176 45 46 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=8.185 $Y=1.01
+ $X2=7.515 $Y2=1.01
r177 41 66 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.39 $Y=0.925
+ $X2=7.39 $Y2=1.01
r178 41 43 3.68782 $w=2.48e-07 $l=8e-08 $layer=LI1_cond $X=7.39 $Y=0.925
+ $X2=7.39 $Y2=0.845
r179 37 65 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.4 $Y=1.935 $X2=7.4
+ $Y2=1.85
r180 37 39 1.57151 $w=3.28e-07 $l=4.5e-08 $layer=LI1_cond $X=7.4 $Y=1.935
+ $X2=7.4 $Y2=1.98
r181 35 66 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.265 $Y=1.01
+ $X2=7.39 $Y2=1.01
r182 35 36 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=7.265 $Y=1.01
+ $X2=6.575 $Y2=1.01
r183 33 65 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.235 $Y=1.85
+ $X2=7.4 $Y2=1.85
r184 33 34 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=7.235 $Y=1.85
+ $X2=6.565 $Y2=1.85
r185 29 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.49 $Y=0.925
+ $X2=6.575 $Y2=1.01
r186 29 31 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=6.49 $Y=0.925
+ $X2=6.49 $Y2=0.845
r187 25 34 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.4 $Y=1.935
+ $X2=6.565 $Y2=1.85
r188 25 27 1.57151 $w=3.28e-07 $l=4.5e-08 $layer=LI1_cond $X=6.4 $Y=1.935
+ $X2=6.4 $Y2=1.98
r189 8 59 300 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=2 $X=9.19
+ $Y=1.835 $X2=9.4 $Y2=1.98
r190 7 51 300 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=2 $X=8.19
+ $Y=1.835 $X2=8.4 $Y2=1.98
r191 6 39 300 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=2 $X=7.19
+ $Y=1.835 $X2=7.4 $Y2=1.98
r192 5 27 300 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=2 $X=6.19
+ $Y=1.835 $X2=6.4 $Y2=1.98
r193 4 74 182 $w=1.7e-07 $l=7.07248e-07 $layer=licon1_NDIFF $count=1 $X=9.14
+ $Y=0.235 $X2=9.35 $Y2=0.845
r194 3 68 182 $w=1.7e-07 $l=6.66783e-07 $layer=licon1_NDIFF $count=1 $X=8.14
+ $Y=0.235 $X2=8.35 $Y2=0.805
r195 2 43 182 $w=1.7e-07 $l=6.76387e-07 $layer=licon1_NDIFF $count=1 $X=7.21
+ $Y=0.235 $X2=7.35 $Y2=0.845
r196 1 31 182 $w=1.7e-07 $l=6.76387e-07 $layer=licon1_NDIFF $count=1 $X=6.35
+ $Y=0.235 $X2=6.49 $Y2=0.845
.ends

.subckt PM_SKY130_FD_SC_LP__BUFLP_8%A_114_47# 1 2 3 10 12 14 15 18 20
c36 10 0 2.10106e-20 $X=1.555 $Y=0.34
r37 20 23 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=0.71 $Y=0.34
+ $X2=0.71 $Y2=0.485
r38 16 18 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=2.5 $Y=0.775
+ $X2=2.5 $Y2=0.42
r39 14 16 7.07017 $w=2.35e-07 $l=2.15708e-07 $layer=LI1_cond $X=2.335 $Y=0.892
+ $X2=2.5 $Y2=0.775
r40 14 15 29.9145 $w=2.33e-07 $l=6.1e-07 $layer=LI1_cond $X=2.335 $Y=0.892
+ $X2=1.725 $Y2=0.892
r41 13 15 7.04737 $w=2.35e-07 $l=1.53734e-07 $layer=LI1_cond $X=1.64 $Y=0.775
+ $X2=1.725 $Y2=0.892
r42 12 26 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.64 $Y=0.425
+ $X2=1.64 $Y2=0.34
r43 12 13 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=1.64 $Y=0.425
+ $X2=1.64 $Y2=0.775
r44 11 20 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.875 $Y=0.34
+ $X2=0.71 $Y2=0.34
r45 10 26 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.555 $Y=0.34
+ $X2=1.64 $Y2=0.34
r46 10 11 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.555 $Y=0.34
+ $X2=0.875 $Y2=0.34
r47 3 18 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=2.36
+ $Y=0.235 $X2=2.5 $Y2=0.42
r48 2 26 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=1.5
+ $Y=0.235 $X2=1.64 $Y2=0.42
r49 1 23 182 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.235 $X2=0.71 $Y2=0.485
.ends

.subckt PM_SKY130_FD_SC_LP__BUFLP_8%VGND 1 2 3 4 5 6 21 25 29 31 35 37 41 43 45
+ 48 49 51 52 53 54 55 70 79 82 86
r144 85 86 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.32 $Y=0
+ $X2=10.32 $Y2=0
r145 82 83 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r146 79 80 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r147 77 86 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.84 $Y=0
+ $X2=10.32 $Y2=0
r148 76 77 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=9.84 $Y=0
+ $X2=9.84 $Y2=0
r149 74 77 1.07034 $w=4.9e-07 $l=3.84e-06 $layer=MET1_cond $X=6 $Y=0 $X2=9.84
+ $Y2=0
r150 74 83 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=5.52
+ $Y2=0
r151 73 76 250.524 $w=1.68e-07 $l=3.84e-06 $layer=LI1_cond $X=6 $Y=0 $X2=9.84
+ $Y2=0
r152 73 74 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=6 $Y=0 $X2=6
+ $Y2=0
r153 71 82 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.715 $Y=0 $X2=5.59
+ $Y2=0
r154 71 73 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=5.715 $Y=0 $X2=6
+ $Y2=0
r155 70 85 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=10.115 $Y=0
+ $X2=10.337 $Y2=0
r156 70 76 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=10.115 $Y=0
+ $X2=9.84 $Y2=0
r157 69 80 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.56
+ $Y2=0
r158 68 69 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r159 66 69 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r160 65 66 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r161 63 66 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r162 62 63 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r163 59 63 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=0.24 $Y=0
+ $X2=1.68 $Y2=0
r164 58 62 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=0.24 $Y=0 $X2=1.68
+ $Y2=0
r165 58 59 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r166 55 83 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=5.28 $Y=0
+ $X2=5.52 $Y2=0
r167 55 80 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=5.28 $Y=0 $X2=4.56
+ $Y2=0
r168 53 68 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=3.625 $Y=0 $X2=3.6
+ $Y2=0
r169 53 54 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.625 $Y=0 $X2=3.75
+ $Y2=0
r170 51 65 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=2.845 $Y=0
+ $X2=2.64 $Y2=0
r171 51 52 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.845 $Y=0 $X2=2.93
+ $Y2=0
r172 50 68 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=3.015 $Y=0 $X2=3.6
+ $Y2=0
r173 50 52 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.015 $Y=0 $X2=2.93
+ $Y2=0
r174 48 62 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=1.905 $Y=0
+ $X2=1.68 $Y2=0
r175 48 49 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.905 $Y=0 $X2=2.03
+ $Y2=0
r176 47 65 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=2.155 $Y=0
+ $X2=2.64 $Y2=0
r177 47 49 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.155 $Y=0 $X2=2.03
+ $Y2=0
r178 43 85 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=10.28 $Y=0.085
+ $X2=10.337 $Y2=0
r179 43 45 13.969 $w=3.28e-07 $l=4e-07 $layer=LI1_cond $X=10.28 $Y=0.085
+ $X2=10.28 $Y2=0.485
r180 39 82 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.59 $Y=0.085
+ $X2=5.59 $Y2=0
r181 39 41 18.4391 $w=2.48e-07 $l=4e-07 $layer=LI1_cond $X=5.59 $Y=0.085
+ $X2=5.59 $Y2=0.485
r182 38 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.815 $Y=0 $X2=4.65
+ $Y2=0
r183 37 82 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.465 $Y=0 $X2=5.59
+ $Y2=0
r184 37 38 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=5.465 $Y=0
+ $X2=4.815 $Y2=0
r185 33 79 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.65 $Y=0.085
+ $X2=4.65 $Y2=0
r186 33 35 13.969 $w=3.28e-07 $l=4e-07 $layer=LI1_cond $X=4.65 $Y=0.085 $X2=4.65
+ $Y2=0.485
r187 32 54 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.875 $Y=0 $X2=3.75
+ $Y2=0
r188 31 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.485 $Y=0 $X2=4.65
+ $Y2=0
r189 31 32 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=4.485 $Y=0
+ $X2=3.875 $Y2=0
r190 27 54 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.75 $Y=0.085
+ $X2=3.75 $Y2=0
r191 27 29 18.4391 $w=2.48e-07 $l=4e-07 $layer=LI1_cond $X=3.75 $Y=0.085
+ $X2=3.75 $Y2=0.485
r192 23 52 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.93 $Y=0.085
+ $X2=2.93 $Y2=0
r193 23 25 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=2.93 $Y=0.085
+ $X2=2.93 $Y2=0.38
r194 19 49 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.03 $Y=0.085
+ $X2=2.03 $Y2=0
r195 19 21 16.3647 $w=2.48e-07 $l=3.55e-07 $layer=LI1_cond $X=2.03 $Y=0.085
+ $X2=2.03 $Y2=0.44
r196 6 45 182 $w=1.7e-07 $l=3.20156e-07 $layer=licon1_NDIFF $count=1 $X=10.12
+ $Y=0.235 $X2=10.28 $Y2=0.485
r197 5 41 182 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=1 $X=5.49
+ $Y=0.235 $X2=5.63 $Y2=0.485
r198 4 35 182 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=1 $X=4.51
+ $Y=0.235 $X2=4.65 $Y2=0.485
r199 3 29 182 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=1 $X=3.65
+ $Y=0.235 $X2=3.79 $Y2=0.485
r200 2 25 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.79
+ $Y=0.235 $X2=2.93 $Y2=0.38
r201 1 21 182 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_NDIFF $count=1 $X=1.93
+ $Y=0.235 $X2=2.07 $Y2=0.44
.ends

.subckt PM_SKY130_FD_SC_LP__BUFLP_8%A_644_47# 1 2 3 4 5 6 7 8 27 29 30 33 35 39
+ 41 43 44 45 47 49 51 55 57 58 61 66 71
c117 47 0 3.3145e-20 $X=7.685 $Y=0.34
c118 45 0 3.31432e-20 $X=6.755 $Y=0.34
c119 43 0 6.55541e-20 $X=6.06 $Y=0.425
c120 41 0 7.33657e-20 $X=5.895 $Y=1.01
r121 71 74 6.46067 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=8.85 $Y=0.34
+ $X2=8.85 $Y2=0.525
r122 66 69 6.46067 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=7.85 $Y=0.34
+ $X2=7.85 $Y2=0.525
r123 61 64 5.76222 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=6.92 $Y=0.34
+ $X2=6.92 $Y2=0.505
r124 53 55 3.68782 $w=2.48e-07 $l=8e-08 $layer=LI1_cond $X=9.82 $Y=0.425
+ $X2=9.82 $Y2=0.505
r125 52 71 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.015 $Y=0.34
+ $X2=8.85 $Y2=0.34
r126 51 53 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=9.695 $Y=0.34
+ $X2=9.82 $Y2=0.425
r127 51 52 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=9.695 $Y=0.34
+ $X2=9.015 $Y2=0.34
r128 50 66 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.015 $Y=0.34
+ $X2=7.85 $Y2=0.34
r129 49 71 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.685 $Y=0.34
+ $X2=8.85 $Y2=0.34
r130 49 50 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=8.685 $Y=0.34
+ $X2=8.015 $Y2=0.34
r131 48 61 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.085 $Y=0.34
+ $X2=6.92 $Y2=0.34
r132 47 66 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.685 $Y=0.34
+ $X2=7.85 $Y2=0.34
r133 47 48 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=7.685 $Y=0.34
+ $X2=7.085 $Y2=0.34
r134 46 60 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.225 $Y=0.34
+ $X2=6.06 $Y2=0.34
r135 45 61 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.755 $Y=0.34
+ $X2=6.92 $Y2=0.34
r136 45 46 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=6.755 $Y=0.34
+ $X2=6.225 $Y2=0.34
r137 43 60 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.06 $Y=0.425
+ $X2=6.06 $Y2=0.34
r138 43 44 17.4613 $w=3.28e-07 $l=5e-07 $layer=LI1_cond $X=6.06 $Y=0.425
+ $X2=6.06 $Y2=0.925
r139 42 58 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.285 $Y=1.01
+ $X2=5.16 $Y2=1.01
r140 41 44 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.895 $Y=1.01
+ $X2=6.06 $Y2=0.925
r141 41 42 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=5.895 $Y=1.01
+ $X2=5.285 $Y2=1.01
r142 37 58 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.16 $Y=0.925
+ $X2=5.16 $Y2=1.01
r143 37 39 23.2793 $w=2.48e-07 $l=5.05e-07 $layer=LI1_cond $X=5.16 $Y=0.925
+ $X2=5.16 $Y2=0.42
r144 36 57 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.305 $Y=1.01
+ $X2=4.18 $Y2=1.01
r145 35 58 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.035 $Y=1.01
+ $X2=5.16 $Y2=1.01
r146 35 36 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=5.035 $Y=1.01
+ $X2=4.305 $Y2=1.01
r147 31 57 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.18 $Y=0.925
+ $X2=4.18 $Y2=1.01
r148 31 33 23.2793 $w=2.48e-07 $l=5.05e-07 $layer=LI1_cond $X=4.18 $Y=0.925
+ $X2=4.18 $Y2=0.42
r149 29 57 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.055 $Y=1.01
+ $X2=4.18 $Y2=1.01
r150 29 30 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=4.055 $Y=1.01
+ $X2=3.445 $Y2=1.01
r151 25 30 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.32 $Y=0.925
+ $X2=3.445 $Y2=1.01
r152 25 27 23.2793 $w=2.48e-07 $l=5.05e-07 $layer=LI1_cond $X=3.32 $Y=0.925
+ $X2=3.32 $Y2=0.42
r153 8 55 182 $w=1.7e-07 $l=3.32716e-07 $layer=licon1_NDIFF $count=1 $X=9.64
+ $Y=0.235 $X2=9.78 $Y2=0.505
r154 7 74 182 $w=1.7e-07 $l=3.80789e-07 $layer=licon1_NDIFF $count=1 $X=8.64
+ $Y=0.235 $X2=8.85 $Y2=0.525
r155 6 69 182 $w=1.7e-07 $l=3.80789e-07 $layer=licon1_NDIFF $count=1 $X=7.64
+ $Y=0.235 $X2=7.85 $Y2=0.525
r156 5 64 182 $w=1.7e-07 $l=3.32716e-07 $layer=licon1_NDIFF $count=1 $X=6.78
+ $Y=0.235 $X2=6.92 $Y2=0.505
r157 4 60 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=5.92
+ $Y=0.235 $X2=6.06 $Y2=0.42
r158 3 39 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=5.06
+ $Y=0.235 $X2=5.2 $Y2=0.42
r159 2 33 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=4.08
+ $Y=0.235 $X2=4.22 $Y2=0.42
r160 1 27 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=3.22
+ $Y=0.235 $X2=3.36 $Y2=0.42
.ends

