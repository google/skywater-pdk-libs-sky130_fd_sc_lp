* File: sky130_fd_sc_lp__o41ai_2.pex.spice
* Created: Fri Aug 28 11:20:26 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O41AI_2%B1 3 7 9 11 12 14 15 16 25
r44 24 26 5.47727 $w=4.84e-07 $l=5.5e-08 $layer=POLY_cond $X=0.9 $Y=1.27
+ $X2=0.955 $Y2=1.27
r45 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.9
+ $Y=1.44 $X2=0.9 $Y2=1.44
r46 22 24 37.345 $w=4.84e-07 $l=3.75e-07 $layer=POLY_cond $X=0.525 $Y=1.27
+ $X2=0.9 $Y2=1.27
r47 20 22 2.48967 $w=4.84e-07 $l=2.5e-08 $layer=POLY_cond $X=0.5 $Y=1.27
+ $X2=0.525 $Y2=1.27
r48 20 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.5 $Y=1.1
+ $X2=0.5 $Y2=1.1
r49 16 25 4.22145 $w=5.08e-07 $l=1.8e-07 $layer=LI1_cond $X=0.72 $Y=1.27 $X2=0.9
+ $Y2=1.27
r50 16 21 5.15955 $w=5.08e-07 $l=2.2e-07 $layer=LI1_cond $X=0.72 $Y=1.27 $X2=0.5
+ $Y2=1.27
r51 15 21 6.09765 $w=5.08e-07 $l=2.6e-07 $layer=LI1_cond $X=0.24 $Y=1.27 $X2=0.5
+ $Y2=1.27
r52 12 14 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.545 $Y=1.185
+ $X2=1.545 $Y2=0.655
r53 9 12 42.8223 $w=4.84e-07 $l=4.3e-07 $layer=POLY_cond $X=1.115 $Y=1.27
+ $X2=1.545 $Y2=1.27
r54 9 26 15.9339 $w=4.84e-07 $l=1.6e-07 $layer=POLY_cond $X=1.115 $Y=1.27
+ $X2=0.955 $Y2=1.27
r55 9 11 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.115 $Y=1.185
+ $X2=1.115 $Y2=0.655
r56 5 26 30.5883 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=0.955 $Y=1.605
+ $X2=0.955 $Y2=1.27
r57 5 7 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=0.955 $Y=1.605
+ $X2=0.955 $Y2=2.465
r58 1 22 30.5883 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=0.525 $Y=1.605
+ $X2=0.525 $Y2=1.27
r59 1 3 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=0.525 $Y=1.605
+ $X2=0.525 $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__O41AI_2%A4 3 7 11 15 17 18 28
c59 28 0 1.06007e-19 $X=2.57 $Y=1.5
c60 11 0 2.40322e-19 $X=2.335 $Y=2.455
r61 26 28 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=2.55 $Y=1.5 $X2=2.57
+ $Y2=1.5
r62 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.55
+ $Y=1.5 $X2=2.55 $Y2=1.5
r63 24 26 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=2.335 $Y=1.5
+ $X2=2.55 $Y2=1.5
r64 23 24 62.9501 $w=3.3e-07 $l=3.6e-07 $layer=POLY_cond $X=1.975 $Y=1.5
+ $X2=2.335 $Y2=1.5
r65 21 23 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=1.905 $Y=1.5 $X2=1.975
+ $Y2=1.5
r66 17 18 13.3295 $w=4.13e-07 $l=4.8e-07 $layer=LI1_cond $X=2.64 $Y=1.542
+ $X2=3.12 $Y2=1.542
r67 17 27 2.49927 $w=4.13e-07 $l=9e-08 $layer=LI1_cond $X=2.64 $Y=1.542 $X2=2.55
+ $Y2=1.542
r68 13 28 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.57 $Y=1.335
+ $X2=2.57 $Y2=1.5
r69 13 15 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=2.57 $Y=1.335
+ $X2=2.57 $Y2=0.655
r70 9 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.335 $Y=1.665
+ $X2=2.335 $Y2=1.5
r71 9 11 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.335 $Y=1.665
+ $X2=2.335 $Y2=2.455
r72 5 23 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.975 $Y=1.335
+ $X2=1.975 $Y2=1.5
r73 5 7 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=1.975 $Y=1.335
+ $X2=1.975 $Y2=0.655
r74 1 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.905 $Y=1.665
+ $X2=1.905 $Y2=1.5
r75 1 3 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.905 $Y=1.665
+ $X2=1.905 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_LP__O41AI_2%A3 3 7 11 15 17 22 23
c53 23 0 1.87136e-19 $X=3.47 $Y=1.5
c54 22 0 1.6433e-19 $X=3.47 $Y=1.5
c55 11 0 1.55482e-19 $X=3.43 $Y=2.455
r56 22 24 2.97531 $w=3.24e-07 $l=2e-08 $layer=POLY_cond $X=3.47 $Y=1.5 $X2=3.49
+ $Y2=1.5
r57 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.47
+ $Y=1.5 $X2=3.47 $Y2=1.5
r58 20 22 5.95062 $w=3.24e-07 $l=4e-08 $layer=POLY_cond $X=3.43 $Y=1.5 $X2=3.47
+ $Y2=1.5
r59 17 23 5.07075 $w=3.73e-07 $l=1.65e-07 $layer=LI1_cond $X=3.572 $Y=1.665
+ $X2=3.572 $Y2=1.5
r60 13 24 20.7868 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.49 $Y=1.335
+ $X2=3.49 $Y2=1.5
r61 13 15 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=3.49 $Y=1.335
+ $X2=3.49 $Y2=0.655
r62 9 20 20.7868 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.43 $Y=1.665
+ $X2=3.43 $Y2=1.5
r63 9 11 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.43 $Y=1.665
+ $X2=3.43 $Y2=2.455
r64 5 20 63.9691 $w=3.24e-07 $l=4.3e-07 $layer=POLY_cond $X=3 $Y=1.5 $X2=3.43
+ $Y2=1.5
r65 5 7 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=3 $Y=1.655 $X2=3
+ $Y2=2.455
r66 1 5 20.7868 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3 $Y=1.335 $X2=3
+ $Y2=1.5
r67 1 3 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=3 $Y=1.335 $X2=3
+ $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__O41AI_2%A2 3 7 9 11 12 13 14 16 17 18 19
c54 19 0 1.55482e-19 $X=5.04 $Y=1.665
c55 12 0 6.58452e-21 $X=4.735 $Y=1.65
c56 9 0 8.11286e-20 $X=4.38 $Y=1.725
r57 27 28 3.92935 $w=3.68e-07 $l=3e-08 $layer=POLY_cond $X=4.35 $Y=1.535
+ $X2=4.38 $Y2=1.535
r58 25 27 27.5054 $w=3.68e-07 $l=2.1e-07 $layer=POLY_cond $X=4.14 $Y=1.535
+ $X2=4.35 $Y2=1.535
r59 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.14
+ $Y=1.51 $X2=4.14 $Y2=1.51
r60 23 25 28.8152 $w=3.68e-07 $l=2.2e-07 $layer=POLY_cond $X=3.92 $Y=1.535
+ $X2=4.14 $Y2=1.535
r61 18 19 13.3295 $w=4.13e-07 $l=4.8e-07 $layer=LI1_cond $X=4.56 $Y=1.542
+ $X2=5.04 $Y2=1.542
r62 18 26 11.6633 $w=4.13e-07 $l=4.2e-07 $layer=LI1_cond $X=4.56 $Y=1.542
+ $X2=4.14 $Y2=1.542
r63 17 26 1.66618 $w=4.13e-07 $l=6e-08 $layer=LI1_cond $X=4.08 $Y=1.542 $X2=4.14
+ $Y2=1.542
r64 14 16 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=4.81 $Y=1.725
+ $X2=4.81 $Y2=2.465
r65 13 28 27.2372 $w=3.68e-07 $l=1.47817e-07 $layer=POLY_cond $X=4.455 $Y=1.65
+ $X2=4.38 $Y2=1.535
r66 12 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.735 $Y=1.65
+ $X2=4.81 $Y2=1.725
r67 12 13 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=4.735 $Y=1.65
+ $X2=4.455 $Y2=1.65
r68 9 28 23.8357 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=4.38 $Y=1.725
+ $X2=4.38 $Y2=1.535
r69 9 11 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=4.38 $Y=1.725
+ $X2=4.38 $Y2=2.465
r70 5 27 23.8357 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=4.35 $Y=1.345
+ $X2=4.35 $Y2=1.535
r71 5 7 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=4.35 $Y=1.345 $X2=4.35
+ $Y2=0.655
r72 1 23 23.8357 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=3.92 $Y=1.345
+ $X2=3.92 $Y2=1.535
r73 1 3 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.92 $Y=1.345 $X2=3.92
+ $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__O41AI_2%A1 1 3 4 5 6 8 11 15 17 18 26
c42 18 0 6.58452e-21 $X=6 $Y=1.665
r43 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.95
+ $Y=1.42 $X2=5.95 $Y2=1.42
r44 26 28 34.4286 $w=3.92e-07 $l=2.8e-07 $layer=POLY_cond $X=5.67 $Y=1.385
+ $X2=5.95 $Y2=1.385
r45 24 26 22.7474 $w=3.92e-07 $l=1.85e-07 $layer=POLY_cond $X=5.485 $Y=1.385
+ $X2=5.67 $Y2=1.385
r46 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.485
+ $Y=1.42 $X2=5.485 $Y2=1.42
r47 22 24 30.125 $w=3.92e-07 $l=2.45e-07 $layer=POLY_cond $X=5.24 $Y=1.385
+ $X2=5.485 $Y2=1.385
r48 21 22 3.68878 $w=3.92e-07 $l=3e-08 $layer=POLY_cond $X=5.21 $Y=1.385
+ $X2=5.24 $Y2=1.385
r49 18 29 1.38849 $w=4.13e-07 $l=5e-08 $layer=LI1_cond $X=6 $Y=1.542 $X2=5.95
+ $Y2=1.542
r50 17 29 11.941 $w=4.13e-07 $l=4.3e-07 $layer=LI1_cond $X=5.52 $Y=1.542
+ $X2=5.95 $Y2=1.542
r51 17 25 0.97194 $w=4.13e-07 $l=3.5e-08 $layer=LI1_cond $X=5.52 $Y=1.542
+ $X2=5.485 $Y2=1.542
r52 13 26 25.3688 $w=1.5e-07 $l=2e-07 $layer=POLY_cond $X=5.67 $Y=1.585 $X2=5.67
+ $Y2=1.385
r53 13 15 451.234 $w=1.5e-07 $l=8.8e-07 $layer=POLY_cond $X=5.67 $Y=1.585
+ $X2=5.67 $Y2=2.465
r54 9 22 25.3688 $w=1.5e-07 $l=2e-07 $layer=POLY_cond $X=5.24 $Y=1.585 $X2=5.24
+ $Y2=1.385
r55 9 11 451.234 $w=1.5e-07 $l=8.8e-07 $layer=POLY_cond $X=5.24 $Y=1.585
+ $X2=5.24 $Y2=2.465
r56 6 21 25.3688 $w=1.5e-07 $l=2e-07 $layer=POLY_cond $X=5.21 $Y=1.185 $X2=5.21
+ $Y2=1.385
r57 6 8 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=5.21 $Y=1.185 $X2=5.21
+ $Y2=0.655
r58 4 21 28.3659 $w=3.92e-07 $l=1.58114e-07 $layer=POLY_cond $X=5.135 $Y=1.26
+ $X2=5.21 $Y2=1.385
r59 4 5 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=5.135 $Y=1.26
+ $X2=4.855 $Y2=1.26
r60 1 5 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.78 $Y=1.185
+ $X2=4.855 $Y2=1.26
r61 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=4.78 $Y=1.185 $X2=4.78
+ $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__O41AI_2%VPWR 1 2 3 10 12 18 24 26 28 33 43 44 50 53
r73 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r74 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r75 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r76 44 54 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=5.52
+ $Y2=3.33
r77 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r78 41 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.62 $Y=3.33
+ $X2=5.455 $Y2=3.33
r79 41 43 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=5.62 $Y=3.33 $X2=6
+ $Y2=3.33
r80 40 54 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=5.52 $Y2=3.33
r81 39 40 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r82 37 51 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r83 36 39 219.209 $w=1.68e-07 $l=3.36e-06 $layer=LI1_cond $X=1.68 $Y=3.33
+ $X2=5.04 $Y2=3.33
r84 36 37 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r85 34 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.335 $Y=3.33
+ $X2=1.17 $Y2=3.33
r86 34 36 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.335 $Y=3.33
+ $X2=1.68 $Y2=3.33
r87 33 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.29 $Y=3.33
+ $X2=5.455 $Y2=3.33
r88 33 39 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=5.29 $Y=3.33
+ $X2=5.04 $Y2=3.33
r89 32 51 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r90 32 48 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r91 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r92 29 47 4.40011 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=3.33
+ $X2=0.222 $Y2=3.33
r93 29 31 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.445 $Y=3.33
+ $X2=0.72 $Y2=3.33
r94 28 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.005 $Y=3.33
+ $X2=1.17 $Y2=3.33
r95 28 31 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.005 $Y=3.33
+ $X2=0.72 $Y2=3.33
r96 26 40 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=5.04 $Y2=3.33
r97 26 37 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=1.68 $Y2=3.33
r98 22 53 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.455 $Y=3.245
+ $X2=5.455 $Y2=3.33
r99 22 24 30.7318 $w=3.28e-07 $l=8.8e-07 $layer=LI1_cond $X=5.455 $Y=3.245
+ $X2=5.455 $Y2=2.365
r100 18 21 28.6365 $w=3.28e-07 $l=8.2e-07 $layer=LI1_cond $X=1.17 $Y=2.13
+ $X2=1.17 $Y2=2.95
r101 16 50 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.17 $Y=3.245
+ $X2=1.17 $Y2=3.33
r102 16 21 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.17 $Y=3.245
+ $X2=1.17 $Y2=2.95
r103 12 15 37.2623 $w=2.98e-07 $l=9.7e-07 $layer=LI1_cond $X=0.295 $Y=1.98
+ $X2=0.295 $Y2=2.95
r104 10 47 3.11756 $w=3e-07 $l=1.15888e-07 $layer=LI1_cond $X=0.295 $Y=3.245
+ $X2=0.222 $Y2=3.33
r105 10 15 11.3324 $w=2.98e-07 $l=2.95e-07 $layer=LI1_cond $X=0.295 $Y=3.245
+ $X2=0.295 $Y2=2.95
r106 3 24 300 $w=1.7e-07 $l=5.95903e-07 $layer=licon1_PDIFF $count=2 $X=5.315
+ $Y=1.835 $X2=5.455 $Y2=2.365
r107 2 21 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=1.03
+ $Y=1.835 $X2=1.17 $Y2=2.95
r108 2 18 400 $w=1.7e-07 $l=3.58225e-07 $layer=licon1_PDIFF $count=1 $X=1.03
+ $Y=1.835 $X2=1.17 $Y2=2.13
r109 1 15 400 $w=1.7e-07 $l=1.17584e-06 $layer=licon1_PDIFF $count=1 $X=0.185
+ $Y=1.835 $X2=0.31 $Y2=2.95
r110 1 12 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.185
+ $Y=1.835 $X2=0.31 $Y2=1.98
.ends

.subckt PM_SKY130_FD_SC_LP__O41AI_2%Y 1 2 3 12 17 20 24 28 29 33
c47 29 0 1.6433e-19 $X=2.16 $Y=1.665
r48 32 33 8.88198 $w=5.38e-07 $l=1.25e-07 $layer=LI1_cond $X=1.36 $Y=1.605
+ $X2=1.235 $Y2=1.605
r49 29 36 0.885984 $w=5.38e-07 $l=4e-08 $layer=LI1_cond $X=2.16 $Y=1.605
+ $X2=2.12 $Y2=1.605
r50 28 36 9.74582 $w=5.38e-07 $l=4.4e-07 $layer=LI1_cond $X=1.68 $Y=1.605
+ $X2=2.12 $Y2=1.605
r51 28 32 7.08787 $w=5.38e-07 $l=3.2e-07 $layer=LI1_cond $X=1.68 $Y=1.605
+ $X2=1.36 $Y2=1.605
r52 24 26 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=2.12 $Y=1.95
+ $X2=2.12 $Y2=2.63
r53 22 36 3.61838 $w=3.3e-07 $l=2.7e-07 $layer=LI1_cond $X=2.12 $Y=1.875
+ $X2=2.12 $Y2=1.605
r54 22 24 2.61919 $w=3.28e-07 $l=7.5e-08 $layer=LI1_cond $X=2.12 $Y=1.875
+ $X2=2.12 $Y2=1.95
r55 18 32 5.26139 $w=2.5e-07 $l=2.7e-07 $layer=LI1_cond $X=1.36 $Y=1.335
+ $X2=1.36 $Y2=1.605
r56 18 20 26.5062 $w=2.48e-07 $l=5.75e-07 $layer=LI1_cond $X=1.36 $Y=1.335
+ $X2=1.36 $Y2=0.76
r57 17 33 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=0.835 $Y=1.79
+ $X2=1.235 $Y2=1.79
r58 12 14 48.7169 $w=2.18e-07 $l=9.3e-07 $layer=LI1_cond $X=0.725 $Y=1.98
+ $X2=0.725 $Y2=2.91
r59 10 17 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=0.725 $Y=1.875
+ $X2=0.835 $Y2=1.79
r60 10 12 5.5003 $w=2.18e-07 $l=1.05e-07 $layer=LI1_cond $X=0.725 $Y=1.875
+ $X2=0.725 $Y2=1.98
r61 3 26 400 $w=1.7e-07 $l=8.72195e-07 $layer=licon1_PDIFF $count=1 $X=1.98
+ $Y=1.825 $X2=2.12 $Y2=2.63
r62 3 24 400 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=1.98
+ $Y=1.825 $X2=2.12 $Y2=1.95
r63 2 14 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=0.6
+ $Y=1.835 $X2=0.74 $Y2=2.91
r64 2 12 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.6
+ $Y=1.835 $X2=0.74 $Y2=1.98
r65 1 20 182 $w=1.7e-07 $l=5.90868e-07 $layer=licon1_NDIFF $count=1 $X=1.19
+ $Y=0.235 $X2=1.33 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_LP__O41AI_2%A_313_365# 1 2 3 10 12 14 16 19 20 22 24
r45 22 31 2.85134 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=3.68 $Y=2.09 $X2=3.68
+ $Y2=2.005
r46 22 24 21.2759 $w=2.58e-07 $l=4.8e-07 $layer=LI1_cond $X=3.68 $Y=2.09
+ $X2=3.68 $Y2=2.57
r47 21 29 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.84 $Y=2.005
+ $X2=2.675 $Y2=2.005
r48 20 31 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.55 $Y=2.005
+ $X2=3.68 $Y2=2.005
r49 20 21 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=3.55 $Y=2.005
+ $X2=2.84 $Y2=2.005
r50 17 19 15.1913 $w=3.28e-07 $l=4.35e-07 $layer=LI1_cond $X=2.675 $Y=2.895
+ $X2=2.675 $Y2=2.46
r51 16 29 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.675 $Y=2.09
+ $X2=2.675 $Y2=2.005
r52 16 19 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=2.675 $Y=2.09
+ $X2=2.675 $Y2=2.46
r53 15 27 4.20357 $w=1.8e-07 $l=1.3e-07 $layer=LI1_cond $X=1.785 $Y=2.985
+ $X2=1.655 $Y2=2.985
r54 14 17 7.61292 $w=1.8e-07 $l=2.05122e-07 $layer=LI1_cond $X=2.51 $Y=2.985
+ $X2=2.675 $Y2=2.895
r55 14 15 44.6717 $w=1.78e-07 $l=7.25e-07 $layer=LI1_cond $X=2.51 $Y=2.985
+ $X2=1.785 $Y2=2.985
r56 10 27 2.91016 $w=2.6e-07 $l=9e-08 $layer=LI1_cond $X=1.655 $Y=2.895
+ $X2=1.655 $Y2=2.985
r57 10 12 30.3624 $w=2.58e-07 $l=6.85e-07 $layer=LI1_cond $X=1.655 $Y=2.895
+ $X2=1.655 $Y2=2.21
r58 3 31 600 $w=1.7e-07 $l=2.4e-07 $layer=licon1_PDIFF $count=1 $X=3.505
+ $Y=1.825 $X2=3.645 $Y2=2.005
r59 3 24 600 $w=1.7e-07 $l=8.11988e-07 $layer=licon1_PDIFF $count=1 $X=3.505
+ $Y=1.825 $X2=3.645 $Y2=2.57
r60 2 29 600 $w=1.7e-07 $l=3.43402e-07 $layer=licon1_PDIFF $count=1 $X=2.41
+ $Y=1.825 $X2=2.675 $Y2=2.005
r61 2 19 300 $w=1.7e-07 $l=7.55976e-07 $layer=licon1_PDIFF $count=2 $X=2.41
+ $Y=1.825 $X2=2.675 $Y2=2.46
r62 1 27 400 $w=1.7e-07 $l=1.1458e-06 $layer=licon1_PDIFF $count=1 $X=1.565
+ $Y=1.825 $X2=1.69 $Y2=2.91
r63 1 12 400 $w=1.7e-07 $l=4.43114e-07 $layer=licon1_PDIFF $count=1 $X=1.565
+ $Y=1.825 $X2=1.69 $Y2=2.21
.ends

.subckt PM_SKY130_FD_SC_LP__O41AI_2%A_615_365# 1 2 9 11 12 15
c27 12 0 1.07931e-19 $X=3.38 $Y=2.99
c28 9 0 1.32391e-19 $X=3.215 $Y=2.365
r29 13 15 18.8582 $w=3.28e-07 $l=5.4e-07 $layer=LI1_cond $X=4.595 $Y=2.905
+ $X2=4.595 $Y2=2.365
r30 11 13 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.43 $Y=2.99
+ $X2=4.595 $Y2=2.905
r31 11 12 68.5027 $w=1.68e-07 $l=1.05e-06 $layer=LI1_cond $X=4.43 $Y=2.99
+ $X2=3.38 $Y2=2.99
r32 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.215 $Y=2.905
+ $X2=3.38 $Y2=2.99
r33 7 9 18.8582 $w=3.28e-07 $l=5.4e-07 $layer=LI1_cond $X=3.215 $Y=2.905
+ $X2=3.215 $Y2=2.365
r34 2 15 300 $w=1.7e-07 $l=5.95903e-07 $layer=licon1_PDIFF $count=2 $X=4.455
+ $Y=1.835 $X2=4.595 $Y2=2.365
r35 1 9 300 $w=1.7e-07 $l=6.0597e-07 $layer=licon1_PDIFF $count=2 $X=3.075
+ $Y=1.825 $X2=3.215 $Y2=2.365
.ends

.subckt PM_SKY130_FD_SC_LP__O41AI_2%A_808_367# 1 2 3 10 12 14 18 20 22 24 29
r32 22 31 2.85134 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=5.92 $Y=2.09 $X2=5.92
+ $Y2=2.005
r33 22 24 15.292 $w=2.58e-07 $l=3.45e-07 $layer=LI1_cond $X=5.92 $Y=2.09
+ $X2=5.92 $Y2=2.435
r34 21 29 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=5.12 $Y=2.005
+ $X2=5.025 $Y2=2.005
r35 20 31 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=5.79 $Y=2.005
+ $X2=5.92 $Y2=2.005
r36 20 21 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.79 $Y=2.005
+ $X2=5.12 $Y2=2.005
r37 16 29 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=5.025 $Y=2.09
+ $X2=5.025 $Y2=2.005
r38 16 18 20.1388 $w=1.88e-07 $l=3.45e-07 $layer=LI1_cond $X=5.025 $Y=2.09
+ $X2=5.025 $Y2=2.435
r39 15 27 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=4.26 $Y=2.005
+ $X2=4.13 $Y2=2.005
r40 14 29 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=4.93 $Y=2.005
+ $X2=5.025 $Y2=2.005
r41 14 15 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.93 $Y=2.005
+ $X2=4.26 $Y2=2.005
r42 10 27 2.85134 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=4.13 $Y=2.09 $X2=4.13
+ $Y2=2.005
r43 10 12 21.2759 $w=2.58e-07 $l=4.8e-07 $layer=LI1_cond $X=4.13 $Y=2.09
+ $X2=4.13 $Y2=2.57
r44 3 31 600 $w=1.7e-07 $l=2.29565e-07 $layer=licon1_PDIFF $count=1 $X=5.745
+ $Y=1.835 $X2=5.885 $Y2=2.005
r45 3 24 300 $w=1.7e-07 $l=6.66333e-07 $layer=licon1_PDIFF $count=2 $X=5.745
+ $Y=1.835 $X2=5.885 $Y2=2.435
r46 2 29 600 $w=1.7e-07 $l=2.29565e-07 $layer=licon1_PDIFF $count=1 $X=4.885
+ $Y=1.835 $X2=5.025 $Y2=2.005
r47 2 18 300 $w=1.7e-07 $l=6.66333e-07 $layer=licon1_PDIFF $count=2 $X=4.885
+ $Y=1.835 $X2=5.025 $Y2=2.435
r48 1 27 600 $w=1.7e-07 $l=2.23942e-07 $layer=licon1_PDIFF $count=1 $X=4.04
+ $Y=1.835 $X2=4.165 $Y2=2.005
r49 1 12 600 $w=1.7e-07 $l=7.95047e-07 $layer=licon1_PDIFF $count=1 $X=4.04
+ $Y=1.835 $X2=4.165 $Y2=2.57
.ends

.subckt PM_SKY130_FD_SC_LP__O41AI_2%A_155_47# 1 2 3 4 5 6 21 23 24 25 26 29 31
+ 35 37 41 43 47 50 53 54 55
r85 45 47 24.5428 $w=2.68e-07 $l=5.75e-07 $layer=LI1_cond $X=5.475 $Y=0.995
+ $X2=5.475 $Y2=0.42
r86 44 55 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=4.66 $Y=1.08
+ $X2=4.565 $Y2=1.08
r87 43 45 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=5.34 $Y=1.08
+ $X2=5.475 $Y2=0.995
r88 43 44 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=5.34 $Y=1.08
+ $X2=4.66 $Y2=1.08
r89 39 55 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=4.565 $Y=0.995
+ $X2=4.565 $Y2=1.08
r90 39 41 33.5646 $w=1.88e-07 $l=5.75e-07 $layer=LI1_cond $X=4.565 $Y=0.995
+ $X2=4.565 $Y2=0.42
r91 38 54 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=3.8 $Y=1.08
+ $X2=3.685 $Y2=1.08
r92 37 55 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=4.47 $Y=1.08
+ $X2=4.565 $Y2=1.08
r93 37 38 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.47 $Y=1.08 $X2=3.8
+ $Y2=1.08
r94 33 54 0.280307 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.685 $Y=0.995
+ $X2=3.685 $Y2=1.08
r95 33 35 28.8111 $w=2.28e-07 $l=5.75e-07 $layer=LI1_cond $X=3.685 $Y=0.995
+ $X2=3.685 $Y2=0.42
r96 32 53 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=2.9 $Y=1.08 $X2=2.76
+ $Y2=1.08
r97 31 54 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=3.57 $Y=1.08
+ $X2=3.685 $Y2=1.08
r98 31 32 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.57 $Y=1.08 $X2=2.9
+ $Y2=1.08
r99 27 53 0.375625 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.76 $Y=0.995
+ $X2=2.76 $Y2=1.08
r100 27 29 23.6662 $w=2.78e-07 $l=5.75e-07 $layer=LI1_cond $X=2.76 $Y=0.995
+ $X2=2.76 $Y2=0.42
r101 25 53 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=2.62 $Y=1.08 $X2=2.76
+ $Y2=1.08
r102 25 26 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=2.62 $Y=1.08
+ $X2=1.925 $Y2=1.08
r103 24 26 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=1.79 $Y=0.995
+ $X2=1.925 $Y2=1.08
r104 23 52 2.81454 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.79 $Y=0.425
+ $X2=1.79 $Y2=0.34
r105 23 24 24.3294 $w=2.68e-07 $l=5.7e-07 $layer=LI1_cond $X=1.79 $Y=0.425
+ $X2=1.79 $Y2=0.995
r106 22 50 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.065 $Y=0.34
+ $X2=0.9 $Y2=0.34
r107 21 52 4.47015 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=1.655 $Y=0.34
+ $X2=1.79 $Y2=0.34
r108 21 22 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=1.655 $Y=0.34
+ $X2=1.065 $Y2=0.34
r109 6 47 91 $w=1.7e-07 $l=2.52636e-07 $layer=licon1_NDIFF $count=2 $X=5.285
+ $Y=0.235 $X2=5.445 $Y2=0.42
r110 5 41 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=4.425
+ $Y=0.235 $X2=4.565 $Y2=0.42
r111 4 35 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=3.565
+ $Y=0.235 $X2=3.705 $Y2=0.42
r112 3 29 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=2.645
+ $Y=0.235 $X2=2.785 $Y2=0.42
r113 2 52 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=1.62
+ $Y=0.235 $X2=1.76 $Y2=0.42
r114 1 50 91 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=2 $X=0.775
+ $Y=0.235 $X2=0.9 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_LP__O41AI_2%VGND 1 2 3 4 15 17 21 25 29 31 33 38 43 50
+ 51 54 57 60 63
r76 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r77 60 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r78 54 55 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r79 51 64 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=0 $X2=5.04
+ $Y2=0
r80 50 51 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=0 $X2=6 $Y2=0
r81 48 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.16 $Y=0 $X2=4.995
+ $Y2=0
r82 48 50 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=5.16 $Y=0 $X2=6
+ $Y2=0
r83 47 64 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.04
+ $Y2=0
r84 47 61 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=4.08
+ $Y2=0
r85 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r86 44 60 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.3 $Y=0 $X2=4.135
+ $Y2=0
r87 44 46 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=4.3 $Y=0 $X2=4.56
+ $Y2=0
r88 43 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.83 $Y=0 $X2=4.995
+ $Y2=0
r89 43 46 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=4.83 $Y=0 $X2=4.56
+ $Y2=0
r90 42 61 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r91 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r92 39 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.4 $Y=0 $X2=3.235
+ $Y2=0
r93 39 41 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=3.4 $Y=0 $X2=3.6 $Y2=0
r94 38 60 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.97 $Y=0 $X2=4.135
+ $Y2=0
r95 38 41 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=3.97 $Y=0 $X2=3.6
+ $Y2=0
r96 36 55 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=0.24 $Y=0 $X2=2.16
+ $Y2=0
r97 35 36 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r98 33 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.1 $Y=0 $X2=2.265
+ $Y2=0
r99 33 35 121.348 $w=1.68e-07 $l=1.86e-06 $layer=LI1_cond $X=2.1 $Y=0 $X2=0.24
+ $Y2=0
r100 31 42 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r101 31 55 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.16
+ $Y2=0
r102 31 57 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r103 27 63 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.995 $Y=0.085
+ $X2=4.995 $Y2=0
r104 27 29 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=4.995 $Y=0.085
+ $X2=4.995 $Y2=0.36
r105 23 60 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.135 $Y=0.085
+ $X2=4.135 $Y2=0
r106 23 25 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=4.135 $Y=0.085
+ $X2=4.135 $Y2=0.36
r107 19 57 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.235 $Y=0.085
+ $X2=3.235 $Y2=0
r108 19 21 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=3.235 $Y=0.085
+ $X2=3.235 $Y2=0.36
r109 18 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.43 $Y=0 $X2=2.265
+ $Y2=0
r110 17 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.07 $Y=0 $X2=3.235
+ $Y2=0
r111 17 18 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=3.07 $Y=0 $X2=2.43
+ $Y2=0
r112 13 54 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.265 $Y=0.085
+ $X2=2.265 $Y2=0
r113 13 15 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.265 $Y=0.085
+ $X2=2.265 $Y2=0.36
r114 4 29 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=4.855
+ $Y=0.235 $X2=4.995 $Y2=0.36
r115 3 25 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=3.995
+ $Y=0.235 $X2=4.135 $Y2=0.36
r116 2 21 91 $w=1.7e-07 $l=2.13542e-07 $layer=licon1_NDIFF $count=2 $X=3.075
+ $Y=0.235 $X2=3.235 $Y2=0.36
r117 1 15 91 $w=1.7e-07 $l=2.7037e-07 $layer=licon1_NDIFF $count=2 $X=2.05
+ $Y=0.235 $X2=2.265 $Y2=0.36
.ends

