* File: sky130_fd_sc_lp__einvp_4.pxi.spice
* Created: Fri Aug 28 10:33:58 2020
* 
x_PM_SKY130_FD_SC_LP__EINVP_4%TE N_TE_c_106_n N_TE_M1016_g N_TE_M1004_g
+ N_TE_c_108_n N_TE_c_109_n N_TE_M1005_g N_TE_c_110_n N_TE_c_111_n N_TE_M1006_g
+ N_TE_c_112_n N_TE_c_113_n N_TE_M1014_g N_TE_c_114_n N_TE_c_115_n N_TE_M1017_g
+ N_TE_c_116_n N_TE_c_117_n N_TE_c_118_n N_TE_c_119_n N_TE_c_120_n N_TE_c_121_n
+ TE TE TE TE N_TE_c_122_n N_TE_c_123_n N_TE_c_124_n
+ PM_SKY130_FD_SC_LP__EINVP_4%TE
x_PM_SKY130_FD_SC_LP__EINVP_4%A_35_47# N_A_35_47#_M1016_s N_A_35_47#_M1004_s
+ N_A_35_47#_c_199_n N_A_35_47#_c_200_n N_A_35_47#_c_213_n N_A_35_47#_M1000_g
+ N_A_35_47#_c_201_n N_A_35_47#_c_215_n N_A_35_47#_M1007_g N_A_35_47#_c_202_n
+ N_A_35_47#_c_217_n N_A_35_47#_M1012_g N_A_35_47#_c_203_n N_A_35_47#_c_219_n
+ N_A_35_47#_M1015_g N_A_35_47#_c_204_n N_A_35_47#_c_205_n N_A_35_47#_c_206_n
+ N_A_35_47#_c_207_n N_A_35_47#_c_208_n N_A_35_47#_c_209_n N_A_35_47#_c_224_n
+ N_A_35_47#_c_225_n N_A_35_47#_c_210_n PM_SKY130_FD_SC_LP__EINVP_4%A_35_47#
x_PM_SKY130_FD_SC_LP__EINVP_4%A N_A_M1003_g N_A_M1001_g N_A_M1008_g N_A_M1002_g
+ N_A_c_291_n N_A_c_292_n N_A_M1011_g N_A_M1009_g N_A_M1013_g N_A_M1010_g
+ N_A_c_295_n A N_A_c_296_n PM_SKY130_FD_SC_LP__EINVP_4%A
x_PM_SKY130_FD_SC_LP__EINVP_4%VPWR N_VPWR_M1004_d N_VPWR_M1000_d N_VPWR_M1012_d
+ N_VPWR_c_381_n N_VPWR_c_382_n N_VPWR_c_383_n N_VPWR_c_384_n N_VPWR_c_385_n
+ N_VPWR_c_386_n N_VPWR_c_387_n VPWR N_VPWR_c_388_n N_VPWR_c_389_n
+ N_VPWR_c_380_n N_VPWR_c_391_n PM_SKY130_FD_SC_LP__EINVP_4%VPWR
x_PM_SKY130_FD_SC_LP__EINVP_4%A_301_367# N_A_301_367#_M1000_s
+ N_A_301_367#_M1007_s N_A_301_367#_M1015_s N_A_301_367#_M1002_d
+ N_A_301_367#_M1010_d N_A_301_367#_c_466_n N_A_301_367#_c_450_n
+ N_A_301_367#_c_451_n N_A_301_367#_c_497_n N_A_301_367#_c_452_n
+ N_A_301_367#_c_501_n N_A_301_367#_c_481_n N_A_301_367#_c_483_n
+ N_A_301_367#_c_484_n N_A_301_367#_c_453_n N_A_301_367#_c_454_n
+ N_A_301_367#_c_455_n N_A_301_367#_c_509_n
+ PM_SKY130_FD_SC_LP__EINVP_4%A_301_367#
x_PM_SKY130_FD_SC_LP__EINVP_4%Z N_Z_M1003_d N_Z_M1008_d N_Z_M1013_d N_Z_M1001_s
+ N_Z_M1009_s N_Z_c_523_n N_Z_c_524_n N_Z_c_525_n N_Z_c_539_n N_Z_c_542_n
+ N_Z_c_526_n N_Z_c_528_n N_Z_c_555_n N_Z_c_527_n N_Z_c_557_n Z Z N_Z_c_560_n
+ PM_SKY130_FD_SC_LP__EINVP_4%Z
x_PM_SKY130_FD_SC_LP__EINVP_4%VGND N_VGND_M1016_d N_VGND_M1006_d N_VGND_M1017_d
+ N_VGND_c_592_n N_VGND_c_593_n N_VGND_c_594_n N_VGND_c_595_n N_VGND_c_596_n
+ N_VGND_c_597_n N_VGND_c_598_n VGND N_VGND_c_599_n N_VGND_c_600_n
+ N_VGND_c_601_n N_VGND_c_602_n PM_SKY130_FD_SC_LP__EINVP_4%VGND
x_PM_SKY130_FD_SC_LP__EINVP_4%A_204_47# N_A_204_47#_M1005_s N_A_204_47#_M1014_s
+ N_A_204_47#_M1003_s N_A_204_47#_M1011_s N_A_204_47#_c_714_n
+ N_A_204_47#_c_667_n N_A_204_47#_c_671_n N_A_204_47#_c_718_n
+ N_A_204_47#_c_660_n N_A_204_47#_c_661_n N_A_204_47#_c_662_n
+ N_A_204_47#_c_663_n N_A_204_47#_c_688_n N_A_204_47#_c_664_n
+ N_A_204_47#_c_665_n N_A_204_47#_c_680_n N_A_204_47#_c_666_n
+ PM_SKY130_FD_SC_LP__EINVP_4%A_204_47#
cc_1 VNB N_TE_c_106_n 0.0192412f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=1.185
cc_2 VNB N_TE_M1004_g 0.0208454f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=2.465
cc_3 VNB N_TE_c_108_n 0.0140981f $X=-0.19 $Y=-0.245 $X2=0.87 $Y2=1.275
cc_4 VNB N_TE_c_109_n 0.0161884f $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=1.185
cc_5 VNB N_TE_c_110_n 0.0121815f $X=-0.19 $Y=-0.245 $X2=1.3 $Y2=1.275
cc_6 VNB N_TE_c_111_n 0.016004f $X=-0.19 $Y=-0.245 $X2=1.375 $Y2=1.185
cc_7 VNB N_TE_c_112_n 0.0109861f $X=-0.19 $Y=-0.245 $X2=1.73 $Y2=1.275
cc_8 VNB N_TE_c_113_n 0.0160063f $X=-0.19 $Y=-0.245 $X2=1.805 $Y2=1.185
cc_9 VNB N_TE_c_114_n 0.0103769f $X=-0.19 $Y=-0.245 $X2=2.16 $Y2=1.275
cc_10 VNB N_TE_c_115_n 0.0190343f $X=-0.19 $Y=-0.245 $X2=2.235 $Y2=1.185
cc_11 VNB N_TE_c_116_n 0.0294793f $X=-0.19 $Y=-0.245 $X2=2.875 $Y2=1.275
cc_12 VNB N_TE_c_117_n 0.0073341f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=1.275
cc_13 VNB N_TE_c_118_n 0.00657097f $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=1.275
cc_14 VNB N_TE_c_119_n 0.00542151f $X=-0.19 $Y=-0.245 $X2=1.375 $Y2=1.275
cc_15 VNB N_TE_c_120_n 0.00438817f $X=-0.19 $Y=-0.245 $X2=1.805 $Y2=1.275
cc_16 VNB N_TE_c_121_n 0.00438817f $X=-0.19 $Y=-0.245 $X2=2.235 $Y2=1.275
cc_17 VNB N_TE_c_122_n 0.0373228f $X=-0.19 $Y=-0.245 $X2=3.04 $Y2=1.17
cc_18 VNB N_TE_c_123_n 0.00762831f $X=-0.19 $Y=-0.245 $X2=3.04 $Y2=1.17
cc_19 VNB N_TE_c_124_n 0.0124019f $X=-0.19 $Y=-0.245 $X2=2.875 $Y2=1.32
cc_20 VNB N_A_35_47#_c_199_n 0.0106044f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_35_47#_c_200_n 0.00765429f $X=-0.19 $Y=-0.245 $X2=0.87 $Y2=1.275
cc_22 VNB N_A_35_47#_c_201_n 0.00692614f $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=0.655
cc_23 VNB N_A_35_47#_c_202_n 0.00699387f $X=-0.19 $Y=-0.245 $X2=1.375 $Y2=0.655
cc_24 VNB N_A_35_47#_c_203_n 0.0130275f $X=-0.19 $Y=-0.245 $X2=1.805 $Y2=0.655
cc_25 VNB N_A_35_47#_c_204_n 0.00381313f $X=-0.19 $Y=-0.245 $X2=2.875 $Y2=1.275
cc_26 VNB N_A_35_47#_c_205_n 0.00381313f $X=-0.19 $Y=-0.245 $X2=2.31 $Y2=1.275
cc_27 VNB N_A_35_47#_c_206_n 0.00381313f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=1.275
cc_28 VNB N_A_35_47#_c_207_n 0.0500299f $X=-0.19 $Y=-0.245 $X2=1.805 $Y2=1.275
cc_29 VNB N_A_35_47#_c_208_n 4.4709e-19 $X=-0.19 $Y=-0.245 $X2=2.555 $Y2=1.21
cc_30 VNB N_A_35_47#_c_209_n 0.020594f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_35_47#_c_210_n 0.0102039f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_M1003_g 0.0223995f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=0.655
cc_33 VNB N_A_M1008_g 0.0190492f $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=0.655
cc_34 VNB N_A_c_291_n 0.0167383f $X=-0.19 $Y=-0.245 $X2=1.375 $Y2=0.655
cc_35 VNB N_A_c_292_n 0.0373728f $X=-0.19 $Y=-0.245 $X2=1.73 $Y2=1.275
cc_36 VNB N_A_M1011_g 0.0190269f $X=-0.19 $Y=-0.245 $X2=1.805 $Y2=0.655
cc_37 VNB N_A_M1013_g 0.0231513f $X=-0.19 $Y=-0.245 $X2=2.31 $Y2=1.275
cc_38 VNB N_A_c_295_n 0.0328194f $X=-0.19 $Y=-0.245 $X2=2.075 $Y2=1.21
cc_39 VNB N_A_c_296_n 0.00726545f $X=-0.19 $Y=-0.245 $X2=3.04 $Y2=1.275
cc_40 VNB N_VPWR_c_380_n 0.243291f $X=-0.19 $Y=-0.245 $X2=2.16 $Y2=1.32
cc_41 VNB N_Z_c_523_n 0.00908751f $X=-0.19 $Y=-0.245 $X2=1.73 $Y2=1.275
cc_42 VNB N_Z_c_524_n 0.00321778f $X=-0.19 $Y=-0.245 $X2=1.805 $Y2=1.185
cc_43 VNB N_Z_c_525_n 0.00638395f $X=-0.19 $Y=-0.245 $X2=1.805 $Y2=0.655
cc_44 VNB N_Z_c_526_n 0.0139722f $X=-0.19 $Y=-0.245 $X2=2.875 $Y2=1.275
cc_45 VNB N_Z_c_527_n 0.0455377f $X=-0.19 $Y=-0.245 $X2=2.075 $Y2=1.21
cc_46 VNB N_VGND_c_592_n 0.00813315f $X=-0.19 $Y=-0.245 $X2=0.945 $Y2=0.655
cc_47 VNB N_VGND_c_593_n 3.15212e-19 $X=-0.19 $Y=-0.245 $X2=1.375 $Y2=0.655
cc_48 VNB N_VGND_c_594_n 0.00737078f $X=-0.19 $Y=-0.245 $X2=1.805 $Y2=1.185
cc_49 VNB N_VGND_c_595_n 0.0147711f $X=-0.19 $Y=-0.245 $X2=2.16 $Y2=1.275
cc_50 VNB N_VGND_c_596_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=1.88 $Y2=1.275
cc_51 VNB N_VGND_c_597_n 0.0122995f $X=-0.19 $Y=-0.245 $X2=2.235 $Y2=0.655
cc_52 VNB N_VGND_c_598_n 0.00510637f $X=-0.19 $Y=-0.245 $X2=2.235 $Y2=0.655
cc_53 VNB N_VGND_c_599_n 0.01848f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=1.275
cc_54 VNB N_VGND_c_600_n 0.0772449f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_601_n 0.310103f $X=-0.19 $Y=-0.245 $X2=3.04 $Y2=1.275
cc_56 VNB N_VGND_c_602_n 0.00500104f $X=-0.19 $Y=-0.245 $X2=1.68 $Y2=1.32
cc_57 VNB N_A_204_47#_c_660_n 0.0182856f $X=-0.19 $Y=-0.245 $X2=2.16 $Y2=1.275
cc_58 VNB N_A_204_47#_c_661_n 0.0108682f $X=-0.19 $Y=-0.245 $X2=2.235 $Y2=0.655
cc_59 VNB N_A_204_47#_c_662_n 0.0156097f $X=-0.19 $Y=-0.245 $X2=2.235 $Y2=0.655
cc_60 VNB N_A_204_47#_c_663_n 0.00617619f $X=-0.19 $Y=-0.245 $X2=2.875 $Y2=1.275
cc_61 VNB N_A_204_47#_c_664_n 0.00556228f $X=-0.19 $Y=-0.245 $X2=1.805 $Y2=1.275
cc_62 VNB N_A_204_47#_c_665_n 0.00229853f $X=-0.19 $Y=-0.245 $X2=2.555 $Y2=1.21
cc_63 VNB N_A_204_47#_c_666_n 0.0020718f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VPB N_TE_M1004_g 0.0269488f $X=-0.19 $Y=1.655 $X2=0.515 $Y2=2.465
cc_65 VPB N_A_35_47#_c_199_n 0.0104044f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_66 VPB N_A_35_47#_c_200_n 0.00422276f $X=-0.19 $Y=1.655 $X2=0.87 $Y2=1.275
cc_67 VPB N_A_35_47#_c_213_n 0.0185007f $X=-0.19 $Y=1.655 $X2=0.59 $Y2=1.275
cc_68 VPB N_A_35_47#_c_201_n 0.00418369f $X=-0.19 $Y=1.655 $X2=0.945 $Y2=0.655
cc_69 VPB N_A_35_47#_c_215_n 0.0153032f $X=-0.19 $Y=1.655 $X2=1.02 $Y2=1.275
cc_70 VPB N_A_35_47#_c_202_n 0.00418344f $X=-0.19 $Y=1.655 $X2=1.375 $Y2=0.655
cc_71 VPB N_A_35_47#_c_217_n 0.0153032f $X=-0.19 $Y=1.655 $X2=1.45 $Y2=1.275
cc_72 VPB N_A_35_47#_c_203_n 0.00739589f $X=-0.19 $Y=1.655 $X2=1.805 $Y2=0.655
cc_73 VPB N_A_35_47#_c_219_n 0.0177738f $X=-0.19 $Y=1.655 $X2=1.88 $Y2=1.275
cc_74 VPB N_A_35_47#_c_204_n 0.00111435f $X=-0.19 $Y=1.655 $X2=2.875 $Y2=1.275
cc_75 VPB N_A_35_47#_c_205_n 0.00111435f $X=-0.19 $Y=1.655 $X2=2.31 $Y2=1.275
cc_76 VPB N_A_35_47#_c_206_n 0.00111435f $X=-0.19 $Y=1.655 $X2=0.515 $Y2=1.275
cc_77 VPB N_A_35_47#_c_208_n 0.0566079f $X=-0.19 $Y=1.655 $X2=2.555 $Y2=1.21
cc_78 VPB N_A_35_47#_c_224_n 0.0113222f $X=-0.19 $Y=1.655 $X2=3.04 $Y2=1.17
cc_79 VPB N_A_35_47#_c_225_n 0.0530631f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_80 VPB N_A_M1001_g 0.0211884f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_81 VPB N_A_M1002_g 0.0192673f $X=-0.19 $Y=1.655 $X2=1.375 $Y2=1.185
cc_82 VPB N_A_c_291_n 0.00576413f $X=-0.19 $Y=1.655 $X2=1.375 $Y2=0.655
cc_83 VPB N_A_c_292_n 0.00863678f $X=-0.19 $Y=1.655 $X2=1.73 $Y2=1.275
cc_84 VPB N_A_M1009_g 0.0182523f $X=-0.19 $Y=1.655 $X2=2.235 $Y2=1.185
cc_85 VPB N_A_M1010_g 0.0249076f $X=-0.19 $Y=1.655 $X2=1.805 $Y2=1.275
cc_86 VPB N_A_c_295_n 0.00519541f $X=-0.19 $Y=1.655 $X2=2.075 $Y2=1.21
cc_87 VPB N_A_c_296_n 0.00652396f $X=-0.19 $Y=1.655 $X2=3.04 $Y2=1.275
cc_88 VPB N_VPWR_c_381_n 0.0260406f $X=-0.19 $Y=1.655 $X2=0.945 $Y2=0.655
cc_89 VPB N_VPWR_c_382_n 3.99129e-19 $X=-0.19 $Y=1.655 $X2=1.73 $Y2=1.275
cc_90 VPB N_VPWR_c_383_n 3.99129e-19 $X=-0.19 $Y=1.655 $X2=1.88 $Y2=1.275
cc_91 VPB N_VPWR_c_384_n 0.0287548f $X=-0.19 $Y=1.655 $X2=2.31 $Y2=1.275
cc_92 VPB N_VPWR_c_385_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0.515 $Y2=1.275
cc_93 VPB N_VPWR_c_386_n 0.0129398f $X=-0.19 $Y=1.655 $X2=1.375 $Y2=1.275
cc_94 VPB N_VPWR_c_387_n 0.00436868f $X=-0.19 $Y=1.655 $X2=1.805 $Y2=1.275
cc_95 VPB N_VPWR_c_388_n 0.01848f $X=-0.19 $Y=1.655 $X2=2.075 $Y2=1.21
cc_96 VPB N_VPWR_c_389_n 0.0630161f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_97 VPB N_VPWR_c_380_n 0.0723964f $X=-0.19 $Y=1.655 $X2=2.16 $Y2=1.32
cc_98 VPB N_VPWR_c_391_n 0.00564836f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_99 VPB N_A_301_367#_c_450_n 0.00298643f $X=-0.19 $Y=1.655 $X2=1.805 $Y2=0.655
cc_100 VPB N_A_301_367#_c_451_n 0.00238957f $X=-0.19 $Y=1.655 $X2=2.16 $Y2=1.275
cc_101 VPB N_A_301_367#_c_452_n 0.0142153f $X=-0.19 $Y=1.655 $X2=0.515 $Y2=1.275
cc_102 VPB N_A_301_367#_c_453_n 0.00746637f $X=-0.19 $Y=1.655 $X2=3.04 $Y2=1.17
cc_103 VPB N_A_301_367#_c_454_n 0.0443905f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_104 VPB N_A_301_367#_c_455_n 0.00151731f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_105 VPB N_Z_c_528_n 0.00139814f $X=-0.19 $Y=1.655 $X2=2.31 $Y2=1.275
cc_106 N_TE_c_110_n N_A_35_47#_c_199_n 0.0177451f $X=1.3 $Y=1.275 $X2=0 $Y2=0
cc_107 N_TE_c_124_n N_A_35_47#_c_199_n 0.0105471f $X=2.875 $Y=1.32 $X2=0 $Y2=0
cc_108 N_TE_M1004_g N_A_35_47#_c_200_n 0.0117796f $X=0.515 $Y=2.465 $X2=0 $Y2=0
cc_109 N_TE_c_118_n N_A_35_47#_c_200_n 0.0177451f $X=0.945 $Y=1.275 $X2=0 $Y2=0
cc_110 N_TE_c_112_n N_A_35_47#_c_201_n 0.0177451f $X=1.73 $Y=1.275 $X2=0 $Y2=0
cc_111 N_TE_c_114_n N_A_35_47#_c_202_n 0.0177451f $X=2.16 $Y=1.275 $X2=0 $Y2=0
cc_112 N_TE_c_116_n N_A_35_47#_c_203_n 0.0177451f $X=2.875 $Y=1.275 $X2=0 $Y2=0
cc_113 N_TE_c_123_n N_A_35_47#_c_203_n 0.00293036f $X=3.04 $Y=1.17 $X2=0 $Y2=0
cc_114 N_TE_c_119_n N_A_35_47#_c_204_n 0.0177451f $X=1.375 $Y=1.275 $X2=0 $Y2=0
cc_115 N_TE_c_120_n N_A_35_47#_c_205_n 0.0177451f $X=1.805 $Y=1.275 $X2=0 $Y2=0
cc_116 N_TE_c_121_n N_A_35_47#_c_206_n 0.0177451f $X=2.235 $Y=1.275 $X2=0 $Y2=0
cc_117 N_TE_c_106_n N_A_35_47#_c_207_n 0.0181448f $X=0.515 $Y=1.185 $X2=0 $Y2=0
cc_118 N_TE_M1004_g N_A_35_47#_c_208_n 0.00868539f $X=0.515 $Y=2.465 $X2=0 $Y2=0
cc_119 N_TE_M1004_g N_A_35_47#_c_209_n 0.0261704f $X=0.515 $Y=2.465 $X2=0 $Y2=0
cc_120 N_TE_c_108_n N_A_35_47#_c_209_n 0.016379f $X=0.87 $Y=1.275 $X2=0 $Y2=0
cc_121 N_TE_c_110_n N_A_35_47#_c_209_n 0.00337305f $X=1.3 $Y=1.275 $X2=0 $Y2=0
cc_122 N_TE_c_124_n N_A_35_47#_c_209_n 7.51347e-19 $X=2.875 $Y=1.32 $X2=0 $Y2=0
cc_123 N_TE_M1004_g N_A_35_47#_c_224_n 7.03757e-19 $X=0.515 $Y=2.465 $X2=0 $Y2=0
cc_124 N_TE_c_122_n N_A_M1003_g 0.00409019f $X=3.04 $Y=1.17 $X2=0 $Y2=0
cc_125 N_TE_c_123_n N_A_M1003_g 0.00186375f $X=3.04 $Y=1.17 $X2=0 $Y2=0
cc_126 N_TE_c_122_n N_A_c_292_n 4.28716e-19 $X=3.04 $Y=1.17 $X2=0 $Y2=0
cc_127 N_TE_c_123_n N_A_c_292_n 0.00240162f $X=3.04 $Y=1.17 $X2=0 $Y2=0
cc_128 N_TE_M1004_g N_VPWR_c_381_n 0.00799836f $X=0.515 $Y=2.465 $X2=0 $Y2=0
cc_129 N_TE_M1004_g N_VPWR_c_388_n 0.00585385f $X=0.515 $Y=2.465 $X2=0 $Y2=0
cc_130 N_TE_M1004_g N_VPWR_c_380_n 0.0127904f $X=0.515 $Y=2.465 $X2=0 $Y2=0
cc_131 N_TE_c_114_n N_A_301_367#_c_450_n 5.70092e-19 $X=2.16 $Y=1.275 $X2=0
+ $Y2=0
cc_132 N_TE_c_124_n N_A_301_367#_c_450_n 0.0315943f $X=2.875 $Y=1.32 $X2=0 $Y2=0
cc_133 N_TE_c_112_n N_A_301_367#_c_451_n 2.28252e-19 $X=1.73 $Y=1.275 $X2=0
+ $Y2=0
cc_134 N_TE_c_124_n N_A_301_367#_c_451_n 0.00983462f $X=2.875 $Y=1.32 $X2=0
+ $Y2=0
cc_135 N_TE_c_116_n N_A_301_367#_c_452_n 5.36783e-19 $X=2.875 $Y=1.275 $X2=0
+ $Y2=0
cc_136 N_TE_c_122_n N_A_301_367#_c_452_n 4.3032e-19 $X=3.04 $Y=1.17 $X2=0 $Y2=0
cc_137 N_TE_c_123_n N_A_301_367#_c_452_n 0.01796f $X=3.04 $Y=1.17 $X2=0 $Y2=0
cc_138 N_TE_c_124_n N_A_301_367#_c_452_n 0.0135969f $X=2.875 $Y=1.32 $X2=0 $Y2=0
cc_139 N_TE_c_116_n N_A_301_367#_c_455_n 3.97078e-19 $X=2.875 $Y=1.275 $X2=0
+ $Y2=0
cc_140 N_TE_c_124_n N_A_301_367#_c_455_n 0.0103848f $X=2.875 $Y=1.32 $X2=0 $Y2=0
cc_141 N_TE_c_122_n N_Z_c_523_n 0.00160514f $X=3.04 $Y=1.17 $X2=0 $Y2=0
cc_142 N_TE_c_123_n N_Z_c_523_n 0.00138814f $X=3.04 $Y=1.17 $X2=0 $Y2=0
cc_143 N_TE_c_122_n N_Z_c_525_n 7.91414e-19 $X=3.04 $Y=1.17 $X2=0 $Y2=0
cc_144 N_TE_c_123_n N_Z_c_525_n 0.0128361f $X=3.04 $Y=1.17 $X2=0 $Y2=0
cc_145 N_TE_c_106_n N_VGND_c_592_n 0.00424645f $X=0.515 $Y=1.185 $X2=0 $Y2=0
cc_146 N_TE_c_108_n N_VGND_c_592_n 0.00259854f $X=0.87 $Y=1.275 $X2=0 $Y2=0
cc_147 N_TE_c_109_n N_VGND_c_592_n 0.00349164f $X=0.945 $Y=1.185 $X2=0 $Y2=0
cc_148 N_TE_c_109_n N_VGND_c_593_n 5.90035e-19 $X=0.945 $Y=1.185 $X2=0 $Y2=0
cc_149 N_TE_c_111_n N_VGND_c_593_n 0.0107111f $X=1.375 $Y=1.185 $X2=0 $Y2=0
cc_150 N_TE_c_113_n N_VGND_c_593_n 0.0106305f $X=1.805 $Y=1.185 $X2=0 $Y2=0
cc_151 N_TE_c_115_n N_VGND_c_593_n 5.75816e-19 $X=2.235 $Y=1.185 $X2=0 $Y2=0
cc_152 N_TE_c_113_n N_VGND_c_594_n 5.34794e-19 $X=1.805 $Y=1.185 $X2=0 $Y2=0
cc_153 N_TE_c_115_n N_VGND_c_594_n 0.00863329f $X=2.235 $Y=1.185 $X2=0 $Y2=0
cc_154 N_TE_c_109_n N_VGND_c_595_n 0.00585385f $X=0.945 $Y=1.185 $X2=0 $Y2=0
cc_155 N_TE_c_111_n N_VGND_c_595_n 0.00486043f $X=1.375 $Y=1.185 $X2=0 $Y2=0
cc_156 N_TE_c_113_n N_VGND_c_597_n 0.00486043f $X=1.805 $Y=1.185 $X2=0 $Y2=0
cc_157 N_TE_c_115_n N_VGND_c_597_n 0.00364083f $X=2.235 $Y=1.185 $X2=0 $Y2=0
cc_158 N_TE_c_106_n N_VGND_c_599_n 0.00585385f $X=0.515 $Y=1.185 $X2=0 $Y2=0
cc_159 N_TE_c_106_n N_VGND_c_601_n 0.0114907f $X=0.515 $Y=1.185 $X2=0 $Y2=0
cc_160 N_TE_c_109_n N_VGND_c_601_n 0.0105224f $X=0.945 $Y=1.185 $X2=0 $Y2=0
cc_161 N_TE_c_111_n N_VGND_c_601_n 0.00824727f $X=1.375 $Y=1.185 $X2=0 $Y2=0
cc_162 N_TE_c_113_n N_VGND_c_601_n 0.00824727f $X=1.805 $Y=1.185 $X2=0 $Y2=0
cc_163 N_TE_c_115_n N_VGND_c_601_n 0.00430165f $X=2.235 $Y=1.185 $X2=0 $Y2=0
cc_164 N_TE_c_111_n N_A_204_47#_c_667_n 0.0128062f $X=1.375 $Y=1.185 $X2=0 $Y2=0
cc_165 N_TE_c_112_n N_A_204_47#_c_667_n 0.00211801f $X=1.73 $Y=1.275 $X2=0 $Y2=0
cc_166 N_TE_c_113_n N_A_204_47#_c_667_n 0.0121284f $X=1.805 $Y=1.185 $X2=0 $Y2=0
cc_167 N_TE_c_124_n N_A_204_47#_c_667_n 0.0230266f $X=2.875 $Y=1.32 $X2=0 $Y2=0
cc_168 N_TE_c_110_n N_A_204_47#_c_671_n 0.00246821f $X=1.3 $Y=1.275 $X2=0 $Y2=0
cc_169 N_TE_c_115_n N_A_204_47#_c_660_n 0.0168721f $X=2.235 $Y=1.185 $X2=0 $Y2=0
cc_170 N_TE_c_116_n N_A_204_47#_c_660_n 0.0112066f $X=2.875 $Y=1.275 $X2=0 $Y2=0
cc_171 N_TE_c_122_n N_A_204_47#_c_660_n 0.00911281f $X=3.04 $Y=1.17 $X2=0 $Y2=0
cc_172 N_TE_c_123_n N_A_204_47#_c_660_n 0.0266238f $X=3.04 $Y=1.17 $X2=0 $Y2=0
cc_173 N_TE_c_124_n N_A_204_47#_c_660_n 0.0479824f $X=2.875 $Y=1.32 $X2=0 $Y2=0
cc_174 N_TE_c_115_n N_A_204_47#_c_661_n 0.00341855f $X=2.235 $Y=1.185 $X2=0
+ $Y2=0
cc_175 N_TE_c_122_n N_A_204_47#_c_662_n 2.52092e-19 $X=3.04 $Y=1.17 $X2=0 $Y2=0
cc_176 N_TE_c_123_n N_A_204_47#_c_662_n 0.00149749f $X=3.04 $Y=1.17 $X2=0 $Y2=0
cc_177 N_TE_c_114_n N_A_204_47#_c_680_n 0.00213216f $X=2.16 $Y=1.275 $X2=0 $Y2=0
cc_178 N_TE_c_124_n N_A_204_47#_c_680_n 0.0141815f $X=2.875 $Y=1.32 $X2=0 $Y2=0
cc_179 N_A_35_47#_c_203_n N_A_M1001_g 0.00566965f $X=3.06 $Y=1.65 $X2=0 $Y2=0
cc_180 N_A_35_47#_c_203_n N_A_c_292_n 0.00220275f $X=3.06 $Y=1.65 $X2=0 $Y2=0
cc_181 N_A_35_47#_c_203_n N_A_c_296_n 0.00227535f $X=3.06 $Y=1.65 $X2=0 $Y2=0
cc_182 N_A_35_47#_c_208_n N_VPWR_c_381_n 0.00155436f $X=0.3 $Y=1.98 $X2=0 $Y2=0
cc_183 N_A_35_47#_c_209_n N_VPWR_c_381_n 0.0252284f $X=1.065 $Y=1.532 $X2=0
+ $Y2=0
cc_184 N_A_35_47#_c_224_n N_VPWR_c_381_n 0.0333256f $X=1.18 $Y=1.74 $X2=0 $Y2=0
cc_185 N_A_35_47#_c_225_n N_VPWR_c_381_n 0.00390561f $X=1.18 $Y=1.74 $X2=0 $Y2=0
cc_186 N_A_35_47#_c_213_n N_VPWR_c_382_n 0.0162094f $X=1.845 $Y=1.725 $X2=0
+ $Y2=0
cc_187 N_A_35_47#_c_215_n N_VPWR_c_382_n 0.0142791f $X=2.275 $Y=1.725 $X2=0
+ $Y2=0
cc_188 N_A_35_47#_c_217_n N_VPWR_c_382_n 7.27171e-19 $X=2.705 $Y=1.725 $X2=0
+ $Y2=0
cc_189 N_A_35_47#_c_215_n N_VPWR_c_383_n 7.24342e-19 $X=2.275 $Y=1.725 $X2=0
+ $Y2=0
cc_190 N_A_35_47#_c_217_n N_VPWR_c_383_n 0.0141279f $X=2.705 $Y=1.725 $X2=0
+ $Y2=0
cc_191 N_A_35_47#_c_219_n N_VPWR_c_383_n 0.0160983f $X=3.135 $Y=1.725 $X2=0
+ $Y2=0
cc_192 N_A_35_47#_c_213_n N_VPWR_c_384_n 0.00486043f $X=1.845 $Y=1.725 $X2=0
+ $Y2=0
cc_193 N_A_35_47#_c_215_n N_VPWR_c_386_n 0.00486043f $X=2.275 $Y=1.725 $X2=0
+ $Y2=0
cc_194 N_A_35_47#_c_217_n N_VPWR_c_386_n 0.00486043f $X=2.705 $Y=1.725 $X2=0
+ $Y2=0
cc_195 N_A_35_47#_c_208_n N_VPWR_c_388_n 0.0190529f $X=0.3 $Y=1.98 $X2=0 $Y2=0
cc_196 N_A_35_47#_c_219_n N_VPWR_c_389_n 0.00486043f $X=3.135 $Y=1.725 $X2=0
+ $Y2=0
cc_197 N_A_35_47#_M1004_s N_VPWR_c_380_n 0.00249946f $X=0.175 $Y=1.835 $X2=0
+ $Y2=0
cc_198 N_A_35_47#_c_213_n N_VPWR_c_380_n 0.00954696f $X=1.845 $Y=1.725 $X2=0
+ $Y2=0
cc_199 N_A_35_47#_c_215_n N_VPWR_c_380_n 0.00824727f $X=2.275 $Y=1.725 $X2=0
+ $Y2=0
cc_200 N_A_35_47#_c_217_n N_VPWR_c_380_n 0.00824727f $X=2.705 $Y=1.725 $X2=0
+ $Y2=0
cc_201 N_A_35_47#_c_219_n N_VPWR_c_380_n 0.00890141f $X=3.135 $Y=1.725 $X2=0
+ $Y2=0
cc_202 N_A_35_47#_c_208_n N_VPWR_c_380_n 0.0113912f $X=0.3 $Y=1.98 $X2=0 $Y2=0
cc_203 N_A_35_47#_c_224_n N_A_301_367#_c_466_n 0.0236661f $X=1.18 $Y=1.74 $X2=0
+ $Y2=0
cc_204 N_A_35_47#_c_225_n N_A_301_367#_c_466_n 0.00257381f $X=1.18 $Y=1.74 $X2=0
+ $Y2=0
cc_205 N_A_35_47#_c_213_n N_A_301_367#_c_450_n 0.0130909f $X=1.845 $Y=1.725
+ $X2=0 $Y2=0
cc_206 N_A_35_47#_c_201_n N_A_301_367#_c_450_n 0.00248966f $X=2.2 $Y=1.65 $X2=0
+ $Y2=0
cc_207 N_A_35_47#_c_215_n N_A_301_367#_c_450_n 0.0129953f $X=2.275 $Y=1.725
+ $X2=0 $Y2=0
cc_208 N_A_35_47#_c_199_n N_A_301_367#_c_451_n 0.00507731f $X=1.77 $Y=1.65 $X2=0
+ $Y2=0
cc_209 N_A_35_47#_c_224_n N_A_301_367#_c_451_n 0.0140196f $X=1.18 $Y=1.74 $X2=0
+ $Y2=0
cc_210 N_A_35_47#_c_225_n N_A_301_367#_c_451_n 0.00149685f $X=1.18 $Y=1.74 $X2=0
+ $Y2=0
cc_211 N_A_35_47#_c_217_n N_A_301_367#_c_452_n 0.0130517f $X=2.705 $Y=1.725
+ $X2=0 $Y2=0
cc_212 N_A_35_47#_c_203_n N_A_301_367#_c_452_n 0.00250337f $X=3.06 $Y=1.65 $X2=0
+ $Y2=0
cc_213 N_A_35_47#_c_219_n N_A_301_367#_c_452_n 0.0134148f $X=3.135 $Y=1.725
+ $X2=0 $Y2=0
cc_214 N_A_35_47#_c_202_n N_A_301_367#_c_455_n 0.00269641f $X=2.63 $Y=1.65 $X2=0
+ $Y2=0
cc_215 N_A_35_47#_c_207_n N_VGND_c_592_n 0.0031603f $X=0.3 $Y=0.42 $X2=0 $Y2=0
cc_216 N_A_35_47#_c_209_n N_VGND_c_592_n 0.014759f $X=1.065 $Y=1.532 $X2=0 $Y2=0
cc_217 N_A_35_47#_c_207_n N_VGND_c_599_n 0.0190529f $X=0.3 $Y=0.42 $X2=0 $Y2=0
cc_218 N_A_35_47#_M1016_s N_VGND_c_601_n 0.00249946f $X=0.175 $Y=0.235 $X2=0
+ $Y2=0
cc_219 N_A_35_47#_c_207_n N_VGND_c_601_n 0.0113912f $X=0.3 $Y=0.42 $X2=0 $Y2=0
cc_220 N_A_35_47#_c_199_n N_A_204_47#_c_667_n 9.70834e-19 $X=1.77 $Y=1.65 $X2=0
+ $Y2=0
cc_221 N_A_35_47#_c_209_n N_A_204_47#_c_667_n 0.00317335f $X=1.065 $Y=1.532
+ $X2=0 $Y2=0
cc_222 N_A_35_47#_c_200_n N_A_204_47#_c_671_n 2.71826e-19 $X=1.345 $Y=1.65 $X2=0
+ $Y2=0
cc_223 N_A_35_47#_c_209_n N_A_204_47#_c_671_n 0.00917453f $X=1.065 $Y=1.532
+ $X2=0 $Y2=0
cc_224 N_A_M1001_g N_VPWR_c_389_n 0.00357877f $X=3.915 $Y=2.465 $X2=0 $Y2=0
cc_225 N_A_M1002_g N_VPWR_c_389_n 0.00357877f $X=4.345 $Y=2.465 $X2=0 $Y2=0
cc_226 N_A_M1009_g N_VPWR_c_389_n 0.00357877f $X=4.855 $Y=2.465 $X2=0 $Y2=0
cc_227 N_A_M1010_g N_VPWR_c_389_n 0.00357877f $X=5.285 $Y=2.465 $X2=0 $Y2=0
cc_228 N_A_M1001_g N_VPWR_c_380_n 0.00600534f $X=3.915 $Y=2.465 $X2=0 $Y2=0
cc_229 N_A_M1002_g N_VPWR_c_380_n 0.00554494f $X=4.345 $Y=2.465 $X2=0 $Y2=0
cc_230 N_A_M1009_g N_VPWR_c_380_n 0.00554494f $X=4.855 $Y=2.465 $X2=0 $Y2=0
cc_231 N_A_M1010_g N_VPWR_c_380_n 0.00628381f $X=5.285 $Y=2.465 $X2=0 $Y2=0
cc_232 N_A_M1001_g N_A_301_367#_c_452_n 0.00415707f $X=3.915 $Y=2.465 $X2=0
+ $Y2=0
cc_233 N_A_c_292_n N_A_301_367#_c_452_n 5.56121e-19 $X=4.42 $Y=1.51 $X2=0 $Y2=0
cc_234 N_A_c_296_n N_A_301_367#_c_452_n 0.00725484f $X=4.21 $Y=1.51 $X2=0 $Y2=0
cc_235 N_A_M1001_g N_A_301_367#_c_481_n 0.0115031f $X=3.915 $Y=2.465 $X2=0 $Y2=0
cc_236 N_A_M1002_g N_A_301_367#_c_481_n 0.012237f $X=4.345 $Y=2.465 $X2=0 $Y2=0
cc_237 N_A_c_291_n N_A_301_367#_c_483_n 5.55133e-19 $X=4.78 $Y=1.51 $X2=0 $Y2=0
cc_238 N_A_M1009_g N_A_301_367#_c_484_n 0.012237f $X=4.855 $Y=2.465 $X2=0 $Y2=0
cc_239 N_A_M1010_g N_A_301_367#_c_484_n 0.0118089f $X=5.285 $Y=2.465 $X2=0 $Y2=0
cc_240 N_A_M1010_g N_A_301_367#_c_454_n 0.00339022f $X=5.285 $Y=2.465 $X2=0
+ $Y2=0
cc_241 N_A_M1003_g N_Z_c_524_n 0.0132611f $X=3.915 $Y=0.765 $X2=0 $Y2=0
cc_242 N_A_M1008_g N_Z_c_524_n 0.0134431f $X=4.345 $Y=0.765 $X2=0 $Y2=0
cc_243 N_A_c_292_n N_Z_c_524_n 0.00381774f $X=4.42 $Y=1.51 $X2=0 $Y2=0
cc_244 N_A_c_296_n N_Z_c_524_n 0.0433001f $X=4.21 $Y=1.51 $X2=0 $Y2=0
cc_245 N_A_c_292_n N_Z_c_525_n 0.00204754f $X=4.42 $Y=1.51 $X2=0 $Y2=0
cc_246 N_A_c_296_n N_Z_c_525_n 0.00671397f $X=4.21 $Y=1.51 $X2=0 $Y2=0
cc_247 N_A_M1002_g N_Z_c_539_n 0.0140951f $X=4.345 $Y=2.465 $X2=0 $Y2=0
cc_248 N_A_c_291_n N_Z_c_539_n 8.63213e-19 $X=4.78 $Y=1.51 $X2=0 $Y2=0
cc_249 N_A_c_296_n N_Z_c_539_n 0.00766292f $X=4.21 $Y=1.51 $X2=0 $Y2=0
cc_250 N_A_M1011_g N_Z_c_542_n 0.00460795f $X=4.855 $Y=0.765 $X2=0 $Y2=0
cc_251 N_A_M1008_g N_Z_c_526_n 0.00220165f $X=4.345 $Y=0.765 $X2=0 $Y2=0
cc_252 N_A_c_291_n N_Z_c_526_n 0.0152035f $X=4.78 $Y=1.51 $X2=0 $Y2=0
cc_253 N_A_M1011_g N_Z_c_526_n 0.00548318f $X=4.855 $Y=0.765 $X2=0 $Y2=0
cc_254 N_A_M1013_g N_Z_c_526_n 4.1391e-19 $X=5.285 $Y=0.765 $X2=0 $Y2=0
cc_255 N_A_c_295_n N_Z_c_526_n 0.0344631f $X=5.285 $Y=1.51 $X2=0 $Y2=0
cc_256 N_A_c_296_n N_Z_c_526_n 0.0109077f $X=4.21 $Y=1.51 $X2=0 $Y2=0
cc_257 N_A_M1002_g N_Z_c_528_n 0.00560779f $X=4.345 $Y=2.465 $X2=0 $Y2=0
cc_258 N_A_c_291_n N_Z_c_528_n 0.00745563f $X=4.78 $Y=1.51 $X2=0 $Y2=0
cc_259 N_A_M1009_g N_Z_c_528_n 0.00877388f $X=4.855 $Y=2.465 $X2=0 $Y2=0
cc_260 N_A_M1010_g N_Z_c_528_n 0.0100889f $X=5.285 $Y=2.465 $X2=0 $Y2=0
cc_261 N_A_c_295_n N_Z_c_528_n 0.0127855f $X=5.285 $Y=1.51 $X2=0 $Y2=0
cc_262 N_A_c_296_n N_Z_c_528_n 0.0165711f $X=4.21 $Y=1.51 $X2=0 $Y2=0
cc_263 N_A_M1010_g N_Z_c_555_n 0.00745759f $X=5.285 $Y=2.465 $X2=0 $Y2=0
cc_264 N_A_M1013_g N_Z_c_527_n 0.00984797f $X=5.285 $Y=0.765 $X2=0 $Y2=0
cc_265 N_A_M1009_g N_Z_c_557_n 0.012618f $X=4.855 $Y=2.465 $X2=0 $Y2=0
cc_266 N_A_M1010_g N_Z_c_557_n 0.00170116f $X=5.285 $Y=2.465 $X2=0 $Y2=0
cc_267 N_A_M1001_g Z 0.00804424f $X=3.915 $Y=2.465 $X2=0 $Y2=0
cc_268 N_A_M1001_g N_Z_c_560_n 0.00216601f $X=3.915 $Y=2.465 $X2=0 $Y2=0
cc_269 N_A_c_292_n N_Z_c_560_n 6.52992e-19 $X=4.42 $Y=1.51 $X2=0 $Y2=0
cc_270 N_A_c_296_n N_Z_c_560_n 0.0208725f $X=4.21 $Y=1.51 $X2=0 $Y2=0
cc_271 N_A_M1003_g N_VGND_c_600_n 0.00292999f $X=3.915 $Y=0.765 $X2=0 $Y2=0
cc_272 N_A_M1008_g N_VGND_c_600_n 0.00292999f $X=4.345 $Y=0.765 $X2=0 $Y2=0
cc_273 N_A_M1011_g N_VGND_c_600_n 0.00293025f $X=4.855 $Y=0.765 $X2=0 $Y2=0
cc_274 N_A_M1013_g N_VGND_c_600_n 0.00482246f $X=5.285 $Y=0.765 $X2=0 $Y2=0
cc_275 N_A_M1003_g N_VGND_c_601_n 0.0042879f $X=3.915 $Y=0.765 $X2=0 $Y2=0
cc_276 N_A_M1008_g N_VGND_c_601_n 0.00403268f $X=4.345 $Y=0.765 $X2=0 $Y2=0
cc_277 N_A_M1011_g N_VGND_c_601_n 0.00403272f $X=4.855 $Y=0.765 $X2=0 $Y2=0
cc_278 N_A_M1013_g N_VGND_c_601_n 0.00976044f $X=5.285 $Y=0.765 $X2=0 $Y2=0
cc_279 N_A_M1003_g N_A_204_47#_c_661_n 0.0040552f $X=3.915 $Y=0.765 $X2=0 $Y2=0
cc_280 N_A_M1003_g N_A_204_47#_c_662_n 0.0103134f $X=3.915 $Y=0.765 $X2=0 $Y2=0
cc_281 N_A_M1003_g N_A_204_47#_c_688_n 0.0108409f $X=3.915 $Y=0.765 $X2=0 $Y2=0
cc_282 N_A_M1008_g N_A_204_47#_c_688_n 0.00680334f $X=4.345 $Y=0.765 $X2=0 $Y2=0
cc_283 N_A_M1011_g N_A_204_47#_c_688_n 3.0466e-19 $X=4.855 $Y=0.765 $X2=0 $Y2=0
cc_284 N_A_M1008_g N_A_204_47#_c_664_n 0.00871648f $X=4.345 $Y=0.765 $X2=0 $Y2=0
cc_285 N_A_M1011_g N_A_204_47#_c_664_n 0.0126895f $X=4.855 $Y=0.765 $X2=0 $Y2=0
cc_286 N_A_M1013_g N_A_204_47#_c_664_n 0.00216665f $X=5.285 $Y=0.765 $X2=0 $Y2=0
cc_287 N_A_M1011_g N_A_204_47#_c_665_n 0.00105493f $X=4.855 $Y=0.765 $X2=0 $Y2=0
cc_288 N_A_M1013_g N_A_204_47#_c_665_n 0.00110088f $X=5.285 $Y=0.765 $X2=0 $Y2=0
cc_289 N_A_c_295_n N_A_204_47#_c_665_n 0.0024431f $X=5.285 $Y=1.51 $X2=0 $Y2=0
cc_290 N_A_M1003_g N_A_204_47#_c_666_n 0.00148464f $X=3.915 $Y=0.765 $X2=0 $Y2=0
cc_291 N_A_M1008_g N_A_204_47#_c_666_n 0.00148464f $X=4.345 $Y=0.765 $X2=0 $Y2=0
cc_292 N_VPWR_c_380_n N_A_301_367#_M1000_s 0.00409968f $X=5.52 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_293 N_VPWR_c_380_n N_A_301_367#_M1007_s 0.00536646f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_294 N_VPWR_c_380_n N_A_301_367#_M1015_s 0.00667163f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_295 N_VPWR_c_380_n N_A_301_367#_M1002_d 0.00287894f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_296 N_VPWR_c_380_n N_A_301_367#_M1010_d 0.0021516f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_297 N_VPWR_c_381_n N_A_301_367#_c_466_n 0.0256071f $X=0.73 $Y=1.98 $X2=0
+ $Y2=0
cc_298 N_VPWR_c_384_n N_A_301_367#_c_466_n 0.0142419f $X=1.895 $Y=3.33 $X2=0
+ $Y2=0
cc_299 N_VPWR_c_380_n N_A_301_367#_c_466_n 0.00808656f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_300 N_VPWR_M1000_d N_A_301_367#_c_450_n 0.00176461f $X=1.92 $Y=1.835 $X2=0
+ $Y2=0
cc_301 N_VPWR_c_382_n N_A_301_367#_c_450_n 0.0170777f $X=2.06 $Y=2.18 $X2=0
+ $Y2=0
cc_302 N_VPWR_c_386_n N_A_301_367#_c_497_n 0.0124525f $X=2.755 $Y=3.33 $X2=0
+ $Y2=0
cc_303 N_VPWR_c_380_n N_A_301_367#_c_497_n 0.00730901f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_304 N_VPWR_M1012_d N_A_301_367#_c_452_n 0.00180746f $X=2.78 $Y=1.835 $X2=0
+ $Y2=0
cc_305 N_VPWR_c_383_n N_A_301_367#_c_452_n 0.0163514f $X=2.92 $Y=2.19 $X2=0
+ $Y2=0
cc_306 N_VPWR_c_389_n N_A_301_367#_c_501_n 0.0371328f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_307 N_VPWR_c_380_n N_A_301_367#_c_501_n 0.020994f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_308 N_VPWR_c_389_n N_A_301_367#_c_481_n 0.035059f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_309 N_VPWR_c_380_n N_A_301_367#_c_481_n 0.0225481f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_310 N_VPWR_c_389_n N_A_301_367#_c_484_n 0.0347063f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_311 N_VPWR_c_380_n N_A_301_367#_c_484_n 0.0221721f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_312 N_VPWR_c_389_n N_A_301_367#_c_453_n 0.0182731f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_313 N_VPWR_c_380_n N_A_301_367#_c_453_n 0.0104917f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_314 N_VPWR_c_389_n N_A_301_367#_c_509_n 0.0202773f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_315 N_VPWR_c_380_n N_A_301_367#_c_509_n 0.0128296f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_316 N_VPWR_c_380_n N_Z_M1001_s 0.00225186f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_317 N_VPWR_c_380_n N_Z_M1009_s 0.00225186f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_318 N_A_301_367#_c_481_n N_Z_M1001_s 0.00332344f $X=4.435 $Y=2.99 $X2=0 $Y2=0
cc_319 N_A_301_367#_c_484_n N_Z_M1009_s 0.00332344f $X=5.395 $Y=2.99 $X2=0 $Y2=0
cc_320 N_A_301_367#_c_452_n N_Z_c_525_n 0.00928287f $X=3.255 $Y=1.84 $X2=0 $Y2=0
cc_321 N_A_301_367#_M1002_d N_Z_c_539_n 0.00186122f $X=4.42 $Y=1.835 $X2=0 $Y2=0
cc_322 N_A_301_367#_c_483_n N_Z_c_539_n 0.0054959f $X=4.6 $Y=2.425 $X2=0 $Y2=0
cc_323 N_A_301_367#_c_454_n N_Z_c_526_n 0.0186268f $X=5.5 $Y=1.98 $X2=0 $Y2=0
cc_324 N_A_301_367#_M1002_d N_Z_c_528_n 0.00112096f $X=4.42 $Y=1.835 $X2=0 $Y2=0
cc_325 N_A_301_367#_c_454_n N_Z_c_528_n 0.00512509f $X=5.5 $Y=1.98 $X2=0 $Y2=0
cc_326 N_A_301_367#_c_484_n N_Z_c_555_n 0.0135951f $X=5.395 $Y=2.99 $X2=0 $Y2=0
cc_327 N_A_301_367#_M1002_d N_Z_c_557_n 0.00195872f $X=4.42 $Y=1.835 $X2=0 $Y2=0
cc_328 N_A_301_367#_c_483_n N_Z_c_557_n 0.0160037f $X=4.6 $Y=2.425 $X2=0 $Y2=0
cc_329 N_A_301_367#_c_481_n Z 0.0143076f $X=4.435 $Y=2.99 $X2=0 $Y2=0
cc_330 N_Z_c_527_n N_VGND_c_600_n 0.0147756f $X=5.5 $Y=0.49 $X2=0 $Y2=0
cc_331 N_Z_c_527_n N_VGND_c_601_n 0.0111688f $X=5.5 $Y=0.49 $X2=0 $Y2=0
cc_332 N_Z_c_524_n N_A_204_47#_M1003_s 0.00184993f $X=4.465 $Y=1.17 $X2=0 $Y2=0
cc_333 N_Z_c_523_n N_A_204_47#_c_660_n 0.0110264f $X=3.62 $Y=0.7 $X2=0 $Y2=0
cc_334 N_Z_c_523_n N_A_204_47#_c_661_n 0.00734006f $X=3.62 $Y=0.7 $X2=0 $Y2=0
cc_335 N_Z_M1003_d N_A_204_47#_c_662_n 0.00387431f $X=3.495 $Y=0.345 $X2=0 $Y2=0
cc_336 N_Z_c_523_n N_A_204_47#_c_662_n 0.0249684f $X=3.62 $Y=0.7 $X2=0 $Y2=0
cc_337 N_Z_c_524_n N_A_204_47#_c_662_n 0.00275981f $X=4.465 $Y=1.17 $X2=0 $Y2=0
cc_338 N_Z_c_524_n N_A_204_47#_c_688_n 0.0155976f $X=4.465 $Y=1.17 $X2=0 $Y2=0
cc_339 N_Z_M1008_d N_A_204_47#_c_664_n 0.00267852f $X=4.42 $Y=0.345 $X2=0 $Y2=0
cc_340 N_Z_c_524_n N_A_204_47#_c_664_n 0.00275981f $X=4.465 $Y=1.17 $X2=0 $Y2=0
cc_341 N_Z_c_542_n N_A_204_47#_c_664_n 0.0187566f $X=4.63 $Y=0.7 $X2=0 $Y2=0
cc_342 N_Z_c_527_n N_A_204_47#_c_664_n 0.00166817f $X=5.5 $Y=0.49 $X2=0 $Y2=0
cc_343 N_Z_c_526_n N_A_204_47#_c_665_n 0.0269525f $X=4.885 $Y=1.555 $X2=0 $Y2=0
cc_344 N_Z_c_527_n N_A_204_47#_c_665_n 0.00233156f $X=5.5 $Y=0.49 $X2=0 $Y2=0
cc_345 N_VGND_c_601_n N_A_204_47#_M1005_s 0.0041489f $X=5.52 $Y=0 $X2=-0.19
+ $Y2=-0.245
cc_346 N_VGND_c_601_n N_A_204_47#_M1014_s 0.00400904f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_347 N_VGND_c_595_n N_A_204_47#_c_714_n 0.0136943f $X=1.425 $Y=0 $X2=0 $Y2=0
cc_348 N_VGND_c_601_n N_A_204_47#_c_714_n 0.00866972f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_349 N_VGND_M1006_d N_A_204_47#_c_667_n 0.00345033f $X=1.45 $Y=0.235 $X2=0
+ $Y2=0
cc_350 N_VGND_c_593_n N_A_204_47#_c_667_n 0.0170777f $X=1.59 $Y=0.58 $X2=0 $Y2=0
cc_351 N_VGND_c_597_n N_A_204_47#_c_718_n 0.0124525f $X=2.285 $Y=0 $X2=0 $Y2=0
cc_352 N_VGND_c_601_n N_A_204_47#_c_718_n 0.00730901f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_353 N_VGND_M1017_d N_A_204_47#_c_660_n 0.00535668f $X=2.31 $Y=0.235 $X2=0
+ $Y2=0
cc_354 N_VGND_c_594_n N_A_204_47#_c_660_n 0.0220323f $X=2.45 $Y=0.44 $X2=0 $Y2=0
cc_355 N_VGND_c_597_n N_A_204_47#_c_660_n 0.0020749f $X=2.285 $Y=0 $X2=0 $Y2=0
cc_356 N_VGND_c_600_n N_A_204_47#_c_660_n 0.00348829f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_357 N_VGND_c_601_n N_A_204_47#_c_660_n 0.0114178f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_358 N_VGND_c_594_n N_A_204_47#_c_661_n 0.00821649f $X=2.45 $Y=0.44 $X2=0
+ $Y2=0
cc_359 N_VGND_c_600_n N_A_204_47#_c_662_n 0.046582f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_360 N_VGND_c_601_n N_A_204_47#_c_662_n 0.0283842f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_361 N_VGND_c_594_n N_A_204_47#_c_663_n 0.0123491f $X=2.45 $Y=0.44 $X2=0 $Y2=0
cc_362 N_VGND_c_600_n N_A_204_47#_c_663_n 0.023463f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_363 N_VGND_c_601_n N_A_204_47#_c_663_n 0.0135145f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_364 N_VGND_c_600_n N_A_204_47#_c_664_n 0.0552933f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_365 N_VGND_c_601_n N_A_204_47#_c_664_n 0.0326727f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_366 N_VGND_c_600_n N_A_204_47#_c_666_n 0.0219516f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_367 N_VGND_c_601_n N_A_204_47#_c_666_n 0.0125121f $X=5.52 $Y=0 $X2=0 $Y2=0
