* File: sky130_fd_sc_lp__o2bb2ai_4.pex.spice
* Created: Wed Sep  2 10:22:24 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O2BB2AI_4%B1 3 7 11 15 19 23 27 31 33 38 42 43 44 45
+ 46 47 64 67 68 71
c123 47 0 1.33268e-19 $X=3.6 $Y=2.035
c124 42 0 2.41113e-20 $X=1.2 $Y=2.035
c125 38 0 1.7747e-19 $X=1.235 $Y=1.645
c126 31 0 1.08037e-19 $X=3.625 $Y=2.465
c127 27 0 1.8603e-19 $X=3.605 $Y=0.745
r128 67 70 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.645 $Y=1.51
+ $X2=3.645 $Y2=1.675
r129 67 69 54.9546 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=3.645 $Y=1.51
+ $X2=3.645 $Y2=1.295
r130 67 68 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.645
+ $Y=1.51 $X2=3.645 $Y2=1.51
r131 63 64 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=1.375 $Y=1.51
+ $X2=1.445 $Y2=1.51
r132 60 61 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=0.945 $Y=1.51
+ $X2=1.015 $Y2=1.51
r133 56 58 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=0.515 $Y=1.51
+ $X2=0.585 $Y2=1.51
r134 47 71 4.92601 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=3.645 $Y=2.04
+ $X2=3.48 $Y2=2.04
r135 47 68 11.9092 $w=4.98e-07 $l=4.4e-07 $layer=LI1_cond $X=3.645 $Y=1.95
+ $X2=3.645 $Y2=1.51
r136 46 71 22.1818 $w=1.78e-07 $l=3.6e-07 $layer=LI1_cond $X=3.12 $Y=2.04
+ $X2=3.48 $Y2=2.04
r137 45 46 29.5758 $w=1.78e-07 $l=4.8e-07 $layer=LI1_cond $X=2.64 $Y=2.04
+ $X2=3.12 $Y2=2.04
r138 44 45 29.5758 $w=1.78e-07 $l=4.8e-07 $layer=LI1_cond $X=2.16 $Y=2.04
+ $X2=2.64 $Y2=2.04
r139 43 44 29.5758 $w=1.78e-07 $l=4.8e-07 $layer=LI1_cond $X=1.68 $Y=2.04
+ $X2=2.16 $Y2=2.04
r140 43 72 16.3283 $w=1.78e-07 $l=2.65e-07 $layer=LI1_cond $X=1.68 $Y=2.04
+ $X2=1.415 $Y2=2.04
r141 42 72 5.2341 $w=1.8e-07 $l=1.8e-07 $layer=LI1_cond $X=1.235 $Y=2.04
+ $X2=1.415 $Y2=2.04
r142 41 63 21.8577 $w=3.3e-07 $l=1.25e-07 $layer=POLY_cond $X=1.25 $Y=1.51
+ $X2=1.375 $Y2=1.51
r143 41 61 41.0924 $w=3.3e-07 $l=2.35e-07 $layer=POLY_cond $X=1.25 $Y=1.51
+ $X2=1.015 $Y2=1.51
r144 40 41 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.25
+ $Y=1.51 $X2=1.25 $Y2=1.51
r145 38 42 7.66235 $w=5.28e-07 $l=3.05e-07 $layer=LI1_cond $X=1.235 $Y=1.645
+ $X2=1.235 $Y2=1.95
r146 38 40 2.78647 $w=3.6e-07 $l=1.1e-07 $layer=LI1_cond $X=1.235 $Y=1.645
+ $X2=1.235 $Y2=1.535
r147 36 60 6.12014 $w=3.3e-07 $l=3.5e-08 $layer=POLY_cond $X=0.91 $Y=1.51
+ $X2=0.945 $Y2=1.51
r148 36 58 56.8299 $w=3.3e-07 $l=3.25e-07 $layer=POLY_cond $X=0.91 $Y=1.51
+ $X2=0.585 $Y2=1.51
r149 35 36 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.91
+ $Y=1.51 $X2=0.91 $Y2=1.51
r150 33 40 4.55968 $w=2.2e-07 $l=1.8e-07 $layer=LI1_cond $X=1.055 $Y=1.535
+ $X2=1.235 $Y2=1.535
r151 33 35 7.59565 $w=2.18e-07 $l=1.45e-07 $layer=LI1_cond $X=1.055 $Y=1.535
+ $X2=0.91 $Y2=1.535
r152 31 70 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.625 $Y=2.465
+ $X2=3.625 $Y2=1.675
r153 27 69 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=3.605 $Y=0.745
+ $X2=3.605 $Y2=1.295
r154 21 64 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.445 $Y=1.675
+ $X2=1.445 $Y2=1.51
r155 21 23 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.445 $Y=1.675
+ $X2=1.445 $Y2=2.465
r156 17 63 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.375 $Y=1.345
+ $X2=1.375 $Y2=1.51
r157 17 19 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=1.375 $Y=1.345
+ $X2=1.375 $Y2=0.745
r158 13 61 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.015 $Y=1.675
+ $X2=1.015 $Y2=1.51
r159 13 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.015 $Y=1.675
+ $X2=1.015 $Y2=2.465
r160 9 60 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.945 $Y=1.345
+ $X2=0.945 $Y2=1.51
r161 9 11 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=0.945 $Y=1.345
+ $X2=0.945 $Y2=0.745
r162 5 58 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.585 $Y=1.675
+ $X2=0.585 $Y2=1.51
r163 5 7 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=0.585 $Y=1.675
+ $X2=0.585 $Y2=2.465
r164 1 56 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.515 $Y=1.345
+ $X2=0.515 $Y2=1.51
r165 1 3 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=0.515 $Y=1.345 $X2=0.515
+ $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_LP__O2BB2AI_4%B2 3 7 11 15 19 23 27 31 33 34 35 36 60
c83 60 0 2.01581e-19 $X=3.195 $Y=1.51
c84 36 0 1.08037e-19 $X=3.12 $Y=1.665
c85 27 0 6.61592e-20 $X=3.095 $Y=0.745
r86 59 60 17.4861 $w=3.3e-07 $l=1e-07 $layer=POLY_cond $X=3.095 $Y=1.51
+ $X2=3.195 $Y2=1.51
r87 57 59 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=2.915 $Y=1.51
+ $X2=3.095 $Y2=1.51
r88 57 58 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.915
+ $Y=1.51 $X2=2.915 $Y2=1.51
r89 55 57 26.2292 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=2.765 $Y=1.51
+ $X2=2.915 $Y2=1.51
r90 54 55 17.4861 $w=3.3e-07 $l=1e-07 $layer=POLY_cond $X=2.665 $Y=1.51
+ $X2=2.765 $Y2=1.51
r91 52 54 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=2.575 $Y=1.51
+ $X2=2.665 $Y2=1.51
r92 52 53 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.575
+ $Y=1.51 $X2=2.575 $Y2=1.51
r93 50 52 41.9667 $w=3.3e-07 $l=2.4e-07 $layer=POLY_cond $X=2.335 $Y=1.51
+ $X2=2.575 $Y2=1.51
r94 49 53 11.0375 $w=3.53e-07 $l=3.4e-07 $layer=LI1_cond $X=2.235 $Y=1.602
+ $X2=2.575 $Y2=1.602
r95 48 50 17.4861 $w=3.3e-07 $l=1e-07 $layer=POLY_cond $X=2.235 $Y=1.51
+ $X2=2.335 $Y2=1.51
r96 48 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.235
+ $Y=1.51 $X2=2.235 $Y2=1.51
r97 46 48 57.7042 $w=3.3e-07 $l=3.3e-07 $layer=POLY_cond $X=1.905 $Y=1.51
+ $X2=2.235 $Y2=1.51
r98 44 46 1.74861 $w=3.3e-07 $l=1e-08 $layer=POLY_cond $X=1.895 $Y=1.51
+ $X2=1.905 $Y2=1.51
r99 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.895
+ $Y=1.51 $X2=1.895 $Y2=1.51
r100 41 44 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=1.805 $Y=1.51
+ $X2=1.895 $Y2=1.51
r101 36 58 6.65495 $w=3.53e-07 $l=2.05e-07 $layer=LI1_cond $X=3.12 $Y=1.602
+ $X2=2.915 $Y2=1.602
r102 35 58 8.92738 $w=3.53e-07 $l=2.75e-07 $layer=LI1_cond $X=2.64 $Y=1.602
+ $X2=2.915 $Y2=1.602
r103 35 53 2.11011 $w=3.53e-07 $l=6.5e-08 $layer=LI1_cond $X=2.64 $Y=1.602
+ $X2=2.575 $Y2=1.602
r104 34 49 2.43474 $w=3.53e-07 $l=7.5e-08 $layer=LI1_cond $X=2.16 $Y=1.602
+ $X2=2.235 $Y2=1.602
r105 34 45 8.60274 $w=3.53e-07 $l=2.65e-07 $layer=LI1_cond $X=2.16 $Y=1.602
+ $X2=1.895 $Y2=1.602
r106 33 45 6.97958 $w=3.53e-07 $l=2.15e-07 $layer=LI1_cond $X=1.68 $Y=1.602
+ $X2=1.895 $Y2=1.602
r107 29 60 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.195 $Y=1.675
+ $X2=3.195 $Y2=1.51
r108 29 31 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.195 $Y=1.675
+ $X2=3.195 $Y2=2.465
r109 25 59 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.095 $Y=1.345
+ $X2=3.095 $Y2=1.51
r110 25 27 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=3.095 $Y=1.345
+ $X2=3.095 $Y2=0.745
r111 21 55 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.765 $Y=1.675
+ $X2=2.765 $Y2=1.51
r112 21 23 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.765 $Y=1.675
+ $X2=2.765 $Y2=2.465
r113 17 54 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.665 $Y=1.345
+ $X2=2.665 $Y2=1.51
r114 17 19 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=2.665 $Y=1.345
+ $X2=2.665 $Y2=0.745
r115 13 50 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.335 $Y=1.675
+ $X2=2.335 $Y2=1.51
r116 13 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.335 $Y=1.675
+ $X2=2.335 $Y2=2.465
r117 9 48 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.235 $Y=1.345
+ $X2=2.235 $Y2=1.51
r118 9 11 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=2.235 $Y=1.345
+ $X2=2.235 $Y2=0.745
r119 5 46 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.905 $Y=1.675
+ $X2=1.905 $Y2=1.51
r120 5 7 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.905 $Y=1.675
+ $X2=1.905 $Y2=2.465
r121 1 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.805 $Y=1.345
+ $X2=1.805 $Y2=1.51
r122 1 3 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=1.805 $Y=1.345 $X2=1.805
+ $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_LP__O2BB2AI_4%A_804_39# 1 2 3 4 5 6 21 25 29 33 37 41 45
+ 49 51 60 61 62 65 69 73 77 81 85 87 91 95 97 100 101 102 104 108 110 115 125
c190 97 0 5.44017e-20 $X=9.815 $Y=1.165
r191 122 123 57.7042 $w=3.3e-07 $l=3.3e-07 $layer=POLY_cond $X=5.055 $Y=1.51
+ $X2=5.385 $Y2=1.51
r192 121 122 17.4861 $w=3.3e-07 $l=1e-07 $layer=POLY_cond $X=4.955 $Y=1.51
+ $X2=5.055 $Y2=1.51
r193 120 121 71.6931 $w=3.3e-07 $l=4.1e-07 $layer=POLY_cond $X=4.545 $Y=1.51
+ $X2=4.955 $Y2=1.51
r194 119 120 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=4.525 $Y=1.51
+ $X2=4.545 $Y2=1.51
r195 112 113 9.01001 $w=3.28e-07 $l=2.58e-07 $layer=LI1_cond $X=9.31 $Y=0.907
+ $X2=9.31 $Y2=1.165
r196 110 112 7.22896 $w=3.28e-07 $l=2.07e-07 $layer=LI1_cond $X=9.31 $Y=0.7
+ $X2=9.31 $Y2=0.907
r197 104 106 5.26282 $w=2.98e-07 $l=1.37e-07 $layer=LI1_cond $X=8.435 $Y=0.77
+ $X2=8.435 $Y2=0.907
r198 99 100 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=9.905 $Y=1.255
+ $X2=9.905 $Y2=1.765
r199 98 113 4.28565 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=9.475 $Y=1.165
+ $X2=9.31 $Y2=1.165
r200 97 99 6.81649 $w=1.8e-07 $l=1.27279e-07 $layer=LI1_cond $X=9.815 $Y=1.165
+ $X2=9.905 $Y2=1.255
r201 97 98 20.9495 $w=1.78e-07 $l=3.4e-07 $layer=LI1_cond $X=9.815 $Y=1.165
+ $X2=9.475 $Y2=1.165
r202 96 115 5.16603 $w=1.8e-07 $l=9e-08 $layer=LI1_cond $X=9.39 $Y=1.855 $X2=9.3
+ $Y2=1.855
r203 95 100 6.81649 $w=1.8e-07 $l=1.27279e-07 $layer=LI1_cond $X=9.815 $Y=1.855
+ $X2=9.905 $Y2=1.765
r204 95 96 26.1869 $w=1.78e-07 $l=4.25e-07 $layer=LI1_cond $X=9.815 $Y=1.855
+ $X2=9.39 $Y2=1.855
r205 91 93 57.303 $w=1.78e-07 $l=9.3e-07 $layer=LI1_cond $X=9.3 $Y=1.98 $X2=9.3
+ $Y2=2.91
r206 89 115 1.34256 $w=1.8e-07 $l=9e-08 $layer=LI1_cond $X=9.3 $Y=1.945 $X2=9.3
+ $Y2=1.855
r207 89 91 2.15657 $w=1.78e-07 $l=3.5e-08 $layer=LI1_cond $X=9.3 $Y=1.945
+ $X2=9.3 $Y2=1.98
r208 88 106 3.58581 $w=1.85e-07 $l=1.5e-07 $layer=LI1_cond $X=8.585 $Y=0.907
+ $X2=8.435 $Y2=0.907
r209 87 112 4.14273 $w=1.85e-07 $l=1.65e-07 $layer=LI1_cond $X=9.145 $Y=0.907
+ $X2=9.31 $Y2=0.907
r210 87 88 33.5725 $w=1.83e-07 $l=5.6e-07 $layer=LI1_cond $X=9.145 $Y=0.907
+ $X2=8.585 $Y2=0.907
r211 86 108 5.40251 $w=1.8e-07 $l=9.5e-08 $layer=LI1_cond $X=8.53 $Y=1.855
+ $X2=8.435 $Y2=1.855
r212 85 115 5.16603 $w=1.8e-07 $l=9e-08 $layer=LI1_cond $X=9.21 $Y=1.855 $X2=9.3
+ $Y2=1.855
r213 85 86 41.899 $w=1.78e-07 $l=6.8e-07 $layer=LI1_cond $X=9.21 $Y=1.855
+ $X2=8.53 $Y2=1.855
r214 81 83 54.2871 $w=1.88e-07 $l=9.3e-07 $layer=LI1_cond $X=8.435 $Y=1.98
+ $X2=8.435 $Y2=2.91
r215 79 108 1.14861 $w=1.9e-07 $l=9e-08 $layer=LI1_cond $X=8.435 $Y=1.945
+ $X2=8.435 $Y2=1.855
r216 79 81 2.04306 $w=1.88e-07 $l=3.5e-08 $layer=LI1_cond $X=8.435 $Y=1.945
+ $X2=8.435 $Y2=1.98
r217 78 102 5.40251 $w=1.8e-07 $l=9.5e-08 $layer=LI1_cond $X=7.33 $Y=1.855
+ $X2=7.235 $Y2=1.855
r218 77 108 5.40251 $w=1.8e-07 $l=9.5e-08 $layer=LI1_cond $X=8.34 $Y=1.855
+ $X2=8.435 $Y2=1.855
r219 77 78 62.2323 $w=1.78e-07 $l=1.01e-06 $layer=LI1_cond $X=8.34 $Y=1.855
+ $X2=7.33 $Y2=1.855
r220 73 75 54.2871 $w=1.88e-07 $l=9.3e-07 $layer=LI1_cond $X=7.235 $Y=1.98
+ $X2=7.235 $Y2=2.91
r221 71 102 1.14861 $w=1.9e-07 $l=9e-08 $layer=LI1_cond $X=7.235 $Y=1.945
+ $X2=7.235 $Y2=1.855
r222 71 73 2.04306 $w=1.88e-07 $l=3.5e-08 $layer=LI1_cond $X=7.235 $Y=1.945
+ $X2=7.235 $Y2=1.98
r223 70 101 5.40251 $w=1.8e-07 $l=9.5e-08 $layer=LI1_cond $X=6.47 $Y=1.855
+ $X2=6.375 $Y2=1.855
r224 69 102 5.40251 $w=1.8e-07 $l=9.5e-08 $layer=LI1_cond $X=7.14 $Y=1.855
+ $X2=7.235 $Y2=1.855
r225 69 70 41.2828 $w=1.78e-07 $l=6.7e-07 $layer=LI1_cond $X=7.14 $Y=1.855
+ $X2=6.47 $Y2=1.855
r226 65 67 54.2871 $w=1.88e-07 $l=9.3e-07 $layer=LI1_cond $X=6.375 $Y=1.98
+ $X2=6.375 $Y2=2.91
r227 63 101 1.14861 $w=1.9e-07 $l=9e-08 $layer=LI1_cond $X=6.375 $Y=1.945
+ $X2=6.375 $Y2=1.855
r228 63 65 2.04306 $w=1.88e-07 $l=3.5e-08 $layer=LI1_cond $X=6.375 $Y=1.945
+ $X2=6.375 $Y2=1.98
r229 61 101 5.40251 $w=1.8e-07 $l=9.5e-08 $layer=LI1_cond $X=6.28 $Y=1.855
+ $X2=6.375 $Y2=1.855
r230 61 62 34.197 $w=1.78e-07 $l=5.55e-07 $layer=LI1_cond $X=6.28 $Y=1.855
+ $X2=5.725 $Y2=1.855
r231 60 62 6.82373 $w=1.8e-07 $l=1.25499e-07 $layer=LI1_cond $X=5.64 $Y=1.765
+ $X2=5.725 $Y2=1.855
r232 59 60 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=5.64 $Y=1.595
+ $X2=5.64 $Y2=1.765
r233 58 125 6.12014 $w=3.3e-07 $l=3.5e-08 $layer=POLY_cond $X=5.53 $Y=1.51
+ $X2=5.565 $Y2=1.51
r234 58 123 25.3549 $w=3.3e-07 $l=1.45e-07 $layer=POLY_cond $X=5.53 $Y=1.51
+ $X2=5.385 $Y2=1.51
r235 57 58 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.53
+ $Y=1.51 $X2=5.53 $Y2=1.51
r236 54 119 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=4.51 $Y=1.51
+ $X2=4.525 $Y2=1.51
r237 54 116 72.5674 $w=3.3e-07 $l=4.15e-07 $layer=POLY_cond $X=4.51 $Y=1.51
+ $X2=4.095 $Y2=1.51
r238 53 57 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=4.51 $Y=1.51
+ $X2=5.53 $Y2=1.51
r239 53 54 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.51
+ $Y=1.51 $X2=4.51 $Y2=1.51
r240 51 59 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.555 $Y=1.51
+ $X2=5.64 $Y2=1.595
r241 51 57 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=5.555 $Y=1.51
+ $X2=5.53 $Y2=1.51
r242 47 125 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.565 $Y=1.345
+ $X2=5.565 $Y2=1.51
r243 47 49 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=5.565 $Y=1.345
+ $X2=5.565 $Y2=0.745
r244 43 123 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.385 $Y=1.675
+ $X2=5.385 $Y2=1.51
r245 43 45 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=5.385 $Y=1.675
+ $X2=5.385 $Y2=2.465
r246 39 122 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.055 $Y=1.345
+ $X2=5.055 $Y2=1.51
r247 39 41 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=5.055 $Y=1.345
+ $X2=5.055 $Y2=0.745
r248 35 121 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.955 $Y=1.675
+ $X2=4.955 $Y2=1.51
r249 35 37 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=4.955 $Y=1.675
+ $X2=4.955 $Y2=2.465
r250 31 120 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.545 $Y=1.345
+ $X2=4.545 $Y2=1.51
r251 31 33 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=4.545 $Y=1.345
+ $X2=4.545 $Y2=0.745
r252 27 119 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.525 $Y=1.675
+ $X2=4.525 $Y2=1.51
r253 27 29 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=4.525 $Y=1.675
+ $X2=4.525 $Y2=2.465
r254 23 116 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.095 $Y=1.675
+ $X2=4.095 $Y2=1.51
r255 23 25 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=4.095 $Y=1.675
+ $X2=4.095 $Y2=2.465
r256 19 116 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.095 $Y=1.345
+ $X2=4.095 $Y2=1.51
r257 19 21 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=4.095 $Y=1.345
+ $X2=4.095 $Y2=0.745
r258 6 93 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=9.155
+ $Y=1.835 $X2=9.295 $Y2=2.91
r259 6 91 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=9.155
+ $Y=1.835 $X2=9.295 $Y2=1.98
r260 5 83 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=8.295
+ $Y=1.835 $X2=8.435 $Y2=2.91
r261 5 81 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=8.295
+ $Y=1.835 $X2=8.435 $Y2=1.98
r262 4 75 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=7.095
+ $Y=1.835 $X2=7.235 $Y2=2.91
r263 4 73 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=7.095
+ $Y=1.835 $X2=7.235 $Y2=1.98
r264 3 67 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=6.235
+ $Y=1.835 $X2=6.375 $Y2=2.91
r265 3 65 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=6.235
+ $Y=1.835 $X2=6.375 $Y2=1.98
r266 2 110 91 $w=1.7e-07 $l=4.3946e-07 $layer=licon1_NDIFF $count=2 $X=9.17
+ $Y=0.325 $X2=9.31 $Y2=0.7
r267 1 104 182 $w=1.7e-07 $l=5.10221e-07 $layer=licon1_NDIFF $count=1 $X=8.31
+ $Y=0.325 $X2=8.45 $Y2=0.77
.ends

.subckt PM_SKY130_FD_SC_LP__O2BB2AI_4%A1_N 3 7 11 15 19 23 27 31 38 41 42 58 60
+ 67
c92 23 0 1.73643e-19 $X=7.375 $Y=0.745
r93 55 56 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=7.375 $Y=1.51
+ $X2=7.45 $Y2=1.51
r94 54 55 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=7.02 $Y=1.51
+ $X2=7.375 $Y2=1.51
r95 53 54 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=6.945 $Y=1.51
+ $X2=7.02 $Y2=1.51
r96 50 51 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=6.515 $Y=1.51
+ $X2=6.59 $Y2=1.51
r97 49 60 1.10754 $w=3.83e-07 $l=3.7e-08 $layer=LI1_cond $X=6.41 $Y=1.402
+ $X2=6.373 $Y2=1.402
r98 48 50 18.3604 $w=3.3e-07 $l=1.05e-07 $layer=POLY_cond $X=6.41 $Y=1.51
+ $X2=6.515 $Y2=1.51
r99 48 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.41
+ $Y=1.51 $X2=6.41 $Y2=1.51
r100 45 48 43.7153 $w=3.3e-07 $l=2.5e-07 $layer=POLY_cond $X=6.16 $Y=1.51
+ $X2=6.41 $Y2=1.51
r101 42 67 6.19425 $w=3.83e-07 $l=8.5e-08 $layer=LI1_cond $X=6.48 $Y=1.402
+ $X2=6.565 $Y2=1.402
r102 42 49 2.09535 $w=3.83e-07 $l=7e-08 $layer=LI1_cond $X=6.48 $Y=1.402
+ $X2=6.41 $Y2=1.402
r103 41 60 11.1652 $w=3.83e-07 $l=3.73e-07 $layer=LI1_cond $X=6 $Y=1.402
+ $X2=6.373 $Y2=1.402
r104 39 58 6.12014 $w=3.3e-07 $l=3.5e-08 $layer=POLY_cond $X=7.77 $Y=1.51
+ $X2=7.805 $Y2=1.51
r105 39 56 55.9556 $w=3.3e-07 $l=3.2e-07 $layer=POLY_cond $X=7.77 $Y=1.51
+ $X2=7.45 $Y2=1.51
r106 38 39 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.77
+ $Y=1.51 $X2=7.77 $Y2=1.51
r107 36 53 34.0979 $w=3.3e-07 $l=1.95e-07 $layer=POLY_cond $X=6.75 $Y=1.51
+ $X2=6.945 $Y2=1.51
r108 36 51 27.9778 $w=3.3e-07 $l=1.6e-07 $layer=POLY_cond $X=6.75 $Y=1.51
+ $X2=6.59 $Y2=1.51
r109 35 38 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=6.75 $Y=1.51
+ $X2=7.77 $Y2=1.51
r110 35 67 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=6.75 $Y=1.51
+ $X2=6.565 $Y2=1.51
r111 35 36 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.75
+ $Y=1.51 $X2=6.75 $Y2=1.51
r112 29 58 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.805 $Y=1.345
+ $X2=7.805 $Y2=1.51
r113 29 31 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=7.805 $Y=1.345
+ $X2=7.805 $Y2=0.745
r114 25 56 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.45 $Y=1.675
+ $X2=7.45 $Y2=1.51
r115 25 27 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=7.45 $Y=1.675
+ $X2=7.45 $Y2=2.465
r116 21 55 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.375 $Y=1.345
+ $X2=7.375 $Y2=1.51
r117 21 23 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=7.375 $Y=1.345
+ $X2=7.375 $Y2=0.745
r118 17 54 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.02 $Y=1.675
+ $X2=7.02 $Y2=1.51
r119 17 19 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=7.02 $Y=1.675
+ $X2=7.02 $Y2=2.465
r120 13 53 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.945 $Y=1.345
+ $X2=6.945 $Y2=1.51
r121 13 15 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=6.945 $Y=1.345
+ $X2=6.945 $Y2=0.745
r122 9 51 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.59 $Y=1.675
+ $X2=6.59 $Y2=1.51
r123 9 11 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=6.59 $Y=1.675
+ $X2=6.59 $Y2=2.465
r124 5 50 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.515 $Y=1.345
+ $X2=6.515 $Y2=1.51
r125 5 7 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=6.515 $Y=1.345 $X2=6.515
+ $Y2=0.745
r126 1 45 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.16 $Y=1.675
+ $X2=6.16 $Y2=1.51
r127 1 3 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=6.16 $Y=1.675
+ $X2=6.16 $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__O2BB2AI_4%A2_N 1 3 6 8 10 13 15 17 20 22 24 27 31 34
+ 35 51 53 61
c85 20 0 1.84104e-19 $X=9.095 $Y=0.745
r86 51 52 1.92287 $w=3.76e-07 $l=1.5e-08 $layer=POLY_cond $X=9.51 $Y=1.535
+ $X2=9.525 $Y2=1.535
r87 48 49 1.92287 $w=3.76e-07 $l=1.5e-08 $layer=POLY_cond $X=9.08 $Y=1.535
+ $X2=9.095 $Y2=1.535
r88 47 53 0.73214 $w=4.23e-07 $l=2.7e-08 $layer=LI1_cond $X=8.79 $Y=1.382
+ $X2=8.763 $Y2=1.382
r89 46 48 37.1755 $w=3.76e-07 $l=2.9e-07 $layer=POLY_cond $X=8.79 $Y=1.535
+ $X2=9.08 $Y2=1.535
r90 46 47 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.79
+ $Y=1.51 $X2=8.79 $Y2=1.51
r91 44 46 16.0239 $w=3.76e-07 $l=1.25e-07 $layer=POLY_cond $X=8.665 $Y=1.535
+ $X2=8.79 $Y2=1.535
r92 43 44 1.92287 $w=3.76e-07 $l=1.5e-08 $layer=POLY_cond $X=8.65 $Y=1.535
+ $X2=8.665 $Y2=1.535
r93 42 53 8.4874 $w=4.23e-07 $l=3.13e-07 $layer=LI1_cond $X=8.45 $Y=1.382
+ $X2=8.763 $Y2=1.382
r94 41 43 25.6383 $w=3.76e-07 $l=2e-07 $layer=POLY_cond $X=8.45 $Y=1.535
+ $X2=8.65 $Y2=1.535
r95 41 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.45
+ $Y=1.51 $X2=8.45 $Y2=1.51
r96 39 41 27.5612 $w=3.76e-07 $l=2.15e-07 $layer=POLY_cond $X=8.235 $Y=1.535
+ $X2=8.45 $Y2=1.535
r97 38 39 1.92287 $w=3.76e-07 $l=1.5e-08 $layer=POLY_cond $X=8.22 $Y=1.535
+ $X2=8.235 $Y2=1.535
r98 35 61 6.86232 $w=4.23e-07 $l=9.5e-08 $layer=LI1_cond $X=8.88 $Y=1.382
+ $X2=8.975 $Y2=1.382
r99 35 47 2.44047 $w=4.23e-07 $l=9e-08 $layer=LI1_cond $X=8.88 $Y=1.382 $X2=8.79
+ $Y2=1.382
r100 34 42 1.35582 $w=4.23e-07 $l=5e-08 $layer=LI1_cond $X=8.4 $Y=1.382 $X2=8.45
+ $Y2=1.382
r101 32 51 5.12766 $w=3.76e-07 $l=4e-08 $layer=POLY_cond $X=9.47 $Y=1.535
+ $X2=9.51 $Y2=1.535
r102 32 49 48.0718 $w=3.76e-07 $l=3.75e-07 $layer=POLY_cond $X=9.47 $Y=1.535
+ $X2=9.095 $Y2=1.535
r103 31 61 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=9.47 $Y=1.51
+ $X2=8.975 $Y2=1.51
r104 31 32 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=9.47
+ $Y=1.51 $X2=9.47 $Y2=1.51
r105 25 52 24.356 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=9.525 $Y=1.345
+ $X2=9.525 $Y2=1.535
r106 25 27 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=9.525 $Y=1.345
+ $X2=9.525 $Y2=0.745
r107 22 51 24.356 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=9.51 $Y=1.725
+ $X2=9.51 $Y2=1.535
r108 22 24 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=9.51 $Y=1.725
+ $X2=9.51 $Y2=2.465
r109 18 49 24.356 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=9.095 $Y=1.345
+ $X2=9.095 $Y2=1.535
r110 18 20 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=9.095 $Y=1.345
+ $X2=9.095 $Y2=0.745
r111 15 48 24.356 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=9.08 $Y=1.725
+ $X2=9.08 $Y2=1.535
r112 15 17 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=9.08 $Y=1.725
+ $X2=9.08 $Y2=2.465
r113 11 44 24.356 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=8.665 $Y=1.345
+ $X2=8.665 $Y2=1.535
r114 11 13 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=8.665 $Y=1.345
+ $X2=8.665 $Y2=0.745
r115 8 43 24.356 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=8.65 $Y=1.725
+ $X2=8.65 $Y2=1.535
r116 8 10 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=8.65 $Y=1.725
+ $X2=8.65 $Y2=2.465
r117 4 39 24.356 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=8.235 $Y=1.345
+ $X2=8.235 $Y2=1.535
r118 4 6 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=8.235 $Y=1.345 $X2=8.235
+ $Y2=0.745
r119 1 38 24.356 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=8.22 $Y=1.725
+ $X2=8.22 $Y2=1.535
r120 1 3 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=8.22 $Y=1.725
+ $X2=8.22 $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__O2BB2AI_4%VPWR 1 2 3 4 5 6 7 8 9 28 30 36 40 44 50
+ 56 62 68 72 74 79 80 82 83 85 86 87 89 104 112 116 121 130 133 136 139 143
r160 142 143 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r161 139 140 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r162 136 137 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r163 133 134 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r164 130 131 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r165 127 128 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r166 125 143 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=9.84 $Y2=3.33
r167 125 140 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=8.88 $Y2=3.33
r168 124 125 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r169 122 139 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.03 $Y=3.33
+ $X2=8.865 $Y2=3.33
r170 122 124 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=9.03 $Y=3.33
+ $X2=9.36 $Y2=3.33
r171 121 142 4.5891 $w=1.7e-07 $l=2.6e-07 $layer=LI1_cond $X=9.56 $Y=3.33
+ $X2=9.82 $Y2=3.33
r172 121 124 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=9.56 $Y=3.33
+ $X2=9.36 $Y2=3.33
r173 120 140 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=8.88 $Y2=3.33
r174 120 137 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=7.92 $Y2=3.33
r175 119 120 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r176 117 136 13.3456 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=8.17 $Y=3.33
+ $X2=7.835 $Y2=3.33
r177 117 119 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=8.17 $Y=3.33
+ $X2=8.4 $Y2=3.33
r178 116 139 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.7 $Y=3.33
+ $X2=8.865 $Y2=3.33
r179 116 119 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=8.7 $Y=3.33 $X2=8.4
+ $Y2=3.33
r180 115 137 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=7.92 $Y2=3.33
r181 114 115 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r182 112 136 13.3456 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=7.5 $Y=3.33
+ $X2=7.835 $Y2=3.33
r183 112 114 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=7.5 $Y=3.33
+ $X2=7.44 $Y2=3.33
r184 111 115 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=7.44 $Y2=3.33
r185 111 134 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=6 $Y2=3.33
r186 110 111 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r187 108 133 13.399 $w=1.7e-07 $l=3.38e-07 $layer=LI1_cond $X=6.11 $Y=3.33
+ $X2=5.772 $Y2=3.33
r188 108 110 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=6.11 $Y=3.33
+ $X2=6.48 $Y2=3.33
r189 104 133 13.399 $w=1.7e-07 $l=3.37e-07 $layer=LI1_cond $X=5.435 $Y=3.33
+ $X2=5.772 $Y2=3.33
r190 104 106 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=5.435 $Y=3.33
+ $X2=5.04 $Y2=3.33
r191 102 103 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r192 100 103 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.56 $Y2=3.33
r193 99 100 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r194 97 100 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=3.6 $Y2=3.33
r195 97 131 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r196 96 99 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=1.68 $Y=3.33
+ $X2=3.6 $Y2=3.33
r197 96 97 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r198 94 130 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.395 $Y=3.33
+ $X2=1.23 $Y2=3.33
r199 94 96 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.395 $Y=3.33
+ $X2=1.68 $Y2=3.33
r200 93 131 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r201 93 128 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r202 92 93 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r203 90 127 3.60924 $w=1.7e-07 $l=2.38e-07 $layer=LI1_cond $X=0.475 $Y=3.33
+ $X2=0.237 $Y2=3.33
r204 90 92 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=0.475 $Y=3.33
+ $X2=0.72 $Y2=3.33
r205 89 130 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.065 $Y=3.33
+ $X2=1.23 $Y2=3.33
r206 89 92 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.065 $Y=3.33
+ $X2=0.72 $Y2=3.33
r207 87 134 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=6 $Y2=3.33
r208 87 103 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=4.56 $Y2=3.33
r209 87 106 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r210 85 110 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=6.64 $Y=3.33
+ $X2=6.48 $Y2=3.33
r211 85 86 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.64 $Y=3.33
+ $X2=6.805 $Y2=3.33
r212 84 114 30.6631 $w=1.68e-07 $l=4.7e-07 $layer=LI1_cond $X=6.97 $Y=3.33
+ $X2=7.44 $Y2=3.33
r213 84 86 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.97 $Y=3.33
+ $X2=6.805 $Y2=3.33
r214 82 102 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=4.575 $Y=3.33
+ $X2=4.56 $Y2=3.33
r215 82 83 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.575 $Y=3.33
+ $X2=4.74 $Y2=3.33
r216 81 106 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=4.905 $Y=3.33
+ $X2=5.04 $Y2=3.33
r217 81 83 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.905 $Y=3.33
+ $X2=4.74 $Y2=3.33
r218 79 99 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=3.745 $Y=3.33
+ $X2=3.6 $Y2=3.33
r219 79 80 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=3.745 $Y=3.33
+ $X2=3.895 $Y2=3.33
r220 78 102 33.5989 $w=1.68e-07 $l=5.15e-07 $layer=LI1_cond $X=4.045 $Y=3.33
+ $X2=4.56 $Y2=3.33
r221 78 80 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=4.045 $Y=3.33
+ $X2=3.895 $Y2=3.33
r222 74 77 26.1919 $w=3.28e-07 $l=7.5e-07 $layer=LI1_cond $X=9.725 $Y=2.2
+ $X2=9.725 $Y2=2.95
r223 72 142 3.17707 $w=3.3e-07 $l=1.30767e-07 $layer=LI1_cond $X=9.725 $Y=3.245
+ $X2=9.82 $Y2=3.33
r224 72 77 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=9.725 $Y=3.245
+ $X2=9.725 $Y2=2.95
r225 68 71 26.5411 $w=3.28e-07 $l=7.6e-07 $layer=LI1_cond $X=8.865 $Y=2.21
+ $X2=8.865 $Y2=2.97
r226 66 139 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.865 $Y=3.245
+ $X2=8.865 $Y2=3.33
r227 66 71 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=8.865 $Y=3.245
+ $X2=8.865 $Y2=2.97
r228 62 65 13.5675 $w=6.68e-07 $l=7.6e-07 $layer=LI1_cond $X=7.835 $Y=2.21
+ $X2=7.835 $Y2=2.97
r229 60 136 2.76849 $w=6.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.835 $Y=3.245
+ $X2=7.835 $Y2=3.33
r230 60 65 4.90928 $w=6.68e-07 $l=2.75e-07 $layer=LI1_cond $X=7.835 $Y=3.245
+ $X2=7.835 $Y2=2.97
r231 56 59 26.5411 $w=3.28e-07 $l=7.6e-07 $layer=LI1_cond $X=6.805 $Y=2.21
+ $X2=6.805 $Y2=2.97
r232 54 86 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.805 $Y=3.245
+ $X2=6.805 $Y2=3.33
r233 54 59 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=6.805 $Y=3.245
+ $X2=6.805 $Y2=2.97
r234 50 53 13.467 $w=6.73e-07 $l=7.6e-07 $layer=LI1_cond $X=5.772 $Y=2.21
+ $X2=5.772 $Y2=2.97
r235 48 133 2.78459 $w=6.75e-07 $l=8.5e-08 $layer=LI1_cond $X=5.772 $Y=3.245
+ $X2=5.772 $Y2=3.33
r236 48 53 4.87291 $w=6.73e-07 $l=2.75e-07 $layer=LI1_cond $X=5.772 $Y=3.245
+ $X2=5.772 $Y2=2.97
r237 44 47 26.5411 $w=3.28e-07 $l=7.6e-07 $layer=LI1_cond $X=4.74 $Y=2.21
+ $X2=4.74 $Y2=2.97
r238 42 83 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.74 $Y=3.245
+ $X2=4.74 $Y2=3.33
r239 42 47 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=4.74 $Y=3.245
+ $X2=4.74 $Y2=2.97
r240 38 80 0.597483 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.895 $Y=3.245
+ $X2=3.895 $Y2=3.33
r241 38 40 10.7561 $w=2.98e-07 $l=2.8e-07 $layer=LI1_cond $X=3.895 $Y=3.245
+ $X2=3.895 $Y2=2.965
r242 34 130 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.23 $Y=3.245
+ $X2=1.23 $Y2=3.33
r243 34 36 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=1.23 $Y=3.245
+ $X2=1.23 $Y2=2.815
r244 30 33 51.2294 $w=2.08e-07 $l=9.7e-07 $layer=LI1_cond $X=0.37 $Y=1.98
+ $X2=0.37 $Y2=2.95
r245 28 127 3.30595 $w=2.1e-07 $l=1.70276e-07 $layer=LI1_cond $X=0.37 $Y=3.245
+ $X2=0.237 $Y2=3.33
r246 28 33 15.5801 $w=2.08e-07 $l=2.95e-07 $layer=LI1_cond $X=0.37 $Y=3.245
+ $X2=0.37 $Y2=2.95
r247 9 77 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=9.585
+ $Y=1.835 $X2=9.725 $Y2=2.95
r248 9 74 400 $w=1.7e-07 $l=4.29331e-07 $layer=licon1_PDIFF $count=1 $X=9.585
+ $Y=1.835 $X2=9.725 $Y2=2.2
r249 8 71 400 $w=1.7e-07 $l=1.20297e-06 $layer=licon1_PDIFF $count=1 $X=8.725
+ $Y=1.835 $X2=8.865 $Y2=2.97
r250 8 68 400 $w=1.7e-07 $l=4.3946e-07 $layer=licon1_PDIFF $count=1 $X=8.725
+ $Y=1.835 $X2=8.865 $Y2=2.21
r251 7 65 200 $w=1.7e-07 $l=1.20297e-06 $layer=licon1_PDIFF $count=3 $X=7.525
+ $Y=1.835 $X2=7.665 $Y2=2.97
r252 7 62 200 $w=1.7e-07 $l=4.3946e-07 $layer=licon1_PDIFF $count=3 $X=7.525
+ $Y=1.835 $X2=7.665 $Y2=2.21
r253 6 59 400 $w=1.7e-07 $l=1.20297e-06 $layer=licon1_PDIFF $count=1 $X=6.665
+ $Y=1.835 $X2=6.805 $Y2=2.97
r254 6 56 400 $w=1.7e-07 $l=4.3946e-07 $layer=licon1_PDIFF $count=1 $X=6.665
+ $Y=1.835 $X2=6.805 $Y2=2.21
r255 5 53 200 $w=1.7e-07 $l=1.20297e-06 $layer=licon1_PDIFF $count=3 $X=5.46
+ $Y=1.835 $X2=5.6 $Y2=2.97
r256 5 50 200 $w=1.7e-07 $l=4.3946e-07 $layer=licon1_PDIFF $count=3 $X=5.46
+ $Y=1.835 $X2=5.6 $Y2=2.21
r257 4 47 400 $w=1.7e-07 $l=1.20297e-06 $layer=licon1_PDIFF $count=1 $X=4.6
+ $Y=1.835 $X2=4.74 $Y2=2.97
r258 4 44 400 $w=1.7e-07 $l=4.3946e-07 $layer=licon1_PDIFF $count=1 $X=4.6
+ $Y=1.835 $X2=4.74 $Y2=2.21
r259 3 40 600 $w=1.7e-07 $l=1.21668e-06 $layer=licon1_PDIFF $count=1 $X=3.7
+ $Y=1.835 $X2=3.88 $Y2=2.965
r260 2 36 600 $w=1.7e-07 $l=1.04766e-06 $layer=licon1_PDIFF $count=1 $X=1.09
+ $Y=1.835 $X2=1.23 $Y2=2.815
r261 1 33 400 $w=1.7e-07 $l=1.17584e-06 $layer=licon1_PDIFF $count=1 $X=0.245
+ $Y=1.835 $X2=0.37 $Y2=2.95
r262 1 30 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.245
+ $Y=1.835 $X2=0.37 $Y2=1.98
.ends

.subckt PM_SKY130_FD_SC_LP__O2BB2AI_4%A_132_367# 1 2 3 4 15 19 21 23 24 29
c41 4 0 1.33268e-19 $X=3.27 $Y=1.835
r42 27 29 36.04 $w=2.73e-07 $l=8.6e-07 $layer=LI1_cond $X=2.55 $Y=2.937 $X2=3.41
+ $Y2=2.937
r43 25 36 3.02719 $w=2.75e-07 $l=1.05e-07 $layer=LI1_cond $X=1.785 $Y=2.937
+ $X2=1.68 $Y2=2.937
r44 25 27 32.0589 $w=2.73e-07 $l=7.65e-07 $layer=LI1_cond $X=1.785 $Y=2.937
+ $X2=2.55 $Y2=2.937
r45 24 36 3.94976 $w=2.1e-07 $l=1.37e-07 $layer=LI1_cond $X=1.68 $Y=2.8 $X2=1.68
+ $Y2=2.937
r46 23 34 3.09364 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=1.68 $Y=2.52 $X2=1.68
+ $Y2=2.435
r47 23 24 14.7879 $w=2.08e-07 $l=2.8e-07 $layer=LI1_cond $X=1.68 $Y=2.52
+ $X2=1.68 $Y2=2.8
r48 22 32 1.84097 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=0.895 $Y=2.435
+ $X2=0.795 $Y2=2.435
r49 21 34 3.82155 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.575 $Y=2.435
+ $X2=1.68 $Y2=2.435
r50 21 22 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.575 $Y=2.435
+ $X2=0.895 $Y2=2.435
r51 17 32 4.60183 $w=1.95e-07 $l=8.5e-08 $layer=LI1_cond $X=0.795 $Y=2.52
+ $X2=0.795 $Y2=2.435
r52 17 19 21.6273 $w=1.98e-07 $l=3.9e-07 $layer=LI1_cond $X=0.795 $Y=2.52
+ $X2=0.795 $Y2=2.91
r53 13 32 4.60183 $w=1.95e-07 $l=8.74643e-08 $layer=LI1_cond $X=0.79 $Y=2.35
+ $X2=0.795 $Y2=2.435
r54 13 15 21.5981 $w=1.88e-07 $l=3.7e-07 $layer=LI1_cond $X=0.79 $Y=2.35
+ $X2=0.79 $Y2=1.98
r55 4 29 600 $w=1.7e-07 $l=1.14787e-06 $layer=licon1_PDIFF $count=1 $X=3.27
+ $Y=1.835 $X2=3.41 $Y2=2.915
r56 3 27 600 $w=1.7e-07 $l=1.14787e-06 $layer=licon1_PDIFF $count=1 $X=2.41
+ $Y=1.835 $X2=2.55 $Y2=2.915
r57 2 36 600 $w=1.7e-07 $l=1.15223e-06 $layer=licon1_PDIFF $count=1 $X=1.52
+ $Y=1.835 $X2=1.68 $Y2=2.91
r58 2 34 600 $w=1.7e-07 $l=7.55778e-07 $layer=licon1_PDIFF $count=1 $X=1.52
+ $Y=1.835 $X2=1.68 $Y2=2.515
r59 1 32 600 $w=1.7e-07 $l=6.66333e-07 $layer=licon1_PDIFF $count=1 $X=0.66
+ $Y=1.835 $X2=0.8 $Y2=2.435
r60 1 19 600 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=0.66
+ $Y=1.835 $X2=0.8 $Y2=2.91
r61 1 15 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.66
+ $Y=1.835 $X2=0.8 $Y2=1.98
.ends

.subckt PM_SKY130_FD_SC_LP__O2BB2AI_4%Y 1 2 3 4 5 6 20 24 27 31 33 35 39 45 47
+ 48 49 50 51 52 53
c85 27 0 1.8603e-19 $X=4.33 $Y=0.7
r86 52 53 10.8327 $w=4.98e-07 $l=3.95e-07 $layer=LI1_cond $X=3.6 $Y=2.465
+ $X2=3.995 $Y2=2.465
r87 51 52 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=3.12 $Y=2.465
+ $X2=3.6 $Y2=2.465
r88 51 68 4.88915 $w=3.28e-07 $l=1.4e-07 $layer=LI1_cond $X=3.12 $Y=2.465
+ $X2=2.98 $Y2=2.465
r89 50 68 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=2.64 $Y=2.465
+ $X2=2.98 $Y2=2.465
r90 49 50 18.1597 $w=3.28e-07 $l=5.2e-07 $layer=LI1_cond $X=2.12 $Y=2.465
+ $X2=2.64 $Y2=2.465
r91 43 45 13.0959 $w=3.28e-07 $l=3.75e-07 $layer=LI1_cond $X=5.35 $Y=1.075
+ $X2=5.35 $Y2=0.7
r92 39 41 54.2871 $w=1.88e-07 $l=9.3e-07 $layer=LI1_cond $X=5.17 $Y=1.98
+ $X2=5.17 $Y2=2.91
r93 37 39 2.04306 $w=1.88e-07 $l=3.5e-08 $layer=LI1_cond $X=5.17 $Y=1.945
+ $X2=5.17 $Y2=1.98
r94 36 47 2.76166 $w=1.7e-07 $l=2.5e-07 $layer=LI1_cond $X=4.495 $Y=1.16
+ $X2=4.245 $Y2=1.16
r95 35 43 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.185 $Y=1.16
+ $X2=5.35 $Y2=1.075
r96 35 36 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=5.185 $Y=1.16
+ $X2=4.495 $Y2=1.16
r97 34 48 3.3199 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=4.405 $Y=1.86 $X2=4.2
+ $Y2=1.86
r98 33 37 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=5.075 $Y=1.86
+ $X2=5.17 $Y2=1.945
r99 33 34 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.075 $Y=1.86
+ $X2=4.405 $Y2=1.86
r100 29 53 5.58832 $w=3e-07 $l=2.13014e-07 $layer=LI1_cond $X=4.31 $Y=2.63
+ $X2=4.2 $Y2=2.465
r101 29 31 16.3445 $w=1.88e-07 $l=2.8e-07 $layer=LI1_cond $X=4.31 $Y=2.63
+ $X2=4.31 $Y2=2.91
r102 25 47 3.70735 $w=2.5e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.33 $Y=1.075
+ $X2=4.245 $Y2=1.16
r103 25 27 13.0959 $w=3.28e-07 $l=3.75e-07 $layer=LI1_cond $X=4.33 $Y=1.075
+ $X2=4.33 $Y2=0.7
r104 22 53 5.58832 $w=3e-07 $l=1.65e-07 $layer=LI1_cond $X=4.2 $Y=2.3 $X2=4.2
+ $Y2=2.465
r105 22 24 8.99468 $w=4.08e-07 $l=3.2e-07 $layer=LI1_cond $X=4.2 $Y=2.3 $X2=4.2
+ $Y2=1.98
r106 21 48 3.24686 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=4.2 $Y=1.945 $X2=4.2
+ $Y2=1.86
r107 21 24 0.983793 $w=4.08e-07 $l=3.5e-08 $layer=LI1_cond $X=4.2 $Y=1.945
+ $X2=4.2 $Y2=1.98
r108 20 48 3.24686 $w=2.9e-07 $l=1.56844e-07 $layer=LI1_cond $X=4.08 $Y=1.775
+ $X2=4.2 $Y2=1.86
r109 19 47 3.70735 $w=2.5e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.08 $Y=1.245
+ $X2=4.245 $Y2=1.16
r110 19 20 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=4.08 $Y=1.245
+ $X2=4.08 $Y2=1.775
r111 6 41 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=5.03
+ $Y=1.835 $X2=5.17 $Y2=2.91
r112 6 39 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=5.03
+ $Y=1.835 $X2=5.17 $Y2=1.98
r113 5 31 600 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=4.17
+ $Y=1.835 $X2=4.31 $Y2=2.91
r114 5 24 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=4.17
+ $Y=1.835 $X2=4.31 $Y2=1.98
r115 4 68 600 $w=1.7e-07 $l=6.96491e-07 $layer=licon1_PDIFF $count=1 $X=2.84
+ $Y=1.835 $X2=2.98 $Y2=2.465
r116 3 49 600 $w=1.7e-07 $l=6.96491e-07 $layer=licon1_PDIFF $count=1 $X=1.98
+ $Y=1.835 $X2=2.12 $Y2=2.465
r117 2 45 91 $w=1.7e-07 $l=4.72361e-07 $layer=licon1_NDIFF $count=2 $X=5.13
+ $Y=0.325 $X2=5.35 $Y2=0.7
r118 1 27 91 $w=1.7e-07 $l=4.47912e-07 $layer=licon1_NDIFF $count=2 $X=4.17
+ $Y=0.325 $X2=4.33 $Y2=0.7
.ends

.subckt PM_SKY130_FD_SC_LP__O2BB2AI_4%A_35_65# 1 2 3 4 5 6 7 24 26 27 30 32 36
+ 38 42 44 49 51 52 53 56 58 62 64 65 66 67 68
c117 53 0 6.61592e-20 $X=3.985 $Y=0.35
r118 60 62 1.55137 $w=2.58e-07 $l=3.5e-08 $layer=LI1_cond $X=5.815 $Y=0.435
+ $X2=5.815 $Y2=0.47
r119 59 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.005 $Y=0.35
+ $X2=4.84 $Y2=0.35
r120 58 60 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=5.685 $Y=0.35
+ $X2=5.815 $Y2=0.435
r121 58 59 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=5.685 $Y=0.35
+ $X2=5.005 $Y2=0.35
r122 54 68 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.84 $Y=0.435
+ $X2=4.84 $Y2=0.35
r123 54 56 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=4.84 $Y=0.435
+ $X2=4.84 $Y2=0.45
r124 52 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.675 $Y=0.35
+ $X2=4.84 $Y2=0.35
r125 52 53 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=4.675 $Y=0.35
+ $X2=3.985 $Y2=0.35
r126 51 67 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=3.74 $Y=1.085
+ $X2=3.74 $Y2=0.905
r127 47 67 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=3.82 $Y=0.74
+ $X2=3.82 $Y2=0.905
r128 47 49 10.1275 $w=3.28e-07 $l=2.9e-07 $layer=LI1_cond $X=3.82 $Y=0.74
+ $X2=3.82 $Y2=0.45
r129 46 53 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.82 $Y=0.435
+ $X2=3.985 $Y2=0.35
r130 46 49 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=3.82 $Y=0.435
+ $X2=3.82 $Y2=0.45
r131 45 66 5.52892 $w=1.75e-07 $l=9.74679e-08 $layer=LI1_cond $X=2.975 $Y=1.17
+ $X2=2.88 $Y2=1.165
r132 44 51 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.655 $Y=1.17
+ $X2=3.74 $Y2=1.085
r133 44 45 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=3.655 $Y=1.17
+ $X2=2.975 $Y2=1.17
r134 40 66 1.04816 $w=1.9e-07 $l=9e-08 $layer=LI1_cond $X=2.88 $Y=1.075 $X2=2.88
+ $Y2=1.165
r135 40 42 35.3158 $w=1.88e-07 $l=6.05e-07 $layer=LI1_cond $X=2.88 $Y=1.075
+ $X2=2.88 $Y2=0.47
r136 39 65 5.40251 $w=1.8e-07 $l=9.5e-08 $layer=LI1_cond $X=2.115 $Y=1.165
+ $X2=2.02 $Y2=1.165
r137 38 66 5.52892 $w=1.75e-07 $l=9.5e-08 $layer=LI1_cond $X=2.785 $Y=1.165
+ $X2=2.88 $Y2=1.165
r138 38 39 41.2828 $w=1.78e-07 $l=6.7e-07 $layer=LI1_cond $X=2.785 $Y=1.165
+ $X2=2.115 $Y2=1.165
r139 34 65 1.14861 $w=1.9e-07 $l=9e-08 $layer=LI1_cond $X=2.02 $Y=1.075 $X2=2.02
+ $Y2=1.165
r140 34 36 35.3158 $w=1.88e-07 $l=6.05e-07 $layer=LI1_cond $X=2.02 $Y=1.075
+ $X2=2.02 $Y2=0.47
r141 33 64 5.40251 $w=1.8e-07 $l=9.5e-08 $layer=LI1_cond $X=1.255 $Y=1.165
+ $X2=1.16 $Y2=1.165
r142 32 65 5.40251 $w=1.8e-07 $l=9.5e-08 $layer=LI1_cond $X=1.925 $Y=1.165
+ $X2=2.02 $Y2=1.165
r143 32 33 41.2828 $w=1.78e-07 $l=6.7e-07 $layer=LI1_cond $X=1.925 $Y=1.165
+ $X2=1.255 $Y2=1.165
r144 28 64 1.14861 $w=1.9e-07 $l=9e-08 $layer=LI1_cond $X=1.16 $Y=1.075 $X2=1.16
+ $Y2=1.165
r145 28 30 35.3158 $w=1.88e-07 $l=6.05e-07 $layer=LI1_cond $X=1.16 $Y=1.075
+ $X2=1.16 $Y2=0.47
r146 26 64 5.40251 $w=1.8e-07 $l=9.5e-08 $layer=LI1_cond $X=1.065 $Y=1.165
+ $X2=1.16 $Y2=1.165
r147 26 27 41.899 $w=1.78e-07 $l=6.8e-07 $layer=LI1_cond $X=1.065 $Y=1.165
+ $X2=0.385 $Y2=1.165
r148 22 27 7.0541 $w=1.8e-07 $l=1.63936e-07 $layer=LI1_cond $X=0.26 $Y=1.075
+ $X2=0.385 $Y2=1.165
r149 22 24 27.8891 $w=2.48e-07 $l=6.05e-07 $layer=LI1_cond $X=0.26 $Y=1.075
+ $X2=0.26 $Y2=0.47
r150 7 62 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.64
+ $Y=0.325 $X2=5.78 $Y2=0.47
r151 6 56 91 $w=1.7e-07 $l=2.755e-07 $layer=licon1_NDIFF $count=2 $X=4.62
+ $Y=0.325 $X2=4.84 $Y2=0.45
r152 5 49 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=3.68
+ $Y=0.325 $X2=3.82 $Y2=0.45
r153 4 42 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.74
+ $Y=0.325 $X2=2.88 $Y2=0.47
r154 3 36 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.88
+ $Y=0.325 $X2=2.02 $Y2=0.47
r155 2 30 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.02
+ $Y=0.325 $X2=1.16 $Y2=0.47
r156 1 24 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.175
+ $Y=0.325 $X2=0.3 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_LP__O2BB2AI_4%VGND 1 2 3 4 5 6 21 25 29 33 37 39 43 46
+ 47 49 50 52 53 54 55 56 58 84 85 88 91
r135 91 92 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r136 88 89 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r137 84 85 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=9.84 $Y=0
+ $X2=9.84 $Y2=0
r138 82 85 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=7.92 $Y=0
+ $X2=9.84 $Y2=0
r139 82 92 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=7.44
+ $Y2=0
r140 81 84 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=7.92 $Y=0 $X2=9.84
+ $Y2=0
r141 81 82 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=7.92 $Y=0
+ $X2=7.92 $Y2=0
r142 79 91 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.755 $Y=0 $X2=7.59
+ $Y2=0
r143 79 81 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=7.755 $Y=0
+ $X2=7.92 $Y2=0
r144 78 92 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=7.44
+ $Y2=0
r145 77 78 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=6.48 $Y=0
+ $X2=6.48 $Y2=0
r146 74 77 187.893 $w=1.68e-07 $l=2.88e-06 $layer=LI1_cond $X=3.6 $Y=0 $X2=6.48
+ $Y2=0
r147 74 75 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=3.6 $Y=0
+ $X2=3.6 $Y2=0
r148 72 75 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r149 71 72 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r150 69 72 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r151 68 69 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r152 66 69 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r153 66 89 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r154 65 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r155 63 88 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.895 $Y=0 $X2=0.73
+ $Y2=0
r156 63 65 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.895 $Y=0 $X2=1.2
+ $Y2=0
r157 61 89 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r158 60 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r159 58 88 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.565 $Y=0 $X2=0.73
+ $Y2=0
r160 58 60 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.565 $Y=0
+ $X2=0.24 $Y2=0
r161 56 78 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=5.04 $Y=0
+ $X2=6.48 $Y2=0
r162 56 75 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=5.04 $Y=0 $X2=3.6
+ $Y2=0
r163 54 77 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=6.565 $Y=0 $X2=6.48
+ $Y2=0
r164 54 55 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.565 $Y=0 $X2=6.73
+ $Y2=0
r165 52 71 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=3.145 $Y=0 $X2=3.12
+ $Y2=0
r166 52 53 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=3.145 $Y=0 $X2=3.315
+ $Y2=0
r167 51 74 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=3.485 $Y=0 $X2=3.6
+ $Y2=0
r168 51 53 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=3.485 $Y=0 $X2=3.315
+ $Y2=0
r169 49 68 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=2.285 $Y=0
+ $X2=2.16 $Y2=0
r170 49 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.285 $Y=0 $X2=2.45
+ $Y2=0
r171 48 71 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=2.615 $Y=0
+ $X2=3.12 $Y2=0
r172 48 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.615 $Y=0 $X2=2.45
+ $Y2=0
r173 46 65 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=1.425 $Y=0 $X2=1.2
+ $Y2=0
r174 46 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.425 $Y=0 $X2=1.59
+ $Y2=0
r175 45 68 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=1.755 $Y=0
+ $X2=2.16 $Y2=0
r176 45 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.755 $Y=0 $X2=1.59
+ $Y2=0
r177 41 91 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.59 $Y=0.085
+ $X2=7.59 $Y2=0
r178 41 43 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=7.59 $Y=0.085
+ $X2=7.59 $Y2=0.45
r179 40 55 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.895 $Y=0 $X2=6.73
+ $Y2=0
r180 39 91 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.425 $Y=0 $X2=7.59
+ $Y2=0
r181 39 40 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=7.425 $Y=0
+ $X2=6.895 $Y2=0
r182 35 55 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.73 $Y=0.085
+ $X2=6.73 $Y2=0
r183 35 37 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=6.73 $Y=0.085
+ $X2=6.73 $Y2=0.58
r184 31 53 0.987631 $w=3.4e-07 $l=8.5e-08 $layer=LI1_cond $X=3.315 $Y=0.085
+ $X2=3.315 $Y2=0
r185 31 33 12.3718 $w=3.38e-07 $l=3.65e-07 $layer=LI1_cond $X=3.315 $Y=0.085
+ $X2=3.315 $Y2=0.45
r186 27 50 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.45 $Y=0.085
+ $X2=2.45 $Y2=0
r187 27 29 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=2.45 $Y=0.085
+ $X2=2.45 $Y2=0.45
r188 23 47 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.59 $Y=0.085
+ $X2=1.59 $Y2=0
r189 23 25 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=1.59 $Y=0.085
+ $X2=1.59 $Y2=0.45
r190 19 88 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=0.085
+ $X2=0.73 $Y2=0
r191 19 21 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=0.73 $Y=0.085
+ $X2=0.73 $Y2=0.45
r192 6 43 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=7.45
+ $Y=0.325 $X2=7.59 $Y2=0.45
r193 5 37 182 $w=1.7e-07 $l=3.17372e-07 $layer=licon1_NDIFF $count=1 $X=6.59
+ $Y=0.325 $X2=6.73 $Y2=0.58
r194 4 33 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=3.17
+ $Y=0.325 $X2=3.31 $Y2=0.45
r195 3 29 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=2.31
+ $Y=0.325 $X2=2.45 $Y2=0.45
r196 2 25 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=1.45
+ $Y=0.325 $X2=1.59 $Y2=0.45
r197 1 21 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=0.59
+ $Y=0.325 $X2=0.73 $Y2=0.45
.ends

.subckt PM_SKY130_FD_SC_LP__O2BB2AI_4%A_1235_65# 1 2 3 4 5 16 18 20 24 26 32 33
+ 34 38 42 48
c72 48 0 1.29702e-19 $X=8.865 $Y=0.35
c73 42 0 1.73643e-19 $X=7.155 $Y=0.955
r74 48 51 6.28605 $w=2.18e-07 $l=1.2e-07 $layer=LI1_cond $X=8.865 $Y=0.35
+ $X2=8.865 $Y2=0.47
r75 45 46 7.76364 $w=1.98e-07 $l=1.4e-07 $layer=LI1_cond $X=7.155 $Y=1.02
+ $X2=7.155 $Y2=1.16
r76 42 45 3.60455 $w=1.98e-07 $l=6.5e-08 $layer=LI1_cond $X=7.155 $Y=0.955
+ $X2=7.155 $Y2=1.02
r77 42 43 4.75232 $w=1.98e-07 $l=8.5e-08 $layer=LI1_cond $X=7.155 $Y=0.955
+ $X2=7.155 $Y2=0.87
r78 36 38 1.22229 $w=3.28e-07 $l=3.5e-08 $layer=LI1_cond $X=9.82 $Y=0.435
+ $X2=9.82 $Y2=0.47
r79 35 48 2.2496 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=8.975 $Y=0.35
+ $X2=8.865 $Y2=0.35
r80 34 36 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=9.655 $Y=0.35
+ $X2=9.82 $Y2=0.435
r81 34 35 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=9.655 $Y=0.35
+ $X2=8.975 $Y2=0.35
r82 32 48 2.2496 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=8.755 $Y=0.35
+ $X2=8.865 $Y2=0.35
r83 32 33 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=8.755 $Y=0.35
+ $X2=8.115 $Y2=0.35
r84 29 31 35.3158 $w=1.88e-07 $l=6.05e-07 $layer=LI1_cond $X=8.02 $Y=1.075
+ $X2=8.02 $Y2=0.47
r85 28 33 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=8.02 $Y=0.435
+ $X2=8.115 $Y2=0.35
r86 28 31 2.04306 $w=1.88e-07 $l=3.5e-08 $layer=LI1_cond $X=8.02 $Y=0.435
+ $X2=8.02 $Y2=0.47
r87 27 46 1.68994 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=7.255 $Y=1.16 $X2=7.155
+ $Y2=1.16
r88 26 29 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=7.925 $Y=1.16
+ $X2=8.02 $Y2=1.075
r89 26 27 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=7.925 $Y=1.16
+ $X2=7.255 $Y2=1.16
r90 24 43 23.3493 $w=1.88e-07 $l=4e-07 $layer=LI1_cond $X=7.16 $Y=0.47 $X2=7.16
+ $Y2=0.87
r91 21 41 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=6.395 $Y=0.955
+ $X2=6.265 $Y2=0.955
r92 20 42 1.68994 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=7.055 $Y=0.955
+ $X2=7.155 $Y2=0.955
r93 20 21 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=7.055 $Y=0.955
+ $X2=6.395 $Y2=0.955
r94 16 41 2.85134 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=6.265 $Y=0.87
+ $X2=6.265 $Y2=0.955
r95 16 18 17.7299 $w=2.58e-07 $l=4e-07 $layer=LI1_cond $X=6.265 $Y=0.87
+ $X2=6.265 $Y2=0.47
r96 5 38 91 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_NDIFF $count=2 $X=9.6
+ $Y=0.325 $X2=9.82 $Y2=0.47
r97 4 51 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=8.74
+ $Y=0.325 $X2=8.88 $Y2=0.47
r98 3 31 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=7.88
+ $Y=0.325 $X2=8.02 $Y2=0.47
r99 2 45 182 $w=1.7e-07 $l=7.61791e-07 $layer=licon1_NDIFF $count=1 $X=7.02
+ $Y=0.325 $X2=7.16 $Y2=1.02
r100 2 24 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=7.02
+ $Y=0.325 $X2=7.16 $Y2=0.47
r101 1 41 182 $w=1.7e-07 $l=6.89674e-07 $layer=licon1_NDIFF $count=1 $X=6.175
+ $Y=0.325 $X2=6.3 $Y2=0.955
r102 1 18 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=6.175
+ $Y=0.325 $X2=6.3 $Y2=0.47
.ends

