* File: sky130_fd_sc_lp__a41oi_2.pex.spice
* Created: Wed Sep  2 09:29:41 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A41OI_2%B1 1 3 6 8 10 13 15 17 30
c45 6 0 3.03319e-20 $X=0.855 $Y=2.465
r46 29 30 53.3327 $w=3.3e-07 $l=3.05e-07 $layer=POLY_cond $X=0.98 $Y=1.35
+ $X2=1.285 $Y2=1.35
r47 28 29 21.8577 $w=3.3e-07 $l=1.25e-07 $layer=POLY_cond $X=0.855 $Y=1.35
+ $X2=0.98 $Y2=1.35
r48 26 28 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=0.64 $Y=1.35
+ $X2=0.855 $Y2=1.35
r49 23 26 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=0.55 $Y=1.35 $X2=0.64
+ $Y2=1.35
r50 17 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.64
+ $Y=1.35 $X2=0.64 $Y2=1.35
r51 15 17 8.85984 $w=5.38e-07 $l=4e-07 $layer=LI1_cond $X=0.24 $Y=1.48 $X2=0.64
+ $Y2=1.48
r52 11 30 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.285 $Y=1.515
+ $X2=1.285 $Y2=1.35
r53 11 13 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=1.285 $Y=1.515
+ $X2=1.285 $Y2=2.465
r54 8 29 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.98 $Y=1.185
+ $X2=0.98 $Y2=1.35
r55 8 10 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.98 $Y=1.185
+ $X2=0.98 $Y2=0.655
r56 4 28 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.855 $Y=1.515
+ $X2=0.855 $Y2=1.35
r57 4 6 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=0.855 $Y=1.515
+ $X2=0.855 $Y2=2.465
r58 1 23 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.55 $Y=1.185
+ $X2=0.55 $Y2=1.35
r59 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.55 $Y=1.185 $X2=0.55
+ $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__A41OI_2%A1 3 5 7 10 12 14 15 16 22 24
c60 24 0 2.48304e-19 $X=2.31 $Y=1.46
c61 12 0 8.67364e-20 $X=2.38 $Y=1.295
c62 3 0 1.56476e-19 $X=1.715 $Y=2.465
r63 24 25 10.7111 $w=3.15e-07 $l=7e-08 $layer=POLY_cond $X=2.31 $Y=1.46 $X2=2.38
+ $Y2=1.46
r64 23 24 55.0857 $w=3.15e-07 $l=3.6e-07 $layer=POLY_cond $X=1.95 $Y=1.46
+ $X2=2.31 $Y2=1.46
r65 21 23 32.8984 $w=3.15e-07 $l=2.15e-07 $layer=POLY_cond $X=1.735 $Y=1.46
+ $X2=1.95 $Y2=1.46
r66 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.735
+ $Y=1.46 $X2=1.735 $Y2=1.46
r67 19 21 3.06032 $w=3.15e-07 $l=2e-08 $layer=POLY_cond $X=1.715 $Y=1.46
+ $X2=1.735 $Y2=1.46
r68 16 22 1.58461 $w=3.98e-07 $l=5.5e-08 $layer=LI1_cond $X=1.68 $Y=1.41
+ $X2=1.735 $Y2=1.41
r69 15 16 13.8293 $w=3.98e-07 $l=4.8e-07 $layer=LI1_cond $X=1.2 $Y=1.41 $X2=1.68
+ $Y2=1.41
r70 12 25 20.1192 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.38 $Y=1.295
+ $X2=2.38 $Y2=1.46
r71 12 14 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.38 $Y=1.295
+ $X2=2.38 $Y2=0.765
r72 8 24 20.1192 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.31 $Y=1.625
+ $X2=2.31 $Y2=1.46
r73 8 10 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=2.31 $Y=1.625
+ $X2=2.31 $Y2=2.465
r74 5 23 20.1192 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.95 $Y=1.295
+ $X2=1.95 $Y2=1.46
r75 5 7 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.95 $Y=1.295 $X2=1.95
+ $Y2=0.765
r76 1 19 20.1192 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.715 $Y=1.625
+ $X2=1.715 $Y2=1.46
r77 1 3 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=1.715 $Y=1.625
+ $X2=1.715 $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__A41OI_2%A2 3 7 11 15 17 22 23 24
c53 24 0 1.94313e-19 $X=3.6 $Y=1.665
c54 22 0 1.29864e-19 $X=3.675 $Y=1.51
r55 28 29 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.52
+ $Y=1.51 $X2=3.52 $Y2=1.51
r56 24 29 2.27643 $w=4.03e-07 $l=8e-08 $layer=LI1_cond $X=3.6 $Y=1.627 $X2=3.52
+ $Y2=1.627
r57 23 29 11.3822 $w=4.03e-07 $l=4e-07 $layer=LI1_cond $X=3.12 $Y=1.627 $X2=3.52
+ $Y2=1.627
r58 22 28 27.1035 $w=3.3e-07 $l=1.55e-07 $layer=POLY_cond $X=3.675 $Y=1.51
+ $X2=3.52 $Y2=1.51
r59 20 21 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=2.81 $Y=1.51
+ $X2=3.24 $Y2=1.51
r60 18 20 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=2.74 $Y=1.51 $X2=2.81
+ $Y2=1.51
r61 17 28 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=3.315 $Y=1.51
+ $X2=3.52 $Y2=1.51
r62 17 21 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=3.315 $Y=1.51
+ $X2=3.24 $Y2=1.51
r63 13 22 32.1775 $w=3.3e-07 $l=1.98997e-07 $layer=POLY_cond $X=3.75 $Y=1.675
+ $X2=3.675 $Y2=1.51
r64 13 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.75 $Y=1.675
+ $X2=3.75 $Y2=2.465
r65 9 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.24 $Y=1.345
+ $X2=3.24 $Y2=1.51
r66 9 11 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=3.24 $Y=1.345
+ $X2=3.24 $Y2=0.765
r67 5 20 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.81 $Y=1.345
+ $X2=2.81 $Y2=1.51
r68 5 7 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=2.81 $Y=1.345 $X2=2.81
+ $Y2=0.765
r69 1 18 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.74 $Y=1.675
+ $X2=2.74 $Y2=1.51
r70 1 3 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.74 $Y=1.675 $X2=2.74
+ $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__A41OI_2%A3 3 5 7 8 10 13 15 20 29
c63 20 0 1.29864e-19 $X=4.56 $Y=1.295
c64 13 0 2.55151e-20 $X=4.78 $Y=2.465
c65 8 0 7.56076e-20 $X=4.78 $Y=1.295
c66 3 0 8.00027e-20 $X=4.18 $Y=2.465
r67 27 29 27.9778 $w=3.3e-07 $l=1.6e-07 $layer=POLY_cond $X=4.62 $Y=1.46
+ $X2=4.78 $Y2=1.46
r68 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.62
+ $Y=1.46 $X2=4.62 $Y2=1.46
r69 25 27 47.2125 $w=3.3e-07 $l=2.7e-07 $layer=POLY_cond $X=4.35 $Y=1.46
+ $X2=4.62 $Y2=1.46
r70 20 28 2.3537 $w=3.11e-07 $l=6e-08 $layer=LI1_cond $X=4.56 $Y=1.377 $X2=4.62
+ $Y2=1.377
r71 18 25 13.9889 $w=3.3e-07 $l=8e-08 $layer=POLY_cond $X=4.27 $Y=1.46 $X2=4.35
+ $Y2=1.46
r72 18 22 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=4.27 $Y=1.46 $X2=4.18
+ $Y2=1.46
r73 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.27
+ $Y=1.46 $X2=4.27 $Y2=1.46
r74 15 20 8.76629 $w=3.11e-07 $l=1.9718e-07 $layer=LI1_cond $X=4.4 $Y=1.46
+ $X2=4.56 $Y2=1.377
r75 15 17 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=4.4 $Y=1.46 $X2=4.27
+ $Y2=1.46
r76 11 29 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.78 $Y=1.625
+ $X2=4.78 $Y2=1.46
r77 11 13 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=4.78 $Y=1.625
+ $X2=4.78 $Y2=2.465
r78 8 29 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.78 $Y=1.295
+ $X2=4.78 $Y2=1.46
r79 8 10 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=4.78 $Y=1.295
+ $X2=4.78 $Y2=0.765
r80 5 25 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.35 $Y=1.295
+ $X2=4.35 $Y2=1.46
r81 5 7 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=4.35 $Y=1.295 $X2=4.35
+ $Y2=0.765
r82 1 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.18 $Y=1.625
+ $X2=4.18 $Y2=1.46
r83 1 3 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=4.18 $Y=1.625 $X2=4.18
+ $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__A41OI_2%A4 3 7 11 15 17 18 26
c41 18 0 2.55151e-20 $X=6 $Y=1.665
r42 24 26 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=5.425 $Y=1.51
+ $X2=5.64 $Y2=1.51
r43 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.425
+ $Y=1.51 $X2=5.425 $Y2=1.51
r44 21 24 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=5.21 $Y=1.51
+ $X2=5.425 $Y2=1.51
r45 17 18 17.0207 $w=3.23e-07 $l=4.8e-07 $layer=LI1_cond $X=5.52 $Y=1.587 $X2=6
+ $Y2=1.587
r46 17 25 3.36868 $w=3.23e-07 $l=9.5e-08 $layer=LI1_cond $X=5.52 $Y=1.587
+ $X2=5.425 $Y2=1.587
r47 13 26 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.64 $Y=1.675
+ $X2=5.64 $Y2=1.51
r48 13 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=5.64 $Y=1.675
+ $X2=5.64 $Y2=2.465
r49 9 26 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.64 $Y=1.345
+ $X2=5.64 $Y2=1.51
r50 9 11 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=5.64 $Y=1.345
+ $X2=5.64 $Y2=0.765
r51 5 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.21 $Y=1.675
+ $X2=5.21 $Y2=1.51
r52 5 7 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=5.21 $Y=1.675 $X2=5.21
+ $Y2=2.465
r53 1 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.21 $Y=1.345
+ $X2=5.21 $Y2=1.51
r54 1 3 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=5.21 $Y=1.345 $X2=5.21
+ $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_LP__A41OI_2%A_103_367# 1 2 3 4 5 6 19 21 23 25 26 27 31
+ 33 38 41 43 44 45 47 49 51 53 62 63
c97 62 0 2.90469e-19 $X=2.525 $Y=2.205
c98 26 0 3.03319e-20 $X=1.535 $Y=2.885
r99 66 67 1.44094 $w=2.54e-07 $l=3e-08 $layer=LI1_cond $X=4.96 $Y=1.98 $X2=4.96
+ $Y2=2.01
r100 64 66 8.64567 $w=2.54e-07 $l=1.8e-07 $layer=LI1_cond $X=4.96 $Y=1.8
+ $X2=4.96 $Y2=1.98
r101 51 69 2.85134 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=5.89 $Y=2.095
+ $X2=5.89 $Y2=2.01
r102 51 53 36.1247 $w=2.58e-07 $l=8.15e-07 $layer=LI1_cond $X=5.89 $Y=2.095
+ $X2=5.89 $Y2=2.91
r103 50 67 3.08766 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=5.09 $Y=2.01
+ $X2=4.96 $Y2=2.01
r104 49 69 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=5.76 $Y=2.01
+ $X2=5.89 $Y2=2.01
r105 49 50 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.76 $Y=2.01
+ $X2=5.09 $Y2=2.01
r106 45 67 3.98846 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=4.96 $Y=2.095
+ $X2=4.96 $Y2=2.01
r107 45 47 15.5137 $w=2.58e-07 $l=3.5e-07 $layer=LI1_cond $X=4.96 $Y=2.095
+ $X2=4.96 $Y2=2.445
r108 43 64 3.08766 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=4.83 $Y=1.8 $X2=4.96
+ $Y2=1.8
r109 43 44 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=4.83 $Y=1.8 $X2=4.13
+ $Y2=1.8
r110 39 63 4.11778 $w=2.67e-07 $l=1.06925e-07 $layer=LI1_cond $X=4 $Y=2.325
+ $X2=3.992 $Y2=2.222
r111 39 41 5.31897 $w=2.58e-07 $l=1.2e-07 $layer=LI1_cond $X=4 $Y=2.325 $X2=4
+ $Y2=2.445
r112 36 63 4.11778 $w=2.67e-07 $l=1.02e-07 $layer=LI1_cond $X=3.992 $Y=2.12
+ $X2=3.992 $Y2=2.222
r113 36 38 5.86698 $w=2.73e-07 $l=1.4e-07 $layer=LI1_cond $X=3.992 $Y=2.12
+ $X2=3.992 $Y2=1.98
r114 35 44 7.32204 $w=1.7e-07 $l=1.75425e-07 $layer=LI1_cond $X=3.992 $Y=1.885
+ $X2=4.13 $Y2=1.8
r115 35 38 3.98117 $w=2.73e-07 $l=9.5e-08 $layer=LI1_cond $X=3.992 $Y=1.885
+ $X2=3.992 $Y2=1.98
r116 34 62 8.03064 $w=1.87e-07 $l=1.65e-07 $layer=LI1_cond $X=2.69 $Y=2.222
+ $X2=2.525 $Y2=2.222
r117 33 63 2.31614 $w=2.05e-07 $l=1.37e-07 $layer=LI1_cond $X=3.855 $Y=2.222
+ $X2=3.992 $Y2=2.222
r118 33 34 63.0288 $w=2.03e-07 $l=1.165e-06 $layer=LI1_cond $X=3.855 $Y=2.222
+ $X2=2.69 $Y2=2.222
r119 29 62 0.588983 $w=3.3e-07 $l=1.03e-07 $layer=LI1_cond $X=2.525 $Y=2.325
+ $X2=2.525 $Y2=2.222
r120 29 31 21.4773 $w=3.28e-07 $l=6.15e-07 $layer=LI1_cond $X=2.525 $Y=2.325
+ $X2=2.525 $Y2=2.94
r121 28 60 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.665 $Y=2.205
+ $X2=1.535 $Y2=2.205
r122 27 62 8.03064 $w=1.87e-07 $l=1.73292e-07 $layer=LI1_cond $X=2.36 $Y=2.205
+ $X2=2.525 $Y2=2.222
r123 27 28 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=2.36 $Y=2.205
+ $X2=1.665 $Y2=2.205
r124 26 58 3.08262 $w=2.6e-07 $l=1.11131e-07 $layer=LI1_cond $X=1.535 $Y=2.885
+ $X2=1.5 $Y2=2.98
r125 25 60 2.85134 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=1.535 $Y=2.29
+ $X2=1.535 $Y2=2.205
r126 25 26 26.3732 $w=2.58e-07 $l=5.95e-07 $layer=LI1_cond $X=1.535 $Y=2.29
+ $X2=1.535 $Y2=2.885
r127 24 56 4.20357 $w=1.8e-07 $l=1.3e-07 $layer=LI1_cond $X=0.735 $Y=2.985
+ $X2=0.605 $Y2=2.985
r128 23 58 4.03111 $w=1.8e-07 $l=1.67481e-07 $layer=LI1_cond $X=1.335 $Y=2.985
+ $X2=1.5 $Y2=2.98
r129 23 24 36.9697 $w=1.78e-07 $l=6e-07 $layer=LI1_cond $X=1.335 $Y=2.985
+ $X2=0.735 $Y2=2.985
r130 19 56 2.91016 $w=2.6e-07 $l=9e-08 $layer=LI1_cond $X=0.605 $Y=2.895
+ $X2=0.605 $Y2=2.985
r131 19 21 35.903 $w=2.58e-07 $l=8.1e-07 $layer=LI1_cond $X=0.605 $Y=2.895
+ $X2=0.605 $Y2=2.085
r132 6 69 400 $w=1.7e-07 $l=3.17372e-07 $layer=licon1_PDIFF $count=1 $X=5.715
+ $Y=1.835 $X2=5.855 $Y2=2.09
r133 6 53 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=5.715
+ $Y=1.835 $X2=5.855 $Y2=2.91
r134 5 66 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=4.855
+ $Y=1.835 $X2=4.995 $Y2=1.98
r135 5 47 300 $w=1.7e-07 $l=6.76387e-07 $layer=licon1_PDIFF $count=2 $X=4.855
+ $Y=1.835 $X2=4.995 $Y2=2.445
r136 4 41 300 $w=1.7e-07 $l=6.76387e-07 $layer=licon1_PDIFF $count=2 $X=3.825
+ $Y=1.835 $X2=3.965 $Y2=2.445
r137 4 38 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=3.825
+ $Y=1.835 $X2=3.965 $Y2=1.98
r138 3 62 400 $w=1.7e-07 $l=4.34396e-07 $layer=licon1_PDIFF $count=1 $X=2.385
+ $Y=1.835 $X2=2.525 $Y2=2.205
r139 3 31 400 $w=1.7e-07 $l=1.17291e-06 $layer=licon1_PDIFF $count=1 $X=2.385
+ $Y=1.835 $X2=2.525 $Y2=2.94
r140 2 60 300 $w=1.7e-07 $l=5.15267e-07 $layer=licon1_PDIFF $count=2 $X=1.36
+ $Y=1.835 $X2=1.5 $Y2=2.285
r141 2 58 600 $w=1.7e-07 $l=1.20297e-06 $layer=licon1_PDIFF $count=1 $X=1.36
+ $Y=1.835 $X2=1.5 $Y2=2.97
r142 1 56 400 $w=1.7e-07 $l=1.13578e-06 $layer=licon1_PDIFF $count=1 $X=0.515
+ $Y=1.835 $X2=0.64 $Y2=2.91
r143 1 21 400 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_PDIFF $count=1 $X=0.515
+ $Y=1.835 $X2=0.64 $Y2=2.085
.ends

.subckt PM_SKY130_FD_SC_LP__A41OI_2%Y 1 2 3 12 14 15 18 23 27 29 33 34 38
r63 33 38 7.96408 $w=5.23e-07 $l=9e-08 $layer=LI1_cond $X=2.16 $Y=1.687 $X2=2.07
+ $Y2=1.687
r64 31 32 3.51899 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=2.165 $Y=0.955
+ $X2=2.165 $Y2=1.04
r65 29 31 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.165 $Y=0.68
+ $X2=2.165 $Y2=0.955
r66 27 32 0.886495 $w=2.58e-07 $l=2e-08 $layer=LI1_cond $X=2.2 $Y=1.06 $X2=2.2
+ $Y2=1.04
r67 25 34 10.0243 $w=5.23e-07 $l=4.4e-07 $layer=LI1_cond $X=2.2 $Y=1.687
+ $X2=2.64 $Y2=1.687
r68 25 33 0.911298 $w=5.23e-07 $l=4e-08 $layer=LI1_cond $X=2.2 $Y=1.687 $X2=2.16
+ $Y2=1.687
r69 25 27 16.1785 $w=2.58e-07 $l=3.65e-07 $layer=LI1_cond $X=2.2 $Y=1.425
+ $X2=2.2 $Y2=1.06
r70 23 38 54.4759 $w=1.68e-07 $l=8.35e-07 $layer=LI1_cond $X=1.235 $Y=1.865
+ $X2=2.07 $Y2=1.865
r71 18 20 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=1.07 $Y=1.96
+ $X2=1.07 $Y2=2.64
r72 16 23 17.4739 $w=1.11e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.07 $Y=1.95
+ $X2=1.235 $Y2=1.865
r73 16 18 0.349225 $w=3.28e-07 $l=1e-08 $layer=LI1_cond $X=1.07 $Y=1.95 $X2=1.07
+ $Y2=1.96
r74 14 31 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2 $Y=0.955 $X2=2.165
+ $Y2=0.955
r75 14 15 74.3743 $w=1.68e-07 $l=1.14e-06 $layer=LI1_cond $X=2 $Y=0.955 $X2=0.86
+ $Y2=0.955
r76 10 15 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=0.765 $Y=0.87
+ $X2=0.86 $Y2=0.955
r77 10 12 26.2679 $w=1.88e-07 $l=4.5e-07 $layer=LI1_cond $X=0.765 $Y=0.87
+ $X2=0.765 $Y2=0.42
r78 3 20 400 $w=1.7e-07 $l=8.72195e-07 $layer=licon1_PDIFF $count=1 $X=0.93
+ $Y=1.835 $X2=1.07 $Y2=2.64
r79 3 18 400 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=0.93
+ $Y=1.835 $X2=1.07 $Y2=1.96
r80 2 29 182 $w=1.7e-07 $l=3.98905e-07 $layer=licon1_NDIFF $count=1 $X=2.025
+ $Y=0.345 $X2=2.165 $Y2=0.68
r81 2 27 182 $w=1.7e-07 $l=7.81873e-07 $layer=licon1_NDIFF $count=1 $X=2.025
+ $Y=0.345 $X2=2.165 $Y2=1.06
r82 1 12 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=0.625
+ $Y=0.235 $X2=0.765 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__A41OI_2%VPWR 1 2 3 4 15 19 25 28 29 31 32 33 42 46
+ 56 57 60 67
r81 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r82 63 64 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r83 60 63 10.2521 $w=8.38e-07 $l=7.2e-07 $layer=LI1_cond $X=3.28 $Y=2.61
+ $X2=3.28 $Y2=3.33
r84 56 57 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r85 54 57 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=3.33 $X2=6
+ $Y2=3.33
r86 54 68 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=4.56 $Y2=3.33
r87 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r88 51 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.645 $Y=3.33
+ $X2=4.48 $Y2=3.33
r89 51 53 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=4.645 $Y=3.33
+ $X2=5.04 $Y2=3.33
r90 50 68 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r91 50 64 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.6 $Y2=3.33
r92 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r93 47 63 10.5369 $w=1.7e-07 $l=4.2e-07 $layer=LI1_cond $X=3.7 $Y=3.33 $X2=3.28
+ $Y2=3.33
r94 47 49 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=3.7 $Y=3.33 $X2=4.08
+ $Y2=3.33
r95 46 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.315 $Y=3.33
+ $X2=4.48 $Y2=3.33
r96 46 49 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=4.315 $Y=3.33
+ $X2=4.08 $Y2=3.33
r97 44 45 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r98 42 63 10.5369 $w=1.7e-07 $l=4.2e-07 $layer=LI1_cond $X=2.86 $Y=3.33 $X2=3.28
+ $Y2=3.33
r99 42 44 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=2.86 $Y=3.33
+ $X2=2.64 $Y2=3.33
r100 41 45 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r101 40 41 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r102 37 41 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.68 $Y2=3.33
r103 36 40 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=0.24 $Y=3.33
+ $X2=1.68 $Y2=3.33
r104 36 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r105 33 64 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r106 33 45 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.64 $Y2=3.33
r107 31 53 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=5.26 $Y=3.33
+ $X2=5.04 $Y2=3.33
r108 31 32 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.26 $Y=3.33
+ $X2=5.425 $Y2=3.33
r109 30 56 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=5.59 $Y=3.33 $X2=6
+ $Y2=3.33
r110 30 32 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.59 $Y=3.33
+ $X2=5.425 $Y2=3.33
r111 28 40 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=1.845 $Y=3.33
+ $X2=1.68 $Y2=3.33
r112 28 29 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.845 $Y=3.33
+ $X2=2.01 $Y2=3.33
r113 27 44 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=2.175 $Y=3.33
+ $X2=2.64 $Y2=3.33
r114 27 29 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.175 $Y=3.33
+ $X2=2.01 $Y2=3.33
r115 23 32 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.425 $Y=3.245
+ $X2=5.425 $Y2=3.33
r116 23 25 30.0334 $w=3.28e-07 $l=8.6e-07 $layer=LI1_cond $X=5.425 $Y=3.245
+ $X2=5.425 $Y2=2.385
r117 19 22 28.2872 $w=3.28e-07 $l=8.1e-07 $layer=LI1_cond $X=4.48 $Y=2.14
+ $X2=4.48 $Y2=2.95
r118 17 67 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.48 $Y=3.245
+ $X2=4.48 $Y2=3.33
r119 17 22 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=4.48 $Y=3.245
+ $X2=4.48 $Y2=2.95
r120 13 29 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.01 $Y=3.245
+ $X2=2.01 $Y2=3.33
r121 13 15 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=2.01 $Y=3.245
+ $X2=2.01 $Y2=2.57
r122 4 25 300 $w=1.7e-07 $l=6.16036e-07 $layer=licon1_PDIFF $count=2 $X=5.285
+ $Y=1.835 $X2=5.425 $Y2=2.385
r123 3 22 400 $w=1.7e-07 $l=1.22233e-06 $layer=licon1_PDIFF $count=1 $X=4.255
+ $Y=1.835 $X2=4.48 $Y2=2.95
r124 3 19 400 $w=1.7e-07 $l=4.02057e-07 $layer=licon1_PDIFF $count=1 $X=4.255
+ $Y=1.835 $X2=4.48 $Y2=2.14
r125 2 60 150 $w=1.7e-07 $l=1.07639e-06 $layer=licon1_PDIFF $count=4 $X=2.815
+ $Y=1.835 $X2=3.535 $Y2=2.61
r126 1 15 300 $w=1.7e-07 $l=8.3781e-07 $layer=licon1_PDIFF $count=2 $X=1.79
+ $Y=1.835 $X2=2.01 $Y2=2.57
.ends

.subckt PM_SKY130_FD_SC_LP__A41OI_2%VGND 1 2 3 10 12 16 20 23 24 25 27 40 41 47
r64 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r65 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r66 40 41 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=0 $X2=6 $Y2=0
r67 38 41 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=6
+ $Y2=0
r68 37 38 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r69 35 48 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r70 34 37 219.209 $w=1.68e-07 $l=3.36e-06 $layer=LI1_cond $X=1.68 $Y=0 $X2=5.04
+ $Y2=0
r71 34 35 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r72 32 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.36 $Y=0 $X2=1.195
+ $Y2=0
r73 32 34 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=1.36 $Y=0 $X2=1.68
+ $Y2=0
r74 31 48 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r75 31 45 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r76 30 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r77 28 44 4.62272 $w=1.7e-07 $l=2.5e-07 $layer=LI1_cond $X=0.5 $Y=0 $X2=0.25
+ $Y2=0
r78 28 30 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=0.5 $Y=0 $X2=0.72
+ $Y2=0
r79 27 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.03 $Y=0 $X2=1.195
+ $Y2=0
r80 27 30 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=1.03 $Y=0 $X2=0.72
+ $Y2=0
r81 25 38 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=3.12 $Y=0 $X2=5.04
+ $Y2=0
r82 25 35 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=3.12 $Y=0 $X2=1.68
+ $Y2=0
r83 23 37 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=5.26 $Y=0 $X2=5.04
+ $Y2=0
r84 23 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.26 $Y=0 $X2=5.425
+ $Y2=0
r85 22 40 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=5.59 $Y=0 $X2=6
+ $Y2=0
r86 22 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.59 $Y=0 $X2=5.425
+ $Y2=0
r87 18 24 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.425 $Y=0.085
+ $X2=5.425 $Y2=0
r88 18 20 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=5.425 $Y=0.085
+ $X2=5.425 $Y2=0.47
r89 14 47 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.195 $Y=0.085
+ $X2=1.195 $Y2=0
r90 14 16 17.112 $w=3.28e-07 $l=4.9e-07 $layer=LI1_cond $X=1.195 $Y=0.085
+ $X2=1.195 $Y2=0.575
r91 10 44 3.14345 $w=3.3e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.335 $Y=0.085
+ $X2=0.25 $Y2=0
r92 10 12 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.335 $Y=0.085
+ $X2=0.335 $Y2=0.38
r93 3 20 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=5.285
+ $Y=0.345 $X2=5.425 $Y2=0.47
r94 2 16 182 $w=1.7e-07 $l=4.0398e-07 $layer=licon1_NDIFF $count=1 $X=1.055
+ $Y=0.235 $X2=1.195 $Y2=0.575
r95 1 12 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.21
+ $Y=0.235 $X2=0.335 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_LP__A41OI_2%A_318_69# 1 2 3 10 16 17 20 22
r39 22 25 8.02594 $w=2.78e-07 $l=1.95e-07 $layer=LI1_cond $X=1.69 $Y=0.34
+ $X2=1.69 $Y2=0.535
r40 18 20 14.1436 $w=3.28e-07 $l=4.05e-07 $layer=LI1_cond $X=3.525 $Y=1.085
+ $X2=3.525 $Y2=0.68
r41 16 18 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.36 $Y=1.17
+ $X2=3.525 $Y2=1.085
r42 16 17 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.36 $Y=1.17
+ $X2=2.69 $Y2=1.17
r43 13 17 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=2.595 $Y=1.085
+ $X2=2.69 $Y2=1.17
r44 13 15 34.7321 $w=1.88e-07 $l=5.95e-07 $layer=LI1_cond $X=2.595 $Y=1.085
+ $X2=2.595 $Y2=0.49
r45 12 15 3.79426 $w=1.88e-07 $l=6.5e-08 $layer=LI1_cond $X=2.595 $Y=0.425
+ $X2=2.595 $Y2=0.49
r46 11 22 3.65648 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=1.83 $Y=0.34 $X2=1.69
+ $Y2=0.34
r47 10 12 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=2.5 $Y=0.34
+ $X2=2.595 $Y2=0.425
r48 10 11 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.5 $Y=0.34 $X2=1.83
+ $Y2=0.34
r49 3 20 91 $w=1.7e-07 $l=4.27288e-07 $layer=licon1_NDIFF $count=2 $X=3.315
+ $Y=0.345 $X2=3.525 $Y2=0.68
r50 2 15 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.455
+ $Y=0.345 $X2=2.595 $Y2=0.49
r51 1 25 182 $w=1.7e-07 $l=2.44643e-07 $layer=licon1_NDIFF $count=1 $X=1.59
+ $Y=0.345 $X2=1.715 $Y2=0.535
.ends

.subckt PM_SKY130_FD_SC_LP__A41OI_2%A_577_69# 1 2 9 11 12 13
c31 12 0 8.67364e-20 $X=3.19 $Y=0.34
c32 11 0 7.56076e-20 $X=4.4 $Y=0.34
r33 13 16 8.20679 $w=3.28e-07 $l=2.35e-07 $layer=LI1_cond $X=4.565 $Y=0.34
+ $X2=4.565 $Y2=0.575
r34 11 13 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.4 $Y=0.34
+ $X2=4.565 $Y2=0.34
r35 11 12 78.9412 $w=1.68e-07 $l=1.21e-06 $layer=LI1_cond $X=4.4 $Y=0.34
+ $X2=3.19 $Y2=0.34
r36 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.025 $Y=0.425
+ $X2=3.19 $Y2=0.34
r37 7 9 1.57151 $w=3.28e-07 $l=4.5e-08 $layer=LI1_cond $X=3.025 $Y=0.425
+ $X2=3.025 $Y2=0.47
r38 2 16 182 $w=1.7e-07 $l=2.91719e-07 $layer=licon1_NDIFF $count=1 $X=4.425
+ $Y=0.345 $X2=4.565 $Y2=0.575
r39 1 9 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=2.885
+ $Y=0.345 $X2=3.025 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_LP__A41OI_2%A_788_69# 1 2 3 10 14 16 20 23 29
r44 29 30 8.61957 $w=1.84e-07 $l=1.3e-07 $layer=LI1_cond $X=4.995 $Y=1.04
+ $X2=4.995 $Y2=1.17
r45 27 29 5.63587 $w=1.84e-07 $l=8.5e-08 $layer=LI1_cond $X=4.995 $Y=0.955
+ $X2=4.995 $Y2=1.04
r46 23 25 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=4.065 $Y=0.68
+ $X2=4.065 $Y2=0.955
r47 18 20 26.3732 $w=2.58e-07 $l=5.95e-07 $layer=LI1_cond $X=5.89 $Y=1.085
+ $X2=5.89 $Y2=0.49
r48 17 30 1.1945 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=5.09 $Y=1.17 $X2=4.995
+ $Y2=1.17
r49 16 18 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=5.76 $Y=1.17
+ $X2=5.89 $Y2=1.085
r50 16 17 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.76 $Y=1.17
+ $X2=5.09 $Y2=1.17
r51 12 27 5.45789 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=4.995 $Y=0.87
+ $X2=4.995 $Y2=0.955
r52 12 14 22.1818 $w=1.88e-07 $l=3.8e-07 $layer=LI1_cond $X=4.995 $Y=0.87
+ $X2=4.995 $Y2=0.49
r53 11 25 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.23 $Y=0.955
+ $X2=4.065 $Y2=0.955
r54 10 27 1.1945 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=4.9 $Y=0.955 $X2=4.995
+ $Y2=0.955
r55 10 11 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.9 $Y=0.955
+ $X2=4.23 $Y2=0.955
r56 3 20 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.715
+ $Y=0.345 $X2=5.855 $Y2=0.49
r57 2 29 182 $w=1.7e-07 $l=7.61791e-07 $layer=licon1_NDIFF $count=1 $X=4.855
+ $Y=0.345 $X2=4.995 $Y2=1.04
r58 2 14 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=4.855
+ $Y=0.345 $X2=4.995 $Y2=0.49
r59 1 23 91 $w=1.7e-07 $l=3.92556e-07 $layer=licon1_NDIFF $count=2 $X=3.94
+ $Y=0.345 $X2=4.065 $Y2=0.68
.ends

