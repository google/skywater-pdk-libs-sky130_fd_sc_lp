* File: sky130_fd_sc_lp__o22ai_1.pex.spice
* Created: Wed Sep  2 10:20:35 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O22AI_1%B1 1 3 6 8 9 16
r27 13 16 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=0.27 $Y=1.46
+ $X2=0.475 $Y2=1.46
r28 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=1.46 $X2=0.27 $Y2=1.46
r29 9 14 8.75003 $w=2.68e-07 $l=2.05e-07 $layer=LI1_cond $X=0.22 $Y=1.665
+ $X2=0.22 $Y2=1.46
r30 8 14 7.04271 $w=2.68e-07 $l=1.65e-07 $layer=LI1_cond $X=0.22 $Y=1.295
+ $X2=0.22 $Y2=1.46
r31 4 16 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=1.625
+ $X2=0.475 $Y2=1.46
r32 4 6 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=0.475 $Y=1.625
+ $X2=0.475 $Y2=2.465
r33 1 16 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=1.295
+ $X2=0.475 $Y2=1.46
r34 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.475 $Y=1.295
+ $X2=0.475 $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_LP__O22AI_1%B2 3 7 9 12
c36 3 0 1.42087e-19 $X=0.835 $Y=2.465
r37 12 15 46.504 $w=3.55e-07 $l=1.65e-07 $layer=POLY_cond $X=0.937 $Y=1.51
+ $X2=0.937 $Y2=1.675
r38 12 14 46.504 $w=3.55e-07 $l=1.65e-07 $layer=POLY_cond $X=0.937 $Y=1.51
+ $X2=0.937 $Y2=1.345
r39 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.95
+ $Y=1.51 $X2=0.95 $Y2=1.51
r40 9 13 7.11385 $w=4.03e-07 $l=2.5e-07 $layer=LI1_cond $X=1.2 $Y=1.547 $X2=0.95
+ $Y2=1.547
r41 7 14 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=0.905 $Y=0.765
+ $X2=0.905 $Y2=1.345
r42 3 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=0.835 $Y=2.465
+ $X2=0.835 $Y2=1.675
.ends

.subckt PM_SKY130_FD_SC_LP__O22AI_1%A2 1 3 6 8 9 17
c37 8 0 1.42087e-19 $X=1.68 $Y=1.295
c38 1 0 1.85841e-19 $X=1.4 $Y=1.295
r39 15 17 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=1.54 $Y=1.46 $X2=1.63
+ $Y2=1.46
r40 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.54
+ $Y=1.46 $X2=1.54 $Y2=1.46
r41 12 15 24.4806 $w=3.3e-07 $l=1.4e-07 $layer=POLY_cond $X=1.4 $Y=1.46 $X2=1.54
+ $Y2=1.46
r42 9 16 7.62099 $w=3.08e-07 $l=2.05e-07 $layer=LI1_cond $X=1.61 $Y=1.665
+ $X2=1.61 $Y2=1.46
r43 8 16 6.13397 $w=3.08e-07 $l=1.65e-07 $layer=LI1_cond $X=1.61 $Y=1.295
+ $X2=1.61 $Y2=1.46
r44 4 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.63 $Y=1.625
+ $X2=1.63 $Y2=1.46
r45 4 6 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=1.63 $Y=1.625 $X2=1.63
+ $Y2=2.465
r46 1 12 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.4 $Y=1.295 $X2=1.4
+ $Y2=1.46
r47 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.4 $Y=1.295 $X2=1.4
+ $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_LP__O22AI_1%A1 3 7 8 10 12 14 21
r30 21 22 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.5 $Y=1.46
+ $X2=2.5 $Y2=1.46
r31 14 22 3.10094 $w=5.38e-07 $l=1.4e-07 $layer=LI1_cond $X=2.64 $Y=1.48 $X2=2.5
+ $Y2=1.48
r32 12 22 7.53086 $w=5.38e-07 $l=3.4e-07 $layer=LI1_cond $X=2.16 $Y=1.48 $X2=2.5
+ $Y2=1.48
r33 9 21 44.5896 $w=3.3e-07 $l=2.55e-07 $layer=POLY_cond $X=2.245 $Y=1.46
+ $X2=2.5 $Y2=1.46
r34 8 11 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.08 $Y=1.46
+ $X2=2.08 $Y2=1.625
r35 8 10 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.08 $Y=1.46
+ $X2=2.08 $Y2=1.295
r36 8 9 2.83073 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.08 $Y=1.46
+ $X2=2.245 $Y2=1.46
r37 7 10 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.17 $Y=0.765
+ $X2=2.17 $Y2=1.295
r38 3 11 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=1.99 $Y=2.465
+ $X2=1.99 $Y2=1.625
.ends

.subckt PM_SKY130_FD_SC_LP__O22AI_1%VPWR 1 2 7 9 15 19 21 31 32 38
r29 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r30 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r31 32 39 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r32 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r33 29 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.37 $Y=3.33
+ $X2=2.205 $Y2=3.33
r34 29 31 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=2.37 $Y=3.33 $X2=2.64
+ $Y2=3.33
r35 28 39 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r36 27 28 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r37 25 36 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r38 24 27 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.72 $Y=3.33 $X2=1.68
+ $Y2=3.33
r39 24 25 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r40 22 35 4.12789 $w=1.7e-07 $l=1.78e-07 $layer=LI1_cond $X=0.355 $Y=3.33
+ $X2=0.177 $Y2=3.33
r41 22 24 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.355 $Y=3.33
+ $X2=0.72 $Y2=3.33
r42 21 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.04 $Y=3.33
+ $X2=2.205 $Y2=3.33
r43 21 27 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=2.04 $Y=3.33
+ $X2=1.68 $Y2=3.33
r44 19 28 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=1.68 $Y2=3.33
r45 19 25 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=0.72 $Y2=3.33
r46 15 18 33.0018 $w=3.28e-07 $l=9.45e-07 $layer=LI1_cond $X=2.205 $Y=2.005
+ $X2=2.205 $Y2=2.95
r47 13 38 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.205 $Y=3.245
+ $X2=2.205 $Y2=3.33
r48 13 18 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.205 $Y=3.245
+ $X2=2.205 $Y2=2.95
r49 9 12 38.3409 $w=2.58e-07 $l=8.65e-07 $layer=LI1_cond $X=0.225 $Y=2.085
+ $X2=0.225 $Y2=2.95
r50 7 35 3.08432 $w=2.6e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.225 $Y=3.245
+ $X2=0.177 $Y2=3.33
r51 7 12 13.0758 $w=2.58e-07 $l=2.95e-07 $layer=LI1_cond $X=0.225 $Y=3.245
+ $X2=0.225 $Y2=2.95
r52 2 18 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=2.065
+ $Y=1.835 $X2=2.205 $Y2=2.95
r53 2 15 400 $w=1.7e-07 $l=2.29565e-07 $layer=licon1_PDIFF $count=1 $X=2.065
+ $Y=1.835 $X2=2.205 $Y2=2.005
r54 1 12 400 $w=1.7e-07 $l=1.17584e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.835 $X2=0.26 $Y2=2.95
r55 1 9 400 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.835 $X2=0.26 $Y2=2.085
.ends

.subckt PM_SKY130_FD_SC_LP__O22AI_1%Y 1 2 9 13 14 15 16 21 22
c31 9 0 1.85841e-19 $X=0.69 $Y=0.695
r32 21 22 12.3534 $w=1.073e-06 $l=8.5e-08 $layer=LI1_cond $X=1.062 $Y=2.015
+ $X2=1.062 $Y2=1.93
r33 16 30 1.53209 $w=1.073e-06 $l=1.35e-07 $layer=LI1_cond $X=1.062 $Y=2.775
+ $X2=1.062 $Y2=2.91
r34 15 16 4.19907 $w=1.073e-06 $l=3.7e-07 $layer=LI1_cond $X=1.062 $Y=2.405
+ $X2=1.062 $Y2=2.775
r35 14 15 4.19907 $w=1.073e-06 $l=3.7e-07 $layer=LI1_cond $X=1.062 $Y=2.035
+ $X2=1.062 $Y2=2.405
r36 14 21 0.226977 $w=1.073e-06 $l=2e-08 $layer=LI1_cond $X=1.062 $Y=2.035
+ $X2=1.062 $Y2=2.015
r37 13 22 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=0.61 $Y=1.175
+ $X2=0.61 $Y2=1.93
r38 7 13 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.69 $Y=1.01
+ $X2=0.69 $Y2=1.175
r39 7 9 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=0.69 $Y=1.01 $X2=0.69
+ $Y2=0.695
r40 2 30 200 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=3 $X=0.91
+ $Y=1.835 $X2=1.05 $Y2=2.91
r41 2 21 200 $w=1.7e-07 $l=2.4e-07 $layer=licon1_PDIFF $count=3 $X=0.91 $Y=1.835
+ $X2=1.05 $Y2=2.015
r42 1 9 91 $w=1.7e-07 $l=4.14126e-07 $layer=licon1_NDIFF $count=2 $X=0.55
+ $Y=0.345 $X2=0.69 $Y2=0.695
.ends

.subckt PM_SKY130_FD_SC_LP__O22AI_1%A_27_69# 1 2 3 12 14 15 20 21 22 24
r33 22 27 2.85134 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=2.42 $Y=0.87 $X2=2.42
+ $Y2=0.955
r34 22 24 16.8434 $w=2.58e-07 $l=3.8e-07 $layer=LI1_cond $X=2.42 $Y=0.87
+ $X2=2.42 $Y2=0.49
r35 20 27 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.29 $Y=0.955
+ $X2=2.42 $Y2=0.955
r36 20 21 65.8931 $w=1.68e-07 $l=1.01e-06 $layer=LI1_cond $X=2.29 $Y=0.955
+ $X2=1.28 $Y2=0.955
r37 17 21 7.17723 $w=1.7e-07 $l=1.65118e-07 $layer=LI1_cond $X=1.152 $Y=0.87
+ $X2=1.28 $Y2=0.955
r38 17 19 17.1737 $w=2.53e-07 $l=3.8e-07 $layer=LI1_cond $X=1.152 $Y=0.87
+ $X2=1.152 $Y2=0.49
r39 16 19 2.9376 $w=2.53e-07 $l=6.5e-08 $layer=LI1_cond $X=1.152 $Y=0.425
+ $X2=1.152 $Y2=0.49
r40 14 16 7.17723 $w=1.7e-07 $l=1.64085e-07 $layer=LI1_cond $X=1.025 $Y=0.34
+ $X2=1.152 $Y2=0.425
r41 14 15 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.025 $Y=0.34
+ $X2=0.355 $Y2=0.34
r42 10 15 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=0.225 $Y=0.425
+ $X2=0.355 $Y2=0.34
r43 10 12 2.88111 $w=2.58e-07 $l=6.5e-08 $layer=LI1_cond $X=0.225 $Y=0.425
+ $X2=0.225 $Y2=0.49
r44 3 27 182 $w=1.7e-07 $l=6.76387e-07 $layer=licon1_NDIFF $count=1 $X=2.245
+ $Y=0.345 $X2=2.385 $Y2=0.955
r45 3 24 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=2.245
+ $Y=0.345 $X2=2.385 $Y2=0.49
r46 2 19 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=0.98
+ $Y=0.345 $X2=1.12 $Y2=0.49
r47 1 12 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.345 $X2=0.26 $Y2=0.49
.ends

.subckt PM_SKY130_FD_SC_LP__O22AI_1%VGND 1 4 6 16 17 21
r25 21 24 10.2649 $w=6.68e-07 $l=5.75e-07 $layer=LI1_cond $X=1.785 $Y=0
+ $X2=1.785 $Y2=0.575
r26 21 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r27 17 22 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=1.68
+ $Y2=0
r28 16 17 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r29 14 21 9.03384 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=2.12 $Y=0 $X2=1.785
+ $Y2=0
r30 14 16 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=2.12 $Y=0 $X2=2.64
+ $Y2=0
r31 12 13 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r32 9 13 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r33 8 12 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r34 8 9 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r35 6 21 9.03384 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=1.45 $Y=0 $X2=1.785
+ $Y2=0
r36 6 12 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=1.45 $Y=0 $X2=1.2
+ $Y2=0
r37 4 22 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=1.68
+ $Y2=0
r38 4 13 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=1.2
+ $Y2=0
r39 1 24 91 $w=1.7e-07 $l=5.83781e-07 $layer=licon1_NDIFF $count=2 $X=1.475
+ $Y=0.345 $X2=1.955 $Y2=0.575
.ends

