* NGSPICE file created from sky130_fd_sc_lp__sdfstp_lp.ext - technology: sky130A

.subckt sky130_fd_sc_lp__sdfstp_lp CLK D SCD SCE SET_B VGND VNB VPB VPWR Q
M1000 a_245_406# SCD VPWR VPB phighvt w=1e+06u l=250000u
+  ad=5.7e+11p pd=5.14e+06u as=3.3553e+12p ps=2.281e+07u
M1001 a_458_406# D a_352_406# VPB phighvt w=1e+06u l=250000u
+  ad=2.4e+11p pd=2.48e+06u as=5.55e+11p ps=5.11e+06u
M1002 VPWR CLK a_750_108# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=2.85e+11p ps=2.57e+06u
M1003 VPWR a_2006_125# a_2767_57# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=2.85e+11p ps=2.57e+06u
M1004 VGND SCE a_144_47# VNB nshort w=420000u l=150000u
+  ad=1.24265e+12p pd=1.281e+07u as=8.82e+10p ps=1.26e+06u
M1005 a_2584_57# a_2006_125# a_2172_40# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=1.197e+11p ps=1.41e+06u
M1006 VPWR SCE a_27_409# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=2.85e+11p ps=2.57e+06u
M1007 VGND a_2006_125# a_2584_57# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_1928_125# a_1199_419# VGND VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1009 VPWR a_1425_99# a_1371_419# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=2.8e+11p ps=2.56e+06u
M1010 VPWR SET_B a_1425_99# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=2.8e+11p ps=2.56e+06u
M1011 a_2006_125# a_750_108# a_1928_419# VPB phighvt w=1e+06u l=250000u
+  ad=9.35e+11p pd=5.87e+06u as=2.4e+11p ps=2.48e+06u
M1012 VGND a_2006_125# a_2854_57# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1013 a_2206_419# a_986_409# a_2006_125# VPB phighvt w=1e+06u l=250000u
+  ad=2.9e+11p pd=2.58e+06u as=0p ps=0u
M1014 VGND SET_B a_1736_125# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1015 VPWR a_2006_125# a_2172_40# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=2.85e+11p ps=2.57e+06u
M1016 a_352_406# a_27_409# a_245_406# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_144_47# SCE a_27_409# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1018 VPWR SCE a_458_406# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_1199_419# a_986_409# a_352_406# VPB phighvt w=1e+06u l=250000u
+  ad=6.1e+11p pd=3.22e+06u as=0p ps=0u
M1020 a_1199_419# a_750_108# a_352_406# VNB nshort w=420000u l=150000u
+  ad=1.722e+11p pd=1.66e+06u as=2.373e+11p ps=2.81e+06u
M1021 a_2006_125# SET_B VPWR VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_368_47# a_27_409# VGND VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1023 a_352_406# D a_368_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 VGND SCD a_532_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1025 a_1736_125# a_1199_419# a_1425_99# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1026 Q a_2767_57# a_3012_57# VNB nshort w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=8.82e+10p ps=1.26e+06u
M1027 a_2854_57# a_2006_125# a_2767_57# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1028 a_1371_419# a_750_108# a_1199_419# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1029 VGND CLK a_837_108# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1030 a_986_409# a_750_108# a_1001_108# VNB nshort w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=8.82e+10p ps=1.26e+06u
M1031 a_1001_108# a_750_108# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 a_3012_57# a_2767_57# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 VPWR a_2172_40# a_2206_419# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1034 VGND a_1425_99# a_1383_125# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1035 a_986_409# a_750_108# VPWR VPB phighvt w=1e+06u l=250000u
+  ad=2.7e+11p pd=2.54e+06u as=0p ps=0u
M1036 a_1425_99# a_1199_419# VPWR VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1037 Q a_2767_57# VPWR VPB phighvt w=1e+06u l=250000u
+  ad=2.85e+11p pd=2.57e+06u as=0p ps=0u
M1038 VGND SET_B a_2202_66# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1039 a_2124_66# a_750_108# a_2006_125# VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=2.7035e+11p ps=2.31e+06u
M1040 a_2202_66# a_2172_40# a_2124_66# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1041 a_837_108# CLK a_750_108# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1042 a_2006_125# a_986_409# a_1928_125# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1043 a_1928_419# a_1199_419# VPWR VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1044 a_532_47# SCE a_352_406# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1045 a_1383_125# a_986_409# a_1199_419# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

