* File: sky130_fd_sc_lp__or3_lp.pex.spice
* Created: Wed Sep  2 10:30:49 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__OR3_LP%A_108_31# 1 2 3 12 14 15 16 18 21 23 25 28 29
+ 31 32 35 37 43 47 49 50 51
r109 49 50 9.3668 $w=4.73e-07 $l=1.65e-07 $layer=LI1_cond $X=3.487 $Y=2.23
+ $X2=3.487 $Y2=2.065
r110 45 51 3.70735 $w=2.5e-07 $l=1.18427e-07 $layer=LI1_cond $X=3.64 $Y=1.035
+ $X2=3.56 $Y2=0.95
r111 45 50 67.1979 $w=1.68e-07 $l=1.03e-06 $layer=LI1_cond $X=3.64 $Y=1.035
+ $X2=3.64 $Y2=2.065
r112 41 51 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.56 $Y=0.865
+ $X2=3.56 $Y2=0.95
r113 41 43 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=3.56 $Y=0.865
+ $X2=3.56 $Y2=0.495
r114 38 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.145 $Y=0.95
+ $X2=1.98 $Y2=0.95
r115 37 51 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.395 $Y=0.95
+ $X2=3.56 $Y2=0.95
r116 37 38 81.5508 $w=1.68e-07 $l=1.25e-06 $layer=LI1_cond $X=3.395 $Y=0.95
+ $X2=2.145 $Y2=0.95
r117 33 47 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.98 $Y=0.865
+ $X2=1.98 $Y2=0.95
r118 33 35 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.98 $Y=0.865
+ $X2=1.98 $Y2=0.495
r119 31 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.815 $Y=0.95
+ $X2=1.98 $Y2=0.95
r120 31 32 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=1.815 $Y=0.95
+ $X2=1.355 $Y2=0.95
r121 28 29 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.19
+ $Y=1.335 $X2=1.19 $Y2=1.335
r122 26 32 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.19 $Y=1.035
+ $X2=1.355 $Y2=0.95
r123 26 28 10.4768 $w=3.28e-07 $l=3e-07 $layer=LI1_cond $X=1.19 $Y=1.035
+ $X2=1.19 $Y2=1.335
r124 24 29 1.83347 $w=4.55e-07 $l=1.5e-08 $layer=POLY_cond $X=1.127 $Y=1.32
+ $X2=1.127 $Y2=1.335
r125 24 25 11.0167 $w=3.02e-07 $l=7.5e-08 $layer=POLY_cond $X=1.127 $Y=1.32
+ $X2=1.127 $Y2=1.245
r126 23 29 33.9804 $w=4.55e-07 $l=2.78e-07 $layer=POLY_cond $X=1.127 $Y=1.613
+ $X2=1.127 $Y2=1.335
r127 19 25 11.0167 $w=3.02e-07 $l=1.85753e-07 $layer=POLY_cond $X=0.975 $Y=1.17
+ $X2=1.127 $Y2=1.245
r128 19 21 346.117 $w=1.5e-07 $l=6.75e-07 $layer=POLY_cond $X=0.975 $Y=1.17
+ $X2=0.975 $Y2=0.495
r129 16 23 44.4147 $w=3.82e-07 $l=4.33553e-07 $layer=POLY_cond $X=0.945 $Y=1.965
+ $X2=1.127 $Y2=1.613
r130 16 18 111.824 $w=2.5e-07 $l=5.8e-07 $layer=POLY_cond $X=0.945 $Y=1.965
+ $X2=0.945 $Y2=2.545
r131 14 25 15.6242 $w=1.5e-07 $l=2.27e-07 $layer=POLY_cond $X=0.9 $Y=1.245
+ $X2=1.127 $Y2=1.245
r132 14 15 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=0.9 $Y=1.245
+ $X2=0.69 $Y2=1.245
r133 10 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.615 $Y=1.17
+ $X2=0.69 $Y2=1.245
r134 10 12 346.117 $w=1.5e-07 $l=6.75e-07 $layer=POLY_cond $X=0.615 $Y=1.17
+ $X2=0.615 $Y2=0.495
r135 3 49 300 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_PDIFF $count=2 $X=3.275
+ $Y=2.045 $X2=3.415 $Y2=2.23
r136 2 43 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=3.42
+ $Y=0.285 $X2=3.56 $Y2=0.495
r137 1 35 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.84
+ $Y=0.285 $X2=1.98 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__OR3_LP%A 1 3 4 5 6 8 12 13 15 16 17 18 19 20 34 35
+ 36
r65 34 36 46.2775 $w=4.25e-07 $l=1.65e-07 $layer=POLY_cond $X=1.902 $Y=1.38
+ $X2=1.902 $Y2=1.215
r66 34 35 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.855
+ $Y=1.38 $X2=1.855 $Y2=1.38
r67 19 20 6.23308 $w=7.08e-07 $l=3.7e-07 $layer=LI1_cond $X=1.92 $Y=2.405
+ $X2=1.92 $Y2=2.775
r68 18 19 6.23308 $w=7.08e-07 $l=3.7e-07 $layer=LI1_cond $X=1.92 $Y=2.035
+ $X2=1.92 $Y2=2.405
r69 17 18 6.23308 $w=7.08e-07 $l=3.7e-07 $layer=LI1_cond $X=1.92 $Y=1.665
+ $X2=1.92 $Y2=2.035
r70 17 35 4.80116 $w=7.08e-07 $l=2.85e-07 $layer=LI1_cond $X=1.92 $Y=1.665
+ $X2=1.92 $Y2=1.38
r71 13 15 103.148 $w=2.5e-07 $l=5.35e-07 $layer=POLY_cond $X=2.09 $Y=2.01
+ $X2=2.09 $Y2=2.545
r72 12 13 45.1206 $w=3.6e-07 $l=4.20625e-07 $layer=POLY_cond $X=1.902 $Y=1.673
+ $X2=2.09 $Y2=2.01
r73 11 34 6.15041 $w=4.25e-07 $l=4.7e-08 $layer=POLY_cond $X=1.902 $Y=1.427
+ $X2=1.902 $Y2=1.38
r74 11 12 32.1915 $w=4.25e-07 $l=2.46e-07 $layer=POLY_cond $X=1.902 $Y=1.427
+ $X2=1.902 $Y2=1.673
r75 9 16 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.765 $Y=0.93
+ $X2=1.765 $Y2=0.855
r76 9 36 146.138 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=1.765 $Y=0.93
+ $X2=1.765 $Y2=1.215
r77 6 16 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.765 $Y=0.78
+ $X2=1.765 $Y2=0.855
r78 6 8 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=1.765 $Y=0.78 $X2=1.765
+ $Y2=0.495
r79 4 16 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.69 $Y=0.855
+ $X2=1.765 $Y2=0.855
r80 4 5 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=1.69 $Y=0.855 $X2=1.48
+ $Y2=0.855
r81 1 5 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.405 $Y=0.78
+ $X2=1.48 $Y2=0.855
r82 1 3 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=1.405 $Y=0.78 $X2=1.405
+ $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__OR3_LP%B 1 3 4 5 10 12 14 15 17 18 19 20 21 22 23 29
+ 30
r60 29 30 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.62
+ $Y=1.38 $X2=2.62 $Y2=1.38
r61 22 23 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=2.62 $Y=2.405
+ $X2=2.62 $Y2=2.775
r62 21 22 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=2.62 $Y=2.035
+ $X2=2.62 $Y2=2.405
r63 20 21 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=2.62 $Y=1.665
+ $X2=2.62 $Y2=2.035
r64 20 30 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=2.62 $Y=1.665
+ $X2=2.62 $Y2=1.38
r65 18 29 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.62 $Y=1.72
+ $X2=2.62 $Y2=1.38
r66 18 19 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.62 $Y=1.72
+ $X2=2.62 $Y2=1.885
r67 17 29 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.62 $Y=1.215
+ $X2=2.62 $Y2=1.38
r68 12 15 20.4101 $w=1.5e-07 $l=8.12404e-08 $layer=POLY_cond $X=2.555 $Y=0.78
+ $X2=2.542 $Y2=0.855
r69 12 14 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.555 $Y=0.78
+ $X2=2.555 $Y2=0.495
r70 10 19 163.979 $w=2.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.58 $Y=2.545
+ $X2=2.58 $Y2=1.885
r71 6 15 20.4101 $w=1.5e-07 $l=8.07775e-08 $layer=POLY_cond $X=2.53 $Y=0.93
+ $X2=2.542 $Y2=0.855
r72 6 17 146.138 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.53 $Y=0.93
+ $X2=2.53 $Y2=1.215
r73 4 15 5.30422 $w=1.5e-07 $l=8.7e-08 $layer=POLY_cond $X=2.455 $Y=0.855
+ $X2=2.542 $Y2=0.855
r74 4 5 94.8617 $w=1.5e-07 $l=1.85e-07 $layer=POLY_cond $X=2.455 $Y=0.855
+ $X2=2.27 $Y2=0.855
r75 1 5 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.195 $Y=0.78
+ $X2=2.27 $Y2=0.855
r76 1 3 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.195 $Y=0.78 $X2=2.195
+ $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__OR3_LP%C 1 3 8 10 12 16 19 20 21 22 25 26
r47 25 26 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.19
+ $Y=1.38 $X2=3.19 $Y2=1.38
r48 22 26 9.38418 $w=3.48e-07 $l=2.85e-07 $layer=LI1_cond $X=3.18 $Y=1.665
+ $X2=3.18 $Y2=1.38
r49 20 25 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=3.19 $Y=1.72
+ $X2=3.19 $Y2=1.38
r50 20 21 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.19 $Y=1.72
+ $X2=3.19 $Y2=1.885
r51 19 25 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.19 $Y=1.215
+ $X2=3.19 $Y2=1.38
r52 15 16 125.628 $w=1.5e-07 $l=2.45e-07 $layer=POLY_cond $X=3.1 $Y=0.855
+ $X2=3.345 $Y2=0.855
r53 13 15 58.9681 $w=1.5e-07 $l=1.15e-07 $layer=POLY_cond $X=2.985 $Y=0.855
+ $X2=3.1 $Y2=0.855
r54 10 16 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.345 $Y=0.78
+ $X2=3.345 $Y2=0.855
r55 10 12 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.345 $Y=0.78
+ $X2=3.345 $Y2=0.495
r56 8 21 163.979 $w=2.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.15 $Y=2.545
+ $X2=3.15 $Y2=1.885
r57 4 15 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.1 $Y=0.93 $X2=3.1
+ $Y2=0.855
r58 4 19 146.138 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.1 $Y=0.93 $X2=3.1
+ $Y2=1.215
r59 1 13 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.985 $Y=0.78
+ $X2=2.985 $Y2=0.855
r60 1 3 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.985 $Y=0.78 $X2=2.985
+ $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__OR3_LP%X 1 2 7 8 9 10 11 12 13 35
r21 13 57 2.07652 $w=7.18e-07 $l=1.25e-07 $layer=LI1_cond $X=0.485 $Y=2.775
+ $X2=0.485 $Y2=2.9
r22 12 13 6.14651 $w=7.18e-07 $l=3.7e-07 $layer=LI1_cond $X=0.485 $Y=2.405
+ $X2=0.485 $Y2=2.775
r23 12 49 3.57162 $w=7.18e-07 $l=2.15e-07 $layer=LI1_cond $X=0.485 $Y=2.405
+ $X2=0.485 $Y2=2.19
r24 11 49 2.57489 $w=7.18e-07 $l=1.55e-07 $layer=LI1_cond $X=0.485 $Y=2.035
+ $X2=0.485 $Y2=2.19
r25 10 11 6.14651 $w=7.18e-07 $l=3.7e-07 $layer=LI1_cond $X=0.485 $Y=1.665
+ $X2=0.485 $Y2=2.035
r26 9 10 6.14651 $w=7.18e-07 $l=3.7e-07 $layer=LI1_cond $X=0.485 $Y=1.295
+ $X2=0.485 $Y2=1.665
r27 8 9 6.14651 $w=7.18e-07 $l=3.7e-07 $layer=LI1_cond $X=0.485 $Y=0.925
+ $X2=0.485 $Y2=1.295
r28 8 35 2.07652 $w=7.18e-07 $l=1.25e-07 $layer=LI1_cond $X=0.485 $Y=0.925
+ $X2=0.485 $Y2=0.8
r29 7 35 4.3828 $w=7.2e-07 $l=2.45e-07 $layer=LI1_cond $X=0.485 $Y=0.555
+ $X2=0.485 $Y2=0.8
r30 7 60 1.16561 $w=6.28e-07 $l=6e-08 $layer=LI1_cond $X=0.485 $Y=0.555
+ $X2=0.485 $Y2=0.495
r31 2 57 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.535
+ $Y=2.045 $X2=0.68 $Y2=2.9
r32 2 49 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.535
+ $Y=2.045 $X2=0.68 $Y2=2.19
r33 1 60 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.255
+ $Y=0.285 $X2=0.4 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__OR3_LP%VPWR 1 6 10 12 22 23 26
r29 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r30 22 23 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r31 20 27 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r32 19 22 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=1.68 $Y=3.33
+ $X2=3.6 $Y2=3.33
r33 19 20 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r34 17 26 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.375 $Y=3.33
+ $X2=1.21 $Y2=3.33
r35 17 19 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.375 $Y=3.33
+ $X2=1.68 $Y2=3.33
r36 15 27 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r37 14 15 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r38 12 26 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.045 $Y=3.33
+ $X2=1.21 $Y2=3.33
r39 12 14 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=1.045 $Y=3.33
+ $X2=0.72 $Y2=3.33
r40 10 23 0.468274 $w=4.9e-07 $l=1.68e-06 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=3.6 $Y2=3.33
r41 10 20 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=1.68 $Y2=3.33
r42 6 9 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=1.21 $Y=2.19 $X2=1.21
+ $Y2=2.9
r43 4 26 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.21 $Y=3.245 $X2=1.21
+ $Y2=3.33
r44 4 9 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=1.21 $Y=3.245
+ $X2=1.21 $Y2=2.9
r45 1 9 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=1.07
+ $Y=2.045 $X2=1.21 $Y2=2.9
r46 1 6 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.07
+ $Y=2.045 $X2=1.21 $Y2=2.19
.ends

.subckt PM_SKY130_FD_SC_LP__OR3_LP%VGND 1 2 9 13 15 17 22 29 30 33 36
r52 36 37 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r53 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r54 30 37 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=2.64
+ $Y2=0
r55 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r56 27 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.935 $Y=0 $X2=2.77
+ $Y2=0
r57 27 29 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=2.935 $Y=0 $X2=3.6
+ $Y2=0
r58 26 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r59 25 26 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r60 23 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.355 $Y=0 $X2=1.19
+ $Y2=0
r61 23 25 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=1.355 $Y=0 $X2=1.68
+ $Y2=0
r62 22 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.605 $Y=0 $X2=2.77
+ $Y2=0
r63 22 25 60.3476 $w=1.68e-07 $l=9.25e-07 $layer=LI1_cond $X=2.605 $Y=0 $X2=1.68
+ $Y2=0
r64 20 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r65 19 20 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r66 17 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.025 $Y=0 $X2=1.19
+ $Y2=0
r67 17 19 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.025 $Y=0 $X2=0.72
+ $Y2=0
r68 15 37 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=2.64
+ $Y2=0
r69 15 26 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=1.68
+ $Y2=0
r70 11 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.77 $Y=0.085
+ $X2=2.77 $Y2=0
r71 11 13 13.6198 $w=3.28e-07 $l=3.9e-07 $layer=LI1_cond $X=2.77 $Y=0.085
+ $X2=2.77 $Y2=0.475
r72 7 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.19 $Y=0.085 $X2=1.19
+ $Y2=0
r73 7 9 13.6198 $w=3.28e-07 $l=3.9e-07 $layer=LI1_cond $X=1.19 $Y=0.085 $X2=1.19
+ $Y2=0.475
r74 2 13 182 $w=1.7e-07 $l=2.504e-07 $layer=licon1_NDIFF $count=1 $X=2.63
+ $Y=0.285 $X2=2.77 $Y2=0.475
r75 1 9 182 $w=1.7e-07 $l=2.504e-07 $layer=licon1_NDIFF $count=1 $X=1.05
+ $Y=0.285 $X2=1.19 $Y2=0.475
.ends

