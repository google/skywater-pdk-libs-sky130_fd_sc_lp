* File: sky130_fd_sc_lp__nor2_2.spice
* Created: Wed Sep  2 10:07:30 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__nor2_2.pex.spice"
.subckt sky130_fd_sc_lp__nor2_2  VNB VPB A B VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1000 N_Y_M1000_d N_A_M1000_g N_VGND_M1000_s VNB NSHORT L=0.15 W=0.84 AD=0.1176
+ AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2 SB=75001.5 A=0.126
+ P=1.98 MULT=1
MM1002 N_Y_M1000_d N_A_M1002_g N_VGND_M1002_s VNB NSHORT L=0.15 W=0.84 AD=0.1176
+ AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6 SB=75001.1 A=0.126
+ P=1.98 MULT=1
MM1001 N_VGND_M1002_s N_B_M1001_g N_Y_M1001_s VNB NSHORT L=0.15 W=0.84 AD=0.1176
+ AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.1 SB=75000.7 A=0.126
+ P=1.98 MULT=1
MM1004 N_VGND_M1004_d N_B_M1004_g N_Y_M1001_s VNB NSHORT L=0.15 W=0.84 AD=0.252
+ AS=0.1176 PD=2.28 PS=1.12 NRD=4.992 NRS=0 M=1 R=5.6 SA=75001.5 SB=75000.2
+ A=0.126 P=1.98 MULT=1
MM1003 N_A_28_367#_M1003_d N_A_M1003_g N_VPWR_M1003_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75001.6 A=0.189 P=2.82 MULT=1
MM1006 N_A_28_367#_M1006_d N_A_M1006_g N_VPWR_M1003_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75001.2 A=0.189 P=2.82 MULT=1
MM1005 N_A_28_367#_M1006_d N_B_M1005_g N_Y_M1005_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75000.8 A=0.189 P=2.82 MULT=1
MM1007 N_A_28_367#_M1007_d N_B_M1007_g N_Y_M1005_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.5166 AS=0.1764 PD=3.34 PS=1.54 NRD=22.655 NRS=0 M=1 R=8.4 SA=75001.5
+ SB=75000.3 A=0.189 P=2.82 MULT=1
DX8_noxref VNB VPB NWDIODE A=5.1847 P=9.29
*
.include "sky130_fd_sc_lp__nor2_2.pxi.spice"
*
.ends
*
*
