* File: sky130_fd_sc_lp__a311o_2.pex.spice
* Created: Fri Aug 28 09:57:38 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A311O_2%A_85_21# 1 2 3 10 12 15 17 19 21 22 24 26 30
+ 33 34 35 36 37 40 42 46 52 54 56
c128 24 0 2.55214e-20 $X=1.005 $Y=2.465
r129 50 52 15.7996 $w=3.08e-07 $l=4.25e-07 $layer=LI1_cond $X=3.905 $Y=0.845
+ $X2=3.905 $Y2=0.42
r130 46 48 33.8748 $w=3.28e-07 $l=9.7e-07 $layer=LI1_cond $X=3.895 $Y=1.98
+ $X2=3.895 $Y2=2.95
r131 44 46 3.66686 $w=3.28e-07 $l=1.05e-07 $layer=LI1_cond $X=3.895 $Y=1.875
+ $X2=3.895 $Y2=1.98
r132 43 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.035 $Y=0.93
+ $X2=2.87 $Y2=0.93
r133 42 50 7.59919 $w=1.7e-07 $l=1.92873e-07 $layer=LI1_cond $X=3.75 $Y=0.93
+ $X2=3.905 $Y2=0.845
r134 42 43 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=3.75 $Y=0.93
+ $X2=3.035 $Y2=0.93
r135 38 56 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.87 $Y=0.845
+ $X2=2.87 $Y2=0.93
r136 38 40 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=2.87 $Y=0.845
+ $X2=2.87 $Y2=0.38
r137 36 44 7.61292 $w=1.8e-07 $l=2.05122e-07 $layer=LI1_cond $X=3.73 $Y=1.785
+ $X2=3.895 $Y2=1.875
r138 36 37 153.116 $w=1.78e-07 $l=2.485e-06 $layer=LI1_cond $X=3.73 $Y=1.785
+ $X2=1.245 $Y2=1.785
r139 34 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.705 $Y=0.93
+ $X2=2.87 $Y2=0.93
r140 34 35 95.2513 $w=1.68e-07 $l=1.46e-06 $layer=LI1_cond $X=2.705 $Y=0.93
+ $X2=1.245 $Y2=0.93
r141 33 37 6.82373 $w=1.8e-07 $l=1.25499e-07 $layer=LI1_cond $X=1.16 $Y=1.695
+ $X2=1.245 $Y2=1.785
r142 33 54 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=1.16 $Y=1.695
+ $X2=1.16 $Y2=1.515
r143 31 57 11.5066 $w=3.77e-07 $l=9e-08 $layer=POLY_cond $X=1.045 $Y=1.35
+ $X2=1.045 $Y2=1.26
r144 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.07
+ $Y=1.35 $X2=1.07 $Y2=1.35
r145 28 54 7.14225 $w=2.58e-07 $l=1.3e-07 $layer=LI1_cond $X=1.115 $Y=1.385
+ $X2=1.115 $Y2=1.515
r146 28 30 1.55137 $w=2.58e-07 $l=3.5e-08 $layer=LI1_cond $X=1.115 $Y=1.385
+ $X2=1.115 $Y2=1.35
r147 27 35 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=1.115 $Y=1.015
+ $X2=1.245 $Y2=0.93
r148 27 30 14.8488 $w=2.58e-07 $l=3.35e-07 $layer=LI1_cond $X=1.115 $Y=1.015
+ $X2=1.115 $Y2=1.35
r149 22 31 39.1678 $w=3.77e-07 $l=1.83916e-07 $layer=POLY_cond $X=1.005 $Y=1.515
+ $X2=1.045 $Y2=1.35
r150 22 24 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=1.005 $Y=1.515
+ $X2=1.005 $Y2=2.465
r151 19 57 27.6612 $w=3.77e-07 $l=1.47817e-07 $layer=POLY_cond $X=0.93 $Y=1.185
+ $X2=1.045 $Y2=1.26
r152 19 21 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.93 $Y=1.185
+ $X2=0.93 $Y2=0.655
r153 18 26 5.30422 $w=1.5e-07 $l=1.13e-07 $layer=POLY_cond $X=0.65 $Y=1.26
+ $X2=0.537 $Y2=1.26
r154 17 57 24.4204 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=0.855 $Y=1.26
+ $X2=1.045 $Y2=1.26
r155 17 18 105.117 $w=1.5e-07 $l=2.05e-07 $layer=POLY_cond $X=0.855 $Y=1.26
+ $X2=0.65 $Y2=1.26
r156 13 26 20.4101 $w=1.5e-07 $l=9.20598e-08 $layer=POLY_cond $X=0.575 $Y=1.335
+ $X2=0.537 $Y2=1.26
r157 13 15 579.426 $w=1.5e-07 $l=1.13e-06 $layer=POLY_cond $X=0.575 $Y=1.335
+ $X2=0.575 $Y2=2.465
r158 10 26 20.4101 $w=1.5e-07 $l=9.16515e-08 $layer=POLY_cond $X=0.5 $Y=1.185
+ $X2=0.537 $Y2=1.26
r159 10 12 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.5 $Y=1.185
+ $X2=0.5 $Y2=0.655
r160 3 48 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=3.755
+ $Y=1.835 $X2=3.895 $Y2=2.95
r161 3 46 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=3.755
+ $Y=1.835 $X2=3.895 $Y2=1.98
r162 2 52 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=3.755
+ $Y=0.235 $X2=3.895 $Y2=0.42
r163 1 56 182 $w=1.7e-07 $l=7.86479e-07 $layer=licon1_NDIFF $count=1 $X=2.675
+ $Y=0.235 $X2=2.87 $Y2=0.93
r164 1 40 182 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_NDIFF $count=1 $X=2.675
+ $Y=0.235 $X2=2.87 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_LP__A311O_2%A3 3 7 8 11 13
c33 8 0 2.55214e-20 $X=1.68 $Y=1.295
c34 3 0 8.61388e-21 $X=1.63 $Y=2.465
r35 11 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.61 $Y=1.35
+ $X2=1.61 $Y2=1.515
r36 11 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.61 $Y=1.35
+ $X2=1.61 $Y2=1.185
r37 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.61
+ $Y=1.35 $X2=1.61 $Y2=1.35
r38 7 13 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.7 $Y=0.655 $X2=1.7
+ $Y2=1.185
r39 3 14 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=1.63 $Y=2.465
+ $X2=1.63 $Y2=1.515
.ends

.subckt PM_SKY130_FD_SC_LP__A311O_2%A2 3 6 8 11 13
c33 13 0 2.35266e-20 $X=2.15 $Y=1.195
c34 8 0 8.61388e-21 $X=2.16 $Y=1.295
r35 11 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.15 $Y=1.36
+ $X2=2.15 $Y2=1.525
r36 11 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.15 $Y=1.36
+ $X2=2.15 $Y2=1.195
r37 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.15
+ $Y=1.36 $X2=2.15 $Y2=1.36
r38 6 14 482 $w=1.5e-07 $l=9.4e-07 $layer=POLY_cond $X=2.06 $Y=2.465 $X2=2.06
+ $Y2=1.525
r39 3 13 173.52 $w=1.5e-07 $l=5.4e-07 $layer=POLY_cond $X=2.06 $Y=0.655 $X2=2.06
+ $Y2=1.195
.ends

.subckt PM_SKY130_FD_SC_LP__A311O_2%A1 3 6 8 11 13
c33 13 0 2.60245e-20 $X=2.69 $Y=1.195
c34 8 0 3.18756e-20 $X=2.64 $Y=1.295
r35 11 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.69 $Y=1.36
+ $X2=2.69 $Y2=1.525
r36 11 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.69 $Y=1.36
+ $X2=2.69 $Y2=1.195
r37 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.69
+ $Y=1.36 $X2=2.69 $Y2=1.36
r38 6 14 482 $w=1.5e-07 $l=9.4e-07 $layer=POLY_cond $X=2.78 $Y=2.465 $X2=2.78
+ $Y2=1.525
r39 3 13 173.52 $w=1.5e-07 $l=5.4e-07 $layer=POLY_cond $X=2.6 $Y=0.655 $X2=2.6
+ $Y2=1.195
.ends

.subckt PM_SKY130_FD_SC_LP__A311O_2%B1 3 6 8 9 13 15
c33 13 0 1.6798e-19 $X=3.23 $Y=1.35
c34 9 0 2.60245e-20 $X=3.6 $Y=1.295
c35 6 0 1.26579e-20 $X=3.21 $Y=2.465
r36 13 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.23 $Y=1.35
+ $X2=3.23 $Y2=1.515
r37 13 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.23 $Y=1.35
+ $X2=3.23 $Y2=1.185
r38 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.23
+ $Y=1.35 $X2=3.23 $Y2=1.35
r39 9 14 12.5413 $w=3.38e-07 $l=3.7e-07 $layer=LI1_cond $X=3.6 $Y=1.355 $X2=3.23
+ $Y2=1.355
r40 8 14 3.72849 $w=3.38e-07 $l=1.1e-07 $layer=LI1_cond $X=3.12 $Y=1.355
+ $X2=3.23 $Y2=1.355
r41 6 16 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=3.21 $Y=2.465
+ $X2=3.21 $Y2=1.515
r42 3 15 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=3.14 $Y=0.655
+ $X2=3.14 $Y2=1.185
.ends

.subckt PM_SKY130_FD_SC_LP__A311O_2%C1 1 3 6 8 13
c26 8 0 1.72289e-19 $X=4.08 $Y=1.295
r27 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.95
+ $Y=1.36 $X2=3.95 $Y2=1.36
r28 10 13 47.2125 $w=3.3e-07 $l=2.7e-07 $layer=POLY_cond $X=3.68 $Y=1.36
+ $X2=3.95 $Y2=1.36
r29 8 14 4.4064 $w=3.38e-07 $l=1.3e-07 $layer=LI1_cond $X=4.08 $Y=1.355 $X2=3.95
+ $Y2=1.355
r30 4 10 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.68 $Y=1.525
+ $X2=3.68 $Y2=1.36
r31 4 6 482 $w=1.5e-07 $l=9.4e-07 $layer=POLY_cond $X=3.68 $Y=1.525 $X2=3.68
+ $Y2=2.465
r32 1 10 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.68 $Y=1.195
+ $X2=3.68 $Y2=1.36
r33 1 3 173.52 $w=1.5e-07 $l=5.4e-07 $layer=POLY_cond $X=3.68 $Y=1.195 $X2=3.68
+ $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__A311O_2%VPWR 1 2 3 10 12 16 20 26 29 30 31 41 42 48
r57 48 49 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r58 46 49 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.2 $Y2=3.33
r59 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r60 41 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r61 39 42 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=4.08 $Y2=3.33
r62 38 41 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=2.64 $Y=3.33
+ $X2=4.08 $Y2=3.33
r63 38 39 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r64 33 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.48 $Y=3.33
+ $X2=1.315 $Y2=3.33
r65 33 35 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.48 $Y=3.33
+ $X2=2.16 $Y2=3.33
r66 31 39 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r67 31 49 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.2 $Y2=3.33
r68 31 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r69 29 35 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=2.26 $Y=3.33 $X2=2.16
+ $Y2=3.33
r70 29 30 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.26 $Y=3.33
+ $X2=2.425 $Y2=3.33
r71 28 38 3.26203 $w=1.68e-07 $l=5e-08 $layer=LI1_cond $X=2.59 $Y=3.33 $X2=2.64
+ $Y2=3.33
r72 28 30 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.59 $Y=3.33
+ $X2=2.425 $Y2=3.33
r73 24 30 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.425 $Y=3.245
+ $X2=2.425 $Y2=3.33
r74 24 26 26.1919 $w=3.28e-07 $l=7.5e-07 $layer=LI1_cond $X=2.425 $Y=3.245
+ $X2=2.425 $Y2=2.495
r75 20 23 28.6365 $w=3.28e-07 $l=8.2e-07 $layer=LI1_cond $X=1.315 $Y=2.13
+ $X2=1.315 $Y2=2.95
r76 18 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.315 $Y=3.245
+ $X2=1.315 $Y2=3.33
r77 18 23 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.315 $Y=3.245
+ $X2=1.315 $Y2=2.95
r78 17 45 4.08013 $w=1.7e-07 $l=2.33e-07 $layer=LI1_cond $X=0.465 $Y=3.33
+ $X2=0.232 $Y2=3.33
r79 16 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.15 $Y=3.33
+ $X2=1.315 $Y2=3.33
r80 16 17 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=1.15 $Y=3.33
+ $X2=0.465 $Y2=3.33
r81 12 15 41.4026 $w=2.68e-07 $l=9.7e-07 $layer=LI1_cond $X=0.33 $Y=1.98
+ $X2=0.33 $Y2=2.95
r82 10 45 3.20456 $w=2.7e-07 $l=1.33918e-07 $layer=LI1_cond $X=0.33 $Y=3.245
+ $X2=0.232 $Y2=3.33
r83 10 15 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.33 $Y=3.245
+ $X2=0.33 $Y2=2.95
r84 3 26 300 $w=1.7e-07 $l=7.91833e-07 $layer=licon1_PDIFF $count=2 $X=2.135
+ $Y=1.835 $X2=2.425 $Y2=2.495
r85 2 23 400 $w=1.7e-07 $l=1.22689e-06 $layer=licon1_PDIFF $count=1 $X=1.08
+ $Y=1.835 $X2=1.315 $Y2=2.95
r86 2 20 400 $w=1.7e-07 $l=3.95411e-07 $layer=licon1_PDIFF $count=1 $X=1.08
+ $Y=1.835 $X2=1.315 $Y2=2.13
r87 1 15 400 $w=1.7e-07 $l=1.17584e-06 $layer=licon1_PDIFF $count=1 $X=0.235
+ $Y=1.835 $X2=0.36 $Y2=2.95
r88 1 12 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.235
+ $Y=1.835 $X2=0.36 $Y2=1.98
.ends

.subckt PM_SKY130_FD_SC_LP__A311O_2%X 1 2 9 10 11 12 13 14 15 16 26 40
r29 37 40 1.28049 $w=2.68e-07 $l=3e-08 $layer=LI1_cond $X=0.77 $Y=1.985 $X2=0.77
+ $Y2=2.015
r30 16 47 5.76222 $w=2.68e-07 $l=1.35e-07 $layer=LI1_cond $X=0.77 $Y=2.775
+ $X2=0.77 $Y2=2.91
r31 15 16 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.77 $Y=2.405
+ $X2=0.77 $Y2=2.775
r32 14 37 0.768295 $w=2.68e-07 $l=1.8e-08 $layer=LI1_cond $X=0.77 $Y=1.967
+ $X2=0.77 $Y2=1.985
r33 14 50 6.41812 $w=2.68e-07 $l=1.17e-07 $layer=LI1_cond $X=0.77 $Y=1.967
+ $X2=0.77 $Y2=1.85
r34 14 15 15.0671 $w=2.68e-07 $l=3.53e-07 $layer=LI1_cond $X=0.77 $Y=2.052
+ $X2=0.77 $Y2=2.405
r35 14 40 1.57927 $w=2.68e-07 $l=3.7e-08 $layer=LI1_cond $X=0.77 $Y=2.052
+ $X2=0.77 $Y2=2.015
r36 13 50 11.7247 $w=1.73e-07 $l=1.85e-07 $layer=LI1_cond $X=0.722 $Y=1.665
+ $X2=0.722 $Y2=1.85
r37 11 12 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.695 $Y=0.925
+ $X2=0.695 $Y2=1.295
r38 10 11 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.695 $Y=0.555
+ $X2=0.695 $Y2=0.925
r39 10 26 6.76434 $w=2.28e-07 $l=1.35e-07 $layer=LI1_cond $X=0.695 $Y=0.555
+ $X2=0.695 $Y2=0.42
r40 9 13 8.23896 $w=1.73e-07 $l=1.3e-07 $layer=LI1_cond $X=0.722 $Y=1.535
+ $X2=0.722 $Y2=1.665
r41 7 12 6.26328 $w=2.28e-07 $l=1.25e-07 $layer=LI1_cond $X=0.695 $Y=1.42
+ $X2=0.695 $Y2=1.295
r42 7 9 6.44922 $w=2.28e-07 $l=1.15e-07 $layer=LI1_cond $X=0.695 $Y=1.42
+ $X2=0.695 $Y2=1.535
r43 2 47 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=0.65
+ $Y=1.835 $X2=0.79 $Y2=2.91
r44 2 40 400 $w=1.7e-07 $l=2.4e-07 $layer=licon1_PDIFF $count=1 $X=0.65 $Y=1.835
+ $X2=0.79 $Y2=2.015
r45 1 26 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=0.575
+ $Y=0.235 $X2=0.715 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__A311O_2%A_341_367# 1 2 7 9 11 13 15
r33 13 20 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.995 $Y=2.215
+ $X2=2.995 $Y2=2.13
r34 13 15 25.668 $w=3.28e-07 $l=7.35e-07 $layer=LI1_cond $X=2.995 $Y=2.215
+ $X2=2.995 $Y2=2.95
r35 12 18 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.01 $Y=2.13
+ $X2=1.845 $Y2=2.13
r36 11 20 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.83 $Y=2.13
+ $X2=2.995 $Y2=2.13
r37 11 12 53.4973 $w=1.68e-07 $l=8.2e-07 $layer=LI1_cond $X=2.83 $Y=2.13
+ $X2=2.01 $Y2=2.13
r38 7 18 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.845 $Y=2.215
+ $X2=1.845 $Y2=2.13
r39 7 9 25.668 $w=3.28e-07 $l=7.35e-07 $layer=LI1_cond $X=1.845 $Y=2.215
+ $X2=1.845 $Y2=2.95
r40 2 20 400 $w=1.7e-07 $l=3.58225e-07 $layer=licon1_PDIFF $count=1 $X=2.855
+ $Y=1.835 $X2=2.995 $Y2=2.13
r41 2 15 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=2.855
+ $Y=1.835 $X2=2.995 $Y2=2.95
r42 1 18 400 $w=1.7e-07 $l=3.58225e-07 $layer=licon1_PDIFF $count=1 $X=1.705
+ $Y=1.835 $X2=1.845 $Y2=2.13
r43 1 9 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=1.705
+ $Y=1.835 $X2=1.845 $Y2=2.95
.ends

.subckt PM_SKY130_FD_SC_LP__A311O_2%VGND 1 2 3 10 12 16 19 20 21 23 36 37 44
r53 44 47 9.81855 $w=6.68e-07 $l=5.5e-07 $layer=LI1_cond $X=1.315 $Y=0 $X2=1.315
+ $Y2=0.55
r54 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r55 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r56 36 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r57 34 37 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=4.08
+ $Y2=0
r58 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r59 31 45 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r60 30 33 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.68 $Y=0 $X2=3.12
+ $Y2=0
r61 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r62 28 44 9.03384 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=1.65 $Y=0 $X2=1.315
+ $Y2=0
r63 28 30 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=1.65 $Y=0 $X2=1.68
+ $Y2=0
r64 27 45 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r65 27 41 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r66 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r67 24 40 4.35645 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=0.41 $Y=0 $X2=0.205
+ $Y2=0
r68 24 26 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=0.41 $Y=0 $X2=0.72
+ $Y2=0
r69 23 44 9.03384 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=0.98 $Y=0 $X2=1.315
+ $Y2=0
r70 23 26 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=0.98 $Y=0 $X2=0.72
+ $Y2=0
r71 21 34 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r72 21 31 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.68
+ $Y2=0
r73 19 33 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=3.25 $Y=0 $X2=3.12
+ $Y2=0
r74 19 20 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.25 $Y=0 $X2=3.415
+ $Y2=0
r75 18 36 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=3.58 $Y=0 $X2=4.08
+ $Y2=0
r76 18 20 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.58 $Y=0 $X2=3.415
+ $Y2=0
r77 14 20 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.415 $Y=0.085
+ $X2=3.415 $Y2=0
r78 14 16 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=3.415 $Y=0.085
+ $X2=3.415 $Y2=0.55
r79 10 40 3.08139 $w=2.9e-07 $l=1.11018e-07 $layer=LI1_cond $X=0.265 $Y=0.085
+ $X2=0.205 $Y2=0
r80 10 12 11.7231 $w=2.88e-07 $l=2.95e-07 $layer=LI1_cond $X=0.265 $Y=0.085
+ $X2=0.265 $Y2=0.38
r81 3 16 182 $w=1.7e-07 $l=4.02772e-07 $layer=licon1_NDIFF $count=1 $X=3.215
+ $Y=0.235 $X2=3.415 $Y2=0.55
r82 2 47 91 $w=1.7e-07 $l=6.17738e-07 $layer=licon1_NDIFF $count=2 $X=1.005
+ $Y=0.235 $X2=1.485 $Y2=0.55
r83 1 12 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.14
+ $Y=0.235 $X2=0.285 $Y2=0.38
.ends

