# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__sdfbbp_1
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__sdfbbp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  15.84000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.465000 1.525000 1.795000 1.855000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.598500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 15.380000 0.265000 15.750000 1.125000 ;
        RECT 15.380000 1.815000 15.750000 3.065000 ;
        RECT 15.580000 1.125000 15.750000 1.815000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.598500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 13.880000 0.265000 14.315000 1.075000 ;
        RECT 13.960000 1.765000 14.315000 3.065000 ;
        RECT 14.145000 1.075000 14.315000 1.765000 ;
    END
  END Q_N
  PIN RESET_B
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 13.065000 1.180000 13.395000 1.515000 ;
    END
  END RESET_B
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.215000 0.550000 1.885000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.760000 1.550000 1.285000 1.880000 ;
    END
  END SCE
  PIN SET_B
    ANTENNAGATEAREA  0.444000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT  6.815000 1.920000  7.105000 1.965000 ;
        RECT  6.815000 1.965000 11.425000 2.105000 ;
        RECT  6.815000 2.105000  7.105000 2.150000 ;
        RECT 11.135000 1.920000 11.425000 1.965000 ;
        RECT 11.135000 2.105000 11.425000 2.150000 ;
    END
  END SET_B
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 3.445000 1.500000 3.775000 2.170000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT  0.000000 -0.085000 15.840000 0.085000 ;
        RECT  0.175000  0.085000  0.505000 1.035000 ;
        RECT  1.785000  0.085000  2.035000 0.995000 ;
        RECT  3.265000  0.085000  3.435000 0.970000 ;
        RECT  5.225000  0.085000  5.475000 0.650000 ;
        RECT  7.005000  0.085000  7.255000 0.845000 ;
        RECT  8.935000  0.085000  9.265000 0.595000 ;
        RECT 10.860000  0.085000 11.190000 0.820000 ;
        RECT 13.450000  0.085000 13.700000 1.000000 ;
        RECT 14.950000  0.085000 15.200000 1.125000 ;
      LAYER mcon ;
        RECT  0.155000 -0.085000  0.325000 0.085000 ;
        RECT  0.635000 -0.085000  0.805000 0.085000 ;
        RECT  1.115000 -0.085000  1.285000 0.085000 ;
        RECT  1.595000 -0.085000  1.765000 0.085000 ;
        RECT  2.075000 -0.085000  2.245000 0.085000 ;
        RECT  2.555000 -0.085000  2.725000 0.085000 ;
        RECT  3.035000 -0.085000  3.205000 0.085000 ;
        RECT  3.515000 -0.085000  3.685000 0.085000 ;
        RECT  3.995000 -0.085000  4.165000 0.085000 ;
        RECT  4.475000 -0.085000  4.645000 0.085000 ;
        RECT  4.955000 -0.085000  5.125000 0.085000 ;
        RECT  5.435000 -0.085000  5.605000 0.085000 ;
        RECT  5.915000 -0.085000  6.085000 0.085000 ;
        RECT  6.395000 -0.085000  6.565000 0.085000 ;
        RECT  6.875000 -0.085000  7.045000 0.085000 ;
        RECT  7.355000 -0.085000  7.525000 0.085000 ;
        RECT  7.835000 -0.085000  8.005000 0.085000 ;
        RECT  8.315000 -0.085000  8.485000 0.085000 ;
        RECT  8.795000 -0.085000  8.965000 0.085000 ;
        RECT  9.275000 -0.085000  9.445000 0.085000 ;
        RECT  9.755000 -0.085000  9.925000 0.085000 ;
        RECT 10.235000 -0.085000 10.405000 0.085000 ;
        RECT 10.715000 -0.085000 10.885000 0.085000 ;
        RECT 11.195000 -0.085000 11.365000 0.085000 ;
        RECT 11.675000 -0.085000 11.845000 0.085000 ;
        RECT 12.155000 -0.085000 12.325000 0.085000 ;
        RECT 12.635000 -0.085000 12.805000 0.085000 ;
        RECT 13.115000 -0.085000 13.285000 0.085000 ;
        RECT 13.595000 -0.085000 13.765000 0.085000 ;
        RECT 14.075000 -0.085000 14.245000 0.085000 ;
        RECT 14.555000 -0.085000 14.725000 0.085000 ;
        RECT 15.035000 -0.085000 15.205000 0.085000 ;
        RECT 15.515000 -0.085000 15.685000 0.085000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 15.840000 0.245000 ;
        RECT 0.000000  0.245000  0.500000 0.500000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.800000  0.500000 3.085000 ;
        RECT 0.000000 3.085000 15.840000 3.575000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT  0.000000 3.245000 15.840000 3.415000 ;
        RECT  0.625000 2.415000  0.955000 3.245000 ;
        RECT  2.555000 2.385000  2.805000 3.245000 ;
        RECT  3.545000 2.350000  3.875000 3.245000 ;
        RECT  5.045000 2.265000  5.375000 3.245000 ;
        RECT  6.955000 2.680000  7.285000 3.245000 ;
        RECT  8.375000 2.310000  8.705000 3.245000 ;
        RECT 11.010000 2.680000 11.340000 3.245000 ;
        RECT 12.370000 2.680000 12.700000 3.245000 ;
        RECT 13.450000 2.680000 13.780000 3.245000 ;
        RECT 14.950000 1.815000 15.200000 3.245000 ;
      LAYER mcon ;
        RECT  0.155000 3.245000  0.325000 3.415000 ;
        RECT  0.635000 3.245000  0.805000 3.415000 ;
        RECT  1.115000 3.245000  1.285000 3.415000 ;
        RECT  1.595000 3.245000  1.765000 3.415000 ;
        RECT  2.075000 3.245000  2.245000 3.415000 ;
        RECT  2.555000 3.245000  2.725000 3.415000 ;
        RECT  3.035000 3.245000  3.205000 3.415000 ;
        RECT  3.515000 3.245000  3.685000 3.415000 ;
        RECT  3.995000 3.245000  4.165000 3.415000 ;
        RECT  4.475000 3.245000  4.645000 3.415000 ;
        RECT  4.955000 3.245000  5.125000 3.415000 ;
        RECT  5.435000 3.245000  5.605000 3.415000 ;
        RECT  5.915000 3.245000  6.085000 3.415000 ;
        RECT  6.395000 3.245000  6.565000 3.415000 ;
        RECT  6.875000 3.245000  7.045000 3.415000 ;
        RECT  7.355000 3.245000  7.525000 3.415000 ;
        RECT  7.835000 3.245000  8.005000 3.415000 ;
        RECT  8.315000 3.245000  8.485000 3.415000 ;
        RECT  8.795000 3.245000  8.965000 3.415000 ;
        RECT  9.275000 3.245000  9.445000 3.415000 ;
        RECT  9.755000 3.245000  9.925000 3.415000 ;
        RECT 10.235000 3.245000 10.405000 3.415000 ;
        RECT 10.715000 3.245000 10.885000 3.415000 ;
        RECT 11.195000 3.245000 11.365000 3.415000 ;
        RECT 11.675000 3.245000 11.845000 3.415000 ;
        RECT 12.155000 3.245000 12.325000 3.415000 ;
        RECT 12.635000 3.245000 12.805000 3.415000 ;
        RECT 13.115000 3.245000 13.285000 3.415000 ;
        RECT 13.595000 3.245000 13.765000 3.415000 ;
        RECT 14.075000 3.245000 14.245000 3.415000 ;
        RECT 14.555000 3.245000 14.725000 3.415000 ;
        RECT 15.035000 3.245000 15.205000 3.415000 ;
        RECT 15.515000 3.245000 15.685000 3.415000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.115000 2.065000  1.305000 2.235000 ;
      RECT  0.115000 2.235000  0.445000 3.065000 ;
      RECT  0.995000 0.575000  1.325000 1.175000 ;
      RECT  0.995000 1.175000  2.385000 1.345000 ;
      RECT  1.135000 2.235000  1.305000 2.895000 ;
      RECT  1.135000 2.895000  2.325000 3.065000 ;
      RECT  1.485000 2.035000  2.145000 2.205000 ;
      RECT  1.485000 2.205000  1.815000 2.715000 ;
      RECT  1.975000 1.345000  2.145000 2.035000 ;
      RECT  1.995000 2.385000  2.325000 2.895000 ;
      RECT  2.215000 0.265000  3.085000 0.435000 ;
      RECT  2.215000 0.435000  2.385000 1.175000 ;
      RECT  2.325000 1.525000  2.735000 1.685000 ;
      RECT  2.325000 1.685000  3.155000 1.855000 ;
      RECT  2.565000 0.615000  2.735000 1.525000 ;
      RECT  2.915000 0.435000  3.085000 1.150000 ;
      RECT  2.915000 1.150000  3.785000 1.320000 ;
      RECT  2.985000 1.855000  3.155000 2.385000 ;
      RECT  2.985000 2.385000  3.315000 3.065000 ;
      RECT  3.615000 0.265000  5.045000 0.435000 ;
      RECT  3.615000 0.435000  3.785000 1.150000 ;
      RECT  3.965000 0.615000  4.345000 1.730000 ;
      RECT  4.055000 1.730000  4.345000 3.030000 ;
      RECT  4.525000 0.615000  4.695000 1.915000 ;
      RECT  4.525000 1.915000  5.560000 2.085000 ;
      RECT  4.525000 2.085000  4.865000 2.945000 ;
      RECT  4.875000 0.435000  5.045000 0.830000 ;
      RECT  4.875000 0.830000  5.955000 1.000000 ;
      RECT  4.925000 1.180000  5.215000 1.410000 ;
      RECT  5.045000 1.410000  5.215000 1.415000 ;
      RECT  5.045000 1.415000  5.560000 1.915000 ;
      RECT  5.625000 2.265000  5.955000 2.725000 ;
      RECT  5.705000 0.265000  5.955000 0.830000 ;
      RECT  5.785000 1.000000  5.955000 2.265000 ;
      RECT  6.135000 0.265000  6.465000 1.025000 ;
      RECT  6.135000 1.025000  7.995000 1.195000 ;
      RECT  6.135000 1.195000  6.305000 2.725000 ;
      RECT  6.485000 1.450000  6.815000 1.770000 ;
      RECT  6.485000 1.770000  6.655000 2.330000 ;
      RECT  6.485000 2.330000  7.795000 2.500000 ;
      RECT  6.845000 1.950000  7.165000 2.150000 ;
      RECT  6.995000 1.375000  7.525000 1.780000 ;
      RECT  6.995000 1.780000  7.165000 1.950000 ;
      RECT  7.435000 0.265000  8.705000 0.465000 ;
      RECT  7.435000 0.465000  7.765000 0.845000 ;
      RECT  7.465000 1.960000  9.360000 2.130000 ;
      RECT  7.465000 2.130000  7.795000 2.330000 ;
      RECT  7.465000 2.500000  7.795000 2.725000 ;
      RECT  7.705000 1.195000  7.995000 1.695000 ;
      RECT  7.945000 0.645000  8.345000 0.815000 ;
      RECT  8.175000 0.815000  8.345000 1.960000 ;
      RECT  8.525000 0.775000  9.615000 0.945000 ;
      RECT  8.525000 0.945000  8.820000 1.315000 ;
      RECT  9.030000 1.125000  9.360000 1.960000 ;
      RECT  9.280000 2.595000 10.395000 2.765000 ;
      RECT  9.280000 2.765000  9.610000 3.015000 ;
      RECT  9.445000 0.265000 10.655000 0.435000 ;
      RECT  9.445000 0.435000  9.615000 0.775000 ;
      RECT  9.610000 1.125000  9.955000 2.085000 ;
      RECT  9.610000 2.085000 10.045000 2.415000 ;
      RECT  9.795000 0.615000 10.305000 0.945000 ;
      RECT 10.135000 0.945000 10.305000 1.350000 ;
      RECT 10.135000 1.350000 11.760000 1.520000 ;
      RECT 10.225000 1.520000 10.395000 2.595000 ;
      RECT 10.485000 0.435000 10.655000 1.000000 ;
      RECT 10.485000 1.000000 11.760000 1.170000 ;
      RECT 10.575000 1.745000 10.870000 2.330000 ;
      RECT 10.575000 2.330000 13.780000 2.500000 ;
      RECT 11.080000 1.765000 11.410000 2.150000 ;
      RECT 11.370000 0.265000 12.650000 0.435000 ;
      RECT 11.370000 0.435000 11.700000 0.650000 ;
      RECT 11.520000 2.500000 11.850000 3.065000 ;
      RECT 11.590000 0.830000 13.270000 1.000000 ;
      RECT 11.590000 1.520000 11.760000 1.715000 ;
      RECT 11.590000 1.715000 11.970000 2.045000 ;
      RECT 11.940000 1.205000 12.320000 1.535000 ;
      RECT 12.150000 1.535000 12.320000 2.330000 ;
      RECT 12.400000 0.435000 12.650000 0.650000 ;
      RECT 12.500000 1.000000 12.800000 1.765000 ;
      RECT 12.500000 1.765000 13.270000 1.935000 ;
      RECT 12.940000 1.935000 13.270000 2.150000 ;
      RECT 13.020000 0.635000 13.270000 0.830000 ;
      RECT 13.610000 1.255000 13.965000 1.585000 ;
      RECT 13.610000 1.585000 13.780000 2.330000 ;
      RECT 14.520000 0.665000 14.770000 1.305000 ;
      RECT 14.520000 1.305000 15.400000 1.635000 ;
      RECT 14.520000 1.635000 14.770000 2.495000 ;
    LAYER mcon ;
      RECT  4.955000 1.210000  5.125000 1.380000 ;
      RECT  6.875000 1.950000  7.045000 2.120000 ;
      RECT  9.755000 1.210000  9.925000 1.380000 ;
      RECT 11.195000 1.950000 11.365000 2.120000 ;
    LAYER met1 ;
      RECT 4.895000 1.180000 5.185000 1.225000 ;
      RECT 4.895000 1.225000 9.985000 1.365000 ;
      RECT 4.895000 1.365000 5.185000 1.410000 ;
      RECT 9.695000 1.180000 9.985000 1.225000 ;
      RECT 9.695000 1.365000 9.985000 1.410000 ;
  END
END sky130_fd_sc_lp__sdfbbp_1
END LIBRARY
