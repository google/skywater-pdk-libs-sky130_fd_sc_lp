* File: sky130_fd_sc_lp__and3_2.pxi.spice
* Created: Wed Sep  2 09:31:40 2020
* 
x_PM_SKY130_FD_SC_LP__AND3_2%A N_A_c_66_n N_A_M1000_g N_A_c_61_n N_A_M1008_g
+ N_A_c_62_n N_A_c_63_n A N_A_c_64_n N_A_c_65_n PM_SKY130_FD_SC_LP__AND3_2%A
x_PM_SKY130_FD_SC_LP__AND3_2%B N_B_M1004_g N_B_M1003_g B N_B_c_98_n N_B_c_99_n
+ PM_SKY130_FD_SC_LP__AND3_2%B
x_PM_SKY130_FD_SC_LP__AND3_2%C N_C_M1005_g N_C_M1006_g C N_C_c_132_n N_C_c_133_n
+ PM_SKY130_FD_SC_LP__AND3_2%C
x_PM_SKY130_FD_SC_LP__AND3_2%A_27_385# N_A_27_385#_M1008_s N_A_27_385#_M1000_s
+ N_A_27_385#_M1003_d N_A_27_385#_M1002_g N_A_27_385#_M1001_g
+ N_A_27_385#_c_171_n N_A_27_385#_M1009_g N_A_27_385#_M1007_g
+ N_A_27_385#_c_174_n N_A_27_385#_c_183_n N_A_27_385#_c_175_n
+ N_A_27_385#_c_184_n N_A_27_385#_c_185_n N_A_27_385#_c_176_n
+ N_A_27_385#_c_177_n N_A_27_385#_c_186_n N_A_27_385#_c_187_n
+ N_A_27_385#_c_178_n N_A_27_385#_c_188_n N_A_27_385#_c_179_n
+ N_A_27_385#_c_180_n PM_SKY130_FD_SC_LP__AND3_2%A_27_385#
x_PM_SKY130_FD_SC_LP__AND3_2%VPWR N_VPWR_M1000_d N_VPWR_M1006_d N_VPWR_M1007_s
+ N_VPWR_c_279_n N_VPWR_c_280_n N_VPWR_c_281_n N_VPWR_c_282_n VPWR
+ N_VPWR_c_283_n N_VPWR_c_284_n N_VPWR_c_285_n N_VPWR_c_286_n N_VPWR_c_287_n
+ N_VPWR_c_278_n PM_SKY130_FD_SC_LP__AND3_2%VPWR
x_PM_SKY130_FD_SC_LP__AND3_2%X N_X_M1002_d N_X_M1001_d N_X_c_316_n N_X_c_312_n X
+ X X X N_X_c_313_n PM_SKY130_FD_SC_LP__AND3_2%X
x_PM_SKY130_FD_SC_LP__AND3_2%VGND N_VGND_M1005_d N_VGND_M1009_s N_VGND_c_346_n
+ N_VGND_c_347_n N_VGND_c_348_n VGND N_VGND_c_349_n N_VGND_c_350_n
+ N_VGND_c_351_n N_VGND_c_352_n PM_SKY130_FD_SC_LP__AND3_2%VGND
cc_1 VNB N_A_c_61_n 0.0190116f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=0.765
cc_2 VNB N_A_c_62_n 0.038555f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=0.84
cc_3 VNB N_A_c_63_n 0.0244202f $X=-0.19 $Y=-0.245 $X2=0.275 $Y2=1.44
cc_4 VNB N_A_c_64_n 0.0429422f $X=-0.19 $Y=-0.245 $X2=0.275 $Y2=1.1
cc_5 VNB N_A_c_65_n 0.0231889f $X=-0.19 $Y=-0.245 $X2=0.275 $Y2=1.1
cc_6 VNB N_B_M1004_g 0.0321007f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.135
cc_7 VNB N_B_M1003_g 0.0117546f $X=-0.19 $Y=-0.245 $X2=0.275 $Y2=0.84
cc_8 VNB N_B_c_98_n 0.0296292f $X=-0.19 $Y=-0.245 $X2=0.275 $Y2=1.44
cc_9 VNB N_B_c_99_n 0.00241713f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_10 VNB N_C_M1005_g 0.0404397f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.135
cc_11 VNB N_C_M1006_g 0.00793387f $X=-0.19 $Y=-0.245 $X2=0.275 $Y2=0.84
cc_12 VNB N_C_c_132_n 0.0307224f $X=-0.19 $Y=-0.245 $X2=0.275 $Y2=1.44
cc_13 VNB N_C_c_133_n 0.00395565f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_14 VNB N_A_27_385#_M1002_g 0.0219288f $X=-0.19 $Y=-0.245 $X2=0.275 $Y2=1.44
cc_15 VNB N_A_27_385#_M1001_g 0.00244699f $X=-0.19 $Y=-0.245 $X2=0.275 $Y2=1.1
cc_16 VNB N_A_27_385#_c_171_n 0.0125902f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.27
cc_17 VNB N_A_27_385#_M1009_g 0.0282033f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_27_385#_M1007_g 0.0170691f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_27_385#_c_174_n 0.0106668f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_27_385#_c_175_n 0.0163748f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_27_385#_c_176_n 0.0206652f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_27_385#_c_177_n 0.00366547f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_27_385#_c_178_n 0.00183732f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_27_385#_c_179_n 0.00309378f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_27_385#_c_180_n 0.0272864f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_VPWR_c_278_n 0.123877f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_X_c_312_n 0.00210619f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_28 VNB N_X_c_313_n 0.00266207f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_346_n 0.00564356f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_347_n 0.0110265f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_348_n 0.0476091f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_32 VNB N_VGND_c_349_n 0.0409936f $X=-0.19 $Y=-0.245 $X2=0.275 $Y2=1.1
cc_33 VNB N_VGND_c_350_n 0.0200381f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_351_n 0.00631679f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_352_n 0.170557f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VPB N_A_c_66_n 0.0232107f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=1.815
cc_37 VPB N_A_c_63_n 0.0215533f $X=-0.19 $Y=1.655 $X2=0.275 $Y2=1.44
cc_38 VPB N_B_M1003_g 0.027154f $X=-0.19 $Y=1.655 $X2=0.275 $Y2=0.84
cc_39 VPB N_C_M1006_g 0.0274056f $X=-0.19 $Y=1.655 $X2=0.275 $Y2=0.84
cc_40 VPB N_A_27_385#_M1001_g 0.02228f $X=-0.19 $Y=1.655 $X2=0.275 $Y2=1.1
cc_41 VPB N_A_27_385#_M1007_g 0.0264958f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_42 VPB N_A_27_385#_c_183_n 0.0180391f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_43 VPB N_A_27_385#_c_184_n 0.00840357f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_44 VPB N_A_27_385#_c_185_n 0.00867164f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_45 VPB N_A_27_385#_c_186_n 8.54762e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_46 VPB N_A_27_385#_c_187_n 0.00914202f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_47 VPB N_A_27_385#_c_188_n 0.00633246f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_48 VPB N_A_27_385#_c_179_n 4.94364e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_49 VPB N_VPWR_c_279_n 0.0454521f $X=-0.19 $Y=1.655 $X2=0.275 $Y2=1.44
cc_50 VPB N_VPWR_c_280_n 0.0161432f $X=-0.19 $Y=1.655 $X2=0.275 $Y2=1.1
cc_51 VPB N_VPWR_c_281_n 0.0110006f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_52 VPB N_VPWR_c_282_n 0.0633729f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_53 VPB N_VPWR_c_283_n 0.0199636f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_54 VPB N_VPWR_c_284_n 0.0203024f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_55 VPB N_VPWR_c_285_n 0.0175247f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_56 VPB N_VPWR_c_286_n 0.00497514f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_57 VPB N_VPWR_c_287_n 0.00757184f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_58 VPB N_VPWR_c_278_n 0.0808088f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_59 VPB X 0.00167405f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_60 VPB N_X_c_313_n 0.00111866f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_61 N_A_c_61_n N_B_M1004_g 0.0521271f $X=0.545 $Y=0.765 $X2=0 $Y2=0
cc_62 N_A_c_64_n N_B_M1004_g 0.00696816f $X=0.275 $Y=1.1 $X2=0 $Y2=0
cc_63 N_A_c_65_n N_B_M1004_g 6.28508e-19 $X=0.275 $Y=1.1 $X2=0 $Y2=0
cc_64 N_A_c_63_n N_B_M1003_g 0.0274166f $X=0.275 $Y=1.44 $X2=0 $Y2=0
cc_65 N_A_c_65_n N_B_M1003_g 2.89988e-19 $X=0.275 $Y=1.1 $X2=0 $Y2=0
cc_66 N_A_c_64_n N_B_c_98_n 0.0213895f $X=0.275 $Y=1.1 $X2=0 $Y2=0
cc_67 N_A_c_65_n N_B_c_98_n 4.00596e-19 $X=0.275 $Y=1.1 $X2=0 $Y2=0
cc_68 N_A_c_64_n N_B_c_99_n 0.00107507f $X=0.275 $Y=1.1 $X2=0 $Y2=0
cc_69 N_A_c_65_n N_B_c_99_n 0.023185f $X=0.275 $Y=1.1 $X2=0 $Y2=0
cc_70 N_A_c_65_n N_C_c_133_n 0.00164786f $X=0.275 $Y=1.1 $X2=0 $Y2=0
cc_71 N_A_c_66_n N_A_27_385#_c_183_n 0.00179199f $X=0.475 $Y=1.815 $X2=0 $Y2=0
cc_72 N_A_c_61_n N_A_27_385#_c_175_n 0.00863804f $X=0.545 $Y=0.765 $X2=0 $Y2=0
cc_73 N_A_c_66_n N_A_27_385#_c_184_n 0.00903735f $X=0.475 $Y=1.815 $X2=0 $Y2=0
cc_74 N_A_c_63_n N_A_27_385#_c_184_n 0.00781205f $X=0.275 $Y=1.44 $X2=0 $Y2=0
cc_75 N_A_c_65_n N_A_27_385#_c_184_n 0.00350165f $X=0.275 $Y=1.1 $X2=0 $Y2=0
cc_76 N_A_c_63_n N_A_27_385#_c_185_n 0.0120703f $X=0.275 $Y=1.44 $X2=0 $Y2=0
cc_77 N_A_c_65_n N_A_27_385#_c_185_n 0.022615f $X=0.275 $Y=1.1 $X2=0 $Y2=0
cc_78 N_A_c_61_n N_A_27_385#_c_176_n 0.00479145f $X=0.545 $Y=0.765 $X2=0 $Y2=0
cc_79 N_A_c_62_n N_A_27_385#_c_176_n 0.00628106f $X=0.545 $Y=0.84 $X2=0 $Y2=0
cc_80 N_A_c_61_n N_A_27_385#_c_177_n 0.00200762f $X=0.545 $Y=0.765 $X2=0 $Y2=0
cc_81 N_A_c_62_n N_A_27_385#_c_177_n 0.0191487f $X=0.545 $Y=0.84 $X2=0 $Y2=0
cc_82 N_A_c_65_n N_A_27_385#_c_177_n 0.0224188f $X=0.275 $Y=1.1 $X2=0 $Y2=0
cc_83 N_A_c_66_n N_VPWR_c_279_n 0.00354012f $X=0.475 $Y=1.815 $X2=0 $Y2=0
cc_84 N_A_c_66_n N_VPWR_c_278_n 0.00380473f $X=0.475 $Y=1.815 $X2=0 $Y2=0
cc_85 N_A_c_61_n N_VGND_c_349_n 0.00420209f $X=0.545 $Y=0.765 $X2=0 $Y2=0
cc_86 N_A_c_62_n N_VGND_c_349_n 0.00175334f $X=0.545 $Y=0.84 $X2=0 $Y2=0
cc_87 N_A_c_61_n N_VGND_c_352_n 0.00675007f $X=0.545 $Y=0.765 $X2=0 $Y2=0
cc_88 N_A_c_62_n N_VGND_c_352_n 0.00148235f $X=0.545 $Y=0.84 $X2=0 $Y2=0
cc_89 N_B_M1004_g N_C_M1005_g 0.0449997f $X=0.905 $Y=0.445 $X2=0 $Y2=0
cc_90 N_B_c_99_n N_C_M1005_g 3.31196e-19 $X=0.815 $Y=1.29 $X2=0 $Y2=0
cc_91 N_B_M1003_g N_C_M1006_g 0.0194406f $X=0.905 $Y=2.135 $X2=0 $Y2=0
cc_92 N_B_c_98_n N_C_c_132_n 0.0449997f $X=0.815 $Y=1.29 $X2=0 $Y2=0
cc_93 N_B_c_99_n N_C_c_132_n 2.6023e-19 $X=0.815 $Y=1.29 $X2=0 $Y2=0
cc_94 N_B_c_98_n N_C_c_133_n 0.00248554f $X=0.815 $Y=1.29 $X2=0 $Y2=0
cc_95 N_B_c_99_n N_C_c_133_n 0.0176348f $X=0.815 $Y=1.29 $X2=0 $Y2=0
cc_96 N_B_M1004_g N_A_27_385#_c_175_n 0.00210343f $X=0.905 $Y=0.445 $X2=0 $Y2=0
cc_97 N_B_M1003_g N_A_27_385#_c_184_n 0.0177819f $X=0.905 $Y=2.135 $X2=0 $Y2=0
cc_98 N_B_c_98_n N_A_27_385#_c_184_n 0.00382224f $X=0.815 $Y=1.29 $X2=0 $Y2=0
cc_99 N_B_c_99_n N_A_27_385#_c_184_n 0.0147224f $X=0.815 $Y=1.29 $X2=0 $Y2=0
cc_100 N_B_M1004_g N_A_27_385#_c_176_n 0.0137744f $X=0.905 $Y=0.445 $X2=0 $Y2=0
cc_101 N_B_c_98_n N_A_27_385#_c_176_n 0.00373994f $X=0.815 $Y=1.29 $X2=0 $Y2=0
cc_102 N_B_c_99_n N_A_27_385#_c_176_n 0.0135177f $X=0.815 $Y=1.29 $X2=0 $Y2=0
cc_103 N_B_M1003_g N_A_27_385#_c_186_n 8.54033e-19 $X=0.905 $Y=2.135 $X2=0 $Y2=0
cc_104 N_B_M1003_g N_VPWR_c_279_n 0.0019248f $X=0.905 $Y=2.135 $X2=0 $Y2=0
cc_105 N_B_M1003_g N_VPWR_c_280_n 5.32474e-19 $X=0.905 $Y=2.135 $X2=0 $Y2=0
cc_106 N_B_M1003_g N_VPWR_c_278_n 0.00380473f $X=0.905 $Y=2.135 $X2=0 $Y2=0
cc_107 N_B_M1004_g N_VGND_c_349_n 0.00430895f $X=0.905 $Y=0.445 $X2=0 $Y2=0
cc_108 N_B_M1004_g N_VGND_c_352_n 0.00578626f $X=0.905 $Y=0.445 $X2=0 $Y2=0
cc_109 N_C_M1005_g N_A_27_385#_M1002_g 0.0205944f $X=1.265 $Y=0.445 $X2=0 $Y2=0
cc_110 N_C_c_132_n N_A_27_385#_M1002_g 0.00294109f $X=1.355 $Y=1.35 $X2=0 $Y2=0
cc_111 N_C_M1006_g N_A_27_385#_M1001_g 0.0170622f $X=1.41 $Y=2.135 $X2=0 $Y2=0
cc_112 N_C_M1005_g N_A_27_385#_c_176_n 0.0134904f $X=1.265 $Y=0.445 $X2=0 $Y2=0
cc_113 N_C_c_132_n N_A_27_385#_c_176_n 0.00497037f $X=1.355 $Y=1.35 $X2=0 $Y2=0
cc_114 N_C_c_133_n N_A_27_385#_c_176_n 0.0143092f $X=1.355 $Y=1.35 $X2=0 $Y2=0
cc_115 N_C_M1006_g N_A_27_385#_c_186_n 0.00143017f $X=1.41 $Y=2.135 $X2=0 $Y2=0
cc_116 N_C_M1006_g N_A_27_385#_c_187_n 0.0162822f $X=1.41 $Y=2.135 $X2=0 $Y2=0
cc_117 N_C_c_132_n N_A_27_385#_c_187_n 0.00245383f $X=1.355 $Y=1.35 $X2=0 $Y2=0
cc_118 N_C_c_133_n N_A_27_385#_c_187_n 0.00993486f $X=1.355 $Y=1.35 $X2=0 $Y2=0
cc_119 N_C_M1005_g N_A_27_385#_c_178_n 0.00620607f $X=1.265 $Y=0.445 $X2=0 $Y2=0
cc_120 N_C_c_132_n N_A_27_385#_c_178_n 7.15825e-19 $X=1.355 $Y=1.35 $X2=0 $Y2=0
cc_121 N_C_c_133_n N_A_27_385#_c_178_n 0.00492191f $X=1.355 $Y=1.35 $X2=0 $Y2=0
cc_122 N_C_c_132_n N_A_27_385#_c_188_n 0.0026786f $X=1.355 $Y=1.35 $X2=0 $Y2=0
cc_123 N_C_c_133_n N_A_27_385#_c_188_n 0.0137403f $X=1.355 $Y=1.35 $X2=0 $Y2=0
cc_124 N_C_M1006_g N_A_27_385#_c_179_n 0.00400022f $X=1.41 $Y=2.135 $X2=0 $Y2=0
cc_125 N_C_c_132_n N_A_27_385#_c_179_n 0.00159564f $X=1.355 $Y=1.35 $X2=0 $Y2=0
cc_126 N_C_c_133_n N_A_27_385#_c_179_n 0.0138962f $X=1.355 $Y=1.35 $X2=0 $Y2=0
cc_127 N_C_M1006_g N_A_27_385#_c_180_n 0.00437689f $X=1.41 $Y=2.135 $X2=0 $Y2=0
cc_128 N_C_c_132_n N_A_27_385#_c_180_n 0.0150508f $X=1.355 $Y=1.35 $X2=0 $Y2=0
cc_129 N_C_c_133_n N_A_27_385#_c_180_n 2.49989e-19 $X=1.355 $Y=1.35 $X2=0 $Y2=0
cc_130 N_C_M1006_g N_VPWR_c_280_n 0.0089984f $X=1.41 $Y=2.135 $X2=0 $Y2=0
cc_131 N_C_M1006_g N_VPWR_c_278_n 0.00319597f $X=1.41 $Y=2.135 $X2=0 $Y2=0
cc_132 N_C_M1005_g N_VGND_c_346_n 0.0103772f $X=1.265 $Y=0.445 $X2=0 $Y2=0
cc_133 N_C_M1005_g N_VGND_c_349_n 0.00430895f $X=1.265 $Y=0.445 $X2=0 $Y2=0
cc_134 N_C_M1005_g N_VGND_c_352_n 0.00649022f $X=1.265 $Y=0.445 $X2=0 $Y2=0
cc_135 N_A_27_385#_c_187_n N_VPWR_M1006_d 0.00108477f $X=1.695 $Y=1.79 $X2=0
+ $Y2=0
cc_136 N_A_27_385#_c_179_n N_VPWR_M1006_d 0.00119515f $X=1.895 $Y=1.44 $X2=0
+ $Y2=0
cc_137 N_A_27_385#_c_184_n N_VPWR_c_279_n 0.0172048f $X=0.99 $Y=1.79 $X2=0 $Y2=0
cc_138 N_A_27_385#_M1001_g N_VPWR_c_280_n 0.00564151f $X=1.935 $Y=2.465 $X2=0
+ $Y2=0
cc_139 N_A_27_385#_c_187_n N_VPWR_c_280_n 0.0164231f $X=1.695 $Y=1.79 $X2=0
+ $Y2=0
cc_140 N_A_27_385#_c_179_n N_VPWR_c_280_n 0.00973747f $X=1.895 $Y=1.44 $X2=0
+ $Y2=0
cc_141 N_A_27_385#_c_180_n N_VPWR_c_280_n 4.48963e-19 $X=1.895 $Y=1.35 $X2=0
+ $Y2=0
cc_142 N_A_27_385#_M1007_g N_VPWR_c_282_n 0.0111001f $X=2.365 $Y=2.465 $X2=0
+ $Y2=0
cc_143 N_A_27_385#_M1001_g N_VPWR_c_285_n 0.00585385f $X=1.935 $Y=2.465 $X2=0
+ $Y2=0
cc_144 N_A_27_385#_M1007_g N_VPWR_c_285_n 0.00526178f $X=2.365 $Y=2.465 $X2=0
+ $Y2=0
cc_145 N_A_27_385#_M1001_g N_VPWR_c_278_n 0.0118084f $X=1.935 $Y=2.465 $X2=0
+ $Y2=0
cc_146 N_A_27_385#_M1007_g N_VPWR_c_278_n 0.0102191f $X=2.365 $Y=2.465 $X2=0
+ $Y2=0
cc_147 N_A_27_385#_M1009_g N_X_c_316_n 0.00967747f $X=2.365 $Y=0.655 $X2=0 $Y2=0
cc_148 N_A_27_385#_M1002_g N_X_c_312_n 6.57003e-19 $X=1.935 $Y=0.655 $X2=0 $Y2=0
cc_149 N_A_27_385#_c_171_n N_X_c_312_n 0.00203333f $X=2.29 $Y=1.35 $X2=0 $Y2=0
cc_150 N_A_27_385#_M1009_g N_X_c_312_n 0.00203342f $X=2.365 $Y=0.655 $X2=0 $Y2=0
cc_151 N_A_27_385#_c_178_n N_X_c_312_n 0.00809133f $X=1.78 $Y=1.275 $X2=0 $Y2=0
cc_152 N_A_27_385#_M1001_g X 8.25265e-19 $X=1.935 $Y=2.465 $X2=0 $Y2=0
cc_153 N_A_27_385#_c_171_n X 0.00314165f $X=2.29 $Y=1.35 $X2=0 $Y2=0
cc_154 N_A_27_385#_M1007_g X 0.00190089f $X=2.365 $Y=2.465 $X2=0 $Y2=0
cc_155 N_A_27_385#_c_179_n X 0.00330789f $X=1.895 $Y=1.44 $X2=0 $Y2=0
cc_156 N_A_27_385#_c_180_n X 0.00111228f $X=1.895 $Y=1.35 $X2=0 $Y2=0
cc_157 N_A_27_385#_M1007_g X 0.0147653f $X=2.365 $Y=2.465 $X2=0 $Y2=0
cc_158 N_A_27_385#_M1002_g N_X_c_313_n 0.00130825f $X=1.935 $Y=0.655 $X2=0 $Y2=0
cc_159 N_A_27_385#_M1001_g N_X_c_313_n 0.00152508f $X=1.935 $Y=2.465 $X2=0 $Y2=0
cc_160 N_A_27_385#_c_171_n N_X_c_313_n 0.00853996f $X=2.29 $Y=1.35 $X2=0 $Y2=0
cc_161 N_A_27_385#_M1009_g N_X_c_313_n 0.00872021f $X=2.365 $Y=0.655 $X2=0 $Y2=0
cc_162 N_A_27_385#_M1007_g N_X_c_313_n 0.0187876f $X=2.365 $Y=2.465 $X2=0 $Y2=0
cc_163 N_A_27_385#_c_174_n N_X_c_313_n 0.00627637f $X=2.365 $Y=1.35 $X2=0 $Y2=0
cc_164 N_A_27_385#_c_178_n N_X_c_313_n 0.00875455f $X=1.78 $Y=1.275 $X2=0 $Y2=0
cc_165 N_A_27_385#_c_179_n N_X_c_313_n 0.0350302f $X=1.895 $Y=1.44 $X2=0 $Y2=0
cc_166 N_A_27_385#_c_180_n N_X_c_313_n 0.00117603f $X=1.895 $Y=1.35 $X2=0 $Y2=0
cc_167 N_A_27_385#_c_176_n N_VGND_M1005_d 0.00696743f $X=1.695 $Y=0.76 $X2=-0.19
+ $Y2=-0.245
cc_168 N_A_27_385#_c_178_n N_VGND_M1005_d 0.00309434f $X=1.78 $Y=1.275 $X2=-0.19
+ $Y2=-0.245
cc_169 N_A_27_385#_M1002_g N_VGND_c_346_n 0.00637914f $X=1.935 $Y=0.655 $X2=0
+ $Y2=0
cc_170 N_A_27_385#_c_176_n N_VGND_c_346_n 0.0260949f $X=1.695 $Y=0.76 $X2=0
+ $Y2=0
cc_171 N_A_27_385#_M1009_g N_VGND_c_348_n 0.0103479f $X=2.365 $Y=0.655 $X2=0
+ $Y2=0
cc_172 N_A_27_385#_c_175_n N_VGND_c_349_n 0.0208498f $X=0.33 $Y=0.42 $X2=0 $Y2=0
cc_173 N_A_27_385#_c_176_n N_VGND_c_349_n 0.0151309f $X=1.695 $Y=0.76 $X2=0
+ $Y2=0
cc_174 N_A_27_385#_M1002_g N_VGND_c_350_n 0.0058023f $X=1.935 $Y=0.655 $X2=0
+ $Y2=0
cc_175 N_A_27_385#_M1009_g N_VGND_c_350_n 0.00526178f $X=2.365 $Y=0.655 $X2=0
+ $Y2=0
cc_176 N_A_27_385#_c_176_n N_VGND_c_350_n 0.00107293f $X=1.695 $Y=0.76 $X2=0
+ $Y2=0
cc_177 N_A_27_385#_M1008_s N_VGND_c_352_n 0.00215158f $X=0.205 $Y=0.235 $X2=0
+ $Y2=0
cc_178 N_A_27_385#_M1002_g N_VGND_c_352_n 0.0112087f $X=1.935 $Y=0.655 $X2=0
+ $Y2=0
cc_179 N_A_27_385#_M1009_g N_VGND_c_352_n 0.0102191f $X=2.365 $Y=0.655 $X2=0
+ $Y2=0
cc_180 N_A_27_385#_c_175_n N_VGND_c_352_n 0.012522f $X=0.33 $Y=0.42 $X2=0 $Y2=0
cc_181 N_A_27_385#_c_176_n N_VGND_c_352_n 0.0283055f $X=1.695 $Y=0.76 $X2=0
+ $Y2=0
cc_182 N_VPWR_c_278_n N_X_M1001_d 0.00310528f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_183 N_VPWR_c_282_n X 0.0952263f $X=2.595 $Y=1.98 $X2=0 $Y2=0
cc_184 N_VPWR_c_285_n X 0.0174203f $X=2.5 $Y=3.33 $X2=0 $Y2=0
cc_185 N_VPWR_c_278_n X 0.0111395f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_186 N_X_c_316_n N_VGND_c_348_n 0.0622128f $X=2.15 $Y=0.42 $X2=0 $Y2=0
cc_187 N_X_c_316_n N_VGND_c_350_n 0.0163558f $X=2.15 $Y=0.42 $X2=0 $Y2=0
cc_188 N_X_M1002_d N_VGND_c_352_n 0.0041489f $X=2.01 $Y=0.235 $X2=0 $Y2=0
cc_189 N_X_c_316_n N_VGND_c_352_n 0.00996792f $X=2.15 $Y=0.42 $X2=0 $Y2=0
cc_190 A_124_47# N_VGND_c_352_n 0.00256433f $X=0.62 $Y=0.235 $X2=2.64 $Y2=0
cc_191 A_196_47# N_VGND_c_352_n 0.00256433f $X=0.98 $Y=0.235 $X2=2.64 $Y2=0
