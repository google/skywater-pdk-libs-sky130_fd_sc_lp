# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__or4b_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_lp__or4b_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.840000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.850000 1.345000 2.275000 1.835000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.445000 0.840000 2.765000 1.835000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.935000 1.125000 3.245000 1.835000 ;
    END
  END C
  PIN D_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.375000 0.480000 1.750000 ;
    END
  END D_N
  PIN X
    ANTENNADIFFAREA  0.588000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.010000 0.985000 1.330000 1.155000 ;
        RECT 1.010000 1.155000 1.180000 1.845000 ;
        RECT 1.010000 1.845000 1.320000 2.185000 ;
        RECT 1.140000 0.255000 1.330000 0.985000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.840000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.840000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.840000 0.085000 ;
      RECT 0.000000  3.245000 3.840000 3.415000 ;
      RECT 0.115000  0.700000 0.445000 0.985000 ;
      RECT 0.115000  0.985000 0.830000 1.155000 ;
      RECT 0.115000  1.920000 0.830000 2.260000 ;
      RECT 0.640000  0.085000 0.970000 0.815000 ;
      RECT 0.640000  2.695000 0.970000 3.245000 ;
      RECT 0.650000  1.155000 0.830000 1.920000 ;
      RECT 0.660000  2.260000 0.830000 2.355000 ;
      RECT 0.660000  2.355000 3.440000 2.525000 ;
      RECT 1.350000  1.335000 1.670000 1.665000 ;
      RECT 1.500000  0.085000 1.890000 0.835000 ;
      RECT 1.500000  1.005000 2.275000 1.175000 ;
      RECT 1.500000  1.175000 1.670000 1.335000 ;
      RECT 1.500000  1.665000 1.670000 2.005000 ;
      RECT 1.500000  2.005000 3.745000 2.185000 ;
      RECT 1.500000  2.695000 1.830000 3.245000 ;
      RECT 2.060000  0.280000 2.275000 1.005000 ;
      RECT 2.455000  0.085000 2.815000 0.610000 ;
      RECT 2.985000  0.255000 3.315000 0.725000 ;
      RECT 2.985000  0.725000 3.745000 0.895000 ;
      RECT 3.100000  2.525000 3.440000 3.045000 ;
      RECT 3.415000  0.895000 3.745000 2.005000 ;
      RECT 3.485000  0.085000 3.745000 0.555000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
  END
END sky130_fd_sc_lp__or4b_2
END LIBRARY
