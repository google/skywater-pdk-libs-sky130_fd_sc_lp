* File: sky130_fd_sc_lp__o41ai_lp.spice
* Created: Wed Sep  2 10:28:35 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__o41ai_lp.pex.spice"
.subckt sky130_fd_sc_lp__o41ai_lp  VNB VPB B1 A4 A3 A2 A1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A1	A1
* A2	A2
* A3	A3
* A4	A4
* B1	B1
* VPB	VPB
* VNB	VNB
MM1007 N_A_153_57#_M1007_d N_B1_M1007_g N_Y_M1007_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.1533 PD=0.7 PS=1.57 NRD=0 NRS=22.848 M=1 R=2.8 SA=75000.3
+ SB=75002.3 A=0.063 P=1.14 MULT=1
MM1003 N_VGND_M1003_d N_A4_M1003_g N_A_153_57#_M1007_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1029 AS=0.0588 PD=0.91 PS=0.7 NRD=22.848 NRS=0 M=1 R=2.8 SA=75000.7
+ SB=75001.9 A=0.063 P=1.14 MULT=1
MM1000 N_A_153_57#_M1000_d N_A3_M1000_g N_VGND_M1003_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.1029 PD=0.7 PS=0.91 NRD=0 NRS=37.14 M=1 R=2.8 SA=75001.4
+ SB=75001.2 A=0.063 P=1.14 MULT=1
MM1004 N_VGND_M1004_d N_A2_M1004_g N_A_153_57#_M1000_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0924 AS=0.0588 PD=0.86 PS=0.7 NRD=22.848 NRS=0 M=1 R=2.8 SA=75001.8
+ SB=75000.8 A=0.063 P=1.14 MULT=1
MM1005 N_A_153_57#_M1005_d N_A1_M1005_g N_VGND_M1004_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0924 PD=1.41 PS=0.86 NRD=0 NRS=22.848 M=1 R=2.8 SA=75002.4
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1002 N_Y_M1002_d N_B1_M1002_g N_VPWR_M1002_s VPB PHIGHVT L=0.25 W=1 AD=0.14
+ AS=0.285 PD=1.28 PS=2.57 NRD=0 NRS=0 M=1 R=4 SA=125000 SB=125002 A=0.25 P=2.5
+ MULT=1
MM1009 A_259_419# N_A4_M1009_g N_Y_M1002_d VPB PHIGHVT L=0.25 W=1 AD=0.125
+ AS=0.14 PD=1.25 PS=1.28 NRD=13.7703 NRS=0 M=1 R=4 SA=125001 SB=125002 A=0.25
+ P=2.5 MULT=1
MM1001 A_359_419# N_A3_M1001_g A_259_419# VPB PHIGHVT L=0.25 W=1 AD=0.16
+ AS=0.125 PD=1.32 PS=1.25 NRD=20.6653 NRS=13.7703 M=1 R=4 SA=125001 SB=125001
+ A=0.25 P=2.5 MULT=1
MM1008 A_473_419# N_A2_M1008_g A_359_419# VPB PHIGHVT L=0.25 W=1 AD=0.16 AS=0.16
+ PD=1.32 PS=1.32 NRD=20.6653 NRS=20.6653 M=1 R=4 SA=125002 SB=125001 A=0.25
+ P=2.5 MULT=1
MM1006 N_VPWR_M1006_d N_A1_M1006_g A_473_419# VPB PHIGHVT L=0.25 W=1 AD=0.285
+ AS=0.16 PD=2.57 PS=1.32 NRD=0 NRS=20.6653 M=1 R=4 SA=125002 SB=125000 A=0.25
+ P=2.5 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9751 P=11.21
*
.include "sky130_fd_sc_lp__o41ai_lp.pxi.spice"
*
.ends
*
*
