# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__einvp_8
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__einvp_8 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.120000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  2.520000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.295000 1.210000 7.245000 1.345000 ;
        RECT 6.295000 1.345000 7.985000 1.595000 ;
    END
  END A
  PIN TE
    ANTENNAGATEAREA  1.323000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.155000 1.210000 0.805000 1.750000 ;
    END
  END TE
  PIN Z
    ANTENNADIFFAREA  2.352000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.685000 1.525000 6.125000 1.765000 ;
        RECT 5.685000 1.765000 8.535000 1.935000 ;
        RECT 5.685000 1.935000 5.915000 2.735000 ;
        RECT 5.755000 0.725000 7.665000 0.995000 ;
        RECT 5.755000 0.995000 6.125000 1.525000 ;
        RECT 6.585000 1.935000 6.775000 2.735000 ;
        RECT 7.415000 0.995000 7.665000 1.005000 ;
        RECT 7.415000 1.005000 8.560000 1.175000 ;
        RECT 7.445000 1.935000 7.635000 2.735000 ;
        RECT 8.155000 1.175000 8.535000 1.765000 ;
        RECT 8.305000 1.935000 8.535000 2.735000 ;
        RECT 8.335000 0.615000 8.560000 1.005000 ;
    END
  END Z
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 9.120000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 9.120000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 9.120000 0.085000 ;
      RECT 0.000000  3.245000 9.120000 3.415000 ;
      RECT 0.455000  1.920000 0.725000 3.245000 ;
      RECT 0.555000  0.085000 0.855000 1.040000 ;
      RECT 0.945000  1.855000 1.315000 1.930000 ;
      RECT 0.945000  1.930000 1.615000 3.075000 ;
      RECT 1.025000  0.255000 1.315000 1.855000 ;
      RECT 1.785000  1.550000 5.515000 1.720000 ;
      RECT 1.785000  1.720000 2.075000 3.075000 ;
      RECT 1.815000  0.255000 2.075000 1.210000 ;
      RECT 1.815000  1.210000 5.585000 1.380000 ;
      RECT 2.245000  0.085000 2.575000 1.040000 ;
      RECT 2.245000  1.890000 2.505000 3.245000 ;
      RECT 2.675000  1.720000 2.935000 3.075000 ;
      RECT 2.745000  0.255000 2.935000 1.210000 ;
      RECT 3.105000  0.085000 3.435000 1.040000 ;
      RECT 3.105000  1.890000 3.370000 3.245000 ;
      RECT 3.540000  1.720000 3.800000 3.075000 ;
      RECT 3.605000  0.255000 3.795000 1.210000 ;
      RECT 3.965000  0.085000 4.295000 1.040000 ;
      RECT 3.970000  1.890000 4.225000 3.245000 ;
      RECT 4.395000  1.720000 4.660000 3.075000 ;
      RECT 4.465000  0.255000 4.685000 1.210000 ;
      RECT 4.830000  1.890000 5.090000 3.245000 ;
      RECT 4.855000  0.085000 5.085000 1.040000 ;
      RECT 5.255000  0.275000 9.025000 0.445000 ;
      RECT 5.255000  0.445000 8.165000 0.555000 ;
      RECT 5.255000  0.555000 5.585000 1.210000 ;
      RECT 5.260000  1.720000 5.515000 2.905000 ;
      RECT 5.260000  2.905000 8.995000 3.075000 ;
      RECT 6.085000  2.105000 6.415000 2.905000 ;
      RECT 6.945000  2.105000 7.275000 2.905000 ;
      RECT 7.805000  2.105000 8.135000 2.905000 ;
      RECT 7.835000  0.555000 8.165000 0.825000 ;
      RECT 8.705000  1.815000 8.995000 2.905000 ;
      RECT 8.730000  0.445000 9.025000 1.095000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
      RECT 8.315000 -0.085000 8.485000 0.085000 ;
      RECT 8.315000  3.245000 8.485000 3.415000 ;
      RECT 8.795000 -0.085000 8.965000 0.085000 ;
      RECT 8.795000  3.245000 8.965000 3.415000 ;
  END
END sky130_fd_sc_lp__einvp_8
