* File: sky130_fd_sc_lp__nand2b_1.pex.spice
* Created: Fri Aug 28 10:47:58 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__NAND2B_1%A_N 3 7 11 13 14 17 18
c31 18 0 3.73553e-20 $X=0.29 $Y=1.1
r32 17 18 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.29 $Y=1.1
+ $X2=0.29 $Y2=1.1
r33 14 18 1.17263 $w=5.08e-07 $l=5e-08 $layer=LI1_cond $X=0.24 $Y=1.27 $X2=0.29
+ $Y2=1.27
r34 12 17 28.3893 $w=4.9e-07 $l=2.6e-07 $layer=POLY_cond $X=0.37 $Y=1.36
+ $X2=0.37 $Y2=1.1
r35 12 13 54.9885 $w=4.9e-07 $l=2.45e-07 $layer=POLY_cond $X=0.37 $Y=1.36
+ $X2=0.37 $Y2=1.605
r36 11 17 16.9244 $w=4.9e-07 $l=1.55e-07 $layer=POLY_cond $X=0.37 $Y=0.945
+ $X2=0.37 $Y2=1.1
r37 10 11 44.6155 $w=4.9e-07 $l=1.5e-07 $layer=POLY_cond $X=0.48 $Y=0.795
+ $X2=0.48 $Y2=0.945
r38 7 10 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=0.76 $Y=0.445
+ $X2=0.76 $Y2=0.795
r39 3 13 225.617 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=0.54 $Y=2.045
+ $X2=0.54 $Y2=1.605
.ends

.subckt PM_SKY130_FD_SC_LP__NAND2B_1%B 3 5 7 8 9 15
c44 3 0 3.73553e-20 $X=1.065 $Y=2.465
r45 13 15 3.48014 $w=2.77e-07 $l=2e-08 $layer=POLY_cond $X=1.045 $Y=1.35
+ $X2=1.065 $Y2=1.35
r46 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.045
+ $Y=1.35 $X2=1.045 $Y2=1.35
r47 9 14 4.25306 $w=4.18e-07 $l=1.55e-07 $layer=LI1_cond $X=1.2 $Y=1.225
+ $X2=1.045 $Y2=1.225
r48 8 14 8.91771 $w=4.18e-07 $l=3.25e-07 $layer=LI1_cond $X=0.72 $Y=1.225
+ $X2=1.045 $Y2=1.225
r49 5 15 35.6715 $w=2.77e-07 $l=2.75409e-07 $layer=POLY_cond $X=1.27 $Y=1.185
+ $X2=1.065 $Y2=1.35
r50 5 7 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.27 $Y=1.185 $X2=1.27
+ $Y2=0.655
r51 1 15 17.1008 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.065 $Y=1.515
+ $X2=1.065 $Y2=1.35
r52 1 3 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=1.065 $Y=1.515
+ $X2=1.065 $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__NAND2B_1%A_40_367# 1 2 9 12 15 16 17 20 24 26 27 28
+ 29 31 34 35
r81 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.735
+ $Y=1.44 $X2=1.735 $Y2=1.44
r82 31 34 8.99492 $w=3.54e-07 $l=2.23226e-07 $layer=LI1_cond $X=1.54 $Y=1.275
+ $X2=1.677 $Y2=1.44
r83 30 31 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=1.54 $Y=0.845
+ $X2=1.54 $Y2=1.275
r84 28 34 8.61582 $w=3.54e-07 $l=3.43511e-07 $layer=LI1_cond $X=1.455 $Y=1.69
+ $X2=1.677 $Y2=1.44
r85 28 29 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=1.455 $Y=1.69
+ $X2=0.78 $Y2=1.69
r86 26 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.455 $Y=0.76
+ $X2=1.54 $Y2=0.845
r87 26 27 53.1711 $w=1.68e-07 $l=8.15e-07 $layer=LI1_cond $X=1.455 $Y=0.76
+ $X2=0.64 $Y2=0.76
r88 22 27 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=0.51 $Y=0.675
+ $X2=0.64 $Y2=0.76
r89 22 24 10.1947 $w=2.58e-07 $l=2.3e-07 $layer=LI1_cond $X=0.51 $Y=0.675
+ $X2=0.51 $Y2=0.445
r90 18 29 28.8317 $w=1.94e-07 $l=4.7697e-07 $layer=LI1_cond $X=0.325 $Y=1.735
+ $X2=0.78 $Y2=1.69
r91 18 20 6.28605 $w=3.28e-07 $l=1.8e-07 $layer=LI1_cond $X=0.325 $Y=1.865
+ $X2=0.325 $Y2=2.045
r92 16 35 13.8825 $w=3.45e-07 $l=8.3e-08 $layer=POLY_cond $X=1.727 $Y=1.357
+ $X2=1.727 $Y2=1.44
r93 16 17 47.5363 $w=3.45e-07 $l=1.72e-07 $layer=POLY_cond $X=1.727 $Y=1.357
+ $X2=1.727 $Y2=1.185
r94 14 35 22.5799 $w=3.45e-07 $l=1.35e-07 $layer=POLY_cond $X=1.727 $Y=1.575
+ $X2=1.727 $Y2=1.44
r95 14 15 43.8566 $w=3.45e-07 $l=1.5e-07 $layer=POLY_cond $X=1.66 $Y=1.575
+ $X2=1.66 $Y2=1.725
r96 12 17 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.63 $Y=0.655
+ $X2=1.63 $Y2=1.185
r97 9 15 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=1.495 $Y=2.465
+ $X2=1.495 $Y2=1.725
r98 2 20 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=0.2
+ $Y=1.835 $X2=0.325 $Y2=2.045
r99 1 24 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.42
+ $Y=0.235 $X2=0.545 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__NAND2B_1%VPWR 1 2 11 17 19 21 28 29 32 35
r25 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r26 32 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r27 29 36 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r28 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r29 26 35 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.875 $Y=3.33
+ $X2=1.71 $Y2=3.33
r30 26 28 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.875 $Y=3.33
+ $X2=2.16 $Y2=3.33
r31 22 32 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.945 $Y=3.33
+ $X2=0.815 $Y2=3.33
r32 22 24 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.945 $Y=3.33
+ $X2=1.2 $Y2=3.33
r33 21 35 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.545 $Y=3.33
+ $X2=1.71 $Y2=3.33
r34 21 24 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.545 $Y=3.33
+ $X2=1.2 $Y2=3.33
r35 19 36 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r36 19 33 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r37 19 24 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r38 15 35 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.71 $Y=3.245
+ $X2=1.71 $Y2=3.33
r39 15 17 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=1.71 $Y=3.245
+ $X2=1.71 $Y2=2.415
r40 11 14 33.2435 $w=2.58e-07 $l=7.5e-07 $layer=LI1_cond $X=0.815 $Y=2.2
+ $X2=0.815 $Y2=2.95
r41 9 32 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=0.815 $Y=3.245
+ $X2=0.815 $Y2=3.33
r42 9 14 13.0758 $w=2.58e-07 $l=2.95e-07 $layer=LI1_cond $X=0.815 $Y=3.245
+ $X2=0.815 $Y2=2.95
r43 2 17 300 $w=1.7e-07 $l=6.4622e-07 $layer=licon1_PDIFF $count=2 $X=1.57
+ $Y=1.835 $X2=1.71 $Y2=2.415
r44 1 14 400 $w=1.7e-07 $l=1.22689e-06 $layer=licon1_PDIFF $count=1 $X=0.615
+ $Y=1.835 $X2=0.85 $Y2=2.95
r45 1 11 400 $w=1.7e-07 $l=4.67974e-07 $layer=licon1_PDIFF $count=1 $X=0.615
+ $Y=1.835 $X2=0.85 $Y2=2.2
.ends

.subckt PM_SKY130_FD_SC_LP__NAND2B_1%Y 1 2 7 11 14 15 18 19 20
r31 19 20 16.4002 $w=2.58e-07 $l=3.7e-07 $layer=LI1_cond $X=1.245 $Y=2.405
+ $X2=1.245 $Y2=2.775
r32 15 19 12.8542 $w=2.58e-07 $l=2.9e-07 $layer=LI1_cond $X=1.245 $Y=2.115
+ $X2=1.245 $Y2=2.405
r33 15 17 2.85134 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=1.245 $Y=2.115
+ $X2=1.245 $Y2=2.03
r34 14 18 39.9827 $w=2.43e-07 $l=8.5e-07 $layer=LI1_cond $X=2.192 $Y=1.945
+ $X2=2.192 $Y2=1.095
r35 9 18 9.34621 $w=5.18e-07 $l=2.6e-07 $layer=LI1_cond $X=2.055 $Y=0.835
+ $X2=2.055 $Y2=1.095
r36 9 11 9.54563 $w=5.18e-07 $l=4.15e-07 $layer=LI1_cond $X=2.055 $Y=0.835
+ $X2=2.055 $Y2=0.42
r37 8 17 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.375 $Y=2.03
+ $X2=1.245 $Y2=2.03
r38 7 14 7.11011 $w=1.7e-07 $l=1.58915e-07 $layer=LI1_cond $X=2.07 $Y=2.03
+ $X2=2.192 $Y2=1.945
r39 7 8 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=2.07 $Y=2.03
+ $X2=1.375 $Y2=2.03
r40 2 19 300 $w=1.7e-07 $l=7.06541e-07 $layer=licon1_PDIFF $count=2 $X=1.14
+ $Y=1.835 $X2=1.28 $Y2=2.475
r41 2 17 600 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_PDIFF $count=1 $X=1.14
+ $Y=1.835 $X2=1.28 $Y2=2.03
r42 1 11 91 $w=1.7e-07 $l=2.5807e-07 $layer=licon1_NDIFF $count=2 $X=1.705
+ $Y=0.235 $X2=1.88 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__NAND2B_1%VGND 1 6 9 10 11 21 22
r27 21 22 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r28 18 21 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r29 14 15 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r30 11 22 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r31 11 15 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r32 11 18 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r33 9 14 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=0.81 $Y=0 $X2=0.72
+ $Y2=0
r34 9 10 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.81 $Y=0 $X2=0.975
+ $Y2=0
r35 8 18 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=1.14 $Y=0 $X2=1.2 $Y2=0
r36 8 10 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.14 $Y=0 $X2=0.975
+ $Y2=0
r37 4 10 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.975 $Y=0.085
+ $X2=0.975 $Y2=0
r38 4 6 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.975 $Y=0.085
+ $X2=0.975 $Y2=0.38
r39 1 6 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=0.835
+ $Y=0.235 $X2=0.975 $Y2=0.38
.ends

