* File: sky130_fd_sc_lp__nor2_lp.pxi.spice
* Created: Fri Aug 28 10:54:05 2020
* 
x_PM_SKY130_FD_SC_LP__NOR2_LP%A N_A_M1000_g N_A_M1004_g N_A_c_38_n N_A_M1002_g
+ N_A_c_40_n N_A_c_44_n A A A N_A_c_42_n PM_SKY130_FD_SC_LP__NOR2_LP%A
x_PM_SKY130_FD_SC_LP__NOR2_LP%B N_B_M1005_g N_B_c_80_n N_B_c_81_n N_B_M1003_g
+ N_B_c_83_n N_B_M1001_g N_B_c_84_n N_B_c_76_n B B B B B N_B_c_78_n
+ PM_SKY130_FD_SC_LP__NOR2_LP%B
x_PM_SKY130_FD_SC_LP__NOR2_LP%VPB__2 N_VPB__2_M1004_s N_VPB__2_c_116_n
+ N_VPB__2_c_117_n VPB__2 N_VPB__2_c_118_n N_VPB__2_c_115_n
+ PM_SKY130_FD_SC_LP__NOR2_LP%VPB__2
x_PM_SKY130_FD_SC_LP__NOR2_LP%Y N_Y_M1002_d N_Y_M1005_d Y Y Y Y Y Y Y
+ PM_SKY130_FD_SC_LP__NOR2_LP%Y
x_PM_SKY130_FD_SC_LP__NOR2_LP%VNB__2 N_VNB__2_M1000_s N_VNB__2_M1001_d
+ N_VNB__2_c_157_n N_VNB__2_c_158_n N_VNB__2_c_159_n N_VNB__2_c_160_n VNB__2
+ N_VNB__2_c_161_n N_VNB__2_c_162_n PM_SKY130_FD_SC_LP__NOR2_LP%VNB__2
cc_1 VNB N_A_M1000_g 0.0274458f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=0.77
cc_2 VNB N_A_c_38_n 0.0215151f $X=-0.19 $Y=-0.245 $X2=0.89 $Y2=1.255
cc_3 VNB N_A_M1002_g 0.0192706f $X=-0.19 $Y=-0.245 $X2=0.965 $Y2=0.77
cc_4 VNB N_A_c_40_n 0.0146721f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=1.255
cc_5 VNB A 0.03032f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_6 VNB N_A_c_42_n 0.0281728f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=1.345
cc_7 VNB N_B_M1003_g 0.0438648f $X=-0.19 $Y=-0.245 $X2=0.89 $Y2=1.255
cc_8 VNB N_B_M1001_g 0.0274458f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=1.33
cc_9 VNB N_B_c_76_n 0.0232141f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_10 VNB B 0.0367255f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.95
cc_11 VNB N_B_c_78_n 0.0175337f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=2.035
cc_12 VNB N_VPB__2_c_115_n 0.103974f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=1.255
cc_13 VNB Y 0.00506809f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=2.66
cc_14 VNB N_VNB__2_c_157_n 0.0147687f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=2.66
cc_15 VNB N_VNB__2_c_158_n 0.0452369f $X=-0.19 $Y=-0.245 $X2=0.89 $Y2=1.255
cc_16 VNB N_VNB__2_c_159_n 0.0160446f $X=-0.19 $Y=-0.245 $X2=0.965 $Y2=1.18
cc_17 VNB N_VNB__2_c_160_n 0.0452369f $X=-0.19 $Y=-0.245 $X2=0.965 $Y2=0.77
cc_18 VNB N_VNB__2_c_161_n 0.039476f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=1.685
cc_19 VNB N_VNB__2_c_162_n 0.18881f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VPB N_A_M1004_g 0.052723f $X=-0.19 $Y=1.655 $X2=0.575 $Y2=2.66
cc_21 VPB N_A_c_44_n 0.0177236f $X=-0.19 $Y=1.655 $X2=0.485 $Y2=1.85
cc_22 VPB A 0.0382317f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_23 VPB N_A_c_42_n 0.00252164f $X=-0.19 $Y=1.655 $X2=0.485 $Y2=1.345
cc_24 VPB N_B_M1005_g 0.0513092f $X=-0.19 $Y=1.655 $X2=0.575 $Y2=0.77
cc_25 VPB N_B_c_80_n 0.020349f $X=-0.19 $Y=1.655 $X2=0.575 $Y2=1.85
cc_26 VPB N_B_c_81_n 0.00846326f $X=-0.19 $Y=1.655 $X2=0.575 $Y2=2.66
cc_27 VPB N_B_M1003_g 0.00241318f $X=-0.19 $Y=1.655 $X2=0.89 $Y2=1.255
cc_28 VPB N_B_c_83_n 0.0338589f $X=-0.19 $Y=1.655 $X2=0.965 $Y2=1.18
cc_29 VPB N_B_c_84_n 0.0100371f $X=-0.19 $Y=1.655 $X2=0.485 $Y2=1.685
cc_30 VPB N_B_c_76_n 0.00330557f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_31 VPB B 0.0895781f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.95
cc_32 VPB N_VPB__2_c_116_n 0.0147428f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_33 VPB N_VPB__2_c_117_n 0.0372899f $X=-0.19 $Y=1.655 $X2=0.575 $Y2=2.66
cc_34 VPB N_VPB__2_c_118_n 0.0550275f $X=-0.19 $Y=1.655 $X2=0.485 $Y2=1.33
cc_35 VPB N_VPB__2_c_115_n 0.0821532f $X=-0.19 $Y=1.655 $X2=0.485 $Y2=1.255
cc_36 VPB Y 0.0162488f $X=-0.19 $Y=1.655 $X2=0.575 $Y2=2.66
cc_37 N_A_M1004_g N_B_M1005_g 0.0330137f $X=0.575 $Y=2.66 $X2=0 $Y2=0
cc_38 N_A_c_38_n N_B_c_81_n 0.00706287f $X=0.89 $Y=1.255 $X2=0 $Y2=0
cc_39 N_A_c_44_n N_B_c_81_n 0.0330137f $X=0.485 $Y=1.85 $X2=0 $Y2=0
cc_40 A N_B_c_81_n 0.00371338f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_41 N_A_M1002_g N_B_M1003_g 0.0230493f $X=0.965 $Y=0.77 $X2=0 $Y2=0
cc_42 A N_B_M1003_g 0.0010466f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_43 N_A_c_42_n N_B_M1003_g 0.00394668f $X=0.485 $Y=1.345 $X2=0 $Y2=0
cc_44 N_A_M1004_g N_VPB__2_c_117_n 0.0141994f $X=0.575 $Y=2.66 $X2=0 $Y2=0
cc_45 N_A_c_44_n N_VPB__2_c_117_n 7.66517e-19 $X=0.485 $Y=1.85 $X2=0 $Y2=0
cc_46 A N_VPB__2_c_117_n 0.0214312f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_47 N_A_M1004_g N_VPB__2_c_118_n 0.00426961f $X=0.575 $Y=2.66 $X2=0 $Y2=0
cc_48 N_A_M1004_g N_VPB__2_c_115_n 0.00434697f $X=0.575 $Y=2.66 $X2=0 $Y2=0
cc_49 N_A_M1000_g Y 0.00247239f $X=0.575 $Y=0.77 $X2=0 $Y2=0
cc_50 N_A_M1004_g Y 0.00268998f $X=0.575 $Y=2.66 $X2=0 $Y2=0
cc_51 N_A_c_38_n Y 0.00466605f $X=0.89 $Y=1.255 $X2=0 $Y2=0
cc_52 N_A_M1002_g Y 0.0167795f $X=0.965 $Y=0.77 $X2=0 $Y2=0
cc_53 N_A_c_44_n Y 3.45973e-19 $X=0.485 $Y=1.85 $X2=0 $Y2=0
cc_54 A Y 0.0791063f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_55 N_A_c_42_n Y 0.00107551f $X=0.485 $Y=1.345 $X2=0 $Y2=0
cc_56 N_A_M1000_g N_VNB__2_c_158_n 0.0140129f $X=0.575 $Y=0.77 $X2=0 $Y2=0
cc_57 N_A_M1002_g N_VNB__2_c_158_n 0.00163467f $X=0.965 $Y=0.77 $X2=0 $Y2=0
cc_58 N_A_c_40_n N_VNB__2_c_158_n 0.00139912f $X=0.485 $Y=1.255 $X2=0 $Y2=0
cc_59 A N_VNB__2_c_158_n 0.028459f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_60 N_A_M1000_g N_VNB__2_c_161_n 0.00375057f $X=0.575 $Y=0.77 $X2=0 $Y2=0
cc_61 N_A_M1002_g N_VNB__2_c_161_n 0.0043233f $X=0.965 $Y=0.77 $X2=0 $Y2=0
cc_62 N_A_M1000_g N_VNB__2_c_162_n 0.00409726f $X=0.575 $Y=0.77 $X2=0 $Y2=0
cc_63 N_A_M1002_g N_VNB__2_c_162_n 0.00487769f $X=0.965 $Y=0.77 $X2=0 $Y2=0
cc_64 N_B_M1005_g N_VPB__2_c_117_n 0.0018473f $X=0.965 $Y=2.66 $X2=0 $Y2=0
cc_65 N_B_M1005_g N_VPB__2_c_118_n 0.00491683f $X=0.965 $Y=2.66 $X2=0 $Y2=0
cc_66 B N_VPB__2_c_118_n 0.0231512f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_67 N_B_M1005_g N_VPB__2_c_115_n 0.00517496f $X=0.965 $Y=2.66 $X2=0 $Y2=0
cc_68 B N_VPB__2_c_115_n 0.0246855f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_69 N_B_M1005_g Y 0.0291017f $X=0.965 $Y=2.66 $X2=0 $Y2=0
cc_70 N_B_c_80_n Y 0.0173207f $X=1.32 $Y=1.775 $X2=0 $Y2=0
cc_71 N_B_c_81_n Y 0.00190972f $X=1.04 $Y=1.775 $X2=0 $Y2=0
cc_72 N_B_M1003_g Y 0.0305535f $X=1.395 $Y=0.77 $X2=0 $Y2=0
cc_73 N_B_M1001_g Y 0.00247533f $X=1.785 $Y=0.77 $X2=0 $Y2=0
cc_74 N_B_c_84_n Y 0.00336398f $X=1.395 $Y=1.775 $X2=0 $Y2=0
cc_75 B Y 0.122588f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_76 N_B_c_78_n Y 4.31827e-19 $X=1.875 $Y=1.345 $X2=0 $Y2=0
cc_77 N_B_M1003_g N_VNB__2_c_160_n 0.00163467f $X=1.395 $Y=0.77 $X2=0 $Y2=0
cc_78 N_B_M1001_g N_VNB__2_c_160_n 0.0140129f $X=1.785 $Y=0.77 $X2=0 $Y2=0
cc_79 B N_VNB__2_c_160_n 0.028459f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_80 N_B_c_78_n N_VNB__2_c_160_n 0.00139912f $X=1.875 $Y=1.345 $X2=0 $Y2=0
cc_81 N_B_M1003_g N_VNB__2_c_161_n 0.0043233f $X=1.395 $Y=0.77 $X2=0 $Y2=0
cc_82 N_B_M1001_g N_VNB__2_c_161_n 0.00375057f $X=1.785 $Y=0.77 $X2=0 $Y2=0
cc_83 N_B_M1003_g N_VNB__2_c_162_n 0.00487769f $X=1.395 $Y=0.77 $X2=0 $Y2=0
cc_84 N_B_M1001_g N_VNB__2_c_162_n 0.00409726f $X=1.785 $Y=0.77 $X2=0 $Y2=0
cc_85 N_VPB__2_c_117_n Y 0.0145731f $X=0.36 $Y=2.66 $X2=0 $Y2=0
cc_86 N_VPB__2_c_118_n Y 0.0106618f $X=2.16 $Y=3.33 $X2=0 $Y2=0
cc_87 N_VPB__2_c_115_n Y 0.0114128f $X=2.16 $Y=3.33 $X2=0 $Y2=0
cc_88 Y N_VNB__2_c_158_n 0.0177412f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_89 Y N_VNB__2_c_160_n 0.0177412f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_90 Y N_VNB__2_c_161_n 0.0105983f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_91 Y N_VNB__2_c_162_n 0.0113894f $X=1.115 $Y=0.47 $X2=0 $Y2=0
