* File: sky130_fd_sc_lp__nor4bb_4.pxi.spice
* Created: Fri Aug 28 10:59:11 2020
* 
x_PM_SKY130_FD_SC_LP__NOR4BB_4%D_N N_D_N_M1015_g N_D_N_M1032_g D_N N_D_N_c_161_n
+ N_D_N_c_162_n PM_SKY130_FD_SC_LP__NOR4BB_4%D_N
x_PM_SKY130_FD_SC_LP__NOR4BB_4%C_N N_C_N_M1028_g N_C_N_M1010_g C_N N_C_N_c_185_n
+ N_C_N_c_186_n PM_SKY130_FD_SC_LP__NOR4BB_4%C_N
x_PM_SKY130_FD_SC_LP__NOR4BB_4%A_37_51# N_A_37_51#_M1015_s N_A_37_51#_M1032_s
+ N_A_37_51#_M1002_g N_A_37_51#_M1005_g N_A_37_51#_M1009_g N_A_37_51#_M1012_g
+ N_A_37_51#_M1019_g N_A_37_51#_M1026_g N_A_37_51#_M1030_g N_A_37_51#_M1029_g
+ N_A_37_51#_c_221_n N_A_37_51#_c_232_n N_A_37_51#_c_222_n N_A_37_51#_c_223_n
+ N_A_37_51#_c_224_n N_A_37_51#_c_234_n N_A_37_51#_c_225_n N_A_37_51#_c_235_n
+ N_A_37_51#_c_226_n N_A_37_51#_c_236_n N_A_37_51#_c_227_n
+ PM_SKY130_FD_SC_LP__NOR4BB_4%A_37_51#
x_PM_SKY130_FD_SC_LP__NOR4BB_4%A_206_51# N_A_206_51#_M1028_d N_A_206_51#_M1010_d
+ N_A_206_51#_M1001_g N_A_206_51#_M1000_g N_A_206_51#_M1007_g
+ N_A_206_51#_M1004_g N_A_206_51#_M1013_g N_A_206_51#_M1022_g
+ N_A_206_51#_M1027_g N_A_206_51#_M1034_g N_A_206_51#_c_369_n
+ N_A_206_51#_c_359_n N_A_206_51#_c_360_n N_A_206_51#_c_361_n
+ N_A_206_51#_c_362_n N_A_206_51#_c_440_p N_A_206_51#_c_363_n
+ N_A_206_51#_c_364_n PM_SKY130_FD_SC_LP__NOR4BB_4%A_206_51#
x_PM_SKY130_FD_SC_LP__NOR4BB_4%B N_B_M1008_g N_B_M1006_g N_B_M1014_g N_B_M1023_g
+ N_B_M1021_g N_B_M1024_g N_B_M1033_g N_B_M1035_g N_B_c_508_n B N_B_c_509_n
+ N_B_c_510_n PM_SKY130_FD_SC_LP__NOR4BB_4%B
x_PM_SKY130_FD_SC_LP__NOR4BB_4%A N_A_M1016_g N_A_M1003_g N_A_M1017_g N_A_M1011_g
+ N_A_M1018_g N_A_M1020_g N_A_M1031_g N_A_M1025_g A A A A N_A_c_616_n
+ N_A_c_617_n PM_SKY130_FD_SC_LP__NOR4BB_4%A
x_PM_SKY130_FD_SC_LP__NOR4BB_4%VPWR N_VPWR_M1032_d N_VPWR_M1003_d N_VPWR_M1020_d
+ N_VPWR_c_685_n N_VPWR_c_686_n N_VPWR_c_687_n VPWR N_VPWR_c_688_n
+ N_VPWR_c_689_n N_VPWR_c_690_n N_VPWR_c_691_n N_VPWR_c_684_n N_VPWR_c_693_n
+ N_VPWR_c_694_n N_VPWR_c_695_n PM_SKY130_FD_SC_LP__NOR4BB_4%VPWR
x_PM_SKY130_FD_SC_LP__NOR4BB_4%A_347_349# N_A_347_349#_M1005_d
+ N_A_347_349#_M1012_d N_A_347_349#_M1030_d N_A_347_349#_M1007_s
+ N_A_347_349#_M1027_s N_A_347_349#_c_789_n N_A_347_349#_c_799_n
+ N_A_347_349#_c_790_n N_A_347_349#_c_833_p N_A_347_349#_c_811_n
+ N_A_347_349#_c_844_p N_A_347_349#_c_813_n N_A_347_349#_c_791_n
+ N_A_347_349#_c_792_n N_A_347_349#_c_836_p N_A_347_349#_c_793_n
+ PM_SKY130_FD_SC_LP__NOR4BB_4%A_347_349#
x_PM_SKY130_FD_SC_LP__NOR4BB_4%Y N_Y_M1002_s N_Y_M1026_s N_Y_M1000_d N_Y_M1022_d
+ N_Y_M1006_s N_Y_M1024_s N_Y_M1016_d N_Y_M1018_d N_Y_M1005_s N_Y_M1019_s
+ N_Y_c_868_n N_Y_c_960_n N_Y_c_871_n N_Y_c_873_n N_Y_c_862_n N_Y_c_863_n
+ N_Y_c_883_n N_Y_c_963_n N_Y_c_864_n N_Y_c_889_n N_Y_c_1003_p N_Y_c_851_n
+ N_Y_c_852_n N_Y_c_1004_p N_Y_c_853_n N_Y_c_854_n N_Y_c_999_p N_Y_c_855_n
+ N_Y_c_995_p N_Y_c_856_n N_Y_c_1005_p N_Y_c_857_n N_Y_c_1006_p N_Y_c_890_n
+ N_Y_c_865_n N_Y_c_858_n N_Y_c_859_n N_Y_c_860_n Y Y N_Y_c_867_n Y
+ PM_SKY130_FD_SC_LP__NOR4BB_4%Y
x_PM_SKY130_FD_SC_LP__NOR4BB_4%A_774_349# N_A_774_349#_M1001_d
+ N_A_774_349#_M1013_d N_A_774_349#_M1008_s N_A_774_349#_M1021_s
+ N_A_774_349#_c_1029_n N_A_774_349#_c_1025_n N_A_774_349#_c_1026_n
+ N_A_774_349#_c_1036_n N_A_774_349#_c_1027_n N_A_774_349#_c_1043_n
+ N_A_774_349#_c_1046_n N_A_774_349#_c_1048_n N_A_774_349#_c_1050_n
+ N_A_774_349#_c_1028_n N_A_774_349#_c_1053_n
+ PM_SKY130_FD_SC_LP__NOR4BB_4%A_774_349#
x_PM_SKY130_FD_SC_LP__NOR4BB_4%A_1139_367# N_A_1139_367#_M1008_d
+ N_A_1139_367#_M1014_d N_A_1139_367#_M1033_d N_A_1139_367#_M1011_s
+ N_A_1139_367#_M1025_s N_A_1139_367#_c_1090_n N_A_1139_367#_c_1091_n
+ N_A_1139_367#_c_1099_n N_A_1139_367#_c_1104_n N_A_1139_367#_c_1155_n
+ N_A_1139_367#_c_1092_n N_A_1139_367#_c_1093_n N_A_1139_367#_c_1094_n
+ N_A_1139_367#_c_1137_n N_A_1139_367#_c_1120_n N_A_1139_367#_c_1141_n
+ N_A_1139_367#_c_1124_n N_A_1139_367#_c_1095_n N_A_1139_367#_c_1096_n
+ N_A_1139_367#_c_1117_n N_A_1139_367#_c_1130_n
+ PM_SKY130_FD_SC_LP__NOR4BB_4%A_1139_367#
x_PM_SKY130_FD_SC_LP__NOR4BB_4%VGND N_VGND_M1015_d N_VGND_M1002_d N_VGND_M1009_d
+ N_VGND_M1029_d N_VGND_M1004_s N_VGND_M1034_s N_VGND_M1023_d N_VGND_M1035_d
+ N_VGND_M1017_s N_VGND_M1031_s N_VGND_c_1158_n N_VGND_c_1159_n N_VGND_c_1160_n
+ N_VGND_c_1161_n N_VGND_c_1162_n N_VGND_c_1163_n N_VGND_c_1164_n
+ N_VGND_c_1165_n N_VGND_c_1166_n N_VGND_c_1167_n N_VGND_c_1168_n
+ N_VGND_c_1169_n N_VGND_c_1170_n N_VGND_c_1171_n N_VGND_c_1172_n VGND
+ N_VGND_c_1173_n N_VGND_c_1174_n N_VGND_c_1175_n N_VGND_c_1176_n
+ N_VGND_c_1177_n N_VGND_c_1178_n N_VGND_c_1179_n N_VGND_c_1180_n
+ N_VGND_c_1181_n N_VGND_c_1182_n N_VGND_c_1183_n N_VGND_c_1184_n
+ N_VGND_c_1185_n N_VGND_c_1186_n N_VGND_c_1187_n N_VGND_c_1188_n
+ PM_SKY130_FD_SC_LP__NOR4BB_4%VGND
cc_1 VNB N_D_N_M1015_g 0.0270926f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=0.675
cc_2 VNB N_D_N_M1032_g 0.00183793f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=2.465
cc_3 VNB N_D_N_c_161_n 0.012893f $X=-0.19 $Y=-0.245 $X2=0.31 $Y2=1.46
cc_4 VNB N_D_N_c_162_n 0.049553f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.46
cc_5 VNB N_C_N_M1028_g 0.0279106f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=0.675
cc_6 VNB N_C_N_c_185_n 0.0319063f $X=-0.19 $Y=-0.245 $X2=0.31 $Y2=1.46
cc_7 VNB N_C_N_c_186_n 0.0060767f $X=-0.19 $Y=-0.245 $X2=0.31 $Y2=1.46
cc_8 VNB N_A_37_51#_M1002_g 0.0234929f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_9 VNB N_A_37_51#_M1009_g 0.0207899f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=1.46
cc_10 VNB N_A_37_51#_M1026_g 0.0208069f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_37_51#_M1029_g 0.0199381f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_37_51#_c_221_n 0.0306079f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_37_51#_c_222_n 0.00270301f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_37_51#_c_223_n 0.00900805f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_37_51#_c_224_n 0.00835541f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_37_51#_c_225_n 0.00141487f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_37_51#_c_226_n 0.00118898f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_37_51#_c_227_n 0.0805856f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_206_51#_M1000_g 0.019586f $X=-0.19 $Y=-0.245 $X2=0.31 $Y2=1.46
cc_20 VNB N_A_206_51#_M1004_g 0.0187554f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_206_51#_M1022_g 0.0187545f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_206_51#_M1034_g 0.0214498f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_206_51#_c_359_n 0.00986993f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_206_51#_c_360_n 0.0102566f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_206_51#_c_361_n 0.0180978f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_206_51#_c_362_n 0.00206836f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_206_51#_c_363_n 0.0181099f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_206_51#_c_364_n 0.0737507f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_B_M1008_g 0.00283446f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=0.675
cc_30 VNB N_B_M1006_g 0.0231921f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=2.465
cc_31 VNB N_B_M1014_g 0.00248075f $X=-0.19 $Y=-0.245 $X2=0.31 $Y2=1.46
cc_32 VNB N_B_M1023_g 0.0197131f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.46
cc_33 VNB N_B_M1021_g 0.00249114f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=1.665
cc_34 VNB N_B_M1024_g 0.0197131f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_B_M1033_g 0.00258021f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_B_M1035_g 0.0198996f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_B_c_508_n 0.00138429f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_B_c_509_n 9.26646e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_B_c_510_n 0.0995349f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_M1016_g 0.0208975f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=0.675
cc_41 VNB N_A_M1003_g 0.00140842f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=2.465
cc_42 VNB N_A_M1017_g 0.0207302f $X=-0.19 $Y=-0.245 $X2=0.31 $Y2=1.46
cc_43 VNB N_A_M1011_g 0.00123234f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.46
cc_44 VNB N_A_M1018_g 0.0207302f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=1.665
cc_45 VNB N_A_M1020_g 0.00123234f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_M1031_g 0.0303822f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_M1025_g 0.00167754f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB A 0.011363f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_c_616_n 0.0717602f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_c_617_n 0.0461398f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_VPWR_c_684_n 0.40251f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_Y_c_851_n 0.00304538f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_Y_c_852_n 0.00203369f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_Y_c_853_n 0.00798225f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_Y_c_854_n 0.00264459f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_Y_c_855_n 0.00310505f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_Y_c_856_n 0.00555338f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_Y_c_857_n 0.00639798f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_Y_c_858_n 0.00145984f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_Y_c_859_n 0.00147023f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_Y_c_860_n 0.00152782f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB Y 0.00572348f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_VGND_c_1158_n 8.4979e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_VGND_c_1159_n 0.0105942f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_VGND_c_1160_n 0.0055866f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_VGND_c_1161_n 0.017028f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_1162_n 0.00269882f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_VGND_c_1163_n 3.0911e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_VGND_c_1164_n 0.00198997f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_VGND_c_1165_n 3.0911e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_VGND_c_1166_n 0.0129398f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_VGND_c_1167_n 3.0911e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_VGND_c_1168_n 3.15212e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_VGND_c_1169_n 0.013298f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_VGND_c_1170_n 0.0398497f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_VGND_c_1171_n 0.0129398f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_VGND_c_1172_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_VGND_c_1173_n 0.0171927f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_VGND_c_1174_n 0.0163237f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_VGND_c_1175_n 0.0174355f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_VGND_c_1176_n 0.0122054f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_VGND_c_1177_n 0.0129398f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_VGND_c_1178_n 0.0129398f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_VGND_c_1179_n 0.0147711f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_VGND_c_1180_n 0.00463869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_VGND_c_1181_n 0.00634414f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_VGND_c_1182_n 0.0063123f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_VGND_c_1183_n 0.00509914f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_VGND_c_1184_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_VGND_c_1185_n 0.0113265f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_VGND_c_1186_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_VGND_c_1187_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_93 VNB N_VGND_c_1188_n 0.468024f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_94 VPB N_D_N_M1032_g 0.0259114f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=2.465
cc_95 VPB N_D_N_c_161_n 0.00907257f $X=-0.19 $Y=1.655 $X2=0.31 $Y2=1.46
cc_96 VPB N_C_N_M1010_g 0.0230553f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=2.465
cc_97 VPB N_C_N_c_185_n 0.00818654f $X=-0.19 $Y=1.655 $X2=0.31 $Y2=1.46
cc_98 VPB N_C_N_c_186_n 0.00333865f $X=-0.19 $Y=1.655 $X2=0.31 $Y2=1.46
cc_99 VPB N_A_37_51#_M1005_g 0.0228713f $X=-0.19 $Y=1.655 $X2=0.31 $Y2=1.46
cc_100 VPB N_A_37_51#_M1012_g 0.0182288f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_101 VPB N_A_37_51#_M1019_g 0.0182361f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_102 VPB N_A_37_51#_M1030_g 0.0184586f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_103 VPB N_A_37_51#_c_232_n 0.0227891f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_104 VPB N_A_37_51#_c_224_n 0.00326617f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_105 VPB N_A_37_51#_c_234_n 0.0165836f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_106 VPB N_A_37_51#_c_235_n 0.00134889f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_107 VPB N_A_37_51#_c_236_n 0.0234997f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_108 VPB N_A_37_51#_c_227_n 0.0187225f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_109 VPB N_A_206_51#_M1001_g 0.0188572f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_110 VPB N_A_206_51#_M1007_g 0.0182361f $X=-0.19 $Y=1.655 $X2=0.28 $Y2=1.46
cc_111 VPB N_A_206_51#_M1013_g 0.0182153f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_112 VPB N_A_206_51#_M1027_g 0.0220207f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_113 VPB N_A_206_51#_c_369_n 0.0128185f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_114 VPB N_A_206_51#_c_360_n 0.00716508f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_115 VPB N_A_206_51#_c_364_n 0.0153611f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_116 VPB N_B_M1008_g 0.0237252f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=0.675
cc_117 VPB N_B_M1014_g 0.0192166f $X=-0.19 $Y=1.655 $X2=0.31 $Y2=1.46
cc_118 VPB N_B_M1021_g 0.018641f $X=-0.19 $Y=1.655 $X2=0.28 $Y2=1.665
cc_119 VPB N_B_M1033_g 0.0189012f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_120 VPB N_B_c_509_n 0.00548176f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_121 VPB N_A_M1003_g 0.0195552f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=2.465
cc_122 VPB N_A_M1011_g 0.0187443f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=1.46
cc_123 VPB N_A_M1020_g 0.0187475f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_124 VPB N_A_M1025_g 0.0252427f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_125 VPB A 0.017364f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_126 VPB N_VPWR_c_685_n 4.89148e-19 $X=-0.19 $Y=1.655 $X2=0.31 $Y2=1.46
cc_127 VPB N_VPWR_c_686_n 3.99129e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_128 VPB N_VPWR_c_687_n 3.99129e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_129 VPB N_VPWR_c_688_n 0.016967f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_130 VPB N_VPWR_c_689_n 0.163262f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_131 VPB N_VPWR_c_690_n 0.0129398f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_132 VPB N_VPWR_c_691_n 0.0177625f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_133 VPB N_VPWR_c_684_n 0.0786764f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_134 VPB N_VPWR_c_693_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_135 VPB N_VPWR_c_694_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_136 VPB N_VPWR_c_695_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_137 VPB N_A_347_349#_c_789_n 0.00199363f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_138 VPB N_A_347_349#_c_790_n 0.00421819f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_139 VPB N_A_347_349#_c_791_n 0.0101958f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_140 VPB N_A_347_349#_c_792_n 0.00203831f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_141 VPB N_A_347_349#_c_793_n 0.00674148f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_142 VPB N_Y_c_862_n 0.00304705f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_143 VPB N_Y_c_863_n 0.00187832f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_144 VPB N_Y_c_864_n 0.010918f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_145 VPB N_Y_c_865_n 0.00181876f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_146 VPB Y 0.00174402f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_147 VPB N_Y_c_867_n 0.00895015f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_148 VPB N_A_774_349#_c_1025_n 0.00199363f $X=-0.19 $Y=1.655 $X2=0.28 $Y2=1.46
cc_149 VPB N_A_774_349#_c_1026_n 0.00203932f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_150 VPB N_A_774_349#_c_1027_n 0.0133143f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_151 VPB N_A_774_349#_c_1028_n 0.00203932f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_152 VPB N_A_1139_367#_c_1090_n 0.00310887f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_153 VPB N_A_1139_367#_c_1091_n 0.00485547f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_154 VPB N_A_1139_367#_c_1092_n 0.00295483f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_155 VPB N_A_1139_367#_c_1093_n 0.00189886f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_156 VPB N_A_1139_367#_c_1094_n 0.00368563f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_157 VPB N_A_1139_367#_c_1095_n 0.00743874f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_158 VPB N_A_1139_367#_c_1096_n 0.0369431f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_159 N_D_N_M1015_g N_C_N_M1028_g 0.0272262f $X=0.525 $Y=0.675 $X2=0 $Y2=0
cc_160 N_D_N_M1032_g N_C_N_M1010_g 0.0272262f $X=0.525 $Y=2.465 $X2=0 $Y2=0
cc_161 N_D_N_c_162_n N_C_N_c_185_n 0.0272262f $X=0.525 $Y=1.46 $X2=0 $Y2=0
cc_162 N_D_N_M1015_g N_A_37_51#_c_222_n 0.0176373f $X=0.525 $Y=0.675 $X2=0 $Y2=0
cc_163 N_D_N_c_161_n N_A_37_51#_c_222_n 0.0056539f $X=0.31 $Y=1.46 $X2=0 $Y2=0
cc_164 N_D_N_c_162_n N_A_37_51#_c_222_n 0.00134357f $X=0.525 $Y=1.46 $X2=0 $Y2=0
cc_165 N_D_N_c_161_n N_A_37_51#_c_223_n 0.0205005f $X=0.31 $Y=1.46 $X2=0 $Y2=0
cc_166 N_D_N_c_162_n N_A_37_51#_c_223_n 0.00638328f $X=0.525 $Y=1.46 $X2=0 $Y2=0
cc_167 N_D_N_M1015_g N_A_37_51#_c_224_n 0.00976034f $X=0.525 $Y=0.675 $X2=0
+ $Y2=0
cc_168 N_D_N_c_161_n N_A_37_51#_c_224_n 0.0293932f $X=0.31 $Y=1.46 $X2=0 $Y2=0
cc_169 N_D_N_M1032_g N_A_37_51#_c_236_n 0.023729f $X=0.525 $Y=2.465 $X2=0 $Y2=0
cc_170 N_D_N_c_161_n N_A_37_51#_c_236_n 0.0257749f $X=0.31 $Y=1.46 $X2=0 $Y2=0
cc_171 N_D_N_c_162_n N_A_37_51#_c_236_n 0.0015691f $X=0.525 $Y=1.46 $X2=0 $Y2=0
cc_172 N_D_N_M1032_g N_VPWR_c_685_n 0.011439f $X=0.525 $Y=2.465 $X2=0 $Y2=0
cc_173 N_D_N_M1032_g N_VPWR_c_688_n 0.00486043f $X=0.525 $Y=2.465 $X2=0 $Y2=0
cc_174 N_D_N_M1032_g N_VPWR_c_684_n 0.00553852f $X=0.525 $Y=2.465 $X2=0 $Y2=0
cc_175 N_D_N_M1015_g N_VGND_c_1158_n 0.0118508f $X=0.525 $Y=0.675 $X2=0 $Y2=0
cc_176 N_D_N_M1015_g N_VGND_c_1173_n 0.00469214f $X=0.525 $Y=0.675 $X2=0 $Y2=0
cc_177 N_D_N_M1015_g N_VGND_c_1188_n 0.0091547f $X=0.525 $Y=0.675 $X2=0 $Y2=0
cc_178 N_C_N_M1028_g N_A_37_51#_c_222_n 0.00139605f $X=0.955 $Y=0.675 $X2=0
+ $Y2=0
cc_179 N_C_N_M1028_g N_A_37_51#_c_224_n 0.00648073f $X=0.955 $Y=0.675 $X2=0
+ $Y2=0
cc_180 N_C_N_c_186_n N_A_37_51#_c_224_n 0.0309802f $X=1.09 $Y=1.51 $X2=0 $Y2=0
cc_181 N_C_N_M1010_g N_A_37_51#_c_234_n 0.0174707f $X=0.955 $Y=2.465 $X2=0 $Y2=0
cc_182 N_C_N_c_186_n N_A_37_51#_c_234_n 2.50215e-19 $X=1.09 $Y=1.51 $X2=0 $Y2=0
cc_183 N_C_N_c_185_n N_A_37_51#_c_227_n 0.00372429f $X=1.09 $Y=1.51 $X2=0 $Y2=0
cc_184 N_C_N_M1010_g N_A_206_51#_c_369_n 0.00281638f $X=0.955 $Y=2.465 $X2=0
+ $Y2=0
cc_185 N_C_N_c_185_n N_A_206_51#_c_369_n 0.00117836f $X=1.09 $Y=1.51 $X2=0 $Y2=0
cc_186 N_C_N_c_186_n N_A_206_51#_c_369_n 0.02024f $X=1.09 $Y=1.51 $X2=0 $Y2=0
cc_187 N_C_N_M1028_g N_A_206_51#_c_360_n 0.00293027f $X=0.955 $Y=0.675 $X2=0
+ $Y2=0
cc_188 N_C_N_M1010_g N_A_206_51#_c_360_n 0.00211812f $X=0.955 $Y=2.465 $X2=0
+ $Y2=0
cc_189 N_C_N_c_185_n N_A_206_51#_c_360_n 0.00145825f $X=1.09 $Y=1.51 $X2=0 $Y2=0
cc_190 N_C_N_c_186_n N_A_206_51#_c_360_n 0.0327007f $X=1.09 $Y=1.51 $X2=0 $Y2=0
cc_191 N_C_N_M1028_g N_A_206_51#_c_363_n 0.00196337f $X=0.955 $Y=0.675 $X2=0
+ $Y2=0
cc_192 N_C_N_c_185_n N_A_206_51#_c_363_n 0.00127412f $X=1.09 $Y=1.51 $X2=0 $Y2=0
cc_193 N_C_N_c_186_n N_A_206_51#_c_363_n 0.0162575f $X=1.09 $Y=1.51 $X2=0 $Y2=0
cc_194 N_C_N_M1010_g N_VPWR_c_685_n 0.0253312f $X=0.955 $Y=2.465 $X2=0 $Y2=0
cc_195 N_C_N_M1010_g N_VPWR_c_689_n 0.00486043f $X=0.955 $Y=2.465 $X2=0 $Y2=0
cc_196 N_C_N_M1010_g N_VPWR_c_684_n 0.00603991f $X=0.955 $Y=2.465 $X2=0 $Y2=0
cc_197 N_C_N_M1010_g N_A_347_349#_c_791_n 0.00946396f $X=0.955 $Y=2.465 $X2=0
+ $Y2=0
cc_198 N_C_N_M1028_g N_VGND_c_1158_n 0.0114818f $X=0.955 $Y=0.675 $X2=0 $Y2=0
cc_199 N_C_N_M1028_g N_VGND_c_1159_n 0.00225739f $X=0.955 $Y=0.675 $X2=0 $Y2=0
cc_200 N_C_N_M1028_g N_VGND_c_1174_n 0.00469214f $X=0.955 $Y=0.675 $X2=0 $Y2=0
cc_201 N_C_N_M1028_g N_VGND_c_1188_n 0.00945295f $X=0.955 $Y=0.675 $X2=0 $Y2=0
cc_202 N_A_37_51#_c_234_n N_A_206_51#_M1010_d 0.00708486f $X=1.82 $Y=2.395 $X2=0
+ $Y2=0
cc_203 N_A_37_51#_M1030_g N_A_206_51#_M1001_g 0.0253942f $X=3.365 $Y=2.375 $X2=0
+ $Y2=0
cc_204 N_A_37_51#_M1029_g N_A_206_51#_M1000_g 0.0326128f $X=3.435 $Y=0.655 $X2=0
+ $Y2=0
cc_205 N_A_37_51#_M1005_g N_A_206_51#_c_369_n 0.00109524f $X=2.075 $Y=2.375
+ $X2=0 $Y2=0
cc_206 N_A_37_51#_c_234_n N_A_206_51#_c_369_n 0.0443538f $X=1.82 $Y=2.395 $X2=0
+ $Y2=0
cc_207 N_A_37_51#_c_235_n N_A_206_51#_c_369_n 0.016518f $X=1.922 $Y=2.31 $X2=0
+ $Y2=0
cc_208 N_A_37_51#_M1002_g N_A_206_51#_c_359_n 0.00502883f $X=1.975 $Y=0.655
+ $X2=0 $Y2=0
cc_209 N_A_37_51#_M1002_g N_A_206_51#_c_360_n 0.00247517f $X=1.975 $Y=0.655
+ $X2=0 $Y2=0
cc_210 N_A_37_51#_M1005_g N_A_206_51#_c_360_n 0.00160339f $X=2.075 $Y=2.375
+ $X2=0 $Y2=0
cc_211 N_A_37_51#_c_222_n N_A_206_51#_c_360_n 6.70846e-19 $X=0.645 $Y=1.11 $X2=0
+ $Y2=0
cc_212 N_A_37_51#_c_224_n N_A_206_51#_c_360_n 0.00818415f $X=0.735 $Y=1.93 $X2=0
+ $Y2=0
cc_213 N_A_37_51#_c_225_n N_A_206_51#_c_360_n 0.0135453f $X=1.922 $Y=1.515 $X2=0
+ $Y2=0
cc_214 N_A_37_51#_c_235_n N_A_206_51#_c_360_n 0.0293902f $X=1.922 $Y=2.31 $X2=0
+ $Y2=0
cc_215 N_A_37_51#_c_227_n N_A_206_51#_c_360_n 0.00477586f $X=3.435 $Y=1.42 $X2=0
+ $Y2=0
cc_216 N_A_37_51#_M1002_g N_A_206_51#_c_361_n 0.0163446f $X=1.975 $Y=0.655 $X2=0
+ $Y2=0
cc_217 N_A_37_51#_M1009_g N_A_206_51#_c_361_n 0.0113322f $X=2.405 $Y=0.655 $X2=0
+ $Y2=0
cc_218 N_A_37_51#_M1026_g N_A_206_51#_c_361_n 0.0113326f $X=3.005 $Y=0.655 $X2=0
+ $Y2=0
cc_219 N_A_37_51#_M1029_g N_A_206_51#_c_361_n 0.0108241f $X=3.435 $Y=0.655 $X2=0
+ $Y2=0
cc_220 N_A_37_51#_c_225_n N_A_206_51#_c_361_n 0.0159146f $X=1.922 $Y=1.515 $X2=0
+ $Y2=0
cc_221 N_A_37_51#_c_226_n N_A_206_51#_c_361_n 0.104851f $X=3.345 $Y=1.42 $X2=0
+ $Y2=0
cc_222 N_A_37_51#_c_227_n N_A_206_51#_c_361_n 0.0150162f $X=3.435 $Y=1.42 $X2=0
+ $Y2=0
cc_223 N_A_37_51#_M1029_g N_A_206_51#_c_362_n 0.00181339f $X=3.435 $Y=0.655
+ $X2=0 $Y2=0
cc_224 N_A_37_51#_c_226_n N_A_206_51#_c_362_n 0.0127007f $X=3.345 $Y=1.42 $X2=0
+ $Y2=0
cc_225 N_A_37_51#_c_227_n N_A_206_51#_c_362_n 8.37465e-19 $X=3.435 $Y=1.42 $X2=0
+ $Y2=0
cc_226 N_A_37_51#_M1002_g N_A_206_51#_c_363_n 3.23195e-19 $X=1.975 $Y=0.655
+ $X2=0 $Y2=0
cc_227 N_A_37_51#_c_222_n N_A_206_51#_c_363_n 0.00555193f $X=0.645 $Y=1.11 $X2=0
+ $Y2=0
cc_228 N_A_37_51#_c_226_n N_A_206_51#_c_364_n 2.20823e-19 $X=3.345 $Y=1.42 $X2=0
+ $Y2=0
cc_229 N_A_37_51#_c_227_n N_A_206_51#_c_364_n 0.0237318f $X=3.435 $Y=1.42 $X2=0
+ $Y2=0
cc_230 N_A_37_51#_c_224_n N_VPWR_M1032_d 6.80144e-19 $X=0.735 $Y=1.93 $X2=-0.19
+ $Y2=-0.245
cc_231 N_A_37_51#_c_236_n N_VPWR_M1032_d 0.00276932f $X=0.825 $Y=2.205 $X2=-0.19
+ $Y2=-0.245
cc_232 N_A_37_51#_c_236_n N_VPWR_c_685_n 0.0179755f $X=0.825 $Y=2.205 $X2=0
+ $Y2=0
cc_233 N_A_37_51#_c_232_n N_VPWR_c_688_n 0.0176409f $X=0.31 $Y=2.49 $X2=0 $Y2=0
cc_234 N_A_37_51#_M1005_g N_VPWR_c_689_n 0.00303788f $X=2.075 $Y=2.375 $X2=0
+ $Y2=0
cc_235 N_A_37_51#_M1012_g N_VPWR_c_689_n 0.00302473f $X=2.505 $Y=2.375 $X2=0
+ $Y2=0
cc_236 N_A_37_51#_M1019_g N_VPWR_c_689_n 0.00302473f $X=2.935 $Y=2.375 $X2=0
+ $Y2=0
cc_237 N_A_37_51#_M1030_g N_VPWR_c_689_n 0.00302501f $X=3.365 $Y=2.375 $X2=0
+ $Y2=0
cc_238 N_A_37_51#_M1032_s N_VPWR_c_684_n 0.00245679f $X=0.185 $Y=1.835 $X2=0
+ $Y2=0
cc_239 N_A_37_51#_M1005_g N_VPWR_c_684_n 0.00483749f $X=2.075 $Y=2.375 $X2=0
+ $Y2=0
cc_240 N_A_37_51#_M1012_g N_VPWR_c_684_n 0.0043467f $X=2.505 $Y=2.375 $X2=0
+ $Y2=0
cc_241 N_A_37_51#_M1019_g N_VPWR_c_684_n 0.0043467f $X=2.935 $Y=2.375 $X2=0
+ $Y2=0
cc_242 N_A_37_51#_M1030_g N_VPWR_c_684_n 0.00435646f $X=3.365 $Y=2.375 $X2=0
+ $Y2=0
cc_243 N_A_37_51#_c_232_n N_VPWR_c_684_n 0.00999551f $X=0.31 $Y=2.49 $X2=0 $Y2=0
cc_244 N_A_37_51#_c_234_n N_VPWR_c_684_n 0.0267738f $X=1.82 $Y=2.395 $X2=0 $Y2=0
cc_245 N_A_37_51#_c_236_n N_VPWR_c_684_n 0.0066936f $X=0.825 $Y=2.205 $X2=0
+ $Y2=0
cc_246 N_A_37_51#_c_234_n N_A_347_349#_M1005_d 0.00620037f $X=1.82 $Y=2.395
+ $X2=-0.19 $Y2=-0.245
cc_247 N_A_37_51#_c_235_n N_A_347_349#_M1005_d 0.0109777f $X=1.922 $Y=2.31
+ $X2=-0.19 $Y2=-0.245
cc_248 N_A_37_51#_M1005_g N_A_347_349#_c_789_n 0.0108332f $X=2.075 $Y=2.375
+ $X2=0 $Y2=0
cc_249 N_A_37_51#_M1012_g N_A_347_349#_c_789_n 0.0102372f $X=2.505 $Y=2.375
+ $X2=0 $Y2=0
cc_250 N_A_37_51#_M1005_g N_A_347_349#_c_799_n 6.35714e-19 $X=2.075 $Y=2.375
+ $X2=0 $Y2=0
cc_251 N_A_37_51#_M1012_g N_A_347_349#_c_799_n 0.0105167f $X=2.505 $Y=2.375
+ $X2=0 $Y2=0
cc_252 N_A_37_51#_M1019_g N_A_347_349#_c_799_n 0.0106252f $X=2.935 $Y=2.375
+ $X2=0 $Y2=0
cc_253 N_A_37_51#_M1030_g N_A_347_349#_c_799_n 6.43964e-19 $X=3.365 $Y=2.375
+ $X2=0 $Y2=0
cc_254 N_A_37_51#_M1019_g N_A_347_349#_c_790_n 0.0101906f $X=2.935 $Y=2.375
+ $X2=0 $Y2=0
cc_255 N_A_37_51#_M1030_g N_A_347_349#_c_790_n 0.0125396f $X=3.365 $Y=2.375
+ $X2=0 $Y2=0
cc_256 N_A_37_51#_M1005_g N_A_347_349#_c_791_n 0.00690072f $X=2.075 $Y=2.375
+ $X2=0 $Y2=0
cc_257 N_A_37_51#_M1012_g N_A_347_349#_c_791_n 5.41136e-19 $X=2.505 $Y=2.375
+ $X2=0 $Y2=0
cc_258 N_A_37_51#_c_234_n N_A_347_349#_c_791_n 0.0218699f $X=1.82 $Y=2.395 $X2=0
+ $Y2=0
cc_259 N_A_37_51#_M1012_g N_A_347_349#_c_792_n 0.00137179f $X=2.505 $Y=2.375
+ $X2=0 $Y2=0
cc_260 N_A_37_51#_M1019_g N_A_347_349#_c_792_n 0.00137179f $X=2.935 $Y=2.375
+ $X2=0 $Y2=0
cc_261 N_A_37_51#_M1002_g N_Y_c_868_n 0.00444742f $X=1.975 $Y=0.655 $X2=0 $Y2=0
cc_262 N_A_37_51#_M1009_g N_Y_c_868_n 0.00647128f $X=2.405 $Y=0.655 $X2=0 $Y2=0
cc_263 N_A_37_51#_M1026_g N_Y_c_868_n 8.17275e-19 $X=3.005 $Y=0.655 $X2=0 $Y2=0
cc_264 N_A_37_51#_M1009_g N_Y_c_871_n 0.00888334f $X=2.405 $Y=0.655 $X2=0 $Y2=0
cc_265 N_A_37_51#_M1026_g N_Y_c_871_n 0.00941278f $X=3.005 $Y=0.655 $X2=0 $Y2=0
cc_266 N_A_37_51#_M1002_g N_Y_c_873_n 0.00251291f $X=1.975 $Y=0.655 $X2=0 $Y2=0
cc_267 N_A_37_51#_M1009_g N_Y_c_873_n 0.00101901f $X=2.405 $Y=0.655 $X2=0 $Y2=0
cc_268 N_A_37_51#_M1012_g N_Y_c_862_n 0.0128162f $X=2.505 $Y=2.375 $X2=0 $Y2=0
cc_269 N_A_37_51#_M1019_g N_Y_c_862_n 0.0129249f $X=2.935 $Y=2.375 $X2=0 $Y2=0
cc_270 N_A_37_51#_c_226_n N_Y_c_862_n 0.0469272f $X=3.345 $Y=1.42 $X2=0 $Y2=0
cc_271 N_A_37_51#_c_227_n N_Y_c_862_n 0.00243542f $X=3.435 $Y=1.42 $X2=0 $Y2=0
cc_272 N_A_37_51#_M1005_g N_Y_c_863_n 4.90985e-19 $X=2.075 $Y=2.375 $X2=0 $Y2=0
cc_273 N_A_37_51#_c_235_n N_Y_c_863_n 0.00870837f $X=1.922 $Y=2.31 $X2=0 $Y2=0
cc_274 N_A_37_51#_c_226_n N_Y_c_863_n 0.0153881f $X=3.345 $Y=1.42 $X2=0 $Y2=0
cc_275 N_A_37_51#_c_227_n N_Y_c_863_n 0.00296179f $X=3.435 $Y=1.42 $X2=0 $Y2=0
cc_276 N_A_37_51#_M1009_g N_Y_c_883_n 8.08771e-19 $X=2.405 $Y=0.655 $X2=0 $Y2=0
cc_277 N_A_37_51#_M1026_g N_Y_c_883_n 0.00620552f $X=3.005 $Y=0.655 $X2=0 $Y2=0
cc_278 N_A_37_51#_M1029_g N_Y_c_883_n 0.00592294f $X=3.435 $Y=0.655 $X2=0 $Y2=0
cc_279 N_A_37_51#_M1030_g N_Y_c_864_n 0.0139648f $X=3.365 $Y=2.375 $X2=0 $Y2=0
cc_280 N_A_37_51#_c_226_n N_Y_c_864_n 0.01563f $X=3.345 $Y=1.42 $X2=0 $Y2=0
cc_281 N_A_37_51#_c_227_n N_Y_c_864_n 0.00200474f $X=3.435 $Y=1.42 $X2=0 $Y2=0
cc_282 N_A_37_51#_M1029_g N_Y_c_889_n 0.0089043f $X=3.435 $Y=0.655 $X2=0 $Y2=0
cc_283 N_A_37_51#_M1026_g N_Y_c_890_n 7.15068e-19 $X=3.005 $Y=0.655 $X2=0 $Y2=0
cc_284 N_A_37_51#_M1029_g N_Y_c_890_n 7.15068e-19 $X=3.435 $Y=0.655 $X2=0 $Y2=0
cc_285 N_A_37_51#_c_226_n N_Y_c_865_n 0.0186283f $X=3.345 $Y=1.42 $X2=0 $Y2=0
cc_286 N_A_37_51#_c_227_n N_Y_c_865_n 0.00283411f $X=3.435 $Y=1.42 $X2=0 $Y2=0
cc_287 N_A_37_51#_c_222_n N_VGND_M1015_d 0.0019798f $X=0.645 $Y=1.11 $X2=-0.19
+ $Y2=-0.245
cc_288 N_A_37_51#_c_222_n N_VGND_c_1158_n 0.0167529f $X=0.645 $Y=1.11 $X2=0
+ $Y2=0
cc_289 N_A_37_51#_M1002_g N_VGND_c_1159_n 0.0158707f $X=1.975 $Y=0.655 $X2=0
+ $Y2=0
cc_290 N_A_37_51#_M1009_g N_VGND_c_1160_n 0.0047103f $X=2.405 $Y=0.655 $X2=0
+ $Y2=0
cc_291 N_A_37_51#_M1026_g N_VGND_c_1160_n 0.00574924f $X=3.005 $Y=0.655 $X2=0
+ $Y2=0
cc_292 N_A_37_51#_M1026_g N_VGND_c_1161_n 0.00417814f $X=3.005 $Y=0.655 $X2=0
+ $Y2=0
cc_293 N_A_37_51#_M1029_g N_VGND_c_1161_n 0.00417814f $X=3.435 $Y=0.655 $X2=0
+ $Y2=0
cc_294 N_A_37_51#_M1029_g N_VGND_c_1162_n 0.00436654f $X=3.435 $Y=0.655 $X2=0
+ $Y2=0
cc_295 N_A_37_51#_c_221_n N_VGND_c_1173_n 0.0174563f $X=0.31 $Y=0.42 $X2=0 $Y2=0
cc_296 N_A_37_51#_M1002_g N_VGND_c_1175_n 0.0054895f $X=1.975 $Y=0.655 $X2=0
+ $Y2=0
cc_297 N_A_37_51#_M1009_g N_VGND_c_1175_n 0.00413124f $X=2.405 $Y=0.655 $X2=0
+ $Y2=0
cc_298 N_A_37_51#_M1002_g N_VGND_c_1188_n 0.0112727f $X=1.975 $Y=0.655 $X2=0
+ $Y2=0
cc_299 N_A_37_51#_M1009_g N_VGND_c_1188_n 0.00612913f $X=2.405 $Y=0.655 $X2=0
+ $Y2=0
cc_300 N_A_37_51#_M1026_g N_VGND_c_1188_n 0.00619988f $X=3.005 $Y=0.655 $X2=0
+ $Y2=0
cc_301 N_A_37_51#_M1029_g N_VGND_c_1188_n 0.00593637f $X=3.435 $Y=0.655 $X2=0
+ $Y2=0
cc_302 N_A_37_51#_c_221_n N_VGND_c_1188_n 0.00963638f $X=0.31 $Y=0.42 $X2=0
+ $Y2=0
cc_303 N_A_206_51#_M1034_g N_B_M1006_g 0.00592444f $X=5.225 $Y=0.655 $X2=0 $Y2=0
cc_304 N_A_206_51#_M1027_g N_B_c_509_n 5.4976e-19 $X=5.085 $Y=2.375 $X2=0 $Y2=0
cc_305 N_A_206_51#_M1027_g N_B_c_510_n 2.25796e-19 $X=5.085 $Y=2.375 $X2=0 $Y2=0
cc_306 N_A_206_51#_c_364_n N_B_c_510_n 0.00629347f $X=5.225 $Y=1.42 $X2=0 $Y2=0
cc_307 N_A_206_51#_M1001_g N_VPWR_c_689_n 0.00466675f $X=3.795 $Y=2.375 $X2=0
+ $Y2=0
cc_308 N_A_206_51#_M1007_g N_VPWR_c_689_n 0.00302473f $X=4.225 $Y=2.375 $X2=0
+ $Y2=0
cc_309 N_A_206_51#_M1013_g N_VPWR_c_689_n 0.00302473f $X=4.655 $Y=2.375 $X2=0
+ $Y2=0
cc_310 N_A_206_51#_M1027_g N_VPWR_c_689_n 0.00302473f $X=5.085 $Y=2.375 $X2=0
+ $Y2=0
cc_311 N_A_206_51#_M1010_d N_VPWR_c_684_n 0.00395695f $X=1.03 $Y=1.835 $X2=0
+ $Y2=0
cc_312 N_A_206_51#_M1001_g N_VPWR_c_684_n 0.00898886f $X=3.795 $Y=2.375 $X2=0
+ $Y2=0
cc_313 N_A_206_51#_M1007_g N_VPWR_c_684_n 0.0043467f $X=4.225 $Y=2.375 $X2=0
+ $Y2=0
cc_314 N_A_206_51#_M1013_g N_VPWR_c_684_n 0.0043467f $X=4.655 $Y=2.375 $X2=0
+ $Y2=0
cc_315 N_A_206_51#_M1027_g N_VPWR_c_684_n 0.00484658f $X=5.085 $Y=2.375 $X2=0
+ $Y2=0
cc_316 N_A_206_51#_M1001_g N_A_347_349#_c_790_n 5.72e-19 $X=3.795 $Y=2.375 $X2=0
+ $Y2=0
cc_317 N_A_206_51#_M1001_g N_A_347_349#_c_811_n 0.0122595f $X=3.795 $Y=2.375
+ $X2=0 $Y2=0
cc_318 N_A_206_51#_M1007_g N_A_347_349#_c_811_n 0.0122129f $X=4.225 $Y=2.375
+ $X2=0 $Y2=0
cc_319 N_A_206_51#_M1013_g N_A_347_349#_c_813_n 0.0122595f $X=4.655 $Y=2.375
+ $X2=0 $Y2=0
cc_320 N_A_206_51#_M1027_g N_A_347_349#_c_813_n 0.0122595f $X=5.085 $Y=2.375
+ $X2=0 $Y2=0
cc_321 N_A_206_51#_c_364_n N_A_347_349#_c_793_n 2.85505e-19 $X=5.225 $Y=1.42
+ $X2=0 $Y2=0
cc_322 N_A_206_51#_c_361_n N_Y_M1002_s 0.00176461f $X=3.72 $Y=1.08 $X2=-0.19
+ $Y2=-0.245
cc_323 N_A_206_51#_c_361_n N_Y_M1026_s 0.00176461f $X=3.72 $Y=1.08 $X2=0 $Y2=0
cc_324 N_A_206_51#_c_361_n N_Y_c_871_n 0.0406043f $X=3.72 $Y=1.08 $X2=0 $Y2=0
cc_325 N_A_206_51#_c_361_n N_Y_c_873_n 0.0177368f $X=3.72 $Y=1.08 $X2=0 $Y2=0
cc_326 N_A_206_51#_M1000_g N_Y_c_883_n 3.68986e-19 $X=3.935 $Y=0.655 $X2=0 $Y2=0
cc_327 N_A_206_51#_M1001_g N_Y_c_864_n 0.0108274f $X=3.795 $Y=2.375 $X2=0 $Y2=0
cc_328 N_A_206_51#_M1007_g N_Y_c_864_n 0.010883f $X=4.225 $Y=2.375 $X2=0 $Y2=0
cc_329 N_A_206_51#_M1013_g N_Y_c_864_n 0.010883f $X=4.655 $Y=2.375 $X2=0 $Y2=0
cc_330 N_A_206_51#_M1027_g N_Y_c_864_n 0.0136603f $X=5.085 $Y=2.375 $X2=0 $Y2=0
cc_331 N_A_206_51#_c_361_n N_Y_c_864_n 0.00730632f $X=3.72 $Y=1.08 $X2=0 $Y2=0
cc_332 N_A_206_51#_c_362_n N_Y_c_864_n 0.0127093f $X=3.805 $Y=1.335 $X2=0 $Y2=0
cc_333 N_A_206_51#_c_440_p N_Y_c_864_n 0.0837539f $X=4.905 $Y=1.42 $X2=0 $Y2=0
cc_334 N_A_206_51#_c_364_n N_Y_c_864_n 0.0115391f $X=5.225 $Y=1.42 $X2=0 $Y2=0
cc_335 N_A_206_51#_M1000_g N_Y_c_889_n 0.0120778f $X=3.935 $Y=0.655 $X2=0 $Y2=0
cc_336 N_A_206_51#_c_361_n N_Y_c_889_n 0.0283574f $X=3.72 $Y=1.08 $X2=0 $Y2=0
cc_337 N_A_206_51#_c_440_p N_Y_c_889_n 0.00393123f $X=4.905 $Y=1.42 $X2=0 $Y2=0
cc_338 N_A_206_51#_c_364_n N_Y_c_889_n 4.62646e-19 $X=5.225 $Y=1.42 $X2=0 $Y2=0
cc_339 N_A_206_51#_M1004_g N_Y_c_851_n 0.0130886f $X=4.365 $Y=0.655 $X2=0 $Y2=0
cc_340 N_A_206_51#_M1022_g N_Y_c_851_n 0.013286f $X=4.795 $Y=0.655 $X2=0 $Y2=0
cc_341 N_A_206_51#_c_440_p N_Y_c_851_n 0.0469271f $X=4.905 $Y=1.42 $X2=0 $Y2=0
cc_342 N_A_206_51#_c_364_n N_Y_c_851_n 0.00289453f $X=5.225 $Y=1.42 $X2=0 $Y2=0
cc_343 N_A_206_51#_M1000_g N_Y_c_852_n 7.28841e-19 $X=3.935 $Y=0.655 $X2=0 $Y2=0
cc_344 N_A_206_51#_c_361_n N_Y_c_852_n 0.011362f $X=3.72 $Y=1.08 $X2=0 $Y2=0
cc_345 N_A_206_51#_c_440_p N_Y_c_852_n 0.0149829f $X=4.905 $Y=1.42 $X2=0 $Y2=0
cc_346 N_A_206_51#_c_364_n N_Y_c_852_n 0.00299787f $X=5.225 $Y=1.42 $X2=0 $Y2=0
cc_347 N_A_206_51#_M1034_g N_Y_c_854_n 0.0160086f $X=5.225 $Y=0.655 $X2=0 $Y2=0
cc_348 N_A_206_51#_c_440_p N_Y_c_854_n 0.0125528f $X=4.905 $Y=1.42 $X2=0 $Y2=0
cc_349 N_A_206_51#_c_364_n N_Y_c_854_n 0.00299787f $X=5.225 $Y=1.42 $X2=0 $Y2=0
cc_350 N_A_206_51#_c_361_n N_Y_c_890_n 0.0169862f $X=3.72 $Y=1.08 $X2=0 $Y2=0
cc_351 N_A_206_51#_M1022_g Y 4.00458e-19 $X=4.795 $Y=0.655 $X2=0 $Y2=0
cc_352 N_A_206_51#_M1027_g Y 0.00385189f $X=5.085 $Y=2.375 $X2=0 $Y2=0
cc_353 N_A_206_51#_M1034_g Y 0.00290061f $X=5.225 $Y=0.655 $X2=0 $Y2=0
cc_354 N_A_206_51#_c_440_p Y 0.0136681f $X=4.905 $Y=1.42 $X2=0 $Y2=0
cc_355 N_A_206_51#_c_364_n Y 0.0172619f $X=5.225 $Y=1.42 $X2=0 $Y2=0
cc_356 N_A_206_51#_M1001_g N_A_774_349#_c_1029_n 0.00567926f $X=3.795 $Y=2.375
+ $X2=0 $Y2=0
cc_357 N_A_206_51#_M1007_g N_A_774_349#_c_1029_n 0.00691995f $X=4.225 $Y=2.375
+ $X2=0 $Y2=0
cc_358 N_A_206_51#_M1013_g N_A_774_349#_c_1029_n 5.36673e-19 $X=4.655 $Y=2.375
+ $X2=0 $Y2=0
cc_359 N_A_206_51#_M1007_g N_A_774_349#_c_1025_n 0.0102372f $X=4.225 $Y=2.375
+ $X2=0 $Y2=0
cc_360 N_A_206_51#_M1013_g N_A_774_349#_c_1025_n 0.0102372f $X=4.655 $Y=2.375
+ $X2=0 $Y2=0
cc_361 N_A_206_51#_M1001_g N_A_774_349#_c_1026_n 0.00268726f $X=3.795 $Y=2.375
+ $X2=0 $Y2=0
cc_362 N_A_206_51#_M1007_g N_A_774_349#_c_1026_n 0.00136552f $X=4.225 $Y=2.375
+ $X2=0 $Y2=0
cc_363 N_A_206_51#_M1007_g N_A_774_349#_c_1036_n 4.7782e-19 $X=4.225 $Y=2.375
+ $X2=0 $Y2=0
cc_364 N_A_206_51#_M1013_g N_A_774_349#_c_1036_n 0.0065713f $X=4.655 $Y=2.375
+ $X2=0 $Y2=0
cc_365 N_A_206_51#_M1027_g N_A_774_349#_c_1036_n 0.0112802f $X=5.085 $Y=2.375
+ $X2=0 $Y2=0
cc_366 N_A_206_51#_M1027_g N_A_774_349#_c_1027_n 0.0130642f $X=5.085 $Y=2.375
+ $X2=0 $Y2=0
cc_367 N_A_206_51#_M1013_g N_A_774_349#_c_1028_n 0.0017155f $X=4.655 $Y=2.375
+ $X2=0 $Y2=0
cc_368 N_A_206_51#_M1027_g N_A_774_349#_c_1028_n 0.00141072f $X=5.085 $Y=2.375
+ $X2=0 $Y2=0
cc_369 N_A_206_51#_c_361_n N_VGND_M1002_d 0.00262118f $X=3.72 $Y=1.08 $X2=0
+ $Y2=0
cc_370 N_A_206_51#_c_363_n N_VGND_M1002_d 0.00106962f $X=1.635 $Y=1.085 $X2=0
+ $Y2=0
cc_371 N_A_206_51#_c_361_n N_VGND_M1009_d 0.00397399f $X=3.72 $Y=1.08 $X2=0
+ $Y2=0
cc_372 N_A_206_51#_c_361_n N_VGND_M1029_d 0.00253298f $X=3.72 $Y=1.08 $X2=0
+ $Y2=0
cc_373 N_A_206_51#_c_359_n N_VGND_c_1159_n 0.0423573f $X=1.17 $Y=0.42 $X2=0
+ $Y2=0
cc_374 N_A_206_51#_c_363_n N_VGND_c_1159_n 0.0248327f $X=1.635 $Y=1.085 $X2=0
+ $Y2=0
cc_375 N_A_206_51#_M1000_g N_VGND_c_1162_n 0.00664552f $X=3.935 $Y=0.655 $X2=0
+ $Y2=0
cc_376 N_A_206_51#_M1004_g N_VGND_c_1162_n 5.14991e-19 $X=4.365 $Y=0.655 $X2=0
+ $Y2=0
cc_377 N_A_206_51#_M1000_g N_VGND_c_1163_n 6.48667e-19 $X=3.935 $Y=0.655 $X2=0
+ $Y2=0
cc_378 N_A_206_51#_M1004_g N_VGND_c_1163_n 0.0100562f $X=4.365 $Y=0.655 $X2=0
+ $Y2=0
cc_379 N_A_206_51#_M1022_g N_VGND_c_1163_n 0.010076f $X=4.795 $Y=0.655 $X2=0
+ $Y2=0
cc_380 N_A_206_51#_M1034_g N_VGND_c_1163_n 6.11179e-19 $X=5.225 $Y=0.655 $X2=0
+ $Y2=0
cc_381 N_A_206_51#_M1022_g N_VGND_c_1164_n 6.2389e-19 $X=4.795 $Y=0.655 $X2=0
+ $Y2=0
cc_382 N_A_206_51#_M1034_g N_VGND_c_1164_n 0.0110426f $X=5.225 $Y=0.655 $X2=0
+ $Y2=0
cc_383 N_A_206_51#_c_359_n N_VGND_c_1174_n 0.0178111f $X=1.17 $Y=0.42 $X2=0
+ $Y2=0
cc_384 N_A_206_51#_M1000_g N_VGND_c_1176_n 0.00355956f $X=3.935 $Y=0.655 $X2=0
+ $Y2=0
cc_385 N_A_206_51#_M1004_g N_VGND_c_1176_n 0.00486043f $X=4.365 $Y=0.655 $X2=0
+ $Y2=0
cc_386 N_A_206_51#_M1022_g N_VGND_c_1177_n 0.00486043f $X=4.795 $Y=0.655 $X2=0
+ $Y2=0
cc_387 N_A_206_51#_M1034_g N_VGND_c_1177_n 0.00486043f $X=5.225 $Y=0.655 $X2=0
+ $Y2=0
cc_388 N_A_206_51#_M1000_g N_VGND_c_1188_n 0.00415754f $X=3.935 $Y=0.655 $X2=0
+ $Y2=0
cc_389 N_A_206_51#_M1004_g N_VGND_c_1188_n 0.00824727f $X=4.365 $Y=0.655 $X2=0
+ $Y2=0
cc_390 N_A_206_51#_M1022_g N_VGND_c_1188_n 0.00824727f $X=4.795 $Y=0.655 $X2=0
+ $Y2=0
cc_391 N_A_206_51#_M1034_g N_VGND_c_1188_n 0.00824727f $X=5.225 $Y=0.655 $X2=0
+ $Y2=0
cc_392 N_A_206_51#_c_359_n N_VGND_c_1188_n 0.0100304f $X=1.17 $Y=0.42 $X2=0
+ $Y2=0
cc_393 N_B_M1035_g N_A_M1016_g 0.0210758f $X=7.33 $Y=0.655 $X2=0 $Y2=0
cc_394 N_B_c_510_n N_A_M1016_g 0.0240911f $X=7.33 $Y=1.44 $X2=0 $Y2=0
cc_395 N_B_M1033_g A 5.33717e-19 $X=7.325 $Y=2.465 $X2=0 $Y2=0
cc_396 N_B_c_508_n A 0.00751696f $X=7.31 $Y=1.44 $X2=0 $Y2=0
cc_397 N_B_c_510_n A 6.38564e-19 $X=7.33 $Y=1.44 $X2=0 $Y2=0
cc_398 N_B_M1033_g N_A_c_616_n 0.0211479f $X=7.325 $Y=2.465 $X2=0 $Y2=0
cc_399 N_B_c_508_n N_A_c_616_n 7.91318e-19 $X=7.31 $Y=1.44 $X2=0 $Y2=0
cc_400 N_B_M1033_g N_VPWR_c_686_n 0.00130952f $X=7.325 $Y=2.465 $X2=0 $Y2=0
cc_401 N_B_M1008_g N_VPWR_c_689_n 0.00357842f $X=6.035 $Y=2.465 $X2=0 $Y2=0
cc_402 N_B_M1014_g N_VPWR_c_689_n 0.00357842f $X=6.465 $Y=2.465 $X2=0 $Y2=0
cc_403 N_B_M1021_g N_VPWR_c_689_n 0.00357842f $X=6.895 $Y=2.465 $X2=0 $Y2=0
cc_404 N_B_M1033_g N_VPWR_c_689_n 0.00547432f $X=7.325 $Y=2.465 $X2=0 $Y2=0
cc_405 N_B_M1008_g N_VPWR_c_684_n 0.00675085f $X=6.035 $Y=2.465 $X2=0 $Y2=0
cc_406 N_B_M1014_g N_VPWR_c_684_n 0.00535118f $X=6.465 $Y=2.465 $X2=0 $Y2=0
cc_407 N_B_M1021_g N_VPWR_c_684_n 0.00535118f $X=6.895 $Y=2.465 $X2=0 $Y2=0
cc_408 N_B_M1033_g N_VPWR_c_684_n 0.00991323f $X=7.325 $Y=2.465 $X2=0 $Y2=0
cc_409 N_B_M1006_g N_Y_c_853_n 0.0156688f $X=6.04 $Y=0.655 $X2=0 $Y2=0
cc_410 N_B_c_509_n N_Y_c_853_n 0.0274366f $X=5.95 $Y=1.44 $X2=0 $Y2=0
cc_411 N_B_c_510_n N_Y_c_853_n 0.00445594f $X=7.33 $Y=1.44 $X2=0 $Y2=0
cc_412 N_B_M1023_g N_Y_c_855_n 0.0135143f $X=6.47 $Y=0.655 $X2=0 $Y2=0
cc_413 N_B_M1024_g N_Y_c_855_n 0.0135143f $X=6.9 $Y=0.655 $X2=0 $Y2=0
cc_414 N_B_c_508_n N_Y_c_855_n 0.0447065f $X=7.31 $Y=1.44 $X2=0 $Y2=0
cc_415 N_B_c_510_n N_Y_c_855_n 0.00247028f $X=7.33 $Y=1.44 $X2=0 $Y2=0
cc_416 N_B_M1035_g N_Y_c_856_n 0.0134678f $X=7.33 $Y=0.655 $X2=0 $Y2=0
cc_417 N_B_c_508_n N_Y_c_856_n 0.0175552f $X=7.31 $Y=1.44 $X2=0 $Y2=0
cc_418 N_B_c_510_n N_Y_c_856_n 0.00171432f $X=7.33 $Y=1.44 $X2=0 $Y2=0
cc_419 N_B_c_508_n N_Y_c_858_n 0.0112077f $X=7.31 $Y=1.44 $X2=0 $Y2=0
cc_420 N_B_c_509_n N_Y_c_858_n 0.0036624f $X=5.95 $Y=1.44 $X2=0 $Y2=0
cc_421 N_B_c_510_n N_Y_c_858_n 0.00257649f $X=7.33 $Y=1.44 $X2=0 $Y2=0
cc_422 N_B_c_508_n N_Y_c_859_n 0.014687f $X=7.31 $Y=1.44 $X2=0 $Y2=0
cc_423 N_B_c_510_n N_Y_c_859_n 0.00257649f $X=7.33 $Y=1.44 $X2=0 $Y2=0
cc_424 N_B_M1008_g Y 3.95178e-19 $X=6.035 $Y=2.465 $X2=0 $Y2=0
cc_425 N_B_M1006_g Y 0.00218583f $X=6.04 $Y=0.655 $X2=0 $Y2=0
cc_426 N_B_c_509_n Y 0.0270911f $X=5.95 $Y=1.44 $X2=0 $Y2=0
cc_427 N_B_c_510_n Y 0.00487102f $X=7.33 $Y=1.44 $X2=0 $Y2=0
cc_428 N_B_M1008_g N_Y_c_867_n 0.00196532f $X=6.035 $Y=2.465 $X2=0 $Y2=0
cc_429 N_B_c_509_n N_Y_c_867_n 0.0130513f $X=5.95 $Y=1.44 $X2=0 $Y2=0
cc_430 N_B_M1008_g N_A_774_349#_c_1027_n 0.0133475f $X=6.035 $Y=2.465 $X2=0
+ $Y2=0
cc_431 N_B_M1008_g N_A_774_349#_c_1043_n 0.0116414f $X=6.035 $Y=2.465 $X2=0
+ $Y2=0
cc_432 N_B_M1014_g N_A_774_349#_c_1043_n 0.00707931f $X=6.465 $Y=2.465 $X2=0
+ $Y2=0
cc_433 N_B_M1021_g N_A_774_349#_c_1043_n 5.31039e-19 $X=6.895 $Y=2.465 $X2=0
+ $Y2=0
cc_434 N_B_M1014_g N_A_774_349#_c_1046_n 0.0110641f $X=6.465 $Y=2.465 $X2=0
+ $Y2=0
cc_435 N_B_M1021_g N_A_774_349#_c_1046_n 0.0110641f $X=6.895 $Y=2.465 $X2=0
+ $Y2=0
cc_436 N_B_M1021_g N_A_774_349#_c_1048_n 6.34972e-19 $X=6.895 $Y=2.465 $X2=0
+ $Y2=0
cc_437 N_B_M1033_g N_A_774_349#_c_1048_n 0.00213579f $X=7.325 $Y=2.465 $X2=0
+ $Y2=0
cc_438 N_B_M1014_g N_A_774_349#_c_1050_n 6.34958e-19 $X=6.465 $Y=2.465 $X2=0
+ $Y2=0
cc_439 N_B_M1021_g N_A_774_349#_c_1050_n 0.00994996f $X=6.895 $Y=2.465 $X2=0
+ $Y2=0
cc_440 N_B_M1033_g N_A_774_349#_c_1050_n 0.00871855f $X=7.325 $Y=2.465 $X2=0
+ $Y2=0
cc_441 N_B_M1008_g N_A_774_349#_c_1053_n 6.26406e-19 $X=6.035 $Y=2.465 $X2=0
+ $Y2=0
cc_442 N_B_M1014_g N_A_774_349#_c_1053_n 6.26406e-19 $X=6.465 $Y=2.465 $X2=0
+ $Y2=0
cc_443 N_B_c_509_n N_A_1139_367#_c_1090_n 0.00959823f $X=5.95 $Y=1.44 $X2=0
+ $Y2=0
cc_444 N_B_c_510_n N_A_1139_367#_c_1090_n 5.90803e-19 $X=7.33 $Y=1.44 $X2=0
+ $Y2=0
cc_445 N_B_M1008_g N_A_1139_367#_c_1099_n 0.0124169f $X=6.035 $Y=2.465 $X2=0
+ $Y2=0
cc_446 N_B_M1014_g N_A_1139_367#_c_1099_n 0.0118226f $X=6.465 $Y=2.465 $X2=0
+ $Y2=0
cc_447 N_B_c_508_n N_A_1139_367#_c_1099_n 0.00805623f $X=7.31 $Y=1.44 $X2=0
+ $Y2=0
cc_448 N_B_c_509_n N_A_1139_367#_c_1099_n 0.0160685f $X=5.95 $Y=1.44 $X2=0 $Y2=0
cc_449 N_B_c_510_n N_A_1139_367#_c_1099_n 0.00183567f $X=7.33 $Y=1.44 $X2=0
+ $Y2=0
cc_450 N_B_M1008_g N_A_1139_367#_c_1104_n 7.77357e-19 $X=6.035 $Y=2.465 $X2=0
+ $Y2=0
cc_451 N_B_M1014_g N_A_1139_367#_c_1104_n 0.0028166f $X=6.465 $Y=2.465 $X2=0
+ $Y2=0
cc_452 N_B_M1021_g N_A_1139_367#_c_1092_n 0.013791f $X=6.895 $Y=2.465 $X2=0
+ $Y2=0
cc_453 N_B_M1033_g N_A_1139_367#_c_1092_n 0.0135329f $X=7.325 $Y=2.465 $X2=0
+ $Y2=0
cc_454 N_B_c_508_n N_A_1139_367#_c_1092_n 0.0447054f $X=7.31 $Y=1.44 $X2=0 $Y2=0
cc_455 N_B_c_510_n N_A_1139_367#_c_1092_n 0.00359093f $X=7.33 $Y=1.44 $X2=0
+ $Y2=0
cc_456 N_B_M1008_g N_A_1139_367#_c_1093_n 3.34568e-19 $X=6.035 $Y=2.465 $X2=0
+ $Y2=0
cc_457 N_B_M1014_g N_A_1139_367#_c_1093_n 0.00447448f $X=6.465 $Y=2.465 $X2=0
+ $Y2=0
cc_458 N_B_c_508_n N_A_1139_367#_c_1093_n 0.0198477f $X=7.31 $Y=1.44 $X2=0 $Y2=0
cc_459 N_B_c_509_n N_A_1139_367#_c_1093_n 0.00681022f $X=5.95 $Y=1.44 $X2=0
+ $Y2=0
cc_460 N_B_c_510_n N_A_1139_367#_c_1093_n 0.00257649f $X=7.33 $Y=1.44 $X2=0
+ $Y2=0
cc_461 N_B_c_508_n N_A_1139_367#_c_1094_n 0.00231855f $X=7.31 $Y=1.44 $X2=0
+ $Y2=0
cc_462 N_B_c_510_n N_A_1139_367#_c_1094_n 7.66562e-19 $X=7.33 $Y=1.44 $X2=0
+ $Y2=0
cc_463 N_B_M1014_g N_A_1139_367#_c_1117_n 0.001918f $X=6.465 $Y=2.465 $X2=0
+ $Y2=0
cc_464 N_B_M1006_g N_VGND_c_1164_n 0.0110436f $X=6.04 $Y=0.655 $X2=0 $Y2=0
cc_465 N_B_M1023_g N_VGND_c_1164_n 6.2389e-19 $X=6.47 $Y=0.655 $X2=0 $Y2=0
cc_466 N_B_M1006_g N_VGND_c_1165_n 6.14008e-19 $X=6.04 $Y=0.655 $X2=0 $Y2=0
cc_467 N_B_M1023_g N_VGND_c_1165_n 0.010177f $X=6.47 $Y=0.655 $X2=0 $Y2=0
cc_468 N_B_M1024_g N_VGND_c_1165_n 0.010177f $X=6.9 $Y=0.655 $X2=0 $Y2=0
cc_469 N_B_M1035_g N_VGND_c_1165_n 6.14008e-19 $X=7.33 $Y=0.655 $X2=0 $Y2=0
cc_470 N_B_M1024_g N_VGND_c_1166_n 0.00486043f $X=6.9 $Y=0.655 $X2=0 $Y2=0
cc_471 N_B_M1035_g N_VGND_c_1166_n 0.00486043f $X=7.33 $Y=0.655 $X2=0 $Y2=0
cc_472 N_B_M1024_g N_VGND_c_1167_n 6.14008e-19 $X=6.9 $Y=0.655 $X2=0 $Y2=0
cc_473 N_B_M1035_g N_VGND_c_1167_n 0.0101412f $X=7.33 $Y=0.655 $X2=0 $Y2=0
cc_474 N_B_M1006_g N_VGND_c_1171_n 0.00486043f $X=6.04 $Y=0.655 $X2=0 $Y2=0
cc_475 N_B_M1023_g N_VGND_c_1171_n 0.00486043f $X=6.47 $Y=0.655 $X2=0 $Y2=0
cc_476 N_B_M1006_g N_VGND_c_1188_n 0.00824727f $X=6.04 $Y=0.655 $X2=0 $Y2=0
cc_477 N_B_M1023_g N_VGND_c_1188_n 0.00824727f $X=6.47 $Y=0.655 $X2=0 $Y2=0
cc_478 N_B_M1024_g N_VGND_c_1188_n 0.00824727f $X=6.9 $Y=0.655 $X2=0 $Y2=0
cc_479 N_B_M1035_g N_VGND_c_1188_n 0.00824727f $X=7.33 $Y=0.655 $X2=0 $Y2=0
cc_480 N_A_M1003_g N_VPWR_c_686_n 0.0158178f $X=7.76 $Y=2.465 $X2=0 $Y2=0
cc_481 N_A_M1011_g N_VPWR_c_686_n 0.0146175f $X=8.19 $Y=2.465 $X2=0 $Y2=0
cc_482 N_A_M1020_g N_VPWR_c_686_n 6.77662e-19 $X=8.62 $Y=2.465 $X2=0 $Y2=0
cc_483 N_A_M1011_g N_VPWR_c_687_n 6.77662e-19 $X=8.19 $Y=2.465 $X2=0 $Y2=0
cc_484 N_A_M1020_g N_VPWR_c_687_n 0.0146175f $X=8.62 $Y=2.465 $X2=0 $Y2=0
cc_485 N_A_M1025_g N_VPWR_c_687_n 0.0165018f $X=9.05 $Y=2.465 $X2=0 $Y2=0
cc_486 N_A_M1003_g N_VPWR_c_689_n 0.00486043f $X=7.76 $Y=2.465 $X2=0 $Y2=0
cc_487 N_A_M1011_g N_VPWR_c_690_n 0.00486043f $X=8.19 $Y=2.465 $X2=0 $Y2=0
cc_488 N_A_M1020_g N_VPWR_c_690_n 0.00486043f $X=8.62 $Y=2.465 $X2=0 $Y2=0
cc_489 N_A_M1025_g N_VPWR_c_691_n 0.00486043f $X=9.05 $Y=2.465 $X2=0 $Y2=0
cc_490 N_A_M1003_g N_VPWR_c_684_n 0.00828469f $X=7.76 $Y=2.465 $X2=0 $Y2=0
cc_491 N_A_M1011_g N_VPWR_c_684_n 0.00824727f $X=8.19 $Y=2.465 $X2=0 $Y2=0
cc_492 N_A_M1020_g N_VPWR_c_684_n 0.00824727f $X=8.62 $Y=2.465 $X2=0 $Y2=0
cc_493 N_A_M1025_g N_VPWR_c_684_n 0.00924348f $X=9.05 $Y=2.465 $X2=0 $Y2=0
cc_494 N_A_M1016_g N_Y_c_856_n 0.0168144f $X=7.76 $Y=0.655 $X2=0 $Y2=0
cc_495 A N_Y_c_856_n 0.00553546f $X=9.275 $Y=1.58 $X2=0 $Y2=0
cc_496 N_A_M1017_g N_Y_c_857_n 0.0135881f $X=8.19 $Y=0.655 $X2=0 $Y2=0
cc_497 N_A_M1018_g N_Y_c_857_n 0.0134347f $X=8.62 $Y=0.655 $X2=0 $Y2=0
cc_498 N_A_M1031_g N_Y_c_857_n 0.00285015f $X=9.05 $Y=0.655 $X2=0 $Y2=0
cc_499 A N_Y_c_857_n 0.0608615f $X=9.275 $Y=1.58 $X2=0 $Y2=0
cc_500 N_A_c_616_n N_Y_c_857_n 0.00494626f $X=9.125 $Y=1.46 $X2=0 $Y2=0
cc_501 A N_Y_c_860_n 0.0143344f $X=9.275 $Y=1.58 $X2=0 $Y2=0
cc_502 N_A_c_616_n N_Y_c_860_n 0.00252923f $X=9.125 $Y=1.46 $X2=0 $Y2=0
cc_503 N_A_M1003_g N_A_1139_367#_c_1094_n 0.00501369f $X=7.76 $Y=2.465 $X2=0
+ $Y2=0
cc_504 A N_A_1139_367#_c_1094_n 0.0048137f $X=9.275 $Y=1.58 $X2=0 $Y2=0
cc_505 N_A_M1003_g N_A_1139_367#_c_1120_n 0.0155885f $X=7.76 $Y=2.465 $X2=0
+ $Y2=0
cc_506 N_A_M1011_g N_A_1139_367#_c_1120_n 0.0122129f $X=8.19 $Y=2.465 $X2=0
+ $Y2=0
cc_507 A N_A_1139_367#_c_1120_n 0.0335837f $X=9.275 $Y=1.58 $X2=0 $Y2=0
cc_508 N_A_c_616_n N_A_1139_367#_c_1120_n 5.04482e-19 $X=9.125 $Y=1.46 $X2=0
+ $Y2=0
cc_509 N_A_M1020_g N_A_1139_367#_c_1124_n 0.0122595f $X=8.62 $Y=2.465 $X2=0
+ $Y2=0
cc_510 N_A_M1025_g N_A_1139_367#_c_1124_n 0.0122595f $X=9.05 $Y=2.465 $X2=0
+ $Y2=0
cc_511 A N_A_1139_367#_c_1124_n 0.0434214f $X=9.275 $Y=1.58 $X2=0 $Y2=0
cc_512 N_A_c_616_n N_A_1139_367#_c_1124_n 5.04482e-19 $X=9.125 $Y=1.46 $X2=0
+ $Y2=0
cc_513 A N_A_1139_367#_c_1095_n 0.0223278f $X=9.275 $Y=1.58 $X2=0 $Y2=0
cc_514 N_A_c_617_n N_A_1139_367#_c_1095_n 0.00145637f $X=9.33 $Y=1.46 $X2=0
+ $Y2=0
cc_515 A N_A_1139_367#_c_1130_n 0.0155814f $X=9.275 $Y=1.58 $X2=0 $Y2=0
cc_516 N_A_c_616_n N_A_1139_367#_c_1130_n 5.70981e-19 $X=9.125 $Y=1.46 $X2=0
+ $Y2=0
cc_517 N_A_M1016_g N_VGND_c_1167_n 0.0101412f $X=7.76 $Y=0.655 $X2=0 $Y2=0
cc_518 N_A_M1017_g N_VGND_c_1167_n 6.14008e-19 $X=8.19 $Y=0.655 $X2=0 $Y2=0
cc_519 N_A_M1016_g N_VGND_c_1168_n 6.14008e-19 $X=7.76 $Y=0.655 $X2=0 $Y2=0
cc_520 N_A_M1017_g N_VGND_c_1168_n 0.010177f $X=8.19 $Y=0.655 $X2=0 $Y2=0
cc_521 N_A_M1018_g N_VGND_c_1168_n 0.0102576f $X=8.62 $Y=0.655 $X2=0 $Y2=0
cc_522 N_A_M1031_g N_VGND_c_1168_n 6.28227e-19 $X=9.05 $Y=0.655 $X2=0 $Y2=0
cc_523 N_A_M1031_g N_VGND_c_1170_n 0.00707768f $X=9.05 $Y=0.655 $X2=0 $Y2=0
cc_524 A N_VGND_c_1170_n 0.0172135f $X=9.275 $Y=1.58 $X2=0 $Y2=0
cc_525 N_A_c_617_n N_VGND_c_1170_n 0.00707122f $X=9.33 $Y=1.46 $X2=0 $Y2=0
cc_526 N_A_M1016_g N_VGND_c_1178_n 0.00486043f $X=7.76 $Y=0.655 $X2=0 $Y2=0
cc_527 N_A_M1017_g N_VGND_c_1178_n 0.00486043f $X=8.19 $Y=0.655 $X2=0 $Y2=0
cc_528 N_A_M1018_g N_VGND_c_1179_n 0.00486043f $X=8.62 $Y=0.655 $X2=0 $Y2=0
cc_529 N_A_M1031_g N_VGND_c_1179_n 0.00585385f $X=9.05 $Y=0.655 $X2=0 $Y2=0
cc_530 N_A_M1016_g N_VGND_c_1188_n 0.00824727f $X=7.76 $Y=0.655 $X2=0 $Y2=0
cc_531 N_A_M1017_g N_VGND_c_1188_n 0.00824727f $X=8.19 $Y=0.655 $X2=0 $Y2=0
cc_532 N_A_M1018_g N_VGND_c_1188_n 0.00824727f $X=8.62 $Y=0.655 $X2=0 $Y2=0
cc_533 N_A_M1031_g N_VGND_c_1188_n 0.0115186f $X=9.05 $Y=0.655 $X2=0 $Y2=0
cc_534 N_VPWR_c_689_n N_A_347_349#_c_789_n 0.0333877f $X=7.81 $Y=3.33 $X2=0
+ $Y2=0
cc_535 N_VPWR_c_684_n N_A_347_349#_c_789_n 0.0187857f $X=9.36 $Y=3.33 $X2=0
+ $Y2=0
cc_536 N_VPWR_c_689_n N_A_347_349#_c_790_n 0.0516336f $X=7.81 $Y=3.33 $X2=0
+ $Y2=0
cc_537 N_VPWR_c_684_n N_A_347_349#_c_790_n 0.0287249f $X=9.36 $Y=3.33 $X2=0
+ $Y2=0
cc_538 N_VPWR_c_689_n N_A_347_349#_c_791_n 0.0226238f $X=7.81 $Y=3.33 $X2=0
+ $Y2=0
cc_539 N_VPWR_c_684_n N_A_347_349#_c_791_n 0.0124909f $X=9.36 $Y=3.33 $X2=0
+ $Y2=0
cc_540 N_VPWR_c_689_n N_A_347_349#_c_792_n 0.0234809f $X=7.81 $Y=3.33 $X2=0
+ $Y2=0
cc_541 N_VPWR_c_684_n N_A_347_349#_c_792_n 0.0126009f $X=9.36 $Y=3.33 $X2=0
+ $Y2=0
cc_542 N_VPWR_c_684_n N_A_774_349#_M1008_s 0.00223559f $X=9.36 $Y=3.33 $X2=0
+ $Y2=0
cc_543 N_VPWR_c_684_n N_A_774_349#_M1021_s 0.00223559f $X=9.36 $Y=3.33 $X2=0
+ $Y2=0
cc_544 N_VPWR_c_689_n N_A_774_349#_c_1025_n 0.0333615f $X=7.81 $Y=3.33 $X2=0
+ $Y2=0
cc_545 N_VPWR_c_684_n N_A_774_349#_c_1025_n 0.0187823f $X=9.36 $Y=3.33 $X2=0
+ $Y2=0
cc_546 N_VPWR_c_689_n N_A_774_349#_c_1026_n 0.0235321f $X=7.81 $Y=3.33 $X2=0
+ $Y2=0
cc_547 N_VPWR_c_684_n N_A_774_349#_c_1026_n 0.0126106f $X=9.36 $Y=3.33 $X2=0
+ $Y2=0
cc_548 N_VPWR_c_689_n N_A_774_349#_c_1027_n 0.0654595f $X=7.81 $Y=3.33 $X2=0
+ $Y2=0
cc_549 N_VPWR_c_684_n N_A_774_349#_c_1027_n 0.0384259f $X=9.36 $Y=3.33 $X2=0
+ $Y2=0
cc_550 N_VPWR_c_689_n N_A_774_349#_c_1046_n 0.0300582f $X=7.81 $Y=3.33 $X2=0
+ $Y2=0
cc_551 N_VPWR_c_684_n N_A_774_349#_c_1046_n 0.0188286f $X=9.36 $Y=3.33 $X2=0
+ $Y2=0
cc_552 N_VPWR_c_689_n N_A_774_349#_c_1048_n 0.01906f $X=7.81 $Y=3.33 $X2=0 $Y2=0
cc_553 N_VPWR_c_684_n N_A_774_349#_c_1048_n 0.0124545f $X=9.36 $Y=3.33 $X2=0
+ $Y2=0
cc_554 N_VPWR_c_689_n N_A_774_349#_c_1028_n 0.0235321f $X=7.81 $Y=3.33 $X2=0
+ $Y2=0
cc_555 N_VPWR_c_684_n N_A_774_349#_c_1028_n 0.0126106f $X=9.36 $Y=3.33 $X2=0
+ $Y2=0
cc_556 N_VPWR_c_689_n N_A_774_349#_c_1053_n 0.0190915f $X=7.81 $Y=3.33 $X2=0
+ $Y2=0
cc_557 N_VPWR_c_684_n N_A_774_349#_c_1053_n 0.0124642f $X=9.36 $Y=3.33 $X2=0
+ $Y2=0
cc_558 N_VPWR_c_684_n N_A_1139_367#_M1008_d 0.0021598f $X=9.36 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_559 N_VPWR_c_684_n N_A_1139_367#_M1014_d 0.00225186f $X=9.36 $Y=3.33 $X2=0
+ $Y2=0
cc_560 N_VPWR_c_684_n N_A_1139_367#_M1033_d 0.00540667f $X=9.36 $Y=3.33 $X2=0
+ $Y2=0
cc_561 N_VPWR_c_684_n N_A_1139_367#_M1011_s 0.00536646f $X=9.36 $Y=3.33 $X2=0
+ $Y2=0
cc_562 N_VPWR_c_684_n N_A_1139_367#_M1025_s 0.00371702f $X=9.36 $Y=3.33 $X2=0
+ $Y2=0
cc_563 N_VPWR_c_689_n N_A_1139_367#_c_1137_n 0.012804f $X=7.81 $Y=3.33 $X2=0
+ $Y2=0
cc_564 N_VPWR_c_684_n N_A_1139_367#_c_1137_n 0.00750339f $X=9.36 $Y=3.33 $X2=0
+ $Y2=0
cc_565 N_VPWR_M1003_d N_A_1139_367#_c_1120_n 0.00334931f $X=7.835 $Y=1.835 $X2=0
+ $Y2=0
cc_566 N_VPWR_c_686_n N_A_1139_367#_c_1120_n 0.0170777f $X=7.975 $Y=2.38 $X2=0
+ $Y2=0
cc_567 N_VPWR_c_690_n N_A_1139_367#_c_1141_n 0.0124525f $X=8.67 $Y=3.33 $X2=0
+ $Y2=0
cc_568 N_VPWR_c_684_n N_A_1139_367#_c_1141_n 0.00730901f $X=9.36 $Y=3.33 $X2=0
+ $Y2=0
cc_569 N_VPWR_M1020_d N_A_1139_367#_c_1124_n 0.00334931f $X=8.695 $Y=1.835 $X2=0
+ $Y2=0
cc_570 N_VPWR_c_687_n N_A_1139_367#_c_1124_n 0.0170777f $X=8.835 $Y=2.38 $X2=0
+ $Y2=0
cc_571 N_VPWR_c_691_n N_A_1139_367#_c_1096_n 0.0178111f $X=9.36 $Y=3.33 $X2=0
+ $Y2=0
cc_572 N_VPWR_c_684_n N_A_1139_367#_c_1096_n 0.0100304f $X=9.36 $Y=3.33 $X2=0
+ $Y2=0
cc_573 N_A_347_349#_c_789_n N_Y_M1005_s 0.00176461f $X=2.555 $Y=2.99 $X2=0 $Y2=0
cc_574 N_A_347_349#_c_790_n N_Y_M1019_s 0.00176461f $X=3.455 $Y=2.99 $X2=0 $Y2=0
cc_575 N_A_347_349#_c_789_n N_Y_c_960_n 0.0126348f $X=2.555 $Y=2.99 $X2=0 $Y2=0
cc_576 N_A_347_349#_M1012_d N_Y_c_862_n 0.00176461f $X=2.58 $Y=1.745 $X2=0 $Y2=0
cc_577 N_A_347_349#_c_799_n N_Y_c_862_n 0.0170777f $X=2.72 $Y=2.11 $X2=0 $Y2=0
cc_578 N_A_347_349#_c_790_n N_Y_c_963_n 0.0126348f $X=3.455 $Y=2.99 $X2=0 $Y2=0
cc_579 N_A_347_349#_M1030_d N_Y_c_864_n 0.00176773f $X=3.44 $Y=1.745 $X2=0 $Y2=0
cc_580 N_A_347_349#_M1007_s N_Y_c_864_n 0.00176773f $X=4.3 $Y=1.745 $X2=0 $Y2=0
cc_581 N_A_347_349#_M1027_s N_Y_c_864_n 3.40767e-19 $X=5.16 $Y=1.745 $X2=0 $Y2=0
cc_582 N_A_347_349#_c_833_p N_Y_c_864_n 0.0135577f $X=3.565 $Y=2.205 $X2=0 $Y2=0
cc_583 N_A_347_349#_c_811_n N_Y_c_864_n 0.0324652f $X=4.345 $Y=2.12 $X2=0 $Y2=0
cc_584 N_A_347_349#_c_813_n N_Y_c_864_n 0.0324652f $X=5.205 $Y=2.12 $X2=0 $Y2=0
cc_585 N_A_347_349#_c_836_p N_Y_c_864_n 0.0135898f $X=4.44 $Y=2.12 $X2=0 $Y2=0
cc_586 N_A_347_349#_c_793_n N_Y_c_864_n 0.00265841f $X=5.3 $Y=2.2 $X2=0 $Y2=0
cc_587 N_A_347_349#_M1027_s N_Y_c_867_n 0.00240707f $X=5.16 $Y=1.745 $X2=0 $Y2=0
cc_588 N_A_347_349#_c_793_n N_Y_c_867_n 0.0195262f $X=5.3 $Y=2.2 $X2=0 $Y2=0
cc_589 N_A_347_349#_c_811_n N_A_774_349#_M1001_d 0.00339939f $X=4.345 $Y=2.12
+ $X2=-0.19 $Y2=1.655
cc_590 N_A_347_349#_c_813_n N_A_774_349#_M1013_d 0.00339939f $X=5.205 $Y=2.12
+ $X2=0 $Y2=0
cc_591 N_A_347_349#_c_811_n N_A_774_349#_c_1029_n 0.0171184f $X=4.345 $Y=2.12
+ $X2=0 $Y2=0
cc_592 N_A_347_349#_M1007_s N_A_774_349#_c_1025_n 0.00176461f $X=4.3 $Y=1.745
+ $X2=0 $Y2=0
cc_593 N_A_347_349#_c_844_p N_A_774_349#_c_1025_n 0.0126631f $X=4.44 $Y=2.57
+ $X2=0 $Y2=0
cc_594 N_A_347_349#_c_790_n N_A_774_349#_c_1026_n 0.0104256f $X=3.455 $Y=2.99
+ $X2=0 $Y2=0
cc_595 N_A_347_349#_c_813_n N_A_774_349#_c_1036_n 0.0171184f $X=5.205 $Y=2.12
+ $X2=0 $Y2=0
cc_596 N_A_347_349#_M1027_s N_A_774_349#_c_1027_n 0.00277855f $X=5.16 $Y=1.745
+ $X2=0 $Y2=0
cc_597 N_A_347_349#_c_793_n N_A_774_349#_c_1027_n 0.0191464f $X=5.3 $Y=2.2 $X2=0
+ $Y2=0
cc_598 N_A_347_349#_c_793_n N_A_1139_367#_c_1090_n 0.0147157f $X=5.3 $Y=2.2
+ $X2=0 $Y2=0
cc_599 N_A_347_349#_c_793_n N_A_1139_367#_c_1091_n 0.0378048f $X=5.3 $Y=2.2
+ $X2=0 $Y2=0
cc_600 N_Y_c_864_n N_A_774_349#_M1001_d 0.00177204f $X=5.25 $Y=1.775 $X2=-0.19
+ $Y2=-0.245
cc_601 N_Y_c_864_n N_A_774_349#_M1013_d 0.00177204f $X=5.25 $Y=1.775 $X2=0 $Y2=0
cc_602 N_Y_c_856_n N_A_1139_367#_c_1094_n 0.00574729f $X=7.88 $Y=1.09 $X2=0
+ $Y2=0
cc_603 N_Y_c_871_n N_VGND_M1009_d 0.00753335f $X=3.055 $Y=0.74 $X2=0 $Y2=0
cc_604 N_Y_c_889_n N_VGND_M1029_d 0.00480725f $X=4.055 $Y=0.74 $X2=0 $Y2=0
cc_605 N_Y_c_851_n N_VGND_M1004_s 0.00176461f $X=4.915 $Y=1.08 $X2=0 $Y2=0
cc_606 N_Y_c_853_n N_VGND_M1034_s 0.00394721f $X=6.16 $Y=1.08 $X2=0 $Y2=0
cc_607 N_Y_c_854_n N_VGND_M1034_s 0.0035276f $X=5.615 $Y=1.08 $X2=0 $Y2=0
cc_608 N_Y_c_855_n N_VGND_M1023_d 0.00176461f $X=7.02 $Y=1.09 $X2=0 $Y2=0
cc_609 N_Y_c_856_n N_VGND_M1035_d 0.00176461f $X=7.88 $Y=1.09 $X2=0 $Y2=0
cc_610 N_Y_c_857_n N_VGND_M1017_s 0.00176461f $X=8.74 $Y=1.09 $X2=0 $Y2=0
cc_611 N_Y_c_871_n N_VGND_c_1160_n 0.0250837f $X=3.055 $Y=0.74 $X2=0 $Y2=0
cc_612 N_Y_c_883_n N_VGND_c_1160_n 0.0163868f $X=3.22 $Y=0.36 $X2=0 $Y2=0
cc_613 N_Y_c_871_n N_VGND_c_1161_n 0.00259694f $X=3.055 $Y=0.74 $X2=0 $Y2=0
cc_614 N_Y_c_883_n N_VGND_c_1161_n 0.0187344f $X=3.22 $Y=0.36 $X2=0 $Y2=0
cc_615 N_Y_c_889_n N_VGND_c_1161_n 0.00235176f $X=4.055 $Y=0.74 $X2=0 $Y2=0
cc_616 N_Y_c_889_n N_VGND_c_1162_n 0.0197854f $X=4.055 $Y=0.74 $X2=0 $Y2=0
cc_617 N_Y_c_851_n N_VGND_c_1163_n 0.0170777f $X=4.915 $Y=1.08 $X2=0 $Y2=0
cc_618 N_Y_c_853_n N_VGND_c_1164_n 0.0257809f $X=6.16 $Y=1.08 $X2=0 $Y2=0
cc_619 N_Y_c_854_n N_VGND_c_1164_n 0.025251f $X=5.615 $Y=1.08 $X2=0 $Y2=0
cc_620 N_Y_c_855_n N_VGND_c_1165_n 0.0170777f $X=7.02 $Y=1.09 $X2=0 $Y2=0
cc_621 N_Y_c_995_p N_VGND_c_1166_n 0.0124525f $X=7.115 $Y=0.42 $X2=0 $Y2=0
cc_622 N_Y_c_856_n N_VGND_c_1167_n 0.0170777f $X=7.88 $Y=1.09 $X2=0 $Y2=0
cc_623 N_Y_c_857_n N_VGND_c_1168_n 0.0170777f $X=8.74 $Y=1.09 $X2=0 $Y2=0
cc_624 N_Y_c_857_n N_VGND_c_1170_n 0.00166618f $X=8.74 $Y=1.09 $X2=0 $Y2=0
cc_625 N_Y_c_999_p N_VGND_c_1171_n 0.0124525f $X=6.255 $Y=0.42 $X2=0 $Y2=0
cc_626 N_Y_c_868_n N_VGND_c_1175_n 0.0194075f $X=2.19 $Y=0.36 $X2=0 $Y2=0
cc_627 N_Y_c_871_n N_VGND_c_1175_n 0.00228867f $X=3.055 $Y=0.74 $X2=0 $Y2=0
cc_628 N_Y_c_889_n N_VGND_c_1176_n 0.00235807f $X=4.055 $Y=0.74 $X2=0 $Y2=0
cc_629 N_Y_c_1003_p N_VGND_c_1176_n 0.0124525f $X=4.15 $Y=0.42 $X2=0 $Y2=0
cc_630 N_Y_c_1004_p N_VGND_c_1177_n 0.0124525f $X=5.01 $Y=0.42 $X2=0 $Y2=0
cc_631 N_Y_c_1005_p N_VGND_c_1178_n 0.0124525f $X=7.975 $Y=0.42 $X2=0 $Y2=0
cc_632 N_Y_c_1006_p N_VGND_c_1179_n 0.0136943f $X=8.835 $Y=0.42 $X2=0 $Y2=0
cc_633 N_Y_M1002_s N_VGND_c_1188_n 0.00223559f $X=2.05 $Y=0.235 $X2=0 $Y2=0
cc_634 N_Y_M1026_s N_VGND_c_1188_n 0.00223559f $X=3.08 $Y=0.235 $X2=0 $Y2=0
cc_635 N_Y_M1000_d N_VGND_c_1188_n 0.00396356f $X=4.01 $Y=0.235 $X2=0 $Y2=0
cc_636 N_Y_M1022_d N_VGND_c_1188_n 0.00536646f $X=4.87 $Y=0.235 $X2=0 $Y2=0
cc_637 N_Y_M1006_s N_VGND_c_1188_n 0.00536646f $X=6.115 $Y=0.235 $X2=0 $Y2=0
cc_638 N_Y_M1024_s N_VGND_c_1188_n 0.00536646f $X=6.975 $Y=0.235 $X2=0 $Y2=0
cc_639 N_Y_M1016_d N_VGND_c_1188_n 0.00536646f $X=7.835 $Y=0.235 $X2=0 $Y2=0
cc_640 N_Y_M1018_d N_VGND_c_1188_n 0.0041489f $X=8.695 $Y=0.235 $X2=0 $Y2=0
cc_641 N_Y_c_868_n N_VGND_c_1188_n 0.0126695f $X=2.19 $Y=0.36 $X2=0 $Y2=0
cc_642 N_Y_c_871_n N_VGND_c_1188_n 0.0103708f $X=3.055 $Y=0.74 $X2=0 $Y2=0
cc_643 N_Y_c_883_n N_VGND_c_1188_n 0.0123282f $X=3.22 $Y=0.36 $X2=0 $Y2=0
cc_644 N_Y_c_889_n N_VGND_c_1188_n 0.00969956f $X=4.055 $Y=0.74 $X2=0 $Y2=0
cc_645 N_Y_c_1003_p N_VGND_c_1188_n 0.00730901f $X=4.15 $Y=0.42 $X2=0 $Y2=0
cc_646 N_Y_c_1004_p N_VGND_c_1188_n 0.00730901f $X=5.01 $Y=0.42 $X2=0 $Y2=0
cc_647 N_Y_c_999_p N_VGND_c_1188_n 0.00730901f $X=6.255 $Y=0.42 $X2=0 $Y2=0
cc_648 N_Y_c_995_p N_VGND_c_1188_n 0.00730901f $X=7.115 $Y=0.42 $X2=0 $Y2=0
cc_649 N_Y_c_1005_p N_VGND_c_1188_n 0.00730901f $X=7.975 $Y=0.42 $X2=0 $Y2=0
cc_650 N_Y_c_1006_p N_VGND_c_1188_n 0.00866972f $X=8.835 $Y=0.42 $X2=0 $Y2=0
cc_651 N_A_774_349#_c_1027_n N_A_1139_367#_M1008_d 0.00506312f $X=6.085 $Y=2.98
+ $X2=-0.19 $Y2=1.655
cc_652 N_A_774_349#_c_1046_n N_A_1139_367#_M1014_d 0.00333487f $X=6.945 $Y=2.98
+ $X2=0 $Y2=0
cc_653 N_A_774_349#_c_1027_n N_A_1139_367#_c_1091_n 0.0191464f $X=6.085 $Y=2.98
+ $X2=0 $Y2=0
cc_654 N_A_774_349#_M1008_s N_A_1139_367#_c_1099_n 0.0042115f $X=6.11 $Y=1.835
+ $X2=0 $Y2=0
cc_655 N_A_774_349#_c_1043_n N_A_1139_367#_c_1099_n 0.0171184f $X=6.25 $Y=2.49
+ $X2=0 $Y2=0
cc_656 N_A_774_349#_c_1046_n N_A_1139_367#_c_1155_n 0.0127906f $X=6.945 $Y=2.98
+ $X2=0 $Y2=0
cc_657 N_A_774_349#_M1021_s N_A_1139_367#_c_1092_n 0.00180746f $X=6.97 $Y=1.835
+ $X2=0 $Y2=0
cc_658 N_A_774_349#_c_1050_n N_A_1139_367#_c_1092_n 0.0163515f $X=7.11 $Y=2.14
+ $X2=0 $Y2=0
