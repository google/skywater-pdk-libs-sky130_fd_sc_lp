* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__sdfsbp_lp CLK D SCD SCE SET_B VGND VNB VPB VPWR Q Q_N
X0 a_1201_419# a_987_409# a_1381_125# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 a_761_113# CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X2 a_2019_419# a_987_409# a_2193_419# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X3 a_1729_125# SET_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 VPWR SCD a_245_409# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X5 a_1423_99# SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X6 a_2220_40# a_2019_419# a_2524_57# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 a_352_409# D a_458_409# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X8 a_458_409# SCE VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X9 a_2193_419# a_2220_40# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X10 a_352_409# SCE a_526_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X11 VPWR a_2019_419# Q_N VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X12 VPWR a_2865_74# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X13 VPWR a_1201_419# a_1423_99# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X14 VGND a_761_113# a_1006_113# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X15 a_352_409# a_761_113# a_1201_419# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X16 VGND a_1201_419# a_1915_125# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X17 a_27_409# SCE a_138_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X18 a_2250_66# SET_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X19 a_27_409# SCE VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X20 a_1373_419# a_1423_99# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X21 a_138_47# SCE VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X22 a_2682_57# a_2019_419# Q_N VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X23 a_2172_66# a_2220_40# a_2250_66# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X24 VPWR a_761_113# a_987_409# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X25 a_362_47# D a_352_409# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X26 a_848_113# CLK VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X27 VGND a_2865_74# a_3109_74# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X28 VPWR SET_B a_2019_419# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X29 a_1915_125# a_987_409# a_2019_419# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X30 a_1921_419# a_761_113# a_2019_419# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X31 a_245_409# a_27_409# a_352_409# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X32 a_352_409# a_987_409# a_1201_419# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X33 a_761_113# CLK a_848_113# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X34 a_1006_113# a_761_113# a_987_409# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X35 a_2865_74# a_2019_419# a_2951_74# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X36 VPWR a_1201_419# a_1921_419# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X37 a_2524_57# a_2019_419# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X38 a_1381_125# a_1423_99# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X39 a_1423_99# a_1201_419# a_1729_125# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X40 VGND a_2019_419# a_2682_57# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X41 a_2951_74# a_2019_419# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X42 a_1201_419# a_761_113# a_1373_419# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X43 VGND a_27_409# a_362_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X44 a_526_47# SCD VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X45 a_2019_419# a_761_113# a_2172_66# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X46 a_2865_74# a_2019_419# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X47 a_2220_40# a_2019_419# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X48 a_3109_74# a_2865_74# Q VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
