* File: sky130_fd_sc_lp__a2bb2o_m.pxi.spice
* Created: Fri Aug 28 09:56:20 2020
* 
x_PM_SKY130_FD_SC_LP__A2BB2O_M%A_85_345# N_A_85_345#_M1002_d N_A_85_345#_M1011_s
+ N_A_85_345#_M1006_g N_A_85_345#_M1000_g N_A_85_345#_c_81_n N_A_85_345#_c_82_n
+ N_A_85_345#_c_83_n N_A_85_345#_c_84_n N_A_85_345#_c_73_n N_A_85_345#_c_74_n
+ N_A_85_345#_c_86_n N_A_85_345#_c_75_n N_A_85_345#_c_76_n N_A_85_345#_c_77_n
+ N_A_85_345#_c_78_n PM_SKY130_FD_SC_LP__A2BB2O_M%A_85_345#
x_PM_SKY130_FD_SC_LP__A2BB2O_M%A1_N N_A1_N_M1004_g N_A1_N_M1003_g A1_N A1_N A1_N
+ N_A1_N_c_154_n N_A1_N_c_155_n PM_SKY130_FD_SC_LP__A2BB2O_M%A1_N
x_PM_SKY130_FD_SC_LP__A2BB2O_M%A2_N N_A2_N_M1007_g N_A2_N_M1001_g A2_N A2_N
+ N_A2_N_c_195_n PM_SKY130_FD_SC_LP__A2BB2O_M%A2_N
x_PM_SKY130_FD_SC_LP__A2BB2O_M%A_210_125# N_A_210_125#_M1004_d
+ N_A_210_125#_M1007_d N_A_210_125#_M1002_g N_A_210_125#_c_231_n
+ N_A_210_125#_c_232_n N_A_210_125#_M1011_g N_A_210_125#_c_234_n
+ N_A_210_125#_c_235_n N_A_210_125#_c_238_n N_A_210_125#_c_239_n
+ N_A_210_125#_c_236_n PM_SKY130_FD_SC_LP__A2BB2O_M%A_210_125#
x_PM_SKY130_FD_SC_LP__A2BB2O_M%B2 N_B2_M1009_g N_B2_M1005_g N_B2_c_297_n
+ N_B2_c_298_n N_B2_c_302_n B2 B2 B2 B2 N_B2_c_300_n
+ PM_SKY130_FD_SC_LP__A2BB2O_M%B2
x_PM_SKY130_FD_SC_LP__A2BB2O_M%B1 N_B1_M1010_g N_B1_M1008_g N_B1_c_341_n
+ N_B1_c_342_n N_B1_c_346_n B1 B1 N_B1_c_344_n PM_SKY130_FD_SC_LP__A2BB2O_M%B1
x_PM_SKY130_FD_SC_LP__A2BB2O_M%X N_X_M1006_s N_X_M1000_s X X X X X X X X
+ PM_SKY130_FD_SC_LP__A2BB2O_M%X
x_PM_SKY130_FD_SC_LP__A2BB2O_M%VPWR N_VPWR_M1000_d N_VPWR_M1005_d N_VPWR_c_389_n
+ N_VPWR_c_390_n N_VPWR_c_391_n N_VPWR_c_392_n VPWR N_VPWR_c_393_n
+ N_VPWR_c_388_n N_VPWR_c_395_n PM_SKY130_FD_SC_LP__A2BB2O_M%VPWR
x_PM_SKY130_FD_SC_LP__A2BB2O_M%A_479_429# N_A_479_429#_M1011_d
+ N_A_479_429#_M1008_d N_A_479_429#_c_429_n N_A_479_429#_c_430_n
+ PM_SKY130_FD_SC_LP__A2BB2O_M%A_479_429#
x_PM_SKY130_FD_SC_LP__A2BB2O_M%VGND N_VGND_M1006_d N_VGND_M1001_d N_VGND_M1010_d
+ N_VGND_c_443_n N_VGND_c_456_n N_VGND_c_444_n N_VGND_c_445_n N_VGND_c_450_n
+ VGND N_VGND_c_446_n N_VGND_c_447_n N_VGND_c_448_n
+ PM_SKY130_FD_SC_LP__A2BB2O_M%VGND
cc_1 VNB N_A_85_345#_M1006_g 0.0475844f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=0.835
cc_2 VNB N_A_85_345#_c_73_n 0.0116397f $X=-0.19 $Y=-0.245 $X2=2 $Y2=1.685
cc_3 VNB N_A_85_345#_c_74_n 0.00100495f $X=-0.19 $Y=-0.245 $X2=0.675 $Y2=1.685
cc_4 VNB N_A_85_345#_c_75_n 7.00475e-19 $X=-0.19 $Y=-0.245 $X2=2.21 $Y2=0.9
cc_5 VNB N_A_85_345#_c_76_n 0.00436326f $X=-0.19 $Y=-0.245 $X2=2.13 $Y2=1.6
cc_6 VNB N_A_85_345#_c_77_n 0.00141507f $X=-0.19 $Y=-0.245 $X2=2.107 $Y2=1.685
cc_7 VNB N_A_85_345#_c_78_n 0.00181173f $X=-0.19 $Y=-0.245 $X2=2.21 $Y2=1.38
cc_8 VNB N_A1_N_M1003_g 0.00952534f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB A1_N 0.0155135f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A1_N_c_154_n 0.0305372f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.89
cc_11 VNB N_A1_N_c_155_n 0.0187846f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=2.23
cc_12 VNB N_A2_N_M1001_g 0.0457741f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=1.725
cc_13 VNB N_A_210_125#_M1002_g 0.0128724f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_210_125#_c_231_n 0.0213861f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=2.395
cc_15 VNB N_A_210_125#_c_232_n 0.00957542f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=2.885
cc_16 VNB N_A_210_125#_M1011_g 0.0204654f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.725
cc_17 VNB N_A_210_125#_c_234_n 0.0190919f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.77
cc_18 VNB N_A_210_125#_c_235_n 0.0488448f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.89
cc_19 VNB N_A_210_125#_c_236_n 0.0108726f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_B2_c_297_n 0.0170294f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=0.835
cc_21 VNB N_B2_c_298_n 0.0206202f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB B2 0.0121343f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=2.885
cc_23 VNB N_B2_c_300_n 0.0174671f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.89
cc_24 VNB N_B1_c_341_n 0.0226332f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=0.835
cc_25 VNB N_B1_c_342_n 0.0246446f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB B1 0.0304524f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_B1_c_344_n 0.0188276f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.89
cc_28 VNB X 0.0199306f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=1.725
cc_29 VNB X 0.0366716f $X=-0.19 $Y=-0.245 $X2=0.675 $Y2=1.685
cc_30 VNB N_VPWR_c_388_n 0.163682f $X=-0.19 $Y=-0.245 $X2=2.21 $Y2=0.9
cc_31 VNB N_VGND_c_443_n 0.0210851f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=2.885
cc_32 VNB N_VGND_c_444_n 0.0162041f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.725
cc_33 VNB N_VGND_c_445_n 0.0413337f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=2.395
cc_34 VNB N_VGND_c_446_n 0.0640863f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_447_n 0.025002f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.89
cc_36 VNB N_VGND_c_448_n 0.258753f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VPB N_A_85_345#_M1006_g 0.00370759f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=0.835
cc_38 VPB N_A_85_345#_M1000_g 0.0304582f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=2.885
cc_39 VPB N_A_85_345#_c_81_n 0.0253766f $X=-0.19 $Y=1.655 $X2=0.59 $Y2=2.23
cc_40 VPB N_A_85_345#_c_82_n 0.0184149f $X=-0.19 $Y=1.655 $X2=0.59 $Y2=2.395
cc_41 VPB N_A_85_345#_c_83_n 0.0011811f $X=-0.19 $Y=1.655 $X2=0.59 $Y2=1.89
cc_42 VPB N_A_85_345#_c_84_n 0.0184008f $X=-0.19 $Y=1.655 $X2=0.59 $Y2=1.89
cc_43 VPB N_A_85_345#_c_73_n 0.0199343f $X=-0.19 $Y=1.655 $X2=2 $Y2=1.685
cc_44 VPB N_A_85_345#_c_86_n 0.00927633f $X=-0.19 $Y=1.655 $X2=2.105 $Y2=2.27
cc_45 VPB N_A_85_345#_c_77_n 0.00177569f $X=-0.19 $Y=1.655 $X2=2.107 $Y2=1.685
cc_46 VPB N_A1_N_M1003_g 0.0575225f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_47 VPB N_A2_N_M1007_g 0.0435068f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_48 VPB N_A2_N_M1001_g 0.0129602f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=1.725
cc_49 VPB A2_N 0.015028f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=2.395
cc_50 VPB N_A2_N_c_195_n 0.0377183f $X=-0.19 $Y=1.655 $X2=0.59 $Y2=2.395
cc_51 VPB N_A_210_125#_M1011_g 0.043922f $X=-0.19 $Y=1.655 $X2=0.59 $Y2=1.725
cc_52 VPB N_A_210_125#_c_238_n 0.0138396f $X=-0.19 $Y=1.655 $X2=2.107 $Y2=1.77
cc_53 VPB N_A_210_125#_c_239_n 0.0421843f $X=-0.19 $Y=1.655 $X2=2.107 $Y2=2.27
cc_54 VPB N_B2_M1005_g 0.0280606f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_55 VPB N_B2_c_302_n 0.0151435f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=2.395
cc_56 VPB B2 0.00271714f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=2.885
cc_57 VPB N_B1_M1008_g 0.0396965f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_58 VPB N_B1_c_346_n 0.0190802f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=2.395
cc_59 VPB B1 0.0112676f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_60 VPB X 0.0191647f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=2.885
cc_61 VPB X 0.0479366f $X=-0.19 $Y=1.655 $X2=0.675 $Y2=1.685
cc_62 VPB N_VPWR_c_389_n 4.89148e-19 $X=-0.19 $Y=1.655 $X2=0.61 $Y2=2.395
cc_63 VPB N_VPWR_c_390_n 0.0307237f $X=-0.19 $Y=1.655 $X2=0.59 $Y2=1.89
cc_64 VPB N_VPWR_c_391_n 0.0491592f $X=-0.19 $Y=1.655 $X2=0.59 $Y2=2.395
cc_65 VPB N_VPWR_c_392_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0.59 $Y2=1.77
cc_66 VPB N_VPWR_c_393_n 0.0241005f $X=-0.19 $Y=1.655 $X2=2.21 $Y2=1.215
cc_67 VPB N_VPWR_c_388_n 0.0885158f $X=-0.19 $Y=1.655 $X2=2.21 $Y2=0.9
cc_68 VPB N_VPWR_c_395_n 0.0238348f $X=-0.19 $Y=1.655 $X2=2.13 $Y2=1.38
cc_69 VPB N_A_479_429#_c_429_n 0.0140737f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=2.395
cc_70 VPB N_A_479_429#_c_430_n 0.00673679f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=2.885
cc_71 N_A_85_345#_M1006_g N_A1_N_M1003_g 0.00863047f $X=0.545 $Y=0.835 $X2=0
+ $Y2=0
cc_72 N_A_85_345#_M1000_g N_A1_N_M1003_g 0.0225396f $X=0.61 $Y=2.885 $X2=0 $Y2=0
cc_73 N_A_85_345#_c_83_n N_A1_N_M1003_g 0.00232652f $X=0.59 $Y=1.89 $X2=0 $Y2=0
cc_74 N_A_85_345#_c_84_n N_A1_N_M1003_g 0.0412509f $X=0.59 $Y=1.89 $X2=0 $Y2=0
cc_75 N_A_85_345#_c_73_n N_A1_N_M1003_g 0.0157734f $X=2 $Y=1.685 $X2=0 $Y2=0
cc_76 N_A_85_345#_M1006_g A1_N 0.00227189f $X=0.545 $Y=0.835 $X2=0 $Y2=0
cc_77 N_A_85_345#_c_84_n A1_N 6.3024e-19 $X=0.59 $Y=1.89 $X2=0 $Y2=0
cc_78 N_A_85_345#_c_73_n A1_N 0.0722612f $X=2 $Y=1.685 $X2=0 $Y2=0
cc_79 N_A_85_345#_c_74_n A1_N 0.00309486f $X=0.675 $Y=1.685 $X2=0 $Y2=0
cc_80 N_A_85_345#_c_75_n A1_N 0.0115262f $X=2.21 $Y=0.9 $X2=0 $Y2=0
cc_81 N_A_85_345#_c_73_n N_A1_N_c_154_n 0.00463702f $X=2 $Y=1.685 $X2=0 $Y2=0
cc_82 N_A_85_345#_M1006_g N_A1_N_c_155_n 0.0258329f $X=0.545 $Y=0.835 $X2=0
+ $Y2=0
cc_83 N_A_85_345#_c_86_n N_A2_N_M1007_g 9.0287e-19 $X=2.105 $Y=2.27 $X2=0 $Y2=0
cc_84 N_A_85_345#_c_73_n N_A2_N_M1001_g 0.0123327f $X=2 $Y=1.685 $X2=0 $Y2=0
cc_85 N_A_85_345#_c_86_n N_A2_N_M1001_g 0.00193269f $X=2.105 $Y=2.27 $X2=0 $Y2=0
cc_86 N_A_85_345#_c_75_n N_A2_N_M1001_g 9.32009e-19 $X=2.21 $Y=0.9 $X2=0 $Y2=0
cc_87 N_A_85_345#_c_76_n N_A2_N_M1001_g 0.00346552f $X=2.13 $Y=1.6 $X2=0 $Y2=0
cc_88 N_A_85_345#_c_78_n N_A2_N_M1001_g 3.33473e-19 $X=2.21 $Y=1.38 $X2=0 $Y2=0
cc_89 N_A_85_345#_M1000_g A2_N 4.32286e-19 $X=0.61 $Y=2.885 $X2=0 $Y2=0
cc_90 N_A_85_345#_c_81_n A2_N 0.00128395f $X=0.59 $Y=2.23 $X2=0 $Y2=0
cc_91 N_A_85_345#_c_83_n A2_N 0.0155435f $X=0.59 $Y=1.89 $X2=0 $Y2=0
cc_92 N_A_85_345#_c_73_n A2_N 0.0492036f $X=2 $Y=1.685 $X2=0 $Y2=0
cc_93 N_A_85_345#_c_86_n A2_N 0.0325385f $X=2.105 $Y=2.27 $X2=0 $Y2=0
cc_94 N_A_85_345#_c_73_n N_A2_N_c_195_n 0.00651536f $X=2 $Y=1.685 $X2=0 $Y2=0
cc_95 N_A_85_345#_c_86_n N_A2_N_c_195_n 0.00267311f $X=2.105 $Y=2.27 $X2=0 $Y2=0
cc_96 N_A_85_345#_c_75_n N_A_210_125#_M1002_g 0.00682393f $X=2.21 $Y=0.9 $X2=0
+ $Y2=0
cc_97 N_A_85_345#_c_75_n N_A_210_125#_c_231_n 0.0076187f $X=2.21 $Y=0.9 $X2=0
+ $Y2=0
cc_98 N_A_85_345#_c_78_n N_A_210_125#_c_231_n 0.00694047f $X=2.21 $Y=1.38 $X2=0
+ $Y2=0
cc_99 N_A_85_345#_c_73_n N_A_210_125#_c_232_n 0.00289003f $X=2 $Y=1.685 $X2=0
+ $Y2=0
cc_100 N_A_85_345#_c_75_n N_A_210_125#_c_232_n 0.00103513f $X=2.21 $Y=0.9 $X2=0
+ $Y2=0
cc_101 N_A_85_345#_c_77_n N_A_210_125#_c_232_n 0.00190498f $X=2.107 $Y=1.685
+ $X2=0 $Y2=0
cc_102 N_A_85_345#_c_78_n N_A_210_125#_c_232_n 0.00174438f $X=2.21 $Y=1.38 $X2=0
+ $Y2=0
cc_103 N_A_85_345#_c_86_n N_A_210_125#_M1011_g 0.00758583f $X=2.105 $Y=2.27
+ $X2=0 $Y2=0
cc_104 N_A_85_345#_c_76_n N_A_210_125#_M1011_g 0.00301503f $X=2.13 $Y=1.6 $X2=0
+ $Y2=0
cc_105 N_A_85_345#_c_77_n N_A_210_125#_M1011_g 0.00270248f $X=2.107 $Y=1.685
+ $X2=0 $Y2=0
cc_106 N_A_85_345#_c_78_n N_A_210_125#_M1011_g 0.00889946f $X=2.21 $Y=1.38 $X2=0
+ $Y2=0
cc_107 N_A_85_345#_c_75_n N_A_210_125#_c_234_n 0.00651818f $X=2.21 $Y=0.9 $X2=0
+ $Y2=0
cc_108 N_A_85_345#_c_75_n N_A_210_125#_c_235_n 0.00177486f $X=2.21 $Y=0.9 $X2=0
+ $Y2=0
cc_109 N_A_85_345#_c_86_n N_A_210_125#_c_238_n 0.0108774f $X=2.105 $Y=2.27 $X2=0
+ $Y2=0
cc_110 N_A_85_345#_c_86_n N_A_210_125#_c_239_n 0.00311674f $X=2.105 $Y=2.27
+ $X2=0 $Y2=0
cc_111 N_A_85_345#_c_75_n N_B2_c_297_n 0.00134852f $X=2.21 $Y=0.9 $X2=0 $Y2=0
cc_112 N_A_85_345#_c_86_n B2 0.0026929f $X=2.105 $Y=2.27 $X2=0 $Y2=0
cc_113 N_A_85_345#_c_75_n B2 0.0351601f $X=2.21 $Y=0.9 $X2=0 $Y2=0
cc_114 N_A_85_345#_c_76_n B2 0.0106358f $X=2.13 $Y=1.6 $X2=0 $Y2=0
cc_115 N_A_85_345#_c_77_n B2 0.00919664f $X=2.107 $Y=1.685 $X2=0 $Y2=0
cc_116 N_A_85_345#_M1006_g X 0.00604901f $X=0.545 $Y=0.835 $X2=0 $Y2=0
cc_117 N_A_85_345#_M1000_g X 8.19663e-19 $X=0.61 $Y=2.885 $X2=0 $Y2=0
cc_118 N_A_85_345#_c_82_n X 0.00216294f $X=0.59 $Y=2.395 $X2=0 $Y2=0
cc_119 N_A_85_345#_M1006_g X 0.0215053f $X=0.545 $Y=0.835 $X2=0 $Y2=0
cc_120 N_A_85_345#_M1000_g X 0.00691671f $X=0.61 $Y=2.885 $X2=0 $Y2=0
cc_121 N_A_85_345#_c_83_n X 0.0429192f $X=0.59 $Y=1.89 $X2=0 $Y2=0
cc_122 N_A_85_345#_c_84_n X 0.0163879f $X=0.59 $Y=1.89 $X2=0 $Y2=0
cc_123 N_A_85_345#_c_74_n X 0.0130204f $X=0.675 $Y=1.685 $X2=0 $Y2=0
cc_124 N_A_85_345#_M1000_g N_VPWR_c_389_n 0.0116476f $X=0.61 $Y=2.885 $X2=0
+ $Y2=0
cc_125 N_A_85_345#_c_82_n N_VPWR_c_389_n 0.00146222f $X=0.59 $Y=2.395 $X2=0
+ $Y2=0
cc_126 N_A_85_345#_c_83_n N_VPWR_c_389_n 4.9066e-19 $X=0.59 $Y=1.89 $X2=0 $Y2=0
cc_127 N_A_85_345#_M1000_g N_VPWR_c_388_n 0.00947252f $X=0.61 $Y=2.885 $X2=0
+ $Y2=0
cc_128 N_A_85_345#_M1000_g N_VPWR_c_395_n 0.00486043f $X=0.61 $Y=2.885 $X2=0
+ $Y2=0
cc_129 N_A_85_345#_c_86_n N_A_479_429#_c_430_n 0.0101002f $X=2.105 $Y=2.27 $X2=0
+ $Y2=0
cc_130 N_A_85_345#_M1006_g N_VGND_c_443_n 0.00118155f $X=0.545 $Y=0.835 $X2=0
+ $Y2=0
cc_131 N_A_85_345#_c_73_n N_VGND_c_450_n 0.00321077f $X=2 $Y=1.685 $X2=0 $Y2=0
cc_132 N_A_85_345#_M1006_g N_VGND_c_447_n 0.00404248f $X=0.545 $Y=0.835 $X2=0
+ $Y2=0
cc_133 N_A_85_345#_M1006_g N_VGND_c_448_n 0.00456913f $X=0.545 $Y=0.835 $X2=0
+ $Y2=0
cc_134 N_A_85_345#_c_75_n N_VGND_c_448_n 0.00579074f $X=2.21 $Y=0.9 $X2=0 $Y2=0
cc_135 N_A1_N_M1003_g N_A2_N_M1001_g 0.0135352f $X=1.04 $Y=2.885 $X2=0 $Y2=0
cc_136 A1_N N_A2_N_M1001_g 0.0110445f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_137 N_A1_N_c_154_n N_A2_N_M1001_g 0.0174877f $X=1.065 $Y=1.32 $X2=0 $Y2=0
cc_138 N_A1_N_c_155_n N_A2_N_M1001_g 0.0160339f $X=1.065 $Y=1.155 $X2=0 $Y2=0
cc_139 N_A1_N_M1003_g A2_N 0.00895434f $X=1.04 $Y=2.885 $X2=0 $Y2=0
cc_140 N_A1_N_M1003_g N_A2_N_c_195_n 0.0865862f $X=1.04 $Y=2.885 $X2=0 $Y2=0
cc_141 A1_N N_A_210_125#_c_232_n 8.86168e-19 $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_142 A1_N N_A_210_125#_M1011_g 2.59163e-19 $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_143 N_A1_N_M1003_g N_A_210_125#_c_238_n 0.00113457f $X=1.04 $Y=2.885 $X2=0
+ $Y2=0
cc_144 N_A1_N_c_155_n N_A_210_125#_c_236_n 0.00171415f $X=1.065 $Y=1.155 $X2=0
+ $Y2=0
cc_145 A1_N X 0.0107423f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_146 N_A1_N_M1003_g N_VPWR_c_389_n 0.00997272f $X=1.04 $Y=2.885 $X2=0 $Y2=0
cc_147 N_A1_N_M1003_g N_VPWR_c_391_n 0.00486043f $X=1.04 $Y=2.885 $X2=0 $Y2=0
cc_148 N_A1_N_M1003_g N_VPWR_c_388_n 0.00818711f $X=1.04 $Y=2.885 $X2=0 $Y2=0
cc_149 A1_N N_VGND_c_443_n 0.0149235f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_150 N_A1_N_c_155_n N_VGND_c_443_n 0.00130366f $X=1.065 $Y=1.155 $X2=0 $Y2=0
cc_151 A1_N N_VGND_c_456_n 0.0490488f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_152 N_A1_N_c_154_n N_VGND_c_456_n 0.0044032f $X=1.065 $Y=1.32 $X2=0 $Y2=0
cc_153 N_A1_N_c_155_n N_VGND_c_456_n 0.0105429f $X=1.065 $Y=1.155 $X2=0 $Y2=0
cc_154 A1_N N_VGND_c_450_n 0.00592622f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_155 N_A1_N_c_155_n N_VGND_c_446_n 0.00415323f $X=1.065 $Y=1.155 $X2=0 $Y2=0
cc_156 N_A1_N_c_155_n N_VGND_c_448_n 0.00469432f $X=1.065 $Y=1.155 $X2=0 $Y2=0
cc_157 N_A2_N_M1001_g N_A_210_125#_M1011_g 0.00673677f $X=1.565 $Y=0.835 $X2=0
+ $Y2=0
cc_158 A2_N N_A_210_125#_M1011_g 0.00208365f $X=1.595 $Y=1.95 $X2=0 $Y2=0
cc_159 N_A2_N_c_195_n N_A_210_125#_M1011_g 0.00464751f $X=1.55 $Y=2.035 $X2=0
+ $Y2=0
cc_160 N_A2_N_M1001_g N_A_210_125#_c_234_n 0.00500639f $X=1.565 $Y=0.835 $X2=0
+ $Y2=0
cc_161 N_A2_N_M1001_g N_A_210_125#_c_235_n 0.0200881f $X=1.565 $Y=0.835 $X2=0
+ $Y2=0
cc_162 N_A2_N_M1007_g N_A_210_125#_c_238_n 0.00674048f $X=1.4 $Y=2.885 $X2=0
+ $Y2=0
cc_163 A2_N N_A_210_125#_c_238_n 0.0173997f $X=1.595 $Y=1.95 $X2=0 $Y2=0
cc_164 N_A2_N_c_195_n N_A_210_125#_c_238_n 8.45508e-19 $X=1.55 $Y=2.035 $X2=0
+ $Y2=0
cc_165 N_A2_N_M1007_g N_A_210_125#_c_239_n 0.00256456f $X=1.4 $Y=2.885 $X2=0
+ $Y2=0
cc_166 N_A2_N_M1001_g N_A_210_125#_c_236_n 0.0040979f $X=1.565 $Y=0.835 $X2=0
+ $Y2=0
cc_167 N_A2_N_M1007_g N_VPWR_c_389_n 0.00188275f $X=1.4 $Y=2.885 $X2=0 $Y2=0
cc_168 N_A2_N_M1007_g N_VPWR_c_391_n 0.00547815f $X=1.4 $Y=2.885 $X2=0 $Y2=0
cc_169 N_A2_N_M1007_g N_VPWR_c_388_n 0.00740955f $X=1.4 $Y=2.885 $X2=0 $Y2=0
cc_170 A2_N N_VPWR_c_388_n 0.012715f $X=1.595 $Y=1.95 $X2=0 $Y2=0
cc_171 N_A2_N_M1001_g N_VGND_c_456_n 0.0100647f $X=1.565 $Y=0.835 $X2=0 $Y2=0
cc_172 N_A_210_125#_M1011_g N_B2_M1005_g 0.0234918f $X=2.32 $Y=2.355 $X2=0 $Y2=0
cc_173 N_A_210_125#_M1002_g N_B2_c_297_n 0.0079426f $X=1.995 $Y=0.835 $X2=0
+ $Y2=0
cc_174 N_A_210_125#_c_235_n N_B2_c_297_n 6.3969e-19 $X=2.085 $Y=0.35 $X2=0 $Y2=0
cc_175 N_A_210_125#_M1011_g N_B2_c_298_n 0.0201167f $X=2.32 $Y=2.355 $X2=0 $Y2=0
cc_176 N_A_210_125#_M1002_g B2 0.00241047f $X=1.995 $Y=0.835 $X2=0 $Y2=0
cc_177 N_A_210_125#_c_231_n B2 0.0045912f $X=2.245 $Y=1.23 $X2=0 $Y2=0
cc_178 N_A_210_125#_c_235_n B2 0.0012842f $X=2.085 $Y=0.35 $X2=0 $Y2=0
cc_179 N_A_210_125#_c_231_n N_B2_c_300_n 0.0201167f $X=2.245 $Y=1.23 $X2=0 $Y2=0
cc_180 N_A_210_125#_c_238_n N_VPWR_c_389_n 0.00777152f $X=2.23 $Y=2.9 $X2=0
+ $Y2=0
cc_181 N_A_210_125#_M1011_g N_VPWR_c_390_n 0.00872446f $X=2.32 $Y=2.355 $X2=0
+ $Y2=0
cc_182 N_A_210_125#_c_238_n N_VPWR_c_390_n 0.0120931f $X=2.23 $Y=2.9 $X2=0 $Y2=0
cc_183 N_A_210_125#_c_238_n N_VPWR_c_391_n 0.052071f $X=2.23 $Y=2.9 $X2=0 $Y2=0
cc_184 N_A_210_125#_c_239_n N_VPWR_c_391_n 0.00870324f $X=2.23 $Y=2.9 $X2=0
+ $Y2=0
cc_185 N_A_210_125#_M1007_d N_VPWR_c_388_n 0.00232217f $X=1.475 $Y=2.675 $X2=0
+ $Y2=0
cc_186 N_A_210_125#_c_238_n N_VPWR_c_388_n 0.0324901f $X=2.23 $Y=2.9 $X2=0 $Y2=0
cc_187 N_A_210_125#_c_239_n N_VPWR_c_388_n 0.0111008f $X=2.23 $Y=2.9 $X2=0 $Y2=0
cc_188 N_A_210_125#_M1011_g N_A_479_429#_c_430_n 0.00130894f $X=2.32 $Y=2.355
+ $X2=0 $Y2=0
cc_189 N_A_210_125#_c_236_n N_VGND_c_443_n 0.022712f $X=1.27 $Y=0.35 $X2=0 $Y2=0
cc_190 N_A_210_125#_M1004_d N_VGND_c_456_n 0.00750174f $X=1.05 $Y=0.625 $X2=0
+ $Y2=0
cc_191 N_A_210_125#_c_234_n N_VGND_c_456_n 0.00648956f $X=2.085 $Y=0.35 $X2=0
+ $Y2=0
cc_192 N_A_210_125#_c_236_n N_VGND_c_456_n 0.0238109f $X=1.27 $Y=0.35 $X2=0
+ $Y2=0
cc_193 N_A_210_125#_c_234_n N_VGND_c_450_n 0.0090638f $X=2.085 $Y=0.35 $X2=0
+ $Y2=0
cc_194 N_A_210_125#_c_234_n N_VGND_c_446_n 0.048472f $X=2.085 $Y=0.35 $X2=0
+ $Y2=0
cc_195 N_A_210_125#_c_235_n N_VGND_c_446_n 0.00651318f $X=2.085 $Y=0.35 $X2=0
+ $Y2=0
cc_196 N_A_210_125#_c_236_n N_VGND_c_446_n 0.021319f $X=1.27 $Y=0.35 $X2=0 $Y2=0
cc_197 N_A_210_125#_c_234_n N_VGND_c_448_n 0.0289483f $X=2.085 $Y=0.35 $X2=0
+ $Y2=0
cc_198 N_A_210_125#_c_235_n N_VGND_c_448_n 0.0101042f $X=2.085 $Y=0.35 $X2=0
+ $Y2=0
cc_199 N_A_210_125#_c_236_n N_VGND_c_448_n 0.0125277f $X=1.27 $Y=0.35 $X2=0
+ $Y2=0
cc_200 N_B2_M1005_g N_B1_M1008_g 0.0192022f $X=2.75 $Y=2.355 $X2=0 $Y2=0
cc_201 N_B2_c_297_n N_B1_c_341_n 0.0173099f $X=2.77 $Y=1.155 $X2=0 $Y2=0
cc_202 B2 N_B1_c_341_n 0.00889831f $X=2.555 $Y=0.47 $X2=0 $Y2=0
cc_203 N_B2_c_298_n N_B1_c_342_n 0.0140837f $X=2.77 $Y=1.66 $X2=0 $Y2=0
cc_204 N_B2_c_302_n N_B1_c_346_n 0.0140837f $X=2.77 $Y=1.825 $X2=0 $Y2=0
cc_205 B2 N_B1_c_346_n 4.50479e-19 $X=2.555 $Y=0.47 $X2=0 $Y2=0
cc_206 B2 B1 0.0429398f $X=2.555 $Y=0.47 $X2=0 $Y2=0
cc_207 N_B2_c_300_n B1 0.00385061f $X=2.77 $Y=1.32 $X2=0 $Y2=0
cc_208 B2 N_B1_c_344_n 8.11098e-19 $X=2.555 $Y=0.47 $X2=0 $Y2=0
cc_209 N_B2_c_300_n N_B1_c_344_n 0.0140837f $X=2.77 $Y=1.32 $X2=0 $Y2=0
cc_210 N_B2_M1005_g N_VPWR_c_390_n 0.00652278f $X=2.75 $Y=2.355 $X2=0 $Y2=0
cc_211 N_B2_M1005_g N_VPWR_c_391_n 0.00336309f $X=2.75 $Y=2.355 $X2=0 $Y2=0
cc_212 N_B2_M1005_g N_VPWR_c_388_n 0.00420878f $X=2.75 $Y=2.355 $X2=0 $Y2=0
cc_213 N_B2_M1005_g N_A_479_429#_c_429_n 0.0142011f $X=2.75 $Y=2.355 $X2=0 $Y2=0
cc_214 N_B2_c_302_n N_A_479_429#_c_429_n 0.00373211f $X=2.77 $Y=1.825 $X2=0
+ $Y2=0
cc_215 B2 N_A_479_429#_c_429_n 0.0157721f $X=2.555 $Y=0.47 $X2=0 $Y2=0
cc_216 N_B2_c_302_n N_A_479_429#_c_430_n 2.60927e-19 $X=2.77 $Y=1.825 $X2=0
+ $Y2=0
cc_217 B2 N_A_479_429#_c_430_n 0.00717074f $X=2.555 $Y=0.47 $X2=0 $Y2=0
cc_218 N_B2_c_297_n N_VGND_c_445_n 3.59935e-19 $X=2.77 $Y=1.155 $X2=0 $Y2=0
cc_219 B2 N_VGND_c_445_n 0.0160467f $X=2.555 $Y=0.47 $X2=0 $Y2=0
cc_220 N_B2_c_297_n N_VGND_c_446_n 6.87871e-19 $X=2.77 $Y=1.155 $X2=0 $Y2=0
cc_221 B2 N_VGND_c_446_n 0.00893474f $X=2.555 $Y=0.47 $X2=0 $Y2=0
cc_222 B2 N_VGND_c_448_n 0.0101801f $X=2.555 $Y=0.47 $X2=0 $Y2=0
cc_223 B2 A_551_125# 0.00557666f $X=2.555 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_224 N_B1_M1008_g N_VPWR_c_390_n 0.0037594f $X=3.25 $Y=2.355 $X2=0 $Y2=0
cc_225 N_B1_M1008_g N_VPWR_c_393_n 0.00348629f $X=3.25 $Y=2.355 $X2=0 $Y2=0
cc_226 N_B1_M1008_g N_VPWR_c_388_n 0.00432409f $X=3.25 $Y=2.355 $X2=0 $Y2=0
cc_227 N_B1_M1008_g N_A_479_429#_c_429_n 0.0161576f $X=3.25 $Y=2.355 $X2=0 $Y2=0
cc_228 N_B1_c_346_n N_A_479_429#_c_429_n 0.00489473f $X=3.31 $Y=1.825 $X2=0
+ $Y2=0
cc_229 B1 N_A_479_429#_c_429_n 0.0321565f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_230 N_B1_c_341_n N_VGND_c_445_n 0.00965695f $X=3.31 $Y=1.155 $X2=0 $Y2=0
cc_231 B1 N_VGND_c_445_n 0.0156438f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_232 N_B1_c_344_n N_VGND_c_445_n 0.00438035f $X=3.31 $Y=1.32 $X2=0 $Y2=0
cc_233 N_B1_c_341_n N_VGND_c_446_n 0.00345209f $X=3.31 $Y=1.155 $X2=0 $Y2=0
cc_234 N_B1_c_341_n N_VGND_c_448_n 0.00394323f $X=3.31 $Y=1.155 $X2=0 $Y2=0
cc_235 N_X_M1000_s N_VPWR_c_388_n 0.0043444f $X=0.25 $Y=2.675 $X2=0 $Y2=0
cc_236 X N_VPWR_c_388_n 0.0121996f $X=0.155 $Y=2.69 $X2=0 $Y2=0
cc_237 X N_VPWR_c_395_n 0.0145388f $X=0.155 $Y=2.69 $X2=0 $Y2=0
cc_238 X N_VGND_c_443_n 0.0198289f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_239 X N_VGND_c_447_n 0.0096722f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_240 X N_VGND_c_448_n 0.0111021f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_241 N_VPWR_c_388_n A_223_535# 0.00308167f $X=3.6 $Y=3.33 $X2=-0.19 $Y2=-0.245
cc_242 N_VPWR_M1005_d N_A_479_429#_c_429_n 0.00256964f $X=2.825 $Y=2.145 $X2=0
+ $Y2=0
cc_243 N_VPWR_c_390_n N_A_479_429#_c_429_n 0.0186478f $X=2.985 $Y=2.44 $X2=0
+ $Y2=0
