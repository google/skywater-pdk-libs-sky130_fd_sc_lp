* NGSPICE file created from sky130_fd_sc_lp__a21bo_m.ext - technology: sky130A

.subckt sky130_fd_sc_lp__a21bo_m A1 A2 B1_N VGND VNB VPB VPWR X
M1000 a_80_72# a_196_98# VGND VNB nshort w=420000u l=150000u
+  ad=1.512e+11p pd=1.56e+06u as=3.549e+11p ps=4.21e+06u
M1001 a_196_98# B1_N VPWR VPB phighvt w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=2.352e+11p ps=2.8e+06u
M1002 VGND a_80_72# X VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1003 a_419_439# a_196_98# a_80_72# VPB phighvt w=420000u l=150000u
+  ad=2.289e+11p pd=2.77e+06u as=1.113e+11p ps=1.37e+06u
M1004 a_499_47# A1 a_80_72# VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1005 VGND A2 a_499_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_196_98# B1_N VGND VNB nshort w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1007 a_419_439# A2 VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPWR a_80_72# X VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1009 VPWR A1 a_419_439# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

