# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__decap_4
  CLASS CORE SPACER ;
  FOREIGN sky130_fd_sc_lp__decap_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  1.920000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 1.920000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 1.920000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 1.920000 0.085000 ;
      RECT 0.000000  3.245000 1.920000 3.415000 ;
      RECT 0.095000  2.105000 0.425000 3.245000 ;
      RECT 0.170000  0.085000 0.500000 1.605000 ;
      RECT 0.170000  1.605000 0.740000 1.935000 ;
      RECT 1.180000  1.340000 1.715000 1.675000 ;
      RECT 1.385000  1.675000 1.715000 3.245000 ;
      RECT 1.450000  0.085000 1.780000 1.125000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
  END
END sky130_fd_sc_lp__decap_4
END LIBRARY
