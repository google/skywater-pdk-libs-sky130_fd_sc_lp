* File: sky130_fd_sc_lp__sdfsbp_1.pex.spice
* Created: Fri Aug 28 11:29:09 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__SDFSBP_1%SCE 2 3 4 7 9 11 14 18 22 26 27 29 39 44
c93 26 0 1.26284e-19 $X=2.29 $Y=1.16
c94 22 0 5.50256e-20 $X=2.125 $Y=2.21
c95 18 0 1.81346e-19 $X=2.315 $Y=0.445
r96 37 39 38.4695 $w=3.3e-07 $l=2.2e-07 $layer=POLY_cond $X=0.72 $Y=2.08
+ $X2=0.94 $Y2=2.08
r97 35 37 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=0.51 $Y=2.08
+ $X2=0.72 $Y2=2.08
r98 33 35 38.4695 $w=3.3e-07 $l=2.2e-07 $layer=POLY_cond $X=0.29 $Y=2.08
+ $X2=0.51 $Y2=2.08
r99 29 44 10.0876 $w=3.78e-07 $l=2.15e-07 $layer=LI1_cond $X=0.72 $Y=2.105
+ $X2=0.935 $Y2=2.105
r100 29 37 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.72
+ $Y=2.08 $X2=0.72 $Y2=2.08
r101 26 27 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.29
+ $Y=1.16 $X2=2.29 $Y2=1.16
r102 24 26 44.4843 $w=2.48e-07 $l=9.65e-07 $layer=LI1_cond $X=2.25 $Y=2.125
+ $X2=2.25 $Y2=1.16
r103 22 24 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.125 $Y=2.21
+ $X2=2.25 $Y2=2.125
r104 22 44 77.6364 $w=1.68e-07 $l=1.19e-06 $layer=LI1_cond $X=2.125 $Y=2.21
+ $X2=0.935 $Y2=2.21
r105 21 27 38.9318 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.29 $Y=0.995
+ $X2=2.29 $Y2=1.16
r106 18 21 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=2.315 $Y=0.445
+ $X2=2.315 $Y2=0.995
r107 12 39 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.94 $Y=2.245
+ $X2=0.94 $Y2=2.08
r108 12 14 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.94 $Y=2.245
+ $X2=0.94 $Y2=2.725
r109 9 11 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.755 $Y=0.765
+ $X2=0.755 $Y2=0.445
r110 5 35 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.51 $Y=2.245
+ $X2=0.51 $Y2=2.08
r111 5 7 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.51 $Y=2.245
+ $X2=0.51 $Y2=2.725
r112 3 9 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.68 $Y=0.84
+ $X2=0.755 $Y2=0.765
r113 3 4 161.521 $w=1.5e-07 $l=3.15e-07 $layer=POLY_cond $X=0.68 $Y=0.84
+ $X2=0.365 $Y2=0.84
r114 2 33 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.29 $Y=1.915
+ $X2=0.29 $Y2=2.08
r115 1 4 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.29 $Y=0.915
+ $X2=0.365 $Y2=0.84
r116 1 2 512.766 $w=1.5e-07 $l=1e-06 $layer=POLY_cond $X=0.29 $Y=0.915 $X2=0.29
+ $Y2=1.915
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSBP_1%D 3 5 7 8 9 10 21 28
c44 28 0 1.89811e-19 $X=1.75 $Y=0.93
r45 25 28 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=1.545 $Y=0.93
+ $X2=1.75 $Y2=0.93
r46 21 24 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.39 $Y=1.86
+ $X2=1.39 $Y2=2.025
r47 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.39
+ $Y=1.86 $X2=1.39 $Y2=1.86
r48 10 22 3.13852 $w=7.58e-07 $l=1.95e-07 $layer=LI1_cond $X=1.51 $Y=1.665
+ $X2=1.51 $Y2=1.86
r49 9 10 5.95514 $w=7.58e-07 $l=3.7e-07 $layer=LI1_cond $X=1.51 $Y=1.295
+ $X2=1.51 $Y2=1.665
r50 8 9 5.95514 $w=7.58e-07 $l=3.7e-07 $layer=LI1_cond $X=1.51 $Y=0.925 $X2=1.51
+ $Y2=1.295
r51 8 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.75
+ $Y=0.93 $X2=1.75 $Y2=0.93
r52 5 25 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.545 $Y=0.765
+ $X2=1.545 $Y2=0.93
r53 5 7 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.545 $Y=0.765
+ $X2=1.545 $Y2=0.445
r54 3 24 358.936 $w=1.5e-07 $l=7e-07 $layer=POLY_cond $X=1.3 $Y=2.725 $X2=1.3
+ $Y2=2.025
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSBP_1%A_34_481# 1 2 9 11 15 17 18 20 23 27 33 35
c67 18 0 5.50256e-20 $X=1.185 $Y=1.29
c68 15 0 7.18248e-20 $X=1.84 $Y=2.725
r69 30 33 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=0.255 $Y=0.445
+ $X2=0.54 $Y2=0.445
r70 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.77
+ $Y=1.29 $X2=0.77 $Y2=1.29
r71 25 35 0.432806 $w=3.3e-07 $l=1.3e-07 $layer=LI1_cond $X=0.39 $Y=1.29
+ $X2=0.26 $Y2=1.29
r72 25 27 13.2706 $w=3.28e-07 $l=3.8e-07 $layer=LI1_cond $X=0.39 $Y=1.29
+ $X2=0.77 $Y2=1.29
r73 21 35 6.36606 $w=2.55e-07 $l=1.65e-07 $layer=LI1_cond $X=0.26 $Y=1.455
+ $X2=0.26 $Y2=1.29
r74 21 23 48.5356 $w=2.58e-07 $l=1.095e-06 $layer=LI1_cond $X=0.26 $Y=1.455
+ $X2=0.26 $Y2=2.55
r75 20 35 6.36606 $w=2.55e-07 $l=1.67481e-07 $layer=LI1_cond $X=0.255 $Y=1.125
+ $X2=0.26 $Y2=1.29
r76 19 30 2.36532 $w=2.5e-07 $l=1.65e-07 $layer=LI1_cond $X=0.255 $Y=0.61
+ $X2=0.255 $Y2=0.445
r77 19 20 23.7403 $w=2.48e-07 $l=5.15e-07 $layer=LI1_cond $X=0.255 $Y=0.61
+ $X2=0.255 $Y2=1.125
r78 17 28 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.11 $Y=1.29
+ $X2=0.77 $Y2=1.29
r79 17 18 13.5877 $w=2.4e-07 $l=7.5e-08 $layer=POLY_cond $X=1.11 $Y=1.29
+ $X2=1.185 $Y2=1.29
r80 13 15 651.213 $w=1.5e-07 $l=1.27e-06 $layer=POLY_cond $X=1.84 $Y=1.455
+ $X2=1.84 $Y2=2.725
r81 12 18 13.5877 $w=2.4e-07 $l=1.21861e-07 $layer=POLY_cond $X=1.26 $Y=1.38
+ $X2=1.185 $Y2=1.29
r82 11 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.765 $Y=1.38
+ $X2=1.84 $Y2=1.455
r83 11 12 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=1.765 $Y=1.38
+ $X2=1.26 $Y2=1.38
r84 7 18 12.1617 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.185 $Y=1.125
+ $X2=1.185 $Y2=1.29
r85 7 9 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=1.185 $Y=1.125
+ $X2=1.185 $Y2=0.445
r86 2 23 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.17
+ $Y=2.405 $X2=0.295 $Y2=2.55
r87 1 33 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.415
+ $Y=0.235 $X2=0.54 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSBP_1%SCD 3 6 9 11 12 13 20 21
c45 11 0 7.18248e-20 $X=2.64 $Y=1.295
r46 18 21 17.4861 $w=3.3e-07 $l=1e-07 $layer=POLY_cond $X=2.64 $Y=2.04 $X2=2.74
+ $Y2=2.04
r47 18 20 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.64 $Y=2.04
+ $X2=2.475 $Y2=2.04
r48 13 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.64
+ $Y=2.04 $X2=2.64 $Y2=2.04
r49 12 13 21.5981 $w=1.88e-07 $l=3.7e-07 $layer=LI1_cond $X=2.64 $Y=1.665
+ $X2=2.64 $Y2=2.035
r50 11 12 21.5981 $w=1.88e-07 $l=3.7e-07 $layer=LI1_cond $X=2.64 $Y=1.295
+ $X2=2.64 $Y2=1.665
r51 7 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.74 $Y=1.875
+ $X2=2.74 $Y2=2.04
r52 7 9 733.255 $w=1.5e-07 $l=1.43e-06 $layer=POLY_cond $X=2.74 $Y=1.875
+ $X2=2.74 $Y2=0.445
r53 6 20 102.553 $w=1.5e-07 $l=2e-07 $layer=POLY_cond $X=2.275 $Y=2.13 $X2=2.475
+ $Y2=2.13
r54 1 6 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.2 $Y=2.205
+ $X2=2.275 $Y2=2.13
r55 1 3 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=2.2 $Y=2.205 $X2=2.2
+ $Y2=2.725
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSBP_1%CLK 1 3 7 9 10 11
c40 7 0 3.14497e-19 $X=3.17 $Y=0.445
r41 16 17 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.44
+ $Y=1.005 $X2=3.44 $Y2=1.005
r42 10 11 9.21977 $w=4.78e-07 $l=3.7e-07 $layer=LI1_cond $X=3.515 $Y=1.295
+ $X2=3.515 $Y2=1.665
r43 10 17 7.22631 $w=4.78e-07 $l=2.9e-07 $layer=LI1_cond $X=3.515 $Y=1.295
+ $X2=3.515 $Y2=1.005
r44 9 17 1.99346 $w=4.78e-07 $l=8e-08 $layer=LI1_cond $X=3.515 $Y=0.925
+ $X2=3.515 $Y2=1.005
r45 5 16 40.728 $w=4.52e-07 $l=2.30499e-07 $layer=POLY_cond $X=3.17 $Y=0.84
+ $X2=3.327 $Y2=1.005
r46 5 7 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=3.17 $Y=0.84 $X2=3.17
+ $Y2=0.445
r47 1 16 92.9802 $w=4.52e-07 $l=7.49223e-07 $layer=POLY_cond $X=3.125 $Y=1.66
+ $X2=3.327 $Y2=1.005
r48 1 3 546.096 $w=1.5e-07 $l=1.065e-06 $layer=POLY_cond $X=3.125 $Y=1.66
+ $X2=3.125 $Y2=2.725
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSBP_1%A_901_441# 1 2 9 13 15 17 20 23 24 25 26 27
+ 30 34 36 39 40 41 43 44 46 50 53
c163 46 0 1.3719e-19 $X=9.625 $Y=1.515
c164 41 0 1.71354e-19 $X=7.985 $Y=1.865
c165 40 0 5.23886e-20 $X=8.955 $Y=1.865
c166 26 0 2.67723e-19 $X=9.6 $Y=1.515
c167 24 0 1.21539e-20 $X=5.655 $Y=1.71
c168 20 0 1.15797e-19 $X=10.05 $Y=2.65
r169 56 57 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.06
+ $Y=1.54 $X2=6.06 $Y2=1.54
r170 53 56 3.54598 $w=2.58e-07 $l=8e-08 $layer=LI1_cond $X=6.095 $Y=1.46
+ $X2=6.095 $Y2=1.54
r171 50 52 6.40426 $w=6.23e-07 $l=1.65e-07 $layer=LI1_cond $X=4.792 $Y=1.54
+ $X2=4.792 $Y2=1.375
r172 50 51 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.01
+ $Y=1.54 $X2=5.01 $Y2=1.54
r173 46 47 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.625
+ $Y=1.515 $X2=9.625 $Y2=1.515
r174 44 46 29.1866 $w=1.88e-07 $l=5e-07 $layer=LI1_cond $X=9.125 $Y=1.515
+ $X2=9.625 $Y2=1.515
r175 42 44 6.84389 $w=1.9e-07 $l=1.30767e-07 $layer=LI1_cond $X=9.04 $Y=1.61
+ $X2=9.125 $Y2=1.515
r176 42 43 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=9.04 $Y=1.61
+ $X2=9.04 $Y2=1.78
r177 40 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.955 $Y=1.865
+ $X2=9.04 $Y2=1.78
r178 40 41 63.2834 $w=1.68e-07 $l=9.7e-07 $layer=LI1_cond $X=8.955 $Y=1.865
+ $X2=7.985 $Y2=1.865
r179 39 41 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.9 $Y=1.78
+ $X2=7.985 $Y2=1.865
r180 38 39 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=7.9 $Y=1.545
+ $X2=7.9 $Y2=1.78
r181 37 53 3.22376 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=6.225 $Y=1.46
+ $X2=6.095 $Y2=1.46
r182 36 38 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.815 $Y=1.46
+ $X2=7.9 $Y2=1.545
r183 36 37 103.733 $w=1.68e-07 $l=1.59e-06 $layer=LI1_cond $X=7.815 $Y=1.46
+ $X2=6.225 $Y2=1.46
r184 34 52 31.116 $w=2.98e-07 $l=8.1e-07 $layer=LI1_cond $X=4.855 $Y=0.565
+ $X2=4.855 $Y2=1.375
r185 28 50 2.81318 $w=6.23e-07 $l=1.47e-07 $layer=LI1_cond $X=4.792 $Y=1.687
+ $X2=4.792 $Y2=1.54
r186 28 30 12.688 $w=6.23e-07 $l=6.63e-07 $layer=LI1_cond $X=4.792 $Y=1.687
+ $X2=4.792 $Y2=2.35
r187 27 47 61.2015 $w=3.3e-07 $l=3.5e-07 $layer=POLY_cond $X=9.975 $Y=1.515
+ $X2=9.625 $Y2=1.515
r188 26 47 4.37153 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=9.6 $Y=1.515
+ $X2=9.625 $Y2=1.515
r189 25 57 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=6.075 $Y=1.54
+ $X2=6.06 $Y2=1.54
r190 23 51 45.5174 $w=6.7e-07 $l=5.7e-07 $layer=POLY_cond $X=5.58 $Y=1.71
+ $X2=5.01 $Y2=1.71
r191 23 24 6.88608 $w=5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.58 $Y=1.71
+ $X2=5.655 $Y2=1.71
r192 22 57 57.7042 $w=3.3e-07 $l=3.3e-07 $layer=POLY_cond $X=5.73 $Y=1.54
+ $X2=6.06 $Y2=1.54
r193 22 24 6.88608 $w=5e-07 $l=2.04083e-07 $layer=POLY_cond $X=5.73 $Y=1.54
+ $X2=5.655 $Y2=1.71
r194 18 27 28.7299 $w=2.68e-07 $l=1.98997e-07 $layer=POLY_cond $X=10.05 $Y=1.68
+ $X2=9.975 $Y2=1.515
r195 18 20 497.383 $w=1.5e-07 $l=9.7e-07 $layer=POLY_cond $X=10.05 $Y=1.68
+ $X2=10.05 $Y2=2.65
r196 15 26 32.1775 $w=3.3e-07 $l=1.98997e-07 $layer=POLY_cond $X=9.525 $Y=1.35
+ $X2=9.6 $Y2=1.515
r197 15 17 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=9.525 $Y=1.35
+ $X2=9.525 $Y2=0.915
r198 11 25 32.1775 $w=3.3e-07 $l=1.98997e-07 $layer=POLY_cond $X=6.15 $Y=1.375
+ $X2=6.075 $Y2=1.54
r199 11 13 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=6.15 $Y=1.375
+ $X2=6.15 $Y2=0.805
r200 7 24 23.237 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=5.655 $Y=2.045
+ $X2=5.655 $Y2=1.71
r201 7 9 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=5.655 $Y=2.045
+ $X2=5.655 $Y2=2.525
r202 2 30 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=4.505
+ $Y=2.205 $X2=4.645 $Y2=2.35
r203 1 34 182 $w=1.7e-07 $l=2.60768e-07 $layer=licon1_NDIFF $count=1 $X=4.7
+ $Y=0.365 $X2=4.84 $Y2=0.565
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSBP_1%A_1274_401# 1 2 9 13 15 20 24 25 27 28 29
+ 31 32 33 35 41
c130 33 0 1.93097e-19 $X=9.475 $Y=1.865
c131 24 0 1.15797e-19 $X=9.305 $Y=2.385
r132 40 41 10.4086 $w=3.01e-07 $l=6.5e-08 $layer=POLY_cond $X=6.445 $Y=1.99
+ $X2=6.51 $Y2=1.99
r133 34 35 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=10.045 $Y=1.25
+ $X2=10.045 $Y2=1.78
r134 32 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.96 $Y=1.865
+ $X2=10.045 $Y2=1.78
r135 32 33 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=9.96 $Y=1.865
+ $X2=9.475 $Y2=1.865
r136 30 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.39 $Y=1.95
+ $X2=9.475 $Y2=1.865
r137 30 31 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=9.39 $Y=1.95
+ $X2=9.39 $Y2=2.3
r138 28 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.96 $Y=1.165
+ $X2=10.045 $Y2=1.25
r139 28 29 83.1818 $w=1.68e-07 $l=1.275e-06 $layer=LI1_cond $X=9.96 $Y=1.165
+ $X2=8.685 $Y2=1.165
r140 27 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.6 $Y=1.08
+ $X2=8.685 $Y2=1.165
r141 26 27 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=8.6 $Y=0.855
+ $X2=8.6 $Y2=1.08
r142 25 39 5.32087 $w=3.21e-07 $l=1.4e-07 $layer=LI1_cond $X=7.327 $Y=2.385
+ $X2=7.327 $Y2=2.525
r143 24 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.305 $Y=2.385
+ $X2=9.39 $Y2=2.3
r144 24 25 119.064 $w=1.68e-07 $l=1.825e-06 $layer=LI1_cond $X=9.305 $Y=2.385
+ $X2=7.48 $Y2=2.385
r145 20 26 6.96323 $w=2.2e-07 $l=1.46458e-07 $layer=LI1_cond $X=8.515 $Y=0.745
+ $X2=8.6 $Y2=0.855
r146 20 22 48.7169 $w=2.18e-07 $l=9.3e-07 $layer=LI1_cond $X=8.515 $Y=0.745
+ $X2=7.585 $Y2=0.745
r147 18 41 17.6146 $w=3.01e-07 $l=1.1e-07 $layer=POLY_cond $X=6.62 $Y=1.99
+ $X2=6.51 $Y2=1.99
r148 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.62
+ $Y=1.99 $X2=6.62 $Y2=1.99
r149 15 25 12.8461 $w=3.21e-07 $l=4.72313e-07 $layer=LI1_cond $X=7.005 $Y=2.047
+ $X2=7.327 $Y2=2.385
r150 15 17 15.5681 $w=2.83e-07 $l=3.85e-07 $layer=LI1_cond $X=7.005 $Y=2.047
+ $X2=6.62 $Y2=2.047
r151 11 41 19.0468 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.51 $Y=1.825
+ $X2=6.51 $Y2=1.99
r152 11 13 523.021 $w=1.5e-07 $l=1.02e-06 $layer=POLY_cond $X=6.51 $Y=1.825
+ $X2=6.51 $Y2=0.805
r153 7 40 19.0468 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.445 $Y=2.155
+ $X2=6.445 $Y2=1.99
r154 7 9 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=6.445 $Y=2.155
+ $X2=6.445 $Y2=2.525
r155 2 39 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=7.175
+ $Y=2.315 $X2=7.315 $Y2=2.525
r156 1 22 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=7.46
+ $Y=0.595 $X2=7.585 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSBP_1%A_1146_463# 1 2 9 11 13 15 16 18 20 22 24
+ 26 31 35 37 38 41 42 44 47 48 50 55 56 57
c140 50 0 7.46252e-20 $X=8.61 $Y=1.515
c141 35 0 2.20475e-19 $X=5.935 $Y=0.805
r142 55 56 8.71257 $w=2.88e-07 $l=1.7e-07 $layer=LI1_cond $X=5.83 $Y=1.885
+ $X2=5.83 $Y2=2.055
r143 50 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.61
+ $Y=1.515 $X2=8.61 $Y2=1.515
r144 48 50 16.0526 $w=1.88e-07 $l=2.75e-07 $layer=LI1_cond $X=8.335 $Y=1.515
+ $X2=8.61 $Y2=1.515
r145 47 48 6.84389 $w=1.9e-07 $l=1.30767e-07 $layer=LI1_cond $X=8.25 $Y=1.42
+ $X2=8.335 $Y2=1.515
r146 46 47 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=8.25 $Y=1.205
+ $X2=8.25 $Y2=1.42
r147 45 57 5.40251 $w=1.8e-07 $l=9.5e-08 $layer=LI1_cond $X=7.25 $Y=1.115
+ $X2=7.155 $Y2=1.115
r148 44 46 6.82373 $w=1.8e-07 $l=1.25499e-07 $layer=LI1_cond $X=8.165 $Y=1.115
+ $X2=8.25 $Y2=1.205
r149 44 45 56.3788 $w=1.78e-07 $l=9.15e-07 $layer=LI1_cond $X=8.165 $Y=1.115
+ $X2=7.25 $Y2=1.115
r150 41 42 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.155
+ $Y=0.69 $X2=7.155 $Y2=0.69
r151 39 57 1.14861 $w=1.9e-07 $l=9e-08 $layer=LI1_cond $X=7.155 $Y=1.025
+ $X2=7.155 $Y2=1.115
r152 39 41 19.555 $w=1.88e-07 $l=3.35e-07 $layer=LI1_cond $X=7.155 $Y=1.025
+ $X2=7.155 $Y2=0.69
r153 37 57 5.40251 $w=1.8e-07 $l=9.5e-08 $layer=LI1_cond $X=7.06 $Y=1.115
+ $X2=7.155 $Y2=1.115
r154 37 38 59.1515 $w=1.78e-07 $l=9.6e-07 $layer=LI1_cond $X=7.06 $Y=1.115
+ $X2=6.1 $Y2=1.115
r155 33 38 8.81111 $w=1.8e-07 $l=1.3e-07 $layer=LI1_cond $X=5.97 $Y=1.115
+ $X2=6.1 $Y2=1.115
r156 33 53 18.1257 $w=1.75e-07 $l=2.6e-07 $layer=LI1_cond $X=5.97 $Y=1.115
+ $X2=5.71 $Y2=1.115
r157 33 35 9.75144 $w=2.58e-07 $l=2.2e-07 $layer=LI1_cond $X=5.97 $Y=1.025
+ $X2=5.97 $Y2=0.805
r158 31 56 18.6775 $w=2.88e-07 $l=4.7e-07 $layer=LI1_cond $X=5.89 $Y=2.525
+ $X2=5.89 $Y2=2.055
r159 27 53 0.89264 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=5.71 $Y=1.205 $X2=5.71
+ $Y2=1.115
r160 27 55 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=5.71 $Y=1.205
+ $X2=5.71 $Y2=1.885
r161 26 51 57.7042 $w=3.3e-07 $l=3.3e-07 $layer=POLY_cond $X=8.94 $Y=1.515
+ $X2=8.61 $Y2=1.515
r162 23 42 76.0647 $w=3.3e-07 $l=4.35e-07 $layer=POLY_cond $X=7.155 $Y=1.125
+ $X2=7.155 $Y2=0.69
r163 23 24 13.5877 $w=2.4e-07 $l=7.5e-08 $layer=POLY_cond $X=7.155 $Y=1.125
+ $X2=7.155 $Y2=1.2
r164 20 26 41.2111 $w=2.18e-07 $l=1.98997e-07 $layer=POLY_cond $X=9.165 $Y=1.35
+ $X2=9.09 $Y2=1.515
r165 20 22 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=9.165 $Y=1.35
+ $X2=9.165 $Y2=0.915
r166 16 26 41.2111 $w=2.18e-07 $l=1.98997e-07 $layer=POLY_cond $X=9.015 $Y=1.68
+ $X2=9.09 $Y2=1.515
r167 16 18 325.606 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=9.015 $Y=1.68
+ $X2=9.015 $Y2=2.315
r168 13 15 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=7.8 $Y=1.125
+ $X2=7.8 $Y2=0.805
r169 12 24 12.1617 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.32 $Y=1.2
+ $X2=7.155 $Y2=1.2
r170 11 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.725 $Y=1.2
+ $X2=7.8 $Y2=1.125
r171 11 12 207.67 $w=1.5e-07 $l=4.05e-07 $layer=POLY_cond $X=7.725 $Y=1.2
+ $X2=7.32 $Y2=1.2
r172 7 24 13.5877 $w=2.4e-07 $l=9.87421e-08 $layer=POLY_cond $X=7.1 $Y=1.275
+ $X2=7.155 $Y2=1.2
r173 7 9 640.957 $w=1.5e-07 $l=1.25e-06 $layer=POLY_cond $X=7.1 $Y=1.275 $X2=7.1
+ $Y2=2.525
r174 2 31 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=5.73
+ $Y=2.315 $X2=5.87 $Y2=2.525
r175 1 35 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=5.795
+ $Y=0.595 $X2=5.935 $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSBP_1%SET_B 1 3 5 9 13 15 16 19 23 24 27 29 35 36
+ 37
r117 36 43 29.8398 $w=2.08e-07 $l=5.65e-07 $layer=LI1_cond $X=11.365 $Y=2.025
+ $X2=10.8 $Y2=2.025
r118 35 38 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=11.365 $Y=2.035
+ $X2=11.365 $Y2=2.2
r119 35 37 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=11.365 $Y=2.035
+ $X2=11.365 $Y2=1.87
r120 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.365
+ $Y=2.035 $X2=11.365 $Y2=2.035
r121 29 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=2.035
+ $X2=10.8 $Y2=2.035
r122 27 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.55
+ $Y=1.955 $X2=7.55 $Y2=1.955
r123 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=2.035
+ $X2=7.44 $Y2=2.035
r124 24 26 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.585 $Y=2.035
+ $X2=7.44 $Y2=2.035
r125 23 29 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=10.655 $Y=2.035
+ $X2=10.8 $Y2=2.035
r126 23 24 3.7995 $w=1.4e-07 $l=3.07e-06 $layer=MET1_cond $X=10.655 $Y=2.035
+ $X2=7.585 $Y2=2.035
r127 21 37 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=11.305 $Y=1.29
+ $X2=11.305 $Y2=1.87
r128 19 38 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=11.275 $Y=2.65
+ $X2=11.275 $Y2=2.2
r129 15 21 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=11.23 $Y=1.215
+ $X2=11.305 $Y2=1.29
r130 15 16 197.415 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=11.23 $Y=1.215
+ $X2=10.845 $Y2=1.215
r131 11 16 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=10.77 $Y=1.14
+ $X2=10.845 $Y2=1.215
r132 11 13 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=10.77 $Y=1.14
+ $X2=10.77 $Y2=0.8
r133 7 9 505.074 $w=1.5e-07 $l=9.85e-07 $layer=POLY_cond $X=8.16 $Y=1.79
+ $X2=8.16 $Y2=0.805
r134 6 32 11.4178 $w=3.3e-07 $l=1.1e-07 $layer=POLY_cond $X=7.605 $Y=1.955
+ $X2=7.495 $Y2=1.955
r135 5 7 32.1775 $w=3.3e-07 $l=1.98997e-07 $layer=POLY_cond $X=8.085 $Y=1.955
+ $X2=8.16 $Y2=1.79
r136 5 6 83.9334 $w=3.3e-07 $l=4.8e-07 $layer=POLY_cond $X=8.085 $Y=1.955
+ $X2=7.605 $Y2=1.955
r137 1 32 20.7597 $w=1.5e-07 $l=1.81659e-07 $layer=POLY_cond $X=7.53 $Y=2.12
+ $X2=7.495 $Y2=1.955
r138 1 3 207.67 $w=1.5e-07 $l=4.05e-07 $layer=POLY_cond $X=7.53 $Y=2.12 $X2=7.53
+ $Y2=2.525
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSBP_1%A_640_481# 1 2 7 8 12 13 14 18 19 20 23 25
+ 29 31 35 39 45 47 48 51 53 57 58 62 63
c136 53 0 1.60744e-19 $X=3.925 $Y=0.495
c137 35 0 1.89578e-19 $X=9.525 $Y=2.44
c138 23 0 1.58686e-19 $X=5.72 $Y=0.805
r139 62 63 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.04
+ $Y=1.06 $X2=4.04 $Y2=1.06
r140 60 62 64.8818 $w=1.98e-07 $l=1.17e-06 $layer=LI1_cond $X=4.025 $Y=2.23
+ $X2=4.025 $Y2=1.06
r141 59 62 22.1818 $w=1.98e-07 $l=4e-07 $layer=LI1_cond $X=4.025 $Y=0.66
+ $X2=4.025 $Y2=1.06
r142 57 60 6.81784 $w=2.05e-07 $l=1.43541e-07 $layer=LI1_cond $X=3.925 $Y=2.332
+ $X2=4.025 $Y2=2.23
r143 57 58 26.51 $w=2.03e-07 $l=4.9e-07 $layer=LI1_cond $X=3.925 $Y=2.332
+ $X2=3.435 $Y2=2.332
r144 53 59 7.36389 $w=3.3e-07 $l=2.09105e-07 $layer=LI1_cond $X=3.925 $Y=0.495
+ $X2=4.025 $Y2=0.66
r145 53 55 18.8582 $w=3.28e-07 $l=5.4e-07 $layer=LI1_cond $X=3.925 $Y=0.495
+ $X2=3.385 $Y2=0.495
r146 49 58 6.82929 $w=2.05e-07 $l=1.42808e-07 $layer=LI1_cond $X=3.34 $Y=2.435
+ $X2=3.435 $Y2=2.332
r147 49 51 7.29665 $w=1.88e-07 $l=1.25e-07 $layer=LI1_cond $X=3.34 $Y=2.435
+ $X2=3.34 $Y2=2.56
r148 43 63 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=4.04 $Y=1.415
+ $X2=4.04 $Y2=1.06
r149 43 45 199.979 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=4.04 $Y=1.49
+ $X2=4.43 $Y2=1.49
r150 41 63 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=4.04 $Y=1.045
+ $X2=4.04 $Y2=1.06
r151 37 39 279.457 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=10.05 $Y=0.255
+ $X2=10.05 $Y2=0.8
r152 33 35 325.606 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=9.525 $Y=3.075
+ $X2=9.525 $Y2=2.44
r153 32 48 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.16 $Y=3.15
+ $X2=6.085 $Y2=3.15
r154 31 33 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.45 $Y=3.15
+ $X2=9.525 $Y2=3.075
r155 31 32 1687 $w=1.5e-07 $l=3.29e-06 $layer=POLY_cond $X=9.45 $Y=3.15 $X2=6.16
+ $Y2=3.15
r156 27 48 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.085 $Y=3.075
+ $X2=6.085 $Y2=3.15
r157 27 29 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=6.085 $Y=3.075
+ $X2=6.085 $Y2=2.525
r158 26 47 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.795 $Y=0.18
+ $X2=5.72 $Y2=0.18
r159 25 37 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.975 $Y=0.18
+ $X2=10.05 $Y2=0.255
r160 25 26 2143.36 $w=1.5e-07 $l=4.18e-06 $layer=POLY_cond $X=9.975 $Y=0.18
+ $X2=5.795 $Y2=0.18
r161 21 47 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.72 $Y=0.255
+ $X2=5.72 $Y2=0.18
r162 21 23 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=5.72 $Y=0.255
+ $X2=5.72 $Y2=0.805
r163 19 47 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.645 $Y=0.18
+ $X2=5.72 $Y2=0.18
r164 19 20 484.564 $w=1.5e-07 $l=9.45e-07 $layer=POLY_cond $X=5.645 $Y=0.18
+ $X2=4.7 $Y2=0.18
r165 16 18 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=4.625 $Y=0.895
+ $X2=4.625 $Y2=0.575
r166 15 20 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.625 $Y=0.255
+ $X2=4.7 $Y2=0.18
r167 15 18 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=4.625 $Y=0.255
+ $X2=4.625 $Y2=0.575
r168 13 48 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.01 $Y=3.15
+ $X2=6.085 $Y2=3.15
r169 13 14 771.713 $w=1.5e-07 $l=1.505e-06 $layer=POLY_cond $X=6.01 $Y=3.15
+ $X2=4.505 $Y2=3.15
r170 10 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.43 $Y=3.075
+ $X2=4.505 $Y2=3.15
r171 10 12 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=4.43 $Y=3.075
+ $X2=4.43 $Y2=2.525
r172 9 45 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.43 $Y=1.565
+ $X2=4.43 $Y2=1.49
r173 9 12 492.255 $w=1.5e-07 $l=9.6e-07 $layer=POLY_cond $X=4.43 $Y=1.565
+ $X2=4.43 $Y2=2.525
r174 8 41 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=4.205 $Y=0.97
+ $X2=4.04 $Y2=1.045
r175 7 16 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.55 $Y=0.97
+ $X2=4.625 $Y2=0.895
r176 7 8 176.904 $w=1.5e-07 $l=3.45e-07 $layer=POLY_cond $X=4.55 $Y=0.97
+ $X2=4.205 $Y2=0.97
r177 2 51 600 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_PDIFF $count=1 $X=3.2
+ $Y=2.405 $X2=3.34 $Y2=2.56
r178 1 55 182 $w=1.7e-07 $l=3.2249e-07 $layer=licon1_NDIFF $count=1 $X=3.245
+ $Y=0.235 $X2=3.385 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSBP_1%A_2067_92# 1 2 9 13 16 17 20 24 27 29 34
c80 29 0 6.55926e-20 $X=12.062 $Y=1.622
c81 20 0 1.86545e-20 $X=10.825 $Y=1.665
r82 31 34 5.0366 $w=2.68e-07 $l=1.18e-07 $layer=LI1_cond $X=12.062 $Y=2.6
+ $X2=12.18 $Y2=2.6
r83 27 31 3.29739 $w=1.75e-07 $l=1.35e-07 $layer=LI1_cond $X=12.062 $Y=2.465
+ $X2=12.062 $Y2=2.6
r84 26 29 2.96557 $w=1.75e-07 $l=1.28e-07 $layer=LI1_cond $X=12.062 $Y=1.75
+ $X2=12.062 $Y2=1.622
r85 26 27 45.3143 $w=1.73e-07 $l=7.15e-07 $layer=LI1_cond $X=12.062 $Y=1.75
+ $X2=12.062 $Y2=2.465
r86 22 29 23.0489 $w=2.53e-07 $l=5.1e-07 $layer=LI1_cond $X=11.552 $Y=1.622
+ $X2=12.062 $Y2=1.622
r87 22 24 17.3678 $w=3.53e-07 $l=5.35e-07 $layer=LI1_cond $X=11.552 $Y=1.495
+ $X2=11.552 $Y2=0.96
r88 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.825
+ $Y=1.665 $X2=10.825 $Y2=1.665
r89 17 22 7.99931 $w=2.53e-07 $l=1.77e-07 $layer=LI1_cond $X=11.375 $Y=1.622
+ $X2=11.552 $Y2=1.622
r90 17 19 24.8566 $w=2.53e-07 $l=5.5e-07 $layer=LI1_cond $X=11.375 $Y=1.622
+ $X2=10.825 $Y2=1.622
r91 15 20 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=10.485 $Y=1.665
+ $X2=10.825 $Y2=1.665
r92 15 16 5.03009 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=10.485 $Y=1.665
+ $X2=10.41 $Y2=1.665
r93 11 16 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.41 $Y=1.83
+ $X2=10.41 $Y2=1.665
r94 11 13 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=10.41 $Y=1.83
+ $X2=10.41 $Y2=2.65
r95 7 16 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.41 $Y=1.5
+ $X2=10.41 $Y2=1.665
r96 7 9 358.936 $w=1.5e-07 $l=7e-07 $layer=POLY_cond $X=10.41 $Y=1.5 $X2=10.41
+ $Y2=0.8
r97 2 34 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=12.055
+ $Y=2.42 $X2=12.18 $Y2=2.63
r98 1 24 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=11.475
+ $Y=0.75 $X2=11.6 $Y2=0.96
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSBP_1%A_1920_119# 1 2 3 12 14 15 18 20 25 26 27
+ 28 30 33 37 40 42 47 48 49 53 54 55 56 57 59 60 61 62 66 67 76 81 82 89 97
c205 81 0 5.14661e-20 $X=13.57 $Y=0.415
c206 76 0 6.55926e-20 $X=12.5 $Y=1.755
c207 60 0 1.66769e-19 $X=13.405 $Y=0.535
r208 87 89 12.5444 $w=3.45e-07 $l=7.5e-08 $layer=POLY_cond $X=12.492 $Y=1.975
+ $X2=12.492 $Y2=2.05
r209 84 85 8.03218 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=13.57 $Y=0.535
+ $X2=13.57 $Y2=0.765
r210 82 94 32.3493 $w=3.3e-07 $l=1.85e-07 $layer=POLY_cond $X=13.57 $Y=0.415
+ $X2=13.57 $Y2=0.6
r211 81 84 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=13.57 $Y=0.415
+ $X2=13.57 $Y2=0.535
r212 81 82 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=13.57
+ $Y=0.415 $X2=13.57 $Y2=0.415
r213 79 91 46.3655 $w=3.45e-07 $l=1.65e-07 $layer=POLY_cond $X=12.492 $Y=2.095
+ $X2=12.492 $Y2=2.26
r214 79 89 7.52664 $w=3.45e-07 $l=4.5e-08 $layer=POLY_cond $X=12.492 $Y=2.095
+ $X2=12.492 $Y2=2.05
r215 78 79 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=12.5
+ $Y=2.095 $X2=12.5 $Y2=2.095
r216 76 87 36.7969 $w=3.45e-07 $l=2.2e-07 $layer=POLY_cond $X=12.492 $Y=1.755
+ $X2=12.492 $Y2=1.975
r217 75 78 9.57968 $w=4.33e-07 $l=3.4e-07 $layer=LI1_cond $X=12.557 $Y=1.755
+ $X2=12.557 $Y2=2.095
r218 75 76 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=12.5
+ $Y=1.755 $X2=12.5 $Y2=1.755
r219 70 72 1.02178 $w=5.97e-07 $l=5e-08 $layer=LI1_cond $X=9.74 $Y=2.5 $X2=9.79
+ $Y2=2.5
r220 67 98 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=14.772 $Y=1.505
+ $X2=14.772 $Y2=1.67
r221 67 97 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=14.772 $Y=1.505
+ $X2=14.772 $Y2=1.34
r222 66 67 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=14.75
+ $Y=1.505 $X2=14.75 $Y2=1.505
r223 64 66 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=14.75 $Y=0.85
+ $X2=14.75 $Y2=1.505
r224 63 85 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.735 $Y=0.765
+ $X2=13.57 $Y2=0.765
r225 62 64 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=14.665 $Y=0.765
+ $X2=14.75 $Y2=0.85
r226 62 63 60.6738 $w=1.68e-07 $l=9.3e-07 $layer=LI1_cond $X=14.665 $Y=0.765
+ $X2=13.735 $Y2=0.765
r227 60 84 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.405 $Y=0.535
+ $X2=13.57 $Y2=0.535
r228 60 61 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=13.405 $Y=0.535
+ $X2=12.795 $Y2=0.535
r229 59 75 9.31566 $w=4.33e-07 $l=2.29063e-07 $layer=LI1_cond $X=12.71 $Y=1.59
+ $X2=12.557 $Y2=1.755
r230 58 61 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=12.71 $Y=0.62
+ $X2=12.795 $Y2=0.535
r231 58 59 63.2834 $w=1.68e-07 $l=9.7e-07 $layer=LI1_cond $X=12.71 $Y=0.62
+ $X2=12.71 $Y2=1.59
r232 56 78 9.31566 $w=4.33e-07 $l=1.85257e-07 $layer=LI1_cond $X=12.6 $Y=2.26
+ $X2=12.557 $Y2=2.095
r233 56 57 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=12.6 $Y=2.26
+ $X2=12.6 $Y2=2.905
r234 54 57 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=12.515 $Y=2.99
+ $X2=12.6 $Y2=2.905
r235 54 55 56.107 $w=1.68e-07 $l=8.6e-07 $layer=LI1_cond $X=12.515 $Y=2.99
+ $X2=11.655 $Y2=2.99
r236 51 55 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=11.525 $Y=2.905
+ $X2=11.655 $Y2=2.99
r237 51 53 11.0812 $w=2.58e-07 $l=2.5e-07 $layer=LI1_cond $X=11.525 $Y=2.905
+ $X2=11.525 $Y2=2.655
r238 50 53 8.20008 $w=2.58e-07 $l=1.85e-07 $layer=LI1_cond $X=11.525 $Y=2.47
+ $X2=11.525 $Y2=2.655
r239 48 50 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=11.395 $Y=2.385
+ $X2=11.525 $Y2=2.47
r240 48 49 59.6952 $w=1.68e-07 $l=9.15e-07 $layer=LI1_cond $X=11.395 $Y=2.385
+ $X2=10.48 $Y2=2.385
r241 47 49 8.70441 $w=5.97e-07 $l=3.04549e-07 $layer=LI1_cond $X=10.395 $Y=2.12
+ $X2=10.48 $Y2=2.385
r242 47 72 12.3635 $w=5.97e-07 $l=7.71962e-07 $layer=LI1_cond $X=10.395 $Y=2.12
+ $X2=9.79 $Y2=2.5
r243 46 47 78.9412 $w=1.68e-07 $l=1.21e-06 $layer=LI1_cond $X=10.395 $Y=0.91
+ $X2=10.395 $Y2=2.12
r244 42 46 7.28469 $w=2.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=10.31 $Y=0.775
+ $X2=10.395 $Y2=0.91
r245 42 44 24.3294 $w=2.68e-07 $l=5.7e-07 $layer=LI1_cond $X=10.31 $Y=0.775
+ $X2=9.74 $Y2=0.775
r246 39 76 2.50888 $w=3.45e-07 $l=1.5e-08 $layer=POLY_cond $X=12.492 $Y=1.74
+ $X2=12.492 $Y2=1.755
r247 39 40 175.879 $w=1.5e-07 $l=3.43e-07 $layer=POLY_cond $X=12.492 $Y=1.665
+ $X2=12.835 $Y2=1.665
r248 37 97 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=14.885 $Y=0.81
+ $X2=14.885 $Y2=1.34
r249 33 98 407.649 $w=1.5e-07 $l=7.95e-07 $layer=POLY_cond $X=14.725 $Y=2.465
+ $X2=14.725 $Y2=1.67
r250 28 30 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=13.165 $Y=2.125
+ $X2=13.165 $Y2=2.52
r251 26 94 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=13.405 $Y=0.6
+ $X2=13.57 $Y2=0.6
r252 26 27 253.819 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=13.405 $Y=0.6
+ $X2=12.91 $Y2=0.6
r253 23 40 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=12.835 $Y=1.59
+ $X2=12.835 $Y2=1.665
r254 23 25 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=12.835 $Y=1.59
+ $X2=12.835 $Y2=0.96
r255 22 27 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=12.835 $Y=0.675
+ $X2=12.91 $Y2=0.6
r256 22 25 146.138 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=12.835 $Y=0.675
+ $X2=12.835 $Y2=0.96
r257 21 89 22.2839 $w=1.5e-07 $l=1.73e-07 $layer=POLY_cond $X=12.665 $Y=2.05
+ $X2=12.492 $Y2=2.05
r258 20 28 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=13.09 $Y=2.05
+ $X2=13.165 $Y2=2.125
r259 20 21 217.926 $w=1.5e-07 $l=4.25e-07 $layer=POLY_cond $X=13.09 $Y=2.05
+ $X2=12.665 $Y2=2.05
r260 18 91 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=12.395 $Y=2.63
+ $X2=12.395 $Y2=2.26
r261 14 39 88.1957 $w=1.5e-07 $l=1.72e-07 $layer=POLY_cond $X=12.32 $Y=1.665
+ $X2=12.492 $Y2=1.665
r262 14 15 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=12.32 $Y=1.665
+ $X2=11.89 $Y2=1.665
r263 10 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=11.815 $Y=1.59
+ $X2=11.89 $Y2=1.665
r264 10 12 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=11.815 $Y=1.59
+ $X2=11.815 $Y2=0.96
r265 3 53 600 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_PDIFF $count=1 $X=11.35
+ $Y=2.44 $X2=11.49 $Y2=2.655
r266 2 72 600 $w=1.7e-07 $l=7.84267e-07 $layer=licon1_PDIFF $count=1 $X=9.6
+ $Y=2.02 $X2=9.79 $Y2=2.715
r267 2 70 600 $w=1.7e-07 $l=3.27605e-07 $layer=licon1_PDIFF $count=1 $X=9.6
+ $Y=2.02 $X2=9.74 $Y2=2.285
r268 1 44 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=9.6
+ $Y=0.595 $X2=9.74 $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSBP_1%A_2582_150# 1 2 9 11 13 16 18 21 23 24 27
+ 33 35
c63 35 0 1.50676e-19 $X=13.475 $Y=1.83
c64 33 0 1.66769e-19 $X=13.56 $Y=1.325
c65 9 0 5.14661e-20 $X=14.22 $Y=1.415
r66 27 35 22.8272 $w=2.58e-07 $l=5.15e-07 $layer=LI1_cond $X=13.415 $Y=2.345
+ $X2=13.415 $Y2=1.83
r67 24 35 6.91979 $w=3.78e-07 $l=1.9e-07 $layer=LI1_cond $X=13.475 $Y=1.64
+ $X2=13.475 $Y2=1.83
r68 23 33 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=13.56
+ $Y=1.325 $X2=13.56 $Y2=1.325
r69 23 24 9.40151 $w=3.78e-07 $l=3.1e-07 $layer=LI1_cond $X=13.475 $Y=1.33
+ $X2=13.475 $Y2=1.64
r70 19 23 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=13.1 $Y=1.245
+ $X2=13.475 $Y2=1.245
r71 19 21 8.75003 $w=2.68e-07 $l=2.05e-07 $layer=LI1_cond $X=13.1 $Y=1.16
+ $X2=13.1 $Y2=0.955
r72 14 18 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=14.295 $Y=1.49
+ $X2=14.295 $Y2=1.415
r73 14 16 499.947 $w=1.5e-07 $l=9.75e-07 $layer=POLY_cond $X=14.295 $Y=1.49
+ $X2=14.295 $Y2=2.465
r74 11 18 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=14.295 $Y=1.34
+ $X2=14.295 $Y2=1.415
r75 11 13 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=14.295 $Y=1.34
+ $X2=14.295 $Y2=0.81
r76 10 33 19.5363 $w=1.5e-07 $l=2.05122e-07 $layer=POLY_cond $X=13.725 $Y=1.415
+ $X2=13.56 $Y2=1.325
r77 9 18 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=14.22 $Y=1.415
+ $X2=14.295 $Y2=1.415
r78 9 10 253.819 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=14.22 $Y=1.415
+ $X2=13.725 $Y2=1.415
r79 2 27 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=13.24
+ $Y=2.2 $X2=13.38 $Y2=2.345
r80 1 21 182 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_NDIFF $count=1 $X=12.91
+ $Y=0.75 $X2=13.05 $Y2=0.955
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSBP_1%VPWR 1 2 3 4 5 6 7 8 27 31 35 39 43 48 49
+ 50 54 56 57 59 60 61 63 68 76 91 95 114 115 118 121 124 135 137
r162 133 135 8.81011 $w=7.73e-07 $l=5e-09 $layer=LI1_cond $X=8.88 $Y=3.027
+ $X2=8.885 $Y2=3.027
r163 133 134 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r164 131 133 2.46932 $w=7.73e-07 $l=1.6e-07 $layer=LI1_cond $X=8.72 $Y=3.027
+ $X2=8.88 $Y2=3.027
r165 127 128 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r166 124 127 9.7783 $w=3.28e-07 $l=2.8e-07 $layer=LI1_cond $X=4.12 $Y=3.05
+ $X2=4.12 $Y2=3.33
r167 121 122 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r168 118 119 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r169 114 115 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=15.12 $Y=3.33
+ $X2=15.12 $Y2=3.33
r170 112 115 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=14.16 $Y=3.33
+ $X2=15.12 $Y2=3.33
r171 111 112 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=14.16 $Y=3.33
+ $X2=14.16 $Y2=3.33
r172 109 112 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=13.2 $Y=3.33
+ $X2=14.16 $Y2=3.33
r173 108 111 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=13.2 $Y=3.33
+ $X2=14.16 $Y2=3.33
r174 108 109 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=13.2 $Y=3.33
+ $X2=13.2 $Y2=3.33
r175 106 109 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.72 $Y=3.33
+ $X2=13.2 $Y2=3.33
r176 105 106 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=12.72 $Y=3.33
+ $X2=12.72 $Y2=3.33
r177 103 106 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=11.28 $Y=3.33
+ $X2=12.72 $Y2=3.33
r178 103 141 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=3.33
+ $X2=10.8 $Y2=3.33
r179 102 105 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=11.28 $Y=3.33
+ $X2=12.72 $Y2=3.33
r180 102 103 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.28 $Y=3.33
+ $X2=11.28 $Y2=3.33
r181 100 102 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=11.225 $Y=3.33
+ $X2=11.28 $Y2=3.33
r182 99 141 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=3.33
+ $X2=10.8 $Y2=3.33
r183 99 134 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=10.32 $Y=3.33
+ $X2=8.88 $Y2=3.33
r184 98 135 93.6203 $w=1.68e-07 $l=1.435e-06 $layer=LI1_cond $X=10.32 $Y=3.33
+ $X2=8.885 $Y2=3.33
r185 98 99 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.32 $Y=3.33
+ $X2=10.32 $Y2=3.33
r186 95 100 9.90988 $w=1.7e-07 $l=3.83e-07 $layer=LI1_cond $X=10.842 $Y=3.33
+ $X2=11.225 $Y2=3.33
r187 95 141 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=3.33
+ $X2=10.8 $Y2=3.33
r188 95 137 9.45918 $w=7.63e-07 $l=6.05e-07 $layer=LI1_cond $X=10.842 $Y=3.33
+ $X2=10.842 $Y2=2.725
r189 95 98 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=10.46 $Y=3.33
+ $X2=10.32 $Y2=3.33
r190 94 134 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=8.88 $Y2=3.33
r191 93 94 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r192 91 131 3.42619 $w=7.73e-07 $l=2.22e-07 $layer=LI1_cond $X=8.498 $Y=3.027
+ $X2=8.72 $Y2=3.027
r193 91 93 1.51246 $w=7.73e-07 $l=9.8e-08 $layer=LI1_cond $X=8.498 $Y=3.027
+ $X2=8.4 $Y2=3.027
r194 89 90 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r195 87 90 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=7.44 $Y2=3.33
r196 86 87 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r197 84 87 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=6.48 $Y2=3.33
r198 84 128 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=4.08 $Y2=3.33
r199 83 86 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=4.56 $Y=3.33
+ $X2=6.48 $Y2=3.33
r200 83 84 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r201 81 127 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.285 $Y=3.33
+ $X2=4.12 $Y2=3.33
r202 81 83 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=4.285 $Y=3.33
+ $X2=4.56 $Y2=3.33
r203 80 128 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r204 80 122 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=2.64 $Y2=3.33
r205 79 80 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r206 77 121 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.735 $Y=3.33
+ $X2=2.57 $Y2=3.33
r207 77 79 56.4332 $w=1.68e-07 $l=8.65e-07 $layer=LI1_cond $X=2.735 $Y=3.33
+ $X2=3.6 $Y2=3.33
r208 76 127 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.955 $Y=3.33
+ $X2=4.12 $Y2=3.33
r209 76 79 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=3.955 $Y=3.33
+ $X2=3.6 $Y2=3.33
r210 75 122 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r211 74 75 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r212 72 75 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r213 72 119 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r214 71 74 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=3.33 $X2=2.16
+ $Y2=3.33
r215 71 72 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r216 69 118 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.89 $Y=3.33
+ $X2=0.725 $Y2=3.33
r217 69 71 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=0.89 $Y=3.33
+ $X2=1.2 $Y2=3.33
r218 68 121 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.405 $Y=3.33
+ $X2=2.57 $Y2=3.33
r219 68 74 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=2.405 $Y=3.33
+ $X2=2.16 $Y2=3.33
r220 66 119 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r221 65 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r222 63 118 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.56 $Y=3.33
+ $X2=0.725 $Y2=3.33
r223 63 65 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=0.56 $Y=3.33
+ $X2=0.24 $Y2=3.33
r224 61 94 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=7.68 $Y=3.33
+ $X2=8.4 $Y2=3.33
r225 61 90 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=7.68 $Y=3.33
+ $X2=7.44 $Y2=3.33
r226 59 111 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=14.425 $Y=3.33
+ $X2=14.16 $Y2=3.33
r227 59 60 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=14.425 $Y=3.33
+ $X2=14.52 $Y2=3.33
r228 58 114 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=14.615 $Y=3.33
+ $X2=15.12 $Y2=3.33
r229 58 60 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=14.615 $Y=3.33
+ $X2=14.52 $Y2=3.33
r230 56 105 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=12.855 $Y=3.33
+ $X2=12.72 $Y2=3.33
r231 56 57 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=12.855 $Y=3.33
+ $X2=12.985 $Y2=3.33
r232 55 108 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=13.115 $Y=3.33
+ $X2=13.2 $Y2=3.33
r233 55 57 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=13.115 $Y=3.33
+ $X2=12.985 $Y2=3.33
r234 54 89 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=7.65 $Y=3.33
+ $X2=7.44 $Y2=3.33
r235 53 54 11.4338 $w=7.73e-07 $l=1.75e-07 $layer=LI1_cond $X=7.825 $Y=3.027
+ $X2=7.65 $Y2=3.027
r236 50 93 5.60228 $w=7.73e-07 $l=3.63e-07 $layer=LI1_cond $X=8.037 $Y=3.027
+ $X2=8.4 $Y2=3.027
r237 50 53 3.27185 $w=7.73e-07 $l=2.12e-07 $layer=LI1_cond $X=8.037 $Y=3.027
+ $X2=7.825 $Y2=3.027
r238 48 86 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=6.505 $Y=3.33
+ $X2=6.48 $Y2=3.33
r239 48 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.505 $Y=3.33
+ $X2=6.67 $Y2=3.33
r240 47 89 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=6.835 $Y=3.33
+ $X2=7.44 $Y2=3.33
r241 47 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.835 $Y=3.33
+ $X2=6.67 $Y2=3.33
r242 43 46 56.3301 $w=1.88e-07 $l=9.65e-07 $layer=LI1_cond $X=14.52 $Y=2.005
+ $X2=14.52 $Y2=2.97
r243 41 60 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=14.52 $Y=3.245
+ $X2=14.52 $Y2=3.33
r244 41 46 16.0526 $w=1.88e-07 $l=2.75e-07 $layer=LI1_cond $X=14.52 $Y=3.245
+ $X2=14.52 $Y2=2.97
r245 37 57 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=12.985 $Y=3.245
+ $X2=12.985 $Y2=3.33
r246 37 39 39.8923 $w=2.58e-07 $l=9e-07 $layer=LI1_cond $X=12.985 $Y=3.245
+ $X2=12.985 $Y2=2.345
r247 33 49 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.67 $Y=3.245
+ $X2=6.67 $Y2=3.33
r248 33 35 25.1442 $w=3.28e-07 $l=7.2e-07 $layer=LI1_cond $X=6.67 $Y=3.245
+ $X2=6.67 $Y2=2.525
r249 29 121 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.57 $Y=3.245
+ $X2=2.57 $Y2=3.33
r250 29 31 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=2.57 $Y=3.245
+ $X2=2.57 $Y2=2.92
r251 25 118 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.725 $Y=3.245
+ $X2=0.725 $Y2=3.33
r252 25 27 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=0.725 $Y=3.245
+ $X2=0.725 $Y2=2.55
r253 8 46 400 $w=1.7e-07 $l=1.20297e-06 $layer=licon1_PDIFF $count=1 $X=14.37
+ $Y=1.835 $X2=14.51 $Y2=2.97
r254 8 43 400 $w=1.7e-07 $l=2.29565e-07 $layer=licon1_PDIFF $count=1 $X=14.37
+ $Y=1.835 $X2=14.51 $Y2=2.005
r255 7 39 300 $w=1.7e-07 $l=5.1614e-07 $layer=licon1_PDIFF $count=2 $X=12.47
+ $Y=2.42 $X2=12.95 $Y2=2.345
r256 6 137 300 $w=1.7e-07 $l=7.03207e-07 $layer=licon1_PDIFF $count=2 $X=10.485
+ $Y=2.44 $X2=11.06 $Y2=2.725
r257 5 131 400 $w=1.7e-07 $l=1.30398e-06 $layer=licon1_PDIFF $count=1 $X=7.605
+ $Y=2.315 $X2=8.72 $Y2=2.725
r258 5 53 400 $w=1.7e-07 $l=5.08232e-07 $layer=licon1_PDIFF $count=1 $X=7.605
+ $Y=2.315 $X2=7.825 $Y2=2.725
r259 4 35 600 $w=1.7e-07 $l=2.74955e-07 $layer=licon1_PDIFF $count=1 $X=6.52
+ $Y=2.315 $X2=6.67 $Y2=2.525
r260 3 124 600 $w=1.7e-07 $l=9.05345e-07 $layer=licon1_PDIFF $count=1 $X=3.995
+ $Y=2.205 $X2=4.12 $Y2=3.05
r261 2 31 600 $w=1.7e-07 $l=6.45872e-07 $layer=licon1_PDIFF $count=1 $X=2.275
+ $Y=2.405 $X2=2.57 $Y2=2.92
r262 1 27 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=0.585
+ $Y=2.405 $X2=0.725 $Y2=2.55
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSBP_1%A_275_481# 1 2 3 4 15 19 21 24 26 27 28 29
+ 31 34 39 40 47 48
c122 31 0 1.21539e-20 $X=5.365 $Y=1.035
c123 21 0 1.81346e-19 $X=2.905 $Y=0.74
c124 15 0 2.1728e-19 $X=2.37 $Y=0.437
r125 47 49 6.72258 $w=2.98e-07 $l=1.75e-07 $layer=LI1_cond $X=5.425 $Y=2.525
+ $X2=5.425 $Y2=2.7
r126 47 48 8.16804 $w=2.98e-07 $l=1.65e-07 $layer=LI1_cond $X=5.425 $Y=2.525
+ $X2=5.425 $Y2=2.36
r127 40 42 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=3.69 $Y=2.7
+ $X2=3.69 $Y2=2.98
r128 31 45 12.9998 $w=3.33e-07 $l=3.29955e-07 $layer=LI1_cond $X=5.365 $Y=1.035
+ $X2=5.462 $Y2=0.75
r129 31 48 81.6414 $w=1.78e-07 $l=1.325e-06 $layer=LI1_cond $X=5.365 $Y=1.035
+ $X2=5.365 $Y2=2.36
r130 30 40 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.775 $Y=2.7
+ $X2=3.69 $Y2=2.7
r131 29 49 4.061 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=5.275 $Y=2.7 $X2=5.425
+ $Y2=2.7
r132 29 30 97.861 $w=1.68e-07 $l=1.5e-06 $layer=LI1_cond $X=5.275 $Y=2.7
+ $X2=3.775 $Y2=2.7
r133 27 42 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.605 $Y=2.98
+ $X2=3.69 $Y2=2.98
r134 27 28 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=3.605 $Y=2.98
+ $X2=3.075 $Y2=2.98
r135 26 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.99 $Y=2.895
+ $X2=3.075 $Y2=2.98
r136 25 39 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.99 $Y=2.645
+ $X2=2.99 $Y2=2.56
r137 25 26 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=2.99 $Y=2.645
+ $X2=2.99 $Y2=2.895
r138 24 39 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.99 $Y=2.475
+ $X2=2.99 $Y2=2.56
r139 23 24 107.647 $w=1.68e-07 $l=1.65e-06 $layer=LI1_cond $X=2.99 $Y=0.825
+ $X2=2.99 $Y2=2.475
r140 22 37 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.54 $Y=0.74
+ $X2=2.455 $Y2=0.74
r141 21 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.905 $Y=0.74
+ $X2=2.99 $Y2=0.825
r142 21 22 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=2.905 $Y=0.74
+ $X2=2.54 $Y2=0.74
r143 20 34 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.79 $Y=2.56
+ $X2=1.625 $Y2=2.56
r144 19 39 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.905 $Y=2.56
+ $X2=2.99 $Y2=2.56
r145 19 20 72.7433 $w=1.68e-07 $l=1.115e-06 $layer=LI1_cond $X=2.905 $Y=2.56
+ $X2=1.79 $Y2=2.56
r146 15 37 19.7679 $w=1.68e-07 $l=3.03e-07 $layer=LI1_cond $X=2.455 $Y=0.437
+ $X2=2.455 $Y2=0.74
r147 15 17 9.87808 $w=3.13e-07 $l=2.7e-07 $layer=LI1_cond $X=2.37 $Y=0.437
+ $X2=2.1 $Y2=0.437
r148 4 47 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=5.315
+ $Y=2.315 $X2=5.44 $Y2=2.525
r149 3 34 300 $w=1.7e-07 $l=3.2596e-07 $layer=licon1_PDIFF $count=2 $X=1.375
+ $Y=2.405 $X2=1.625 $Y2=2.58
r150 2 45 182 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=1 $X=5.38
+ $Y=0.595 $X2=5.505 $Y2=0.75
r151 1 17 91 $w=1.7e-07 $l=5.755e-07 $layer=licon1_NDIFF $count=2 $X=1.62
+ $Y=0.235 $X2=2.1 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSBP_1%Q 1 2 7 8 9 10 11 18
r20 11 32 4.64417 $w=3.33e-07 $l=1.35e-07 $layer=LI1_cond $X=14.082 $Y=2.775
+ $X2=14.082 $Y2=2.91
r21 10 11 12.7285 $w=3.33e-07 $l=3.7e-07 $layer=LI1_cond $X=14.082 $Y=2.405
+ $X2=14.082 $Y2=2.775
r22 9 10 14.6205 $w=3.33e-07 $l=4.25e-07 $layer=LI1_cond $X=14.082 $Y=1.98
+ $X2=14.082 $Y2=2.405
r23 8 9 10.8364 $w=3.33e-07 $l=3.15e-07 $layer=LI1_cond $X=14.082 $Y=1.665
+ $X2=14.082 $Y2=1.98
r24 7 8 12.7285 $w=3.33e-07 $l=3.7e-07 $layer=LI1_cond $X=14.082 $Y=1.295
+ $X2=14.082 $Y2=1.665
r25 7 18 6.53624 $w=3.33e-07 $l=1.9e-07 $layer=LI1_cond $X=14.082 $Y=1.295
+ $X2=14.082 $Y2=1.105
r26 2 32 400 $w=1.7e-07 $l=1.13578e-06 $layer=licon1_PDIFF $count=1 $X=13.955
+ $Y=1.835 $X2=14.08 $Y2=2.91
r27 2 9 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=13.955
+ $Y=1.835 $X2=14.08 $Y2=1.98
r28 1 18 182 $w=1.7e-07 $l=7.84156e-07 $layer=licon1_NDIFF $count=1 $X=13.935
+ $Y=0.39 $X2=14.08 $Y2=1.105
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSBP_1%Q_N 1 2 7 8 9 10 11 12 13 46
r13 33 46 0.654797 $w=4.38e-07 $l=2.5e-08 $layer=LI1_cond $X=15.055 $Y=2.06
+ $X2=15.055 $Y2=2.035
r14 13 40 3.5359 $w=4.38e-07 $l=1.35e-07 $layer=LI1_cond $X=15.055 $Y=2.775
+ $X2=15.055 $Y2=2.91
r15 12 13 9.691 $w=4.38e-07 $l=3.7e-07 $layer=LI1_cond $X=15.055 $Y=2.405
+ $X2=15.055 $Y2=2.775
r16 11 46 0.785757 $w=4.38e-07 $l=3e-08 $layer=LI1_cond $X=15.055 $Y=2.005
+ $X2=15.055 $Y2=2.035
r17 11 44 6.03044 $w=4.38e-07 $l=1.65e-07 $layer=LI1_cond $X=15.055 $Y=2.005
+ $X2=15.055 $Y2=1.84
r18 11 12 8.25044 $w=4.38e-07 $l=3.15e-07 $layer=LI1_cond $X=15.055 $Y=2.09
+ $X2=15.055 $Y2=2.405
r19 11 33 0.785757 $w=4.38e-07 $l=3e-08 $layer=LI1_cond $X=15.055 $Y=2.09
+ $X2=15.055 $Y2=2.06
r20 10 44 7.46954 $w=2.68e-07 $l=1.75e-07 $layer=LI1_cond $X=15.14 $Y=1.665
+ $X2=15.14 $Y2=1.84
r21 9 10 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=15.14 $Y=1.295
+ $X2=15.14 $Y2=1.665
r22 8 9 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=15.14 $Y=0.925
+ $X2=15.14 $Y2=1.295
r23 7 8 16.2196 $w=2.68e-07 $l=3.8e-07 $layer=LI1_cond $X=15.14 $Y=0.545
+ $X2=15.14 $Y2=0.925
r24 2 11 400 $w=1.7e-07 $l=2.29565e-07 $layer=licon1_PDIFF $count=1 $X=14.8
+ $Y=1.835 $X2=14.94 $Y2=2.005
r25 2 40 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=14.8
+ $Y=1.835 $X2=14.94 $Y2=2.91
r26 1 7 91 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=2 $X=14.96
+ $Y=0.39 $X2=15.1 $Y2=0.545
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSBP_1%VGND 1 2 3 4 5 6 7 8 27 31 35 39 43 47 51
+ 55 58 59 61 62 64 65 67 68 70 71 72 96 107 111 121 122 125 128 131
c166 47 0 1.86545e-20 $X=10.985 $Y=0.795
r167 131 132 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.64 $Y=0
+ $X2=14.64 $Y2=0
r168 128 129 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.24 $Y=0
+ $X2=12.24 $Y2=0
r169 125 126 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=8.88 $Y=0
+ $X2=8.88 $Y2=0
r170 122 132 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=15.12 $Y=0
+ $X2=14.64 $Y2=0
r171 121 122 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=15.12 $Y=0
+ $X2=15.12 $Y2=0
r172 119 131 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=14.755 $Y=0
+ $X2=14.59 $Y2=0
r173 119 121 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=14.755 $Y=0
+ $X2=15.12 $Y2=0
r174 118 132 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=14.16 $Y=0
+ $X2=14.64 $Y2=0
r175 117 118 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=14.16 $Y=0
+ $X2=14.16 $Y2=0
r176 115 118 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=12.72 $Y=0
+ $X2=14.16 $Y2=0
r177 115 129 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.72 $Y=0
+ $X2=12.24 $Y2=0
r178 114 117 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=12.72 $Y=0
+ $X2=14.16 $Y2=0
r179 114 115 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=12.72 $Y=0
+ $X2=12.72 $Y2=0
r180 112 128 12.0118 $w=1.7e-07 $l=2.78e-07 $layer=LI1_cond $X=12.455 $Y=0
+ $X2=12.177 $Y2=0
r181 112 114 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=12.455 $Y=0
+ $X2=12.72 $Y2=0
r182 111 131 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=14.425 $Y=0
+ $X2=14.59 $Y2=0
r183 111 117 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=14.425 $Y=0
+ $X2=14.16 $Y2=0
r184 110 129 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.76 $Y=0
+ $X2=12.24 $Y2=0
r185 109 110 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.76 $Y=0
+ $X2=11.76 $Y2=0
r186 107 128 12.0118 $w=1.7e-07 $l=2.77e-07 $layer=LI1_cond $X=11.9 $Y=0
+ $X2=12.177 $Y2=0
r187 107 109 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=11.9 $Y=0
+ $X2=11.76 $Y2=0
r188 106 110 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=10.8 $Y=0
+ $X2=11.76 $Y2=0
r189 105 106 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.8 $Y=0
+ $X2=10.8 $Y2=0
r190 103 106 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=9.36 $Y=0
+ $X2=10.8 $Y2=0
r191 103 126 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=0
+ $X2=8.88 $Y2=0
r192 102 105 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=9.36 $Y=0
+ $X2=10.8 $Y2=0
r193 102 103 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.36 $Y=0
+ $X2=9.36 $Y2=0
r194 100 125 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=9.055 $Y=0 $X2=8.955
+ $Y2=0
r195 100 102 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=9.055 $Y=0
+ $X2=9.36 $Y2=0
r196 98 99 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.96 $Y=0
+ $X2=6.96 $Y2=0
r197 96 125 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=8.855 $Y=0 $X2=8.955
+ $Y2=0
r198 96 98 123.631 $w=1.68e-07 $l=1.895e-06 $layer=LI1_cond $X=8.855 $Y=0
+ $X2=6.96 $Y2=0
r199 95 99 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6.96
+ $Y2=0
r200 94 95 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.48 $Y=0
+ $X2=6.48 $Y2=0
r201 92 95 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=4.56 $Y=0
+ $X2=6.48 $Y2=0
r202 91 94 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=4.56 $Y=0 $X2=6.48
+ $Y2=0
r203 91 92 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.56 $Y=0
+ $X2=4.56 $Y2=0
r204 89 92 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=4.56
+ $Y2=0
r205 88 89 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r206 86 89 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=4.08
+ $Y2=0
r207 85 88 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=3.12 $Y=0 $X2=4.08
+ $Y2=0
r208 85 86 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r209 83 86 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r210 82 83 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r211 80 83 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.64
+ $Y2=0
r212 79 82 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.64
+ $Y2=0
r213 79 80 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r214 76 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r215 75 76 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r216 72 126 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=7.68 $Y=0
+ $X2=8.88 $Y2=0
r217 72 99 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=7.68 $Y=0 $X2=6.96
+ $Y2=0
r218 70 105 1.30481 $w=1.68e-07 $l=2e-08 $layer=LI1_cond $X=10.82 $Y=0 $X2=10.8
+ $Y2=0
r219 70 71 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.82 $Y=0
+ $X2=10.985 $Y2=0
r220 69 109 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=11.15 $Y=0
+ $X2=11.76 $Y2=0
r221 69 71 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.15 $Y=0
+ $X2=10.985 $Y2=0
r222 67 94 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=6.56 $Y=0 $X2=6.48
+ $Y2=0
r223 67 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.56 $Y=0 $X2=6.725
+ $Y2=0
r224 66 98 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=6.89 $Y=0 $X2=6.96
+ $Y2=0
r225 66 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.89 $Y=0 $X2=6.725
+ $Y2=0
r226 64 88 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=4.295 $Y=0
+ $X2=4.08 $Y2=0
r227 64 65 6.81202 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=4.295 $Y=0 $X2=4.415
+ $Y2=0
r228 63 91 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=4.535 $Y=0 $X2=4.56
+ $Y2=0
r229 63 65 6.81202 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=4.535 $Y=0 $X2=4.415
+ $Y2=0
r230 62 85 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.955 $Y=0 $X2=3.12
+ $Y2=0
r231 61 82 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=2.79 $Y=0 $X2=2.64
+ $Y2=0
r232 61 62 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.79 $Y=0 $X2=2.955
+ $Y2=0
r233 58 75 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=0.805 $Y=0 $X2=0.72
+ $Y2=0
r234 58 59 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.805 $Y=0 $X2=0.97
+ $Y2=0
r235 57 79 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=1.135 $Y=0 $X2=1.2
+ $Y2=0
r236 57 59 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.135 $Y=0 $X2=0.97
+ $Y2=0
r237 53 131 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=14.59 $Y=0.085
+ $X2=14.59 $Y2=0
r238 53 55 11.1752 $w=3.28e-07 $l=3.2e-07 $layer=LI1_cond $X=14.59 $Y=0.085
+ $X2=14.59 $Y2=0.405
r239 49 128 2.33542 $w=5.55e-07 $l=8.5e-08 $layer=LI1_cond $X=12.177 $Y=0.085
+ $X2=12.177 $Y2=0
r240 49 51 17.8873 $w=5.53e-07 $l=8.3e-07 $layer=LI1_cond $X=12.177 $Y=0.085
+ $X2=12.177 $Y2=0.915
r241 45 71 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.985 $Y=0.085
+ $X2=10.985 $Y2=0
r242 45 47 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=10.985 $Y=0.085
+ $X2=10.985 $Y2=0.795
r243 41 125 0.764409 $w=2e-07 $l=8.5e-08 $layer=LI1_cond $X=8.955 $Y=0.085
+ $X2=8.955 $Y2=0
r244 41 43 36.6 $w=1.98e-07 $l=6.6e-07 $layer=LI1_cond $X=8.955 $Y=0.085
+ $X2=8.955 $Y2=0.745
r245 37 68 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.725 $Y=0.085
+ $X2=6.725 $Y2=0
r246 37 39 22.8742 $w=3.28e-07 $l=6.55e-07 $layer=LI1_cond $X=6.725 $Y=0.085
+ $X2=6.725 $Y2=0.74
r247 33 65 0.135687 $w=2.4e-07 $l=8.5e-08 $layer=LI1_cond $X=4.415 $Y=0.085
+ $X2=4.415 $Y2=0
r248 33 35 23.0489 $w=2.38e-07 $l=4.8e-07 $layer=LI1_cond $X=4.415 $Y=0.085
+ $X2=4.415 $Y2=0.565
r249 29 62 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.955 $Y=0.085
+ $X2=2.955 $Y2=0
r250 29 31 10.1275 $w=3.28e-07 $l=2.9e-07 $layer=LI1_cond $X=2.955 $Y=0.085
+ $X2=2.955 $Y2=0.375
r251 25 59 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.97 $Y=0.085
+ $X2=0.97 $Y2=0
r252 25 27 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=0.97 $Y=0.085
+ $X2=0.97 $Y2=0.445
r253 8 55 182 $w=1.7e-07 $l=2.27376e-07 $layer=licon1_NDIFF $count=1 $X=14.37
+ $Y=0.39 $X2=14.59 $Y2=0.405
r254 7 51 91 $w=1.7e-07 $l=5.56417e-07 $layer=licon1_NDIFF $count=2 $X=11.89
+ $Y=0.75 $X2=12.37 $Y2=0.915
r255 6 47 182 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_NDIFF $count=1 $X=10.845
+ $Y=0.59 $X2=10.985 $Y2=0.795
r256 5 43 182 $w=1.7e-07 $l=7.86432e-07 $layer=licon1_NDIFF $count=1 $X=8.235
+ $Y=0.595 $X2=8.95 $Y2=0.745
r257 4 39 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=6.585
+ $Y=0.595 $X2=6.725 $Y2=0.74
r258 3 35 182 $w=1.7e-07 $l=2.54951e-07 $layer=licon1_NDIFF $count=1 $X=4.285
+ $Y=0.365 $X2=4.41 $Y2=0.565
r259 2 31 182 $w=1.7e-07 $l=1.9799e-07 $layer=licon1_NDIFF $count=1 $X=2.815
+ $Y=0.235 $X2=2.955 $Y2=0.375
r260 1 27 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.83
+ $Y=0.235 $X2=0.97 $Y2=0.445
.ends

