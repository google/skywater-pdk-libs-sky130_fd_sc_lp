* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__a31o_m A1 A2 A3 B1 VGND VNB VPB VPWR X
X0 VPWR A1 a_274_512# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X1 a_274_512# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X2 X a_86_172# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 a_274_512# B1 a_86_172# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X4 a_282_66# A2 a_354_66# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 X a_86_172# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X6 a_354_66# A1 a_86_172# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 a_86_172# B1 VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 VPWR A3 a_274_512# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X9 VGND A3 a_282_66# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
