* NGSPICE file created from sky130_fd_sc_lp__a221oi_0.ext - technology: sky130A

.subckt sky130_fd_sc_lp__a221oi_0 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
M1000 a_228_47# B2 VGND VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=2.856e+11p ps=3.04e+06u
M1001 Y B1 a_228_47# VNB nshort w=420000u l=150000u
+  ad=2.625e+11p pd=2.93e+06u as=0p ps=0u
M1002 a_242_487# B2 a_156_487# VPB phighvt w=640000u l=150000u
+  ad=4.864e+11p pd=4.08e+06u as=3.936e+11p ps=3.79e+06u
M1003 VPWR A1 a_242_487# VPB phighvt w=640000u l=150000u
+  ad=2.24e+11p pd=1.98e+06u as=0p ps=0u
M1004 a_242_487# A2 VPWR VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VGND A2 a_408_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1006 a_408_47# A1 Y VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_156_487# C1 Y VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.696e+11p ps=1.81e+06u
M1008 a_156_487# B1 a_242_487# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND C1 Y VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

