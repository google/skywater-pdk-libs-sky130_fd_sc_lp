* File: sky130_fd_sc_lp__nand4bb_2.spice
* Created: Wed Sep  2 10:06:46 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__nand4bb_2.pex.spice"
.subckt sky130_fd_sc_lp__nand4bb_2  VNB VPB B_N A_N C D VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* D	D
* C	C
* A_N	A_N
* B_N	B_N
* VPB	VPB
* VNB	VNB
MM1015 N_VGND_M1015_d N_B_N_M1015_g N_A_27_373#_M1015_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1016 N_A_223_49#_M1016_d N_A_N_M1016_g N_VGND_M1015_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1008 N_Y_M1008_d N_A_223_49#_M1008_g N_A_357_47#_M1008_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75001.6 A=0.126 P=1.98 MULT=1
MM1013 N_Y_M1008_d N_A_223_49#_M1013_g N_A_357_47#_M1013_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1218 PD=1.12 PS=1.13 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1005 N_A_357_47#_M1013_s N_A_27_373#_M1005_g N_A_614_47#_M1005_s VNB NSHORT
+ L=0.15 W=0.84 AD=0.1218 AS=0.147 PD=1.13 PS=1.19 NRD=1.428 NRS=9.996 M=1 R=5.6
+ SA=75001.1 SB=75000.7 A=0.126 P=1.98 MULT=1
MM1009 N_A_357_47#_M1009_d N_A_27_373#_M1009_g N_A_614_47#_M1005_s VNB NSHORT
+ L=0.15 W=0.84 AD=0.2226 AS=0.147 PD=2.21 PS=1.19 NRD=0 NRS=0 M=1 R=5.6
+ SA=75001.6 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1007 N_A_614_47#_M1007_d N_C_M1007_g N_A_821_47#_M1007_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75001.5 A=0.126 P=1.98 MULT=1
MM1017 N_A_614_47#_M1007_d N_C_M1017_g N_A_821_47#_M1017_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1002 N_VGND_M1002_d N_D_M1002_g N_A_821_47#_M1017_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.1
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1010 N_VGND_M1002_d N_D_M1010_g N_A_821_47#_M1010_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75001.5
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1000 N_VPWR_M1000_d N_B_N_M1000_g N_A_27_373#_M1000_s VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1155 AS=0.1113 PD=0.97 PS=1.37 NRD=9.3772 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.9 A=0.063 P=1.14 MULT=1
MM1006 N_A_223_49#_M1006_d N_A_N_M1006_g N_VPWR_M1000_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1113 AS=0.1155 PD=1.37 PS=0.97 NRD=0 NRS=117.254 M=1 R=2.8
+ SA=75000.9 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1003 N_Y_M1003_d N_A_223_49#_M1003_g N_VPWR_M1003_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75003.6 A=0.189 P=2.82 MULT=1
MM1018 N_Y_M1003_d N_A_223_49#_M1018_g N_VPWR_M1018_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75003.1 A=0.189 P=2.82 MULT=1
MM1001 N_Y_M1001_d N_A_27_373#_M1001_g N_VPWR_M1018_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75002.7 A=0.189 P=2.82 MULT=1
MM1012 N_Y_M1001_d N_A_27_373#_M1012_g N_VPWR_M1012_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.5
+ SB=75002.3 A=0.189 P=2.82 MULT=1
MM1004 N_Y_M1004_d N_C_M1004_g N_VPWR_M1012_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.9
+ SB=75001.9 A=0.189 P=2.82 MULT=1
MM1019 N_Y_M1004_d N_C_M1019_g N_VPWR_M1019_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.3
+ SB=75001.4 A=0.189 P=2.82 MULT=1
MM1011 N_Y_M1011_d N_D_M1011_g N_VPWR_M1019_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.4158 AS=0.1764 PD=1.92 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.8 SB=75001
+ A=0.189 P=2.82 MULT=1
MM1014 N_Y_M1011_d N_D_M1014_g N_VPWR_M1014_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.4158 AS=0.3339 PD=1.92 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75003.6
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX20_noxref VNB VPB NWDIODE A=12.3463 P=16.97
c_63 VNB 0 1.27355e-19 $X=0 $Y=0
*
.include "sky130_fd_sc_lp__nand4bb_2.pxi.spice"
*
.ends
*
*
