* File: sky130_fd_sc_lp__o31a_4.pxi.spice
* Created: Fri Aug 28 11:15:40 2020
* 
x_PM_SKY130_FD_SC_LP__O31A_4%A_101_23# N_A_101_23#_M1014_d N_A_101_23#_M1006_s
+ N_A_101_23#_M1015_s N_A_101_23#_M1001_g N_A_101_23#_M1000_g
+ N_A_101_23#_M1012_g N_A_101_23#_M1009_g N_A_101_23#_M1016_g
+ N_A_101_23#_M1010_g N_A_101_23#_M1017_g N_A_101_23#_M1019_g
+ N_A_101_23#_c_121_n N_A_101_23#_c_122_n N_A_101_23#_c_123_n
+ N_A_101_23#_c_124_n N_A_101_23#_c_125_n N_A_101_23#_c_133_n
+ N_A_101_23#_c_147_p N_A_101_23#_c_126_n N_A_101_23#_c_179_p
+ N_A_101_23#_c_159_p N_A_101_23#_c_127_n PM_SKY130_FD_SC_LP__O31A_4%A_101_23#
x_PM_SKY130_FD_SC_LP__O31A_4%B1 N_B1_M1006_g N_B1_c_247_n N_B1_c_248_n
+ N_B1_M1013_g N_B1_M1014_g N_B1_M1021_g B1 B1 N_B1_c_251_n N_B1_c_255_n
+ PM_SKY130_FD_SC_LP__O31A_4%B1
x_PM_SKY130_FD_SC_LP__O31A_4%A3 N_A3_M1003_g N_A3_M1015_g N_A3_M1018_g
+ N_A3_M1023_g A3 A3 A3 N_A3_c_308_n PM_SKY130_FD_SC_LP__O31A_4%A3
x_PM_SKY130_FD_SC_LP__O31A_4%A2 N_A2_M1002_g N_A2_M1007_g N_A2_M1004_g
+ N_A2_M1020_g N_A2_c_366_n N_A2_c_360_n N_A2_c_361_n A2 N_A2_c_362_n
+ N_A2_c_363_n N_A2_c_370_n A2 PM_SKY130_FD_SC_LP__O31A_4%A2
x_PM_SKY130_FD_SC_LP__O31A_4%A1 N_A1_c_433_n N_A1_M1008_g N_A1_M1005_g
+ N_A1_c_435_n N_A1_M1022_g N_A1_M1011_g A1 A1 N_A1_c_438_n
+ PM_SKY130_FD_SC_LP__O31A_4%A1
x_PM_SKY130_FD_SC_LP__O31A_4%VPWR N_VPWR_M1000_d N_VPWR_M1009_d N_VPWR_M1019_d
+ N_VPWR_M1013_d N_VPWR_M1005_s N_VPWR_c_488_n N_VPWR_c_489_n N_VPWR_c_490_n
+ N_VPWR_c_491_n N_VPWR_c_492_n N_VPWR_c_493_n N_VPWR_c_494_n N_VPWR_c_495_n
+ N_VPWR_c_496_n N_VPWR_c_497_n N_VPWR_c_498_n VPWR N_VPWR_c_499_n
+ N_VPWR_c_500_n N_VPWR_c_501_n N_VPWR_c_502_n N_VPWR_c_487_n
+ PM_SKY130_FD_SC_LP__O31A_4%VPWR
x_PM_SKY130_FD_SC_LP__O31A_4%X N_X_M1001_d N_X_M1016_d N_X_M1000_s N_X_M1010_s
+ N_X_c_588_n N_X_c_593_n N_X_c_594_n N_X_c_640_p N_X_c_589_n N_X_c_626_n
+ N_X_c_595_n N_X_c_641_p N_X_c_631_n N_X_c_590_n N_X_c_596_n X X N_X_c_591_n X
+ PM_SKY130_FD_SC_LP__O31A_4%X
x_PM_SKY130_FD_SC_LP__O31A_4%A_720_367# N_A_720_367#_M1015_d
+ N_A_720_367#_M1023_d N_A_720_367#_M1020_s N_A_720_367#_c_646_n
+ N_A_720_367#_c_658_n N_A_720_367#_c_647_n N_A_720_367#_c_660_n
+ PM_SKY130_FD_SC_LP__O31A_4%A_720_367#
x_PM_SKY130_FD_SC_LP__O31A_4%A_975_367# N_A_975_367#_M1007_d
+ N_A_975_367#_M1011_d N_A_975_367#_c_698_n N_A_975_367#_c_706_n
+ N_A_975_367#_c_692_n PM_SKY130_FD_SC_LP__O31A_4%A_975_367#
x_PM_SKY130_FD_SC_LP__O31A_4%VGND N_VGND_M1001_s N_VGND_M1012_s N_VGND_M1017_s
+ N_VGND_M1003_d N_VGND_M1002_d N_VGND_M1022_s N_VGND_c_708_n N_VGND_c_709_n
+ N_VGND_c_710_n N_VGND_c_711_n N_VGND_c_712_n N_VGND_c_713_n N_VGND_c_714_n
+ VGND N_VGND_c_715_n N_VGND_c_716_n N_VGND_c_717_n N_VGND_c_718_n
+ N_VGND_c_719_n N_VGND_c_720_n N_VGND_c_721_n N_VGND_c_722_n N_VGND_c_723_n
+ N_VGND_c_724_n N_VGND_c_725_n N_VGND_c_726_n PM_SKY130_FD_SC_LP__O31A_4%VGND
x_PM_SKY130_FD_SC_LP__O31A_4%A_528_65# N_A_528_65#_M1014_s N_A_528_65#_M1021_s
+ N_A_528_65#_M1018_s N_A_528_65#_M1008_d N_A_528_65#_M1004_s
+ N_A_528_65#_c_808_n N_A_528_65#_c_809_n N_A_528_65#_c_810_n
+ N_A_528_65#_c_811_n N_A_528_65#_c_812_n N_A_528_65#_c_813_n
+ N_A_528_65#_c_841_n N_A_528_65#_c_814_n N_A_528_65#_c_815_n
+ N_A_528_65#_c_816_n N_A_528_65#_c_817_n N_A_528_65#_c_860_n
+ PM_SKY130_FD_SC_LP__O31A_4%A_528_65#
cc_1 VNB N_A_101_23#_M1001_g 0.0259723f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=0.665
cc_2 VNB N_A_101_23#_M1012_g 0.0213935f $X=-0.19 $Y=-0.245 $X2=1.01 $Y2=0.665
cc_3 VNB N_A_101_23#_M1016_g 0.0214129f $X=-0.19 $Y=-0.245 $X2=1.44 $Y2=0.665
cc_4 VNB N_A_101_23#_M1017_g 0.0278929f $X=-0.19 $Y=-0.245 $X2=1.87 $Y2=0.665
cc_5 VNB N_A_101_23#_c_121_n 0.0129176f $X=-0.19 $Y=-0.245 $X2=2.635 $Y2=1.49
cc_6 VNB N_A_101_23#_c_122_n 0.00242998f $X=-0.19 $Y=-0.245 $X2=2.735 $Y2=1.405
cc_7 VNB N_A_101_23#_c_123_n 0.00118309f $X=-0.19 $Y=-0.245 $X2=2.74 $Y2=1.98
cc_8 VNB N_A_101_23#_c_124_n 0.00671633f $X=-0.19 $Y=-0.245 $X2=3.13 $Y2=1.16
cc_9 VNB N_A_101_23#_c_125_n 0.00288238f $X=-0.19 $Y=-0.245 $X2=2.835 $Y2=1.16
cc_10 VNB N_A_101_23#_c_126_n 8.64934e-19 $X=-0.19 $Y=-0.245 $X2=2.735 $Y2=1.49
cc_11 VNB N_A_101_23#_c_127_n 0.087855f $X=-0.19 $Y=-0.245 $X2=2.095 $Y2=1.49
cc_12 VNB N_B1_M1006_g 0.00737266f $X=-0.19 $Y=-0.245 $X2=4.015 $Y2=1.835
cc_13 VNB N_B1_c_247_n 0.0156451f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_B1_c_248_n 0.012929f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_B1_M1014_g 0.023132f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_B1_M1021_g 0.0197604f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_B1_c_251_n 0.0459421f $X=-0.19 $Y=-0.245 $X2=1.44 $Y2=1.325
cc_18 VNB N_A3_M1003_g 0.0194944f $X=-0.19 $Y=-0.245 $X2=4.015 $Y2=1.835
cc_19 VNB N_A3_M1018_g 0.0195091f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=0.665
cc_20 VNB A3 0.00886055f $X=-0.19 $Y=-0.245 $X2=1.01 $Y2=0.665
cc_21 VNB N_A3_c_308_n 0.0319393f $X=-0.19 $Y=-0.245 $X2=1.44 $Y2=0.665
cc_22 VNB N_A2_M1002_g 0.02274f $X=-0.19 $Y=-0.245 $X2=4.015 $Y2=1.835
cc_23 VNB N_A2_M1004_g 0.0242392f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=0.665
cc_24 VNB N_A2_M1020_g 0.0018481f $X=-0.19 $Y=-0.245 $X2=0.805 $Y2=2.465
cc_25 VNB N_A2_c_360_n 0.00409935f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A2_c_361_n 0.054269f $X=-0.19 $Y=-0.245 $X2=1.235 $Y2=1.655
cc_27 VNB N_A2_c_362_n 0.0279412f $X=-0.19 $Y=-0.245 $X2=1.44 $Y2=0.665
cc_28 VNB N_A2_c_363_n 0.00620331f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A1_c_433_n 0.0180359f $X=-0.19 $Y=-0.245 $X2=3.155 $Y2=0.325
cc_30 VNB N_A1_M1005_g 0.00242879f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A1_c_435_n 0.0158864f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A1_M1011_g 0.00256904f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB A1 0.00892449f $X=-0.19 $Y=-0.245 $X2=0.805 $Y2=2.465
cc_34 VNB N_A1_c_438_n 0.0365224f $X=-0.19 $Y=-0.245 $X2=1.235 $Y2=2.465
cc_35 VNB N_VPWR_c_487_n 0.283096f $X=-0.19 $Y=-0.245 $X2=1.87 $Y2=1.49
cc_36 VNB N_X_c_588_n 0.00262291f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_X_c_589_n 0.00621437f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_X_c_590_n 0.00147023f $X=-0.19 $Y=-0.245 $X2=2.635 $Y2=1.49
cc_39 VNB N_X_c_591_n 0.0134283f $X=-0.19 $Y=-0.245 $X2=2.03 $Y2=1.49
cc_40 VNB X 0.0228864f $X=-0.19 $Y=-0.245 $X2=2.735 $Y2=1.405
cc_41 VNB N_VGND_c_708_n 0.0137908f $X=-0.19 $Y=-0.245 $X2=1.01 $Y2=0.665
cc_42 VNB N_VGND_c_709_n 0.0281524f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_710_n 4.71799e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_711_n 0.0222109f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_712_n 0.00236188f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_713_n 0.00688794f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_714_n 0.00236631f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_715_n 0.0130715f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.49
cc_49 VNB N_VGND_c_716_n 0.0130715f $X=-0.19 $Y=-0.245 $X2=2.735 $Y2=1.245
cc_50 VNB N_VGND_c_717_n 0.0432975f $X=-0.19 $Y=-0.245 $X2=2.74 $Y2=1.98
cc_51 VNB N_VGND_c_718_n 0.0165332f $X=-0.19 $Y=-0.245 $X2=3.295 $Y2=0.69
cc_52 VNB N_VGND_c_719_n 0.0166924f $X=-0.19 $Y=-0.245 $X2=2.735 $Y2=1.49
cc_53 VNB N_VGND_c_720_n 0.0161944f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.49
cc_54 VNB N_VGND_c_721_n 0.370406f $X=-0.19 $Y=-0.245 $X2=0.805 $Y2=1.49
cc_55 VNB N_VGND_c_722_n 0.00451663f $X=-0.19 $Y=-0.245 $X2=2.03 $Y2=1.49
cc_56 VNB N_VGND_c_723_n 0.00521013f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_VGND_c_724_n 0.00549308f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_725_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_726_n 0.00549308f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_528_65#_c_808_n 0.00535789f $X=-0.19 $Y=-0.245 $X2=1.01 $Y2=1.325
cc_61 VNB N_A_528_65#_c_809_n 0.00460382f $X=-0.19 $Y=-0.245 $X2=1.01 $Y2=0.665
cc_62 VNB N_A_528_65#_c_810_n 0.0048949f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_A_528_65#_c_811_n 0.00310505f $X=-0.19 $Y=-0.245 $X2=1.44 $Y2=1.325
cc_64 VNB N_A_528_65#_c_812_n 0.00241833f $X=-0.19 $Y=-0.245 $X2=1.44 $Y2=0.665
cc_65 VNB N_A_528_65#_c_813_n 0.00200301f $X=-0.19 $Y=-0.245 $X2=1.665 $Y2=1.655
cc_66 VNB N_A_528_65#_c_814_n 0.00200301f $X=-0.19 $Y=-0.245 $X2=1.87 $Y2=0.665
cc_67 VNB N_A_528_65#_c_815_n 0.00850359f $X=-0.19 $Y=-0.245 $X2=2.095 $Y2=1.655
cc_68 VNB N_A_528_65#_c_816_n 0.0235434f $X=-0.19 $Y=-0.245 $X2=2.635 $Y2=1.49
cc_69 VNB N_A_528_65#_c_817_n 0.00319622f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VPB N_A_101_23#_M1000_g 0.022883f $X=-0.19 $Y=1.655 $X2=0.805 $Y2=2.465
cc_71 VPB N_A_101_23#_M1009_g 0.0188632f $X=-0.19 $Y=1.655 $X2=1.235 $Y2=2.465
cc_72 VPB N_A_101_23#_M1010_g 0.0188632f $X=-0.19 $Y=1.655 $X2=1.665 $Y2=2.465
cc_73 VPB N_A_101_23#_M1019_g 0.0197141f $X=-0.19 $Y=1.655 $X2=2.095 $Y2=2.465
cc_74 VPB N_A_101_23#_c_123_n 0.00328487f $X=-0.19 $Y=1.655 $X2=2.74 $Y2=1.98
cc_75 VPB N_A_101_23#_c_133_n 0.0189477f $X=-0.19 $Y=1.655 $X2=3.99 $Y2=2.375
cc_76 VPB N_A_101_23#_c_127_n 0.0138863f $X=-0.19 $Y=1.655 $X2=2.095 $Y2=1.49
cc_77 VPB N_B1_M1006_g 0.0197397f $X=-0.19 $Y=1.655 $X2=4.015 $Y2=1.835
cc_78 VPB N_B1_M1013_g 0.0222235f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_79 VPB N_B1_c_251_n 0.0105341f $X=-0.19 $Y=1.655 $X2=1.44 $Y2=1.325
cc_80 VPB N_B1_c_255_n 0.00535433f $X=-0.19 $Y=1.655 $X2=1.44 $Y2=0.665
cc_81 VPB N_A3_M1015_g 0.022883f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_82 VPB N_A3_M1023_g 0.0183189f $X=-0.19 $Y=1.655 $X2=0.805 $Y2=2.465
cc_83 VPB A3 0.0101297f $X=-0.19 $Y=1.655 $X2=1.01 $Y2=0.665
cc_84 VPB N_A3_c_308_n 0.00477272f $X=-0.19 $Y=1.655 $X2=1.44 $Y2=0.665
cc_85 VPB N_A2_M1007_g 0.0203869f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_86 VPB N_A2_M1020_g 0.0239978f $X=-0.19 $Y=1.655 $X2=0.805 $Y2=2.465
cc_87 VPB N_A2_c_366_n 0.0142451f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_88 VPB N_A2_c_360_n 0.00182616f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_89 VPB N_A2_c_362_n 0.00781826f $X=-0.19 $Y=1.655 $X2=1.44 $Y2=0.665
cc_90 VPB N_A2_c_363_n 4.95949e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_91 VPB N_A2_c_370_n 0.00142005f $X=-0.19 $Y=1.655 $X2=1.87 $Y2=0.665
cc_92 VPB N_A1_M1005_g 0.020248f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_93 VPB N_A1_M1011_g 0.0188011f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_94 VPB N_VPWR_c_488_n 0.0415892f $X=-0.19 $Y=1.655 $X2=1.01 $Y2=1.325
cc_95 VPB N_VPWR_c_489_n 3.0911e-19 $X=-0.19 $Y=1.655 $X2=1.235 $Y2=2.465
cc_96 VPB N_VPWR_c_490_n 0.0130339f $X=-0.19 $Y=1.655 $X2=1.44 $Y2=0.665
cc_97 VPB N_VPWR_c_491_n 0.00319877f $X=-0.19 $Y=1.655 $X2=1.665 $Y2=2.465
cc_98 VPB N_VPWR_c_492_n 0.0095672f $X=-0.19 $Y=1.655 $X2=2.095 $Y2=1.655
cc_99 VPB N_VPWR_c_493_n 0.0100738f $X=-0.19 $Y=1.655 $X2=2.095 $Y2=2.465
cc_100 VPB N_VPWR_c_494_n 0.0313042f $X=-0.19 $Y=1.655 $X2=0.67 $Y2=1.49
cc_101 VPB N_VPWR_c_495_n 0.0156676f $X=-0.19 $Y=1.655 $X2=2.03 $Y2=1.49
cc_102 VPB N_VPWR_c_496_n 0.00510842f $X=-0.19 $Y=1.655 $X2=2.03 $Y2=1.49
cc_103 VPB N_VPWR_c_497_n 0.0129398f $X=-0.19 $Y=1.655 $X2=2.03 $Y2=1.49
cc_104 VPB N_VPWR_c_498_n 0.00436868f $X=-0.19 $Y=1.655 $X2=2.735 $Y2=1.245
cc_105 VPB N_VPWR_c_499_n 0.0130339f $X=-0.19 $Y=1.655 $X2=3.99 $Y2=2.375
cc_106 VPB N_VPWR_c_500_n 0.0774826f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_107 VPB N_VPWR_c_501_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_108 VPB N_VPWR_c_502_n 0.00510842f $X=-0.19 $Y=1.655 $X2=1.01 $Y2=1.49
cc_109 VPB N_VPWR_c_487_n 0.068806f $X=-0.19 $Y=1.655 $X2=1.87 $Y2=1.49
cc_110 VPB N_X_c_593_n 0.00846128f $X=-0.19 $Y=1.655 $X2=0.805 $Y2=2.465
cc_111 VPB N_X_c_594_n 0.018596f $X=-0.19 $Y=1.655 $X2=0.805 $Y2=2.465
cc_112 VPB N_X_c_595_n 0.00540935f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_113 VPB N_X_c_596_n 0.00147023f $X=-0.19 $Y=1.655 $X2=0.67 $Y2=1.49
cc_114 VPB X 0.00565f $X=-0.19 $Y=1.655 $X2=2.735 $Y2=1.405
cc_115 VPB N_A_720_367#_c_646_n 0.00258644f $X=-0.19 $Y=1.655 $X2=0.58 $Y2=1.325
cc_116 VPB N_A_720_367#_c_647_n 0.0106954f $X=-0.19 $Y=1.655 $X2=1.01 $Y2=0.665
cc_117 N_A_101_23#_M1019_g N_B1_M1006_g 0.0224156f $X=2.095 $Y=2.465 $X2=0 $Y2=0
cc_118 N_A_101_23#_c_121_n N_B1_M1006_g 0.00863021f $X=2.635 $Y=1.49 $X2=0 $Y2=0
cc_119 N_A_101_23#_c_123_n N_B1_M1006_g 0.00561163f $X=2.74 $Y=1.98 $X2=0 $Y2=0
cc_120 N_A_101_23#_c_121_n N_B1_c_247_n 0.00121584f $X=2.635 $Y=1.49 $X2=0 $Y2=0
cc_121 N_A_101_23#_c_122_n N_B1_c_247_n 0.00859058f $X=2.735 $Y=1.405 $X2=0
+ $Y2=0
cc_122 N_A_101_23#_c_124_n N_B1_c_247_n 0.00756898f $X=3.13 $Y=1.16 $X2=0 $Y2=0
cc_123 N_A_101_23#_c_126_n N_B1_c_247_n 0.0061425f $X=2.735 $Y=1.49 $X2=0 $Y2=0
cc_124 N_A_101_23#_c_121_n N_B1_c_248_n 0.00782791f $X=2.635 $Y=1.49 $X2=0 $Y2=0
cc_125 N_A_101_23#_c_127_n N_B1_c_248_n 0.0171487f $X=2.095 $Y=1.49 $X2=0 $Y2=0
cc_126 N_A_101_23#_c_133_n N_B1_M1013_g 0.0181167f $X=3.99 $Y=2.375 $X2=0 $Y2=0
cc_127 N_A_101_23#_c_122_n N_B1_M1014_g 0.00345499f $X=2.735 $Y=1.405 $X2=0
+ $Y2=0
cc_128 N_A_101_23#_c_124_n N_B1_M1014_g 0.0124292f $X=3.13 $Y=1.16 $X2=0 $Y2=0
cc_129 N_A_101_23#_c_147_p N_B1_M1014_g 0.0109256f $X=3.295 $Y=0.69 $X2=0 $Y2=0
cc_130 N_A_101_23#_c_124_n N_B1_M1021_g 0.00376278f $X=3.13 $Y=1.16 $X2=0 $Y2=0
cc_131 N_A_101_23#_c_147_p N_B1_M1021_g 0.00506691f $X=3.295 $Y=0.69 $X2=0 $Y2=0
cc_132 N_A_101_23#_c_123_n N_B1_c_251_n 0.00222432f $X=2.74 $Y=1.98 $X2=0 $Y2=0
cc_133 N_A_101_23#_c_124_n N_B1_c_251_n 0.00274768f $X=3.13 $Y=1.16 $X2=0 $Y2=0
cc_134 N_A_101_23#_c_133_n N_B1_c_251_n 8.05999e-19 $X=3.99 $Y=2.375 $X2=0 $Y2=0
cc_135 N_A_101_23#_c_126_n N_B1_c_251_n 7.59131e-19 $X=2.735 $Y=1.49 $X2=0 $Y2=0
cc_136 N_A_101_23#_c_123_n N_B1_c_255_n 0.0302846f $X=2.74 $Y=1.98 $X2=0 $Y2=0
cc_137 N_A_101_23#_c_124_n N_B1_c_255_n 0.0262508f $X=3.13 $Y=1.16 $X2=0 $Y2=0
cc_138 N_A_101_23#_c_133_n N_B1_c_255_n 0.0220843f $X=3.99 $Y=2.375 $X2=0 $Y2=0
cc_139 N_A_101_23#_c_126_n N_B1_c_255_n 0.0123333f $X=2.735 $Y=1.49 $X2=0 $Y2=0
cc_140 N_A_101_23#_c_133_n N_A3_M1015_g 0.0131906f $X=3.99 $Y=2.375 $X2=0 $Y2=0
cc_141 N_A_101_23#_c_159_p N_A3_M1015_g 0.0185264f $X=4.155 $Y=2.455 $X2=0 $Y2=0
cc_142 N_A_101_23#_c_133_n A3 0.00159973f $X=3.99 $Y=2.375 $X2=0 $Y2=0
cc_143 N_A_101_23#_c_133_n N_VPWR_M1013_d 0.00503106f $X=3.99 $Y=2.375 $X2=0
+ $Y2=0
cc_144 N_A_101_23#_M1000_g N_VPWR_c_488_n 0.0152824f $X=0.805 $Y=2.465 $X2=0
+ $Y2=0
cc_145 N_A_101_23#_M1009_g N_VPWR_c_488_n 7.27171e-19 $X=1.235 $Y=2.465 $X2=0
+ $Y2=0
cc_146 N_A_101_23#_M1000_g N_VPWR_c_489_n 7.27171e-19 $X=0.805 $Y=2.465 $X2=0
+ $Y2=0
cc_147 N_A_101_23#_M1009_g N_VPWR_c_489_n 0.0142189f $X=1.235 $Y=2.465 $X2=0
+ $Y2=0
cc_148 N_A_101_23#_M1010_g N_VPWR_c_489_n 0.0144441f $X=1.665 $Y=2.465 $X2=0
+ $Y2=0
cc_149 N_A_101_23#_M1019_g N_VPWR_c_489_n 7.42371e-19 $X=2.095 $Y=2.465 $X2=0
+ $Y2=0
cc_150 N_A_101_23#_M1010_g N_VPWR_c_490_n 0.00486043f $X=1.665 $Y=2.465 $X2=0
+ $Y2=0
cc_151 N_A_101_23#_M1019_g N_VPWR_c_490_n 0.00486043f $X=2.095 $Y=2.465 $X2=0
+ $Y2=0
cc_152 N_A_101_23#_M1010_g N_VPWR_c_491_n 8.15296e-19 $X=1.665 $Y=2.465 $X2=0
+ $Y2=0
cc_153 N_A_101_23#_M1019_g N_VPWR_c_491_n 0.0195453f $X=2.095 $Y=2.465 $X2=0
+ $Y2=0
cc_154 N_A_101_23#_c_121_n N_VPWR_c_491_n 0.0212432f $X=2.635 $Y=1.49 $X2=0
+ $Y2=0
cc_155 N_A_101_23#_c_123_n N_VPWR_c_491_n 0.0185502f $X=2.74 $Y=1.98 $X2=0 $Y2=0
cc_156 N_A_101_23#_c_127_n N_VPWR_c_491_n 6.18324e-19 $X=2.095 $Y=1.49 $X2=0
+ $Y2=0
cc_157 N_A_101_23#_c_133_n N_VPWR_c_492_n 0.0220026f $X=3.99 $Y=2.375 $X2=0
+ $Y2=0
cc_158 N_A_101_23#_c_159_p N_VPWR_c_492_n 0.0124704f $X=4.155 $Y=2.455 $X2=0
+ $Y2=0
cc_159 N_A_101_23#_M1000_g N_VPWR_c_497_n 0.00486043f $X=0.805 $Y=2.465 $X2=0
+ $Y2=0
cc_160 N_A_101_23#_M1009_g N_VPWR_c_497_n 0.00486043f $X=1.235 $Y=2.465 $X2=0
+ $Y2=0
cc_161 N_A_101_23#_c_179_p N_VPWR_c_499_n 0.0120977f $X=2.74 $Y=2.425 $X2=0
+ $Y2=0
cc_162 N_A_101_23#_c_159_p N_VPWR_c_500_n 0.0160429f $X=4.155 $Y=2.455 $X2=0
+ $Y2=0
cc_163 N_A_101_23#_M1006_s N_VPWR_c_487_n 0.00571434f $X=2.6 $Y=1.835 $X2=0
+ $Y2=0
cc_164 N_A_101_23#_M1015_s N_VPWR_c_487_n 0.00345315f $X=4.015 $Y=1.835 $X2=0
+ $Y2=0
cc_165 N_A_101_23#_M1000_g N_VPWR_c_487_n 0.00824727f $X=0.805 $Y=2.465 $X2=0
+ $Y2=0
cc_166 N_A_101_23#_M1009_g N_VPWR_c_487_n 0.00824727f $X=1.235 $Y=2.465 $X2=0
+ $Y2=0
cc_167 N_A_101_23#_M1010_g N_VPWR_c_487_n 0.00824727f $X=1.665 $Y=2.465 $X2=0
+ $Y2=0
cc_168 N_A_101_23#_M1019_g N_VPWR_c_487_n 0.00824727f $X=2.095 $Y=2.465 $X2=0
+ $Y2=0
cc_169 N_A_101_23#_c_179_p N_VPWR_c_487_n 0.00691495f $X=2.74 $Y=2.425 $X2=0
+ $Y2=0
cc_170 N_A_101_23#_c_159_p N_VPWR_c_487_n 0.0102362f $X=4.155 $Y=2.455 $X2=0
+ $Y2=0
cc_171 N_A_101_23#_M1001_g N_X_c_588_n 0.0156387f $X=0.58 $Y=0.665 $X2=0 $Y2=0
cc_172 N_A_101_23#_c_121_n N_X_c_588_n 0.0127595f $X=2.635 $Y=1.49 $X2=0 $Y2=0
cc_173 N_A_101_23#_M1000_g N_X_c_593_n 0.0152201f $X=0.805 $Y=2.465 $X2=0 $Y2=0
cc_174 N_A_101_23#_c_121_n N_X_c_593_n 0.0281744f $X=2.635 $Y=1.49 $X2=0 $Y2=0
cc_175 N_A_101_23#_c_127_n N_X_c_593_n 0.00646686f $X=2.095 $Y=1.49 $X2=0 $Y2=0
cc_176 N_A_101_23#_M1012_g N_X_c_589_n 0.0139493f $X=1.01 $Y=0.665 $X2=0 $Y2=0
cc_177 N_A_101_23#_M1016_g N_X_c_589_n 0.0136265f $X=1.44 $Y=0.665 $X2=0 $Y2=0
cc_178 N_A_101_23#_M1017_g N_X_c_589_n 0.00400533f $X=1.87 $Y=0.665 $X2=0 $Y2=0
cc_179 N_A_101_23#_c_121_n N_X_c_589_n 0.0593934f $X=2.635 $Y=1.49 $X2=0 $Y2=0
cc_180 N_A_101_23#_c_127_n N_X_c_589_n 0.00585496f $X=2.095 $Y=1.49 $X2=0 $Y2=0
cc_181 N_A_101_23#_M1009_g N_X_c_595_n 0.013227f $X=1.235 $Y=2.465 $X2=0 $Y2=0
cc_182 N_A_101_23#_M1010_g N_X_c_595_n 0.0130648f $X=1.665 $Y=2.465 $X2=0 $Y2=0
cc_183 N_A_101_23#_M1019_g N_X_c_595_n 0.00117174f $X=2.095 $Y=2.465 $X2=0 $Y2=0
cc_184 N_A_101_23#_c_121_n N_X_c_595_n 0.0593056f $X=2.635 $Y=1.49 $X2=0 $Y2=0
cc_185 N_A_101_23#_c_123_n N_X_c_595_n 0.00191072f $X=2.74 $Y=1.98 $X2=0 $Y2=0
cc_186 N_A_101_23#_c_127_n N_X_c_595_n 0.00585496f $X=2.095 $Y=1.49 $X2=0 $Y2=0
cc_187 N_A_101_23#_c_121_n N_X_c_590_n 0.014687f $X=2.635 $Y=1.49 $X2=0 $Y2=0
cc_188 N_A_101_23#_c_127_n N_X_c_590_n 0.00298081f $X=2.095 $Y=1.49 $X2=0 $Y2=0
cc_189 N_A_101_23#_c_121_n N_X_c_596_n 0.014687f $X=2.635 $Y=1.49 $X2=0 $Y2=0
cc_190 N_A_101_23#_c_127_n N_X_c_596_n 0.00298081f $X=2.095 $Y=1.49 $X2=0 $Y2=0
cc_191 N_A_101_23#_M1001_g X 0.00704142f $X=0.58 $Y=0.665 $X2=0 $Y2=0
cc_192 N_A_101_23#_M1000_g X 0.00279639f $X=0.805 $Y=2.465 $X2=0 $Y2=0
cc_193 N_A_101_23#_c_121_n X 0.0138088f $X=2.635 $Y=1.49 $X2=0 $Y2=0
cc_194 N_A_101_23#_c_127_n X 0.00469505f $X=2.095 $Y=1.49 $X2=0 $Y2=0
cc_195 N_A_101_23#_c_133_n N_A_720_367#_M1015_d 0.0109432f $X=3.99 $Y=2.375
+ $X2=-0.19 $Y2=-0.245
cc_196 N_A_101_23#_M1015_s N_A_720_367#_c_646_n 0.00334509f $X=4.015 $Y=1.835
+ $X2=0 $Y2=0
cc_197 N_A_101_23#_c_133_n N_A_720_367#_c_646_n 0.0268549f $X=3.99 $Y=2.375
+ $X2=0 $Y2=0
cc_198 N_A_101_23#_c_159_p N_A_720_367#_c_646_n 0.0155387f $X=4.155 $Y=2.455
+ $X2=0 $Y2=0
cc_199 N_A_101_23#_M1001_g N_VGND_c_709_n 0.0120262f $X=0.58 $Y=0.665 $X2=0
+ $Y2=0
cc_200 N_A_101_23#_M1012_g N_VGND_c_709_n 6.10117e-19 $X=1.01 $Y=0.665 $X2=0
+ $Y2=0
cc_201 N_A_101_23#_M1001_g N_VGND_c_710_n 6.10117e-19 $X=0.58 $Y=0.665 $X2=0
+ $Y2=0
cc_202 N_A_101_23#_M1012_g N_VGND_c_710_n 0.0110386f $X=1.01 $Y=0.665 $X2=0
+ $Y2=0
cc_203 N_A_101_23#_M1016_g N_VGND_c_710_n 0.0110386f $X=1.44 $Y=0.665 $X2=0
+ $Y2=0
cc_204 N_A_101_23#_M1017_g N_VGND_c_710_n 6.10117e-19 $X=1.87 $Y=0.665 $X2=0
+ $Y2=0
cc_205 N_A_101_23#_M1016_g N_VGND_c_711_n 6.8136e-19 $X=1.44 $Y=0.665 $X2=0
+ $Y2=0
cc_206 N_A_101_23#_M1017_g N_VGND_c_711_n 0.017606f $X=1.87 $Y=0.665 $X2=0 $Y2=0
cc_207 N_A_101_23#_c_121_n N_VGND_c_711_n 0.0174641f $X=2.635 $Y=1.49 $X2=0
+ $Y2=0
cc_208 N_A_101_23#_c_125_n N_VGND_c_711_n 0.00150507f $X=2.835 $Y=1.16 $X2=0
+ $Y2=0
cc_209 N_A_101_23#_c_127_n N_VGND_c_711_n 0.00679686f $X=2.095 $Y=1.49 $X2=0
+ $Y2=0
cc_210 N_A_101_23#_M1001_g N_VGND_c_715_n 0.00477554f $X=0.58 $Y=0.665 $X2=0
+ $Y2=0
cc_211 N_A_101_23#_M1012_g N_VGND_c_715_n 0.00477554f $X=1.01 $Y=0.665 $X2=0
+ $Y2=0
cc_212 N_A_101_23#_M1016_g N_VGND_c_716_n 0.00477554f $X=1.44 $Y=0.665 $X2=0
+ $Y2=0
cc_213 N_A_101_23#_M1017_g N_VGND_c_716_n 0.00477554f $X=1.87 $Y=0.665 $X2=0
+ $Y2=0
cc_214 N_A_101_23#_M1001_g N_VGND_c_721_n 0.00825815f $X=0.58 $Y=0.665 $X2=0
+ $Y2=0
cc_215 N_A_101_23#_M1012_g N_VGND_c_721_n 0.00825815f $X=1.01 $Y=0.665 $X2=0
+ $Y2=0
cc_216 N_A_101_23#_M1016_g N_VGND_c_721_n 0.00825815f $X=1.44 $Y=0.665 $X2=0
+ $Y2=0
cc_217 N_A_101_23#_M1017_g N_VGND_c_721_n 0.00825815f $X=1.87 $Y=0.665 $X2=0
+ $Y2=0
cc_218 N_A_101_23#_c_124_n N_A_528_65#_M1014_s 0.00119058f $X=3.13 $Y=1.16
+ $X2=-0.19 $Y2=-0.245
cc_219 N_A_101_23#_c_125_n N_A_528_65#_M1014_s 0.00307898f $X=2.835 $Y=1.16
+ $X2=-0.19 $Y2=-0.245
cc_220 N_A_101_23#_M1017_g N_A_528_65#_c_808_n 0.00128166f $X=1.87 $Y=0.665
+ $X2=0 $Y2=0
cc_221 N_A_101_23#_c_121_n N_A_528_65#_c_808_n 4.89368e-19 $X=2.635 $Y=1.49
+ $X2=0 $Y2=0
cc_222 N_A_101_23#_c_124_n N_A_528_65#_c_808_n 0.00912321f $X=3.13 $Y=1.16 $X2=0
+ $Y2=0
cc_223 N_A_101_23#_c_125_n N_A_528_65#_c_808_n 0.0179692f $X=2.835 $Y=1.16 $X2=0
+ $Y2=0
cc_224 N_A_101_23#_M1014_d N_A_528_65#_c_809_n 0.00176773f $X=3.155 $Y=0.325
+ $X2=0 $Y2=0
cc_225 N_A_101_23#_c_124_n N_A_528_65#_c_809_n 0.00281285f $X=3.13 $Y=1.16 $X2=0
+ $Y2=0
cc_226 N_A_101_23#_c_147_p N_A_528_65#_c_809_n 0.0160064f $X=3.295 $Y=0.69 $X2=0
+ $Y2=0
cc_227 N_A_101_23#_c_124_n N_A_528_65#_c_812_n 0.0108938f $X=3.13 $Y=1.16 $X2=0
+ $Y2=0
cc_228 N_B1_M1021_g N_A3_M1003_g 0.0139331f $X=3.51 $Y=0.745 $X2=0 $Y2=0
cc_229 N_B1_c_255_n N_A3_M1015_g 0.00364557f $X=3.17 $Y=1.51 $X2=0 $Y2=0
cc_230 N_B1_M1013_g A3 3.07252e-19 $X=2.955 $Y=2.465 $X2=0 $Y2=0
cc_231 N_B1_c_251_n A3 0.00888341f $X=3.17 $Y=1.51 $X2=0 $Y2=0
cc_232 N_B1_c_255_n A3 0.0260862f $X=3.17 $Y=1.51 $X2=0 $Y2=0
cc_233 N_B1_c_251_n N_A3_c_308_n 0.0169716f $X=3.17 $Y=1.51 $X2=0 $Y2=0
cc_234 N_B1_c_255_n N_VPWR_M1013_d 0.00355574f $X=3.17 $Y=1.51 $X2=0 $Y2=0
cc_235 N_B1_M1006_g N_VPWR_c_491_n 0.019536f $X=2.525 $Y=2.465 $X2=0 $Y2=0
cc_236 N_B1_M1013_g N_VPWR_c_491_n 6.24191e-19 $X=2.955 $Y=2.465 $X2=0 $Y2=0
cc_237 N_B1_M1006_g N_VPWR_c_492_n 5.82718e-19 $X=2.525 $Y=2.465 $X2=0 $Y2=0
cc_238 N_B1_M1013_g N_VPWR_c_492_n 0.0130411f $X=2.955 $Y=2.465 $X2=0 $Y2=0
cc_239 N_B1_M1006_g N_VPWR_c_499_n 0.00486043f $X=2.525 $Y=2.465 $X2=0 $Y2=0
cc_240 N_B1_M1013_g N_VPWR_c_499_n 0.00486043f $X=2.955 $Y=2.465 $X2=0 $Y2=0
cc_241 N_B1_M1006_g N_VPWR_c_487_n 0.00824727f $X=2.525 $Y=2.465 $X2=0 $Y2=0
cc_242 N_B1_M1013_g N_VPWR_c_487_n 0.00824727f $X=2.955 $Y=2.465 $X2=0 $Y2=0
cc_243 N_B1_M1013_g N_A_720_367#_c_646_n 8.43086e-19 $X=2.955 $Y=2.465 $X2=0
+ $Y2=0
cc_244 N_B1_c_255_n N_A_720_367#_c_646_n 0.0143828f $X=3.17 $Y=1.51 $X2=0 $Y2=0
cc_245 N_B1_M1021_g N_VGND_c_712_n 5.18213e-19 $X=3.51 $Y=0.745 $X2=0 $Y2=0
cc_246 N_B1_M1014_g N_VGND_c_717_n 0.00302501f $X=3.08 $Y=0.745 $X2=0 $Y2=0
cc_247 N_B1_M1021_g N_VGND_c_717_n 0.00302501f $X=3.51 $Y=0.745 $X2=0 $Y2=0
cc_248 N_B1_M1014_g N_VGND_c_721_n 0.0048466f $X=3.08 $Y=0.745 $X2=0 $Y2=0
cc_249 N_B1_M1021_g N_VGND_c_721_n 0.00435646f $X=3.51 $Y=0.745 $X2=0 $Y2=0
cc_250 N_B1_c_247_n N_A_528_65#_c_808_n 0.00142201f $X=2.88 $Y=1.42 $X2=0 $Y2=0
cc_251 N_B1_M1014_g N_A_528_65#_c_809_n 0.0131978f $X=3.08 $Y=0.745 $X2=0 $Y2=0
cc_252 N_B1_M1021_g N_A_528_65#_c_809_n 0.0121029f $X=3.51 $Y=0.745 $X2=0 $Y2=0
cc_253 N_B1_M1021_g N_A_528_65#_c_812_n 6.54275e-19 $X=3.51 $Y=0.745 $X2=0 $Y2=0
cc_254 N_A3_M1018_g N_A2_M1002_g 0.0181721f $X=4.37 $Y=0.745 $X2=0 $Y2=0
cc_255 N_A3_M1023_g N_A2_M1007_g 0.0181721f $X=4.37 $Y=2.465 $X2=0 $Y2=0
cc_256 A3 N_A2_c_362_n 0.00290837f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_257 N_A3_c_308_n N_A2_c_362_n 0.0181721f $X=4.37 $Y=1.51 $X2=0 $Y2=0
cc_258 A3 N_A2_c_363_n 0.0235673f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_259 N_A3_c_308_n N_A2_c_363_n 6.58083e-19 $X=4.37 $Y=1.51 $X2=0 $Y2=0
cc_260 A3 N_A2_c_370_n 0.00392223f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_261 N_A3_M1015_g N_VPWR_c_492_n 0.0094741f $X=3.94 $Y=2.465 $X2=0 $Y2=0
cc_262 N_A3_M1015_g N_VPWR_c_500_n 0.0054895f $X=3.94 $Y=2.465 $X2=0 $Y2=0
cc_263 N_A3_M1023_g N_VPWR_c_500_n 0.00564131f $X=4.37 $Y=2.465 $X2=0 $Y2=0
cc_264 N_A3_M1015_g N_VPWR_c_487_n 0.0114203f $X=3.94 $Y=2.465 $X2=0 $Y2=0
cc_265 N_A3_M1023_g N_VPWR_c_487_n 0.0103088f $X=4.37 $Y=2.465 $X2=0 $Y2=0
cc_266 N_A3_M1015_g N_A_720_367#_c_646_n 0.00925001f $X=3.94 $Y=2.465 $X2=0
+ $Y2=0
cc_267 N_A3_M1023_g N_A_720_367#_c_646_n 0.01275f $X=4.37 $Y=2.465 $X2=0 $Y2=0
cc_268 A3 N_A_720_367#_c_646_n 0.060264f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_269 N_A3_c_308_n N_A_720_367#_c_646_n 5.8554e-19 $X=4.37 $Y=1.51 $X2=0 $Y2=0
cc_270 N_A3_M1015_g N_A_720_367#_c_658_n 2.44839e-19 $X=3.94 $Y=2.465 $X2=0
+ $Y2=0
cc_271 N_A3_M1023_g N_A_720_367#_c_658_n 0.0089023f $X=4.37 $Y=2.465 $X2=0 $Y2=0
cc_272 N_A3_M1015_g N_A_720_367#_c_660_n 6.77146e-19 $X=3.94 $Y=2.465 $X2=0
+ $Y2=0
cc_273 N_A3_M1023_g N_A_720_367#_c_660_n 0.00369808f $X=4.37 $Y=2.465 $X2=0
+ $Y2=0
cc_274 A3 N_A_720_367#_c_660_n 0.0184068f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_275 N_A3_M1003_g N_VGND_c_712_n 0.0100743f $X=3.94 $Y=0.745 $X2=0 $Y2=0
cc_276 N_A3_M1018_g N_VGND_c_712_n 0.0101563f $X=4.37 $Y=0.745 $X2=0 $Y2=0
cc_277 N_A3_M1003_g N_VGND_c_717_n 0.00414769f $X=3.94 $Y=0.745 $X2=0 $Y2=0
cc_278 N_A3_M1018_g N_VGND_c_718_n 0.00414769f $X=4.37 $Y=0.745 $X2=0 $Y2=0
cc_279 N_A3_M1003_g N_VGND_c_721_n 0.0078848f $X=3.94 $Y=0.745 $X2=0 $Y2=0
cc_280 N_A3_M1018_g N_VGND_c_721_n 0.0078848f $X=4.37 $Y=0.745 $X2=0 $Y2=0
cc_281 N_A3_M1003_g N_A_528_65#_c_809_n 5.73473e-19 $X=3.94 $Y=0.745 $X2=0 $Y2=0
cc_282 N_A3_M1003_g N_A_528_65#_c_811_n 0.0130281f $X=3.94 $Y=0.745 $X2=0 $Y2=0
cc_283 N_A3_M1018_g N_A_528_65#_c_811_n 0.0130709f $X=4.37 $Y=0.745 $X2=0 $Y2=0
cc_284 A3 N_A_528_65#_c_811_n 0.0473477f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_285 N_A3_c_308_n N_A_528_65#_c_811_n 0.00244902f $X=4.37 $Y=1.51 $X2=0 $Y2=0
cc_286 A3 N_A_528_65#_c_812_n 0.0161224f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_287 N_A3_M1018_g N_A_528_65#_c_813_n 8.32918e-19 $X=4.37 $Y=0.745 $X2=0 $Y2=0
cc_288 A3 N_A_528_65#_c_817_n 0.0161224f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_289 N_A2_M1002_g N_A1_c_433_n 0.0268432f $X=4.8 $Y=0.745 $X2=-0.19 $Y2=-0.245
cc_290 N_A2_M1007_g N_A1_M1005_g 0.0366562f $X=4.8 $Y=2.465 $X2=0 $Y2=0
cc_291 N_A2_c_366_n N_A1_M1005_g 0.0119949f $X=6.265 $Y=1.79 $X2=0 $Y2=0
cc_292 N_A2_M1004_g N_A1_c_435_n 0.0363037f $X=6.245 $Y=0.745 $X2=0 $Y2=0
cc_293 N_A2_M1020_g N_A1_M1011_g 0.0363037f $X=6.245 $Y=2.465 $X2=0 $Y2=0
cc_294 N_A2_c_366_n N_A1_M1011_g 0.010446f $X=6.265 $Y=1.79 $X2=0 $Y2=0
cc_295 N_A2_M1002_g A1 6.09533e-19 $X=4.8 $Y=0.745 $X2=0 $Y2=0
cc_296 N_A2_M1004_g A1 0.00470067f $X=6.245 $Y=0.745 $X2=0 $Y2=0
cc_297 N_A2_c_366_n A1 0.0540168f $X=6.265 $Y=1.79 $X2=0 $Y2=0
cc_298 N_A2_c_360_n A1 0.0202492f $X=6.43 $Y=1.46 $X2=0 $Y2=0
cc_299 N_A2_c_363_n A1 0.0160159f $X=4.935 $Y=1.51 $X2=0 $Y2=0
cc_300 N_A2_c_366_n N_A1_c_438_n 0.00243542f $X=6.265 $Y=1.79 $X2=0 $Y2=0
cc_301 N_A2_c_360_n N_A1_c_438_n 0.00111997f $X=6.43 $Y=1.46 $X2=0 $Y2=0
cc_302 N_A2_c_361_n N_A1_c_438_n 0.0363037f $X=6.43 $Y=1.46 $X2=0 $Y2=0
cc_303 N_A2_c_362_n N_A1_c_438_n 0.0208961f $X=4.935 $Y=1.51 $X2=0 $Y2=0
cc_304 N_A2_c_363_n N_A1_c_438_n 0.00571114f $X=4.935 $Y=1.51 $X2=0 $Y2=0
cc_305 N_A2_c_366_n N_VPWR_M1005_s 0.00176891f $X=6.265 $Y=1.79 $X2=0 $Y2=0
cc_306 N_A2_M1020_g N_VPWR_c_493_n 0.0158617f $X=6.245 $Y=2.465 $X2=0 $Y2=0
cc_307 N_A2_M1020_g N_VPWR_c_494_n 0.0128934f $X=6.245 $Y=2.465 $X2=0 $Y2=0
cc_308 N_A2_M1007_g N_VPWR_c_500_n 0.0054895f $X=4.8 $Y=2.465 $X2=0 $Y2=0
cc_309 N_A2_M1020_g N_VPWR_c_500_n 0.00417534f $X=6.245 $Y=2.465 $X2=0 $Y2=0
cc_310 N_A2_M1007_g N_VPWR_c_487_n 0.0104266f $X=4.8 $Y=2.465 $X2=0 $Y2=0
cc_311 N_A2_M1020_g N_VPWR_c_487_n 0.0067963f $X=6.245 $Y=2.465 $X2=0 $Y2=0
cc_312 N_A2_c_366_n N_A_720_367#_M1020_s 0.00248446f $X=6.265 $Y=1.79 $X2=0
+ $Y2=0
cc_313 N_A2_M1007_g N_A_720_367#_c_658_n 0.0113228f $X=4.8 $Y=2.465 $X2=0 $Y2=0
cc_314 N_A2_M1007_g N_A_720_367#_c_647_n 0.016678f $X=4.8 $Y=2.465 $X2=0 $Y2=0
cc_315 N_A2_M1020_g N_A_720_367#_c_647_n 0.00971117f $X=6.245 $Y=2.465 $X2=0
+ $Y2=0
cc_316 N_A2_c_366_n N_A_720_367#_c_647_n 0.0773291f $X=6.265 $Y=1.79 $X2=0 $Y2=0
cc_317 N_A2_c_361_n N_A_720_367#_c_647_n 0.00103682f $X=6.43 $Y=1.46 $X2=0 $Y2=0
cc_318 N_A2_c_362_n N_A_720_367#_c_647_n 9.21299e-19 $X=4.935 $Y=1.51 $X2=0
+ $Y2=0
cc_319 N_A2_c_370_n N_A_720_367#_c_647_n 0.0246518f $X=5.027 $Y=1.705 $X2=0
+ $Y2=0
cc_320 N_A2_M1007_g N_A_720_367#_c_660_n 0.00499989f $X=4.8 $Y=2.465 $X2=0 $Y2=0
cc_321 N_A2_c_366_n N_A_975_367#_M1007_d 5.00837e-19 $X=6.265 $Y=1.79 $X2=-0.19
+ $Y2=-0.245
cc_322 N_A2_c_370_n N_A_975_367#_M1007_d 0.00307759f $X=5.027 $Y=1.705 $X2=-0.19
+ $Y2=-0.245
cc_323 N_A2_c_366_n N_A_975_367#_M1011_d 0.00176891f $X=6.265 $Y=1.79 $X2=0
+ $Y2=0
cc_324 N_A2_M1020_g N_A_975_367#_c_692_n 0.0030857f $X=6.245 $Y=2.465 $X2=0
+ $Y2=0
cc_325 N_A2_M1002_g N_VGND_c_712_n 6.04191e-19 $X=4.8 $Y=0.745 $X2=0 $Y2=0
cc_326 N_A2_M1002_g N_VGND_c_713_n 0.00410592f $X=4.8 $Y=0.745 $X2=0 $Y2=0
cc_327 N_A2_M1004_g N_VGND_c_714_n 0.010633f $X=6.245 $Y=0.745 $X2=0 $Y2=0
cc_328 N_A2_M1002_g N_VGND_c_718_n 0.0046928f $X=4.8 $Y=0.745 $X2=0 $Y2=0
cc_329 N_A2_M1004_g N_VGND_c_720_n 0.00414769f $X=6.245 $Y=0.745 $X2=0 $Y2=0
cc_330 N_A2_M1002_g N_VGND_c_721_n 0.009055f $X=4.8 $Y=0.745 $X2=0 $Y2=0
cc_331 N_A2_M1004_g N_VGND_c_721_n 0.00823375f $X=6.245 $Y=0.745 $X2=0 $Y2=0
cc_332 N_A2_M1002_g N_A_528_65#_c_813_n 0.00940481f $X=4.8 $Y=0.745 $X2=0 $Y2=0
cc_333 N_A2_M1002_g N_A_528_65#_c_841_n 0.014872f $X=4.8 $Y=0.745 $X2=0 $Y2=0
cc_334 N_A2_c_366_n N_A_528_65#_c_841_n 0.00354498f $X=6.265 $Y=1.79 $X2=0 $Y2=0
cc_335 N_A2_c_362_n N_A_528_65#_c_841_n 0.00123765f $X=4.935 $Y=1.51 $X2=0 $Y2=0
cc_336 N_A2_c_363_n N_A_528_65#_c_841_n 0.0163082f $X=4.935 $Y=1.51 $X2=0 $Y2=0
cc_337 N_A2_M1002_g N_A_528_65#_c_814_n 8.50177e-19 $X=4.8 $Y=0.745 $X2=0 $Y2=0
cc_338 N_A2_M1004_g N_A_528_65#_c_815_n 0.0136418f $X=6.245 $Y=0.745 $X2=0 $Y2=0
cc_339 N_A2_c_366_n N_A_528_65#_c_815_n 0.00337347f $X=6.265 $Y=1.79 $X2=0 $Y2=0
cc_340 N_A2_c_360_n N_A_528_65#_c_815_n 0.018314f $X=6.43 $Y=1.46 $X2=0 $Y2=0
cc_341 N_A2_c_361_n N_A_528_65#_c_815_n 0.00168047f $X=6.43 $Y=1.46 $X2=0 $Y2=0
cc_342 N_A2_M1004_g N_A_528_65#_c_816_n 7.37323e-19 $X=6.245 $Y=0.745 $X2=0
+ $Y2=0
cc_343 N_A2_M1002_g N_A_528_65#_c_817_n 0.00373571f $X=4.8 $Y=0.745 $X2=0 $Y2=0
cc_344 N_A1_M1005_g N_VPWR_c_493_n 0.00345954f $X=5.385 $Y=2.465 $X2=0 $Y2=0
cc_345 N_A1_M1011_g N_VPWR_c_493_n 0.00997209f $X=5.815 $Y=2.465 $X2=0 $Y2=0
cc_346 N_A1_M1005_g N_VPWR_c_500_n 0.00357877f $X=5.385 $Y=2.465 $X2=0 $Y2=0
cc_347 N_A1_M1011_g N_VPWR_c_500_n 0.00357877f $X=5.815 $Y=2.465 $X2=0 $Y2=0
cc_348 N_A1_M1005_g N_VPWR_c_487_n 0.00580255f $X=5.385 $Y=2.465 $X2=0 $Y2=0
cc_349 N_A1_M1011_g N_VPWR_c_487_n 0.00537654f $X=5.815 $Y=2.465 $X2=0 $Y2=0
cc_350 N_A1_M1005_g N_A_720_367#_c_658_n 0.00100584f $X=5.385 $Y=2.465 $X2=0
+ $Y2=0
cc_351 N_A1_M1005_g N_A_720_367#_c_647_n 0.0148595f $X=5.385 $Y=2.465 $X2=0
+ $Y2=0
cc_352 N_A1_M1011_g N_A_720_367#_c_647_n 0.0123792f $X=5.815 $Y=2.465 $X2=0
+ $Y2=0
cc_353 N_A1_M1005_g N_A_720_367#_c_660_n 5.61804e-19 $X=5.385 $Y=2.465 $X2=0
+ $Y2=0
cc_354 N_A1_M1005_g N_A_975_367#_c_692_n 0.0145913f $X=5.385 $Y=2.465 $X2=0
+ $Y2=0
cc_355 N_A1_M1011_g N_A_975_367#_c_692_n 0.0095355f $X=5.815 $Y=2.465 $X2=0
+ $Y2=0
cc_356 N_A1_c_433_n N_VGND_c_713_n 0.00407067f $X=5.385 $Y=1.275 $X2=0 $Y2=0
cc_357 N_A1_c_433_n N_VGND_c_714_n 4.8425e-19 $X=5.385 $Y=1.275 $X2=0 $Y2=0
cc_358 N_A1_c_435_n N_VGND_c_714_n 0.00857476f $X=5.815 $Y=1.275 $X2=0 $Y2=0
cc_359 N_A1_c_433_n N_VGND_c_719_n 0.0046928f $X=5.385 $Y=1.275 $X2=0 $Y2=0
cc_360 N_A1_c_435_n N_VGND_c_719_n 0.00414769f $X=5.815 $Y=1.275 $X2=0 $Y2=0
cc_361 N_A1_c_433_n N_VGND_c_721_n 0.00905646f $X=5.385 $Y=1.275 $X2=0 $Y2=0
cc_362 N_A1_c_435_n N_VGND_c_721_n 0.00787505f $X=5.815 $Y=1.275 $X2=0 $Y2=0
cc_363 N_A1_c_433_n N_A_528_65#_c_813_n 8.48075e-19 $X=5.385 $Y=1.275 $X2=0
+ $Y2=0
cc_364 N_A1_c_433_n N_A_528_65#_c_841_n 0.0126765f $X=5.385 $Y=1.275 $X2=0 $Y2=0
cc_365 A1 N_A_528_65#_c_841_n 0.00424561f $X=5.915 $Y=1.21 $X2=0 $Y2=0
cc_366 N_A1_c_433_n N_A_528_65#_c_814_n 0.00809758f $X=5.385 $Y=1.275 $X2=0
+ $Y2=0
cc_367 N_A1_c_435_n N_A_528_65#_c_814_n 2.09864e-19 $X=5.815 $Y=1.275 $X2=0
+ $Y2=0
cc_368 N_A1_c_435_n N_A_528_65#_c_815_n 0.0120489f $X=5.815 $Y=1.275 $X2=0 $Y2=0
cc_369 A1 N_A_528_65#_c_815_n 0.0264244f $X=5.915 $Y=1.21 $X2=0 $Y2=0
cc_370 A1 N_A_528_65#_c_817_n 0.00105878f $X=5.915 $Y=1.21 $X2=0 $Y2=0
cc_371 N_A1_c_433_n N_A_528_65#_c_860_n 7.32094e-19 $X=5.385 $Y=1.275 $X2=0
+ $Y2=0
cc_372 A1 N_A_528_65#_c_860_n 0.019204f $X=5.915 $Y=1.21 $X2=0 $Y2=0
cc_373 N_A1_c_438_n N_A_528_65#_c_860_n 6.68767e-19 $X=5.815 $Y=1.44 $X2=0 $Y2=0
cc_374 N_VPWR_c_487_n N_X_M1000_s 0.00536646f $X=6.48 $Y=3.33 $X2=0 $Y2=0
cc_375 N_VPWR_c_487_n N_X_M1010_s 0.00571434f $X=6.48 $Y=3.33 $X2=0 $Y2=0
cc_376 N_VPWR_M1000_d N_X_c_593_n 0.00262981f $X=0.465 $Y=1.835 $X2=0 $Y2=0
cc_377 N_VPWR_c_488_n N_X_c_593_n 0.0220026f $X=0.59 $Y=2.18 $X2=0 $Y2=0
cc_378 N_VPWR_c_497_n N_X_c_626_n 0.0124525f $X=1.285 $Y=3.33 $X2=0 $Y2=0
cc_379 N_VPWR_c_487_n N_X_c_626_n 0.00730901f $X=6.48 $Y=3.33 $X2=0 $Y2=0
cc_380 N_VPWR_M1009_d N_X_c_595_n 0.00176461f $X=1.31 $Y=1.835 $X2=0 $Y2=0
cc_381 N_VPWR_c_489_n N_X_c_595_n 0.0170777f $X=1.45 $Y=2.18 $X2=0 $Y2=0
cc_382 N_VPWR_c_491_n N_X_c_595_n 0.00503283f $X=2.31 $Y=1.98 $X2=0 $Y2=0
cc_383 N_VPWR_c_490_n N_X_c_631_n 0.0120977f $X=2.145 $Y=3.33 $X2=0 $Y2=0
cc_384 N_VPWR_c_487_n N_X_c_631_n 0.00691495f $X=6.48 $Y=3.33 $X2=0 $Y2=0
cc_385 N_VPWR_c_487_n N_A_720_367#_M1015_d 0.0113783f $X=6.48 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_386 N_VPWR_c_487_n N_A_720_367#_M1023_d 0.00223559f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_387 N_VPWR_c_493_n N_A_720_367#_M1020_s 0.00338954f $X=6.365 $Y=2.55 $X2=0
+ $Y2=0
cc_388 N_VPWR_c_494_n N_A_720_367#_M1020_s 0.00372718f $X=6.495 $Y=3.245 $X2=0
+ $Y2=0
cc_389 N_VPWR_c_487_n N_A_720_367#_M1020_s 5.30836e-19 $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_390 N_VPWR_c_500_n N_A_720_367#_c_658_n 0.0182419f $X=6.365 $Y=3.33 $X2=0
+ $Y2=0
cc_391 N_VPWR_c_487_n N_A_720_367#_c_658_n 0.0120429f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_392 N_VPWR_M1005_s N_A_720_367#_c_647_n 0.00342759f $X=5.46 $Y=1.835 $X2=0
+ $Y2=0
cc_393 N_VPWR_c_493_n N_A_720_367#_c_647_n 0.0694076f $X=6.365 $Y=2.55 $X2=0
+ $Y2=0
cc_394 N_VPWR_c_487_n N_A_975_367#_M1007_d 0.00526276f $X=6.48 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_395 N_VPWR_c_493_n N_A_975_367#_M1011_d 0.00351073f $X=6.365 $Y=2.55 $X2=0
+ $Y2=0
cc_396 N_VPWR_c_487_n N_A_975_367#_M1011_d 0.00223577f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_397 N_VPWR_c_500_n N_A_975_367#_c_698_n 0.0227896f $X=6.365 $Y=3.33 $X2=0
+ $Y2=0
cc_398 N_VPWR_c_487_n N_A_975_367#_c_698_n 0.0127935f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_399 N_VPWR_M1005_s N_A_975_367#_c_692_n 0.00336331f $X=5.46 $Y=1.835 $X2=0
+ $Y2=0
cc_400 N_VPWR_c_493_n N_A_975_367#_c_692_n 0.0382539f $X=6.365 $Y=2.55 $X2=0
+ $Y2=0
cc_401 N_VPWR_c_500_n N_A_975_367#_c_692_n 0.0519195f $X=6.365 $Y=3.33 $X2=0
+ $Y2=0
cc_402 N_VPWR_c_487_n N_A_975_367#_c_692_n 0.0339791f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_403 N_X_c_588_n N_VGND_M1001_s 0.00119058f $X=0.7 $Y=1.14 $X2=-0.19
+ $Y2=-0.245
cc_404 N_X_c_591_n N_VGND_M1001_s 0.00119244f $X=0.21 $Y=1.225 $X2=-0.19
+ $Y2=-0.245
cc_405 N_X_c_589_n N_VGND_M1012_s 0.00176461f $X=1.56 $Y=1.14 $X2=0 $Y2=0
cc_406 N_X_c_588_n N_VGND_c_709_n 0.0109431f $X=0.7 $Y=1.14 $X2=0 $Y2=0
cc_407 N_X_c_591_n N_VGND_c_709_n 0.0122196f $X=0.21 $Y=1.225 $X2=0 $Y2=0
cc_408 N_X_c_589_n N_VGND_c_710_n 0.0170777f $X=1.56 $Y=1.14 $X2=0 $Y2=0
cc_409 N_X_c_589_n N_VGND_c_711_n 0.0027708f $X=1.56 $Y=1.14 $X2=0 $Y2=0
cc_410 N_X_c_640_p N_VGND_c_715_n 0.0124525f $X=0.795 $Y=0.42 $X2=0 $Y2=0
cc_411 N_X_c_641_p N_VGND_c_716_n 0.0124525f $X=1.655 $Y=0.42 $X2=0 $Y2=0
cc_412 N_X_M1001_d N_VGND_c_721_n 0.00536646f $X=0.655 $Y=0.245 $X2=0 $Y2=0
cc_413 N_X_M1016_d N_VGND_c_721_n 0.00536646f $X=1.515 $Y=0.245 $X2=0 $Y2=0
cc_414 N_X_c_640_p N_VGND_c_721_n 0.00730901f $X=0.795 $Y=0.42 $X2=0 $Y2=0
cc_415 N_X_c_641_p N_VGND_c_721_n 0.00730901f $X=1.655 $Y=0.42 $X2=0 $Y2=0
cc_416 N_A_720_367#_c_647_n N_A_975_367#_M1007_d 0.00751329f $X=6.46 $Y=2.16
+ $X2=-0.19 $Y2=1.655
cc_417 N_A_720_367#_c_647_n N_A_975_367#_M1011_d 0.00356607f $X=6.46 $Y=2.16
+ $X2=0 $Y2=0
cc_418 N_A_720_367#_c_647_n N_A_975_367#_c_706_n 0.0264484f $X=6.46 $Y=2.16
+ $X2=0 $Y2=0
cc_419 N_A_720_367#_c_647_n N_A_975_367#_c_692_n 0.00301506f $X=6.46 $Y=2.16
+ $X2=0 $Y2=0
cc_420 N_VGND_c_711_n N_A_528_65#_c_808_n 0.0228401f $X=2.085 $Y=0.39 $X2=0
+ $Y2=0
cc_421 N_VGND_c_712_n N_A_528_65#_c_809_n 0.0100029f $X=4.155 $Y=0.45 $X2=0
+ $Y2=0
cc_422 N_VGND_c_717_n N_A_528_65#_c_809_n 0.0566591f $X=3.99 $Y=0 $X2=0 $Y2=0
cc_423 N_VGND_c_721_n N_A_528_65#_c_809_n 0.0316105f $X=6.48 $Y=0 $X2=0 $Y2=0
cc_424 N_VGND_c_711_n N_A_528_65#_c_810_n 0.00928107f $X=2.085 $Y=0.39 $X2=0
+ $Y2=0
cc_425 N_VGND_c_717_n N_A_528_65#_c_810_n 0.0235763f $X=3.99 $Y=0 $X2=0 $Y2=0
cc_426 N_VGND_c_721_n N_A_528_65#_c_810_n 0.0128145f $X=6.48 $Y=0 $X2=0 $Y2=0
cc_427 N_VGND_M1003_d N_A_528_65#_c_811_n 0.00180746f $X=4.015 $Y=0.325 $X2=0
+ $Y2=0
cc_428 N_VGND_c_712_n N_A_528_65#_c_811_n 0.0163515f $X=4.155 $Y=0.45 $X2=0
+ $Y2=0
cc_429 N_VGND_c_712_n N_A_528_65#_c_813_n 0.0219626f $X=4.155 $Y=0.45 $X2=0
+ $Y2=0
cc_430 N_VGND_c_713_n N_A_528_65#_c_813_n 0.0147356f $X=5.09 $Y=0.565 $X2=0
+ $Y2=0
cc_431 N_VGND_c_718_n N_A_528_65#_c_813_n 0.0139581f $X=4.925 $Y=0 $X2=0 $Y2=0
cc_432 N_VGND_c_721_n N_A_528_65#_c_813_n 0.00966529f $X=6.48 $Y=0 $X2=0 $Y2=0
cc_433 N_VGND_M1002_d N_A_528_65#_c_841_n 0.00845026f $X=4.875 $Y=0.325 $X2=0
+ $Y2=0
cc_434 N_VGND_c_713_n N_A_528_65#_c_841_n 0.0261161f $X=5.09 $Y=0.565 $X2=0
+ $Y2=0
cc_435 N_VGND_c_713_n N_A_528_65#_c_814_n 0.0144087f $X=5.09 $Y=0.565 $X2=0
+ $Y2=0
cc_436 N_VGND_c_714_n N_A_528_65#_c_814_n 0.0155838f $X=6.03 $Y=0.47 $X2=0 $Y2=0
cc_437 N_VGND_c_719_n N_A_528_65#_c_814_n 0.0139581f $X=5.865 $Y=0 $X2=0 $Y2=0
cc_438 N_VGND_c_721_n N_A_528_65#_c_814_n 0.00966529f $X=6.48 $Y=0 $X2=0 $Y2=0
cc_439 N_VGND_M1022_s N_A_528_65#_c_815_n 0.0037201f $X=5.89 $Y=0.325 $X2=0
+ $Y2=0
cc_440 N_VGND_c_714_n N_A_528_65#_c_815_n 0.0171619f $X=6.03 $Y=0.47 $X2=0 $Y2=0
cc_441 N_VGND_c_714_n N_A_528_65#_c_816_n 0.0155838f $X=6.03 $Y=0.47 $X2=0 $Y2=0
cc_442 N_VGND_c_720_n N_A_528_65#_c_816_n 0.0140356f $X=6.48 $Y=0 $X2=0 $Y2=0
cc_443 N_VGND_c_721_n N_A_528_65#_c_816_n 0.00977851f $X=6.48 $Y=0 $X2=0 $Y2=0
