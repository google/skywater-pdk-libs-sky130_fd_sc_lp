* File: sky130_fd_sc_lp__dlrtp_lp2.pxi.spice
* Created: Fri Aug 28 10:27:29 2020
* 
x_PM_SKY130_FD_SC_LP__DLRTP_LP2%D N_D_c_156_n N_D_M1016_g N_D_M1022_g
+ N_D_c_157_n N_D_M1004_g N_D_c_158_n N_D_c_159_n D N_D_c_160_n N_D_c_161_n
+ PM_SKY130_FD_SC_LP__DLRTP_LP2%D
x_PM_SKY130_FD_SC_LP__DLRTP_LP2%GATE N_GATE_M1014_g N_GATE_M1017_g
+ N_GATE_c_200_n N_GATE_M1008_g GATE N_GATE_c_202_n
+ PM_SKY130_FD_SC_LP__DLRTP_LP2%GATE
x_PM_SKY130_FD_SC_LP__DLRTP_LP2%A_256_405# N_A_256_405#_M1008_d
+ N_A_256_405#_M1014_d N_A_256_405#_c_245_n N_A_256_405#_M1021_g
+ N_A_256_405#_c_264_n N_A_256_405#_M1001_g N_A_256_405#_c_246_n
+ N_A_256_405#_c_247_n N_A_256_405#_M1023_g N_A_256_405#_c_248_n
+ N_A_256_405#_M1019_g N_A_256_405#_c_249_n N_A_256_405#_M1018_g
+ N_A_256_405#_c_250_n N_A_256_405#_c_251_n N_A_256_405#_c_252_n
+ N_A_256_405#_c_253_n N_A_256_405#_c_254_n N_A_256_405#_c_255_n
+ N_A_256_405#_c_256_n N_A_256_405#_c_257_n N_A_256_405#_c_258_n
+ N_A_256_405#_c_259_n N_A_256_405#_c_270_n N_A_256_405#_c_260_n
+ N_A_256_405#_c_261_n N_A_256_405#_c_262_n N_A_256_405#_c_263_n
+ PM_SKY130_FD_SC_LP__DLRTP_LP2%A_256_405#
x_PM_SKY130_FD_SC_LP__DLRTP_LP2%A_27_122# N_A_27_122#_M1016_s
+ N_A_27_122#_M1022_s N_A_27_122#_M1010_g N_A_27_122#_c_401_n
+ N_A_27_122#_M1005_g N_A_27_122#_c_396_n N_A_27_122#_c_397_n
+ N_A_27_122#_c_404_n N_A_27_122#_c_405_n N_A_27_122#_c_406_n
+ N_A_27_122#_c_407_n N_A_27_122#_c_408_n N_A_27_122#_c_409_n
+ N_A_27_122#_c_398_n N_A_27_122#_c_399_n N_A_27_122#_c_411_n
+ N_A_27_122#_c_400_n N_A_27_122#_c_413_n
+ PM_SKY130_FD_SC_LP__DLRTP_LP2%A_27_122#
x_PM_SKY130_FD_SC_LP__DLRTP_LP2%A_413_47# N_A_413_47#_M1021_s
+ N_A_413_47#_M1001_s N_A_413_47#_M1011_g N_A_413_47#_c_509_n
+ N_A_413_47#_M1006_g N_A_413_47#_c_519_n N_A_413_47#_c_499_n
+ N_A_413_47#_c_511_n N_A_413_47#_c_500_n N_A_413_47#_c_512_n
+ N_A_413_47#_c_513_n N_A_413_47#_c_501_n N_A_413_47#_c_502_n
+ N_A_413_47#_c_551_n N_A_413_47#_c_503_n N_A_413_47#_c_504_n
+ N_A_413_47#_c_505_n N_A_413_47#_c_506_n N_A_413_47#_c_507_n
+ N_A_413_47#_c_508_n PM_SKY130_FD_SC_LP__DLRTP_LP2%A_413_47#
x_PM_SKY130_FD_SC_LP__DLRTP_LP2%A_898_21# N_A_898_21#_M1002_s
+ N_A_898_21#_M1020_d N_A_898_21#_M1015_g N_A_898_21#_c_641_n
+ N_A_898_21#_c_642_n N_A_898_21#_c_643_n N_A_898_21#_M1009_g
+ N_A_898_21#_M1012_g N_A_898_21#_M1000_g N_A_898_21#_M1013_g
+ N_A_898_21#_c_648_n N_A_898_21#_c_649_n N_A_898_21#_c_650_n
+ N_A_898_21#_c_659_n N_A_898_21#_c_651_n N_A_898_21#_c_652_n
+ N_A_898_21#_c_653_n N_A_898_21#_c_654_n N_A_898_21#_c_655_n
+ N_A_898_21#_c_656_n PM_SKY130_FD_SC_LP__DLRTP_LP2%A_898_21#
x_PM_SKY130_FD_SC_LP__DLRTP_LP2%A_736_47# N_A_736_47#_M1011_d
+ N_A_736_47#_M1019_d N_A_736_47#_M1020_g N_A_736_47#_c_765_n
+ N_A_736_47#_M1002_g N_A_736_47#_c_767_n N_A_736_47#_c_779_n
+ N_A_736_47#_c_787_n N_A_736_47#_c_768_n N_A_736_47#_c_769_n
+ N_A_736_47#_c_775_n N_A_736_47#_c_770_n N_A_736_47#_c_780_n
+ N_A_736_47#_c_771_n N_A_736_47#_c_772_n N_A_736_47#_c_773_n
+ PM_SKY130_FD_SC_LP__DLRTP_LP2%A_736_47#
x_PM_SKY130_FD_SC_LP__DLRTP_LP2%RESET_B N_RESET_B_c_874_n N_RESET_B_M1007_g
+ N_RESET_B_M1003_g N_RESET_B_c_880_n RESET_B N_RESET_B_c_876_n
+ N_RESET_B_c_877_n PM_SKY130_FD_SC_LP__DLRTP_LP2%RESET_B
x_PM_SKY130_FD_SC_LP__DLRTP_LP2%VPWR N_VPWR_M1022_d N_VPWR_M1001_d
+ N_VPWR_M1009_d N_VPWR_M1007_d N_VPWR_c_915_n N_VPWR_c_916_n N_VPWR_c_917_n
+ N_VPWR_c_918_n N_VPWR_c_919_n VPWR N_VPWR_c_920_n N_VPWR_c_921_n
+ N_VPWR_c_922_n N_VPWR_c_914_n N_VPWR_c_924_n N_VPWR_c_925_n N_VPWR_c_926_n
+ N_VPWR_c_927_n PM_SKY130_FD_SC_LP__DLRTP_LP2%VPWR
x_PM_SKY130_FD_SC_LP__DLRTP_LP2%Q N_Q_M1013_d N_Q_M1000_d Q Q Q Q Q Q Q Q Q
+ PM_SKY130_FD_SC_LP__DLRTP_LP2%Q
x_PM_SKY130_FD_SC_LP__DLRTP_LP2%VGND N_VGND_M1004_d N_VGND_M1023_d
+ N_VGND_M1015_d N_VGND_M1003_d N_VGND_c_1019_n N_VGND_c_1020_n N_VGND_c_1021_n
+ N_VGND_c_1022_n N_VGND_c_1023_n N_VGND_c_1024_n VGND N_VGND_c_1025_n
+ N_VGND_c_1026_n N_VGND_c_1027_n N_VGND_c_1028_n N_VGND_c_1029_n
+ N_VGND_c_1030_n N_VGND_c_1031_n N_VGND_c_1032_n
+ PM_SKY130_FD_SC_LP__DLRTP_LP2%VGND
cc_1 VNB N_D_c_156_n 0.0192939f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.105
cc_2 VNB N_D_c_157_n 0.0163095f $X=-0.19 $Y=-0.245 $X2=0.885 $Y2=1.105
cc_3 VNB N_D_c_158_n 0.0287344f $X=-0.19 $Y=-0.245 $X2=0.885 $Y2=1.18
cc_4 VNB N_D_c_159_n 0.00226072f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=1.865
cc_5 VNB N_D_c_160_n 0.0316575f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.36
cc_6 VNB N_D_c_161_n 0.00558412f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.36
cc_7 VNB N_GATE_M1014_g 0.00130545f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.82
cc_8 VNB N_GATE_M1017_g 0.0214923f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_GATE_c_200_n 0.0192859f $X=-0.19 $Y=-0.245 $X2=0.885 $Y2=0.82
cc_10 VNB N_GATE_M1008_g 0.0208342f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=1.18
cc_11 VNB N_GATE_c_202_n 0.0463701f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.36
cc_12 VNB N_A_256_405#_c_245_n 0.0171816f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_256_405#_c_246_n 0.0176764f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=1.69
cc_14 VNB N_A_256_405#_c_247_n 0.013607f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_15 VNB N_A_256_405#_c_248_n 0.0283076f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.36
cc_16 VNB N_A_256_405#_c_249_n 0.0264693f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_256_405#_c_250_n 0.00599687f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_256_405#_c_251_n 0.0031851f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_256_405#_c_252_n 0.0153497f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_256_405#_c_253_n 0.00970791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_256_405#_c_254_n 0.00257354f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_256_405#_c_255_n 0.0145478f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_256_405#_c_256_n 0.00270166f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_256_405#_c_257_n 0.0162903f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_256_405#_c_258_n 2.44051e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_256_405#_c_259_n 0.0054559f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_256_405#_c_260_n 0.0313653f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_256_405#_c_261_n 0.0203322f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_256_405#_c_262_n 0.00484309f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_256_405#_c_263_n 0.0381692f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_27_122#_M1010_g 0.0562436f $X=-0.19 $Y=-0.245 $X2=0.885 $Y2=0.82
cc_32 VNB N_A_27_122#_c_396_n 0.0232862f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_27_122#_c_397_n 0.0217692f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=1.865
cc_34 VNB N_A_27_122#_c_398_n 0.00254612f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_27_122#_c_399_n 0.020836f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_27_122#_c_400_n 0.0300931f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_413_47#_c_499_n 0.016162f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_38 VNB N_A_413_47#_c_500_n 0.012695f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.36
cc_39 VNB N_A_413_47#_c_501_n 0.00114335f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_413_47#_c_502_n 0.0307061f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_413_47#_c_503_n 0.00553223f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_413_47#_c_504_n 0.0345786f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_413_47#_c_505_n 0.00416923f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_413_47#_c_506_n 0.029529f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_413_47#_c_507_n 0.00320283f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_413_47#_c_508_n 0.0169775f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_898_21#_M1015_g 0.024054f $X=-0.19 $Y=-0.245 $X2=0.885 $Y2=0.82
cc_48 VNB N_A_898_21#_c_641_n 0.0229094f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.18
cc_49 VNB N_A_898_21#_c_642_n 0.00741149f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_898_21#_c_643_n 0.00742906f $X=-0.19 $Y=-0.245 $X2=0.885 $Y2=1.18
cc_51 VNB N_A_898_21#_M1009_g 0.00487747f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=1.69
cc_52 VNB N_A_898_21#_M1012_g 0.0185918f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=1.36
cc_53 VNB N_A_898_21#_M1000_g 0.0075825f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_898_21#_M1013_g 0.0218067f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_898_21#_c_648_n 0.0156293f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_898_21#_c_649_n 0.0152308f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_898_21#_c_650_n 0.0139186f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_898_21#_c_651_n 0.022626f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_898_21#_c_652_n 0.0116338f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_898_21#_c_653_n 0.0438897f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_A_898_21#_c_654_n 0.00441683f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_A_898_21#_c_655_n 0.00235538f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_A_898_21#_c_656_n 0.0730798f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_A_736_47#_c_765_n 0.0234549f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_A_736_47#_M1002_g 0.0210978f $X=-0.19 $Y=-0.245 $X2=0.885 $Y2=1.18
cc_66 VNB N_A_736_47#_c_767_n 0.0135238f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_67 VNB N_A_736_47#_c_768_n 0.00822778f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_A_736_47#_c_769_n 0.00422455f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_736_47#_c_770_n 0.00175204f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_A_736_47#_c_771_n 0.00688339f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_A_736_47#_c_772_n 0.00144345f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_A_736_47#_c_773_n 0.0279818f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_RESET_B_c_874_n 0.0166382f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.82
cc_74 VNB N_RESET_B_M1003_g 0.0366269f $X=-0.19 $Y=-0.245 $X2=0.885 $Y2=0.82
cc_75 VNB N_RESET_B_c_876_n 0.0156836f $X=-0.19 $Y=-0.245 $X2=0.885 $Y2=1.18
cc_76 VNB N_RESET_B_c_877_n 0.0049783f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_VPWR_c_914_n 0.322901f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB Q 0.0682573f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_VGND_c_1019_n 0.0388411f $X=-0.19 $Y=-0.245 $X2=0.885 $Y2=1.18
cc_80 VNB N_VGND_c_1020_n 4.89148e-19 $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_81 VNB N_VGND_c_1021_n 0.0131641f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.36
cc_82 VNB N_VGND_c_1022_n 0.00177638f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_VGND_c_1023_n 0.0471905f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_VGND_c_1024_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_VGND_c_1025_n 0.0301785f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_VGND_c_1026_n 0.043495f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_VGND_c_1027_n 0.0290222f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_VGND_c_1028_n 0.0279366f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_VGND_c_1029_n 0.439627f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_VGND_c_1030_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_VGND_c_1031_n 0.00436611f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_VGND_c_1032_n 0.00500486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_93 VPB N_D_M1022_g 0.0370908f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=2.595
cc_94 VPB N_D_c_159_n 0.013177f $X=-0.19 $Y=1.655 $X2=0.595 $Y2=1.865
cc_95 VPB N_D_c_160_n 0.00194062f $X=-0.19 $Y=1.655 $X2=0.605 $Y2=1.36
cc_96 VPB N_D_c_161_n 0.00234335f $X=-0.19 $Y=1.655 $X2=0.605 $Y2=1.36
cc_97 VPB N_GATE_M1014_g 0.0328197f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=0.82
cc_98 VPB N_A_256_405#_c_264_n 0.0358958f $X=-0.19 $Y=1.655 $X2=0.595 $Y2=1.255
cc_99 VPB N_A_256_405#_c_248_n 0.0152949f $X=-0.19 $Y=1.655 $X2=0.605 $Y2=1.36
cc_100 VPB N_A_256_405#_M1019_g 0.0284307f $X=-0.19 $Y=1.655 $X2=0.622 $Y2=1.36
cc_101 VPB N_A_256_405#_c_251_n 0.0120968f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_102 VPB N_A_256_405#_c_254_n 0.00653217f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_103 VPB N_A_256_405#_c_259_n 0.00326046f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_104 VPB N_A_256_405#_c_270_n 0.00592028f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_105 VPB N_A_256_405#_c_260_n 0.00301928f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_106 VPB N_A_256_405#_c_261_n 9.62611e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_107 VPB N_A_27_122#_c_401_n 0.0342814f $X=-0.19 $Y=1.655 $X2=0.595 $Y2=1.18
cc_108 VPB N_A_27_122#_c_396_n 0.0172471f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_109 VPB N_A_27_122#_c_397_n 0.0172806f $X=-0.19 $Y=1.655 $X2=0.595 $Y2=1.865
cc_110 VPB N_A_27_122#_c_404_n 0.00941382f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_111 VPB N_A_27_122#_c_405_n 0.00710076f $X=-0.19 $Y=1.655 $X2=0.622 $Y2=1.36
cc_112 VPB N_A_27_122#_c_406_n 0.0134814f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_113 VPB N_A_27_122#_c_407_n 0.0080362f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_114 VPB N_A_27_122#_c_408_n 0.0151521f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_115 VPB N_A_27_122#_c_409_n 0.0039324f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_116 VPB N_A_27_122#_c_398_n 0.00496059f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_117 VPB N_A_27_122#_c_411_n 0.0135379f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_118 VPB N_A_27_122#_c_400_n 0.0199876f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_119 VPB N_A_27_122#_c_413_n 0.0255395f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_120 VPB N_A_413_47#_c_509_n 0.0121238f $X=-0.19 $Y=1.655 $X2=0.885 $Y2=0.82
cc_121 VPB N_A_413_47#_M1006_g 0.0246112f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_122 VPB N_A_413_47#_c_511_n 7.33997e-19 $X=-0.19 $Y=1.655 $X2=0.605 $Y2=1.36
cc_123 VPB N_A_413_47#_c_512_n 0.00885883f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_124 VPB N_A_413_47#_c_513_n 0.00278214f $X=-0.19 $Y=1.655 $X2=0.622 $Y2=1.665
cc_125 VPB N_A_413_47#_c_501_n 0.00197679f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_126 VPB N_A_413_47#_c_506_n 0.00726743f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_127 VPB N_A_898_21#_M1009_g 0.0422317f $X=-0.19 $Y=1.655 $X2=0.595 $Y2=1.69
cc_128 VPB N_A_898_21#_M1000_g 0.0497053f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_129 VPB N_A_898_21#_c_659_n 0.00549821f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_130 VPB N_A_898_21#_c_654_n 0.00312646f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_131 VPB N_A_736_47#_M1020_g 0.0384096f $X=-0.19 $Y=1.655 $X2=0.885 $Y2=0.82
cc_132 VPB N_A_736_47#_c_775_n 0.00238489f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_133 VPB N_A_736_47#_c_770_n 0.00429752f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_134 VPB N_A_736_47#_c_772_n 6.27587e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_135 VPB N_A_736_47#_c_773_n 0.0174171f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_136 VPB N_RESET_B_c_874_n 0.0046318f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=0.82
cc_137 VPB N_RESET_B_M1007_g 0.0285571f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=2.595
cc_138 VPB N_RESET_B_c_880_n 0.013451f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=1.18
cc_139 VPB N_RESET_B_c_877_n 0.00386701f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_140 VPB N_VPWR_c_915_n 0.00360509f $X=-0.19 $Y=1.655 $X2=0.595 $Y2=1.69
cc_141 VPB N_VPWR_c_916_n 0.00284591f $X=-0.19 $Y=1.655 $X2=0.595 $Y2=1.36
cc_142 VPB N_VPWR_c_917_n 0.00936359f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_143 VPB N_VPWR_c_918_n 0.0216394f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_144 VPB N_VPWR_c_919_n 0.0105893f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_145 VPB N_VPWR_c_920_n 0.0450419f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_146 VPB N_VPWR_c_921_n 0.071533f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_147 VPB N_VPWR_c_922_n 0.0262716f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_148 VPB N_VPWR_c_914_n 0.0627065f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_149 VPB N_VPWR_c_924_n 0.0227192f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_150 VPB N_VPWR_c_925_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_151 VPB N_VPWR_c_926_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_152 VPB N_VPWR_c_927_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_153 VPB Q 0.0235588f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_154 VPB Q 0.019313f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=1.18
cc_155 VPB Q 0.0365561f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_156 N_D_M1022_g N_GATE_M1014_g 0.0401043f $X=0.545 $Y=2.595 $X2=0 $Y2=0
cc_157 N_D_c_159_n N_GATE_M1014_g 0.00186043f $X=0.595 $Y=1.865 $X2=0 $Y2=0
cc_158 N_D_c_161_n N_GATE_M1014_g 4.26954e-19 $X=0.605 $Y=1.36 $X2=0 $Y2=0
cc_159 N_D_c_157_n N_GATE_M1017_g 0.0130197f $X=0.885 $Y=1.105 $X2=0 $Y2=0
cc_160 N_D_c_160_n N_GATE_M1017_g 0.00390982f $X=0.605 $Y=1.36 $X2=0 $Y2=0
cc_161 N_D_c_161_n N_GATE_M1017_g 0.00412172f $X=0.605 $Y=1.36 $X2=0 $Y2=0
cc_162 N_D_c_160_n GATE 3.80404e-19 $X=0.605 $Y=1.36 $X2=0 $Y2=0
cc_163 N_D_c_161_n GATE 0.0250138f $X=0.605 $Y=1.36 $X2=0 $Y2=0
cc_164 N_D_c_160_n N_GATE_c_202_n 0.0215187f $X=0.605 $Y=1.36 $X2=0 $Y2=0
cc_165 N_D_c_161_n N_GATE_c_202_n 0.00205442f $X=0.605 $Y=1.36 $X2=0 $Y2=0
cc_166 N_D_c_161_n N_A_256_405#_c_254_n 0.00124999f $X=0.605 $Y=1.36 $X2=0 $Y2=0
cc_167 N_D_M1022_g N_A_256_405#_c_270_n 0.0010478f $X=0.545 $Y=2.595 $X2=0 $Y2=0
cc_168 N_D_c_161_n N_A_256_405#_c_261_n 0.00118273f $X=0.605 $Y=1.36 $X2=0 $Y2=0
cc_169 N_D_M1022_g N_A_27_122#_c_405_n 0.00392461f $X=0.545 $Y=2.595 $X2=0 $Y2=0
cc_170 N_D_M1022_g N_A_27_122#_c_406_n 0.0172714f $X=0.545 $Y=2.595 $X2=0 $Y2=0
cc_171 N_D_c_159_n N_A_27_122#_c_406_n 3.34149e-19 $X=0.595 $Y=1.865 $X2=0 $Y2=0
cc_172 N_D_c_161_n N_A_27_122#_c_406_n 0.00965431f $X=0.605 $Y=1.36 $X2=0 $Y2=0
cc_173 N_D_c_156_n N_A_27_122#_c_399_n 0.00940551f $X=0.495 $Y=1.105 $X2=0 $Y2=0
cc_174 N_D_c_157_n N_A_27_122#_c_399_n 0.00120234f $X=0.885 $Y=1.105 $X2=0 $Y2=0
cc_175 N_D_M1022_g N_A_27_122#_c_411_n 0.00547636f $X=0.545 $Y=2.595 $X2=0 $Y2=0
cc_176 N_D_c_156_n N_A_27_122#_c_400_n 0.0264126f $X=0.495 $Y=1.105 $X2=0 $Y2=0
cc_177 N_D_c_161_n N_A_27_122#_c_400_n 0.0485314f $X=0.605 $Y=1.36 $X2=0 $Y2=0
cc_178 N_D_M1022_g N_A_27_122#_c_413_n 0.0147858f $X=0.545 $Y=2.595 $X2=0 $Y2=0
cc_179 N_D_M1022_g N_VPWR_c_915_n 0.0119258f $X=0.545 $Y=2.595 $X2=0 $Y2=0
cc_180 N_D_M1022_g N_VPWR_c_914_n 0.00813366f $X=0.545 $Y=2.595 $X2=0 $Y2=0
cc_181 N_D_M1022_g N_VPWR_c_924_n 0.00644473f $X=0.545 $Y=2.595 $X2=0 $Y2=0
cc_182 N_D_c_156_n N_VGND_c_1019_n 0.00174824f $X=0.495 $Y=1.105 $X2=0 $Y2=0
cc_183 N_D_c_157_n N_VGND_c_1019_n 0.0135192f $X=0.885 $Y=1.105 $X2=0 $Y2=0
cc_184 N_D_c_156_n N_VGND_c_1025_n 0.00407419f $X=0.495 $Y=1.105 $X2=0 $Y2=0
cc_185 N_D_c_157_n N_VGND_c_1025_n 0.00351846f $X=0.885 $Y=1.105 $X2=0 $Y2=0
cc_186 N_D_c_156_n N_VGND_c_1029_n 0.00473597f $X=0.495 $Y=1.105 $X2=0 $Y2=0
cc_187 N_D_c_157_n N_VGND_c_1029_n 0.00397821f $X=0.885 $Y=1.105 $X2=0 $Y2=0
cc_188 N_GATE_M1008_g N_A_256_405#_c_250_n 0.00773833f $X=1.755 $Y=1.135 $X2=0
+ $Y2=0
cc_189 N_GATE_M1014_g N_A_256_405#_c_254_n 0.0060063f $X=1.155 $Y=2.525 $X2=0
+ $Y2=0
cc_190 N_GATE_c_200_n N_A_256_405#_c_254_n 8.81407e-19 $X=1.68 $Y=1.57 $X2=0
+ $Y2=0
cc_191 GATE N_A_256_405#_c_254_n 0.00265328f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_192 N_GATE_c_202_n N_A_256_405#_c_254_n 0.00124184f $X=1.47 $Y=1.66 $X2=0
+ $Y2=0
cc_193 N_GATE_M1017_g N_A_256_405#_c_255_n 0.00251958f $X=1.395 $Y=1.135 $X2=0
+ $Y2=0
cc_194 N_GATE_M1008_g N_A_256_405#_c_255_n 0.0134533f $X=1.755 $Y=1.135 $X2=0
+ $Y2=0
cc_195 N_GATE_M1014_g N_A_256_405#_c_270_n 0.00651758f $X=1.155 $Y=2.525 $X2=0
+ $Y2=0
cc_196 GATE N_A_256_405#_c_270_n 0.00212558f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_197 N_GATE_c_202_n N_A_256_405#_c_270_n 0.00768067f $X=1.47 $Y=1.66 $X2=0
+ $Y2=0
cc_198 N_GATE_M1008_g N_A_256_405#_c_260_n 0.00572505f $X=1.755 $Y=1.135 $X2=0
+ $Y2=0
cc_199 N_GATE_M1017_g N_A_256_405#_c_261_n 0.00130238f $X=1.395 $Y=1.135 $X2=0
+ $Y2=0
cc_200 N_GATE_c_200_n N_A_256_405#_c_261_n 0.0138845f $X=1.68 $Y=1.57 $X2=0
+ $Y2=0
cc_201 N_GATE_M1008_g N_A_256_405#_c_261_n 0.00739271f $X=1.755 $Y=1.135 $X2=0
+ $Y2=0
cc_202 GATE N_A_256_405#_c_261_n 0.0219118f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_203 N_GATE_c_202_n N_A_256_405#_c_261_n 0.00778243f $X=1.47 $Y=1.66 $X2=0
+ $Y2=0
cc_204 N_GATE_M1014_g N_A_27_122#_c_406_n 0.0231227f $X=1.155 $Y=2.525 $X2=0
+ $Y2=0
cc_205 GATE N_A_27_122#_c_406_n 0.0061624f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_206 N_GATE_M1014_g N_A_27_122#_c_407_n 0.00303902f $X=1.155 $Y=2.525 $X2=0
+ $Y2=0
cc_207 N_GATE_M1014_g N_A_27_122#_c_409_n 3.47799e-19 $X=1.155 $Y=2.525 $X2=0
+ $Y2=0
cc_208 N_GATE_M1014_g N_A_27_122#_c_411_n 0.0015159f $X=1.155 $Y=2.525 $X2=0
+ $Y2=0
cc_209 N_GATE_M1014_g N_A_27_122#_c_413_n 8.16956e-19 $X=1.155 $Y=2.525 $X2=0
+ $Y2=0
cc_210 N_GATE_M1008_g N_A_413_47#_c_502_n 0.00206431f $X=1.755 $Y=1.135 $X2=0
+ $Y2=0
cc_211 N_GATE_M1014_g N_VPWR_c_915_n 0.00471971f $X=1.155 $Y=2.525 $X2=0 $Y2=0
cc_212 N_GATE_M1014_g N_VPWR_c_920_n 0.00635322f $X=1.155 $Y=2.525 $X2=0 $Y2=0
cc_213 N_GATE_M1014_g N_VPWR_c_914_n 0.00925143f $X=1.155 $Y=2.525 $X2=0 $Y2=0
cc_214 N_GATE_M1017_g N_VGND_c_1019_n 0.00383559f $X=1.395 $Y=1.135 $X2=0 $Y2=0
cc_215 GATE N_VGND_c_1019_n 0.00961786f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_216 N_GATE_c_202_n N_VGND_c_1019_n 0.00590166f $X=1.47 $Y=1.66 $X2=0 $Y2=0
cc_217 N_GATE_M1017_g N_VGND_c_1029_n 0.00393927f $X=1.395 $Y=1.135 $X2=0 $Y2=0
cc_218 N_GATE_M1008_g N_VGND_c_1029_n 0.00393927f $X=1.755 $Y=1.135 $X2=0 $Y2=0
cc_219 N_A_256_405#_c_247_n N_A_27_122#_M1010_g 0.0200122f $X=2.785 $Y=0.73
+ $X2=0 $Y2=0
cc_220 N_A_256_405#_c_248_n N_A_27_122#_M1010_g 0.00145715f $X=4.065 $Y=1.85
+ $X2=0 $Y2=0
cc_221 N_A_256_405#_c_256_n N_A_27_122#_M1010_g 0.00256391f $X=2.455 $Y=1.455
+ $X2=0 $Y2=0
cc_222 N_A_256_405#_c_257_n N_A_27_122#_M1010_g 0.00960662f $X=3.22 $Y=1.16
+ $X2=0 $Y2=0
cc_223 N_A_256_405#_c_259_n N_A_27_122#_M1010_g 2.20407e-19 $X=4.005 $Y=1.5
+ $X2=0 $Y2=0
cc_224 N_A_256_405#_c_262_n N_A_27_122#_M1010_g 0.0155292f $X=3.305 $Y=1.16
+ $X2=0 $Y2=0
cc_225 N_A_256_405#_c_263_n N_A_27_122#_M1010_g 0.00876746f $X=2.375 $Y=1.455
+ $X2=0 $Y2=0
cc_226 N_A_256_405#_M1019_g N_A_27_122#_c_401_n 0.0741153f $X=4.065 $Y=2.595
+ $X2=0 $Y2=0
cc_227 N_A_256_405#_c_259_n N_A_27_122#_c_401_n 0.0029558f $X=4.005 $Y=1.5 $X2=0
+ $Y2=0
cc_228 N_A_256_405#_c_246_n N_A_27_122#_c_396_n 0.00183352f $X=2.71 $Y=0.805
+ $X2=0 $Y2=0
cc_229 N_A_256_405#_c_257_n N_A_27_122#_c_396_n 0.00540299f $X=3.22 $Y=1.16
+ $X2=0 $Y2=0
cc_230 N_A_256_405#_c_260_n N_A_27_122#_c_396_n 0.0200273f $X=2.375 $Y=1.62
+ $X2=0 $Y2=0
cc_231 N_A_256_405#_c_261_n N_A_27_122#_c_396_n 0.00120538f $X=2.455 $Y=1.62
+ $X2=0 $Y2=0
cc_232 N_A_256_405#_c_263_n N_A_27_122#_c_396_n 0.00156916f $X=2.375 $Y=1.455
+ $X2=0 $Y2=0
cc_233 N_A_256_405#_c_248_n N_A_27_122#_c_397_n 0.0184282f $X=4.065 $Y=1.85
+ $X2=0 $Y2=0
cc_234 N_A_256_405#_c_259_n N_A_27_122#_c_397_n 0.016945f $X=4.005 $Y=1.5 $X2=0
+ $Y2=0
cc_235 N_A_256_405#_c_262_n N_A_27_122#_c_397_n 0.0130715f $X=3.305 $Y=1.16
+ $X2=0 $Y2=0
cc_236 N_A_256_405#_M1019_g N_A_27_122#_c_404_n 0.00515706f $X=4.065 $Y=2.595
+ $X2=0 $Y2=0
cc_237 N_A_256_405#_M1014_d N_A_27_122#_c_406_n 0.00770714f $X=1.28 $Y=2.025
+ $X2=0 $Y2=0
cc_238 N_A_256_405#_c_270_n N_A_27_122#_c_406_n 0.0231542f $X=1.55 $Y=2.13 $X2=0
+ $Y2=0
cc_239 N_A_256_405#_c_261_n N_A_27_122#_c_406_n 0.00558517f $X=2.455 $Y=1.62
+ $X2=0 $Y2=0
cc_240 N_A_256_405#_c_264_n N_A_27_122#_c_407_n 0.00464127f $X=2.515 $Y=2.09
+ $X2=0 $Y2=0
cc_241 N_A_256_405#_c_270_n N_A_27_122#_c_407_n 0.00916854f $X=1.55 $Y=2.13
+ $X2=0 $Y2=0
cc_242 N_A_256_405#_c_264_n N_A_27_122#_c_408_n 0.0205122f $X=2.515 $Y=2.09
+ $X2=0 $Y2=0
cc_243 N_A_256_405#_c_260_n N_A_27_122#_c_408_n 0.00416569f $X=2.375 $Y=1.62
+ $X2=0 $Y2=0
cc_244 N_A_256_405#_c_261_n N_A_27_122#_c_408_n 0.0402886f $X=2.455 $Y=1.62
+ $X2=0 $Y2=0
cc_245 N_A_256_405#_c_254_n N_A_27_122#_c_409_n 0.00324419f $X=1.55 $Y=2.005
+ $X2=0 $Y2=0
cc_246 N_A_256_405#_c_270_n N_A_27_122#_c_409_n 0.0111178f $X=1.55 $Y=2.13 $X2=0
+ $Y2=0
cc_247 N_A_256_405#_c_261_n N_A_27_122#_c_409_n 0.0143719f $X=2.455 $Y=1.62
+ $X2=0 $Y2=0
cc_248 N_A_256_405#_c_256_n N_A_27_122#_c_398_n 0.0019055f $X=2.455 $Y=1.455
+ $X2=0 $Y2=0
cc_249 N_A_256_405#_c_257_n N_A_27_122#_c_398_n 0.0221127f $X=3.22 $Y=1.16 $X2=0
+ $Y2=0
cc_250 N_A_256_405#_c_260_n N_A_27_122#_c_398_n 0.00686394f $X=2.375 $Y=1.62
+ $X2=0 $Y2=0
cc_251 N_A_256_405#_c_261_n N_A_27_122#_c_398_n 0.0220051f $X=2.455 $Y=1.62
+ $X2=0 $Y2=0
cc_252 N_A_256_405#_c_262_n N_A_27_122#_c_398_n 0.0162026f $X=3.305 $Y=1.16
+ $X2=0 $Y2=0
cc_253 N_A_256_405#_M1019_g N_A_413_47#_c_509_n 0.00554309f $X=4.065 $Y=2.595
+ $X2=0 $Y2=0
cc_254 N_A_256_405#_M1019_g N_A_413_47#_M1006_g 0.0245482f $X=4.065 $Y=2.595
+ $X2=0 $Y2=0
cc_255 N_A_256_405#_c_264_n N_A_413_47#_c_519_n 0.0159733f $X=2.515 $Y=2.09
+ $X2=0 $Y2=0
cc_256 N_A_256_405#_M1019_g N_A_413_47#_c_519_n 0.00613887f $X=4.065 $Y=2.595
+ $X2=0 $Y2=0
cc_257 N_A_256_405#_c_259_n N_A_413_47#_c_519_n 0.0096365f $X=4.005 $Y=1.5 $X2=0
+ $Y2=0
cc_258 N_A_256_405#_c_262_n N_A_413_47#_c_519_n 0.00448562f $X=3.305 $Y=1.16
+ $X2=0 $Y2=0
cc_259 N_A_256_405#_c_245_n N_A_413_47#_c_499_n 3.54547e-19 $X=2.425 $Y=0.73
+ $X2=0 $Y2=0
cc_260 N_A_256_405#_c_246_n N_A_413_47#_c_499_n 0.0114266f $X=2.71 $Y=0.805
+ $X2=0 $Y2=0
cc_261 N_A_256_405#_c_247_n N_A_413_47#_c_499_n 0.00354303f $X=2.785 $Y=0.73
+ $X2=0 $Y2=0
cc_262 N_A_256_405#_c_257_n N_A_413_47#_c_499_n 0.0485349f $X=3.22 $Y=1.16 $X2=0
+ $Y2=0
cc_263 N_A_256_405#_c_258_n N_A_413_47#_c_499_n 0.00410463f $X=2.54 $Y=1.16
+ $X2=0 $Y2=0
cc_264 N_A_256_405#_c_259_n N_A_413_47#_c_499_n 0.00724109f $X=4.005 $Y=1.5
+ $X2=0 $Y2=0
cc_265 N_A_256_405#_c_262_n N_A_413_47#_c_499_n 0.0128956f $X=3.305 $Y=1.16
+ $X2=0 $Y2=0
cc_266 N_A_256_405#_c_263_n N_A_413_47#_c_499_n 4.55432e-19 $X=2.375 $Y=1.455
+ $X2=0 $Y2=0
cc_267 N_A_256_405#_M1019_g N_A_413_47#_c_511_n 0.00748099f $X=4.065 $Y=2.595
+ $X2=0 $Y2=0
cc_268 N_A_256_405#_c_248_n N_A_413_47#_c_500_n 0.00504024f $X=4.065 $Y=1.85
+ $X2=0 $Y2=0
cc_269 N_A_256_405#_c_249_n N_A_413_47#_c_500_n 0.0128363f $X=4.145 $Y=1.335
+ $X2=0 $Y2=0
cc_270 N_A_256_405#_c_253_n N_A_413_47#_c_500_n 0.00100378f $X=4.16 $Y=0.88
+ $X2=0 $Y2=0
cc_271 N_A_256_405#_c_259_n N_A_413_47#_c_500_n 0.0176156f $X=4.005 $Y=1.5 $X2=0
+ $Y2=0
cc_272 N_A_256_405#_c_248_n N_A_413_47#_c_512_n 0.00409261f $X=4.065 $Y=1.85
+ $X2=0 $Y2=0
cc_273 N_A_256_405#_M1019_g N_A_413_47#_c_512_n 0.0131907f $X=4.065 $Y=2.595
+ $X2=0 $Y2=0
cc_274 N_A_256_405#_c_259_n N_A_413_47#_c_512_n 0.0125871f $X=4.005 $Y=1.5 $X2=0
+ $Y2=0
cc_275 N_A_256_405#_c_248_n N_A_413_47#_c_513_n 0.00302044f $X=4.065 $Y=1.85
+ $X2=0 $Y2=0
cc_276 N_A_256_405#_M1019_g N_A_413_47#_c_513_n 0.00177177f $X=4.065 $Y=2.595
+ $X2=0 $Y2=0
cc_277 N_A_256_405#_c_259_n N_A_413_47#_c_513_n 0.0135646f $X=4.005 $Y=1.5 $X2=0
+ $Y2=0
cc_278 N_A_256_405#_c_248_n N_A_413_47#_c_501_n 0.00508972f $X=4.065 $Y=1.85
+ $X2=0 $Y2=0
cc_279 N_A_256_405#_c_245_n N_A_413_47#_c_502_n 0.0132432f $X=2.425 $Y=0.73
+ $X2=0 $Y2=0
cc_280 N_A_256_405#_c_247_n N_A_413_47#_c_502_n 0.00206982f $X=2.785 $Y=0.73
+ $X2=0 $Y2=0
cc_281 N_A_256_405#_c_250_n N_A_413_47#_c_502_n 0.00358482f $X=2.425 $Y=0.805
+ $X2=0 $Y2=0
cc_282 N_A_256_405#_c_255_n N_A_413_47#_c_502_n 0.00638371f $X=1.97 $Y=1.09
+ $X2=0 $Y2=0
cc_283 N_A_256_405#_c_258_n N_A_413_47#_c_502_n 0.00884952f $X=2.54 $Y=1.16
+ $X2=0 $Y2=0
cc_284 N_A_256_405#_c_260_n N_A_413_47#_c_502_n 6.21605e-19 $X=2.375 $Y=1.62
+ $X2=0 $Y2=0
cc_285 N_A_256_405#_c_261_n N_A_413_47#_c_502_n 0.00180461f $X=2.455 $Y=1.62
+ $X2=0 $Y2=0
cc_286 N_A_256_405#_c_263_n N_A_413_47#_c_502_n 0.00256282f $X=2.375 $Y=1.455
+ $X2=0 $Y2=0
cc_287 N_A_256_405#_c_264_n N_A_413_47#_c_551_n 0.0161819f $X=2.515 $Y=2.09
+ $X2=0 $Y2=0
cc_288 N_A_256_405#_c_253_n N_A_413_47#_c_503_n 0.00189314f $X=4.16 $Y=0.88
+ $X2=0 $Y2=0
cc_289 N_A_256_405#_c_259_n N_A_413_47#_c_503_n 0.0177517f $X=4.005 $Y=1.5 $X2=0
+ $Y2=0
cc_290 N_A_256_405#_c_262_n N_A_413_47#_c_503_n 0.00142563f $X=3.305 $Y=1.16
+ $X2=0 $Y2=0
cc_291 N_A_256_405#_c_248_n N_A_413_47#_c_504_n 0.00107992f $X=4.065 $Y=1.85
+ $X2=0 $Y2=0
cc_292 N_A_256_405#_c_253_n N_A_413_47#_c_504_n 0.0213211f $X=4.16 $Y=0.88 $X2=0
+ $Y2=0
cc_293 N_A_256_405#_c_259_n N_A_413_47#_c_504_n 0.00223255f $X=4.005 $Y=1.5
+ $X2=0 $Y2=0
cc_294 N_A_256_405#_c_248_n N_A_413_47#_c_505_n 0.00438844f $X=4.065 $Y=1.85
+ $X2=0 $Y2=0
cc_295 N_A_256_405#_c_259_n N_A_413_47#_c_505_n 0.0267533f $X=4.005 $Y=1.5 $X2=0
+ $Y2=0
cc_296 N_A_256_405#_c_248_n N_A_413_47#_c_506_n 0.0172882f $X=4.065 $Y=1.85
+ $X2=0 $Y2=0
cc_297 N_A_256_405#_c_249_n N_A_413_47#_c_506_n 0.0135117f $X=4.145 $Y=1.335
+ $X2=0 $Y2=0
cc_298 N_A_256_405#_c_259_n N_A_413_47#_c_506_n 3.43945e-19 $X=4.005 $Y=1.5
+ $X2=0 $Y2=0
cc_299 N_A_256_405#_c_249_n N_A_413_47#_c_507_n 0.00438844f $X=4.145 $Y=1.335
+ $X2=0 $Y2=0
cc_300 N_A_256_405#_c_252_n N_A_413_47#_c_508_n 0.0134789f $X=4.16 $Y=0.73 $X2=0
+ $Y2=0
cc_301 N_A_256_405#_c_253_n N_A_413_47#_c_508_n 8.9655e-19 $X=4.16 $Y=0.88 $X2=0
+ $Y2=0
cc_302 N_A_256_405#_c_252_n N_A_898_21#_M1015_g 0.0214586f $X=4.16 $Y=0.73 $X2=0
+ $Y2=0
cc_303 N_A_256_405#_c_249_n N_A_898_21#_c_642_n 0.00608154f $X=4.145 $Y=1.335
+ $X2=0 $Y2=0
cc_304 N_A_256_405#_c_253_n N_A_898_21#_c_642_n 0.0214586f $X=4.16 $Y=0.88 $X2=0
+ $Y2=0
cc_305 N_A_256_405#_c_252_n N_A_736_47#_c_779_n 0.0106686f $X=4.16 $Y=0.73 $X2=0
+ $Y2=0
cc_306 N_A_256_405#_M1019_g N_A_736_47#_c_780_n 0.0183851f $X=4.065 $Y=2.595
+ $X2=0 $Y2=0
cc_307 N_A_256_405#_c_249_n N_A_736_47#_c_771_n 3.12531e-19 $X=4.145 $Y=1.335
+ $X2=0 $Y2=0
cc_308 N_A_256_405#_c_264_n N_VPWR_c_916_n 0.0155327f $X=2.515 $Y=2.09 $X2=0
+ $Y2=0
cc_309 N_A_256_405#_c_264_n N_VPWR_c_920_n 0.00840199f $X=2.515 $Y=2.09 $X2=0
+ $Y2=0
cc_310 N_A_256_405#_M1019_g N_VPWR_c_921_n 0.00939541f $X=4.065 $Y=2.595 $X2=0
+ $Y2=0
cc_311 N_A_256_405#_c_264_n N_VPWR_c_914_n 0.00890821f $X=2.515 $Y=2.09 $X2=0
+ $Y2=0
cc_312 N_A_256_405#_M1019_g N_VPWR_c_914_n 0.0148209f $X=4.065 $Y=2.595 $X2=0
+ $Y2=0
cc_313 N_A_256_405#_c_255_n N_VGND_c_1019_n 0.00194949f $X=1.97 $Y=1.09 $X2=0
+ $Y2=0
cc_314 N_A_256_405#_c_245_n N_VGND_c_1020_n 0.00199396f $X=2.425 $Y=0.73 $X2=0
+ $Y2=0
cc_315 N_A_256_405#_c_247_n N_VGND_c_1020_n 0.00952074f $X=2.785 $Y=0.73 $X2=0
+ $Y2=0
cc_316 N_A_256_405#_c_252_n N_VGND_c_1023_n 0.00366111f $X=4.16 $Y=0.73 $X2=0
+ $Y2=0
cc_317 N_A_256_405#_c_245_n N_VGND_c_1026_n 0.00367566f $X=2.425 $Y=0.73 $X2=0
+ $Y2=0
cc_318 N_A_256_405#_c_247_n N_VGND_c_1026_n 0.00364083f $X=2.785 $Y=0.73 $X2=0
+ $Y2=0
cc_319 N_A_256_405#_c_245_n N_VGND_c_1029_n 0.00669453f $X=2.425 $Y=0.73 $X2=0
+ $Y2=0
cc_320 N_A_256_405#_c_247_n N_VGND_c_1029_n 0.00416707f $X=2.785 $Y=0.73 $X2=0
+ $Y2=0
cc_321 N_A_256_405#_c_252_n N_VGND_c_1029_n 0.00560843f $X=4.16 $Y=0.73 $X2=0
+ $Y2=0
cc_322 N_A_27_122#_c_408_n N_A_413_47#_M1001_s 0.00434523f $X=2.75 $Y=2.05 $X2=0
+ $Y2=0
cc_323 N_A_27_122#_c_401_n N_A_413_47#_c_519_n 0.0225509f $X=3.575 $Y=2.03 $X2=0
+ $Y2=0
cc_324 N_A_27_122#_c_396_n N_A_413_47#_c_519_n 0.00954944f $X=3.14 $Y=1.59 $X2=0
+ $Y2=0
cc_325 N_A_27_122#_c_408_n N_A_413_47#_c_519_n 0.0408756f $X=2.75 $Y=2.05 $X2=0
+ $Y2=0
cc_326 N_A_27_122#_M1010_g N_A_413_47#_c_499_n 0.01171f $X=3.215 $Y=0.445 $X2=0
+ $Y2=0
cc_327 N_A_27_122#_c_397_n N_A_413_47#_c_499_n 0.00104421f $X=3.525 $Y=1.59
+ $X2=0 $Y2=0
cc_328 N_A_27_122#_c_401_n N_A_413_47#_c_511_n 0.00657478f $X=3.575 $Y=2.03
+ $X2=0 $Y2=0
cc_329 N_A_27_122#_c_401_n N_A_413_47#_c_513_n 0.00322665f $X=3.575 $Y=2.03
+ $X2=0 $Y2=0
cc_330 N_A_27_122#_c_404_n N_A_413_47#_c_513_n 0.00159794f $X=3.575 $Y=1.905
+ $X2=0 $Y2=0
cc_331 N_A_27_122#_c_406_n N_A_413_47#_c_551_n 0.0141898f $X=1.815 $Y=2.52 $X2=0
+ $Y2=0
cc_332 N_A_27_122#_c_407_n N_A_413_47#_c_551_n 0.00948056f $X=1.9 $Y=2.435 $X2=0
+ $Y2=0
cc_333 N_A_27_122#_c_408_n N_A_413_47#_c_551_n 0.0148745f $X=2.75 $Y=2.05 $X2=0
+ $Y2=0
cc_334 N_A_27_122#_M1010_g N_A_413_47#_c_503_n 0.00118825f $X=3.215 $Y=0.445
+ $X2=0 $Y2=0
cc_335 N_A_27_122#_c_397_n N_A_413_47#_c_504_n 0.00259646f $X=3.525 $Y=1.59
+ $X2=0 $Y2=0
cc_336 N_A_27_122#_M1010_g N_A_413_47#_c_508_n 0.0544409f $X=3.215 $Y=0.445
+ $X2=0 $Y2=0
cc_337 N_A_27_122#_c_401_n N_A_736_47#_c_780_n 0.00257902f $X=3.575 $Y=2.03
+ $X2=0 $Y2=0
cc_338 N_A_27_122#_c_406_n N_VPWR_M1022_d 0.0104293f $X=1.815 $Y=2.52 $X2=-0.19
+ $Y2=-0.245
cc_339 N_A_27_122#_c_408_n N_VPWR_M1001_d 0.00500324f $X=2.75 $Y=2.05 $X2=0
+ $Y2=0
cc_340 N_A_27_122#_c_406_n N_VPWR_c_915_n 0.0199416f $X=1.815 $Y=2.52 $X2=0
+ $Y2=0
cc_341 N_A_27_122#_c_413_n N_VPWR_c_915_n 0.0185531f $X=0.267 $Y=2.52 $X2=0
+ $Y2=0
cc_342 N_A_27_122#_c_401_n N_VPWR_c_916_n 0.0138456f $X=3.575 $Y=2.03 $X2=0
+ $Y2=0
cc_343 N_A_27_122#_c_406_n N_VPWR_c_920_n 0.0141615f $X=1.815 $Y=2.52 $X2=0
+ $Y2=0
cc_344 N_A_27_122#_c_401_n N_VPWR_c_921_n 0.00975641f $X=3.575 $Y=2.03 $X2=0
+ $Y2=0
cc_345 N_A_27_122#_M1022_s N_VPWR_c_914_n 0.0023218f $X=0.135 $Y=2.095 $X2=0
+ $Y2=0
cc_346 N_A_27_122#_c_401_n N_VPWR_c_914_n 0.0111162f $X=3.575 $Y=2.03 $X2=0
+ $Y2=0
cc_347 N_A_27_122#_c_406_n N_VPWR_c_914_n 0.0316137f $X=1.815 $Y=2.52 $X2=0
+ $Y2=0
cc_348 N_A_27_122#_c_413_n N_VPWR_c_914_n 0.0134754f $X=0.267 $Y=2.52 $X2=0
+ $Y2=0
cc_349 N_A_27_122#_c_406_n N_VPWR_c_924_n 0.00265901f $X=1.815 $Y=2.52 $X2=0
+ $Y2=0
cc_350 N_A_27_122#_c_413_n N_VPWR_c_924_n 0.0214436f $X=0.267 $Y=2.52 $X2=0
+ $Y2=0
cc_351 N_A_27_122#_c_399_n N_VGND_c_1019_n 0.01354f $X=0.28 $Y=0.8 $X2=0 $Y2=0
cc_352 N_A_27_122#_M1010_g N_VGND_c_1020_n 0.0108487f $X=3.215 $Y=0.445 $X2=0
+ $Y2=0
cc_353 N_A_27_122#_M1010_g N_VGND_c_1023_n 0.00364083f $X=3.215 $Y=0.445 $X2=0
+ $Y2=0
cc_354 N_A_27_122#_c_399_n N_VGND_c_1025_n 0.007677f $X=0.28 $Y=0.8 $X2=0 $Y2=0
cc_355 N_A_27_122#_M1010_g N_VGND_c_1029_n 0.00429664f $X=3.215 $Y=0.445 $X2=0
+ $Y2=0
cc_356 N_A_27_122#_c_399_n N_VGND_c_1029_n 0.010926f $X=0.28 $Y=0.8 $X2=0 $Y2=0
cc_357 N_A_413_47#_c_500_n N_A_898_21#_c_642_n 0.00333086f $X=4.35 $Y=1.01 $X2=0
+ $Y2=0
cc_358 N_A_413_47#_c_505_n N_A_898_21#_c_642_n 0.00126928f $X=4.595 $Y=1.43
+ $X2=0 $Y2=0
cc_359 N_A_413_47#_c_506_n N_A_898_21#_c_642_n 0.0134161f $X=4.595 $Y=1.43 $X2=0
+ $Y2=0
cc_360 N_A_413_47#_c_509_n N_A_898_21#_c_643_n 0.0209814f $X=4.595 $Y=1.935
+ $X2=0 $Y2=0
cc_361 N_A_413_47#_c_501_n N_A_898_21#_c_643_n 3.42921e-19 $X=4.555 $Y=1.845
+ $X2=0 $Y2=0
cc_362 N_A_413_47#_M1006_g N_A_898_21#_M1009_g 0.0681554f $X=4.595 $Y=2.595
+ $X2=0 $Y2=0
cc_363 N_A_413_47#_c_512_n N_A_898_21#_M1009_g 4.03281e-19 $X=4.35 $Y=1.93 $X2=0
+ $Y2=0
cc_364 N_A_413_47#_c_500_n N_A_898_21#_c_648_n 5.37086e-19 $X=4.35 $Y=1.01 $X2=0
+ $Y2=0
cc_365 N_A_413_47#_c_507_n N_A_898_21#_c_648_n 9.19002e-19 $X=4.555 $Y=1.265
+ $X2=0 $Y2=0
cc_366 N_A_413_47#_c_505_n N_A_898_21#_c_649_n 3.42921e-19 $X=4.595 $Y=1.43
+ $X2=0 $Y2=0
cc_367 N_A_413_47#_c_506_n N_A_898_21#_c_649_n 0.0209814f $X=4.595 $Y=1.43 $X2=0
+ $Y2=0
cc_368 N_A_413_47#_c_500_n N_A_736_47#_c_779_n 0.0243339f $X=4.35 $Y=1.01 $X2=0
+ $Y2=0
cc_369 N_A_413_47#_c_503_n N_A_736_47#_c_779_n 0.00475921f $X=3.715 $Y=0.81
+ $X2=0 $Y2=0
cc_370 N_A_413_47#_c_504_n N_A_736_47#_c_779_n 4.12436e-19 $X=3.695 $Y=0.93
+ $X2=0 $Y2=0
cc_371 N_A_413_47#_c_508_n N_A_736_47#_c_779_n 0.00391466f $X=3.695 $Y=0.765
+ $X2=0 $Y2=0
cc_372 N_A_413_47#_M1006_g N_A_736_47#_c_787_n 0.018389f $X=4.595 $Y=2.595 $X2=0
+ $Y2=0
cc_373 N_A_413_47#_c_512_n N_A_736_47#_c_787_n 0.0181265f $X=4.35 $Y=1.93 $X2=0
+ $Y2=0
cc_374 N_A_413_47#_c_500_n N_A_736_47#_c_769_n 0.00314842f $X=4.35 $Y=1.01 $X2=0
+ $Y2=0
cc_375 N_A_413_47#_c_505_n N_A_736_47#_c_769_n 0.0116756f $X=4.595 $Y=1.43 $X2=0
+ $Y2=0
cc_376 N_A_413_47#_c_506_n N_A_736_47#_c_769_n 8.4353e-19 $X=4.595 $Y=1.43 $X2=0
+ $Y2=0
cc_377 N_A_413_47#_c_507_n N_A_736_47#_c_769_n 0.00681083f $X=4.555 $Y=1.265
+ $X2=0 $Y2=0
cc_378 N_A_413_47#_c_509_n N_A_736_47#_c_775_n 2.6691e-19 $X=4.595 $Y=1.935
+ $X2=0 $Y2=0
cc_379 N_A_413_47#_M1006_g N_A_736_47#_c_775_n 0.00207511f $X=4.595 $Y=2.595
+ $X2=0 $Y2=0
cc_380 N_A_413_47#_c_512_n N_A_736_47#_c_775_n 0.0133724f $X=4.35 $Y=1.93 $X2=0
+ $Y2=0
cc_381 N_A_413_47#_c_501_n N_A_736_47#_c_775_n 0.00647763f $X=4.555 $Y=1.845
+ $X2=0 $Y2=0
cc_382 N_A_413_47#_c_506_n N_A_736_47#_c_775_n 4.70475e-19 $X=4.595 $Y=1.43
+ $X2=0 $Y2=0
cc_383 N_A_413_47#_M1006_g N_A_736_47#_c_780_n 0.0165729f $X=4.595 $Y=2.595
+ $X2=0 $Y2=0
cc_384 N_A_413_47#_c_519_n N_A_736_47#_c_780_n 0.013152f $X=3.815 $Y=2.4 $X2=0
+ $Y2=0
cc_385 N_A_413_47#_c_511_n N_A_736_47#_c_780_n 0.00869659f $X=3.9 $Y=2.315 $X2=0
+ $Y2=0
cc_386 N_A_413_47#_c_512_n N_A_736_47#_c_780_n 0.022033f $X=4.35 $Y=1.93 $X2=0
+ $Y2=0
cc_387 N_A_413_47#_c_500_n N_A_736_47#_c_771_n 0.00785373f $X=4.35 $Y=1.01 $X2=0
+ $Y2=0
cc_388 N_A_413_47#_c_505_n N_A_736_47#_c_771_n 0.00363449f $X=4.595 $Y=1.43
+ $X2=0 $Y2=0
cc_389 N_A_413_47#_c_505_n N_A_736_47#_c_772_n 0.0270215f $X=4.595 $Y=1.43 $X2=0
+ $Y2=0
cc_390 N_A_413_47#_c_506_n N_A_736_47#_c_772_n 0.0020377f $X=4.595 $Y=1.43 $X2=0
+ $Y2=0
cc_391 N_A_413_47#_c_519_n N_VPWR_M1001_d 0.0251919f $X=3.815 $Y=2.4 $X2=0 $Y2=0
cc_392 N_A_413_47#_c_519_n N_VPWR_c_916_n 0.0204264f $X=3.815 $Y=2.4 $X2=0 $Y2=0
cc_393 N_A_413_47#_c_551_n N_VPWR_c_916_n 0.0258074f $X=2.25 $Y=2.48 $X2=0 $Y2=0
cc_394 N_A_413_47#_c_551_n N_VPWR_c_920_n 0.014447f $X=2.25 $Y=2.48 $X2=0 $Y2=0
cc_395 N_A_413_47#_M1006_g N_VPWR_c_921_n 0.00939541f $X=4.595 $Y=2.595 $X2=0
+ $Y2=0
cc_396 N_A_413_47#_M1001_s N_VPWR_c_914_n 0.00444327f $X=2.105 $Y=2.095 $X2=0
+ $Y2=0
cc_397 N_A_413_47#_M1006_g N_VPWR_c_914_n 0.0161801f $X=4.595 $Y=2.595 $X2=0
+ $Y2=0
cc_398 N_A_413_47#_c_519_n N_VPWR_c_914_n 0.0409575f $X=3.815 $Y=2.4 $X2=0 $Y2=0
cc_399 N_A_413_47#_c_551_n N_VPWR_c_914_n 0.00941258f $X=2.25 $Y=2.48 $X2=0
+ $Y2=0
cc_400 N_A_413_47#_c_519_n A_740_419# 0.00392117f $X=3.815 $Y=2.4 $X2=-0.19
+ $Y2=-0.245
cc_401 N_A_413_47#_c_511_n A_740_419# 0.0024603f $X=3.9 $Y=2.315 $X2=-0.19
+ $Y2=-0.245
cc_402 N_A_413_47#_c_499_n N_VGND_c_1020_n 0.0195998f $X=3.57 $Y=0.81 $X2=0
+ $Y2=0
cc_403 N_A_413_47#_c_502_n N_VGND_c_1020_n 0.0120699f $X=2.21 $Y=0.47 $X2=0
+ $Y2=0
cc_404 N_A_413_47#_c_508_n N_VGND_c_1020_n 0.00214335f $X=3.695 $Y=0.765 $X2=0
+ $Y2=0
cc_405 N_A_413_47#_c_499_n N_VGND_c_1023_n 0.00584617f $X=3.57 $Y=0.81 $X2=0
+ $Y2=0
cc_406 N_A_413_47#_c_503_n N_VGND_c_1023_n 0.00339779f $X=3.715 $Y=0.81 $X2=0
+ $Y2=0
cc_407 N_A_413_47#_c_504_n N_VGND_c_1023_n 4.15653e-19 $X=3.695 $Y=0.93 $X2=0
+ $Y2=0
cc_408 N_A_413_47#_c_508_n N_VGND_c_1023_n 0.00438737f $X=3.695 $Y=0.765 $X2=0
+ $Y2=0
cc_409 N_A_413_47#_c_499_n N_VGND_c_1026_n 0.00505036f $X=3.57 $Y=0.81 $X2=0
+ $Y2=0
cc_410 N_A_413_47#_c_502_n N_VGND_c_1026_n 0.0263217f $X=2.21 $Y=0.47 $X2=0
+ $Y2=0
cc_411 N_A_413_47#_M1021_s N_VGND_c_1029_n 0.00232985f $X=2.065 $Y=0.235 $X2=0
+ $Y2=0
cc_412 N_A_413_47#_c_499_n N_VGND_c_1029_n 0.0199216f $X=3.57 $Y=0.81 $X2=0
+ $Y2=0
cc_413 N_A_413_47#_c_502_n N_VGND_c_1029_n 0.0162517f $X=2.21 $Y=0.47 $X2=0
+ $Y2=0
cc_414 N_A_413_47#_c_503_n N_VGND_c_1029_n 0.00575652f $X=3.715 $Y=0.81 $X2=0
+ $Y2=0
cc_415 N_A_413_47#_c_508_n N_VGND_c_1029_n 0.00649907f $X=3.695 $Y=0.765 $X2=0
+ $Y2=0
cc_416 N_A_898_21#_M1009_g N_A_736_47#_M1020_g 0.0303836f $X=5.095 $Y=2.595
+ $X2=0 $Y2=0
cc_417 N_A_898_21#_c_659_n N_A_736_47#_M1020_g 0.0188022f $X=6.065 $Y=2.24 $X2=0
+ $Y2=0
cc_418 N_A_898_21#_c_654_n N_A_736_47#_M1020_g 0.00916492f $X=6.065 $Y=2.075
+ $X2=0 $Y2=0
cc_419 N_A_898_21#_c_649_n N_A_736_47#_c_765_n 0.00510146f $X=5.095 $Y=1.425
+ $X2=0 $Y2=0
cc_420 N_A_898_21#_c_652_n N_A_736_47#_c_765_n 0.00617577f $X=6.07 $Y=0.96 $X2=0
+ $Y2=0
cc_421 N_A_898_21#_c_654_n N_A_736_47#_c_765_n 0.0151164f $X=6.065 $Y=2.075
+ $X2=0 $Y2=0
cc_422 N_A_898_21#_c_650_n N_A_736_47#_M1002_g 0.0179332f $X=5.79 $Y=0.495 $X2=0
+ $Y2=0
cc_423 N_A_898_21#_c_650_n N_A_736_47#_c_767_n 0.00335137f $X=5.79 $Y=0.495
+ $X2=0 $Y2=0
cc_424 N_A_898_21#_c_651_n N_A_736_47#_c_767_n 0.00174617f $X=6.775 $Y=0.96
+ $X2=0 $Y2=0
cc_425 N_A_898_21#_c_652_n N_A_736_47#_c_767_n 0.00666812f $X=6.07 $Y=0.96 $X2=0
+ $Y2=0
cc_426 N_A_898_21#_c_653_n N_A_736_47#_c_767_n 0.0205728f $X=5.455 $Y=1.02 $X2=0
+ $Y2=0
cc_427 N_A_898_21#_M1015_g N_A_736_47#_c_779_n 0.0181307f $X=4.565 $Y=0.445
+ $X2=0 $Y2=0
cc_428 N_A_898_21#_M1009_g N_A_736_47#_c_787_n 0.0126256f $X=5.095 $Y=2.595
+ $X2=0 $Y2=0
cc_429 N_A_898_21#_M1015_g N_A_736_47#_c_768_n 0.011927f $X=4.565 $Y=0.445 $X2=0
+ $Y2=0
cc_430 N_A_898_21#_c_641_n N_A_736_47#_c_768_n 0.00342787f $X=4.97 $Y=0.93 $X2=0
+ $Y2=0
cc_431 N_A_898_21#_c_641_n N_A_736_47#_c_769_n 4.05506e-19 $X=4.97 $Y=0.93 $X2=0
+ $Y2=0
cc_432 N_A_898_21#_c_648_n N_A_736_47#_c_769_n 0.00751998f $X=5.045 $Y=1.02
+ $X2=0 $Y2=0
cc_433 N_A_898_21#_c_649_n N_A_736_47#_c_769_n 0.0133006f $X=5.095 $Y=1.425
+ $X2=0 $Y2=0
cc_434 N_A_898_21#_c_652_n N_A_736_47#_c_769_n 0.0109683f $X=6.07 $Y=0.96 $X2=0
+ $Y2=0
cc_435 N_A_898_21#_M1009_g N_A_736_47#_c_775_n 0.0133137f $X=5.095 $Y=2.595
+ $X2=0 $Y2=0
cc_436 N_A_898_21#_c_643_n N_A_736_47#_c_770_n 0.00413648f $X=5.095 $Y=1.55
+ $X2=0 $Y2=0
cc_437 N_A_898_21#_M1009_g N_A_736_47#_c_770_n 0.00912162f $X=5.095 $Y=2.595
+ $X2=0 $Y2=0
cc_438 N_A_898_21#_c_652_n N_A_736_47#_c_770_n 0.0239011f $X=6.07 $Y=0.96 $X2=0
+ $Y2=0
cc_439 N_A_898_21#_c_653_n N_A_736_47#_c_770_n 0.00454086f $X=5.455 $Y=1.02
+ $X2=0 $Y2=0
cc_440 N_A_898_21#_c_654_n N_A_736_47#_c_770_n 0.0238596f $X=6.065 $Y=2.075
+ $X2=0 $Y2=0
cc_441 N_A_898_21#_M1009_g N_A_736_47#_c_780_n 0.00302099f $X=5.095 $Y=2.595
+ $X2=0 $Y2=0
cc_442 N_A_898_21#_c_641_n N_A_736_47#_c_771_n 0.0122391f $X=4.97 $Y=0.93 $X2=0
+ $Y2=0
cc_443 N_A_898_21#_c_648_n N_A_736_47#_c_771_n 0.00739286f $X=5.045 $Y=1.02
+ $X2=0 $Y2=0
cc_444 N_A_898_21#_c_652_n N_A_736_47#_c_771_n 0.0130737f $X=6.07 $Y=0.96 $X2=0
+ $Y2=0
cc_445 N_A_898_21#_c_643_n N_A_736_47#_c_772_n 0.00191634f $X=5.095 $Y=1.55
+ $X2=0 $Y2=0
cc_446 N_A_898_21#_M1009_g N_A_736_47#_c_772_n 0.00312747f $X=5.095 $Y=2.595
+ $X2=0 $Y2=0
cc_447 N_A_898_21#_c_643_n N_A_736_47#_c_773_n 0.0214256f $X=5.095 $Y=1.55 $X2=0
+ $Y2=0
cc_448 N_A_898_21#_c_652_n N_A_736_47#_c_773_n 0.00702355f $X=6.07 $Y=0.96 $X2=0
+ $Y2=0
cc_449 N_A_898_21#_c_653_n N_A_736_47#_c_773_n 0.0101411f $X=5.455 $Y=1.02 $X2=0
+ $Y2=0
cc_450 N_A_898_21#_c_654_n N_A_736_47#_c_773_n 0.00979551f $X=6.065 $Y=2.075
+ $X2=0 $Y2=0
cc_451 N_A_898_21#_M1000_g N_RESET_B_c_874_n 0.0180746f $X=6.905 $Y=2.595 $X2=0
+ $Y2=0
cc_452 N_A_898_21#_M1000_g N_RESET_B_M1007_g 0.0145253f $X=6.905 $Y=2.595 $X2=0
+ $Y2=0
cc_453 N_A_898_21#_c_659_n N_RESET_B_M1007_g 0.0215506f $X=6.065 $Y=2.24 $X2=0
+ $Y2=0
cc_454 N_A_898_21#_M1012_g N_RESET_B_M1003_g 0.0313868f $X=6.825 $Y=0.495 $X2=0
+ $Y2=0
cc_455 N_A_898_21#_c_650_n N_RESET_B_M1003_g 0.0024651f $X=5.79 $Y=0.495 $X2=0
+ $Y2=0
cc_456 N_A_898_21#_c_651_n N_RESET_B_M1003_g 0.0142652f $X=6.775 $Y=0.96 $X2=0
+ $Y2=0
cc_457 N_A_898_21#_c_654_n N_RESET_B_M1003_g 0.00345813f $X=6.065 $Y=2.075 $X2=0
+ $Y2=0
cc_458 N_A_898_21#_c_655_n N_RESET_B_M1003_g 0.00106337f $X=6.94 $Y=1.04 $X2=0
+ $Y2=0
cc_459 N_A_898_21#_c_651_n N_RESET_B_c_876_n 0.00284447f $X=6.775 $Y=0.96 $X2=0
+ $Y2=0
cc_460 N_A_898_21#_c_654_n N_RESET_B_c_876_n 0.0080708f $X=6.065 $Y=2.075 $X2=0
+ $Y2=0
cc_461 N_A_898_21#_c_655_n N_RESET_B_c_876_n 3.4421e-19 $X=6.94 $Y=1.04 $X2=0
+ $Y2=0
cc_462 N_A_898_21#_c_656_n N_RESET_B_c_876_n 0.0205815f $X=6.94 $Y=1.04 $X2=0
+ $Y2=0
cc_463 N_A_898_21#_M1000_g N_RESET_B_c_877_n 0.00813402f $X=6.905 $Y=2.595 $X2=0
+ $Y2=0
cc_464 N_A_898_21#_c_651_n N_RESET_B_c_877_n 0.0258951f $X=6.775 $Y=0.96 $X2=0
+ $Y2=0
cc_465 N_A_898_21#_c_654_n N_RESET_B_c_877_n 0.0483207f $X=6.065 $Y=2.075 $X2=0
+ $Y2=0
cc_466 N_A_898_21#_c_655_n N_RESET_B_c_877_n 0.0243457f $X=6.94 $Y=1.04 $X2=0
+ $Y2=0
cc_467 N_A_898_21#_c_656_n N_RESET_B_c_877_n 0.00201853f $X=6.94 $Y=1.04 $X2=0
+ $Y2=0
cc_468 N_A_898_21#_M1009_g N_VPWR_c_917_n 0.0274295f $X=5.095 $Y=2.595 $X2=0
+ $Y2=0
cc_469 N_A_898_21#_c_659_n N_VPWR_c_917_n 0.0254641f $X=6.065 $Y=2.24 $X2=0
+ $Y2=0
cc_470 N_A_898_21#_c_659_n N_VPWR_c_918_n 0.0177952f $X=6.065 $Y=2.24 $X2=0
+ $Y2=0
cc_471 N_A_898_21#_M1000_g N_VPWR_c_919_n 0.00343102f $X=6.905 $Y=2.595 $X2=0
+ $Y2=0
cc_472 N_A_898_21#_c_659_n N_VPWR_c_919_n 0.0651988f $X=6.065 $Y=2.24 $X2=0
+ $Y2=0
cc_473 N_A_898_21#_c_656_n N_VPWR_c_919_n 2.98866e-19 $X=6.94 $Y=1.04 $X2=0
+ $Y2=0
cc_474 N_A_898_21#_M1009_g N_VPWR_c_921_n 0.00975641f $X=5.095 $Y=2.595 $X2=0
+ $Y2=0
cc_475 N_A_898_21#_M1000_g N_VPWR_c_922_n 0.00939541f $X=6.905 $Y=2.595 $X2=0
+ $Y2=0
cc_476 N_A_898_21#_M1020_d N_VPWR_c_914_n 0.00223819f $X=5.925 $Y=2.095 $X2=0
+ $Y2=0
cc_477 N_A_898_21#_M1009_g N_VPWR_c_914_n 0.0174579f $X=5.095 $Y=2.595 $X2=0
+ $Y2=0
cc_478 N_A_898_21#_M1000_g N_VPWR_c_914_n 0.0171101f $X=6.905 $Y=2.595 $X2=0
+ $Y2=0
cc_479 N_A_898_21#_c_659_n N_VPWR_c_914_n 0.0123247f $X=6.065 $Y=2.24 $X2=0
+ $Y2=0
cc_480 N_A_898_21#_M1000_g Q 0.017745f $X=6.905 $Y=2.595 $X2=0 $Y2=0
cc_481 N_A_898_21#_M1013_g Q 0.0274103f $X=7.185 $Y=0.495 $X2=0 $Y2=0
cc_482 N_A_898_21#_c_655_n Q 0.044913f $X=6.94 $Y=1.04 $X2=0 $Y2=0
cc_483 N_A_898_21#_M1000_g Q 0.0050851f $X=6.905 $Y=2.595 $X2=0 $Y2=0
cc_484 N_A_898_21#_c_655_n Q 0.00358608f $X=6.94 $Y=1.04 $X2=0 $Y2=0
cc_485 N_A_898_21#_c_656_n Q 0.00566388f $X=6.94 $Y=1.04 $X2=0 $Y2=0
cc_486 N_A_898_21#_M1000_g Q 0.0165125f $X=6.905 $Y=2.595 $X2=0 $Y2=0
cc_487 N_A_898_21#_M1015_g N_VGND_c_1021_n 0.00538803f $X=4.565 $Y=0.445 $X2=0
+ $Y2=0
cc_488 N_A_898_21#_c_648_n N_VGND_c_1021_n 0.00953038f $X=5.045 $Y=1.02 $X2=0
+ $Y2=0
cc_489 N_A_898_21#_c_650_n N_VGND_c_1021_n 0.027074f $X=5.79 $Y=0.495 $X2=0
+ $Y2=0
cc_490 N_A_898_21#_c_652_n N_VGND_c_1021_n 0.00704863f $X=6.07 $Y=0.96 $X2=0
+ $Y2=0
cc_491 N_A_898_21#_c_653_n N_VGND_c_1021_n 6.99172e-19 $X=5.455 $Y=1.02 $X2=0
+ $Y2=0
cc_492 N_A_898_21#_M1012_g N_VGND_c_1022_n 0.0122592f $X=6.825 $Y=0.495 $X2=0
+ $Y2=0
cc_493 N_A_898_21#_M1013_g N_VGND_c_1022_n 0.00208237f $X=7.185 $Y=0.495 $X2=0
+ $Y2=0
cc_494 N_A_898_21#_c_650_n N_VGND_c_1022_n 0.0174827f $X=5.79 $Y=0.495 $X2=0
+ $Y2=0
cc_495 N_A_898_21#_c_651_n N_VGND_c_1022_n 0.0207959f $X=6.775 $Y=0.96 $X2=0
+ $Y2=0
cc_496 N_A_898_21#_M1015_g N_VGND_c_1023_n 0.00366111f $X=4.565 $Y=0.445 $X2=0
+ $Y2=0
cc_497 N_A_898_21#_c_650_n N_VGND_c_1027_n 0.0293877f $X=5.79 $Y=0.495 $X2=0
+ $Y2=0
cc_498 N_A_898_21#_M1012_g N_VGND_c_1028_n 0.00445056f $X=6.825 $Y=0.495 $X2=0
+ $Y2=0
cc_499 N_A_898_21#_M1013_g N_VGND_c_1028_n 0.0053602f $X=7.185 $Y=0.495 $X2=0
+ $Y2=0
cc_500 N_A_898_21#_M1015_g N_VGND_c_1029_n 0.00675335f $X=4.565 $Y=0.445 $X2=0
+ $Y2=0
cc_501 N_A_898_21#_c_641_n N_VGND_c_1029_n 0.00408348f $X=4.97 $Y=0.93 $X2=0
+ $Y2=0
cc_502 N_A_898_21#_M1012_g N_VGND_c_1029_n 0.00796275f $X=6.825 $Y=0.495 $X2=0
+ $Y2=0
cc_503 N_A_898_21#_M1013_g N_VGND_c_1029_n 0.0109508f $X=7.185 $Y=0.495 $X2=0
+ $Y2=0
cc_504 N_A_898_21#_c_650_n N_VGND_c_1029_n 0.0165008f $X=5.79 $Y=0.495 $X2=0
+ $Y2=0
cc_505 N_A_898_21#_c_652_n N_VGND_c_1029_n 0.00831524f $X=6.07 $Y=0.96 $X2=0
+ $Y2=0
cc_506 N_A_736_47#_c_773_n N_RESET_B_c_874_n 0.0150673f $X=5.905 $Y=1.59 $X2=0
+ $Y2=0
cc_507 N_A_736_47#_c_765_n N_RESET_B_M1003_g 0.00776937f $X=5.905 $Y=1.425 $X2=0
+ $Y2=0
cc_508 N_A_736_47#_M1002_g N_RESET_B_M1003_g 0.0422714f $X=6.005 $Y=0.495 $X2=0
+ $Y2=0
cc_509 N_A_736_47#_M1020_g N_RESET_B_c_880_n 0.0332613f $X=5.8 $Y=2.595 $X2=0
+ $Y2=0
cc_510 N_A_736_47#_c_765_n N_RESET_B_c_876_n 0.0150673f $X=5.905 $Y=1.425 $X2=0
+ $Y2=0
cc_511 N_A_736_47#_c_765_n N_RESET_B_c_877_n 5.22268e-19 $X=5.905 $Y=1.425 $X2=0
+ $Y2=0
cc_512 N_A_736_47#_M1020_g N_VPWR_c_917_n 0.0105636f $X=5.8 $Y=2.595 $X2=0 $Y2=0
cc_513 N_A_736_47#_c_787_n N_VPWR_c_917_n 0.0133991f $X=4.94 $Y=2.28 $X2=0 $Y2=0
cc_514 N_A_736_47#_c_775_n N_VPWR_c_917_n 0.00849477f $X=5.025 $Y=2.195 $X2=0
+ $Y2=0
cc_515 N_A_736_47#_c_770_n N_VPWR_c_917_n 0.0178782f $X=5.595 $Y=1.59 $X2=0
+ $Y2=0
cc_516 N_A_736_47#_c_773_n N_VPWR_c_917_n 0.00403174f $X=5.905 $Y=1.59 $X2=0
+ $Y2=0
cc_517 N_A_736_47#_M1020_g N_VPWR_c_918_n 0.00939541f $X=5.8 $Y=2.595 $X2=0
+ $Y2=0
cc_518 N_A_736_47#_M1020_g N_VPWR_c_919_n 0.001289f $X=5.8 $Y=2.595 $X2=0 $Y2=0
cc_519 N_A_736_47#_c_780_n N_VPWR_c_921_n 0.0177952f $X=4.33 $Y=2.36 $X2=0 $Y2=0
cc_520 N_A_736_47#_M1019_d N_VPWR_c_914_n 0.00223819f $X=4.19 $Y=2.095 $X2=0
+ $Y2=0
cc_521 N_A_736_47#_M1020_g N_VPWR_c_914_n 0.0165358f $X=5.8 $Y=2.595 $X2=0 $Y2=0
cc_522 N_A_736_47#_c_780_n N_VPWR_c_914_n 0.0123247f $X=4.33 $Y=2.36 $X2=0 $Y2=0
cc_523 N_A_736_47#_c_787_n A_944_419# 0.0103783f $X=4.94 $Y=2.28 $X2=-0.19
+ $Y2=-0.245
cc_524 N_A_736_47#_c_779_n N_VGND_M1015_d 0.00531208f $X=4.7 $Y=0.42 $X2=0 $Y2=0
cc_525 N_A_736_47#_c_768_n N_VGND_M1015_d 0.00268423f $X=4.785 $Y=0.855 $X2=0
+ $Y2=0
cc_526 N_A_736_47#_c_779_n N_VGND_c_1020_n 0.00725122f $X=4.7 $Y=0.42 $X2=0
+ $Y2=0
cc_527 N_A_736_47#_M1002_g N_VGND_c_1021_n 0.00261211f $X=6.005 $Y=0.495 $X2=0
+ $Y2=0
cc_528 N_A_736_47#_c_779_n N_VGND_c_1021_n 0.0203998f $X=4.7 $Y=0.42 $X2=0 $Y2=0
cc_529 N_A_736_47#_c_768_n N_VGND_c_1021_n 0.00954491f $X=4.785 $Y=0.855 $X2=0
+ $Y2=0
cc_530 N_A_736_47#_c_771_n N_VGND_c_1021_n 0.00445552f $X=5.025 $Y=0.94 $X2=0
+ $Y2=0
cc_531 N_A_736_47#_M1002_g N_VGND_c_1022_n 0.00197525f $X=6.005 $Y=0.495 $X2=0
+ $Y2=0
cc_532 N_A_736_47#_c_779_n N_VGND_c_1023_n 0.0503659f $X=4.7 $Y=0.42 $X2=0 $Y2=0
cc_533 N_A_736_47#_M1002_g N_VGND_c_1027_n 0.00342832f $X=6.005 $Y=0.495 $X2=0
+ $Y2=0
cc_534 N_A_736_47#_M1011_d N_VGND_c_1029_n 0.00396812f $X=3.68 $Y=0.235 $X2=0
+ $Y2=0
cc_535 N_A_736_47#_M1002_g N_VGND_c_1029_n 0.00612558f $X=6.005 $Y=0.495 $X2=0
+ $Y2=0
cc_536 N_A_736_47#_c_779_n N_VGND_c_1029_n 0.0384731f $X=4.7 $Y=0.42 $X2=0 $Y2=0
cc_537 N_A_736_47#_c_771_n N_VGND_c_1029_n 0.00574849f $X=5.025 $Y=0.94 $X2=0
+ $Y2=0
cc_538 N_A_736_47#_c_779_n A_850_47# 0.00329503f $X=4.7 $Y=0.42 $X2=-0.19
+ $Y2=-0.245
cc_539 N_RESET_B_M1007_g N_VPWR_c_918_n 0.00840199f $X=6.33 $Y=2.595 $X2=0 $Y2=0
cc_540 N_RESET_B_M1007_g N_VPWR_c_919_n 0.0226999f $X=6.33 $Y=2.595 $X2=0 $Y2=0
cc_541 N_RESET_B_c_880_n N_VPWR_c_919_n 6.60569e-19 $X=6.372 $Y=1.895 $X2=0
+ $Y2=0
cc_542 N_RESET_B_c_877_n N_VPWR_c_919_n 0.0140375f $X=6.375 $Y=1.39 $X2=0 $Y2=0
cc_543 N_RESET_B_M1007_g N_VPWR_c_914_n 0.0136033f $X=6.33 $Y=2.595 $X2=0 $Y2=0
cc_544 N_RESET_B_M1007_g Q 2.76905e-19 $X=6.33 $Y=2.595 $X2=0 $Y2=0
cc_545 N_RESET_B_M1003_g N_VGND_c_1022_n 0.0110754f $X=6.395 $Y=0.495 $X2=0
+ $Y2=0
cc_546 N_RESET_B_M1003_g N_VGND_c_1027_n 0.00445056f $X=6.395 $Y=0.495 $X2=0
+ $Y2=0
cc_547 N_RESET_B_M1003_g N_VGND_c_1029_n 0.00804604f $X=6.395 $Y=0.495 $X2=0
+ $Y2=0
cc_548 N_VPWR_c_914_n A_740_419# 0.00353798f $X=7.44 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_549 N_VPWR_c_914_n A_944_419# 0.0107073f $X=7.44 $Y=3.33 $X2=-0.19 $Y2=-0.245
cc_550 N_VPWR_c_914_n N_Q_M1000_d 0.0023218f $X=7.44 $Y=3.33 $X2=0 $Y2=0
cc_551 N_VPWR_c_919_n Q 0.0306587f $X=6.595 $Y=2.24 $X2=0 $Y2=0
cc_552 N_VPWR_c_922_n Q 0.0352317f $X=7.44 $Y=3.33 $X2=0 $Y2=0
cc_553 N_VPWR_c_914_n Q 0.021402f $X=7.44 $Y=3.33 $X2=0 $Y2=0
cc_554 Q N_VGND_c_1022_n 0.00658623f $X=7.355 $Y=0.47 $X2=0 $Y2=0
cc_555 Q N_VGND_c_1028_n 0.0167213f $X=7.355 $Y=0.47 $X2=0 $Y2=0
cc_556 Q N_VGND_c_1029_n 0.0095959f $X=7.355 $Y=0.47 $X2=0 $Y2=0
cc_557 N_VGND_c_1029_n A_500_47# 0.00271994f $X=7.44 $Y=0 $X2=-0.19 $Y2=-0.245
cc_558 N_VGND_c_1029_n A_658_47# 0.0031085f $X=7.44 $Y=0 $X2=-0.19 $Y2=-0.245
cc_559 N_VGND_c_1029_n A_850_47# 0.00194865f $X=7.44 $Y=0 $X2=-0.19 $Y2=-0.245
