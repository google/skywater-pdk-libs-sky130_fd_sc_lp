* File: sky130_fd_sc_lp__a31o_m.pxi.spice
* Created: Wed Sep  2 09:26:43 2020
* 
x_PM_SKY130_FD_SC_LP__A31O_M%A_86_172# N_A_86_172#_M1001_d N_A_86_172#_M1007_d
+ N_A_86_172#_c_86_n N_A_86_172#_c_98_n N_A_86_172#_c_99_n N_A_86_172#_M1005_g
+ N_A_86_172#_M1000_g N_A_86_172#_c_87_n N_A_86_172#_c_88_n N_A_86_172#_c_89_n
+ N_A_86_172#_c_90_n N_A_86_172#_c_91_n N_A_86_172#_c_92_n N_A_86_172#_c_93_n
+ N_A_86_172#_c_94_n N_A_86_172#_c_95_n N_A_86_172#_c_96_n N_A_86_172#_c_102_n
+ PM_SKY130_FD_SC_LP__A31O_M%A_86_172#
x_PM_SKY130_FD_SC_LP__A31O_M%A3 N_A3_M1008_g N_A3_c_174_n N_A3_M1003_g
+ N_A3_c_175_n N_A3_c_176_n N_A3_c_182_n N_A3_c_177_n N_A3_c_183_n N_A3_c_184_n
+ A3 A3 A3 A3 N_A3_c_179_n PM_SKY130_FD_SC_LP__A31O_M%A3
x_PM_SKY130_FD_SC_LP__A31O_M%A2 N_A2_M1004_g N_A2_M1002_g N_A2_c_237_n
+ N_A2_c_242_n A2 A2 A2 N_A2_c_239_n PM_SKY130_FD_SC_LP__A31O_M%A2
x_PM_SKY130_FD_SC_LP__A31O_M%A1 N_A1_M1001_g N_A1_M1009_g N_A1_c_283_n
+ N_A1_c_284_n N_A1_c_285_n N_A1_c_286_n N_A1_c_291_n A1 A1 A1 N_A1_c_288_n
+ PM_SKY130_FD_SC_LP__A31O_M%A1
x_PM_SKY130_FD_SC_LP__A31O_M%B1 N_B1_c_336_n N_B1_M1006_g N_B1_M1007_g
+ N_B1_c_337_n N_B1_c_342_n N_B1_c_343_n N_B1_c_338_n B1 B1 B1 B1 N_B1_c_340_n
+ PM_SKY130_FD_SC_LP__A31O_M%B1
x_PM_SKY130_FD_SC_LP__A31O_M%X N_X_M1005_s N_X_M1000_s N_X_c_385_n N_X_c_386_n
+ N_X_c_387_n N_X_c_383_n X PM_SKY130_FD_SC_LP__A31O_M%X
x_PM_SKY130_FD_SC_LP__A31O_M%VPWR N_VPWR_M1000_d N_VPWR_M1002_d N_VPWR_c_412_n
+ N_VPWR_c_413_n N_VPWR_c_414_n N_VPWR_c_415_n N_VPWR_c_416_n N_VPWR_c_417_n
+ VPWR N_VPWR_c_418_n N_VPWR_c_411_n PM_SKY130_FD_SC_LP__A31O_M%VPWR
x_PM_SKY130_FD_SC_LP__A31O_M%A_274_512# N_A_274_512#_M1008_d
+ N_A_274_512#_M1009_d N_A_274_512#_c_451_n N_A_274_512#_c_452_n
+ N_A_274_512#_c_453_n N_A_274_512#_c_454_n N_A_274_512#_c_455_n
+ N_A_274_512#_c_471_n PM_SKY130_FD_SC_LP__A31O_M%A_274_512#
x_PM_SKY130_FD_SC_LP__A31O_M%VGND N_VGND_M1005_d N_VGND_M1006_d N_VGND_c_484_n
+ N_VGND_c_485_n N_VGND_c_486_n VGND N_VGND_c_487_n N_VGND_c_488_n
+ N_VGND_c_489_n N_VGND_c_490_n N_VGND_c_491_n PM_SKY130_FD_SC_LP__A31O_M%VGND
cc_1 VNB N_A_86_172#_c_86_n 0.00750025f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.16
cc_2 VNB N_A_86_172#_c_87_n 0.0216271f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=0.86
cc_3 VNB N_A_86_172#_c_88_n 0.0267019f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.01
cc_4 VNB N_A_86_172#_c_89_n 0.0169161f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=1.53
cc_5 VNB N_A_86_172#_c_90_n 0.0343755f $X=-0.19 $Y=-0.245 $X2=2.165 $Y2=0.945
cc_6 VNB N_A_86_172#_c_91_n 0.00200489f $X=-0.19 $Y=-0.245 $X2=2.27 $Y2=0.605
cc_7 VNB N_A_86_172#_c_92_n 0.0293025f $X=-0.19 $Y=-0.245 $X2=3.05 $Y2=0.945
cc_8 VNB N_A_86_172#_c_93_n 0.03006f $X=-0.19 $Y=-0.245 $X2=3.135 $Y2=2.67
cc_9 VNB N_A_86_172#_c_94_n 0.00231391f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=1.025
cc_10 VNB N_A_86_172#_c_95_n 0.027801f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=1.025
cc_11 VNB N_A_86_172#_c_96_n 0.00150062f $X=-0.19 $Y=-0.245 $X2=2.27 $Y2=0.945
cc_12 VNB N_A3_c_174_n 0.0174785f $X=-0.19 $Y=-0.245 $X2=0.79 $Y2=2.235
cc_13 VNB N_A3_c_175_n 0.0135151f $X=-0.19 $Y=-0.245 $X2=0.835 $Y2=0.54
cc_14 VNB N_A3_c_176_n 0.0171951f $X=-0.19 $Y=-0.245 $X2=0.865 $Y2=2.31
cc_15 VNB N_A3_c_177_n 0.0154511f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=1.01
cc_16 VNB A3 0.00140938f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=1.53
cc_17 VNB N_A3_c_179_n 0.0158229f $X=-0.19 $Y=-0.245 $X2=3.05 $Y2=0.945
cc_18 VNB N_A2_M1004_g 0.0348461f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A2_c_237_n 0.0163111f $X=-0.19 $Y=-0.245 $X2=0.835 $Y2=0.86
cc_20 VNB A2 5.95155e-19 $X=-0.19 $Y=-0.245 $X2=0.835 $Y2=0.54
cc_21 VNB N_A2_c_239_n 0.016141f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.01
cc_22 VNB N_A1_c_283_n 0.0168681f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=2.235
cc_23 VNB N_A1_c_284_n 0.0110092f $X=-0.19 $Y=-0.245 $X2=0.835 $Y2=0.86
cc_24 VNB N_A1_c_285_n 0.0136258f $X=-0.19 $Y=-0.245 $X2=0.835 $Y2=0.54
cc_25 VNB N_A1_c_286_n 0.0166021f $X=-0.19 $Y=-0.245 $X2=0.865 $Y2=2.31
cc_26 VNB A1 0.00124485f $X=-0.19 $Y=-0.245 $X2=0.865 $Y2=2.77
cc_27 VNB N_A1_c_288_n 0.0164567f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_B1_c_336_n 0.0216648f $X=-0.19 $Y=-0.245 $X2=2.13 $Y2=0.33
cc_29 VNB N_B1_c_337_n 0.0232971f $X=-0.19 $Y=-0.245 $X2=0.835 $Y2=0.54
cc_30 VNB N_B1_c_338_n 0.0370487f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=1.01
cc_31 VNB B1 0.00854373f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=0.86
cc_32 VNB N_B1_c_340_n 0.00674266f $X=-0.19 $Y=-0.245 $X2=2.27 $Y2=0.605
cc_33 VNB N_X_c_383_n 0.0251938f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB X 0.0470173f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.01
cc_35 VNB N_VPWR_c_411_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=0.945
cc_36 VNB N_VGND_c_484_n 0.00563551f $X=-0.19 $Y=-0.245 $X2=0.79 $Y2=2.235
cc_37 VNB N_VGND_c_485_n 0.0418526f $X=-0.19 $Y=-0.245 $X2=0.835 $Y2=0.86
cc_38 VNB N_VGND_c_486_n 0.00973164f $X=-0.19 $Y=-0.245 $X2=0.865 $Y2=2.77
cc_39 VNB N_VGND_c_487_n 0.0260718f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=0.86
cc_40 VNB N_VGND_c_488_n 0.0198045f $X=-0.19 $Y=-0.245 $X2=0.68 $Y2=0.945
cc_41 VNB N_VGND_c_489_n 0.211982f $X=-0.19 $Y=-0.245 $X2=2.27 $Y2=0.86
cc_42 VNB N_VGND_c_490_n 0.00587606f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_491_n 0.0040393f $X=-0.19 $Y=-0.245 $X2=3.135 $Y2=1.03
cc_44 VPB N_A_86_172#_c_86_n 0.037268f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=2.16
cc_45 VPB N_A_86_172#_c_98_n 0.0290759f $X=-0.19 $Y=1.655 $X2=0.79 $Y2=2.235
cc_46 VPB N_A_86_172#_c_99_n 0.0177735f $X=-0.19 $Y=1.655 $X2=0.58 $Y2=2.235
cc_47 VPB N_A_86_172#_M1000_g 0.0284917f $X=-0.19 $Y=1.655 $X2=0.865 $Y2=2.77
cc_48 VPB N_A_86_172#_c_93_n 0.0483019f $X=-0.19 $Y=1.655 $X2=3.135 $Y2=2.67
cc_49 VPB N_A_86_172#_c_102_n 0.0179461f $X=-0.19 $Y=1.655 $X2=2.8 $Y2=2.835
cc_50 VPB N_A3_M1008_g 0.0234632f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=1.53
cc_51 VPB N_A3_c_176_n 0.00743361f $X=-0.19 $Y=1.655 $X2=0.865 $Y2=2.31
cc_52 VPB N_A3_c_182_n 0.0196236f $X=-0.19 $Y=1.655 $X2=0.865 $Y2=2.77
cc_53 VPB N_A3_c_183_n 0.0140719f $X=-0.19 $Y=1.655 $X2=0.67 $Y2=1.01
cc_54 VPB N_A3_c_184_n 0.0138042f $X=-0.19 $Y=1.655 $X2=0.595 $Y2=1.365
cc_55 VPB A3 0.00620894f $X=-0.19 $Y=1.655 $X2=0.595 $Y2=1.53
cc_56 VPB N_A2_M1002_g 0.0438998f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=1.53
cc_57 VPB N_A2_c_237_n 0.00675646f $X=-0.19 $Y=1.655 $X2=0.835 $Y2=0.86
cc_58 VPB N_A2_c_242_n 0.0166436f $X=-0.19 $Y=1.655 $X2=0.835 $Y2=0.54
cc_59 VPB A2 0.00214549f $X=-0.19 $Y=1.655 $X2=0.835 $Y2=0.54
cc_60 VPB N_A1_M1009_g 0.0426935f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=2.16
cc_61 VPB N_A1_c_286_n 0.00687703f $X=-0.19 $Y=1.655 $X2=0.865 $Y2=2.31
cc_62 VPB N_A1_c_291_n 0.0168293f $X=-0.19 $Y=1.655 $X2=0.865 $Y2=2.77
cc_63 VPB A1 0.00374143f $X=-0.19 $Y=1.655 $X2=0.865 $Y2=2.77
cc_64 VPB N_B1_M1007_g 0.0304143f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_65 VPB N_B1_c_342_n 0.0260585f $X=-0.19 $Y=1.655 $X2=0.865 $Y2=2.77
cc_66 VPB N_B1_c_343_n 0.0263162f $X=-0.19 $Y=1.655 $X2=0.865 $Y2=2.77
cc_67 VPB B1 0.00804311f $X=-0.19 $Y=1.655 $X2=0.67 $Y2=0.86
cc_68 VPB N_B1_c_340_n 0.0104988f $X=-0.19 $Y=1.655 $X2=2.27 $Y2=0.605
cc_69 VPB N_X_c_385_n 0.00973547f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=1.53
cc_70 VPB N_X_c_386_n 0.0142304f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=2.16
cc_71 VPB N_X_c_387_n 0.0134524f $X=-0.19 $Y=1.655 $X2=0.835 $Y2=0.86
cc_72 VPB X 0.00254216f $X=-0.19 $Y=1.655 $X2=0.67 $Y2=1.01
cc_73 VPB N_VPWR_c_412_n 0.0028869f $X=-0.19 $Y=1.655 $X2=0.79 $Y2=2.235
cc_74 VPB N_VPWR_c_413_n 0.00700763f $X=-0.19 $Y=1.655 $X2=0.835 $Y2=0.54
cc_75 VPB N_VPWR_c_414_n 0.0297875f $X=-0.19 $Y=1.655 $X2=0.865 $Y2=2.77
cc_76 VPB N_VPWR_c_415_n 0.00577257f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_77 VPB N_VPWR_c_416_n 0.0167318f $X=-0.19 $Y=1.655 $X2=0.67 $Y2=0.86
cc_78 VPB N_VPWR_c_417_n 0.00362871f $X=-0.19 $Y=1.655 $X2=0.67 $Y2=1.01
cc_79 VPB N_VPWR_c_418_n 0.0390861f $X=-0.19 $Y=1.655 $X2=3.135 $Y2=2.67
cc_80 VPB N_VPWR_c_411_n 0.0809097f $X=-0.19 $Y=1.655 $X2=0.595 $Y2=0.945
cc_81 VPB N_A_274_512#_c_451_n 0.0140862f $X=-0.19 $Y=1.655 $X2=0.79 $Y2=2.235
cc_82 VPB N_A_274_512#_c_452_n 0.00433353f $X=-0.19 $Y=1.655 $X2=0.58 $Y2=2.235
cc_83 VPB N_A_274_512#_c_453_n 6.74103e-19 $X=-0.19 $Y=1.655 $X2=0.835 $Y2=0.54
cc_84 VPB N_A_274_512#_c_454_n 0.00210031f $X=-0.19 $Y=1.655 $X2=0.865 $Y2=2.31
cc_85 VPB N_A_274_512#_c_455_n 0.00118134f $X=-0.19 $Y=1.655 $X2=0.865 $Y2=2.77
cc_86 N_A_86_172#_M1000_g N_A3_M1008_g 0.0193886f $X=0.865 $Y=2.77 $X2=0 $Y2=0
cc_87 N_A_86_172#_c_87_n N_A3_c_174_n 0.0119323f $X=0.67 $Y=0.86 $X2=0 $Y2=0
cc_88 N_A_86_172#_c_90_n N_A3_c_175_n 0.00286917f $X=2.165 $Y=0.945 $X2=0 $Y2=0
cc_89 N_A_86_172#_c_94_n N_A3_c_175_n 9.63156e-19 $X=0.595 $Y=1.025 $X2=0 $Y2=0
cc_90 N_A_86_172#_c_95_n N_A3_c_175_n 0.00859942f $X=0.595 $Y=1.025 $X2=0 $Y2=0
cc_91 N_A_86_172#_c_86_n N_A3_c_176_n 0.0110703f $X=0.505 $Y=2.16 $X2=0 $Y2=0
cc_92 N_A_86_172#_c_89_n N_A3_c_176_n 0.00875151f $X=0.595 $Y=1.53 $X2=0 $Y2=0
cc_93 N_A_86_172#_c_88_n N_A3_c_177_n 0.00975607f $X=0.67 $Y=1.01 $X2=0 $Y2=0
cc_94 N_A_86_172#_c_90_n N_A3_c_177_n 0.0133494f $X=2.165 $Y=0.945 $X2=0 $Y2=0
cc_95 N_A_86_172#_c_86_n N_A3_c_183_n 0.00358572f $X=0.505 $Y=2.16 $X2=0 $Y2=0
cc_96 N_A_86_172#_c_98_n N_A3_c_184_n 0.00958522f $X=0.79 $Y=2.235 $X2=0 $Y2=0
cc_97 N_A_86_172#_c_86_n A3 0.00184691f $X=0.505 $Y=2.16 $X2=0 $Y2=0
cc_98 N_A_86_172#_c_98_n A3 0.00277992f $X=0.79 $Y=2.235 $X2=0 $Y2=0
cc_99 N_A_86_172#_c_90_n A3 0.0176418f $X=2.165 $Y=0.945 $X2=0 $Y2=0
cc_100 N_A_86_172#_c_94_n A3 0.0120293f $X=0.595 $Y=1.025 $X2=0 $Y2=0
cc_101 N_A_86_172#_c_95_n A3 0.00121806f $X=0.595 $Y=1.025 $X2=0 $Y2=0
cc_102 N_A_86_172#_c_90_n N_A3_c_179_n 0.00394381f $X=2.165 $Y=0.945 $X2=0 $Y2=0
cc_103 N_A_86_172#_c_94_n N_A3_c_179_n 9.09175e-19 $X=0.595 $Y=1.025 $X2=0 $Y2=0
cc_104 N_A_86_172#_c_95_n N_A3_c_179_n 0.00875151f $X=0.595 $Y=1.025 $X2=0 $Y2=0
cc_105 N_A_86_172#_c_90_n N_A2_M1004_g 0.0113707f $X=2.165 $Y=0.945 $X2=0 $Y2=0
cc_106 N_A_86_172#_c_90_n A2 0.0128266f $X=2.165 $Y=0.945 $X2=0 $Y2=0
cc_107 N_A_86_172#_c_90_n N_A2_c_239_n 0.0060732f $X=2.165 $Y=0.945 $X2=0 $Y2=0
cc_108 N_A_86_172#_c_91_n N_A1_c_283_n 0.00275684f $X=2.27 $Y=0.605 $X2=0 $Y2=0
cc_109 N_A_86_172#_c_90_n N_A1_c_284_n 0.00915793f $X=2.165 $Y=0.945 $X2=0 $Y2=0
cc_110 N_A_86_172#_c_96_n N_A1_c_284_n 0.00258457f $X=2.27 $Y=0.945 $X2=0 $Y2=0
cc_111 N_A_86_172#_c_90_n N_A1_c_285_n 0.00279016f $X=2.165 $Y=0.945 $X2=0 $Y2=0
cc_112 N_A_86_172#_c_96_n N_A1_c_285_n 8.66006e-19 $X=2.27 $Y=0.945 $X2=0 $Y2=0
cc_113 N_A_86_172#_c_90_n A1 0.00644157f $X=2.165 $Y=0.945 $X2=0 $Y2=0
cc_114 N_A_86_172#_c_96_n A1 0.0116089f $X=2.27 $Y=0.945 $X2=0 $Y2=0
cc_115 N_A_86_172#_c_96_n N_A1_c_288_n 0.00406005f $X=2.27 $Y=0.945 $X2=0 $Y2=0
cc_116 N_A_86_172#_c_91_n N_B1_c_336_n 0.00275684f $X=2.27 $Y=0.605 $X2=-0.19
+ $Y2=-0.245
cc_117 N_A_86_172#_c_93_n N_B1_M1007_g 0.00366515f $X=3.135 $Y=2.67 $X2=0 $Y2=0
cc_118 N_A_86_172#_c_102_n N_B1_M1007_g 7.68056e-19 $X=2.8 $Y=2.835 $X2=0 $Y2=0
cc_119 N_A_86_172#_c_92_n N_B1_c_337_n 0.0179466f $X=3.05 $Y=0.945 $X2=0 $Y2=0
cc_120 N_A_86_172#_c_102_n N_B1_c_343_n 0.00354466f $X=2.8 $Y=2.835 $X2=0 $Y2=0
cc_121 N_A_86_172#_c_92_n N_B1_c_338_n 0.00304397f $X=3.05 $Y=0.945 $X2=0 $Y2=0
cc_122 N_A_86_172#_c_93_n N_B1_c_338_n 0.0078232f $X=3.135 $Y=2.67 $X2=0 $Y2=0
cc_123 N_A_86_172#_c_92_n B1 0.0241304f $X=3.05 $Y=0.945 $X2=0 $Y2=0
cc_124 N_A_86_172#_c_93_n B1 0.0942646f $X=3.135 $Y=2.67 $X2=0 $Y2=0
cc_125 N_A_86_172#_c_102_n B1 0.0124276f $X=2.8 $Y=2.835 $X2=0 $Y2=0
cc_126 N_A_86_172#_c_92_n N_B1_c_340_n 0.00239773f $X=3.05 $Y=0.945 $X2=0 $Y2=0
cc_127 N_A_86_172#_c_93_n N_B1_c_340_n 0.0165869f $X=3.135 $Y=2.67 $X2=0 $Y2=0
cc_128 N_A_86_172#_c_86_n N_X_c_385_n 0.016618f $X=0.505 $Y=2.16 $X2=0 $Y2=0
cc_129 N_A_86_172#_c_89_n N_X_c_385_n 0.00234037f $X=0.595 $Y=1.53 $X2=0 $Y2=0
cc_130 N_A_86_172#_c_94_n N_X_c_385_n 0.0137049f $X=0.595 $Y=1.025 $X2=0 $Y2=0
cc_131 N_A_86_172#_c_86_n N_X_c_387_n 0.0149878f $X=0.505 $Y=2.16 $X2=0 $Y2=0
cc_132 N_A_86_172#_c_98_n N_X_c_387_n 0.0103878f $X=0.79 $Y=2.235 $X2=0 $Y2=0
cc_133 N_A_86_172#_c_99_n N_X_c_387_n 0.00703363f $X=0.58 $Y=2.235 $X2=0 $Y2=0
cc_134 N_A_86_172#_M1000_g N_X_c_387_n 0.00705012f $X=0.865 $Y=2.77 $X2=0 $Y2=0
cc_135 N_A_86_172#_c_88_n N_X_c_383_n 0.00586231f $X=0.67 $Y=1.01 $X2=0 $Y2=0
cc_136 N_A_86_172#_c_90_n N_X_c_383_n 0.00223064f $X=2.165 $Y=0.945 $X2=0 $Y2=0
cc_137 N_A_86_172#_c_94_n N_X_c_383_n 0.0130164f $X=0.595 $Y=1.025 $X2=0 $Y2=0
cc_138 N_A_86_172#_c_87_n X 0.00426332f $X=0.67 $Y=0.86 $X2=0 $Y2=0
cc_139 N_A_86_172#_c_88_n X 0.0231769f $X=0.67 $Y=1.01 $X2=0 $Y2=0
cc_140 N_A_86_172#_c_94_n X 0.0461949f $X=0.595 $Y=1.025 $X2=0 $Y2=0
cc_141 N_A_86_172#_M1000_g N_VPWR_c_412_n 0.0145198f $X=0.865 $Y=2.77 $X2=0
+ $Y2=0
cc_142 N_A_86_172#_M1000_g N_VPWR_c_414_n 0.00396895f $X=0.865 $Y=2.77 $X2=0
+ $Y2=0
cc_143 N_A_86_172#_c_102_n N_VPWR_c_418_n 0.0172889f $X=2.8 $Y=2.835 $X2=0 $Y2=0
cc_144 N_A_86_172#_M1000_g N_VPWR_c_411_n 0.00796233f $X=0.865 $Y=2.77 $X2=0
+ $Y2=0
cc_145 N_A_86_172#_c_102_n N_VPWR_c_411_n 0.0173002f $X=2.8 $Y=2.835 $X2=0 $Y2=0
cc_146 N_A_86_172#_c_93_n N_A_274_512#_c_453_n 0.00492616f $X=3.135 $Y=2.67
+ $X2=0 $Y2=0
cc_147 N_A_86_172#_c_87_n N_VGND_c_484_n 0.00909339f $X=0.67 $Y=0.86 $X2=0 $Y2=0
cc_148 N_A_86_172#_c_90_n N_VGND_c_484_n 0.0144194f $X=2.165 $Y=0.945 $X2=0
+ $Y2=0
cc_149 N_A_86_172#_c_91_n N_VGND_c_485_n 0.00590978f $X=2.27 $Y=0.605 $X2=0
+ $Y2=0
cc_150 N_A_86_172#_c_92_n N_VGND_c_486_n 0.0122803f $X=3.05 $Y=0.945 $X2=0 $Y2=0
cc_151 N_A_86_172#_c_87_n N_VGND_c_487_n 0.00477152f $X=0.67 $Y=0.86 $X2=0 $Y2=0
cc_152 N_A_86_172#_c_87_n N_VGND_c_489_n 0.00524756f $X=0.67 $Y=0.86 $X2=0 $Y2=0
cc_153 N_A_86_172#_c_88_n N_VGND_c_489_n 8.74901e-19 $X=0.67 $Y=1.01 $X2=0 $Y2=0
cc_154 N_A_86_172#_c_90_n N_VGND_c_489_n 0.0344595f $X=2.165 $Y=0.945 $X2=0
+ $Y2=0
cc_155 N_A_86_172#_c_91_n N_VGND_c_489_n 0.00721211f $X=2.27 $Y=0.605 $X2=0
+ $Y2=0
cc_156 N_A_86_172#_c_92_n N_VGND_c_489_n 0.0218844f $X=3.05 $Y=0.945 $X2=0 $Y2=0
cc_157 N_A3_c_174_n N_A2_M1004_g 0.0519416f $X=1.335 $Y=0.86 $X2=0 $Y2=0
cc_158 N_A3_c_175_n N_A2_M1004_g 0.00944401f $X=1.135 $Y=1.25 $X2=0 $Y2=0
cc_159 N_A3_c_183_n N_A2_M1002_g 0.00750819f $X=1.26 $Y=2.16 $X2=0 $Y2=0
cc_160 N_A3_c_184_n N_A2_M1002_g 0.0249544f $X=1.26 $Y=2.31 $X2=0 $Y2=0
cc_161 A3 N_A2_M1002_g 0.001448f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_162 N_A3_c_176_n N_A2_c_237_n 0.013805f $X=1.135 $Y=1.755 $X2=0 $Y2=0
cc_163 N_A3_c_182_n N_A2_c_242_n 0.013805f $X=1.135 $Y=1.92 $X2=0 $Y2=0
cc_164 N_A3_c_183_n A2 0.00124265f $X=1.26 $Y=2.16 $X2=0 $Y2=0
cc_165 A3 A2 0.0406968f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_166 N_A3_c_179_n A2 0.00209143f $X=1.135 $Y=1.415 $X2=0 $Y2=0
cc_167 A3 N_A2_c_239_n 0.0024142f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_168 N_A3_c_179_n N_A2_c_239_n 0.013805f $X=1.135 $Y=1.415 $X2=0 $Y2=0
cc_169 N_A3_c_176_n N_X_c_385_n 0.00156152f $X=1.135 $Y=1.755 $X2=0 $Y2=0
cc_170 A3 N_X_c_385_n 0.00871808f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_171 N_A3_c_182_n N_X_c_387_n 3.24239e-19 $X=1.135 $Y=1.92 $X2=0 $Y2=0
cc_172 N_A3_c_183_n N_X_c_387_n 7.96664e-19 $X=1.26 $Y=2.16 $X2=0 $Y2=0
cc_173 A3 N_X_c_387_n 0.0301555f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_174 N_A3_M1008_g N_VPWR_c_412_n 0.00710401f $X=1.295 $Y=2.77 $X2=0 $Y2=0
cc_175 N_A3_c_184_n N_VPWR_c_412_n 2.15039e-19 $X=1.26 $Y=2.31 $X2=0 $Y2=0
cc_176 A3 N_VPWR_c_412_n 0.0108099f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_177 N_A3_M1008_g N_VPWR_c_416_n 0.00396895f $X=1.295 $Y=2.77 $X2=0 $Y2=0
cc_178 N_A3_M1008_g N_VPWR_c_411_n 0.00653065f $X=1.295 $Y=2.77 $X2=0 $Y2=0
cc_179 A3 N_VPWR_c_411_n 0.0020961f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_180 N_A3_M1008_g N_A_274_512#_c_452_n 0.00129652f $X=1.295 $Y=2.77 $X2=0
+ $Y2=0
cc_181 A3 N_A_274_512#_c_452_n 0.0134205f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_182 N_A3_M1008_g N_A_274_512#_c_455_n 0.00393028f $X=1.295 $Y=2.77 $X2=0
+ $Y2=0
cc_183 N_A3_c_174_n N_VGND_c_484_n 0.00352506f $X=1.335 $Y=0.86 $X2=0 $Y2=0
cc_184 N_A3_c_177_n N_VGND_c_484_n 0.00276894f $X=1.335 $Y=0.935 $X2=0 $Y2=0
cc_185 N_A3_c_174_n N_VGND_c_485_n 0.00495161f $X=1.335 $Y=0.86 $X2=0 $Y2=0
cc_186 N_A3_c_174_n N_VGND_c_489_n 0.00527891f $X=1.335 $Y=0.86 $X2=0 $Y2=0
cc_187 N_A3_c_177_n N_VGND_c_489_n 6.57583e-19 $X=1.335 $Y=0.935 $X2=0 $Y2=0
cc_188 N_A2_M1002_g N_A1_M1009_g 0.0371223f $X=1.725 $Y=2.77 $X2=0 $Y2=0
cc_189 A2 N_A1_M1009_g 2.44944e-19 $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_190 N_A2_M1004_g N_A1_c_283_n 0.0516143f $X=1.695 $Y=0.54 $X2=0 $Y2=0
cc_191 N_A2_M1004_g N_A1_c_285_n 0.0115219f $X=1.695 $Y=0.54 $X2=0 $Y2=0
cc_192 A2 N_A1_c_285_n 0.00225314f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_193 N_A2_c_237_n N_A1_c_286_n 0.0138165f $X=1.675 $Y=1.755 $X2=0 $Y2=0
cc_194 N_A2_c_242_n N_A1_c_291_n 0.0138165f $X=1.675 $Y=1.92 $X2=0 $Y2=0
cc_195 N_A2_M1002_g A1 0.00120362f $X=1.725 $Y=2.77 $X2=0 $Y2=0
cc_196 A2 A1 0.0397158f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_197 N_A2_c_239_n A1 0.00236757f $X=1.675 $Y=1.415 $X2=0 $Y2=0
cc_198 N_A2_c_239_n N_A1_c_288_n 0.0138165f $X=1.675 $Y=1.415 $X2=0 $Y2=0
cc_199 N_A2_M1002_g N_VPWR_c_412_n 4.22719e-19 $X=1.725 $Y=2.77 $X2=0 $Y2=0
cc_200 N_A2_M1002_g N_VPWR_c_413_n 0.00153144f $X=1.725 $Y=2.77 $X2=0 $Y2=0
cc_201 N_A2_M1002_g N_VPWR_c_416_n 0.00478016f $X=1.725 $Y=2.77 $X2=0 $Y2=0
cc_202 N_A2_M1002_g N_VPWR_c_411_n 0.00494571f $X=1.725 $Y=2.77 $X2=0 $Y2=0
cc_203 N_A2_M1002_g N_A_274_512#_c_451_n 0.0124784f $X=1.725 $Y=2.77 $X2=0 $Y2=0
cc_204 N_A2_c_242_n N_A_274_512#_c_451_n 0.00135248f $X=1.675 $Y=1.92 $X2=0
+ $Y2=0
cc_205 A2 N_A_274_512#_c_451_n 0.00871491f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_206 N_A2_c_242_n N_A_274_512#_c_452_n 0.00324522f $X=1.675 $Y=1.92 $X2=0
+ $Y2=0
cc_207 A2 N_A_274_512#_c_452_n 0.00367309f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_208 N_A2_M1002_g N_A_274_512#_c_453_n 4.75542e-19 $X=1.725 $Y=2.77 $X2=0
+ $Y2=0
cc_209 N_A2_M1002_g N_A_274_512#_c_455_n 0.00142278f $X=1.725 $Y=2.77 $X2=0
+ $Y2=0
cc_210 N_A2_M1004_g N_VGND_c_485_n 0.00495161f $X=1.695 $Y=0.54 $X2=0 $Y2=0
cc_211 N_A2_M1004_g N_VGND_c_489_n 0.0053101f $X=1.695 $Y=0.54 $X2=0 $Y2=0
cc_212 N_A1_c_283_n N_B1_c_336_n 0.0136837f $X=2.09 $Y=0.86 $X2=-0.19 $Y2=-0.245
cc_213 N_A1_c_284_n N_B1_c_337_n 0.00972223f $X=2.09 $Y=1.01 $X2=0 $Y2=0
cc_214 N_A1_M1009_g N_B1_c_342_n 0.00680517f $X=2.155 $Y=2.77 $X2=0 $Y2=0
cc_215 N_A1_c_291_n N_B1_c_342_n 0.0117132f $X=2.215 $Y=1.92 $X2=0 $Y2=0
cc_216 A1 N_B1_c_342_n 6.61674e-19 $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_217 N_A1_M1009_g N_B1_c_343_n 0.0247701f $X=2.155 $Y=2.77 $X2=0 $Y2=0
cc_218 N_A1_c_285_n N_B1_c_338_n 0.00783838f $X=2.215 $Y=1.25 $X2=0 $Y2=0
cc_219 A1 N_B1_c_338_n 8.20913e-19 $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_220 N_A1_c_288_n N_B1_c_338_n 0.0117132f $X=2.215 $Y=1.415 $X2=0 $Y2=0
cc_221 N_A1_M1009_g B1 0.00257873f $X=2.155 $Y=2.77 $X2=0 $Y2=0
cc_222 A1 B1 0.0525447f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_223 N_A1_c_288_n B1 0.00472782f $X=2.215 $Y=1.415 $X2=0 $Y2=0
cc_224 N_A1_c_286_n N_B1_c_340_n 0.0117132f $X=2.215 $Y=1.755 $X2=0 $Y2=0
cc_225 N_A1_M1009_g N_VPWR_c_413_n 0.0030534f $X=2.155 $Y=2.77 $X2=0 $Y2=0
cc_226 N_A1_M1009_g N_VPWR_c_418_n 0.00451107f $X=2.155 $Y=2.77 $X2=0 $Y2=0
cc_227 N_A1_M1009_g N_VPWR_c_411_n 0.00480605f $X=2.155 $Y=2.77 $X2=0 $Y2=0
cc_228 N_A1_M1009_g N_A_274_512#_c_451_n 0.0106452f $X=2.155 $Y=2.77 $X2=0 $Y2=0
cc_229 N_A1_c_291_n N_A_274_512#_c_451_n 0.00380923f $X=2.215 $Y=1.92 $X2=0
+ $Y2=0
cc_230 A1 N_A_274_512#_c_451_n 0.0158818f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_231 N_A1_M1009_g N_A_274_512#_c_453_n 0.00403149f $X=2.155 $Y=2.77 $X2=0
+ $Y2=0
cc_232 N_A1_M1009_g N_A_274_512#_c_471_n 0.00258817f $X=2.155 $Y=2.77 $X2=0
+ $Y2=0
cc_233 N_A1_c_283_n N_VGND_c_485_n 0.00495161f $X=2.09 $Y=0.86 $X2=0 $Y2=0
cc_234 N_A1_c_283_n N_VGND_c_489_n 0.00537285f $X=2.09 $Y=0.86 $X2=0 $Y2=0
cc_235 N_A1_c_284_n N_VGND_c_489_n 8.97103e-19 $X=2.09 $Y=1.01 $X2=0 $Y2=0
cc_236 N_B1_M1007_g N_VPWR_c_418_n 0.00451107f $X=2.585 $Y=2.77 $X2=0 $Y2=0
cc_237 N_B1_M1007_g N_VPWR_c_411_n 0.00569702f $X=2.585 $Y=2.77 $X2=0 $Y2=0
cc_238 B1 N_VPWR_c_411_n 0.00576653f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_239 N_B1_M1007_g N_A_274_512#_c_451_n 0.00119549f $X=2.585 $Y=2.77 $X2=0
+ $Y2=0
cc_240 B1 N_A_274_512#_c_451_n 0.0136882f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_241 N_B1_M1007_g N_A_274_512#_c_453_n 0.00168828f $X=2.585 $Y=2.77 $X2=0
+ $Y2=0
cc_242 N_B1_M1007_g N_A_274_512#_c_471_n 0.00365784f $X=2.585 $Y=2.77 $X2=0
+ $Y2=0
cc_243 N_B1_c_336_n N_VGND_c_485_n 0.00495161f $X=2.485 $Y=0.86 $X2=0 $Y2=0
cc_244 N_B1_c_336_n N_VGND_c_486_n 0.00500444f $X=2.485 $Y=0.86 $X2=0 $Y2=0
cc_245 N_B1_c_337_n N_VGND_c_486_n 0.00435962f $X=2.695 $Y=0.935 $X2=0 $Y2=0
cc_246 N_B1_c_336_n N_VGND_c_489_n 0.00574769f $X=2.485 $Y=0.86 $X2=0 $Y2=0
cc_247 N_B1_c_337_n N_VGND_c_489_n 7.25333e-19 $X=2.695 $Y=0.935 $X2=0 $Y2=0
cc_248 N_X_c_387_n N_VPWR_c_414_n 0.0055846f $X=0.65 $Y=2.705 $X2=0 $Y2=0
cc_249 N_X_c_387_n N_VPWR_c_411_n 0.00645943f $X=0.65 $Y=2.705 $X2=0 $Y2=0
cc_250 N_X_c_383_n N_VGND_c_487_n 0.0234097f $X=0.62 $Y=0.515 $X2=0 $Y2=0
cc_251 N_X_c_383_n N_VGND_c_489_n 0.0205489f $X=0.62 $Y=0.515 $X2=0 $Y2=0
cc_252 N_VPWR_c_413_n N_A_274_512#_c_451_n 0.01357f $X=1.94 $Y=2.835 $X2=0 $Y2=0
cc_253 N_VPWR_c_411_n N_A_274_512#_c_451_n 0.0118197f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_254 N_VPWR_c_412_n N_A_274_512#_c_454_n 0.0103861f $X=1.08 $Y=2.835 $X2=0
+ $Y2=0
cc_255 N_VPWR_c_413_n N_A_274_512#_c_454_n 0.0013068f $X=1.94 $Y=2.835 $X2=0
+ $Y2=0
cc_256 N_VPWR_c_416_n N_A_274_512#_c_454_n 0.00999378f $X=1.835 $Y=3.33 $X2=0
+ $Y2=0
cc_257 N_VPWR_c_411_n N_A_274_512#_c_454_n 0.00774102f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_258 N_VPWR_c_418_n N_A_274_512#_c_471_n 0.00789072f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_259 N_VPWR_c_411_n N_A_274_512#_c_471_n 0.0106694f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
