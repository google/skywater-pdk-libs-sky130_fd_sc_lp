* File: sky130_fd_sc_lp__a21o_m.pxi.spice
* Created: Fri Aug 28 09:51:23 2020
* 
x_PM_SKY130_FD_SC_LP__A21O_M%A_80_153# N_A_80_153#_M1001_d N_A_80_153#_M1005_s
+ N_A_80_153#_c_68_n N_A_80_153#_M1004_g N_A_80_153#_c_62_n N_A_80_153#_M1007_g
+ N_A_80_153#_c_63_n N_A_80_153#_c_70_n N_A_80_153#_c_64_n N_A_80_153#_c_72_n
+ N_A_80_153#_c_65_n N_A_80_153#_c_104_p N_A_80_153#_c_73_n N_A_80_153#_c_74_n
+ N_A_80_153#_c_75_n N_A_80_153#_c_66_n N_A_80_153#_c_67_n
+ PM_SKY130_FD_SC_LP__A21O_M%A_80_153#
x_PM_SKY130_FD_SC_LP__A21O_M%B1 N_B1_M1001_g N_B1_M1005_g N_B1_c_136_n
+ N_B1_c_141_n B1 B1 B1 N_B1_c_138_n PM_SKY130_FD_SC_LP__A21O_M%B1
x_PM_SKY130_FD_SC_LP__A21O_M%A1 N_A1_M1006_g N_A1_M1002_g A1 A1 A1 A1
+ N_A1_c_184_n PM_SKY130_FD_SC_LP__A21O_M%A1
x_PM_SKY130_FD_SC_LP__A21O_M%A2 N_A2_c_227_n N_A2_M1003_g N_A2_c_228_n
+ N_A2_c_229_n N_A2_M1000_g N_A2_c_231_n A2 A2 A2 A2 A2 N_A2_c_233_n
+ PM_SKY130_FD_SC_LP__A21O_M%A2
x_PM_SKY130_FD_SC_LP__A21O_M%X N_X_M1007_s N_X_M1004_s X X X X X X X N_X_c_262_n
+ PM_SKY130_FD_SC_LP__A21O_M%X
x_PM_SKY130_FD_SC_LP__A21O_M%VPWR N_VPWR_M1004_d N_VPWR_M1002_d N_VPWR_c_280_n
+ N_VPWR_c_281_n VPWR N_VPWR_c_282_n N_VPWR_c_283_n N_VPWR_c_284_n
+ N_VPWR_c_279_n N_VPWR_c_286_n N_VPWR_c_287_n PM_SKY130_FD_SC_LP__A21O_M%VPWR
x_PM_SKY130_FD_SC_LP__A21O_M%A_324_508# N_A_324_508#_M1005_d
+ N_A_324_508#_M1000_d N_A_324_508#_c_317_n N_A_324_508#_c_318_n
+ N_A_324_508#_c_319_n N_A_324_508#_c_320_n
+ PM_SKY130_FD_SC_LP__A21O_M%A_324_508#
x_PM_SKY130_FD_SC_LP__A21O_M%VGND N_VGND_M1007_d N_VGND_M1003_d N_VGND_c_340_n
+ N_VGND_c_341_n N_VGND_c_342_n N_VGND_c_343_n VGND N_VGND_c_344_n
+ N_VGND_c_345_n N_VGND_c_346_n N_VGND_c_347_n PM_SKY130_FD_SC_LP__A21O_M%VGND
cc_1 VNB N_A_80_153#_c_62_n 0.0197916f $X=-0.19 $Y=-0.245 $X2=0.745 $Y2=0.765
cc_2 VNB N_A_80_153#_c_63_n 0.0272277f $X=-0.19 $Y=-0.245 $X2=0.745 $Y2=0.84
cc_3 VNB N_A_80_153#_c_64_n 0.00600621f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=2.01
cc_4 VNB N_A_80_153#_c_65_n 0.0248718f $X=-0.19 $Y=-0.245 $X2=1.285 $Y2=0.945
cc_5 VNB N_A_80_153#_c_66_n 0.00434797f $X=-0.19 $Y=-0.245 $X2=1.39 $Y2=0.495
cc_6 VNB N_A_80_153#_c_67_n 0.0411125f $X=-0.19 $Y=-0.245 $X2=0.587 $Y2=1.845
cc_7 VNB N_B1_M1001_g 0.053953f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_B1_c_136_n 0.00298644f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.885
cc_9 VNB B1 0.00516995f $X=-0.19 $Y=-0.245 $X2=0.745 $Y2=0.445
cc_10 VNB N_B1_c_138_n 0.01806f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.03
cc_11 VNB N_A1_M1006_g 0.0388458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB A1 0.00995783f $X=-0.19 $Y=-0.245 $X2=0.587 $Y2=2.032
cc_13 VNB N_A1_c_184_n 0.054544f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.84
cc_14 VNB N_A2_c_227_n 0.0186666f $X=-0.19 $Y=-0.245 $X2=1.25 $Y2=0.235
cc_15 VNB N_A2_c_228_n 0.0511701f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A2_c_229_n 0.00616447f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A2_M1000_g 0.0122616f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.845
cc_18 VNB N_A2_c_231_n 0.0374543f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.885
cc_19 VNB A2 0.0264813f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.885
cc_20 VNB N_A2_c_233_n 0.0377282f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=2.345
cc_21 VNB X 0.0480026f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.845
cc_22 VNB N_X_c_262_n 0.0228066f $X=-0.19 $Y=-0.245 $X2=0.587 $Y2=1.845
cc_23 VNB N_VPWR_c_279_n 0.123877f $X=-0.19 $Y=-0.245 $X2=1.225 $Y2=2.43
cc_24 VNB N_VGND_c_340_n 0.00494119f $X=-0.19 $Y=-0.245 $X2=0.587 $Y2=2.032
cc_25 VNB N_VGND_c_341_n 0.0123364f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.885
cc_26 VNB N_VGND_c_342_n 0.0255669f $X=-0.19 $Y=-0.245 $X2=0.745 $Y2=0.445
cc_27 VNB N_VGND_c_343_n 0.00401177f $X=-0.19 $Y=-0.245 $X2=0.745 $Y2=0.445
cc_28 VNB N_VGND_c_344_n 0.0274307f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=2.345
cc_29 VNB N_VGND_c_345_n 0.0179462f $X=-0.19 $Y=-0.245 $X2=1.225 $Y2=2.43
cc_30 VNB N_VGND_c_346_n 0.178943f $X=-0.19 $Y=-0.245 $X2=0.695 $Y2=2.43
cc_31 VNB N_VGND_c_347_n 0.00510247f $X=-0.19 $Y=-0.245 $X2=1.33 $Y2=2.685
cc_32 VPB N_A_80_153#_c_68_n 0.0252814f $X=-0.19 $Y=1.655 $X2=0.587 $Y2=2.328
cc_33 VPB N_A_80_153#_M1004_g 0.0260263f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.885
cc_34 VPB N_A_80_153#_c_70_n 0.0228317f $X=-0.19 $Y=1.655 $X2=0.587 $Y2=2.515
cc_35 VPB N_A_80_153#_c_64_n 0.0016077f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=2.01
cc_36 VPB N_A_80_153#_c_72_n 0.0235292f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=2.01
cc_37 VPB N_A_80_153#_c_73_n 0.0223003f $X=-0.19 $Y=1.655 $X2=1.225 $Y2=2.43
cc_38 VPB N_A_80_153#_c_74_n 0.00164639f $X=-0.19 $Y=1.655 $X2=0.695 $Y2=2.43
cc_39 VPB N_A_80_153#_c_75_n 6.94659e-19 $X=-0.19 $Y=1.655 $X2=1.33 $Y2=2.685
cc_40 VPB N_A_80_153#_c_67_n 0.00923156f $X=-0.19 $Y=1.655 $X2=0.587 $Y2=1.845
cc_41 VPB N_B1_M1005_g 0.0344459f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.915
cc_42 VPB N_B1_c_136_n 0.0326408f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.885
cc_43 VPB N_B1_c_141_n 0.0402369f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_44 VPB N_A1_M1002_g 0.0474009f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.915
cc_45 VPB A1 0.00942861f $X=-0.19 $Y=1.655 $X2=0.587 $Y2=2.032
cc_46 VPB N_A1_c_184_n 0.0256449f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.84
cc_47 VPB N_A2_M1000_g 0.0702391f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=1.845
cc_48 VPB A2 0.0247697f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.885
cc_49 VPB X 0.0491517f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=1.845
cc_50 VPB N_VPWR_c_280_n 0.00747396f $X=-0.19 $Y=1.655 $X2=0.587 $Y2=2.032
cc_51 VPB N_VPWR_c_281_n 0.00856386f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.885
cc_52 VPB N_VPWR_c_282_n 0.0163199f $X=-0.19 $Y=1.655 $X2=0.745 $Y2=0.445
cc_53 VPB N_VPWR_c_283_n 0.0365605f $X=-0.19 $Y=1.655 $X2=0.587 $Y2=2.515
cc_54 VPB N_VPWR_c_284_n 0.0195007f $X=-0.19 $Y=1.655 $X2=0.695 $Y2=0.945
cc_55 VPB N_VPWR_c_279_n 0.0631636f $X=-0.19 $Y=1.655 $X2=1.225 $Y2=2.43
cc_56 VPB N_VPWR_c_286_n 0.00510247f $X=-0.19 $Y=1.655 $X2=1.33 $Y2=2.685
cc_57 VPB N_VPWR_c_287_n 0.00401341f $X=-0.19 $Y=1.655 $X2=1.39 $Y2=0.86
cc_58 VPB N_A_324_508#_c_317_n 0.00116345f $X=-0.19 $Y=1.655 $X2=0.587 $Y2=2.032
cc_59 VPB N_A_324_508#_c_318_n 0.020104f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.515
cc_60 VPB N_A_324_508#_c_319_n 0.00425042f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.885
cc_61 VPB N_A_324_508#_c_320_n 0.00317049f $X=-0.19 $Y=1.655 $X2=0.745 $Y2=0.765
cc_62 N_A_80_153#_c_62_n N_B1_M1001_g 0.0220544f $X=0.745 $Y=0.765 $X2=0 $Y2=0
cc_63 N_A_80_153#_c_64_n N_B1_M1001_g 0.00401547f $X=0.61 $Y=2.01 $X2=0 $Y2=0
cc_64 N_A_80_153#_c_65_n N_B1_M1001_g 0.0129809f $X=1.285 $Y=0.945 $X2=0 $Y2=0
cc_65 N_A_80_153#_c_66_n N_B1_M1001_g 0.00497181f $X=1.39 $Y=0.495 $X2=0 $Y2=0
cc_66 N_A_80_153#_c_67_n N_B1_M1001_g 0.00709221f $X=0.587 $Y=1.845 $X2=0 $Y2=0
cc_67 N_A_80_153#_c_68_n N_B1_M1005_g 0.0045766f $X=0.587 $Y=2.328 $X2=0 $Y2=0
cc_68 N_A_80_153#_c_73_n N_B1_M1005_g 0.00242153f $X=1.225 $Y=2.43 $X2=0 $Y2=0
cc_69 N_A_80_153#_c_75_n N_B1_M1005_g 5.77961e-19 $X=1.33 $Y=2.685 $X2=0 $Y2=0
cc_70 N_A_80_153#_c_64_n N_B1_c_136_n 0.00152629f $X=0.61 $Y=2.01 $X2=0 $Y2=0
cc_71 N_A_80_153#_c_72_n N_B1_c_136_n 0.0118864f $X=0.61 $Y=2.01 $X2=0 $Y2=0
cc_72 N_A_80_153#_c_68_n N_B1_c_141_n 0.0118864f $X=0.587 $Y=2.328 $X2=0 $Y2=0
cc_73 N_A_80_153#_c_73_n N_B1_c_141_n 0.0160494f $X=1.225 $Y=2.43 $X2=0 $Y2=0
cc_74 N_A_80_153#_c_64_n B1 0.0365834f $X=0.61 $Y=2.01 $X2=0 $Y2=0
cc_75 N_A_80_153#_c_72_n B1 9.19168e-19 $X=0.61 $Y=2.01 $X2=0 $Y2=0
cc_76 N_A_80_153#_c_65_n B1 0.0160209f $X=1.285 $Y=0.945 $X2=0 $Y2=0
cc_77 N_A_80_153#_c_73_n B1 0.0140828f $X=1.225 $Y=2.43 $X2=0 $Y2=0
cc_78 N_A_80_153#_c_67_n B1 0.001042f $X=0.587 $Y=1.845 $X2=0 $Y2=0
cc_79 N_A_80_153#_c_64_n N_B1_c_138_n 0.0044118f $X=0.61 $Y=2.01 $X2=0 $Y2=0
cc_80 N_A_80_153#_c_65_n N_B1_c_138_n 0.00413135f $X=1.285 $Y=0.945 $X2=0 $Y2=0
cc_81 N_A_80_153#_c_67_n N_B1_c_138_n 0.00704451f $X=0.587 $Y=1.845 $X2=0 $Y2=0
cc_82 N_A_80_153#_c_65_n N_A1_M1006_g 0.00190264f $X=1.285 $Y=0.945 $X2=0 $Y2=0
cc_83 N_A_80_153#_c_66_n N_A1_M1006_g 0.00487883f $X=1.39 $Y=0.495 $X2=0 $Y2=0
cc_84 N_A_80_153#_c_65_n A1 0.0102014f $X=1.285 $Y=0.945 $X2=0 $Y2=0
cc_85 N_A_80_153#_c_66_n A1 0.00107079f $X=1.39 $Y=0.495 $X2=0 $Y2=0
cc_86 N_A_80_153#_c_62_n X 0.00263206f $X=0.745 $Y=0.765 $X2=0 $Y2=0
cc_87 N_A_80_153#_c_63_n X 0.0517809f $X=0.745 $Y=0.84 $X2=0 $Y2=0
cc_88 N_A_80_153#_c_64_n X 0.0907352f $X=0.61 $Y=2.01 $X2=0 $Y2=0
cc_89 N_A_80_153#_c_104_p X 0.0130705f $X=0.695 $Y=0.945 $X2=0 $Y2=0
cc_90 N_A_80_153#_c_74_n X 0.0131107f $X=0.695 $Y=2.43 $X2=0 $Y2=0
cc_91 N_A_80_153#_c_62_n N_X_c_262_n 5.77639e-19 $X=0.745 $Y=0.765 $X2=0 $Y2=0
cc_92 N_A_80_153#_c_63_n N_X_c_262_n 0.00863138f $X=0.745 $Y=0.84 $X2=0 $Y2=0
cc_93 N_A_80_153#_c_104_p N_X_c_262_n 0.00840428f $X=0.695 $Y=0.945 $X2=0 $Y2=0
cc_94 N_A_80_153#_c_66_n N_X_c_262_n 5.74754e-19 $X=1.39 $Y=0.495 $X2=0 $Y2=0
cc_95 N_A_80_153#_M1004_g N_VPWR_c_280_n 0.0123931f $X=0.475 $Y=2.885 $X2=0
+ $Y2=0
cc_96 N_A_80_153#_c_70_n N_VPWR_c_280_n 0.00271264f $X=0.587 $Y=2.515 $X2=0
+ $Y2=0
cc_97 N_A_80_153#_c_73_n N_VPWR_c_280_n 0.00702913f $X=1.225 $Y=2.43 $X2=0 $Y2=0
cc_98 N_A_80_153#_c_74_n N_VPWR_c_280_n 0.00618126f $X=0.695 $Y=2.43 $X2=0 $Y2=0
cc_99 N_A_80_153#_c_75_n N_VPWR_c_280_n 2.27411e-19 $X=1.33 $Y=2.685 $X2=0 $Y2=0
cc_100 N_A_80_153#_M1004_g N_VPWR_c_282_n 0.00486043f $X=0.475 $Y=2.885 $X2=0
+ $Y2=0
cc_101 N_A_80_153#_c_75_n N_VPWR_c_283_n 0.00546891f $X=1.33 $Y=2.685 $X2=0
+ $Y2=0
cc_102 N_A_80_153#_M1004_g N_VPWR_c_279_n 0.0093594f $X=0.475 $Y=2.885 $X2=0
+ $Y2=0
cc_103 N_A_80_153#_c_73_n N_VPWR_c_279_n 0.0137674f $X=1.225 $Y=2.43 $X2=0 $Y2=0
cc_104 N_A_80_153#_c_74_n N_VPWR_c_279_n 8.01572e-19 $X=0.695 $Y=2.43 $X2=0
+ $Y2=0
cc_105 N_A_80_153#_c_75_n N_VPWR_c_279_n 0.00697209f $X=1.33 $Y=2.685 $X2=0
+ $Y2=0
cc_106 N_A_80_153#_c_73_n N_A_324_508#_c_317_n 0.00317988f $X=1.225 $Y=2.43
+ $X2=0 $Y2=0
cc_107 N_A_80_153#_c_75_n N_A_324_508#_c_317_n 0.00152375f $X=1.33 $Y=2.685
+ $X2=0 $Y2=0
cc_108 N_A_80_153#_c_73_n N_A_324_508#_c_319_n 0.00974692f $X=1.225 $Y=2.43
+ $X2=0 $Y2=0
cc_109 N_A_80_153#_c_62_n N_VGND_c_340_n 0.00288714f $X=0.745 $Y=0.765 $X2=0
+ $Y2=0
cc_110 N_A_80_153#_c_65_n N_VGND_c_340_n 0.0088326f $X=1.285 $Y=0.945 $X2=0
+ $Y2=0
cc_111 N_A_80_153#_c_62_n N_VGND_c_342_n 0.00585385f $X=0.745 $Y=0.765 $X2=0
+ $Y2=0
cc_112 N_A_80_153#_c_63_n N_VGND_c_342_n 7.12021e-19 $X=0.745 $Y=0.84 $X2=0
+ $Y2=0
cc_113 N_A_80_153#_c_66_n N_VGND_c_344_n 0.00890272f $X=1.39 $Y=0.495 $X2=0
+ $Y2=0
cc_114 N_A_80_153#_M1001_d N_VGND_c_346_n 0.00378408f $X=1.25 $Y=0.235 $X2=0
+ $Y2=0
cc_115 N_A_80_153#_c_62_n N_VGND_c_346_n 0.00754763f $X=0.745 $Y=0.765 $X2=0
+ $Y2=0
cc_116 N_A_80_153#_c_63_n N_VGND_c_346_n 7.45101e-19 $X=0.745 $Y=0.84 $X2=0
+ $Y2=0
cc_117 N_A_80_153#_c_65_n N_VGND_c_346_n 0.0117102f $X=1.285 $Y=0.945 $X2=0
+ $Y2=0
cc_118 N_A_80_153#_c_104_p N_VGND_c_346_n 0.00216827f $X=0.695 $Y=0.945 $X2=0
+ $Y2=0
cc_119 N_A_80_153#_c_66_n N_VGND_c_346_n 0.00778069f $X=1.39 $Y=0.495 $X2=0
+ $Y2=0
cc_120 N_B1_M1001_g N_A1_M1006_g 0.0430198f $X=1.175 $Y=0.445 $X2=0 $Y2=0
cc_121 N_B1_c_136_n N_A1_M1002_g 0.00372299f $X=1.155 $Y=2.065 $X2=0 $Y2=0
cc_122 N_B1_c_141_n N_A1_M1002_g 0.0311308f $X=1.545 $Y=2.14 $X2=0 $Y2=0
cc_123 B1 N_A1_M1002_g 2.78042e-19 $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_124 N_B1_M1001_g A1 4.10536e-19 $X=1.175 $Y=0.445 $X2=0 $Y2=0
cc_125 N_B1_c_136_n A1 0.00203588f $X=1.155 $Y=2.065 $X2=0 $Y2=0
cc_126 N_B1_c_141_n A1 6.40048e-19 $X=1.545 $Y=2.14 $X2=0 $Y2=0
cc_127 B1 A1 0.0295221f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_128 N_B1_c_138_n A1 8.85865e-19 $X=1.155 $Y=1.615 $X2=0 $Y2=0
cc_129 N_B1_c_141_n N_A1_c_184_n 0.00666414f $X=1.545 $Y=2.14 $X2=0 $Y2=0
cc_130 B1 N_A1_c_184_n 0.00377067f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_131 N_B1_c_138_n N_A1_c_184_n 0.0249104f $X=1.155 $Y=1.615 $X2=0 $Y2=0
cc_132 N_B1_M1005_g N_VPWR_c_280_n 0.00525322f $X=1.545 $Y=2.75 $X2=0 $Y2=0
cc_133 N_B1_M1005_g N_VPWR_c_283_n 0.00461464f $X=1.545 $Y=2.75 $X2=0 $Y2=0
cc_134 N_B1_M1005_g N_VPWR_c_279_n 0.00914415f $X=1.545 $Y=2.75 $X2=0 $Y2=0
cc_135 N_B1_M1005_g N_A_324_508#_c_317_n 5.67832e-19 $X=1.545 $Y=2.75 $X2=0
+ $Y2=0
cc_136 N_B1_M1005_g N_A_324_508#_c_319_n 0.00264313f $X=1.545 $Y=2.75 $X2=0
+ $Y2=0
cc_137 N_B1_M1001_g N_VGND_c_340_n 0.00288714f $X=1.175 $Y=0.445 $X2=0 $Y2=0
cc_138 N_B1_M1001_g N_VGND_c_344_n 0.00585385f $X=1.175 $Y=0.445 $X2=0 $Y2=0
cc_139 N_B1_M1001_g N_VGND_c_346_n 0.0063829f $X=1.175 $Y=0.445 $X2=0 $Y2=0
cc_140 N_A1_M1006_g N_A2_c_227_n 0.0507187f $X=1.605 $Y=0.445 $X2=-0.19
+ $Y2=-0.245
cc_141 A1 N_A2_c_228_n 0.00998468f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_142 A1 N_A2_c_229_n 0.00699874f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_143 N_A1_c_184_n N_A2_c_229_n 0.00883959f $X=1.885 $Y=1.32 $X2=0 $Y2=0
cc_144 N_A1_M1002_g N_A2_c_231_n 0.0336748f $X=1.975 $Y=2.75 $X2=0 $Y2=0
cc_145 A1 A2 0.0714941f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_146 N_A1_c_184_n A2 2.08627e-19 $X=1.885 $Y=1.32 $X2=0 $Y2=0
cc_147 N_A1_M1006_g N_A2_c_233_n 0.00243334f $X=1.605 $Y=0.445 $X2=0 $Y2=0
cc_148 A1 N_A2_c_233_n 0.0126907f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_149 N_A1_c_184_n N_A2_c_233_n 0.0336748f $X=1.885 $Y=1.32 $X2=0 $Y2=0
cc_150 N_A1_M1002_g N_VPWR_c_281_n 0.00327258f $X=1.975 $Y=2.75 $X2=0 $Y2=0
cc_151 N_A1_M1002_g N_VPWR_c_283_n 0.00461464f $X=1.975 $Y=2.75 $X2=0 $Y2=0
cc_152 N_A1_M1002_g N_VPWR_c_279_n 0.00468324f $X=1.975 $Y=2.75 $X2=0 $Y2=0
cc_153 N_A1_M1002_g N_A_324_508#_c_317_n 9.4709e-19 $X=1.975 $Y=2.75 $X2=0 $Y2=0
cc_154 N_A1_M1002_g N_A_324_508#_c_318_n 0.0115629f $X=1.975 $Y=2.75 $X2=0 $Y2=0
cc_155 A1 N_A_324_508#_c_318_n 0.0294481f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_156 A1 N_A_324_508#_c_319_n 0.00566793f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_157 N_A1_c_184_n N_A_324_508#_c_319_n 0.0051995f $X=1.885 $Y=1.32 $X2=0 $Y2=0
cc_158 N_A1_M1006_g N_VGND_c_341_n 0.00204405f $X=1.605 $Y=0.445 $X2=0 $Y2=0
cc_159 A1 N_VGND_c_341_n 0.00831697f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_160 N_A1_M1006_g N_VGND_c_344_n 0.00585385f $X=1.605 $Y=0.445 $X2=0 $Y2=0
cc_161 N_A1_M1006_g N_VGND_c_346_n 0.0108402f $X=1.605 $Y=0.445 $X2=0 $Y2=0
cc_162 A1 N_VGND_c_346_n 0.00858622f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_163 N_A2_M1000_g N_VPWR_c_281_n 0.00327258f $X=2.405 $Y=2.75 $X2=0 $Y2=0
cc_164 N_A2_M1000_g N_VPWR_c_284_n 0.00461464f $X=2.405 $Y=2.75 $X2=0 $Y2=0
cc_165 N_A2_M1000_g N_VPWR_c_279_n 0.00471813f $X=2.405 $Y=2.75 $X2=0 $Y2=0
cc_166 N_A2_M1000_g N_A_324_508#_c_318_n 0.0177285f $X=2.405 $Y=2.75 $X2=0 $Y2=0
cc_167 A2 N_A_324_508#_c_318_n 0.017531f $X=2.555 $Y=0.47 $X2=0 $Y2=0
cc_168 N_A2_M1000_g N_A_324_508#_c_320_n 0.0020107f $X=2.405 $Y=2.75 $X2=0 $Y2=0
cc_169 N_A2_c_227_n N_VGND_c_341_n 0.0106247f $X=1.965 $Y=0.765 $X2=0 $Y2=0
cc_170 N_A2_c_228_n N_VGND_c_341_n 0.00733883f $X=2.33 $Y=0.84 $X2=0 $Y2=0
cc_171 A2 N_VGND_c_341_n 0.00115588f $X=2.555 $Y=0.47 $X2=0 $Y2=0
cc_172 N_A2_c_227_n N_VGND_c_344_n 0.00486043f $X=1.965 $Y=0.765 $X2=0 $Y2=0
cc_173 N_A2_c_228_n N_VGND_c_345_n 0.00511017f $X=2.33 $Y=0.84 $X2=0 $Y2=0
cc_174 A2 N_VGND_c_345_n 0.0059365f $X=2.555 $Y=0.47 $X2=0 $Y2=0
cc_175 N_A2_c_227_n N_VGND_c_346_n 0.00444929f $X=1.965 $Y=0.765 $X2=0 $Y2=0
cc_176 N_A2_c_228_n N_VGND_c_346_n 0.00619634f $X=2.33 $Y=0.84 $X2=0 $Y2=0
cc_177 A2 N_VGND_c_346_n 0.00676397f $X=2.555 $Y=0.47 $X2=0 $Y2=0
cc_178 X N_VPWR_c_282_n 0.00831216f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_179 N_X_M1004_s N_VPWR_c_279_n 0.00489501f $X=0.135 $Y=2.675 $X2=0 $Y2=0
cc_180 X N_VPWR_c_279_n 0.0069578f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_181 N_X_c_262_n N_VGND_c_342_n 0.0200121f $X=0.53 $Y=0.51 $X2=0 $Y2=0
cc_182 N_X_M1007_s N_VGND_c_346_n 0.00247251f $X=0.405 $Y=0.235 $X2=0 $Y2=0
cc_183 N_X_c_262_n N_VGND_c_346_n 0.0173604f $X=0.53 $Y=0.51 $X2=0 $Y2=0
cc_184 N_VPWR_c_283_n N_A_324_508#_c_317_n 0.00523228f $X=2.085 $Y=3.33 $X2=0
+ $Y2=0
cc_185 N_VPWR_c_279_n N_A_324_508#_c_317_n 0.00699584f $X=2.64 $Y=3.33 $X2=0
+ $Y2=0
cc_186 N_VPWR_c_281_n N_A_324_508#_c_318_n 0.0142847f $X=2.19 $Y=2.815 $X2=0
+ $Y2=0
cc_187 N_VPWR_c_279_n N_A_324_508#_c_318_n 0.0135041f $X=2.64 $Y=3.33 $X2=0
+ $Y2=0
cc_188 N_VPWR_c_284_n N_A_324_508#_c_320_n 0.00549876f $X=2.64 $Y=3.33 $X2=0
+ $Y2=0
cc_189 N_VPWR_c_279_n N_A_324_508#_c_320_n 0.00699584f $X=2.64 $Y=3.33 $X2=0
+ $Y2=0
cc_190 N_VGND_c_346_n A_336_47# 0.00648704f $X=2.64 $Y=0 $X2=-0.19 $Y2=-0.245
