* NGSPICE file created from sky130_fd_sc_lp__o41ai_m.ext - technology: sky130A

.subckt sky130_fd_sc_lp__o41ai_m A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
M1000 Y B1 VPWR VPB phighvt w=420000u l=150000u
+  ad=1.911e+11p pd=1.75e+06u as=2.226e+11p ps=2.74e+06u
M1001 a_463_371# A2 a_355_371# VPB phighvt w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=1.638e+11p ps=1.62e+06u
M1002 a_175_47# A1 VGND VNB nshort w=420000u l=150000u
+  ad=3.696e+11p pd=4.28e+06u as=2.835e+11p ps=3.03e+06u
M1003 VPWR A1 a_463_371# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VGND A4 a_175_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_247_371# A4 Y VPB phighvt w=420000u l=150000u
+  ad=1.638e+11p pd=1.62e+06u as=0p ps=0u
M1006 a_175_47# B1 Y VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=2.058e+11p ps=1.82e+06u
M1007 a_175_47# A3 VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_355_371# A3 a_247_371# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND A2 a_175_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

