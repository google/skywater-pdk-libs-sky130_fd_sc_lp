* File: sky130_fd_sc_lp__and3b_m.spice
* Created: Fri Aug 28 10:07:15 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__and3b_m.pex.spice"
.subckt sky130_fd_sc_lp__and3b_m  VNB VPB A_N B C VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* C	C
* B	B
* A_N	A_N
* VPB	VPB
* VNB	VNB
MM1006 N_A_110_53#_M1006_d N_A_N_M1006_g N_VGND_M1006_s VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.1113 PD=1.37 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1002 A_304_53# N_A_110_53#_M1002_g N_A_220_53#_M1002_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.1134 PD=0.63 PS=1.38 NRD=14.28 NRS=1.428 M=1 R=2.8
+ SA=75000.2 SB=75001.5 A=0.063 P=1.14 MULT=1
MM1003 A_376_53# N_B_M1003_g A_304_53# VNB NSHORT L=0.15 W=0.42 AD=0.0819
+ AS=0.0441 PD=0.81 PS=0.63 NRD=39.996 NRS=14.28 M=1 R=2.8 SA=75000.6 SB=75001.2
+ A=0.063 P=1.14 MULT=1
MM1005 N_VGND_M1005_d N_C_M1005_g A_376_53# VNB NSHORT L=0.15 W=0.42 AD=0.0588
+ AS=0.0819 PD=0.7 PS=0.81 NRD=0 NRS=39.996 M=1 R=2.8 SA=75001.1 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1009 N_X_M1009_d N_A_220_53#_M1009_g N_VGND_M1005_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.5 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1008 N_A_110_53#_M1008_d N_A_N_M1008_g N_VPWR_M1008_s VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1113 AS=0.1113 PD=1.37 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1004 N_VPWR_M1004_d N_A_110_53#_M1004_g N_A_220_53#_M1004_s VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.6 A=0.063 P=1.14 MULT=1
MM1000 N_A_220_53#_M1000_d N_B_M1000_g N_VPWR_M1004_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6 SB=75001.2
+ A=0.063 P=1.14 MULT=1
MM1007 N_VPWR_M1007_d N_C_M1007_g N_A_220_53#_M1000_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.09135 AS=0.0588 PD=0.855 PS=0.7 NRD=37.5088 NRS=0 M=1 R=2.8 SA=75001.1
+ SB=75000.8 A=0.063 P=1.14 MULT=1
MM1001 N_X_M1001_d N_A_220_53#_M1001_g N_VPWR_M1007_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.1113 AS=0.09135 PD=1.37 PS=0.855 NRD=0 NRS=35.1645 M=1 R=2.8 SA=75001.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9751 P=11.21
*
.include "sky130_fd_sc_lp__and3b_m.pxi.spice"
*
.ends
*
*
