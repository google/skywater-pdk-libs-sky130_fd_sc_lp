* File: sky130_fd_sc_lp__fa_m.spice
* Created: Wed Sep  2 09:53:36 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__fa_m.pex.spice"
.subckt sky130_fd_sc_lp__fa_m  VNB VPB B CIN A COUT VPWR SUM VGND
* 
* VGND	VGND
* SUM	SUM
* VPWR	VPWR
* COUT	COUT
* A	A
* CIN	CIN
* B	B
* VPB	VPB
* VNB	VNB
MM1021 N_VGND_M1021_d N_A_80_241#_M1021_g N_COUT_M1021_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.5 A=0.063 P=1.14 MULT=1
MM1013 A_227_125# N_A_M1013_g N_VGND_M1021_d VNB NSHORT L=0.15 W=0.42 AD=0.0441
+ AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.6 SB=75002.1
+ A=0.063 P=1.14 MULT=1
MM1007 N_A_80_241#_M1007_d N_B_M1007_g A_227_125# VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001
+ SB=75001.7 A=0.063 P=1.14 MULT=1
MM1008 N_A_385_125#_M1008_d N_CIN_M1008_g N_A_80_241#_M1007_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0756 AS=0.0588 PD=0.78 PS=0.7 NRD=22.848 NRS=0 M=1 R=2.8
+ SA=75001.4 SB=75001.3 A=0.063 P=1.14 MULT=1
MM1026 N_VGND_M1026_d N_A_M1026_g N_A_385_125#_M1008_d VNB NSHORT L=0.15 W=0.42
+ AD=0.09135 AS=0.0756 PD=0.855 PS=0.78 NRD=30 NRS=0 M=1 R=2.8 SA=75001.9
+ SB=75000.8 A=0.063 P=1.14 MULT=1
MM1009 N_A_385_125#_M1009_d N_B_M1009_g N_VGND_M1026_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.09135 PD=1.37 PS=0.855 NRD=0 NRS=14.28 M=1 R=2.8 SA=75002.5
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1023 N_A_843_119#_M1023_d N_B_M1023_g N_VGND_M1023_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75003.1
+ A=0.063 P=1.14 MULT=1
MM1017 N_VGND_M1017_d N_CIN_M1017_g N_A_843_119#_M1023_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75002.7 A=0.063 P=1.14 MULT=1
MM1018 N_A_843_119#_M1018_d N_A_M1018_g N_VGND_M1017_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.1 SB=75002.2
+ A=0.063 P=1.14 MULT=1
MM1027 N_A_1101_119#_M1027_d N_A_80_241#_M1027_g N_A_843_119#_M1018_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.0672 AS=0.0588 PD=0.74 PS=0.7 NRD=11.424 NRS=0 M=1 R=2.8
+ SA=75001.5 SB=75001.8 A=0.063 P=1.14 MULT=1
MM1000 A_1195_119# N_CIN_M1000_g N_A_1101_119#_M1027_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0672 PD=0.63 PS=0.74 NRD=14.28 NRS=0 M=1 R=2.8 SA=75001.9
+ SB=75001.3 A=0.063 P=1.14 MULT=1
MM1022 A_1267_119# N_B_M1022_g A_1195_119# VNB NSHORT L=0.15 W=0.42 AD=0.0441
+ AS=0.0441 PD=0.63 PS=0.63 NRD=14.28 NRS=14.28 M=1 R=2.8 SA=75002.3 SB=75001
+ A=0.063 P=1.14 MULT=1
MM1012 N_VGND_M1012_d N_A_M1012_g A_1267_119# VNB NSHORT L=0.15 W=0.42 AD=0.0588
+ AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75002.7 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1019 N_SUM_M1019_d N_A_1101_119#_M1019_g N_VGND_M1012_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75003.1
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1024 N_VPWR_M1024_d N_A_80_241#_M1024_g N_COUT_M1024_s VPB PHIGHVT L=0.15
+ W=0.42 AD=0.09135 AS=0.1113 PD=0.855 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.6 A=0.063 P=1.14 MULT=1
MM1002 A_227_367# N_A_M1002_g N_VPWR_M1024_d VPB PHIGHVT L=0.15 W=0.42 AD=0.0441
+ AS=0.09135 PD=0.63 PS=0.855 NRD=23.443 NRS=72.693 M=1 R=2.8 SA=75000.8
+ SB=75002 A=0.063 P=1.14 MULT=1
MM1005 N_A_80_241#_M1005_d N_B_M1005_g A_227_367# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=23.443 M=1 R=2.8 SA=75001.1
+ SB=75001.6 A=0.063 P=1.14 MULT=1
MM1025 N_A_385_367#_M1025_d N_CIN_M1025_g N_A_80_241#_M1005_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.6
+ SB=75001.2 A=0.063 P=1.14 MULT=1
MM1010 N_VPWR_M1010_d N_A_M1010_g N_A_385_367#_M1025_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.11975 AS=0.0588 PD=1.015 PS=0.7 NRD=72.693 NRS=0 M=1 R=2.8 SA=75002
+ SB=75000.8 A=0.063 P=1.14 MULT=1
MM1004 N_A_385_367#_M1004_d N_B_M1004_g N_VPWR_M1010_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.1113 AS=0.11975 PD=1.37 PS=1.015 NRD=0 NRS=39.8531 M=1 R=2.8 SA=75002.3
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1006 N_A_843_391#_M1006_d N_B_M1006_g N_VPWR_M1006_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75003.3
+ A=0.063 P=1.14 MULT=1
MM1014 N_VPWR_M1014_d N_CIN_M1014_g N_A_843_391#_M1006_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75002.8 A=0.063 P=1.14 MULT=1
MM1003 N_A_843_391#_M1003_d N_A_M1003_g N_VPWR_M1014_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.1 SB=75002.4
+ A=0.063 P=1.14 MULT=1
MM1016 N_A_1101_119#_M1016_d N_A_80_241#_M1016_g N_A_843_391#_M1003_d VPB
+ PHIGHVT L=0.15 W=0.42 AD=0.0672 AS=0.0588 PD=0.74 PS=0.7 NRD=18.7544 NRS=0 M=1
+ R=2.8 SA=75001.5 SB=75002 A=0.063 P=1.14 MULT=1
MM1011 A_1195_391# N_CIN_M1011_g N_A_1101_119#_M1016_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0441 AS=0.0672 PD=0.63 PS=0.74 NRD=23.443 NRS=0 M=1 R=2.8 SA=75001.9
+ SB=75001.5 A=0.063 P=1.14 MULT=1
MM1015 A_1267_391# N_B_M1015_g A_1195_391# VPB PHIGHVT L=0.15 W=0.42 AD=0.0441
+ AS=0.0441 PD=0.63 PS=0.63 NRD=23.443 NRS=23.443 M=1 R=2.8 SA=75002.3
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1020 N_VPWR_M1020_d N_A_M1020_g A_1267_391# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.09135 AS=0.0441 PD=0.855 PS=0.63 NRD=0 NRS=23.443 M=1 R=2.8 SA=75002.7
+ SB=75000.8 A=0.063 P=1.14 MULT=1
MM1001 N_SUM_M1001_d N_A_1101_119#_M1001_g N_VPWR_M1020_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1113 AS=0.09135 PD=1.37 PS=0.855 NRD=0 NRS=72.693 M=1 R=2.8
+ SA=75003.3 SB=75000.2 A=0.063 P=1.14 MULT=1
DX28_noxref VNB VPB NWDIODE A=15.1003 P=19.97
*
.include "sky130_fd_sc_lp__fa_m.pxi.spice"
*
.ends
*
*
