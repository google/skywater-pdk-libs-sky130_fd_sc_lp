* File: sky130_fd_sc_lp__a311oi_1.pxi.spice
* Created: Fri Aug 28 09:58:14 2020
* 
x_PM_SKY130_FD_SC_LP__A311OI_1%A3 N_A3_M1003_g N_A3_M1009_g A3 A3 N_A3_c_53_n
+ N_A3_c_54_n PM_SKY130_FD_SC_LP__A311OI_1%A3
x_PM_SKY130_FD_SC_LP__A311OI_1%A2 N_A2_M1008_g N_A2_M1000_g A2 N_A2_c_76_n
+ N_A2_c_77_n PM_SKY130_FD_SC_LP__A311OI_1%A2
x_PM_SKY130_FD_SC_LP__A311OI_1%A1 N_A1_c_108_n N_A1_M1007_g N_A1_M1001_g A1
+ N_A1_c_110_n N_A1_c_111_n PM_SKY130_FD_SC_LP__A311OI_1%A1
x_PM_SKY130_FD_SC_LP__A311OI_1%B1 N_B1_c_138_n N_B1_M1002_g N_B1_M1005_g B1
+ N_B1_c_140_n N_B1_c_141_n PM_SKY130_FD_SC_LP__A311OI_1%B1
x_PM_SKY130_FD_SC_LP__A311OI_1%C1 N_C1_c_170_n N_C1_M1004_g N_C1_M1006_g C1
+ N_C1_c_173_n PM_SKY130_FD_SC_LP__A311OI_1%C1
x_PM_SKY130_FD_SC_LP__A311OI_1%VPWR N_VPWR_M1009_s N_VPWR_M1000_d N_VPWR_c_197_n
+ N_VPWR_c_198_n N_VPWR_c_199_n N_VPWR_c_200_n VPWR N_VPWR_c_201_n
+ N_VPWR_c_202_n N_VPWR_c_196_n N_VPWR_c_204_n PM_SKY130_FD_SC_LP__A311OI_1%VPWR
x_PM_SKY130_FD_SC_LP__A311OI_1%A_181_367# N_A_181_367#_M1009_d
+ N_A_181_367#_M1001_d N_A_181_367#_c_239_n N_A_181_367#_c_236_n
+ N_A_181_367#_c_237_n N_A_181_367#_c_250_n
+ PM_SKY130_FD_SC_LP__A311OI_1%A_181_367#
x_PM_SKY130_FD_SC_LP__A311OI_1%Y N_Y_M1007_d N_Y_M1004_d N_Y_M1006_d N_Y_c_271_n
+ N_Y_c_275_n N_Y_c_276_n Y Y Y Y Y N_Y_c_277_n N_Y_c_290_n Y N_Y_c_273_n
+ PM_SKY130_FD_SC_LP__A311OI_1%Y
x_PM_SKY130_FD_SC_LP__A311OI_1%VGND N_VGND_M1003_s N_VGND_M1002_d N_VGND_c_328_n
+ N_VGND_c_329_n VGND N_VGND_c_330_n N_VGND_c_331_n N_VGND_c_332_n
+ N_VGND_c_333_n N_VGND_c_334_n N_VGND_c_335_n PM_SKY130_FD_SC_LP__A311OI_1%VGND
cc_1 VNB N_A3_M1009_g 0.0111375f $X=-0.19 $Y=-0.245 $X2=0.83 $Y2=2.465
cc_2 VNB A3 0.0469715f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_3 VNB N_A3_c_53_n 0.0354612f $X=-0.19 $Y=-0.245 $X2=0.74 $Y2=1.355
cc_4 VNB N_A3_c_54_n 0.0219466f $X=-0.19 $Y=-0.245 $X2=0.74 $Y2=1.19
cc_5 VNB N_A2_M1000_g 0.00839614f $X=-0.19 $Y=-0.245 $X2=0.83 $Y2=2.465
cc_6 VNB A2 0.00406629f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_7 VNB N_A2_c_76_n 0.0295459f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A2_c_77_n 0.0172093f $X=-0.19 $Y=-0.245 $X2=0.74 $Y2=1.355
cc_9 VNB N_A1_c_108_n 0.0182485f $X=-0.19 $Y=-0.245 $X2=0.83 $Y2=1.19
cc_10 VNB N_A1_M1001_g 0.008981f $X=-0.19 $Y=-0.245 $X2=0.83 $Y2=2.465
cc_11 VNB N_A1_c_110_n 0.00491115f $X=-0.19 $Y=-0.245 $X2=0.74 $Y2=1.355
cc_12 VNB N_A1_c_111_n 0.0325675f $X=-0.19 $Y=-0.245 $X2=0.74 $Y2=1.19
cc_13 VNB N_B1_c_138_n 0.0190798f $X=-0.19 $Y=-0.245 $X2=0.83 $Y2=1.19
cc_14 VNB N_B1_M1005_g 0.00786958f $X=-0.19 $Y=-0.245 $X2=0.83 $Y2=2.465
cc_15 VNB N_B1_c_140_n 0.0046968f $X=-0.19 $Y=-0.245 $X2=0.74 $Y2=1.355
cc_16 VNB N_B1_c_141_n 0.034597f $X=-0.19 $Y=-0.245 $X2=0.74 $Y2=1.19
cc_17 VNB N_C1_c_170_n 0.0229316f $X=-0.19 $Y=-0.245 $X2=0.83 $Y2=1.19
cc_18 VNB N_C1_M1006_g 0.0101754f $X=-0.19 $Y=-0.245 $X2=0.83 $Y2=2.465
cc_19 VNB C1 0.00469037f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_20 VNB N_C1_c_173_n 0.0509468f $X=-0.19 $Y=-0.245 $X2=0.74 $Y2=1.355
cc_21 VNB N_VPWR_c_196_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_Y_c_271_n 0.00428887f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB Y 0.00851864f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_Y_c_273_n 0.0230339f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_328_n 0.0333434f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_26 VNB N_VGND_c_329_n 0.00561756f $X=-0.19 $Y=-0.245 $X2=0.74 $Y2=1.355
cc_27 VNB N_VGND_c_330_n 0.0164632f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.355
cc_28 VNB N_VGND_c_331_n 0.039478f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_332_n 0.0181824f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_333_n 0.202657f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_334_n 0.00513431f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_335_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VPB N_A3_M1009_g 0.0271235f $X=-0.19 $Y=1.655 $X2=0.83 $Y2=2.465
cc_34 VPB N_A2_M1000_g 0.021327f $X=-0.19 $Y=1.655 $X2=0.83 $Y2=2.465
cc_35 VPB N_A1_M1001_g 0.0226445f $X=-0.19 $Y=1.655 $X2=0.83 $Y2=2.465
cc_36 VPB N_B1_M1005_g 0.0211255f $X=-0.19 $Y=1.655 $X2=0.83 $Y2=2.465
cc_37 VPB N_C1_M1006_g 0.0237058f $X=-0.19 $Y=1.655 $X2=0.83 $Y2=2.465
cc_38 VPB N_VPWR_c_197_n 0.05508f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_39 VPB N_VPWR_c_198_n 0.00564356f $X=-0.19 $Y=1.655 $X2=0.74 $Y2=1.19
cc_40 VPB N_VPWR_c_199_n 0.0164632f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=1.355
cc_41 VPB N_VPWR_c_200_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_42 VPB N_VPWR_c_201_n 0.0177387f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_43 VPB N_VPWR_c_202_n 0.0462617f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_44 VPB N_VPWR_c_196_n 0.058938f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_45 VPB N_VPWR_c_204_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_46 VPB N_A_181_367#_c_236_n 0.011045f $X=-0.19 $Y=1.655 $X2=0.74 $Y2=1.355
cc_47 VPB N_A_181_367#_c_237_n 0.00680871f $X=-0.19 $Y=1.655 $X2=0.74 $Y2=1.355
cc_48 VPB N_Y_c_271_n 8.75531e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_49 VPB N_Y_c_275_n 0.0117131f $X=-0.19 $Y=1.655 $X2=0.74 $Y2=1.355
cc_50 VPB N_Y_c_276_n 0.0462319f $X=-0.19 $Y=1.655 $X2=0.74 $Y2=1.355
cc_51 N_A3_M1009_g N_A2_M1000_g 0.024397f $X=0.83 $Y=2.465 $X2=0 $Y2=0
cc_52 A3 A2 0.0275639f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_53 N_A3_c_54_n A2 0.00200674f $X=0.74 $Y=1.19 $X2=0 $Y2=0
cc_54 A3 N_A2_c_76_n 3.54112e-19 $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_55 N_A3_c_53_n N_A2_c_76_n 0.0205934f $X=0.74 $Y=1.355 $X2=0 $Y2=0
cc_56 N_A3_c_54_n N_A2_c_77_n 0.0440308f $X=0.74 $Y=1.19 $X2=0 $Y2=0
cc_57 N_A3_M1009_g N_VPWR_c_197_n 0.023736f $X=0.83 $Y=2.465 $X2=0 $Y2=0
cc_58 A3 N_VPWR_c_197_n 0.0187744f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_59 N_A3_c_53_n N_VPWR_c_197_n 0.00390317f $X=0.74 $Y=1.355 $X2=0 $Y2=0
cc_60 N_A3_M1009_g N_VPWR_c_201_n 0.00486043f $X=0.83 $Y=2.465 $X2=0 $Y2=0
cc_61 N_A3_M1009_g N_VPWR_c_196_n 0.00833196f $X=0.83 $Y=2.465 $X2=0 $Y2=0
cc_62 N_A3_M1009_g N_A_181_367#_c_237_n 0.00421401f $X=0.83 $Y=2.465 $X2=0 $Y2=0
cc_63 N_A3_c_54_n N_Y_c_277_n 0.0064984f $X=0.74 $Y=1.19 $X2=0 $Y2=0
cc_64 A3 N_VGND_c_328_n 0.0249987f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_65 N_A3_c_53_n N_VGND_c_328_n 0.00401953f $X=0.74 $Y=1.355 $X2=0 $Y2=0
cc_66 N_A3_c_54_n N_VGND_c_328_n 0.0189915f $X=0.74 $Y=1.19 $X2=0 $Y2=0
cc_67 N_A3_c_54_n N_VGND_c_331_n 0.00486043f $X=0.74 $Y=1.19 $X2=0 $Y2=0
cc_68 N_A3_c_54_n N_VGND_c_333_n 0.00842105f $X=0.74 $Y=1.19 $X2=0 $Y2=0
cc_69 N_A2_c_77_n N_A1_c_108_n 0.0457139f $X=1.28 $Y=1.19 $X2=-0.19 $Y2=-0.245
cc_70 N_A2_M1000_g N_A1_M1001_g 0.0309823f $X=1.285 $Y=2.465 $X2=0 $Y2=0
cc_71 A2 N_A1_c_110_n 0.0267228f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_72 N_A2_c_76_n N_A1_c_110_n 0.00215024f $X=1.28 $Y=1.355 $X2=0 $Y2=0
cc_73 A2 N_A1_c_111_n 2.9608e-19 $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_74 N_A2_c_76_n N_A1_c_111_n 0.0204667f $X=1.28 $Y=1.355 $X2=0 $Y2=0
cc_75 N_A2_M1000_g N_VPWR_c_197_n 0.00146708f $X=1.285 $Y=2.465 $X2=0 $Y2=0
cc_76 N_A2_M1000_g N_VPWR_c_198_n 0.0139526f $X=1.285 $Y=2.465 $X2=0 $Y2=0
cc_77 N_A2_M1000_g N_VPWR_c_201_n 0.0054895f $X=1.285 $Y=2.465 $X2=0 $Y2=0
cc_78 N_A2_M1000_g N_VPWR_c_196_n 0.0106157f $X=1.285 $Y=2.465 $X2=0 $Y2=0
cc_79 N_A2_M1000_g N_A_181_367#_c_239_n 0.0176367f $X=1.285 $Y=2.465 $X2=0 $Y2=0
cc_80 N_A2_M1000_g N_A_181_367#_c_236_n 0.0121117f $X=1.285 $Y=2.465 $X2=0 $Y2=0
cc_81 A2 N_A_181_367#_c_236_n 0.0100321f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_82 N_A2_c_76_n N_A_181_367#_c_236_n 0.00225326f $X=1.28 $Y=1.355 $X2=0 $Y2=0
cc_83 N_A2_M1000_g N_A_181_367#_c_237_n 0.00224409f $X=1.285 $Y=2.465 $X2=0
+ $Y2=0
cc_84 A2 N_A_181_367#_c_237_n 0.0148883f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_85 N_A2_c_76_n N_A_181_367#_c_237_n 0.00225253f $X=1.28 $Y=1.355 $X2=0 $Y2=0
cc_86 A2 N_Y_c_277_n 0.0225243f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_87 N_A2_c_76_n N_Y_c_277_n 0.00227547f $X=1.28 $Y=1.355 $X2=0 $Y2=0
cc_88 N_A2_c_77_n N_Y_c_277_n 0.0298304f $X=1.28 $Y=1.19 $X2=0 $Y2=0
cc_89 N_A2_c_77_n N_VGND_c_328_n 0.00178646f $X=1.28 $Y=1.19 $X2=0 $Y2=0
cc_90 N_A2_c_77_n N_VGND_c_331_n 0.00357877f $X=1.28 $Y=1.19 $X2=0 $Y2=0
cc_91 N_A2_c_77_n N_VGND_c_333_n 0.00557914f $X=1.28 $Y=1.19 $X2=0 $Y2=0
cc_92 N_A1_c_108_n N_B1_c_138_n 0.020843f $X=1.73 $Y=1.19 $X2=-0.19 $Y2=-0.245
cc_93 N_A1_c_111_n N_B1_M1005_g 0.0350821f $X=1.94 $Y=1.355 $X2=0 $Y2=0
cc_94 N_A1_c_110_n N_B1_c_140_n 0.0267973f $X=1.82 $Y=1.355 $X2=0 $Y2=0
cc_95 N_A1_c_111_n N_B1_c_140_n 0.00235219f $X=1.94 $Y=1.355 $X2=0 $Y2=0
cc_96 N_A1_c_110_n N_B1_c_141_n 2.56571e-19 $X=1.82 $Y=1.355 $X2=0 $Y2=0
cc_97 N_A1_c_111_n N_B1_c_141_n 0.0202195f $X=1.94 $Y=1.355 $X2=0 $Y2=0
cc_98 N_A1_M1001_g N_VPWR_c_198_n 0.0156311f $X=1.94 $Y=2.465 $X2=0 $Y2=0
cc_99 N_A1_M1001_g N_VPWR_c_202_n 0.00585385f $X=1.94 $Y=2.465 $X2=0 $Y2=0
cc_100 N_A1_M1001_g N_VPWR_c_196_n 0.0118061f $X=1.94 $Y=2.465 $X2=0 $Y2=0
cc_101 N_A1_M1001_g N_A_181_367#_c_239_n 9.6303e-19 $X=1.94 $Y=2.465 $X2=0 $Y2=0
cc_102 N_A1_M1001_g N_A_181_367#_c_236_n 0.0178523f $X=1.94 $Y=2.465 $X2=0 $Y2=0
cc_103 N_A1_c_110_n N_A_181_367#_c_236_n 0.0273929f $X=1.82 $Y=1.355 $X2=0 $Y2=0
cc_104 N_A1_c_111_n N_A_181_367#_c_236_n 0.0052993f $X=1.94 $Y=1.355 $X2=0 $Y2=0
cc_105 N_A1_M1001_g N_A_181_367#_c_250_n 0.0165359f $X=1.94 $Y=2.465 $X2=0 $Y2=0
cc_106 N_A1_c_111_n Y 0.00432747f $X=1.94 $Y=1.355 $X2=0 $Y2=0
cc_107 N_A1_c_108_n N_Y_c_277_n 0.0356487f $X=1.73 $Y=1.19 $X2=0 $Y2=0
cc_108 N_A1_c_110_n N_Y_c_277_n 0.024849f $X=1.82 $Y=1.355 $X2=0 $Y2=0
cc_109 N_A1_c_108_n N_VGND_c_331_n 0.00357877f $X=1.73 $Y=1.19 $X2=0 $Y2=0
cc_110 N_A1_c_108_n N_VGND_c_333_n 0.00586375f $X=1.73 $Y=1.19 $X2=0 $Y2=0
cc_111 N_B1_c_138_n N_C1_c_170_n 0.023955f $X=2.3 $Y=1.185 $X2=-0.19 $Y2=-0.245
cc_112 N_B1_M1005_g N_C1_M1006_g 0.0605135f $X=2.525 $Y=2.465 $X2=0 $Y2=0
cc_113 N_B1_c_140_n N_C1_c_173_n 2.48192e-19 $X=2.39 $Y=1.35 $X2=0 $Y2=0
cc_114 N_B1_c_141_n N_C1_c_173_n 0.0605135f $X=2.525 $Y=1.35 $X2=0 $Y2=0
cc_115 N_B1_M1005_g N_VPWR_c_202_n 0.00585385f $X=2.525 $Y=2.465 $X2=0 $Y2=0
cc_116 N_B1_M1005_g N_VPWR_c_196_n 0.0111935f $X=2.525 $Y=2.465 $X2=0 $Y2=0
cc_117 N_B1_M1005_g N_A_181_367#_c_236_n 0.00186079f $X=2.525 $Y=2.465 $X2=0
+ $Y2=0
cc_118 N_B1_c_140_n N_A_181_367#_c_236_n 0.0278508f $X=2.39 $Y=1.35 $X2=0 $Y2=0
cc_119 N_B1_c_141_n N_A_181_367#_c_236_n 0.0047714f $X=2.525 $Y=1.35 $X2=0 $Y2=0
cc_120 N_B1_c_138_n N_Y_c_271_n 0.00333524f $X=2.3 $Y=1.185 $X2=0 $Y2=0
cc_121 N_B1_c_140_n N_Y_c_271_n 0.0251371f $X=2.39 $Y=1.35 $X2=0 $Y2=0
cc_122 N_B1_c_141_n N_Y_c_271_n 0.00648031f $X=2.525 $Y=1.35 $X2=0 $Y2=0
cc_123 N_B1_M1005_g N_Y_c_275_n 0.00122356f $X=2.525 $Y=2.465 $X2=0 $Y2=0
cc_124 N_B1_c_138_n Y 0.00960032f $X=2.3 $Y=1.185 $X2=0 $Y2=0
cc_125 N_B1_c_140_n Y 0.0265379f $X=2.39 $Y=1.35 $X2=0 $Y2=0
cc_126 N_B1_c_138_n N_Y_c_290_n 0.00977985f $X=2.3 $Y=1.185 $X2=0 $Y2=0
cc_127 N_B1_c_141_n N_Y_c_290_n 0.00741896f $X=2.525 $Y=1.35 $X2=0 $Y2=0
cc_128 N_B1_c_138_n N_Y_c_273_n 8.53709e-19 $X=2.3 $Y=1.185 $X2=0 $Y2=0
cc_129 N_B1_c_138_n N_VGND_c_329_n 0.00583946f $X=2.3 $Y=1.185 $X2=0 $Y2=0
cc_130 N_B1_c_138_n N_VGND_c_331_n 0.0055505f $X=2.3 $Y=1.185 $X2=0 $Y2=0
cc_131 N_B1_c_138_n N_VGND_c_333_n 0.00698258f $X=2.3 $Y=1.185 $X2=0 $Y2=0
cc_132 N_C1_M1006_g N_VPWR_c_202_n 0.00585385f $X=2.885 $Y=2.465 $X2=0 $Y2=0
cc_133 N_C1_M1006_g N_VPWR_c_196_n 0.0116377f $X=2.885 $Y=2.465 $X2=0 $Y2=0
cc_134 N_C1_c_170_n N_Y_c_271_n 0.00837922f $X=2.885 $Y=1.185 $X2=0 $Y2=0
cc_135 N_C1_M1006_g N_Y_c_271_n 0.00845104f $X=2.885 $Y=2.465 $X2=0 $Y2=0
cc_136 C1 N_Y_c_271_n 0.0230504f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_137 N_C1_c_173_n N_Y_c_271_n 0.00660618f $X=3.07 $Y=1.35 $X2=0 $Y2=0
cc_138 N_C1_M1006_g N_Y_c_275_n 0.0188364f $X=2.885 $Y=2.465 $X2=0 $Y2=0
cc_139 C1 N_Y_c_275_n 0.0172186f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_140 N_C1_c_173_n N_Y_c_275_n 0.00266267f $X=3.07 $Y=1.35 $X2=0 $Y2=0
cc_141 N_C1_c_170_n Y 8.38887e-19 $X=2.885 $Y=1.185 $X2=0 $Y2=0
cc_142 N_C1_c_170_n Y 0.0147726f $X=2.885 $Y=1.185 $X2=0 $Y2=0
cc_143 C1 Y 0.0173199f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_144 N_C1_c_173_n Y 0.00168381f $X=3.07 $Y=1.35 $X2=0 $Y2=0
cc_145 N_C1_c_170_n N_Y_c_273_n 0.0111986f $X=2.885 $Y=1.185 $X2=0 $Y2=0
cc_146 N_C1_c_170_n N_VGND_c_329_n 0.00578173f $X=2.885 $Y=1.185 $X2=0 $Y2=0
cc_147 N_C1_c_170_n N_VGND_c_332_n 0.0054895f $X=2.885 $Y=1.185 $X2=0 $Y2=0
cc_148 N_C1_c_170_n N_VGND_c_333_n 0.00747785f $X=2.885 $Y=1.185 $X2=0 $Y2=0
cc_149 N_VPWR_c_196_n N_A_181_367#_M1009_d 0.00400207f $X=3.12 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_150 N_VPWR_c_196_n N_A_181_367#_M1001_d 0.00724561f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_151 N_VPWR_c_198_n N_A_181_367#_c_239_n 0.064709f $X=1.625 $Y=2.115 $X2=0
+ $Y2=0
cc_152 N_VPWR_c_201_n N_A_181_367#_c_239_n 0.0174459f $X=1.46 $Y=3.33 $X2=0
+ $Y2=0
cc_153 N_VPWR_c_196_n N_A_181_367#_c_239_n 0.0108194f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_154 N_VPWR_M1000_d N_A_181_367#_c_236_n 0.00608312f $X=1.36 $Y=1.835 $X2=0
+ $Y2=0
cc_155 N_VPWR_c_198_n N_A_181_367#_c_236_n 0.0266856f $X=1.625 $Y=2.115 $X2=0
+ $Y2=0
cc_156 N_VPWR_c_197_n N_A_181_367#_c_237_n 0.0025823f $X=0.615 $Y=1.98 $X2=0
+ $Y2=0
cc_157 N_VPWR_c_198_n N_A_181_367#_c_250_n 0.0572855f $X=1.625 $Y=2.115 $X2=0
+ $Y2=0
cc_158 N_VPWR_c_202_n N_A_181_367#_c_250_n 0.0226794f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_159 N_VPWR_c_196_n N_A_181_367#_c_250_n 0.0127519f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_160 N_VPWR_c_196_n A_520_367# 0.00899413f $X=3.12 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_161 N_VPWR_c_196_n N_Y_M1006_d 0.00249946f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_162 N_VPWR_c_202_n N_Y_c_276_n 0.0190529f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_163 N_VPWR_c_196_n N_Y_c_276_n 0.0113912f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_164 N_A_181_367#_c_236_n N_Y_c_271_n 9.93198e-19 $X=2.075 $Y=1.775 $X2=0
+ $Y2=0
cc_165 N_A_181_367#_c_236_n N_Y_c_275_n 0.00932535f $X=2.075 $Y=1.775 $X2=0
+ $Y2=0
cc_166 N_A_181_367#_c_236_n N_Y_c_277_n 0.0092948f $X=2.075 $Y=1.775 $X2=0 $Y2=0
cc_167 N_A_181_367#_c_237_n N_Y_c_277_n 8.39264e-19 $X=1.235 $Y=1.775 $X2=0
+ $Y2=0
cc_168 A_520_367# N_Y_c_275_n 0.00366293f $X=2.6 $Y=1.835 $X2=0.615 $Y2=2.95
cc_169 N_Y_c_271_n N_VGND_M1002_d 0.00106811f $X=2.73 $Y=1.705 $X2=0 $Y2=0
cc_170 Y N_VGND_M1002_d 0.0014499f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_171 N_Y_c_290_n N_VGND_M1002_d 0.00640984f $X=2.645 $Y=0.927 $X2=0 $Y2=0
cc_172 N_Y_c_277_n N_VGND_c_328_n 0.0458265f $X=1.865 $Y=0.635 $X2=0 $Y2=0
cc_173 N_Y_c_290_n N_VGND_c_329_n 0.0255576f $X=2.645 $Y=0.927 $X2=0 $Y2=0
cc_174 N_Y_c_277_n N_VGND_c_331_n 0.0738892f $X=1.865 $Y=0.635 $X2=0 $Y2=0
cc_175 N_Y_c_273_n N_VGND_c_332_n 0.0208381f $X=3.1 $Y=0.38 $X2=0 $Y2=0
cc_176 N_Y_M1007_d N_VGND_c_333_n 0.00339796f $X=1.805 $Y=0.235 $X2=0 $Y2=0
cc_177 N_Y_M1004_d N_VGND_c_333_n 0.00215158f $X=2.96 $Y=0.235 $X2=0 $Y2=0
cc_178 Y N_VGND_c_333_n 0.00540037f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_179 N_Y_c_277_n N_VGND_c_333_n 0.0455389f $X=1.865 $Y=0.635 $X2=0 $Y2=0
cc_180 N_Y_c_290_n N_VGND_c_333_n 0.00634013f $X=2.645 $Y=0.927 $X2=0 $Y2=0
cc_181 N_Y_c_273_n N_VGND_c_333_n 0.0125193f $X=3.1 $Y=0.38 $X2=0 $Y2=0
cc_182 N_Y_c_277_n A_181_47# 0.0101476f $X=1.865 $Y=0.635 $X2=-0.19 $Y2=-0.245
cc_183 N_Y_c_277_n A_270_47# 0.00528158f $X=1.865 $Y=0.635 $X2=-0.19 $Y2=-0.245
cc_184 N_VGND_c_333_n A_181_47# 0.00689478f $X=3.12 $Y=0 $X2=-0.19 $Y2=-0.245
cc_185 N_VGND_c_333_n A_270_47# 0.00245291f $X=3.12 $Y=0 $X2=-0.19 $Y2=-0.245
