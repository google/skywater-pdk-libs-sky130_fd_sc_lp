* File: sky130_fd_sc_lp__nand4_m.pex.spice
* Created: Fri Aug 28 10:51:21 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__NAND4_M%D 3 7 12 13 14 15 16 17 23
r33 23 24 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.63
+ $Y=1.32 $X2=0.63 $Y2=1.32
r34 16 17 7.90266 $w=5.58e-07 $l=3.7e-07 $layer=LI1_cond $X=0.435 $Y=1.665
+ $X2=0.435 $Y2=2.035
r35 16 24 7.3687 $w=5.58e-07 $l=3.45e-07 $layer=LI1_cond $X=0.435 $Y=1.665
+ $X2=0.435 $Y2=1.32
r36 15 24 0.533964 $w=5.58e-07 $l=2.5e-08 $layer=LI1_cond $X=0.435 $Y=1.295
+ $X2=0.435 $Y2=1.32
r37 14 15 7.90266 $w=5.58e-07 $l=3.7e-07 $layer=LI1_cond $X=0.435 $Y=0.925
+ $X2=0.435 $Y2=1.295
r38 12 23 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=0.63 $Y=1.675
+ $X2=0.63 $Y2=1.32
r39 12 13 43.5886 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=0.7 $Y=1.675 $X2=0.7
+ $Y2=1.825
r40 10 23 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.63 $Y=1.155
+ $X2=0.63 $Y2=1.32
r41 7 13 356.372 $w=1.5e-07 $l=6.95e-07 $layer=POLY_cond $X=0.86 $Y=2.52
+ $X2=0.86 $Y2=1.825
r42 3 10 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=0.72 $Y=0.445
+ $X2=0.72 $Y2=1.155
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4_M%C 3 6 9 10 11 12 13 14 15 21
c47 11 0 1.22132e-19 $X=1.2 $Y=1.435
r48 14 15 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=1.2 $Y=1.295 $X2=1.2
+ $Y2=1.665
r49 13 14 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=1.2 $Y=0.925 $X2=1.2
+ $Y2=1.295
r50 13 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.2 $Y=0.93
+ $X2=1.2 $Y2=0.93
r51 12 13 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=1.2 $Y=0.555 $X2=1.2
+ $Y2=0.925
r52 10 21 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.2 $Y=1.27 $X2=1.2
+ $Y2=0.93
r53 10 11 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.2 $Y=1.27 $X2=1.2
+ $Y2=1.435
r54 9 21 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.2 $Y=0.765 $X2=1.2
+ $Y2=0.93
r55 6 11 556.351 $w=1.5e-07 $l=1.085e-06 $layer=POLY_cond $X=1.29 $Y=2.52
+ $X2=1.29 $Y2=1.435
r56 3 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.11 $Y=0.445 $X2=1.11
+ $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4_M%B 3 6 9 10 11 12 13 14 15 21
r49 21 22 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.77
+ $Y=0.93 $X2=1.77 $Y2=0.93
r50 14 15 16.4002 $w=2.58e-07 $l=3.7e-07 $layer=LI1_cond $X=1.725 $Y=1.295
+ $X2=1.725 $Y2=1.665
r51 14 22 16.1785 $w=2.58e-07 $l=3.65e-07 $layer=LI1_cond $X=1.725 $Y=1.295
+ $X2=1.725 $Y2=0.93
r52 13 22 0.221624 $w=2.58e-07 $l=5e-09 $layer=LI1_cond $X=1.725 $Y=0.925
+ $X2=1.725 $Y2=0.93
r53 12 13 16.4002 $w=2.58e-07 $l=3.7e-07 $layer=LI1_cond $X=1.725 $Y=0.555
+ $X2=1.725 $Y2=0.925
r54 10 21 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.77 $Y=1.27
+ $X2=1.77 $Y2=0.93
r55 10 11 40.8701 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.77 $Y=1.27
+ $X2=1.77 $Y2=1.435
r56 9 21 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.77 $Y=0.765
+ $X2=1.77 $Y2=0.93
r57 6 11 556.351 $w=1.5e-07 $l=1.085e-06 $layer=POLY_cond $X=1.72 $Y=2.52
+ $X2=1.72 $Y2=1.435
r58 3 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.68 $Y=0.445 $X2=1.68
+ $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4_M%A 3 7 10 13 17 18 19 20 21 26
c43 7 0 1.03456e-19 $X=2.25 $Y=0.445
r44 26 27 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.34
+ $Y=1.005 $X2=2.34 $Y2=1.005
r45 20 21 12.183 $w=3.48e-07 $l=3.7e-07 $layer=LI1_cond $X=2.25 $Y=1.295
+ $X2=2.25 $Y2=1.665
r46 20 27 9.54881 $w=3.48e-07 $l=2.9e-07 $layer=LI1_cond $X=2.25 $Y=1.295
+ $X2=2.25 $Y2=1.005
r47 19 27 2.63416 $w=3.48e-07 $l=8e-08 $layer=LI1_cond $X=2.25 $Y=0.925 $X2=2.25
+ $Y2=1.005
r48 17 26 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.34 $Y=1.345
+ $X2=2.34 $Y2=1.005
r49 17 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.34 $Y=1.345
+ $X2=2.34 $Y2=1.51
r50 16 26 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.34 $Y=0.84
+ $X2=2.34 $Y2=1.005
r51 11 13 51.2766 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=2.15 $Y=1.75 $X2=2.25
+ $Y2=1.75
r52 10 13 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.25 $Y=1.675
+ $X2=2.25 $Y2=1.75
r53 10 18 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.25 $Y=1.675
+ $X2=2.25 $Y2=1.51
r54 7 16 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=2.25 $Y=0.445
+ $X2=2.25 $Y2=0.84
r55 1 11 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.15 $Y=1.825
+ $X2=2.15 $Y2=1.75
r56 1 3 356.372 $w=1.5e-07 $l=6.95e-07 $layer=POLY_cond $X=2.15 $Y=1.825
+ $X2=2.15 $Y2=2.52
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4_M%VPWR 1 2 3 12 16 18 20 23 24 26 27 28 37 43
r34 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r35 40 43 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r36 39 40 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r37 37 42 3.61693 $w=1.7e-07 $l=2.27e-07 $layer=LI1_cond $X=2.425 $Y=3.33
+ $X2=2.652 $Y2=3.33
r38 37 39 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=2.425 $Y=3.33
+ $X2=2.16 $Y2=3.33
r39 35 36 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r40 32 36 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.2 $Y2=3.33
r41 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r42 28 40 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=2.16 $Y2=3.33
r43 28 36 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=1.2 $Y2=3.33
r44 26 35 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=1.4 $Y=3.33 $X2=1.2
+ $Y2=3.33
r45 26 27 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.4 $Y=3.33
+ $X2=1.505 $Y2=3.33
r46 25 39 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=1.61 $Y=3.33
+ $X2=2.16 $Y2=3.33
r47 25 27 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.61 $Y=3.33
+ $X2=1.505 $Y2=3.33
r48 23 31 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=0.54 $Y=3.33 $X2=0.24
+ $Y2=3.33
r49 23 24 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=0.54 $Y=3.33
+ $X2=0.645 $Y2=3.33
r50 22 35 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=0.75 $Y=3.33 $X2=1.2
+ $Y2=3.33
r51 22 24 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=0.75 $Y=3.33
+ $X2=0.645 $Y2=3.33
r52 18 42 3.29826 $w=2.1e-07 $l=1.58915e-07 $layer=LI1_cond $X=2.53 $Y=3.245
+ $X2=2.652 $Y2=3.33
r53 18 20 38.026 $w=2.08e-07 $l=7.2e-07 $layer=LI1_cond $X=2.53 $Y=3.245
+ $X2=2.53 $Y2=2.525
r54 14 27 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=1.505 $Y=3.245
+ $X2=1.505 $Y2=3.33
r55 14 16 38.026 $w=2.08e-07 $l=7.2e-07 $layer=LI1_cond $X=1.505 $Y=3.245
+ $X2=1.505 $Y2=2.525
r56 10 24 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=0.645 $Y=3.245
+ $X2=0.645 $Y2=3.33
r57 10 12 38.026 $w=2.08e-07 $l=7.2e-07 $layer=LI1_cond $X=0.645 $Y=3.245
+ $X2=0.645 $Y2=2.525
r58 3 20 600 $w=1.7e-07 $l=3.98246e-07 $layer=licon1_PDIFF $count=1 $X=2.225
+ $Y=2.31 $X2=2.53 $Y2=2.525
r59 2 16 600 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_PDIFF $count=1 $X=1.365
+ $Y=2.31 $X2=1.505 $Y2=2.525
r60 1 12 600 $w=1.7e-07 $l=2.7037e-07 $layer=licon1_PDIFF $count=1 $X=0.52
+ $Y=2.31 $X2=0.645 $Y2=2.525
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4_M%Y 1 2 3 11 15 17 18 19 20 28 31 37 42
c52 28 0 1.22132e-19 $X=1.83 $Y=2.035
c53 15 0 1.03456e-19 $X=2.69 $Y=0.495
r54 29 31 1.30481 $w=1.68e-07 $l=2e-08 $layer=LI1_cond $X=1.18 $Y=2.035 $X2=1.2
+ $Y2=2.035
r55 20 28 10.0494 $w=1.7e-07 $l=2.07e-07 $layer=LI1_cond $X=2.037 $Y=2.035
+ $X2=1.83 $Y2=2.035
r56 20 42 9.10246 $w=5.83e-07 $l=3.95e-07 $layer=LI1_cond $X=2.037 $Y=2.12
+ $X2=2.037 $Y2=2.515
r57 19 28 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=1.68 $Y=2.035
+ $X2=1.83 $Y2=2.035
r58 18 29 3.82155 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.075 $Y=2.035
+ $X2=1.18 $Y2=2.035
r59 18 37 17.2256 $w=2.73e-07 $l=3.95e-07 $layer=LI1_cond $X=1.075 $Y=2.12
+ $X2=1.075 $Y2=2.515
r60 18 19 29.2278 $w=1.68e-07 $l=4.48e-07 $layer=LI1_cond $X=1.232 $Y=2.035
+ $X2=1.68 $Y2=2.035
r61 18 31 2.0877 $w=1.68e-07 $l=3.2e-08 $layer=LI1_cond $X=1.232 $Y=2.035
+ $X2=1.2 $Y2=2.035
r62 17 20 13.6419 $w=3.38e-07 $l=3.6e-07 $layer=LI1_cond $X=2.605 $Y=2.035
+ $X2=2.245 $Y2=2.035
r63 13 15 7.15912 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=2.485 $Y=0.495
+ $X2=2.69 $Y2=0.495
r64 11 17 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.69 $Y=1.95
+ $X2=2.605 $Y2=2.035
r65 10 15 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.69 $Y=0.66
+ $X2=2.69 $Y2=0.495
r66 10 11 84.1604 $w=1.68e-07 $l=1.29e-06 $layer=LI1_cond $X=2.69 $Y=0.66
+ $X2=2.69 $Y2=1.95
r67 3 42 600 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=1 $X=1.795
+ $Y=2.31 $X2=1.935 $Y2=2.515
r68 2 37 600 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=1 $X=0.935
+ $Y=2.31 $X2=1.075 $Y2=2.515
r69 1 13 182 $w=1.7e-07 $l=3.30454e-07 $layer=licon1_NDIFF $count=1 $X=2.325
+ $Y=0.235 $X2=2.485 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4_M%VGND 1 6 9 10 11 21 22
r34 21 22 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r35 18 21 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=0.72 $Y=0 $X2=2.64
+ $Y2=0
r36 18 19 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r37 15 19 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r38 14 15 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r39 11 22 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=1.44 $Y=0 $X2=2.64
+ $Y2=0
r40 11 19 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=0.72
+ $Y2=0
r41 9 14 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=0.34 $Y=0 $X2=0.24
+ $Y2=0
r42 9 10 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.34 $Y=0 $X2=0.505
+ $Y2=0
r43 8 18 3.26203 $w=1.68e-07 $l=5e-08 $layer=LI1_cond $X=0.67 $Y=0 $X2=0.72
+ $Y2=0
r44 8 10 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.67 $Y=0 $X2=0.505
+ $Y2=0
r45 4 10 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.505 $Y=0.085
+ $X2=0.505 $Y2=0
r46 4 6 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.505 $Y=0.085
+ $X2=0.505 $Y2=0.38
r47 1 6 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.38
+ $Y=0.235 $X2=0.505 $Y2=0.38
.ends

