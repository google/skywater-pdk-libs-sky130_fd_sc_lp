* File: sky130_fd_sc_lp__a311o_0.pxi.spice
* Created: Fri Aug 28 09:57:20 2020
* 
x_PM_SKY130_FD_SC_LP__A311O_0%A_72_312# N_A_72_312#_M1001_d N_A_72_312#_M1003_d
+ N_A_72_312#_M1000_d N_A_72_312#_M1006_g N_A_72_312#_M1004_g N_A_72_312#_c_96_n
+ N_A_72_312#_c_97_n N_A_72_312#_c_86_n N_A_72_312#_c_87_n N_A_72_312#_c_99_n
+ N_A_72_312#_c_100_n N_A_72_312#_c_88_n N_A_72_312#_c_89_n N_A_72_312#_c_90_n
+ N_A_72_312#_c_91_n N_A_72_312#_c_92_n N_A_72_312#_c_93_n N_A_72_312#_c_94_n
+ N_A_72_312#_c_102_n N_A_72_312#_c_103_n N_A_72_312#_c_104_n
+ PM_SKY130_FD_SC_LP__A311O_0%A_72_312#
x_PM_SKY130_FD_SC_LP__A311O_0%A3 N_A3_M1008_g N_A3_M1011_g N_A3_c_194_n
+ N_A3_c_195_n N_A3_c_196_n A3 A3 A3 N_A3_c_198_n PM_SKY130_FD_SC_LP__A311O_0%A3
x_PM_SKY130_FD_SC_LP__A311O_0%A2 N_A2_c_234_n N_A2_M1005_g N_A2_M1009_g
+ N_A2_c_236_n A2 A2 A2 A2 N_A2_c_238_n N_A2_c_239_n
+ PM_SKY130_FD_SC_LP__A311O_0%A2
x_PM_SKY130_FD_SC_LP__A311O_0%A1 N_A1_M1001_g N_A1_M1007_g N_A1_c_281_n
+ N_A1_c_282_n A1 A1 A1 A1 N_A1_c_284_n PM_SKY130_FD_SC_LP__A311O_0%A1
x_PM_SKY130_FD_SC_LP__A311O_0%B1 N_B1_M1002_g N_B1_M1010_g N_B1_c_328_n
+ N_B1_c_329_n B1 B1 N_B1_c_330_n N_B1_c_331_n PM_SKY130_FD_SC_LP__A311O_0%B1
x_PM_SKY130_FD_SC_LP__A311O_0%C1 N_C1_M1000_g N_C1_M1003_g N_C1_c_377_n
+ N_C1_c_378_n C1 C1 C1 N_C1_c_375_n PM_SKY130_FD_SC_LP__A311O_0%C1
x_PM_SKY130_FD_SC_LP__A311O_0%X N_X_M1006_s N_X_M1004_s N_X_c_416_n N_X_c_413_n
+ X X X N_X_c_415_n PM_SKY130_FD_SC_LP__A311O_0%X
x_PM_SKY130_FD_SC_LP__A311O_0%VPWR N_VPWR_M1004_d N_VPWR_M1005_d N_VPWR_c_441_n
+ N_VPWR_c_442_n N_VPWR_c_443_n N_VPWR_c_444_n VPWR N_VPWR_c_445_n
+ N_VPWR_c_440_n N_VPWR_c_447_n PM_SKY130_FD_SC_LP__A311O_0%VPWR
x_PM_SKY130_FD_SC_LP__A311O_0%A_224_486# N_A_224_486#_M1008_d
+ N_A_224_486#_M1007_d N_A_224_486#_c_482_n N_A_224_486#_c_483_n
+ N_A_224_486#_c_484_n N_A_224_486#_c_488_n
+ PM_SKY130_FD_SC_LP__A311O_0%A_224_486#
x_PM_SKY130_FD_SC_LP__A311O_0%VGND N_VGND_M1006_d N_VGND_M1010_d N_VGND_c_511_n
+ N_VGND_c_512_n N_VGND_c_513_n N_VGND_c_514_n VGND N_VGND_c_515_n
+ N_VGND_c_516_n N_VGND_c_517_n N_VGND_c_518_n PM_SKY130_FD_SC_LP__A311O_0%VGND
cc_1 VNB N_A_72_312#_M1006_g 0.0699527f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=0.45
cc_2 VNB N_A_72_312#_c_86_n 0.00102128f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.725
cc_3 VNB N_A_72_312#_c_87_n 0.0123496f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.725
cc_4 VNB N_A_72_312#_c_88_n 0.00147406f $X=-0.19 $Y=-0.245 $X2=2.595 $Y2=0.45
cc_5 VNB N_A_72_312#_c_89_n 0.00451211f $X=-0.19 $Y=-0.245 $X2=3 $Y2=0.825
cc_6 VNB N_A_72_312#_c_90_n 0.00354932f $X=-0.19 $Y=-0.245 $X2=2.725 $Y2=0.825
cc_7 VNB N_A_72_312#_c_91_n 0.00494788f $X=-0.19 $Y=-0.245 $X2=3.1 $Y2=2.035
cc_8 VNB N_A_72_312#_c_92_n 0.0106785f $X=-0.19 $Y=-0.245 $X2=3.375 $Y2=0.825
cc_9 VNB N_A_72_312#_c_93_n 0.0183697f $X=-0.19 $Y=-0.245 $X2=3.48 $Y2=0.45
cc_10 VNB N_A_72_312#_c_94_n 0.00165317f $X=-0.19 $Y=-0.245 $X2=3.1 $Y2=0.825
cc_11 VNB N_A3_M1008_g 0.0106863f $X=-0.19 $Y=-0.245 $X2=3.15 $Y2=2.43
cc_12 VNB N_A3_c_194_n 0.0175038f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A3_c_195_n 0.0209097f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=1.56
cc_14 VNB N_A3_c_196_n 0.0158044f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=0.45
cc_15 VNB A3 0.00888846f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=0.45
cc_16 VNB N_A3_c_198_n 0.0151095f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.56
cc_17 VNB N_A2_c_234_n 0.0204428f $X=-0.19 $Y=-0.245 $X2=3.34 $Y2=0.24
cc_18 VNB N_A2_M1005_g 0.0117991f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A2_c_236_n 0.017941f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=1.56
cc_20 VNB A2 0.00622804f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=0.45
cc_21 VNB N_A2_c_238_n 0.0184657f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=2.065
cc_22 VNB N_A2_c_239_n 0.0168667f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=2.035
cc_23 VNB N_A1_M1001_g 0.0336295f $X=-0.19 $Y=-0.245 $X2=3.15 $Y2=2.43
cc_24 VNB N_A1_c_281_n 0.022407f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=0.45
cc_25 VNB N_A1_c_282_n 0.00493621f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=0.45
cc_26 VNB A1 0.0104257f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A1_c_284_n 0.0177193f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=2.035
cc_28 VNB N_B1_M1010_g 0.0359256f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_B1_c_328_n 0.0216166f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=0.45
cc_30 VNB N_B1_c_329_n 0.00440602f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=0.45
cc_31 VNB N_B1_c_330_n 0.0157747f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.725
cc_32 VNB N_B1_c_331_n 0.00679839f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.56
cc_33 VNB N_C1_M1003_g 0.0601096f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB C1 0.0339548f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_C1_c_375_n 0.0258537f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=2.065
cc_36 VNB N_X_c_413_n 0.0128368f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=0.45
cc_37 VNB X 0.0173041f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=2.75
cc_38 VNB N_X_c_415_n 0.0427377f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=2.23
cc_39 VNB N_VPWR_c_440_n 0.163682f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.725
cc_40 VNB N_VGND_c_511_n 0.00576562f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_512_n 6.17563e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_513_n 0.0212916f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=2.75
cc_43 VNB N_VGND_c_514_n 0.00632182f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_515_n 0.0500149f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.725
cc_45 VNB N_VGND_c_516_n 0.0183369f $X=-0.19 $Y=-0.245 $X2=3 $Y2=0.825
cc_46 VNB N_VGND_c_517_n 0.213833f $X=-0.19 $Y=-0.245 $X2=2.725 $Y2=0.825
cc_47 VNB N_VGND_c_518_n 0.00415849f $X=-0.19 $Y=-0.245 $X2=3.11 $Y2=2.23
cc_48 VPB N_A_72_312#_M1004_g 0.0263637f $X=-0.19 $Y=1.655 $X2=0.615 $Y2=2.75
cc_49 VPB N_A_72_312#_c_96_n 0.0261608f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=2.065
cc_50 VPB N_A_72_312#_c_97_n 0.0168024f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=2.23
cc_51 VPB N_A_72_312#_c_87_n 0.00544883f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=1.725
cc_52 VPB N_A_72_312#_c_99_n 0.0559901f $X=-0.19 $Y=1.655 $X2=3 $Y2=2.132
cc_53 VPB N_A_72_312#_c_100_n 0.00104146f $X=-0.19 $Y=1.655 $X2=0.69 $Y2=2.132
cc_54 VPB N_A_72_312#_c_91_n 0.00252205f $X=-0.19 $Y=1.655 $X2=3.1 $Y2=2.035
cc_55 VPB N_A_72_312#_c_102_n 0.00115851f $X=-0.19 $Y=1.655 $X2=3.1 $Y2=2.132
cc_56 VPB N_A_72_312#_c_103_n 0.0323084f $X=-0.19 $Y=1.655 $X2=3.29 $Y2=2.575
cc_57 VPB N_A_72_312#_c_104_n 0.0054662f $X=-0.19 $Y=1.655 $X2=3.237 $Y2=2.39
cc_58 VPB N_A3_M1008_g 0.0508152f $X=-0.19 $Y=1.655 $X2=3.15 $Y2=2.43
cc_59 VPB A3 0.00393855f $X=-0.19 $Y=1.655 $X2=0.615 $Y2=0.45
cc_60 VPB N_A2_M1005_g 0.0588136f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_61 VPB A2 0.00407091f $X=-0.19 $Y=1.655 $X2=0.615 $Y2=0.45
cc_62 VPB N_A1_M1007_g 0.0523661f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_63 VPB N_A1_c_282_n 0.0118314f $X=-0.19 $Y=1.655 $X2=0.615 $Y2=0.45
cc_64 VPB A1 0.00341207f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_65 VPB N_B1_M1002_g 0.0429126f $X=-0.19 $Y=1.655 $X2=3.15 $Y2=2.43
cc_66 VPB N_B1_c_329_n 0.0110942f $X=-0.19 $Y=1.655 $X2=0.615 $Y2=0.45
cc_67 VPB N_B1_c_331_n 0.00404871f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=1.56
cc_68 VPB N_C1_M1000_g 0.0299631f $X=-0.19 $Y=1.655 $X2=3.15 $Y2=2.43
cc_69 VPB N_C1_c_377_n 0.0266007f $X=-0.19 $Y=1.655 $X2=0.615 $Y2=0.45
cc_70 VPB N_C1_c_378_n 0.0334744f $X=-0.19 $Y=1.655 $X2=0.615 $Y2=0.45
cc_71 VPB C1 0.0349525f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_72 VPB N_C1_c_375_n 0.00450168f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=2.065
cc_73 VPB N_X_c_416_n 0.0390468f $X=-0.19 $Y=1.655 $X2=0.615 $Y2=1.56
cc_74 VPB N_X_c_413_n 0.0356129f $X=-0.19 $Y=1.655 $X2=0.615 $Y2=0.45
cc_75 VPB N_VPWR_c_441_n 0.00767633f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_76 VPB N_VPWR_c_442_n 0.0174259f $X=-0.19 $Y=1.655 $X2=0.615 $Y2=0.45
cc_77 VPB N_VPWR_c_443_n 0.0209111f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_78 VPB N_VPWR_c_444_n 0.00439477f $X=-0.19 $Y=1.655 $X2=0.615 $Y2=2.23
cc_79 VPB N_VPWR_c_445_n 0.0478554f $X=-0.19 $Y=1.655 $X2=0.56 $Y2=1.725
cc_80 VPB N_VPWR_c_440_n 0.0777675f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=1.725
cc_81 VPB N_VPWR_c_447_n 0.0172789f $X=-0.19 $Y=1.655 $X2=3 $Y2=2.132
cc_82 VPB N_A_224_486#_c_482_n 0.00223416f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_83 VPB N_A_224_486#_c_483_n 0.00822909f $X=-0.19 $Y=1.655 $X2=0.615 $Y2=0.45
cc_84 VPB N_A_224_486#_c_484_n 0.00316877f $X=-0.19 $Y=1.655 $X2=0.615 $Y2=0.45
cc_85 N_A_72_312#_M1006_g N_A3_M1008_g 0.0506443f $X=0.615 $Y=0.45 $X2=0 $Y2=0
cc_86 N_A_72_312#_c_86_n N_A3_M1008_g 0.00210994f $X=0.525 $Y=1.725 $X2=0 $Y2=0
cc_87 N_A_72_312#_c_99_n N_A3_M1008_g 0.0166602f $X=3 $Y=2.132 $X2=0 $Y2=0
cc_88 N_A_72_312#_M1006_g N_A3_c_194_n 0.0134526f $X=0.615 $Y=0.45 $X2=0 $Y2=0
cc_89 N_A_72_312#_c_99_n N_A3_c_196_n 0.0022036f $X=3 $Y=2.132 $X2=0 $Y2=0
cc_90 N_A_72_312#_M1006_g A3 0.00395818f $X=0.615 $Y=0.45 $X2=0 $Y2=0
cc_91 N_A_72_312#_c_86_n A3 0.0145779f $X=0.525 $Y=1.725 $X2=0 $Y2=0
cc_92 N_A_72_312#_c_99_n A3 0.0308211f $X=3 $Y=2.132 $X2=0 $Y2=0
cc_93 N_A_72_312#_M1006_g N_A3_c_198_n 0.0402207f $X=0.615 $Y=0.45 $X2=0 $Y2=0
cc_94 N_A_72_312#_c_99_n N_A2_M1005_g 0.0161417f $X=3 $Y=2.132 $X2=0 $Y2=0
cc_95 N_A_72_312#_c_99_n N_A2_c_236_n 6.19858e-19 $X=3 $Y=2.132 $X2=0 $Y2=0
cc_96 N_A_72_312#_c_99_n A2 0.0245292f $X=3 $Y=2.132 $X2=0 $Y2=0
cc_97 N_A_72_312#_c_88_n N_A1_M1001_g 0.00303499f $X=2.595 $Y=0.45 $X2=0 $Y2=0
cc_98 N_A_72_312#_c_90_n N_A1_M1001_g 6.55135e-19 $X=2.725 $Y=0.825 $X2=0 $Y2=0
cc_99 N_A_72_312#_c_99_n N_A1_M1007_g 0.0151028f $X=3 $Y=2.132 $X2=0 $Y2=0
cc_100 N_A_72_312#_c_99_n N_A1_c_282_n 0.00126102f $X=3 $Y=2.132 $X2=0 $Y2=0
cc_101 N_A_72_312#_M1001_d A1 0.00340609f $X=2.19 $Y=0.24 $X2=0 $Y2=0
cc_102 N_A_72_312#_c_99_n A1 0.0238929f $X=3 $Y=2.132 $X2=0 $Y2=0
cc_103 N_A_72_312#_c_88_n A1 0.0266745f $X=2.595 $Y=0.45 $X2=0 $Y2=0
cc_104 N_A_72_312#_c_90_n A1 0.0137713f $X=2.725 $Y=0.825 $X2=0 $Y2=0
cc_105 N_A_72_312#_c_99_n N_B1_M1002_g 0.0147264f $X=3 $Y=2.132 $X2=0 $Y2=0
cc_106 N_A_72_312#_c_91_n N_B1_M1002_g 0.00329697f $X=3.1 $Y=2.035 $X2=0 $Y2=0
cc_107 N_A_72_312#_c_104_n N_B1_M1002_g 0.0034246f $X=3.237 $Y=2.39 $X2=0 $Y2=0
cc_108 N_A_72_312#_c_88_n N_B1_M1010_g 0.00151093f $X=2.595 $Y=0.45 $X2=0 $Y2=0
cc_109 N_A_72_312#_c_89_n N_B1_M1010_g 0.0150585f $X=3 $Y=0.825 $X2=0 $Y2=0
cc_110 N_A_72_312#_c_91_n N_B1_M1010_g 0.00874057f $X=3.1 $Y=2.035 $X2=0 $Y2=0
cc_111 N_A_72_312#_c_99_n N_B1_c_329_n 0.00353282f $X=3 $Y=2.132 $X2=0 $Y2=0
cc_112 N_A_72_312#_c_89_n N_B1_c_330_n 2.41254e-19 $X=3 $Y=0.825 $X2=0 $Y2=0
cc_113 N_A_72_312#_c_90_n N_B1_c_330_n 0.0011206f $X=2.725 $Y=0.825 $X2=0 $Y2=0
cc_114 N_A_72_312#_c_99_n N_B1_c_331_n 0.0301207f $X=3 $Y=2.132 $X2=0 $Y2=0
cc_115 N_A_72_312#_c_89_n N_B1_c_331_n 0.00801536f $X=3 $Y=0.825 $X2=0 $Y2=0
cc_116 N_A_72_312#_c_90_n N_B1_c_331_n 0.0221537f $X=2.725 $Y=0.825 $X2=0 $Y2=0
cc_117 N_A_72_312#_c_91_n N_B1_c_331_n 0.0606557f $X=3.1 $Y=2.035 $X2=0 $Y2=0
cc_118 N_A_72_312#_c_102_n N_C1_M1000_g 0.00443004f $X=3.1 $Y=2.132 $X2=0 $Y2=0
cc_119 N_A_72_312#_c_103_n N_C1_M1000_g 0.0164275f $X=3.29 $Y=2.575 $X2=0 $Y2=0
cc_120 N_A_72_312#_c_104_n N_C1_M1000_g 0.00625193f $X=3.237 $Y=2.39 $X2=0 $Y2=0
cc_121 N_A_72_312#_c_91_n N_C1_M1003_g 0.015161f $X=3.1 $Y=2.035 $X2=0 $Y2=0
cc_122 N_A_72_312#_c_92_n N_C1_M1003_g 0.0150743f $X=3.375 $Y=0.825 $X2=0 $Y2=0
cc_123 N_A_72_312#_c_93_n N_C1_M1003_g 0.00263805f $X=3.48 $Y=0.45 $X2=0 $Y2=0
cc_124 N_A_72_312#_c_94_n N_C1_M1003_g 0.00228713f $X=3.1 $Y=0.825 $X2=0 $Y2=0
cc_125 N_A_72_312#_c_91_n N_C1_c_377_n 0.00766925f $X=3.1 $Y=2.035 $X2=0 $Y2=0
cc_126 N_A_72_312#_c_91_n N_C1_c_378_n 0.00571315f $X=3.1 $Y=2.035 $X2=0 $Y2=0
cc_127 N_A_72_312#_c_102_n N_C1_c_378_n 0.00571597f $X=3.1 $Y=2.132 $X2=0 $Y2=0
cc_128 N_A_72_312#_c_103_n N_C1_c_378_n 0.0080654f $X=3.29 $Y=2.575 $X2=0 $Y2=0
cc_129 N_A_72_312#_c_91_n C1 0.0712833f $X=3.1 $Y=2.035 $X2=0 $Y2=0
cc_130 N_A_72_312#_c_92_n C1 0.0251401f $X=3.375 $Y=0.825 $X2=0 $Y2=0
cc_131 N_A_72_312#_c_102_n C1 0.0156309f $X=3.1 $Y=2.132 $X2=0 $Y2=0
cc_132 N_A_72_312#_c_103_n C1 0.00778028f $X=3.29 $Y=2.575 $X2=0 $Y2=0
cc_133 N_A_72_312#_c_91_n N_C1_c_375_n 0.00683643f $X=3.1 $Y=2.035 $X2=0 $Y2=0
cc_134 N_A_72_312#_c_92_n N_C1_c_375_n 0.00169782f $X=3.375 $Y=0.825 $X2=0 $Y2=0
cc_135 N_A_72_312#_M1004_g N_X_c_416_n 0.00769015f $X=0.615 $Y=2.75 $X2=0 $Y2=0
cc_136 N_A_72_312#_c_97_n N_X_c_416_n 0.00414205f $X=0.525 $Y=2.23 $X2=0 $Y2=0
cc_137 N_A_72_312#_c_100_n N_X_c_416_n 0.0112975f $X=0.69 $Y=2.132 $X2=0 $Y2=0
cc_138 N_A_72_312#_M1006_g N_X_c_413_n 0.00364948f $X=0.615 $Y=0.45 $X2=0 $Y2=0
cc_139 N_A_72_312#_M1004_g N_X_c_413_n 0.00395485f $X=0.615 $Y=2.75 $X2=0 $Y2=0
cc_140 N_A_72_312#_c_86_n N_X_c_413_n 0.0350635f $X=0.525 $Y=1.725 $X2=0 $Y2=0
cc_141 N_A_72_312#_c_87_n N_X_c_413_n 0.0162824f $X=0.525 $Y=1.725 $X2=0 $Y2=0
cc_142 N_A_72_312#_c_100_n N_X_c_413_n 0.0155727f $X=0.69 $Y=2.132 $X2=0 $Y2=0
cc_143 N_A_72_312#_M1006_g X 0.00929683f $X=0.615 $Y=0.45 $X2=0 $Y2=0
cc_144 N_A_72_312#_c_86_n X 0.0117368f $X=0.525 $Y=1.725 $X2=0 $Y2=0
cc_145 N_A_72_312#_c_87_n X 0.00426075f $X=0.525 $Y=1.725 $X2=0 $Y2=0
cc_146 N_A_72_312#_M1006_g N_X_c_415_n 0.023887f $X=0.615 $Y=0.45 $X2=0 $Y2=0
cc_147 N_A_72_312#_M1004_g N_VPWR_c_441_n 0.00289192f $X=0.615 $Y=2.75 $X2=0
+ $Y2=0
cc_148 N_A_72_312#_c_99_n N_VPWR_c_441_n 0.0186665f $X=3 $Y=2.132 $X2=0 $Y2=0
cc_149 N_A_72_312#_M1004_g N_VPWR_c_443_n 0.00525141f $X=0.615 $Y=2.75 $X2=0
+ $Y2=0
cc_150 N_A_72_312#_c_103_n N_VPWR_c_445_n 0.0305971f $X=3.29 $Y=2.575 $X2=0
+ $Y2=0
cc_151 N_A_72_312#_M1004_g N_VPWR_c_440_n 0.0106115f $X=0.615 $Y=2.75 $X2=0
+ $Y2=0
cc_152 N_A_72_312#_c_103_n N_VPWR_c_440_n 0.0162457f $X=3.29 $Y=2.575 $X2=0
+ $Y2=0
cc_153 N_A_72_312#_c_99_n N_A_224_486#_c_483_n 0.0917454f $X=3 $Y=2.132 $X2=0
+ $Y2=0
cc_154 N_A_72_312#_c_103_n N_A_224_486#_c_483_n 0.00764979f $X=3.29 $Y=2.575
+ $X2=0 $Y2=0
cc_155 N_A_72_312#_c_99_n N_A_224_486#_c_484_n 0.0279092f $X=3 $Y=2.132 $X2=0
+ $Y2=0
cc_156 N_A_72_312#_c_103_n N_A_224_486#_c_488_n 0.019063f $X=3.29 $Y=2.575 $X2=0
+ $Y2=0
cc_157 N_A_72_312#_M1006_g N_VGND_c_511_n 0.00513243f $X=0.615 $Y=0.45 $X2=0
+ $Y2=0
cc_158 N_A_72_312#_c_89_n N_VGND_c_512_n 0.00558637f $X=3 $Y=0.825 $X2=0 $Y2=0
cc_159 N_A_72_312#_c_94_n N_VGND_c_512_n 0.0150119f $X=3.1 $Y=0.825 $X2=0 $Y2=0
cc_160 N_A_72_312#_M1006_g N_VGND_c_513_n 0.00545083f $X=0.615 $Y=0.45 $X2=0
+ $Y2=0
cc_161 N_A_72_312#_c_88_n N_VGND_c_515_n 0.0136323f $X=2.595 $Y=0.45 $X2=0 $Y2=0
cc_162 N_A_72_312#_c_89_n N_VGND_c_515_n 0.0022495f $X=3 $Y=0.825 $X2=0 $Y2=0
cc_163 N_A_72_312#_c_92_n N_VGND_c_516_n 0.0022495f $X=3.375 $Y=0.825 $X2=0
+ $Y2=0
cc_164 N_A_72_312#_c_93_n N_VGND_c_516_n 0.0151469f $X=3.48 $Y=0.45 $X2=0 $Y2=0
cc_165 N_A_72_312#_M1001_d N_VGND_c_517_n 0.0115275f $X=2.19 $Y=0.24 $X2=0 $Y2=0
cc_166 N_A_72_312#_M1003_d N_VGND_c_517_n 0.0023277f $X=3.34 $Y=0.24 $X2=0 $Y2=0
cc_167 N_A_72_312#_M1006_g N_VGND_c_517_n 0.0112487f $X=0.615 $Y=0.45 $X2=0
+ $Y2=0
cc_168 N_A_72_312#_c_88_n N_VGND_c_517_n 0.00928586f $X=2.595 $Y=0.45 $X2=0
+ $Y2=0
cc_169 N_A_72_312#_c_89_n N_VGND_c_517_n 0.00421113f $X=3 $Y=0.825 $X2=0 $Y2=0
cc_170 N_A_72_312#_c_92_n N_VGND_c_517_n 0.0038286f $X=3.375 $Y=0.825 $X2=0
+ $Y2=0
cc_171 N_A_72_312#_c_93_n N_VGND_c_517_n 0.0102412f $X=3.48 $Y=0.45 $X2=0 $Y2=0
cc_172 N_A_72_312#_c_94_n N_VGND_c_517_n 8.45664e-19 $X=3.1 $Y=0.825 $X2=0 $Y2=0
cc_173 N_A3_c_195_n N_A2_c_234_n 0.0138518f $X=1.065 $Y=1.275 $X2=0 $Y2=0
cc_174 N_A3_M1008_g N_A2_M1005_g 0.0434026f $X=1.045 $Y=2.75 $X2=0 $Y2=0
cc_175 N_A3_c_196_n N_A2_c_236_n 0.0138518f $X=1.065 $Y=1.44 $X2=0 $Y2=0
cc_176 N_A3_M1008_g A2 3.50201e-19 $X=1.045 $Y=2.75 $X2=0 $Y2=0
cc_177 N_A3_c_194_n A2 0.00178322f $X=1.065 $Y=0.77 $X2=0 $Y2=0
cc_178 A3 A2 0.0865138f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_179 N_A3_c_198_n A2 5.57284e-19 $X=1.065 $Y=0.935 $X2=0 $Y2=0
cc_180 A3 N_A2_c_238_n 0.00795045f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_181 N_A3_c_198_n N_A2_c_238_n 0.0138518f $X=1.065 $Y=0.935 $X2=0 $Y2=0
cc_182 N_A3_c_194_n N_A2_c_239_n 0.030481f $X=1.065 $Y=0.77 $X2=0 $Y2=0
cc_183 N_A3_c_195_n X 9.31673e-19 $X=1.065 $Y=1.275 $X2=0 $Y2=0
cc_184 N_A3_c_194_n N_X_c_415_n 7.76119e-19 $X=1.065 $Y=0.77 $X2=0 $Y2=0
cc_185 A3 N_X_c_415_n 0.0235187f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_186 N_A3_c_198_n N_X_c_415_n 9.31673e-19 $X=1.065 $Y=0.935 $X2=0 $Y2=0
cc_187 N_A3_M1008_g N_VPWR_c_441_n 0.00184008f $X=1.045 $Y=2.75 $X2=0 $Y2=0
cc_188 N_A3_M1008_g N_VPWR_c_442_n 0.00560159f $X=1.045 $Y=2.75 $X2=0 $Y2=0
cc_189 N_A3_M1008_g N_VPWR_c_440_n 0.0105762f $X=1.045 $Y=2.75 $X2=0 $Y2=0
cc_190 N_A3_M1008_g N_A_224_486#_c_484_n 5.21028e-19 $X=1.045 $Y=2.75 $X2=0
+ $Y2=0
cc_191 N_A3_c_194_n N_VGND_c_511_n 0.00326685f $X=1.065 $Y=0.77 $X2=0 $Y2=0
cc_192 A3 N_VGND_c_511_n 0.00518778f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_193 N_A3_c_198_n N_VGND_c_511_n 0.00439289f $X=1.065 $Y=0.935 $X2=0 $Y2=0
cc_194 N_A3_c_194_n N_VGND_c_515_n 0.0058025f $X=1.065 $Y=0.77 $X2=0 $Y2=0
cc_195 N_A3_c_194_n N_VGND_c_517_n 0.006294f $X=1.065 $Y=0.77 $X2=0 $Y2=0
cc_196 A3 N_VGND_c_517_n 0.011579f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_197 A2 N_A1_M1001_g 0.00448597f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_198 N_A2_c_238_n N_A1_M1001_g 0.0122301f $X=1.635 $Y=0.935 $X2=0 $Y2=0
cc_199 N_A2_c_239_n N_A1_M1001_g 0.0208403f $X=1.62 $Y=0.77 $X2=0 $Y2=0
cc_200 N_A2_M1005_g N_A1_M1007_g 0.0200914f $X=1.515 $Y=2.75 $X2=0 $Y2=0
cc_201 A2 N_A1_M1007_g 3.02763e-19 $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_202 N_A2_M1005_g N_A1_c_281_n 0.00713419f $X=1.515 $Y=2.75 $X2=0 $Y2=0
cc_203 N_A2_c_236_n N_A1_c_281_n 0.0122301f $X=1.62 $Y=1.44 $X2=0 $Y2=0
cc_204 N_A2_M1005_g A1 9.85136e-19 $X=1.515 $Y=2.75 $X2=0 $Y2=0
cc_205 A2 A1 0.109895f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_206 N_A2_c_238_n A1 0.00205984f $X=1.635 $Y=0.935 $X2=0 $Y2=0
cc_207 N_A2_c_239_n A1 4.75512e-19 $X=1.62 $Y=0.77 $X2=0 $Y2=0
cc_208 N_A2_c_234_n N_A1_c_284_n 0.0122301f $X=1.62 $Y=1.26 $X2=0 $Y2=0
cc_209 N_A2_M1005_g N_VPWR_c_442_n 0.00409234f $X=1.515 $Y=2.75 $X2=0 $Y2=0
cc_210 N_A2_M1005_g N_VPWR_c_440_n 0.00642206f $X=1.515 $Y=2.75 $X2=0 $Y2=0
cc_211 N_A2_M1005_g N_VPWR_c_447_n 0.0020956f $X=1.515 $Y=2.75 $X2=0 $Y2=0
cc_212 N_A2_M1005_g N_A_224_486#_c_482_n 0.0110851f $X=1.515 $Y=2.75 $X2=0 $Y2=0
cc_213 N_A2_M1005_g N_A_224_486#_c_483_n 0.0101847f $X=1.515 $Y=2.75 $X2=0 $Y2=0
cc_214 N_A2_M1005_g N_A_224_486#_c_484_n 0.00106507f $X=1.515 $Y=2.75 $X2=0
+ $Y2=0
cc_215 A2 N_VGND_c_515_n 0.0104893f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_216 N_A2_c_238_n N_VGND_c_515_n 0.00154767f $X=1.635 $Y=0.935 $X2=0 $Y2=0
cc_217 N_A2_c_239_n N_VGND_c_515_n 0.00425722f $X=1.62 $Y=0.77 $X2=0 $Y2=0
cc_218 A2 N_VGND_c_517_n 0.0101356f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_219 N_A2_c_238_n N_VGND_c_517_n 0.00159874f $X=1.635 $Y=0.935 $X2=0 $Y2=0
cc_220 N_A2_c_239_n N_VGND_c_517_n 0.00703954f $X=1.62 $Y=0.77 $X2=0 $Y2=0
cc_221 A2 A_330_48# 0.00400584f $X=1.595 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_222 N_A1_M1007_g N_B1_M1002_g 0.0373947f $X=2.285 $Y=2.75 $X2=0 $Y2=0
cc_223 N_A1_M1001_g N_B1_M1010_g 0.012458f $X=2.115 $Y=0.45 $X2=0 $Y2=0
cc_224 A1 N_B1_M1010_g 0.00401949f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_225 N_A1_c_281_n N_B1_c_328_n 0.0137828f $X=2.205 $Y=1.585 $X2=0 $Y2=0
cc_226 N_A1_c_282_n N_B1_c_329_n 0.0137828f $X=2.205 $Y=1.75 $X2=0 $Y2=0
cc_227 A1 N_B1_c_330_n 5.8438e-19 $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_228 N_A1_c_284_n N_B1_c_330_n 0.0137828f $X=2.205 $Y=1.245 $X2=0 $Y2=0
cc_229 N_A1_M1007_g N_B1_c_331_n 7.85348e-19 $X=2.285 $Y=2.75 $X2=0 $Y2=0
cc_230 A1 N_B1_c_331_n 0.0620003f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_231 N_A1_c_284_n N_B1_c_331_n 0.00448642f $X=2.205 $Y=1.245 $X2=0 $Y2=0
cc_232 N_A1_M1007_g N_VPWR_c_445_n 0.00410918f $X=2.285 $Y=2.75 $X2=0 $Y2=0
cc_233 N_A1_M1007_g N_VPWR_c_440_n 0.00634261f $X=2.285 $Y=2.75 $X2=0 $Y2=0
cc_234 N_A1_M1007_g N_VPWR_c_447_n 0.00355844f $X=2.285 $Y=2.75 $X2=0 $Y2=0
cc_235 N_A1_M1007_g N_A_224_486#_c_483_n 0.0112566f $X=2.285 $Y=2.75 $X2=0 $Y2=0
cc_236 N_A1_M1007_g N_A_224_486#_c_488_n 0.0105488f $X=2.285 $Y=2.75 $X2=0 $Y2=0
cc_237 N_A1_M1001_g N_VGND_c_515_n 0.00376923f $X=2.115 $Y=0.45 $X2=0 $Y2=0
cc_238 A1 N_VGND_c_515_n 0.0094923f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_239 N_A1_M1001_g N_VGND_c_517_n 0.00631815f $X=2.115 $Y=0.45 $X2=0 $Y2=0
cc_240 A1 N_VGND_c_517_n 0.00977804f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_241 N_B1_M1010_g N_C1_M1003_g 0.0426021f $X=2.835 $Y=0.45 $X2=0 $Y2=0
cc_242 N_B1_c_331_n N_C1_M1003_g 3.24328e-19 $X=2.745 $Y=1.245 $X2=0 $Y2=0
cc_243 N_B1_M1002_g N_C1_c_377_n 0.00733604f $X=2.715 $Y=2.75 $X2=0 $Y2=0
cc_244 N_B1_c_329_n N_C1_c_377_n 0.00728272f $X=2.745 $Y=1.75 $X2=0 $Y2=0
cc_245 N_B1_c_331_n N_C1_c_377_n 3.06993e-19 $X=2.745 $Y=1.245 $X2=0 $Y2=0
cc_246 N_B1_M1002_g N_C1_c_378_n 0.0722268f $X=2.715 $Y=2.75 $X2=0 $Y2=0
cc_247 N_B1_c_328_n N_C1_c_375_n 0.00728272f $X=2.745 $Y=1.585 $X2=0 $Y2=0
cc_248 N_B1_c_331_n N_C1_c_375_n 2.36439e-19 $X=2.745 $Y=1.245 $X2=0 $Y2=0
cc_249 N_B1_M1002_g N_VPWR_c_445_n 0.00526824f $X=2.715 $Y=2.75 $X2=0 $Y2=0
cc_250 N_B1_M1002_g N_VPWR_c_440_n 0.00970393f $X=2.715 $Y=2.75 $X2=0 $Y2=0
cc_251 N_B1_M1002_g N_A_224_486#_c_483_n 0.00306928f $X=2.715 $Y=2.75 $X2=0
+ $Y2=0
cc_252 N_B1_M1002_g N_A_224_486#_c_488_n 0.00651011f $X=2.715 $Y=2.75 $X2=0
+ $Y2=0
cc_253 N_B1_M1010_g N_VGND_c_512_n 0.00928184f $X=2.835 $Y=0.45 $X2=0 $Y2=0
cc_254 N_B1_M1010_g N_VGND_c_515_n 0.00391173f $X=2.835 $Y=0.45 $X2=0 $Y2=0
cc_255 N_B1_M1010_g N_VGND_c_517_n 0.00528383f $X=2.835 $Y=0.45 $X2=0 $Y2=0
cc_256 N_C1_M1000_g N_VPWR_c_445_n 0.00371938f $X=3.075 $Y=2.75 $X2=0 $Y2=0
cc_257 N_C1_M1000_g N_VPWR_c_440_n 0.00677341f $X=3.075 $Y=2.75 $X2=0 $Y2=0
cc_258 N_C1_M1000_g N_A_224_486#_c_483_n 4.32374e-19 $X=3.075 $Y=2.75 $X2=0
+ $Y2=0
cc_259 N_C1_M1000_g N_A_224_486#_c_488_n 0.00114807f $X=3.075 $Y=2.75 $X2=0
+ $Y2=0
cc_260 N_C1_M1003_g N_VGND_c_512_n 0.00922356f $X=3.265 $Y=0.45 $X2=0 $Y2=0
cc_261 N_C1_M1003_g N_VGND_c_516_n 0.00391173f $X=3.265 $Y=0.45 $X2=0 $Y2=0
cc_262 N_C1_M1003_g N_VGND_c_517_n 0.00574249f $X=3.265 $Y=0.45 $X2=0 $Y2=0
cc_263 N_X_c_416_n N_VPWR_c_441_n 0.0273301f $X=0.4 $Y=2.575 $X2=0 $Y2=0
cc_264 N_X_c_416_n N_VPWR_c_443_n 0.0341453f $X=0.4 $Y=2.575 $X2=0 $Y2=0
cc_265 N_X_c_416_n N_VPWR_c_440_n 0.0184668f $X=0.4 $Y=2.575 $X2=0 $Y2=0
cc_266 N_X_c_415_n N_VGND_c_513_n 0.026696f $X=0.4 $Y=0.45 $X2=0 $Y2=0
cc_267 N_X_M1006_s N_VGND_c_517_n 0.00215771f $X=0.275 $Y=0.24 $X2=0 $Y2=0
cc_268 N_X_c_415_n N_VGND_c_517_n 0.018188f $X=0.4 $Y=0.45 $X2=0 $Y2=0
cc_269 N_VPWR_c_441_n N_A_224_486#_c_482_n 3.23977e-19 $X=0.83 $Y=2.575 $X2=0
+ $Y2=0
cc_270 N_VPWR_c_442_n N_A_224_486#_c_482_n 0.0234158f $X=1.635 $Y=3.33 $X2=0
+ $Y2=0
cc_271 N_VPWR_c_440_n N_A_224_486#_c_482_n 0.0126396f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_272 N_VPWR_c_447_n N_A_224_486#_c_482_n 0.0127488f $X=2.07 $Y=2.905 $X2=0
+ $Y2=0
cc_273 N_VPWR_M1005_d N_A_224_486#_c_483_n 0.00726743f $X=1.59 $Y=2.43 $X2=0
+ $Y2=0
cc_274 N_VPWR_c_442_n N_A_224_486#_c_483_n 0.00186514f $X=1.635 $Y=3.33 $X2=0
+ $Y2=0
cc_275 N_VPWR_c_445_n N_A_224_486#_c_483_n 0.00186514f $X=3.6 $Y=3.33 $X2=0
+ $Y2=0
cc_276 N_VPWR_c_440_n N_A_224_486#_c_483_n 0.00954917f $X=3.6 $Y=3.33 $X2=0
+ $Y2=0
cc_277 N_VPWR_c_447_n N_A_224_486#_c_483_n 0.0399249f $X=2.07 $Y=2.905 $X2=0
+ $Y2=0
cc_278 N_VPWR_c_441_n N_A_224_486#_c_484_n 0.0016373f $X=0.83 $Y=2.575 $X2=0
+ $Y2=0
cc_279 N_VPWR_c_445_n N_A_224_486#_c_488_n 0.013951f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_280 N_VPWR_c_440_n N_A_224_486#_c_488_n 0.0121125f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_281 N_VGND_c_517_n A_246_48# 0.00626785f $X=3.6 $Y=0 $X2=-0.19 $Y2=-0.245
cc_282 N_VGND_c_517_n A_330_48# 0.0092215f $X=3.6 $Y=0 $X2=-0.19 $Y2=-0.245
