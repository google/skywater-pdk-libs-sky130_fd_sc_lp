* NGSPICE file created from sky130_fd_sc_lp__o211a_m.ext - technology: sky130A

.subckt sky130_fd_sc_lp__o211a_m A1 A2 B1 C1 VGND VNB VPB VPWR X
M1000 VGND A1 a_217_49# VNB nshort w=420000u l=150000u
+  ad=2.625e+11p pd=2.93e+06u as=2.289e+11p ps=2.77e+06u
M1001 a_80_60# C1 VPWR VPB phighvt w=420000u l=150000u
+  ad=2.751e+11p pd=2.99e+06u as=3.36e+11p ps=3.28e+06u
M1002 VGND a_80_60# X VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1003 VPWR a_80_60# X VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1004 VPWR B1 a_80_60# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_217_49# A2 VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_80_60# C1 a_488_49# VNB nshort w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=8.82e+10p ps=1.26e+06u
M1007 a_300_371# A1 VPWR VPB phighvt w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1008 a_488_49# B1 a_217_49# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_80_60# A2 a_300_371# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

