* File: sky130_fd_sc_lp__dfxtp_4.pxi.spice
* Created: Fri Aug 28 10:24:29 2020
* 
x_PM_SKY130_FD_SC_LP__DFXTP_4%CLK N_CLK_c_188_n N_CLK_M1004_g N_CLK_M1023_g
+ N_CLK_c_190_n CLK CLK CLK CLK CLK N_CLK_c_192_n N_CLK_c_193_n
+ PM_SKY130_FD_SC_LP__DFXTP_4%CLK
x_PM_SKY130_FD_SC_LP__DFXTP_4%D N_D_M1019_g N_D_M1027_g N_D_c_217_n N_D_c_218_n
+ N_D_c_219_n D D N_D_c_220_n N_D_c_221_n PM_SKY130_FD_SC_LP__DFXTP_4%D
x_PM_SKY130_FD_SC_LP__DFXTP_4%A_217_413# N_A_217_413#_M1011_s
+ N_A_217_413#_M1015_s N_A_217_413#_M1008_g N_A_217_413#_c_258_n
+ N_A_217_413#_M1005_g N_A_217_413#_M1007_g N_A_217_413#_c_261_n
+ N_A_217_413#_c_271_n N_A_217_413#_c_272_n N_A_217_413#_M1006_g
+ N_A_217_413#_c_262_n N_A_217_413#_c_275_n N_A_217_413#_c_276_n
+ N_A_217_413#_c_277_n N_A_217_413#_c_278_n N_A_217_413#_c_263_n
+ N_A_217_413#_c_280_n N_A_217_413#_c_298_p N_A_217_413#_c_264_n
+ N_A_217_413#_c_282_n N_A_217_413#_c_336_p N_A_217_413#_c_283_n
+ N_A_217_413#_c_284_n N_A_217_413#_c_265_n N_A_217_413#_c_266_n
+ N_A_217_413#_c_267_n PM_SKY130_FD_SC_LP__DFXTP_4%A_217_413#
x_PM_SKY130_FD_SC_LP__DFXTP_4%A_684_93# N_A_684_93#_M1016_d N_A_684_93#_M1003_d
+ N_A_684_93#_M1001_g N_A_684_93#_M1024_g N_A_684_93#_c_431_n
+ N_A_684_93#_c_427_n N_A_684_93#_c_433_n N_A_684_93#_c_434_n
+ N_A_684_93#_c_428_n N_A_684_93#_c_429_n PM_SKY130_FD_SC_LP__DFXTP_4%A_684_93#
x_PM_SKY130_FD_SC_LP__DFXTP_4%A_526_413# N_A_526_413#_M1000_d
+ N_A_526_413#_M1008_d N_A_526_413#_M1003_g N_A_526_413#_M1016_g
+ N_A_526_413#_c_495_n N_A_526_413#_c_496_n N_A_526_413#_c_497_n
+ N_A_526_413#_c_498_n N_A_526_413#_c_499_n N_A_526_413#_c_500_n
+ N_A_526_413#_c_501_n PM_SKY130_FD_SC_LP__DFXTP_4%A_526_413#
x_PM_SKY130_FD_SC_LP__DFXTP_4%A_110_70# N_A_110_70#_M1004_d N_A_110_70#_M1023_d
+ N_A_110_70#_c_567_n N_A_110_70#_c_568_n N_A_110_70#_M1015_g
+ N_A_110_70#_M1011_g N_A_110_70#_c_583_n N_A_110_70#_c_584_n
+ N_A_110_70#_c_571_n N_A_110_70#_c_572_n N_A_110_70#_M1000_g
+ N_A_110_70#_c_574_n N_A_110_70#_M1022_g N_A_110_70#_c_586_n
+ N_A_110_70#_M1021_g N_A_110_70#_M1017_g N_A_110_70#_c_576_n
+ N_A_110_70#_c_577_n N_A_110_70#_c_588_n N_A_110_70#_c_578_n
+ N_A_110_70#_c_579_n N_A_110_70#_c_589_n N_A_110_70#_c_580_n
+ N_A_110_70#_c_581_n N_A_110_70#_c_591_n PM_SKY130_FD_SC_LP__DFXTP_4%A_110_70#
x_PM_SKY130_FD_SC_LP__DFXTP_4%A_1112_93# N_A_1112_93#_M1026_d
+ N_A_1112_93#_M1028_d N_A_1112_93#_M1010_g N_A_1112_93#_M1012_g
+ N_A_1112_93#_M1013_g N_A_1112_93#_M1002_g N_A_1112_93#_M1014_g
+ N_A_1112_93#_M1009_g N_A_1112_93#_M1020_g N_A_1112_93#_M1018_g
+ N_A_1112_93#_M1029_g N_A_1112_93#_M1025_g N_A_1112_93#_c_708_n
+ N_A_1112_93#_c_722_n N_A_1112_93#_c_723_n N_A_1112_93#_c_709_n
+ N_A_1112_93#_c_725_n N_A_1112_93#_c_710_n N_A_1112_93#_c_711_n
+ N_A_1112_93#_c_712_n N_A_1112_93#_c_713_n N_A_1112_93#_c_714_n
+ N_A_1112_93#_c_715_n PM_SKY130_FD_SC_LP__DFXTP_4%A_1112_93#
x_PM_SKY130_FD_SC_LP__DFXTP_4%A_941_379# N_A_941_379#_M1007_d
+ N_A_941_379#_M1021_d N_A_941_379#_M1026_g N_A_941_379#_M1028_g
+ N_A_941_379#_c_850_n N_A_941_379#_c_851_n N_A_941_379#_c_852_n
+ N_A_941_379#_c_853_n N_A_941_379#_c_854_n N_A_941_379#_c_855_n
+ PM_SKY130_FD_SC_LP__DFXTP_4%A_941_379#
x_PM_SKY130_FD_SC_LP__DFXTP_4%VPWR N_VPWR_M1023_s N_VPWR_M1015_d N_VPWR_M1024_d
+ N_VPWR_M1012_d N_VPWR_M1002_d N_VPWR_M1009_d N_VPWR_M1025_d N_VPWR_c_929_n
+ N_VPWR_c_930_n N_VPWR_c_931_n N_VPWR_c_932_n N_VPWR_c_933_n N_VPWR_c_934_n
+ N_VPWR_c_935_n N_VPWR_c_936_n N_VPWR_c_937_n N_VPWR_c_938_n N_VPWR_c_939_n
+ N_VPWR_c_940_n VPWR N_VPWR_c_941_n N_VPWR_c_942_n N_VPWR_c_943_n
+ N_VPWR_c_944_n N_VPWR_c_945_n N_VPWR_c_946_n N_VPWR_c_947_n N_VPWR_c_948_n
+ N_VPWR_c_928_n PM_SKY130_FD_SC_LP__DFXTP_4%VPWR
x_PM_SKY130_FD_SC_LP__DFXTP_4%A_431_119# N_A_431_119#_M1019_d
+ N_A_431_119#_M1027_d N_A_431_119#_c_1047_n N_A_431_119#_c_1048_n
+ N_A_431_119#_c_1051_n N_A_431_119#_c_1046_n
+ PM_SKY130_FD_SC_LP__DFXTP_4%A_431_119#
x_PM_SKY130_FD_SC_LP__DFXTP_4%Q N_Q_M1013_d N_Q_M1020_d N_Q_M1002_s N_Q_M1018_s
+ N_Q_c_1124_p N_Q_c_1108_n N_Q_c_1071_n N_Q_c_1075_n N_Q_c_1076_n N_Q_c_1125_p
+ N_Q_c_1113_n N_Q_c_1077_n Q Q Q Q Q Q N_Q_c_1073_n N_Q_c_1074_n
+ PM_SKY130_FD_SC_LP__DFXTP_4%Q
x_PM_SKY130_FD_SC_LP__DFXTP_4%VGND N_VGND_M1004_s N_VGND_M1011_d N_VGND_M1001_d
+ N_VGND_M1010_d N_VGND_M1013_s N_VGND_M1014_s N_VGND_M1029_s N_VGND_c_1131_n
+ N_VGND_c_1132_n N_VGND_c_1133_n N_VGND_c_1134_n N_VGND_c_1135_n
+ N_VGND_c_1136_n N_VGND_c_1137_n N_VGND_c_1138_n N_VGND_c_1139_n
+ N_VGND_c_1140_n N_VGND_c_1141_n N_VGND_c_1142_n VGND N_VGND_c_1143_n
+ N_VGND_c_1144_n N_VGND_c_1145_n N_VGND_c_1146_n N_VGND_c_1147_n
+ N_VGND_c_1148_n N_VGND_c_1149_n N_VGND_c_1150_n N_VGND_c_1151_n
+ PM_SKY130_FD_SC_LP__DFXTP_4%VGND
cc_1 VNB N_CLK_c_188_n 0.024794f $X=-0.19 $Y=-0.245 $X2=0.352 $Y2=1.353
cc_2 VNB N_CLK_M1023_g 0.00639683f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.66
cc_3 VNB N_CLK_c_190_n 0.0243131f $X=-0.19 $Y=-0.245 $X2=0.352 $Y2=1.55
cc_4 VNB CLK 0.0333978f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_5 VNB N_CLK_c_192_n 0.025499f $X=-0.19 $Y=-0.245 $X2=0.32 $Y2=1.045
cc_6 VNB N_CLK_c_193_n 0.0249498f $X=-0.19 $Y=-0.245 $X2=0.352 $Y2=0.88
cc_7 VNB N_D_c_217_n 0.0171588f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_D_c_218_n 0.0175675f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_9 VNB N_D_c_219_n 0.0114296f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_10 VNB N_D_c_220_n 0.0164255f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_D_c_221_n 0.00770037f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_217_413#_c_258_n 0.0112368f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_13 VNB N_A_217_413#_M1005_g 0.0397652f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=2.32
cc_14 VNB N_A_217_413#_M1007_g 0.023759f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_217_413#_c_261_n 0.00560896f $X=-0.19 $Y=-0.245 $X2=0.32 $Y2=1.045
cc_16 VNB N_A_217_413#_c_262_n 0.005023f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_217_413#_c_263_n 0.00322053f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_217_413#_c_264_n 0.001321f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_217_413#_c_265_n 0.0034738f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_217_413#_c_266_n 0.0534494f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_217_413#_c_267_n 0.0160664f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_684_93#_M1001_g 0.029198f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_684_93#_c_427_n 0.024219f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_684_93#_c_428_n 0.00808095f $X=-0.19 $Y=-0.245 $X2=0.32 $Y2=1.045
cc_25 VNB N_A_684_93#_c_429_n 0.00226342f $X=-0.19 $Y=-0.245 $X2=0.255 $Y2=0.925
cc_26 VNB N_A_526_413#_c_495_n 0.00198257f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_526_413#_c_496_n 0.00290482f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_526_413#_c_497_n 0.0230975f $X=-0.19 $Y=-0.245 $X2=0.32 $Y2=1.045
cc_29 VNB N_A_526_413#_c_498_n 8.42564e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_526_413#_c_499_n 0.028858f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_526_413#_c_500_n 0.00634745f $X=-0.19 $Y=-0.245 $X2=0.255
+ $Y2=1.295
cc_32 VNB N_A_526_413#_c_501_n 0.0175366f $X=-0.19 $Y=-0.245 $X2=0.255 $Y2=2.035
cc_33 VNB N_A_110_70#_c_567_n 0.0146274f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.66
cc_34 VNB N_A_110_70#_c_568_n 0.0184716f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.66
cc_35 VNB N_A_110_70#_M1015_g 0.0147788f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_36 VNB N_A_110_70#_M1011_g 0.0352568f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_110_70#_c_571_n 0.0642759f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_110_70#_c_572_n 0.012806f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_110_70#_M1000_g 0.0387206f $X=-0.19 $Y=-0.245 $X2=0.32 $Y2=1.045
cc_40 VNB N_A_110_70#_c_574_n 0.205137f $X=-0.19 $Y=-0.245 $X2=0.255 $Y2=0.925
cc_41 VNB N_A_110_70#_M1017_g 0.0348281f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_110_70#_c_576_n 0.0143713f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_110_70#_c_577_n 0.00749069f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_110_70#_c_578_n 0.0149542f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_110_70#_c_579_n 0.00137438f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_110_70#_c_580_n 0.00834834f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_110_70#_c_581_n 0.0190456f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_1112_93#_M1010_g 0.0267704f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_1112_93#_M1012_g 0.00120551f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_50 VNB N_A_1112_93#_M1013_g 0.027912f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_1112_93#_M1002_g 5.57101e-19 $X=-0.19 $Y=-0.245 $X2=0.352
+ $Y2=1.045
cc_52 VNB N_A_1112_93#_M1014_g 0.0213292f $X=-0.19 $Y=-0.245 $X2=0.255 $Y2=0.925
cc_53 VNB N_A_1112_93#_M1009_g 4.57707e-19 $X=-0.19 $Y=-0.245 $X2=0.255
+ $Y2=1.295
cc_54 VNB N_A_1112_93#_M1020_g 0.0213088f $X=-0.19 $Y=-0.245 $X2=0.255 $Y2=2.035
cc_55 VNB N_A_1112_93#_M1018_g 4.57404e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_1112_93#_M1029_g 0.0259216f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_1112_93#_M1025_g 4.93851e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_1112_93#_c_708_n 2.86442e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_1112_93#_c_709_n 0.0018533f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_1112_93#_c_710_n 0.0105987f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_A_1112_93#_c_711_n 0.00649282f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_A_1112_93#_c_712_n 0.00905732f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_A_1112_93#_c_713_n 0.0383373f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_A_1112_93#_c_714_n 0.0372674f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_A_1112_93#_c_715_n 0.0727247f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_A_941_379#_M1028_g 0.00182145f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_67 VNB N_A_941_379#_c_850_n 0.00169389f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.95
cc_68 VNB N_A_941_379#_c_851_n 0.00517363f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_941_379#_c_852_n 0.0185498f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_A_941_379#_c_853_n 0.00156209f $X=-0.19 $Y=-0.245 $X2=0.352 $Y2=0.88
cc_71 VNB N_A_941_379#_c_854_n 0.0360596f $X=-0.19 $Y=-0.245 $X2=0.255 $Y2=0.925
cc_72 VNB N_A_941_379#_c_855_n 0.0227923f $X=-0.19 $Y=-0.245 $X2=0.255 $Y2=1.665
cc_73 VNB N_VPWR_c_928_n 0.382608f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_A_431_119#_c_1046_n 0.0134295f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_Q_c_1071_n 0.00369191f $X=-0.19 $Y=-0.245 $X2=0.352 $Y2=0.88
cc_76 VNB Q 0.022474f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_Q_c_1073_n 0.00304538f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_Q_c_1074_n 0.021559f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_VGND_c_1131_n 0.0112376f $X=-0.19 $Y=-0.245 $X2=0.32 $Y2=1.045
cc_80 VNB N_VGND_c_1132_n 0.0216486f $X=-0.19 $Y=-0.245 $X2=0.352 $Y2=0.88
cc_81 VNB N_VGND_c_1133_n 0.010047f $X=-0.19 $Y=-0.245 $X2=0.255 $Y2=1.045
cc_82 VNB N_VGND_c_1134_n 0.0206848f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_VGND_c_1135_n 0.0104512f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_VGND_c_1136_n 0.0227912f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_VGND_c_1137_n 0.0159764f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_VGND_c_1138_n 3.16049e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_VGND_c_1139_n 0.0108441f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_VGND_c_1140_n 0.0197175f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_VGND_c_1141_n 0.0498005f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_VGND_c_1142_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_VGND_c_1143_n 0.0345113f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_VGND_c_1144_n 0.0515635f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_93 VNB N_VGND_c_1145_n 0.0148832f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_94 VNB N_VGND_c_1146_n 0.0129398f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_95 VNB N_VGND_c_1147_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_96 VNB N_VGND_c_1148_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_97 VNB N_VGND_c_1149_n 0.00557808f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_98 VNB N_VGND_c_1150_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_99 VNB N_VGND_c_1151_n 0.472108f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_100 VPB N_CLK_M1023_g 0.0603647f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.66
cc_101 VPB CLK 0.0350833f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_102 VPB N_D_M1027_g 0.026317f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=1.55
cc_103 VPB N_D_c_219_n 0.0168082f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_104 VPB N_D_c_221_n 0.00619922f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_105 VPB N_A_217_413#_M1008_g 0.0206607f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_106 VPB N_A_217_413#_c_258_n 0.0145904f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_107 VPB N_A_217_413#_c_261_n 0.0100553f $X=-0.19 $Y=1.655 $X2=0.32 $Y2=1.045
cc_108 VPB N_A_217_413#_c_271_n 0.0283922f $X=-0.19 $Y=1.655 $X2=0.32 $Y2=1.045
cc_109 VPB N_A_217_413#_c_272_n 0.0119087f $X=-0.19 $Y=1.655 $X2=0.352 $Y2=0.88
cc_110 VPB N_A_217_413#_M1006_g 0.0255974f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_111 VPB N_A_217_413#_c_262_n 0.00300491f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_112 VPB N_A_217_413#_c_275_n 0.00710388f $X=-0.19 $Y=1.655 $X2=0.255
+ $Y2=2.035
cc_113 VPB N_A_217_413#_c_276_n 3.40079e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_114 VPB N_A_217_413#_c_277_n 0.0096403f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_115 VPB N_A_217_413#_c_278_n 0.00271588f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_116 VPB N_A_217_413#_c_263_n 0.00189472f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_117 VPB N_A_217_413#_c_280_n 0.0124088f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_118 VPB N_A_217_413#_c_264_n 0.00402248f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_119 VPB N_A_217_413#_c_282_n 0.0140188f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_120 VPB N_A_217_413#_c_283_n 0.00159986f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_121 VPB N_A_217_413#_c_284_n 0.00383404f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_122 VPB N_A_217_413#_c_267_n 0.0252621f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_123 VPB N_A_684_93#_M1024_g 0.0312426f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_124 VPB N_A_684_93#_c_431_n 0.0029759f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_125 VPB N_A_684_93#_c_427_n 0.00791434f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_126 VPB N_A_684_93#_c_433_n 0.00784958f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_127 VPB N_A_684_93#_c_434_n 0.00176458f $X=-0.19 $Y=1.655 $X2=0.352 $Y2=1.045
cc_128 VPB N_A_684_93#_c_428_n 0.00246451f $X=-0.19 $Y=1.655 $X2=0.32 $Y2=1.045
cc_129 VPB N_A_526_413#_M1003_g 0.0224934f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_130 VPB N_A_526_413#_c_496_n 0.00641718f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_131 VPB N_A_526_413#_c_498_n 0.00156562f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_132 VPB N_A_526_413#_c_499_n 0.00686781f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_133 VPB N_A_110_70#_M1015_g 0.0504359f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_134 VPB N_A_110_70#_c_583_n 0.124953f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_135 VPB N_A_110_70#_c_584_n 0.012806f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_136 VPB N_A_110_70#_M1022_g 0.0587785f $X=-0.19 $Y=1.655 $X2=0.255 $Y2=1.295
cc_137 VPB N_A_110_70#_c_586_n 0.099865f $X=-0.19 $Y=1.655 $X2=0.255 $Y2=1.665
cc_138 VPB N_A_110_70#_M1021_g 0.0423797f $X=-0.19 $Y=1.655 $X2=0.255 $Y2=2.405
cc_139 VPB N_A_110_70#_c_588_n 0.00749069f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_140 VPB N_A_110_70#_c_589_n 0.019077f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_141 VPB N_A_110_70#_c_581_n 0.0226415f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_142 VPB N_A_110_70#_c_591_n 0.00830723f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_143 VPB N_A_1112_93#_M1012_g 0.0429565f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_144 VPB N_A_1112_93#_M1002_g 0.0242718f $X=-0.19 $Y=1.655 $X2=0.352 $Y2=1.045
cc_145 VPB N_A_1112_93#_M1009_g 0.0187468f $X=-0.19 $Y=1.655 $X2=0.255 $Y2=1.295
cc_146 VPB N_A_1112_93#_M1018_g 0.0187266f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_147 VPB N_A_1112_93#_M1025_g 0.0225355f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_148 VPB N_A_1112_93#_c_708_n 2.79281e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_149 VPB N_A_1112_93#_c_722_n 0.00803288f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_150 VPB N_A_1112_93#_c_723_n 0.00919925f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_151 VPB N_A_1112_93#_c_709_n 0.00848735f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_152 VPB N_A_1112_93#_c_725_n 0.0118759f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_153 VPB N_A_1112_93#_c_711_n 0.00546222f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_154 VPB N_A_1112_93#_c_714_n 0.00214235f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_155 VPB N_A_941_379#_M1028_g 0.0254049f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_156 VPB N_A_941_379#_c_851_n 0.00536555f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_157 VPB N_VPWR_c_929_n 0.0112117f $X=-0.19 $Y=1.655 $X2=0.32 $Y2=1.045
cc_158 VPB N_VPWR_c_930_n 0.0214587f $X=-0.19 $Y=1.655 $X2=0.352 $Y2=0.88
cc_159 VPB N_VPWR_c_931_n 0.0180505f $X=-0.19 $Y=1.655 $X2=0.255 $Y2=1.045
cc_160 VPB N_VPWR_c_932_n 0.0113065f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_161 VPB N_VPWR_c_933_n 0.02069f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_162 VPB N_VPWR_c_934_n 0.0173908f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_163 VPB N_VPWR_c_935_n 0.0184865f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_164 VPB N_VPWR_c_936_n 3.15212e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_165 VPB N_VPWR_c_937_n 0.0108182f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_166 VPB N_VPWR_c_938_n 0.0197167f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_167 VPB N_VPWR_c_939_n 0.0588727f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_168 VPB N_VPWR_c_940_n 0.00594246f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_169 VPB N_VPWR_c_941_n 0.0306255f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_170 VPB N_VPWR_c_942_n 0.055386f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_171 VPB N_VPWR_c_943_n 0.0147711f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_172 VPB N_VPWR_c_944_n 0.0129398f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_173 VPB N_VPWR_c_945_n 0.00250432f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_174 VPB N_VPWR_c_946_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_175 VPB N_VPWR_c_947_n 0.00564836f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_176 VPB N_VPWR_c_948_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_177 VPB N_VPWR_c_928_n 0.111905f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_178 VPB N_A_431_119#_c_1047_n 0.00222478f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_179 VPB N_A_431_119#_c_1048_n 8.39791e-19 $X=-0.19 $Y=1.655 $X2=0.155
+ $Y2=0.84
cc_180 VPB N_A_431_119#_c_1046_n 0.0052586f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_181 VPB N_Q_c_1075_n 0.00304538f $X=-0.19 $Y=1.655 $X2=0.255 $Y2=0.925
cc_182 VPB N_Q_c_1076_n 0.00296628f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_183 VPB N_Q_c_1077_n 0.00144145f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_184 VPB Q 0.0109235f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_185 VPB Q 0.0216433f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_186 VPB Q 0.00402406f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_187 N_CLK_c_188_n N_A_110_70#_c_568_n 0.018028f $X=0.352 $Y=1.353 $X2=0 $Y2=0
cc_188 CLK N_A_110_70#_c_568_n 5.05264e-19 $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_189 CLK N_A_110_70#_c_578_n 0.12421f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_190 N_CLK_c_193_n N_A_110_70#_c_578_n 0.00571717f $X=0.352 $Y=0.88 $X2=0
+ $Y2=0
cc_191 N_CLK_c_188_n N_A_110_70#_c_579_n 0.00571717f $X=0.352 $Y=1.353 $X2=0
+ $Y2=0
cc_192 N_CLK_M1023_g N_A_110_70#_c_589_n 0.00571717f $X=0.475 $Y=2.66 $X2=0
+ $Y2=0
cc_193 N_CLK_c_192_n N_A_110_70#_c_580_n 0.00571717f $X=0.32 $Y=1.045 $X2=0
+ $Y2=0
cc_194 N_CLK_c_190_n N_A_110_70#_c_581_n 0.018028f $X=0.352 $Y=1.55 $X2=0 $Y2=0
cc_195 N_CLK_c_190_n N_A_110_70#_c_591_n 0.00571717f $X=0.352 $Y=1.55 $X2=0
+ $Y2=0
cc_196 CLK N_VPWR_M1023_s 0.00300356f $X=0.155 $Y=0.84 $X2=-0.19 $Y2=-0.245
cc_197 N_CLK_M1023_g N_VPWR_c_930_n 0.0115546f $X=0.475 $Y=2.66 $X2=0 $Y2=0
cc_198 CLK N_VPWR_c_930_n 0.0232425f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_199 N_CLK_M1023_g N_VPWR_c_941_n 0.00396895f $X=0.475 $Y=2.66 $X2=0 $Y2=0
cc_200 N_CLK_M1023_g N_VPWR_c_928_n 0.00796233f $X=0.475 $Y=2.66 $X2=0 $Y2=0
cc_201 CLK N_VPWR_c_928_n 0.00159622f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_202 CLK N_VGND_c_1132_n 0.0266997f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_203 N_CLK_c_192_n N_VGND_c_1132_n 0.00156152f $X=0.32 $Y=1.045 $X2=0 $Y2=0
cc_204 N_CLK_c_193_n N_VGND_c_1132_n 0.0134006f $X=0.352 $Y=0.88 $X2=0 $Y2=0
cc_205 N_CLK_c_193_n N_VGND_c_1143_n 0.00396895f $X=0.352 $Y=0.88 $X2=0 $Y2=0
cc_206 CLK N_VGND_c_1151_n 0.0015796f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_207 N_CLK_c_193_n N_VGND_c_1151_n 0.00796233f $X=0.352 $Y=0.88 $X2=0 $Y2=0
cc_208 N_D_M1027_g N_A_217_413#_M1008_g 0.0148077f $X=2.125 $Y=2.275 $X2=0 $Y2=0
cc_209 N_D_M1027_g N_A_217_413#_c_262_n 0.00111981f $X=2.125 $Y=2.275 $X2=0
+ $Y2=0
cc_210 N_D_c_220_n N_A_217_413#_c_262_n 4.38778e-19 $X=1.99 $Y=1.29 $X2=0 $Y2=0
cc_211 N_D_c_221_n N_A_217_413#_c_262_n 0.05234f $X=1.99 $Y=1.29 $X2=0 $Y2=0
cc_212 N_D_M1027_g N_A_217_413#_c_275_n 0.0053131f $X=2.125 $Y=2.275 $X2=0 $Y2=0
cc_213 N_D_c_219_n N_A_217_413#_c_275_n 0.00158631f $X=2.012 $Y=1.795 $X2=0
+ $Y2=0
cc_214 N_D_c_221_n N_A_217_413#_c_275_n 0.0315771f $X=1.99 $Y=1.29 $X2=0 $Y2=0
cc_215 N_D_M1027_g N_A_217_413#_c_276_n 0.0083829f $X=2.125 $Y=2.275 $X2=0 $Y2=0
cc_216 N_D_M1027_g N_A_217_413#_c_277_n 0.00848284f $X=2.125 $Y=2.275 $X2=0
+ $Y2=0
cc_217 N_D_M1027_g N_A_217_413#_c_278_n 0.00139353f $X=2.125 $Y=2.275 $X2=0
+ $Y2=0
cc_218 N_D_M1027_g N_A_217_413#_c_263_n 7.18735e-19 $X=2.125 $Y=2.275 $X2=0
+ $Y2=0
cc_219 N_D_c_219_n N_A_217_413#_c_267_n 0.0148077f $X=2.012 $Y=1.795 $X2=0 $Y2=0
cc_220 N_D_M1027_g N_A_110_70#_M1015_g 0.012766f $X=2.125 $Y=2.275 $X2=0 $Y2=0
cc_221 N_D_c_218_n N_A_110_70#_M1015_g 0.0147499f $X=2.012 $Y=1.535 $X2=0 $Y2=0
cc_222 N_D_c_221_n N_A_110_70#_M1015_g 0.00356161f $X=1.99 $Y=1.29 $X2=0 $Y2=0
cc_223 N_D_c_217_n N_A_110_70#_M1011_g 0.0109826f $X=1.99 $Y=1.125 $X2=0 $Y2=0
cc_224 N_D_c_220_n N_A_110_70#_M1011_g 0.00711562f $X=1.99 $Y=1.29 $X2=0 $Y2=0
cc_225 N_D_c_221_n N_A_110_70#_M1011_g 0.00316885f $X=1.99 $Y=1.29 $X2=0 $Y2=0
cc_226 N_D_M1027_g N_A_110_70#_c_583_n 0.00316148f $X=2.125 $Y=2.275 $X2=0 $Y2=0
cc_227 N_D_c_217_n N_A_110_70#_c_571_n 0.0104164f $X=1.99 $Y=1.125 $X2=0 $Y2=0
cc_228 N_D_c_217_n N_A_110_70#_M1000_g 0.0125895f $X=1.99 $Y=1.125 $X2=0 $Y2=0
cc_229 N_D_c_218_n N_A_110_70#_c_576_n 0.00711562f $X=2.012 $Y=1.535 $X2=0 $Y2=0
cc_230 N_D_c_221_n N_A_110_70#_c_576_n 0.00475747f $X=1.99 $Y=1.29 $X2=0 $Y2=0
cc_231 N_D_M1027_g N_VPWR_c_931_n 6.15821e-19 $X=2.125 $Y=2.275 $X2=0 $Y2=0
cc_232 N_D_M1027_g N_A_431_119#_c_1047_n 0.00423488f $X=2.125 $Y=2.275 $X2=0
+ $Y2=0
cc_233 N_D_c_217_n N_A_431_119#_c_1051_n 0.00319919f $X=1.99 $Y=1.125 $X2=0
+ $Y2=0
cc_234 N_D_c_217_n N_A_431_119#_c_1046_n 0.0138015f $X=1.99 $Y=1.125 $X2=0 $Y2=0
cc_235 N_D_c_219_n N_A_431_119#_c_1046_n 0.00423488f $X=2.012 $Y=1.795 $X2=0
+ $Y2=0
cc_236 N_D_c_221_n N_A_431_119#_c_1046_n 0.0518775f $X=1.99 $Y=1.29 $X2=0 $Y2=0
cc_237 N_D_c_217_n N_VGND_c_1133_n 0.00391586f $X=1.99 $Y=1.125 $X2=0 $Y2=0
cc_238 N_D_c_220_n N_VGND_c_1133_n 0.00111171f $X=1.99 $Y=1.29 $X2=0 $Y2=0
cc_239 N_D_c_221_n N_VGND_c_1133_n 0.0270791f $X=1.99 $Y=1.29 $X2=0 $Y2=0
cc_240 N_D_c_217_n N_VGND_c_1151_n 9.39239e-19 $X=1.99 $Y=1.125 $X2=0 $Y2=0
cc_241 N_A_217_413#_c_298_p N_A_684_93#_M1003_d 0.00529129f $X=4.76 $Y=2.37
+ $X2=0 $Y2=0
cc_242 N_A_217_413#_M1005_g N_A_684_93#_M1001_g 0.0379268f $X=3.135 $Y=0.805
+ $X2=0 $Y2=0
cc_243 N_A_217_413#_c_298_p N_A_684_93#_M1024_g 0.0102944f $X=4.76 $Y=2.37 $X2=0
+ $Y2=0
cc_244 N_A_217_413#_c_284_n N_A_684_93#_M1024_g 0.00309856f $X=3.41 $Y=2.37
+ $X2=0 $Y2=0
cc_245 N_A_217_413#_c_267_n N_A_684_93#_M1024_g 0.00178452f $X=2.855 $Y=1.71
+ $X2=0 $Y2=0
cc_246 N_A_217_413#_M1005_g N_A_684_93#_c_431_n 9.48507e-19 $X=3.135 $Y=0.805
+ $X2=0 $Y2=0
cc_247 N_A_217_413#_c_258_n N_A_684_93#_c_427_n 0.0379268f $X=3.06 $Y=1.62 $X2=0
+ $Y2=0
cc_248 N_A_217_413#_c_284_n N_A_684_93#_c_427_n 2.18062e-19 $X=3.41 $Y=2.37
+ $X2=0 $Y2=0
cc_249 N_A_217_413#_c_298_p N_A_684_93#_c_433_n 0.0386036f $X=4.76 $Y=2.37 $X2=0
+ $Y2=0
cc_250 N_A_217_413#_c_298_p N_A_684_93#_c_434_n 0.0116559f $X=4.76 $Y=2.37 $X2=0
+ $Y2=0
cc_251 N_A_217_413#_c_284_n N_A_684_93#_c_434_n 0.00547817f $X=3.41 $Y=2.37
+ $X2=0 $Y2=0
cc_252 N_A_217_413#_c_298_p N_A_684_93#_c_428_n 0.0105058f $X=4.76 $Y=2.37 $X2=0
+ $Y2=0
cc_253 N_A_217_413#_c_264_n N_A_684_93#_c_428_n 0.0232735f $X=4.845 $Y=2.285
+ $X2=0 $Y2=0
cc_254 N_A_217_413#_c_265_n N_A_684_93#_c_428_n 0.023884f $X=4.825 $Y=1.39 $X2=0
+ $Y2=0
cc_255 N_A_217_413#_c_266_n N_A_684_93#_c_428_n 0.0028159f $X=4.825 $Y=1.39
+ $X2=0 $Y2=0
cc_256 N_A_217_413#_M1007_g N_A_684_93#_c_429_n 0.00735362f $X=4.77 $Y=0.805
+ $X2=0 $Y2=0
cc_257 N_A_217_413#_c_263_n N_A_526_413#_M1008_d 0.00451021f $X=2.69 $Y=1.71
+ $X2=0 $Y2=0
cc_258 N_A_217_413#_c_298_p N_A_526_413#_M1003_g 0.0119921f $X=4.76 $Y=2.37
+ $X2=0 $Y2=0
cc_259 N_A_217_413#_c_284_n N_A_526_413#_M1003_g 6.84237e-19 $X=3.41 $Y=2.37
+ $X2=0 $Y2=0
cc_260 N_A_217_413#_M1005_g N_A_526_413#_c_495_n 0.00274127f $X=3.135 $Y=0.805
+ $X2=0 $Y2=0
cc_261 N_A_217_413#_M1008_g N_A_526_413#_c_496_n 0.00146724f $X=2.555 $Y=2.275
+ $X2=0 $Y2=0
cc_262 N_A_217_413#_c_258_n N_A_526_413#_c_496_n 0.0134803f $X=3.06 $Y=1.62
+ $X2=0 $Y2=0
cc_263 N_A_217_413#_M1005_g N_A_526_413#_c_496_n 0.00681316f $X=3.135 $Y=0.805
+ $X2=0 $Y2=0
cc_264 N_A_217_413#_c_263_n N_A_526_413#_c_496_n 0.0593984f $X=2.69 $Y=1.71
+ $X2=0 $Y2=0
cc_265 N_A_217_413#_c_280_n N_A_526_413#_c_496_n 0.0148002f $X=3.325 $Y=2.62
+ $X2=0 $Y2=0
cc_266 N_A_217_413#_c_267_n N_A_526_413#_c_496_n 0.00229229f $X=2.855 $Y=1.71
+ $X2=0 $Y2=0
cc_267 N_A_217_413#_M1005_g N_A_526_413#_c_497_n 0.007872f $X=3.135 $Y=0.805
+ $X2=0 $Y2=0
cc_268 N_A_217_413#_M1005_g N_A_526_413#_c_500_n 0.0124827f $X=3.135 $Y=0.805
+ $X2=0 $Y2=0
cc_269 N_A_217_413#_c_263_n N_A_526_413#_c_500_n 0.00427303f $X=2.69 $Y=1.71
+ $X2=0 $Y2=0
cc_270 N_A_217_413#_c_267_n N_A_526_413#_c_500_n 0.00748768f $X=2.855 $Y=1.71
+ $X2=0 $Y2=0
cc_271 N_A_217_413#_M1007_g N_A_526_413#_c_501_n 0.0137007f $X=4.77 $Y=0.805
+ $X2=0 $Y2=0
cc_272 N_A_217_413#_c_266_n N_A_526_413#_c_501_n 0.00901731f $X=4.825 $Y=1.39
+ $X2=0 $Y2=0
cc_273 N_A_217_413#_c_262_n N_A_110_70#_c_567_n 0.00892691f $X=1.305 $Y=2.045
+ $X2=0 $Y2=0
cc_274 N_A_217_413#_c_262_n N_A_110_70#_M1015_g 0.0180764f $X=1.305 $Y=2.045
+ $X2=0 $Y2=0
cc_275 N_A_217_413#_c_275_n N_A_110_70#_M1015_g 0.0123887f $X=1.905 $Y=2.13
+ $X2=0 $Y2=0
cc_276 N_A_217_413#_c_276_n N_A_110_70#_M1015_g 0.00155565f $X=1.99 $Y=2.535
+ $X2=0 $Y2=0
cc_277 N_A_217_413#_c_282_n N_A_110_70#_M1015_g 0.00457378f $X=1.21 $Y=2.21
+ $X2=0 $Y2=0
cc_278 N_A_217_413#_c_262_n N_A_110_70#_M1011_g 0.00616984f $X=1.305 $Y=2.045
+ $X2=0 $Y2=0
cc_279 N_A_217_413#_c_336_p N_A_110_70#_M1011_g 0.00403215f $X=1.325 $Y=0.805
+ $X2=0 $Y2=0
cc_280 N_A_217_413#_M1008_g N_A_110_70#_c_583_n 0.00316141f $X=2.555 $Y=2.275
+ $X2=0 $Y2=0
cc_281 N_A_217_413#_c_277_n N_A_110_70#_c_583_n 0.00686109f $X=2.595 $Y=2.62
+ $X2=0 $Y2=0
cc_282 N_A_217_413#_c_278_n N_A_110_70#_c_583_n 0.00304989f $X=2.075 $Y=2.62
+ $X2=0 $Y2=0
cc_283 N_A_217_413#_c_280_n N_A_110_70#_c_583_n 0.00562499f $X=3.325 $Y=2.62
+ $X2=0 $Y2=0
cc_284 N_A_217_413#_c_283_n N_A_110_70#_c_583_n 0.00316385f $X=2.685 $Y=2.62
+ $X2=0 $Y2=0
cc_285 N_A_217_413#_M1005_g N_A_110_70#_M1000_g 0.0137363f $X=3.135 $Y=0.805
+ $X2=0 $Y2=0
cc_286 N_A_217_413#_c_263_n N_A_110_70#_M1000_g 6.2237e-19 $X=2.69 $Y=1.71 $X2=0
+ $Y2=0
cc_287 N_A_217_413#_c_267_n N_A_110_70#_M1000_g 0.00539331f $X=2.855 $Y=1.71
+ $X2=0 $Y2=0
cc_288 N_A_217_413#_M1005_g N_A_110_70#_c_574_n 0.0104164f $X=3.135 $Y=0.805
+ $X2=0 $Y2=0
cc_289 N_A_217_413#_M1007_g N_A_110_70#_c_574_n 0.0104164f $X=4.77 $Y=0.805
+ $X2=0 $Y2=0
cc_290 N_A_217_413#_M1008_g N_A_110_70#_M1022_g 0.00806439f $X=2.555 $Y=2.275
+ $X2=0 $Y2=0
cc_291 N_A_217_413#_c_258_n N_A_110_70#_M1022_g 0.00212758f $X=3.06 $Y=1.62
+ $X2=0 $Y2=0
cc_292 N_A_217_413#_c_263_n N_A_110_70#_M1022_g 0.00191521f $X=2.69 $Y=1.71
+ $X2=0 $Y2=0
cc_293 N_A_217_413#_c_280_n N_A_110_70#_M1022_g 0.0158389f $X=3.325 $Y=2.62
+ $X2=0 $Y2=0
cc_294 N_A_217_413#_c_284_n N_A_110_70#_M1022_g 0.00798039f $X=3.41 $Y=2.37
+ $X2=0 $Y2=0
cc_295 N_A_217_413#_c_298_p N_A_110_70#_c_586_n 0.00638427f $X=4.76 $Y=2.37
+ $X2=0 $Y2=0
cc_296 N_A_217_413#_c_284_n N_A_110_70#_c_586_n 0.00139589f $X=3.41 $Y=2.37
+ $X2=0 $Y2=0
cc_297 N_A_217_413#_c_261_n N_A_110_70#_M1021_g 0.00638636f $X=5.105 $Y=1.825
+ $X2=0 $Y2=0
cc_298 N_A_217_413#_c_298_p N_A_110_70#_M1021_g 0.0194848f $X=4.76 $Y=2.37 $X2=0
+ $Y2=0
cc_299 N_A_217_413#_c_264_n N_A_110_70#_M1021_g 0.00735955f $X=4.845 $Y=2.285
+ $X2=0 $Y2=0
cc_300 N_A_217_413#_c_266_n N_A_110_70#_M1021_g 0.00359963f $X=4.825 $Y=1.39
+ $X2=0 $Y2=0
cc_301 N_A_217_413#_M1007_g N_A_110_70#_M1017_g 0.0152311f $X=4.77 $Y=0.805
+ $X2=0 $Y2=0
cc_302 N_A_217_413#_c_271_n N_A_110_70#_M1017_g 0.00155915f $X=5.43 $Y=1.9 $X2=0
+ $Y2=0
cc_303 N_A_217_413#_c_262_n N_A_110_70#_c_576_n 0.00413091f $X=1.305 $Y=2.045
+ $X2=0 $Y2=0
cc_304 N_A_217_413#_c_336_p N_A_110_70#_c_578_n 0.026572f $X=1.325 $Y=0.805
+ $X2=0 $Y2=0
cc_305 N_A_217_413#_c_262_n N_A_110_70#_c_589_n 0.0086706f $X=1.305 $Y=2.045
+ $X2=0 $Y2=0
cc_306 N_A_217_413#_c_282_n N_A_110_70#_c_589_n 0.0508726f $X=1.21 $Y=2.21 $X2=0
+ $Y2=0
cc_307 N_A_217_413#_c_262_n N_A_110_70#_c_580_n 0.0515636f $X=1.305 $Y=2.045
+ $X2=0 $Y2=0
cc_308 N_A_217_413#_c_262_n N_A_110_70#_c_581_n 0.00352999f $X=1.305 $Y=2.045
+ $X2=0 $Y2=0
cc_309 N_A_217_413#_c_282_n N_A_110_70#_c_581_n 0.003061f $X=1.21 $Y=2.21 $X2=0
+ $Y2=0
cc_310 N_A_217_413#_M1007_g N_A_1112_93#_M1010_g 7.02146e-19 $X=4.77 $Y=0.805
+ $X2=0 $Y2=0
cc_311 N_A_217_413#_c_266_n N_A_1112_93#_M1010_g 0.00241023f $X=4.825 $Y=1.39
+ $X2=0 $Y2=0
cc_312 N_A_217_413#_c_261_n N_A_1112_93#_M1012_g 0.0027368f $X=5.105 $Y=1.825
+ $X2=0 $Y2=0
cc_313 N_A_217_413#_c_271_n N_A_1112_93#_M1012_g 0.0562535f $X=5.43 $Y=1.9 $X2=0
+ $Y2=0
cc_314 N_A_217_413#_c_261_n N_A_1112_93#_c_708_n 2.34177e-19 $X=5.105 $Y=1.825
+ $X2=0 $Y2=0
cc_315 N_A_217_413#_c_266_n N_A_1112_93#_c_708_n 2.04674e-19 $X=4.825 $Y=1.39
+ $X2=0 $Y2=0
cc_316 N_A_217_413#_c_261_n N_A_1112_93#_c_723_n 4.3326e-19 $X=5.105 $Y=1.825
+ $X2=0 $Y2=0
cc_317 N_A_217_413#_c_271_n N_A_1112_93#_c_723_n 0.00221046f $X=5.43 $Y=1.9
+ $X2=0 $Y2=0
cc_318 N_A_217_413#_c_271_n N_A_1112_93#_c_714_n 0.00131728f $X=5.43 $Y=1.9
+ $X2=0 $Y2=0
cc_319 N_A_217_413#_c_266_n N_A_1112_93#_c_714_n 0.00598403f $X=4.825 $Y=1.39
+ $X2=0 $Y2=0
cc_320 N_A_217_413#_c_298_p N_A_941_379#_M1021_d 0.00967097f $X=4.76 $Y=2.37
+ $X2=0 $Y2=0
cc_321 N_A_217_413#_c_264_n N_A_941_379#_M1021_d 0.00604697f $X=4.845 $Y=2.285
+ $X2=0 $Y2=0
cc_322 N_A_217_413#_M1007_g N_A_941_379#_c_850_n 0.00208291f $X=4.77 $Y=0.805
+ $X2=0 $Y2=0
cc_323 N_A_217_413#_c_265_n N_A_941_379#_c_850_n 0.00200937f $X=4.825 $Y=1.39
+ $X2=0 $Y2=0
cc_324 N_A_217_413#_c_266_n N_A_941_379#_c_850_n 0.00642055f $X=4.825 $Y=1.39
+ $X2=0 $Y2=0
cc_325 N_A_217_413#_M1007_g N_A_941_379#_c_851_n 4.5825e-19 $X=4.77 $Y=0.805
+ $X2=0 $Y2=0
cc_326 N_A_217_413#_c_261_n N_A_941_379#_c_851_n 0.00719655f $X=5.105 $Y=1.825
+ $X2=0 $Y2=0
cc_327 N_A_217_413#_c_271_n N_A_941_379#_c_851_n 0.0129093f $X=5.43 $Y=1.9 $X2=0
+ $Y2=0
cc_328 N_A_217_413#_c_272_n N_A_941_379#_c_851_n 0.0037533f $X=5.18 $Y=1.9 $X2=0
+ $Y2=0
cc_329 N_A_217_413#_M1006_g N_A_941_379#_c_851_n 0.0210015f $X=5.505 $Y=2.415
+ $X2=0 $Y2=0
cc_330 N_A_217_413#_c_298_p N_A_941_379#_c_851_n 0.0136054f $X=4.76 $Y=2.37
+ $X2=0 $Y2=0
cc_331 N_A_217_413#_c_265_n N_A_941_379#_c_851_n 0.0746923f $X=4.825 $Y=1.39
+ $X2=0 $Y2=0
cc_332 N_A_217_413#_c_266_n N_A_941_379#_c_851_n 0.00832869f $X=4.825 $Y=1.39
+ $X2=0 $Y2=0
cc_333 N_A_217_413#_c_271_n N_A_941_379#_c_852_n 0.00478132f $X=5.43 $Y=1.9
+ $X2=0 $Y2=0
cc_334 N_A_217_413#_c_275_n N_VPWR_M1015_d 0.0102533f $X=1.905 $Y=2.13 $X2=0
+ $Y2=0
cc_335 N_A_217_413#_c_276_n N_VPWR_M1015_d 0.00348377f $X=1.99 $Y=2.535 $X2=0
+ $Y2=0
cc_336 N_A_217_413#_c_298_p N_VPWR_M1024_d 0.00722879f $X=4.76 $Y=2.37 $X2=0
+ $Y2=0
cc_337 N_A_217_413#_c_275_n N_VPWR_c_931_n 0.0130182f $X=1.905 $Y=2.13 $X2=0
+ $Y2=0
cc_338 N_A_217_413#_c_276_n N_VPWR_c_931_n 0.00985916f $X=1.99 $Y=2.535 $X2=0
+ $Y2=0
cc_339 N_A_217_413#_c_278_n N_VPWR_c_931_n 0.0136569f $X=2.075 $Y=2.62 $X2=0
+ $Y2=0
cc_340 N_A_217_413#_c_282_n N_VPWR_c_931_n 5.90496e-19 $X=1.21 $Y=2.21 $X2=0
+ $Y2=0
cc_341 N_A_217_413#_c_298_p N_VPWR_c_932_n 0.0250461f $X=4.76 $Y=2.37 $X2=0
+ $Y2=0
cc_342 N_A_217_413#_c_284_n N_VPWR_c_932_n 0.00465758f $X=3.41 $Y=2.37 $X2=0
+ $Y2=0
cc_343 N_A_217_413#_M1006_g N_VPWR_c_939_n 0.00375548f $X=5.505 $Y=2.415 $X2=0
+ $Y2=0
cc_344 N_A_217_413#_c_282_n N_VPWR_c_941_n 0.00565673f $X=1.21 $Y=2.21 $X2=0
+ $Y2=0
cc_345 N_A_217_413#_c_277_n N_VPWR_c_942_n 0.00965489f $X=2.595 $Y=2.62 $X2=0
+ $Y2=0
cc_346 N_A_217_413#_c_278_n N_VPWR_c_942_n 0.00350151f $X=2.075 $Y=2.62 $X2=0
+ $Y2=0
cc_347 N_A_217_413#_c_280_n N_VPWR_c_942_n 0.00995092f $X=3.325 $Y=2.62 $X2=0
+ $Y2=0
cc_348 N_A_217_413#_c_283_n N_VPWR_c_942_n 0.003716f $X=2.685 $Y=2.62 $X2=0
+ $Y2=0
cc_349 N_A_217_413#_c_284_n N_VPWR_c_942_n 0.00333843f $X=3.41 $Y=2.37 $X2=0
+ $Y2=0
cc_350 N_A_217_413#_M1006_g N_VPWR_c_928_n 0.00447875f $X=5.505 $Y=2.415 $X2=0
+ $Y2=0
cc_351 N_A_217_413#_c_277_n N_VPWR_c_928_n 0.0129146f $X=2.595 $Y=2.62 $X2=0
+ $Y2=0
cc_352 N_A_217_413#_c_278_n N_VPWR_c_928_n 0.0045202f $X=2.075 $Y=2.62 $X2=0
+ $Y2=0
cc_353 N_A_217_413#_c_280_n N_VPWR_c_928_n 0.0134921f $X=3.325 $Y=2.62 $X2=0
+ $Y2=0
cc_354 N_A_217_413#_c_282_n N_VPWR_c_928_n 0.00825004f $X=1.21 $Y=2.21 $X2=0
+ $Y2=0
cc_355 N_A_217_413#_c_283_n N_VPWR_c_928_n 0.00479376f $X=2.685 $Y=2.62 $X2=0
+ $Y2=0
cc_356 N_A_217_413#_c_284_n N_VPWR_c_928_n 0.00433963f $X=3.41 $Y=2.37 $X2=0
+ $Y2=0
cc_357 N_A_217_413#_M1008_g N_A_431_119#_c_1047_n 9.42626e-19 $X=2.555 $Y=2.275
+ $X2=0 $Y2=0
cc_358 N_A_217_413#_c_263_n N_A_431_119#_c_1047_n 0.0195783f $X=2.69 $Y=1.71
+ $X2=0 $Y2=0
cc_359 N_A_217_413#_c_275_n N_A_431_119#_c_1048_n 0.00788521f $X=1.905 $Y=2.13
+ $X2=0 $Y2=0
cc_360 N_A_217_413#_c_277_n N_A_431_119#_c_1048_n 0.0135779f $X=2.595 $Y=2.62
+ $X2=0 $Y2=0
cc_361 N_A_217_413#_M1005_g N_A_431_119#_c_1046_n 0.00159792f $X=3.135 $Y=0.805
+ $X2=0 $Y2=0
cc_362 N_A_217_413#_c_263_n N_A_431_119#_c_1046_n 0.0264168f $X=2.69 $Y=1.71
+ $X2=0 $Y2=0
cc_363 N_A_217_413#_c_267_n N_A_431_119#_c_1046_n 0.00312234f $X=2.855 $Y=1.71
+ $X2=0 $Y2=0
cc_364 N_A_217_413#_c_284_n A_666_413# 0.0020218f $X=3.41 $Y=2.37 $X2=-0.19
+ $Y2=-0.245
cc_365 N_A_217_413#_c_336_p N_VGND_c_1143_n 0.00472802f $X=1.325 $Y=0.805 $X2=0
+ $Y2=0
cc_366 N_A_217_413#_M1005_g N_VGND_c_1151_n 9.39239e-19 $X=3.135 $Y=0.805 $X2=0
+ $Y2=0
cc_367 N_A_217_413#_M1007_g N_VGND_c_1151_n 9.39239e-19 $X=4.77 $Y=0.805 $X2=0
+ $Y2=0
cc_368 N_A_217_413#_c_336_p N_VGND_c_1151_n 0.00825355f $X=1.325 $Y=0.805 $X2=0
+ $Y2=0
cc_369 N_A_684_93#_M1024_g N_A_526_413#_M1003_g 0.0246286f $X=3.615 $Y=2.275
+ $X2=0 $Y2=0
cc_370 N_A_684_93#_c_431_n N_A_526_413#_M1003_g 0.00150266f $X=3.585 $Y=1.53
+ $X2=0 $Y2=0
cc_371 N_A_684_93#_c_427_n N_A_526_413#_M1003_g 5.9872e-19 $X=3.585 $Y=1.53
+ $X2=0 $Y2=0
cc_372 N_A_684_93#_c_433_n N_A_526_413#_M1003_g 0.0142623f $X=4.39 $Y=1.985
+ $X2=0 $Y2=0
cc_373 N_A_684_93#_c_428_n N_A_526_413#_M1003_g 0.00329392f $X=4.475 $Y=1.855
+ $X2=0 $Y2=0
cc_374 N_A_684_93#_M1024_g N_A_526_413#_c_496_n 9.74239e-19 $X=3.615 $Y=2.275
+ $X2=0 $Y2=0
cc_375 N_A_684_93#_c_431_n N_A_526_413#_c_496_n 0.0214371f $X=3.585 $Y=1.53
+ $X2=0 $Y2=0
cc_376 N_A_684_93#_c_427_n N_A_526_413#_c_496_n 8.98363e-19 $X=3.585 $Y=1.53
+ $X2=0 $Y2=0
cc_377 N_A_684_93#_c_434_n N_A_526_413#_c_496_n 0.0143458f $X=3.75 $Y=1.985
+ $X2=0 $Y2=0
cc_378 N_A_684_93#_M1001_g N_A_526_413#_c_497_n 0.0155105f $X=3.495 $Y=0.805
+ $X2=0 $Y2=0
cc_379 N_A_684_93#_c_431_n N_A_526_413#_c_497_n 0.0256226f $X=3.585 $Y=1.53
+ $X2=0 $Y2=0
cc_380 N_A_684_93#_c_427_n N_A_526_413#_c_497_n 0.00496611f $X=3.585 $Y=1.53
+ $X2=0 $Y2=0
cc_381 N_A_684_93#_c_433_n N_A_526_413#_c_497_n 0.00693547f $X=4.39 $Y=1.985
+ $X2=0 $Y2=0
cc_382 N_A_684_93#_c_428_n N_A_526_413#_c_497_n 0.0134141f $X=4.475 $Y=1.855
+ $X2=0 $Y2=0
cc_383 N_A_684_93#_M1001_g N_A_526_413#_c_498_n 0.00145132f $X=3.495 $Y=0.805
+ $X2=0 $Y2=0
cc_384 N_A_684_93#_c_431_n N_A_526_413#_c_498_n 0.0143145f $X=3.585 $Y=1.53
+ $X2=0 $Y2=0
cc_385 N_A_684_93#_c_427_n N_A_526_413#_c_498_n 0.00137486f $X=3.585 $Y=1.53
+ $X2=0 $Y2=0
cc_386 N_A_684_93#_c_433_n N_A_526_413#_c_498_n 0.019714f $X=4.39 $Y=1.985 $X2=0
+ $Y2=0
cc_387 N_A_684_93#_c_428_n N_A_526_413#_c_498_n 0.0294488f $X=4.475 $Y=1.855
+ $X2=0 $Y2=0
cc_388 N_A_684_93#_M1001_g N_A_526_413#_c_499_n 6.66966e-19 $X=3.495 $Y=0.805
+ $X2=0 $Y2=0
cc_389 N_A_684_93#_c_431_n N_A_526_413#_c_499_n 8.05543e-19 $X=3.585 $Y=1.53
+ $X2=0 $Y2=0
cc_390 N_A_684_93#_c_427_n N_A_526_413#_c_499_n 0.0194714f $X=3.585 $Y=1.53
+ $X2=0 $Y2=0
cc_391 N_A_684_93#_c_433_n N_A_526_413#_c_499_n 0.00225044f $X=4.39 $Y=1.985
+ $X2=0 $Y2=0
cc_392 N_A_684_93#_M1001_g N_A_526_413#_c_500_n 9.84651e-19 $X=3.495 $Y=0.805
+ $X2=0 $Y2=0
cc_393 N_A_684_93#_M1001_g N_A_526_413#_c_501_n 0.0132918f $X=3.495 $Y=0.805
+ $X2=0 $Y2=0
cc_394 N_A_684_93#_c_428_n N_A_526_413#_c_501_n 0.010517f $X=4.475 $Y=1.855
+ $X2=0 $Y2=0
cc_395 N_A_684_93#_c_429_n N_A_526_413#_c_501_n 0.00475773f $X=4.455 $Y=0.77
+ $X2=0 $Y2=0
cc_396 N_A_684_93#_M1001_g N_A_110_70#_c_574_n 0.0104164f $X=3.495 $Y=0.805
+ $X2=0 $Y2=0
cc_397 N_A_684_93#_c_429_n N_A_110_70#_c_574_n 0.00516589f $X=4.455 $Y=0.77
+ $X2=0 $Y2=0
cc_398 N_A_684_93#_M1024_g N_A_110_70#_M1022_g 0.0412556f $X=3.615 $Y=2.275
+ $X2=0 $Y2=0
cc_399 N_A_684_93#_c_434_n N_A_110_70#_M1022_g 0.00154303f $X=3.75 $Y=1.985
+ $X2=0 $Y2=0
cc_400 N_A_684_93#_M1024_g N_A_110_70#_c_586_n 0.00391504f $X=3.615 $Y=2.275
+ $X2=0 $Y2=0
cc_401 N_A_684_93#_c_428_n N_A_110_70#_M1021_g 0.00579595f $X=4.475 $Y=1.855
+ $X2=0 $Y2=0
cc_402 N_A_684_93#_c_428_n N_A_941_379#_c_850_n 0.00675366f $X=4.475 $Y=1.855
+ $X2=0 $Y2=0
cc_403 N_A_684_93#_c_428_n N_A_941_379#_c_851_n 0.00134528f $X=4.475 $Y=1.855
+ $X2=0 $Y2=0
cc_404 N_A_684_93#_c_433_n N_VPWR_M1024_d 0.00433164f $X=4.39 $Y=1.985 $X2=0
+ $Y2=0
cc_405 N_A_684_93#_M1024_g N_VPWR_c_928_n 9.7053e-19 $X=3.615 $Y=2.275 $X2=0
+ $Y2=0
cc_406 N_A_684_93#_c_434_n A_666_413# 0.00120338f $X=3.75 $Y=1.985 $X2=-0.19
+ $Y2=-0.245
cc_407 N_A_684_93#_M1001_g N_VGND_c_1134_n 0.00934084f $X=3.495 $Y=0.805 $X2=0
+ $Y2=0
cc_408 N_A_684_93#_c_429_n N_VGND_c_1134_n 0.0196363f $X=4.455 $Y=0.77 $X2=0
+ $Y2=0
cc_409 N_A_684_93#_c_429_n N_VGND_c_1144_n 0.00590721f $X=4.455 $Y=0.77 $X2=0
+ $Y2=0
cc_410 N_A_684_93#_M1001_g N_VGND_c_1151_n 9.39239e-19 $X=3.495 $Y=0.805 $X2=0
+ $Y2=0
cc_411 N_A_684_93#_c_429_n N_VGND_c_1151_n 0.00727686f $X=4.455 $Y=0.77 $X2=0
+ $Y2=0
cc_412 N_A_526_413#_c_495_n N_A_110_70#_M1000_g 0.00358963f $X=2.885 $Y=0.805
+ $X2=0 $Y2=0
cc_413 N_A_526_413#_c_495_n N_A_110_70#_c_574_n 0.0050195f $X=2.885 $Y=0.805
+ $X2=0 $Y2=0
cc_414 N_A_526_413#_c_501_n N_A_110_70#_c_574_n 0.0103738f $X=4.13 $Y=1.345
+ $X2=0 $Y2=0
cc_415 N_A_526_413#_c_496_n N_A_110_70#_M1022_g 0.00159443f $X=3.03 $Y=2.19
+ $X2=0 $Y2=0
cc_416 N_A_526_413#_c_497_n N_A_110_70#_M1022_g 0.00311047f $X=3.96 $Y=1.19
+ $X2=0 $Y2=0
cc_417 N_A_526_413#_M1003_g N_A_110_70#_c_586_n 0.0100858f $X=4.2 $Y=2.315 $X2=0
+ $Y2=0
cc_418 N_A_526_413#_M1003_g N_A_110_70#_M1021_g 0.0360516f $X=4.2 $Y=2.315 $X2=0
+ $Y2=0
cc_419 N_A_526_413#_M1003_g N_VPWR_c_932_n 0.00771933f $X=4.2 $Y=2.315 $X2=0
+ $Y2=0
cc_420 N_A_526_413#_M1003_g N_VPWR_c_928_n 9.39239e-19 $X=4.2 $Y=2.315 $X2=0
+ $Y2=0
cc_421 N_A_526_413#_c_495_n N_A_431_119#_c_1046_n 0.0192974f $X=2.885 $Y=0.805
+ $X2=0 $Y2=0
cc_422 N_A_526_413#_c_496_n N_A_431_119#_c_1046_n 0.00674484f $X=3.03 $Y=2.19
+ $X2=0 $Y2=0
cc_423 N_A_526_413#_c_497_n N_VGND_M1001_d 0.00447087f $X=3.96 $Y=1.19 $X2=0
+ $Y2=0
cc_424 N_A_526_413#_c_497_n N_VGND_c_1134_n 0.0274538f $X=3.96 $Y=1.19 $X2=0
+ $Y2=0
cc_425 N_A_526_413#_c_499_n N_VGND_c_1134_n 3.3741e-19 $X=4.125 $Y=1.51 $X2=0
+ $Y2=0
cc_426 N_A_526_413#_c_501_n N_VGND_c_1134_n 0.00724078f $X=4.13 $Y=1.345 $X2=0
+ $Y2=0
cc_427 N_A_526_413#_c_495_n N_VGND_c_1141_n 0.00563533f $X=2.885 $Y=0.805 $X2=0
+ $Y2=0
cc_428 N_A_526_413#_c_495_n N_VGND_c_1151_n 0.00864182f $X=2.885 $Y=0.805 $X2=0
+ $Y2=0
cc_429 N_A_526_413#_c_501_n N_VGND_c_1151_n 9.39239e-19 $X=4.13 $Y=1.345 $X2=0
+ $Y2=0
cc_430 N_A_110_70#_M1017_g N_A_1112_93#_M1010_g 0.0412772f $X=5.275 $Y=0.805
+ $X2=0 $Y2=0
cc_431 N_A_110_70#_c_574_n N_A_941_379#_c_850_n 0.00393009f $X=5.2 $Y=0.18 $X2=0
+ $Y2=0
cc_432 N_A_110_70#_M1017_g N_A_941_379#_c_850_n 0.020545f $X=5.275 $Y=0.805
+ $X2=0 $Y2=0
cc_433 N_A_110_70#_M1021_g N_A_941_379#_c_851_n 0.00811873f $X=4.63 $Y=2.315
+ $X2=0 $Y2=0
cc_434 N_A_110_70#_c_589_n N_VPWR_c_930_n 0.0125559f $X=0.69 $Y=2.485 $X2=0
+ $Y2=0
cc_435 N_A_110_70#_M1015_g N_VPWR_c_931_n 0.0146817f $X=1.425 $Y=2.385 $X2=0
+ $Y2=0
cc_436 N_A_110_70#_c_583_n N_VPWR_c_931_n 0.0162871f $X=3.18 $Y=3.15 $X2=0 $Y2=0
cc_437 N_A_110_70#_M1022_g N_VPWR_c_932_n 0.0108186f $X=3.255 $Y=2.275 $X2=0
+ $Y2=0
cc_438 N_A_110_70#_c_586_n N_VPWR_c_932_n 0.0253901f $X=4.555 $Y=3.15 $X2=0
+ $Y2=0
cc_439 N_A_110_70#_M1021_g N_VPWR_c_932_n 0.00616623f $X=4.63 $Y=2.315 $X2=0
+ $Y2=0
cc_440 N_A_110_70#_c_586_n N_VPWR_c_939_n 0.0225642f $X=4.555 $Y=3.15 $X2=0
+ $Y2=0
cc_441 N_A_110_70#_c_584_n N_VPWR_c_941_n 0.00718072f $X=1.5 $Y=3.15 $X2=0 $Y2=0
cc_442 N_A_110_70#_c_589_n N_VPWR_c_941_n 0.0119929f $X=0.69 $Y=2.485 $X2=0
+ $Y2=0
cc_443 N_A_110_70#_c_583_n N_VPWR_c_942_n 0.0558531f $X=3.18 $Y=3.15 $X2=0 $Y2=0
cc_444 N_A_110_70#_c_583_n N_VPWR_c_928_n 0.0456536f $X=3.18 $Y=3.15 $X2=0 $Y2=0
cc_445 N_A_110_70#_c_584_n N_VPWR_c_928_n 0.0114291f $X=1.5 $Y=3.15 $X2=0 $Y2=0
cc_446 N_A_110_70#_c_586_n N_VPWR_c_928_n 0.0497629f $X=4.555 $Y=3.15 $X2=0
+ $Y2=0
cc_447 N_A_110_70#_c_588_n N_VPWR_c_928_n 0.0042224f $X=3.255 $Y=3.15 $X2=0
+ $Y2=0
cc_448 N_A_110_70#_c_589_n N_VPWR_c_928_n 0.00958569f $X=0.69 $Y=2.485 $X2=0
+ $Y2=0
cc_449 N_A_110_70#_c_571_n N_A_431_119#_c_1051_n 0.00432573f $X=2.535 $Y=0.18
+ $X2=0 $Y2=0
cc_450 N_A_110_70#_M1000_g N_A_431_119#_c_1051_n 0.00384091f $X=2.61 $Y=0.805
+ $X2=0 $Y2=0
cc_451 N_A_110_70#_M1000_g N_A_431_119#_c_1046_n 0.0015453f $X=2.61 $Y=0.805
+ $X2=0 $Y2=0
cc_452 N_A_110_70#_M1011_g N_VGND_c_1133_n 0.0148841f $X=1.54 $Y=0.805 $X2=0
+ $Y2=0
cc_453 N_A_110_70#_c_571_n N_VGND_c_1133_n 0.0241992f $X=2.535 $Y=0.18 $X2=0
+ $Y2=0
cc_454 N_A_110_70#_M1000_g N_VGND_c_1133_n 0.00548981f $X=2.61 $Y=0.805 $X2=0
+ $Y2=0
cc_455 N_A_110_70#_c_574_n N_VGND_c_1134_n 0.0260329f $X=5.2 $Y=0.18 $X2=0 $Y2=0
cc_456 N_A_110_70#_c_574_n N_VGND_c_1135_n 0.00954179f $X=5.2 $Y=0.18 $X2=0
+ $Y2=0
cc_457 N_A_110_70#_c_571_n N_VGND_c_1141_n 0.0550093f $X=2.535 $Y=0.18 $X2=0
+ $Y2=0
cc_458 N_A_110_70#_c_572_n N_VGND_c_1143_n 0.00703166f $X=1.615 $Y=0.18 $X2=0
+ $Y2=0
cc_459 N_A_110_70#_c_578_n N_VGND_c_1143_n 0.00930971f $X=0.69 $Y=0.56 $X2=0
+ $Y2=0
cc_460 N_A_110_70#_c_574_n N_VGND_c_1144_n 0.0401726f $X=5.2 $Y=0.18 $X2=0 $Y2=0
cc_461 N_A_110_70#_c_571_n N_VGND_c_1151_n 0.0201867f $X=2.535 $Y=0.18 $X2=0
+ $Y2=0
cc_462 N_A_110_70#_c_572_n N_VGND_c_1151_n 0.0109674f $X=1.615 $Y=0.18 $X2=0
+ $Y2=0
cc_463 N_A_110_70#_c_574_n N_VGND_c_1151_n 0.0900349f $X=5.2 $Y=0.18 $X2=0 $Y2=0
cc_464 N_A_110_70#_c_577_n N_VGND_c_1151_n 0.00880231f $X=2.61 $Y=0.18 $X2=0
+ $Y2=0
cc_465 N_A_110_70#_c_578_n N_VGND_c_1151_n 0.00926582f $X=0.69 $Y=0.56 $X2=0
+ $Y2=0
cc_466 N_A_1112_93#_c_708_n N_A_941_379#_M1028_g 9.50988e-19 $X=5.725 $Y=1.45
+ $X2=0 $Y2=0
cc_467 N_A_1112_93#_c_722_n N_A_941_379#_M1028_g 0.0148544f $X=6.51 $Y=1.78
+ $X2=0 $Y2=0
cc_468 N_A_1112_93#_c_709_n N_A_941_379#_M1028_g 0.00532036f $X=6.63 $Y=1.865
+ $X2=0 $Y2=0
cc_469 N_A_1112_93#_c_725_n N_A_941_379#_M1028_g 0.00412549f $X=6.605 $Y=1.87
+ $X2=0 $Y2=0
cc_470 N_A_1112_93#_c_713_n N_A_941_379#_M1028_g 0.00252445f $X=7.265 $Y=1.48
+ $X2=0 $Y2=0
cc_471 N_A_1112_93#_c_714_n N_A_941_379#_M1028_g 0.0232797f $X=5.865 $Y=1.45
+ $X2=0 $Y2=0
cc_472 N_A_1112_93#_M1010_g N_A_941_379#_c_850_n 0.00160737f $X=5.635 $Y=0.805
+ $X2=0 $Y2=0
cc_473 N_A_1112_93#_M1010_g N_A_941_379#_c_851_n 0.00632635f $X=5.635 $Y=0.805
+ $X2=0 $Y2=0
cc_474 N_A_1112_93#_M1012_g N_A_941_379#_c_851_n 0.00102382f $X=5.865 $Y=2.415
+ $X2=0 $Y2=0
cc_475 N_A_1112_93#_c_708_n N_A_941_379#_c_851_n 0.0236047f $X=5.725 $Y=1.45
+ $X2=0 $Y2=0
cc_476 N_A_1112_93#_c_723_n N_A_941_379#_c_851_n 0.0127992f $X=5.89 $Y=1.78
+ $X2=0 $Y2=0
cc_477 N_A_1112_93#_M1026_d N_A_941_379#_c_852_n 0.00123568f $X=6.3 $Y=0.235
+ $X2=0 $Y2=0
cc_478 N_A_1112_93#_M1010_g N_A_941_379#_c_852_n 0.0153473f $X=5.635 $Y=0.805
+ $X2=0 $Y2=0
cc_479 N_A_1112_93#_c_708_n N_A_941_379#_c_852_n 0.025062f $X=5.725 $Y=1.45
+ $X2=0 $Y2=0
cc_480 N_A_1112_93#_c_722_n N_A_941_379#_c_852_n 0.00892364f $X=6.51 $Y=1.78
+ $X2=0 $Y2=0
cc_481 N_A_1112_93#_c_710_n N_A_941_379#_c_852_n 0.0141714f $X=6.665 $Y=1.395
+ $X2=0 $Y2=0
cc_482 N_A_1112_93#_c_712_n N_A_941_379#_c_852_n 0.00489107f $X=6.46 $Y=0.39
+ $X2=0 $Y2=0
cc_483 N_A_1112_93#_c_714_n N_A_941_379#_c_852_n 0.00645478f $X=5.865 $Y=1.45
+ $X2=0 $Y2=0
cc_484 N_A_1112_93#_M1010_g N_A_941_379#_c_853_n 5.54372e-19 $X=5.635 $Y=0.805
+ $X2=0 $Y2=0
cc_485 N_A_1112_93#_c_708_n N_A_941_379#_c_853_n 0.00839748f $X=5.725 $Y=1.45
+ $X2=0 $Y2=0
cc_486 N_A_1112_93#_c_722_n N_A_941_379#_c_853_n 0.0189119f $X=6.51 $Y=1.78
+ $X2=0 $Y2=0
cc_487 N_A_1112_93#_c_709_n N_A_941_379#_c_853_n 0.00995671f $X=6.63 $Y=1.865
+ $X2=0 $Y2=0
cc_488 N_A_1112_93#_c_710_n N_A_941_379#_c_853_n 0.015425f $X=6.665 $Y=1.395
+ $X2=0 $Y2=0
cc_489 N_A_1112_93#_c_714_n N_A_941_379#_c_853_n 0.00110243f $X=5.865 $Y=1.45
+ $X2=0 $Y2=0
cc_490 N_A_1112_93#_c_708_n N_A_941_379#_c_854_n 5.17151e-19 $X=5.725 $Y=1.45
+ $X2=0 $Y2=0
cc_491 N_A_1112_93#_c_722_n N_A_941_379#_c_854_n 0.00168569f $X=6.51 $Y=1.78
+ $X2=0 $Y2=0
cc_492 N_A_1112_93#_c_709_n N_A_941_379#_c_854_n 0.00124336f $X=6.63 $Y=1.865
+ $X2=0 $Y2=0
cc_493 N_A_1112_93#_c_710_n N_A_941_379#_c_854_n 0.00391264f $X=6.665 $Y=1.395
+ $X2=0 $Y2=0
cc_494 N_A_1112_93#_c_712_n N_A_941_379#_c_854_n 0.00313877f $X=6.46 $Y=0.39
+ $X2=0 $Y2=0
cc_495 N_A_1112_93#_c_713_n N_A_941_379#_c_854_n 0.00432716f $X=7.265 $Y=1.48
+ $X2=0 $Y2=0
cc_496 N_A_1112_93#_c_714_n N_A_941_379#_c_854_n 0.0147235f $X=5.865 $Y=1.45
+ $X2=0 $Y2=0
cc_497 N_A_1112_93#_M1010_g N_A_941_379#_c_855_n 0.0194781f $X=5.635 $Y=0.805
+ $X2=0 $Y2=0
cc_498 N_A_1112_93#_c_710_n N_A_941_379#_c_855_n 0.0044191f $X=6.665 $Y=1.395
+ $X2=0 $Y2=0
cc_499 N_A_1112_93#_c_712_n N_A_941_379#_c_855_n 0.00521075f $X=6.46 $Y=0.39
+ $X2=0 $Y2=0
cc_500 N_A_1112_93#_c_722_n N_VPWR_M1012_d 0.00232649f $X=6.51 $Y=1.78 $X2=0
+ $Y2=0
cc_501 N_A_1112_93#_M1012_g N_VPWR_c_933_n 0.0115147f $X=5.865 $Y=2.415 $X2=0
+ $Y2=0
cc_502 N_A_1112_93#_c_722_n N_VPWR_c_933_n 0.0220026f $X=6.51 $Y=1.78 $X2=0
+ $Y2=0
cc_503 N_A_1112_93#_c_725_n N_VPWR_c_933_n 0.03715f $X=6.605 $Y=1.87 $X2=0 $Y2=0
cc_504 N_A_1112_93#_c_725_n N_VPWR_c_934_n 0.0118006f $X=6.605 $Y=1.87 $X2=0
+ $Y2=0
cc_505 N_A_1112_93#_M1002_g N_VPWR_c_935_n 0.00768161f $X=7.34 $Y=2.465 $X2=0
+ $Y2=0
cc_506 N_A_1112_93#_c_709_n N_VPWR_c_935_n 0.0037807f $X=6.63 $Y=1.865 $X2=0
+ $Y2=0
cc_507 N_A_1112_93#_c_725_n N_VPWR_c_935_n 0.0792111f $X=6.605 $Y=1.87 $X2=0
+ $Y2=0
cc_508 N_A_1112_93#_c_711_n N_VPWR_c_935_n 0.0177424f $X=8.45 $Y=1.48 $X2=0
+ $Y2=0
cc_509 N_A_1112_93#_c_713_n N_VPWR_c_935_n 0.0072038f $X=7.265 $Y=1.48 $X2=0
+ $Y2=0
cc_510 N_A_1112_93#_M1002_g N_VPWR_c_936_n 7.47048e-19 $X=7.34 $Y=2.465 $X2=0
+ $Y2=0
cc_511 N_A_1112_93#_M1009_g N_VPWR_c_936_n 0.0148627f $X=7.77 $Y=2.465 $X2=0
+ $Y2=0
cc_512 N_A_1112_93#_M1018_g N_VPWR_c_936_n 0.0147822f $X=8.2 $Y=2.465 $X2=0
+ $Y2=0
cc_513 N_A_1112_93#_M1025_g N_VPWR_c_936_n 7.32829e-19 $X=8.63 $Y=2.465 $X2=0
+ $Y2=0
cc_514 N_A_1112_93#_M1018_g N_VPWR_c_938_n 5.67328e-19 $X=8.2 $Y=2.465 $X2=0
+ $Y2=0
cc_515 N_A_1112_93#_M1025_g N_VPWR_c_938_n 0.0125837f $X=8.63 $Y=2.465 $X2=0
+ $Y2=0
cc_516 N_A_1112_93#_M1012_g N_VPWR_c_939_n 0.00375548f $X=5.865 $Y=2.415 $X2=0
+ $Y2=0
cc_517 N_A_1112_93#_M1002_g N_VPWR_c_943_n 0.00585385f $X=7.34 $Y=2.465 $X2=0
+ $Y2=0
cc_518 N_A_1112_93#_M1009_g N_VPWR_c_943_n 0.00486043f $X=7.77 $Y=2.465 $X2=0
+ $Y2=0
cc_519 N_A_1112_93#_M1018_g N_VPWR_c_944_n 0.00486043f $X=8.2 $Y=2.465 $X2=0
+ $Y2=0
cc_520 N_A_1112_93#_M1025_g N_VPWR_c_944_n 0.00486043f $X=8.63 $Y=2.465 $X2=0
+ $Y2=0
cc_521 N_A_1112_93#_M1012_g N_VPWR_c_928_n 0.00447875f $X=5.865 $Y=2.415 $X2=0
+ $Y2=0
cc_522 N_A_1112_93#_M1002_g N_VPWR_c_928_n 0.0118221f $X=7.34 $Y=2.465 $X2=0
+ $Y2=0
cc_523 N_A_1112_93#_M1009_g N_VPWR_c_928_n 0.00824727f $X=7.77 $Y=2.465 $X2=0
+ $Y2=0
cc_524 N_A_1112_93#_M1018_g N_VPWR_c_928_n 0.00824727f $X=8.2 $Y=2.465 $X2=0
+ $Y2=0
cc_525 N_A_1112_93#_M1025_g N_VPWR_c_928_n 0.00824727f $X=8.63 $Y=2.465 $X2=0
+ $Y2=0
cc_526 N_A_1112_93#_c_725_n N_VPWR_c_928_n 0.00892005f $X=6.605 $Y=1.87 $X2=0
+ $Y2=0
cc_527 N_A_1112_93#_M1013_g N_Q_c_1071_n 0.00254528f $X=7.34 $Y=0.655 $X2=0
+ $Y2=0
cc_528 N_A_1112_93#_c_710_n N_Q_c_1071_n 0.00414334f $X=6.665 $Y=1.395 $X2=0
+ $Y2=0
cc_529 N_A_1112_93#_c_711_n N_Q_c_1071_n 0.0185589f $X=8.45 $Y=1.48 $X2=0 $Y2=0
cc_530 N_A_1112_93#_c_715_n N_Q_c_1071_n 0.00256759f $X=8.63 $Y=1.48 $X2=0 $Y2=0
cc_531 N_A_1112_93#_M1009_g N_Q_c_1075_n 0.013253f $X=7.77 $Y=2.465 $X2=0 $Y2=0
cc_532 N_A_1112_93#_M1018_g N_Q_c_1075_n 0.0134064f $X=8.2 $Y=2.465 $X2=0 $Y2=0
cc_533 N_A_1112_93#_c_711_n N_Q_c_1075_n 0.0467265f $X=8.45 $Y=1.48 $X2=0 $Y2=0
cc_534 N_A_1112_93#_c_715_n N_Q_c_1075_n 0.00246472f $X=8.63 $Y=1.48 $X2=0 $Y2=0
cc_535 N_A_1112_93#_M1002_g N_Q_c_1076_n 0.00162204f $X=7.34 $Y=2.465 $X2=0
+ $Y2=0
cc_536 N_A_1112_93#_c_709_n N_Q_c_1076_n 0.00280662f $X=6.63 $Y=1.865 $X2=0
+ $Y2=0
cc_537 N_A_1112_93#_c_711_n N_Q_c_1076_n 0.0181554f $X=8.45 $Y=1.48 $X2=0 $Y2=0
cc_538 N_A_1112_93#_c_715_n N_Q_c_1076_n 0.00256759f $X=8.63 $Y=1.48 $X2=0 $Y2=0
cc_539 N_A_1112_93#_c_711_n N_Q_c_1077_n 0.0153308f $X=8.45 $Y=1.48 $X2=0 $Y2=0
cc_540 N_A_1112_93#_c_715_n N_Q_c_1077_n 0.00256759f $X=8.63 $Y=1.48 $X2=0 $Y2=0
cc_541 N_A_1112_93#_M1025_g Q 0.018142f $X=8.63 $Y=2.465 $X2=0 $Y2=0
cc_542 N_A_1112_93#_c_711_n Q 0.00736973f $X=8.45 $Y=1.48 $X2=0 $Y2=0
cc_543 N_A_1112_93#_M1025_g Q 0.0124658f $X=8.63 $Y=2.465 $X2=0 $Y2=0
cc_544 N_A_1112_93#_M1029_g Q 0.0194571f $X=8.63 $Y=0.655 $X2=0 $Y2=0
cc_545 N_A_1112_93#_c_711_n Q 0.0131807f $X=8.45 $Y=1.48 $X2=0 $Y2=0
cc_546 N_A_1112_93#_M1014_g N_Q_c_1073_n 0.0137655f $X=7.77 $Y=0.655 $X2=0 $Y2=0
cc_547 N_A_1112_93#_M1020_g N_Q_c_1073_n 0.0140083f $X=8.2 $Y=0.655 $X2=0 $Y2=0
cc_548 N_A_1112_93#_c_711_n N_Q_c_1073_n 0.0690414f $X=8.45 $Y=1.48 $X2=0 $Y2=0
cc_549 N_A_1112_93#_c_715_n N_Q_c_1073_n 0.00246472f $X=8.63 $Y=1.48 $X2=0 $Y2=0
cc_550 N_A_1112_93#_M1029_g N_Q_c_1074_n 0.0217121f $X=8.63 $Y=0.655 $X2=0 $Y2=0
cc_551 N_A_1112_93#_c_715_n N_Q_c_1074_n 0.00251812f $X=8.63 $Y=1.48 $X2=0 $Y2=0
cc_552 N_A_1112_93#_M1010_g N_VGND_c_1135_n 0.00780896f $X=5.635 $Y=0.805 $X2=0
+ $Y2=0
cc_553 N_A_1112_93#_c_712_n N_VGND_c_1136_n 0.0250466f $X=6.46 $Y=0.39 $X2=0
+ $Y2=0
cc_554 N_A_1112_93#_M1013_g N_VGND_c_1137_n 0.00702716f $X=7.34 $Y=0.655 $X2=0
+ $Y2=0
cc_555 N_A_1112_93#_c_711_n N_VGND_c_1137_n 0.0152469f $X=8.45 $Y=1.48 $X2=0
+ $Y2=0
cc_556 N_A_1112_93#_c_712_n N_VGND_c_1137_n 0.0577107f $X=6.46 $Y=0.39 $X2=0
+ $Y2=0
cc_557 N_A_1112_93#_c_713_n N_VGND_c_1137_n 0.00686121f $X=7.265 $Y=1.48 $X2=0
+ $Y2=0
cc_558 N_A_1112_93#_M1013_g N_VGND_c_1138_n 6.44378e-19 $X=7.34 $Y=0.655 $X2=0
+ $Y2=0
cc_559 N_A_1112_93#_M1014_g N_VGND_c_1138_n 0.011376f $X=7.77 $Y=0.655 $X2=0
+ $Y2=0
cc_560 N_A_1112_93#_M1020_g N_VGND_c_1138_n 0.0112752f $X=8.2 $Y=0.655 $X2=0
+ $Y2=0
cc_561 N_A_1112_93#_M1029_g N_VGND_c_1138_n 6.18138e-19 $X=8.63 $Y=0.655 $X2=0
+ $Y2=0
cc_562 N_A_1112_93#_M1020_g N_VGND_c_1140_n 5.67328e-19 $X=8.2 $Y=0.655 $X2=0
+ $Y2=0
cc_563 N_A_1112_93#_M1029_g N_VGND_c_1140_n 0.0118244f $X=8.63 $Y=0.655 $X2=0
+ $Y2=0
cc_564 N_A_1112_93#_M1010_g N_VGND_c_1144_n 0.00431487f $X=5.635 $Y=0.805 $X2=0
+ $Y2=0
cc_565 N_A_1112_93#_M1013_g N_VGND_c_1145_n 0.00585385f $X=7.34 $Y=0.655 $X2=0
+ $Y2=0
cc_566 N_A_1112_93#_M1014_g N_VGND_c_1145_n 0.00486043f $X=7.77 $Y=0.655 $X2=0
+ $Y2=0
cc_567 N_A_1112_93#_M1020_g N_VGND_c_1146_n 0.00486043f $X=8.2 $Y=0.655 $X2=0
+ $Y2=0
cc_568 N_A_1112_93#_M1029_g N_VGND_c_1146_n 0.00486043f $X=8.63 $Y=0.655 $X2=0
+ $Y2=0
cc_569 N_A_1112_93#_M1026_d N_VGND_c_1151_n 0.00233241f $X=6.3 $Y=0.235 $X2=0
+ $Y2=0
cc_570 N_A_1112_93#_M1010_g N_VGND_c_1151_n 0.00477801f $X=5.635 $Y=0.805 $X2=0
+ $Y2=0
cc_571 N_A_1112_93#_M1013_g N_VGND_c_1151_n 0.0118358f $X=7.34 $Y=0.655 $X2=0
+ $Y2=0
cc_572 N_A_1112_93#_M1014_g N_VGND_c_1151_n 0.00824727f $X=7.77 $Y=0.655 $X2=0
+ $Y2=0
cc_573 N_A_1112_93#_M1020_g N_VGND_c_1151_n 0.00824727f $X=8.2 $Y=0.655 $X2=0
+ $Y2=0
cc_574 N_A_1112_93#_M1029_g N_VGND_c_1151_n 0.00454119f $X=8.63 $Y=0.655 $X2=0
+ $Y2=0
cc_575 N_A_1112_93#_c_712_n N_VGND_c_1151_n 0.0172024f $X=6.46 $Y=0.39 $X2=0
+ $Y2=0
cc_576 N_A_941_379#_M1028_g N_VPWR_c_933_n 0.0159049f $X=6.39 $Y=2.355 $X2=0
+ $Y2=0
cc_577 N_A_941_379#_c_851_n N_VPWR_c_933_n 0.0195971f $X=5.195 $Y=2.195 $X2=0
+ $Y2=0
cc_578 N_A_941_379#_M1028_g N_VPWR_c_934_n 0.00400407f $X=6.39 $Y=2.355 $X2=0
+ $Y2=0
cc_579 N_A_941_379#_M1028_g N_VPWR_c_935_n 0.0035114f $X=6.39 $Y=2.355 $X2=0
+ $Y2=0
cc_580 N_A_941_379#_c_851_n N_VPWR_c_939_n 0.00487078f $X=5.195 $Y=2.195 $X2=0
+ $Y2=0
cc_581 N_A_941_379#_M1028_g N_VPWR_c_928_n 0.00804497f $X=6.39 $Y=2.355 $X2=0
+ $Y2=0
cc_582 N_A_941_379#_c_851_n N_VPWR_c_928_n 0.00755367f $X=5.195 $Y=2.195 $X2=0
+ $Y2=0
cc_583 N_A_941_379#_c_852_n N_VGND_M1010_d 0.00311014f $X=6.15 $Y=1.1 $X2=0
+ $Y2=0
cc_584 N_A_941_379#_c_850_n N_VGND_c_1135_n 0.0069029f $X=5.235 $Y=1.185 $X2=0
+ $Y2=0
cc_585 N_A_941_379#_c_852_n N_VGND_c_1135_n 0.025029f $X=6.15 $Y=1.1 $X2=0 $Y2=0
cc_586 N_A_941_379#_c_855_n N_VGND_c_1135_n 0.0116717f $X=6.315 $Y=1.185 $X2=0
+ $Y2=0
cc_587 N_A_941_379#_c_855_n N_VGND_c_1136_n 0.00579478f $X=6.315 $Y=1.185 $X2=0
+ $Y2=0
cc_588 N_A_941_379#_c_855_n N_VGND_c_1137_n 0.00207168f $X=6.315 $Y=1.185 $X2=0
+ $Y2=0
cc_589 N_A_941_379#_c_850_n N_VGND_c_1144_n 0.00644329f $X=5.235 $Y=1.185 $X2=0
+ $Y2=0
cc_590 N_A_941_379#_c_850_n N_VGND_c_1151_n 0.00980982f $X=5.235 $Y=1.185 $X2=0
+ $Y2=0
cc_591 N_A_941_379#_c_855_n N_VGND_c_1151_n 0.013259f $X=6.315 $Y=1.185 $X2=0
+ $Y2=0
cc_592 N_A_941_379#_c_850_n A_1070_119# 4.51105e-19 $X=5.235 $Y=1.185 $X2=-0.19
+ $Y2=-0.245
cc_593 N_VPWR_c_928_n N_Q_M1002_s 0.0041489f $X=8.88 $Y=3.33 $X2=0 $Y2=0
cc_594 N_VPWR_c_928_n N_Q_M1018_s 0.00536646f $X=8.88 $Y=3.33 $X2=0 $Y2=0
cc_595 N_VPWR_c_943_n N_Q_c_1108_n 0.0136943f $X=7.82 $Y=3.33 $X2=0 $Y2=0
cc_596 N_VPWR_c_928_n N_Q_c_1108_n 0.00866972f $X=8.88 $Y=3.33 $X2=0 $Y2=0
cc_597 N_VPWR_M1009_d N_Q_c_1075_n 0.00176461f $X=7.845 $Y=1.835 $X2=0 $Y2=0
cc_598 N_VPWR_c_936_n N_Q_c_1075_n 0.0170777f $X=7.985 $Y=2.16 $X2=0 $Y2=0
cc_599 N_VPWR_c_935_n N_Q_c_1076_n 0.00166618f $X=7.125 $Y=1.98 $X2=0 $Y2=0
cc_600 N_VPWR_c_944_n N_Q_c_1113_n 0.0124525f $X=8.68 $Y=3.33 $X2=0 $Y2=0
cc_601 N_VPWR_c_928_n N_Q_c_1113_n 0.00730901f $X=8.88 $Y=3.33 $X2=0 $Y2=0
cc_602 N_VPWR_M1025_d Q 0.00177014f $X=8.705 $Y=1.835 $X2=0 $Y2=0
cc_603 N_VPWR_M1025_d Q 0.0109009f $X=8.705 $Y=1.835 $X2=0 $Y2=0
cc_604 N_VPWR_c_938_n Q 0.0188763f $X=8.845 $Y=2.795 $X2=0 $Y2=0
cc_605 N_VPWR_c_928_n Q 0.00176098f $X=8.88 $Y=3.33 $X2=0 $Y2=0
cc_606 N_A_431_119#_c_1051_n N_VGND_c_1141_n 0.0057866f $X=2.385 $Y=0.79 $X2=0
+ $Y2=0
cc_607 N_A_431_119#_c_1051_n N_VGND_c_1151_n 0.0085359f $X=2.385 $Y=0.79 $X2=0
+ $Y2=0
cc_608 N_Q_c_1073_n N_VGND_M1014_s 0.00176461f $X=8.32 $Y=1.032 $X2=0 $Y2=0
cc_609 N_Q_c_1074_n N_VGND_M1029_s 0.00333756f $X=8.915 $Y=1.032 $X2=0 $Y2=0
cc_610 N_Q_c_1071_n N_VGND_c_1137_n 0.00166417f $X=7.65 $Y=1.14 $X2=0 $Y2=0
cc_611 N_Q_c_1073_n N_VGND_c_1138_n 0.0170777f $X=8.32 $Y=1.032 $X2=0 $Y2=0
cc_612 N_Q_c_1074_n N_VGND_c_1140_n 0.0227469f $X=8.915 $Y=1.032 $X2=0 $Y2=0
cc_613 N_Q_c_1124_p N_VGND_c_1145_n 0.0138717f $X=7.555 $Y=0.42 $X2=0 $Y2=0
cc_614 N_Q_c_1125_p N_VGND_c_1146_n 0.0123249f $X=8.415 $Y=0.42 $X2=0 $Y2=0
cc_615 N_Q_M1013_d N_VGND_c_1151_n 0.00397496f $X=7.415 $Y=0.235 $X2=0 $Y2=0
cc_616 N_Q_M1020_d N_VGND_c_1151_n 0.00405668f $X=8.275 $Y=0.235 $X2=0 $Y2=0
cc_617 N_Q_c_1124_p N_VGND_c_1151_n 0.00886411f $X=7.555 $Y=0.42 $X2=0 $Y2=0
cc_618 N_Q_c_1125_p N_VGND_c_1151_n 0.00728036f $X=8.415 $Y=0.42 $X2=0 $Y2=0
cc_619 N_Q_c_1074_n N_VGND_c_1151_n 0.00752816f $X=8.915 $Y=1.032 $X2=0 $Y2=0
