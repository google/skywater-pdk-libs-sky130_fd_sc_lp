* File: sky130_fd_sc_lp__o41ai_lp.pex.spice
* Created: Fri Aug 28 11:20:43 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O41AI_LP%B1 3 7 11 12 13 14 18 19
r36 18 19 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.63
+ $Y=1.29 $X2=0.63 $Y2=1.29
r37 13 14 11.8446 $w=3.58e-07 $l=3.7e-07 $layer=LI1_cond $X=0.645 $Y=1.295
+ $X2=0.645 $Y2=1.665
r38 13 19 0.160062 $w=3.58e-07 $l=5e-09 $layer=LI1_cond $X=0.645 $Y=1.295
+ $X2=0.645 $Y2=1.29
r39 11 18 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.63 $Y=1.63
+ $X2=0.63 $Y2=1.29
r40 11 12 30.8683 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.63 $Y=1.63
+ $X2=0.63 $Y2=1.795
r41 10 18 41.8716 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.63 $Y=1.125
+ $X2=0.63 $Y2=1.29
r42 7 10 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=0.69 $Y=0.495
+ $X2=0.69 $Y2=1.125
r43 3 12 198.763 $w=2.5e-07 $l=8e-07 $layer=POLY_cond $X=0.64 $Y=2.595 $X2=0.64
+ $Y2=1.795
.ends

.subckt PM_SKY130_FD_SC_LP__O41AI_LP%A4 3 5 7 11 12 13 17
r46 12 13 13.0959 $w=3.28e-07 $l=3.75e-07 $layer=LI1_cond $X=1.17 $Y=1.29
+ $X2=1.17 $Y2=1.665
r47 12 17 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.17
+ $Y=1.29 $X2=1.17 $Y2=1.29
r48 11 17 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.17 $Y=1.63
+ $X2=1.17 $Y2=1.29
r49 10 17 40.8701 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.17 $Y=1.125
+ $X2=1.17 $Y2=1.29
r50 5 11 30.6163 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.17 $Y=1.795
+ $X2=1.17 $Y2=1.63
r51 5 7 198.763 $w=2.5e-07 $l=8e-07 $layer=POLY_cond $X=1.17 $Y=1.795 $X2=1.17
+ $Y2=2.595
r52 3 10 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=1.12 $Y=0.495
+ $X2=1.12 $Y2=1.125
.ends

.subckt PM_SKY130_FD_SC_LP__O41AI_LP%A3 3 7 11 12 13 14 15 16 22 23
r49 22 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.71
+ $Y=1.43 $X2=1.71 $Y2=1.43
r50 15 16 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.71 $Y=2.405
+ $X2=1.71 $Y2=2.775
r51 14 15 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.71 $Y=2.035
+ $X2=1.71 $Y2=2.405
r52 13 14 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.71 $Y=1.665
+ $X2=1.71 $Y2=2.035
r53 13 23 8.20679 $w=3.28e-07 $l=2.35e-07 $layer=LI1_cond $X=1.71 $Y=1.665
+ $X2=1.71 $Y2=1.43
r54 11 22 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.71 $Y=1.77
+ $X2=1.71 $Y2=1.43
r55 11 12 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.71 $Y=1.77
+ $X2=1.71 $Y2=1.935
r56 10 22 40.8701 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.71 $Y=1.265
+ $X2=1.71 $Y2=1.43
r57 7 10 394.83 $w=1.5e-07 $l=7.7e-07 $layer=POLY_cond $X=1.76 $Y=0.495 $X2=1.76
+ $Y2=1.265
r58 3 12 163.979 $w=2.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.67 $Y=2.595
+ $X2=1.67 $Y2=1.935
.ends

.subckt PM_SKY130_FD_SC_LP__O41AI_LP%A2 3 7 11 12 13 14 15 16 22 23
c45 3 0 1.75272e-19 $X=2.19 $Y=0.495
r46 22 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.28
+ $Y=1.43 $X2=2.28 $Y2=1.43
r47 15 16 10.9334 $w=3.88e-07 $l=3.7e-07 $layer=LI1_cond $X=2.25 $Y=2.405
+ $X2=2.25 $Y2=2.775
r48 14 15 10.9334 $w=3.88e-07 $l=3.7e-07 $layer=LI1_cond $X=2.25 $Y=2.035
+ $X2=2.25 $Y2=2.405
r49 13 14 10.9334 $w=3.88e-07 $l=3.7e-07 $layer=LI1_cond $X=2.25 $Y=1.665
+ $X2=2.25 $Y2=2.035
r50 13 23 6.94421 $w=3.88e-07 $l=2.35e-07 $layer=LI1_cond $X=2.25 $Y=1.665
+ $X2=2.25 $Y2=1.43
r51 11 22 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.28 $Y=1.77
+ $X2=2.28 $Y2=1.43
r52 11 12 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.28 $Y=1.77
+ $X2=2.28 $Y2=1.935
r53 10 22 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.28 $Y=1.265
+ $X2=2.28 $Y2=1.43
r54 7 12 163.979 $w=2.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.24 $Y=2.595
+ $X2=2.24 $Y2=1.935
r55 3 10 394.83 $w=1.5e-07 $l=7.7e-07 $layer=POLY_cond $X=2.19 $Y=0.495 $X2=2.19
+ $Y2=1.265
.ends

.subckt PM_SKY130_FD_SC_LP__O41AI_LP%A1 3 7 9 12
c29 9 0 1.75272e-19 $X=3.12 $Y=1.665
r30 12 15 72.9334 $w=4.55e-07 $l=5.05e-07 $layer=POLY_cond $X=2.912 $Y=1.39
+ $X2=2.912 $Y2=1.895
r31 12 14 47.0767 $w=4.55e-07 $l=1.65e-07 $layer=POLY_cond $X=2.912 $Y=1.39
+ $X2=2.912 $Y2=1.225
r32 12 13 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.975
+ $Y=1.39 $X2=2.975 $Y2=1.39
r33 9 13 2.58853 $w=6.68e-07 $l=1.45e-07 $layer=LI1_cond $X=3.12 $Y=1.56
+ $X2=2.975 $Y2=1.56
r34 7 14 374.319 $w=1.5e-07 $l=7.3e-07 $layer=POLY_cond $X=2.78 $Y=0.495
+ $X2=2.78 $Y2=1.225
r35 3 15 173.918 $w=2.5e-07 $l=7e-07 $layer=POLY_cond $X=2.81 $Y=2.595 $X2=2.81
+ $Y2=1.895
.ends

.subckt PM_SKY130_FD_SC_LP__O41AI_LP%VPWR 1 2 7 9 11 13 17 19 32
r39 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r40 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r41 26 32 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r42 25 26 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r43 23 29 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r44 22 25 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=0.72 $Y=3.33
+ $X2=2.64 $Y2=3.33
r45 22 23 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r46 20 28 4.55841 $w=1.7e-07 $l=2.7e-07 $layer=LI1_cond $X=0.54 $Y=3.33 $X2=0.27
+ $Y2=3.33
r47 20 22 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=0.54 $Y=3.33
+ $X2=0.72 $Y2=3.33
r48 19 31 4.72267 $w=1.7e-07 $l=2.25e-07 $layer=LI1_cond $X=2.91 $Y=3.33
+ $X2=3.135 $Y2=3.33
r49 19 25 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=2.91 $Y=3.33 $X2=2.64
+ $Y2=3.33
r50 17 26 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r51 17 23 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.72 $Y2=3.33
r52 13 16 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=3.075 $Y=2.24
+ $X2=3.075 $Y2=2.95
r53 11 31 3.0435 $w=3.3e-07 $l=1.11018e-07 $layer=LI1_cond $X=3.075 $Y=3.245
+ $X2=3.135 $Y2=3.33
r54 11 16 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=3.075 $Y=3.245
+ $X2=3.075 $Y2=2.95
r55 7 28 3.20777 $w=3.3e-07 $l=1.41244e-07 $layer=LI1_cond $X=0.375 $Y=3.245
+ $X2=0.27 $Y2=3.33
r56 7 9 26.3665 $w=3.28e-07 $l=7.55e-07 $layer=LI1_cond $X=0.375 $Y=3.245
+ $X2=0.375 $Y2=2.49
r57 2 16 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=2.935
+ $Y=2.095 $X2=3.075 $Y2=2.95
r58 2 13 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.935
+ $Y=2.095 $X2=3.075 $Y2=2.24
r59 1 9 300 $w=1.7e-07 $l=4.61844e-07 $layer=licon1_PDIFF $count=2 $X=0.23
+ $Y=2.095 $X2=0.375 $Y2=2.49
.ends

.subckt PM_SKY130_FD_SC_LP__O41AI_LP%Y 1 2 8 9 10 13 15 18
r37 15 22 8.99073 $w=4.43e-07 $l=1.7e-07 $layer=LI1_cond $X=0.337 $Y=0.555
+ $X2=0.337 $Y2=0.725
r38 15 18 1.55386 $w=4.43e-07 $l=6e-08 $layer=LI1_cond $X=0.337 $Y=0.555
+ $X2=0.337 $Y2=0.495
r39 11 13 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=0.905 $Y=2.145
+ $X2=0.905 $Y2=2.24
r40 9 11 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.74 $Y=2.06
+ $X2=0.905 $Y2=2.145
r41 9 10 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=0.74 $Y=2.06
+ $X2=0.285 $Y2=2.06
r42 8 10 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.2 $Y=1.975
+ $X2=0.285 $Y2=2.06
r43 8 22 81.5508 $w=1.68e-07 $l=1.25e-06 $layer=LI1_cond $X=0.2 $Y=1.975 $X2=0.2
+ $Y2=0.725
r44 2 13 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=0.765
+ $Y=2.095 $X2=0.905 $Y2=2.24
r45 1 18 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.25
+ $Y=0.285 $X2=0.395 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__O41AI_LP%A_153_57# 1 2 3 12 14 15 18 20 24 26
r57 22 24 13.2706 $w=3.28e-07 $l=3.8e-07 $layer=LI1_cond $X=2.995 $Y=0.875
+ $X2=2.995 $Y2=0.495
r58 21 26 8.61065 $w=1.7e-07 $l=1.88348e-07 $layer=LI1_cond $X=2.14 $Y=0.96
+ $X2=1.975 $Y2=0.91
r59 20 22 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.83 $Y=0.96
+ $X2=2.995 $Y2=0.875
r60 20 21 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.83 $Y=0.96 $X2=2.14
+ $Y2=0.96
r61 16 26 0.89609 $w=3.3e-07 $l=1.35e-07 $layer=LI1_cond $X=1.975 $Y=0.775
+ $X2=1.975 $Y2=0.91
r62 16 18 9.7783 $w=3.28e-07 $l=2.8e-07 $layer=LI1_cond $X=1.975 $Y=0.775
+ $X2=1.975 $Y2=0.495
r63 14 26 8.61065 $w=1.7e-07 $l=1.88348e-07 $layer=LI1_cond $X=1.81 $Y=0.86
+ $X2=1.975 $Y2=0.91
r64 14 15 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=1.81 $Y=0.86
+ $X2=1.07 $Y2=0.86
r65 10 15 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.905 $Y=0.775
+ $X2=1.07 $Y2=0.86
r66 10 12 9.7783 $w=3.28e-07 $l=2.8e-07 $layer=LI1_cond $X=0.905 $Y=0.775
+ $X2=0.905 $Y2=0.495
r67 3 24 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.855
+ $Y=0.285 $X2=2.995 $Y2=0.495
r68 2 18 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.835
+ $Y=0.285 $X2=1.975 $Y2=0.495
r69 1 12 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.765
+ $Y=0.285 $X2=0.905 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__O41AI_LP%VGND 1 2 9 13 16 17 19 20 21 34 35
r37 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r38 32 35 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r39 31 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r40 28 29 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r41 25 29 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r42 24 28 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r43 24 25 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r44 21 32 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r45 21 29 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r46 19 31 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=2.32 $Y=0 $X2=2.16
+ $Y2=0
r47 19 20 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.32 $Y=0 $X2=2.485
+ $Y2=0
r48 18 34 30.6631 $w=1.68e-07 $l=4.7e-07 $layer=LI1_cond $X=2.65 $Y=0 $X2=3.12
+ $Y2=0
r49 18 20 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.65 $Y=0 $X2=2.485
+ $Y2=0
r50 16 28 3.26203 $w=1.68e-07 $l=5e-08 $layer=LI1_cond $X=1.25 $Y=0 $X2=1.2
+ $Y2=0
r51 16 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.25 $Y=0 $X2=1.415
+ $Y2=0
r52 15 31 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=1.58 $Y=0 $X2=2.16
+ $Y2=0
r53 15 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.58 $Y=0 $X2=1.415
+ $Y2=0
r54 11 20 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.485 $Y=0.085
+ $X2=2.485 $Y2=0
r55 11 13 13.7944 $w=3.28e-07 $l=3.95e-07 $layer=LI1_cond $X=2.485 $Y=0.085
+ $X2=2.485 $Y2=0.48
r56 7 17 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.415 $Y=0.085
+ $X2=1.415 $Y2=0
r57 7 9 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=1.415 $Y=0.085
+ $X2=1.415 $Y2=0.43
r58 2 13 182 $w=1.7e-07 $l=3.02159e-07 $layer=licon1_NDIFF $count=1 $X=2.265
+ $Y=0.285 $X2=2.485 $Y2=0.48
r59 1 9 182 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_NDIFF $count=1 $X=1.195
+ $Y=0.285 $X2=1.415 $Y2=0.43
.ends

