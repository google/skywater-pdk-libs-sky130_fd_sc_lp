* File: sky130_fd_sc_lp__dlrtn_lp.pex.spice
* Created: Fri Aug 28 10:26:49 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__DLRTN_LP%D 1 3 7 10 12 14 16 17 18 19 20 24 25 26
c44 25 0 1.96767e-19 $X=0.625 $Y=1.275
c45 10 0 6.50813e-20 $X=0.665 $Y=2.575
r46 24 26 46.7569 $w=3.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.605 $Y=1.275
+ $X2=0.605 $Y2=1.11
r47 24 25 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.625
+ $Y=1.275 $X2=0.625 $Y2=1.275
r48 19 20 11.3708 $w=3.73e-07 $l=3.7e-07 $layer=LI1_cond $X=0.647 $Y=1.295
+ $X2=0.647 $Y2=1.665
r49 19 25 0.614636 $w=3.73e-07 $l=2e-08 $layer=LI1_cond $X=0.647 $Y=1.295
+ $X2=0.647 $Y2=1.275
r50 14 16 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.855 $Y=0.73
+ $X2=0.855 $Y2=0.445
r51 13 17 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.57 $Y=0.805
+ $X2=0.495 $Y2=0.805
r52 12 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.78 $Y=0.805
+ $X2=0.855 $Y2=0.73
r53 12 13 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=0.78 $Y=0.805
+ $X2=0.57 $Y2=0.805
r54 10 18 197.521 $w=2.5e-07 $l=7.95e-07 $layer=POLY_cond $X=0.665 $Y=2.575
+ $X2=0.665 $Y2=1.78
r55 7 18 34.9505 $w=3.7e-07 $l=1.85e-07 $layer=POLY_cond $X=0.605 $Y=1.595
+ $X2=0.605 $Y2=1.78
r56 6 24 3.11915 $w=3.7e-07 $l=2e-08 $layer=POLY_cond $X=0.605 $Y=1.295
+ $X2=0.605 $Y2=1.275
r57 6 7 46.7872 $w=3.7e-07 $l=3e-07 $layer=POLY_cond $X=0.605 $Y=1.295 $X2=0.605
+ $Y2=1.595
r58 4 17 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.495 $Y=0.88
+ $X2=0.495 $Y2=0.805
r59 4 26 117.936 $w=1.5e-07 $l=2.3e-07 $layer=POLY_cond $X=0.495 $Y=0.88
+ $X2=0.495 $Y2=1.11
r60 1 17 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.495 $Y=0.73
+ $X2=0.495 $Y2=0.805
r61 1 3 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.495 $Y=0.73 $X2=0.495
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__DLRTN_LP%GATE_N 1 3 7 9 13 16 18 19 23
c53 18 0 6.50813e-20 $X=1.2 $Y=1.295
c54 7 0 1.96767e-19 $X=1.285 $Y=0.445
r55 18 19 13.2706 $w=3.28e-07 $l=3.8e-07 $layer=LI1_cond $X=1.195 $Y=1.285
+ $X2=1.195 $Y2=1.665
r56 18 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.195
+ $Y=1.285 $X2=1.195 $Y2=1.285
r57 17 23 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.195 $Y=1.625
+ $X2=1.195 $Y2=1.285
r58 15 23 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=1.195 $Y=1.27
+ $X2=1.195 $Y2=1.285
r59 15 16 13.5877 $w=2.4e-07 $l=7.5e-08 $layer=POLY_cond $X=1.195 $Y=1.27
+ $X2=1.195 $Y2=1.195
r60 11 13 346.117 $w=1.5e-07 $l=6.75e-07 $layer=POLY_cond $X=1.675 $Y=1.12
+ $X2=1.675 $Y2=0.445
r61 10 16 12.1617 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.36 $Y=1.195
+ $X2=1.195 $Y2=1.195
r62 9 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.6 $Y=1.195
+ $X2=1.675 $Y2=1.12
r63 9 10 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=1.6 $Y=1.195 $X2=1.36
+ $Y2=1.195
r64 5 16 13.5877 $w=2.4e-07 $l=1.21861e-07 $layer=POLY_cond $X=1.285 $Y=1.12
+ $X2=1.195 $Y2=1.195
r65 5 7 346.117 $w=1.5e-07 $l=6.75e-07 $layer=POLY_cond $X=1.285 $Y=1.12
+ $X2=1.285 $Y2=0.445
r66 1 17 30.6163 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.195 $Y=1.79
+ $X2=1.195 $Y2=1.625
r67 1 3 195.036 $w=2.5e-07 $l=7.85e-07 $layer=POLY_cond $X=1.195 $Y=1.79
+ $X2=1.195 $Y2=2.575
.ends

.subckt PM_SKY130_FD_SC_LP__DLRTN_LP%A_264_415# 1 2 7 11 13 14 17 19 23 27 30 31
+ 33 35 40 47 54 55 60 62
c134 31 0 1.26497e-19 $X=4.38 $Y=1.825
c135 30 0 1.06304e-19 $X=4.055 $Y=1.675
r136 55 70 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.965 $Y=1.18
+ $X2=3.965 $Y2=1.345
r137 55 69 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.965 $Y=1.18
+ $X2=3.965 $Y2=1.015
r138 54 55 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.965
+ $Y=1.18 $X2=3.965 $Y2=1.18
r139 50 54 47.4946 $w=3.28e-07 $l=1.36e-06 $layer=LI1_cond $X=2.605 $Y=1.18
+ $X2=3.965 $Y2=1.18
r140 50 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.605
+ $Y=1.18 $X2=2.605 $Y2=1.18
r141 48 62 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=1.735 $Y=1.75
+ $X2=1.735 $Y2=1.66
r142 47 48 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.735
+ $Y=1.75 $X2=1.735 $Y2=1.75
r143 45 47 11.5244 $w=3.03e-07 $l=3.05e-07 $layer=LI1_cond $X=1.722 $Y=2.055
+ $X2=1.722 $Y2=1.75
r144 44 60 9.8067 $w=1.88e-07 $l=1.68e-07 $layer=LI1_cond $X=1.722 $Y=0.39
+ $X2=1.89 $Y2=0.39
r145 44 47 47.798 $w=3.03e-07 $l=1.265e-06 $layer=LI1_cond $X=1.722 $Y=0.485
+ $X2=1.722 $Y2=1.75
r146 40 45 6.87288 $w=2.6e-07 $l=2.07036e-07 $layer=LI1_cond $X=1.57 $Y=2.185
+ $X2=1.722 $Y2=2.055
r147 40 42 4.87572 $w=2.58e-07 $l=1.1e-07 $layer=LI1_cond $X=1.57 $Y=2.185
+ $X2=1.46 $Y2=2.185
r148 31 36 166.649 $w=1.5e-07 $l=3.25e-07 $layer=POLY_cond $X=4.38 $Y=1.75
+ $X2=4.055 $Y2=1.75
r149 31 33 186.34 $w=2.5e-07 $l=7.5e-07 $layer=POLY_cond $X=4.38 $Y=1.825
+ $X2=4.38 $Y2=2.575
r150 30 36 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.055 $Y=1.675
+ $X2=4.055 $Y2=1.75
r151 30 70 169.213 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=4.055 $Y=1.675
+ $X2=4.055 $Y2=1.345
r152 27 69 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=3.875 $Y=0.445
+ $X2=3.875 $Y2=1.015
r153 21 23 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=3.055 $Y=0.805
+ $X2=3.055 $Y2=0.445
r154 20 51 48.8514 $w=2.96e-07 $l=3.85357e-07 $layer=POLY_cond $X=2.77 $Y=0.88
+ $X2=2.575 $Y2=1.18
r155 19 21 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.98 $Y=0.88
+ $X2=3.055 $Y2=0.805
r156 19 20 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=2.98 $Y=0.88
+ $X2=2.77 $Y2=0.88
r157 15 20 23.9164 $w=2.96e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.695 $Y=0.805
+ $X2=2.77 $Y2=0.88
r158 15 17 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=2.695 $Y=0.805
+ $X2=2.695 $Y2=0.445
r159 14 35 15.9654 $w=2e-07 $l=9.68246e-08 $layer=POLY_cond $X=2.455 $Y=1.585
+ $X2=2.405 $Y2=1.66
r160 13 51 38.5718 $w=2.96e-07 $l=2.16852e-07 $layer=POLY_cond $X=2.455 $Y=1.345
+ $X2=2.575 $Y2=1.18
r161 13 14 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=2.455 $Y=1.345
+ $X2=2.455 $Y2=1.585
r162 9 35 15.9654 $w=2e-07 $l=7.5e-08 $layer=POLY_cond $X=2.405 $Y=1.735
+ $X2=2.405 $Y2=1.66
r163 9 11 208.701 $w=2.5e-07 $l=8.4e-07 $layer=POLY_cond $X=2.405 $Y=1.735
+ $X2=2.405 $Y2=2.575
r164 8 62 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.9 $Y=1.66
+ $X2=1.735 $Y2=1.66
r165 7 35 9.46703 $w=1.5e-07 $l=1.25e-07 $layer=POLY_cond $X=2.28 $Y=1.66
+ $X2=2.405 $Y2=1.66
r166 7 8 194.851 $w=1.5e-07 $l=3.8e-07 $layer=POLY_cond $X=2.28 $Y=1.66 $X2=1.9
+ $Y2=1.66
r167 2 42 600 $w=1.7e-07 $l=2.08567e-07 $layer=licon1_PDIFF $count=1 $X=1.32
+ $Y=2.075 $X2=1.46 $Y2=2.225
r168 1 60 182 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=1 $X=1.75
+ $Y=0.235 $X2=1.89 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_LP__DLRTN_LP%A_27_47# 1 2 9 13 14 17 21 23 26 27 29 30
+ 33 37 38 43 48
c93 30 0 6.88529e-20 $X=3.065 $Y=1.75
r94 43 45 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.36 $Y=2.58
+ $X2=1.36 $Y2=2.75
r95 39 41 8.41198 $w=4.53e-07 $l=3.2e-07 $layer=LI1_cond $X=0.337 $Y=2.58
+ $X2=0.337 $Y2=2.9
r96 37 39 9.46348 $w=4.53e-07 $l=3.6e-07 $layer=LI1_cond $X=0.337 $Y=2.22
+ $X2=0.337 $Y2=2.58
r97 37 38 9.25191 $w=4.53e-07 $l=1.65e-07 $layer=LI1_cond $X=0.337 $Y=2.22
+ $X2=0.337 $Y2=2.055
r98 35 38 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=0.195 $Y=0.675
+ $X2=0.195 $Y2=2.055
r99 33 35 9.84219 $w=3.33e-07 $l=2.05e-07 $layer=LI1_cond $X=0.277 $Y=0.47
+ $X2=0.277 $Y2=0.675
r100 30 49 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.065 $Y=1.75
+ $X2=3.065 $Y2=1.915
r101 30 48 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.065 $Y=1.75
+ $X2=3.065 $Y2=1.585
r102 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.065
+ $Y=1.75 $X2=3.065 $Y2=1.75
r103 27 29 17.112 $w=3.28e-07 $l=4.9e-07 $layer=LI1_cond $X=2.575 $Y=1.75
+ $X2=3.065 $Y2=1.75
r104 25 27 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.49 $Y=1.915
+ $X2=2.575 $Y2=1.75
r105 25 26 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=2.49 $Y=1.915
+ $X2=2.49 $Y2=2.665
r106 24 45 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.445 $Y=2.75
+ $X2=1.36 $Y2=2.75
r107 23 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.405 $Y=2.75
+ $X2=2.49 $Y2=2.665
r108 23 24 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.405 $Y=2.75
+ $X2=1.445 $Y2=2.75
r109 22 39 6.56868 $w=1.7e-07 $l=2.28e-07 $layer=LI1_cond $X=0.565 $Y=2.58
+ $X2=0.337 $Y2=2.58
r110 21 43 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.275 $Y=2.58
+ $X2=1.36 $Y2=2.58
r111 21 22 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=1.275 $Y=2.58
+ $X2=0.565 $Y2=2.58
r112 15 17 384.574 $w=1.5e-07 $l=7.5e-07 $layer=POLY_cond $X=3.485 $Y=1.195
+ $X2=3.485 $Y2=0.445
r113 13 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.41 $Y=1.27
+ $X2=3.485 $Y2=1.195
r114 13 14 92.2979 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=3.41 $Y=1.27
+ $X2=3.23 $Y2=1.27
r115 11 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.155 $Y=1.345
+ $X2=3.23 $Y2=1.27
r116 11 48 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=3.155 $Y=1.345
+ $X2=3.155 $Y2=1.585
r117 9 49 163.979 $w=2.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.105 $Y=2.575
+ $X2=3.105 $Y2=1.915
r118 2 41 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=0.255
+ $Y=2.075 $X2=0.4 $Y2=2.9
r119 2 37 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.255
+ $Y=2.075 $X2=0.4 $Y2=2.22
r120 1 33 182 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.28 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_LP__DLRTN_LP%A_399_415# 1 2 9 13 15 18 22 24 25 26 31 32
+ 34 38 42 44
c113 44 0 1.26497e-19 $X=4.477 $Y=1.435
c114 38 0 1.06304e-19 $X=3.605 $Y=1.67
c115 32 0 6.90166e-20 $X=4.505 $Y=0.93
c116 18 0 6.88529e-20 $X=2.14 $Y=2.27
r117 42 49 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.605 $Y=1.75
+ $X2=3.605 $Y2=1.915
r118 41 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.605
+ $Y=1.75 $X2=3.605 $Y2=1.75
r119 38 41 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=3.605 $Y=1.67
+ $X2=3.605 $Y2=1.75
r120 34 44 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=4.395 $Y=1.585
+ $X2=4.395 $Y2=1.435
r121 31 32 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.505
+ $Y=0.93 $X2=4.505 $Y2=0.93
r122 29 44 8.53494 $w=3.33e-07 $l=1.67e-07 $layer=LI1_cond $X=4.477 $Y=1.268
+ $X2=4.477 $Y2=1.435
r123 29 31 11.6276 $w=3.33e-07 $l=3.38e-07 $layer=LI1_cond $X=4.477 $Y=1.268
+ $X2=4.477 $Y2=0.93
r124 28 31 3.26812 $w=3.33e-07 $l=9.5e-08 $layer=LI1_cond $X=4.477 $Y=0.835
+ $X2=4.477 $Y2=0.93
r125 27 38 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.77 $Y=1.67
+ $X2=3.605 $Y2=1.67
r126 26 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.31 $Y=1.67
+ $X2=4.395 $Y2=1.585
r127 26 27 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=4.31 $Y=1.67
+ $X2=3.77 $Y2=1.67
r128 24 28 7.80856 $w=1.7e-07 $l=2.05144e-07 $layer=LI1_cond $X=4.31 $Y=0.75
+ $X2=4.477 $Y2=0.835
r129 24 25 108.626 $w=1.68e-07 $l=1.665e-06 $layer=LI1_cond $X=4.31 $Y=0.75
+ $X2=2.645 $Y2=0.75
r130 20 25 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=2.48 $Y=0.75
+ $X2=2.645 $Y2=0.75
r131 20 35 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=2.48 $Y=0.75
+ $X2=2.14 $Y2=0.75
r132 20 22 6.80989 $w=3.28e-07 $l=1.95e-07 $layer=LI1_cond $X=2.48 $Y=0.665
+ $X2=2.48 $Y2=0.47
r133 16 35 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.14 $Y=0.835
+ $X2=2.14 $Y2=0.75
r134 16 18 93.6203 $w=1.68e-07 $l=1.435e-06 $layer=LI1_cond $X=2.14 $Y=0.835
+ $X2=2.14 $Y2=2.27
r135 15 32 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.505 $Y=0.765
+ $X2=4.505 $Y2=0.93
r136 13 15 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=4.415 $Y=0.445
+ $X2=4.415 $Y2=0.765
r137 9 49 163.979 $w=2.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.595 $Y=2.575
+ $X2=3.595 $Y2=1.915
r138 2 18 600 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_PDIFF $count=1 $X=1.995
+ $Y=2.075 $X2=2.14 $Y2=2.27
r139 1 22 182 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_NDIFF $count=1 $X=2.335
+ $Y=0.235 $X2=2.48 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_LP__DLRTN_LP%A_949_335# 1 2 9 13 19 23 27 29 30 32 37 40
+ 43 45 47 49 50 51 53 54 56 59 65 66
r135 64 65 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.875
+ $Y=1.02 $X2=6.875 $Y2=1.02
r136 58 59 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.34
+ $Y=1.02 $X2=5.34 $Y2=1.02
r137 56 66 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=6.765 $Y=2.055
+ $X2=6.765 $Y2=1.525
r138 54 66 8.99121 $w=3.58e-07 $l=1.8e-07 $layer=LI1_cond $X=6.86 $Y=1.345
+ $X2=6.86 $Y2=1.525
r139 53 64 2.57345 $w=3.6e-07 $l=8.5e-08 $layer=LI1_cond $X=6.86 $Y=1.025
+ $X2=6.86 $Y2=0.94
r140 53 54 10.2439 $w=3.58e-07 $l=3.2e-07 $layer=LI1_cond $X=6.86 $Y=1.025
+ $X2=6.86 $Y2=1.345
r141 52 62 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.195 $Y=2.14
+ $X2=6.03 $Y2=2.14
r142 51 56 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.68 $Y=2.14
+ $X2=6.765 $Y2=2.055
r143 51 52 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=6.68 $Y=2.14
+ $X2=6.195 $Y2=2.14
r144 49 64 5.44966 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=6.68 $Y=0.94
+ $X2=6.86 $Y2=0.94
r145 49 50 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=6.68 $Y=0.94
+ $X2=5.985 $Y2=0.94
r146 45 62 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.03 $Y=2.225
+ $X2=6.03 $Y2=2.14
r147 45 47 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=6.03 $Y=2.225
+ $X2=6.03 $Y2=2.9
r148 41 50 9.52 $w=2.35e-07 $l=2.0106e-07 $layer=LI1_cond $X=5.82 $Y=1.02
+ $X2=5.985 $Y2=0.94
r149 41 58 24.9191 $w=2.35e-07 $l=4.8e-07 $layer=LI1_cond $X=5.82 $Y=1.02
+ $X2=5.34 $Y2=1.02
r150 41 43 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=5.82 $Y=0.855
+ $X2=5.82 $Y2=0.495
r151 39 65 55.6971 $w=3.45e-07 $l=3.33e-07 $layer=POLY_cond $X=6.882 $Y=1.353
+ $X2=6.882 $Y2=1.02
r152 39 40 33.2433 $w=3.45e-07 $l=1.72e-07 $layer=POLY_cond $X=6.882 $Y=1.353
+ $X2=6.882 $Y2=1.525
r153 36 65 2.50888 $w=3.45e-07 $l=1.5e-08 $layer=POLY_cond $X=6.882 $Y=1.005
+ $X2=6.882 $Y2=1.02
r154 36 37 155.368 $w=1.5e-07 $l=3.03e-07 $layer=POLY_cond $X=6.882 $Y=0.93
+ $X2=7.185 $Y2=0.93
r155 33 36 29.2277 $w=1.5e-07 $l=5.7e-08 $layer=POLY_cond $X=6.825 $Y=0.93
+ $X2=6.882 $Y2=0.93
r156 31 59 48.9612 $w=3.3e-07 $l=2.8e-07 $layer=POLY_cond $X=5.06 $Y=1.02
+ $X2=5.34 $Y2=1.02
r157 31 32 5.03009 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=5.06 $Y=1.02
+ $X2=4.985 $Y2=1.02
r158 29 30 47.1291 $w=2.5e-07 $l=1.5e-07 $layer=POLY_cond $X=4.902 $Y=1.675
+ $X2=4.902 $Y2=1.825
r159 25 37 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.185 $Y=0.855
+ $X2=7.185 $Y2=0.93
r160 25 27 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=7.185 $Y=0.855
+ $X2=7.185 $Y2=0.495
r161 23 40 260.876 $w=2.5e-07 $l=1.05e-06 $layer=POLY_cond $X=6.93 $Y=2.575
+ $X2=6.93 $Y2=1.525
r162 17 33 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.825 $Y=0.855
+ $X2=6.825 $Y2=0.93
r163 17 19 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=6.825 $Y=0.855
+ $X2=6.825 $Y2=0.495
r164 15 32 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.985 $Y=1.185
+ $X2=4.985 $Y2=1.02
r165 15 29 251.255 $w=1.5e-07 $l=4.9e-07 $layer=POLY_cond $X=4.985 $Y=1.185
+ $X2=4.985 $Y2=1.675
r166 11 32 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.985 $Y=0.855
+ $X2=4.985 $Y2=1.02
r167 11 13 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=4.985 $Y=0.855
+ $X2=4.985 $Y2=0.445
r168 9 30 186.34 $w=2.5e-07 $l=7.5e-07 $layer=POLY_cond $X=4.87 $Y=2.575
+ $X2=4.87 $Y2=1.825
r169 2 62 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=5.89
+ $Y=2.075 $X2=6.03 $Y2=2.22
r170 2 47 400 $w=1.7e-07 $l=8.92258e-07 $layer=licon1_PDIFF $count=1 $X=5.89
+ $Y=2.075 $X2=6.03 $Y2=2.9
r171 1 43 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=5.675
+ $Y=0.285 $X2=5.82 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__DLRTN_LP%A_744_415# 1 2 9 12 13 15 18 20 22 24 28 31
+ 33 36 41 45
c99 41 0 6.90166e-20 $X=4.91 $Y=1.59
c100 36 0 1.77071e-19 $X=5.54 $Y=1.59
r101 44 45 20.9834 $w=3.3e-07 $l=1.2e-07 $layer=POLY_cond $X=5.765 $Y=1.59
+ $X2=5.885 $Y2=1.59
r102 37 44 39.3438 $w=3.3e-07 $l=2.25e-07 $layer=POLY_cond $X=5.54 $Y=1.59
+ $X2=5.765 $Y2=1.59
r103 36 37 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.54
+ $Y=1.59 $X2=5.54 $Y2=1.59
r104 34 41 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.995 $Y=1.59
+ $X2=4.91 $Y2=1.59
r105 34 36 19.0328 $w=3.28e-07 $l=5.45e-07 $layer=LI1_cond $X=4.995 $Y=1.59
+ $X2=5.54 $Y2=1.59
r106 32 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.91 $Y=1.755
+ $X2=4.91 $Y2=1.59
r107 32 33 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=4.91 $Y=1.755
+ $X2=4.91 $Y2=2.055
r108 31 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.91 $Y=1.425
+ $X2=4.91 $Y2=1.59
r109 30 31 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=4.91 $Y=0.485
+ $X2=4.91 $Y2=1.425
r110 29 40 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.28 $Y=2.14
+ $X2=4.115 $Y2=2.14
r111 28 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.825 $Y=2.14
+ $X2=4.91 $Y2=2.055
r112 28 29 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=4.825 $Y=2.14
+ $X2=4.28 $Y2=2.14
r113 24 30 6.84389 $w=1.9e-07 $l=1.30767e-07 $layer=LI1_cond $X=4.825 $Y=0.39
+ $X2=4.91 $Y2=0.485
r114 24 26 36.4833 $w=1.88e-07 $l=6.25e-07 $layer=LI1_cond $X=4.825 $Y=0.39
+ $X2=4.2 $Y2=0.39
r115 20 40 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.115 $Y=2.225
+ $X2=4.115 $Y2=2.14
r116 20 22 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=4.115 $Y=2.225
+ $X2=4.115 $Y2=2.9
r117 16 18 76.9149 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=5.885 $Y=0.89
+ $X2=6.035 $Y2=0.89
r118 13 18 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.035 $Y=0.815
+ $X2=6.035 $Y2=0.89
r119 13 15 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=6.035 $Y=0.815
+ $X2=6.035 $Y2=0.495
r120 12 45 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.885 $Y=1.425
+ $X2=5.885 $Y2=1.59
r121 11 16 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.885 $Y=0.965
+ $X2=5.885 $Y2=0.89
r122 11 12 235.872 $w=1.5e-07 $l=4.6e-07 $layer=POLY_cond $X=5.885 $Y=0.965
+ $X2=5.885 $Y2=1.425
r123 7 44 9.34494 $w=2.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.765 $Y=1.755
+ $X2=5.765 $Y2=1.59
r124 7 9 203.732 $w=2.5e-07 $l=8.2e-07 $layer=POLY_cond $X=5.765 $Y=1.755
+ $X2=5.765 $Y2=2.575
r125 2 40 400 $w=1.7e-07 $l=4.61844e-07 $layer=licon1_PDIFF $count=1 $X=3.72
+ $Y=2.075 $X2=4.115 $Y2=2.22
r126 2 22 400 $w=1.7e-07 $l=1.00324e-06 $layer=licon1_PDIFF $count=1 $X=3.72
+ $Y=2.075 $X2=4.115 $Y2=2.9
r127 1 26 182 $w=1.7e-07 $l=3.18198e-07 $layer=licon1_NDIFF $count=1 $X=3.95
+ $Y=0.235 $X2=4.2 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_LP__DLRTN_LP%RESET_B 3 7 11 12 13 16 17
c50 11 0 1.77071e-19 $X=6.335 $Y=1.71
r51 16 17 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.335
+ $Y=1.37 $X2=6.335 $Y2=1.37
r52 13 17 5.98039 $w=6.68e-07 $l=3.35e-07 $layer=LI1_cond $X=6 $Y=1.54 $X2=6.335
+ $Y2=1.54
r53 11 16 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=6.335 $Y=1.71
+ $X2=6.335 $Y2=1.37
r54 11 12 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.335 $Y=1.71
+ $X2=6.335 $Y2=1.875
r55 10 16 41.8716 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.335 $Y=1.205
+ $X2=6.335 $Y2=1.37
r56 7 10 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=6.395 $Y=0.495
+ $X2=6.395 $Y2=1.205
r57 3 12 173.918 $w=2.5e-07 $l=7e-07 $layer=POLY_cond $X=6.295 $Y=2.575
+ $X2=6.295 $Y2=1.875
.ends

.subckt PM_SKY130_FD_SC_LP__DLRTN_LP%VPWR 1 2 3 4 15 19 23 29 32 33 35 36 38 39
+ 40 58 64 65 68
r74 68 69 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r75 65 69 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=6.48 $Y2=3.33
r76 64 65 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r77 62 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.725 $Y=3.33
+ $X2=6.56 $Y2=3.33
r78 62 64 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=6.725 $Y=3.33
+ $X2=7.44 $Y2=3.33
r79 61 69 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=6.48
+ $Y2=3.33
r80 60 61 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r81 58 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.395 $Y=3.33
+ $X2=6.56 $Y2=3.33
r82 58 60 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=6.395 $Y=3.33 $X2=6
+ $Y2=3.33
r83 57 61 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=3.33 $X2=6
+ $Y2=3.33
r84 56 57 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r85 53 56 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=3.12 $Y=3.33
+ $X2=5.04 $Y2=3.33
r86 53 54 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r87 51 54 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r88 50 51 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r89 48 51 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r90 47 50 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r91 47 48 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r92 44 48 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r93 43 44 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r94 40 57 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=3.84 $Y=3.33
+ $X2=5.04 $Y2=3.33
r95 40 54 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=3.84 $Y=3.33
+ $X2=3.12 $Y2=3.33
r96 38 56 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=5.175 $Y=3.33
+ $X2=5.04 $Y2=3.33
r97 38 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.175 $Y=3.33
+ $X2=5.34 $Y2=3.33
r98 37 60 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=5.505 $Y=3.33 $X2=6
+ $Y2=3.33
r99 37 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.505 $Y=3.33
+ $X2=5.34 $Y2=3.33
r100 35 50 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=2.755 $Y=3.33
+ $X2=2.64 $Y2=3.33
r101 35 36 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.755 $Y=3.33
+ $X2=2.88 $Y2=3.33
r102 34 53 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=3.005 $Y=3.33
+ $X2=3.12 $Y2=3.33
r103 34 36 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.005 $Y=3.33
+ $X2=2.88 $Y2=3.33
r104 32 43 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=0.765 $Y=3.33
+ $X2=0.72 $Y2=3.33
r105 32 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.765 $Y=3.33
+ $X2=0.93 $Y2=3.33
r106 31 47 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=1.095 $Y=3.33
+ $X2=1.2 $Y2=3.33
r107 31 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.095 $Y=3.33
+ $X2=0.93 $Y2=3.33
r108 27 68 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.56 $Y=3.245
+ $X2=6.56 $Y2=3.33
r109 27 29 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=6.56 $Y=3.245
+ $X2=6.56 $Y2=2.57
r110 23 26 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=5.34 $Y=2.22
+ $X2=5.34 $Y2=2.93
r111 21 39 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.34 $Y=3.245
+ $X2=5.34 $Y2=3.33
r112 21 26 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=5.34 $Y=3.245
+ $X2=5.34 $Y2=2.93
r113 17 36 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.88 $Y=3.245
+ $X2=2.88 $Y2=3.33
r114 17 19 45.4063 $w=2.48e-07 $l=9.85e-07 $layer=LI1_cond $X=2.88 $Y=3.245
+ $X2=2.88 $Y2=2.26
r115 13 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.93 $Y=3.245
+ $X2=0.93 $Y2=3.33
r116 13 15 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=0.93 $Y=3.245
+ $X2=0.93 $Y2=2.93
r117 4 29 300 $w=1.7e-07 $l=5.60647e-07 $layer=licon1_PDIFF $count=2 $X=6.42
+ $Y=2.075 $X2=6.56 $Y2=2.57
r118 3 26 400 $w=1.7e-07 $l=1.01292e-06 $layer=licon1_PDIFF $count=1 $X=4.995
+ $Y=2.075 $X2=5.34 $Y2=2.93
r119 3 23 400 $w=1.7e-07 $l=4.11157e-07 $layer=licon1_PDIFF $count=1 $X=4.995
+ $Y=2.075 $X2=5.34 $Y2=2.22
r120 2 19 300 $w=1.7e-07 $l=3.91727e-07 $layer=licon1_PDIFF $count=2 $X=2.53
+ $Y=2.075 $X2=2.84 $Y2=2.26
r121 1 15 600 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=0.79
+ $Y=2.075 $X2=0.93 $Y2=2.93
.ends

.subckt PM_SKY130_FD_SC_LP__DLRTN_LP%Q 1 2 7 8 9 10 11 12 13 36 39
r22 37 39 1.8556 $w=5.33e-07 $l=8.3e-08 $layer=LI1_cond $X=7.297 $Y=2.322
+ $X2=7.297 $Y2=2.405
r23 36 47 0.69845 $w=3.28e-07 $l=2e-08 $layer=LI1_cond $X=7.4 $Y=2.035 $X2=7.4
+ $Y2=2.055
r24 13 44 2.79458 $w=5.33e-07 $l=1.25e-07 $layer=LI1_cond $X=7.297 $Y=2.775
+ $X2=7.297 $Y2=2.9
r25 12 37 0.0223566 $w=5.33e-07 $l=1e-09 $layer=LI1_cond $X=7.297 $Y=2.321
+ $X2=7.297 $Y2=2.322
r26 12 49 2.25802 $w=5.33e-07 $l=1.01e-07 $layer=LI1_cond $X=7.297 $Y=2.321
+ $X2=7.297 $Y2=2.22
r27 12 13 8.24959 $w=5.33e-07 $l=3.69e-07 $layer=LI1_cond $X=7.297 $Y=2.406
+ $X2=7.297 $Y2=2.775
r28 12 39 0.0223566 $w=5.33e-07 $l=1e-09 $layer=LI1_cond $X=7.297 $Y=2.406
+ $X2=7.297 $Y2=2.405
r29 11 49 2.97343 $w=5.33e-07 $l=1.33e-07 $layer=LI1_cond $X=7.297 $Y=2.087
+ $X2=7.297 $Y2=2.22
r30 11 47 2.46032 $w=5.33e-07 $l=3.2e-08 $layer=LI1_cond $X=7.297 $Y=2.087
+ $X2=7.297 $Y2=2.055
r31 11 36 1.15244 $w=3.28e-07 $l=3.3e-08 $layer=LI1_cond $X=7.4 $Y=2.002 $X2=7.4
+ $Y2=2.035
r32 10 11 11.7689 $w=3.28e-07 $l=3.37e-07 $layer=LI1_cond $X=7.4 $Y=1.665
+ $X2=7.4 $Y2=2.002
r33 9 10 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=7.4 $Y=1.295 $X2=7.4
+ $Y2=1.665
r34 8 9 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=7.4 $Y=0.925 $X2=7.4
+ $Y2=1.295
r35 7 8 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=7.4 $Y=0.495 $X2=7.4
+ $Y2=0.925
r36 2 49 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=7.055
+ $Y=2.075 $X2=7.195 $Y2=2.22
r37 2 44 400 $w=1.7e-07 $l=8.92258e-07 $layer=licon1_PDIFF $count=1 $X=7.055
+ $Y=2.075 $X2=7.195 $Y2=2.9
r38 1 7 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=7.26
+ $Y=0.285 $X2=7.4 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__DLRTN_LP%VGND 1 2 3 4 15 17 21 25 29 32 33 34 36 48
+ 54 55 58 61 64
r103 64 65 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r104 61 62 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=0
+ $X2=3.12 $Y2=0
r105 59 62 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=1.2 $Y=0 $X2=3.12
+ $Y2=0
r106 58 59 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r107 55 65 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.44 $Y=0 $X2=6.48
+ $Y2=0
r108 54 55 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r109 52 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.775 $Y=0 $X2=6.61
+ $Y2=0
r110 52 54 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=6.775 $Y=0 $X2=7.44
+ $Y2=0
r111 51 65 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=6.48
+ $Y2=0
r112 50 51 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r113 48 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.445 $Y=0 $X2=6.61
+ $Y2=0
r114 48 50 60.3476 $w=1.68e-07 $l=9.25e-07 $layer=LI1_cond $X=6.445 $Y=0
+ $X2=5.52 $Y2=0
r115 47 51 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=5.52
+ $Y2=0
r116 46 47 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r117 44 62 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=3.12
+ $Y2=0
r118 43 46 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=3.6 $Y=0 $X2=5.04
+ $Y2=0
r119 43 44 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r120 41 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.435 $Y=0 $X2=3.27
+ $Y2=0
r121 41 43 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=3.435 $Y=0 $X2=3.6
+ $Y2=0
r122 39 59 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r123 38 39 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r124 36 58 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.905 $Y=0 $X2=1.07
+ $Y2=0
r125 36 38 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=0.905 $Y=0
+ $X2=0.72 $Y2=0
r126 34 47 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=3.84 $Y=0 $X2=5.04
+ $Y2=0
r127 34 44 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.84 $Y=0 $X2=3.6
+ $Y2=0
r128 32 46 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=5.175 $Y=0
+ $X2=5.04 $Y2=0
r129 32 33 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.175 $Y=0 $X2=5.3
+ $Y2=0
r130 31 50 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=5.425 $Y=0 $X2=5.52
+ $Y2=0
r131 31 33 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.425 $Y=0 $X2=5.3
+ $Y2=0
r132 27 64 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.61 $Y=0.085
+ $X2=6.61 $Y2=0
r133 27 29 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=6.61 $Y=0.085
+ $X2=6.61 $Y2=0.47
r134 23 33 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.3 $Y=0.085
+ $X2=5.3 $Y2=0
r135 23 25 16.5952 $w=2.48e-07 $l=3.6e-07 $layer=LI1_cond $X=5.3 $Y=0.085
+ $X2=5.3 $Y2=0.445
r136 19 61 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.27 $Y=0.085
+ $X2=3.27 $Y2=0
r137 19 21 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=3.27 $Y=0.085
+ $X2=3.27 $Y2=0.39
r138 18 58 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.235 $Y=0 $X2=1.07
+ $Y2=0
r139 17 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.105 $Y=0 $X2=3.27
+ $Y2=0
r140 17 18 122 $w=1.68e-07 $l=1.87e-06 $layer=LI1_cond $X=3.105 $Y=0 $X2=1.235
+ $Y2=0
r141 13 58 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.07 $Y=0.085
+ $X2=1.07 $Y2=0
r142 13 15 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=1.07 $Y=0.085
+ $X2=1.07 $Y2=0.445
r143 4 29 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=6.47
+ $Y=0.285 $X2=6.61 $Y2=0.47
r144 3 25 182 $w=1.7e-07 $l=2.93428e-07 $layer=licon1_NDIFF $count=1 $X=5.06
+ $Y=0.235 $X2=5.26 $Y2=0.445
r145 2 21 182 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=1 $X=3.13
+ $Y=0.235 $X2=3.27 $Y2=0.39
r146 1 15 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.93
+ $Y=0.235 $X2=1.07 $Y2=0.445
.ends

