* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__o311a_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
X0 a_355_367# A2 a_427_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X1 a_85_21# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X2 X a_85_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X3 X a_85_21# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X4 a_679_47# C1 a_85_21# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X5 VGND A1 a_355_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X6 VPWR a_85_21# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X7 VPWR C1 a_85_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X8 VGND A3 a_355_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X9 a_427_367# A3 a_85_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X10 VPWR A1 a_355_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X11 a_355_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X12 a_355_47# B1 a_679_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X13 VGND a_85_21# X VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
.ends
