* File: sky130_fd_sc_lp__sleep_pargate_plv_7.pex.spice
* Created: Fri Aug 28 11:32:28 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__SLEEP_PARGATE_PLV_7%SLEEP 1 3 5 6 7 8 9 16
c23 16 0 4.0798e-20 $X=8.42 $Y=1.985
r24 20 21 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=8.42
+ $Y=2.665 $X2=8.42 $Y2=2.665
r25 16 20 91.1288 $w=4.15e-07 $l=6.8e-07 $layer=POLY_cond $X=8.377 $Y=1.985
+ $X2=8.377 $Y2=2.665
r26 9 21 5.86755 $w=5.28e-07 $l=2.6e-07 $layer=LI1_cond $X=8.52 $Y=2.405
+ $X2=8.52 $Y2=2.665
r27 8 9 9.47836 $w=5.28e-07 $l=4.2e-07 $layer=LI1_cond $X=8.52 $Y=1.985 $X2=8.52
+ $Y2=2.405
r28 8 16 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=8.42
+ $Y=1.985 $X2=8.42 $Y2=1.985
r29 7 8 7.22161 $w=5.28e-07 $l=3.2e-07 $layer=LI1_cond $X=8.52 $Y=1.665 $X2=8.52
+ $Y2=1.985
r30 6 7 8.34998 $w=5.28e-07 $l=3.7e-07 $layer=LI1_cond $X=8.52 $Y=1.295 $X2=8.52
+ $Y2=1.665
r31 5 6 8.34998 $w=5.28e-07 $l=3.7e-07 $layer=LI1_cond $X=8.52 $Y=0.925 $X2=8.52
+ $Y2=1.295
r32 4 20 2.01019 $w=4.15e-07 $l=1.5e-08 $layer=POLY_cond $X=8.377 $Y=2.68
+ $X2=8.377 $Y2=2.665
r33 1 4 35.4752 $w=1.5e-07 $l=2.41607e-07 $layer=POLY_cond $X=8.17 $Y=2.755
+ $X2=8.377 $Y2=2.68
r34 1 3 1161.62 $w=1.5e-07 $l=3.615e-06 $layer=POLY_cond $X=8.17 $Y=2.755
+ $X2=4.555 $Y2=2.755
.ends

.subckt PM_SKY130_FD_SC_LP__SLEEP_PARGATE_PLV_7%VPWR 1 4 22 27 32 37 42 47 48
c48 47 0 4.0798e-20 $X=7.775 $Y=2.54
r49 47 48 2.25 $w=1.5e-07 $l=3e-07 $layer=via $count=2 $X=7.775 $Y=2.54
+ $X2=7.775 $Y2=2.54
r50 43 48 0.0591216 $w=3.33e-06 $l=1.575e-06 $layer=MET2_cond $X=6.2 $Y=1.665
+ $X2=7.775 $Y2=1.665
r51 42 43 2.25 $w=1.5e-07 $l=3e-07 $layer=via $count=2 $X=6.2 $Y=2.54 $X2=6.2
+ $Y2=2.54
r52 38 43 0.0583709 $w=3.33e-06 $l=1.555e-06 $layer=MET2_cond $X=4.645 $Y=1.665
+ $X2=6.2 $Y2=1.665
r53 37 38 2.25 $w=1.5e-07 $l=3e-07 $layer=via $count=2 $X=4.645 $Y=2.54
+ $X2=4.645 $Y2=2.54
r54 32 33 2.25 $w=1.5e-07 $l=3e-07 $layer=via $count=2 $X=3.09 $Y=2.54 $X2=3.09
+ $Y2=2.54
r55 28 33 0.0579955 $w=3.33e-06 $l=1.545e-06 $layer=MET2_cond $X=1.545 $Y=1.665
+ $X2=3.09 $Y2=1.665
r56 27 28 2.25 $w=1.5e-07 $l=3e-07 $layer=via $count=2 $X=1.545 $Y=2.54
+ $X2=1.545 $Y2=2.54
r57 22 47 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.8 $Y=2.54 $X2=7.8
+ $Y2=2.54
r58 19 22 69.1466 $w=2.58e-07 $l=1.56e-06 $layer=LI1_cond $X=6.225 $Y=2.54
+ $X2=7.785 $Y2=2.54
r59 19 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.225 $Y=2.54
+ $X2=6.225 $Y2=2.54
r60 16 19 68.925 $w=2.58e-07 $l=1.555e-06 $layer=LI1_cond $X=4.67 $Y=2.54
+ $X2=6.225 $Y2=2.54
r61 16 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.67 $Y=2.54
+ $X2=4.67 $Y2=2.54
r62 13 16 68.925 $w=2.58e-07 $l=1.555e-06 $layer=LI1_cond $X=3.115 $Y=2.54
+ $X2=4.67 $Y2=2.54
r63 13 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.115 $Y=2.54
+ $X2=3.115 $Y2=2.54
r64 10 13 68.925 $w=2.58e-07 $l=1.555e-06 $layer=LI1_cond $X=1.56 $Y=2.54
+ $X2=3.115 $Y2=2.54
r65 10 27 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.56 $Y=2.54
+ $X2=1.56 $Y2=2.54
r66 7 10 10.4163 $w=2.58e-07 $l=2.35e-07 $layer=LI1_cond $X=1.325 $Y=2.54
+ $X2=1.56 $Y2=2.54
r67 4 38 0.00319069 $w=3.33e-06 $l=8.5e-08 $layer=MET2_cond $X=4.56 $Y=1.665
+ $X2=4.645 $Y2=1.665
r68 4 33 0.0551802 $w=3.33e-06 $l=1.47e-06 $layer=MET2_cond $X=4.56 $Y=1.665
+ $X2=3.09 $Y2=1.665
r69 1 22 60 $w=1.7e-07 $l=6.79221e-06 $layer=licon1_PDIFF $count=10 $X=1.055
+ $Y=2.415 $X2=7.785 $Y2=2.54
r70 1 7 60 $w=1.7e-07 $l=3.26573e-07 $layer=licon1_PDIFF $count=10 $X=1.055
+ $Y=2.415 $X2=1.325 $Y2=2.54
.ends

.subckt PM_SKY130_FD_SC_LP__SLEEP_PARGATE_PLV_7%VIRTPWR 1 4 8 9 23 29 38 44 53
+ 56 57 64 65 70 74 79 80
c59 80 0 1.43534e-19 $X=6.51 $Y=3.33
c60 74 0 1.43534e-19 $X=4.955 $Y=3.33
c61 70 0 1.43534e-19 $X=3.4 $Y=3.33
c62 53 0 9.97624e-20 $X=7.005 $Y=2.97
c63 44 0 9.6669e-20 $X=5.45 $Y=2.97
c64 38 0 9.6669e-20 $X=3.895 $Y=2.97
c65 29 0 9.6669e-20 $X=1.98 $Y=2.97
r66 80 84 0.024068 $w=4.9e-07 $l=3.23e-07 $layer=MET1_cond $X=6.832 $Y=3.33
+ $X2=7.155 $Y2=3.33
r67 74 81 0.022181 $w=4.9e-07 $l=3.13e-07 $layer=MET1_cond $X=5.267 $Y=3.33
+ $X2=5.58 $Y2=3.33
r68 74 79 0.0432039 $w=4.9e-07 $l=1.55e-07 $layer=MET1_cond $X=4.955 $Y=3.33
+ $X2=4.8 $Y2=3.33
r69 70 75 0.022181 $w=4.9e-07 $l=3.13e-07 $layer=MET1_cond $X=3.712 $Y=3.33
+ $X2=4.025 $Y2=3.33
r70 65 71 0.022181 $w=4.9e-07 $l=3.13e-07 $layer=MET1_cond $X=2.157 $Y=3.33
+ $X2=2.47 $Y2=3.33
r71 63 84 0.213232 $w=4.9e-07 $l=7.65e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=7.155 $Y2=3.33
r72 62 64 9.36939 $w=5.73e-07 $l=1.35e-07 $layer=LI1_cond $X=7.92 $Y=3.127
+ $X2=8.055 $Y2=3.127
r73 62 63 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r74 60 62 2.80818 $w=5.73e-07 $l=1.35e-07 $layer=LI1_cond $X=7.785 $Y=3.127
+ $X2=7.92 $Y2=3.127
r75 56 64 53.8235 $w=1.68e-07 $l=8.25e-07 $layer=LI1_cond $X=8.88 $Y=3.33
+ $X2=8.055 $Y2=3.33
r76 56 57 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r77 52 53 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=7.005 $Y=2.97
+ $X2=7.005 $Y2=2.97
r78 50 80 0.00836204 $w=4.9e-07 $l=3e-08 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=6.51 $Y2=3.33
r79 49 52 10.9207 $w=5.73e-07 $l=5.25e-07 $layer=LI1_cond $X=6.48 $Y=3.127
+ $X2=7.005 $Y2=3.127
r80 49 50 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r81 46 49 19.9693 $w=5.73e-07 $l=9.6e-07 $layer=LI1_cond $X=5.52 $Y=3.127
+ $X2=6.48 $Y2=3.127
r82 46 74 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r83 43 46 1.4561 $w=5.73e-07 $l=7e-08 $layer=LI1_cond $X=5.45 $Y=3.127 $X2=5.52
+ $Y2=3.127
r84 43 44 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=5.45 $Y=2.97
+ $X2=5.45 $Y2=2.97
r85 41 79 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=4.8 $Y2=3.33
r86 40 43 18.5132 $w=5.73e-07 $l=8.9e-07 $layer=LI1_cond $X=4.56 $Y=3.127
+ $X2=5.45 $Y2=3.127
r87 40 41 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r88 37 40 13.8329 $w=5.73e-07 $l=6.65e-07 $layer=LI1_cond $X=3.895 $Y=3.127
+ $X2=4.56 $Y2=3.127
r89 37 38 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.895 $Y=2.97
+ $X2=3.895 $Y2=2.97
r90 35 70 0.0780457 $w=4.9e-07 $l=2.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.4 $Y2=3.33
r91 34 37 16.1211 $w=5.73e-07 $l=7.75e-07 $layer=LI1_cond $X=3.12 $Y=3.127
+ $X2=3.895 $Y2=3.127
r92 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r93 31 34 16.2251 $w=5.73e-07 $l=7.8e-07 $layer=LI1_cond $X=2.34 $Y=3.127
+ $X2=3.12 $Y2=3.127
r94 29 31 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.34 $Y=2.97
+ $X2=2.34 $Y2=2.97
r95 28 31 7.48849 $w=5.73e-07 $l=3.6e-07 $layer=LI1_cond $X=1.98 $Y=3.127
+ $X2=2.34 $Y2=3.127
r96 28 29 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.98 $Y=2.97
+ $X2=1.98 $Y2=2.97
r97 26 65 0.0459912 $w=4.9e-07 $l=1.65e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.845 $Y2=3.33
r98 25 28 6.24041 $w=5.73e-07 $l=3e-07 $layer=LI1_cond $X=1.68 $Y=3.127 $X2=1.98
+ $Y2=3.127
r99 25 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r100 23 60 0.353623 $w=5.73e-07 $l=1.7e-08 $layer=LI1_cond $X=7.768 $Y=3.127
+ $X2=7.785 $Y2=3.127
r101 23 52 15.8714 $w=5.73e-07 $l=7.63e-07 $layer=LI1_cond $X=7.768 $Y=3.127
+ $X2=7.005 $Y2=3.127
r102 20 21 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r103 9 80 0.0250352 $w=6.45e-07 $l=1.23e-07 $layer=MET1_cond $X=6.832 $Y=3.207
+ $X2=6.832 $Y2=3.33
r104 9 53 0.0482385 $w=6.45e-07 $l=2.37e-07 $layer=MET1_cond $X=6.832 $Y=3.207
+ $X2=6.832 $Y2=2.97
r105 9 74 0.0258363 $w=6.25e-07 $l=1.23e-07 $layer=MET1_cond $X=5.267 $Y=3.207
+ $X2=5.267 $Y2=3.33
r106 9 44 0.0497821 $w=6.25e-07 $l=2.37e-07 $layer=MET1_cond $X=5.267 $Y=3.207
+ $X2=5.267 $Y2=2.97
r107 9 70 0.0258363 $w=6.25e-07 $l=1.23e-07 $layer=MET1_cond $X=3.712 $Y=3.207
+ $X2=3.712 $Y2=3.33
r108 9 38 0.0497821 $w=6.25e-07 $l=2.37e-07 $layer=MET1_cond $X=3.712 $Y=3.207
+ $X2=3.712 $Y2=2.97
r109 9 65 0.0258363 $w=6.25e-07 $l=1.23e-07 $layer=MET1_cond $X=2.157 $Y=3.207
+ $X2=2.157 $Y2=3.33
r110 9 29 0.0497821 $w=6.25e-07 $l=2.37e-07 $layer=MET1_cond $X=2.157 $Y=3.207
+ $X2=2.157 $Y2=2.97
r111 9 57 0.2071 $w=4.9e-07 $l=7.43e-07 $layer=MET1_cond $X=8.137 $Y=3.33
+ $X2=8.88 $Y2=3.33
r112 9 63 0.0604854 $w=4.9e-07 $l=2.17e-07 $layer=MET1_cond $X=8.137 $Y=3.33
+ $X2=7.92 $Y2=3.33
r113 9 50 0.12125 $w=4.9e-07 $l=4.35e-07 $layer=MET1_cond $X=6.045 $Y=3.33
+ $X2=6.48 $Y2=3.33
r114 9 81 0.129612 $w=4.9e-07 $l=4.65e-07 $layer=MET1_cond $X=6.045 $Y=3.33
+ $X2=5.58 $Y2=3.33
r115 9 41 0.0195114 $w=4.9e-07 $l=7e-08 $layer=MET1_cond $X=4.49 $Y=3.33
+ $X2=4.56 $Y2=3.33
r116 9 75 0.129612 $w=4.9e-07 $l=4.65e-07 $layer=MET1_cond $X=4.49 $Y=3.33
+ $X2=4.025 $Y2=3.33
r117 9 35 0.0515659 $w=4.9e-07 $l=1.85e-07 $layer=MET1_cond $X=2.935 $Y=3.33
+ $X2=3.12 $Y2=3.33
r118 9 71 0.129612 $w=4.9e-07 $l=4.65e-07 $layer=MET1_cond $X=2.935 $Y=3.33
+ $X2=2.47 $Y2=3.33
r119 9 26 0.211281 $w=4.9e-07 $l=7.58e-07 $layer=MET1_cond $X=0.922 $Y=3.33
+ $X2=1.68 $Y2=3.33
r120 9 21 0.0563044 $w=4.9e-07 $l=2.02e-07 $layer=MET1_cond $X=0.922 $Y=3.33
+ $X2=0.72 $Y2=3.33
r121 8 20 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.055 $Y=3.33
+ $X2=0.72 $Y2=3.33
r122 7 8 12.1776 $w=5.73e-07 $l=2.7e-07 $layer=LI1_cond $X=1.325 $Y=3.127
+ $X2=1.055 $Y2=3.127
r123 4 25 7.03086 $w=5.73e-07 $l=3.38e-07 $layer=LI1_cond $X=1.342 $Y=3.127
+ $X2=1.68 $Y2=3.127
r124 4 7 0.353623 $w=5.73e-07 $l=1.7e-08 $layer=LI1_cond $X=1.342 $Y=3.127
+ $X2=1.325 $Y2=3.127
r125 1 60 60 $w=1.7e-07 $l=6.79964e-06 $layer=licon1_PDIFF $count=10 $X=1.055
+ $Y=2.83 $X2=7.785 $Y2=2.97
r126 1 7 60 $w=1.7e-07 $l=3.32716e-07 $layer=licon1_PDIFF $count=10 $X=1.055
+ $Y=2.83 $X2=1.325 $Y2=2.97
.ends

