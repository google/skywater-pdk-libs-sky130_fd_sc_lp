* File: sky130_fd_sc_lp__sdfxtp_2.pxi.spice
* Created: Fri Aug 28 11:30:48 2020
* 
x_PM_SKY130_FD_SC_LP__SDFXTP_2%A_55_119# N_A_55_119#_M1008_s N_A_55_119#_M1029_s
+ N_A_55_119#_M1007_g N_A_55_119#_M1005_g N_A_55_119#_c_229_n
+ N_A_55_119#_c_235_n N_A_55_119#_c_258_p N_A_55_119#_c_236_n
+ N_A_55_119#_c_230_n N_A_55_119#_c_231_n N_A_55_119#_c_238_n
+ N_A_55_119#_c_239_n N_A_55_119#_c_232_n N_A_55_119#_c_240_n
+ PM_SKY130_FD_SC_LP__SDFXTP_2%A_55_119#
x_PM_SKY130_FD_SC_LP__SDFXTP_2%D N_D_M1004_g N_D_M1018_g D D D N_D_c_316_n
+ N_D_c_317_n PM_SKY130_FD_SC_LP__SDFXTP_2%D
x_PM_SKY130_FD_SC_LP__SDFXTP_2%SCE N_SCE_c_363_n N_SCE_M1008_g N_SCE_c_364_n
+ N_SCE_M1029_g N_SCE_c_357_n N_SCE_c_358_n N_SCE_c_365_n N_SCE_c_366_n
+ N_SCE_M1030_g N_SCE_M1017_g N_SCE_c_360_n N_SCE_c_368_n N_SCE_c_369_n SCE SCE
+ SCE N_SCE_c_362_n PM_SKY130_FD_SC_LP__SDFXTP_2%SCE
x_PM_SKY130_FD_SC_LP__SDFXTP_2%SCD N_SCD_M1001_g N_SCD_M1009_g SCD SCD
+ N_SCD_c_430_n PM_SKY130_FD_SC_LP__SDFXTP_2%SCD
x_PM_SKY130_FD_SC_LP__SDFXTP_2%CLK N_CLK_M1031_g N_CLK_M1023_g N_CLK_c_480_n
+ N_CLK_c_481_n CLK CLK CLK N_CLK_c_478_n PM_SKY130_FD_SC_LP__SDFXTP_2%CLK
x_PM_SKY130_FD_SC_LP__SDFXTP_2%A_610_487# N_A_610_487#_M1023_d
+ N_A_610_487#_M1031_d N_A_610_487#_M1032_g N_A_610_487#_c_539_n
+ N_A_610_487#_M1006_g N_A_610_487#_M1012_g N_A_610_487#_M1011_g
+ N_A_610_487#_M1019_g N_A_610_487#_M1026_g N_A_610_487#_c_528_n
+ N_A_610_487#_c_543_n N_A_610_487#_c_529_n N_A_610_487#_c_544_n
+ N_A_610_487#_c_545_n N_A_610_487#_c_530_n N_A_610_487#_c_531_n
+ N_A_610_487#_c_603_p N_A_610_487#_c_547_n N_A_610_487#_c_548_n
+ N_A_610_487#_c_549_n N_A_610_487#_c_550_n N_A_610_487#_c_551_n
+ N_A_610_487#_c_635_p N_A_610_487#_c_627_p N_A_610_487#_c_709_p
+ N_A_610_487#_c_552_n N_A_610_487#_c_532_n N_A_610_487#_c_533_n
+ N_A_610_487#_c_585_p N_A_610_487#_c_534_n N_A_610_487#_c_535_n
+ N_A_610_487#_c_605_p N_A_610_487#_c_536_n N_A_610_487#_c_670_p
+ N_A_610_487#_c_555_n N_A_610_487#_c_556_n N_A_610_487#_c_537_n
+ N_A_610_487#_c_538_n PM_SKY130_FD_SC_LP__SDFXTP_2%A_610_487#
x_PM_SKY130_FD_SC_LP__SDFXTP_2%A_831_47# N_A_831_47#_M1032_d N_A_831_47#_M1006_d
+ N_A_831_47#_c_780_n N_A_831_47#_c_781_n N_A_831_47#_c_782_n
+ N_A_831_47#_c_783_n N_A_831_47#_M1021_g N_A_831_47#_M1027_g
+ N_A_831_47#_M1033_g N_A_831_47#_c_762_n N_A_831_47#_c_763_n
+ N_A_831_47#_c_764_n N_A_831_47#_M1016_g N_A_831_47#_c_785_n
+ N_A_831_47#_c_766_n N_A_831_47#_c_767_n N_A_831_47#_c_768_n
+ N_A_831_47#_c_769_n N_A_831_47#_c_770_n N_A_831_47#_c_771_n
+ N_A_831_47#_c_843_p N_A_831_47#_c_860_p N_A_831_47#_c_844_p
+ N_A_831_47#_c_772_n N_A_831_47#_c_773_n N_A_831_47#_c_774_n
+ N_A_831_47#_c_775_n N_A_831_47#_c_776_n N_A_831_47#_c_777_n
+ N_A_831_47#_c_778_n N_A_831_47#_c_779_n PM_SKY130_FD_SC_LP__SDFXTP_2%A_831_47#
x_PM_SKY130_FD_SC_LP__SDFXTP_2%A_1178_399# N_A_1178_399#_M1015_d
+ N_A_1178_399#_M1014_d N_A_1178_399#_M1002_g N_A_1178_399#_M1020_g
+ N_A_1178_399#_c_935_n N_A_1178_399#_c_942_n N_A_1178_399#_c_936_n
+ N_A_1178_399#_c_937_n N_A_1178_399#_c_945_n N_A_1178_399#_c_938_n
+ N_A_1178_399#_c_939_n N_A_1178_399#_c_940_n
+ PM_SKY130_FD_SC_LP__SDFXTP_2%A_1178_399#
x_PM_SKY130_FD_SC_LP__SDFXTP_2%A_1047_125# N_A_1047_125#_M1012_d
+ N_A_1047_125#_M1021_d N_A_1047_125#_M1014_g N_A_1047_125#_c_1012_n
+ N_A_1047_125#_M1015_g N_A_1047_125#_c_1013_n N_A_1047_125#_c_1014_n
+ N_A_1047_125#_c_1021_n N_A_1047_125#_c_1015_n N_A_1047_125#_c_1022_n
+ N_A_1047_125#_c_1016_n N_A_1047_125#_c_1017_n N_A_1047_125#_c_1018_n
+ PM_SKY130_FD_SC_LP__SDFXTP_2%A_1047_125#
x_PM_SKY130_FD_SC_LP__SDFXTP_2%A_1665_381# N_A_1665_381#_M1025_d
+ N_A_1665_381#_M1000_d N_A_1665_381#_M1022_g N_A_1665_381#_M1028_g
+ N_A_1665_381#_c_1107_n N_A_1665_381#_M1003_g N_A_1665_381#_M1013_g
+ N_A_1665_381#_c_1108_n N_A_1665_381#_M1010_g N_A_1665_381#_M1024_g
+ N_A_1665_381#_c_1119_n N_A_1665_381#_c_1109_n N_A_1665_381#_c_1120_n
+ N_A_1665_381#_c_1110_n N_A_1665_381#_c_1121_n N_A_1665_381#_c_1111_n
+ N_A_1665_381#_c_1112_n N_A_1665_381#_c_1123_n N_A_1665_381#_c_1113_n
+ N_A_1665_381#_c_1125_n N_A_1665_381#_c_1114_n
+ PM_SKY130_FD_SC_LP__SDFXTP_2%A_1665_381#
x_PM_SKY130_FD_SC_LP__SDFXTP_2%A_1517_63# N_A_1517_63#_M1033_d
+ N_A_1517_63#_M1019_d N_A_1517_63#_M1025_g N_A_1517_63#_M1000_g
+ N_A_1517_63#_c_1210_n N_A_1517_63#_c_1211_n N_A_1517_63#_c_1224_n
+ N_A_1517_63#_c_1212_n N_A_1517_63#_c_1213_n N_A_1517_63#_c_1220_n
+ N_A_1517_63#_c_1221_n N_A_1517_63#_c_1214_n N_A_1517_63#_c_1215_n
+ N_A_1517_63#_c_1216_n PM_SKY130_FD_SC_LP__SDFXTP_2%A_1517_63#
x_PM_SKY130_FD_SC_LP__SDFXTP_2%VPWR N_VPWR_M1029_d N_VPWR_M1001_d N_VPWR_M1006_s
+ N_VPWR_M1002_d N_VPWR_M1022_d N_VPWR_M1013_s N_VPWR_M1024_s N_VPWR_c_1308_n
+ N_VPWR_c_1309_n N_VPWR_c_1310_n N_VPWR_c_1311_n N_VPWR_c_1312_n
+ N_VPWR_c_1313_n N_VPWR_c_1314_n N_VPWR_c_1315_n N_VPWR_c_1316_n
+ N_VPWR_c_1317_n N_VPWR_c_1318_n N_VPWR_c_1319_n N_VPWR_c_1320_n VPWR
+ N_VPWR_c_1321_n N_VPWR_c_1322_n N_VPWR_c_1323_n N_VPWR_c_1324_n
+ N_VPWR_c_1325_n N_VPWR_c_1326_n N_VPWR_c_1327_n N_VPWR_c_1328_n
+ N_VPWR_c_1307_n PM_SKY130_FD_SC_LP__SDFXTP_2%VPWR
x_PM_SKY130_FD_SC_LP__SDFXTP_2%A_328_119# N_A_328_119#_M1004_d
+ N_A_328_119#_M1012_s N_A_328_119#_M1018_d N_A_328_119#_M1021_s
+ N_A_328_119#_c_1447_n N_A_328_119#_c_1462_n N_A_328_119#_c_1448_n
+ N_A_328_119#_c_1449_n N_A_328_119#_c_1453_n N_A_328_119#_c_1454_n
+ N_A_328_119#_c_1450_n N_A_328_119#_c_1451_n N_A_328_119#_c_1452_n
+ N_A_328_119#_c_1457_n N_A_328_119#_c_1458_n N_A_328_119#_c_1459_n
+ N_A_328_119#_c_1460_n N_A_328_119#_c_1534_n N_A_328_119#_c_1461_n
+ PM_SKY130_FD_SC_LP__SDFXTP_2%A_328_119#
x_PM_SKY130_FD_SC_LP__SDFXTP_2%Q N_Q_M1003_d N_Q_M1013_d Q Q Q Q Q Q Q
+ PM_SKY130_FD_SC_LP__SDFXTP_2%Q
x_PM_SKY130_FD_SC_LP__SDFXTP_2%VGND N_VGND_M1008_d N_VGND_M1009_d N_VGND_M1032_s
+ N_VGND_M1020_d N_VGND_M1028_d N_VGND_M1003_s N_VGND_M1010_s N_VGND_c_1596_n
+ N_VGND_c_1597_n N_VGND_c_1598_n N_VGND_c_1599_n N_VGND_c_1600_n
+ N_VGND_c_1601_n N_VGND_c_1602_n N_VGND_c_1603_n N_VGND_c_1604_n
+ N_VGND_c_1605_n N_VGND_c_1606_n N_VGND_c_1607_n N_VGND_c_1608_n
+ N_VGND_c_1609_n N_VGND_c_1610_n VGND N_VGND_c_1611_n N_VGND_c_1612_n
+ N_VGND_c_1613_n N_VGND_c_1614_n N_VGND_c_1615_n N_VGND_c_1616_n
+ N_VGND_c_1617_n PM_SKY130_FD_SC_LP__SDFXTP_2%VGND
cc_1 VNB N_A_55_119#_M1007_g 0.0366998f $X=-0.19 $Y=-0.245 $X2=1.205 $Y2=0.805
cc_2 VNB N_A_55_119#_c_229_n 0.0324232f $X=-0.19 $Y=-0.245 $X2=0.195 $Y2=2.3
cc_3 VNB N_A_55_119#_c_230_n 0.00481746f $X=-0.19 $Y=-0.245 $X2=1.085 $Y2=1.8
cc_4 VNB N_A_55_119#_c_231_n 0.00884453f $X=-0.19 $Y=-0.245 $X2=1.085 $Y2=1.8
cc_5 VNB N_A_55_119#_c_232_n 0.0173222f $X=-0.19 $Y=-0.245 $X2=0.42 $Y2=0.805
cc_6 VNB N_D_M1018_g 0.0125615f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB D 0.0181786f $X=-0.19 $Y=-0.245 $X2=1.205 $Y2=0.805
cc_8 VNB N_D_c_316_n 0.0364292f $X=-0.19 $Y=-0.245 $X2=1 $Y2=2.385
cc_9 VNB N_D_c_317_n 0.012663f $X=-0.19 $Y=-0.245 $X2=1.125 $Y2=1.945
cc_10 VNB N_SCE_M1008_g 0.0411022f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_SCE_c_357_n 0.120351f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_SCE_c_358_n 0.012806f $X=-0.19 $Y=-0.245 $X2=1.995 $Y2=2.275
cc_13 VNB N_SCE_M1017_g 0.0359959f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=2.56
cc_14 VNB N_SCE_c_360_n 0.0211933f $X=-0.19 $Y=-0.245 $X2=1.125 $Y2=1.945
cc_15 VNB SCE 0.00813091f $X=-0.19 $Y=-0.245 $X2=1.085 $Y2=1.8
cc_16 VNB N_SCE_c_362_n 0.0176677f $X=-0.19 $Y=-0.245 $X2=0.195 $Y2=0.805
cc_17 VNB N_SCD_M1009_g 0.0324328f $X=-0.19 $Y=-0.245 $X2=1.205 $Y2=1.635
cc_18 VNB SCD 0.00802221f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_SCD_c_430_n 0.0263858f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_CLK_M1023_g 0.041342f $X=-0.19 $Y=-0.245 $X2=1.205 $Y2=1.635
cc_21 VNB CLK 0.0100624f $X=-0.19 $Y=-0.245 $X2=1.995 $Y2=2.755
cc_22 VNB N_CLK_c_478_n 0.0275321f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_610_487#_M1032_g 0.0646175f $X=-0.19 $Y=-0.245 $X2=1.205 $Y2=0.805
cc_24 VNB N_A_610_487#_M1012_g 0.0361715f $X=-0.19 $Y=-0.245 $X2=0.195 $Y2=2.3
cc_25 VNB N_A_610_487#_c_528_n 0.00462692f $X=-0.19 $Y=-0.245 $X2=2.015 $Y2=2.11
cc_26 VNB N_A_610_487#_c_529_n 0.0206539f $X=-0.19 $Y=-0.245 $X2=0.42 $Y2=0.805
cc_27 VNB N_A_610_487#_c_530_n 0.00813654f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_610_487#_c_531_n 0.0171902f $X=-0.19 $Y=-0.245 $X2=2.015 $Y2=2.275
cc_29 VNB N_A_610_487#_c_532_n 0.00211762f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_610_487#_c_533_n 0.0100368f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_610_487#_c_534_n 0.0033081f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_610_487#_c_535_n 0.0356013f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_610_487#_c_536_n 0.00234234f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_610_487#_c_537_n 0.0361233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_610_487#_c_538_n 0.019074f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_831_47#_c_762_n 0.0299486f $X=-0.19 $Y=-0.245 $X2=1 $Y2=2.385
cc_37 VNB N_A_831_47#_c_763_n 0.0196383f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=2.385
cc_38 VNB N_A_831_47#_c_764_n 0.01815f $X=-0.19 $Y=-0.245 $X2=1.125 $Y2=1.945
cc_39 VNB N_A_831_47#_M1016_g 0.00772025f $X=-0.19 $Y=-0.245 $X2=1.085 $Y2=1.8
cc_40 VNB N_A_831_47#_c_766_n 0.00456154f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_831_47#_c_767_n 0.00195821f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_831_47#_c_768_n 0.0427691f $X=-0.19 $Y=-0.245 $X2=0.42 $Y2=0.805
cc_43 VNB N_A_831_47#_c_769_n 0.0280353f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_831_47#_c_770_n 0.0476232f $X=-0.19 $Y=-0.245 $X2=1.205 $Y2=1.8
cc_45 VNB N_A_831_47#_c_771_n 0.00117389f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_831_47#_c_772_n 0.00513335f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_831_47#_c_773_n 0.00201478f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_831_47#_c_774_n 0.0014026f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_831_47#_c_775_n 0.020026f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_831_47#_c_776_n 0.00349975f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_831_47#_c_777_n 0.0112294f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_831_47#_c_778_n 0.0132198f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_831_47#_c_779_n 0.019017f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_1178_399#_M1020_g 0.030873f $X=-0.19 $Y=-0.245 $X2=1.995 $Y2=2.755
cc_55 VNB N_A_1178_399#_c_935_n 0.00919998f $X=-0.19 $Y=-0.245 $X2=0.195 $Y2=2.3
cc_56 VNB N_A_1178_399#_c_936_n 0.00362566f $X=-0.19 $Y=-0.245 $X2=0.462
+ $Y2=2.56
cc_57 VNB N_A_1178_399#_c_937_n 0.00591493f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_1178_399#_c_938_n 0.0114283f $X=-0.19 $Y=-0.245 $X2=1.085 $Y2=1.8
cc_59 VNB N_A_1178_399#_c_939_n 0.0208809f $X=-0.19 $Y=-0.245 $X2=2.015 $Y2=2.11
cc_60 VNB N_A_1178_399#_c_940_n 8.6333e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_A_1047_125#_M1014_g 0.0160399f $X=-0.19 $Y=-0.245 $X2=1.205
+ $Y2=0.805
cc_62 VNB N_A_1047_125#_c_1012_n 0.0226521f $X=-0.19 $Y=-0.245 $X2=1.995
+ $Y2=2.275
cc_63 VNB N_A_1047_125#_c_1013_n 0.00265201f $X=-0.19 $Y=-0.245 $X2=0.195
+ $Y2=0.97
cc_64 VNB N_A_1047_125#_c_1014_n 4.74114e-19 $X=-0.19 $Y=-0.245 $X2=0.462
+ $Y2=2.56
cc_65 VNB N_A_1047_125#_c_1015_n 0.00247535f $X=-0.19 $Y=-0.245 $X2=1.085
+ $Y2=1.8
cc_66 VNB N_A_1047_125#_c_1016_n 0.00106972f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_A_1047_125#_c_1017_n 0.0197369f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_A_1047_125#_c_1018_n 0.045112f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_1665_381#_M1028_g 0.0567343f $X=-0.19 $Y=-0.245 $X2=1.995
+ $Y2=2.755
cc_70 VNB N_A_1665_381#_c_1107_n 0.0185197f $X=-0.19 $Y=-0.245 $X2=0.195
+ $Y2=0.97
cc_71 VNB N_A_1665_381#_c_1108_n 0.0192418f $X=-0.19 $Y=-0.245 $X2=0.61
+ $Y2=2.385
cc_72 VNB N_A_1665_381#_c_1109_n 0.00478064f $X=-0.19 $Y=-0.245 $X2=0.42
+ $Y2=0.805
cc_73 VNB N_A_1665_381#_c_1110_n 0.0100767f $X=-0.19 $Y=-0.245 $X2=1.205 $Y2=1.8
cc_74 VNB N_A_1665_381#_c_1111_n 0.00866028f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_A_1665_381#_c_1112_n 0.0062369f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_A_1665_381#_c_1113_n 0.00367887f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_A_1665_381#_c_1114_n 0.0594528f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_A_1517_63#_M1025_g 0.0308613f $X=-0.19 $Y=-0.245 $X2=1.205 $Y2=0.805
cc_79 VNB N_A_1517_63#_c_1210_n 0.024581f $X=-0.19 $Y=-0.245 $X2=0.462 $Y2=2.47
cc_80 VNB N_A_1517_63#_c_1211_n 0.00109937f $X=-0.19 $Y=-0.245 $X2=0.462
+ $Y2=2.56
cc_81 VNB N_A_1517_63#_c_1212_n 0.00111963f $X=-0.19 $Y=-0.245 $X2=1.25 $Y2=2.11
cc_82 VNB N_A_1517_63#_c_1213_n 0.00295336f $X=-0.19 $Y=-0.245 $X2=2.015
+ $Y2=2.11
cc_83 VNB N_A_1517_63#_c_1214_n 0.00668664f $X=-0.19 $Y=-0.245 $X2=0.42
+ $Y2=0.805
cc_84 VNB N_A_1517_63#_c_1215_n 0.0113029f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_A_1517_63#_c_1216_n 0.0177183f $X=-0.19 $Y=-0.245 $X2=0.195
+ $Y2=2.385
cc_86 VNB N_VPWR_c_1307_n 0.462217f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_A_328_119#_c_1447_n 0.0017092f $X=-0.19 $Y=-0.245 $X2=0.462 $Y2=2.47
cc_88 VNB N_A_328_119#_c_1448_n 0.0190865f $X=-0.19 $Y=-0.245 $X2=1 $Y2=2.385
cc_89 VNB N_A_328_119#_c_1449_n 0.00342293f $X=-0.19 $Y=-0.245 $X2=0.61
+ $Y2=2.385
cc_90 VNB N_A_328_119#_c_1450_n 0.00294697f $X=-0.19 $Y=-0.245 $X2=1.085 $Y2=1.8
cc_91 VNB N_A_328_119#_c_1451_n 0.0045634f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_A_328_119#_c_1452_n 0.0119432f $X=-0.19 $Y=-0.245 $X2=1.25 $Y2=2.11
cc_93 VNB Q 0.00451818f $X=-0.19 $Y=-0.245 $X2=1.205 $Y2=1.635
cc_94 VNB N_VGND_c_1596_n 0.0110712f $X=-0.19 $Y=-0.245 $X2=1.125 $Y2=1.8
cc_95 VNB N_VGND_c_1597_n 0.0182157f $X=-0.19 $Y=-0.245 $X2=1.25 $Y2=2.11
cc_96 VNB N_VGND_c_1598_n 0.00726878f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_97 VNB N_VGND_c_1599_n 0.0106398f $X=-0.19 $Y=-0.245 $X2=0.42 $Y2=0.805
cc_98 VNB N_VGND_c_1600_n 0.0560351f $X=-0.19 $Y=-0.245 $X2=0.195 $Y2=2.385
cc_99 VNB N_VGND_c_1601_n 0.0070026f $X=-0.19 $Y=-0.245 $X2=1.085 $Y2=1.8
cc_100 VNB N_VGND_c_1602_n 0.0137f $X=-0.19 $Y=-0.245 $X2=2.015 $Y2=2.275
cc_101 VNB N_VGND_c_1603_n 0.0113208f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_102 VNB N_VGND_c_1604_n 0.0515222f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_103 VNB N_VGND_c_1605_n 0.0222099f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_104 VNB N_VGND_c_1606_n 0.00292972f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_105 VNB N_VGND_c_1607_n 0.0489704f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_106 VNB N_VGND_c_1608_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_107 VNB N_VGND_c_1609_n 0.0194265f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_108 VNB N_VGND_c_1610_n 0.00513462f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_109 VNB N_VGND_c_1611_n 0.0510706f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_110 VNB N_VGND_c_1612_n 0.0190669f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_111 VNB N_VGND_c_1613_n 0.0165716f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_112 VNB N_VGND_c_1614_n 0.00651182f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_113 VNB N_VGND_c_1615_n 0.00403597f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_114 VNB N_VGND_c_1616_n 0.00596278f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_115 VNB N_VGND_c_1617_n 0.587618f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_116 VPB N_A_55_119#_M1005_g 0.0198688f $X=-0.19 $Y=1.655 $X2=1.995 $Y2=2.755
cc_117 VPB N_A_55_119#_c_229_n 0.0311407f $X=-0.19 $Y=1.655 $X2=0.195 $Y2=2.3
cc_118 VPB N_A_55_119#_c_235_n 0.0245138f $X=-0.19 $Y=1.655 $X2=0.48 $Y2=2.56
cc_119 VPB N_A_55_119#_c_236_n 0.0172998f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=2.385
cc_120 VPB N_A_55_119#_c_231_n 0.0263798f $X=-0.19 $Y=1.655 $X2=1.085 $Y2=1.8
cc_121 VPB N_A_55_119#_c_238_n 0.0163026f $X=-0.19 $Y=1.655 $X2=2.015 $Y2=2.11
cc_122 VPB N_A_55_119#_c_239_n 0.0363526f $X=-0.19 $Y=1.655 $X2=2.015 $Y2=2.11
cc_123 VPB N_A_55_119#_c_240_n 0.00167526f $X=-0.19 $Y=1.655 $X2=1 $Y2=1.945
cc_124 VPB N_D_M1018_g 0.0554059f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_125 VPB N_SCE_c_363_n 0.0196169f $X=-0.19 $Y=1.655 $X2=0.335 $Y2=2.435
cc_126 VPB N_SCE_c_364_n 0.020451f $X=-0.19 $Y=1.655 $X2=1.205 $Y2=1.635
cc_127 VPB N_SCE_c_365_n 0.0253957f $X=-0.19 $Y=1.655 $X2=1.995 $Y2=2.755
cc_128 VPB N_SCE_c_366_n 0.016092f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_129 VPB N_SCE_c_360_n 0.00404552f $X=-0.19 $Y=1.655 $X2=1.125 $Y2=1.945
cc_130 VPB N_SCE_c_368_n 0.0161901f $X=-0.19 $Y=1.655 $X2=1.125 $Y2=1.8
cc_131 VPB N_SCE_c_369_n 0.0124885f $X=-0.19 $Y=1.655 $X2=1.085 $Y2=1.8
cc_132 VPB SCE 0.00706126f $X=-0.19 $Y=1.655 $X2=1.085 $Y2=1.8
cc_133 VPB N_SCD_M1001_g 0.0526767f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_134 VPB SCD 0.00852514f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_135 VPB N_SCD_c_430_n 0.00891619f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_136 VPB N_CLK_M1031_g 0.0388405f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_137 VPB N_CLK_c_480_n 0.0239612f $X=-0.19 $Y=1.655 $X2=1.995 $Y2=2.275
cc_138 VPB N_CLK_c_481_n 0.0312804f $X=-0.19 $Y=1.655 $X2=1.995 $Y2=2.755
cc_139 VPB CLK 0.00741917f $X=-0.19 $Y=1.655 $X2=1.995 $Y2=2.755
cc_140 VPB N_A_610_487#_c_539_n 0.0232422f $X=-0.19 $Y=1.655 $X2=1.995 $Y2=2.275
cc_141 VPB N_A_610_487#_M1011_g 0.0337141f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_142 VPB N_A_610_487#_M1019_g 0.0238688f $X=-0.19 $Y=1.655 $X2=1.125 $Y2=1.8
cc_143 VPB N_A_610_487#_c_528_n 0.059415f $X=-0.19 $Y=1.655 $X2=2.015 $Y2=2.11
cc_144 VPB N_A_610_487#_c_543_n 0.00728249f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_145 VPB N_A_610_487#_c_544_n 0.0113928f $X=-0.19 $Y=1.655 $X2=0.462 $Y2=2.385
cc_146 VPB N_A_610_487#_c_545_n 0.00357272f $X=-0.19 $Y=1.655 $X2=1 $Y2=1.945
cc_147 VPB N_A_610_487#_c_530_n 0.00664666f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_148 VPB N_A_610_487#_c_547_n 0.0319986f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_149 VPB N_A_610_487#_c_548_n 0.0013797f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_150 VPB N_A_610_487#_c_549_n 0.00297982f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_151 VPB N_A_610_487#_c_550_n 0.0021469f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_152 VPB N_A_610_487#_c_551_n 0.00649404f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_153 VPB N_A_610_487#_c_552_n 0.00129583f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_154 VPB N_A_610_487#_c_532_n 0.00221916f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_155 VPB N_A_610_487#_c_536_n 8.85708e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_156 VPB N_A_610_487#_c_555_n 0.0384193f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_157 VPB N_A_610_487#_c_556_n 0.00327944f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_158 VPB N_A_610_487#_c_537_n 0.0226748f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_159 VPB N_A_831_47#_c_780_n 0.00808408f $X=-0.19 $Y=1.655 $X2=1.205 $Y2=0.805
cc_160 VPB N_A_831_47#_c_781_n 0.0394805f $X=-0.19 $Y=1.655 $X2=1.205 $Y2=0.805
cc_161 VPB N_A_831_47#_c_782_n 0.00963269f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_162 VPB N_A_831_47#_c_783_n 0.0205762f $X=-0.19 $Y=1.655 $X2=1.995 $Y2=2.275
cc_163 VPB N_A_831_47#_M1016_g 0.052182f $X=-0.19 $Y=1.655 $X2=1.085 $Y2=1.8
cc_164 VPB N_A_831_47#_c_785_n 0.0164234f $X=-0.19 $Y=1.655 $X2=2.015 $Y2=2.11
cc_165 VPB N_A_831_47#_c_767_n 0.0101405f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_166 VPB N_A_831_47#_c_768_n 0.00163661f $X=-0.19 $Y=1.655 $X2=0.42 $Y2=0.805
cc_167 VPB N_A_1178_399#_c_935_n 0.0259948f $X=-0.19 $Y=1.655 $X2=0.195 $Y2=2.3
cc_168 VPB N_A_1178_399#_c_942_n 0.0454128f $X=-0.19 $Y=1.655 $X2=0.462 $Y2=2.47
cc_169 VPB N_A_1178_399#_c_936_n 0.00458567f $X=-0.19 $Y=1.655 $X2=0.462
+ $Y2=2.56
cc_170 VPB N_A_1178_399#_c_937_n 0.0100006f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_171 VPB N_A_1178_399#_c_945_n 0.00251048f $X=-0.19 $Y=1.655 $X2=0.61
+ $Y2=2.385
cc_172 VPB N_A_1047_125#_M1014_g 0.0491506f $X=-0.19 $Y=1.655 $X2=1.205
+ $Y2=0.805
cc_173 VPB N_A_1047_125#_c_1013_n 0.00308289f $X=-0.19 $Y=1.655 $X2=0.195
+ $Y2=0.97
cc_174 VPB N_A_1047_125#_c_1021_n 0.0027162f $X=-0.19 $Y=1.655 $X2=0.61
+ $Y2=2.385
cc_175 VPB N_A_1047_125#_c_1022_n 0.0063264f $X=-0.19 $Y=1.655 $X2=2.015
+ $Y2=2.11
cc_176 VPB N_A_1665_381#_M1022_g 0.0243723f $X=-0.19 $Y=1.655 $X2=1.205
+ $Y2=0.805
cc_177 VPB N_A_1665_381#_M1028_g 0.0132394f $X=-0.19 $Y=1.655 $X2=1.995
+ $Y2=2.755
cc_178 VPB N_A_1665_381#_M1013_g 0.0221874f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_179 VPB N_A_1665_381#_M1024_g 0.0255345f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_180 VPB N_A_1665_381#_c_1119_n 0.00633239f $X=-0.19 $Y=1.655 $X2=2.015
+ $Y2=2.11
cc_181 VPB N_A_1665_381#_c_1120_n 0.00931335f $X=-0.19 $Y=1.655 $X2=0.462
+ $Y2=2.385
cc_182 VPB N_A_1665_381#_c_1121_n 0.00683224f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_183 VPB N_A_1665_381#_c_1111_n 0.00786655f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_184 VPB N_A_1665_381#_c_1123_n 0.00529195f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_185 VPB N_A_1665_381#_c_1113_n 2.31763e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_186 VPB N_A_1665_381#_c_1125_n 0.0360055f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_187 VPB N_A_1665_381#_c_1114_n 0.0120264f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_188 VPB N_A_1517_63#_M1000_g 0.0271207f $X=-0.19 $Y=1.655 $X2=1.995 $Y2=2.755
cc_189 VPB N_A_1517_63#_c_1211_n 0.0152325f $X=-0.19 $Y=1.655 $X2=0.462 $Y2=2.56
cc_190 VPB N_A_1517_63#_c_1212_n 0.00130493f $X=-0.19 $Y=1.655 $X2=1.25 $Y2=2.11
cc_191 VPB N_A_1517_63#_c_1220_n 0.00517514f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_192 VPB N_A_1517_63#_c_1221_n 0.00291193f $X=-0.19 $Y=1.655 $X2=0.195
+ $Y2=0.805
cc_193 VPB N_A_1517_63#_c_1214_n 0.00861702f $X=-0.19 $Y=1.655 $X2=0.42
+ $Y2=0.805
cc_194 VPB N_A_1517_63#_c_1215_n 0.00267681f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_195 VPB N_VPWR_c_1308_n 0.00631679f $X=-0.19 $Y=1.655 $X2=1.125 $Y2=1.8
cc_196 VPB N_VPWR_c_1309_n 0.00562178f $X=-0.19 $Y=1.655 $X2=1.25 $Y2=2.11
cc_197 VPB N_VPWR_c_1310_n 0.0197316f $X=-0.19 $Y=1.655 $X2=2.015 $Y2=2.11
cc_198 VPB N_VPWR_c_1311_n 0.0118301f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_199 VPB N_VPWR_c_1312_n 0.0116949f $X=-0.19 $Y=1.655 $X2=0.195 $Y2=2.385
cc_200 VPB N_VPWR_c_1313_n 0.0131805f $X=-0.19 $Y=1.655 $X2=1.085 $Y2=1.8
cc_201 VPB N_VPWR_c_1314_n 0.0145625f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_202 VPB N_VPWR_c_1315_n 0.0112949f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_203 VPB N_VPWR_c_1316_n 0.0585851f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_204 VPB N_VPWR_c_1317_n 0.024208f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_205 VPB N_VPWR_c_1318_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_206 VPB N_VPWR_c_1319_n 0.0574825f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_207 VPB N_VPWR_c_1320_n 0.00535984f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_208 VPB N_VPWR_c_1321_n 0.0427666f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_209 VPB N_VPWR_c_1322_n 0.0563127f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_210 VPB N_VPWR_c_1323_n 0.0179602f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_211 VPB N_VPWR_c_1324_n 0.0150561f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_212 VPB N_VPWR_c_1325_n 0.00420575f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_213 VPB N_VPWR_c_1326_n 0.0047828f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_214 VPB N_VPWR_c_1327_n 0.0129576f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_215 VPB N_VPWR_c_1328_n 0.00484208f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_216 VPB N_VPWR_c_1307_n 0.126303f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_217 VPB N_A_328_119#_c_1453_n 0.0050896f $X=-0.19 $Y=1.655 $X2=1.125
+ $Y2=1.945
cc_218 VPB N_A_328_119#_c_1454_n 0.00321318f $X=-0.19 $Y=1.655 $X2=1.125 $Y2=1.8
cc_219 VPB N_A_328_119#_c_1450_n 0.00271698f $X=-0.19 $Y=1.655 $X2=1.085 $Y2=1.8
cc_220 VPB N_A_328_119#_c_1452_n 0.00718361f $X=-0.19 $Y=1.655 $X2=1.25 $Y2=2.11
cc_221 VPB N_A_328_119#_c_1457_n 0.00120685f $X=-0.19 $Y=1.655 $X2=2.015
+ $Y2=2.11
cc_222 VPB N_A_328_119#_c_1458_n 0.0136945f $X=-0.19 $Y=1.655 $X2=0.42 $Y2=0.805
cc_223 VPB N_A_328_119#_c_1459_n 8.59522e-19 $X=-0.19 $Y=1.655 $X2=0.42
+ $Y2=0.805
cc_224 VPB N_A_328_119#_c_1460_n 0.00541849f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_225 VPB N_A_328_119#_c_1461_n 0.00259008f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_226 VPB Q 0.0029492f $X=-0.19 $Y=1.655 $X2=1.205 $Y2=1.635
cc_227 N_A_55_119#_M1005_g N_D_M1018_g 0.0140934f $X=1.995 $Y=2.755 $X2=0 $Y2=0
cc_228 N_A_55_119#_c_230_n N_D_M1018_g 0.0019693f $X=1.085 $Y=1.8 $X2=0 $Y2=0
cc_229 N_A_55_119#_c_231_n N_D_M1018_g 0.0100355f $X=1.085 $Y=1.8 $X2=0 $Y2=0
cc_230 N_A_55_119#_c_238_n N_D_M1018_g 0.023429f $X=2.015 $Y=2.11 $X2=0 $Y2=0
cc_231 N_A_55_119#_c_239_n N_D_M1018_g 0.021335f $X=2.015 $Y=2.11 $X2=0 $Y2=0
cc_232 N_A_55_119#_c_240_n N_D_M1018_g 9.39703e-19 $X=1 $Y=1.945 $X2=0 $Y2=0
cc_233 N_A_55_119#_M1007_g D 0.0319129f $X=1.205 $Y=0.805 $X2=0 $Y2=0
cc_234 N_A_55_119#_c_230_n D 0.0107826f $X=1.085 $Y=1.8 $X2=0 $Y2=0
cc_235 N_A_55_119#_c_238_n D 0.0197429f $X=2.015 $Y=2.11 $X2=0 $Y2=0
cc_236 N_A_55_119#_c_231_n N_D_c_316_n 0.0424878f $X=1.085 $Y=1.8 $X2=0 $Y2=0
cc_237 N_A_55_119#_c_238_n N_D_c_316_n 0.0023618f $X=2.015 $Y=2.11 $X2=0 $Y2=0
cc_238 N_A_55_119#_M1007_g N_D_c_317_n 0.0424878f $X=1.205 $Y=0.805 $X2=0 $Y2=0
cc_239 N_A_55_119#_c_229_n N_SCE_c_363_n 0.00760356f $X=0.195 $Y=2.3 $X2=0 $Y2=0
cc_240 N_A_55_119#_c_231_n N_SCE_c_363_n 0.00438282f $X=1.085 $Y=1.8 $X2=0 $Y2=0
cc_241 N_A_55_119#_c_240_n N_SCE_c_363_n 0.00250258f $X=1 $Y=1.945 $X2=0 $Y2=0
cc_242 N_A_55_119#_M1007_g N_SCE_M1008_g 0.023975f $X=1.205 $Y=0.805 $X2=0 $Y2=0
cc_243 N_A_55_119#_c_229_n N_SCE_M1008_g 0.00509765f $X=0.195 $Y=2.3 $X2=0 $Y2=0
cc_244 N_A_55_119#_c_258_p N_SCE_c_364_n 0.0101881f $X=1 $Y=2.385 $X2=0 $Y2=0
cc_245 N_A_55_119#_M1007_g N_SCE_c_357_n 0.00886244f $X=1.205 $Y=0.805 $X2=0
+ $Y2=0
cc_246 N_A_55_119#_c_258_p N_SCE_c_365_n 0.00797451f $X=1 $Y=2.385 $X2=0 $Y2=0
cc_247 N_A_55_119#_c_231_n N_SCE_c_365_n 0.0223217f $X=1.085 $Y=1.8 $X2=0 $Y2=0
cc_248 N_A_55_119#_c_238_n N_SCE_c_365_n 0.00289614f $X=2.015 $Y=2.11 $X2=0
+ $Y2=0
cc_249 N_A_55_119#_c_240_n N_SCE_c_365_n 0.016824f $X=1 $Y=1.945 $X2=0 $Y2=0
cc_250 N_A_55_119#_c_240_n N_SCE_c_366_n 0.00603805f $X=1 $Y=1.945 $X2=0 $Y2=0
cc_251 N_A_55_119#_c_230_n N_SCE_c_360_n 2.14219e-19 $X=1.085 $Y=1.8 $X2=0 $Y2=0
cc_252 N_A_55_119#_c_231_n N_SCE_c_360_n 0.0151913f $X=1.085 $Y=1.8 $X2=0 $Y2=0
cc_253 N_A_55_119#_c_236_n N_SCE_c_368_n 0.0025538f $X=0.61 $Y=2.385 $X2=0 $Y2=0
cc_254 N_A_55_119#_c_235_n N_SCE_c_369_n 4.15226e-19 $X=0.48 $Y=2.56 $X2=0 $Y2=0
cc_255 N_A_55_119#_c_258_p N_SCE_c_369_n 0.00220199f $X=1 $Y=2.385 $X2=0 $Y2=0
cc_256 N_A_55_119#_c_236_n N_SCE_c_369_n 0.00315535f $X=0.61 $Y=2.385 $X2=0
+ $Y2=0
cc_257 N_A_55_119#_M1007_g SCE 0.0052521f $X=1.205 $Y=0.805 $X2=0 $Y2=0
cc_258 N_A_55_119#_c_229_n SCE 0.0764783f $X=0.195 $Y=2.3 $X2=0 $Y2=0
cc_259 N_A_55_119#_c_236_n SCE 0.0300504f $X=0.61 $Y=2.385 $X2=0 $Y2=0
cc_260 N_A_55_119#_c_230_n SCE 0.0242882f $X=1.085 $Y=1.8 $X2=0 $Y2=0
cc_261 N_A_55_119#_c_231_n SCE 0.00226971f $X=1.085 $Y=1.8 $X2=0 $Y2=0
cc_262 N_A_55_119#_c_232_n SCE 0.00694649f $X=0.42 $Y=0.805 $X2=0 $Y2=0
cc_263 N_A_55_119#_c_240_n SCE 0.0164401f $X=1 $Y=1.945 $X2=0 $Y2=0
cc_264 N_A_55_119#_c_229_n N_SCE_c_362_n 0.0162737f $X=0.195 $Y=2.3 $X2=0 $Y2=0
cc_265 N_A_55_119#_c_232_n N_SCE_c_362_n 0.00341357f $X=0.42 $Y=0.805 $X2=0
+ $Y2=0
cc_266 N_A_55_119#_M1005_g N_SCD_M1001_g 0.0344379f $X=1.995 $Y=2.755 $X2=0
+ $Y2=0
cc_267 N_A_55_119#_c_238_n N_SCD_M1001_g 2.99193e-19 $X=2.015 $Y=2.11 $X2=0
+ $Y2=0
cc_268 N_A_55_119#_c_239_n N_SCD_M1001_g 0.0204068f $X=2.015 $Y=2.11 $X2=0 $Y2=0
cc_269 N_A_55_119#_c_238_n SCD 0.00631569f $X=2.015 $Y=2.11 $X2=0 $Y2=0
cc_270 N_A_55_119#_c_239_n SCD 0.00380896f $X=2.015 $Y=2.11 $X2=0 $Y2=0
cc_271 N_A_55_119#_c_258_p N_VPWR_M1029_d 0.00180618f $X=1 $Y=2.385 $X2=-0.19
+ $Y2=-0.245
cc_272 N_A_55_119#_c_240_n N_VPWR_M1029_d 7.98001e-19 $X=1 $Y=1.945 $X2=-0.19
+ $Y2=-0.245
cc_273 N_A_55_119#_c_258_p N_VPWR_c_1308_n 0.0137545f $X=1 $Y=2.385 $X2=0 $Y2=0
cc_274 N_A_55_119#_c_240_n N_VPWR_c_1308_n 0.00643497f $X=1 $Y=1.945 $X2=0 $Y2=0
cc_275 N_A_55_119#_c_235_n N_VPWR_c_1317_n 0.018877f $X=0.48 $Y=2.56 $X2=0 $Y2=0
cc_276 N_A_55_119#_M1005_g N_VPWR_c_1321_n 0.00405136f $X=1.995 $Y=2.755 $X2=0
+ $Y2=0
cc_277 N_A_55_119#_M1005_g N_VPWR_c_1307_n 0.00593005f $X=1.995 $Y=2.755 $X2=0
+ $Y2=0
cc_278 N_A_55_119#_c_235_n N_VPWR_c_1307_n 0.0113564f $X=0.48 $Y=2.56 $X2=0
+ $Y2=0
cc_279 N_A_55_119#_c_258_p N_VPWR_c_1307_n 6.80523e-19 $X=1 $Y=2.385 $X2=0 $Y2=0
cc_280 N_A_55_119#_c_236_n N_VPWR_c_1307_n 0.0117121f $X=0.61 $Y=2.385 $X2=0
+ $Y2=0
cc_281 N_A_55_119#_c_240_n N_VPWR_c_1307_n 0.00244199f $X=1 $Y=1.945 $X2=0 $Y2=0
cc_282 N_A_55_119#_M1005_g N_A_328_119#_c_1462_n 0.00958872f $X=1.995 $Y=2.755
+ $X2=0 $Y2=0
cc_283 N_A_55_119#_c_238_n N_A_328_119#_c_1462_n 0.0106876f $X=2.015 $Y=2.11
+ $X2=0 $Y2=0
cc_284 N_A_55_119#_c_239_n N_A_328_119#_c_1462_n 0.00261661f $X=2.015 $Y=2.11
+ $X2=0 $Y2=0
cc_285 N_A_55_119#_c_238_n N_A_328_119#_c_1449_n 0.00300212f $X=2.015 $Y=2.11
+ $X2=0 $Y2=0
cc_286 N_A_55_119#_c_239_n N_A_328_119#_c_1449_n 0.00200612f $X=2.015 $Y=2.11
+ $X2=0 $Y2=0
cc_287 N_A_55_119#_c_238_n N_A_328_119#_c_1454_n 0.0151549f $X=2.015 $Y=2.11
+ $X2=0 $Y2=0
cc_288 N_A_55_119#_c_239_n N_A_328_119#_c_1454_n 0.00118566f $X=2.015 $Y=2.11
+ $X2=0 $Y2=0
cc_289 N_A_55_119#_M1005_g N_A_328_119#_c_1457_n 0.0090591f $X=1.995 $Y=2.755
+ $X2=0 $Y2=0
cc_290 N_A_55_119#_c_238_n N_A_328_119#_c_1457_n 0.02267f $X=2.015 $Y=2.11 $X2=0
+ $Y2=0
cc_291 N_A_55_119#_c_239_n N_A_328_119#_c_1457_n 0.00145582f $X=2.015 $Y=2.11
+ $X2=0 $Y2=0
cc_292 N_A_55_119#_c_240_n N_A_328_119#_c_1457_n 9.65141e-19 $X=1 $Y=1.945 $X2=0
+ $Y2=0
cc_293 N_A_55_119#_M1005_g N_A_328_119#_c_1460_n 0.00405675f $X=1.995 $Y=2.755
+ $X2=0 $Y2=0
cc_294 N_A_55_119#_c_238_n N_A_328_119#_c_1460_n 0.0131642f $X=2.015 $Y=2.11
+ $X2=0 $Y2=0
cc_295 N_A_55_119#_c_239_n N_A_328_119#_c_1460_n 0.00104107f $X=2.015 $Y=2.11
+ $X2=0 $Y2=0
cc_296 N_A_55_119#_M1007_g N_VGND_c_1596_n 0.00180401f $X=1.205 $Y=0.805 $X2=0
+ $Y2=0
cc_297 N_A_55_119#_c_231_n N_VGND_c_1596_n 6.40196e-19 $X=1.085 $Y=1.8 $X2=0
+ $Y2=0
cc_298 N_A_55_119#_c_232_n N_VGND_c_1605_n 0.00774495f $X=0.42 $Y=0.805 $X2=0
+ $Y2=0
cc_299 N_A_55_119#_c_232_n N_VGND_c_1617_n 0.0130121f $X=0.42 $Y=0.805 $X2=0
+ $Y2=0
cc_300 D N_SCE_M1008_g 0.00428957f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_301 D N_SCE_c_357_n 0.0105633f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_302 N_D_c_317_n N_SCE_c_357_n 0.00886244f $X=1.655 $Y=1.125 $X2=0 $Y2=0
cc_303 N_D_M1018_g N_SCE_c_365_n 0.0628746f $X=1.565 $Y=2.755 $X2=0 $Y2=0
cc_304 D N_SCE_M1017_g 0.00716974f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_305 N_D_c_316_n N_SCE_M1017_g 6.23435e-19 $X=1.655 $Y=1.29 $X2=0 $Y2=0
cc_306 N_D_c_317_n N_SCE_M1017_g 0.00769648f $X=1.655 $Y=1.125 $X2=0 $Y2=0
cc_307 N_D_M1018_g SCE 4.79853e-19 $X=1.565 $Y=2.755 $X2=0 $Y2=0
cc_308 D SCE 0.0195009f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_309 N_D_c_316_n N_SCD_M1009_g 0.00332848f $X=1.655 $Y=1.29 $X2=0 $Y2=0
cc_310 N_D_M1018_g SCD 0.00814246f $X=1.565 $Y=2.755 $X2=0 $Y2=0
cc_311 N_D_M1018_g N_SCD_c_430_n 0.00240956f $X=1.565 $Y=2.755 $X2=0 $Y2=0
cc_312 D N_SCD_c_430_n 4.25105e-19 $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_313 N_D_c_316_n N_SCD_c_430_n 0.00210068f $X=1.655 $Y=1.29 $X2=0 $Y2=0
cc_314 N_D_M1018_g N_VPWR_c_1321_n 0.00529818f $X=1.565 $Y=2.755 $X2=0 $Y2=0
cc_315 N_D_M1018_g N_VPWR_c_1307_n 0.00975072f $X=1.565 $Y=2.755 $X2=0 $Y2=0
cc_316 D N_A_328_119#_M1004_d 0.00429435f $X=1.115 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_317 D N_A_328_119#_c_1447_n 0.039432f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_318 N_D_c_317_n N_A_328_119#_c_1447_n 0.00137824f $X=1.655 $Y=1.125 $X2=0
+ $Y2=0
cc_319 D N_A_328_119#_c_1449_n 0.0150804f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_320 N_D_c_316_n N_A_328_119#_c_1449_n 0.00199586f $X=1.655 $Y=1.29 $X2=0
+ $Y2=0
cc_321 N_D_M1018_g N_A_328_119#_c_1457_n 0.0113301f $X=1.565 $Y=2.755 $X2=0
+ $Y2=0
cc_322 D N_VGND_c_1596_n 0.0320145f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_323 D N_VGND_c_1607_n 0.0253171f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_324 D N_VGND_c_1617_n 0.0208218f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_325 N_SCE_M1017_g N_SCD_M1009_g 0.0408067f $X=2.245 $Y=0.805 $X2=0 $Y2=0
cc_326 N_SCE_M1017_g SCD 7.78388e-19 $X=2.245 $Y=0.805 $X2=0 $Y2=0
cc_327 N_SCE_c_364_n N_VPWR_c_1308_n 0.00387218f $X=0.695 $Y=2.325 $X2=0 $Y2=0
cc_328 N_SCE_c_365_n N_VPWR_c_1308_n 0.0010287f $X=1.13 $Y=2.25 $X2=0 $Y2=0
cc_329 N_SCE_c_366_n N_VPWR_c_1308_n 0.00379803f $X=1.205 $Y=2.325 $X2=0 $Y2=0
cc_330 N_SCE_c_364_n N_VPWR_c_1317_n 0.00565115f $X=0.695 $Y=2.325 $X2=0 $Y2=0
cc_331 N_SCE_c_366_n N_VPWR_c_1321_n 0.00565115f $X=1.205 $Y=2.325 $X2=0 $Y2=0
cc_332 N_SCE_c_364_n N_VPWR_c_1307_n 0.00730004f $X=0.695 $Y=2.325 $X2=0 $Y2=0
cc_333 N_SCE_c_366_n N_VPWR_c_1307_n 0.00940631f $X=1.205 $Y=2.325 $X2=0 $Y2=0
cc_334 N_SCE_c_357_n N_A_328_119#_c_1447_n 0.00277252f $X=2.17 $Y=0.18 $X2=0
+ $Y2=0
cc_335 N_SCE_M1017_g N_A_328_119#_c_1447_n 0.00290323f $X=2.245 $Y=0.805 $X2=0
+ $Y2=0
cc_336 N_SCE_M1017_g N_A_328_119#_c_1448_n 0.0102129f $X=2.245 $Y=0.805 $X2=0
+ $Y2=0
cc_337 N_SCE_c_366_n N_A_328_119#_c_1457_n 0.00212409f $X=1.205 $Y=2.325 $X2=0
+ $Y2=0
cc_338 N_SCE_M1008_g N_VGND_c_1596_n 0.0125111f $X=0.635 $Y=0.805 $X2=0 $Y2=0
cc_339 N_SCE_c_357_n N_VGND_c_1596_n 0.0174837f $X=2.17 $Y=0.18 $X2=0 $Y2=0
cc_340 SCE N_VGND_c_1596_n 0.00762044f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_341 N_SCE_c_357_n N_VGND_c_1597_n 0.0104863f $X=2.17 $Y=0.18 $X2=0 $Y2=0
cc_342 N_SCE_c_358_n N_VGND_c_1605_n 0.0064002f $X=0.71 $Y=0.18 $X2=0 $Y2=0
cc_343 N_SCE_c_357_n N_VGND_c_1607_n 0.0385467f $X=2.17 $Y=0.18 $X2=0 $Y2=0
cc_344 N_SCE_c_357_n N_VGND_c_1617_n 0.0539738f $X=2.17 $Y=0.18 $X2=0 $Y2=0
cc_345 N_SCE_c_358_n N_VGND_c_1617_n 0.0110282f $X=0.71 $Y=0.18 $X2=0 $Y2=0
cc_346 N_SCD_M1009_g N_CLK_M1023_g 0.012838f $X=2.605 $Y=0.805 $X2=0 $Y2=0
cc_347 N_SCD_M1001_g N_CLK_c_480_n 0.00429345f $X=2.465 $Y=2.755 $X2=0 $Y2=0
cc_348 N_SCD_M1001_g N_CLK_c_481_n 0.0325457f $X=2.465 $Y=2.755 $X2=0 $Y2=0
cc_349 SCD N_CLK_c_478_n 9.93011e-19 $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_350 N_SCD_c_430_n N_CLK_c_478_n 0.012838f $X=2.515 $Y=1.54 $X2=0 $Y2=0
cc_351 N_SCD_M1001_g N_A_610_487#_c_543_n 7.17552e-19 $X=2.465 $Y=2.755 $X2=0
+ $Y2=0
cc_352 N_SCD_M1001_g N_A_610_487#_c_545_n 2.24983e-19 $X=2.465 $Y=2.755 $X2=0
+ $Y2=0
cc_353 N_SCD_M1001_g N_VPWR_c_1309_n 0.0123798f $X=2.465 $Y=2.755 $X2=0 $Y2=0
cc_354 N_SCD_M1001_g N_VPWR_c_1321_n 0.00500222f $X=2.465 $Y=2.755 $X2=0 $Y2=0
cc_355 N_SCD_M1001_g N_VPWR_c_1307_n 0.00636283f $X=2.465 $Y=2.755 $X2=0 $Y2=0
cc_356 N_SCD_M1001_g N_A_328_119#_c_1462_n 0.0107911f $X=2.465 $Y=2.755 $X2=0
+ $Y2=0
cc_357 SCD N_A_328_119#_c_1462_n 0.00475847f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_358 N_SCD_M1009_g N_A_328_119#_c_1448_n 0.0163316f $X=2.605 $Y=0.805 $X2=0
+ $Y2=0
cc_359 SCD N_A_328_119#_c_1448_n 0.0447059f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_360 N_SCD_c_430_n N_A_328_119#_c_1448_n 0.00503823f $X=2.515 $Y=1.54 $X2=0
+ $Y2=0
cc_361 SCD N_A_328_119#_c_1449_n 0.0087955f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_362 N_SCD_M1001_g N_A_328_119#_c_1454_n 0.00777866f $X=2.465 $Y=2.755 $X2=0
+ $Y2=0
cc_363 SCD N_A_328_119#_c_1454_n 0.0358032f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_364 N_SCD_c_430_n N_A_328_119#_c_1454_n 0.00115729f $X=2.515 $Y=1.54 $X2=0
+ $Y2=0
cc_365 N_SCD_M1001_g N_A_328_119#_c_1450_n 0.0032767f $X=2.465 $Y=2.755 $X2=0
+ $Y2=0
cc_366 N_SCD_M1009_g N_A_328_119#_c_1450_n 0.0034931f $X=2.605 $Y=0.805 $X2=0
+ $Y2=0
cc_367 SCD N_A_328_119#_c_1450_n 0.0258176f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_368 N_SCD_c_430_n N_A_328_119#_c_1450_n 7.60996e-19 $X=2.515 $Y=1.54 $X2=0
+ $Y2=0
cc_369 N_SCD_M1001_g N_A_328_119#_c_1457_n 0.00205794f $X=2.465 $Y=2.755 $X2=0
+ $Y2=0
cc_370 N_SCD_M1001_g N_A_328_119#_c_1459_n 0.00193606f $X=2.465 $Y=2.755 $X2=0
+ $Y2=0
cc_371 SCD N_A_328_119#_c_1459_n 8.9813e-19 $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_372 N_SCD_M1001_g N_A_328_119#_c_1460_n 0.00965657f $X=2.465 $Y=2.755 $X2=0
+ $Y2=0
cc_373 N_SCD_M1009_g N_VGND_c_1597_n 0.00392993f $X=2.605 $Y=0.805 $X2=0 $Y2=0
cc_374 N_SCD_M1009_g N_VGND_c_1607_n 0.00431487f $X=2.605 $Y=0.805 $X2=0 $Y2=0
cc_375 N_SCD_M1009_g N_VGND_c_1617_n 0.00477801f $X=2.605 $Y=0.805 $X2=0 $Y2=0
cc_376 CLK N_A_610_487#_M1032_g 0.00134903f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_377 N_CLK_c_480_n N_A_610_487#_c_528_n 0.011862f $X=3.202 $Y=1.945 $X2=0
+ $Y2=0
cc_378 N_CLK_M1031_g N_A_610_487#_c_543_n 0.00751422f $X=2.975 $Y=2.755 $X2=0
+ $Y2=0
cc_379 N_CLK_M1023_g N_A_610_487#_c_529_n 6.46038e-19 $X=3.125 $Y=0.805 $X2=0
+ $Y2=0
cc_380 CLK N_A_610_487#_c_529_n 0.0422841f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_381 N_CLK_c_478_n N_A_610_487#_c_529_n 0.00216518f $X=3.34 $Y=1.59 $X2=0
+ $Y2=0
cc_382 N_CLK_c_481_n N_A_610_487#_c_544_n 9.61242e-19 $X=3.202 $Y=2.095 $X2=0
+ $Y2=0
cc_383 CLK N_A_610_487#_c_544_n 0.0275105f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_384 N_CLK_M1031_g N_A_610_487#_c_545_n 0.00529442f $X=2.975 $Y=2.755 $X2=0
+ $Y2=0
cc_385 N_CLK_c_481_n N_A_610_487#_c_545_n 0.00931384f $X=3.202 $Y=2.095 $X2=0
+ $Y2=0
cc_386 CLK N_A_610_487#_c_545_n 0.00807478f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_387 CLK N_A_610_487#_c_530_n 0.0743043f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_388 N_CLK_c_478_n N_A_610_487#_c_530_n 5.30074e-19 $X=3.34 $Y=1.59 $X2=0
+ $Y2=0
cc_389 CLK N_A_610_487#_c_531_n 0.0057211f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_390 N_CLK_c_478_n N_A_610_487#_c_531_n 0.011862f $X=3.34 $Y=1.59 $X2=0 $Y2=0
cc_391 N_CLK_M1031_g N_VPWR_c_1309_n 0.00298127f $X=2.975 $Y=2.755 $X2=0 $Y2=0
cc_392 N_CLK_M1031_g N_VPWR_c_1310_n 0.00531373f $X=2.975 $Y=2.755 $X2=0 $Y2=0
cc_393 N_CLK_M1031_g N_VPWR_c_1311_n 0.00276607f $X=2.975 $Y=2.755 $X2=0 $Y2=0
cc_394 N_CLK_M1031_g N_VPWR_c_1307_n 0.0111439f $X=2.975 $Y=2.755 $X2=0 $Y2=0
cc_395 N_CLK_M1031_g N_A_328_119#_c_1462_n 9.48441e-19 $X=2.975 $Y=2.755 $X2=0
+ $Y2=0
cc_396 N_CLK_M1023_g N_A_328_119#_c_1448_n 0.00865939f $X=3.125 $Y=0.805 $X2=0
+ $Y2=0
cc_397 CLK N_A_328_119#_c_1448_n 0.00702775f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_398 N_CLK_M1031_g N_A_328_119#_c_1453_n 0.00365821f $X=2.975 $Y=2.755 $X2=0
+ $Y2=0
cc_399 N_CLK_c_481_n N_A_328_119#_c_1453_n 0.0069929f $X=3.202 $Y=2.095 $X2=0
+ $Y2=0
cc_400 CLK N_A_328_119#_c_1453_n 0.0135426f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_401 N_CLK_M1023_g N_A_328_119#_c_1450_n 0.00278718f $X=3.125 $Y=0.805 $X2=0
+ $Y2=0
cc_402 N_CLK_c_480_n N_A_328_119#_c_1450_n 0.00798191f $X=3.202 $Y=1.945 $X2=0
+ $Y2=0
cc_403 N_CLK_c_481_n N_A_328_119#_c_1450_n 0.00368309f $X=3.202 $Y=2.095 $X2=0
+ $Y2=0
cc_404 CLK N_A_328_119#_c_1450_n 0.0471363f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_405 N_CLK_c_478_n N_A_328_119#_c_1450_n 0.00579954f $X=3.34 $Y=1.59 $X2=0
+ $Y2=0
cc_406 N_CLK_M1031_g N_A_328_119#_c_1458_n 0.00746626f $X=2.975 $Y=2.755 $X2=0
+ $Y2=0
cc_407 CLK N_A_328_119#_c_1458_n 0.00378238f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_408 N_CLK_M1031_g N_A_328_119#_c_1459_n 0.0014777f $X=2.975 $Y=2.755 $X2=0
+ $Y2=0
cc_409 N_CLK_M1031_g N_A_328_119#_c_1460_n 0.00548623f $X=2.975 $Y=2.755 $X2=0
+ $Y2=0
cc_410 N_CLK_M1023_g N_VGND_c_1597_n 0.00304762f $X=3.125 $Y=0.805 $X2=0 $Y2=0
cc_411 N_CLK_M1023_g N_VGND_c_1598_n 0.0010895f $X=3.125 $Y=0.805 $X2=0 $Y2=0
cc_412 N_CLK_M1023_g N_VGND_c_1609_n 0.00431487f $X=3.125 $Y=0.805 $X2=0 $Y2=0
cc_413 N_CLK_M1023_g N_VGND_c_1617_n 0.00477801f $X=3.125 $Y=0.805 $X2=0 $Y2=0
cc_414 N_A_610_487#_c_547_n N_A_831_47#_M1006_d 0.00281332f $X=5.675 $Y=2.92
+ $X2=0 $Y2=0
cc_415 N_A_610_487#_c_528_n N_A_831_47#_c_780_n 0.00641574f $X=3.99 $Y=2.085
+ $X2=0 $Y2=0
cc_416 N_A_610_487#_c_530_n N_A_831_47#_c_780_n 2.57906e-19 $X=3.99 $Y=1.59
+ $X2=0 $Y2=0
cc_417 N_A_610_487#_M1011_g N_A_831_47#_c_781_n 0.0170084f $X=5.605 $Y=2.465
+ $X2=0 $Y2=0
cc_418 N_A_610_487#_c_537_n N_A_831_47#_c_781_n 0.0098848f $X=5.605 $Y=1.59
+ $X2=0 $Y2=0
cc_419 N_A_610_487#_c_528_n N_A_831_47#_c_782_n 0.00260659f $X=3.99 $Y=2.085
+ $X2=0 $Y2=0
cc_420 N_A_610_487#_c_547_n N_A_831_47#_c_782_n 0.00393176f $X=5.675 $Y=2.92
+ $X2=0 $Y2=0
cc_421 N_A_610_487#_c_547_n N_A_831_47#_c_783_n 0.00669047f $X=5.675 $Y=2.92
+ $X2=0 $Y2=0
cc_422 N_A_610_487#_c_550_n N_A_831_47#_c_783_n 8.66444e-19 $X=5.76 $Y=2.835
+ $X2=0 $Y2=0
cc_423 N_A_610_487#_c_533_n N_A_831_47#_c_762_n 0.00629299f $X=8.02 $Y=1.36
+ $X2=0 $Y2=0
cc_424 N_A_610_487#_c_585_p N_A_831_47#_c_762_n 0.00480691f $X=7.635 $Y=1.36
+ $X2=0 $Y2=0
cc_425 N_A_610_487#_c_534_n N_A_831_47#_c_762_n 0.00378873f $X=8.185 $Y=1.01
+ $X2=0 $Y2=0
cc_426 N_A_610_487#_c_533_n N_A_831_47#_c_763_n 0.0111434f $X=8.02 $Y=1.36 $X2=0
+ $Y2=0
cc_427 N_A_610_487#_c_535_n N_A_831_47#_c_763_n 0.00619375f $X=8.185 $Y=1.01
+ $X2=0 $Y2=0
cc_428 N_A_610_487#_c_532_n N_A_831_47#_c_764_n 0.00724954f $X=7.55 $Y=1.835
+ $X2=0 $Y2=0
cc_429 N_A_610_487#_c_533_n N_A_831_47#_c_764_n 0.0068713f $X=8.02 $Y=1.36 $X2=0
+ $Y2=0
cc_430 N_A_610_487#_c_585_p N_A_831_47#_c_764_n 0.00128885f $X=7.635 $Y=1.36
+ $X2=0 $Y2=0
cc_431 N_A_610_487#_c_555_n N_A_831_47#_c_764_n 0.0117242f $X=7.465 $Y=1.93
+ $X2=0 $Y2=0
cc_432 N_A_610_487#_c_556_n N_A_831_47#_c_764_n 2.84171e-19 $X=7.55 $Y=1.95
+ $X2=0 $Y2=0
cc_433 N_A_610_487#_M1019_g N_A_831_47#_M1016_g 0.0172615f $X=7.515 $Y=2.675
+ $X2=0 $Y2=0
cc_434 N_A_610_487#_c_552_n N_A_831_47#_M1016_g 5.07137e-19 $X=7.38 $Y=2.745
+ $X2=0 $Y2=0
cc_435 N_A_610_487#_c_532_n N_A_831_47#_M1016_g 0.00368051f $X=7.55 $Y=1.835
+ $X2=0 $Y2=0
cc_436 N_A_610_487#_c_555_n N_A_831_47#_M1016_g 0.011739f $X=7.465 $Y=1.93 $X2=0
+ $Y2=0
cc_437 N_A_610_487#_c_556_n N_A_831_47#_M1016_g 6.05019e-19 $X=7.55 $Y=1.95
+ $X2=0 $Y2=0
cc_438 N_A_610_487#_c_531_n N_A_831_47#_c_785_n 0.0204446f $X=3.99 $Y=1.59 $X2=0
+ $Y2=0
cc_439 N_A_610_487#_c_537_n N_A_831_47#_c_785_n 0.00711564f $X=5.605 $Y=1.59
+ $X2=0 $Y2=0
cc_440 N_A_610_487#_c_531_n N_A_831_47#_c_766_n 0.0059912f $X=3.99 $Y=1.59 $X2=0
+ $Y2=0
cc_441 N_A_610_487#_c_528_n N_A_831_47#_c_767_n 0.0114191f $X=3.99 $Y=2.085
+ $X2=0 $Y2=0
cc_442 N_A_610_487#_c_603_p N_A_831_47#_c_767_n 0.00665878f $X=4.06 $Y=2.835
+ $X2=0 $Y2=0
cc_443 N_A_610_487#_c_547_n N_A_831_47#_c_767_n 0.0219518f $X=5.675 $Y=2.92
+ $X2=0 $Y2=0
cc_444 N_A_610_487#_c_605_p N_A_831_47#_c_767_n 0.0099866f $X=4.025 $Y=2.385
+ $X2=0 $Y2=0
cc_445 N_A_610_487#_M1032_g N_A_831_47#_c_768_n 0.0204446f $X=4.08 $Y=0.445
+ $X2=0 $Y2=0
cc_446 N_A_610_487#_M1012_g N_A_831_47#_c_768_n 0.00711564f $X=5.16 $Y=0.835
+ $X2=0 $Y2=0
cc_447 N_A_610_487#_c_530_n N_A_831_47#_c_768_n 7.476e-19 $X=3.99 $Y=1.59 $X2=0
+ $Y2=0
cc_448 N_A_610_487#_M1012_g N_A_831_47#_c_769_n 0.00637649f $X=5.16 $Y=0.835
+ $X2=0 $Y2=0
cc_449 N_A_610_487#_M1012_g N_A_831_47#_c_770_n 0.00132716f $X=5.16 $Y=0.835
+ $X2=0 $Y2=0
cc_450 N_A_610_487#_M1012_g N_A_831_47#_c_771_n 8.01841e-19 $X=5.16 $Y=0.835
+ $X2=0 $Y2=0
cc_451 N_A_610_487#_c_538_n N_A_831_47#_c_772_n 0.00178565f $X=8.185 $Y=0.845
+ $X2=0 $Y2=0
cc_452 N_A_610_487#_c_533_n N_A_831_47#_c_774_n 0.0115335f $X=8.02 $Y=1.36 $X2=0
+ $Y2=0
cc_453 N_A_610_487#_c_585_p N_A_831_47#_c_774_n 0.0134599f $X=7.635 $Y=1.36
+ $X2=0 $Y2=0
cc_454 N_A_610_487#_c_534_n N_A_831_47#_c_774_n 0.0148564f $X=8.185 $Y=1.01
+ $X2=0 $Y2=0
cc_455 N_A_610_487#_c_535_n N_A_831_47#_c_774_n 8.96194e-19 $X=8.185 $Y=1.01
+ $X2=0 $Y2=0
cc_456 N_A_610_487#_c_538_n N_A_831_47#_c_774_n 0.00348955f $X=8.185 $Y=0.845
+ $X2=0 $Y2=0
cc_457 N_A_610_487#_c_534_n N_A_831_47#_c_775_n 0.00147886f $X=8.185 $Y=1.01
+ $X2=0 $Y2=0
cc_458 N_A_610_487#_c_535_n N_A_831_47#_c_775_n 0.0191321f $X=8.185 $Y=1.01
+ $X2=0 $Y2=0
cc_459 N_A_610_487#_M1012_g N_A_831_47#_c_776_n 0.0035956f $X=5.16 $Y=0.835
+ $X2=0 $Y2=0
cc_460 N_A_610_487#_M1032_g N_A_831_47#_c_777_n 0.0059912f $X=4.08 $Y=0.445
+ $X2=0 $Y2=0
cc_461 N_A_610_487#_c_529_n N_A_831_47#_c_777_n 0.0212735f $X=3.74 $Y=0.865
+ $X2=0 $Y2=0
cc_462 N_A_610_487#_c_530_n N_A_831_47#_c_777_n 0.0971382f $X=3.99 $Y=1.59 $X2=0
+ $Y2=0
cc_463 N_A_610_487#_M1012_g N_A_831_47#_c_778_n 0.0135686f $X=5.16 $Y=0.835
+ $X2=0 $Y2=0
cc_464 N_A_610_487#_c_537_n N_A_831_47#_c_778_n 0.00779577f $X=5.605 $Y=1.59
+ $X2=0 $Y2=0
cc_465 N_A_610_487#_c_538_n N_A_831_47#_c_779_n 0.00647209f $X=8.185 $Y=0.845
+ $X2=0 $Y2=0
cc_466 N_A_610_487#_c_627_p N_A_1178_399#_M1014_d 0.0157206f $X=7.295 $Y=2.83
+ $X2=0 $Y2=0
cc_467 N_A_610_487#_c_552_n N_A_1178_399#_M1014_d 0.00540356f $X=7.38 $Y=2.745
+ $X2=0 $Y2=0
cc_468 N_A_610_487#_M1011_g N_A_1178_399#_c_935_n 0.00915183f $X=5.605 $Y=2.465
+ $X2=0 $Y2=0
cc_469 N_A_610_487#_c_549_n N_A_1178_399#_c_935_n 0.00249765f $X=5.76 $Y=2.115
+ $X2=0 $Y2=0
cc_470 N_A_610_487#_M1011_g N_A_1178_399#_c_942_n 0.0487188f $X=5.605 $Y=2.465
+ $X2=0 $Y2=0
cc_471 N_A_610_487#_c_549_n N_A_1178_399#_c_942_n 0.002881f $X=5.76 $Y=2.115
+ $X2=0 $Y2=0
cc_472 N_A_610_487#_c_550_n N_A_1178_399#_c_942_n 0.00224534f $X=5.76 $Y=2.835
+ $X2=0 $Y2=0
cc_473 N_A_610_487#_c_551_n N_A_1178_399#_c_942_n 0.0295254f $X=6.545 $Y=2.2
+ $X2=0 $Y2=0
cc_474 N_A_610_487#_c_635_p N_A_1178_399#_c_942_n 0.00309101f $X=6.63 $Y=2.745
+ $X2=0 $Y2=0
cc_475 N_A_610_487#_c_551_n N_A_1178_399#_c_936_n 0.0153796f $X=6.545 $Y=2.2
+ $X2=0 $Y2=0
cc_476 N_A_610_487#_c_532_n N_A_1178_399#_c_937_n 0.0228012f $X=7.55 $Y=1.835
+ $X2=0 $Y2=0
cc_477 N_A_610_487#_c_555_n N_A_1178_399#_c_937_n 0.0012826f $X=7.465 $Y=1.93
+ $X2=0 $Y2=0
cc_478 N_A_610_487#_c_556_n N_A_1178_399#_c_937_n 0.00970533f $X=7.55 $Y=1.95
+ $X2=0 $Y2=0
cc_479 N_A_610_487#_M1019_g N_A_1178_399#_c_945_n 0.00136764f $X=7.515 $Y=2.675
+ $X2=0 $Y2=0
cc_480 N_A_610_487#_c_551_n N_A_1178_399#_c_945_n 0.0125838f $X=6.545 $Y=2.2
+ $X2=0 $Y2=0
cc_481 N_A_610_487#_c_627_p N_A_1178_399#_c_945_n 0.0141188f $X=7.295 $Y=2.83
+ $X2=0 $Y2=0
cc_482 N_A_610_487#_c_552_n N_A_1178_399#_c_945_n 0.0385488f $X=7.38 $Y=2.745
+ $X2=0 $Y2=0
cc_483 N_A_610_487#_c_555_n N_A_1178_399#_c_945_n 5.42286e-19 $X=7.465 $Y=1.93
+ $X2=0 $Y2=0
cc_484 N_A_610_487#_c_556_n N_A_1178_399#_c_945_n 0.00970121f $X=7.55 $Y=1.95
+ $X2=0 $Y2=0
cc_485 N_A_610_487#_c_532_n N_A_1178_399#_c_938_n 0.003536f $X=7.55 $Y=1.835
+ $X2=0 $Y2=0
cc_486 N_A_610_487#_c_585_p N_A_1178_399#_c_938_n 0.0136526f $X=7.635 $Y=1.36
+ $X2=0 $Y2=0
cc_487 N_A_610_487#_c_536_n N_A_1178_399#_c_939_n 0.00219246f $X=5.76 $Y=1.59
+ $X2=0 $Y2=0
cc_488 N_A_610_487#_c_537_n N_A_1178_399#_c_939_n 0.0175132f $X=5.605 $Y=1.59
+ $X2=0 $Y2=0
cc_489 N_A_610_487#_c_549_n N_A_1178_399#_c_940_n 0.0144605f $X=5.76 $Y=2.115
+ $X2=0 $Y2=0
cc_490 N_A_610_487#_c_551_n N_A_1178_399#_c_940_n 0.0398204f $X=6.545 $Y=2.2
+ $X2=0 $Y2=0
cc_491 N_A_610_487#_c_536_n N_A_1178_399#_c_940_n 0.0263218f $X=5.76 $Y=1.59
+ $X2=0 $Y2=0
cc_492 N_A_610_487#_c_537_n N_A_1178_399#_c_940_n 3.18259e-19 $X=5.605 $Y=1.59
+ $X2=0 $Y2=0
cc_493 N_A_610_487#_M1019_g N_A_1047_125#_M1014_g 0.0180702f $X=7.515 $Y=2.675
+ $X2=0 $Y2=0
cc_494 N_A_610_487#_c_551_n N_A_1047_125#_M1014_g 0.00206395f $X=6.545 $Y=2.2
+ $X2=0 $Y2=0
cc_495 N_A_610_487#_c_627_p N_A_1047_125#_M1014_g 0.0171215f $X=7.295 $Y=2.83
+ $X2=0 $Y2=0
cc_496 N_A_610_487#_c_552_n N_A_1047_125#_M1014_g 0.00212636f $X=7.38 $Y=2.745
+ $X2=0 $Y2=0
cc_497 N_A_610_487#_c_532_n N_A_1047_125#_M1014_g 8.89372e-19 $X=7.55 $Y=1.835
+ $X2=0 $Y2=0
cc_498 N_A_610_487#_c_555_n N_A_1047_125#_M1014_g 0.00870381f $X=7.465 $Y=1.93
+ $X2=0 $Y2=0
cc_499 N_A_610_487#_c_556_n N_A_1047_125#_M1014_g 5.23253e-19 $X=7.55 $Y=1.95
+ $X2=0 $Y2=0
cc_500 N_A_610_487#_M1012_g N_A_1047_125#_c_1013_n 0.00546045f $X=5.16 $Y=0.835
+ $X2=0 $Y2=0
cc_501 N_A_610_487#_M1011_g N_A_1047_125#_c_1013_n 0.00359131f $X=5.605 $Y=2.465
+ $X2=0 $Y2=0
cc_502 N_A_610_487#_c_549_n N_A_1047_125#_c_1013_n 0.00734639f $X=5.76 $Y=2.115
+ $X2=0 $Y2=0
cc_503 N_A_610_487#_c_536_n N_A_1047_125#_c_1013_n 0.023711f $X=5.76 $Y=1.59
+ $X2=0 $Y2=0
cc_504 N_A_610_487#_c_537_n N_A_1047_125#_c_1013_n 0.015455f $X=5.605 $Y=1.59
+ $X2=0 $Y2=0
cc_505 N_A_610_487#_M1012_g N_A_1047_125#_c_1014_n 3.9023e-19 $X=5.16 $Y=0.835
+ $X2=0 $Y2=0
cc_506 N_A_610_487#_M1011_g N_A_1047_125#_c_1021_n 0.00118873f $X=5.605 $Y=2.465
+ $X2=0 $Y2=0
cc_507 N_A_610_487#_c_547_n N_A_1047_125#_c_1021_n 0.0116818f $X=5.675 $Y=2.92
+ $X2=0 $Y2=0
cc_508 N_A_610_487#_c_549_n N_A_1047_125#_c_1021_n 6.5885e-19 $X=5.76 $Y=2.115
+ $X2=0 $Y2=0
cc_509 N_A_610_487#_c_670_p N_A_1047_125#_c_1021_n 0.0119668f $X=5.76 $Y=2.2
+ $X2=0 $Y2=0
cc_510 N_A_610_487#_M1012_g N_A_1047_125#_c_1015_n 0.00794792f $X=5.16 $Y=0.835
+ $X2=0 $Y2=0
cc_511 N_A_610_487#_c_536_n N_A_1047_125#_c_1015_n 3.99442e-19 $X=5.76 $Y=1.59
+ $X2=0 $Y2=0
cc_512 N_A_610_487#_c_537_n N_A_1047_125#_c_1015_n 0.0073857f $X=5.605 $Y=1.59
+ $X2=0 $Y2=0
cc_513 N_A_610_487#_M1011_g N_A_1047_125#_c_1022_n 0.00224082f $X=5.605 $Y=2.465
+ $X2=0 $Y2=0
cc_514 N_A_610_487#_c_549_n N_A_1047_125#_c_1022_n 0.0122683f $X=5.76 $Y=2.115
+ $X2=0 $Y2=0
cc_515 N_A_610_487#_c_536_n N_A_1047_125#_c_1022_n 7.19884e-19 $X=5.76 $Y=1.59
+ $X2=0 $Y2=0
cc_516 N_A_610_487#_c_537_n N_A_1047_125#_c_1022_n 0.00696318f $X=5.605 $Y=1.59
+ $X2=0 $Y2=0
cc_517 N_A_610_487#_c_536_n N_A_1047_125#_c_1017_n 0.0259364f $X=5.76 $Y=1.59
+ $X2=0 $Y2=0
cc_518 N_A_610_487#_c_537_n N_A_1047_125#_c_1017_n 0.00351984f $X=5.605 $Y=1.59
+ $X2=0 $Y2=0
cc_519 N_A_610_487#_c_533_n N_A_1665_381#_M1028_g 9.60041e-19 $X=8.02 $Y=1.36
+ $X2=0 $Y2=0
cc_520 N_A_610_487#_c_534_n N_A_1665_381#_M1028_g 9.60468e-19 $X=8.185 $Y=1.01
+ $X2=0 $Y2=0
cc_521 N_A_610_487#_c_538_n N_A_1665_381#_M1028_g 0.0620219f $X=8.185 $Y=0.845
+ $X2=0 $Y2=0
cc_522 N_A_610_487#_c_533_n N_A_1517_63#_c_1224_n 0.00137487f $X=8.02 $Y=1.36
+ $X2=0 $Y2=0
cc_523 N_A_610_487#_c_534_n N_A_1517_63#_c_1224_n 0.0200485f $X=8.185 $Y=1.01
+ $X2=0 $Y2=0
cc_524 N_A_610_487#_c_535_n N_A_1517_63#_c_1224_n 0.00116306f $X=8.185 $Y=1.01
+ $X2=0 $Y2=0
cc_525 N_A_610_487#_c_538_n N_A_1517_63#_c_1224_n 0.0122069f $X=8.185 $Y=0.845
+ $X2=0 $Y2=0
cc_526 N_A_610_487#_c_532_n N_A_1517_63#_c_1212_n 0.0137863f $X=7.55 $Y=1.835
+ $X2=0 $Y2=0
cc_527 N_A_610_487#_c_533_n N_A_1517_63#_c_1212_n 0.0124948f $X=8.02 $Y=1.36
+ $X2=0 $Y2=0
cc_528 N_A_610_487#_c_534_n N_A_1517_63#_c_1213_n 0.0216369f $X=8.185 $Y=1.01
+ $X2=0 $Y2=0
cc_529 N_A_610_487#_c_538_n N_A_1517_63#_c_1213_n 0.00531897f $X=8.185 $Y=0.845
+ $X2=0 $Y2=0
cc_530 N_A_610_487#_M1019_g N_A_1517_63#_c_1220_n 8.37386e-19 $X=7.515 $Y=2.675
+ $X2=0 $Y2=0
cc_531 N_A_610_487#_c_552_n N_A_1517_63#_c_1220_n 0.0180477f $X=7.38 $Y=2.745
+ $X2=0 $Y2=0
cc_532 N_A_610_487#_M1019_g N_A_1517_63#_c_1221_n 0.00106533f $X=7.515 $Y=2.675
+ $X2=0 $Y2=0
cc_533 N_A_610_487#_c_552_n N_A_1517_63#_c_1221_n 0.0070626f $X=7.38 $Y=2.745
+ $X2=0 $Y2=0
cc_534 N_A_610_487#_c_532_n N_A_1517_63#_c_1221_n 0.00213305f $X=7.55 $Y=1.835
+ $X2=0 $Y2=0
cc_535 N_A_610_487#_c_555_n N_A_1517_63#_c_1221_n 0.00112789f $X=7.465 $Y=1.93
+ $X2=0 $Y2=0
cc_536 N_A_610_487#_c_556_n N_A_1517_63#_c_1221_n 0.0174762f $X=7.55 $Y=1.95
+ $X2=0 $Y2=0
cc_537 N_A_610_487#_c_533_n N_A_1517_63#_c_1214_n 0.0244958f $X=8.02 $Y=1.36
+ $X2=0 $Y2=0
cc_538 N_A_610_487#_c_535_n N_A_1517_63#_c_1214_n 0.00177208f $X=8.185 $Y=1.01
+ $X2=0 $Y2=0
cc_539 N_A_610_487#_c_533_n N_A_1517_63#_c_1215_n 0.0159951f $X=8.02 $Y=1.36
+ $X2=0 $Y2=0
cc_540 N_A_610_487#_c_534_n N_A_1517_63#_c_1215_n 0.0120675f $X=8.185 $Y=1.01
+ $X2=0 $Y2=0
cc_541 N_A_610_487#_c_535_n N_A_1517_63#_c_1215_n 2.53979e-19 $X=8.185 $Y=1.01
+ $X2=0 $Y2=0
cc_542 N_A_610_487#_c_544_n N_VPWR_M1006_s 0.004503f $X=3.905 $Y=2.385 $X2=0
+ $Y2=0
cc_543 N_A_610_487#_c_603_p N_VPWR_M1006_s 0.0052183f $X=4.06 $Y=2.835 $X2=0
+ $Y2=0
cc_544 N_A_610_487#_c_548_n N_VPWR_M1006_s 0.00166402f $X=4.145 $Y=2.92 $X2=0
+ $Y2=0
cc_545 N_A_610_487#_c_605_p N_VPWR_M1006_s 0.00130486f $X=4.025 $Y=2.385 $X2=0
+ $Y2=0
cc_546 N_A_610_487#_c_551_n N_VPWR_M1002_d 0.0096746f $X=6.545 $Y=2.2 $X2=0
+ $Y2=0
cc_547 N_A_610_487#_c_635_p N_VPWR_M1002_d 0.00761723f $X=6.63 $Y=2.745 $X2=0
+ $Y2=0
cc_548 N_A_610_487#_c_709_p N_VPWR_M1002_d 0.00379224f $X=6.715 $Y=2.83 $X2=0
+ $Y2=0
cc_549 N_A_610_487#_c_543_n N_VPWR_c_1310_n 0.0159421f $X=3.19 $Y=2.58 $X2=0
+ $Y2=0
cc_550 N_A_610_487#_c_539_n N_VPWR_c_1311_n 0.00499394f $X=4.195 $Y=2.235 $X2=0
+ $Y2=0
cc_551 N_A_610_487#_c_543_n N_VPWR_c_1311_n 0.0280135f $X=3.19 $Y=2.58 $X2=0
+ $Y2=0
cc_552 N_A_610_487#_c_544_n N_VPWR_c_1311_n 0.0176815f $X=3.905 $Y=2.385 $X2=0
+ $Y2=0
cc_553 N_A_610_487#_c_603_p N_VPWR_c_1311_n 0.0145482f $X=4.06 $Y=2.835 $X2=0
+ $Y2=0
cc_554 N_A_610_487#_c_548_n N_VPWR_c_1311_n 0.0142638f $X=4.145 $Y=2.92 $X2=0
+ $Y2=0
cc_555 N_A_610_487#_c_547_n N_VPWR_c_1312_n 0.0113459f $X=5.675 $Y=2.92 $X2=0
+ $Y2=0
cc_556 N_A_610_487#_c_550_n N_VPWR_c_1312_n 0.00946973f $X=5.76 $Y=2.835 $X2=0
+ $Y2=0
cc_557 N_A_610_487#_c_551_n N_VPWR_c_1312_n 0.0225362f $X=6.545 $Y=2.2 $X2=0
+ $Y2=0
cc_558 N_A_610_487#_c_635_p N_VPWR_c_1312_n 0.0218441f $X=6.63 $Y=2.745 $X2=0
+ $Y2=0
cc_559 N_A_610_487#_c_709_p N_VPWR_c_1312_n 0.0143119f $X=6.715 $Y=2.83 $X2=0
+ $Y2=0
cc_560 N_A_610_487#_c_539_n N_VPWR_c_1319_n 0.00302068f $X=4.195 $Y=2.235 $X2=0
+ $Y2=0
cc_561 N_A_610_487#_c_547_n N_VPWR_c_1319_n 0.076577f $X=5.675 $Y=2.92 $X2=0
+ $Y2=0
cc_562 N_A_610_487#_c_548_n N_VPWR_c_1319_n 0.00832985f $X=4.145 $Y=2.92 $X2=0
+ $Y2=0
cc_563 N_A_610_487#_M1019_g N_VPWR_c_1322_n 0.00552635f $X=7.515 $Y=2.675 $X2=0
+ $Y2=0
cc_564 N_A_610_487#_c_627_p N_VPWR_c_1322_n 0.0216368f $X=7.295 $Y=2.83 $X2=0
+ $Y2=0
cc_565 N_A_610_487#_c_709_p N_VPWR_c_1322_n 0.00531125f $X=6.715 $Y=2.83 $X2=0
+ $Y2=0
cc_566 N_A_610_487#_c_539_n N_VPWR_c_1307_n 0.00461941f $X=4.195 $Y=2.235 $X2=0
+ $Y2=0
cc_567 N_A_610_487#_M1019_g N_VPWR_c_1307_n 0.0118552f $X=7.515 $Y=2.675 $X2=0
+ $Y2=0
cc_568 N_A_610_487#_c_543_n N_VPWR_c_1307_n 0.0123071f $X=3.19 $Y=2.58 $X2=0
+ $Y2=0
cc_569 N_A_610_487#_c_544_n N_VPWR_c_1307_n 0.00670306f $X=3.905 $Y=2.385 $X2=0
+ $Y2=0
cc_570 N_A_610_487#_c_547_n N_VPWR_c_1307_n 0.0608018f $X=5.675 $Y=2.92 $X2=0
+ $Y2=0
cc_571 N_A_610_487#_c_548_n N_VPWR_c_1307_n 0.0062468f $X=4.145 $Y=2.92 $X2=0
+ $Y2=0
cc_572 N_A_610_487#_c_627_p N_VPWR_c_1307_n 0.0247346f $X=7.295 $Y=2.83 $X2=0
+ $Y2=0
cc_573 N_A_610_487#_c_709_p N_VPWR_c_1307_n 0.00602664f $X=6.715 $Y=2.83 $X2=0
+ $Y2=0
cc_574 N_A_610_487#_c_605_p N_VPWR_c_1307_n 0.001433f $X=4.025 $Y=2.385 $X2=0
+ $Y2=0
cc_575 N_A_610_487#_c_543_n N_A_328_119#_c_1462_n 0.00541383f $X=3.19 $Y=2.58
+ $X2=0 $Y2=0
cc_576 N_A_610_487#_c_545_n N_A_328_119#_c_1462_n 9.21149e-19 $X=3.355 $Y=2.385
+ $X2=0 $Y2=0
cc_577 N_A_610_487#_c_545_n N_A_328_119#_c_1453_n 0.00387139f $X=3.355 $Y=2.385
+ $X2=0 $Y2=0
cc_578 N_A_610_487#_M1012_g N_A_328_119#_c_1451_n 0.00240486f $X=5.16 $Y=0.835
+ $X2=0 $Y2=0
cc_579 N_A_610_487#_M1012_g N_A_328_119#_c_1452_n 0.00911449f $X=5.16 $Y=0.835
+ $X2=0 $Y2=0
cc_580 N_A_610_487#_M1011_g N_A_328_119#_c_1452_n 3.32245e-19 $X=5.605 $Y=2.465
+ $X2=0 $Y2=0
cc_581 N_A_610_487#_c_539_n N_A_328_119#_c_1458_n 0.00614388f $X=4.195 $Y=2.235
+ $X2=0 $Y2=0
cc_582 N_A_610_487#_c_543_n N_A_328_119#_c_1458_n 0.0164217f $X=3.19 $Y=2.58
+ $X2=0 $Y2=0
cc_583 N_A_610_487#_c_544_n N_A_328_119#_c_1458_n 0.0231958f $X=3.905 $Y=2.385
+ $X2=0 $Y2=0
cc_584 N_A_610_487#_c_545_n N_A_328_119#_c_1458_n 0.0125531f $X=3.355 $Y=2.385
+ $X2=0 $Y2=0
cc_585 N_A_610_487#_c_603_p N_A_328_119#_c_1458_n 0.00837914f $X=4.06 $Y=2.835
+ $X2=0 $Y2=0
cc_586 N_A_610_487#_c_547_n N_A_328_119#_c_1458_n 0.0140339f $X=5.675 $Y=2.92
+ $X2=0 $Y2=0
cc_587 N_A_610_487#_c_605_p N_A_328_119#_c_1458_n 0.0127948f $X=4.025 $Y=2.385
+ $X2=0 $Y2=0
cc_588 N_A_610_487#_c_543_n N_A_328_119#_c_1459_n 0.0012632f $X=3.19 $Y=2.58
+ $X2=0 $Y2=0
cc_589 N_A_610_487#_c_545_n N_A_328_119#_c_1459_n 0.00100834f $X=3.355 $Y=2.385
+ $X2=0 $Y2=0
cc_590 N_A_610_487#_c_545_n N_A_328_119#_c_1460_n 0.00547814f $X=3.355 $Y=2.385
+ $X2=0 $Y2=0
cc_591 N_A_610_487#_c_547_n N_A_328_119#_c_1534_n 0.00337947f $X=5.675 $Y=2.92
+ $X2=0 $Y2=0
cc_592 N_A_610_487#_c_547_n N_A_328_119#_c_1461_n 0.0147308f $X=5.675 $Y=2.92
+ $X2=0 $Y2=0
cc_593 N_A_610_487#_M1032_g N_VGND_c_1598_n 0.00987638f $X=4.08 $Y=0.445 $X2=0
+ $Y2=0
cc_594 N_A_610_487#_c_529_n N_VGND_c_1598_n 0.021701f $X=3.74 $Y=0.865 $X2=0
+ $Y2=0
cc_595 N_A_610_487#_c_538_n N_VGND_c_1600_n 0.00321258f $X=8.185 $Y=0.845 $X2=0
+ $Y2=0
cc_596 N_A_610_487#_c_529_n N_VGND_c_1609_n 0.00742794f $X=3.74 $Y=0.865 $X2=0
+ $Y2=0
cc_597 N_A_610_487#_M1032_g N_VGND_c_1611_n 0.00505556f $X=4.08 $Y=0.445 $X2=0
+ $Y2=0
cc_598 N_A_610_487#_M1032_g N_VGND_c_1617_n 0.00651427f $X=4.08 $Y=0.445 $X2=0
+ $Y2=0
cc_599 N_A_610_487#_c_529_n N_VGND_c_1617_n 0.0184067f $X=3.74 $Y=0.865 $X2=0
+ $Y2=0
cc_600 N_A_610_487#_c_538_n N_VGND_c_1617_n 0.0047895f $X=8.185 $Y=0.845 $X2=0
+ $Y2=0
cc_601 N_A_831_47#_c_772_n N_A_1178_399#_M1015_d 0.00517711f $X=7.465 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_602 N_A_831_47#_c_770_n N_A_1178_399#_M1020_g 0.00116728f $X=5.61 $Y=0.35
+ $X2=0 $Y2=0
cc_603 N_A_831_47#_c_771_n N_A_1178_399#_M1020_g 0.00279273f $X=5.812 $Y=0.725
+ $X2=0 $Y2=0
cc_604 N_A_831_47#_c_843_p N_A_1178_399#_M1020_g 0.0133933f $X=6.715 $Y=0.81
+ $X2=0 $Y2=0
cc_605 N_A_831_47#_c_844_p N_A_1178_399#_M1020_g 0.00397169f $X=6.825 $Y=0.725
+ $X2=0 $Y2=0
cc_606 N_A_831_47#_c_778_n N_A_1178_399#_M1020_g 0.0348186f $X=5.61 $Y=0.515
+ $X2=0 $Y2=0
cc_607 N_A_831_47#_c_764_n N_A_1178_399#_c_937_n 4.81982e-19 $X=7.795 $Y=1.46
+ $X2=0 $Y2=0
cc_608 N_A_831_47#_c_772_n N_A_1178_399#_c_938_n 0.013472f $X=7.465 $Y=0.34
+ $X2=0 $Y2=0
cc_609 N_A_831_47#_c_774_n N_A_1178_399#_c_938_n 0.0373376f $X=7.63 $Y=1.01
+ $X2=0 $Y2=0
cc_610 N_A_831_47#_c_779_n N_A_1178_399#_c_938_n 0.0101122f $X=7.615 $Y=0.845
+ $X2=0 $Y2=0
cc_611 N_A_831_47#_c_764_n N_A_1047_125#_M1014_g 0.00212034f $X=7.795 $Y=1.46
+ $X2=0 $Y2=0
cc_612 N_A_831_47#_c_843_p N_A_1047_125#_c_1012_n 0.00623452f $X=6.715 $Y=0.81
+ $X2=0 $Y2=0
cc_613 N_A_831_47#_c_844_p N_A_1047_125#_c_1012_n 0.00981877f $X=6.825 $Y=0.725
+ $X2=0 $Y2=0
cc_614 N_A_831_47#_c_772_n N_A_1047_125#_c_1012_n 0.0107238f $X=7.465 $Y=0.34
+ $X2=0 $Y2=0
cc_615 N_A_831_47#_c_773_n N_A_1047_125#_c_1012_n 0.00367264f $X=6.935 $Y=0.34
+ $X2=0 $Y2=0
cc_616 N_A_831_47#_c_774_n N_A_1047_125#_c_1012_n 6.6666e-19 $X=7.63 $Y=1.01
+ $X2=0 $Y2=0
cc_617 N_A_831_47#_c_779_n N_A_1047_125#_c_1012_n 0.0139565f $X=7.615 $Y=0.845
+ $X2=0 $Y2=0
cc_618 N_A_831_47#_c_769_n N_A_1047_125#_c_1014_n 0.0151213f $X=5.66 $Y=0.375
+ $X2=0 $Y2=0
cc_619 N_A_831_47#_c_770_n N_A_1047_125#_c_1014_n 0.00104745f $X=5.61 $Y=0.35
+ $X2=0 $Y2=0
cc_620 N_A_831_47#_c_771_n N_A_1047_125#_c_1014_n 0.00407788f $X=5.812 $Y=0.725
+ $X2=0 $Y2=0
cc_621 N_A_831_47#_c_860_p N_A_1047_125#_c_1014_n 0.013606f $X=5.965 $Y=0.81
+ $X2=0 $Y2=0
cc_622 N_A_831_47#_c_778_n N_A_1047_125#_c_1014_n 0.00604613f $X=5.61 $Y=0.515
+ $X2=0 $Y2=0
cc_623 N_A_831_47#_c_781_n N_A_1047_125#_c_1021_n 0.00154706f $X=5.1 $Y=2.07
+ $X2=0 $Y2=0
cc_624 N_A_831_47#_c_769_n N_A_1047_125#_c_1015_n 0.00407835f $X=5.66 $Y=0.375
+ $X2=0 $Y2=0
cc_625 N_A_831_47#_c_781_n N_A_1047_125#_c_1022_n 0.00760366f $X=5.1 $Y=2.07
+ $X2=0 $Y2=0
cc_626 N_A_831_47#_c_843_p N_A_1047_125#_c_1016_n 0.0144679f $X=6.715 $Y=0.81
+ $X2=0 $Y2=0
cc_627 N_A_831_47#_c_769_n N_A_1047_125#_c_1017_n 0.00456842f $X=5.66 $Y=0.375
+ $X2=0 $Y2=0
cc_628 N_A_831_47#_c_770_n N_A_1047_125#_c_1017_n 0.00185377f $X=5.61 $Y=0.35
+ $X2=0 $Y2=0
cc_629 N_A_831_47#_c_843_p N_A_1047_125#_c_1017_n 0.0493424f $X=6.715 $Y=0.81
+ $X2=0 $Y2=0
cc_630 N_A_831_47#_c_860_p N_A_1047_125#_c_1017_n 0.0194485f $X=5.965 $Y=0.81
+ $X2=0 $Y2=0
cc_631 N_A_831_47#_c_778_n N_A_1047_125#_c_1017_n 0.00742143f $X=5.61 $Y=0.515
+ $X2=0 $Y2=0
cc_632 N_A_831_47#_c_762_n N_A_1047_125#_c_1018_n 0.0139565f $X=7.615 $Y=1.385
+ $X2=0 $Y2=0
cc_633 N_A_831_47#_c_843_p N_A_1047_125#_c_1018_n 0.00744872f $X=6.715 $Y=0.81
+ $X2=0 $Y2=0
cc_634 N_A_831_47#_c_763_n N_A_1665_381#_M1028_g 0.0126551f $X=7.965 $Y=1.46
+ $X2=0 $Y2=0
cc_635 N_A_831_47#_M1016_g N_A_1665_381#_c_1119_n 5.95094e-19 $X=8.04 $Y=2.675
+ $X2=0 $Y2=0
cc_636 N_A_831_47#_M1016_g N_A_1665_381#_c_1125_n 0.0651711f $X=8.04 $Y=2.675
+ $X2=0 $Y2=0
cc_637 N_A_831_47#_c_772_n N_A_1517_63#_M1033_d 0.00139981f $X=7.465 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_638 N_A_831_47#_c_774_n N_A_1517_63#_M1033_d 0.00374298f $X=7.63 $Y=1.01
+ $X2=-0.19 $Y2=-0.245
cc_639 N_A_831_47#_c_772_n N_A_1517_63#_c_1224_n 0.00769068f $X=7.465 $Y=0.34
+ $X2=0 $Y2=0
cc_640 N_A_831_47#_c_774_n N_A_1517_63#_c_1224_n 0.0194748f $X=7.63 $Y=1.01
+ $X2=0 $Y2=0
cc_641 N_A_831_47#_c_779_n N_A_1517_63#_c_1224_n 9.981e-19 $X=7.615 $Y=0.845
+ $X2=0 $Y2=0
cc_642 N_A_831_47#_c_763_n N_A_1517_63#_c_1212_n 0.00330333f $X=7.965 $Y=1.46
+ $X2=0 $Y2=0
cc_643 N_A_831_47#_M1016_g N_A_1517_63#_c_1212_n 0.00323005f $X=8.04 $Y=2.675
+ $X2=0 $Y2=0
cc_644 N_A_831_47#_c_764_n N_A_1517_63#_c_1220_n 0.00490871f $X=7.795 $Y=1.46
+ $X2=0 $Y2=0
cc_645 N_A_831_47#_M1016_g N_A_1517_63#_c_1220_n 0.0227219f $X=8.04 $Y=2.675
+ $X2=0 $Y2=0
cc_646 N_A_831_47#_M1016_g N_A_1517_63#_c_1221_n 0.0104484f $X=8.04 $Y=2.675
+ $X2=0 $Y2=0
cc_647 N_A_831_47#_M1016_g N_A_1517_63#_c_1214_n 0.0122767f $X=8.04 $Y=2.675
+ $X2=0 $Y2=0
cc_648 N_A_831_47#_c_762_n N_A_1517_63#_c_1215_n 4.42883e-19 $X=7.615 $Y=1.385
+ $X2=0 $Y2=0
cc_649 N_A_831_47#_c_763_n N_A_1517_63#_c_1215_n 0.00464261f $X=7.965 $Y=1.46
+ $X2=0 $Y2=0
cc_650 N_A_831_47#_M1016_g N_VPWR_c_1313_n 0.00187295f $X=8.04 $Y=2.675 $X2=0
+ $Y2=0
cc_651 N_A_831_47#_M1016_g N_VPWR_c_1322_n 0.00467948f $X=8.04 $Y=2.675 $X2=0
+ $Y2=0
cc_652 N_A_831_47#_M1016_g N_VPWR_c_1307_n 0.00455984f $X=8.04 $Y=2.675 $X2=0
+ $Y2=0
cc_653 N_A_831_47#_c_769_n N_A_328_119#_c_1451_n 0.0235197f $X=5.66 $Y=0.375
+ $X2=0 $Y2=0
cc_654 N_A_831_47#_c_771_n N_A_328_119#_c_1451_n 4.139e-19 $X=5.812 $Y=0.725
+ $X2=0 $Y2=0
cc_655 N_A_831_47#_c_777_n N_A_328_119#_c_1451_n 0.0198763f $X=4.47 $Y=1.175
+ $X2=0 $Y2=0
cc_656 N_A_831_47#_c_781_n N_A_328_119#_c_1452_n 0.0133347f $X=5.1 $Y=2.07 $X2=0
+ $Y2=0
cc_657 N_A_831_47#_c_783_n N_A_328_119#_c_1452_n 0.0024821f $X=5.175 $Y=2.145
+ $X2=0 $Y2=0
cc_658 N_A_831_47#_c_766_n N_A_328_119#_c_1452_n 0.0820953f $X=4.47 $Y=1.33
+ $X2=0 $Y2=0
cc_659 N_A_831_47#_c_768_n N_A_328_119#_c_1452_n 0.0102814f $X=4.53 $Y=1.34
+ $X2=0 $Y2=0
cc_660 N_A_831_47#_c_777_n N_A_328_119#_c_1452_n 0.0125148f $X=4.47 $Y=1.175
+ $X2=0 $Y2=0
cc_661 N_A_831_47#_M1006_d N_A_328_119#_c_1458_n 4.27751e-19 $X=4.27 $Y=2.345
+ $X2=0 $Y2=0
cc_662 N_A_831_47#_c_782_n N_A_328_119#_c_1458_n 0.00404824f $X=4.695 $Y=2.07
+ $X2=0 $Y2=0
cc_663 N_A_831_47#_c_767_n N_A_328_119#_c_1458_n 0.0218537f $X=4.53 $Y=1.34
+ $X2=0 $Y2=0
cc_664 N_A_831_47#_c_783_n N_A_328_119#_c_1534_n 0.00285653f $X=5.175 $Y=2.145
+ $X2=0 $Y2=0
cc_665 N_A_831_47#_c_767_n N_A_328_119#_c_1534_n 5.52072e-19 $X=4.53 $Y=1.34
+ $X2=0 $Y2=0
cc_666 N_A_831_47#_c_781_n N_A_328_119#_c_1461_n 0.00500414f $X=5.1 $Y=2.07
+ $X2=0 $Y2=0
cc_667 N_A_831_47#_c_783_n N_A_328_119#_c_1461_n 0.0036846f $X=5.175 $Y=2.145
+ $X2=0 $Y2=0
cc_668 N_A_831_47#_c_767_n N_A_328_119#_c_1461_n 0.0240264f $X=4.53 $Y=1.34
+ $X2=0 $Y2=0
cc_669 N_A_831_47#_c_843_p N_VGND_M1020_d 0.0172838f $X=6.715 $Y=0.81 $X2=0
+ $Y2=0
cc_670 N_A_831_47#_c_844_p N_VGND_M1020_d 0.00443395f $X=6.825 $Y=0.725 $X2=0
+ $Y2=0
cc_671 N_A_831_47#_c_773_n N_VGND_M1020_d 0.00131161f $X=6.935 $Y=0.34 $X2=0
+ $Y2=0
cc_672 N_A_831_47#_c_769_n N_VGND_c_1599_n 0.015313f $X=5.66 $Y=0.375 $X2=0
+ $Y2=0
cc_673 N_A_831_47#_c_770_n N_VGND_c_1599_n 0.00285653f $X=5.61 $Y=0.35 $X2=0
+ $Y2=0
cc_674 N_A_831_47#_c_771_n N_VGND_c_1599_n 0.00452738f $X=5.812 $Y=0.725 $X2=0
+ $Y2=0
cc_675 N_A_831_47#_c_843_p N_VGND_c_1599_n 0.0265079f $X=6.715 $Y=0.81 $X2=0
+ $Y2=0
cc_676 N_A_831_47#_c_844_p N_VGND_c_1599_n 0.0101063f $X=6.825 $Y=0.725 $X2=0
+ $Y2=0
cc_677 N_A_831_47#_c_773_n N_VGND_c_1599_n 0.0147066f $X=6.935 $Y=0.34 $X2=0
+ $Y2=0
cc_678 N_A_831_47#_c_843_p N_VGND_c_1600_n 0.00244165f $X=6.715 $Y=0.81 $X2=0
+ $Y2=0
cc_679 N_A_831_47#_c_772_n N_VGND_c_1600_n 0.0568729f $X=7.465 $Y=0.34 $X2=0
+ $Y2=0
cc_680 N_A_831_47#_c_773_n N_VGND_c_1600_n 0.0156117f $X=6.935 $Y=0.34 $X2=0
+ $Y2=0
cc_681 N_A_831_47#_c_779_n N_VGND_c_1600_n 0.00308045f $X=7.615 $Y=0.845 $X2=0
+ $Y2=0
cc_682 N_A_831_47#_c_769_n N_VGND_c_1611_n 0.0888305f $X=5.66 $Y=0.375 $X2=0
+ $Y2=0
cc_683 N_A_831_47#_c_770_n N_VGND_c_1611_n 0.0065119f $X=5.61 $Y=0.35 $X2=0
+ $Y2=0
cc_684 N_A_831_47#_c_843_p N_VGND_c_1611_n 0.00278148f $X=6.715 $Y=0.81 $X2=0
+ $Y2=0
cc_685 N_A_831_47#_c_776_n N_VGND_c_1611_n 0.0215408f $X=4.365 $Y=0.375 $X2=0
+ $Y2=0
cc_686 N_A_831_47#_M1032_d N_VGND_c_1617_n 0.00421706f $X=4.155 $Y=0.235 $X2=0
+ $Y2=0
cc_687 N_A_831_47#_c_769_n N_VGND_c_1617_n 0.0525457f $X=5.66 $Y=0.375 $X2=0
+ $Y2=0
cc_688 N_A_831_47#_c_770_n N_VGND_c_1617_n 0.010104f $X=5.61 $Y=0.35 $X2=0 $Y2=0
cc_689 N_A_831_47#_c_843_p N_VGND_c_1617_n 0.0121176f $X=6.715 $Y=0.81 $X2=0
+ $Y2=0
cc_690 N_A_831_47#_c_772_n N_VGND_c_1617_n 0.0314951f $X=7.465 $Y=0.34 $X2=0
+ $Y2=0
cc_691 N_A_831_47#_c_773_n N_VGND_c_1617_n 0.00842509f $X=6.935 $Y=0.34 $X2=0
+ $Y2=0
cc_692 N_A_831_47#_c_776_n N_VGND_c_1617_n 0.0129981f $X=4.365 $Y=0.375 $X2=0
+ $Y2=0
cc_693 N_A_831_47#_c_779_n N_VGND_c_1617_n 0.00492879f $X=7.615 $Y=0.845 $X2=0
+ $Y2=0
cc_694 N_A_831_47#_c_860_p A_1149_125# 0.00142858f $X=5.965 $Y=0.81 $X2=-0.19
+ $Y2=-0.245
cc_695 N_A_1178_399#_c_942_n N_A_1047_125#_M1014_g 0.00573053f $X=6.122 $Y=2.145
+ $X2=0 $Y2=0
cc_696 N_A_1178_399#_c_936_n N_A_1047_125#_M1014_g 0.0219359f $X=6.885 $Y=1.72
+ $X2=0 $Y2=0
cc_697 N_A_1178_399#_c_937_n N_A_1047_125#_M1014_g 0.00779034f $X=7.005 $Y=1.945
+ $X2=0 $Y2=0
cc_698 N_A_1178_399#_c_945_n N_A_1047_125#_M1014_g 0.0112605f $X=7.03 $Y=2.41
+ $X2=0 $Y2=0
cc_699 N_A_1178_399#_c_938_n N_A_1047_125#_M1014_g 0.00221461f $X=7.2 $Y=0.76
+ $X2=0 $Y2=0
cc_700 N_A_1178_399#_c_939_n N_A_1047_125#_M1014_g 0.0231857f $X=6.19 $Y=1.51
+ $X2=0 $Y2=0
cc_701 N_A_1178_399#_c_940_n N_A_1047_125#_M1014_g 4.01167e-19 $X=6.355 $Y=1.685
+ $X2=0 $Y2=0
cc_702 N_A_1178_399#_c_938_n N_A_1047_125#_c_1012_n 0.00756446f $X=7.2 $Y=0.76
+ $X2=0 $Y2=0
cc_703 N_A_1178_399#_M1020_g N_A_1047_125#_c_1013_n 0.00384555f $X=6.06 $Y=0.835
+ $X2=0 $Y2=0
cc_704 N_A_1178_399#_M1020_g N_A_1047_125#_c_1016_n 4.32719e-19 $X=6.06 $Y=0.835
+ $X2=0 $Y2=0
cc_705 N_A_1178_399#_c_936_n N_A_1047_125#_c_1016_n 0.0216213f $X=6.885 $Y=1.72
+ $X2=0 $Y2=0
cc_706 N_A_1178_399#_c_937_n N_A_1047_125#_c_1016_n 0.00411523f $X=7.005
+ $Y=1.945 $X2=0 $Y2=0
cc_707 N_A_1178_399#_c_938_n N_A_1047_125#_c_1016_n 0.0196296f $X=7.2 $Y=0.76
+ $X2=0 $Y2=0
cc_708 N_A_1178_399#_M1020_g N_A_1047_125#_c_1017_n 0.0133249f $X=6.06 $Y=0.835
+ $X2=0 $Y2=0
cc_709 N_A_1178_399#_c_936_n N_A_1047_125#_c_1017_n 0.0154711f $X=6.885 $Y=1.72
+ $X2=0 $Y2=0
cc_710 N_A_1178_399#_c_939_n N_A_1047_125#_c_1017_n 0.00632315f $X=6.19 $Y=1.51
+ $X2=0 $Y2=0
cc_711 N_A_1178_399#_c_940_n N_A_1047_125#_c_1017_n 0.0241908f $X=6.355 $Y=1.685
+ $X2=0 $Y2=0
cc_712 N_A_1178_399#_M1020_g N_A_1047_125#_c_1018_n 0.00638849f $X=6.06 $Y=0.835
+ $X2=0 $Y2=0
cc_713 N_A_1178_399#_c_936_n N_A_1047_125#_c_1018_n 0.00337342f $X=6.885 $Y=1.72
+ $X2=0 $Y2=0
cc_714 N_A_1178_399#_c_937_n N_A_1047_125#_c_1018_n 0.007774f $X=7.005 $Y=1.945
+ $X2=0 $Y2=0
cc_715 N_A_1178_399#_c_939_n N_A_1047_125#_c_1018_n 0.00327734f $X=6.19 $Y=1.51
+ $X2=0 $Y2=0
cc_716 N_A_1178_399#_c_942_n N_VPWR_c_1312_n 0.00511209f $X=6.122 $Y=2.145 $X2=0
+ $Y2=0
cc_717 N_A_1178_399#_c_942_n N_VPWR_c_1319_n 0.00399858f $X=6.122 $Y=2.145 $X2=0
+ $Y2=0
cc_718 N_A_1178_399#_M1014_d N_VPWR_c_1307_n 0.00495263f $X=6.89 $Y=2.255 $X2=0
+ $Y2=0
cc_719 N_A_1178_399#_c_942_n N_VPWR_c_1307_n 0.0046122f $X=6.122 $Y=2.145 $X2=0
+ $Y2=0
cc_720 N_A_1178_399#_M1020_g N_VGND_c_1599_n 0.00138928f $X=6.06 $Y=0.835 $X2=0
+ $Y2=0
cc_721 N_A_1178_399#_M1020_g N_VGND_c_1611_n 0.00326244f $X=6.06 $Y=0.835 $X2=0
+ $Y2=0
cc_722 N_A_1178_399#_M1020_g N_VGND_c_1617_n 0.00469432f $X=6.06 $Y=0.835 $X2=0
+ $Y2=0
cc_723 N_A_1047_125#_M1014_g N_VPWR_c_1312_n 0.00899169f $X=6.815 $Y=2.675 $X2=0
+ $Y2=0
cc_724 N_A_1047_125#_M1014_g N_VPWR_c_1322_n 0.00389067f $X=6.815 $Y=2.675 $X2=0
+ $Y2=0
cc_725 N_A_1047_125#_M1014_g N_VPWR_c_1307_n 0.00750974f $X=6.815 $Y=2.675 $X2=0
+ $Y2=0
cc_726 N_A_1047_125#_c_1013_n N_A_328_119#_c_1452_n 0.0478953f $X=5.23 $Y=1.935
+ $X2=0 $Y2=0
cc_727 N_A_1047_125#_c_1014_n N_A_328_119#_c_1452_n 0.00358238f $X=5.375
+ $Y=0.835 $X2=0 $Y2=0
cc_728 N_A_1047_125#_c_1021_n N_A_328_119#_c_1452_n 0.007289f $X=5.39 $Y=2.465
+ $X2=0 $Y2=0
cc_729 N_A_1047_125#_c_1015_n N_A_328_119#_c_1452_n 0.0130065f $X=5.317 $Y=1.16
+ $X2=0 $Y2=0
cc_730 N_A_1047_125#_c_1022_n N_A_328_119#_c_1452_n 0.0120414f $X=5.4 $Y=2.02
+ $X2=0 $Y2=0
cc_731 N_A_1047_125#_c_1021_n N_A_328_119#_c_1534_n 0.00673357f $X=5.39 $Y=2.465
+ $X2=0 $Y2=0
cc_732 N_A_1047_125#_c_1022_n N_A_328_119#_c_1534_n 0.0015766f $X=5.4 $Y=2.02
+ $X2=0 $Y2=0
cc_733 N_A_1047_125#_c_1012_n N_VGND_c_1599_n 0.00295017f $X=6.985 $Y=1.065
+ $X2=0 $Y2=0
cc_734 N_A_1047_125#_c_1012_n N_VGND_c_1600_n 0.00308152f $X=6.985 $Y=1.065
+ $X2=0 $Y2=0
cc_735 N_A_1047_125#_c_1012_n N_VGND_c_1617_n 0.00523582f $X=6.985 $Y=1.065
+ $X2=0 $Y2=0
cc_736 N_A_1665_381#_M1028_g N_A_1517_63#_M1025_g 0.01678f $X=8.635 $Y=0.525
+ $X2=0 $Y2=0
cc_737 N_A_1665_381#_c_1109_n N_A_1517_63#_M1025_g 0.00500635f $X=9.375 $Y=0.39
+ $X2=0 $Y2=0
cc_738 N_A_1665_381#_c_1110_n N_A_1517_63#_M1025_g 0.00840708f $X=9.465 $Y=1.345
+ $X2=0 $Y2=0
cc_739 N_A_1665_381#_c_1112_n N_A_1517_63#_M1025_g 0.00344879f $X=9.38 $Y=0.895
+ $X2=0 $Y2=0
cc_740 N_A_1665_381#_M1022_g N_A_1517_63#_M1000_g 0.00375273f $X=8.4 $Y=2.675
+ $X2=0 $Y2=0
cc_741 N_A_1665_381#_M1028_g N_A_1517_63#_M1000_g 0.0134922f $X=8.635 $Y=0.525
+ $X2=0 $Y2=0
cc_742 N_A_1665_381#_c_1119_n N_A_1517_63#_M1000_g 0.0157338f $X=9.295 $Y=2.065
+ $X2=0 $Y2=0
cc_743 N_A_1665_381#_c_1120_n N_A_1517_63#_M1000_g 0.0035453f $X=9.39 $Y=2.19
+ $X2=0 $Y2=0
cc_744 N_A_1665_381#_c_1121_n N_A_1517_63#_M1000_g 0.00604242f $X=9.465 $Y=1.975
+ $X2=0 $Y2=0
cc_745 N_A_1665_381#_c_1113_n N_A_1517_63#_c_1210_n 0.00371197f $X=9.465 $Y=1.51
+ $X2=0 $Y2=0
cc_746 N_A_1665_381#_c_1114_n N_A_1517_63#_c_1210_n 0.00545418f $X=10.555
+ $Y=1.51 $X2=0 $Y2=0
cc_747 N_A_1665_381#_c_1119_n N_A_1517_63#_c_1211_n 0.0051456f $X=9.295 $Y=2.065
+ $X2=0 $Y2=0
cc_748 N_A_1665_381#_c_1121_n N_A_1517_63#_c_1211_n 0.00317795f $X=9.465
+ $Y=1.975 $X2=0 $Y2=0
cc_749 N_A_1665_381#_M1028_g N_A_1517_63#_c_1224_n 0.00904053f $X=8.635 $Y=0.525
+ $X2=0 $Y2=0
cc_750 N_A_1665_381#_M1028_g N_A_1517_63#_c_1213_n 0.0112941f $X=8.635 $Y=0.525
+ $X2=0 $Y2=0
cc_751 N_A_1665_381#_c_1112_n N_A_1517_63#_c_1213_n 2.72919e-19 $X=9.38 $Y=0.895
+ $X2=0 $Y2=0
cc_752 N_A_1665_381#_M1022_g N_A_1517_63#_c_1220_n 0.00137274f $X=8.4 $Y=2.675
+ $X2=0 $Y2=0
cc_753 N_A_1665_381#_M1028_g N_A_1517_63#_c_1221_n 4.45537e-19 $X=8.635 $Y=0.525
+ $X2=0 $Y2=0
cc_754 N_A_1665_381#_c_1119_n N_A_1517_63#_c_1221_n 0.00776052f $X=9.295
+ $Y=2.065 $X2=0 $Y2=0
cc_755 N_A_1665_381#_c_1125_n N_A_1517_63#_c_1221_n 0.00194869f $X=8.635 $Y=2.07
+ $X2=0 $Y2=0
cc_756 N_A_1665_381#_c_1119_n N_A_1517_63#_c_1214_n 0.0694087f $X=9.295 $Y=2.065
+ $X2=0 $Y2=0
cc_757 N_A_1665_381#_c_1125_n N_A_1517_63#_c_1214_n 0.00642392f $X=8.635 $Y=2.07
+ $X2=0 $Y2=0
cc_758 N_A_1665_381#_M1028_g N_A_1517_63#_c_1215_n 0.0296575f $X=8.635 $Y=0.525
+ $X2=0 $Y2=0
cc_759 N_A_1665_381#_c_1110_n N_A_1517_63#_c_1215_n 0.0166976f $X=9.465 $Y=1.345
+ $X2=0 $Y2=0
cc_760 N_A_1665_381#_c_1121_n N_A_1517_63#_c_1215_n 0.0102705f $X=9.465 $Y=1.975
+ $X2=0 $Y2=0
cc_761 N_A_1665_381#_c_1113_n N_A_1517_63#_c_1215_n 0.0294661f $X=9.465 $Y=1.51
+ $X2=0 $Y2=0
cc_762 N_A_1665_381#_c_1114_n N_A_1517_63#_c_1215_n 2.14833e-19 $X=10.555
+ $Y=1.51 $X2=0 $Y2=0
cc_763 N_A_1665_381#_M1028_g N_A_1517_63#_c_1216_n 0.0366586f $X=8.635 $Y=0.525
+ $X2=0 $Y2=0
cc_764 N_A_1665_381#_c_1110_n N_A_1517_63#_c_1216_n 0.00510337f $X=9.465
+ $Y=1.345 $X2=0 $Y2=0
cc_765 N_A_1665_381#_c_1112_n N_A_1517_63#_c_1216_n 0.00198188f $X=9.38 $Y=0.895
+ $X2=0 $Y2=0
cc_766 N_A_1665_381#_c_1119_n N_VPWR_M1022_d 0.00260896f $X=9.295 $Y=2.065 $X2=0
+ $Y2=0
cc_767 N_A_1665_381#_M1022_g N_VPWR_c_1313_n 0.0178417f $X=8.4 $Y=2.675 $X2=0
+ $Y2=0
cc_768 N_A_1665_381#_c_1119_n N_VPWR_c_1313_n 0.0501823f $X=9.295 $Y=2.065 $X2=0
+ $Y2=0
cc_769 N_A_1665_381#_c_1120_n N_VPWR_c_1313_n 0.0250385f $X=9.39 $Y=2.19 $X2=0
+ $Y2=0
cc_770 N_A_1665_381#_c_1125_n N_VPWR_c_1313_n 0.00667926f $X=8.635 $Y=2.07 $X2=0
+ $Y2=0
cc_771 N_A_1665_381#_M1013_g N_VPWR_c_1314_n 0.0184853f $X=10.125 $Y=2.465 $X2=0
+ $Y2=0
cc_772 N_A_1665_381#_M1024_g N_VPWR_c_1314_n 7.76434e-19 $X=10.555 $Y=2.465
+ $X2=0 $Y2=0
cc_773 N_A_1665_381#_c_1120_n N_VPWR_c_1314_n 0.0553227f $X=9.39 $Y=2.19 $X2=0
+ $Y2=0
cc_774 N_A_1665_381#_c_1121_n N_VPWR_c_1314_n 0.00927918f $X=9.465 $Y=1.975
+ $X2=0 $Y2=0
cc_775 N_A_1665_381#_c_1111_n N_VPWR_c_1314_n 0.0231351f $X=9.97 $Y=1.51 $X2=0
+ $Y2=0
cc_776 N_A_1665_381#_c_1123_n N_VPWR_c_1314_n 0.0143868f $X=9.422 $Y=2.065 $X2=0
+ $Y2=0
cc_777 N_A_1665_381#_c_1114_n N_VPWR_c_1314_n 0.00553375f $X=10.555 $Y=1.51
+ $X2=0 $Y2=0
cc_778 N_A_1665_381#_M1024_g N_VPWR_c_1316_n 0.00776505f $X=10.555 $Y=2.465
+ $X2=0 $Y2=0
cc_779 N_A_1665_381#_M1022_g N_VPWR_c_1322_n 0.00435433f $X=8.4 $Y=2.675 $X2=0
+ $Y2=0
cc_780 N_A_1665_381#_c_1120_n N_VPWR_c_1323_n 0.00866243f $X=9.39 $Y=2.19 $X2=0
+ $Y2=0
cc_781 N_A_1665_381#_M1013_g N_VPWR_c_1324_n 0.00564095f $X=10.125 $Y=2.465
+ $X2=0 $Y2=0
cc_782 N_A_1665_381#_M1024_g N_VPWR_c_1324_n 0.00585385f $X=10.555 $Y=2.465
+ $X2=0 $Y2=0
cc_783 N_A_1665_381#_M1022_g N_VPWR_c_1307_n 0.0043858f $X=8.4 $Y=2.675 $X2=0
+ $Y2=0
cc_784 N_A_1665_381#_M1013_g N_VPWR_c_1307_n 0.00948291f $X=10.125 $Y=2.465
+ $X2=0 $Y2=0
cc_785 N_A_1665_381#_M1024_g N_VPWR_c_1307_n 0.0114507f $X=10.555 $Y=2.465 $X2=0
+ $Y2=0
cc_786 N_A_1665_381#_c_1120_n N_VPWR_c_1307_n 0.00891007f $X=9.39 $Y=2.19 $X2=0
+ $Y2=0
cc_787 N_A_1665_381#_c_1107_n Q 0.00246421f $X=10.125 $Y=1.345 $X2=0 $Y2=0
cc_788 N_A_1665_381#_M1013_g Q 0.00300131f $X=10.125 $Y=2.465 $X2=0 $Y2=0
cc_789 N_A_1665_381#_c_1108_n Q 0.00344894f $X=10.555 $Y=1.345 $X2=0 $Y2=0
cc_790 N_A_1665_381#_M1024_g Q 0.00459033f $X=10.555 $Y=2.465 $X2=0 $Y2=0
cc_791 N_A_1665_381#_c_1110_n Q 0.00403326f $X=9.465 $Y=1.345 $X2=0 $Y2=0
cc_792 N_A_1665_381#_c_1121_n Q 0.0047731f $X=9.465 $Y=1.975 $X2=0 $Y2=0
cc_793 N_A_1665_381#_c_1111_n Q 0.0255779f $X=9.97 $Y=1.51 $X2=0 $Y2=0
cc_794 N_A_1665_381#_c_1114_n Q 0.0301163f $X=10.555 $Y=1.51 $X2=0 $Y2=0
cc_795 N_A_1665_381#_M1028_g N_VGND_c_1600_n 0.0038354f $X=8.635 $Y=0.525 $X2=0
+ $Y2=0
cc_796 N_A_1665_381#_M1028_g N_VGND_c_1601_n 0.00732354f $X=8.635 $Y=0.525 $X2=0
+ $Y2=0
cc_797 N_A_1665_381#_c_1109_n N_VGND_c_1601_n 0.0240593f $X=9.375 $Y=0.39 $X2=0
+ $Y2=0
cc_798 N_A_1665_381#_c_1107_n N_VGND_c_1602_n 0.0130756f $X=10.125 $Y=1.345
+ $X2=0 $Y2=0
cc_799 N_A_1665_381#_c_1108_n N_VGND_c_1602_n 5.32672e-19 $X=10.555 $Y=1.345
+ $X2=0 $Y2=0
cc_800 N_A_1665_381#_c_1109_n N_VGND_c_1602_n 0.0682632f $X=9.375 $Y=0.39 $X2=0
+ $Y2=0
cc_801 N_A_1665_381#_c_1111_n N_VGND_c_1602_n 0.0231351f $X=9.97 $Y=1.51 $X2=0
+ $Y2=0
cc_802 N_A_1665_381#_c_1114_n N_VGND_c_1602_n 0.00553375f $X=10.555 $Y=1.51
+ $X2=0 $Y2=0
cc_803 N_A_1665_381#_c_1108_n N_VGND_c_1604_n 0.00750453f $X=10.555 $Y=1.345
+ $X2=0 $Y2=0
cc_804 N_A_1665_381#_c_1109_n N_VGND_c_1612_n 0.0217292f $X=9.375 $Y=0.39 $X2=0
+ $Y2=0
cc_805 N_A_1665_381#_c_1107_n N_VGND_c_1613_n 0.00539704f $X=10.125 $Y=1.345
+ $X2=0 $Y2=0
cc_806 N_A_1665_381#_c_1108_n N_VGND_c_1613_n 0.00559701f $X=10.555 $Y=1.345
+ $X2=0 $Y2=0
cc_807 N_A_1665_381#_M1025_d N_VGND_c_1617_n 0.00215158f $X=9.235 $Y=0.235 $X2=0
+ $Y2=0
cc_808 N_A_1665_381#_M1028_g N_VGND_c_1617_n 0.00644442f $X=8.635 $Y=0.525 $X2=0
+ $Y2=0
cc_809 N_A_1665_381#_c_1107_n N_VGND_c_1617_n 0.0052351f $X=10.125 $Y=1.345
+ $X2=0 $Y2=0
cc_810 N_A_1665_381#_c_1108_n N_VGND_c_1617_n 0.00537853f $X=10.555 $Y=1.345
+ $X2=0 $Y2=0
cc_811 N_A_1665_381#_c_1109_n N_VGND_c_1617_n 0.0129473f $X=9.375 $Y=0.39 $X2=0
+ $Y2=0
cc_812 N_A_1517_63#_M1000_g N_VPWR_c_1313_n 0.0119292f $X=9.175 $Y=2.465 $X2=0
+ $Y2=0
cc_813 N_A_1517_63#_c_1220_n N_VPWR_c_1313_n 0.0269263f $X=7.73 $Y=2.4 $X2=0
+ $Y2=0
cc_814 N_A_1517_63#_M1000_g N_VPWR_c_1314_n 0.00364217f $X=9.175 $Y=2.465 $X2=0
+ $Y2=0
cc_815 N_A_1517_63#_c_1220_n N_VPWR_c_1322_n 0.0242629f $X=7.73 $Y=2.4 $X2=0
+ $Y2=0
cc_816 N_A_1517_63#_M1000_g N_VPWR_c_1323_n 0.00435433f $X=9.175 $Y=2.465 $X2=0
+ $Y2=0
cc_817 N_A_1517_63#_M1019_d N_VPWR_c_1307_n 0.00371702f $X=7.59 $Y=2.255 $X2=0
+ $Y2=0
cc_818 N_A_1517_63#_M1000_g N_VPWR_c_1307_n 0.0043858f $X=9.175 $Y=2.465 $X2=0
+ $Y2=0
cc_819 N_A_1517_63#_c_1220_n N_VPWR_c_1307_n 0.0135294f $X=7.73 $Y=2.4 $X2=0
+ $Y2=0
cc_820 N_A_1517_63#_c_1224_n N_VGND_c_1600_n 0.0264561f $X=8.49 $Y=0.5 $X2=0
+ $Y2=0
cc_821 N_A_1517_63#_M1025_g N_VGND_c_1601_n 0.00401127f $X=9.16 $Y=0.555 $X2=0
+ $Y2=0
cc_822 N_A_1517_63#_c_1224_n N_VGND_c_1601_n 0.0263403f $X=8.49 $Y=0.5 $X2=0
+ $Y2=0
cc_823 N_A_1517_63#_c_1213_n N_VGND_c_1601_n 0.015682f $X=8.575 $Y=1.135 $X2=0
+ $Y2=0
cc_824 N_A_1517_63#_c_1215_n N_VGND_c_1601_n 0.0143746f $X=9.115 $Y=1.3 $X2=0
+ $Y2=0
cc_825 N_A_1517_63#_c_1216_n N_VGND_c_1601_n 0.00227468f $X=9.115 $Y=1.3 $X2=0
+ $Y2=0
cc_826 N_A_1517_63#_M1025_g N_VGND_c_1602_n 0.00325638f $X=9.16 $Y=0.555 $X2=0
+ $Y2=0
cc_827 N_A_1517_63#_M1025_g N_VGND_c_1612_n 0.0054895f $X=9.16 $Y=0.555 $X2=0
+ $Y2=0
cc_828 N_A_1517_63#_M1025_g N_VGND_c_1617_n 0.0119564f $X=9.16 $Y=0.555 $X2=0
+ $Y2=0
cc_829 N_A_1517_63#_c_1224_n N_VGND_c_1617_n 0.0238703f $X=8.49 $Y=0.5 $X2=0
+ $Y2=0
cc_830 N_A_1517_63#_c_1224_n A_1670_63# 0.00446575f $X=8.49 $Y=0.5 $X2=-0.19
+ $Y2=-0.245
cc_831 N_A_1517_63#_c_1213_n A_1670_63# 7.85546e-19 $X=8.575 $Y=1.135 $X2=-0.19
+ $Y2=-0.245
cc_832 N_VPWR_M1001_d N_A_328_119#_c_1462_n 0.00157134f $X=2.54 $Y=2.435 $X2=0
+ $Y2=0
cc_833 N_VPWR_c_1309_n N_A_328_119#_c_1462_n 0.00712673f $X=2.74 $Y=2.855 $X2=0
+ $Y2=0
cc_834 N_VPWR_c_1321_n N_A_328_119#_c_1462_n 0.00718384f $X=2.625 $Y=3.33 $X2=0
+ $Y2=0
cc_835 N_VPWR_c_1307_n N_A_328_119#_c_1462_n 0.0178551f $X=10.8 $Y=3.33 $X2=0
+ $Y2=0
cc_836 N_VPWR_c_1309_n N_A_328_119#_c_1453_n 0.00163704f $X=2.74 $Y=2.855 $X2=0
+ $Y2=0
cc_837 N_VPWR_c_1321_n N_A_328_119#_c_1457_n 0.0188411f $X=2.625 $Y=3.33 $X2=0
+ $Y2=0
cc_838 N_VPWR_c_1307_n N_A_328_119#_c_1457_n 0.0124871f $X=10.8 $Y=3.33 $X2=0
+ $Y2=0
cc_839 N_VPWR_M1001_d N_A_328_119#_c_1458_n 0.00261095f $X=2.54 $Y=2.435 $X2=0
+ $Y2=0
cc_840 N_VPWR_M1006_s N_A_328_119#_c_1458_n 0.00826046f $X=3.585 $Y=2.345 $X2=0
+ $Y2=0
cc_841 N_VPWR_c_1309_n N_A_328_119#_c_1458_n 0.00182684f $X=2.74 $Y=2.855 $X2=0
+ $Y2=0
cc_842 N_VPWR_c_1311_n N_A_328_119#_c_1458_n 0.00652244f $X=3.72 $Y=2.805 $X2=0
+ $Y2=0
cc_843 N_VPWR_M1001_d N_A_328_119#_c_1459_n 0.00288316f $X=2.54 $Y=2.435 $X2=0
+ $Y2=0
cc_844 N_VPWR_c_1309_n N_A_328_119#_c_1459_n 0.00298356f $X=2.74 $Y=2.855 $X2=0
+ $Y2=0
cc_845 N_VPWR_c_1307_n N_Q_M1013_d 0.00362709f $X=10.8 $Y=3.33 $X2=0 $Y2=0
cc_846 N_VPWR_c_1316_n Q 0.00153242f $X=10.77 $Y=1.98 $X2=0 $Y2=0
cc_847 N_VPWR_c_1324_n Q 0.0142265f $X=10.635 $Y=3.33 $X2=0 $Y2=0
cc_848 N_VPWR_c_1307_n Q 0.00925289f $X=10.8 $Y=3.33 $X2=0 $Y2=0
cc_849 N_VPWR_c_1316_n N_VGND_c_1604_n 0.0121422f $X=10.77 $Y=1.98 $X2=0 $Y2=0
cc_850 N_A_328_119#_c_1462_n A_414_487# 0.00680966f $X=2.285 $Y=2.545 $X2=-0.19
+ $Y2=-0.245
cc_851 N_A_328_119#_c_1448_n N_VGND_c_1597_n 0.0249463f $X=2.905 $Y=1.2 $X2=0
+ $Y2=0
cc_852 N_A_328_119#_c_1447_n N_VGND_c_1607_n 0.00360499f $X=2.02 $Y=0.805 $X2=0
+ $Y2=0
cc_853 N_A_328_119#_c_1447_n N_VGND_c_1617_n 0.00521714f $X=2.02 $Y=0.805 $X2=0
+ $Y2=0
cc_854 Q N_VGND_c_1602_n 0.0304851f $X=10.235 $Y=0.47 $X2=0 $Y2=0
cc_855 Q N_VGND_c_1604_n 0.00306484f $X=10.235 $Y=0.47 $X2=0 $Y2=0
cc_856 Q N_VGND_c_1613_n 0.00964975f $X=10.235 $Y=0.47 $X2=0 $Y2=0
cc_857 Q N_VGND_c_1617_n 0.00865647f $X=10.235 $Y=0.47 $X2=0 $Y2=0
