* File: sky130_fd_sc_lp__o22ai_1.spice
* Created: Wed Sep  2 10:20:35 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__o22ai_1.pex.spice"
.subckt sky130_fd_sc_lp__o22ai_1  VNB VPB B1 B2 A2 A1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A1	A1
* A2	A2
* B2	B2
* B1	B1
* VPB	VPB
* VNB	VNB
MM1003 N_Y_M1003_d N_B1_M1003_g N_A_27_69#_M1003_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75001.9 A=0.126 P=1.98 MULT=1
MM1005 N_A_27_69#_M1005_d N_B2_M1005_g N_Y_M1003_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1449 AS=0.1176 PD=1.185 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75001.5 A=0.126 P=1.98 MULT=1
MM1001 N_VGND_M1001_d N_A2_M1001_g N_A_27_69#_M1005_d VNB NSHORT L=0.15 W=0.84
+ AD=0.2604 AS=0.1449 PD=1.46 PS=1.185 NRD=0 NRS=9.276 M=1 R=5.6 SA=75001.1
+ SB=75001 A=0.126 P=1.98 MULT=1
MM1006 N_A_27_69#_M1006_d N_A1_M1006_g N_VGND_M1001_d VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.2604 PD=2.21 PS=1.46 NRD=0 NRS=0 M=1 R=5.6 SA=75001.9
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1007 A_110_367# N_B1_M1007_g N_VPWR_M1007_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1323 AS=0.3339 PD=1.47 PS=3.05 NRD=7.8012 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75001.7 A=0.189 P=2.82 MULT=1
MM1004 N_Y_M1004_d N_B2_M1004_g A_110_367# VPB PHIGHVT L=0.15 W=1.26 AD=0.40635
+ AS=0.1323 PD=1.905 PS=1.47 NRD=0 NRS=7.8012 M=1 R=8.4 SA=75000.6 SB=75001.3
+ A=0.189 P=2.82 MULT=1
MM1002 A_341_367# N_A2_M1002_g N_Y_M1004_d VPB PHIGHVT L=0.15 W=1.26 AD=0.1323
+ AS=0.40635 PD=1.47 PS=1.905 NRD=7.8012 NRS=0 M=1 R=8.4 SA=75001.3 SB=75000.6
+ A=0.189 P=2.82 MULT=1
MM1000 N_VPWR_M1000_d N_A1_M1000_g A_341_367# VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.1323 PD=3.05 PS=1.47 NRD=0 NRS=7.8012 M=1 R=8.4 SA=75001.7
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX8_noxref VNB VPB NWDIODE A=6.0799 P=10.25
*
.include "sky130_fd_sc_lp__o22ai_1.pxi.spice"
*
.ends
*
*
