* File: sky130_fd_sc_lp__mux2_lp.spice
* Created: Wed Sep  2 10:00:40 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__mux2_lp.pex.spice"
.subckt sky130_fd_sc_lp__mux2_lp  VNB VPB A1 A0 S X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* S	S
* A0	A0
* A1	A1
* VPB	VPB
* VNB	VNB
MM1009 A_114_55# N_A_84_29#_M1009_g N_X_M1009_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1197 PD=0.63 PS=1.41 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75003.5 A=0.063 P=1.14 MULT=1
MM1002 N_VGND_M1002_d N_A_84_29#_M1002_g A_114_55# VNB NSHORT L=0.15 W=0.42
+ AD=0.09555 AS=0.0441 PD=0.875 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6
+ SB=75003.2 A=0.063 P=1.14 MULT=1
MM1005 A_307_55# N_A_200_367#_M1005_g N_VGND_M1002_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.09555 PD=0.66 PS=0.875 NRD=18.564 NRS=49.992 M=1 R=2.8
+ SA=75001.2 SB=75002.6 A=0.063 P=1.14 MULT=1
MM1006 N_A_84_29#_M1006_d N_A0_M1006_g A_307_55# VNB NSHORT L=0.15 W=0.42
+ AD=0.10605 AS=0.0504 PD=0.925 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75001.6
+ SB=75002.2 A=0.063 P=1.14 MULT=1
MM1003 A_516_55# N_A1_M1003_g N_A_84_29#_M1006_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0756 AS=0.10605 PD=0.78 PS=0.925 NRD=35.712 NRS=64.284 M=1 R=2.8
+ SA=75002.2 SB=75001.5 A=0.063 P=1.14 MULT=1
MM1008 N_VGND_M1008_d N_S_M1008_g A_516_55# VNB NSHORT L=0.15 W=0.42 AD=0.0588
+ AS=0.0756 PD=0.7 PS=0.78 NRD=0 NRS=35.712 M=1 R=2.8 SA=75002.7 SB=75001
+ A=0.063 P=1.14 MULT=1
MM1013 A_704_55# N_S_M1013_g N_VGND_M1008_d VNB NSHORT L=0.15 W=0.42 AD=0.0441
+ AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75003.2 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1014 N_A_200_367#_M1014_d N_S_M1014_g A_704_55# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75003.5
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1000 A_123_527# N_A_84_29#_M1000_g N_X_M1000_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0441 AS=0.1197 PD=0.63 PS=1.41 NRD=23.443 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75003.5 A=0.063 P=1.14 MULT=1
MM1015 N_VPWR_M1015_d N_A_84_29#_M1015_g A_123_527# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=23.443 M=1 R=2.8 SA=75000.6
+ SB=75003.1 A=0.063 P=1.14 MULT=1
MM1010 A_281_527# N_A_200_367#_M1010_g N_VPWR_M1015_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0504 AS=0.0588 PD=0.66 PS=0.7 NRD=30.4759 NRS=0 M=1 R=2.8 SA=75001
+ SB=75002.7 A=0.063 P=1.14 MULT=1
MM1001 N_A_84_29#_M1001_d N_A1_M1001_g A_281_527# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0588 AS=0.0504 PD=0.7 PS=0.66 NRD=0 NRS=30.4759 M=1 R=2.8 SA=75001.4
+ SB=75002.3 A=0.063 P=1.14 MULT=1
MM1011 A_445_527# N_A0_M1011_g N_A_84_29#_M1001_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0504 AS=0.0588 PD=0.66 PS=0.7 NRD=30.4759 NRS=0 M=1 R=2.8 SA=75001.8
+ SB=75001.9 A=0.063 P=1.14 MULT=1
MM1012 N_VPWR_M1012_d N_S_M1012_g A_445_527# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.15645 AS=0.0504 PD=1.165 PS=0.66 NRD=0 NRS=30.4759 M=1 R=2.8 SA=75002.2
+ SB=75001.5 A=0.063 P=1.14 MULT=1
MM1004 A_702_527# N_S_M1004_g N_VPWR_M1012_d VPB PHIGHVT L=0.15 W=0.42 AD=0.0441
+ AS=0.15645 PD=0.63 PS=1.165 NRD=23.443 NRS=218.099 M=1 R=2.8 SA=75003.1
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1007 N_A_200_367#_M1007_d N_S_M1007_g A_702_527# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=23.443 M=1 R=2.8 SA=75003.5
+ SB=75000.2 A=0.063 P=1.14 MULT=1
DX16_noxref VNB VPB NWDIODE A=8.7655 P=13.13
*
.include "sky130_fd_sc_lp__mux2_lp.pxi.spice"
*
.ends
*
*
