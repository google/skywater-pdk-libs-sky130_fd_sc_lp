* File: sky130_fd_sc_lp__sdlclkp_1.pxi.spice
* Created: Wed Sep  2 10:37:03 2020
* 
x_PM_SKY130_FD_SC_LP__SDLCLKP_1%SCE N_SCE_M1020_g N_SCE_M1011_g N_SCE_c_161_n
+ N_SCE_c_162_n N_SCE_c_163_n SCE SCE SCE SCE SCE N_SCE_c_165_n
+ PM_SKY130_FD_SC_LP__SDLCLKP_1%SCE
x_PM_SKY130_FD_SC_LP__SDLCLKP_1%GATE N_GATE_M1015_g N_GATE_M1018_g
+ N_GATE_c_198_n N_GATE_c_199_n GATE GATE GATE N_GATE_c_201_n
+ PM_SKY130_FD_SC_LP__SDLCLKP_1%GATE
x_PM_SKY130_FD_SC_LP__SDLCLKP_1%A_334_69# N_A_334_69#_M1016_d
+ N_A_334_69#_M1004_d N_A_334_69#_c_249_n N_A_334_69#_c_259_n
+ N_A_334_69#_M1001_g N_A_334_69#_c_250_n N_A_334_69#_M1006_g
+ N_A_334_69#_c_252_n N_A_334_69#_c_253_n N_A_334_69#_c_254_n
+ N_A_334_69#_c_262_n N_A_334_69#_c_255_n N_A_334_69#_c_256_n
+ N_A_334_69#_c_257_n PM_SKY130_FD_SC_LP__SDLCLKP_1%A_334_69#
x_PM_SKY130_FD_SC_LP__SDLCLKP_1%A_254_357# N_A_254_357#_M1003_s
+ N_A_254_357#_M1007_s N_A_254_357#_c_345_n N_A_254_357#_c_346_n
+ N_A_254_357#_c_347_n N_A_254_357#_c_348_n N_A_254_357#_c_349_n
+ N_A_254_357#_M1016_g N_A_254_357#_c_331_n N_A_254_357#_c_332_n
+ N_A_254_357#_c_333_n N_A_254_357#_c_351_n N_A_254_357#_M1004_g
+ N_A_254_357#_c_334_n N_A_254_357#_c_335_n N_A_254_357#_M1019_g
+ N_A_254_357#_M1017_g N_A_254_357#_c_336_n N_A_254_357#_c_353_n
+ N_A_254_357#_c_337_n N_A_254_357#_c_338_n N_A_254_357#_c_339_n
+ N_A_254_357#_c_340_n N_A_254_357#_c_341_n N_A_254_357#_c_342_n
+ N_A_254_357#_c_343_n N_A_254_357#_c_354_n N_A_254_357#_c_344_n
+ PM_SKY130_FD_SC_LP__SDLCLKP_1%A_254_357#
x_PM_SKY130_FD_SC_LP__SDLCLKP_1%A_737_329# N_A_737_329#_M1021_d
+ N_A_737_329#_M1014_d N_A_737_329#_M1000_g N_A_737_329#_M1009_g
+ N_A_737_329#_c_482_n N_A_737_329#_M1013_g N_A_737_329#_M1008_g
+ N_A_737_329#_c_483_n N_A_737_329#_c_495_n N_A_737_329#_c_496_n
+ N_A_737_329#_c_497_n N_A_737_329#_c_484_n N_A_737_329#_c_499_n
+ N_A_737_329#_c_500_n N_A_737_329#_c_485_n N_A_737_329#_c_486_n
+ N_A_737_329#_c_487_n N_A_737_329#_c_488_n N_A_737_329#_c_489_n
+ N_A_737_329#_c_505_n N_A_737_329#_c_506_n N_A_737_329#_c_490_n
+ N_A_737_329#_c_491_n N_A_737_329#_c_492_n
+ PM_SKY130_FD_SC_LP__SDLCLKP_1%A_737_329#
x_PM_SKY130_FD_SC_LP__SDLCLKP_1%A_623_133# N_A_623_133#_M1019_d
+ N_A_623_133#_M1001_d N_A_623_133#_M1021_g N_A_623_133#_M1014_g
+ N_A_623_133#_c_616_n N_A_623_133#_c_617_n N_A_623_133#_c_618_n
+ N_A_623_133#_c_619_n N_A_623_133#_c_620_n N_A_623_133#_c_621_n
+ PM_SKY130_FD_SC_LP__SDLCLKP_1%A_623_133#
x_PM_SKY130_FD_SC_LP__SDLCLKP_1%CLK N_CLK_c_682_n N_CLK_M1003_g N_CLK_M1007_g
+ N_CLK_c_684_n N_CLK_M1012_g N_CLK_M1002_g CLK CLK N_CLK_c_687_n
+ PM_SKY130_FD_SC_LP__SDLCLKP_1%CLK
x_PM_SKY130_FD_SC_LP__SDLCLKP_1%A_1231_367# N_A_1231_367#_M1013_d
+ N_A_1231_367#_M1002_d N_A_1231_367#_M1010_g N_A_1231_367#_c_738_n
+ N_A_1231_367#_M1005_g N_A_1231_367#_c_739_n N_A_1231_367#_c_752_n
+ N_A_1231_367#_c_740_n N_A_1231_367#_c_758_n N_A_1231_367#_c_741_n
+ N_A_1231_367#_c_742_n PM_SKY130_FD_SC_LP__SDLCLKP_1%A_1231_367#
x_PM_SKY130_FD_SC_LP__SDLCLKP_1%VPWR N_VPWR_M1020_s N_VPWR_M1004_s
+ N_VPWR_M1009_d N_VPWR_M1007_d N_VPWR_M1008_d N_VPWR_c_795_n N_VPWR_c_796_n
+ N_VPWR_c_797_n N_VPWR_c_798_n N_VPWR_c_799_n N_VPWR_c_800_n N_VPWR_c_801_n
+ N_VPWR_c_802_n N_VPWR_c_803_n N_VPWR_c_804_n N_VPWR_c_805_n N_VPWR_c_806_n
+ VPWR N_VPWR_c_807_n N_VPWR_c_808_n N_VPWR_c_794_n N_VPWR_c_810_n
+ PM_SKY130_FD_SC_LP__SDLCLKP_1%VPWR
x_PM_SKY130_FD_SC_LP__SDLCLKP_1%A_154_69# N_A_154_69#_M1011_d
+ N_A_154_69#_M1019_s N_A_154_69#_M1015_d N_A_154_69#_M1001_s
+ N_A_154_69#_c_879_n N_A_154_69#_c_884_n N_A_154_69#_c_885_n
+ N_A_154_69#_c_886_n N_A_154_69#_c_887_n N_A_154_69#_c_888_n
+ N_A_154_69#_c_880_n N_A_154_69#_c_889_n N_A_154_69#_c_897_n
+ N_A_154_69#_c_890_n N_A_154_69#_c_881_n N_A_154_69#_c_882_n
+ PM_SKY130_FD_SC_LP__SDLCLKP_1%A_154_69#
x_PM_SKY130_FD_SC_LP__SDLCLKP_1%GCLK N_GCLK_M1005_d N_GCLK_M1010_d GCLK GCLK
+ GCLK GCLK GCLK GCLK GCLK N_GCLK_c_978_n GCLK
+ PM_SKY130_FD_SC_LP__SDLCLKP_1%GCLK
x_PM_SKY130_FD_SC_LP__SDLCLKP_1%VGND N_VGND_M1011_s N_VGND_M1018_d
+ N_VGND_M1000_d N_VGND_M1003_d N_VGND_M1005_s N_VGND_c_992_n N_VGND_c_993_n
+ N_VGND_c_994_n N_VGND_c_995_n N_VGND_c_996_n N_VGND_c_997_n N_VGND_c_998_n
+ N_VGND_c_999_n N_VGND_c_1000_n N_VGND_c_1001_n VGND N_VGND_c_1002_n
+ N_VGND_c_1003_n N_VGND_c_1004_n N_VGND_c_1005_n N_VGND_c_1006_n
+ N_VGND_c_1007_n PM_SKY130_FD_SC_LP__SDLCLKP_1%VGND
cc_1 VNB N_SCE_M1020_g 0.00662351f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.66
cc_2 VNB N_SCE_c_161_n 0.0201091f $X=-0.19 $Y=-0.245 $X2=0.437 $Y2=0.875
cc_3 VNB N_SCE_c_162_n 0.0415552f $X=-0.19 $Y=-0.245 $X2=0.437 $Y2=1.025
cc_4 VNB N_SCE_c_163_n 0.0295179f $X=-0.19 $Y=-0.245 $X2=0.327 $Y2=1.545
cc_5 VNB SCE 0.0368679f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_6 VNB N_SCE_c_165_n 0.0296875f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.04
cc_7 VNB N_GATE_M1015_g 0.00525076f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.66
cc_8 VNB N_GATE_c_198_n 0.058406f $X=-0.19 $Y=-0.245 $X2=0.327 $Y2=1.323
cc_9 VNB N_GATE_c_199_n 0.0178277f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_10 VNB GATE 0.00927397f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_11 VNB N_GATE_c_201_n 0.0152987f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_334_69#_c_249_n 0.0181763f $X=-0.19 $Y=-0.245 $X2=0.695 $Y2=0.555
cc_13 VNB N_A_334_69#_c_250_n 0.0104758f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.95
cc_14 VNB N_A_334_69#_M1006_g 0.0191606f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_334_69#_c_252_n 0.0161373f $X=-0.19 $Y=-0.245 $X2=0.327 $Y2=1.04
cc_16 VNB N_A_334_69#_c_253_n 0.0139628f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_334_69#_c_254_n 0.00182058f $X=-0.19 $Y=-0.245 $X2=0.275 $Y2=1.295
cc_18 VNB N_A_334_69#_c_255_n 7.63129e-19 $X=-0.19 $Y=-0.245 $X2=0.275 $Y2=2.405
cc_19 VNB N_A_334_69#_c_256_n 9.58179e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_334_69#_c_257_n 0.0108823f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_254_357#_M1016_g 0.036311f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_22 VNB N_A_254_357#_c_331_n 0.016415f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=2.32
cc_23 VNB N_A_254_357#_c_332_n 0.00831967f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_254_357#_c_333_n 0.0191456f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_254_357#_c_334_n 0.0354508f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.04
cc_26 VNB N_A_254_357#_c_335_n 0.0190456f $X=-0.19 $Y=-0.245 $X2=0.275 $Y2=0.925
cc_27 VNB N_A_254_357#_c_336_n 0.0126275f $X=-0.19 $Y=-0.245 $X2=0.275 $Y2=2.035
cc_28 VNB N_A_254_357#_c_337_n 0.00521871f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_254_357#_c_338_n 0.0576782f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_254_357#_c_339_n 0.027738f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_254_357#_c_340_n 0.00483992f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_254_357#_c_341_n 0.0127813f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_254_357#_c_342_n 0.00522365f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_254_357#_c_343_n 0.00551685f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_254_357#_c_344_n 0.0240147f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_737_329#_M1000_g 0.0390251f $X=-0.19 $Y=-0.245 $X2=0.437 $Y2=0.875
cc_37 VNB N_A_737_329#_c_482_n 0.0188007f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_38 VNB N_A_737_329#_c_483_n 0.0221803f $X=-0.19 $Y=-0.245 $X2=0.275 $Y2=0.925
cc_39 VNB N_A_737_329#_c_484_n 0.0117102f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_737_329#_c_485_n 0.00442471f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_737_329#_c_486_n 0.00297749f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_737_329#_c_487_n 0.00119649f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_737_329#_c_488_n 0.00496835f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_737_329#_c_489_n 0.00636607f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_737_329#_c_490_n 0.00109958f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_737_329#_c_491_n 0.0256418f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_737_329#_c_492_n 0.0237193f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_623_133#_M1014_g 0.00633319f $X=-0.19 $Y=-0.245 $X2=0.327
+ $Y2=1.545
cc_49 VNB N_A_623_133#_c_616_n 0.00109786f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.95
cc_50 VNB N_A_623_133#_c_617_n 0.00296423f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_623_133#_c_618_n 0.0190482f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.04
cc_52 VNB N_A_623_133#_c_619_n 0.0353744f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.04
cc_53 VNB N_A_623_133#_c_620_n 0.00328946f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_623_133#_c_621_n 0.0229238f $X=-0.19 $Y=-0.245 $X2=0.275 $Y2=1.04
cc_55 VNB N_CLK_c_682_n 0.0195149f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.545
cc_56 VNB N_CLK_M1007_g 0.0116889f $X=-0.19 $Y=-0.245 $X2=0.695 $Y2=0.555
cc_57 VNB N_CLK_c_684_n 0.0158776f $X=-0.19 $Y=-0.245 $X2=0.327 $Y2=1.025
cc_58 VNB N_CLK_M1002_g 0.00976873f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_59 VNB CLK 0.00790795f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_60 VNB N_CLK_c_687_n 0.0857659f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.04
cc_61 VNB N_A_1231_367#_M1010_g 0.00710968f $X=-0.19 $Y=-0.245 $X2=0.437
+ $Y2=0.875
cc_62 VNB N_A_1231_367#_c_738_n 0.0222054f $X=-0.19 $Y=-0.245 $X2=0.327
+ $Y2=1.323
cc_63 VNB N_A_1231_367#_c_739_n 0.00788311f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_A_1231_367#_c_740_n 8.1447e-19 $X=-0.19 $Y=-0.245 $X2=0.327 $Y2=1.04
cc_65 VNB N_A_1231_367#_c_741_n 0.0216572f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_A_1231_367#_c_742_n 0.0382631f $X=-0.19 $Y=-0.245 $X2=0.275
+ $Y2=2.035
cc_67 VNB N_VPWR_c_794_n 0.322901f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_A_154_69#_c_879_n 0.00832814f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_69 VNB N_A_154_69#_c_880_n 0.0028358f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_A_154_69#_c_881_n 0.00287077f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_A_154_69#_c_882_n 0.00445045f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_GCLK_c_978_n 0.0621704f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.04
cc_73 VNB N_VGND_c_992_n 0.0232135f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_VGND_c_993_n 0.00804296f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_VGND_c_994_n 0.00567558f $X=-0.19 $Y=-0.245 $X2=0.275 $Y2=0.925
cc_76 VNB N_VGND_c_995_n 0.00880887f $X=-0.19 $Y=-0.245 $X2=0.275 $Y2=1.295
cc_77 VNB N_VGND_c_996_n 0.0113717f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_VGND_c_997_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0.275 $Y2=2.035
cc_79 VNB N_VGND_c_998_n 0.0197343f $X=-0.19 $Y=-0.245 $X2=0.275 $Y2=2.405
cc_80 VNB N_VGND_c_999_n 0.00442399f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_VGND_c_1000_n 0.0325898f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_VGND_c_1001_n 0.00401463f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_VGND_c_1002_n 0.0648162f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_VGND_c_1003_n 0.0307448f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_VGND_c_1004_n 0.0152818f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_VGND_c_1005_n 0.420513f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_VGND_c_1006_n 0.0155415f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_VGND_c_1007_n 0.00513431f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VPB N_SCE_M1020_g 0.0542753f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.66
cc_90 VPB SCE 0.0355329f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_91 VPB N_GATE_M1015_g 0.0429245f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.66
cc_92 VPB GATE 0.00454115f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_93 VPB N_A_334_69#_c_249_n 0.0213427f $X=-0.19 $Y=1.655 $X2=0.695 $Y2=0.555
cc_94 VPB N_A_334_69#_c_259_n 0.0341341f $X=-0.19 $Y=1.655 $X2=0.437 $Y2=0.875
cc_95 VPB N_A_334_69#_M1001_g 0.0209905f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_96 VPB N_A_334_69#_c_254_n 0.00378976f $X=-0.19 $Y=1.655 $X2=0.275 $Y2=1.295
cc_97 VPB N_A_334_69#_c_262_n 0.0110306f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_98 VPB N_A_334_69#_c_255_n 0.0024462f $X=-0.19 $Y=1.655 $X2=0.275 $Y2=2.405
cc_99 VPB N_A_334_69#_c_256_n 0.00166771f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_100 VPB N_A_334_69#_c_257_n 0.0361894f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_101 VPB N_A_254_357#_c_345_n 0.0662041f $X=-0.19 $Y=1.655 $X2=0.327 $Y2=1.025
cc_102 VPB N_A_254_357#_c_346_n 0.0376205f $X=-0.19 $Y=1.655 $X2=0.437 $Y2=0.875
cc_103 VPB N_A_254_357#_c_347_n 0.0108767f $X=-0.19 $Y=1.655 $X2=0.437 $Y2=1.025
cc_104 VPB N_A_254_357#_c_348_n 0.16279f $X=-0.19 $Y=1.655 $X2=0.327 $Y2=1.323
cc_105 VPB N_A_254_357#_c_349_n 0.0120529f $X=-0.19 $Y=1.655 $X2=0.327 $Y2=1.545
cc_106 VPB N_A_254_357#_c_333_n 0.00466223f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_107 VPB N_A_254_357#_c_351_n 0.0182455f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_108 VPB N_A_254_357#_M1017_g 0.0368957f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_109 VPB N_A_254_357#_c_353_n 0.00523508f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_110 VPB N_A_254_357#_c_354_n 0.00400385f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_111 VPB N_A_254_357#_c_344_n 0.00259502f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_112 VPB N_A_737_329#_M1009_g 0.0331038f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_113 VPB N_A_737_329#_M1008_g 0.0212131f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_114 VPB N_A_737_329#_c_495_n 0.0075095f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_115 VPB N_A_737_329#_c_496_n 0.00515223f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_116 VPB N_A_737_329#_c_497_n 0.0242295f $X=-0.19 $Y=1.655 $X2=0.275 $Y2=2.405
cc_117 VPB N_A_737_329#_c_484_n 4.31638e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_118 VPB N_A_737_329#_c_499_n 0.0144307f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_119 VPB N_A_737_329#_c_500_n 0.0023353f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_120 VPB N_A_737_329#_c_485_n 0.00950897f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_121 VPB N_A_737_329#_c_486_n 9.85269e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_122 VPB N_A_737_329#_c_487_n 0.00760842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_123 VPB N_A_737_329#_c_488_n 0.0331357f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_124 VPB N_A_737_329#_c_505_n 0.00388552f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_125 VPB N_A_737_329#_c_506_n 4.71579e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_126 VPB N_A_737_329#_c_490_n 0.00153624f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_127 VPB N_A_737_329#_c_491_n 0.00615591f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_128 VPB N_A_623_133#_M1014_g 0.0262133f $X=-0.19 $Y=1.655 $X2=0.327 $Y2=1.545
cc_129 VPB N_A_623_133#_c_617_n 0.0130651f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_130 VPB N_CLK_M1007_g 0.0251958f $X=-0.19 $Y=1.655 $X2=0.695 $Y2=0.555
cc_131 VPB N_CLK_M1002_g 0.0226252f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_132 VPB N_A_1231_367#_M1010_g 0.0249424f $X=-0.19 $Y=1.655 $X2=0.437
+ $Y2=0.875
cc_133 VPB N_A_1231_367#_c_740_n 0.00149024f $X=-0.19 $Y=1.655 $X2=0.327
+ $Y2=1.04
cc_134 VPB N_VPWR_c_795_n 0.0112117f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.95
cc_135 VPB N_VPWR_c_796_n 0.0216486f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_136 VPB N_VPWR_c_797_n 0.0133731f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_137 VPB N_VPWR_c_798_n 0.012156f $X=-0.19 $Y=1.655 $X2=0.275 $Y2=0.925
cc_138 VPB N_VPWR_c_799_n 0.0474826f $X=-0.19 $Y=1.655 $X2=0.275 $Y2=2.035
cc_139 VPB N_VPWR_c_800_n 0.0230288f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_140 VPB N_VPWR_c_801_n 0.0642124f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_141 VPB N_VPWR_c_802_n 0.00533588f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_142 VPB N_VPWR_c_803_n 0.033085f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_143 VPB N_VPWR_c_804_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_144 VPB N_VPWR_c_805_n 0.0218935f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_145 VPB N_VPWR_c_806_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_146 VPB N_VPWR_c_807_n 0.0273694f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_147 VPB N_VPWR_c_808_n 0.0195225f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_148 VPB N_VPWR_c_794_n 0.122834f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_149 VPB N_VPWR_c_810_n 0.0034365f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_150 VPB N_A_154_69#_c_879_n 0.00184303f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_151 VPB N_A_154_69#_c_884_n 0.0121216f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=2.32
cc_152 VPB N_A_154_69#_c_885_n 0.00381301f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_153 VPB N_A_154_69#_c_886_n 0.0033576f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_154 VPB N_A_154_69#_c_887_n 0.0296175f $X=-0.19 $Y=1.655 $X2=0.327 $Y2=1.04
cc_155 VPB N_A_154_69#_c_888_n 0.0024662f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.04
cc_156 VPB N_A_154_69#_c_889_n 0.0178063f $X=-0.19 $Y=1.655 $X2=0.275 $Y2=1.295
cc_157 VPB N_A_154_69#_c_890_n 0.00429331f $X=-0.19 $Y=1.655 $X2=0.275 $Y2=2.405
cc_158 VPB GCLK 0.0596136f $X=-0.19 $Y=1.655 $X2=0.327 $Y2=1.323
cc_159 VPB N_GCLK_c_978_n 0.0103961f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.04
cc_160 N_SCE_M1020_g N_GATE_M1015_g 0.0510162f $X=0.475 $Y=2.66 $X2=0 $Y2=0
cc_161 N_SCE_c_162_n N_GATE_c_198_n 3.15153e-19 $X=0.437 $Y=1.025 $X2=0 $Y2=0
cc_162 N_SCE_c_163_n N_GATE_c_198_n 0.0549978f $X=0.327 $Y=1.545 $X2=0 $Y2=0
cc_163 SCE N_GATE_c_198_n 0.00111964f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_164 N_SCE_c_161_n N_GATE_c_199_n 0.011377f $X=0.437 $Y=0.875 $X2=0 $Y2=0
cc_165 N_SCE_c_162_n N_GATE_c_201_n 0.00932899f $X=0.437 $Y=1.025 $X2=0 $Y2=0
cc_166 N_SCE_c_165_n N_GATE_c_201_n 0.00398159f $X=0.27 $Y=1.04 $X2=0 $Y2=0
cc_167 SCE N_VPWR_M1020_s 0.00297624f $X=0.155 $Y=0.84 $X2=-0.19 $Y2=-0.245
cc_168 N_SCE_M1020_g N_VPWR_c_796_n 0.00974346f $X=0.475 $Y=2.66 $X2=0 $Y2=0
cc_169 SCE N_VPWR_c_796_n 0.0238082f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_170 N_SCE_M1020_g N_VPWR_c_807_n 0.00396895f $X=0.475 $Y=2.66 $X2=0 $Y2=0
cc_171 N_SCE_M1020_g N_VPWR_c_794_n 0.00649579f $X=0.475 $Y=2.66 $X2=0 $Y2=0
cc_172 SCE N_VPWR_c_794_n 0.00284863f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_173 N_SCE_c_161_n N_A_154_69#_c_879_n 0.00899626f $X=0.437 $Y=0.875 $X2=0
+ $Y2=0
cc_174 N_SCE_c_162_n N_A_154_69#_c_879_n 0.00539782f $X=0.437 $Y=1.025 $X2=0
+ $Y2=0
cc_175 SCE N_A_154_69#_c_879_n 0.0622824f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_176 N_SCE_c_165_n N_A_154_69#_c_879_n 0.00666517f $X=0.27 $Y=1.04 $X2=0 $Y2=0
cc_177 N_SCE_M1020_g N_A_154_69#_c_884_n 0.00333099f $X=0.475 $Y=2.66 $X2=0
+ $Y2=0
cc_178 SCE N_A_154_69#_c_884_n 0.019348f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_179 N_SCE_c_161_n N_A_154_69#_c_897_n 0.00454085f $X=0.437 $Y=0.875 $X2=0
+ $Y2=0
cc_180 N_SCE_M1020_g N_A_154_69#_c_890_n 0.0011855f $X=0.475 $Y=2.66 $X2=0 $Y2=0
cc_181 SCE N_A_154_69#_c_890_n 0.0110156f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_182 N_SCE_c_161_n N_VGND_c_992_n 0.00670895f $X=0.437 $Y=0.875 $X2=0 $Y2=0
cc_183 N_SCE_c_162_n N_VGND_c_992_n 0.00472518f $X=0.437 $Y=1.025 $X2=0 $Y2=0
cc_184 SCE N_VGND_c_992_n 0.0155639f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_185 N_SCE_c_161_n N_VGND_c_998_n 0.00413918f $X=0.437 $Y=0.875 $X2=0 $Y2=0
cc_186 N_SCE_c_161_n N_VGND_c_1005_n 0.00758488f $X=0.437 $Y=0.875 $X2=0 $Y2=0
cc_187 N_SCE_c_162_n N_VGND_c_1005_n 0.001674f $X=0.437 $Y=1.025 $X2=0 $Y2=0
cc_188 SCE N_VGND_c_1005_n 0.00871281f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_189 N_GATE_c_198_n N_A_334_69#_c_253_n 9.95255e-19 $X=1.145 $Y=1.395 $X2=0
+ $Y2=0
cc_190 N_GATE_c_199_n N_A_334_69#_c_253_n 8.47434e-19 $X=1.145 $Y=0.875 $X2=0
+ $Y2=0
cc_191 GATE N_A_334_69#_c_253_n 0.0396198f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_192 N_GATE_c_201_n N_A_334_69#_c_253_n 4.50743e-19 $X=1.145 $Y=1.04 $X2=0
+ $Y2=0
cc_193 GATE N_A_334_69#_c_254_n 0.01273f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_194 N_GATE_M1015_g N_A_254_357#_c_347_n 0.0306919f $X=0.835 $Y=2.66 $X2=0
+ $Y2=0
cc_195 N_GATE_c_198_n N_A_254_357#_c_347_n 0.00220505f $X=1.145 $Y=1.395 $X2=0
+ $Y2=0
cc_196 GATE N_A_254_357#_c_347_n 0.00214183f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_197 N_GATE_c_199_n N_A_254_357#_M1016_g 0.0103936f $X=1.145 $Y=0.875 $X2=0
+ $Y2=0
cc_198 GATE N_A_254_357#_M1016_g 0.00360157f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_199 N_GATE_c_201_n N_A_254_357#_M1016_g 0.0143719f $X=1.145 $Y=1.04 $X2=0
+ $Y2=0
cc_200 N_GATE_c_198_n N_A_254_357#_c_332_n 0.0143719f $X=1.145 $Y=1.395 $X2=0
+ $Y2=0
cc_201 N_GATE_c_198_n N_A_254_357#_c_333_n 9.79693e-19 $X=1.145 $Y=1.395 $X2=0
+ $Y2=0
cc_202 GATE N_A_254_357#_c_333_n 7.07916e-19 $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_203 N_GATE_M1015_g N_VPWR_c_796_n 0.00101028f $X=0.835 $Y=2.66 $X2=0 $Y2=0
cc_204 N_GATE_M1015_g N_VPWR_c_797_n 0.00151575f $X=0.835 $Y=2.66 $X2=0 $Y2=0
cc_205 N_GATE_M1015_g N_VPWR_c_807_n 0.0030129f $X=0.835 $Y=2.66 $X2=0 $Y2=0
cc_206 N_GATE_M1015_g N_VPWR_c_794_n 0.00395156f $X=0.835 $Y=2.66 $X2=0 $Y2=0
cc_207 N_GATE_M1015_g N_A_154_69#_c_879_n 0.00961802f $X=0.835 $Y=2.66 $X2=0
+ $Y2=0
cc_208 N_GATE_c_198_n N_A_154_69#_c_879_n 0.00710253f $X=1.145 $Y=1.395 $X2=0
+ $Y2=0
cc_209 N_GATE_c_199_n N_A_154_69#_c_879_n 0.0034428f $X=1.145 $Y=0.875 $X2=0
+ $Y2=0
cc_210 GATE N_A_154_69#_c_879_n 0.0651909f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_211 N_GATE_c_201_n N_A_154_69#_c_879_n 0.00436266f $X=1.145 $Y=1.04 $X2=0
+ $Y2=0
cc_212 N_GATE_M1015_g N_A_154_69#_c_884_n 0.0194704f $X=0.835 $Y=2.66 $X2=0
+ $Y2=0
cc_213 N_GATE_c_198_n N_A_154_69#_c_885_n 2.59179e-19 $X=1.145 $Y=1.395 $X2=0
+ $Y2=0
cc_214 GATE N_A_154_69#_c_885_n 0.0121904f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_215 N_GATE_c_199_n N_A_154_69#_c_897_n 0.00380045f $X=1.145 $Y=0.875 $X2=0
+ $Y2=0
cc_216 GATE N_A_154_69#_c_897_n 0.0010755f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_217 N_GATE_c_201_n N_A_154_69#_c_897_n 0.00184604f $X=1.145 $Y=1.04 $X2=0
+ $Y2=0
cc_218 N_GATE_M1015_g N_A_154_69#_c_890_n 0.00676977f $X=0.835 $Y=2.66 $X2=0
+ $Y2=0
cc_219 N_GATE_c_198_n N_A_154_69#_c_890_n 0.00612733f $X=1.145 $Y=1.395 $X2=0
+ $Y2=0
cc_220 GATE N_A_154_69#_c_890_n 0.014429f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_221 N_GATE_c_199_n N_VGND_c_993_n 0.00324738f $X=1.145 $Y=0.875 $X2=0 $Y2=0
cc_222 GATE N_VGND_c_993_n 0.0100853f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_223 N_GATE_c_201_n N_VGND_c_993_n 4.24321e-19 $X=1.145 $Y=1.04 $X2=0 $Y2=0
cc_224 N_GATE_c_199_n N_VGND_c_998_n 0.00453776f $X=1.145 $Y=0.875 $X2=0 $Y2=0
cc_225 N_GATE_c_199_n N_VGND_c_1005_n 0.00488897f $X=1.145 $Y=0.875 $X2=0 $Y2=0
cc_226 GATE N_VGND_c_1005_n 0.00622984f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_227 N_A_334_69#_c_254_n N_A_254_357#_c_346_n 0.00368438f $X=1.975 $Y=1.657
+ $X2=0 $Y2=0
cc_228 N_A_334_69#_c_255_n N_A_254_357#_c_346_n 4.24076e-19 $X=2.225 $Y=1.72
+ $X2=0 $Y2=0
cc_229 N_A_334_69#_M1001_g N_A_254_357#_c_348_n 0.0104164f $X=3.175 $Y=2.525
+ $X2=0 $Y2=0
cc_230 N_A_334_69#_c_253_n N_A_254_357#_M1016_g 0.0160044f $X=1.81 $Y=0.555
+ $X2=0 $Y2=0
cc_231 N_A_334_69#_c_253_n N_A_254_357#_c_331_n 0.0148445f $X=1.81 $Y=0.555
+ $X2=0 $Y2=0
cc_232 N_A_334_69#_c_255_n N_A_254_357#_c_331_n 8.12529e-19 $X=2.225 $Y=1.72
+ $X2=0 $Y2=0
cc_233 N_A_334_69#_c_253_n N_A_254_357#_c_332_n 0.00223986f $X=1.81 $Y=0.555
+ $X2=0 $Y2=0
cc_234 N_A_334_69#_c_253_n N_A_254_357#_c_333_n 0.00399301f $X=1.81 $Y=0.555
+ $X2=0 $Y2=0
cc_235 N_A_334_69#_c_255_n N_A_254_357#_c_333_n 0.0193539f $X=2.225 $Y=1.72
+ $X2=0 $Y2=0
cc_236 N_A_334_69#_c_256_n N_A_254_357#_c_333_n 0.00351134f $X=2.535 $Y=1.72
+ $X2=0 $Y2=0
cc_237 N_A_334_69#_c_257_n N_A_254_357#_c_333_n 0.0215127f $X=2.535 $Y=1.72
+ $X2=0 $Y2=0
cc_238 N_A_334_69#_c_249_n N_A_254_357#_c_334_n 0.0231623f $X=3.325 $Y=1.66
+ $X2=0 $Y2=0
cc_239 N_A_334_69#_c_252_n N_A_254_357#_c_334_n 0.00588184f $X=3.53 $Y=1.33
+ $X2=0 $Y2=0
cc_240 N_A_334_69#_M1006_g N_A_254_357#_c_335_n 0.0166444f $X=3.53 $Y=0.875
+ $X2=0 $Y2=0
cc_241 N_A_334_69#_M1001_g N_A_254_357#_M1017_g 0.0117194f $X=3.175 $Y=2.525
+ $X2=0 $Y2=0
cc_242 N_A_334_69#_c_255_n N_A_254_357#_c_336_n 0.00146249f $X=2.225 $Y=1.72
+ $X2=0 $Y2=0
cc_243 N_A_334_69#_c_256_n N_A_254_357#_c_336_n 0.00163893f $X=2.535 $Y=1.72
+ $X2=0 $Y2=0
cc_244 N_A_334_69#_c_257_n N_A_254_357#_c_336_n 0.0224538f $X=2.535 $Y=1.72
+ $X2=0 $Y2=0
cc_245 N_A_334_69#_c_262_n N_A_254_357#_c_353_n 0.00440751f $X=2.31 $Y=2.19
+ $X2=0 $Y2=0
cc_246 N_A_334_69#_c_257_n N_A_254_357#_c_353_n 0.00509248f $X=2.535 $Y=1.72
+ $X2=0 $Y2=0
cc_247 N_A_334_69#_c_253_n N_A_254_357#_c_337_n 0.0624668f $X=1.81 $Y=0.555
+ $X2=0 $Y2=0
cc_248 N_A_334_69#_c_255_n N_A_254_357#_c_337_n 0.0180293f $X=2.225 $Y=1.72
+ $X2=0 $Y2=0
cc_249 N_A_334_69#_c_253_n N_A_254_357#_c_338_n 0.00511677f $X=1.81 $Y=0.555
+ $X2=0 $Y2=0
cc_250 N_A_334_69#_M1006_g N_A_254_357#_c_339_n 0.008147f $X=3.53 $Y=0.875 $X2=0
+ $Y2=0
cc_251 N_A_334_69#_c_253_n N_A_254_357#_c_340_n 0.0132691f $X=1.81 $Y=0.555
+ $X2=0 $Y2=0
cc_252 N_A_334_69#_M1006_g N_A_254_357#_c_342_n 0.00348636f $X=3.53 $Y=0.875
+ $X2=0 $Y2=0
cc_253 N_A_334_69#_c_250_n N_A_737_329#_M1000_g 0.00790292f $X=3.4 $Y=1.585
+ $X2=0 $Y2=0
cc_254 N_A_334_69#_M1006_g N_A_737_329#_M1000_g 0.0533039f $X=3.53 $Y=0.875
+ $X2=0 $Y2=0
cc_255 N_A_334_69#_c_259_n N_A_737_329#_M1009_g 0.00239704f $X=3.1 $Y=2.05 $X2=0
+ $Y2=0
cc_256 N_A_334_69#_c_249_n N_A_737_329#_c_488_n 0.00569746f $X=3.325 $Y=1.66
+ $X2=0 $Y2=0
cc_257 N_A_334_69#_M1006_g N_A_623_133#_c_616_n 0.0128596f $X=3.53 $Y=0.875
+ $X2=0 $Y2=0
cc_258 N_A_334_69#_c_252_n N_A_623_133#_c_616_n 0.00368501f $X=3.53 $Y=1.33
+ $X2=0 $Y2=0
cc_259 N_A_334_69#_c_249_n N_A_623_133#_c_617_n 0.0126207f $X=3.325 $Y=1.66
+ $X2=0 $Y2=0
cc_260 N_A_334_69#_c_259_n N_A_623_133#_c_617_n 0.00429944f $X=3.1 $Y=2.05 $X2=0
+ $Y2=0
cc_261 N_A_334_69#_c_250_n N_A_623_133#_c_617_n 0.00357996f $X=3.4 $Y=1.585
+ $X2=0 $Y2=0
cc_262 N_A_334_69#_c_252_n N_A_623_133#_c_618_n 0.009093f $X=3.53 $Y=1.33 $X2=0
+ $Y2=0
cc_263 N_A_334_69#_c_249_n N_A_623_133#_c_620_n 0.00423096f $X=3.325 $Y=1.66
+ $X2=0 $Y2=0
cc_264 N_A_334_69#_c_250_n N_A_623_133#_c_620_n 0.00298601f $X=3.4 $Y=1.585
+ $X2=0 $Y2=0
cc_265 N_A_334_69#_c_252_n N_A_623_133#_c_620_n 0.00392272f $X=3.53 $Y=1.33
+ $X2=0 $Y2=0
cc_266 N_A_334_69#_M1001_g N_VPWR_c_794_n 9.39239e-19 $X=3.175 $Y=2.525 $X2=0
+ $Y2=0
cc_267 N_A_334_69#_c_254_n N_A_154_69#_c_885_n 0.0273494f $X=1.975 $Y=1.657
+ $X2=0 $Y2=0
cc_268 N_A_334_69#_c_262_n N_A_154_69#_c_885_n 0.0138513f $X=2.31 $Y=2.19 $X2=0
+ $Y2=0
cc_269 N_A_334_69#_c_255_n N_A_154_69#_c_885_n 0.00622648f $X=2.225 $Y=1.72
+ $X2=0 $Y2=0
cc_270 N_A_334_69#_c_262_n N_A_154_69#_c_886_n 0.0430365f $X=2.31 $Y=2.19 $X2=0
+ $Y2=0
cc_271 N_A_334_69#_c_262_n N_A_154_69#_c_887_n 0.0188197f $X=2.31 $Y=2.19 $X2=0
+ $Y2=0
cc_272 N_A_334_69#_c_249_n N_A_154_69#_c_880_n 0.00534584f $X=3.325 $Y=1.66
+ $X2=0 $Y2=0
cc_273 N_A_334_69#_c_250_n N_A_154_69#_c_880_n 4.47176e-19 $X=3.4 $Y=1.585 $X2=0
+ $Y2=0
cc_274 N_A_334_69#_c_256_n N_A_154_69#_c_880_n 0.0261898f $X=2.535 $Y=1.72 $X2=0
+ $Y2=0
cc_275 N_A_334_69#_c_257_n N_A_154_69#_c_880_n 3.71683e-19 $X=2.535 $Y=1.72
+ $X2=0 $Y2=0
cc_276 N_A_334_69#_c_249_n N_A_154_69#_c_889_n 0.00786071f $X=3.325 $Y=1.66
+ $X2=0 $Y2=0
cc_277 N_A_334_69#_c_259_n N_A_154_69#_c_889_n 0.017341f $X=3.1 $Y=2.05 $X2=0
+ $Y2=0
cc_278 N_A_334_69#_M1001_g N_A_154_69#_c_889_n 0.0106163f $X=3.175 $Y=2.525
+ $X2=0 $Y2=0
cc_279 N_A_334_69#_c_262_n N_A_154_69#_c_889_n 0.0410629f $X=2.31 $Y=2.19 $X2=0
+ $Y2=0
cc_280 N_A_334_69#_c_257_n N_A_154_69#_c_889_n 0.00149774f $X=2.535 $Y=1.72
+ $X2=0 $Y2=0
cc_281 N_A_334_69#_M1006_g N_A_154_69#_c_881_n 2.06904e-19 $X=3.53 $Y=0.875
+ $X2=0 $Y2=0
cc_282 N_A_334_69#_c_252_n N_A_154_69#_c_882_n 9.30357e-19 $X=3.53 $Y=1.33 $X2=0
+ $Y2=0
cc_283 N_A_334_69#_M1006_g N_VGND_c_1002_n 5.69678e-19 $X=3.53 $Y=0.875 $X2=0
+ $Y2=0
cc_284 N_A_334_69#_c_253_n N_VGND_c_1002_n 0.0112286f $X=1.81 $Y=0.555 $X2=0
+ $Y2=0
cc_285 N_A_334_69#_c_253_n N_VGND_c_1005_n 0.0116871f $X=1.81 $Y=0.555 $X2=0
+ $Y2=0
cc_286 N_A_254_357#_c_341_n N_A_737_329#_M1021_d 0.00685357f $X=5.085 $Y=0.61
+ $X2=-0.19 $Y2=-0.245
cc_287 N_A_254_357#_c_341_n N_A_737_329#_M1000_g 0.00945341f $X=5.085 $Y=0.61
+ $X2=0 $Y2=0
cc_288 N_A_254_357#_c_342_n N_A_737_329#_M1000_g 0.00338302f $X=3.765 $Y=0.455
+ $X2=0 $Y2=0
cc_289 N_A_254_357#_M1017_g N_A_737_329#_M1009_g 0.0404219f $X=3.605 $Y=2.525
+ $X2=0 $Y2=0
cc_290 N_A_254_357#_c_354_n N_A_737_329#_c_496_n 0.0189946f $X=5.275 $Y=1.97
+ $X2=0 $Y2=0
cc_291 N_A_254_357#_c_344_n N_A_737_329#_c_484_n 0.0401343f $X=5.275 $Y=1.795
+ $X2=0 $Y2=0
cc_292 N_A_254_357#_M1007_s N_A_737_329#_c_499_n 0.0120995f $X=5.13 $Y=1.835
+ $X2=0 $Y2=0
cc_293 N_A_254_357#_c_354_n N_A_737_329#_c_499_n 0.0217908f $X=5.275 $Y=1.97
+ $X2=0 $Y2=0
cc_294 N_A_254_357#_c_354_n N_A_737_329#_c_500_n 0.010728f $X=5.275 $Y=1.97
+ $X2=0 $Y2=0
cc_295 N_A_254_357#_c_344_n N_A_737_329#_c_500_n 0.00363285f $X=5.275 $Y=1.795
+ $X2=0 $Y2=0
cc_296 N_A_254_357#_c_344_n N_A_737_329#_c_486_n 0.0107753f $X=5.275 $Y=1.795
+ $X2=0 $Y2=0
cc_297 N_A_254_357#_c_341_n N_A_737_329#_c_489_n 0.0256635f $X=5.085 $Y=0.61
+ $X2=0 $Y2=0
cc_298 N_A_254_357#_c_344_n N_A_737_329#_c_489_n 0.0189781f $X=5.275 $Y=1.795
+ $X2=0 $Y2=0
cc_299 N_A_254_357#_c_344_n N_A_737_329#_c_505_n 0.0141369f $X=5.275 $Y=1.795
+ $X2=0 $Y2=0
cc_300 N_A_254_357#_c_344_n N_A_623_133#_M1014_g 0.00118696f $X=5.275 $Y=1.795
+ $X2=0 $Y2=0
cc_301 N_A_254_357#_c_335_n N_A_623_133#_c_616_n 0.00377898f $X=3.04 $Y=1.195
+ $X2=0 $Y2=0
cc_302 N_A_254_357#_c_339_n N_A_623_133#_c_616_n 0.0239654f $X=3.68 $Y=0.455
+ $X2=0 $Y2=0
cc_303 N_A_254_357#_c_348_n N_A_623_133#_c_617_n 0.00325534f $X=3.53 $Y=3.15
+ $X2=0 $Y2=0
cc_304 N_A_254_357#_M1017_g N_A_623_133#_c_617_n 0.00187398f $X=3.605 $Y=2.525
+ $X2=0 $Y2=0
cc_305 N_A_254_357#_c_341_n N_A_623_133#_c_618_n 0.0173751f $X=5.085 $Y=0.61
+ $X2=0 $Y2=0
cc_306 N_A_254_357#_c_342_n N_A_623_133#_c_618_n 0.00433841f $X=3.765 $Y=0.455
+ $X2=0 $Y2=0
cc_307 N_A_254_357#_c_341_n N_A_623_133#_c_619_n 0.00256984f $X=5.085 $Y=0.61
+ $X2=0 $Y2=0
cc_308 N_A_254_357#_c_334_n N_A_623_133#_c_620_n 6.359e-19 $X=2.965 $Y=1.27
+ $X2=0 $Y2=0
cc_309 N_A_254_357#_c_341_n N_A_623_133#_c_621_n 0.015576f $X=5.085 $Y=0.61
+ $X2=0 $Y2=0
cc_310 N_A_254_357#_c_342_n N_A_623_133#_c_621_n 0.00366893f $X=3.765 $Y=0.455
+ $X2=0 $Y2=0
cc_311 N_A_254_357#_c_343_n N_A_623_133#_c_621_n 0.00586097f $X=5.25 $Y=0.47
+ $X2=0 $Y2=0
cc_312 N_A_254_357#_c_344_n N_A_623_133#_c_621_n 0.00329656f $X=5.275 $Y=1.795
+ $X2=0 $Y2=0
cc_313 N_A_254_357#_c_343_n N_CLK_c_682_n 0.0138228f $X=5.25 $Y=0.47 $X2=-0.19
+ $Y2=-0.245
cc_314 N_A_254_357#_c_354_n N_CLK_M1007_g 0.00497728f $X=5.275 $Y=1.97 $X2=0
+ $Y2=0
cc_315 N_A_254_357#_c_344_n N_CLK_M1007_g 0.00953007f $X=5.275 $Y=1.795 $X2=0
+ $Y2=0
cc_316 N_A_254_357#_c_344_n CLK 0.031951f $X=5.275 $Y=1.795 $X2=0 $Y2=0
cc_317 N_A_254_357#_c_354_n N_CLK_c_687_n 9.09473e-19 $X=5.275 $Y=1.97 $X2=0
+ $Y2=0
cc_318 N_A_254_357#_c_344_n N_CLK_c_687_n 0.0138228f $X=5.275 $Y=1.795 $X2=0
+ $Y2=0
cc_319 N_A_254_357#_c_345_n N_VPWR_c_797_n 0.0108675f $X=1.345 $Y=3.075 $X2=0
+ $Y2=0
cc_320 N_A_254_357#_c_346_n N_VPWR_c_797_n 0.00110701f $X=2.01 $Y=1.86 $X2=0
+ $Y2=0
cc_321 N_A_254_357#_c_348_n N_VPWR_c_797_n 0.0200844f $X=3.53 $Y=3.15 $X2=0
+ $Y2=0
cc_322 N_A_254_357#_c_351_n N_VPWR_c_797_n 0.00168178f $X=2.085 $Y=1.935 $X2=0
+ $Y2=0
cc_323 N_A_254_357#_M1017_g N_VPWR_c_798_n 0.00975547f $X=3.605 $Y=2.525 $X2=0
+ $Y2=0
cc_324 N_A_254_357#_c_348_n N_VPWR_c_801_n 0.0499731f $X=3.53 $Y=3.15 $X2=0
+ $Y2=0
cc_325 N_A_254_357#_c_349_n N_VPWR_c_807_n 0.00718072f $X=1.42 $Y=3.15 $X2=0
+ $Y2=0
cc_326 N_A_254_357#_c_348_n N_VPWR_c_794_n 0.0654157f $X=3.53 $Y=3.15 $X2=0
+ $Y2=0
cc_327 N_A_254_357#_c_349_n N_VPWR_c_794_n 0.0112079f $X=1.42 $Y=3.15 $X2=0
+ $Y2=0
cc_328 N_A_254_357#_c_347_n N_A_154_69#_c_879_n 9.86556e-19 $X=1.42 $Y=1.86
+ $X2=0 $Y2=0
cc_329 N_A_254_357#_c_345_n N_A_154_69#_c_884_n 0.0100891f $X=1.345 $Y=3.075
+ $X2=0 $Y2=0
cc_330 N_A_254_357#_c_345_n N_A_154_69#_c_885_n 0.0127405f $X=1.345 $Y=3.075
+ $X2=0 $Y2=0
cc_331 N_A_254_357#_c_346_n N_A_154_69#_c_885_n 0.0167831f $X=2.01 $Y=1.86 $X2=0
+ $Y2=0
cc_332 N_A_254_357#_c_347_n N_A_154_69#_c_885_n 0.0030216f $X=1.42 $Y=1.86 $X2=0
+ $Y2=0
cc_333 N_A_254_357#_c_332_n N_A_154_69#_c_885_n 8.29285e-19 $X=1.67 $Y=1.27
+ $X2=0 $Y2=0
cc_334 N_A_254_357#_c_351_n N_A_154_69#_c_885_n 0.00554896f $X=2.085 $Y=1.935
+ $X2=0 $Y2=0
cc_335 N_A_254_357#_c_353_n N_A_154_69#_c_885_n 6.89983e-19 $X=2.085 $Y=1.86
+ $X2=0 $Y2=0
cc_336 N_A_254_357#_c_345_n N_A_154_69#_c_886_n 0.00212535f $X=1.345 $Y=3.075
+ $X2=0 $Y2=0
cc_337 N_A_254_357#_c_351_n N_A_154_69#_c_886_n 0.0212731f $X=2.085 $Y=1.935
+ $X2=0 $Y2=0
cc_338 N_A_254_357#_c_348_n N_A_154_69#_c_887_n 0.0225257f $X=3.53 $Y=3.15 $X2=0
+ $Y2=0
cc_339 N_A_254_357#_c_351_n N_A_154_69#_c_887_n 0.00261886f $X=2.085 $Y=1.935
+ $X2=0 $Y2=0
cc_340 N_A_254_357#_M1017_g N_A_154_69#_c_887_n 0.00522941f $X=3.605 $Y=2.525
+ $X2=0 $Y2=0
cc_341 N_A_254_357#_c_348_n N_A_154_69#_c_888_n 0.00345419f $X=3.53 $Y=3.15
+ $X2=0 $Y2=0
cc_342 N_A_254_357#_c_334_n N_A_154_69#_c_880_n 0.00329221f $X=2.965 $Y=1.27
+ $X2=0 $Y2=0
cc_343 N_A_254_357#_c_333_n N_A_154_69#_c_889_n 2.7765e-19 $X=2.085 $Y=1.785
+ $X2=0 $Y2=0
cc_344 N_A_254_357#_c_351_n N_A_154_69#_c_889_n 0.0037956f $X=2.085 $Y=1.935
+ $X2=0 $Y2=0
cc_345 N_A_254_357#_M1017_g N_A_154_69#_c_889_n 5.50134e-19 $X=3.605 $Y=2.525
+ $X2=0 $Y2=0
cc_346 N_A_254_357#_c_334_n N_A_154_69#_c_881_n 0.00600575f $X=2.965 $Y=1.27
+ $X2=0 $Y2=0
cc_347 N_A_254_357#_c_335_n N_A_154_69#_c_881_n 0.00291183f $X=3.04 $Y=1.195
+ $X2=0 $Y2=0
cc_348 N_A_254_357#_c_337_n N_A_154_69#_c_881_n 0.0201699f $X=2.24 $Y=0.84 $X2=0
+ $Y2=0
cc_349 N_A_254_357#_c_338_n N_A_154_69#_c_881_n 0.00319826f $X=2.24 $Y=0.84
+ $X2=0 $Y2=0
cc_350 N_A_254_357#_c_339_n N_A_154_69#_c_881_n 0.0228938f $X=3.68 $Y=0.455
+ $X2=0 $Y2=0
cc_351 N_A_254_357#_c_333_n N_A_154_69#_c_882_n 0.00487509f $X=2.085 $Y=1.785
+ $X2=0 $Y2=0
cc_352 N_A_254_357#_c_334_n N_A_154_69#_c_882_n 0.0102542f $X=2.965 $Y=1.27
+ $X2=0 $Y2=0
cc_353 N_A_254_357#_c_335_n N_A_154_69#_c_882_n 0.00294066f $X=3.04 $Y=1.195
+ $X2=0 $Y2=0
cc_354 N_A_254_357#_c_337_n N_A_154_69#_c_882_n 0.0113258f $X=2.24 $Y=0.84 $X2=0
+ $Y2=0
cc_355 N_A_254_357#_c_338_n N_A_154_69#_c_882_n 0.0012501f $X=2.24 $Y=0.84 $X2=0
+ $Y2=0
cc_356 N_A_254_357#_c_341_n N_VGND_M1000_d 0.00986502f $X=5.085 $Y=0.61 $X2=0
+ $Y2=0
cc_357 N_A_254_357#_M1016_g N_VGND_c_993_n 0.00324738f $X=1.595 $Y=0.555 $X2=0
+ $Y2=0
cc_358 N_A_254_357#_c_341_n N_VGND_c_1000_n 0.0156199f $X=5.085 $Y=0.61 $X2=0
+ $Y2=0
cc_359 N_A_254_357#_c_343_n N_VGND_c_1000_n 0.0136958f $X=5.25 $Y=0.47 $X2=0
+ $Y2=0
cc_360 N_A_254_357#_M1016_g N_VGND_c_1002_n 0.00454892f $X=1.595 $Y=0.555 $X2=0
+ $Y2=0
cc_361 N_A_254_357#_c_335_n N_VGND_c_1002_n 5.69678e-19 $X=3.04 $Y=1.195 $X2=0
+ $Y2=0
cc_362 N_A_254_357#_c_338_n N_VGND_c_1002_n 0.00374823f $X=2.24 $Y=0.84 $X2=0
+ $Y2=0
cc_363 N_A_254_357#_c_339_n N_VGND_c_1002_n 0.0476345f $X=3.68 $Y=0.455 $X2=0
+ $Y2=0
cc_364 N_A_254_357#_c_340_n N_VGND_c_1002_n 0.0107383f $X=2.405 $Y=0.455 $X2=0
+ $Y2=0
cc_365 N_A_254_357#_c_341_n N_VGND_c_1002_n 0.00399169f $X=5.085 $Y=0.61 $X2=0
+ $Y2=0
cc_366 N_A_254_357#_c_342_n N_VGND_c_1002_n 0.00658579f $X=3.765 $Y=0.455 $X2=0
+ $Y2=0
cc_367 N_A_254_357#_M1016_g N_VGND_c_1005_n 0.00892734f $X=1.595 $Y=0.555 $X2=0
+ $Y2=0
cc_368 N_A_254_357#_c_338_n N_VGND_c_1005_n 0.00383128f $X=2.24 $Y=0.84 $X2=0
+ $Y2=0
cc_369 N_A_254_357#_c_339_n N_VGND_c_1005_n 0.0444579f $X=3.68 $Y=0.455 $X2=0
+ $Y2=0
cc_370 N_A_254_357#_c_340_n N_VGND_c_1005_n 0.00948613f $X=2.405 $Y=0.455 $X2=0
+ $Y2=0
cc_371 N_A_254_357#_c_341_n N_VGND_c_1005_n 0.0292736f $X=5.085 $Y=0.61 $X2=0
+ $Y2=0
cc_372 N_A_254_357#_c_342_n N_VGND_c_1005_n 0.00597965f $X=3.765 $Y=0.455 $X2=0
+ $Y2=0
cc_373 N_A_254_357#_c_343_n N_VGND_c_1005_n 0.0101427f $X=5.25 $Y=0.47 $X2=0
+ $Y2=0
cc_374 N_A_254_357#_c_341_n N_VGND_c_1006_n 0.0240258f $X=5.085 $Y=0.61 $X2=0
+ $Y2=0
cc_375 N_A_254_357#_c_342_n A_721_133# 0.00187054f $X=3.765 $Y=0.455 $X2=-0.19
+ $Y2=-0.245
cc_376 N_A_737_329#_M1000_g N_A_623_133#_M1014_g 0.00373808f $X=3.89 $Y=0.875
+ $X2=0 $Y2=0
cc_377 N_A_737_329#_c_495_n N_A_623_133#_M1014_g 0.0162178f $X=4.635 $Y=1.73
+ $X2=0 $Y2=0
cc_378 N_A_737_329#_c_497_n N_A_623_133#_M1014_g 0.00206255f $X=4.73 $Y=2.91
+ $X2=0 $Y2=0
cc_379 N_A_737_329#_c_487_n N_A_623_133#_M1014_g 3.79499e-19 $X=3.825 $Y=1.73
+ $X2=0 $Y2=0
cc_380 N_A_737_329#_c_488_n N_A_623_133#_M1014_g 0.0182313f $X=3.85 $Y=1.81
+ $X2=0 $Y2=0
cc_381 N_A_737_329#_M1000_g N_A_623_133#_c_616_n 0.00291332f $X=3.89 $Y=0.875
+ $X2=0 $Y2=0
cc_382 N_A_737_329#_M1000_g N_A_623_133#_c_617_n 0.00320989f $X=3.89 $Y=0.875
+ $X2=0 $Y2=0
cc_383 N_A_737_329#_M1009_g N_A_623_133#_c_617_n 0.00294285f $X=3.965 $Y=2.525
+ $X2=0 $Y2=0
cc_384 N_A_737_329#_c_487_n N_A_623_133#_c_617_n 0.0231468f $X=3.825 $Y=1.73
+ $X2=0 $Y2=0
cc_385 N_A_737_329#_c_488_n N_A_623_133#_c_617_n 0.00593617f $X=3.85 $Y=1.81
+ $X2=0 $Y2=0
cc_386 N_A_737_329#_M1000_g N_A_623_133#_c_618_n 0.0132957f $X=3.89 $Y=0.875
+ $X2=0 $Y2=0
cc_387 N_A_737_329#_c_495_n N_A_623_133#_c_618_n 0.044807f $X=4.635 $Y=1.73
+ $X2=0 $Y2=0
cc_388 N_A_737_329#_c_484_n N_A_623_133#_c_618_n 0.0151498f $X=4.845 $Y=1.645
+ $X2=0 $Y2=0
cc_389 N_A_737_329#_c_487_n N_A_623_133#_c_618_n 0.0206547f $X=3.825 $Y=1.73
+ $X2=0 $Y2=0
cc_390 N_A_737_329#_c_488_n N_A_623_133#_c_618_n 0.00290345f $X=3.85 $Y=1.81
+ $X2=0 $Y2=0
cc_391 N_A_737_329#_c_489_n N_A_623_133#_c_618_n 0.00362202f $X=4.845 $Y=0.985
+ $X2=0 $Y2=0
cc_392 N_A_737_329#_M1000_g N_A_623_133#_c_619_n 0.0157865f $X=3.89 $Y=0.875
+ $X2=0 $Y2=0
cc_393 N_A_737_329#_c_495_n N_A_623_133#_c_619_n 0.00466401f $X=4.635 $Y=1.73
+ $X2=0 $Y2=0
cc_394 N_A_737_329#_c_484_n N_A_623_133#_c_619_n 0.0135389f $X=4.845 $Y=1.645
+ $X2=0 $Y2=0
cc_395 N_A_737_329#_c_489_n N_A_623_133#_c_619_n 0.00106843f $X=4.845 $Y=0.985
+ $X2=0 $Y2=0
cc_396 N_A_737_329#_M1000_g N_A_623_133#_c_621_n 0.0194717f $X=3.89 $Y=0.875
+ $X2=0 $Y2=0
cc_397 N_A_737_329#_c_484_n N_A_623_133#_c_621_n 0.00295101f $X=4.845 $Y=1.645
+ $X2=0 $Y2=0
cc_398 N_A_737_329#_c_489_n N_A_623_133#_c_621_n 0.00610114f $X=4.845 $Y=0.985
+ $X2=0 $Y2=0
cc_399 N_A_737_329#_c_496_n N_CLK_M1007_g 0.00351628f $X=4.73 $Y=1.95 $X2=0
+ $Y2=0
cc_400 N_A_737_329#_c_497_n N_CLK_M1007_g 0.00550456f $X=4.73 $Y=2.91 $X2=0
+ $Y2=0
cc_401 N_A_737_329#_c_499_n N_CLK_M1007_g 0.0202451f $X=5.62 $Y=2.31 $X2=0 $Y2=0
cc_402 N_A_737_329#_c_500_n N_CLK_M1007_g 0.0034404f $X=5.705 $Y=2.225 $X2=0
+ $Y2=0
cc_403 N_A_737_329#_c_486_n N_CLK_M1007_g 0.00203338f $X=5.79 $Y=1.645 $X2=0
+ $Y2=0
cc_404 N_A_737_329#_c_482_n N_CLK_c_684_n 0.0250823f $X=6.255 $Y=0.79 $X2=0
+ $Y2=0
cc_405 N_A_737_329#_M1008_g N_CLK_M1002_g 0.0129731f $X=6.51 $Y=2.155 $X2=0
+ $Y2=0
cc_406 N_A_737_329#_c_499_n N_CLK_M1002_g 0.00166196f $X=5.62 $Y=2.31 $X2=0
+ $Y2=0
cc_407 N_A_737_329#_c_500_n N_CLK_M1002_g 0.00638178f $X=5.705 $Y=2.225 $X2=0
+ $Y2=0
cc_408 N_A_737_329#_c_485_n N_CLK_M1002_g 0.0142826f $X=6.365 $Y=1.645 $X2=0
+ $Y2=0
cc_409 N_A_737_329#_c_491_n N_CLK_M1002_g 0.011851f $X=6.53 $Y=1.51 $X2=0 $Y2=0
cc_410 N_A_737_329#_c_483_n CLK 0.00401972f $X=6.44 $Y=0.865 $X2=0 $Y2=0
cc_411 N_A_737_329#_c_485_n CLK 0.0314762f $X=6.365 $Y=1.645 $X2=0 $Y2=0
cc_412 N_A_737_329#_c_486_n CLK 0.0131404f $X=5.79 $Y=1.645 $X2=0 $Y2=0
cc_413 N_A_737_329#_c_490_n CLK 0.00365848f $X=6.53 $Y=1.51 $X2=0 $Y2=0
cc_414 N_A_737_329#_c_492_n CLK 0.00373426f $X=6.53 $Y=1.345 $X2=0 $Y2=0
cc_415 N_A_737_329#_c_483_n N_CLK_c_687_n 0.0250823f $X=6.44 $Y=0.865 $X2=0
+ $Y2=0
cc_416 N_A_737_329#_c_485_n N_CLK_c_687_n 0.00357147f $X=6.365 $Y=1.645 $X2=0
+ $Y2=0
cc_417 N_A_737_329#_c_486_n N_CLK_c_687_n 0.00396396f $X=5.79 $Y=1.645 $X2=0
+ $Y2=0
cc_418 N_A_737_329#_c_490_n N_CLK_c_687_n 0.00126484f $X=6.53 $Y=1.51 $X2=0
+ $Y2=0
cc_419 N_A_737_329#_c_492_n N_CLK_c_687_n 0.0217019f $X=6.53 $Y=1.345 $X2=0
+ $Y2=0
cc_420 N_A_737_329#_M1008_g N_A_1231_367#_M1010_g 0.0215058f $X=6.51 $Y=2.155
+ $X2=0 $Y2=0
cc_421 N_A_737_329#_c_490_n N_A_1231_367#_M1010_g 2.84548e-19 $X=6.53 $Y=1.51
+ $X2=0 $Y2=0
cc_422 N_A_737_329#_c_491_n N_A_1231_367#_M1010_g 0.00785851f $X=6.53 $Y=1.51
+ $X2=0 $Y2=0
cc_423 N_A_737_329#_c_483_n N_A_1231_367#_c_738_n 0.00398895f $X=6.44 $Y=0.865
+ $X2=0 $Y2=0
cc_424 N_A_737_329#_c_482_n N_A_1231_367#_c_739_n 0.00486474f $X=6.255 $Y=0.79
+ $X2=0 $Y2=0
cc_425 N_A_737_329#_c_483_n N_A_1231_367#_c_739_n 0.00928613f $X=6.44 $Y=0.865
+ $X2=0 $Y2=0
cc_426 N_A_737_329#_c_492_n N_A_1231_367#_c_739_n 0.00132441f $X=6.53 $Y=1.345
+ $X2=0 $Y2=0
cc_427 N_A_737_329#_M1008_g N_A_1231_367#_c_752_n 0.0112949f $X=6.51 $Y=2.155
+ $X2=0 $Y2=0
cc_428 N_A_737_329#_c_490_n N_A_1231_367#_c_752_n 0.0104529f $X=6.53 $Y=1.51
+ $X2=0 $Y2=0
cc_429 N_A_737_329#_c_491_n N_A_1231_367#_c_752_n 0.0021019f $X=6.53 $Y=1.51
+ $X2=0 $Y2=0
cc_430 N_A_737_329#_M1008_g N_A_1231_367#_c_740_n 0.00381105f $X=6.51 $Y=2.155
+ $X2=0 $Y2=0
cc_431 N_A_737_329#_c_490_n N_A_1231_367#_c_740_n 0.0160729f $X=6.53 $Y=1.51
+ $X2=0 $Y2=0
cc_432 N_A_737_329#_c_491_n N_A_1231_367#_c_740_n 0.00105567f $X=6.53 $Y=1.51
+ $X2=0 $Y2=0
cc_433 N_A_737_329#_M1008_g N_A_1231_367#_c_758_n 0.00701244f $X=6.51 $Y=2.155
+ $X2=0 $Y2=0
cc_434 N_A_737_329#_c_499_n N_A_1231_367#_c_758_n 0.00824032f $X=5.62 $Y=2.31
+ $X2=0 $Y2=0
cc_435 N_A_737_329#_c_500_n N_A_1231_367#_c_758_n 0.0140552f $X=5.705 $Y=2.225
+ $X2=0 $Y2=0
cc_436 N_A_737_329#_c_485_n N_A_1231_367#_c_758_n 0.0157089f $X=6.365 $Y=1.645
+ $X2=0 $Y2=0
cc_437 N_A_737_329#_c_490_n N_A_1231_367#_c_758_n 0.00520993f $X=6.53 $Y=1.51
+ $X2=0 $Y2=0
cc_438 N_A_737_329#_c_491_n N_A_1231_367#_c_758_n 3.02524e-19 $X=6.53 $Y=1.51
+ $X2=0 $Y2=0
cc_439 N_A_737_329#_c_490_n N_A_1231_367#_c_741_n 0.0334087f $X=6.53 $Y=1.51
+ $X2=0 $Y2=0
cc_440 N_A_737_329#_c_491_n N_A_1231_367#_c_741_n 0.0044561f $X=6.53 $Y=1.51
+ $X2=0 $Y2=0
cc_441 N_A_737_329#_c_492_n N_A_1231_367#_c_741_n 0.00965108f $X=6.53 $Y=1.345
+ $X2=0 $Y2=0
cc_442 N_A_737_329#_c_491_n N_A_1231_367#_c_742_n 0.0105445f $X=6.53 $Y=1.51
+ $X2=0 $Y2=0
cc_443 N_A_737_329#_c_492_n N_A_1231_367#_c_742_n 0.00420545f $X=6.53 $Y=1.345
+ $X2=0 $Y2=0
cc_444 N_A_737_329#_c_495_n N_VPWR_M1009_d 0.00223101f $X=4.635 $Y=1.73 $X2=0
+ $Y2=0
cc_445 N_A_737_329#_c_499_n N_VPWR_M1007_d 0.00428227f $X=5.62 $Y=2.31 $X2=0
+ $Y2=0
cc_446 N_A_737_329#_c_500_n N_VPWR_M1007_d 0.006836f $X=5.705 $Y=2.225 $X2=0
+ $Y2=0
cc_447 N_A_737_329#_M1009_g N_VPWR_c_798_n 0.0149689f $X=3.965 $Y=2.525 $X2=0
+ $Y2=0
cc_448 N_A_737_329#_c_495_n N_VPWR_c_798_n 0.0220026f $X=4.635 $Y=1.73 $X2=0
+ $Y2=0
cc_449 N_A_737_329#_c_497_n N_VPWR_c_798_n 0.0258834f $X=4.73 $Y=2.91 $X2=0
+ $Y2=0
cc_450 N_A_737_329#_c_499_n N_VPWR_c_799_n 0.0151808f $X=5.62 $Y=2.31 $X2=0
+ $Y2=0
cc_451 N_A_737_329#_M1008_g N_VPWR_c_800_n 0.00481097f $X=6.51 $Y=2.155 $X2=0
+ $Y2=0
cc_452 N_A_737_329#_M1009_g N_VPWR_c_801_n 0.00431487f $X=3.965 $Y=2.525 $X2=0
+ $Y2=0
cc_453 N_A_737_329#_c_497_n N_VPWR_c_803_n 0.0210042f $X=4.73 $Y=2.91 $X2=0
+ $Y2=0
cc_454 N_A_737_329#_M1008_g N_VPWR_c_805_n 0.00312414f $X=6.51 $Y=2.155 $X2=0
+ $Y2=0
cc_455 N_A_737_329#_M1009_g N_VPWR_c_794_n 0.00477801f $X=3.965 $Y=2.525 $X2=0
+ $Y2=0
cc_456 N_A_737_329#_M1008_g N_VPWR_c_794_n 0.00410284f $X=6.51 $Y=2.155 $X2=0
+ $Y2=0
cc_457 N_A_737_329#_c_497_n N_VPWR_c_794_n 0.0113912f $X=4.73 $Y=2.91 $X2=0
+ $Y2=0
cc_458 N_A_737_329#_c_482_n N_VGND_c_995_n 0.00381028f $X=6.255 $Y=0.79 $X2=0
+ $Y2=0
cc_459 N_A_737_329#_M1000_g N_VGND_c_1002_n 6.38981e-19 $X=3.89 $Y=0.875 $X2=0
+ $Y2=0
cc_460 N_A_737_329#_c_482_n N_VGND_c_1003_n 0.00560159f $X=6.255 $Y=0.79 $X2=0
+ $Y2=0
cc_461 N_A_737_329#_M1021_d N_VGND_c_1005_n 0.00288526f $X=4.555 $Y=0.245 $X2=0
+ $Y2=0
cc_462 N_A_737_329#_c_482_n N_VGND_c_1005_n 0.0112938f $X=6.255 $Y=0.79 $X2=0
+ $Y2=0
cc_463 N_A_737_329#_c_483_n N_VGND_c_1005_n 7.60701e-19 $X=6.44 $Y=0.865 $X2=0
+ $Y2=0
cc_464 N_A_623_133#_M1014_g N_VPWR_c_798_n 0.0187145f $X=4.515 $Y=2.435 $X2=0
+ $Y2=0
cc_465 N_A_623_133#_c_617_n N_VPWR_c_798_n 0.0159835f $X=3.39 $Y=2.525 $X2=0
+ $Y2=0
cc_466 N_A_623_133#_c_617_n N_VPWR_c_801_n 0.00386107f $X=3.39 $Y=2.525 $X2=0
+ $Y2=0
cc_467 N_A_623_133#_M1014_g N_VPWR_c_803_n 0.00461019f $X=4.515 $Y=2.435 $X2=0
+ $Y2=0
cc_468 N_A_623_133#_M1014_g N_VPWR_c_794_n 0.00930161f $X=4.515 $Y=2.435 $X2=0
+ $Y2=0
cc_469 N_A_623_133#_c_617_n N_VPWR_c_794_n 0.00626052f $X=3.39 $Y=2.525 $X2=0
+ $Y2=0
cc_470 N_A_623_133#_c_617_n N_A_154_69#_c_880_n 0.0635885f $X=3.39 $Y=2.525
+ $X2=0 $Y2=0
cc_471 N_A_623_133#_c_616_n N_A_154_69#_c_881_n 0.0281873f $X=3.315 $Y=0.875
+ $X2=0 $Y2=0
cc_472 N_A_623_133#_c_617_n N_A_154_69#_c_882_n 0.00129623f $X=3.39 $Y=2.525
+ $X2=0 $Y2=0
cc_473 N_A_623_133#_c_620_n N_A_154_69#_c_882_n 0.0129171f $X=3.14 $Y=1.275
+ $X2=0 $Y2=0
cc_474 N_A_623_133#_c_621_n N_VGND_c_1000_n 0.00400062f $X=4.42 $Y=1.195 $X2=0
+ $Y2=0
cc_475 N_A_623_133#_c_621_n N_VGND_c_1005_n 0.00814141f $X=4.42 $Y=1.195 $X2=0
+ $Y2=0
cc_476 N_A_623_133#_c_621_n N_VGND_c_1006_n 0.00659856f $X=4.42 $Y=1.195 $X2=0
+ $Y2=0
cc_477 CLK N_A_1231_367#_c_739_n 0.0139872f $X=5.915 $Y=0.84 $X2=0 $Y2=0
cc_478 N_CLK_c_687_n N_A_1231_367#_c_739_n 2.0249e-19 $X=5.895 $Y=1.125 $X2=0
+ $Y2=0
cc_479 N_CLK_M1007_g N_A_1231_367#_c_758_n 3.98283e-19 $X=5.49 $Y=2.155 $X2=0
+ $Y2=0
cc_480 N_CLK_M1002_g N_A_1231_367#_c_758_n 0.00920214f $X=6.08 $Y=2.155 $X2=0
+ $Y2=0
cc_481 CLK N_A_1231_367#_c_741_n 0.0214538f $X=5.915 $Y=0.84 $X2=0 $Y2=0
cc_482 N_CLK_M1007_g N_VPWR_c_799_n 0.00116328f $X=5.49 $Y=2.155 $X2=0 $Y2=0
cc_483 N_CLK_M1002_g N_VPWR_c_799_n 0.00116328f $X=6.08 $Y=2.155 $X2=0 $Y2=0
cc_484 N_CLK_M1007_g N_VPWR_c_803_n 0.00312414f $X=5.49 $Y=2.155 $X2=0 $Y2=0
cc_485 N_CLK_M1002_g N_VPWR_c_805_n 0.00312414f $X=6.08 $Y=2.155 $X2=0 $Y2=0
cc_486 N_CLK_M1007_g N_VPWR_c_794_n 0.00410284f $X=5.49 $Y=2.155 $X2=0 $Y2=0
cc_487 N_CLK_M1002_g N_VPWR_c_794_n 0.00410284f $X=6.08 $Y=2.155 $X2=0 $Y2=0
cc_488 N_CLK_c_682_n N_VGND_c_994_n 0.00291027f $X=5.465 $Y=0.79 $X2=0 $Y2=0
cc_489 N_CLK_c_684_n N_VGND_c_994_n 0.00291027f $X=5.895 $Y=0.79 $X2=0 $Y2=0
cc_490 CLK N_VGND_c_994_n 0.0111362f $X=5.915 $Y=0.84 $X2=0 $Y2=0
cc_491 N_CLK_c_687_n N_VGND_c_994_n 0.00297724f $X=5.895 $Y=1.125 $X2=0 $Y2=0
cc_492 N_CLK_c_682_n N_VGND_c_1000_n 0.00560159f $X=5.465 $Y=0.79 $X2=0 $Y2=0
cc_493 N_CLK_c_684_n N_VGND_c_1003_n 0.00560159f $X=5.895 $Y=0.79 $X2=0 $Y2=0
cc_494 N_CLK_c_682_n N_VGND_c_1005_n 0.0116802f $X=5.465 $Y=0.79 $X2=0 $Y2=0
cc_495 N_CLK_c_684_n N_VGND_c_1005_n 0.00585539f $X=5.895 $Y=0.79 $X2=0 $Y2=0
cc_496 CLK N_VGND_c_1005_n 0.0155107f $X=5.915 $Y=0.84 $X2=0 $Y2=0
cc_497 N_A_1231_367#_c_752_n N_VPWR_M1008_d 0.00724486f $X=6.8 $Y=1.995 $X2=0
+ $Y2=0
cc_498 N_A_1231_367#_c_740_n N_VPWR_M1008_d 8.86476e-19 $X=6.885 $Y=1.91 $X2=0
+ $Y2=0
cc_499 N_A_1231_367#_M1010_g N_VPWR_c_800_n 0.0189772f $X=7.02 $Y=2.465 $X2=0
+ $Y2=0
cc_500 N_A_1231_367#_c_752_n N_VPWR_c_800_n 0.0226966f $X=6.8 $Y=1.995 $X2=0
+ $Y2=0
cc_501 N_A_1231_367#_M1010_g N_VPWR_c_808_n 0.00486043f $X=7.02 $Y=2.465 $X2=0
+ $Y2=0
cc_502 N_A_1231_367#_M1010_g N_VPWR_c_794_n 0.00931409f $X=7.02 $Y=2.465 $X2=0
+ $Y2=0
cc_503 N_A_1231_367#_c_742_n GCLK 0.0050733f $X=7.205 $Y=1.35 $X2=0 $Y2=0
cc_504 N_A_1231_367#_M1010_g N_GCLK_c_978_n 0.00646059f $X=7.02 $Y=2.465 $X2=0
+ $Y2=0
cc_505 N_A_1231_367#_c_738_n N_GCLK_c_978_n 0.0140065f $X=7.205 $Y=1.185 $X2=0
+ $Y2=0
cc_506 N_A_1231_367#_c_740_n N_GCLK_c_978_n 0.0143382f $X=6.885 $Y=1.91 $X2=0
+ $Y2=0
cc_507 N_A_1231_367#_c_741_n N_GCLK_c_978_n 0.0337815f $X=6.885 $Y=1.335 $X2=0
+ $Y2=0
cc_508 N_A_1231_367#_c_741_n N_VGND_M1005_s 0.002326f $X=6.885 $Y=1.335 $X2=0
+ $Y2=0
cc_509 N_A_1231_367#_c_738_n N_VGND_c_995_n 0.0129663f $X=7.205 $Y=1.185 $X2=0
+ $Y2=0
cc_510 N_A_1231_367#_c_739_n N_VGND_c_995_n 0.0386836f $X=6.47 $Y=0.47 $X2=0
+ $Y2=0
cc_511 N_A_1231_367#_c_741_n N_VGND_c_995_n 0.0199639f $X=6.885 $Y=1.335 $X2=0
+ $Y2=0
cc_512 N_A_1231_367#_c_742_n N_VGND_c_995_n 0.00121852f $X=7.205 $Y=1.35 $X2=0
+ $Y2=0
cc_513 N_A_1231_367#_c_739_n N_VGND_c_1003_n 0.0137476f $X=6.47 $Y=0.47 $X2=0
+ $Y2=0
cc_514 N_A_1231_367#_c_738_n N_VGND_c_1004_n 0.00486043f $X=7.205 $Y=1.185 $X2=0
+ $Y2=0
cc_515 N_A_1231_367#_c_738_n N_VGND_c_1005_n 0.00917987f $X=7.205 $Y=1.185 $X2=0
+ $Y2=0
cc_516 N_A_1231_367#_c_739_n N_VGND_c_1005_n 0.0101575f $X=6.47 $Y=0.47 $X2=0
+ $Y2=0
cc_517 N_VPWR_c_796_n N_A_154_69#_c_884_n 0.00847177f $X=0.26 $Y=2.785 $X2=0
+ $Y2=0
cc_518 N_VPWR_c_797_n N_A_154_69#_c_884_n 0.0477901f $X=1.63 $Y=2.435 $X2=0
+ $Y2=0
cc_519 N_VPWR_c_807_n N_A_154_69#_c_884_n 0.0229256f $X=1.455 $Y=3.33 $X2=0
+ $Y2=0
cc_520 N_VPWR_c_794_n N_A_154_69#_c_884_n 0.0179682f $X=7.44 $Y=3.33 $X2=0 $Y2=0
cc_521 N_VPWR_M1004_s N_A_154_69#_c_885_n 0.00881446f $X=1.495 $Y=2.045 $X2=0
+ $Y2=0
cc_522 N_VPWR_c_797_n N_A_154_69#_c_885_n 0.0211114f $X=1.63 $Y=2.435 $X2=0
+ $Y2=0
cc_523 N_VPWR_M1004_s N_A_154_69#_c_886_n 0.0066212f $X=1.495 $Y=2.045 $X2=0
+ $Y2=0
cc_524 N_VPWR_c_797_n N_A_154_69#_c_886_n 0.0458779f $X=1.63 $Y=2.435 $X2=0
+ $Y2=0
cc_525 N_VPWR_c_801_n N_A_154_69#_c_887_n 0.0575051f $X=4.135 $Y=3.33 $X2=0
+ $Y2=0
cc_526 N_VPWR_c_794_n N_A_154_69#_c_887_n 0.0342937f $X=7.44 $Y=3.33 $X2=0 $Y2=0
cc_527 N_VPWR_c_797_n N_A_154_69#_c_888_n 0.0147864f $X=1.63 $Y=2.435 $X2=0
+ $Y2=0
cc_528 N_VPWR_c_801_n N_A_154_69#_c_888_n 0.0102342f $X=4.135 $Y=3.33 $X2=0
+ $Y2=0
cc_529 N_VPWR_c_794_n N_A_154_69#_c_888_n 0.00583289f $X=7.44 $Y=3.33 $X2=0
+ $Y2=0
cc_530 N_VPWR_c_794_n N_GCLK_M1010_d 0.0040649f $X=7.44 $Y=3.33 $X2=0 $Y2=0
cc_531 N_VPWR_c_808_n GCLK 0.0314352f $X=7.44 $Y=3.33 $X2=0 $Y2=0
cc_532 N_VPWR_c_794_n GCLK 0.0172175f $X=7.44 $Y=3.33 $X2=0 $Y2=0
cc_533 N_A_154_69#_c_897_n N_VGND_c_992_n 0.0213953f $X=0.91 $Y=0.555 $X2=0
+ $Y2=0
cc_534 N_A_154_69#_c_897_n N_VGND_c_998_n 0.010891f $X=0.91 $Y=0.555 $X2=0 $Y2=0
cc_535 N_A_154_69#_c_897_n N_VGND_c_1005_n 0.0123102f $X=0.91 $Y=0.555 $X2=0
+ $Y2=0
cc_536 N_GCLK_c_978_n N_VGND_c_1004_n 0.018528f $X=7.42 $Y=0.42 $X2=0 $Y2=0
cc_537 N_GCLK_M1005_d N_VGND_c_1005_n 0.00371702f $X=7.28 $Y=0.235 $X2=0 $Y2=0
cc_538 N_GCLK_c_978_n N_VGND_c_1005_n 0.0104192f $X=7.42 $Y=0.42 $X2=0 $Y2=0
