* File: sky130_fd_sc_lp__sdfxtp_lp.pex.spice
* Created: Fri Aug 28 11:31:09 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__SDFXTP_LP%A_27_409# 1 2 9 13 15 16 17 20 24 28 32 34
+ 35
c66 35 0 1.50941e-19 $X=1.59 $Y=1.33
c67 9 0 4.91194e-20 $X=1.63 $Y=2.585
r68 34 35 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.59
+ $Y=1.33 $X2=1.59 $Y2=1.33
r69 29 32 4.56719 $w=1.7e-07 $l=2.78e-07 $layer=LI1_cond $X=0.67 $Y=1.25
+ $X2=0.392 $Y2=1.25
r70 28 34 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.425 $Y=1.25
+ $X2=1.59 $Y2=1.25
r71 28 29 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=1.425 $Y=1.25
+ $X2=0.67 $Y2=1.25
r72 24 26 32.7294 $w=2.48e-07 $l=7.1e-07 $layer=LI1_cond $X=0.24 $Y=2.19
+ $X2=0.24 $Y2=2.9
r73 22 32 2.40447 $w=4.02e-07 $l=1.898e-07 $layer=LI1_cond $X=0.24 $Y=1.335
+ $X2=0.392 $Y2=1.25
r74 22 24 39.4136 $w=2.48e-07 $l=8.55e-07 $layer=LI1_cond $X=0.24 $Y=1.335
+ $X2=0.24 $Y2=2.19
r75 18 32 2.40447 $w=4.02e-07 $l=8.5e-08 $layer=LI1_cond $X=0.392 $Y=1.165
+ $X2=0.392 $Y2=1.25
r76 18 20 7.11182 $w=5.53e-07 $l=3.3e-07 $layer=LI1_cond $X=0.392 $Y=1.165
+ $X2=0.392 $Y2=0.835
r77 16 35 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.59 $Y=1.67
+ $X2=1.59 $Y2=1.33
r78 16 17 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.59 $Y=1.67
+ $X2=1.59 $Y2=1.835
r79 15 35 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.59 $Y=1.165
+ $X2=1.59 $Y2=1.33
r80 13 15 106.04 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=1.68 $Y=0.835
+ $X2=1.68 $Y2=1.165
r81 9 17 186.34 $w=2.5e-07 $l=7.5e-07 $layer=POLY_cond $X=1.63 $Y=2.585 $X2=1.63
+ $Y2=1.835
r82 2 26 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.045 $X2=0.28 $Y2=2.9
r83 2 24 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.045 $X2=0.28 $Y2=2.19
r84 1 20 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.36
+ $Y=0.625 $X2=0.505 $Y2=0.835
.ends

.subckt PM_SKY130_FD_SC_LP__SDFXTP_LP%D 3 7 11 12 13 16 17
c40 17 0 1.50941e-19 $X=2.13 $Y=1.38
r41 16 17 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.13
+ $Y=1.38 $X2=2.13 $Y2=1.38
r42 13 17 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=2.13 $Y=1.665
+ $X2=2.13 $Y2=1.38
r43 11 16 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.13 $Y=1.72
+ $X2=2.13 $Y2=1.38
r44 11 12 31.6748 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.13 $Y=1.72
+ $X2=2.13 $Y2=1.885
r45 10 16 41.8716 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.13 $Y=1.215
+ $X2=2.13 $Y2=1.38
r46 7 12 173.918 $w=2.5e-07 $l=7e-07 $layer=POLY_cond $X=2.16 $Y=2.585 $X2=2.16
+ $Y2=1.885
r47 3 10 194.851 $w=1.5e-07 $l=3.8e-07 $layer=POLY_cond $X=2.07 $Y=0.835
+ $X2=2.07 $Y2=1.215
.ends

.subckt PM_SKY130_FD_SC_LP__SDFXTP_LP%SCE 3 7 9 14 15 16 20 21 23 26 34
c79 26 0 4.91194e-20 $X=0.72 $Y=1.665
r80 33 34 44.4629 $w=3.3e-07 $l=1.55e-07 $layer=POLY_cond $X=0.72 $Y=1.68
+ $X2=0.875 $Y2=1.68
r81 31 33 1.74861 $w=3.3e-07 $l=1e-08 $layer=POLY_cond $X=0.71 $Y=1.68 $X2=0.72
+ $Y2=1.68
r82 28 31 28.8521 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.545 $Y=1.68
+ $X2=0.71 $Y2=1.68
r83 26 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.71
+ $Y=1.68 $X2=0.71 $Y2=1.68
r84 21 25 40.9178 $w=2.5e-07 $l=1.25e-07 $layer=POLY_cond $X=2.63 $Y=1.245
+ $X2=2.63 $Y2=1.12
r85 21 23 332.928 $w=2.5e-07 $l=1.34e-06 $layer=POLY_cond $X=2.63 $Y=1.245
+ $X2=2.63 $Y2=2.585
r86 20 25 146.138 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.58 $Y=0.835
+ $X2=2.58 $Y2=1.12
r87 17 20 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=2.58 $Y=0.255
+ $X2=2.58 $Y2=0.835
r88 15 17 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.505 $Y=0.18
+ $X2=2.58 $Y2=0.255
r89 15 16 676.851 $w=1.5e-07 $l=1.32e-06 $layer=POLY_cond $X=2.505 $Y=0.18
+ $X2=1.185 $Y2=0.18
r90 12 14 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=1.11 $Y=1.515
+ $X2=1.11 $Y2=0.835
r91 11 16 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.11 $Y=0.255
+ $X2=1.185 $Y2=0.18
r92 11 14 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=1.11 $Y=0.255
+ $X2=1.11 $Y2=0.835
r93 9 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.035 $Y=1.59
+ $X2=1.11 $Y2=1.515
r94 9 34 82.0426 $w=1.5e-07 $l=1.6e-07 $layer=POLY_cond $X=1.035 $Y=1.59
+ $X2=0.875 $Y2=1.59
r95 5 33 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.72 $Y=1.515
+ $X2=0.72 $Y2=1.68
r96 5 7 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=0.72 $Y=1.515 $X2=0.72
+ $Y2=0.835
r97 1 28 9.34494 $w=2.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.545 $Y=1.845
+ $X2=0.545 $Y2=1.68
r98 1 3 173.918 $w=2.5e-07 $l=7e-07 $layer=POLY_cond $X=0.545 $Y=1.845 $X2=0.545
+ $Y2=2.545
.ends

.subckt PM_SKY130_FD_SC_LP__SDFXTP_LP%SCD 3 6 9 11 12 13 17
r41 17 19 46.7569 $w=3.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.15 $Y=1.41
+ $X2=3.15 $Y2=1.245
r42 17 18 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.17
+ $Y=1.41 $X2=3.17 $Y2=1.41
r43 13 18 7.67632 $w=6.68e-07 $l=4.3e-07 $layer=LI1_cond $X=3.6 $Y=1.58 $X2=3.17
+ $Y2=1.58
r44 12 18 0.892596 $w=6.68e-07 $l=5e-08 $layer=LI1_cond $X=3.12 $Y=1.58 $X2=3.17
+ $Y2=1.58
r45 9 11 166.464 $w=2.5e-07 $l=6.7e-07 $layer=POLY_cond $X=3.16 $Y=2.585
+ $X2=3.16 $Y2=1.915
r46 6 11 32.1785 $w=3.7e-07 $l=1.85e-07 $layer=POLY_cond $X=3.15 $Y=1.73
+ $X2=3.15 $Y2=1.915
r47 5 17 3.11915 $w=3.7e-07 $l=2e-08 $layer=POLY_cond $X=3.15 $Y=1.43 $X2=3.15
+ $Y2=1.41
r48 5 6 46.7872 $w=3.7e-07 $l=3e-07 $layer=POLY_cond $X=3.15 $Y=1.43 $X2=3.15
+ $Y2=1.73
r49 3 19 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=3.04 $Y=0.835
+ $X2=3.04 $Y2=1.245
.ends

.subckt PM_SKY130_FD_SC_LP__SDFXTP_LP%CLK 3 7 11 13 21
c42 7 0 1.93089e-19 $X=4.335 $Y=2.235
r43 20 21 8.74306 $w=3.3e-07 $l=5e-08 $layer=POLY_cond $X=4.335 $Y=1.345
+ $X2=4.385 $Y2=1.345
r44 18 20 38.4695 $w=3.3e-07 $l=2.2e-07 $layer=POLY_cond $X=4.115 $Y=1.345
+ $X2=4.335 $Y2=1.345
r45 15 18 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=4.025 $Y=1.345
+ $X2=4.115 $Y2=1.345
r46 13 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.115
+ $Y=1.345 $X2=4.115 $Y2=1.345
r47 9 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.385 $Y=1.18
+ $X2=4.385 $Y2=1.345
r48 9 11 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=4.385 $Y=1.18
+ $X2=4.385 $Y2=0.54
r49 5 20 9.34494 $w=2.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.335 $Y=1.51
+ $X2=4.335 $Y2=1.345
r50 5 7 180.129 $w=2.5e-07 $l=7.25e-07 $layer=POLY_cond $X=4.335 $Y=1.51
+ $X2=4.335 $Y2=2.235
r51 1 15 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.025 $Y=1.18
+ $X2=4.025 $Y2=1.345
r52 1 3 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=4.025 $Y=1.18 $X2=4.025
+ $Y2=0.54
.ends

.subckt PM_SKY130_FD_SC_LP__SDFXTP_LP%A_1576_99# 1 2 3 12 15 17 22 27 29 31 33
+ 35 38 39 40 42
c96 38 0 1.11746e-19 $X=8.045 $Y=1.32
r97 38 43 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.045 $Y=1.32
+ $X2=8.045 $Y2=1.485
r98 38 42 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.045 $Y=1.32
+ $X2=8.045 $Y2=1.155
r99 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.045
+ $Y=1.32 $X2=8.045 $Y2=1.32
r100 35 37 16.0154 $w=2.59e-07 $l=3.4e-07 $layer=LI1_cond $X=8.045 $Y=0.98
+ $X2=8.045 $Y2=1.32
r101 31 33 81.2246 $w=1.68e-07 $l=1.245e-06 $layer=LI1_cond $X=9.275 $Y=0.35
+ $X2=10.52 $Y2=0.35
r102 27 40 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=9.27 $Y=1.88
+ $X2=9.27 $Y2=1.715
r103 27 29 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=9.27 $Y=1.88
+ $X2=9.27 $Y2=2.59
r104 23 39 3.70735 $w=2.5e-07 $l=1.18427e-07 $layer=LI1_cond $X=9.19 $Y=1.065
+ $X2=9.11 $Y2=0.98
r105 23 40 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=9.19 $Y=1.065
+ $X2=9.19 $Y2=1.715
r106 20 39 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=9.11 $Y=0.895
+ $X2=9.11 $Y2=0.98
r107 20 22 2.09535 $w=3.28e-07 $l=6e-08 $layer=LI1_cond $X=9.11 $Y=0.895
+ $X2=9.11 $Y2=0.835
r108 19 31 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=9.11 $Y=0.435
+ $X2=9.275 $Y2=0.35
r109 19 22 13.969 $w=3.28e-07 $l=4e-07 $layer=LI1_cond $X=9.11 $Y=0.435 $X2=9.11
+ $Y2=0.835
r110 18 35 3.20129 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.21 $Y=0.98
+ $X2=8.045 $Y2=0.98
r111 17 39 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.945 $Y=0.98
+ $X2=9.11 $Y2=0.98
r112 17 18 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=8.945 $Y=0.98
+ $X2=8.21 $Y2=0.98
r113 15 43 186.34 $w=2.5e-07 $l=7.5e-07 $layer=POLY_cond $X=8.005 $Y=2.235
+ $X2=8.005 $Y2=1.485
r114 12 42 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=7.955 $Y=0.835
+ $X2=7.955 $Y2=1.155
r115 3 29 400 $w=1.7e-07 $l=9.42974e-07 $layer=licon1_PDIFF $count=1 $X=9.085
+ $Y=1.735 $X2=9.27 $Y2=2.59
r116 3 27 400 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_PDIFF $count=1 $X=9.085
+ $Y=1.735 $X2=9.27 $Y2=1.88
r117 2 33 182 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=1 $X=10.375
+ $Y=0.205 $X2=10.52 $Y2=0.35
r118 1 22 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=8.97
+ $Y=0.625 $X2=9.11 $Y2=0.835
.ends

.subckt PM_SKY130_FD_SC_LP__SDFXTP_LP%A_1263_155# 1 2 9 13 17 21 23 24 27 31 35
+ 38 45
c84 38 0 1.11746e-19 $X=7.25 $Y=1.45
c85 31 0 4.17108e-20 $X=8.46 $Y=1.75
r86 44 45 11.366 $w=3.3e-07 $l=6.5e-08 $layer=POLY_cond $X=8.895 $Y=1.41
+ $X2=8.96 $Y2=1.41
r87 38 40 10.4768 $w=3.28e-07 $l=3e-07 $layer=LI1_cond $X=7.25 $Y=1.45 $X2=7.25
+ $Y2=1.75
r88 36 44 47.2125 $w=3.3e-07 $l=2.7e-07 $layer=POLY_cond $X=8.625 $Y=1.41
+ $X2=8.895 $Y2=1.41
r89 36 41 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=8.625 $Y=1.41
+ $X2=8.535 $Y2=1.41
r90 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.625
+ $Y=1.41 $X2=8.625 $Y2=1.41
r91 33 35 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=8.625 $Y=1.665
+ $X2=8.625 $Y2=1.41
r92 32 40 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.415 $Y=1.75
+ $X2=7.25 $Y2=1.75
r93 31 33 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=8.46 $Y=1.75
+ $X2=8.625 $Y2=1.665
r94 31 32 68.1765 $w=1.68e-07 $l=1.045e-06 $layer=LI1_cond $X=8.46 $Y=1.75
+ $X2=7.415 $Y2=1.75
r95 27 29 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=7.25 $Y=1.88 $X2=7.25
+ $Y2=2.59
r96 25 40 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=7.25 $Y=1.835
+ $X2=7.25 $Y2=1.75
r97 25 27 1.57151 $w=3.28e-07 $l=4.5e-08 $layer=LI1_cond $X=7.25 $Y=1.835
+ $X2=7.25 $Y2=1.88
r98 23 38 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.085 $Y=1.45
+ $X2=7.25 $Y2=1.45
r99 23 24 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=7.085 $Y=1.45
+ $X2=6.89 $Y2=1.45
r100 19 24 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.725 $Y=1.365
+ $X2=6.89 $Y2=1.45
r101 19 21 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=6.725 $Y=1.365
+ $X2=6.725 $Y2=1.05
r102 15 45 9.34494 $w=2.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.96 $Y=1.575
+ $X2=8.96 $Y2=1.41
r103 15 17 163.979 $w=2.5e-07 $l=6.6e-07 $layer=POLY_cond $X=8.96 $Y=1.575
+ $X2=8.96 $Y2=2.235
r104 11 44 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.895 $Y=1.245
+ $X2=8.895 $Y2=1.41
r105 11 13 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=8.895 $Y=1.245
+ $X2=8.895 $Y2=0.835
r106 7 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.535 $Y=1.245
+ $X2=8.535 $Y2=1.41
r107 7 9 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=8.535 $Y=1.245
+ $X2=8.535 $Y2=0.835
r108 2 29 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=7.11
+ $Y=1.735 $X2=7.25 $Y2=2.59
r109 2 27 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=7.11
+ $Y=1.735 $X2=7.25 $Y2=1.88
r110 1 21 182 $w=1.7e-07 $l=5.29953e-07 $layer=licon1_NDIFF $count=1 $X=6.315
+ $Y=0.775 $X2=6.725 $Y2=1.05
.ends

.subckt PM_SKY130_FD_SC_LP__SDFXTP_LP%A_733_66# 1 2 7 9 12 17 18 19 22 24 30 32
+ 35 38 40 42 47 50 51 52 53 54 58 62 64 68 69 71 76
c166 68 0 1.92223e-19 $X=4.46 $Y=0.915
c167 30 0 2.74949e-19 $X=7.515 $Y=2.235
c168 22 0 1.51839e-20 $X=6.94 $Y=0.985
r169 75 77 17.01 $w=5.83e-07 $l=5.05e-07 $layer=LI1_cond $X=4.752 $Y=1.025
+ $X2=4.752 $Y2=1.53
r170 75 76 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.88
+ $Y=1.025 $X2=4.88 $Y2=1.025
r171 71 77 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=4.545 $Y=1.715
+ $X2=4.545 $Y2=1.53
r172 68 75 2.24904 $w=5.83e-07 $l=1.1e-07 $layer=LI1_cond $X=4.752 $Y=0.915
+ $X2=4.752 $Y2=1.025
r173 68 69 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=4.46 $Y=0.915
+ $X2=3.975 $Y2=0.915
r174 64 71 7.21222 $w=2.6e-07 $l=1.67183e-07 $layer=LI1_cond $X=4.46 $Y=1.845
+ $X2=4.545 $Y2=1.715
r175 64 66 17.2866 $w=2.58e-07 $l=3.9e-07 $layer=LI1_cond $X=4.46 $Y=1.845
+ $X2=4.07 $Y2=1.845
r176 60 69 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.81 $Y=0.83
+ $X2=3.975 $Y2=0.915
r177 60 62 10.1275 $w=3.28e-07 $l=2.9e-07 $layer=LI1_cond $X=3.81 $Y=0.83
+ $X2=3.81 $Y2=0.54
r178 53 54 47.1291 $w=2.5e-07 $l=1.5e-07 $layer=POLY_cond $X=7.505 $Y=1.12
+ $X2=7.505 $Y2=1.27
r179 49 76 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=4.88 $Y=1.365
+ $X2=4.88 $Y2=1.025
r180 49 50 31.0234 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.88 $Y=1.365
+ $X2=4.88 $Y2=1.53
r181 46 76 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=4.88 $Y=1.01
+ $X2=4.88 $Y2=1.025
r182 46 47 151.266 $w=1.5e-07 $l=2.95e-07 $layer=POLY_cond $X=4.88 $Y=0.935
+ $X2=5.175 $Y2=0.935
r183 43 46 33.3298 $w=1.5e-07 $l=6.5e-08 $layer=POLY_cond $X=4.815 $Y=0.935
+ $X2=4.88 $Y2=0.935
r184 40 58 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.89 $Y=1.27
+ $X2=9.89 $Y2=1.345
r185 40 42 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=9.89 $Y=1.27
+ $X2=9.89 $Y2=0.985
r186 36 58 117.936 $w=1.5e-07 $l=2.3e-07 $layer=POLY_cond $X=9.66 $Y=1.345
+ $X2=9.89 $Y2=1.345
r187 36 55 133.319 $w=1.5e-07 $l=2.6e-07 $layer=POLY_cond $X=9.66 $Y=1.345
+ $X2=9.4 $Y2=1.345
r188 36 38 202.49 $w=2.5e-07 $l=8.15e-07 $layer=POLY_cond $X=9.66 $Y=1.42
+ $X2=9.66 $Y2=2.235
r189 35 55 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.4 $Y=1.27 $X2=9.4
+ $Y2=1.345
r190 34 35 520.457 $w=1.5e-07 $l=1.015e-06 $layer=POLY_cond $X=9.4 $Y=0.255
+ $X2=9.4 $Y2=1.27
r191 33 52 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.52 $Y=0.18
+ $X2=7.445 $Y2=0.18
r192 32 34 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.325 $Y=0.18
+ $X2=9.4 $Y2=0.255
r193 32 33 925.543 $w=1.5e-07 $l=1.805e-06 $layer=POLY_cond $X=9.325 $Y=0.18
+ $X2=7.52 $Y2=0.18
r194 30 54 239.758 $w=2.5e-07 $l=9.65e-07 $layer=POLY_cond $X=7.515 $Y=2.235
+ $X2=7.515 $Y2=1.27
r195 26 52 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.445 $Y=0.255
+ $X2=7.445 $Y2=0.18
r196 26 53 443.543 $w=1.5e-07 $l=8.65e-07 $layer=POLY_cond $X=7.445 $Y=0.255
+ $X2=7.445 $Y2=1.12
r197 25 51 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.015 $Y=0.18
+ $X2=6.94 $Y2=0.18
r198 24 52 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.37 $Y=0.18
+ $X2=7.445 $Y2=0.18
r199 24 25 182.032 $w=1.5e-07 $l=3.55e-07 $layer=POLY_cond $X=7.37 $Y=0.18
+ $X2=7.015 $Y2=0.18
r200 20 51 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.94 $Y=0.255
+ $X2=6.94 $Y2=0.18
r201 20 22 374.319 $w=1.5e-07 $l=7.3e-07 $layer=POLY_cond $X=6.94 $Y=0.255
+ $X2=6.94 $Y2=0.985
r202 18 51 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.865 $Y=0.18
+ $X2=6.94 $Y2=0.18
r203 18 19 828.117 $w=1.5e-07 $l=1.615e-06 $layer=POLY_cond $X=6.865 $Y=0.18
+ $X2=5.25 $Y2=0.18
r204 15 47 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.175 $Y=0.86
+ $X2=5.175 $Y2=0.935
r205 15 17 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=5.175 $Y=0.86
+ $X2=5.175 $Y2=0.54
r206 14 19 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.175 $Y=0.255
+ $X2=5.25 $Y2=0.18
r207 14 17 146.138 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=5.175 $Y=0.255
+ $X2=5.175 $Y2=0.54
r208 12 50 175.16 $w=2.5e-07 $l=7.05e-07 $layer=POLY_cond $X=4.865 $Y=2.235
+ $X2=4.865 $Y2=1.53
r209 7 43 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.815 $Y=0.86
+ $X2=4.815 $Y2=0.935
r210 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=4.815 $Y=0.86
+ $X2=4.815 $Y2=0.54
r211 2 66 600 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=3.925
+ $Y=1.735 $X2=4.07 $Y2=1.885
r212 1 62 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=3.665
+ $Y=0.33 $X2=3.81 $Y2=0.54
.ends

.subckt PM_SKY130_FD_SC_LP__SDFXTP_LP%A_998_347# 1 2 8 9 10 11 12 13 15 18 20 25
+ 26 28 32 33 36 40 43
c103 40 0 1.93089e-19 $X=5.39 $Y=1.64
c104 18 0 2.1035e-19 $X=6.985 $Y=2.235
c105 10 0 1.92223e-19 $X=5.82 $Y=1.38
r106 42 43 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.655
+ $Y=1.47 $X2=5.655 $Y2=1.47
r107 40 42 5.93211 $w=5.45e-07 $l=2.65e-07 $layer=LI1_cond $X=5.39 $Y=1.64
+ $X2=5.655 $Y2=1.64
r108 39 40 5.82018 $w=5.45e-07 $l=3.62353e-07 $layer=LI1_cond $X=5.13 $Y=1.885
+ $X2=5.39 $Y2=1.64
r109 34 40 3.67229 $w=3.3e-07 $l=3.35e-07 $layer=LI1_cond $X=5.39 $Y=1.305
+ $X2=5.39 $Y2=1.64
r110 34 36 26.7157 $w=3.28e-07 $l=7.65e-07 $layer=LI1_cond $X=5.39 $Y=1.305
+ $X2=5.39 $Y2=0.54
r111 31 43 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=5.655 $Y=1.81
+ $X2=5.655 $Y2=1.47
r112 31 32 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.655 $Y=1.81
+ $X2=5.655 $Y2=1.975
r113 30 43 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=5.655 $Y=1.455
+ $X2=5.655 $Y2=1.47
r114 26 28 340.989 $w=1.5e-07 $l=6.65e-07 $layer=POLY_cond $X=10.32 $Y=1.65
+ $X2=10.32 $Y2=0.985
r115 23 25 191.309 $w=2.5e-07 $l=7.7e-07 $layer=POLY_cond $X=10.35 $Y=3.075
+ $X2=10.35 $Y2=2.305
r116 22 26 29.3902 $w=2.46e-07 $l=1.64317e-07 $layer=POLY_cond $X=10.35 $Y=1.8
+ $X2=10.32 $Y2=1.65
r117 22 25 125.469 $w=2.5e-07 $l=5.05e-07 $layer=POLY_cond $X=10.35 $Y=1.8
+ $X2=10.35 $Y2=2.305
r118 21 33 30.4925 $w=1.5e-07 $l=1.25e-07 $layer=POLY_cond $X=7.11 $Y=3.15
+ $X2=6.985 $Y2=3.15
r119 20 23 29.1797 $w=1.5e-07 $l=1.58114e-07 $layer=POLY_cond $X=10.225 $Y=3.15
+ $X2=10.35 $Y2=3.075
r120 20 21 1597.27 $w=1.5e-07 $l=3.115e-06 $layer=POLY_cond $X=10.225 $Y=3.15
+ $X2=7.11 $Y2=3.15
r121 16 33 1.63566 $w=2.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.985 $Y=3.075
+ $X2=6.985 $Y2=3.15
r122 16 18 208.701 $w=2.5e-07 $l=8.4e-07 $layer=POLY_cond $X=6.985 $Y=3.075
+ $X2=6.985 $Y2=2.235
r123 13 15 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=6.24 $Y=1.305
+ $X2=6.24 $Y2=0.985
r124 11 33 30.4925 $w=1.5e-07 $l=1.25e-07 $layer=POLY_cond $X=6.86 $Y=3.15
+ $X2=6.985 $Y2=3.15
r125 11 12 533.277 $w=1.5e-07 $l=1.04e-06 $layer=POLY_cond $X=6.86 $Y=3.15
+ $X2=5.82 $Y2=3.15
r126 10 30 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=5.82 $Y=1.38
+ $X2=5.655 $Y2=1.455
r127 9 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.165 $Y=1.38
+ $X2=6.24 $Y2=1.305
r128 9 10 176.904 $w=1.5e-07 $l=3.45e-07 $layer=POLY_cond $X=6.165 $Y=1.38
+ $X2=5.82 $Y2=1.38
r129 8 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.745 $Y=3.075
+ $X2=5.82 $Y2=3.15
r130 8 32 564.043 $w=1.5e-07 $l=1.1e-06 $layer=POLY_cond $X=5.745 $Y=3.075
+ $X2=5.745 $Y2=1.975
r131 2 39 600 $w=1.7e-07 $l=2.08567e-07 $layer=licon1_PDIFF $count=1 $X=4.99
+ $Y=1.735 $X2=5.13 $Y2=1.885
r132 1 36 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=5.25
+ $Y=0.33 $X2=5.39 $Y2=0.54
.ends

.subckt PM_SKY130_FD_SC_LP__SDFXTP_LP%A_2148_185# 1 2 9 13 15 16 19 23 27 32 34
+ 41 44 48 51 52 56 57 60
c102 48 0 2.13067e-20 $X=10.94 $Y=1.13
r103 60 62 10.7321 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=12.295 $Y=0.555
+ $X2=12.295 $Y2=0.785
r104 56 57 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=12.56
+ $Y=1.13 $X2=12.56 $Y2=1.13
r105 54 56 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=12.215 $Y=1.05
+ $X2=12.56 $Y2=1.05
r106 53 54 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=11.94 $Y=1.05
+ $X2=12.215 $Y2=1.05
r107 51 52 9.25191 $w=4.53e-07 $l=1.65e-07 $layer=LI1_cond $X=11.797 $Y=1.99
+ $X2=11.797 $Y2=1.825
r108 48 65 13.0036 $w=2.78e-07 $l=7.5e-08 $layer=POLY_cond $X=10.94 $Y=1.11
+ $X2=10.865 $Y2=1.11
r109 47 48 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.94
+ $Y=1.13 $X2=10.94 $Y2=1.13
r110 44 47 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=10.94 $Y=1.05
+ $X2=10.94 $Y2=1.13
r111 41 54 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=12.215 $Y=0.965
+ $X2=12.215 $Y2=1.05
r112 41 62 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=12.215 $Y=0.965
+ $X2=12.215 $Y2=0.785
r113 38 53 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.94 $Y=1.135
+ $X2=11.94 $Y2=1.05
r114 38 52 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=11.94 $Y=1.135
+ $X2=11.94 $Y2=1.825
r115 35 44 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.105 $Y=1.05
+ $X2=10.94 $Y2=1.05
r116 34 53 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=11.855 $Y=1.05
+ $X2=11.94 $Y2=1.05
r117 34 35 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=11.855 $Y=1.05
+ $X2=11.105 $Y2=1.05
r118 29 57 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=12.56 $Y=1.115
+ $X2=12.56 $Y2=1.13
r119 25 32 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=13.425 $Y=0.965
+ $X2=13.425 $Y2=1.04
r120 25 27 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=13.425 $Y=0.965
+ $X2=13.425 $Y2=0.555
r121 21 32 25.6383 $w=1.5e-07 $l=5e-08 $layer=POLY_cond $X=13.375 $Y=1.04
+ $X2=13.425 $Y2=1.04
r122 21 30 158.957 $w=1.5e-07 $l=3.1e-07 $layer=POLY_cond $X=13.375 $Y=1.04
+ $X2=13.065 $Y2=1.04
r123 21 23 329.201 $w=2.5e-07 $l=1.325e-06 $layer=POLY_cond $X=13.375 $Y=1.115
+ $X2=13.375 $Y2=2.44
r124 17 30 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=13.065 $Y=0.965
+ $X2=13.065 $Y2=1.04
r125 17 19 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=13.065 $Y=0.965
+ $X2=13.065 $Y2=0.555
r126 16 29 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=12.725 $Y=1.04
+ $X2=12.56 $Y2=1.115
r127 15 30 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=12.99 $Y=1.04
+ $X2=13.065 $Y2=1.04
r128 15 16 135.883 $w=1.5e-07 $l=2.65e-07 $layer=POLY_cond $X=12.99 $Y=1.04
+ $X2=12.725 $Y2=1.04
r129 11 48 60.6835 $w=2.78e-07 $l=4.32724e-07 $layer=POLY_cond $X=11.29 $Y=0.925
+ $X2=10.94 $Y2=1.11
r130 11 13 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=11.29 $Y=0.925
+ $X2=11.29 $Y2=0.555
r131 7 65 5.35669 $w=2.5e-07 $l=1.85e-07 $layer=POLY_cond $X=10.865 $Y=1.295
+ $X2=10.865 $Y2=1.11
r132 7 9 250.938 $w=2.5e-07 $l=1.01e-06 $layer=POLY_cond $X=10.865 $Y=1.295
+ $X2=10.865 $Y2=2.305
r133 2 51 300 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_PDIFF $count=2 $X=11.595
+ $Y=1.805 $X2=11.735 $Y2=1.99
r134 1 60 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=12.155
+ $Y=0.345 $X2=12.295 $Y2=0.555
.ends

.subckt PM_SKY130_FD_SC_LP__SDFXTP_LP%A_1957_347# 1 2 7 9 13 15 19 23 31 33 35
+ 37
c82 37 0 2.13067e-20 $X=11.51 $Y=1.48
r83 37 40 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=11.51 $Y=1.48 $X2=11.51
+ $Y2=1.56
r84 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.51
+ $Y=1.48 $X2=11.51 $Y2=1.48
r85 34 35 3.80956 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=10.27 $Y=1.56
+ $X2=10.055 $Y2=1.56
r86 33 40 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.345 $Y=1.56
+ $X2=11.51 $Y2=1.56
r87 33 34 70.1337 $w=1.68e-07 $l=1.075e-06 $layer=LI1_cond $X=11.345 $Y=1.56
+ $X2=10.27 $Y2=1.56
r88 29 35 2.88756 $w=3.3e-07 $l=1.07121e-07 $layer=LI1_cond $X=10.105 $Y=1.475
+ $X2=10.055 $Y2=1.56
r89 29 31 14.8421 $w=3.28e-07 $l=4.25e-07 $layer=LI1_cond $X=10.105 $Y=1.475
+ $X2=10.105 $Y2=1.05
r90 25 27 13.6198 $w=3.28e-07 $l=3.9e-07 $layer=LI1_cond $X=10.005 $Y=2.27
+ $X2=10.005 $Y2=2.66
r91 23 25 13.6198 $w=3.28e-07 $l=3.9e-07 $layer=LI1_cond $X=10.005 $Y=1.88
+ $X2=10.005 $Y2=2.27
r92 21 35 2.88756 $w=3.3e-07 $l=1.07121e-07 $layer=LI1_cond $X=10.005 $Y=1.645
+ $X2=10.055 $Y2=1.56
r93 21 23 8.20679 $w=3.28e-07 $l=2.35e-07 $layer=LI1_cond $X=10.005 $Y=1.645
+ $X2=10.005 $Y2=1.88
r94 17 19 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=12.08 $Y=1.165
+ $X2=12.08 $Y2=0.555
r95 16 38 32.4944 $w=3.56e-07 $l=3.34066e-07 $layer=POLY_cond $X=11.795 $Y=1.24
+ $X2=11.57 $Y2=1.48
r96 15 17 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=12.005 $Y=1.24
+ $X2=12.08 $Y2=1.165
r97 15 16 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=12.005 $Y=1.24
+ $X2=11.795 $Y2=1.24
r98 11 16 26.6719 $w=3.56e-07 $l=1.06066e-07 $layer=POLY_cond $X=11.72 $Y=1.165
+ $X2=11.795 $Y2=1.24
r99 11 13 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=11.72 $Y=1.165
+ $X2=11.72 $Y2=0.555
r100 7 38 26.6704 $w=3.56e-07 $l=2.09105e-07 $layer=POLY_cond $X=11.47 $Y=1.645
+ $X2=11.57 $Y2=1.48
r101 7 9 163.979 $w=2.5e-07 $l=6.6e-07 $layer=POLY_cond $X=11.47 $Y=1.645
+ $X2=11.47 $Y2=2.305
r102 2 27 600 $w=1.7e-07 $l=1.02914e-06 $layer=licon1_PDIFF $count=1 $X=9.785
+ $Y=1.735 $X2=10.005 $Y2=2.66
r103 2 25 600 $w=1.7e-07 $l=6.35551e-07 $layer=licon1_PDIFF $count=1 $X=9.785
+ $Y=1.735 $X2=10.005 $Y2=2.27
r104 2 23 600 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_PDIFF $count=1 $X=9.785
+ $Y=1.735 $X2=10.005 $Y2=1.88
r105 1 31 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=9.965
+ $Y=0.775 $X2=10.105 $Y2=1.05
.ends

.subckt PM_SKY130_FD_SC_LP__SDFXTP_LP%VPWR 1 2 3 4 5 6 23 29 33 37 41 43 45 50
+ 51 52 61 68 76 81 87 90 93 96 100
r108 99 100 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.68 $Y=3.33
+ $X2=13.68 $Y2=3.33
r109 96 97 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=11.28 $Y=3.33
+ $X2=11.28 $Y2=3.33
r110 93 94 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=8.4 $Y=3.33 $X2=8.4
+ $Y2=3.33
r111 90 91 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r112 87 88 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r113 85 100 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.2 $Y=3.33
+ $X2=13.68 $Y2=3.33
r114 85 97 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=13.2 $Y=3.33
+ $X2=11.28 $Y2=3.33
r115 84 85 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=13.2 $Y=3.33
+ $X2=13.2 $Y2=3.33
r116 82 96 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.295 $Y=3.33
+ $X2=11.13 $Y2=3.33
r117 82 84 124.283 $w=1.68e-07 $l=1.905e-06 $layer=LI1_cond $X=11.295 $Y=3.33
+ $X2=13.2 $Y2=3.33
r118 81 99 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=13.475 $Y=3.33
+ $X2=13.697 $Y2=3.33
r119 81 84 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=13.475 $Y=3.33
+ $X2=13.2 $Y2=3.33
r120 80 97 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.8 $Y=3.33
+ $X2=11.28 $Y2=3.33
r121 80 94 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=10.8 $Y=3.33
+ $X2=8.4 $Y2=3.33
r122 79 80 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=10.8 $Y=3.33
+ $X2=10.8 $Y2=3.33
r123 77 93 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.435 $Y=3.33
+ $X2=8.27 $Y2=3.33
r124 77 79 154.294 $w=1.68e-07 $l=2.365e-06 $layer=LI1_cond $X=8.435 $Y=3.33
+ $X2=10.8 $Y2=3.33
r125 76 96 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.965 $Y=3.33
+ $X2=11.13 $Y2=3.33
r126 76 79 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=10.965 $Y=3.33
+ $X2=10.8 $Y2=3.33
r127 75 94 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=8.4 $Y2=3.33
r128 74 75 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r129 72 91 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=4.56 $Y2=3.33
r130 71 74 187.893 $w=1.68e-07 $l=2.88e-06 $layer=LI1_cond $X=5.04 $Y=3.33
+ $X2=7.92 $Y2=3.33
r131 71 72 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r132 69 90 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.765 $Y=3.33
+ $X2=4.6 $Y2=3.33
r133 69 71 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=4.765 $Y=3.33
+ $X2=5.04 $Y2=3.33
r134 68 93 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.105 $Y=3.33
+ $X2=8.27 $Y2=3.33
r135 68 74 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=8.105 $Y=3.33
+ $X2=7.92 $Y2=3.33
r136 67 91 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r137 66 67 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r138 64 67 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=4.08 $Y2=3.33
r139 63 66 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=3.12 $Y=3.33
+ $X2=4.08 $Y2=3.33
r140 63 64 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r141 61 90 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.435 $Y=3.33
+ $X2=4.6 $Y2=3.33
r142 61 66 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=4.435 $Y=3.33
+ $X2=4.08 $Y2=3.33
r143 60 64 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r144 59 60 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r145 57 60 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r146 57 88 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r147 56 59 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r148 56 57 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r149 54 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.975 $Y=3.33
+ $X2=0.81 $Y2=3.33
r150 54 56 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=0.975 $Y=3.33
+ $X2=1.2 $Y2=3.33
r151 52 75 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=7.92 $Y2=3.33
r152 52 72 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=5.04 $Y2=3.33
r153 50 59 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=2.73 $Y=3.33 $X2=2.64
+ $Y2=3.33
r154 50 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.73 $Y=3.33
+ $X2=2.895 $Y2=3.33
r155 49 63 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=3.06 $Y=3.33 $X2=3.12
+ $Y2=3.33
r156 49 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.06 $Y=3.33
+ $X2=2.895 $Y2=3.33
r157 45 48 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=13.64 $Y=2.085
+ $X2=13.64 $Y2=2.795
r158 43 99 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=13.64 $Y=3.245
+ $X2=13.697 $Y2=3.33
r159 43 48 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=13.64 $Y=3.245
+ $X2=13.64 $Y2=2.795
r160 39 96 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=11.13 $Y=3.245
+ $X2=11.13 $Y2=3.33
r161 39 41 43.8278 $w=3.28e-07 $l=1.255e-06 $layer=LI1_cond $X=11.13 $Y=3.245
+ $X2=11.13 $Y2=1.99
r162 35 93 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.27 $Y=3.245
+ $X2=8.27 $Y2=3.33
r163 35 37 37.1925 $w=3.28e-07 $l=1.065e-06 $layer=LI1_cond $X=8.27 $Y=3.245
+ $X2=8.27 $Y2=2.18
r164 31 90 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.6 $Y=3.245 $X2=4.6
+ $Y2=3.33
r165 31 33 22.8742 $w=3.28e-07 $l=6.55e-07 $layer=LI1_cond $X=4.6 $Y=3.245
+ $X2=4.6 $Y2=2.59
r166 27 51 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.895 $Y=3.245
+ $X2=2.895 $Y2=3.33
r167 27 29 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=2.895 $Y=3.245
+ $X2=2.895 $Y2=2.94
r168 23 26 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=0.81 $Y=2.19
+ $X2=0.81 $Y2=2.9
r169 21 87 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.81 $Y=3.245
+ $X2=0.81 $Y2=3.33
r170 21 26 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=0.81 $Y=3.245
+ $X2=0.81 $Y2=2.9
r171 6 48 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=13.5
+ $Y=1.94 $X2=13.64 $Y2=2.795
r172 6 45 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=13.5
+ $Y=1.94 $X2=13.64 $Y2=2.085
r173 5 41 300 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_PDIFF $count=2 $X=10.99
+ $Y=1.805 $X2=11.13 $Y2=1.99
r174 4 37 300 $w=1.7e-07 $l=5.10221e-07 $layer=licon1_PDIFF $count=2 $X=8.13
+ $Y=1.735 $X2=8.27 $Y2=2.18
r175 3 33 600 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=4.46
+ $Y=1.735 $X2=4.6 $Y2=2.59
r176 2 29 600 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=2.755
+ $Y=2.085 $X2=2.895 $Y2=2.94
r177 1 26 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=0.67
+ $Y=2.045 $X2=0.81 $Y2=2.9
r178 1 23 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.67
+ $Y=2.045 $X2=0.81 $Y2=2.19
.ends

.subckt PM_SKY130_FD_SC_LP__SDFXTP_LP%A_244_417# 1 2 9 13 17 19
r41 15 17 3.84148 $w=3.28e-07 $l=1.1e-07 $layer=LI1_cond $X=3.425 $Y=2.675
+ $X2=3.425 $Y2=2.785
r42 14 19 3.80956 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.53 $Y=2.59
+ $X2=1.365 $Y2=2.59
r43 13 15 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.26 $Y=2.59
+ $X2=3.425 $Y2=2.675
r44 13 14 112.866 $w=1.68e-07 $l=1.73e-06 $layer=LI1_cond $X=3.26 $Y=2.59
+ $X2=1.53 $Y2=2.59
r45 7 19 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.365 $Y=2.505
+ $X2=1.365 $Y2=2.59
r46 7 9 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=1.365 $Y=2.505
+ $X2=1.365 $Y2=2.23
r47 2 17 600 $w=1.7e-07 $l=7.66812e-07 $layer=licon1_PDIFF $count=1 $X=3.285
+ $Y=2.085 $X2=3.425 $Y2=2.785
r48 1 9 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=1.22
+ $Y=2.085 $X2=1.365 $Y2=2.23
.ends

.subckt PM_SKY130_FD_SC_LP__SDFXTP_LP%A_351_417# 1 2 3 4 13 18 22 23 24 27 31 36
+ 38 40 42
c101 42 0 1.73585e-19 $X=6.72 $Y=1.88
c102 31 0 1.68639e-19 $X=7.155 $Y=0.97
c103 27 0 1.16549e-19 $X=6.72 $Y=2.59
r104 39 42 8.33333 $w=6.08e-07 $l=4.25e-07 $layer=LI1_cond $X=6.295 $Y=2.02
+ $X2=6.72 $Y2=2.02
r105 39 40 8.65265 $w=6.08e-07 $l=8.5e-08 $layer=LI1_cond $X=6.295 $Y=2.02
+ $X2=6.21 $Y2=2.02
r106 34 36 5.22619 $w=4.28e-07 $l=1.95e-07 $layer=LI1_cond $X=2.365 $Y=0.82
+ $X2=2.56 $Y2=0.82
r107 29 31 8.52808 $w=2.48e-07 $l=1.85e-07 $layer=LI1_cond $X=7.195 $Y=0.785
+ $X2=7.195 $Y2=0.97
r108 25 42 4.33422 $w=3.3e-07 $l=3.05e-07 $layer=LI1_cond $X=6.72 $Y=2.325
+ $X2=6.72 $Y2=2.02
r109 25 27 9.25447 $w=3.28e-07 $l=2.65e-07 $layer=LI1_cond $X=6.72 $Y=2.325
+ $X2=6.72 $Y2=2.59
r110 23 29 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=7.07 $Y=0.7
+ $X2=7.195 $Y2=0.785
r111 23 24 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=7.07 $Y=0.7 $X2=6.38
+ $Y2=0.7
r112 22 39 8.42348 $w=1.7e-07 $l=3.05e-07 $layer=LI1_cond $X=6.295 $Y=1.715
+ $X2=6.295 $Y2=2.02
r113 21 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.295 $Y=0.785
+ $X2=6.38 $Y2=0.7
r114 21 22 60.6738 $w=1.68e-07 $l=9.3e-07 $layer=LI1_cond $X=6.295 $Y=0.785
+ $X2=6.295 $Y2=1.715
r115 20 38 4.23118 $w=2.15e-07 $l=1.05119e-07 $layer=LI1_cond $X=2.645 $Y=2.24
+ $X2=2.56 $Y2=2.195
r116 20 40 232.583 $w=1.68e-07 $l=3.565e-06 $layer=LI1_cond $X=2.645 $Y=2.24
+ $X2=6.21 $Y2=2.24
r117 18 38 2.20034 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.56 $Y=2.065
+ $X2=2.56 $Y2=2.195
r118 17 36 6.22023 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=2.56 $Y=1.035
+ $X2=2.56 $Y2=0.82
r119 17 18 67.1979 $w=1.68e-07 $l=1.03e-06 $layer=LI1_cond $X=2.56 $Y=1.035
+ $X2=2.56 $Y2=2.065
r120 13 38 4.23118 $w=2.15e-07 $l=8.5e-08 $layer=LI1_cond $X=2.475 $Y=2.195
+ $X2=2.56 $Y2=2.195
r121 13 15 25.7083 $w=2.58e-07 $l=5.8e-07 $layer=LI1_cond $X=2.475 $Y=2.195
+ $X2=1.895 $Y2=2.195
r122 4 42 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=6.575
+ $Y=1.735 $X2=6.72 $Y2=1.88
r123 4 27 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=6.575
+ $Y=1.735 $X2=6.72 $Y2=2.59
r124 3 15 600 $w=1.7e-07 $l=2.08567e-07 $layer=licon1_PDIFF $count=1 $X=1.755
+ $Y=2.085 $X2=1.895 $Y2=2.235
r125 2 31 182 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_NDIFF $count=1 $X=7.015
+ $Y=0.775 $X2=7.155 $Y2=0.97
r126 1 34 182 $w=1.7e-07 $l=3.02159e-07 $layer=licon1_NDIFF $count=1 $X=2.145
+ $Y=0.625 $X2=2.365 $Y2=0.82
.ends

.subckt PM_SKY130_FD_SC_LP__SDFXTP_LP%Q 1 2 10 13 14 15 28
r30 19 31 3.03483 $w=6.68e-07 $l=1.7e-07 $layer=LI1_cond $X=12.94 $Y=2.255
+ $X2=12.94 $Y2=2.085
r31 15 25 0.357038 $w=6.68e-07 $l=2e-08 $layer=LI1_cond $X=12.94 $Y=2.775
+ $X2=12.94 $Y2=2.795
r32 14 15 6.60521 $w=6.68e-07 $l=3.7e-07 $layer=LI1_cond $X=12.94 $Y=2.405
+ $X2=12.94 $Y2=2.775
r33 14 19 2.67779 $w=6.68e-07 $l=1.5e-07 $layer=LI1_cond $X=12.94 $Y=2.405
+ $X2=12.94 $Y2=2.255
r34 13 31 0.892596 $w=6.68e-07 $l=5e-08 $layer=LI1_cond $X=12.94 $Y=2.035
+ $X2=12.94 $Y2=2.085
r35 13 28 9.71911 $w=6.68e-07 $l=1.15e-07 $layer=LI1_cond $X=12.94 $Y=2.035
+ $X2=12.94 $Y2=1.92
r36 12 28 74.0481 $w=1.68e-07 $l=1.135e-06 $layer=LI1_cond $X=12.99 $Y=0.785
+ $X2=12.99 $Y2=1.92
r37 10 12 10.5284 $w=3.88e-07 $l=2.3e-07 $layer=LI1_cond $X=12.88 $Y=0.555
+ $X2=12.88 $Y2=0.785
r38 2 31 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=12.965
+ $Y=1.94 $X2=13.11 $Y2=2.085
r39 2 25 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=12.965
+ $Y=1.94 $X2=13.11 $Y2=2.795
r40 1 10 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=12.705
+ $Y=0.345 $X2=12.85 $Y2=0.555
.ends

.subckt PM_SKY130_FD_SC_LP__SDFXTP_LP%VGND 1 2 3 4 5 6 21 25 29 33 37 39 41 44
+ 45 46 48 53 58 63 75 83 86 89 92 96
r132 95 96 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.68 $Y=0
+ $X2=13.68 $Y2=0
r133 92 93 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=8.4 $Y=0
+ $X2=8.4 $Y2=0
r134 89 90 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r135 86 87 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r136 83 84 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r137 81 96 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.2 $Y=0
+ $X2=13.68 $Y2=0
r138 80 81 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=13.2 $Y=0 $X2=13.2
+ $Y2=0
r139 78 81 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=11.76 $Y=0
+ $X2=13.2 $Y2=0
r140 77 80 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=11.76 $Y=0
+ $X2=13.2 $Y2=0
r141 77 78 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.76 $Y=0
+ $X2=11.76 $Y2=0
r142 75 95 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=13.475 $Y=0
+ $X2=13.697 $Y2=0
r143 75 80 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=13.475 $Y=0
+ $X2=13.2 $Y2=0
r144 74 78 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=0
+ $X2=11.76 $Y2=0
r145 74 93 0.802756 $w=4.9e-07 $l=2.88e-06 $layer=MET1_cond $X=11.28 $Y=0
+ $X2=8.4 $Y2=0
r146 73 74 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=11.28 $Y=0
+ $X2=11.28 $Y2=0
r147 71 92 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.41 $Y=0 $X2=8.245
+ $Y2=0
r148 71 73 187.241 $w=1.68e-07 $l=2.87e-06 $layer=LI1_cond $X=8.41 $Y=0
+ $X2=11.28 $Y2=0
r149 70 93 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=8.4
+ $Y2=0
r150 69 70 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=7.92 $Y=0
+ $X2=7.92 $Y2=0
r151 67 90 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=4.56
+ $Y2=0
r152 66 69 187.893 $w=1.68e-07 $l=2.88e-06 $layer=LI1_cond $X=5.04 $Y=0 $X2=7.92
+ $Y2=0
r153 66 67 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=5.04 $Y=0
+ $X2=5.04 $Y2=0
r154 64 89 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.765 $Y=0 $X2=4.6
+ $Y2=0
r155 64 66 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=4.765 $Y=0
+ $X2=5.04 $Y2=0
r156 63 92 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.08 $Y=0 $X2=8.245
+ $Y2=0
r157 63 69 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=8.08 $Y=0 $X2=7.92
+ $Y2=0
r158 62 90 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=4.56
+ $Y2=0
r159 62 87 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.12
+ $Y2=0
r160 61 62 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r161 59 86 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.42 $Y=0 $X2=3.255
+ $Y2=0
r162 59 61 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=3.42 $Y=0 $X2=4.08
+ $Y2=0
r163 58 89 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.435 $Y=0 $X2=4.6
+ $Y2=0
r164 58 61 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=4.435 $Y=0
+ $X2=4.08 $Y2=0
r165 57 87 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.68 $Y=0
+ $X2=3.12 $Y2=0
r166 57 84 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r167 56 57 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r168 54 83 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.49 $Y=0 $X2=1.325
+ $Y2=0
r169 54 56 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=1.49 $Y=0 $X2=1.68
+ $Y2=0
r170 53 86 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.09 $Y=0 $X2=3.255
+ $Y2=0
r171 53 56 91.9893 $w=1.68e-07 $l=1.41e-06 $layer=LI1_cond $X=3.09 $Y=0 $X2=1.68
+ $Y2=0
r172 51 84 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r173 50 51 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r174 48 83 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.16 $Y=0 $X2=1.325
+ $Y2=0
r175 48 50 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=1.16 $Y=0 $X2=0.24
+ $Y2=0
r176 46 70 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=7.92
+ $Y2=0
r177 46 67 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=6.96 $Y=0
+ $X2=5.04 $Y2=0
r178 44 73 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=11.34 $Y=0 $X2=11.28
+ $Y2=0
r179 44 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.34 $Y=0
+ $X2=11.505 $Y2=0
r180 43 77 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=11.67 $Y=0 $X2=11.76
+ $Y2=0
r181 43 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.67 $Y=0
+ $X2=11.505 $Y2=0
r182 39 95 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=13.64 $Y=0.085
+ $X2=13.697 $Y2=0
r183 39 41 16.4136 $w=3.28e-07 $l=4.7e-07 $layer=LI1_cond $X=13.64 $Y=0.085
+ $X2=13.64 $Y2=0.555
r184 35 45 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=11.505 $Y=0.085
+ $X2=11.505 $Y2=0
r185 35 37 16.4136 $w=3.28e-07 $l=4.7e-07 $layer=LI1_cond $X=11.505 $Y=0.085
+ $X2=11.505 $Y2=0.555
r186 31 92 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.245 $Y=0.085
+ $X2=8.245 $Y2=0
r187 31 33 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=8.245 $Y=0.085
+ $X2=8.245 $Y2=0.55
r188 27 89 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.6 $Y=0.085 $X2=4.6
+ $Y2=0
r189 27 29 13.7944 $w=3.28e-07 $l=3.95e-07 $layer=LI1_cond $X=4.6 $Y=0.085
+ $X2=4.6 $Y2=0.48
r190 23 86 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.255 $Y=0.085
+ $X2=3.255 $Y2=0
r191 23 25 26.1919 $w=3.28e-07 $l=7.5e-07 $layer=LI1_cond $X=3.255 $Y=0.085
+ $X2=3.255 $Y2=0.835
r192 19 83 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.325 $Y=0.085
+ $X2=1.325 $Y2=0
r193 19 21 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=1.325 $Y=0.085
+ $X2=1.325 $Y2=0.795
r194 6 41 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=13.5
+ $Y=0.345 $X2=13.64 $Y2=0.555
r195 5 37 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=11.365
+ $Y=0.345 $X2=11.505 $Y2=0.555
r196 4 33 182 $w=1.7e-07 $l=2.497e-07 $layer=licon1_NDIFF $count=1 $X=8.03
+ $Y=0.625 $X2=8.245 $Y2=0.55
r197 3 29 182 $w=1.7e-07 $l=2.08567e-07 $layer=licon1_NDIFF $count=1 $X=4.46
+ $Y=0.33 $X2=4.6 $Y2=0.48
r198 2 25 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=3.115
+ $Y=0.625 $X2=3.255 $Y2=0.835
r199 1 21 182 $w=1.7e-07 $l=2.29565e-07 $layer=licon1_NDIFF $count=1 $X=1.185
+ $Y=0.625 $X2=1.325 $Y2=0.795
.ends

.subckt PM_SKY130_FD_SC_LP__SDFXTP_LP%A_1160_155# 1 2 9 11 12 15
r35 13 15 16.3647 $w=2.48e-07 $l=3.55e-07 $layer=LI1_cond $X=7.7 $Y=0.435
+ $X2=7.7 $Y2=0.79
r36 11 13 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=7.575 $Y=0.35
+ $X2=7.7 $Y2=0.435
r37 11 12 100.797 $w=1.68e-07 $l=1.545e-06 $layer=LI1_cond $X=7.575 $Y=0.35
+ $X2=6.03 $Y2=0.35
r38 7 12 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=5.905 $Y=0.435
+ $X2=6.03 $Y2=0.35
r39 7 9 23.2793 $w=2.48e-07 $l=5.05e-07 $layer=LI1_cond $X=5.905 $Y=0.435
+ $X2=5.905 $Y2=0.94
r40 2 15 182 $w=1.7e-07 $l=2.26164e-07 $layer=licon1_NDIFF $count=1 $X=7.595
+ $Y=0.625 $X2=7.74 $Y2=0.79
r41 1 9 182 $w=1.7e-07 $l=2.26164e-07 $layer=licon1_NDIFF $count=1 $X=5.8
+ $Y=0.775 $X2=5.945 $Y2=0.94
.ends

.subckt PM_SKY130_FD_SC_LP__SDFXTP_LP%A_1910_155# 1 2 9 11 12 15
r32 13 15 2.76586 $w=2.48e-07 $l=6e-08 $layer=LI1_cond $X=11.035 $Y=0.615
+ $X2=11.035 $Y2=0.555
r33 11 13 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=10.91 $Y=0.7
+ $X2=11.035 $Y2=0.615
r34 11 12 74.3743 $w=1.68e-07 $l=1.14e-06 $layer=LI1_cond $X=10.91 $Y=0.7
+ $X2=9.77 $Y2=0.7
r35 7 12 7.07814 $w=1.7e-07 $l=1.56844e-07 $layer=LI1_cond $X=9.65 $Y=0.785
+ $X2=9.77 $Y2=0.7
r36 7 9 9.60369 $w=2.38e-07 $l=2e-07 $layer=LI1_cond $X=9.65 $Y=0.785 $X2=9.65
+ $Y2=0.985
r37 2 15 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=10.935
+ $Y=0.345 $X2=11.075 $Y2=0.555
r38 1 9 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=9.55
+ $Y=0.775 $X2=9.675 $Y2=0.985
.ends

