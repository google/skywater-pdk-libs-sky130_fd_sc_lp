* File: sky130_fd_sc_lp__mux2_m.pxi.spice
* Created: Fri Aug 28 10:44:36 2020
* 
x_PM_SKY130_FD_SC_LP__MUX2_M%A_123_269# N_A_123_269#_M1004_d
+ N_A_123_269#_M1001_d N_A_123_269#_M1010_g N_A_123_269#_M1000_g
+ N_A_123_269#_c_81_n N_A_123_269#_c_90_n N_A_123_269#_c_82_n
+ N_A_123_269#_c_83_n N_A_123_269#_c_84_n N_A_123_269#_c_85_n
+ N_A_123_269#_c_86_n N_A_123_269#_c_87_n N_A_123_269#_c_100_p
+ PM_SKY130_FD_SC_LP__MUX2_M%A_123_269#
x_PM_SKY130_FD_SC_LP__MUX2_M%S N_S_M1007_g N_S_M1003_g N_S_M1002_g N_S_M1006_g
+ N_S_c_161_n N_S_c_162_n N_S_c_163_n N_S_c_164_n N_S_c_165_n N_S_c_214_p
+ N_S_c_166_n N_S_c_167_n N_S_c_168_n S S S N_S_c_157_n N_S_c_172_n
+ PM_SKY130_FD_SC_LP__MUX2_M%S
x_PM_SKY130_FD_SC_LP__MUX2_M%A1 N_A1_M1004_g N_A1_M1011_g N_A1_c_260_n
+ N_A1_c_261_n N_A1_c_262_n A1 N_A1_c_263_n N_A1_c_267_n
+ PM_SKY130_FD_SC_LP__MUX2_M%A1
x_PM_SKY130_FD_SC_LP__MUX2_M%A0 N_A0_M1001_g N_A0_M1009_g N_A0_c_320_n
+ N_A0_c_321_n A0 A0 PM_SKY130_FD_SC_LP__MUX2_M%A0
x_PM_SKY130_FD_SC_LP__MUX2_M%A_483_99# N_A_483_99#_M1002_d N_A_483_99#_M1006_d
+ N_A_483_99#_c_362_n N_A_483_99#_M1008_g N_A_483_99#_M1005_g
+ N_A_483_99#_c_364_n N_A_483_99#_c_365_n N_A_483_99#_c_366_n
+ N_A_483_99#_c_367_n N_A_483_99#_c_368_n N_A_483_99#_c_371_n
+ PM_SKY130_FD_SC_LP__MUX2_M%A_483_99#
x_PM_SKY130_FD_SC_LP__MUX2_M%X N_X_M1010_s N_X_M1000_s N_X_c_419_n X X X X X
+ N_X_c_422_n PM_SKY130_FD_SC_LP__MUX2_M%X
x_PM_SKY130_FD_SC_LP__MUX2_M%VPWR N_VPWR_M1000_d N_VPWR_M1005_d N_VPWR_c_437_n
+ N_VPWR_c_438_n VPWR N_VPWR_c_439_n N_VPWR_c_440_n N_VPWR_c_441_n
+ N_VPWR_c_436_n N_VPWR_c_443_n N_VPWR_c_444_n PM_SKY130_FD_SC_LP__MUX2_M%VPWR
x_PM_SKY130_FD_SC_LP__MUX2_M%VGND N_VGND_M1010_d N_VGND_M1008_d N_VGND_c_482_n
+ N_VGND_c_483_n N_VGND_c_484_n N_VGND_c_485_n N_VGND_c_486_n N_VGND_c_487_n
+ VGND N_VGND_c_488_n N_VGND_c_489_n PM_SKY130_FD_SC_LP__MUX2_M%VGND
cc_1 VNB N_A_123_269#_M1010_g 0.0310882f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=0.835
cc_2 VNB N_A_123_269#_c_81_n 0.0112017f $X=-0.19 $Y=-0.245 $X2=0.78 $Y2=1.85
cc_3 VNB N_A_123_269#_c_82_n 8.34889e-19 $X=-0.19 $Y=-0.245 $X2=0.78 $Y2=1.51
cc_4 VNB N_A_123_269#_c_83_n 0.0184605f $X=-0.19 $Y=-0.245 $X2=0.78 $Y2=1.51
cc_5 VNB N_A_123_269#_c_84_n 0.0206598f $X=-0.19 $Y=-0.245 $X2=1.64 $Y2=1.18
cc_6 VNB N_A_123_269#_c_85_n 7.20038e-19 $X=-0.19 $Y=-0.245 $X2=0.865 $Y2=1.18
cc_7 VNB N_A_123_269#_c_86_n 0.00305491f $X=-0.19 $Y=-0.245 $X2=2.03 $Y2=2.525
cc_8 VNB N_A_123_269#_c_87_n 0.00482358f $X=-0.19 $Y=-0.245 $X2=1.805 $Y2=0.9
cc_9 VNB N_S_M1007_g 0.0426173f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_S_M1002_g 0.0478461f $X=-0.19 $Y=-0.245 $X2=0.87 $Y2=2.015
cc_11 VNB S 0.00263926f $X=-0.19 $Y=-0.245 $X2=2.145 $Y2=2.62
cc_12 VNB N_S_c_157_n 0.0102036f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A1_c_260_n 0.0175036f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=0.835
cc_14 VNB N_A1_c_261_n 0.0469489f $X=-0.19 $Y=-0.245 $X2=0.87 $Y2=2.015
cc_15 VNB N_A1_c_262_n 0.0100883f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A1_c_263_n 0.0138832f $X=-0.19 $Y=-0.245 $X2=0.78 $Y2=1.265
cc_17 VNB N_A0_M1009_g 0.0345471f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.345
cc_18 VNB N_A0_c_320_n 0.0171146f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=0.835
cc_19 VNB N_A0_c_321_n 0.0258488f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB A0 0.00382325f $X=-0.19 $Y=-0.245 $X2=0.87 $Y2=2.715
cc_21 VNB N_A_483_99#_c_362_n 0.0172251f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.345
cc_22 VNB N_A_483_99#_M1005_g 0.0098499f $X=-0.19 $Y=-0.245 $X2=0.87 $Y2=2.715
cc_23 VNB N_A_483_99#_c_364_n 0.0109497f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_483_99#_c_365_n 0.0356632f $X=-0.19 $Y=-0.245 $X2=0.78 $Y2=1.345
cc_25 VNB N_A_483_99#_c_366_n 0.0164698f $X=-0.19 $Y=-0.245 $X2=0.78 $Y2=1.85
cc_26 VNB N_A_483_99#_c_367_n 0.00385342f $X=-0.19 $Y=-0.245 $X2=0.78 $Y2=1.51
cc_27 VNB N_A_483_99#_c_368_n 0.0448136f $X=-0.19 $Y=-0.245 $X2=0.78 $Y2=1.51
cc_28 VNB N_X_c_419_n 0.0231748f $X=-0.19 $Y=-0.245 $X2=0.87 $Y2=2.015
cc_29 VNB X 0.0371901f $X=-0.19 $Y=-0.245 $X2=0.87 $Y2=2.715
cc_30 VNB N_VPWR_c_436_n 0.163682f $X=-0.19 $Y=-0.245 $X2=2.03 $Y2=1.265
cc_31 VNB N_VGND_c_482_n 0.0216998f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=0.835
cc_32 VNB N_VGND_c_483_n 0.0249774f $X=-0.19 $Y=-0.245 $X2=0.87 $Y2=2.715
cc_33 VNB N_VGND_c_484_n 0.0250501f $X=-0.19 $Y=-0.245 $X2=0.78 $Y2=1.345
cc_34 VNB N_VGND_c_485_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0.78 $Y2=1.85
cc_35 VNB N_VGND_c_486_n 0.039711f $X=-0.19 $Y=-0.245 $X2=0.78 $Y2=1.265
cc_36 VNB N_VGND_c_487_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0.78 $Y2=1.51
cc_37 VNB N_VGND_c_488_n 0.0296693f $X=-0.19 $Y=-0.245 $X2=2.145 $Y2=2.63
cc_38 VNB N_VGND_c_489_n 0.26107f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VPB N_A_123_269#_M1000_g 0.0458668f $X=-0.19 $Y=1.655 $X2=0.87 $Y2=2.715
cc_40 VPB N_A_123_269#_c_81_n 0.0150862f $X=-0.19 $Y=1.655 $X2=0.78 $Y2=1.85
cc_41 VPB N_A_123_269#_c_90_n 0.0183919f $X=-0.19 $Y=1.655 $X2=0.78 $Y2=2.015
cc_42 VPB N_A_123_269#_c_82_n 0.00239474f $X=-0.19 $Y=1.655 $X2=0.78 $Y2=1.51
cc_43 VPB N_A_123_269#_c_86_n 0.00632834f $X=-0.19 $Y=1.655 $X2=2.03 $Y2=2.525
cc_44 VPB N_S_M1007_g 0.0186813f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_45 VPB N_S_M1003_g 0.0188421f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=1.345
cc_46 VPB N_S_M1006_g 0.0287707f $X=-0.19 $Y=1.655 $X2=0.78 $Y2=1.51
cc_47 VPB N_S_c_161_n 0.023181f $X=-0.19 $Y=1.655 $X2=0.78 $Y2=1.265
cc_48 VPB N_S_c_162_n 0.016409f $X=-0.19 $Y=1.655 $X2=0.78 $Y2=1.51
cc_49 VPB N_S_c_163_n 0.00203614f $X=-0.19 $Y=1.655 $X2=0.78 $Y2=1.51
cc_50 VPB N_S_c_164_n 0.00872809f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_51 VPB N_S_c_165_n 0.0023193f $X=-0.19 $Y=1.655 $X2=1.64 $Y2=1.18
cc_52 VPB N_S_c_166_n 0.00681702f $X=-0.19 $Y=1.655 $X2=1.805 $Y2=1.03
cc_53 VPB N_S_c_167_n 0.0464646f $X=-0.19 $Y=1.655 $X2=1.805 $Y2=0.9
cc_54 VPB N_S_c_168_n 0.00319185f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_55 VPB S 0.00588731f $X=-0.19 $Y=1.655 $X2=2.145 $Y2=2.62
cc_56 VPB S 0.0060616f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_57 VPB N_S_c_157_n 0.00617517f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_58 VPB N_S_c_172_n 0.00125681f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_59 VPB N_A1_M1011_g 0.0287141f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_60 VPB N_A1_c_262_n 0.00296412f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_61 VPB A1 0.00605864f $X=-0.19 $Y=1.655 $X2=0.78 $Y2=1.51
cc_62 VPB N_A1_c_267_n 0.0372942f $X=-0.19 $Y=1.655 $X2=0.78 $Y2=1.51
cc_63 VPB N_A0_M1001_g 0.0453768f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_64 VPB N_A0_c_320_n 0.0187172f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=0.835
cc_65 VPB N_A0_c_321_n 0.00533794f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_66 VPB A0 0.00403547f $X=-0.19 $Y=1.655 $X2=0.87 $Y2=2.715
cc_67 VPB N_A_483_99#_M1005_g 0.0543191f $X=-0.19 $Y=1.655 $X2=0.87 $Y2=2.715
cc_68 VPB N_A_483_99#_c_366_n 0.0456087f $X=-0.19 $Y=1.655 $X2=0.78 $Y2=1.85
cc_69 VPB N_A_483_99#_c_371_n 0.00856322f $X=-0.19 $Y=1.655 $X2=1.805 $Y2=0.9
cc_70 VPB X 0.0454062f $X=-0.19 $Y=1.655 $X2=0.87 $Y2=2.715
cc_71 VPB N_X_c_422_n 0.0297367f $X=-0.19 $Y=1.655 $X2=0.78 $Y2=1.51
cc_72 VPB N_VPWR_c_437_n 0.00863591f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=0.835
cc_73 VPB N_VPWR_c_438_n 0.00886042f $X=-0.19 $Y=1.655 $X2=0.87 $Y2=2.715
cc_74 VPB N_VPWR_c_439_n 0.0283233f $X=-0.19 $Y=1.655 $X2=0.78 $Y2=1.85
cc_75 VPB N_VPWR_c_440_n 0.0400224f $X=-0.19 $Y=1.655 $X2=0.78 $Y2=1.51
cc_76 VPB N_VPWR_c_441_n 0.0200707f $X=-0.19 $Y=1.655 $X2=1.805 $Y2=0.9
cc_77 VPB N_VPWR_c_436_n 0.0834331f $X=-0.19 $Y=1.655 $X2=2.03 $Y2=1.265
cc_78 VPB N_VPWR_c_443_n 0.00632158f $X=-0.19 $Y=1.655 $X2=2.145 $Y2=2.62
cc_79 VPB N_VPWR_c_444_n 0.0063235f $X=-0.19 $Y=1.655 $X2=0.78 $Y2=1.51
cc_80 N_A_123_269#_M1010_g N_S_M1007_g 0.0214014f $X=0.72 $Y=0.835 $X2=0 $Y2=0
cc_81 N_A_123_269#_c_82_n N_S_M1007_g 0.00371897f $X=0.78 $Y=1.51 $X2=0 $Y2=0
cc_82 N_A_123_269#_c_83_n N_S_M1007_g 0.0325448f $X=0.78 $Y=1.51 $X2=0 $Y2=0
cc_83 N_A_123_269#_c_84_n N_S_M1007_g 0.0160967f $X=1.64 $Y=1.18 $X2=0 $Y2=0
cc_84 N_A_123_269#_c_86_n N_S_M1007_g 0.00498144f $X=2.03 $Y=2.525 $X2=0 $Y2=0
cc_85 N_A_123_269#_c_87_n N_S_M1007_g 0.00133101f $X=1.805 $Y=0.9 $X2=0 $Y2=0
cc_86 N_A_123_269#_M1000_g N_S_M1003_g 0.00872137f $X=0.87 $Y=2.715 $X2=0 $Y2=0
cc_87 N_A_123_269#_c_100_p N_S_M1003_g 5.07427e-19 $X=2.145 $Y=2.63 $X2=0 $Y2=0
cc_88 N_A_123_269#_M1000_g N_S_c_163_n 0.00272239f $X=0.87 $Y=2.715 $X2=0 $Y2=0
cc_89 N_A_123_269#_c_100_p N_S_c_163_n 0.00807903f $X=2.145 $Y=2.63 $X2=0 $Y2=0
cc_90 N_A_123_269#_M1001_d N_S_c_164_n 0.00181172f $X=2.005 $Y=2.505 $X2=0 $Y2=0
cc_91 N_A_123_269#_c_100_p N_S_c_164_n 0.0160334f $X=2.145 $Y=2.63 $X2=0 $Y2=0
cc_92 N_A_123_269#_M1000_g N_S_c_165_n 3.07046e-19 $X=0.87 $Y=2.715 $X2=0 $Y2=0
cc_93 N_A_123_269#_M1000_g N_S_c_166_n 0.00140682f $X=0.87 $Y=2.715 $X2=0 $Y2=0
cc_94 N_A_123_269#_c_86_n N_S_c_166_n 0.0217113f $X=2.03 $Y=2.525 $X2=0 $Y2=0
cc_95 N_A_123_269#_c_90_n N_S_c_167_n 0.0325448f $X=0.78 $Y=2.015 $X2=0 $Y2=0
cc_96 N_A_123_269#_c_86_n N_S_c_167_n 0.00118604f $X=2.03 $Y=2.525 $X2=0 $Y2=0
cc_97 N_A_123_269#_c_86_n N_S_c_168_n 0.00795073f $X=2.03 $Y=2.525 $X2=0 $Y2=0
cc_98 N_A_123_269#_c_86_n N_A1_M1011_g 0.00505242f $X=2.03 $Y=2.525 $X2=0 $Y2=0
cc_99 N_A_123_269#_c_100_p N_A1_M1011_g 0.00301393f $X=2.145 $Y=2.63 $X2=0 $Y2=0
cc_100 N_A_123_269#_c_84_n N_A1_c_260_n 0.00272017f $X=1.64 $Y=1.18 $X2=0 $Y2=0
cc_101 N_A_123_269#_c_87_n N_A1_c_260_n 0.0159609f $X=1.805 $Y=0.9 $X2=0 $Y2=0
cc_102 N_A_123_269#_c_87_n N_A1_c_261_n 0.00378298f $X=1.805 $Y=0.9 $X2=0 $Y2=0
cc_103 N_A_123_269#_c_86_n N_A1_c_262_n 0.0399004f $X=2.03 $Y=2.525 $X2=0 $Y2=0
cc_104 N_A_123_269#_c_87_n N_A1_c_262_n 0.0274244f $X=1.805 $Y=0.9 $X2=0 $Y2=0
cc_105 N_A_123_269#_c_86_n A1 0.0242054f $X=2.03 $Y=2.525 $X2=0 $Y2=0
cc_106 N_A_123_269#_c_100_p A1 5.9134e-19 $X=2.145 $Y=2.63 $X2=0 $Y2=0
cc_107 N_A_123_269#_c_84_n N_A1_c_263_n 0.00587197f $X=1.64 $Y=1.18 $X2=0 $Y2=0
cc_108 N_A_123_269#_c_87_n N_A1_c_263_n 0.00785555f $X=1.805 $Y=0.9 $X2=0 $Y2=0
cc_109 N_A_123_269#_c_86_n N_A1_c_267_n 0.00207715f $X=2.03 $Y=2.525 $X2=0 $Y2=0
cc_110 N_A_123_269#_c_100_p N_A1_c_267_n 0.00134601f $X=2.145 $Y=2.63 $X2=0
+ $Y2=0
cc_111 N_A_123_269#_c_86_n N_A0_M1001_g 0.0185114f $X=2.03 $Y=2.525 $X2=0 $Y2=0
cc_112 N_A_123_269#_c_100_p N_A0_M1001_g 0.00395635f $X=2.145 $Y=2.63 $X2=0
+ $Y2=0
cc_113 N_A_123_269#_c_86_n N_A0_M1009_g 0.00522081f $X=2.03 $Y=2.525 $X2=0 $Y2=0
cc_114 N_A_123_269#_c_87_n N_A0_M1009_g 0.0103327f $X=1.805 $Y=0.9 $X2=0 $Y2=0
cc_115 N_A_123_269#_c_84_n N_A0_c_320_n 7.55478e-19 $X=1.64 $Y=1.18 $X2=0 $Y2=0
cc_116 N_A_123_269#_c_87_n N_A0_c_320_n 0.0103006f $X=1.805 $Y=0.9 $X2=0 $Y2=0
cc_117 N_A_123_269#_c_86_n N_A0_c_321_n 0.0169681f $X=2.03 $Y=2.525 $X2=0 $Y2=0
cc_118 N_A_123_269#_c_82_n A0 0.0197579f $X=0.78 $Y=1.51 $X2=0 $Y2=0
cc_119 N_A_123_269#_c_83_n A0 0.00239893f $X=0.78 $Y=1.51 $X2=0 $Y2=0
cc_120 N_A_123_269#_c_84_n A0 0.0382331f $X=1.64 $Y=1.18 $X2=0 $Y2=0
cc_121 N_A_123_269#_c_86_n A0 0.0237693f $X=2.03 $Y=2.525 $X2=0 $Y2=0
cc_122 N_A_123_269#_c_87_n A0 0.00979518f $X=1.805 $Y=0.9 $X2=0 $Y2=0
cc_123 N_A_123_269#_c_86_n N_A_483_99#_M1005_g 5.39447e-19 $X=2.03 $Y=2.525
+ $X2=0 $Y2=0
cc_124 N_A_123_269#_M1010_g N_X_c_419_n 9.09816e-19 $X=0.72 $Y=0.835 $X2=0 $Y2=0
cc_125 N_A_123_269#_M1010_g X 0.00923556f $X=0.72 $Y=0.835 $X2=0 $Y2=0
cc_126 N_A_123_269#_M1000_g X 0.0125408f $X=0.87 $Y=2.715 $X2=0 $Y2=0
cc_127 N_A_123_269#_c_82_n X 0.0300059f $X=0.78 $Y=1.51 $X2=0 $Y2=0
cc_128 N_A_123_269#_c_83_n X 0.0142383f $X=0.78 $Y=1.51 $X2=0 $Y2=0
cc_129 N_A_123_269#_c_85_n X 0.00756562f $X=0.865 $Y=1.18 $X2=0 $Y2=0
cc_130 N_A_123_269#_c_90_n N_X_c_422_n 0.00278999f $X=0.78 $Y=2.015 $X2=0 $Y2=0
cc_131 N_A_123_269#_c_82_n N_X_c_422_n 0.00182811f $X=0.78 $Y=1.51 $X2=0 $Y2=0
cc_132 N_A_123_269#_M1000_g N_VPWR_c_437_n 0.011947f $X=0.87 $Y=2.715 $X2=0
+ $Y2=0
cc_133 N_A_123_269#_M1000_g N_VPWR_c_439_n 0.00532616f $X=0.87 $Y=2.715 $X2=0
+ $Y2=0
cc_134 N_A_123_269#_M1000_g N_VPWR_c_436_n 0.00520409f $X=0.87 $Y=2.715 $X2=0
+ $Y2=0
cc_135 N_A_123_269#_M1010_g N_VGND_c_482_n 0.00816798f $X=0.72 $Y=0.835 $X2=0
+ $Y2=0
cc_136 N_A_123_269#_c_83_n N_VGND_c_482_n 3.86999e-19 $X=0.78 $Y=1.51 $X2=0
+ $Y2=0
cc_137 N_A_123_269#_c_84_n N_VGND_c_482_n 0.0166127f $X=1.64 $Y=1.18 $X2=0 $Y2=0
cc_138 N_A_123_269#_c_85_n N_VGND_c_482_n 0.00345655f $X=0.865 $Y=1.18 $X2=0
+ $Y2=0
cc_139 N_A_123_269#_M1010_g N_VGND_c_484_n 0.00400585f $X=0.72 $Y=0.835 $X2=0
+ $Y2=0
cc_140 N_A_123_269#_M1010_g N_VGND_c_489_n 0.00456913f $X=0.72 $Y=0.835 $X2=0
+ $Y2=0
cc_141 N_S_c_164_n N_A1_M1011_g 0.0136626f $X=2.49 $Y=2.98 $X2=0 $Y2=0
cc_142 N_S_c_168_n N_A1_M1011_g 0.00204216f $X=2.66 $Y=2.43 $X2=0 $Y2=0
cc_143 N_S_M1007_g N_A1_c_261_n 0.0418195f $X=1.23 $Y=0.835 $X2=0 $Y2=0
cc_144 N_S_M1002_g N_A1_c_262_n 0.00130589f $X=3.19 $Y=0.835 $X2=0 $Y2=0
cc_145 S N_A1_c_262_n 0.00864873f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_146 N_S_c_168_n A1 0.0142776f $X=2.66 $Y=2.43 $X2=0 $Y2=0
cc_147 S A1 0.0183776f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_148 S A1 0.0049139f $X=3.035 $Y=2.32 $X2=0 $Y2=0
cc_149 N_S_c_168_n N_A1_c_267_n 0.00127495f $X=2.66 $Y=2.43 $X2=0 $Y2=0
cc_150 N_S_M1007_g N_A0_M1001_g 0.00540716f $X=1.23 $Y=0.835 $X2=0 $Y2=0
cc_151 N_S_c_164_n N_A0_M1001_g 0.0124319f $X=2.49 $Y=2.98 $X2=0 $Y2=0
cc_152 N_S_c_166_n N_A0_M1001_g 0.00391891f $X=1.45 $Y=2.18 $X2=0 $Y2=0
cc_153 N_S_c_167_n N_A0_M1001_g 0.0597606f $X=1.45 $Y=2.18 $X2=0 $Y2=0
cc_154 N_S_M1007_g N_A0_c_320_n 0.0214021f $X=1.23 $Y=0.835 $X2=0 $Y2=0
cc_155 N_S_c_166_n N_A0_c_320_n 3.67457e-19 $X=1.45 $Y=2.18 $X2=0 $Y2=0
cc_156 N_S_c_167_n N_A0_c_320_n 0.00638866f $X=1.45 $Y=2.18 $X2=0 $Y2=0
cc_157 N_S_M1007_g A0 0.0173882f $X=1.23 $Y=0.835 $X2=0 $Y2=0
cc_158 N_S_c_166_n A0 0.0156793f $X=1.45 $Y=2.18 $X2=0 $Y2=0
cc_159 N_S_c_167_n A0 0.00363454f $X=1.45 $Y=2.18 $X2=0 $Y2=0
cc_160 N_S_M1002_g N_A_483_99#_c_362_n 0.00980193f $X=3.19 $Y=0.835 $X2=0 $Y2=0
cc_161 N_S_M1006_g N_A_483_99#_M1005_g 0.0185157f $X=3.34 $Y=2.715 $X2=0 $Y2=0
cc_162 N_S_c_161_n N_A_483_99#_M1005_g 0.0331052f $X=3.28 $Y=2.085 $X2=0 $Y2=0
cc_163 N_S_c_164_n N_A_483_99#_M1005_g 0.00141792f $X=2.49 $Y=2.98 $X2=0 $Y2=0
cc_164 N_S_c_214_p N_A_483_99#_M1005_g 0.00566712f $X=2.575 $Y=2.895 $X2=0 $Y2=0
cc_165 S N_A_483_99#_M1005_g 0.00967861f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_166 S N_A_483_99#_M1005_g 0.0163057f $X=3.035 $Y=2.32 $X2=0 $Y2=0
cc_167 N_S_M1002_g N_A_483_99#_c_364_n 0.0108813f $X=3.19 $Y=0.835 $X2=0 $Y2=0
cc_168 S N_A_483_99#_c_364_n 0.0118756f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_169 N_S_M1002_g N_A_483_99#_c_365_n 0.0146856f $X=3.19 $Y=0.835 $X2=0 $Y2=0
cc_170 S N_A_483_99#_c_365_n 0.00787497f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_171 N_S_c_157_n N_A_483_99#_c_365_n 0.00415972f $X=3.28 $Y=1.745 $X2=0 $Y2=0
cc_172 N_S_M1002_g N_A_483_99#_c_366_n 0.0076894f $X=3.19 $Y=0.835 $X2=0 $Y2=0
cc_173 N_S_M1006_g N_A_483_99#_c_366_n 0.00928484f $X=3.34 $Y=2.715 $X2=0 $Y2=0
cc_174 S N_A_483_99#_c_366_n 0.053802f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_175 N_S_c_157_n N_A_483_99#_c_366_n 0.0163119f $X=3.28 $Y=1.745 $X2=0 $Y2=0
cc_176 N_S_c_172_n N_A_483_99#_c_366_n 0.012125f $X=3.2 $Y=2.345 $X2=0 $Y2=0
cc_177 N_S_M1002_g N_A_483_99#_c_367_n 9.79826e-19 $X=3.19 $Y=0.835 $X2=0 $Y2=0
cc_178 N_S_M1002_g N_A_483_99#_c_368_n 0.0331052f $X=3.19 $Y=0.835 $X2=0 $Y2=0
cc_179 N_S_M1006_g N_A_483_99#_c_371_n 0.00382191f $X=3.34 $Y=2.715 $X2=0 $Y2=0
cc_180 S N_VPWR_M1005_d 7.71375e-19 $X=3.035 $Y=2.32 $X2=0 $Y2=0
cc_181 N_S_c_172_n N_VPWR_M1005_d 0.00201013f $X=3.2 $Y=2.345 $X2=0 $Y2=0
cc_182 N_S_M1003_g N_VPWR_c_437_n 0.00145676f $X=1.57 $Y=2.715 $X2=0 $Y2=0
cc_183 N_S_c_165_n N_VPWR_c_437_n 0.0130038f $X=1.62 $Y=2.98 $X2=0 $Y2=0
cc_184 N_S_c_167_n N_VPWR_c_437_n 0.0046512f $X=1.45 $Y=2.18 $X2=0 $Y2=0
cc_185 N_S_M1006_g N_VPWR_c_438_n 0.00483713f $X=3.34 $Y=2.715 $X2=0 $Y2=0
cc_186 N_S_c_162_n N_VPWR_c_438_n 4.58839e-19 $X=3.28 $Y=2.25 $X2=0 $Y2=0
cc_187 N_S_c_164_n N_VPWR_c_438_n 0.0118055f $X=2.49 $Y=2.98 $X2=0 $Y2=0
cc_188 N_S_c_214_p N_VPWR_c_438_n 0.0120785f $X=2.575 $Y=2.895 $X2=0 $Y2=0
cc_189 S N_VPWR_c_438_n 0.00718783f $X=3.035 $Y=2.32 $X2=0 $Y2=0
cc_190 N_S_c_172_n N_VPWR_c_438_n 0.0142864f $X=3.2 $Y=2.345 $X2=0 $Y2=0
cc_191 N_S_M1003_g N_VPWR_c_440_n 9.47275e-19 $X=1.57 $Y=2.715 $X2=0 $Y2=0
cc_192 N_S_c_164_n N_VPWR_c_440_n 0.0642094f $X=2.49 $Y=2.98 $X2=0 $Y2=0
cc_193 N_S_c_165_n N_VPWR_c_440_n 0.0114622f $X=1.62 $Y=2.98 $X2=0 $Y2=0
cc_194 N_S_M1006_g N_VPWR_c_441_n 0.00527534f $X=3.34 $Y=2.715 $X2=0 $Y2=0
cc_195 N_S_M1006_g N_VPWR_c_436_n 0.00534666f $X=3.34 $Y=2.715 $X2=0 $Y2=0
cc_196 N_S_c_164_n N_VPWR_c_436_n 0.0390945f $X=2.49 $Y=2.98 $X2=0 $Y2=0
cc_197 N_S_c_165_n N_VPWR_c_436_n 0.00657784f $X=1.62 $Y=2.98 $X2=0 $Y2=0
cc_198 S N_VPWR_c_436_n 0.00787748f $X=3.035 $Y=2.32 $X2=0 $Y2=0
cc_199 N_S_c_172_n N_VPWR_c_436_n 0.00640354f $X=3.2 $Y=2.345 $X2=0 $Y2=0
cc_200 N_S_c_164_n A_329_501# 0.00366293f $X=2.49 $Y=2.98 $X2=-0.19 $Y2=-0.245
cc_201 N_S_c_164_n A_487_501# 3.57886e-19 $X=2.49 $Y=2.98 $X2=-0.19 $Y2=-0.245
cc_202 N_S_c_214_p A_487_501# 0.0052497f $X=2.575 $Y=2.895 $X2=-0.19 $Y2=-0.245
cc_203 S A_487_501# 7.27958e-19 $X=3.035 $Y=2.32 $X2=-0.19 $Y2=-0.245
cc_204 N_S_M1007_g N_VGND_c_482_n 0.00509061f $X=1.23 $Y=0.835 $X2=0 $Y2=0
cc_205 N_S_M1002_g N_VGND_c_483_n 0.00896845f $X=3.19 $Y=0.835 $X2=0 $Y2=0
cc_206 N_S_M1007_g N_VGND_c_486_n 0.00415323f $X=1.23 $Y=0.835 $X2=0 $Y2=0
cc_207 N_S_M1002_g N_VGND_c_488_n 0.00415323f $X=3.19 $Y=0.835 $X2=0 $Y2=0
cc_208 N_S_M1007_g N_VGND_c_489_n 0.00469432f $X=1.23 $Y=0.835 $X2=0 $Y2=0
cc_209 N_S_M1002_g N_VGND_c_489_n 0.00469432f $X=3.19 $Y=0.835 $X2=0 $Y2=0
cc_210 N_A1_M1011_g N_A0_M1001_g 0.0240221f $X=2.36 $Y=2.715 $X2=0 $Y2=0
cc_211 A1 N_A0_M1001_g 2.96039e-19 $X=2.555 $Y=1.95 $X2=0 $Y2=0
cc_212 N_A1_c_267_n N_A0_M1001_g 0.0203599f $X=2.38 $Y=2 $X2=0 $Y2=0
cc_213 N_A1_c_260_n N_A0_M1009_g 0.00636409f $X=2.295 $Y=0.35 $X2=0 $Y2=0
cc_214 N_A1_c_261_n N_A0_M1009_g 0.00132287f $X=1.68 $Y=0.35 $X2=0 $Y2=0
cc_215 N_A1_c_262_n N_A0_M1009_g 0.0129117f $X=2.38 $Y=1.835 $X2=0 $Y2=0
cc_216 N_A1_c_263_n N_A0_M1009_g 0.0142479f $X=1.68 $Y=0.515 $X2=0 $Y2=0
cc_217 N_A1_c_263_n N_A0_c_320_n 0.00681988f $X=1.68 $Y=0.515 $X2=0 $Y2=0
cc_218 N_A1_c_262_n N_A0_c_321_n 0.00126829f $X=2.38 $Y=1.835 $X2=0 $Y2=0
cc_219 N_A1_c_262_n N_A_483_99#_c_362_n 0.0152283f $X=2.38 $Y=1.835 $X2=0 $Y2=0
cc_220 N_A1_M1011_g N_A_483_99#_M1005_g 0.0287143f $X=2.36 $Y=2.715 $X2=0 $Y2=0
cc_221 N_A1_c_262_n N_A_483_99#_M1005_g 0.00682487f $X=2.38 $Y=1.835 $X2=0 $Y2=0
cc_222 A1 N_A_483_99#_M1005_g 0.00315776f $X=2.555 $Y=1.95 $X2=0 $Y2=0
cc_223 N_A1_c_267_n N_A_483_99#_M1005_g 0.0192839f $X=2.38 $Y=2 $X2=0 $Y2=0
cc_224 N_A1_c_262_n N_A_483_99#_c_367_n 0.0211429f $X=2.38 $Y=1.835 $X2=0 $Y2=0
cc_225 A1 N_A_483_99#_c_367_n 0.00320098f $X=2.555 $Y=1.95 $X2=0 $Y2=0
cc_226 N_A1_c_262_n N_A_483_99#_c_368_n 0.00596033f $X=2.38 $Y=1.835 $X2=0 $Y2=0
cc_227 A1 N_A_483_99#_c_368_n 0.00457733f $X=2.555 $Y=1.95 $X2=0 $Y2=0
cc_228 N_A1_c_267_n N_A_483_99#_c_368_n 0.00305689f $X=2.38 $Y=2 $X2=0 $Y2=0
cc_229 N_A1_M1011_g N_VPWR_c_440_n 9.29198e-19 $X=2.36 $Y=2.715 $X2=0 $Y2=0
cc_230 N_A1_c_260_n N_VGND_c_482_n 0.00748978f $X=2.295 $Y=0.35 $X2=0 $Y2=0
cc_231 N_A1_c_261_n N_VGND_c_482_n 0.0055216f $X=1.68 $Y=0.35 $X2=0 $Y2=0
cc_232 N_A1_c_260_n N_VGND_c_483_n 0.0144411f $X=2.295 $Y=0.35 $X2=0 $Y2=0
cc_233 N_A1_c_262_n N_VGND_c_483_n 0.0316377f $X=2.38 $Y=1.835 $X2=0 $Y2=0
cc_234 N_A1_c_260_n N_VGND_c_486_n 0.0577846f $X=2.295 $Y=0.35 $X2=0 $Y2=0
cc_235 N_A1_c_261_n N_VGND_c_486_n 0.00651318f $X=1.68 $Y=0.35 $X2=0 $Y2=0
cc_236 N_A1_c_260_n N_VGND_c_489_n 0.0342139f $X=2.295 $Y=0.35 $X2=0 $Y2=0
cc_237 N_A1_c_261_n N_VGND_c_489_n 0.0101042f $X=1.68 $Y=0.35 $X2=0 $Y2=0
cc_238 N_A1_c_262_n A_441_125# 0.00454897f $X=2.38 $Y=1.835 $X2=-0.19 $Y2=-0.245
cc_239 N_A0_M1009_g N_A_483_99#_c_362_n 0.0472711f $X=2.13 $Y=0.835 $X2=0 $Y2=0
cc_240 N_A0_c_321_n N_A_483_99#_M1005_g 0.00161603f $X=1.93 $Y=1.595 $X2=0 $Y2=0
cc_241 N_A0_M1009_g N_A_483_99#_c_368_n 0.00458879f $X=2.13 $Y=0.835 $X2=0 $Y2=0
cc_242 N_A0_M1001_g N_VPWR_c_440_n 9.29198e-19 $X=1.93 $Y=2.715 $X2=0 $Y2=0
cc_243 N_A_483_99#_M1005_g N_VPWR_c_438_n 0.00650319f $X=2.83 $Y=2.715 $X2=0
+ $Y2=0
cc_244 N_A_483_99#_M1005_g N_VPWR_c_440_n 0.0045897f $X=2.83 $Y=2.715 $X2=0
+ $Y2=0
cc_245 N_A_483_99#_c_371_n N_VPWR_c_441_n 0.00863584f $X=3.635 $Y=2.775 $X2=0
+ $Y2=0
cc_246 N_A_483_99#_M1005_g N_VPWR_c_436_n 0.0044912f $X=2.83 $Y=2.715 $X2=0
+ $Y2=0
cc_247 N_A_483_99#_c_371_n N_VPWR_c_436_n 0.0108974f $X=3.635 $Y=2.775 $X2=0
+ $Y2=0
cc_248 N_A_483_99#_c_362_n N_VGND_c_483_n 0.0039041f $X=2.49 $Y=1.155 $X2=0
+ $Y2=0
cc_249 N_A_483_99#_c_364_n N_VGND_c_483_n 0.00829044f $X=3.24 $Y=1.24 $X2=0
+ $Y2=0
cc_250 N_A_483_99#_c_365_n N_VGND_c_483_n 0.00443335f $X=3.635 $Y=1.325 $X2=0
+ $Y2=0
cc_251 N_A_483_99#_c_367_n N_VGND_c_483_n 0.00948609f $X=2.74 $Y=1.32 $X2=0
+ $Y2=0
cc_252 N_A_483_99#_c_368_n N_VGND_c_483_n 0.00371641f $X=2.74 $Y=1.32 $X2=0
+ $Y2=0
cc_253 N_A_483_99#_c_362_n N_VGND_c_486_n 0.00296546f $X=2.49 $Y=1.155 $X2=0
+ $Y2=0
cc_254 N_A_483_99#_c_362_n N_VGND_c_489_n 0.00314612f $X=2.49 $Y=1.155 $X2=0
+ $Y2=0
cc_255 N_A_483_99#_c_365_n N_VGND_c_489_n 0.0130955f $X=3.635 $Y=1.325 $X2=0
+ $Y2=0
cc_256 N_X_c_422_n N_VPWR_c_439_n 0.0166896f $X=0.655 $Y=2.695 $X2=0 $Y2=0
cc_257 N_X_c_422_n N_VPWR_c_436_n 0.0200711f $X=0.655 $Y=2.695 $X2=0 $Y2=0
cc_258 N_X_c_419_n N_VGND_c_482_n 0.0120057f $X=0.505 $Y=0.75 $X2=0 $Y2=0
cc_259 N_X_c_419_n N_VGND_c_484_n 0.00970146f $X=0.505 $Y=0.75 $X2=0 $Y2=0
cc_260 N_X_c_419_n N_VGND_c_489_n 0.0138689f $X=0.505 $Y=0.75 $X2=0 $Y2=0
