* File: sky130_fd_sc_lp__nor3_0.pex.spice
* Created: Wed Sep  2 10:08:49 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__NOR3_0%A 2 5 6 8 10 11 13 16 18 19 20 21 27
r41 27 28 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.27
+ $Y=1.02 $X2=0.27 $Y2=1.02
r42 20 21 13.3251 $w=3.18e-07 $l=3.7e-07 $layer=LI1_cond $X=0.245 $Y=1.665
+ $X2=0.245 $Y2=2.035
r43 19 20 13.3251 $w=3.18e-07 $l=3.7e-07 $layer=LI1_cond $X=0.245 $Y=1.295
+ $X2=0.245 $Y2=1.665
r44 19 28 9.90381 $w=3.18e-07 $l=2.75e-07 $layer=LI1_cond $X=0.245 $Y=1.295
+ $X2=0.245 $Y2=1.02
r45 18 28 3.42132 $w=3.18e-07 $l=9.5e-08 $layer=LI1_cond $X=0.245 $Y=0.925
+ $X2=0.245 $Y2=1.02
r46 14 16 92.2979 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=0.36 $Y=2.23
+ $X2=0.54 $Y2=2.23
r47 12 27 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.27 $Y=1.36
+ $X2=0.27 $Y2=1.02
r48 12 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.27 $Y=1.36
+ $X2=0.27 $Y2=1.525
r49 11 27 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=0.27 $Y=1.005
+ $X2=0.27 $Y2=1.02
r50 10 11 43.5886 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=0.34 $Y=0.855
+ $X2=0.34 $Y2=1.005
r51 6 16 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.54 $Y=2.305
+ $X2=0.54 $Y2=2.23
r52 6 8 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=0.54 $Y=2.305 $X2=0.54
+ $Y2=2.735
r53 5 10 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.5 $Y=0.535 $X2=0.5
+ $Y2=0.855
r54 2 14 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.36 $Y=2.155
+ $X2=0.36 $Y2=2.23
r55 2 13 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=0.36 $Y=2.155
+ $X2=0.36 $Y2=1.525
.ends

.subckt PM_SKY130_FD_SC_LP__NOR3_0%B 3 7 11 12 13 14 15 16 17 25 36
r54 27 36 0.164635 $w=3.48e-07 $l=5e-09 $layer=LI1_cond $X=0.75 $Y=2.04 $X2=0.75
+ $Y2=2.035
r55 25 26 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.84
+ $Y=1.41 $X2=0.84 $Y2=1.41
r56 16 17 14.7036 $w=2.88e-07 $l=3.7e-07 $layer=LI1_cond $X=0.78 $Y=2.405
+ $X2=0.78 $Y2=2.775
r57 16 44 7.55049 $w=2.88e-07 $l=1.9e-07 $layer=LI1_cond $X=0.78 $Y=2.405
+ $X2=0.78 $Y2=2.215
r58 15 44 4.81789 $w=3.48e-07 $l=1.35e-07 $layer=LI1_cond $X=0.75 $Y=2.08
+ $X2=0.75 $Y2=2.215
r59 15 27 1.31708 $w=3.48e-07 $l=4e-08 $layer=LI1_cond $X=0.75 $Y=2.08 $X2=0.75
+ $Y2=2.04
r60 15 36 1.31708 $w=3.48e-07 $l=4e-08 $layer=LI1_cond $X=0.75 $Y=1.995 $X2=0.75
+ $Y2=2.035
r61 14 15 10.8659 $w=3.48e-07 $l=3.3e-07 $layer=LI1_cond $X=0.75 $Y=1.665
+ $X2=0.75 $Y2=1.995
r62 14 26 8.39637 $w=3.48e-07 $l=2.55e-07 $layer=LI1_cond $X=0.75 $Y=1.665
+ $X2=0.75 $Y2=1.41
r63 13 26 3.7866 $w=3.48e-07 $l=1.15e-07 $layer=LI1_cond $X=0.75 $Y=1.295
+ $X2=0.75 $Y2=1.41
r64 11 25 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.84 $Y=1.75
+ $X2=0.84 $Y2=1.41
r65 11 12 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.84 $Y=1.75
+ $X2=0.84 $Y2=1.915
r66 10 25 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.84 $Y=1.245
+ $X2=0.84 $Y2=1.41
r67 7 12 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=0.93 $Y=2.735
+ $X2=0.93 $Y2=1.915
r68 3 10 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=0.93 $Y=0.535
+ $X2=0.93 $Y2=1.245
.ends

.subckt PM_SKY130_FD_SC_LP__NOR3_0%C 3 7 11 12 13 14 15 20
r35 20 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.38
+ $Y=1.375 $X2=1.38 $Y2=1.375
r36 14 15 11.5244 $w=3.68e-07 $l=3.7e-07 $layer=LI1_cond $X=1.28 $Y=1.665
+ $X2=1.28 $Y2=2.035
r37 14 21 9.03266 $w=3.68e-07 $l=2.9e-07 $layer=LI1_cond $X=1.28 $Y=1.665
+ $X2=1.28 $Y2=1.375
r38 13 21 2.49177 $w=3.68e-07 $l=8e-08 $layer=LI1_cond $X=1.28 $Y=1.295 $X2=1.28
+ $Y2=1.375
r39 11 20 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.38 $Y=1.715
+ $X2=1.38 $Y2=1.375
r40 11 12 41.8716 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.38 $Y=1.715
+ $X2=1.38 $Y2=1.88
r41 10 20 38.6168 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.38 $Y=1.21
+ $X2=1.38 $Y2=1.375
r42 7 10 346.117 $w=1.5e-07 $l=6.75e-07 $layer=POLY_cond $X=1.36 $Y=0.535
+ $X2=1.36 $Y2=1.21
r43 3 12 438.415 $w=1.5e-07 $l=8.55e-07 $layer=POLY_cond $X=1.32 $Y=2.735
+ $X2=1.32 $Y2=1.88
.ends

.subckt PM_SKY130_FD_SC_LP__NOR3_0%VPWR 1 4 6 8 15 16
r19 19 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r20 15 16 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r21 13 20 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r22 12 15 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.72 $Y=3.33 $X2=1.68
+ $Y2=3.33
r23 12 13 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r24 10 19 4.4248 $w=1.7e-07 $l=2.33e-07 $layer=LI1_cond $X=0.465 $Y=3.33
+ $X2=0.232 $Y2=3.33
r25 10 12 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.465 $Y=3.33
+ $X2=0.72 $Y2=3.33
r26 8 16 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=0.96 $Y=3.33
+ $X2=1.68 $Y2=3.33
r27 8 13 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=0.96 $Y=3.33
+ $X2=0.72 $Y2=3.33
r28 4 19 3.13344 $w=3.05e-07 $l=1.18427e-07 $layer=LI1_cond $X=0.312 $Y=3.245
+ $X2=0.232 $Y2=3.33
r29 4 6 25.5049 $w=3.03e-07 $l=6.75e-07 $layer=LI1_cond $X=0.312 $Y=3.245
+ $X2=0.312 $Y2=2.57
r30 1 6 300 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_PDIFF $count=2 $X=0.2
+ $Y=2.415 $X2=0.325 $Y2=2.57
.ends

.subckt PM_SKY130_FD_SC_LP__NOR3_0%Y 1 2 3 10 12 17 18 20 21 22 27 33
r42 22 27 2.54441 $w=2e-07 $l=1.77e-07 $layer=LI1_cond $X=1.657 $Y=0.94 $X2=1.48
+ $Y2=0.94
r43 22 33 8.32279 $w=5.23e-07 $l=3.1e-07 $layer=LI1_cond $X=1.657 $Y=0.84
+ $X2=1.657 $Y2=0.53
r44 21 27 15.5273 $w=1.98e-07 $l=2.8e-07 $layer=LI1_cond $X=1.2 $Y=0.94 $X2=1.48
+ $Y2=0.94
r45 21 28 21.6273 $w=1.98e-07 $l=3.9e-07 $layer=LI1_cond $X=1.2 $Y=0.94 $X2=0.81
+ $Y2=0.94
r46 20 28 3.35255 $w=2e-07 $l=1.299e-07 $layer=LI1_cond $X=0.692 $Y=0.915
+ $X2=0.81 $Y2=0.94
r47 17 18 8.20593 $w=4.63e-07 $l=1.65e-07 $layer=LI1_cond $X=1.602 $Y=2.56
+ $X2=1.602 $Y2=2.395
r48 14 22 3.90249 $w=2.77e-07 $l=1.33417e-07 $layer=LI1_cond $X=1.735 $Y=1.04
+ $X2=1.657 $Y2=0.94
r49 14 18 75.1409 $w=1.98e-07 $l=1.355e-06 $layer=LI1_cond $X=1.735 $Y=1.04
+ $X2=1.735 $Y2=2.395
r50 10 20 3.46977 $w=1.9e-07 $l=1.36015e-07 $layer=LI1_cond $X=0.715 $Y=0.79
+ $X2=0.692 $Y2=0.915
r51 10 12 15.177 $w=1.88e-07 $l=2.6e-07 $layer=LI1_cond $X=0.715 $Y=0.79
+ $X2=0.715 $Y2=0.53
r52 3 17 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=1.395
+ $Y=2.415 $X2=1.535 $Y2=2.56
r53 2 33 182 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_NDIFF $count=1 $X=1.435
+ $Y=0.325 $X2=1.575 $Y2=0.53
r54 1 12 182 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_NDIFF $count=1 $X=0.575
+ $Y=0.325 $X2=0.715 $Y2=0.53
.ends

.subckt PM_SKY130_FD_SC_LP__NOR3_0%VGND 1 2 7 9 13 15 17 24 25 31
r28 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r29 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r30 25 32 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r31 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r32 22 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.31 $Y=0 $X2=1.145
+ $Y2=0
r33 22 24 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=1.31 $Y=0 $X2=1.68
+ $Y2=0
r34 21 29 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r35 20 21 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r36 18 28 4.72267 $w=1.7e-07 $l=2.25e-07 $layer=LI1_cond $X=0.45 $Y=0 $X2=0.225
+ $Y2=0
r37 18 20 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=0.45 $Y=0 $X2=0.72
+ $Y2=0
r38 17 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.98 $Y=0 $X2=1.145
+ $Y2=0
r39 17 20 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=0.98 $Y=0 $X2=0.72
+ $Y2=0
r40 15 32 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=0.96 $Y=0 $X2=1.2
+ $Y2=0
r41 15 21 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=0.96 $Y=0 $X2=0.72
+ $Y2=0
r42 11 31 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.145 $Y=0.085
+ $X2=1.145 $Y2=0
r43 11 13 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=1.145 $Y=0.085
+ $X2=1.145 $Y2=0.53
r44 7 28 3.0435 $w=3.3e-07 $l=1.11018e-07 $layer=LI1_cond $X=0.285 $Y=0.085
+ $X2=0.225 $Y2=0
r45 7 9 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=0.285 $Y=0.085
+ $X2=0.285 $Y2=0.53
r46 2 13 182 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_NDIFF $count=1 $X=1.005
+ $Y=0.325 $X2=1.145 $Y2=0.53
r47 1 9 182 $w=1.7e-07 $l=2.60096e-07 $layer=licon1_NDIFF $count=1 $X=0.16
+ $Y=0.325 $X2=0.285 $Y2=0.53
.ends

