* File: sky130_fd_sc_lp__o2bb2a_0.pex.spice
* Created: Fri Aug 28 11:11:29 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O2BB2A_0%A_80_176# 1 2 8 11 15 16 19 20 23 24 25 27
+ 28 29 31 32 33 36 39 40 44 47 48 50
c128 50 0 7.35861e-20 $X=0.58 $Y=0.88
c129 39 0 5.23505e-20 $X=2.29 $Y=2.175
c130 24 0 3.84136e-20 $X=1.005 $Y=2.385
r131 42 44 11.127 $w=2.88e-07 $l=2.8e-07 $layer=LI1_cond $X=2.72 $Y=2.345
+ $X2=2.72 $Y2=2.625
r132 41 48 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.375 $Y=2.26
+ $X2=2.29 $Y2=2.26
r133 40 42 7.43784 $w=1.7e-07 $l=1.8262e-07 $layer=LI1_cond $X=2.575 $Y=2.26
+ $X2=2.72 $Y2=2.345
r134 40 41 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=2.575 $Y=2.26
+ $X2=2.375 $Y2=2.26
r135 39 48 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.29 $Y=2.175
+ $X2=2.29 $Y2=2.26
r136 39 47 97.861 $w=1.68e-07 $l=1.5e-06 $layer=LI1_cond $X=2.29 $Y=2.175
+ $X2=2.29 $Y2=0.675
r137 34 47 6.82988 $w=2.43e-07 $l=1.22e-07 $layer=LI1_cond $X=2.252 $Y=0.553
+ $X2=2.252 $Y2=0.675
r138 34 36 5.08016 $w=2.43e-07 $l=1.08e-07 $layer=LI1_cond $X=2.252 $Y=0.553
+ $X2=2.252 $Y2=0.445
r139 32 48 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.205 $Y=2.26
+ $X2=2.29 $Y2=2.26
r140 32 33 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=2.205 $Y=2.26
+ $X2=1.975 $Y2=2.26
r141 30 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.89 $Y=2.345
+ $X2=1.975 $Y2=2.26
r142 30 31 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=1.89 $Y=2.345
+ $X2=1.89 $Y2=2.905
r143 28 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.805 $Y=2.99
+ $X2=1.89 $Y2=2.905
r144 28 29 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=1.805 $Y=2.99
+ $X2=1.175 $Y2=2.99
r145 27 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.09 $Y=2.905
+ $X2=1.175 $Y2=2.99
r146 26 27 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=1.09 $Y=2.47
+ $X2=1.09 $Y2=2.905
r147 24 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.005 $Y=2.385
+ $X2=1.09 $Y2=2.47
r148 24 25 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=1.005 $Y=2.385
+ $X2=0.715 $Y2=2.385
r149 23 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.63 $Y=2.3
+ $X2=0.715 $Y2=2.385
r150 23 46 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=0.63 $Y=2.3
+ $X2=0.63 $Y2=1.55
r151 20 50 46.5827 $w=3.6e-07 $l=1.65e-07 $layer=POLY_cond $X=0.58 $Y=1.045
+ $X2=0.58 $Y2=0.88
r152 19 20 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.595
+ $Y=1.045 $X2=0.595 $Y2=1.045
r153 17 46 6.3875 $w=2.18e-07 $l=1.1e-07 $layer=LI1_cond $X=0.605 $Y=1.44
+ $X2=0.605 $Y2=1.55
r154 17 19 20.6916 $w=2.18e-07 $l=3.95e-07 $layer=LI1_cond $X=0.605 $Y=1.44
+ $X2=0.605 $Y2=1.045
r155 15 50 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.615 $Y=0.56
+ $X2=0.615 $Y2=0.88
r156 11 16 607.628 $w=1.5e-07 $l=1.185e-06 $layer=POLY_cond $X=0.475 $Y=2.735
+ $X2=0.475 $Y2=1.55
r157 8 16 48.987 $w=3.6e-07 $l=1.8e-07 $layer=POLY_cond $X=0.58 $Y=1.37 $X2=0.58
+ $Y2=1.55
r158 7 20 2.40434 $w=3.6e-07 $l=1.5e-08 $layer=POLY_cond $X=0.58 $Y=1.06
+ $X2=0.58 $Y2=1.045
r159 7 8 49.6898 $w=3.6e-07 $l=3.1e-07 $layer=POLY_cond $X=0.58 $Y=1.06 $X2=0.58
+ $Y2=1.37
r160 2 44 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=2.56
+ $Y=2.415 $X2=2.7 $Y2=2.625
r161 1 36 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=2.145
+ $Y=0.235 $X2=2.27 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__O2BB2A_0%A1_N 3 7 9 10 14
c42 14 0 4.04207e-19 $X=0.98 $Y=1.955
c43 3 0 3.73452e-20 $X=1.045 $Y=0.56
r44 14 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.98 $Y=1.955
+ $X2=0.98 $Y2=2.12
r45 14 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.98 $Y=1.955
+ $X2=0.98 $Y2=1.79
r46 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.98
+ $Y=1.955 $X2=0.98 $Y2=1.955
r47 10 15 2.24867 $w=4.08e-07 $l=8e-08 $layer=LI1_cond $X=1.09 $Y=2.035 $X2=1.09
+ $Y2=1.955
r48 9 15 8.15143 $w=4.08e-07 $l=2.9e-07 $layer=LI1_cond $X=1.09 $Y=1.665
+ $X2=1.09 $Y2=1.955
r49 7 17 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=1.07 $Y=2.625
+ $X2=1.07 $Y2=2.12
r50 3 16 630.702 $w=1.5e-07 $l=1.23e-06 $layer=POLY_cond $X=1.045 $Y=0.56
+ $X2=1.045 $Y2=1.79
.ends

.subckt PM_SKY130_FD_SC_LP__O2BB2A_0%A2_N 3 6 7 9 12 14 15 22 34
c59 34 0 1.87835e-19 $X=1.227 $Y=1.12
c60 12 0 9.07641e-20 $X=1.645 $Y=2.23
r61 26 34 4.34926 $w=2.45e-07 $l=2.6e-07 $layer=LI1_cond $X=1.227 $Y=0.86
+ $X2=1.227 $Y2=1.12
r62 23 34 8.02561 $w=4.53e-07 $l=2.98e-07 $layer=LI1_cond $X=1.525 $Y=1.12
+ $X2=1.227 $Y2=1.12
r63 22 25 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.525 $Y=1.18
+ $X2=1.525 $Y2=1.345
r64 22 24 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.525 $Y=1.18
+ $X2=1.525 $Y2=1.015
r65 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.525
+ $Y=1.18 $X2=1.525 $Y2=1.18
r66 15 34 0.727152 $w=4.53e-07 $l=2.7e-08 $layer=LI1_cond $X=1.2 $Y=1.12
+ $X2=1.227 $Y2=1.12
r67 15 26 0.470385 $w=2.43e-07 $l=1e-08 $layer=LI1_cond $X=1.227 $Y=0.85
+ $X2=1.227 $Y2=0.86
r68 14 15 13.8764 $w=2.43e-07 $l=2.95e-07 $layer=LI1_cond $X=1.227 $Y=0.555
+ $X2=1.227 $Y2=0.85
r69 10 12 94.8617 $w=1.5e-07 $l=1.85e-07 $layer=POLY_cond $X=1.46 $Y=2.23
+ $X2=1.645 $Y2=2.23
r70 7 12 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.645 $Y=2.305
+ $X2=1.645 $Y2=2.23
r71 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.645 $Y=2.305
+ $X2=1.645 $Y2=2.625
r72 6 10 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.46 $Y=2.155
+ $X2=1.46 $Y2=2.23
r73 6 25 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=1.46 $Y=2.155 $X2=1.46
+ $Y2=1.345
r74 3 24 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=1.435 $Y=0.56
+ $X2=1.435 $Y2=1.015
.ends

.subckt PM_SKY130_FD_SC_LP__O2BB2A_0%A_229_483# 1 2 10 11 12 13 14 15 17 20 23
+ 25 29 32 35 39 42
c89 32 0 1.43406e-19 $X=1.875 $Y=1.75
c90 23 0 1.83897e-19 $X=1.55 $Y=2.405
c91 11 0 9.75757e-20 $X=2.41 $Y=0.84
r92 37 39 7.85757 $w=3.28e-07 $l=2.25e-07 $layer=LI1_cond $X=1.65 $Y=0.56
+ $X2=1.875 $Y2=0.56
r93 35 43 46.255 $w=3.35e-07 $l=1.65e-07 $layer=POLY_cond $X=1.942 $Y=1.75
+ $X2=1.942 $Y2=1.915
r94 35 42 46.255 $w=3.35e-07 $l=1.65e-07 $layer=POLY_cond $X=1.942 $Y=1.75
+ $X2=1.942 $Y2=1.585
r95 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.94
+ $Y=1.75 $X2=1.94 $Y2=1.75
r96 32 34 3.33193 $w=2.38e-07 $l=6.5e-08 $layer=LI1_cond $X=1.875 $Y=1.75
+ $X2=1.94 $Y2=1.75
r97 31 32 16.6597 $w=2.38e-07 $l=3.25e-07 $layer=LI1_cond $X=1.55 $Y=1.75
+ $X2=1.875 $Y2=1.75
r98 27 29 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=1.43 $Y=2.57 $X2=1.55
+ $Y2=2.57
r99 25 32 2.70854 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.875 $Y=1.585
+ $X2=1.875 $Y2=1.75
r100 24 39 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.875 $Y=0.725
+ $X2=1.875 $Y2=0.56
r101 24 25 56.107 $w=1.68e-07 $l=8.6e-07 $layer=LI1_cond $X=1.875 $Y=0.725
+ $X2=1.875 $Y2=1.585
r102 23 29 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.55 $Y=2.405
+ $X2=1.55 $Y2=2.57
r103 22 31 2.70854 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.55 $Y=1.915
+ $X2=1.55 $Y2=1.75
r104 22 23 31.9679 $w=1.68e-07 $l=4.9e-07 $layer=LI1_cond $X=1.55 $Y=1.915
+ $X2=1.55 $Y2=2.405
r105 18 20 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=2.485 $Y=2.215
+ $X2=2.485 $Y2=2.625
r106 15 17 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.485 $Y=0.765
+ $X2=2.485 $Y2=0.445
r107 13 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.41 $Y=2.14
+ $X2=2.485 $Y2=2.215
r108 13 14 153.83 $w=1.5e-07 $l=3e-07 $layer=POLY_cond $X=2.41 $Y=2.14 $X2=2.11
+ $Y2=2.14
r109 11 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.41 $Y=0.84
+ $X2=2.485 $Y2=0.765
r110 11 12 153.83 $w=1.5e-07 $l=3e-07 $layer=POLY_cond $X=2.41 $Y=0.84 $X2=2.11
+ $Y2=0.84
r111 10 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.035 $Y=2.065
+ $X2=2.11 $Y2=2.14
r112 10 43 76.9149 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=2.035 $Y=2.065
+ $X2=2.035 $Y2=1.915
r113 7 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.035 $Y=0.915
+ $X2=2.11 $Y2=0.84
r114 7 42 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=2.035 $Y=0.915
+ $X2=2.035 $Y2=1.585
r115 2 27 600 $w=1.7e-07 $l=3.54119e-07 $layer=licon1_PDIFF $count=1 $X=1.145
+ $Y=2.415 $X2=1.43 $Y2=2.57
r116 1 37 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.51
+ $Y=0.35 $X2=1.65 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_LP__O2BB2A_0%B2 3 7 11 12 13 14 18
c40 18 0 6.45449e-20 $X=2.825 $Y=1.32
c41 13 0 9.75757e-20 $X=2.64 $Y=1.295
c42 11 0 1.4009e-19 $X=2.825 $Y=1.66
r43 18 19 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.825
+ $Y=1.32 $X2=2.825 $Y2=1.32
r44 14 19 8.93467 $w=4.43e-07 $l=3.45e-07 $layer=LI1_cond $X=2.767 $Y=1.665
+ $X2=2.767 $Y2=1.32
r45 13 19 0.64744 $w=4.43e-07 $l=2.5e-08 $layer=LI1_cond $X=2.767 $Y=1.295
+ $X2=2.767 $Y2=1.32
r46 11 18 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.825 $Y=1.66
+ $X2=2.825 $Y2=1.32
r47 11 12 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.825 $Y=1.66
+ $X2=2.825 $Y2=1.825
r48 10 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.825 $Y=1.155
+ $X2=2.825 $Y2=1.32
r49 7 12 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=2.915 $Y=2.625
+ $X2=2.915 $Y2=1.825
r50 3 10 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=2.915 $Y=0.445
+ $X2=2.915 $Y2=1.155
.ends

.subckt PM_SKY130_FD_SC_LP__O2BB2A_0%B1 3 7 11 12 13 14 15 20
r32 20 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.365
+ $Y=1.71 $X2=3.365 $Y2=1.71
r33 15 21 7.00406 $w=5.53e-07 $l=3.25e-07 $layer=LI1_cond $X=3.477 $Y=2.035
+ $X2=3.477 $Y2=1.71
r34 14 21 0.969793 $w=5.53e-07 $l=4.5e-08 $layer=LI1_cond $X=3.477 $Y=1.665
+ $X2=3.477 $Y2=1.71
r35 13 14 7.97386 $w=5.53e-07 $l=3.7e-07 $layer=LI1_cond $X=3.477 $Y=1.295
+ $X2=3.477 $Y2=1.665
r36 11 20 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=3.365 $Y=2.05
+ $X2=3.365 $Y2=1.71
r37 11 12 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.365 $Y=2.05
+ $X2=3.365 $Y2=2.215
r38 10 20 38.6168 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.365 $Y=1.545
+ $X2=3.365 $Y2=1.71
r39 7 10 564.043 $w=1.5e-07 $l=1.1e-06 $layer=POLY_cond $X=3.345 $Y=0.445
+ $X2=3.345 $Y2=1.545
r40 3 12 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=3.275 $Y=2.625
+ $X2=3.275 $Y2=2.215
.ends

.subckt PM_SKY130_FD_SC_LP__O2BB2A_0%X 1 2 9 11 12 13 14 15 16 40 43
r19 43 44 0.625011 $w=2.58e-07 $l=1e-08 $layer=LI1_cond $X=0.225 $Y=2.405
+ $X2=0.225 $Y2=2.395
r20 24 35 2.85155 $w=2.3e-07 $l=1.65e-07 $layer=LI1_cond $X=0.21 $Y=0.71
+ $X2=0.21 $Y2=0.545
r21 16 43 1.64002 $w=2.58e-07 $l=3.7e-08 $layer=LI1_cond $X=0.225 $Y=2.442
+ $X2=0.225 $Y2=2.405
r22 16 44 1.90404 $w=2.28e-07 $l=3.8e-08 $layer=LI1_cond $X=0.21 $Y=2.357
+ $X2=0.21 $Y2=2.395
r23 15 16 16.1342 $w=2.28e-07 $l=3.22e-07 $layer=LI1_cond $X=0.21 $Y=2.035
+ $X2=0.21 $Y2=2.357
r24 14 15 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.21 $Y=1.665
+ $X2=0.21 $Y2=2.035
r25 13 14 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.21 $Y=1.295
+ $X2=0.21 $Y2=1.665
r26 12 13 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.21 $Y=0.925
+ $X2=0.21 $Y2=1.295
r27 12 24 10.7728 $w=2.28e-07 $l=2.15e-07 $layer=LI1_cond $X=0.21 $Y=0.925
+ $X2=0.21 $Y2=0.71
r28 11 40 5.5876 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=0.24 $Y=0.545 $X2=0.4
+ $Y2=0.545
r29 11 35 1.04768 $w=3.28e-07 $l=3e-08 $layer=LI1_cond $X=0.24 $Y=0.545 $X2=0.21
+ $Y2=0.545
r30 7 16 3.67895 $w=2.58e-07 $l=8.3e-08 $layer=LI1_cond $X=0.225 $Y=2.525
+ $X2=0.225 $Y2=2.442
r31 7 9 1.55137 $w=2.58e-07 $l=3.5e-08 $layer=LI1_cond $X=0.225 $Y=2.525
+ $X2=0.225 $Y2=2.56
r32 2 9 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.415 $X2=0.26 $Y2=2.56
r33 1 40 182 $w=1.7e-07 $l=2.498e-07 $layer=licon1_NDIFF $count=1 $X=0.275
+ $Y=0.35 $X2=0.4 $Y2=0.545
.ends

.subckt PM_SKY130_FD_SC_LP__O2BB2A_0%VPWR 1 2 3 12 16 18 20 22 24 29 34 40 43 47
r54 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r55 43 44 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r56 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r57 38 47 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r58 38 44 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.16 $Y2=3.33
r59 37 38 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r60 35 43 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.405 $Y=3.33
+ $X2=2.275 $Y2=3.33
r61 35 37 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=2.405 $Y=3.33
+ $X2=3.12 $Y2=3.33
r62 34 46 4.59886 $w=1.7e-07 $l=2.57e-07 $layer=LI1_cond $X=3.325 $Y=3.33
+ $X2=3.582 $Y2=3.33
r63 34 37 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=3.325 $Y=3.33
+ $X2=3.12 $Y2=3.33
r64 33 41 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r65 32 33 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r66 30 40 8.23795 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=0.835 $Y=3.33
+ $X2=0.68 $Y2=3.33
r67 30 32 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.835 $Y=3.33
+ $X2=1.2 $Y2=3.33
r68 29 43 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.145 $Y=3.33
+ $X2=2.275 $Y2=3.33
r69 29 32 61.6524 $w=1.68e-07 $l=9.45e-07 $layer=LI1_cond $X=2.145 $Y=3.33
+ $X2=1.2 $Y2=3.33
r70 27 41 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r71 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r72 24 40 8.23795 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=0.525 $Y=3.33
+ $X2=0.68 $Y2=3.33
r73 24 26 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.525 $Y=3.33
+ $X2=0.24 $Y2=3.33
r74 22 44 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=2.16 $Y2=3.33
r75 22 33 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=1.2 $Y2=3.33
r76 18 46 3.16731 $w=3.3e-07 $l=1.27609e-07 $layer=LI1_cond $X=3.49 $Y=3.245
+ $X2=3.582 $Y2=3.33
r77 18 20 21.652 $w=3.28e-07 $l=6.2e-07 $layer=LI1_cond $X=3.49 $Y=3.245
+ $X2=3.49 $Y2=2.625
r78 14 43 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=2.275 $Y=3.245
+ $X2=2.275 $Y2=3.33
r79 14 16 24.6002 $w=2.58e-07 $l=5.55e-07 $layer=LI1_cond $X=2.275 $Y=3.245
+ $X2=2.275 $Y2=2.69
r80 10 40 0.701276 $w=3.1e-07 $l=8.5e-08 $layer=LI1_cond $X=0.68 $Y=3.245
+ $X2=0.68 $Y2=3.33
r81 10 12 16.3573 $w=3.08e-07 $l=4.4e-07 $layer=LI1_cond $X=0.68 $Y=3.245
+ $X2=0.68 $Y2=2.805
r82 3 20 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=3.35
+ $Y=2.415 $X2=3.49 $Y2=2.625
r83 2 16 600 $w=1.7e-07 $l=6.42962e-07 $layer=licon1_PDIFF $count=1 $X=1.72
+ $Y=2.415 $X2=2.24 $Y2=2.69
r84 1 12 600 $w=1.7e-07 $l=4.54643e-07 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=2.415 $X2=0.69 $Y2=2.805
.ends

.subckt PM_SKY130_FD_SC_LP__O2BB2A_0%VGND 1 2 11 15 17 19 29 30 33 36
r46 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r47 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r48 30 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=3.12
+ $Y2=0
r49 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r50 27 36 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.26 $Y=0 $X2=3.13
+ $Y2=0
r51 27 29 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=3.26 $Y=0 $X2=3.6
+ $Y2=0
r52 26 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r53 25 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r54 23 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r55 22 25 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.64
+ $Y2=0
r56 22 23 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r57 20 33 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.935 $Y=0 $X2=0.805
+ $Y2=0
r58 20 22 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.935 $Y=0 $X2=1.2
+ $Y2=0
r59 19 36 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3 $Y=0 $X2=3.13 $Y2=0
r60 19 25 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=3 $Y=0 $X2=2.64
+ $Y2=0
r61 17 26 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=2.64
+ $Y2=0
r62 17 23 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=1.2
+ $Y2=0
r63 13 36 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=3.13 $Y=0.085
+ $X2=3.13 $Y2=0
r64 13 15 15.9569 $w=2.58e-07 $l=3.6e-07 $layer=LI1_cond $X=3.13 $Y=0.085
+ $X2=3.13 $Y2=0.445
r65 9 33 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=0.805 $Y=0.085
+ $X2=0.805 $Y2=0
r66 9 11 19.5029 $w=2.58e-07 $l=4.4e-07 $layer=LI1_cond $X=0.805 $Y=0.085
+ $X2=0.805 $Y2=0.525
r67 2 15 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.99
+ $Y=0.235 $X2=3.13 $Y2=0.445
r68 1 11 182 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=1 $X=0.69
+ $Y=0.35 $X2=0.83 $Y2=0.525
.ends

.subckt PM_SKY130_FD_SC_LP__O2BB2A_0%A_512_47# 1 2 9 11 12 15
c26 11 0 6.45449e-20 $X=3.43 $Y=0.865
r27 13 15 13.0871 $w=2.93e-07 $l=3.35e-07 $layer=LI1_cond $X=3.577 $Y=0.78
+ $X2=3.577 $Y2=0.445
r28 11 13 7.47753 $w=1.7e-07 $l=1.84673e-07 $layer=LI1_cond $X=3.43 $Y=0.865
+ $X2=3.577 $Y2=0.78
r29 11 12 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=3.43 $Y=0.865 $X2=2.83
+ $Y2=0.865
r30 7 12 7.39867 $w=1.7e-07 $l=1.80566e-07 $layer=LI1_cond $X=2.687 $Y=0.78
+ $X2=2.83 $Y2=0.865
r31 7 9 13.5463 $w=2.83e-07 $l=3.35e-07 $layer=LI1_cond $X=2.687 $Y=0.78
+ $X2=2.687 $Y2=0.445
r32 2 15 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=3.42
+ $Y=0.235 $X2=3.56 $Y2=0.445
r33 1 9 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.56
+ $Y=0.235 $X2=2.7 $Y2=0.445
.ends

