* File: sky130_fd_sc_lp__a211o_4.pxi.spice
* Created: Fri Aug 28 09:47:39 2020
* 
x_PM_SKY130_FD_SC_LP__A211O_4%A_103_263# N_A_103_263#_M1002_s
+ N_A_103_263#_M1019_s N_A_103_263#_M1009_s N_A_103_263#_M1000_s
+ N_A_103_263#_M1001_g N_A_103_263#_M1006_g N_A_103_263#_M1007_g
+ N_A_103_263#_M1014_g N_A_103_263#_M1008_g N_A_103_263#_M1021_g
+ N_A_103_263#_M1013_g N_A_103_263#_M1023_g N_A_103_263#_c_123_n
+ N_A_103_263#_c_124_n N_A_103_263#_c_125_n N_A_103_263#_c_126_n
+ N_A_103_263#_c_221_p N_A_103_263#_c_137_n N_A_103_263#_c_263_p
+ N_A_103_263#_c_167_p N_A_103_263#_c_264_p N_A_103_263#_c_127_n
+ N_A_103_263#_c_278_p N_A_103_263#_c_128_n N_A_103_263#_c_129_n
+ N_A_103_263#_c_142_p N_A_103_263#_c_143_p N_A_103_263#_c_130_n
+ N_A_103_263#_c_131_n PM_SKY130_FD_SC_LP__A211O_4%A_103_263#
x_PM_SKY130_FD_SC_LP__A211O_4%B1 N_B1_M1002_g N_B1_M1015_g N_B1_M1016_g
+ N_B1_c_283_n N_B1_M1022_g N_B1_c_289_n N_B1_c_290_n B1 N_B1_c_284_n
+ N_B1_c_285_n PM_SKY130_FD_SC_LP__A211O_4%B1
x_PM_SKY130_FD_SC_LP__A211O_4%C1 N_C1_c_381_n N_C1_M1004_g N_C1_M1000_g
+ N_C1_c_383_n N_C1_M1019_g N_C1_M1010_g C1 N_C1_c_386_n
+ PM_SKY130_FD_SC_LP__A211O_4%C1
x_PM_SKY130_FD_SC_LP__A211O_4%A2 N_A2_M1005_g N_A2_M1012_g N_A2_M1017_g
+ N_A2_M1018_g N_A2_c_440_n N_A2_c_441_n A2 A2 A2 N_A2_c_444_n N_A2_c_450_n
+ PM_SKY130_FD_SC_LP__A211O_4%A2
x_PM_SKY130_FD_SC_LP__A211O_4%A1 N_A1_M1009_g N_A1_M1003_g N_A1_M1020_g
+ N_A1_M1011_g A1 N_A1_c_519_n N_A1_c_516_n PM_SKY130_FD_SC_LP__A211O_4%A1
x_PM_SKY130_FD_SC_LP__A211O_4%VPWR N_VPWR_M1001_d N_VPWR_M1006_d N_VPWR_M1021_d
+ N_VPWR_M1005_d N_VPWR_M1011_d N_VPWR_c_564_n N_VPWR_c_565_n N_VPWR_c_566_n
+ N_VPWR_c_567_n N_VPWR_c_568_n N_VPWR_c_569_n VPWR N_VPWR_c_570_n
+ N_VPWR_c_571_n N_VPWR_c_572_n N_VPWR_c_573_n N_VPWR_c_574_n N_VPWR_c_563_n
+ N_VPWR_c_576_n N_VPWR_c_577_n N_VPWR_c_578_n N_VPWR_c_579_n
+ PM_SKY130_FD_SC_LP__A211O_4%VPWR
x_PM_SKY130_FD_SC_LP__A211O_4%X N_X_M1007_d N_X_M1013_d N_X_M1001_s N_X_M1014_s
+ N_X_c_672_n N_X_c_673_n N_X_c_666_n N_X_c_709_n N_X_c_674_n N_X_c_720_p
+ N_X_c_667_n N_X_c_714_n N_X_c_694_n N_X_c_675_n N_X_c_668_n X X X X X
+ PM_SKY130_FD_SC_LP__A211O_4%X
x_PM_SKY130_FD_SC_LP__A211O_4%A_527_367# N_A_527_367#_M1015_s
+ N_A_527_367#_M1022_s N_A_527_367#_M1003_s N_A_527_367#_M1018_s
+ N_A_527_367#_c_735_n N_A_527_367#_c_738_n N_A_527_367#_c_784_n
+ N_A_527_367#_c_757_n N_A_527_367#_c_761_n N_A_527_367#_c_762_n
+ N_A_527_367#_c_730_n N_A_527_367#_c_731_n N_A_527_367#_c_769_n
+ N_A_527_367#_c_732_n PM_SKY130_FD_SC_LP__A211O_4%A_527_367#
x_PM_SKY130_FD_SC_LP__A211O_4%A_610_367# N_A_610_367#_M1015_d
+ N_A_610_367#_M1010_d N_A_610_367#_c_802_n
+ PM_SKY130_FD_SC_LP__A211O_4%A_610_367#
x_PM_SKY130_FD_SC_LP__A211O_4%VGND N_VGND_M1007_s N_VGND_M1008_s N_VGND_M1023_s
+ N_VGND_M1004_d N_VGND_M1016_d N_VGND_M1017_s N_VGND_c_817_n N_VGND_c_818_n
+ N_VGND_c_819_n N_VGND_c_820_n N_VGND_c_821_n N_VGND_c_822_n N_VGND_c_823_n
+ N_VGND_c_824_n N_VGND_c_825_n N_VGND_c_826_n VGND N_VGND_c_827_n
+ N_VGND_c_828_n N_VGND_c_829_n N_VGND_c_830_n N_VGND_c_831_n N_VGND_c_832_n
+ N_VGND_c_833_n N_VGND_c_834_n N_VGND_c_835_n PM_SKY130_FD_SC_LP__A211O_4%VGND
x_PM_SKY130_FD_SC_LP__A211O_4%A_1006_47# N_A_1006_47#_M1012_d
+ N_A_1006_47#_M1020_d N_A_1006_47#_c_920_n N_A_1006_47#_c_923_n
+ N_A_1006_47#_c_918_n PM_SKY130_FD_SC_LP__A211O_4%A_1006_47#
cc_1 VNB N_A_103_263#_M1001_g 5.01157e-19 $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=2.465
cc_2 VNB N_A_103_263#_M1006_g 4.57539e-19 $X=-0.19 $Y=-0.245 $X2=1.02 $Y2=2.465
cc_3 VNB N_A_103_263#_M1007_g 0.0282473f $X=-0.19 $Y=-0.245 $X2=1.145 $Y2=0.655
cc_4 VNB N_A_103_263#_M1014_g 4.57707e-19 $X=-0.19 $Y=-0.245 $X2=1.45 $Y2=2.465
cc_5 VNB N_A_103_263#_M1008_g 0.0213292f $X=-0.19 $Y=-0.245 $X2=1.575 $Y2=0.655
cc_6 VNB N_A_103_263#_M1021_g 5.58168e-19 $X=-0.19 $Y=-0.245 $X2=1.88 $Y2=2.465
cc_7 VNB N_A_103_263#_M1013_g 0.0215477f $X=-0.19 $Y=-0.245 $X2=2.005 $Y2=0.655
cc_8 VNB N_A_103_263#_M1023_g 0.0217747f $X=-0.19 $Y=-0.245 $X2=2.45 $Y2=0.655
cc_9 VNB N_A_103_263#_c_123_n 0.00176541f $X=-0.19 $Y=-0.245 $X2=2.475 $Y2=1.49
cc_10 VNB N_A_103_263#_c_124_n 0.00208789f $X=-0.19 $Y=-0.245 $X2=2.56 $Y2=1.395
cc_11 VNB N_A_103_263#_c_125_n 5.33145e-19 $X=-0.19 $Y=-0.245 $X2=2.56 $Y2=2.035
cc_12 VNB N_A_103_263#_c_126_n 0.00416957f $X=-0.19 $Y=-0.245 $X2=3 $Y2=1.07
cc_13 VNB N_A_103_263#_c_127_n 0.0271349f $X=-0.19 $Y=-0.245 $X2=5.505 $Y2=1.15
cc_14 VNB N_A_103_263#_c_128_n 0.00113298f $X=-0.19 $Y=-0.245 $X2=2.56 $Y2=1.49
cc_15 VNB N_A_103_263#_c_129_n 0.0026419f $X=-0.19 $Y=-0.245 $X2=3.095 $Y2=0.93
cc_16 VNB N_A_103_263#_c_130_n 0.00462043f $X=-0.19 $Y=-0.245 $X2=3.97 $Y2=0.93
cc_17 VNB N_A_103_263#_c_131_n 0.132907f $X=-0.19 $Y=-0.245 $X2=2.45 $Y2=1.48
cc_18 VNB N_B1_M1002_g 0.0243938f $X=-0.19 $Y=-0.245 $X2=5.46 $Y2=0.235
cc_19 VNB N_B1_M1016_g 0.0267011f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_B1_c_283_n 0.0285324f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.645
cc_21 VNB N_B1_c_284_n 0.0243819f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_B1_c_285_n 0.00485426f $X=-0.19 $Y=-0.245 $X2=1.575 $Y2=1.315
cc_23 VNB N_C1_c_381_n 0.0144921f $X=-0.19 $Y=-0.245 $X2=2.955 $Y2=0.235
cc_24 VNB N_C1_M1000_g 0.00718504f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_C1_c_383_n 0.0143761f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_C1_M1010_g 0.00689411f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.645
cc_27 VNB C1 9.45698e-19 $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=2.465
cc_28 VNB N_C1_c_386_n 0.0464291f $X=-0.19 $Y=-0.245 $X2=1.145 $Y2=0.655
cc_29 VNB N_A2_M1012_g 0.0273285f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A2_M1017_g 0.0348112f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A2_c_440_n 0.0191683f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A2_c_441_n 0.0298578f $X=-0.19 $Y=-0.245 $X2=1.145 $Y2=1.315
cc_33 VNB A2 0.00339782f $X=-0.19 $Y=-0.245 $X2=1.145 $Y2=0.655
cc_34 VNB A2 7.81979e-19 $X=-0.19 $Y=-0.245 $X2=1.45 $Y2=1.645
cc_35 VNB N_A2_c_444_n 0.0241109f $X=-0.19 $Y=-0.245 $X2=1.88 $Y2=1.645
cc_36 VNB N_A1_M1009_g 0.0232219f $X=-0.19 $Y=-0.245 $X2=5.46 $Y2=0.235
cc_37 VNB N_A1_M1020_g 0.0246694f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A1_c_516_n 0.0326901f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_VPWR_c_563_n 0.283096f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_X_c_666_n 0.0205973f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=2.465
cc_41 VNB N_X_c_667_n 0.00541042f $X=-0.19 $Y=-0.245 $X2=1.575 $Y2=1.315
cc_42 VNB N_X_c_668_n 0.00144145f $X=-0.19 $Y=-0.245 $X2=2.45 $Y2=0.655
cc_43 VNB X 0.0429221f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB X 0.00966496f $X=-0.19 $Y=-0.245 $X2=0.68 $Y2=1.49
cc_45 VNB X 0.025245f $X=-0.19 $Y=-0.245 $X2=3.102 $Y2=0.845
cc_46 VNB N_VGND_c_817_n 0.0157139f $X=-0.19 $Y=-0.245 $X2=1.145 $Y2=1.315
cc_47 VNB N_VGND_c_818_n 0.0129398f $X=-0.19 $Y=-0.245 $X2=1.145 $Y2=0.655
cc_48 VNB N_VGND_c_819_n 3.11777e-19 $X=-0.19 $Y=-0.245 $X2=1.45 $Y2=2.465
cc_49 VNB N_VGND_c_820_n 3.14445e-19 $X=-0.19 $Y=-0.245 $X2=1.575 $Y2=0.655
cc_50 VNB N_VGND_c_821_n 3.19546e-19 $X=-0.19 $Y=-0.245 $X2=1.88 $Y2=2.465
cc_51 VNB N_VGND_c_822_n 0.00617402f $X=-0.19 $Y=-0.245 $X2=2.005 $Y2=0.655
cc_52 VNB N_VGND_c_823_n 0.0102287f $X=-0.19 $Y=-0.245 $X2=2.45 $Y2=1.315
cc_53 VNB N_VGND_c_824_n 0.0436121f $X=-0.19 $Y=-0.245 $X2=2.45 $Y2=0.655
cc_54 VNB N_VGND_c_825_n 0.0242265f $X=-0.19 $Y=-0.245 $X2=2.475 $Y2=1.49
cc_55 VNB N_VGND_c_826_n 0.00513431f $X=-0.19 $Y=-0.245 $X2=0.68 $Y2=1.49
cc_56 VNB N_VGND_c_827_n 0.0135112f $X=-0.19 $Y=-0.245 $X2=2.56 $Y2=1.155
cc_57 VNB N_VGND_c_828_n 0.013276f $X=-0.19 $Y=-0.245 $X2=2.645 $Y2=1.07
cc_58 VNB N_VGND_c_829_n 0.0149824f $X=-0.19 $Y=-0.245 $X2=3.095 $Y2=0.42
cc_59 VNB N_VGND_c_830_n 0.0369363f $X=-0.19 $Y=-0.245 $X2=3.992 $Y2=0.42
cc_60 VNB N_VGND_c_831_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=2.56 $Y2=1.49
cc_61 VNB N_VGND_c_832_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=3.102 $Y2=1.07
cc_62 VNB N_VGND_c_833_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=3.62 $Y2=2.15
cc_63 VNB N_VGND_c_834_n 0.0106716f $X=-0.19 $Y=-0.245 $X2=3.992 $Y2=0.93
cc_64 VNB N_VGND_c_835_n 0.344736f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_A_1006_47#_c_918_n 0.00377124f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VPB N_A_103_263#_M1001_g 0.0225572f $X=-0.19 $Y=1.655 $X2=0.59 $Y2=2.465
cc_67 VPB N_A_103_263#_M1006_g 0.0188947f $X=-0.19 $Y=1.655 $X2=1.02 $Y2=2.465
cc_68 VPB N_A_103_263#_M1014_g 0.018914f $X=-0.19 $Y=1.655 $X2=1.45 $Y2=2.465
cc_69 VPB N_A_103_263#_M1021_g 0.0235499f $X=-0.19 $Y=1.655 $X2=1.88 $Y2=2.465
cc_70 VPB N_A_103_263#_c_125_n 0.0061487f $X=-0.19 $Y=1.655 $X2=2.56 $Y2=2.035
cc_71 VPB N_A_103_263#_c_137_n 0.00758484f $X=-0.19 $Y=1.655 $X2=2.645 $Y2=2.12
cc_72 VPB N_B1_M1015_g 0.0225139f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_73 VPB N_B1_c_283_n 0.00581045f $X=-0.19 $Y=1.655 $X2=0.59 $Y2=1.645
cc_74 VPB N_B1_M1022_g 0.0195668f $X=-0.19 $Y=1.655 $X2=0.59 $Y2=2.465
cc_75 VPB N_B1_c_289_n 0.00201358f $X=-0.19 $Y=1.655 $X2=1.02 $Y2=2.465
cc_76 VPB N_B1_c_290_n 0.00935624f $X=-0.19 $Y=1.655 $X2=1.145 $Y2=0.655
cc_77 VPB N_B1_c_284_n 0.00650746f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_78 VPB N_B1_c_285_n 0.00217978f $X=-0.19 $Y=1.655 $X2=1.575 $Y2=1.315
cc_79 VPB N_C1_M1000_g 0.0187202f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_80 VPB N_C1_M1010_g 0.0191658f $X=-0.19 $Y=1.655 $X2=0.59 $Y2=1.645
cc_81 VPB N_A2_M1018_g 0.0257297f $X=-0.19 $Y=1.655 $X2=0.59 $Y2=2.465
cc_82 VPB N_A2_c_441_n 0.00638499f $X=-0.19 $Y=1.655 $X2=1.145 $Y2=1.315
cc_83 VPB A2 0.00279787f $X=-0.19 $Y=1.655 $X2=1.145 $Y2=0.655
cc_84 VPB A2 0.0032815f $X=-0.19 $Y=1.655 $X2=1.45 $Y2=1.645
cc_85 VPB N_A2_c_444_n 0.00948774f $X=-0.19 $Y=1.655 $X2=1.88 $Y2=1.645
cc_86 VPB N_A2_c_450_n 0.0171125f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_87 VPB N_A1_M1003_g 0.0193842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_88 VPB N_A1_M1011_g 0.018741f $X=-0.19 $Y=1.655 $X2=0.59 $Y2=2.465
cc_89 VPB N_A1_c_519_n 0.00239041f $X=-0.19 $Y=1.655 $X2=1.145 $Y2=0.655
cc_90 VPB N_A1_c_516_n 0.00478891f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_91 VPB N_VPWR_c_564_n 0.0140081f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_92 VPB N_VPWR_c_565_n 0.0415885f $X=-0.19 $Y=1.655 $X2=1.02 $Y2=2.465
cc_93 VPB N_VPWR_c_566_n 3.0911e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_94 VPB N_VPWR_c_567_n 0.0197947f $X=-0.19 $Y=1.655 $X2=1.575 $Y2=0.655
cc_95 VPB N_VPWR_c_568_n 0.00227979f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_96 VPB N_VPWR_c_569_n 4.16958e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_97 VPB N_VPWR_c_570_n 0.0129398f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_98 VPB N_VPWR_c_571_n 0.0129398f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_99 VPB N_VPWR_c_572_n 0.0651247f $X=-0.19 $Y=1.655 $X2=2.56 $Y2=1.395
cc_100 VPB N_VPWR_c_573_n 0.016701f $X=-0.19 $Y=1.655 $X2=3.102 $Y2=0.42
cc_101 VPB N_VPWR_c_574_n 0.0153759f $X=-0.19 $Y=1.655 $X2=3.97 $Y2=0.42
cc_102 VPB N_VPWR_c_563_n 0.0636775f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_103 VPB N_VPWR_c_576_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_104 VPB N_VPWR_c_577_n 0.00510842f $X=-0.19 $Y=1.655 $X2=3.095 $Y2=0.93
cc_105 VPB N_VPWR_c_578_n 0.00510842f $X=-0.19 $Y=1.655 $X2=3.62 $Y2=2.145
cc_106 VPB N_VPWR_c_579_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_107 VPB N_X_c_672_n 0.0026141f $X=-0.19 $Y=1.655 $X2=0.59 $Y2=1.645
cc_108 VPB N_X_c_673_n 0.013434f $X=-0.19 $Y=1.655 $X2=0.59 $Y2=2.465
cc_109 VPB N_X_c_674_n 0.00537118f $X=-0.19 $Y=1.655 $X2=1.145 $Y2=0.655
cc_110 VPB N_X_c_675_n 0.00144499f $X=-0.19 $Y=1.655 $X2=2.45 $Y2=0.655
cc_111 VPB X 0.00546699f $X=-0.19 $Y=1.655 $X2=3.102 $Y2=0.845
cc_112 VPB N_A_527_367#_c_730_n 0.0245119f $X=-0.19 $Y=1.655 $X2=1.575 $Y2=0.655
cc_113 VPB N_A_527_367#_c_731_n 0.00854714f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_114 VPB N_A_527_367#_c_732_n 0.0305687f $X=-0.19 $Y=1.655 $X2=2.45 $Y2=0.655
cc_115 N_A_103_263#_M1023_g N_B1_M1002_g 0.0243197f $X=2.45 $Y=0.655 $X2=0 $Y2=0
cc_116 N_A_103_263#_c_124_n N_B1_M1002_g 0.00395652f $X=2.56 $Y=1.395 $X2=0
+ $Y2=0
cc_117 N_A_103_263#_c_126_n N_B1_M1002_g 0.0130324f $X=3 $Y=1.07 $X2=0 $Y2=0
cc_118 N_A_103_263#_c_125_n N_B1_M1015_g 0.00638055f $X=2.56 $Y=2.035 $X2=0
+ $Y2=0
cc_119 N_A_103_263#_c_142_p N_B1_M1015_g 2.39364e-19 $X=3.62 $Y=2.15 $X2=0 $Y2=0
cc_120 N_A_103_263#_c_143_p N_B1_M1015_g 0.0123401f $X=3.455 $Y=2.145 $X2=0
+ $Y2=0
cc_121 N_A_103_263#_c_127_n N_B1_M1016_g 0.0143444f $X=5.505 $Y=1.15 $X2=0 $Y2=0
cc_122 N_A_103_263#_c_130_n N_B1_M1016_g 0.00143368f $X=3.97 $Y=0.93 $X2=0 $Y2=0
cc_123 N_A_103_263#_c_127_n N_B1_c_283_n 0.00517679f $X=5.505 $Y=1.15 $X2=0
+ $Y2=0
cc_124 N_A_103_263#_c_142_p N_B1_M1022_g 6.58072e-19 $X=3.62 $Y=2.15 $X2=0 $Y2=0
cc_125 N_A_103_263#_c_127_n N_B1_c_289_n 0.0237676f $X=5.505 $Y=1.15 $X2=0 $Y2=0
cc_126 N_A_103_263#_M1000_s N_B1_c_290_n 0.00176891f $X=3.48 $Y=1.835 $X2=0
+ $Y2=0
cc_127 N_A_103_263#_c_127_n N_B1_c_290_n 3.24709e-19 $X=5.505 $Y=1.15 $X2=0
+ $Y2=0
cc_128 N_A_103_263#_c_143_p N_B1_c_290_n 0.0290594f $X=3.455 $Y=2.145 $X2=0
+ $Y2=0
cc_129 N_A_103_263#_c_130_n N_B1_c_290_n 0.00942786f $X=3.97 $Y=0.93 $X2=0 $Y2=0
cc_130 N_A_103_263#_c_124_n N_B1_c_284_n 3.07481e-19 $X=2.56 $Y=1.395 $X2=0
+ $Y2=0
cc_131 N_A_103_263#_c_125_n N_B1_c_284_n 0.00110891f $X=2.56 $Y=2.035 $X2=0
+ $Y2=0
cc_132 N_A_103_263#_c_126_n N_B1_c_284_n 0.00287925f $X=3 $Y=1.07 $X2=0 $Y2=0
cc_133 N_A_103_263#_c_128_n N_B1_c_284_n 0.00137052f $X=2.56 $Y=1.49 $X2=0 $Y2=0
cc_134 N_A_103_263#_c_129_n N_B1_c_284_n 4.95034e-19 $X=3.095 $Y=0.93 $X2=0
+ $Y2=0
cc_135 N_A_103_263#_c_143_p N_B1_c_284_n 0.00280793f $X=3.455 $Y=2.145 $X2=0
+ $Y2=0
cc_136 N_A_103_263#_c_131_n N_B1_c_284_n 0.0186521f $X=2.45 $Y=1.48 $X2=0 $Y2=0
cc_137 N_A_103_263#_c_124_n N_B1_c_285_n 0.0037684f $X=2.56 $Y=1.395 $X2=0 $Y2=0
cc_138 N_A_103_263#_c_125_n N_B1_c_285_n 0.0219909f $X=2.56 $Y=2.035 $X2=0 $Y2=0
cc_139 N_A_103_263#_c_126_n N_B1_c_285_n 0.0127021f $X=3 $Y=1.07 $X2=0 $Y2=0
cc_140 N_A_103_263#_c_128_n N_B1_c_285_n 0.016207f $X=2.56 $Y=1.49 $X2=0 $Y2=0
cc_141 N_A_103_263#_c_129_n N_B1_c_285_n 0.0169397f $X=3.095 $Y=0.93 $X2=0 $Y2=0
cc_142 N_A_103_263#_c_143_p N_B1_c_285_n 0.0210449f $X=3.455 $Y=2.145 $X2=0
+ $Y2=0
cc_143 N_A_103_263#_c_131_n N_B1_c_285_n 2.63286e-19 $X=2.45 $Y=1.48 $X2=0 $Y2=0
cc_144 N_A_103_263#_c_167_p N_C1_c_381_n 0.0132682f $X=3.875 $Y=0.93 $X2=-0.19
+ $Y2=-0.245
cc_145 N_A_103_263#_c_129_n N_C1_c_381_n 0.00200282f $X=3.095 $Y=0.93 $X2=-0.19
+ $Y2=-0.245
cc_146 N_A_103_263#_c_142_p N_C1_M1000_g 0.0019458f $X=3.62 $Y=2.15 $X2=0 $Y2=0
cc_147 N_A_103_263#_c_143_p N_C1_M1000_g 0.00756348f $X=3.455 $Y=2.145 $X2=0
+ $Y2=0
cc_148 N_A_103_263#_c_167_p N_C1_c_383_n 0.0133671f $X=3.875 $Y=0.93 $X2=0 $Y2=0
cc_149 N_A_103_263#_c_130_n N_C1_c_383_n 0.00398777f $X=3.97 $Y=0.93 $X2=0 $Y2=0
cc_150 N_A_103_263#_c_142_p N_C1_M1010_g 0.00466225f $X=3.62 $Y=2.15 $X2=0 $Y2=0
cc_151 N_A_103_263#_c_167_p C1 0.0204255f $X=3.875 $Y=0.93 $X2=0 $Y2=0
cc_152 N_A_103_263#_c_130_n C1 0.0041291f $X=3.97 $Y=0.93 $X2=0 $Y2=0
cc_153 N_A_103_263#_c_167_p N_C1_c_386_n 0.00267212f $X=3.875 $Y=0.93 $X2=0
+ $Y2=0
cc_154 N_A_103_263#_c_130_n N_C1_c_386_n 7.62829e-19 $X=3.97 $Y=0.93 $X2=0 $Y2=0
cc_155 N_A_103_263#_c_127_n N_A2_M1012_g 0.0156975f $X=5.505 $Y=1.15 $X2=0 $Y2=0
cc_156 N_A_103_263#_c_127_n A2 0.0232932f $X=5.505 $Y=1.15 $X2=0 $Y2=0
cc_157 N_A_103_263#_c_127_n N_A2_c_444_n 0.00488923f $X=5.505 $Y=1.15 $X2=0
+ $Y2=0
cc_158 N_A_103_263#_c_127_n N_A1_M1009_g 0.0118992f $X=5.505 $Y=1.15 $X2=0 $Y2=0
cc_159 N_A_103_263#_c_127_n N_A1_M1020_g 0.00468911f $X=5.505 $Y=1.15 $X2=0
+ $Y2=0
cc_160 N_A_103_263#_c_127_n N_A1_c_519_n 0.0233837f $X=5.505 $Y=1.15 $X2=0 $Y2=0
cc_161 N_A_103_263#_c_127_n N_A1_c_516_n 0.00276639f $X=5.505 $Y=1.15 $X2=0
+ $Y2=0
cc_162 N_A_103_263#_M1001_g N_VPWR_c_565_n 0.0152824f $X=0.59 $Y=2.465 $X2=0
+ $Y2=0
cc_163 N_A_103_263#_M1006_g N_VPWR_c_565_n 7.27171e-19 $X=1.02 $Y=2.465 $X2=0
+ $Y2=0
cc_164 N_A_103_263#_M1001_g N_VPWR_c_566_n 7.24342e-19 $X=0.59 $Y=2.465 $X2=0
+ $Y2=0
cc_165 N_A_103_263#_M1006_g N_VPWR_c_566_n 0.0141279f $X=1.02 $Y=2.465 $X2=0
+ $Y2=0
cc_166 N_A_103_263#_M1014_g N_VPWR_c_566_n 0.0141279f $X=1.45 $Y=2.465 $X2=0
+ $Y2=0
cc_167 N_A_103_263#_M1021_g N_VPWR_c_566_n 7.24342e-19 $X=1.88 $Y=2.465 $X2=0
+ $Y2=0
cc_168 N_A_103_263#_M1014_g N_VPWR_c_567_n 8.15296e-19 $X=1.45 $Y=2.465 $X2=0
+ $Y2=0
cc_169 N_A_103_263#_M1021_g N_VPWR_c_567_n 0.0224158f $X=1.88 $Y=2.465 $X2=0
+ $Y2=0
cc_170 N_A_103_263#_c_123_n N_VPWR_c_567_n 0.0211642f $X=2.475 $Y=1.49 $X2=0
+ $Y2=0
cc_171 N_A_103_263#_c_125_n N_VPWR_c_567_n 0.0147661f $X=2.56 $Y=2.035 $X2=0
+ $Y2=0
cc_172 N_A_103_263#_c_137_n N_VPWR_c_567_n 0.0127464f $X=2.645 $Y=2.12 $X2=0
+ $Y2=0
cc_173 N_A_103_263#_c_131_n N_VPWR_c_567_n 0.00822646f $X=2.45 $Y=1.48 $X2=0
+ $Y2=0
cc_174 N_A_103_263#_M1001_g N_VPWR_c_570_n 0.00486043f $X=0.59 $Y=2.465 $X2=0
+ $Y2=0
cc_175 N_A_103_263#_M1006_g N_VPWR_c_570_n 0.00486043f $X=1.02 $Y=2.465 $X2=0
+ $Y2=0
cc_176 N_A_103_263#_M1014_g N_VPWR_c_571_n 0.00486043f $X=1.45 $Y=2.465 $X2=0
+ $Y2=0
cc_177 N_A_103_263#_M1021_g N_VPWR_c_571_n 0.00486043f $X=1.88 $Y=2.465 $X2=0
+ $Y2=0
cc_178 N_A_103_263#_M1000_s N_VPWR_c_563_n 0.00225919f $X=3.48 $Y=1.835 $X2=0
+ $Y2=0
cc_179 N_A_103_263#_M1001_g N_VPWR_c_563_n 0.00824727f $X=0.59 $Y=2.465 $X2=0
+ $Y2=0
cc_180 N_A_103_263#_M1006_g N_VPWR_c_563_n 0.00824727f $X=1.02 $Y=2.465 $X2=0
+ $Y2=0
cc_181 N_A_103_263#_M1014_g N_VPWR_c_563_n 0.00824727f $X=1.45 $Y=2.465 $X2=0
+ $Y2=0
cc_182 N_A_103_263#_M1021_g N_VPWR_c_563_n 0.00824727f $X=1.88 $Y=2.465 $X2=0
+ $Y2=0
cc_183 N_A_103_263#_M1001_g N_X_c_672_n 0.0148644f $X=0.59 $Y=2.465 $X2=0 $Y2=0
cc_184 N_A_103_263#_c_123_n N_X_c_672_n 0.0134628f $X=2.475 $Y=1.49 $X2=0 $Y2=0
cc_185 N_A_103_263#_M1007_g N_X_c_666_n 0.0160954f $X=1.145 $Y=0.655 $X2=0 $Y2=0
cc_186 N_A_103_263#_c_123_n N_X_c_666_n 0.0534793f $X=2.475 $Y=1.49 $X2=0 $Y2=0
cc_187 N_A_103_263#_c_131_n N_X_c_666_n 0.0156348f $X=2.45 $Y=1.48 $X2=0 $Y2=0
cc_188 N_A_103_263#_M1006_g N_X_c_674_n 0.0131755f $X=1.02 $Y=2.465 $X2=0 $Y2=0
cc_189 N_A_103_263#_M1014_g N_X_c_674_n 0.0130133f $X=1.45 $Y=2.465 $X2=0 $Y2=0
cc_190 N_A_103_263#_M1021_g N_X_c_674_n 0.00208318f $X=1.88 $Y=2.465 $X2=0 $Y2=0
cc_191 N_A_103_263#_c_123_n N_X_c_674_n 0.0625613f $X=2.475 $Y=1.49 $X2=0 $Y2=0
cc_192 N_A_103_263#_c_131_n N_X_c_674_n 0.00575333f $X=2.45 $Y=1.48 $X2=0 $Y2=0
cc_193 N_A_103_263#_M1008_g N_X_c_667_n 0.014308f $X=1.575 $Y=0.655 $X2=0 $Y2=0
cc_194 N_A_103_263#_M1013_g N_X_c_667_n 0.0139541f $X=2.005 $Y=0.655 $X2=0 $Y2=0
cc_195 N_A_103_263#_M1023_g N_X_c_667_n 0.00131302f $X=2.45 $Y=0.655 $X2=0 $Y2=0
cc_196 N_A_103_263#_c_123_n N_X_c_667_n 0.0619584f $X=2.475 $Y=1.49 $X2=0 $Y2=0
cc_197 N_A_103_263#_c_124_n N_X_c_667_n 0.00561303f $X=2.56 $Y=1.395 $X2=0 $Y2=0
cc_198 N_A_103_263#_c_221_p N_X_c_667_n 0.00957547f $X=2.645 $Y=1.07 $X2=0 $Y2=0
cc_199 N_A_103_263#_c_131_n N_X_c_667_n 0.00585069f $X=2.45 $Y=1.48 $X2=0 $Y2=0
cc_200 N_A_103_263#_M1023_g N_X_c_694_n 0.00589948f $X=2.45 $Y=0.655 $X2=0 $Y2=0
cc_201 N_A_103_263#_c_221_p N_X_c_694_n 0.00460201f $X=2.645 $Y=1.07 $X2=0 $Y2=0
cc_202 N_A_103_263#_c_123_n N_X_c_675_n 0.0154427f $X=2.475 $Y=1.49 $X2=0 $Y2=0
cc_203 N_A_103_263#_c_131_n N_X_c_675_n 0.00250529f $X=2.45 $Y=1.48 $X2=0 $Y2=0
cc_204 N_A_103_263#_c_123_n N_X_c_668_n 0.0154425f $X=2.475 $Y=1.49 $X2=0 $Y2=0
cc_205 N_A_103_263#_c_131_n N_X_c_668_n 0.00299787f $X=2.45 $Y=1.48 $X2=0 $Y2=0
cc_206 N_A_103_263#_M1007_g X 0.00376785f $X=1.145 $Y=0.655 $X2=0 $Y2=0
cc_207 N_A_103_263#_c_123_n X 0.0154753f $X=2.475 $Y=1.49 $X2=0 $Y2=0
cc_208 N_A_103_263#_c_131_n X 0.0113995f $X=2.45 $Y=1.48 $X2=0 $Y2=0
cc_209 N_A_103_263#_c_125_n N_A_527_367#_M1015_s 0.00243147f $X=2.56 $Y=2.035
+ $X2=-0.19 $Y2=-0.245
cc_210 N_A_103_263#_c_143_p N_A_527_367#_M1015_s 0.00752032f $X=3.455 $Y=2.145
+ $X2=-0.19 $Y2=-0.245
cc_211 N_A_103_263#_M1000_s N_A_527_367#_c_735_n 0.00349583f $X=3.48 $Y=1.835
+ $X2=0 $Y2=0
cc_212 N_A_103_263#_c_142_p N_A_527_367#_c_735_n 0.0156817f $X=3.62 $Y=2.15
+ $X2=0 $Y2=0
cc_213 N_A_103_263#_c_143_p N_A_527_367#_c_735_n 0.0236386f $X=3.455 $Y=2.145
+ $X2=0 $Y2=0
cc_214 N_A_103_263#_c_142_p N_A_527_367#_c_738_n 0.00639668f $X=3.62 $Y=2.15
+ $X2=0 $Y2=0
cc_215 N_A_103_263#_M1021_g N_A_527_367#_c_731_n 0.00111119f $X=1.88 $Y=2.465
+ $X2=0 $Y2=0
cc_216 N_A_103_263#_c_137_n N_A_527_367#_c_731_n 0.00461436f $X=2.645 $Y=2.12
+ $X2=0 $Y2=0
cc_217 N_A_103_263#_c_143_p N_A_527_367#_c_731_n 0.0178135f $X=3.455 $Y=2.145
+ $X2=0 $Y2=0
cc_218 N_A_103_263#_c_143_p N_A_610_367#_M1015_d 0.00372302f $X=3.455 $Y=2.145
+ $X2=-0.19 $Y2=-0.245
cc_219 N_A_103_263#_M1000_s N_A_610_367#_c_802_n 0.00345347f $X=3.48 $Y=1.835
+ $X2=0 $Y2=0
cc_220 N_A_103_263#_c_126_n N_VGND_M1023_s 0.00111061f $X=3 $Y=1.07 $X2=0 $Y2=0
cc_221 N_A_103_263#_c_221_p N_VGND_M1023_s 7.14262e-19 $X=2.645 $Y=1.07 $X2=0
+ $Y2=0
cc_222 N_A_103_263#_c_167_p N_VGND_M1004_d 0.0032689f $X=3.875 $Y=0.93 $X2=0
+ $Y2=0
cc_223 N_A_103_263#_c_127_n N_VGND_M1016_d 0.005639f $X=5.505 $Y=1.15 $X2=0
+ $Y2=0
cc_224 N_A_103_263#_M1007_g N_VGND_c_817_n 0.0122528f $X=1.145 $Y=0.655 $X2=0
+ $Y2=0
cc_225 N_A_103_263#_M1008_g N_VGND_c_817_n 6.28154e-19 $X=1.575 $Y=0.655 $X2=0
+ $Y2=0
cc_226 N_A_103_263#_M1007_g N_VGND_c_818_n 0.00486043f $X=1.145 $Y=0.655 $X2=0
+ $Y2=0
cc_227 N_A_103_263#_M1008_g N_VGND_c_818_n 0.00486043f $X=1.575 $Y=0.655 $X2=0
+ $Y2=0
cc_228 N_A_103_263#_M1007_g N_VGND_c_819_n 6.25324e-19 $X=1.145 $Y=0.655 $X2=0
+ $Y2=0
cc_229 N_A_103_263#_M1008_g N_VGND_c_819_n 0.0110025f $X=1.575 $Y=0.655 $X2=0
+ $Y2=0
cc_230 N_A_103_263#_M1013_g N_VGND_c_819_n 0.0110542f $X=2.005 $Y=0.655 $X2=0
+ $Y2=0
cc_231 N_A_103_263#_M1023_g N_VGND_c_819_n 6.16843e-19 $X=2.45 $Y=0.655 $X2=0
+ $Y2=0
cc_232 N_A_103_263#_M1013_g N_VGND_c_820_n 6.18223e-19 $X=2.005 $Y=0.655 $X2=0
+ $Y2=0
cc_233 N_A_103_263#_M1023_g N_VGND_c_820_n 0.0102149f $X=2.45 $Y=0.655 $X2=0
+ $Y2=0
cc_234 N_A_103_263#_c_126_n N_VGND_c_820_n 0.00969985f $X=3 $Y=1.07 $X2=0 $Y2=0
cc_235 N_A_103_263#_c_221_p N_VGND_c_820_n 0.00734015f $X=2.645 $Y=1.07 $X2=0
+ $Y2=0
cc_236 N_A_103_263#_c_167_p N_VGND_c_821_n 0.016709f $X=3.875 $Y=0.93 $X2=0
+ $Y2=0
cc_237 N_A_103_263#_c_127_n N_VGND_c_822_n 0.0394444f $X=5.505 $Y=1.15 $X2=0
+ $Y2=0
cc_238 N_A_103_263#_M1013_g N_VGND_c_827_n 0.00486043f $X=2.005 $Y=0.655 $X2=0
+ $Y2=0
cc_239 N_A_103_263#_M1023_g N_VGND_c_827_n 0.00486043f $X=2.45 $Y=0.655 $X2=0
+ $Y2=0
cc_240 N_A_103_263#_c_263_p N_VGND_c_828_n 0.0135072f $X=3.095 $Y=0.42 $X2=0
+ $Y2=0
cc_241 N_A_103_263#_c_264_p N_VGND_c_829_n 0.0140491f $X=3.97 $Y=0.42 $X2=0
+ $Y2=0
cc_242 N_A_103_263#_M1002_s N_VGND_c_835_n 0.00420875f $X=2.955 $Y=0.235 $X2=0
+ $Y2=0
cc_243 N_A_103_263#_M1019_s N_VGND_c_835_n 0.00252268f $X=3.83 $Y=0.235 $X2=0
+ $Y2=0
cc_244 N_A_103_263#_M1009_s N_VGND_c_835_n 0.00225186f $X=5.46 $Y=0.235 $X2=0
+ $Y2=0
cc_245 N_A_103_263#_M1007_g N_VGND_c_835_n 0.00824727f $X=1.145 $Y=0.655 $X2=0
+ $Y2=0
cc_246 N_A_103_263#_M1008_g N_VGND_c_835_n 0.00824727f $X=1.575 $Y=0.655 $X2=0
+ $Y2=0
cc_247 N_A_103_263#_M1013_g N_VGND_c_835_n 0.0082859f $X=2.005 $Y=0.655 $X2=0
+ $Y2=0
cc_248 N_A_103_263#_M1023_g N_VGND_c_835_n 0.0082859f $X=2.45 $Y=0.655 $X2=0
+ $Y2=0
cc_249 N_A_103_263#_c_263_p N_VGND_c_835_n 0.00789217f $X=3.095 $Y=0.42 $X2=0
+ $Y2=0
cc_250 N_A_103_263#_c_167_p N_VGND_c_835_n 0.0108383f $X=3.875 $Y=0.93 $X2=0
+ $Y2=0
cc_251 N_A_103_263#_c_264_p N_VGND_c_835_n 0.0090585f $X=3.97 $Y=0.42 $X2=0
+ $Y2=0
cc_252 N_A_103_263#_c_127_n N_A_1006_47#_M1012_d 0.00176461f $X=5.505 $Y=1.15
+ $X2=-0.19 $Y2=-0.245
cc_253 N_A_103_263#_M1009_s N_A_1006_47#_c_920_n 0.00332344f $X=5.46 $Y=0.235
+ $X2=0 $Y2=0
cc_254 N_A_103_263#_c_127_n N_A_1006_47#_c_920_n 0.00280043f $X=5.505 $Y=1.15
+ $X2=0 $Y2=0
cc_255 N_A_103_263#_c_278_p N_A_1006_47#_c_920_n 0.0125759f $X=5.6 $Y=0.76 $X2=0
+ $Y2=0
cc_256 N_A_103_263#_c_127_n N_A_1006_47#_c_923_n 0.0169932f $X=5.505 $Y=1.15
+ $X2=0 $Y2=0
cc_257 N_A_103_263#_c_127_n N_A_1006_47#_c_918_n 0.00201679f $X=5.505 $Y=1.15
+ $X2=0 $Y2=0
cc_258 N_B1_M1002_g N_C1_c_381_n 0.0169646f $X=2.88 $Y=0.655 $X2=-0.19
+ $Y2=-0.245
cc_259 N_B1_M1015_g N_C1_M1000_g 0.0542405f $X=2.975 $Y=2.465 $X2=0 $Y2=0
cc_260 N_B1_c_290_n N_C1_M1000_g 0.0110226f $X=4.12 $Y=1.78 $X2=0 $Y2=0
cc_261 N_B1_c_284_n N_C1_M1000_g 0.00694594f $X=2.9 $Y=1.51 $X2=0 $Y2=0
cc_262 N_B1_c_285_n N_C1_M1000_g 0.004825f $X=2.9 $Y=1.51 $X2=0 $Y2=0
cc_263 N_B1_M1016_g N_C1_c_383_n 0.0124779f $X=4.185 $Y=0.655 $X2=0 $Y2=0
cc_264 N_B1_M1022_g N_C1_M1010_g 0.0459953f $X=4.305 $Y=2.465 $X2=0 $Y2=0
cc_265 N_B1_c_289_n N_C1_M1010_g 8.68178e-19 $X=4.285 $Y=1.5 $X2=0 $Y2=0
cc_266 N_B1_c_290_n N_C1_M1010_g 0.0153573f $X=4.12 $Y=1.78 $X2=0 $Y2=0
cc_267 N_B1_M1002_g C1 7.88883e-19 $X=2.88 $Y=0.655 $X2=0 $Y2=0
cc_268 N_B1_M1016_g C1 8.19068e-19 $X=4.185 $Y=0.655 $X2=0 $Y2=0
cc_269 N_B1_c_283_n C1 3.86588e-19 $X=4.305 $Y=1.665 $X2=0 $Y2=0
cc_270 N_B1_c_289_n C1 0.0036926f $X=4.285 $Y=1.5 $X2=0 $Y2=0
cc_271 N_B1_c_290_n C1 0.0236937f $X=4.12 $Y=1.78 $X2=0 $Y2=0
cc_272 N_B1_c_285_n C1 0.0136476f $X=2.9 $Y=1.51 $X2=0 $Y2=0
cc_273 N_B1_M1002_g N_C1_c_386_n 0.00421268f $X=2.88 $Y=0.655 $X2=0 $Y2=0
cc_274 N_B1_c_283_n N_C1_c_386_n 0.0307316f $X=4.305 $Y=1.665 $X2=0 $Y2=0
cc_275 N_B1_c_289_n N_C1_c_386_n 0.00144437f $X=4.285 $Y=1.5 $X2=0 $Y2=0
cc_276 N_B1_c_290_n N_C1_c_386_n 0.00372279f $X=4.12 $Y=1.78 $X2=0 $Y2=0
cc_277 N_B1_c_284_n N_C1_c_386_n 0.0109874f $X=2.9 $Y=1.51 $X2=0 $Y2=0
cc_278 N_B1_c_285_n N_C1_c_386_n 0.00129105f $X=2.9 $Y=1.51 $X2=0 $Y2=0
cc_279 N_B1_M1016_g N_A2_M1012_g 0.0106458f $X=4.185 $Y=0.655 $X2=0 $Y2=0
cc_280 N_B1_c_283_n N_A2_M1012_g 3.4974e-19 $X=4.305 $Y=1.665 $X2=0 $Y2=0
cc_281 N_B1_c_283_n A2 9.70956e-19 $X=4.305 $Y=1.665 $X2=0 $Y2=0
cc_282 N_B1_M1022_g A2 7.40806e-19 $X=4.305 $Y=2.465 $X2=0 $Y2=0
cc_283 N_B1_c_289_n A2 0.0201708f $X=4.285 $Y=1.5 $X2=0 $Y2=0
cc_284 N_B1_c_283_n N_A2_c_444_n 0.0129341f $X=4.305 $Y=1.665 $X2=0 $Y2=0
cc_285 N_B1_M1022_g N_A2_c_444_n 0.0263082f $X=4.305 $Y=2.465 $X2=0 $Y2=0
cc_286 N_B1_c_289_n N_A2_c_444_n 0.00101935f $X=4.285 $Y=1.5 $X2=0 $Y2=0
cc_287 N_B1_c_289_n N_A2_c_450_n 3.58185e-19 $X=4.285 $Y=1.5 $X2=0 $Y2=0
cc_288 N_B1_M1015_g N_VPWR_c_567_n 0.00714887f $X=2.975 $Y=2.465 $X2=0 $Y2=0
cc_289 N_B1_M1022_g N_VPWR_c_568_n 0.00103262f $X=4.305 $Y=2.465 $X2=0 $Y2=0
cc_290 N_B1_M1015_g N_VPWR_c_572_n 0.00426321f $X=2.975 $Y=2.465 $X2=0 $Y2=0
cc_291 N_B1_M1022_g N_VPWR_c_572_n 0.00439183f $X=4.305 $Y=2.465 $X2=0 $Y2=0
cc_292 N_B1_M1015_g N_VPWR_c_563_n 0.00737132f $X=2.975 $Y=2.465 $X2=0 $Y2=0
cc_293 N_B1_M1022_g N_VPWR_c_563_n 0.0065752f $X=4.305 $Y=2.465 $X2=0 $Y2=0
cc_294 N_B1_c_285_n N_A_527_367#_M1015_s 6.25038e-19 $X=2.9 $Y=1.51 $X2=-0.19
+ $Y2=-0.245
cc_295 N_B1_c_289_n N_A_527_367#_M1022_s 5.42701e-19 $X=4.285 $Y=1.5 $X2=0 $Y2=0
cc_296 N_B1_M1015_g N_A_527_367#_c_735_n 0.0087385f $X=2.975 $Y=2.465 $X2=0
+ $Y2=0
cc_297 N_B1_M1022_g N_A_527_367#_c_735_n 0.010579f $X=4.305 $Y=2.465 $X2=0 $Y2=0
cc_298 N_B1_c_289_n N_A_527_367#_c_735_n 0.00510868f $X=4.285 $Y=1.5 $X2=0 $Y2=0
cc_299 N_B1_c_290_n N_A_527_367#_c_735_n 0.0077539f $X=4.12 $Y=1.78 $X2=0 $Y2=0
cc_300 N_B1_c_283_n N_A_527_367#_c_738_n 2.2623e-19 $X=4.305 $Y=1.665 $X2=0
+ $Y2=0
cc_301 N_B1_M1022_g N_A_527_367#_c_738_n 0.0087874f $X=4.305 $Y=2.465 $X2=0
+ $Y2=0
cc_302 N_B1_c_289_n N_A_527_367#_c_738_n 0.00302975f $X=4.285 $Y=1.5 $X2=0 $Y2=0
cc_303 N_B1_M1015_g N_A_527_367#_c_731_n 0.00224658f $X=2.975 $Y=2.465 $X2=0
+ $Y2=0
cc_304 N_B1_c_290_n N_A_610_367#_M1015_d 7.94385e-19 $X=4.12 $Y=1.78 $X2=-0.19
+ $Y2=-0.245
cc_305 N_B1_c_285_n N_A_610_367#_M1015_d 0.00113653f $X=2.9 $Y=1.51 $X2=-0.19
+ $Y2=-0.245
cc_306 N_B1_c_289_n N_A_610_367#_M1010_d 0.00110246f $X=4.285 $Y=1.5 $X2=0 $Y2=0
cc_307 N_B1_c_290_n N_A_610_367#_M1010_d 0.00300496f $X=4.12 $Y=1.78 $X2=0 $Y2=0
cc_308 N_B1_M1015_g N_A_610_367#_c_802_n 0.00364494f $X=2.975 $Y=2.465 $X2=0
+ $Y2=0
cc_309 N_B1_M1002_g N_VGND_c_820_n 0.00989798f $X=2.88 $Y=0.655 $X2=0 $Y2=0
cc_310 N_B1_M1002_g N_VGND_c_821_n 5.62492e-19 $X=2.88 $Y=0.655 $X2=0 $Y2=0
cc_311 N_B1_M1016_g N_VGND_c_821_n 5.86967e-19 $X=4.185 $Y=0.655 $X2=0 $Y2=0
cc_312 N_B1_M1016_g N_VGND_c_822_n 0.002133f $X=4.185 $Y=0.655 $X2=0 $Y2=0
cc_313 N_B1_M1002_g N_VGND_c_828_n 0.00486043f $X=2.88 $Y=0.655 $X2=0 $Y2=0
cc_314 N_B1_M1016_g N_VGND_c_829_n 0.00585385f $X=4.185 $Y=0.655 $X2=0 $Y2=0
cc_315 N_B1_M1002_g N_VGND_c_835_n 0.00830854f $X=2.88 $Y=0.655 $X2=0 $Y2=0
cc_316 N_B1_M1016_g N_VGND_c_835_n 0.0112163f $X=4.185 $Y=0.655 $X2=0 $Y2=0
cc_317 N_C1_M1000_g N_VPWR_c_572_n 0.00362032f $X=3.405 $Y=2.465 $X2=0 $Y2=0
cc_318 N_C1_M1010_g N_VPWR_c_572_n 0.00362032f $X=3.835 $Y=2.465 $X2=0 $Y2=0
cc_319 N_C1_M1000_g N_VPWR_c_563_n 0.00544452f $X=3.405 $Y=2.465 $X2=0 $Y2=0
cc_320 N_C1_M1010_g N_VPWR_c_563_n 0.00554543f $X=3.835 $Y=2.465 $X2=0 $Y2=0
cc_321 N_C1_M1000_g N_A_527_367#_c_735_n 0.0106828f $X=3.405 $Y=2.465 $X2=0
+ $Y2=0
cc_322 N_C1_M1010_g N_A_527_367#_c_735_n 0.0122377f $X=3.835 $Y=2.465 $X2=0
+ $Y2=0
cc_323 N_C1_M1010_g N_A_527_367#_c_738_n 0.00147872f $X=3.835 $Y=2.465 $X2=0
+ $Y2=0
cc_324 N_C1_M1000_g N_A_527_367#_c_731_n 2.44249e-19 $X=3.405 $Y=2.465 $X2=0
+ $Y2=0
cc_325 N_C1_M1000_g N_A_610_367#_c_802_n 0.0109861f $X=3.405 $Y=2.465 $X2=0
+ $Y2=0
cc_326 N_C1_M1010_g N_A_610_367#_c_802_n 0.0109861f $X=3.835 $Y=2.465 $X2=0
+ $Y2=0
cc_327 N_C1_c_381_n N_VGND_c_820_n 5.9782e-19 $X=3.325 $Y=1.15 $X2=0 $Y2=0
cc_328 N_C1_c_381_n N_VGND_c_821_n 0.00982249f $X=3.325 $Y=1.15 $X2=0 $Y2=0
cc_329 N_C1_c_383_n N_VGND_c_821_n 0.00987906f $X=3.755 $Y=1.15 $X2=0 $Y2=0
cc_330 N_C1_c_381_n N_VGND_c_828_n 0.00486043f $X=3.325 $Y=1.15 $X2=0 $Y2=0
cc_331 N_C1_c_383_n N_VGND_c_829_n 0.00486043f $X=3.755 $Y=1.15 $X2=0 $Y2=0
cc_332 N_C1_c_381_n N_VGND_c_835_n 0.00461284f $X=3.325 $Y=1.15 $X2=0 $Y2=0
cc_333 N_C1_c_383_n N_VGND_c_835_n 0.0045769f $X=3.755 $Y=1.15 $X2=0 $Y2=0
cc_334 N_A2_M1012_g N_A1_M1009_g 0.0243456f $X=4.955 $Y=0.655 $X2=0 $Y2=0
cc_335 A2 N_A1_M1003_g 0.00411507f $X=4.955 $Y=1.95 $X2=0 $Y2=0
cc_336 A2 N_A1_M1003_g 0.0109315f $X=5.915 $Y=1.95 $X2=0 $Y2=0
cc_337 N_A2_c_450_n N_A1_M1003_g 0.0361806f $X=4.935 $Y=1.725 $X2=0 $Y2=0
cc_338 N_A2_M1017_g N_A1_M1020_g 0.0298582f $X=6.245 $Y=0.655 $X2=0 $Y2=0
cc_339 N_A2_M1018_g N_A1_M1011_g 0.0298582f $X=6.245 $Y=2.465 $X2=0 $Y2=0
cc_340 A2 N_A1_M1011_g 0.0146242f $X=5.915 $Y=1.95 $X2=0 $Y2=0
cc_341 N_A2_c_440_n N_A1_c_519_n 0.0127345f $X=6.335 $Y=1.51 $X2=0 $Y2=0
cc_342 A2 N_A1_c_519_n 0.0227931f $X=4.955 $Y=1.95 $X2=0 $Y2=0
cc_343 A2 N_A1_c_519_n 0.0304217f $X=5.915 $Y=1.95 $X2=0 $Y2=0
cc_344 N_A2_c_444_n N_A1_c_519_n 3.78294e-19 $X=4.935 $Y=1.51 $X2=0 $Y2=0
cc_345 N_A2_c_440_n N_A1_c_516_n 0.00528202f $X=6.335 $Y=1.51 $X2=0 $Y2=0
cc_346 N_A2_c_441_n N_A1_c_516_n 0.0298582f $X=6.335 $Y=1.51 $X2=0 $Y2=0
cc_347 A2 N_A1_c_516_n 0.00111845f $X=4.955 $Y=1.95 $X2=0 $Y2=0
cc_348 A2 N_A1_c_516_n 0.00405643f $X=5.915 $Y=1.95 $X2=0 $Y2=0
cc_349 N_A2_c_444_n N_A1_c_516_n 0.0255596f $X=4.935 $Y=1.51 $X2=0 $Y2=0
cc_350 A2 N_VPWR_M1005_d 0.00276569f $X=4.955 $Y=1.95 $X2=0 $Y2=0
cc_351 A2 N_VPWR_M1005_d 0.00768904f $X=5.915 $Y=1.95 $X2=0 $Y2=0
cc_352 A2 N_VPWR_M1011_d 0.00247599f $X=5.915 $Y=1.95 $X2=0 $Y2=0
cc_353 N_A2_c_450_n N_VPWR_c_568_n 0.0118341f $X=4.935 $Y=1.725 $X2=0 $Y2=0
cc_354 N_A2_M1018_g N_VPWR_c_569_n 0.0118284f $X=6.245 $Y=2.465 $X2=0 $Y2=0
cc_355 N_A2_c_450_n N_VPWR_c_572_n 0.00486043f $X=4.935 $Y=1.725 $X2=0 $Y2=0
cc_356 N_A2_M1018_g N_VPWR_c_574_n 0.00486043f $X=6.245 $Y=2.465 $X2=0 $Y2=0
cc_357 N_A2_M1018_g N_VPWR_c_563_n 0.00917987f $X=6.245 $Y=2.465 $X2=0 $Y2=0
cc_358 N_A2_c_450_n N_VPWR_c_563_n 0.00864313f $X=4.935 $Y=1.725 $X2=0 $Y2=0
cc_359 A2 N_A_527_367#_M1003_s 0.00428624f $X=5.915 $Y=1.95 $X2=0 $Y2=0
cc_360 A2 N_A_527_367#_c_757_n 0.0156847f $X=4.955 $Y=1.95 $X2=0 $Y2=0
cc_361 A2 N_A_527_367#_c_757_n 0.0194475f $X=5.915 $Y=1.95 $X2=0 $Y2=0
cc_362 N_A2_c_444_n N_A_527_367#_c_757_n 4.93198e-19 $X=4.935 $Y=1.51 $X2=0
+ $Y2=0
cc_363 N_A2_c_450_n N_A_527_367#_c_757_n 0.0167081f $X=4.935 $Y=1.725 $X2=0
+ $Y2=0
cc_364 N_A2_c_450_n N_A_527_367#_c_761_n 8.22713e-19 $X=4.935 $Y=1.725 $X2=0
+ $Y2=0
cc_365 N_A2_M1018_g N_A_527_367#_c_762_n 0.0121849f $X=6.245 $Y=2.465 $X2=0
+ $Y2=0
cc_366 N_A2_c_440_n N_A_527_367#_c_762_n 0.00366836f $X=6.335 $Y=1.51 $X2=0
+ $Y2=0
cc_367 A2 N_A_527_367#_c_762_n 0.0232526f $X=5.915 $Y=1.95 $X2=0 $Y2=0
cc_368 N_A2_M1018_g N_A_527_367#_c_730_n 0.00799783f $X=6.245 $Y=2.465 $X2=0
+ $Y2=0
cc_369 N_A2_c_440_n N_A_527_367#_c_730_n 0.016959f $X=6.335 $Y=1.51 $X2=0 $Y2=0
cc_370 N_A2_c_441_n N_A_527_367#_c_730_n 0.0043441f $X=6.335 $Y=1.51 $X2=0 $Y2=0
cc_371 A2 N_A_527_367#_c_730_n 0.00580369f $X=5.915 $Y=1.95 $X2=0 $Y2=0
cc_372 A2 N_A_527_367#_c_769_n 0.0153678f $X=5.915 $Y=1.95 $X2=0 $Y2=0
cc_373 N_A2_M1018_g N_A_527_367#_c_732_n 0.00157103f $X=6.245 $Y=2.465 $X2=0
+ $Y2=0
cc_374 N_A2_M1012_g N_VGND_c_822_n 0.00357731f $X=4.955 $Y=0.655 $X2=0 $Y2=0
cc_375 N_A2_M1017_g N_VGND_c_824_n 0.00813703f $X=6.245 $Y=0.655 $X2=0 $Y2=0
cc_376 N_A2_c_440_n N_VGND_c_824_n 0.00842153f $X=6.335 $Y=1.51 $X2=0 $Y2=0
cc_377 N_A2_c_441_n N_VGND_c_824_n 0.00298821f $X=6.335 $Y=1.51 $X2=0 $Y2=0
cc_378 N_A2_M1012_g N_VGND_c_830_n 0.00547432f $X=4.955 $Y=0.655 $X2=0 $Y2=0
cc_379 N_A2_M1017_g N_VGND_c_830_n 0.00547432f $X=6.245 $Y=0.655 $X2=0 $Y2=0
cc_380 N_A2_M1012_g N_VGND_c_835_n 0.0103951f $X=4.955 $Y=0.655 $X2=0 $Y2=0
cc_381 N_A2_M1017_g N_VGND_c_835_n 0.0106866f $X=6.245 $Y=0.655 $X2=0 $Y2=0
cc_382 N_A2_M1012_g N_A_1006_47#_c_923_n 0.00790597f $X=4.955 $Y=0.655 $X2=0
+ $Y2=0
cc_383 N_A2_M1017_g N_A_1006_47#_c_918_n 0.0117427f $X=6.245 $Y=0.655 $X2=0
+ $Y2=0
cc_384 N_A2_c_440_n N_A_1006_47#_c_918_n 0.0184983f $X=6.335 $Y=1.51 $X2=0 $Y2=0
cc_385 N_A1_M1003_g N_VPWR_c_568_n 0.00577291f $X=5.385 $Y=2.465 $X2=0 $Y2=0
cc_386 N_A1_M1003_g N_VPWR_c_569_n 6.44428e-19 $X=5.385 $Y=2.465 $X2=0 $Y2=0
cc_387 N_A1_M1011_g N_VPWR_c_569_n 0.0103844f $X=5.815 $Y=2.465 $X2=0 $Y2=0
cc_388 N_A1_M1003_g N_VPWR_c_573_n 0.0054895f $X=5.385 $Y=2.465 $X2=0 $Y2=0
cc_389 N_A1_M1011_g N_VPWR_c_573_n 0.00486043f $X=5.815 $Y=2.465 $X2=0 $Y2=0
cc_390 N_A1_M1003_g N_VPWR_c_563_n 0.0102704f $X=5.385 $Y=2.465 $X2=0 $Y2=0
cc_391 N_A1_M1011_g N_VPWR_c_563_n 0.00824727f $X=5.815 $Y=2.465 $X2=0 $Y2=0
cc_392 N_A1_M1003_g N_A_527_367#_c_757_n 0.0116122f $X=5.385 $Y=2.465 $X2=0
+ $Y2=0
cc_393 N_A1_M1003_g N_A_527_367#_c_761_n 0.00898828f $X=5.385 $Y=2.465 $X2=0
+ $Y2=0
cc_394 N_A1_M1011_g N_A_527_367#_c_762_n 0.0122129f $X=5.815 $Y=2.465 $X2=0
+ $Y2=0
cc_395 N_A1_M1011_g N_A_527_367#_c_730_n 9.9288e-19 $X=5.815 $Y=2.465 $X2=0
+ $Y2=0
cc_396 N_A1_M1003_g N_A_527_367#_c_769_n 7.32094e-19 $X=5.385 $Y=2.465 $X2=0
+ $Y2=0
cc_397 N_A1_M1009_g N_VGND_c_830_n 0.00357842f $X=5.385 $Y=0.655 $X2=0 $Y2=0
cc_398 N_A1_M1020_g N_VGND_c_830_n 0.00357842f $X=5.815 $Y=0.655 $X2=0 $Y2=0
cc_399 N_A1_M1009_g N_VGND_c_835_n 0.00537652f $X=5.385 $Y=0.655 $X2=0 $Y2=0
cc_400 N_A1_M1020_g N_VGND_c_835_n 0.00537652f $X=5.815 $Y=0.655 $X2=0 $Y2=0
cc_401 N_A1_M1009_g N_A_1006_47#_c_920_n 0.00853491f $X=5.385 $Y=0.655 $X2=0
+ $Y2=0
cc_402 N_A1_M1020_g N_A_1006_47#_c_920_n 0.0105205f $X=5.815 $Y=0.655 $X2=0
+ $Y2=0
cc_403 N_A1_M1009_g N_A_1006_47#_c_923_n 0.00712911f $X=5.385 $Y=0.655 $X2=0
+ $Y2=0
cc_404 N_A1_M1020_g N_A_1006_47#_c_923_n 5.19723e-19 $X=5.815 $Y=0.655 $X2=0
+ $Y2=0
cc_405 N_A1_M1009_g N_A_1006_47#_c_918_n 5.91586e-19 $X=5.385 $Y=0.655 $X2=0
+ $Y2=0
cc_406 N_A1_M1020_g N_A_1006_47#_c_918_n 0.0119924f $X=5.815 $Y=0.655 $X2=0
+ $Y2=0
cc_407 N_VPWR_c_563_n N_X_M1001_s 0.00536646f $X=6.48 $Y=3.33 $X2=0 $Y2=0
cc_408 N_VPWR_c_563_n N_X_M1014_s 0.00536646f $X=6.48 $Y=3.33 $X2=0 $Y2=0
cc_409 N_VPWR_M1001_d N_X_c_672_n 0.00119058f $X=0.25 $Y=1.835 $X2=0 $Y2=0
cc_410 N_VPWR_c_565_n N_X_c_672_n 0.0109431f $X=0.375 $Y=2.18 $X2=0 $Y2=0
cc_411 N_VPWR_M1001_d N_X_c_673_n 0.00147472f $X=0.25 $Y=1.835 $X2=0 $Y2=0
cc_412 N_VPWR_c_565_n N_X_c_673_n 0.0122196f $X=0.375 $Y=2.18 $X2=0 $Y2=0
cc_413 N_VPWR_c_570_n N_X_c_709_n 0.0124525f $X=1.07 $Y=3.33 $X2=0 $Y2=0
cc_414 N_VPWR_c_563_n N_X_c_709_n 0.00730901f $X=6.48 $Y=3.33 $X2=0 $Y2=0
cc_415 N_VPWR_M1006_d N_X_c_674_n 0.00180746f $X=1.095 $Y=1.835 $X2=0 $Y2=0
cc_416 N_VPWR_c_566_n N_X_c_674_n 0.0163515f $X=1.235 $Y=2.19 $X2=0 $Y2=0
cc_417 N_VPWR_c_567_n N_X_c_674_n 0.00503283f $X=2.095 $Y=1.98 $X2=0 $Y2=0
cc_418 N_VPWR_c_571_n N_X_c_714_n 0.0124525f $X=1.93 $Y=3.33 $X2=0 $Y2=0
cc_419 N_VPWR_c_563_n N_X_c_714_n 0.00730901f $X=6.48 $Y=3.33 $X2=0 $Y2=0
cc_420 N_VPWR_c_563_n N_A_527_367#_M1015_s 0.00236551f $X=6.48 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_421 N_VPWR_c_563_n N_A_527_367#_M1022_s 0.00469832f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_422 N_VPWR_c_563_n N_A_527_367#_M1003_s 0.00380103f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_423 N_VPWR_c_563_n N_A_527_367#_M1018_s 0.00371702f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_424 N_VPWR_c_572_n N_A_527_367#_c_735_n 0.00304528f $X=4.895 $Y=3.33 $X2=0
+ $Y2=0
cc_425 N_VPWR_c_563_n N_A_527_367#_c_735_n 0.00704301f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_426 N_VPWR_c_572_n N_A_527_367#_c_738_n 3.86733e-19 $X=4.895 $Y=3.33 $X2=0
+ $Y2=0
cc_427 N_VPWR_c_563_n N_A_527_367#_c_738_n 6.58305e-19 $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_428 N_VPWR_c_572_n N_A_527_367#_c_784_n 0.0216061f $X=4.895 $Y=3.33 $X2=0
+ $Y2=0
cc_429 N_VPWR_c_563_n N_A_527_367#_c_784_n 0.0131407f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_430 N_VPWR_M1005_d N_A_527_367#_c_757_n 0.00682624f $X=4.92 $Y=1.835 $X2=0
+ $Y2=0
cc_431 N_VPWR_c_568_n N_A_527_367#_c_757_n 0.0218816f $X=5.06 $Y=2.77 $X2=0
+ $Y2=0
cc_432 N_VPWR_c_568_n N_A_527_367#_c_761_n 0.0288558f $X=5.06 $Y=2.77 $X2=0
+ $Y2=0
cc_433 N_VPWR_c_573_n N_A_527_367#_c_761_n 0.015688f $X=5.865 $Y=3.33 $X2=0
+ $Y2=0
cc_434 N_VPWR_c_563_n N_A_527_367#_c_761_n 0.00984745f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_435 N_VPWR_M1011_d N_A_527_367#_c_762_n 0.00352922f $X=5.89 $Y=1.835 $X2=0
+ $Y2=0
cc_436 N_VPWR_c_569_n N_A_527_367#_c_762_n 0.0170777f $X=6.03 $Y=2.785 $X2=0
+ $Y2=0
cc_437 N_VPWR_c_567_n N_A_527_367#_c_731_n 0.0365236f $X=2.095 $Y=1.98 $X2=0
+ $Y2=0
cc_438 N_VPWR_c_572_n N_A_527_367#_c_731_n 0.0185173f $X=4.895 $Y=3.33 $X2=0
+ $Y2=0
cc_439 N_VPWR_c_563_n N_A_527_367#_c_731_n 0.011737f $X=6.48 $Y=3.33 $X2=0 $Y2=0
cc_440 N_VPWR_c_574_n N_A_527_367#_c_732_n 0.0178111f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_441 N_VPWR_c_563_n N_A_527_367#_c_732_n 0.0100304f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_442 N_VPWR_c_563_n N_A_610_367#_M1015_d 0.00224306f $X=6.48 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_443 N_VPWR_c_563_n N_A_610_367#_M1010_d 0.00263626f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_444 N_VPWR_c_572_n N_A_610_367#_c_802_n 0.0598996f $X=4.895 $Y=3.33 $X2=0
+ $Y2=0
cc_445 N_VPWR_c_563_n N_A_610_367#_c_802_n 0.0430426f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_446 N_X_c_666_n N_VGND_M1007_s 0.00230047f $X=1.265 $Y=1.14 $X2=-0.19
+ $Y2=-0.245
cc_447 N_X_c_667_n N_VGND_M1008_s 0.00176773f $X=2.125 $Y=1.135 $X2=0 $Y2=0
cc_448 N_X_c_666_n N_VGND_c_817_n 0.0220025f $X=1.265 $Y=1.14 $X2=0 $Y2=0
cc_449 X N_VGND_c_817_n 0.0244516f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_450 N_X_c_720_p N_VGND_c_818_n 0.0124525f $X=1.36 $Y=0.42 $X2=0 $Y2=0
cc_451 N_X_c_667_n N_VGND_c_819_n 0.0171443f $X=2.125 $Y=1.135 $X2=0 $Y2=0
cc_452 N_X_c_694_n N_VGND_c_820_n 0.036685f $X=2.22 $Y=0.42 $X2=0 $Y2=0
cc_453 X N_VGND_c_825_n 0.0120288f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_454 N_X_c_694_n N_VGND_c_827_n 0.0121325f $X=2.22 $Y=0.42 $X2=0 $Y2=0
cc_455 N_X_M1007_d N_VGND_c_835_n 0.00536646f $X=1.22 $Y=0.235 $X2=0 $Y2=0
cc_456 N_X_M1013_d N_VGND_c_835_n 0.00635678f $X=2.08 $Y=0.235 $X2=0 $Y2=0
cc_457 N_X_c_720_p N_VGND_c_835_n 0.00730901f $X=1.36 $Y=0.42 $X2=0 $Y2=0
cc_458 N_X_c_694_n N_VGND_c_835_n 0.00692023f $X=2.22 $Y=0.42 $X2=0 $Y2=0
cc_459 X N_VGND_c_835_n 0.0112771f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_460 N_A_527_367#_c_735_n N_A_610_367#_M1015_d 0.00368379f $X=4.355 $Y=2.51
+ $X2=-0.19 $Y2=1.655
cc_461 N_A_527_367#_c_735_n N_A_610_367#_M1010_d 0.00606553f $X=4.355 $Y=2.51
+ $X2=0 $Y2=0
cc_462 N_A_527_367#_c_735_n N_A_610_367#_c_802_n 0.0611746f $X=4.355 $Y=2.51
+ $X2=0 $Y2=0
cc_463 N_VGND_c_835_n N_A_1006_47#_M1012_d 0.00223559f $X=6.48 $Y=0 $X2=-0.19
+ $Y2=-0.245
cc_464 N_VGND_c_835_n N_A_1006_47#_M1020_d 0.00223559f $X=6.48 $Y=0 $X2=0 $Y2=0
cc_465 N_VGND_c_830_n N_A_1006_47#_c_920_n 0.0298674f $X=6.365 $Y=0 $X2=0 $Y2=0
cc_466 N_VGND_c_835_n N_A_1006_47#_c_920_n 0.0187823f $X=6.48 $Y=0 $X2=0 $Y2=0
cc_467 N_VGND_c_830_n N_A_1006_47#_c_923_n 0.0189944f $X=6.365 $Y=0 $X2=0 $Y2=0
cc_468 N_VGND_c_835_n N_A_1006_47#_c_923_n 0.0124345f $X=6.48 $Y=0 $X2=0 $Y2=0
cc_469 N_VGND_c_824_n N_A_1006_47#_c_918_n 0.0258649f $X=6.46 $Y=0.38 $X2=0
+ $Y2=0
cc_470 N_VGND_c_830_n N_A_1006_47#_c_918_n 0.01906f $X=6.365 $Y=0 $X2=0 $Y2=0
cc_471 N_VGND_c_835_n N_A_1006_47#_c_918_n 0.0124545f $X=6.48 $Y=0 $X2=0 $Y2=0
