* File: sky130_fd_sc_lp__nand2_m.pxi.spice
* Created: Fri Aug 28 10:47:49 2020
* 
x_PM_SKY130_FD_SC_LP__NAND2_M%B N_B_c_31_n N_B_M1000_g N_B_M1003_g N_B_c_34_n B
+ B B B N_B_c_36_n PM_SKY130_FD_SC_LP__NAND2_M%B
x_PM_SKY130_FD_SC_LP__NAND2_M%A N_A_M1001_g N_A_c_64_n N_A_M1002_g N_A_c_66_n A
+ A A A N_A_c_68_n PM_SKY130_FD_SC_LP__NAND2_M%A
x_PM_SKY130_FD_SC_LP__NAND2_M%VPWR N_VPWR_M1000_s N_VPWR_M1002_d N_VPWR_c_90_n
+ N_VPWR_c_91_n N_VPWR_c_92_n N_VPWR_c_93_n VPWR N_VPWR_c_94_n N_VPWR_c_89_n
+ PM_SKY130_FD_SC_LP__NAND2_M%VPWR
x_PM_SKY130_FD_SC_LP__NAND2_M%Y N_Y_M1001_d N_Y_M1000_d Y Y Y Y Y Y Y
+ N_Y_c_117_n N_Y_c_109_n PM_SKY130_FD_SC_LP__NAND2_M%Y
x_PM_SKY130_FD_SC_LP__NAND2_M%VGND N_VGND_M1003_s N_VGND_c_133_n N_VGND_c_134_n
+ VGND N_VGND_c_135_n N_VGND_c_136_n PM_SKY130_FD_SC_LP__NAND2_M%VGND
cc_1 VNB N_B_c_31_n 0.0202004f $X=-0.19 $Y=-0.245 $X2=0.402 $Y2=1.293
cc_2 VNB N_B_M1000_g 0.00912584f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.52
cc_3 VNB N_B_M1003_g 0.0268086f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=0.445
cc_4 VNB N_B_c_34_n 0.0277158f $X=-0.19 $Y=-0.245 $X2=0.402 $Y2=1.51
cc_5 VNB B 0.0334658f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_6 VNB N_B_c_36_n 0.0272544f $X=-0.19 $Y=-0.245 $X2=0.35 $Y2=1.005
cc_7 VNB N_A_M1001_g 0.0276393f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.51
cc_8 VNB N_A_c_64_n 0.0253353f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_M1002_g 0.00912683f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=0.445
cc_10 VNB N_A_c_66_n 0.0225369f $X=-0.19 $Y=-0.245 $X2=0.402 $Y2=1.51
cc_11 VNB A 0.0328414f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_12 VNB N_A_c_68_n 0.0225369f $X=-0.19 $Y=-0.245 $X2=0.35 $Y2=1.005
cc_13 VNB N_VPWR_c_89_n 0.0641695f $X=-0.19 $Y=-0.245 $X2=0.295 $Y2=1.005
cc_14 VNB Y 0.00742946f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=0.445
cc_15 VNB N_Y_c_109_n 0.00360633f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_VGND_c_133_n 0.0133899f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.52
cc_17 VNB N_VGND_c_134_n 0.00495479f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_VGND_c_135_n 0.0289321f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_19 VNB N_VGND_c_136_n 0.113477f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_20 VPB N_B_M1000_g 0.0565969f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=2.52
cc_21 VPB B 0.0231554f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_22 VPB N_A_M1002_g 0.0566023f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=0.445
cc_23 VPB A 0.0232996f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_24 VPB N_VPWR_c_90_n 0.0121156f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=0.84
cc_25 VPB N_VPWR_c_91_n 0.0260741f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=0.445
cc_26 VPB N_VPWR_c_92_n 0.0121156f $X=-0.19 $Y=1.655 $X2=0.402 $Y2=1.51
cc_27 VPB N_VPWR_c_93_n 0.026138f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_28 VPB N_VPWR_c_94_n 0.0191805f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_29 VPB N_VPWR_c_89_n 0.0640933f $X=-0.19 $Y=1.655 $X2=0.295 $Y2=1.005
cc_30 VPB Y 0.0204255f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=0.445
cc_31 N_B_M1003_g N_A_M1001_g 0.018697f $X=0.545 $Y=0.445 $X2=0 $Y2=0
cc_32 N_B_c_31_n N_A_c_64_n 0.018697f $X=0.402 $Y=1.293 $X2=0 $Y2=0
cc_33 N_B_M1000_g N_A_M1002_g 0.0334758f $X=0.505 $Y=2.52 $X2=0 $Y2=0
cc_34 N_B_c_34_n N_A_c_66_n 0.018697f $X=0.402 $Y=1.51 $X2=0 $Y2=0
cc_35 N_B_c_36_n A 5.09445e-19 $X=0.35 $Y=1.005 $X2=0 $Y2=0
cc_36 N_B_c_36_n N_A_c_68_n 0.018697f $X=0.35 $Y=1.005 $X2=0 $Y2=0
cc_37 N_B_M1000_g N_VPWR_c_91_n 0.00385941f $X=0.505 $Y=2.52 $X2=0 $Y2=0
cc_38 B N_VPWR_c_91_n 0.0187102f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_39 N_B_M1000_g N_VPWR_c_94_n 0.00428744f $X=0.505 $Y=2.52 $X2=0 $Y2=0
cc_40 N_B_M1000_g N_VPWR_c_89_n 0.00476395f $X=0.505 $Y=2.52 $X2=0 $Y2=0
cc_41 N_B_c_31_n Y 0.00509613f $X=0.402 $Y=1.293 $X2=0 $Y2=0
cc_42 N_B_M1000_g Y 0.0103489f $X=0.505 $Y=2.52 $X2=0 $Y2=0
cc_43 N_B_M1003_g Y 0.00826999f $X=0.545 $Y=0.445 $X2=0 $Y2=0
cc_44 N_B_c_34_n Y 0.0047259f $X=0.402 $Y=1.51 $X2=0 $Y2=0
cc_45 B Y 0.0890472f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_46 N_B_c_36_n Y 0.0047259f $X=0.35 $Y=1.005 $X2=0 $Y2=0
cc_47 N_B_M1003_g N_Y_c_117_n 0.0105942f $X=0.545 $Y=0.445 $X2=0 $Y2=0
cc_48 N_B_M1003_g N_VGND_c_134_n 0.00460896f $X=0.545 $Y=0.445 $X2=0 $Y2=0
cc_49 B N_VGND_c_134_n 0.0101959f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_50 N_B_c_36_n N_VGND_c_134_n 0.0014208f $X=0.35 $Y=1.005 $X2=0 $Y2=0
cc_51 N_B_M1003_g N_VGND_c_135_n 0.00578301f $X=0.545 $Y=0.445 $X2=0 $Y2=0
cc_52 N_B_M1003_g N_VGND_c_136_n 0.0114256f $X=0.545 $Y=0.445 $X2=0 $Y2=0
cc_53 B N_VGND_c_136_n 0.0034919f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_54 N_B_c_36_n N_VGND_c_136_n 8.84992e-19 $X=0.35 $Y=1.005 $X2=0 $Y2=0
cc_55 N_A_M1002_g N_VPWR_c_93_n 0.00390217f $X=0.935 $Y=2.52 $X2=0 $Y2=0
cc_56 A N_VPWR_c_93_n 0.0187102f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_57 N_A_M1002_g N_VPWR_c_94_n 0.00428744f $X=0.935 $Y=2.52 $X2=0 $Y2=0
cc_58 N_A_M1002_g N_VPWR_c_89_n 0.00476395f $X=0.935 $Y=2.52 $X2=0 $Y2=0
cc_59 N_A_M1001_g Y 0.0193358f $X=0.935 $Y=0.445 $X2=0 $Y2=0
cc_60 A Y 0.0921479f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_61 N_A_M1001_g N_Y_c_109_n 0.0160498f $X=0.935 $Y=0.445 $X2=0 $Y2=0
cc_62 A N_Y_c_109_n 0.0209761f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_63 N_A_c_68_n N_Y_c_109_n 0.00163158f $X=1.07 $Y=1.005 $X2=0 $Y2=0
cc_64 N_A_M1001_g N_VGND_c_135_n 0.00373071f $X=0.935 $Y=0.445 $X2=0 $Y2=0
cc_65 N_A_M1001_g N_VGND_c_136_n 0.00641194f $X=0.935 $Y=0.445 $X2=0 $Y2=0
cc_66 A N_VGND_c_136_n 0.0015741f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_67 N_VPWR_c_91_n Y 0.0159684f $X=0.29 $Y=2.525 $X2=0 $Y2=0
cc_68 N_VPWR_c_93_n Y 0.0150336f $X=1.15 $Y=2.525 $X2=0 $Y2=0
cc_69 N_VPWR_c_94_n Y 0.00806491f $X=1.045 $Y=3.33 $X2=0 $Y2=0
cc_70 N_VPWR_c_89_n Y 0.00690154f $X=1.2 $Y=3.33 $X2=0 $Y2=0
cc_71 N_Y_c_117_n N_VGND_c_135_n 0.00764381f $X=0.71 $Y=0.66 $X2=0 $Y2=0
cc_72 N_Y_c_109_n N_VGND_c_135_n 0.0176173f $X=1.15 $Y=0.495 $X2=0 $Y2=0
cc_73 N_Y_M1001_d N_VGND_c_136_n 0.00234684f $X=1.01 $Y=0.235 $X2=0 $Y2=0
cc_74 N_Y_c_117_n N_VGND_c_136_n 0.00706408f $X=0.71 $Y=0.66 $X2=0 $Y2=0
cc_75 N_Y_c_109_n N_VGND_c_136_n 0.0157023f $X=1.15 $Y=0.495 $X2=0 $Y2=0
cc_76 N_Y_c_117_n A_124_47# 0.00143918f $X=0.71 $Y=0.66 $X2=-0.19 $Y2=-0.245
cc_77 N_VGND_c_136_n A_124_47# 0.00198279f $X=1.2 $Y=0 $X2=-0.19 $Y2=-0.245
