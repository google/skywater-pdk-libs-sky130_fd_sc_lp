* NGSPICE file created from sky130_fd_sc_lp__a2bb2oi_2.ext - technology: sky130A

.subckt sky130_fd_sc_lp__a2bb2oi_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
M1000 VGND A2_N a_459_39# VNB nshort w=840000u l=150000u
+  ad=1.7262e+12p pd=1.251e+07u as=4.704e+11p ps=4.48e+06u
M1001 VPWR A1_N a_699_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=1.26e+12p pd=9.56e+06u as=1.0206e+12p ps=9.18e+06u
M1002 a_30_367# B1 VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=1.3734e+12p pd=1.226e+07u as=0p ps=0u
M1003 Y a_459_39# VGND VNB nshort w=840000u l=150000u
+  ad=4.704e+11p pd=4.48e+06u as=0p ps=0u
M1004 Y B2 a_113_65# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=5.376e+11p ps=4.64e+06u
M1005 a_30_367# B2 VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_459_39# A2_N a_699_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=3.528e+11p pd=3.08e+06u as=0p ps=0u
M1007 a_30_367# a_459_39# Y VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=3.528e+11p ps=3.08e+06u
M1008 a_113_65# B2 Y VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND a_459_39# Y VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND A1_N a_459_39# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR B1 a_30_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VPWR B2 a_30_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_699_367# A1_N VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_699_367# A2_N a_459_39# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VGND B1 a_113_65# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 Y a_459_39# a_30_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_459_39# A2_N VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_113_65# B1 VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_459_39# A1_N VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

