* File: sky130_fd_sc_lp__a2111oi_lp.spice
* Created: Wed Sep  2 09:17:08 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__a2111oi_lp.pex.spice"
.subckt sky130_fd_sc_lp__a2111oi_lp  VNB VPB A1 A2 B1 C1 D1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* D1	D1
* C1	C1
* B1	B1
* A2	A2
* A1	A1
* VPB	VPB
* VNB	VNB
MM1008 A_125_57# N_A1_M1008_g N_Y_M1008_s VNB NSHORT L=0.15 W=0.42 AD=0.0504
+ AS=0.1197 PD=0.66 PS=1.41 NRD=18.564 NRS=0 M=1 R=2.8 SA=75000.2 SB=75001.4
+ A=0.063 P=1.14 MULT=1
MM1005 N_VGND_M1005_d N_A2_M1005_g A_125_57# VNB NSHORT L=0.15 W=0.42 AD=0.0588
+ AS=0.0504 PD=0.7 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75000.6 SB=75001
+ A=0.063 P=1.14 MULT=1
MM1000 A_289_57# N_B1_M1000_g N_VGND_M1005_d VNB NSHORT L=0.15 W=0.42 AD=0.0441
+ AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75001 SB=75000.6 A=0.063
+ P=1.14 MULT=1
MM1009 N_Y_M1009_d N_B1_M1009_g A_289_57# VNB NSHORT L=0.15 W=0.42 AD=0.1134
+ AS=0.0441 PD=1.38 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.4 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1001 A_553_47# N_C1_M1001_g N_VGND_M1001_s VNB NSHORT L=0.15 W=0.42 AD=0.0441
+ AS=0.1134 PD=0.63 PS=1.38 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2 SB=75001.3
+ A=0.063 P=1.14 MULT=1
MM1010 N_Y_M1010_d N_C1_M1010_g A_553_47# VNB NSHORT L=0.15 W=0.42 AD=0.0588
+ AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6 SB=75001 A=0.063
+ P=1.14 MULT=1
MM1002 A_711_47# N_D1_M1002_g N_Y_M1010_d VNB NSHORT L=0.15 W=0.42 AD=0.0441
+ AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75001 SB=75000.6 A=0.063
+ P=1.14 MULT=1
MM1003 N_VGND_M1003_d N_D1_M1003_g A_711_47# VNB NSHORT L=0.15 W=0.42 AD=0.1134
+ AS=0.0441 PD=1.38 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.3 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1006 N_A_131_409#_M1006_d N_A1_M1006_g N_VPWR_M1006_s VPB PHIGHVT L=0.25 W=1
+ AD=0.14 AS=0.27 PD=1.28 PS=2.54 NRD=0 NRS=0 M=1 R=4 SA=125000 SB=125001 A=0.25
+ P=2.5 MULT=1
MM1012 N_VPWR_M1012_d N_A2_M1012_g N_A_131_409#_M1006_d VPB PHIGHVT L=0.25 W=1
+ AD=0.285 AS=0.14 PD=2.57 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125001 SB=125000
+ A=0.25 P=2.5 MULT=1
MM1004 A_539_409# N_B1_M1004_g N_A_131_409#_M1004_s VPB PHIGHVT L=0.25 W=1
+ AD=0.12 AS=0.285 PD=1.24 PS=2.57 NRD=12.7853 NRS=0 M=1 R=4 SA=125000 SB=125001
+ A=0.25 P=2.5 MULT=1
MM1007 A_637_409# N_C1_M1007_g A_539_409# VPB PHIGHVT L=0.25 W=1 AD=0.16 AS=0.12
+ PD=1.32 PS=1.24 NRD=20.6653 NRS=12.7853 M=1 R=4 SA=125001 SB=125001 A=0.25
+ P=2.5 MULT=1
MM1011 N_Y_M1011_d N_D1_M1011_g A_637_409# VPB PHIGHVT L=0.25 W=1 AD=0.285
+ AS=0.16 PD=2.57 PS=1.32 NRD=0 NRS=20.6653 M=1 R=4 SA=125001 SB=125000 A=0.25
+ P=2.5 MULT=1
DX13_noxref VNB VPB NWDIODE A=8.7655 P=13.13
*
.include "sky130_fd_sc_lp__a2111oi_lp.pxi.spice"
*
.ends
*
*
