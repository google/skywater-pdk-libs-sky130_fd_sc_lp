* NGSPICE file created from sky130_fd_sc_lp__srdlrtp_1.ext - technology: sky130A

.subckt sky130_fd_sc_lp__srdlrtp_1 D GATE RESET_B SLEEP_B KAPWR VGND VNB VPB VPWR
+ Q
M1000 a_393_335# GATE KAPWR VPB phighvt w=640000u l=150000u
+  ad=5.439e+11p pd=3.8e+06u as=1.1128e+12p ps=9.79e+06u
M1001 VGND SLEEP_B a_1147_97# VNB nshort w=420000u l=150000u
+  ad=1.19685e+12p pd=1.055e+07u as=8.82e+10p ps=1.26e+06u
M1002 a_366_97# a_336_71# a_280_97# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=1.176e+11p ps=1.4e+06u
M1003 a_1344_97# SLEEP_B VGND VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1004 KAPWR a_438_97# a_612_71# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=5.1e+11p ps=3.02e+06u
M1005 a_114_97# D a_27_97# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=1.197e+11p ps=1.41e+06u
M1006 a_336_71# a_393_335# VGND VNB nshort w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=0p ps=0u
M1007 VGND a_1324_394# a_1624_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=2.415e+11p ps=2.83e+06u
M1008 a_280_97# a_27_97# VPWR VPB phighvt w=640000u l=150000u
+  ad=1.792e+11p pd=1.84e+06u as=1.3453e+12p ps=1.069e+07u
M1009 a_1765_419# a_1324_394# KAPWR VPB phighvt w=1e+06u l=250000u
+  ad=2.1e+11p pd=2.42e+06u as=0p ps=0u
M1010 a_438_97# a_336_71# a_366_97# VNB nshort w=420000u l=150000u
+  ad=2.142e+11p pd=1.86e+06u as=0p ps=0u
M1011 a_1917_47# a_438_97# a_1624_47# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1012 Q a_2120_55# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=3.591e+11p pd=3.09e+06u as=0p ps=0u
M1013 a_612_71# a_438_97# a_1917_47# VNB nshort w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=0p ps=0u
M1014 a_612_71# RESET_B a_1765_419# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VGND a_612_71# a_642_97# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1016 Q a_2120_55# VGND VNB nshort w=840000u l=150000u
+  ad=2.394e+11p pd=2.25e+06u as=0p ps=0u
M1017 VGND a_438_97# a_2120_55# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1018 a_423_487# a_393_335# a_280_97# VPB phighvt w=640000u l=150000u
+  ad=1.344e+11p pd=1.7e+06u as=0p ps=0u
M1019 a_1069_97# GATE a_393_335# VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=1.197e+11p ps=1.41e+06u
M1020 a_1147_97# SLEEP_B a_1069_97# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_438_97# a_393_335# a_423_487# VPB phighvt w=640000u l=150000u
+  ad=4.674e+11p pd=4.42e+06u as=0p ps=0u
M1022 a_1624_47# RESET_B VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_1324_394# SLEEP_B KAPWR VPB phighvt w=1e+06u l=250000u
+  ad=5.131e+11p pd=3.58e+06u as=0p ps=0u
M1024 a_570_97# a_393_335# a_438_97# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1025 a_280_97# a_27_97# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_642_97# a_612_71# a_570_97# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_1565_419# a_336_71# a_438_97# VPB phighvt w=1e+06u l=250000u
+  ad=2.1e+11p pd=2.42e+06u as=0p ps=0u
M1028 KAPWR a_612_71# a_1565_419# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1029 a_1324_394# SLEEP_B a_1344_97# VNB nshort w=420000u l=150000u
+  ad=1.68e+11p pd=1.64e+06u as=0p ps=0u
M1030 VGND RESET_B a_114_97# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 VPWR RESET_B a_27_97# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=2.24e+11p ps=1.98e+06u
M1032 a_27_97# D VPWR VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 VPWR a_393_335# a_336_71# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=2.6615e+11p ps=2.15e+06u
M1034 VPWR a_438_97# a_2120_55# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.824e+11p ps=1.85e+06u
M1035 KAPWR SLEEP_B a_393_335# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

