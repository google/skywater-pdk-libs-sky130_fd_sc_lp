* File: sky130_fd_sc_lp__o21ba_0.spice
* Created: Wed Sep  2 10:16:35 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__o21ba_0.pex.spice"
.subckt sky130_fd_sc_lp__o21ba_0  VNB VPB B1_N A2 A1 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* A1	A1
* A2	A2
* B1_N	B1_N
* VPB	VPB
* VNB	VNB
MM1002 N_VGND_M1002_d N_A_80_225#_M1002_g N_X_M1002_s VNB NSHORT L=0.15 W=0.42
+ AD=0.1302 AS=0.1113 PD=1.04 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75001
+ A=0.063 P=1.14 MULT=1
MM1006 N_A_258_397#_M1006_d N_B1_N_M1006_g N_VGND_M1002_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1113 AS=0.1302 PD=1.37 PS=1.04 NRD=0 NRS=0 M=1 R=2.8 SA=75001
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1004 N_A_499_47#_M1004_d N_A_258_397#_M1004_g N_A_80_225#_M1004_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1008 N_VGND_M1008_d N_A2_M1008_g N_A_499_47#_M1004_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1000 N_A_499_47#_M1000_d N_A1_M1000_g N_VGND_M1008_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.1 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1001 N_VPWR_M1001_d N_A_80_225#_M1001_g N_X_M1001_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.184815 AS=0.1696 PD=1.48528 PS=1.81 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75000.7 A=0.096 P=1.58 MULT=1
MM1007 N_A_258_397#_M1007_d N_B1_N_M1007_g N_VPWR_M1001_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1113 AS=0.121285 PD=1.37 PS=0.974717 NRD=0 NRS=146.568 M=1 R=2.8
+ SA=75000.9 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1005 N_A_80_225#_M1005_d N_A_258_397#_M1005_g N_VPWR_M1005_s VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.0896 AS=0.1824 PD=0.92 PS=1.85 NRD=0 NRS=6.1464 M=1
+ R=4.26667 SA=75000.2 SB=75001 A=0.096 P=1.58 MULT=1
MM1003 A_557_487# N_A2_M1003_g N_A_80_225#_M1005_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0768 AS=0.0896 PD=0.88 PS=0.92 NRD=19.9955 NRS=0 M=1 R=4.26667 SA=75000.6
+ SB=75000.6 A=0.096 P=1.58 MULT=1
MM1009 N_VPWR_M1009_d N_A1_M1009_g A_557_487# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1696 AS=0.0768 PD=1.81 PS=0.88 NRD=0 NRS=19.9955 M=1 R=4.26667 SA=75001
+ SB=75000.2 A=0.096 P=1.58 MULT=1
DX10_noxref VNB VPB NWDIODE A=7.8703 P=12.17
c_76 VPB 0 1.4009e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_lp__o21ba_0.pxi.spice"
*
.ends
*
*
