* File: sky130_fd_sc_lp__nor4bb_1.spice
* Created: Fri Aug 28 10:58:54 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__nor4bb_1.pex.spice"
.subckt sky130_fd_sc_lp__nor4bb_1  VNB VPB D_N B A C_N VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* C_N	C_N
* A	A
* B	B
* D_N	D_N
* VPB	VPB
* VNB	VNB
MM1006 N_VGND_M1006_d N_D_N_M1006_g N_A_27_508#_M1006_s VNB NSHORT L=0.15 W=0.42
+ AD=0.1253 AS=0.1113 PD=0.98 PS=1.37 NRD=85.704 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75003.2 A=0.063 P=1.14 MULT=1
MM1009 N_Y_M1009_d N_A_27_508#_M1009_g N_VGND_M1006_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2506 PD=1.12 PS=1.96 NRD=0 NRS=3.564 M=1 R=5.6 SA=75000.6
+ SB=75002 A=0.126 P=1.98 MULT=1
MM1001 N_VGND_M1001_d N_A_375_269#_M1001_g N_Y_M1009_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1617 AS=0.1176 PD=1.225 PS=1.12 NRD=6.42 NRS=0 M=1 R=5.6 SA=75001
+ SB=75001.6 A=0.126 P=1.98 MULT=1
MM1007 N_Y_M1007_d N_B_M1007_g N_VGND_M1001_d VNB NSHORT L=0.15 W=0.84 AD=0.1365
+ AS=0.1617 PD=1.165 PS=1.225 NRD=0 NRS=8.568 M=1 R=5.6 SA=75001.5 SB=75001
+ A=0.126 P=1.98 MULT=1
MM1000 N_VGND_M1000_d N_A_M1000_g N_Y_M1007_d VNB NSHORT L=0.15 W=0.84 AD=0.2478
+ AS=0.1365 PD=1.94667 PS=1.165 NRD=0 NRS=6.42 M=1 R=5.6 SA=75002 SB=75000.6
+ A=0.126 P=1.98 MULT=1
MM1010 N_A_375_269#_M1010_d N_C_N_M1010_g N_VGND_M1000_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1113 AS=0.1239 PD=1.37 PS=0.973333 NRD=0 NRS=0 M=1 R=2.8
+ SA=75003.2 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1002 N_VPWR_M1002_d N_D_N_M1002_g N_A_27_508#_M1002_s VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1113 AS=0.1113 PD=1.37 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1004 A_333_367# N_A_27_508#_M1004_g N_Y_M1004_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1323 AS=0.3339 PD=1.47 PS=3.05 NRD=7.8012 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75001.8 A=0.189 P=2.82 MULT=1
MM1011 A_405_367# N_A_375_269#_M1011_g A_333_367# VPB PHIGHVT L=0.15 W=1.26
+ AD=0.2457 AS=0.1323 PD=1.65 PS=1.47 NRD=21.8867 NRS=7.8012 M=1 R=8.4
+ SA=75000.6 SB=75001.4 A=0.189 P=2.82 MULT=1
MM1005 A_513_367# N_B_M1005_g A_405_367# VPB PHIGHVT L=0.15 W=1.26 AD=0.2457
+ AS=0.2457 PD=1.65 PS=1.65 NRD=21.8867 NRS=21.8867 M=1 R=8.4 SA=75001.1
+ SB=75000.9 A=0.189 P=2.82 MULT=1
MM1008 N_VPWR_M1008_d N_A_M1008_g A_513_367# VPB PHIGHVT L=0.15 W=1.26 AD=0.2898
+ AS=0.2457 PD=2.475 PS=1.65 NRD=0 NRS=21.8867 M=1 R=8.4 SA=75001.6 SB=75000.4
+ A=0.189 P=2.82 MULT=1
MM1003 N_A_375_269#_M1003_d N_C_N_M1003_g N_VPWR_M1008_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1113 AS=0.0966 PD=1.37 PS=0.825 NRD=0 NRS=82.0702 M=1 R=2.8
+ SA=75002.2 SB=75000.2 A=0.063 P=1.14 MULT=1
DX12_noxref VNB VPB NWDIODE A=8.7655 P=13.13
c_40 VNB 0 1.01016e-19 $X=0 $Y=0
*
.include "sky130_fd_sc_lp__nor4bb_1.pxi.spice"
*
.ends
*
*
