* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__dfsbp_1 CLK D SET_B VGND VNB VPB VPWR Q Q_N
X0 VGND a_1331_151# a_2005_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 VPWR CLK a_111_156# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X2 a_494_119# a_111_156# a_580_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 a_1331_151# a_161_21# a_1141_125# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X4 a_1472_449# a_1535_177# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X5 a_1248_151# a_1535_177# a_1657_71# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 VGND CLK a_111_156# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 VPWR a_1331_151# Q_N VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X8 Q a_2005_119# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X9 a_1657_71# SET_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 Q a_2005_119# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X11 VPWR SET_B a_1331_151# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X12 VPWR D a_494_119# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X13 VGND a_1331_151# Q_N VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X14 a_708_93# a_580_119# a_964_169# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X15 a_1331_151# a_161_21# a_1472_449# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X16 a_666_119# a_708_93# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X17 VPWR a_580_119# a_708_93# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X18 a_1535_177# a_1331_151# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X19 a_580_119# a_111_156# a_687_533# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X20 a_687_533# a_708_93# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X21 VPWR a_1331_151# a_2005_119# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X22 a_161_21# a_111_156# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X23 a_494_119# a_161_21# a_580_119# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X24 a_1535_177# a_1331_151# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X25 VGND D a_494_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X26 a_1259_449# a_111_156# a_1331_151# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X27 a_580_119# a_161_21# a_666_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X28 VGND a_580_119# a_1141_125# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X29 a_1248_151# a_111_156# a_1331_151# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X30 a_708_93# SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X31 VPWR a_580_119# a_1259_449# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X32 a_161_21# a_111_156# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X33 a_964_169# SET_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
