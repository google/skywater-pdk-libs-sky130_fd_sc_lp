* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__iso1p_lp2 A SLEEP KAPWR VGND VNB VPB VPWR X
X0 a_137_409# A a_240_409# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X1 VGND A a_147_57# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 VGND a_137_409# a_469_57# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 a_147_57# A a_137_409# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 a_137_409# SLEEP a_311_57# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 a_240_409# SLEEP KAPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X6 a_469_57# a_137_409# X VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 KAPWR a_137_409# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X8 a_311_57# SLEEP VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
