* File: sky130_fd_sc_lp__a22o_2.spice
* Created: Fri Aug 28 09:54:07 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__a22o_2.pex.spice"
.subckt sky130_fd_sc_lp__a22o_2  VNB VPB A2 A1 B2 B1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* B1	B1
* B2	B2
* A1	A1
* A2	A2
* VPB	VPB
* VNB	VNB
MM1001 N_X_M1001_d N_A_94_249#_M1001_g N_VGND_M1001_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.315 PD=1.12 PS=2.43 NRD=0 NRS=15.708 M=1 R=5.6 SA=75000.3
+ SB=75001.6 A=0.126 P=1.98 MULT=1
MM1002 N_X_M1001_d N_A_94_249#_M1002_g N_VGND_M1002_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1785 PD=1.12 PS=1.265 NRD=0 NRS=11.424 M=1 R=5.6 SA=75000.7
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1005 A_340_49# N_A2_M1005_g N_VGND_M1002_s VNB NSHORT L=0.15 W=0.84 AD=0.0882
+ AS=0.1785 PD=1.05 PS=1.265 NRD=7.14 NRS=9.276 M=1 R=5.6 SA=75001.3 SB=75000.6
+ A=0.126 P=1.98 MULT=1
MM1000 N_A_94_249#_M1000_d N_A1_M1000_g A_340_49# VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.0882 PD=2.21 PS=1.05 NRD=0 NRS=7.14 M=1 R=5.6 SA=75001.7
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1006 A_610_49# N_B2_M1006_g N_VGND_M1006_s VNB NSHORT L=0.15 W=0.84 AD=0.0882
+ AS=0.2394 PD=1.05 PS=2.25 NRD=7.14 NRS=0 M=1 R=5.6 SA=75000.2 SB=75000.6
+ A=0.126 P=1.98 MULT=1
MM1007 N_A_94_249#_M1007_d N_B1_M1007_g A_610_49# VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.0882 PD=2.21 PS=1.05 NRD=0 NRS=7.14 M=1 R=5.6 SA=75000.6
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1008 N_X_M1008_d N_A_94_249#_M1008_g N_VPWR_M1008_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75001.6 A=0.189 P=2.82 MULT=1
MM1011 N_X_M1008_d N_A_94_249#_M1011_g N_VPWR_M1011_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.2709 PD=1.54 PS=1.69 NRD=0 NRS=11.7215 M=1 R=8.4 SA=75000.6
+ SB=75001.2 A=0.189 P=2.82 MULT=1
MM1009 N_A_326_367#_M1009_d N_A2_M1009_g N_VPWR_M1011_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.2709 PD=1.54 PS=1.69 NRD=0 NRS=11.7215 M=1 R=8.4
+ SA=75001.2 SB=75000.6 A=0.189 P=2.82 MULT=1
MM1003 N_VPWR_M1003_d N_A1_M1003_g N_A_326_367#_M1009_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.6
+ SB=75000.2 A=0.189 P=2.82 MULT=1
MM1010 N_A_326_367#_M1010_d N_B2_M1010_g N_A_94_249#_M1010_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1004 N_A_94_249#_M1004_d N_B1_M1004_g N_A_326_367#_M1010_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX12_noxref VNB VPB NWDIODE A=7.8703 P=12.17
*
.include "sky130_fd_sc_lp__a22o_2.pxi.spice"
*
.ends
*
*
