* NGSPICE file created from sky130_fd_sc_lp__a211oi_1.ext - technology: sky130A

.subckt sky130_fd_sc_lp__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
M1000 a_27_367# A1 VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=8.253e+11p pd=6.35e+06u as=4.914e+11p ps=3.3e+06u
M1001 VGND B1 Y VNB nshort w=840000u l=150000u
+  ad=5.502e+11p pd=4.67e+06u as=5.502e+11p ps=4.67e+06u
M1002 a_110_49# A2 VGND VNB nshort w=840000u l=150000u
+  ad=1.764e+11p pd=2.1e+06u as=0p ps=0u
M1003 a_326_367# B1 a_27_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=2.646e+11p pd=2.94e+06u as=0p ps=0u
M1004 Y C1 a_326_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=3.339e+11p pd=3.05e+06u as=0p ps=0u
M1005 Y C1 VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR A2 a_27_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 Y A1 a_110_49# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

