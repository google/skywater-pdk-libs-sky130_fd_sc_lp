* File: sky130_fd_sc_lp__nand3_2.spice
* Created: Wed Sep  2 10:04:16 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__nand3_2.pex.spice"
.subckt sky130_fd_sc_lp__nand3_2  VNB VPB A B C VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* C	C
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1009 N_Y_M1009_d N_A_M1009_g N_A_43_65#_M1009_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75002.5 A=0.126 P=1.98 MULT=1
MM1010 N_Y_M1009_d N_A_M1010_g N_A_43_65#_M1010_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75002.1 A=0.126 P=1.98 MULT=1
MM1002 N_A_43_65#_M1010_s N_B_M1002_g N_A_298_65#_M1002_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1344 PD=1.12 PS=1.16 NRD=0 NRS=2.856 M=1 R=5.6
+ SA=75001.1 SB=75001.6 A=0.126 P=1.98 MULT=1
MM1000 N_VGND_M1000_d N_C_M1000_g N_A_298_65#_M1002_s VNB NSHORT L=0.15 W=0.84
+ AD=0.168 AS=0.1344 PD=1.24 PS=1.16 NRD=7.14 NRS=2.856 M=1 R=5.6 SA=75001.5
+ SB=75001.2 A=0.126 P=1.98 MULT=1
MM1007 N_VGND_M1000_d N_C_M1007_g N_A_298_65#_M1007_s VNB NSHORT L=0.15 W=0.84
+ AD=0.168 AS=0.1176 PD=1.24 PS=1.12 NRD=9.996 NRS=0 M=1 R=5.6 SA=75002.1
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1003 N_A_43_65#_M1003_d N_B_M1003_g N_A_298_65#_M1007_s VNB NSHORT L=0.15
+ W=0.84 AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002.5
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1004 N_Y_M1004_d N_A_M1004_g N_VPWR_M1004_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75002.4 A=0.189 P=2.82 MULT=1
MM1008 N_Y_M1004_d N_A_M1008_g N_VPWR_M1008_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.2016 PD=1.54 PS=1.58 NRD=0 NRS=3.1126 M=1 R=8.4 SA=75000.6
+ SB=75002 A=0.189 P=2.82 MULT=1
MM1005 N_VPWR_M1008_s N_B_M1005_g N_Y_M1005_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.2016 AS=0.1764 PD=1.58 PS=1.54 NRD=3.1126 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75001.5 A=0.189 P=2.82 MULT=1
MM1001 N_VPWR_M1001_d N_C_M1001_g N_Y_M1005_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.2079 AS=0.1764 PD=1.59 PS=1.54 NRD=3.1126 NRS=0 M=1 R=8.4 SA=75001.5
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1011 N_VPWR_M1001_d N_C_M1011_g N_Y_M1011_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.2079 AS=0.1764 PD=1.59 PS=1.54 NRD=4.6886 NRS=0 M=1 R=8.4 SA=75002
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1006 N_VPWR_M1006_d N_B_M1006_g N_Y_M1011_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.4
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX12_noxref VNB VPB NWDIODE A=6.9751 P=11.21
c_35 VNB 0 5.23255e-20 $X=0 $Y=0
*
.include "sky130_fd_sc_lp__nand3_2.pxi.spice"
*
.ends
*
*
