* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__sdlclkp_lp CLK GATE SCE VGND VNB VPB VPWR GCLK
X0 VPWR a_1384_416# GCLK VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X1 a_114_101# GATE a_93_376# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 a_93_376# GATE a_200_376# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X3 a_1016_47# a_698_405# a_860_21# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 a_804_405# a_860_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X5 a_1384_416# a_860_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X6 a_278_101# SCE VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 a_436_101# a_356_278# a_447_376# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 VPWR a_698_405# a_860_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X9 VGND CLK a_1392_192# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 a_698_405# a_356_278# a_804_405# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X11 VPWR CLK a_1384_416# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X12 a_812_47# a_860_21# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X13 a_93_376# a_447_376# a_698_405# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X14 a_356_278# CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X15 a_1392_192# a_860_21# a_1384_416# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X16 a_1548_48# a_1384_416# GCLK VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X17 a_356_278# CLK a_1234_192# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X18 a_93_376# a_356_278# a_698_405# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X19 VGND GATE a_114_101# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X20 a_698_405# a_447_376# a_812_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X21 VGND a_1384_416# a_1548_48# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X22 a_93_376# SCE a_278_101# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X23 VGND a_356_278# a_436_101# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X24 VGND a_698_405# a_1016_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X25 a_200_376# SCE VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X26 VPWR a_356_278# a_447_376# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X27 a_1234_192# CLK VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
