* File: sky130_fd_sc_lp__sdfrtp_1.pxi.spice
* Created: Wed Sep  2 10:34:35 2020
* 
x_PM_SKY130_FD_SC_LP__SDFRTP_1%A_35_74# N_A_35_74#_M1026_s N_A_35_74#_M1021_s
+ N_A_35_74#_c_268_n N_A_35_74#_M1006_g N_A_35_74#_M1015_g N_A_35_74#_c_269_n
+ N_A_35_74#_c_270_n N_A_35_74#_c_271_n N_A_35_74#_c_272_n N_A_35_74#_c_276_n
+ N_A_35_74#_c_273_n N_A_35_74#_c_277_n N_A_35_74#_c_278_n N_A_35_74#_c_279_n
+ PM_SKY130_FD_SC_LP__SDFRTP_1%A_35_74#
x_PM_SKY130_FD_SC_LP__SDFRTP_1%SCE N_SCE_M1026_g N_SCE_c_342_n N_SCE_c_348_n
+ N_SCE_c_349_n N_SCE_M1021_g N_SCE_c_351_n N_SCE_M1001_g N_SCE_M1038_g
+ N_SCE_c_353_n SCE SCE SCE SCE SCE N_SCE_c_345_n N_SCE_c_346_n
+ PM_SKY130_FD_SC_LP__SDFRTP_1%SCE
x_PM_SKY130_FD_SC_LP__SDFRTP_1%D N_D_M1033_g N_D_M1028_g D D D D N_D_c_414_n
+ PM_SKY130_FD_SC_LP__SDFRTP_1%D
x_PM_SKY130_FD_SC_LP__SDFRTP_1%SCD N_SCD_M1000_g N_SCD_M1008_g N_SCD_c_448_n
+ N_SCD_c_452_n SCD SCD SCD N_SCD_c_450_n PM_SKY130_FD_SC_LP__SDFRTP_1%SCD
x_PM_SKY130_FD_SC_LP__SDFRTP_1%A_757_317# N_A_757_317#_M1010_s
+ N_A_757_317#_M1035_s N_A_757_317#_M1019_g N_A_757_317#_M1034_g
+ N_A_757_317#_c_493_n N_A_757_317#_M1004_g N_A_757_317#_M1022_g
+ N_A_757_317#_c_494_n N_A_757_317#_c_495_n N_A_757_317#_c_512_n
+ N_A_757_317#_c_513_n N_A_757_317#_c_496_n N_A_757_317#_c_497_n
+ N_A_757_317#_c_498_n N_A_757_317#_c_499_n N_A_757_317#_c_500_n
+ N_A_757_317#_c_501_n N_A_757_317#_c_631_p N_A_757_317#_c_502_n
+ N_A_757_317#_c_503_n N_A_757_317#_c_504_n N_A_757_317#_c_505_n
+ N_A_757_317#_c_506_n N_A_757_317#_c_507_n N_A_757_317#_c_508_n
+ PM_SKY130_FD_SC_LP__SDFRTP_1%A_757_317#
x_PM_SKY130_FD_SC_LP__SDFRTP_1%A_937_333# N_A_937_333#_M1030_d
+ N_A_937_333#_M1029_d N_A_937_333#_M1002_g N_A_937_333#_c_706_n
+ N_A_937_333#_M1011_g N_A_937_333#_c_700_n N_A_937_333#_c_701_n
+ N_A_937_333#_c_702_n N_A_937_333#_c_703_n N_A_937_333#_c_709_n
+ N_A_937_333#_c_747_p N_A_937_333#_c_728_n N_A_937_333#_c_704_n
+ N_A_937_333#_c_733_n N_A_937_333#_c_758_p N_A_937_333#_c_711_n
+ PM_SKY130_FD_SC_LP__SDFRTP_1%A_937_333#
x_PM_SKY130_FD_SC_LP__SDFRTP_1%RESET_B N_RESET_B_M1027_g N_RESET_B_M1025_g
+ N_RESET_B_c_798_n N_RESET_B_c_799_n N_RESET_B_c_800_n N_RESET_B_c_801_n
+ N_RESET_B_c_802_n N_RESET_B_c_803_n N_RESET_B_c_810_n N_RESET_B_M1013_g
+ N_RESET_B_c_811_n N_RESET_B_c_812_n N_RESET_B_M1036_g N_RESET_B_M1005_g
+ N_RESET_B_M1023_g N_RESET_B_c_806_n N_RESET_B_c_816_n N_RESET_B_c_807_n
+ N_RESET_B_c_808_n N_RESET_B_c_817_n N_RESET_B_c_818_n N_RESET_B_c_819_n
+ N_RESET_B_c_820_n N_RESET_B_c_821_n N_RESET_B_c_822_n N_RESET_B_c_823_n
+ N_RESET_B_c_824_n RESET_B RESET_B N_RESET_B_c_826_n N_RESET_B_c_809_n
+ N_RESET_B_c_828_n PM_SKY130_FD_SC_LP__SDFRTP_1%RESET_B
x_PM_SKY130_FD_SC_LP__SDFRTP_1%A_809_463# N_A_809_463#_M1032_d
+ N_A_809_463#_M1019_d N_A_809_463#_M1013_d N_A_809_463#_M1030_g
+ N_A_809_463#_M1029_g N_A_809_463#_c_1010_n N_A_809_463#_c_1011_n
+ N_A_809_463#_c_1072_n N_A_809_463#_c_1016_n N_A_809_463#_c_1055_n
+ N_A_809_463#_c_1012_n N_A_809_463#_c_1017_n N_A_809_463#_c_1013_n
+ PM_SKY130_FD_SC_LP__SDFRTP_1%A_809_463#
x_PM_SKY130_FD_SC_LP__SDFRTP_1%A_865_255# N_A_865_255#_M1007_d
+ N_A_865_255#_M1018_d N_A_865_255#_M1037_g N_A_865_255#_M1032_g
+ N_A_865_255#_c_1139_n N_A_865_255#_c_1140_n N_A_865_255#_M1017_g
+ N_A_865_255#_c_1125_n N_A_865_255#_c_1126_n N_A_865_255#_M1012_g
+ N_A_865_255#_M1010_g N_A_865_255#_M1035_g N_A_865_255#_c_1129_n
+ N_A_865_255#_c_1130_n N_A_865_255#_c_1131_n N_A_865_255#_c_1147_n
+ N_A_865_255#_c_1148_n N_A_865_255#_c_1149_n N_A_865_255#_c_1150_n
+ N_A_865_255#_c_1132_n N_A_865_255#_c_1133_n N_A_865_255#_c_1134_n
+ N_A_865_255#_c_1135_n N_A_865_255#_c_1136_n N_A_865_255#_c_1154_n
+ N_A_865_255#_c_1137_n PM_SKY130_FD_SC_LP__SDFRTP_1%A_865_255#
x_PM_SKY130_FD_SC_LP__SDFRTP_1%A_1445_69# N_A_1445_69#_M1004_d
+ N_A_1445_69#_M1017_d N_A_1445_69#_c_1324_n N_A_1445_69#_M1009_g
+ N_A_1445_69#_M1014_g N_A_1445_69#_M1003_g N_A_1445_69#_M1039_g
+ N_A_1445_69#_c_1328_n N_A_1445_69#_c_1329_n N_A_1445_69#_c_1330_n
+ N_A_1445_69#_c_1331_n N_A_1445_69#_c_1332_n N_A_1445_69#_c_1347_n
+ N_A_1445_69#_c_1363_n N_A_1445_69#_c_1365_n N_A_1445_69#_c_1333_n
+ N_A_1445_69#_c_1334_n N_A_1445_69#_c_1335_n N_A_1445_69#_c_1336_n
+ N_A_1445_69#_c_1337_n N_A_1445_69#_c_1338_n N_A_1445_69#_c_1339_n
+ N_A_1445_69#_c_1340_n N_A_1445_69#_c_1341_n N_A_1445_69#_c_1342_n
+ N_A_1445_69#_c_1343_n PM_SKY130_FD_SC_LP__SDFRTP_1%A_1445_69#
x_PM_SKY130_FD_SC_LP__SDFRTP_1%A_1641_21# N_A_1641_21#_M1009_d
+ N_A_1641_21#_M1023_d N_A_1641_21#_M1020_g N_A_1641_21#_M1031_g
+ N_A_1641_21#_c_1529_n N_A_1641_21#_c_1530_n N_A_1641_21#_c_1531_n
+ N_A_1641_21#_c_1532_n N_A_1641_21#_c_1533_n N_A_1641_21#_c_1540_n
+ N_A_1641_21#_c_1534_n N_A_1641_21#_c_1535_n N_A_1641_21#_c_1536_n
+ N_A_1641_21#_c_1541_n N_A_1641_21#_c_1613_n N_A_1641_21#_c_1542_n
+ N_A_1641_21#_c_1543_n N_A_1641_21#_c_1537_n
+ PM_SKY130_FD_SC_LP__SDFRTP_1%A_1641_21#
x_PM_SKY130_FD_SC_LP__SDFRTP_1%CLK N_CLK_M1007_g N_CLK_M1018_g N_CLK_c_1643_n
+ N_CLK_c_1644_n CLK CLK CLK N_CLK_c_1645_n N_CLK_c_1648_n
+ PM_SKY130_FD_SC_LP__SDFRTP_1%CLK
x_PM_SKY130_FD_SC_LP__SDFRTP_1%A_2408_367# N_A_2408_367#_M1039_s
+ N_A_2408_367#_M1003_s N_A_2408_367#_M1016_g N_A_2408_367#_M1024_g
+ N_A_2408_367#_c_1692_n N_A_2408_367#_c_1699_n N_A_2408_367#_c_1693_n
+ N_A_2408_367#_c_1694_n N_A_2408_367#_c_1687_n N_A_2408_367#_c_1688_n
+ N_A_2408_367#_c_1689_n N_A_2408_367#_c_1690_n
+ PM_SKY130_FD_SC_LP__SDFRTP_1%A_2408_367#
x_PM_SKY130_FD_SC_LP__SDFRTP_1%VPWR N_VPWR_M1021_d N_VPWR_M1008_d N_VPWR_M1002_d
+ N_VPWR_M1029_s N_VPWR_M1031_d N_VPWR_M1014_d N_VPWR_M1035_d N_VPWR_M1003_d
+ N_VPWR_c_1743_n N_VPWR_c_1744_n N_VPWR_c_1745_n N_VPWR_c_1746_n
+ N_VPWR_c_1747_n N_VPWR_c_1748_n N_VPWR_c_1749_n N_VPWR_c_1750_n
+ N_VPWR_c_1751_n N_VPWR_c_1752_n VPWR N_VPWR_c_1753_n N_VPWR_c_1754_n
+ N_VPWR_c_1755_n N_VPWR_c_1756_n N_VPWR_c_1757_n N_VPWR_c_1758_n
+ N_VPWR_c_1742_n N_VPWR_c_1760_n N_VPWR_c_1761_n N_VPWR_c_1762_n
+ N_VPWR_c_1763_n N_VPWR_c_1764_n N_VPWR_c_1765_n N_VPWR_c_1766_n
+ N_VPWR_c_1767_n PM_SKY130_FD_SC_LP__SDFRTP_1%VPWR
x_PM_SKY130_FD_SC_LP__SDFRTP_1%A_380_50# N_A_380_50#_M1033_d N_A_380_50#_M1032_s
+ N_A_380_50#_M1028_d N_A_380_50#_M1025_d N_A_380_50#_c_1892_n
+ N_A_380_50#_c_1899_n N_A_380_50#_c_1893_n N_A_380_50#_c_1894_n
+ N_A_380_50#_c_1895_n N_A_380_50#_c_1897_n N_A_380_50#_c_1949_n
+ N_A_380_50#_c_1898_n N_A_380_50#_c_1936_n
+ PM_SKY130_FD_SC_LP__SDFRTP_1%A_380_50#
x_PM_SKY130_FD_SC_LP__SDFRTP_1%Q N_Q_M1016_d N_Q_M1024_d Q Q Q Q Q Q
+ N_Q_c_1994_n PM_SKY130_FD_SC_LP__SDFRTP_1%Q
x_PM_SKY130_FD_SC_LP__SDFRTP_1%VGND N_VGND_M1026_d N_VGND_M1027_d N_VGND_M1036_d
+ N_VGND_M1020_d N_VGND_M1010_d N_VGND_M1039_d N_VGND_c_2005_n N_VGND_c_2006_n
+ N_VGND_c_2007_n N_VGND_c_2008_n N_VGND_c_2009_n N_VGND_c_2010_n
+ N_VGND_c_2011_n N_VGND_c_2012_n N_VGND_c_2013_n N_VGND_c_2014_n VGND
+ N_VGND_c_2015_n N_VGND_c_2016_n N_VGND_c_2017_n N_VGND_c_2018_n
+ N_VGND_c_2019_n N_VGND_c_2020_n N_VGND_c_2021_n N_VGND_c_2022_n
+ N_VGND_c_2023_n N_VGND_c_2024_n PM_SKY130_FD_SC_LP__SDFRTP_1%VGND
x_PM_SKY130_FD_SC_LP__SDFRTP_1%noxref_24 N_noxref_24_M1006_s N_noxref_24_M1000_d
+ N_noxref_24_c_2144_n N_noxref_24_c_2148_n N_noxref_24_c_2145_n
+ PM_SKY130_FD_SC_LP__SDFRTP_1%noxref_24
cc_1 VNB N_A_35_74#_c_268_n 0.0212422f $X=-0.19 $Y=-0.245 $X2=1.465 $Y2=0.78
cc_2 VNB N_A_35_74#_c_269_n 0.0196756f $X=-0.19 $Y=-0.245 $X2=0.3 $Y2=0.58
cc_3 VNB N_A_35_74#_c_270_n 0.0334154f $X=-0.19 $Y=-0.245 $X2=0.23 $Y2=1.975
cc_4 VNB N_A_35_74#_c_271_n 0.0147265f $X=-0.19 $Y=-0.245 $X2=1.345 $Y2=0.945
cc_5 VNB N_A_35_74#_c_272_n 0.0396124f $X=-0.19 $Y=-0.245 $X2=1.345 $Y2=0.945
cc_6 VNB N_A_35_74#_c_273_n 0.0103663f $X=-0.19 $Y=-0.245 $X2=0.26 $Y2=0.945
cc_7 VNB N_SCE_M1026_g 0.0388402f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_SCE_c_342_n 0.0337585f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_SCE_M1038_g 0.0262093f $X=-0.19 $Y=-0.245 $X2=1.345 $Y2=0.945
cc_10 VNB SCE 0.0371674f $X=-0.19 $Y=-0.245 $X2=0.23 $Y2=2.47
cc_11 VNB N_SCE_c_345_n 0.0343692f $X=-0.19 $Y=-0.245 $X2=2.51 $Y2=1.98
cc_12 VNB N_SCE_c_346_n 0.0348128f $X=-0.19 $Y=-0.245 $X2=1.465 $Y2=0.945
cc_13 VNB N_D_M1033_g 0.0636509f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB D 0.011249f $X=-0.19 $Y=-0.245 $X2=2.49 $Y2=2.635
cc_15 VNB N_D_c_414_n 0.0269442f $X=-0.19 $Y=-0.245 $X2=0.23 $Y2=1.03
cc_16 VNB N_SCD_M1000_g 0.0281694f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_SCD_c_448_n 0.0246895f $X=-0.19 $Y=-0.245 $X2=2.49 $Y2=2.635
cc_18 VNB SCD 0.00606287f $X=-0.19 $Y=-0.245 $X2=0.26 $Y2=0.86
cc_19 VNB N_SCD_c_450_n 0.0260714f $X=-0.19 $Y=-0.245 $X2=1.345 $Y2=0.945
cc_20 VNB N_A_757_317#_c_493_n 0.0673991f $X=-0.19 $Y=-0.245 $X2=0.26 $Y2=0.86
cc_21 VNB N_A_757_317#_c_494_n 0.00320236f $X=-0.19 $Y=-0.245 $X2=1.345
+ $Y2=0.945
cc_22 VNB N_A_757_317#_c_495_n 0.00402985f $X=-0.19 $Y=-0.245 $X2=1.345
+ $Y2=0.945
cc_23 VNB N_A_757_317#_c_496_n 0.00235833f $X=-0.19 $Y=-0.245 $X2=1.15 $Y2=2.47
cc_24 VNB N_A_757_317#_c_497_n 0.0154208f $X=-0.19 $Y=-0.245 $X2=2.51 $Y2=1.98
cc_25 VNB N_A_757_317#_c_498_n 0.00147433f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_757_317#_c_499_n 0.0200417f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_757_317#_c_500_n 0.00221522f $X=-0.19 $Y=-0.245 $X2=1.345
+ $Y2=0.945
cc_28 VNB N_A_757_317#_c_501_n 0.0156731f $X=-0.19 $Y=-0.245 $X2=1.465 $Y2=0.945
cc_29 VNB N_A_757_317#_c_502_n 0.00766905f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_757_317#_c_503_n 0.00276218f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_757_317#_c_504_n 0.0114317f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_757_317#_c_505_n 0.0118801f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_757_317#_c_506_n 0.0289705f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_757_317#_c_507_n 0.00541985f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_757_317#_c_508_n 0.0158609f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_937_333#_M1011_g 0.0240061f $X=-0.19 $Y=-0.245 $X2=0.26 $Y2=0.58
cc_37 VNB N_A_937_333#_c_700_n 0.0167487f $X=-0.19 $Y=-0.245 $X2=0.23 $Y2=1.03
cc_38 VNB N_A_937_333#_c_701_n 0.0088579f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=0.945
cc_39 VNB N_A_937_333#_c_702_n 0.0093328f $X=-0.19 $Y=-0.245 $X2=1.345 $Y2=0.945
cc_40 VNB N_A_937_333#_c_703_n 0.00775597f $X=-0.19 $Y=-0.245 $X2=1.15 $Y2=2.06
cc_41 VNB N_A_937_333#_c_704_n 0.00196286f $X=-0.19 $Y=-0.245 $X2=2.55 $Y2=1.98
cc_42 VNB N_RESET_B_M1027_g 0.0191999f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_RESET_B_c_798_n 0.0223657f $X=-0.19 $Y=-0.245 $X2=1.465 $Y2=0.46
cc_44 VNB N_RESET_B_c_799_n 0.012806f $X=-0.19 $Y=-0.245 $X2=1.465 $Y2=0.46
cc_45 VNB N_RESET_B_c_800_n 0.0232079f $X=-0.19 $Y=-0.245 $X2=2.49 $Y2=2.635
cc_46 VNB N_RESET_B_c_801_n 0.00905619f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_RESET_B_c_802_n 0.0579791f $X=-0.19 $Y=-0.245 $X2=0.26 $Y2=0.58
cc_48 VNB N_RESET_B_c_803_n 0.150151f $X=-0.19 $Y=-0.245 $X2=0.3 $Y2=0.58
cc_49 VNB N_RESET_B_M1036_g 0.0318232f $X=-0.19 $Y=-0.245 $X2=0.23 $Y2=2.47
cc_50 VNB N_RESET_B_M1005_g 0.0418154f $X=-0.19 $Y=-0.245 $X2=1.055 $Y2=2.46
cc_51 VNB N_RESET_B_c_806_n 0.0174786f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_RESET_B_c_807_n 0.00749069f $X=-0.19 $Y=-0.245 $X2=1.465 $Y2=0.945
cc_53 VNB N_RESET_B_c_808_n 0.0104803f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_RESET_B_c_809_n 0.0203079f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_809_463#_M1030_g 0.0240625f $X=-0.19 $Y=-0.245 $X2=2.49 $Y2=2.635
cc_56 VNB N_A_809_463#_M1029_g 0.00120569f $X=-0.19 $Y=-0.245 $X2=0.3 $Y2=0.58
cc_57 VNB N_A_809_463#_c_1010_n 0.00842474f $X=-0.19 $Y=-0.245 $X2=0.23
+ $Y2=1.975
cc_58 VNB N_A_809_463#_c_1011_n 0.0037754f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=0.945
cc_59 VNB N_A_809_463#_c_1012_n 0.00186512f $X=-0.19 $Y=-0.245 $X2=1.15 $Y2=2.47
cc_60 VNB N_A_809_463#_c_1013_n 0.0768283f $X=-0.19 $Y=-0.245 $X2=1.465
+ $Y2=0.945
cc_61 VNB N_A_865_255#_M1037_g 0.0142822f $X=-0.19 $Y=-0.245 $X2=2.49 $Y2=2.145
cc_62 VNB N_A_865_255#_M1032_g 0.0236551f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_A_865_255#_c_1125_n 0.00970066f $X=-0.19 $Y=-0.245 $X2=1.345
+ $Y2=0.945
cc_64 VNB N_A_865_255#_c_1126_n 0.00316727f $X=-0.19 $Y=-0.245 $X2=1.345
+ $Y2=0.945
cc_65 VNB N_A_865_255#_M1012_g 0.0403327f $X=-0.19 $Y=-0.245 $X2=2.425 $Y2=2.06
cc_66 VNB N_A_865_255#_M1010_g 0.022001f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_A_865_255#_c_1129_n 0.011132f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_A_865_255#_c_1130_n 0.0078841f $X=-0.19 $Y=-0.245 $X2=1.345
+ $Y2=0.945
cc_69 VNB N_A_865_255#_c_1131_n 0.0101702f $X=-0.19 $Y=-0.245 $X2=1.465
+ $Y2=0.945
cc_70 VNB N_A_865_255#_c_1132_n 0.0173687f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_A_865_255#_c_1133_n 7.18436e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_A_865_255#_c_1134_n 0.00803792f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_A_865_255#_c_1135_n 0.0317378f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_A_865_255#_c_1136_n 0.00477428f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_A_865_255#_c_1137_n 0.00198139f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_A_1445_69#_c_1324_n 0.0160971f $X=-0.19 $Y=-0.245 $X2=1.465 $Y2=0.78
cc_77 VNB N_A_1445_69#_M1014_g 0.0134434f $X=-0.19 $Y=-0.245 $X2=2.49 $Y2=2.635
cc_78 VNB N_A_1445_69#_M1003_g 0.00403029f $X=-0.19 $Y=-0.245 $X2=0.3 $Y2=0.58
cc_79 VNB N_A_1445_69#_M1039_g 0.0297229f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=0.945
cc_80 VNB N_A_1445_69#_c_1328_n 0.0235788f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_A_1445_69#_c_1329_n 0.016002f $X=-0.19 $Y=-0.245 $X2=1.15 $Y2=2.06
cc_82 VNB N_A_1445_69#_c_1330_n 0.00747602f $X=-0.19 $Y=-0.245 $X2=0.23 $Y2=2.47
cc_83 VNB N_A_1445_69#_c_1331_n 0.0059897f $X=-0.19 $Y=-0.245 $X2=1.055 $Y2=2.46
cc_84 VNB N_A_1445_69#_c_1332_n 0.00249583f $X=-0.19 $Y=-0.245 $X2=2.55 $Y2=1.98
cc_85 VNB N_A_1445_69#_c_1333_n 0.00127275f $X=-0.19 $Y=-0.245 $X2=2.51
+ $Y2=2.145
cc_86 VNB N_A_1445_69#_c_1334_n 0.00154969f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_A_1445_69#_c_1335_n 0.00791001f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_A_1445_69#_c_1336_n 0.0166602f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_A_1445_69#_c_1337_n 0.00311823f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_A_1445_69#_c_1338_n 0.00522363f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_A_1445_69#_c_1339_n 0.0481702f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_A_1445_69#_c_1340_n 0.0162262f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_93 VNB N_A_1445_69#_c_1341_n 0.00619485f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_94 VNB N_A_1445_69#_c_1342_n 0.0159329f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_95 VNB N_A_1445_69#_c_1343_n 0.0325072f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_96 VNB N_A_1641_21#_M1020_g 0.0232098f $X=-0.19 $Y=-0.245 $X2=2.49 $Y2=2.145
cc_97 VNB N_A_1641_21#_c_1529_n 0.111065f $X=-0.19 $Y=-0.245 $X2=0.26 $Y2=0.58
cc_98 VNB N_A_1641_21#_c_1530_n 0.012806f $X=-0.19 $Y=-0.245 $X2=0.3 $Y2=0.58
cc_99 VNB N_A_1641_21#_c_1531_n 0.0260094f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_100 VNB N_A_1641_21#_c_1532_n 0.00562617f $X=-0.19 $Y=-0.245 $X2=0.23
+ $Y2=1.03
cc_101 VNB N_A_1641_21#_c_1533_n 0.0181522f $X=-0.19 $Y=-0.245 $X2=0.43
+ $Y2=0.945
cc_102 VNB N_A_1641_21#_c_1534_n 0.00337432f $X=-0.19 $Y=-0.245 $X2=2.425
+ $Y2=2.06
cc_103 VNB N_A_1641_21#_c_1535_n 0.00380415f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_104 VNB N_A_1641_21#_c_1536_n 0.00482238f $X=-0.19 $Y=-0.245 $X2=1.055
+ $Y2=2.46
cc_105 VNB N_A_1641_21#_c_1537_n 0.0506687f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_106 VNB N_CLK_M1007_g 0.0260597f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_107 VNB N_CLK_M1018_g 0.00586985f $X=-0.19 $Y=-0.245 $X2=1.465 $Y2=0.78
cc_108 VNB N_CLK_c_1643_n 0.0183597f $X=-0.19 $Y=-0.245 $X2=1.465 $Y2=0.46
cc_109 VNB N_CLK_c_1644_n 0.00391068f $X=-0.19 $Y=-0.245 $X2=2.49 $Y2=2.635
cc_110 VNB N_CLK_c_1645_n 0.0286132f $X=-0.19 $Y=-0.245 $X2=0.23 $Y2=1.03
cc_111 VNB N_A_2408_367#_M1016_g 0.026228f $X=-0.19 $Y=-0.245 $X2=1.465 $Y2=0.46
cc_112 VNB N_A_2408_367#_M1024_g 0.00105913f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_113 VNB N_A_2408_367#_c_1687_n 0.00377889f $X=-0.19 $Y=-0.245 $X2=2.425
+ $Y2=2.06
cc_114 VNB N_A_2408_367#_c_1688_n 0.00314278f $X=-0.19 $Y=-0.245 $X2=1.15
+ $Y2=2.06
cc_115 VNB N_A_2408_367#_c_1689_n 0.00179584f $X=-0.19 $Y=-0.245 $X2=1.055
+ $Y2=2.47
cc_116 VNB N_A_2408_367#_c_1690_n 0.0391508f $X=-0.19 $Y=-0.245 $X2=1.055
+ $Y2=2.46
cc_117 VNB N_VPWR_c_1742_n 0.561729f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_118 VNB N_A_380_50#_c_1892_n 0.010443f $X=-0.19 $Y=-0.245 $X2=0.26 $Y2=0.58
cc_119 VNB N_A_380_50#_c_1893_n 0.00710712f $X=-0.19 $Y=-0.245 $X2=0.43
+ $Y2=0.945
cc_120 VNB N_A_380_50#_c_1894_n 0.0037567f $X=-0.19 $Y=-0.245 $X2=1.345
+ $Y2=0.945
cc_121 VNB N_A_380_50#_c_1895_n 0.00754278f $X=-0.19 $Y=-0.245 $X2=1.15 $Y2=2.06
cc_122 VNB N_Q_c_1994_n 0.0616899f $X=-0.19 $Y=-0.245 $X2=0.43 $Y2=0.945
cc_123 VNB N_VGND_c_2005_n 0.0133739f $X=-0.19 $Y=-0.245 $X2=1.345 $Y2=0.945
cc_124 VNB N_VGND_c_2006_n 0.0081923f $X=-0.19 $Y=-0.245 $X2=2.425 $Y2=2.06
cc_125 VNB N_VGND_c_2007_n 0.00864254f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_126 VNB N_VGND_c_2008_n 0.0123546f $X=-0.19 $Y=-0.245 $X2=2.55 $Y2=1.98
cc_127 VNB N_VGND_c_2009_n 0.0086016f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_128 VNB N_VGND_c_2010_n 0.00284713f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_129 VNB N_VGND_c_2011_n 0.0747335f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_130 VNB N_VGND_c_2012_n 0.00594344f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_131 VNB N_VGND_c_2013_n 0.0536204f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_132 VNB N_VGND_c_2014_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_133 VNB N_VGND_c_2015_n 0.0189123f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_134 VNB N_VGND_c_2016_n 0.0596124f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_135 VNB N_VGND_c_2017_n 0.0507927f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_136 VNB N_VGND_c_2018_n 0.0404181f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_137 VNB N_VGND_c_2019_n 0.0152818f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_138 VNB N_VGND_c_2020_n 0.665682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_139 VNB N_VGND_c_2021_n 0.00567425f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_140 VNB N_VGND_c_2022_n 0.00437061f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_141 VNB N_VGND_c_2023_n 0.00631504f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_142 VNB N_VGND_c_2024_n 0.00529402f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_143 VNB N_noxref_24_c_2144_n 0.00433f $X=-0.19 $Y=-0.245 $X2=1.465 $Y2=0.78
cc_144 VNB N_noxref_24_c_2145_n 0.00389564f $X=-0.19 $Y=-0.245 $X2=0.26 $Y2=0.86
cc_145 VPB N_A_35_74#_M1015_g 0.0214579f $X=-0.19 $Y=1.655 $X2=2.49 $Y2=2.635
cc_146 VPB N_A_35_74#_c_270_n 0.0177161f $X=-0.19 $Y=1.655 $X2=0.23 $Y2=1.975
cc_147 VPB N_A_35_74#_c_276_n 0.0178423f $X=-0.19 $Y=1.655 $X2=2.425 $Y2=2.06
cc_148 VPB N_A_35_74#_c_277_n 0.0707236f $X=-0.19 $Y=1.655 $X2=1.15 $Y2=2.47
cc_149 VPB N_A_35_74#_c_278_n 0.00379253f $X=-0.19 $Y=1.655 $X2=2.51 $Y2=1.98
cc_150 VPB N_A_35_74#_c_279_n 0.0334861f $X=-0.19 $Y=1.655 $X2=2.51 $Y2=1.98
cc_151 VPB N_SCE_c_342_n 0.0429361f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_152 VPB N_SCE_c_348_n 0.0211321f $X=-0.19 $Y=1.655 $X2=1.465 $Y2=0.78
cc_153 VPB N_SCE_c_349_n 0.0253985f $X=-0.19 $Y=1.655 $X2=1.465 $Y2=0.46
cc_154 VPB N_SCE_M1021_g 0.021905f $X=-0.19 $Y=1.655 $X2=2.49 $Y2=2.635
cc_155 VPB N_SCE_c_351_n 0.0208673f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_156 VPB N_SCE_M1001_g 0.0174836f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_157 VPB N_SCE_c_353_n 0.00666874f $X=-0.19 $Y=1.655 $X2=1.345 $Y2=0.945
cc_158 VPB N_D_M1028_g 0.0396785f $X=-0.19 $Y=1.655 $X2=1.465 $Y2=0.78
cc_159 VPB D 0.0103884f $X=-0.19 $Y=1.655 $X2=2.49 $Y2=2.635
cc_160 VPB N_D_c_414_n 0.0294423f $X=-0.19 $Y=1.655 $X2=0.23 $Y2=1.03
cc_161 VPB N_SCD_M1008_g 0.0368956f $X=-0.19 $Y=1.655 $X2=1.465 $Y2=0.78
cc_162 VPB N_SCD_c_452_n 0.0177855f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_163 VPB SCD 0.00583342f $X=-0.19 $Y=1.655 $X2=0.26 $Y2=0.86
cc_164 VPB N_SCD_c_450_n 0.00188422f $X=-0.19 $Y=1.655 $X2=1.345 $Y2=0.945
cc_165 VPB N_A_757_317#_M1019_g 0.0329176f $X=-0.19 $Y=1.655 $X2=1.465 $Y2=0.46
cc_166 VPB N_A_757_317#_M1022_g 0.0304198f $X=-0.19 $Y=1.655 $X2=0.23 $Y2=1.975
cc_167 VPB N_A_757_317#_c_494_n 0.00549079f $X=-0.19 $Y=1.655 $X2=1.345
+ $Y2=0.945
cc_168 VPB N_A_757_317#_c_512_n 0.00181042f $X=-0.19 $Y=1.655 $X2=0.26 $Y2=0.945
cc_169 VPB N_A_757_317#_c_513_n 0.0379395f $X=-0.19 $Y=1.655 $X2=0.23 $Y2=2.47
cc_170 VPB N_A_757_317#_c_502_n 0.00471801f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_171 VPB N_A_757_317#_c_504_n 0.0095548f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_172 VPB N_A_757_317#_c_505_n 0.0218702f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_173 VPB N_A_937_333#_M1002_g 0.0268755f $X=-0.19 $Y=1.655 $X2=1.465 $Y2=0.46
cc_174 VPB N_A_937_333#_c_706_n 0.0255598f $X=-0.19 $Y=1.655 $X2=2.49 $Y2=2.635
cc_175 VPB N_A_937_333#_c_700_n 0.00185687f $X=-0.19 $Y=1.655 $X2=0.23 $Y2=1.03
cc_176 VPB N_A_937_333#_c_702_n 0.0119618f $X=-0.19 $Y=1.655 $X2=1.345 $Y2=0.945
cc_177 VPB N_A_937_333#_c_709_n 0.00384903f $X=-0.19 $Y=1.655 $X2=0.23 $Y2=2.47
cc_178 VPB N_A_937_333#_c_704_n 0.00174904f $X=-0.19 $Y=1.655 $X2=2.55 $Y2=1.98
cc_179 VPB N_A_937_333#_c_711_n 0.0348684f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_180 VPB N_RESET_B_c_810_n 0.0190796f $X=-0.19 $Y=1.655 $X2=0.23 $Y2=1.03
cc_181 VPB N_RESET_B_c_811_n 0.0213189f $X=-0.19 $Y=1.655 $X2=1.345 $Y2=0.945
cc_182 VPB N_RESET_B_c_812_n 0.00826772f $X=-0.19 $Y=1.655 $X2=1.345 $Y2=0.945
cc_183 VPB N_RESET_B_M1005_g 0.02749f $X=-0.19 $Y=1.655 $X2=1.055 $Y2=2.46
cc_184 VPB N_RESET_B_M1023_g 0.0213087f $X=-0.19 $Y=1.655 $X2=2.51 $Y2=1.98
cc_185 VPB N_RESET_B_c_806_n 0.0188514f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_186 VPB N_RESET_B_c_816_n 0.0347854f $X=-0.19 $Y=1.655 $X2=1.345 $Y2=0.945
cc_187 VPB N_RESET_B_c_817_n 0.00308581f $X=-0.19 $Y=1.655 $X2=2.51 $Y2=2.145
cc_188 VPB N_RESET_B_c_818_n 0.00199211f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_189 VPB N_RESET_B_c_819_n 0.00974949f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_190 VPB N_RESET_B_c_820_n 0.00177503f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_191 VPB N_RESET_B_c_821_n 4.13207e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_192 VPB N_RESET_B_c_822_n 0.0100613f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_193 VPB N_RESET_B_c_823_n 0.00488283f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_194 VPB N_RESET_B_c_824_n 0.00444283f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_195 VPB RESET_B 0.00301217f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_196 VPB N_RESET_B_c_826_n 0.0746688f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_197 VPB N_RESET_B_c_809_n 0.0161894f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_198 VPB N_RESET_B_c_828_n 0.0364626f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_199 VPB N_A_809_463#_M1029_g 0.0236856f $X=-0.19 $Y=1.655 $X2=0.3 $Y2=0.58
cc_200 VPB N_A_809_463#_c_1010_n 0.00287554f $X=-0.19 $Y=1.655 $X2=0.23
+ $Y2=1.975
cc_201 VPB N_A_809_463#_c_1016_n 0.00816459f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_202 VPB N_A_809_463#_c_1017_n 0.00667316f $X=-0.19 $Y=1.655 $X2=2.51 $Y2=1.98
cc_203 VPB N_A_865_255#_M1037_g 0.0513141f $X=-0.19 $Y=1.655 $X2=2.49 $Y2=2.145
cc_204 VPB N_A_865_255#_c_1139_n 0.20739f $X=-0.19 $Y=1.655 $X2=0.26 $Y2=0.58
cc_205 VPB N_A_865_255#_c_1140_n 0.012806f $X=-0.19 $Y=1.655 $X2=0.3 $Y2=0.58
cc_206 VPB N_A_865_255#_M1017_g 0.0272974f $X=-0.19 $Y=1.655 $X2=0.43 $Y2=0.945
cc_207 VPB N_A_865_255#_c_1125_n 0.0250775f $X=-0.19 $Y=1.655 $X2=1.345
+ $Y2=0.945
cc_208 VPB N_A_865_255#_c_1126_n 0.00379873f $X=-0.19 $Y=1.655 $X2=1.345
+ $Y2=0.945
cc_209 VPB N_A_865_255#_M1035_g 0.0225996f $X=-0.19 $Y=1.655 $X2=2.55 $Y2=1.98
cc_210 VPB N_A_865_255#_c_1130_n 0.00615094f $X=-0.19 $Y=1.655 $X2=1.345
+ $Y2=0.945
cc_211 VPB N_A_865_255#_c_1131_n 0.0110075f $X=-0.19 $Y=1.655 $X2=1.465
+ $Y2=0.945
cc_212 VPB N_A_865_255#_c_1147_n 0.0147975f $X=-0.19 $Y=1.655 $X2=2.51 $Y2=2.145
cc_213 VPB N_A_865_255#_c_1148_n 0.0131195f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_214 VPB N_A_865_255#_c_1149_n 0.00472322f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_215 VPB N_A_865_255#_c_1150_n 0.00146718f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_216 VPB N_A_865_255#_c_1132_n 0.0180207f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_217 VPB N_A_865_255#_c_1133_n 9.26678e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_218 VPB N_A_865_255#_c_1135_n 0.00948575f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_219 VPB N_A_865_255#_c_1154_n 0.0114992f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_220 VPB N_A_1445_69#_M1014_g 0.0728655f $X=-0.19 $Y=1.655 $X2=2.49 $Y2=2.635
cc_221 VPB N_A_1445_69#_M1003_g 0.0264637f $X=-0.19 $Y=1.655 $X2=0.3 $Y2=0.58
cc_222 VPB N_A_1445_69#_c_1332_n 0.00419055f $X=-0.19 $Y=1.655 $X2=2.55 $Y2=1.98
cc_223 VPB N_A_1445_69#_c_1347_n 0.00268862f $X=-0.19 $Y=1.655 $X2=2.51 $Y2=1.98
cc_224 VPB N_A_1641_21#_M1031_g 0.0295996f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_225 VPB N_A_1641_21#_c_1533_n 0.0181846f $X=-0.19 $Y=1.655 $X2=0.43 $Y2=0.945
cc_226 VPB N_A_1641_21#_c_1540_n 0.0137908f $X=-0.19 $Y=1.655 $X2=1.345
+ $Y2=0.945
cc_227 VPB N_A_1641_21#_c_1541_n 0.00682421f $X=-0.19 $Y=1.655 $X2=2.51 $Y2=1.98
cc_228 VPB N_A_1641_21#_c_1542_n 0.00444026f $X=-0.19 $Y=1.655 $X2=2.51 $Y2=1.98
cc_229 VPB N_A_1641_21#_c_1543_n 0.0362486f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_230 VPB N_CLK_M1018_g 0.0246943f $X=-0.19 $Y=1.655 $X2=1.465 $Y2=0.78
cc_231 VPB N_CLK_c_1645_n 0.0108727f $X=-0.19 $Y=1.655 $X2=0.23 $Y2=1.03
cc_232 VPB N_CLK_c_1648_n 0.0190443f $X=-0.19 $Y=1.655 $X2=1.345 $Y2=0.945
cc_233 VPB N_A_2408_367#_M1024_g 0.0250849f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_234 VPB N_A_2408_367#_c_1692_n 0.00467014f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_235 VPB N_A_2408_367#_c_1693_n 0.00597292f $X=-0.19 $Y=1.655 $X2=1.345
+ $Y2=0.945
cc_236 VPB N_A_2408_367#_c_1694_n 0.00379656f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_237 VPB N_VPWR_c_1743_n 0.00531831f $X=-0.19 $Y=1.655 $X2=0.26 $Y2=0.945
cc_238 VPB N_VPWR_c_1744_n 0.0100613f $X=-0.19 $Y=1.655 $X2=1.055 $Y2=2.46
cc_239 VPB N_VPWR_c_1745_n 0.0153847f $X=-0.19 $Y=1.655 $X2=2.51 $Y2=1.98
cc_240 VPB N_VPWR_c_1746_n 0.0181487f $X=-0.19 $Y=1.655 $X2=1.465 $Y2=0.945
cc_241 VPB N_VPWR_c_1747_n 0.0152043f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_242 VPB N_VPWR_c_1748_n 0.00936972f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_243 VPB N_VPWR_c_1749_n 0.00274115f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_244 VPB N_VPWR_c_1750_n 0.0248121f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_245 VPB N_VPWR_c_1751_n 0.0359931f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_246 VPB N_VPWR_c_1752_n 0.00607747f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_247 VPB N_VPWR_c_1753_n 0.0413539f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_248 VPB N_VPWR_c_1754_n 0.0427079f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_249 VPB N_VPWR_c_1755_n 0.0308922f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_250 VPB N_VPWR_c_1756_n 0.0200512f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_251 VPB N_VPWR_c_1757_n 0.0411356f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_252 VPB N_VPWR_c_1758_n 0.0152818f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_253 VPB N_VPWR_c_1742_n 0.107535f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_254 VPB N_VPWR_c_1760_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_255 VPB N_VPWR_c_1761_n 0.00435574f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_256 VPB N_VPWR_c_1762_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_257 VPB N_VPWR_c_1763_n 0.0417153f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_258 VPB N_VPWR_c_1764_n 0.0143949f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_259 VPB N_VPWR_c_1765_n 0.00492097f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_260 VPB N_VPWR_c_1766_n 0.00501344f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_261 VPB N_VPWR_c_1767_n 0.0080898f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_262 VPB N_A_380_50#_c_1893_n 0.00486276f $X=-0.19 $Y=1.655 $X2=0.43 $Y2=0.945
cc_263 VPB N_A_380_50#_c_1897_n 0.00385785f $X=-0.19 $Y=1.655 $X2=1.055 $Y2=2.46
cc_264 VPB N_A_380_50#_c_1898_n 0.0103533f $X=-0.19 $Y=1.655 $X2=2.51 $Y2=1.98
cc_265 VPB N_Q_c_1994_n 0.0569993f $X=-0.19 $Y=1.655 $X2=0.43 $Y2=0.945
cc_266 N_A_35_74#_c_269_n N_SCE_M1026_g 0.00335876f $X=0.3 $Y=0.58 $X2=0 $Y2=0
cc_267 N_A_35_74#_c_270_n N_SCE_M1026_g 0.0353252f $X=0.23 $Y=1.975 $X2=0 $Y2=0
cc_268 N_A_35_74#_c_271_n N_SCE_M1026_g 0.0177356f $X=1.345 $Y=0.945 $X2=0 $Y2=0
cc_269 N_A_35_74#_c_272_n N_SCE_M1026_g 0.00679574f $X=1.345 $Y=0.945 $X2=0
+ $Y2=0
cc_270 N_A_35_74#_c_277_n N_SCE_c_342_n 0.0167718f $X=1.15 $Y=2.47 $X2=0 $Y2=0
cc_271 N_A_35_74#_c_276_n N_SCE_c_348_n 0.00269987f $X=2.425 $Y=2.06 $X2=0 $Y2=0
cc_272 N_A_35_74#_c_277_n N_SCE_c_348_n 0.0142219f $X=1.15 $Y=2.47 $X2=0 $Y2=0
cc_273 N_A_35_74#_c_277_n N_SCE_c_349_n 0.0217777f $X=1.15 $Y=2.47 $X2=0 $Y2=0
cc_274 N_A_35_74#_c_277_n N_SCE_M1021_g 0.00651992f $X=1.15 $Y=2.47 $X2=0 $Y2=0
cc_275 N_A_35_74#_c_276_n N_SCE_c_351_n 0.0196347f $X=2.425 $Y=2.06 $X2=0 $Y2=0
cc_276 N_A_35_74#_c_276_n N_SCE_c_353_n 0.00977985f $X=2.425 $Y=2.06 $X2=0 $Y2=0
cc_277 N_A_35_74#_c_270_n SCE 0.0159535f $X=0.23 $Y=1.975 $X2=0 $Y2=0
cc_278 N_A_35_74#_c_271_n SCE 0.0709307f $X=1.345 $Y=0.945 $X2=0 $Y2=0
cc_279 N_A_35_74#_c_272_n SCE 0.00981046f $X=1.345 $Y=0.945 $X2=0 $Y2=0
cc_280 N_A_35_74#_c_277_n SCE 0.00720962f $X=1.15 $Y=2.47 $X2=0 $Y2=0
cc_281 N_A_35_74#_c_278_n SCE 0.00908298f $X=2.51 $Y=1.98 $X2=0 $Y2=0
cc_282 N_A_35_74#_c_279_n SCE 0.00114784f $X=2.51 $Y=1.98 $X2=0 $Y2=0
cc_283 N_A_35_74#_c_271_n N_SCE_c_345_n 0.0092968f $X=1.345 $Y=0.945 $X2=0 $Y2=0
cc_284 N_A_35_74#_c_276_n N_SCE_c_346_n 0.00188542f $X=2.425 $Y=2.06 $X2=0 $Y2=0
cc_285 N_A_35_74#_c_278_n N_SCE_c_346_n 6.59891e-19 $X=2.51 $Y=1.98 $X2=0 $Y2=0
cc_286 N_A_35_74#_c_279_n N_SCE_c_346_n 0.00748415f $X=2.51 $Y=1.98 $X2=0 $Y2=0
cc_287 N_A_35_74#_c_268_n N_D_M1033_g 0.0520003f $X=1.465 $Y=0.78 $X2=0 $Y2=0
cc_288 N_A_35_74#_c_271_n N_D_M1033_g 7.20839e-19 $X=1.345 $Y=0.945 $X2=0 $Y2=0
cc_289 N_A_35_74#_c_272_n N_D_M1033_g 0.010027f $X=1.345 $Y=0.945 $X2=0 $Y2=0
cc_290 N_A_35_74#_M1015_g N_D_M1028_g 0.0149331f $X=2.49 $Y=2.635 $X2=0 $Y2=0
cc_291 N_A_35_74#_c_276_n N_D_M1028_g 0.0141229f $X=2.425 $Y=2.06 $X2=0 $Y2=0
cc_292 N_A_35_74#_c_270_n D 0.0141229f $X=0.23 $Y=1.975 $X2=0 $Y2=0
cc_293 N_A_35_74#_c_277_n D 0.124943f $X=1.15 $Y=2.47 $X2=0 $Y2=0
cc_294 N_A_35_74#_c_276_n N_D_c_414_n 0.00597341f $X=2.425 $Y=2.06 $X2=0 $Y2=0
cc_295 N_A_35_74#_c_278_n N_D_c_414_n 8.93124e-19 $X=2.51 $Y=1.98 $X2=0 $Y2=0
cc_296 N_A_35_74#_c_279_n N_D_c_414_n 0.0213899f $X=2.51 $Y=1.98 $X2=0 $Y2=0
cc_297 N_A_35_74#_M1015_g N_SCD_M1008_g 0.0362823f $X=2.49 $Y=2.635 $X2=0 $Y2=0
cc_298 N_A_35_74#_c_278_n N_SCD_c_452_n 0.00107917f $X=2.51 $Y=1.98 $X2=0 $Y2=0
cc_299 N_A_35_74#_c_279_n N_SCD_c_452_n 0.019352f $X=2.51 $Y=1.98 $X2=0 $Y2=0
cc_300 N_A_35_74#_c_278_n SCD 0.0158523f $X=2.51 $Y=1.98 $X2=0 $Y2=0
cc_301 N_A_35_74#_c_279_n SCD 0.00101891f $X=2.51 $Y=1.98 $X2=0 $Y2=0
cc_302 N_A_35_74#_c_276_n N_VPWR_c_1743_n 0.0204885f $X=2.425 $Y=2.06 $X2=0
+ $Y2=0
cc_303 N_A_35_74#_c_277_n N_VPWR_c_1743_n 0.0248406f $X=1.15 $Y=2.47 $X2=0 $Y2=0
cc_304 N_A_35_74#_c_277_n N_VPWR_c_1751_n 0.0444212f $X=1.15 $Y=2.47 $X2=0 $Y2=0
cc_305 N_A_35_74#_M1015_g N_VPWR_c_1753_n 0.00430111f $X=2.49 $Y=2.635 $X2=0
+ $Y2=0
cc_306 N_A_35_74#_M1015_g N_VPWR_c_1742_n 0.00544287f $X=2.49 $Y=2.635 $X2=0
+ $Y2=0
cc_307 N_A_35_74#_c_277_n N_VPWR_c_1742_n 0.0387633f $X=1.15 $Y=2.47 $X2=0 $Y2=0
cc_308 N_A_35_74#_M1015_g N_A_380_50#_c_1899_n 0.00871523f $X=2.49 $Y=2.635
+ $X2=0 $Y2=0
cc_309 N_A_35_74#_c_278_n N_A_380_50#_c_1899_n 0.0149491f $X=2.51 $Y=1.98 $X2=0
+ $Y2=0
cc_310 N_A_35_74#_c_279_n N_A_380_50#_c_1899_n 6.44022e-19 $X=2.51 $Y=1.98 $X2=0
+ $Y2=0
cc_311 N_A_35_74#_c_271_n N_A_380_50#_c_1895_n 0.00473769f $X=1.345 $Y=0.945
+ $X2=0 $Y2=0
cc_312 N_A_35_74#_M1015_g N_A_380_50#_c_1897_n 0.0109461f $X=2.49 $Y=2.635 $X2=0
+ $Y2=0
cc_313 N_A_35_74#_c_276_n N_A_380_50#_c_1897_n 0.0203555f $X=2.425 $Y=2.06 $X2=0
+ $Y2=0
cc_314 N_A_35_74#_c_278_n N_A_380_50#_c_1897_n 0.00112338f $X=2.51 $Y=1.98 $X2=0
+ $Y2=0
cc_315 N_A_35_74#_c_279_n N_A_380_50#_c_1897_n 0.0014565f $X=2.51 $Y=1.98 $X2=0
+ $Y2=0
cc_316 N_A_35_74#_c_268_n N_VGND_c_2005_n 0.00474635f $X=1.465 $Y=0.78 $X2=0
+ $Y2=0
cc_317 N_A_35_74#_c_271_n N_VGND_c_2005_n 0.0217311f $X=1.345 $Y=0.945 $X2=0
+ $Y2=0
cc_318 N_A_35_74#_c_269_n N_VGND_c_2015_n 0.0109303f $X=0.3 $Y=0.58 $X2=0 $Y2=0
cc_319 N_A_35_74#_c_268_n N_VGND_c_2016_n 0.00349953f $X=1.465 $Y=0.78 $X2=0
+ $Y2=0
cc_320 N_A_35_74#_c_268_n N_VGND_c_2020_n 0.00635843f $X=1.465 $Y=0.78 $X2=0
+ $Y2=0
cc_321 N_A_35_74#_c_269_n N_VGND_c_2020_n 0.0119744f $X=0.3 $Y=0.58 $X2=0 $Y2=0
cc_322 N_A_35_74#_c_271_n N_VGND_c_2020_n 0.0149568f $X=1.345 $Y=0.945 $X2=0
+ $Y2=0
cc_323 N_A_35_74#_c_268_n N_noxref_24_c_2144_n 0.00910876f $X=1.465 $Y=0.78
+ $X2=0 $Y2=0
cc_324 N_A_35_74#_c_271_n N_noxref_24_c_2144_n 0.00370401f $X=1.345 $Y=0.945
+ $X2=0 $Y2=0
cc_325 N_A_35_74#_c_271_n N_noxref_24_c_2148_n 0.00982261f $X=1.345 $Y=0.945
+ $X2=0 $Y2=0
cc_326 N_A_35_74#_c_272_n N_noxref_24_c_2148_n 0.00403509f $X=1.345 $Y=0.945
+ $X2=0 $Y2=0
cc_327 N_SCE_M1038_g N_D_M1033_g 0.0180968f $X=2.485 $Y=0.615 $X2=0 $Y2=0
cc_328 SCE N_D_M1033_g 0.0187428f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_329 N_SCE_c_346_n N_D_M1033_g 0.013401f $X=2.395 $Y=1.295 $X2=0 $Y2=0
cc_330 N_SCE_c_351_n N_D_M1028_g 0.0629716f $X=1.625 $Y=2.105 $X2=0 $Y2=0
cc_331 N_SCE_c_342_n D 0.0229603f $X=0.677 $Y=2.03 $X2=0 $Y2=0
cc_332 N_SCE_c_348_n D 0.00464512f $X=1.195 $Y=2.105 $X2=0 $Y2=0
cc_333 SCE D 0.122399f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_334 N_SCE_c_346_n D 6.10408e-19 $X=2.395 $Y=1.295 $X2=0 $Y2=0
cc_335 N_SCE_c_351_n N_D_c_414_n 0.00733278f $X=1.625 $Y=2.105 $X2=0 $Y2=0
cc_336 SCE N_D_c_414_n 0.00546922f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_337 N_SCE_M1038_g N_SCD_M1000_g 0.0336146f $X=2.485 $Y=0.615 $X2=0 $Y2=0
cc_338 SCE N_SCD_c_448_n 0.00394382f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_339 N_SCE_c_346_n N_SCD_c_448_n 0.0336146f $X=2.395 $Y=1.295 $X2=0 $Y2=0
cc_340 SCE SCD 0.0157283f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_341 N_SCE_c_346_n SCD 6.27939e-19 $X=2.395 $Y=1.295 $X2=0 $Y2=0
cc_342 SCE N_SCD_c_450_n 6.11537e-19 $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_343 N_SCE_c_346_n N_SCD_c_450_n 0.00525736f $X=2.395 $Y=1.295 $X2=0 $Y2=0
cc_344 N_SCE_M1021_g N_VPWR_c_1743_n 0.0145212f $X=1.27 $Y=2.635 $X2=0 $Y2=0
cc_345 N_SCE_c_351_n N_VPWR_c_1743_n 0.00208388f $X=1.625 $Y=2.105 $X2=0 $Y2=0
cc_346 N_SCE_M1001_g N_VPWR_c_1743_n 0.0147584f $X=1.7 $Y=2.635 $X2=0 $Y2=0
cc_347 N_SCE_M1021_g N_VPWR_c_1751_n 0.00379792f $X=1.27 $Y=2.635 $X2=0 $Y2=0
cc_348 N_SCE_M1001_g N_VPWR_c_1753_n 0.00379792f $X=1.7 $Y=2.635 $X2=0 $Y2=0
cc_349 N_SCE_M1021_g N_VPWR_c_1742_n 0.00457201f $X=1.27 $Y=2.635 $X2=0 $Y2=0
cc_350 N_SCE_M1001_g N_VPWR_c_1742_n 0.00457201f $X=1.7 $Y=2.635 $X2=0 $Y2=0
cc_351 N_SCE_M1038_g N_A_380_50#_c_1892_n 0.0110587f $X=2.485 $Y=0.615 $X2=0
+ $Y2=0
cc_352 SCE N_A_380_50#_c_1892_n 0.0289468f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_353 N_SCE_c_346_n N_A_380_50#_c_1892_n 0.00212768f $X=2.395 $Y=1.295 $X2=0
+ $Y2=0
cc_354 N_SCE_M1038_g N_A_380_50#_c_1895_n 0.00588568f $X=2.485 $Y=0.615 $X2=0
+ $Y2=0
cc_355 SCE N_A_380_50#_c_1895_n 0.0222162f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_356 N_SCE_c_346_n N_A_380_50#_c_1895_n 0.00215559f $X=2.395 $Y=1.295 $X2=0
+ $Y2=0
cc_357 N_SCE_M1001_g N_A_380_50#_c_1897_n 0.00184794f $X=1.7 $Y=2.635 $X2=0
+ $Y2=0
cc_358 N_SCE_M1026_g N_VGND_c_2005_n 0.00561055f $X=0.515 $Y=0.58 $X2=0 $Y2=0
cc_359 N_SCE_M1026_g N_VGND_c_2015_n 0.00461464f $X=0.515 $Y=0.58 $X2=0 $Y2=0
cc_360 N_SCE_M1038_g N_VGND_c_2016_n 9.29198e-19 $X=2.485 $Y=0.615 $X2=0 $Y2=0
cc_361 N_SCE_M1026_g N_VGND_c_2020_n 0.00476292f $X=0.515 $Y=0.58 $X2=0 $Y2=0
cc_362 N_SCE_M1038_g N_noxref_24_c_2144_n 0.0117791f $X=2.485 $Y=0.615 $X2=0
+ $Y2=0
cc_363 N_SCE_M1038_g N_noxref_24_c_2145_n 0.00103346f $X=2.485 $Y=0.615 $X2=0
+ $Y2=0
cc_364 D N_SCD_c_450_n 0.00655784f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_365 N_D_M1028_g N_VPWR_c_1743_n 0.00230199f $X=2.06 $Y=2.635 $X2=0 $Y2=0
cc_366 N_D_M1028_g N_VPWR_c_1753_n 0.00430111f $X=2.06 $Y=2.635 $X2=0 $Y2=0
cc_367 N_D_M1028_g N_VPWR_c_1742_n 0.00544287f $X=2.06 $Y=2.635 $X2=0 $Y2=0
cc_368 N_D_M1033_g N_A_380_50#_c_1895_n 0.00874656f $X=1.825 $Y=0.46 $X2=0 $Y2=0
cc_369 N_D_M1028_g N_A_380_50#_c_1897_n 0.0118256f $X=2.06 $Y=2.635 $X2=0 $Y2=0
cc_370 N_D_M1033_g N_VGND_c_2016_n 0.00349953f $X=1.825 $Y=0.46 $X2=0 $Y2=0
cc_371 N_D_M1033_g N_VGND_c_2020_n 0.00635843f $X=1.825 $Y=0.46 $X2=0 $Y2=0
cc_372 N_D_M1033_g N_noxref_24_c_2144_n 0.0148629f $X=1.825 $Y=0.46 $X2=0 $Y2=0
cc_373 N_SCD_M1000_g N_RESET_B_M1027_g 0.0134292f $X=2.845 $Y=0.615 $X2=0 $Y2=0
cc_374 SCD N_RESET_B_M1027_g 4.58115e-19 $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_375 N_SCD_c_448_n N_RESET_B_c_801_n 0.0194382f $X=2.992 $Y=1.325 $X2=0 $Y2=0
cc_376 SCD N_RESET_B_c_801_n 0.00551862f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_377 N_SCD_M1008_g N_RESET_B_c_806_n 0.00526854f $X=2.96 $Y=2.635 $X2=0 $Y2=0
cc_378 N_SCD_c_450_n N_RESET_B_c_806_n 0.0194382f $X=3.05 $Y=1.34 $X2=0 $Y2=0
cc_379 N_SCD_M1008_g N_RESET_B_c_816_n 0.0223279f $X=2.96 $Y=2.635 $X2=0 $Y2=0
cc_380 SCD N_RESET_B_c_816_n 7.61824e-19 $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_381 N_SCD_M1008_g N_VPWR_c_1744_n 0.00329429f $X=2.96 $Y=2.635 $X2=0 $Y2=0
cc_382 N_SCD_M1008_g N_VPWR_c_1753_n 0.00457417f $X=2.96 $Y=2.635 $X2=0 $Y2=0
cc_383 N_SCD_M1008_g N_VPWR_c_1742_n 0.00544287f $X=2.96 $Y=2.635 $X2=0 $Y2=0
cc_384 N_SCD_M1000_g N_A_380_50#_c_1892_n 0.0149041f $X=2.845 $Y=0.615 $X2=0
+ $Y2=0
cc_385 N_SCD_c_448_n N_A_380_50#_c_1892_n 0.00356171f $X=2.992 $Y=1.325 $X2=0
+ $Y2=0
cc_386 SCD N_A_380_50#_c_1892_n 0.0256245f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_387 N_SCD_M1008_g N_A_380_50#_c_1899_n 0.0148253f $X=2.96 $Y=2.635 $X2=0
+ $Y2=0
cc_388 N_SCD_c_452_n N_A_380_50#_c_1899_n 5.78718e-19 $X=3.05 $Y=1.845 $X2=0
+ $Y2=0
cc_389 SCD N_A_380_50#_c_1899_n 0.0259543f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_390 N_SCD_M1000_g N_A_380_50#_c_1893_n 0.00440568f $X=2.845 $Y=0.615 $X2=0
+ $Y2=0
cc_391 N_SCD_M1008_g N_A_380_50#_c_1893_n 9.68145e-19 $X=2.96 $Y=2.635 $X2=0
+ $Y2=0
cc_392 N_SCD_c_448_n N_A_380_50#_c_1893_n 7.28965e-19 $X=2.992 $Y=1.325 $X2=0
+ $Y2=0
cc_393 SCD N_A_380_50#_c_1893_n 0.0744761f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_394 N_SCD_M1008_g N_A_380_50#_c_1897_n 0.00185213f $X=2.96 $Y=2.635 $X2=0
+ $Y2=0
cc_395 N_SCD_M1000_g N_VGND_c_2016_n 9.22791e-19 $X=2.845 $Y=0.615 $X2=0 $Y2=0
cc_396 N_SCD_M1000_g N_noxref_24_c_2144_n 0.00817472f $X=2.845 $Y=0.615 $X2=0
+ $Y2=0
cc_397 N_SCD_M1000_g N_noxref_24_c_2145_n 0.00646685f $X=2.845 $Y=0.615 $X2=0
+ $Y2=0
cc_398 N_A_757_317#_c_506_n N_A_937_333#_c_706_n 0.00258545f $X=4.9 $Y=1.29
+ $X2=0 $Y2=0
cc_399 N_A_757_317#_c_507_n N_A_937_333#_c_706_n 3.98058e-19 $X=4.9 $Y=1.29
+ $X2=0 $Y2=0
cc_400 N_A_757_317#_c_499_n N_A_937_333#_M1011_g 0.00235861f $X=7.295 $Y=1.295
+ $X2=0 $Y2=0
cc_401 N_A_757_317#_c_500_n N_A_937_333#_M1011_g 7.02072e-19 $X=5.185 $Y=1.295
+ $X2=0 $Y2=0
cc_402 N_A_757_317#_c_506_n N_A_937_333#_M1011_g 0.019307f $X=4.9 $Y=1.29 $X2=0
+ $Y2=0
cc_403 N_A_757_317#_c_507_n N_A_937_333#_M1011_g 0.0048667f $X=4.9 $Y=1.29 $X2=0
+ $Y2=0
cc_404 N_A_757_317#_c_508_n N_A_937_333#_M1011_g 0.028208f $X=4.9 $Y=1.125 $X2=0
+ $Y2=0
cc_405 N_A_757_317#_c_506_n N_A_937_333#_c_700_n 0.00181244f $X=4.9 $Y=1.29
+ $X2=0 $Y2=0
cc_406 N_A_757_317#_c_499_n N_A_937_333#_c_701_n 0.00359355f $X=7.295 $Y=1.295
+ $X2=0 $Y2=0
cc_407 N_A_757_317#_c_500_n N_A_937_333#_c_701_n 7.06875e-19 $X=5.185 $Y=1.295
+ $X2=0 $Y2=0
cc_408 N_A_757_317#_c_499_n N_A_937_333#_c_702_n 0.0341345f $X=7.295 $Y=1.295
+ $X2=0 $Y2=0
cc_409 N_A_757_317#_c_500_n N_A_937_333#_c_702_n 0.00274791f $X=5.185 $Y=1.295
+ $X2=0 $Y2=0
cc_410 N_A_757_317#_c_506_n N_A_937_333#_c_702_n 2.98125e-19 $X=4.9 $Y=1.29
+ $X2=0 $Y2=0
cc_411 N_A_757_317#_c_507_n N_A_937_333#_c_702_n 0.00761856f $X=4.9 $Y=1.29
+ $X2=0 $Y2=0
cc_412 N_A_757_317#_c_493_n N_A_937_333#_c_703_n 0.00271203f $X=7.15 $Y=1.095
+ $X2=0 $Y2=0
cc_413 N_A_757_317#_c_499_n N_A_937_333#_c_703_n 0.020689f $X=7.295 $Y=1.295
+ $X2=0 $Y2=0
cc_414 N_A_757_317#_c_499_n N_A_937_333#_c_728_n 0.00519041f $X=7.295 $Y=1.295
+ $X2=0 $Y2=0
cc_415 N_A_757_317#_c_497_n N_A_937_333#_c_704_n 0.00139051f $X=4.895 $Y=1.295
+ $X2=0 $Y2=0
cc_416 N_A_757_317#_c_500_n N_A_937_333#_c_704_n 9.21312e-19 $X=5.185 $Y=1.295
+ $X2=0 $Y2=0
cc_417 N_A_757_317#_c_506_n N_A_937_333#_c_704_n 0.00177905f $X=4.9 $Y=1.29
+ $X2=0 $Y2=0
cc_418 N_A_757_317#_c_507_n N_A_937_333#_c_704_n 0.0201225f $X=4.9 $Y=1.29 $X2=0
+ $Y2=0
cc_419 N_A_757_317#_c_493_n N_A_937_333#_c_733_n 0.00292155f $X=7.15 $Y=1.095
+ $X2=0 $Y2=0
cc_420 N_A_757_317#_c_497_n N_A_937_333#_c_711_n 0.00105794f $X=4.895 $Y=1.295
+ $X2=0 $Y2=0
cc_421 N_A_757_317#_c_506_n N_A_937_333#_c_711_n 0.0180362f $X=4.9 $Y=1.29 $X2=0
+ $Y2=0
cc_422 N_A_757_317#_c_507_n N_A_937_333#_c_711_n 2.92334e-19 $X=4.9 $Y=1.29
+ $X2=0 $Y2=0
cc_423 N_A_757_317#_c_502_n N_RESET_B_c_800_n 0.00563574f $X=4.08 $Y=1.295 $X2=0
+ $Y2=0
cc_424 N_A_757_317#_c_505_n N_RESET_B_c_800_n 0.00827426f $X=3.95 $Y=1.75 $X2=0
+ $Y2=0
cc_425 N_A_757_317#_c_502_n N_RESET_B_c_802_n 0.00224282f $X=4.08 $Y=1.295 $X2=0
+ $Y2=0
cc_426 N_A_757_317#_c_508_n N_RESET_B_c_803_n 0.0099884f $X=4.9 $Y=1.125 $X2=0
+ $Y2=0
cc_427 N_A_757_317#_c_501_n N_RESET_B_M1005_g 0.00216111f $X=10.175 $Y=1.295
+ $X2=0 $Y2=0
cc_428 N_A_757_317#_M1019_g N_RESET_B_c_806_n 0.00987775f $X=3.97 $Y=2.525 $X2=0
+ $Y2=0
cc_429 N_A_757_317#_c_502_n N_RESET_B_c_806_n 0.00167349f $X=4.08 $Y=1.295 $X2=0
+ $Y2=0
cc_430 N_A_757_317#_c_505_n N_RESET_B_c_806_n 0.0203599f $X=3.95 $Y=1.75 $X2=0
+ $Y2=0
cc_431 N_A_757_317#_M1019_g N_RESET_B_c_816_n 0.0092933f $X=3.97 $Y=2.525 $X2=0
+ $Y2=0
cc_432 N_A_757_317#_c_499_n N_RESET_B_c_808_n 0.00223746f $X=7.295 $Y=1.295
+ $X2=0 $Y2=0
cc_433 N_A_757_317#_c_507_n N_RESET_B_c_808_n 3.89064e-19 $X=4.9 $Y=1.29 $X2=0
+ $Y2=0
cc_434 N_A_757_317#_M1022_g N_RESET_B_c_819_n 0.0135884f $X=7.815 $Y=2.875 $X2=0
+ $Y2=0
cc_435 N_A_757_317#_c_512_n N_RESET_B_c_819_n 0.00600854f $X=7.955 $Y=2.22 $X2=0
+ $Y2=0
cc_436 N_A_757_317#_c_513_n N_RESET_B_c_819_n 0.00234434f $X=7.955 $Y=2.22 $X2=0
+ $Y2=0
cc_437 N_A_757_317#_M1022_g N_RESET_B_c_821_n 0.00517733f $X=7.815 $Y=2.875
+ $X2=0 $Y2=0
cc_438 N_A_757_317#_M1022_g N_RESET_B_c_823_n 0.00219577f $X=7.815 $Y=2.875
+ $X2=0 $Y2=0
cc_439 N_A_757_317#_c_512_n N_RESET_B_c_823_n 0.00696017f $X=7.955 $Y=2.22 $X2=0
+ $Y2=0
cc_440 N_A_757_317#_c_513_n N_RESET_B_c_823_n 0.00217003f $X=7.955 $Y=2.22 $X2=0
+ $Y2=0
cc_441 N_A_757_317#_c_499_n N_RESET_B_c_809_n 0.00371297f $X=7.295 $Y=1.295
+ $X2=0 $Y2=0
cc_442 N_A_757_317#_c_493_n N_A_809_463#_M1030_g 0.00703541f $X=7.15 $Y=1.095
+ $X2=0 $Y2=0
cc_443 N_A_757_317#_M1019_g N_A_809_463#_c_1010_n 9.43263e-19 $X=3.97 $Y=2.525
+ $X2=0 $Y2=0
cc_444 N_A_757_317#_c_497_n N_A_809_463#_c_1010_n 0.0225166f $X=4.895 $Y=1.295
+ $X2=0 $Y2=0
cc_445 N_A_757_317#_c_498_n N_A_809_463#_c_1010_n 0.00256146f $X=4.225 $Y=1.295
+ $X2=0 $Y2=0
cc_446 N_A_757_317#_c_500_n N_A_809_463#_c_1010_n 4.63228e-19 $X=5.185 $Y=1.295
+ $X2=0 $Y2=0
cc_447 N_A_757_317#_c_502_n N_A_809_463#_c_1010_n 0.055587f $X=4.08 $Y=1.295
+ $X2=0 $Y2=0
cc_448 N_A_757_317#_c_505_n N_A_809_463#_c_1010_n 3.10013e-19 $X=3.95 $Y=1.75
+ $X2=0 $Y2=0
cc_449 N_A_757_317#_c_506_n N_A_809_463#_c_1010_n 0.00208004f $X=4.9 $Y=1.29
+ $X2=0 $Y2=0
cc_450 N_A_757_317#_c_507_n N_A_809_463#_c_1010_n 0.0173174f $X=4.9 $Y=1.29
+ $X2=0 $Y2=0
cc_451 N_A_757_317#_c_508_n N_A_809_463#_c_1010_n 0.00204678f $X=4.9 $Y=1.125
+ $X2=0 $Y2=0
cc_452 N_A_757_317#_c_497_n N_A_809_463#_c_1011_n 0.00874156f $X=4.895 $Y=1.295
+ $X2=0 $Y2=0
cc_453 N_A_757_317#_c_499_n N_A_809_463#_c_1011_n 0.0264322f $X=7.295 $Y=1.295
+ $X2=0 $Y2=0
cc_454 N_A_757_317#_c_500_n N_A_809_463#_c_1011_n 0.00367252f $X=5.185 $Y=1.295
+ $X2=0 $Y2=0
cc_455 N_A_757_317#_c_506_n N_A_809_463#_c_1011_n 0.00396693f $X=4.9 $Y=1.29
+ $X2=0 $Y2=0
cc_456 N_A_757_317#_c_507_n N_A_809_463#_c_1011_n 0.0225689f $X=4.9 $Y=1.29
+ $X2=0 $Y2=0
cc_457 N_A_757_317#_c_508_n N_A_809_463#_c_1011_n 0.00895602f $X=4.9 $Y=1.125
+ $X2=0 $Y2=0
cc_458 N_A_757_317#_c_499_n N_A_809_463#_c_1012_n 0.0205864f $X=7.295 $Y=1.295
+ $X2=0 $Y2=0
cc_459 N_A_757_317#_M1019_g N_A_809_463#_c_1017_n 0.0109189f $X=3.97 $Y=2.525
+ $X2=0 $Y2=0
cc_460 N_A_757_317#_c_502_n N_A_809_463#_c_1017_n 0.0174766f $X=4.08 $Y=1.295
+ $X2=0 $Y2=0
cc_461 N_A_757_317#_c_505_n N_A_809_463#_c_1017_n 5.45775e-19 $X=3.95 $Y=1.75
+ $X2=0 $Y2=0
cc_462 N_A_757_317#_c_493_n N_A_809_463#_c_1013_n 0.00959833f $X=7.15 $Y=1.095
+ $X2=0 $Y2=0
cc_463 N_A_757_317#_c_499_n N_A_809_463#_c_1013_n 0.0097991f $X=7.295 $Y=1.295
+ $X2=0 $Y2=0
cc_464 N_A_757_317#_M1019_g N_A_865_255#_M1037_g 0.0248559f $X=3.97 $Y=2.525
+ $X2=0 $Y2=0
cc_465 N_A_757_317#_c_505_n N_A_865_255#_M1037_g 0.0193707f $X=3.95 $Y=1.75
+ $X2=0 $Y2=0
cc_466 N_A_757_317#_c_506_n N_A_865_255#_M1037_g 0.00140529f $X=4.9 $Y=1.29
+ $X2=0 $Y2=0
cc_467 N_A_757_317#_c_497_n N_A_865_255#_M1032_g 7.81925e-19 $X=4.895 $Y=1.295
+ $X2=0 $Y2=0
cc_468 N_A_757_317#_c_498_n N_A_865_255#_M1032_g 7.4672e-19 $X=4.225 $Y=1.295
+ $X2=0 $Y2=0
cc_469 N_A_757_317#_c_502_n N_A_865_255#_M1032_g 8.17515e-19 $X=4.08 $Y=1.295
+ $X2=0 $Y2=0
cc_470 N_A_757_317#_c_506_n N_A_865_255#_M1032_g 0.019276f $X=4.9 $Y=1.29 $X2=0
+ $Y2=0
cc_471 N_A_757_317#_c_507_n N_A_865_255#_M1032_g 3.96187e-19 $X=4.9 $Y=1.29
+ $X2=0 $Y2=0
cc_472 N_A_757_317#_c_508_n N_A_865_255#_M1032_g 0.0160598f $X=4.9 $Y=1.125
+ $X2=0 $Y2=0
cc_473 N_A_757_317#_M1022_g N_A_865_255#_c_1139_n 0.0100862f $X=7.815 $Y=2.875
+ $X2=0 $Y2=0
cc_474 N_A_757_317#_c_494_n N_A_865_255#_M1017_g 3.74979e-19 $X=7.855 $Y=2.055
+ $X2=0 $Y2=0
cc_475 N_A_757_317#_c_513_n N_A_865_255#_M1017_g 0.0100862f $X=7.955 $Y=2.22
+ $X2=0 $Y2=0
cc_476 N_A_757_317#_c_493_n N_A_865_255#_c_1125_n 0.0206748f $X=7.15 $Y=1.095
+ $X2=0 $Y2=0
cc_477 N_A_757_317#_c_494_n N_A_865_255#_c_1125_n 0.00427538f $X=7.855 $Y=2.055
+ $X2=0 $Y2=0
cc_478 N_A_757_317#_c_495_n N_A_865_255#_c_1125_n 0.00632784f $X=7.77 $Y=1.26
+ $X2=0 $Y2=0
cc_479 N_A_757_317#_c_513_n N_A_865_255#_c_1125_n 0.00379337f $X=7.955 $Y=2.22
+ $X2=0 $Y2=0
cc_480 N_A_757_317#_c_493_n N_A_865_255#_c_1126_n 0.00482177f $X=7.15 $Y=1.095
+ $X2=0 $Y2=0
cc_481 N_A_757_317#_c_493_n N_A_865_255#_M1012_g 0.0214394f $X=7.15 $Y=1.095
+ $X2=0 $Y2=0
cc_482 N_A_757_317#_c_494_n N_A_865_255#_M1012_g 0.0024479f $X=7.855 $Y=2.055
+ $X2=0 $Y2=0
cc_483 N_A_757_317#_c_495_n N_A_865_255#_M1012_g 0.0109534f $X=7.77 $Y=1.26
+ $X2=0 $Y2=0
cc_484 N_A_757_317#_c_501_n N_A_865_255#_M1012_g 0.00449207f $X=10.175 $Y=1.295
+ $X2=0 $Y2=0
cc_485 N_A_757_317#_c_496_n N_A_865_255#_M1010_g 0.0048505f $X=10.41 $Y=1.08
+ $X2=0 $Y2=0
cc_486 N_A_757_317#_c_504_n N_A_865_255#_M1010_g 0.0139758f $X=10.32 $Y=1.295
+ $X2=0 $Y2=0
cc_487 N_A_757_317#_c_504_n N_A_865_255#_M1035_g 0.00370192f $X=10.32 $Y=1.295
+ $X2=0 $Y2=0
cc_488 N_A_757_317#_c_497_n N_A_865_255#_c_1129_n 0.00361569f $X=4.895 $Y=1.295
+ $X2=0 $Y2=0
cc_489 N_A_757_317#_c_498_n N_A_865_255#_c_1129_n 0.00116424f $X=4.225 $Y=1.295
+ $X2=0 $Y2=0
cc_490 N_A_757_317#_c_502_n N_A_865_255#_c_1129_n 0.00738931f $X=4.08 $Y=1.295
+ $X2=0 $Y2=0
cc_491 N_A_757_317#_c_494_n N_A_865_255#_c_1130_n 0.012357f $X=7.855 $Y=2.055
+ $X2=0 $Y2=0
cc_492 N_A_757_317#_c_512_n N_A_865_255#_c_1130_n 0.00134387f $X=7.955 $Y=2.22
+ $X2=0 $Y2=0
cc_493 N_A_757_317#_c_513_n N_A_865_255#_c_1130_n 0.0175786f $X=7.955 $Y=2.22
+ $X2=0 $Y2=0
cc_494 N_A_757_317#_c_501_n N_A_865_255#_c_1131_n 0.031721f $X=10.175 $Y=1.295
+ $X2=0 $Y2=0
cc_495 N_A_757_317#_c_504_n N_A_865_255#_c_1131_n 0.0150382f $X=10.32 $Y=1.295
+ $X2=0 $Y2=0
cc_496 N_A_757_317#_c_504_n N_A_865_255#_c_1147_n 0.0386407f $X=10.32 $Y=1.295
+ $X2=0 $Y2=0
cc_497 N_A_757_317#_M1035_s N_A_865_255#_c_1148_n 0.0070032f $X=10.325 $Y=1.835
+ $X2=0 $Y2=0
cc_498 N_A_757_317#_c_504_n N_A_865_255#_c_1148_n 0.0261288f $X=10.32 $Y=1.295
+ $X2=0 $Y2=0
cc_499 N_A_757_317#_c_501_n N_A_865_255#_c_1132_n 0.00740588f $X=10.175 $Y=1.295
+ $X2=0 $Y2=0
cc_500 N_A_757_317#_c_494_n N_A_865_255#_c_1133_n 0.0240796f $X=7.855 $Y=2.055
+ $X2=0 $Y2=0
cc_501 N_A_757_317#_c_512_n N_A_865_255#_c_1133_n 5.57841e-19 $X=7.955 $Y=2.22
+ $X2=0 $Y2=0
cc_502 N_A_757_317#_c_501_n N_A_865_255#_c_1133_n 0.00696043f $X=10.175 $Y=1.295
+ $X2=0 $Y2=0
cc_503 N_A_757_317#_c_503_n N_A_865_255#_c_1134_n 4.12674e-19 $X=10.32 $Y=1.295
+ $X2=0 $Y2=0
cc_504 N_A_757_317#_c_504_n N_A_865_255#_c_1134_n 0.0554998f $X=10.32 $Y=1.295
+ $X2=0 $Y2=0
cc_505 N_A_757_317#_c_504_n N_A_865_255#_c_1136_n 0.00397447f $X=10.32 $Y=1.295
+ $X2=0 $Y2=0
cc_506 N_A_757_317#_c_496_n N_A_865_255#_c_1137_n 0.00468987f $X=10.41 $Y=1.08
+ $X2=0 $Y2=0
cc_507 N_A_757_317#_c_504_n N_A_1445_69#_M1014_g 0.00407257f $X=10.32 $Y=1.295
+ $X2=0 $Y2=0
cc_508 N_A_757_317#_c_493_n N_A_1445_69#_c_1330_n 0.0149622f $X=7.15 $Y=1.095
+ $X2=0 $Y2=0
cc_509 N_A_757_317#_c_494_n N_A_1445_69#_c_1330_n 0.00613023f $X=7.855 $Y=2.055
+ $X2=0 $Y2=0
cc_510 N_A_757_317#_c_495_n N_A_1445_69#_c_1330_n 0.0225079f $X=7.77 $Y=1.26
+ $X2=0 $Y2=0
cc_511 N_A_757_317#_c_499_n N_A_1445_69#_c_1330_n 0.00989909f $X=7.295 $Y=1.295
+ $X2=0 $Y2=0
cc_512 N_A_757_317#_c_631_p N_A_1445_69#_c_1330_n 0.00234811f $X=7.585 $Y=1.295
+ $X2=0 $Y2=0
cc_513 N_A_757_317#_c_493_n N_A_1445_69#_c_1331_n 8.0378e-19 $X=7.15 $Y=1.095
+ $X2=0 $Y2=0
cc_514 N_A_757_317#_c_493_n N_A_1445_69#_c_1332_n 0.00441379f $X=7.15 $Y=1.095
+ $X2=0 $Y2=0
cc_515 N_A_757_317#_c_494_n N_A_1445_69#_c_1332_n 0.0114408f $X=7.855 $Y=2.055
+ $X2=0 $Y2=0
cc_516 N_A_757_317#_c_495_n N_A_1445_69#_c_1332_n 0.0138867f $X=7.77 $Y=1.26
+ $X2=0 $Y2=0
cc_517 N_A_757_317#_c_499_n N_A_1445_69#_c_1332_n 0.0055921f $X=7.295 $Y=1.295
+ $X2=0 $Y2=0
cc_518 N_A_757_317#_c_631_p N_A_1445_69#_c_1332_n 0.00375708f $X=7.585 $Y=1.295
+ $X2=0 $Y2=0
cc_519 N_A_757_317#_c_494_n N_A_1445_69#_c_1347_n 0.0184824f $X=7.855 $Y=2.055
+ $X2=0 $Y2=0
cc_520 N_A_757_317#_c_512_n N_A_1445_69#_c_1347_n 0.0171568f $X=7.955 $Y=2.22
+ $X2=0 $Y2=0
cc_521 N_A_757_317#_c_513_n N_A_1445_69#_c_1347_n 0.00950837f $X=7.955 $Y=2.22
+ $X2=0 $Y2=0
cc_522 N_A_757_317#_c_495_n N_A_1445_69#_c_1363_n 0.0103241f $X=7.77 $Y=1.26
+ $X2=0 $Y2=0
cc_523 N_A_757_317#_c_501_n N_A_1445_69#_c_1363_n 0.00825826f $X=10.175 $Y=1.295
+ $X2=0 $Y2=0
cc_524 N_A_757_317#_c_493_n N_A_1445_69#_c_1365_n 0.0175576f $X=7.15 $Y=1.095
+ $X2=0 $Y2=0
cc_525 N_A_757_317#_c_495_n N_A_1445_69#_c_1365_n 0.0282502f $X=7.77 $Y=1.26
+ $X2=0 $Y2=0
cc_526 N_A_757_317#_c_499_n N_A_1445_69#_c_1365_n 0.00466612f $X=7.295 $Y=1.295
+ $X2=0 $Y2=0
cc_527 N_A_757_317#_c_631_p N_A_1445_69#_c_1365_n 0.00344018f $X=7.585 $Y=1.295
+ $X2=0 $Y2=0
cc_528 N_A_757_317#_c_495_n N_A_1445_69#_c_1333_n 0.00317367f $X=7.77 $Y=1.26
+ $X2=0 $Y2=0
cc_529 N_A_757_317#_c_495_n N_A_1445_69#_c_1334_n 0.013455f $X=7.77 $Y=1.26
+ $X2=0 $Y2=0
cc_530 N_A_757_317#_c_501_n N_A_1445_69#_c_1334_n 0.013738f $X=10.175 $Y=1.295
+ $X2=0 $Y2=0
cc_531 N_A_757_317#_c_496_n N_A_1445_69#_c_1335_n 0.0119754f $X=10.41 $Y=1.08
+ $X2=0 $Y2=0
cc_532 N_A_757_317#_c_501_n N_A_1445_69#_c_1335_n 0.0012493f $X=10.175 $Y=1.295
+ $X2=0 $Y2=0
cc_533 N_A_757_317#_M1010_s N_A_1445_69#_c_1336_n 0.00729219f $X=10.265 $Y=0.365
+ $X2=0 $Y2=0
cc_534 N_A_757_317#_c_496_n N_A_1445_69#_c_1336_n 0.023281f $X=10.41 $Y=1.08
+ $X2=0 $Y2=0
cc_535 N_A_757_317#_c_501_n N_A_1445_69#_c_1336_n 0.00464062f $X=10.175 $Y=1.295
+ $X2=0 $Y2=0
cc_536 N_A_757_317#_c_503_n N_A_1445_69#_c_1336_n 0.00281974f $X=10.32 $Y=1.295
+ $X2=0 $Y2=0
cc_537 N_A_757_317#_c_496_n N_A_1445_69#_c_1339_n 9.97596e-19 $X=10.41 $Y=1.08
+ $X2=0 $Y2=0
cc_538 N_A_757_317#_c_501_n N_A_1445_69#_c_1339_n 4.95075e-19 $X=10.175 $Y=1.295
+ $X2=0 $Y2=0
cc_539 N_A_757_317#_c_503_n N_A_1445_69#_c_1339_n 6.2081e-19 $X=10.32 $Y=1.295
+ $X2=0 $Y2=0
cc_540 N_A_757_317#_c_504_n N_A_1445_69#_c_1339_n 0.00208332f $X=10.32 $Y=1.295
+ $X2=0 $Y2=0
cc_541 N_A_757_317#_c_501_n N_A_1445_69#_c_1340_n 0.0551477f $X=10.175 $Y=1.295
+ $X2=0 $Y2=0
cc_542 N_A_757_317#_c_496_n N_A_1445_69#_c_1341_n 0.0187977f $X=10.41 $Y=1.08
+ $X2=0 $Y2=0
cc_543 N_A_757_317#_c_501_n N_A_1445_69#_c_1341_n 0.0300027f $X=10.175 $Y=1.295
+ $X2=0 $Y2=0
cc_544 N_A_757_317#_c_503_n N_A_1445_69#_c_1341_n 0.00197618f $X=10.32 $Y=1.295
+ $X2=0 $Y2=0
cc_545 N_A_757_317#_M1022_g N_A_1641_21#_M1031_g 0.0189174f $X=7.815 $Y=2.875
+ $X2=0 $Y2=0
cc_546 N_A_757_317#_c_494_n N_A_1641_21#_c_1533_n 0.0025582f $X=7.855 $Y=2.055
+ $X2=0 $Y2=0
cc_547 N_A_757_317#_c_495_n N_A_1641_21#_c_1533_n 4.5529e-19 $X=7.77 $Y=1.26
+ $X2=0 $Y2=0
cc_548 N_A_757_317#_c_501_n N_A_1641_21#_c_1533_n 0.00199366f $X=10.175 $Y=1.295
+ $X2=0 $Y2=0
cc_549 N_A_757_317#_c_501_n N_A_1641_21#_c_1534_n 0.00191482f $X=10.175 $Y=1.295
+ $X2=0 $Y2=0
cc_550 N_A_757_317#_c_494_n N_A_1641_21#_c_1541_n 0.00513121f $X=7.855 $Y=2.055
+ $X2=0 $Y2=0
cc_551 N_A_757_317#_c_512_n N_A_1641_21#_c_1541_n 0.0126864f $X=7.955 $Y=2.22
+ $X2=0 $Y2=0
cc_552 N_A_757_317#_c_513_n N_A_1641_21#_c_1541_n 2.81621e-19 $X=7.955 $Y=2.22
+ $X2=0 $Y2=0
cc_553 N_A_757_317#_c_512_n N_A_1641_21#_c_1543_n 9.42755e-19 $X=7.955 $Y=2.22
+ $X2=0 $Y2=0
cc_554 N_A_757_317#_c_513_n N_A_1641_21#_c_1543_n 0.0220833f $X=7.955 $Y=2.22
+ $X2=0 $Y2=0
cc_555 N_A_757_317#_c_496_n N_CLK_M1007_g 5.53004e-19 $X=10.41 $Y=1.08 $X2=0
+ $Y2=0
cc_556 N_A_757_317#_M1019_g N_VPWR_c_1754_n 0.00415095f $X=3.97 $Y=2.525 $X2=0
+ $Y2=0
cc_557 N_A_757_317#_M1035_s N_VPWR_c_1742_n 0.00371882f $X=10.325 $Y=1.835 $X2=0
+ $Y2=0
cc_558 N_A_757_317#_M1019_g N_VPWR_c_1742_n 0.00477801f $X=3.97 $Y=2.525 $X2=0
+ $Y2=0
cc_559 N_A_757_317#_M1022_g N_VPWR_c_1742_n 0.00609018f $X=7.815 $Y=2.875 $X2=0
+ $Y2=0
cc_560 N_A_757_317#_M1022_g N_VPWR_c_1763_n 0.00351226f $X=7.815 $Y=2.875 $X2=0
+ $Y2=0
cc_561 N_A_757_317#_M1022_g N_VPWR_c_1764_n 0.00102088f $X=7.815 $Y=2.875 $X2=0
+ $Y2=0
cc_562 N_A_757_317#_M1019_g N_A_380_50#_c_1893_n 0.00512793f $X=3.97 $Y=2.525
+ $X2=0 $Y2=0
cc_563 N_A_757_317#_c_498_n N_A_380_50#_c_1893_n 0.00133446f $X=4.225 $Y=1.295
+ $X2=0 $Y2=0
cc_564 N_A_757_317#_c_502_n N_A_380_50#_c_1893_n 0.0573999f $X=4.08 $Y=1.295
+ $X2=0 $Y2=0
cc_565 N_A_757_317#_c_505_n N_A_380_50#_c_1893_n 0.00204143f $X=3.95 $Y=1.75
+ $X2=0 $Y2=0
cc_566 N_A_757_317#_c_498_n N_A_380_50#_c_1894_n 5.68965e-19 $X=4.225 $Y=1.295
+ $X2=0 $Y2=0
cc_567 N_A_757_317#_c_502_n N_A_380_50#_c_1894_n 0.0123499f $X=4.08 $Y=1.295
+ $X2=0 $Y2=0
cc_568 N_A_757_317#_c_505_n N_A_380_50#_c_1894_n 5.55021e-19 $X=3.95 $Y=1.75
+ $X2=0 $Y2=0
cc_569 N_A_757_317#_M1019_g N_A_380_50#_c_1898_n 0.00650632f $X=3.97 $Y=2.525
+ $X2=0 $Y2=0
cc_570 N_A_757_317#_c_505_n N_A_380_50#_c_1898_n 0.00141034f $X=3.95 $Y=1.75
+ $X2=0 $Y2=0
cc_571 N_A_757_317#_c_498_n N_A_380_50#_c_1936_n 0.00148592f $X=4.225 $Y=1.295
+ $X2=0 $Y2=0
cc_572 N_A_757_317#_c_502_n N_A_380_50#_c_1936_n 0.0158792f $X=4.08 $Y=1.295
+ $X2=0 $Y2=0
cc_573 N_A_757_317#_c_505_n N_A_380_50#_c_1936_n 3.05411e-19 $X=3.95 $Y=1.75
+ $X2=0 $Y2=0
cc_574 N_A_757_317#_c_493_n N_VGND_c_2007_n 6.4099e-19 $X=7.15 $Y=1.095 $X2=0
+ $Y2=0
cc_575 N_A_757_317#_c_499_n N_VGND_c_2007_n 0.00121302f $X=7.295 $Y=1.295 $X2=0
+ $Y2=0
cc_576 N_A_757_317#_c_501_n N_VGND_c_2008_n 0.00227525f $X=10.175 $Y=1.295 $X2=0
+ $Y2=0
cc_577 N_A_757_317#_c_493_n N_VGND_c_2013_n 0.00346493f $X=7.15 $Y=1.095 $X2=0
+ $Y2=0
cc_578 N_A_757_317#_c_493_n N_VGND_c_2020_n 0.00512292f $X=7.15 $Y=1.095 $X2=0
+ $Y2=0
cc_579 N_A_757_317#_c_508_n N_VGND_c_2020_n 9.39239e-19 $X=4.9 $Y=1.125 $X2=0
+ $Y2=0
cc_580 N_A_937_333#_M1011_g N_RESET_B_c_803_n 0.0099884f $X=5.35 $Y=0.805 $X2=0
+ $Y2=0
cc_581 N_A_937_333#_c_702_n N_RESET_B_c_811_n 0.00767548f $X=6.645 $Y=1.685
+ $X2=0 $Y2=0
cc_582 N_A_937_333#_M1002_g N_RESET_B_c_812_n 0.0144004f $X=4.76 $Y=2.525 $X2=0
+ $Y2=0
cc_583 N_A_937_333#_c_706_n N_RESET_B_c_812_n 0.0156065f $X=5.305 $Y=1.77 $X2=0
+ $Y2=0
cc_584 N_A_937_333#_c_702_n N_RESET_B_c_812_n 8.75404e-19 $X=6.645 $Y=1.685
+ $X2=0 $Y2=0
cc_585 N_A_937_333#_M1011_g N_RESET_B_M1036_g 0.0237671f $X=5.35 $Y=0.805 $X2=0
+ $Y2=0
cc_586 N_A_937_333#_M1011_g N_RESET_B_c_808_n 0.00759536f $X=5.35 $Y=0.805 $X2=0
+ $Y2=0
cc_587 N_A_937_333#_c_702_n N_RESET_B_c_808_n 2.63199e-19 $X=6.645 $Y=1.685
+ $X2=0 $Y2=0
cc_588 N_A_937_333#_M1029_d N_RESET_B_c_817_n 0.00262667f $X=6.84 $Y=1.895 $X2=0
+ $Y2=0
cc_589 N_A_937_333#_c_702_n N_RESET_B_c_817_n 0.0164271f $X=6.645 $Y=1.685 $X2=0
+ $Y2=0
cc_590 N_A_937_333#_c_747_p N_RESET_B_c_817_n 0.0114776f $X=6.835 $Y=2.055 $X2=0
+ $Y2=0
cc_591 N_A_937_333#_c_728_n N_RESET_B_c_817_n 0.00465906f $X=6.98 $Y=2.055 $X2=0
+ $Y2=0
cc_592 N_A_937_333#_M1029_d N_RESET_B_c_818_n 0.00280564f $X=6.84 $Y=1.895 $X2=0
+ $Y2=0
cc_593 N_A_937_333#_c_702_n RESET_B 0.02486f $X=6.645 $Y=1.685 $X2=0 $Y2=0
cc_594 N_A_937_333#_c_702_n N_RESET_B_c_826_n 0.00586558f $X=6.645 $Y=1.685
+ $X2=0 $Y2=0
cc_595 N_A_937_333#_c_709_n N_RESET_B_c_826_n 5.70856e-19 $X=6.745 $Y=1.96 $X2=0
+ $Y2=0
cc_596 N_A_937_333#_c_701_n N_RESET_B_c_809_n 0.0261016f $X=5.365 $Y=1.425 $X2=0
+ $Y2=0
cc_597 N_A_937_333#_c_702_n N_RESET_B_c_809_n 0.0151386f $X=6.645 $Y=1.685 $X2=0
+ $Y2=0
cc_598 N_A_937_333#_c_703_n N_A_809_463#_M1030_g 0.00802211f $X=6.74 $Y=0.86
+ $X2=0 $Y2=0
cc_599 N_A_937_333#_c_709_n N_A_809_463#_M1029_g 0.00676302f $X=6.745 $Y=1.96
+ $X2=0 $Y2=0
cc_600 N_A_937_333#_c_747_p N_A_809_463#_M1029_g 0.0064097f $X=6.835 $Y=2.055
+ $X2=0 $Y2=0
cc_601 N_A_937_333#_c_758_p N_A_809_463#_M1029_g 0.00564862f $X=6.74 $Y=1.685
+ $X2=0 $Y2=0
cc_602 N_A_937_333#_c_704_n N_A_809_463#_c_1010_n 0.0296582f $X=4.87 $Y=1.685
+ $X2=0 $Y2=0
cc_603 N_A_937_333#_c_711_n N_A_809_463#_c_1010_n 0.00384259f $X=5.015 $Y=1.83
+ $X2=0 $Y2=0
cc_604 N_A_937_333#_M1011_g N_A_809_463#_c_1011_n 0.013664f $X=5.35 $Y=0.805
+ $X2=0 $Y2=0
cc_605 N_A_937_333#_c_702_n N_A_809_463#_c_1011_n 0.0110571f $X=6.645 $Y=1.685
+ $X2=0 $Y2=0
cc_606 N_A_937_333#_c_703_n N_A_809_463#_c_1011_n 0.0091919f $X=6.74 $Y=0.86
+ $X2=0 $Y2=0
cc_607 N_A_937_333#_c_711_n N_A_809_463#_c_1011_n 0.00107984f $X=5.015 $Y=1.83
+ $X2=0 $Y2=0
cc_608 N_A_937_333#_M1002_g N_A_809_463#_c_1016_n 0.0159032f $X=4.76 $Y=2.525
+ $X2=0 $Y2=0
cc_609 N_A_937_333#_c_706_n N_A_809_463#_c_1016_n 0.00448954f $X=5.305 $Y=1.77
+ $X2=0 $Y2=0
cc_610 N_A_937_333#_c_702_n N_A_809_463#_c_1016_n 0.0234167f $X=6.645 $Y=1.685
+ $X2=0 $Y2=0
cc_611 N_A_937_333#_c_704_n N_A_809_463#_c_1016_n 0.0216455f $X=4.87 $Y=1.685
+ $X2=0 $Y2=0
cc_612 N_A_937_333#_c_711_n N_A_809_463#_c_1016_n 0.00126186f $X=5.015 $Y=1.83
+ $X2=0 $Y2=0
cc_613 N_A_937_333#_M1002_g N_A_809_463#_c_1055_n 5.94484e-19 $X=4.76 $Y=2.525
+ $X2=0 $Y2=0
cc_614 N_A_937_333#_c_702_n N_A_809_463#_c_1012_n 0.0230666f $X=6.645 $Y=1.685
+ $X2=0 $Y2=0
cc_615 N_A_937_333#_c_703_n N_A_809_463#_c_1012_n 0.0318053f $X=6.74 $Y=0.86
+ $X2=0 $Y2=0
cc_616 N_A_937_333#_M1002_g N_A_809_463#_c_1017_n 0.0035809f $X=4.76 $Y=2.525
+ $X2=0 $Y2=0
cc_617 N_A_937_333#_c_702_n N_A_809_463#_c_1013_n 0.0175228f $X=6.645 $Y=1.685
+ $X2=0 $Y2=0
cc_618 N_A_937_333#_c_703_n N_A_809_463#_c_1013_n 0.0120823f $X=6.74 $Y=0.86
+ $X2=0 $Y2=0
cc_619 N_A_937_333#_c_758_p N_A_809_463#_c_1013_n 0.00175482f $X=6.74 $Y=1.685
+ $X2=0 $Y2=0
cc_620 N_A_937_333#_c_704_n N_A_865_255#_M1037_g 7.25643e-19 $X=4.87 $Y=1.685
+ $X2=0 $Y2=0
cc_621 N_A_937_333#_c_711_n N_A_865_255#_M1037_g 0.0735464f $X=5.015 $Y=1.83
+ $X2=0 $Y2=0
cc_622 N_A_937_333#_M1002_g N_A_865_255#_c_1139_n 0.0104164f $X=4.76 $Y=2.525
+ $X2=0 $Y2=0
cc_623 N_A_937_333#_c_709_n N_A_865_255#_M1017_g 4.6226e-19 $X=6.745 $Y=1.96
+ $X2=0 $Y2=0
cc_624 N_A_937_333#_c_728_n N_A_865_255#_M1017_g 0.00338071f $X=6.98 $Y=2.055
+ $X2=0 $Y2=0
cc_625 N_A_937_333#_M1030_d N_A_1445_69#_c_1330_n 6.77055e-19 $X=6.6 $Y=0.345
+ $X2=0 $Y2=0
cc_626 N_A_937_333#_c_703_n N_A_1445_69#_c_1330_n 0.0503335f $X=6.74 $Y=0.86
+ $X2=0 $Y2=0
cc_627 N_A_937_333#_c_758_p N_A_1445_69#_c_1330_n 0.00159831f $X=6.74 $Y=1.685
+ $X2=0 $Y2=0
cc_628 N_A_937_333#_c_709_n N_A_1445_69#_c_1332_n 0.00148115f $X=6.745 $Y=1.96
+ $X2=0 $Y2=0
cc_629 N_A_937_333#_c_728_n N_A_1445_69#_c_1332_n 0.00799859f $X=6.98 $Y=2.055
+ $X2=0 $Y2=0
cc_630 N_A_937_333#_c_758_p N_A_1445_69#_c_1332_n 0.0130589f $X=6.74 $Y=1.685
+ $X2=0 $Y2=0
cc_631 N_A_937_333#_c_709_n N_A_1445_69#_c_1347_n 0.00450102f $X=6.745 $Y=1.96
+ $X2=0 $Y2=0
cc_632 N_A_937_333#_M1030_d N_A_1445_69#_c_1365_n 0.00177231f $X=6.6 $Y=0.345
+ $X2=0 $Y2=0
cc_633 N_A_937_333#_c_703_n N_A_1445_69#_c_1365_n 0.0137712f $X=6.74 $Y=0.86
+ $X2=0 $Y2=0
cc_634 N_A_937_333#_c_733_n N_A_1445_69#_c_1365_n 0.00256296f $X=6.935 $Y=0.47
+ $X2=0 $Y2=0
cc_635 N_A_937_333#_M1002_g N_VPWR_c_1745_n 0.00380191f $X=4.76 $Y=2.525 $X2=0
+ $Y2=0
cc_636 N_A_937_333#_M1002_g N_VPWR_c_1742_n 9.39239e-19 $X=4.76 $Y=2.525 $X2=0
+ $Y2=0
cc_637 N_A_937_333#_c_733_n N_VGND_c_2013_n 0.016655f $X=6.935 $Y=0.47 $X2=0
+ $Y2=0
cc_638 N_A_937_333#_M1011_g N_VGND_c_2020_n 9.39239e-19 $X=5.35 $Y=0.805 $X2=0
+ $Y2=0
cc_639 N_A_937_333#_c_733_n N_VGND_c_2020_n 0.0160226f $X=6.935 $Y=0.47 $X2=0
+ $Y2=0
cc_640 N_RESET_B_c_803_n N_A_809_463#_M1030_g 0.0145776f $X=5.785 $Y=0.18 $X2=0
+ $Y2=0
cc_641 N_RESET_B_c_817_n N_A_809_463#_M1029_g 0.00946683f $X=6.77 $Y=2.405 $X2=0
+ $Y2=0
cc_642 N_RESET_B_c_818_n N_A_809_463#_M1029_g 0.0121932f $X=6.86 $Y=2.905 $X2=0
+ $Y2=0
cc_643 RESET_B N_A_809_463#_M1029_g 0.00110489f $X=5.915 $Y=1.95 $X2=0 $Y2=0
cc_644 RESET_B N_A_809_463#_M1029_g 2.03955e-19 $X=5.915 $Y=2.32 $X2=0 $Y2=0
cc_645 N_RESET_B_c_826_n N_A_809_463#_M1029_g 0.0124519f $X=5.965 $Y=2.04 $X2=0
+ $Y2=0
cc_646 N_RESET_B_c_802_n N_A_809_463#_c_1010_n 0.00112426f $X=3.845 $Y=1.195
+ $X2=0 $Y2=0
cc_647 N_RESET_B_c_803_n N_A_809_463#_c_1011_n 0.0181063f $X=5.785 $Y=0.18 $X2=0
+ $Y2=0
cc_648 N_RESET_B_M1036_g N_A_809_463#_c_1011_n 0.0167315f $X=5.86 $Y=0.775 $X2=0
+ $Y2=0
cc_649 N_RESET_B_c_808_n N_A_809_463#_c_1011_n 0.00101861f $X=5.845 $Y=1.245
+ $X2=0 $Y2=0
cc_650 N_RESET_B_c_803_n N_A_809_463#_c_1072_n 4.8253e-19 $X=5.785 $Y=0.18 $X2=0
+ $Y2=0
cc_651 N_RESET_B_c_810_n N_A_809_463#_c_1016_n 0.0110165f $X=5.3 $Y=2.205 $X2=0
+ $Y2=0
cc_652 N_RESET_B_c_811_n N_A_809_463#_c_1016_n 0.00856615f $X=5.755 $Y=2.13
+ $X2=0 $Y2=0
cc_653 N_RESET_B_c_812_n N_A_809_463#_c_1016_n 0.00295121f $X=5.375 $Y=2.13
+ $X2=0 $Y2=0
cc_654 RESET_B N_A_809_463#_c_1016_n 0.0128442f $X=5.915 $Y=1.95 $X2=0 $Y2=0
cc_655 RESET_B N_A_809_463#_c_1016_n 0.00131106f $X=5.915 $Y=2.32 $X2=0 $Y2=0
cc_656 N_RESET_B_c_826_n N_A_809_463#_c_1016_n 0.00119816f $X=5.965 $Y=2.04
+ $X2=0 $Y2=0
cc_657 N_RESET_B_c_810_n N_A_809_463#_c_1055_n 0.00493669f $X=5.3 $Y=2.205 $X2=0
+ $Y2=0
cc_658 RESET_B N_A_809_463#_c_1055_n 0.0167518f $X=5.915 $Y=2.32 $X2=0 $Y2=0
cc_659 N_RESET_B_c_826_n N_A_809_463#_c_1055_n 0.0017859f $X=5.965 $Y=2.04 $X2=0
+ $Y2=0
cc_660 N_RESET_B_M1036_g N_A_809_463#_c_1012_n 0.0042921f $X=5.86 $Y=0.775 $X2=0
+ $Y2=0
cc_661 N_RESET_B_c_808_n N_A_809_463#_c_1012_n 5.90867e-19 $X=5.845 $Y=1.245
+ $X2=0 $Y2=0
cc_662 N_RESET_B_c_809_n N_A_809_463#_c_1012_n 0.0016726f $X=5.942 $Y=1.875
+ $X2=0 $Y2=0
cc_663 N_RESET_B_c_816_n N_A_809_463#_c_1017_n 2.15626e-19 $X=3.472 $Y=2.205
+ $X2=0 $Y2=0
cc_664 N_RESET_B_c_808_n N_A_809_463#_c_1013_n 0.00508646f $X=5.845 $Y=1.245
+ $X2=0 $Y2=0
cc_665 N_RESET_B_c_817_n N_A_809_463#_c_1013_n 0.00217187f $X=6.77 $Y=2.405
+ $X2=0 $Y2=0
cc_666 N_RESET_B_c_809_n N_A_809_463#_c_1013_n 0.0240233f $X=5.942 $Y=1.875
+ $X2=0 $Y2=0
cc_667 N_RESET_B_c_802_n N_A_865_255#_M1032_g 0.0182413f $X=3.845 $Y=1.195 $X2=0
+ $Y2=0
cc_668 N_RESET_B_c_803_n N_A_865_255#_M1032_g 0.0100158f $X=5.785 $Y=0.18 $X2=0
+ $Y2=0
cc_669 N_RESET_B_c_810_n N_A_865_255#_c_1139_n 0.0103788f $X=5.3 $Y=2.205 $X2=0
+ $Y2=0
cc_670 N_RESET_B_c_817_n N_A_865_255#_c_1139_n 0.00576009f $X=6.77 $Y=2.405
+ $X2=0 $Y2=0
cc_671 N_RESET_B_c_819_n N_A_865_255#_c_1139_n 0.00187555f $X=8.035 $Y=2.99
+ $X2=0 $Y2=0
cc_672 N_RESET_B_c_820_n N_A_865_255#_c_1139_n 0.0032804f $X=6.95 $Y=2.99 $X2=0
+ $Y2=0
cc_673 RESET_B N_A_865_255#_c_1139_n 0.00172171f $X=5.915 $Y=2.32 $X2=0 $Y2=0
cc_674 N_RESET_B_c_826_n N_A_865_255#_c_1139_n 0.00705851f $X=5.965 $Y=2.04
+ $X2=0 $Y2=0
cc_675 N_RESET_B_c_817_n N_A_865_255#_M1017_g 0.00159845f $X=6.77 $Y=2.405 $X2=0
+ $Y2=0
cc_676 N_RESET_B_c_818_n N_A_865_255#_M1017_g 0.00597242f $X=6.86 $Y=2.905 $X2=0
+ $Y2=0
cc_677 N_RESET_B_c_819_n N_A_865_255#_M1017_g 0.0166502f $X=8.035 $Y=2.99 $X2=0
+ $Y2=0
cc_678 N_RESET_B_c_800_n N_A_865_255#_c_1129_n 0.00212649f $X=3.77 $Y=1.27 $X2=0
+ $Y2=0
cc_679 N_RESET_B_M1005_g N_A_865_255#_c_1131_n 0.0113657f $X=9.015 $Y=0.805
+ $X2=0 $Y2=0
cc_680 N_RESET_B_c_822_n N_A_865_255#_c_1132_n 7.65304e-19 $X=8.94 $Y=2.56 $X2=0
+ $Y2=0
cc_681 N_RESET_B_c_823_n N_A_865_255#_c_1132_n 0.00270012f $X=8.285 $Y=2.56
+ $X2=0 $Y2=0
cc_682 N_RESET_B_c_822_n N_A_865_255#_c_1133_n 0.0021052f $X=8.94 $Y=2.56 $X2=0
+ $Y2=0
cc_683 N_RESET_B_c_823_n N_A_865_255#_c_1133_n 0.00491794f $X=8.285 $Y=2.56
+ $X2=0 $Y2=0
cc_684 N_RESET_B_c_819_n N_A_1445_69#_M1017_d 0.0100894f $X=8.035 $Y=2.99 $X2=0
+ $Y2=0
cc_685 N_RESET_B_M1005_g N_A_1445_69#_c_1324_n 0.0493291f $X=9.015 $Y=0.805
+ $X2=0 $Y2=0
cc_686 N_RESET_B_M1005_g N_A_1445_69#_M1014_g 0.0165272f $X=9.015 $Y=0.805 $X2=0
+ $Y2=0
cc_687 N_RESET_B_c_824_n N_A_1445_69#_M1014_g 3.63139e-19 $X=9.105 $Y=2.34 $X2=0
+ $Y2=0
cc_688 N_RESET_B_c_828_n N_A_1445_69#_M1014_g 0.0291857f $X=9.24 $Y=2.34 $X2=0
+ $Y2=0
cc_689 N_RESET_B_c_819_n N_A_1445_69#_c_1347_n 0.0192863f $X=8.035 $Y=2.99 $X2=0
+ $Y2=0
cc_690 N_RESET_B_c_821_n N_A_1445_69#_c_1347_n 0.00333259f $X=8.16 $Y=2.905
+ $X2=0 $Y2=0
cc_691 N_RESET_B_c_823_n N_A_1445_69#_c_1347_n 0.00710145f $X=8.285 $Y=2.56
+ $X2=0 $Y2=0
cc_692 N_RESET_B_M1005_g N_A_1445_69#_c_1333_n 0.00144176f $X=9.015 $Y=0.805
+ $X2=0 $Y2=0
cc_693 N_RESET_B_M1005_g N_A_1445_69#_c_1339_n 0.00612997f $X=9.015 $Y=0.805
+ $X2=0 $Y2=0
cc_694 N_RESET_B_M1005_g N_A_1445_69#_c_1340_n 0.0136325f $X=9.015 $Y=0.805
+ $X2=0 $Y2=0
cc_695 N_RESET_B_M1005_g N_A_1445_69#_c_1341_n 6.37894e-19 $X=9.015 $Y=0.805
+ $X2=0 $Y2=0
cc_696 N_RESET_B_M1005_g N_A_1641_21#_M1020_g 0.00650034f $X=9.015 $Y=0.805
+ $X2=0 $Y2=0
cc_697 N_RESET_B_M1023_g N_A_1641_21#_M1031_g 0.00539753f $X=9.24 $Y=2.875 $X2=0
+ $Y2=0
cc_698 N_RESET_B_c_821_n N_A_1641_21#_M1031_g 0.00203145f $X=8.16 $Y=2.905 $X2=0
+ $Y2=0
cc_699 N_RESET_B_c_822_n N_A_1641_21#_M1031_g 0.014631f $X=8.94 $Y=2.56 $X2=0
+ $Y2=0
cc_700 N_RESET_B_c_824_n N_A_1641_21#_M1031_g 4.93381e-19 $X=9.105 $Y=2.34 $X2=0
+ $Y2=0
cc_701 N_RESET_B_c_828_n N_A_1641_21#_M1031_g 0.00260658f $X=9.24 $Y=2.34 $X2=0
+ $Y2=0
cc_702 N_RESET_B_M1005_g N_A_1641_21#_c_1529_n 0.0104164f $X=9.015 $Y=0.805
+ $X2=0 $Y2=0
cc_703 N_RESET_B_M1005_g N_A_1641_21#_c_1531_n 0.0416539f $X=9.015 $Y=0.805
+ $X2=0 $Y2=0
cc_704 N_RESET_B_c_828_n N_A_1641_21#_c_1533_n 0.0416539f $X=9.24 $Y=2.34 $X2=0
+ $Y2=0
cc_705 N_RESET_B_M1005_g N_A_1641_21#_c_1540_n 0.0110596f $X=9.015 $Y=0.805
+ $X2=0 $Y2=0
cc_706 N_RESET_B_c_822_n N_A_1641_21#_c_1540_n 0.00871457f $X=8.94 $Y=2.56 $X2=0
+ $Y2=0
cc_707 N_RESET_B_c_824_n N_A_1641_21#_c_1540_n 0.0235408f $X=9.105 $Y=2.34 $X2=0
+ $Y2=0
cc_708 N_RESET_B_c_828_n N_A_1641_21#_c_1540_n 0.0068676f $X=9.24 $Y=2.34 $X2=0
+ $Y2=0
cc_709 N_RESET_B_M1005_g N_A_1641_21#_c_1534_n 0.00143992f $X=9.015 $Y=0.805
+ $X2=0 $Y2=0
cc_710 N_RESET_B_M1005_g N_A_1641_21#_c_1541_n 0.00124496f $X=9.015 $Y=0.805
+ $X2=0 $Y2=0
cc_711 N_RESET_B_c_822_n N_A_1641_21#_c_1541_n 0.0245636f $X=8.94 $Y=2.56 $X2=0
+ $Y2=0
cc_712 N_RESET_B_c_824_n N_A_1641_21#_c_1541_n 0.00319592f $X=9.105 $Y=2.34
+ $X2=0 $Y2=0
cc_713 N_RESET_B_M1005_g N_A_1641_21#_c_1542_n 0.00179189f $X=9.015 $Y=0.805
+ $X2=0 $Y2=0
cc_714 N_RESET_B_c_824_n N_A_1641_21#_c_1542_n 0.027831f $X=9.105 $Y=2.34 $X2=0
+ $Y2=0
cc_715 N_RESET_B_c_828_n N_A_1641_21#_c_1542_n 0.0064406f $X=9.24 $Y=2.34 $X2=0
+ $Y2=0
cc_716 N_RESET_B_c_822_n N_A_1641_21#_c_1543_n 0.00680303f $X=8.94 $Y=2.56 $X2=0
+ $Y2=0
cc_717 N_RESET_B_c_824_n N_A_1641_21#_c_1543_n 6.45583e-19 $X=9.105 $Y=2.34
+ $X2=0 $Y2=0
cc_718 N_RESET_B_c_817_n N_VPWR_M1029_s 0.0109208f $X=6.77 $Y=2.405 $X2=0 $Y2=0
cc_719 N_RESET_B_c_816_n N_VPWR_c_1744_n 0.00366409f $X=3.472 $Y=2.205 $X2=0
+ $Y2=0
cc_720 N_RESET_B_c_810_n N_VPWR_c_1745_n 0.00380191f $X=5.3 $Y=2.205 $X2=0 $Y2=0
cc_721 N_RESET_B_c_817_n N_VPWR_c_1746_n 0.0261586f $X=6.77 $Y=2.405 $X2=0 $Y2=0
cc_722 N_RESET_B_c_818_n N_VPWR_c_1746_n 0.0185722f $X=6.86 $Y=2.905 $X2=0 $Y2=0
cc_723 N_RESET_B_c_820_n N_VPWR_c_1746_n 0.0150384f $X=6.95 $Y=2.99 $X2=0 $Y2=0
cc_724 N_RESET_B_M1023_g N_VPWR_c_1747_n 0.00401442f $X=9.24 $Y=2.875 $X2=0
+ $Y2=0
cc_725 N_RESET_B_c_824_n N_VPWR_c_1747_n 0.00109044f $X=9.105 $Y=2.34 $X2=0
+ $Y2=0
cc_726 N_RESET_B_c_816_n N_VPWR_c_1754_n 0.00456028f $X=3.472 $Y=2.205 $X2=0
+ $Y2=0
cc_727 N_RESET_B_c_810_n N_VPWR_c_1742_n 9.39239e-19 $X=5.3 $Y=2.205 $X2=0 $Y2=0
cc_728 N_RESET_B_M1023_g N_VPWR_c_1742_n 0.00572364f $X=9.24 $Y=2.875 $X2=0
+ $Y2=0
cc_729 N_RESET_B_c_816_n N_VPWR_c_1742_n 0.00544287f $X=3.472 $Y=2.205 $X2=0
+ $Y2=0
cc_730 N_RESET_B_c_817_n N_VPWR_c_1742_n 0.0103534f $X=6.77 $Y=2.405 $X2=0 $Y2=0
cc_731 N_RESET_B_c_819_n N_VPWR_c_1742_n 0.0483908f $X=8.035 $Y=2.99 $X2=0 $Y2=0
cc_732 N_RESET_B_c_820_n N_VPWR_c_1742_n 0.00617437f $X=6.95 $Y=2.99 $X2=0 $Y2=0
cc_733 N_RESET_B_c_822_n N_VPWR_c_1742_n 0.00621154f $X=8.94 $Y=2.56 $X2=0 $Y2=0
cc_734 N_RESET_B_c_824_n N_VPWR_c_1742_n 0.00298381f $X=9.105 $Y=2.34 $X2=0
+ $Y2=0
cc_735 RESET_B N_VPWR_c_1742_n 0.0109472f $X=5.915 $Y=2.32 $X2=0 $Y2=0
cc_736 N_RESET_B_c_826_n N_VPWR_c_1742_n 2.88589e-19 $X=5.965 $Y=2.04 $X2=0
+ $Y2=0
cc_737 N_RESET_B_c_819_n N_VPWR_c_1763_n 0.0822086f $X=8.035 $Y=2.99 $X2=0 $Y2=0
cc_738 N_RESET_B_c_820_n N_VPWR_c_1763_n 0.012271f $X=6.95 $Y=2.99 $X2=0 $Y2=0
cc_739 N_RESET_B_c_822_n N_VPWR_c_1763_n 0.00254602f $X=8.94 $Y=2.56 $X2=0 $Y2=0
cc_740 N_RESET_B_M1023_g N_VPWR_c_1764_n 0.00774085f $X=9.24 $Y=2.875 $X2=0
+ $Y2=0
cc_741 N_RESET_B_c_822_n N_VPWR_c_1764_n 0.0292342f $X=8.94 $Y=2.56 $X2=0 $Y2=0
cc_742 N_RESET_B_c_824_n N_VPWR_c_1764_n 0.0149618f $X=9.105 $Y=2.34 $X2=0 $Y2=0
cc_743 N_RESET_B_c_828_n N_VPWR_c_1764_n 0.00109075f $X=9.24 $Y=2.34 $X2=0 $Y2=0
cc_744 N_RESET_B_M1027_g N_A_380_50#_c_1892_n 0.0115341f $X=3.32 $Y=0.615 $X2=0
+ $Y2=0
cc_745 N_RESET_B_c_801_n N_A_380_50#_c_1892_n 0.00216999f $X=3.575 $Y=1.27 $X2=0
+ $Y2=0
cc_746 N_RESET_B_c_816_n N_A_380_50#_c_1899_n 0.0110849f $X=3.472 $Y=2.205 $X2=0
+ $Y2=0
cc_747 N_RESET_B_c_800_n N_A_380_50#_c_1893_n 0.00838538f $X=3.77 $Y=1.27 $X2=0
+ $Y2=0
cc_748 N_RESET_B_c_801_n N_A_380_50#_c_1893_n 0.00421167f $X=3.575 $Y=1.27 $X2=0
+ $Y2=0
cc_749 N_RESET_B_c_802_n N_A_380_50#_c_1893_n 0.00458732f $X=3.845 $Y=1.195
+ $X2=0 $Y2=0
cc_750 N_RESET_B_c_806_n N_A_380_50#_c_1893_n 0.0169624f $X=3.472 $Y=2.055 $X2=0
+ $Y2=0
cc_751 N_RESET_B_c_816_n N_A_380_50#_c_1893_n 0.00788658f $X=3.472 $Y=2.205
+ $X2=0 $Y2=0
cc_752 N_RESET_B_c_800_n N_A_380_50#_c_1894_n 0.00275463f $X=3.77 $Y=1.27 $X2=0
+ $Y2=0
cc_753 N_RESET_B_c_802_n N_A_380_50#_c_1894_n 0.0130583f $X=3.845 $Y=1.195 $X2=0
+ $Y2=0
cc_754 N_RESET_B_c_798_n N_A_380_50#_c_1949_n 7.16211e-19 $X=3.77 $Y=0.18 $X2=0
+ $Y2=0
cc_755 N_RESET_B_c_816_n N_A_380_50#_c_1898_n 0.005409f $X=3.472 $Y=2.205 $X2=0
+ $Y2=0
cc_756 N_RESET_B_c_802_n N_A_380_50#_c_1936_n 0.00445987f $X=3.845 $Y=1.195
+ $X2=0 $Y2=0
cc_757 N_RESET_B_c_803_n N_A_380_50#_c_1936_n 0.00359058f $X=5.785 $Y=0.18 $X2=0
+ $Y2=0
cc_758 N_RESET_B_c_819_n A_1578_533# 0.00648492f $X=8.035 $Y=2.99 $X2=-0.19
+ $Y2=-0.245
cc_759 N_RESET_B_c_821_n A_1578_533# 0.00463087f $X=8.16 $Y=2.905 $X2=-0.19
+ $Y2=-0.245
cc_760 N_RESET_B_M1027_g N_VGND_c_2006_n 0.00291064f $X=3.32 $Y=0.615 $X2=0
+ $Y2=0
cc_761 N_RESET_B_c_798_n N_VGND_c_2006_n 0.0217677f $X=3.77 $Y=0.18 $X2=0 $Y2=0
cc_762 N_RESET_B_c_801_n N_VGND_c_2006_n 7.97771e-19 $X=3.575 $Y=1.27 $X2=0
+ $Y2=0
cc_763 N_RESET_B_c_802_n N_VGND_c_2006_n 0.00842416f $X=3.845 $Y=1.195 $X2=0
+ $Y2=0
cc_764 N_RESET_B_c_803_n N_VGND_c_2007_n 0.0128616f $X=5.785 $Y=0.18 $X2=0 $Y2=0
cc_765 N_RESET_B_M1005_g N_VGND_c_2008_n 0.00762837f $X=9.015 $Y=0.805 $X2=0
+ $Y2=0
cc_766 N_RESET_B_c_798_n N_VGND_c_2011_n 0.0774159f $X=3.77 $Y=0.18 $X2=0 $Y2=0
cc_767 N_RESET_B_c_799_n N_VGND_c_2016_n 0.00620508f $X=3.395 $Y=0.18 $X2=0
+ $Y2=0
cc_768 N_RESET_B_c_798_n N_VGND_c_2020_n 0.00127851f $X=3.77 $Y=0.18 $X2=0 $Y2=0
cc_769 N_RESET_B_c_799_n N_VGND_c_2020_n 0.0068511f $X=3.395 $Y=0.18 $X2=0 $Y2=0
cc_770 N_RESET_B_c_803_n N_VGND_c_2020_n 0.0647347f $X=5.785 $Y=0.18 $X2=0 $Y2=0
cc_771 N_RESET_B_M1005_g N_VGND_c_2020_n 9.39239e-19 $X=9.015 $Y=0.805 $X2=0
+ $Y2=0
cc_772 N_RESET_B_c_807_n N_VGND_c_2020_n 0.00458272f $X=3.845 $Y=0.18 $X2=0
+ $Y2=0
cc_773 N_RESET_B_M1027_g N_noxref_24_c_2145_n 0.00137979f $X=3.32 $Y=0.615 $X2=0
+ $Y2=0
cc_774 N_A_809_463#_c_1010_n N_A_865_255#_M1037_g 0.0158999f $X=4.47 $Y=2.085
+ $X2=0 $Y2=0
cc_775 N_A_809_463#_c_1017_n N_A_865_255#_M1037_g 0.0241535f $X=4.287 $Y=2.25
+ $X2=0 $Y2=0
cc_776 N_A_809_463#_c_1010_n N_A_865_255#_M1032_g 0.00713908f $X=4.47 $Y=2.085
+ $X2=0 $Y2=0
cc_777 N_A_809_463#_c_1072_n N_A_865_255#_M1032_g 0.00535849f $X=4.555 $Y=0.89
+ $X2=0 $Y2=0
cc_778 N_A_809_463#_M1029_g N_A_865_255#_c_1139_n 0.00990589f $X=6.765 $Y=2.315
+ $X2=0 $Y2=0
cc_779 N_A_809_463#_c_1055_n N_A_865_255#_c_1139_n 0.00451434f $X=5.515 $Y=2.525
+ $X2=0 $Y2=0
cc_780 N_A_809_463#_M1029_g N_A_865_255#_c_1126_n 0.0358468f $X=6.765 $Y=2.315
+ $X2=0 $Y2=0
cc_781 N_A_809_463#_c_1010_n N_A_865_255#_c_1129_n 0.00415492f $X=4.47 $Y=2.085
+ $X2=0 $Y2=0
cc_782 N_A_809_463#_c_1013_n N_A_1445_69#_c_1330_n 0.00355274f $X=6.525 $Y=1.402
+ $X2=0 $Y2=0
cc_783 N_A_809_463#_c_1013_n N_A_1445_69#_c_1332_n 0.00134266f $X=6.525 $Y=1.402
+ $X2=0 $Y2=0
cc_784 N_A_809_463#_c_1016_n N_VPWR_M1002_d 0.00296548f $X=5.365 $Y=2.25 $X2=0
+ $Y2=0
cc_785 N_A_809_463#_c_1016_n N_VPWR_c_1745_n 0.022455f $X=5.365 $Y=2.25 $X2=0
+ $Y2=0
cc_786 N_A_809_463#_M1029_g N_VPWR_c_1746_n 0.00439533f $X=6.765 $Y=2.315 $X2=0
+ $Y2=0
cc_787 N_A_809_463#_c_1055_n N_VPWR_c_1746_n 9.26185e-19 $X=5.515 $Y=2.525 $X2=0
+ $Y2=0
cc_788 N_A_809_463#_c_1017_n N_VPWR_c_1754_n 0.00572098f $X=4.287 $Y=2.25 $X2=0
+ $Y2=0
cc_789 N_A_809_463#_c_1055_n N_VPWR_c_1755_n 0.00438561f $X=5.515 $Y=2.525 $X2=0
+ $Y2=0
cc_790 N_A_809_463#_M1029_g N_VPWR_c_1742_n 5.03388e-19 $X=6.765 $Y=2.315 $X2=0
+ $Y2=0
cc_791 N_A_809_463#_c_1055_n N_VPWR_c_1742_n 0.00679974f $X=5.515 $Y=2.525 $X2=0
+ $Y2=0
cc_792 N_A_809_463#_c_1017_n N_VPWR_c_1742_n 0.0106108f $X=4.287 $Y=2.25 $X2=0
+ $Y2=0
cc_793 N_A_809_463#_c_1017_n N_A_380_50#_c_1893_n 0.0101187f $X=4.287 $Y=2.25
+ $X2=0 $Y2=0
cc_794 N_A_809_463#_c_1017_n N_A_380_50#_c_1898_n 0.028653f $X=4.287 $Y=2.25
+ $X2=0 $Y2=0
cc_795 N_A_809_463#_c_1072_n N_A_380_50#_c_1936_n 0.0158998f $X=4.555 $Y=0.89
+ $X2=0 $Y2=0
cc_796 N_A_809_463#_c_1016_n A_895_463# 0.0027472f $X=5.365 $Y=2.25 $X2=-0.19
+ $Y2=-0.245
cc_797 N_A_809_463#_c_1017_n A_895_463# 0.00103754f $X=4.287 $Y=2.25 $X2=-0.19
+ $Y2=-0.245
cc_798 N_A_809_463#_c_1011_n N_VGND_M1036_d 0.00736874f $X=6.145 $Y=0.89 $X2=0
+ $Y2=0
cc_799 N_A_809_463#_M1030_g N_VGND_c_2007_n 0.00840693f $X=6.525 $Y=0.665 $X2=0
+ $Y2=0
cc_800 N_A_809_463#_c_1011_n N_VGND_c_2007_n 0.0229474f $X=6.145 $Y=0.89 $X2=0
+ $Y2=0
cc_801 N_A_809_463#_c_1013_n N_VGND_c_2007_n 9.9456e-19 $X=6.525 $Y=1.402 $X2=0
+ $Y2=0
cc_802 N_A_809_463#_M1030_g N_VGND_c_2013_n 0.00400407f $X=6.525 $Y=0.665 $X2=0
+ $Y2=0
cc_803 N_A_809_463#_M1030_g N_VGND_c_2020_n 0.00784291f $X=6.525 $Y=0.665 $X2=0
+ $Y2=0
cc_804 N_A_809_463#_c_1011_n N_VGND_c_2020_n 0.0531105f $X=6.145 $Y=0.89 $X2=0
+ $Y2=0
cc_805 N_A_809_463#_c_1072_n N_VGND_c_2020_n 0.0057931f $X=4.555 $Y=0.89 $X2=0
+ $Y2=0
cc_806 N_A_809_463#_c_1011_n A_991_119# 0.0042163f $X=6.145 $Y=0.89 $X2=-0.19
+ $Y2=-0.245
cc_807 N_A_809_463#_c_1011_n A_1085_119# 0.00569011f $X=6.145 $Y=0.89 $X2=-0.19
+ $Y2=-0.245
cc_808 N_A_865_255#_c_1131_n N_A_1445_69#_M1014_g 0.0165829f $X=9.8 $Y=1.64
+ $X2=0 $Y2=0
cc_809 N_A_865_255#_c_1147_n N_A_1445_69#_M1014_g 0.0176576f $X=9.922 $Y=2.37
+ $X2=0 $Y2=0
cc_810 N_A_865_255#_c_1149_n N_A_1445_69#_M1014_g 0.00395151f $X=10.045 $Y=2.455
+ $X2=0 $Y2=0
cc_811 N_A_865_255#_c_1137_n N_A_1445_69#_c_1328_n 6.84226e-19 $X=11.465 $Y=1.08
+ $X2=0 $Y2=0
cc_812 N_A_865_255#_c_1126_n N_A_1445_69#_c_1330_n 2.60926e-19 $X=7.27 $Y=1.71
+ $X2=0 $Y2=0
cc_813 N_A_865_255#_M1012_g N_A_1445_69#_c_1330_n 0.00161093f $X=7.92 $Y=0.775
+ $X2=0 $Y2=0
cc_814 N_A_865_255#_M1012_g N_A_1445_69#_c_1331_n 0.00608452f $X=7.92 $Y=0.775
+ $X2=0 $Y2=0
cc_815 N_A_865_255#_M1017_g N_A_1445_69#_c_1332_n 0.00591326f $X=7.195 $Y=2.315
+ $X2=0 $Y2=0
cc_816 N_A_865_255#_c_1125_n N_A_1445_69#_c_1332_n 0.0112761f $X=7.815 $Y=1.71
+ $X2=0 $Y2=0
cc_817 N_A_865_255#_c_1126_n N_A_1445_69#_c_1332_n 0.00394125f $X=7.27 $Y=1.71
+ $X2=0 $Y2=0
cc_818 N_A_865_255#_M1017_g N_A_1445_69#_c_1347_n 0.00346759f $X=7.195 $Y=2.315
+ $X2=0 $Y2=0
cc_819 N_A_865_255#_c_1125_n N_A_1445_69#_c_1347_n 0.00692494f $X=7.815 $Y=1.71
+ $X2=0 $Y2=0
cc_820 N_A_865_255#_M1012_g N_A_1445_69#_c_1363_n 0.00953108f $X=7.92 $Y=0.775
+ $X2=0 $Y2=0
cc_821 N_A_865_255#_c_1132_n N_A_1445_69#_c_1363_n 0.00217205f $X=8.205 $Y=1.65
+ $X2=0 $Y2=0
cc_822 N_A_865_255#_M1012_g N_A_1445_69#_c_1333_n 0.00419106f $X=7.92 $Y=0.775
+ $X2=0 $Y2=0
cc_823 N_A_865_255#_M1012_g N_A_1445_69#_c_1334_n 0.00169264f $X=7.92 $Y=0.775
+ $X2=0 $Y2=0
cc_824 N_A_865_255#_c_1132_n N_A_1445_69#_c_1334_n 0.00272642f $X=8.205 $Y=1.65
+ $X2=0 $Y2=0
cc_825 N_A_865_255#_c_1133_n N_A_1445_69#_c_1334_n 0.0131781f $X=8.37 $Y=1.65
+ $X2=0 $Y2=0
cc_826 N_A_865_255#_M1010_g N_A_1445_69#_c_1335_n 0.00289536f $X=10.625 $Y=0.785
+ $X2=0 $Y2=0
cc_827 N_A_865_255#_M1007_d N_A_1445_69#_c_1336_n 0.00717153f $X=11.325 $Y=0.365
+ $X2=0 $Y2=0
cc_828 N_A_865_255#_M1010_g N_A_1445_69#_c_1336_n 0.0184046f $X=10.625 $Y=0.785
+ $X2=0 $Y2=0
cc_829 N_A_865_255#_c_1134_n N_A_1445_69#_c_1336_n 0.0149579f $X=10.8 $Y=1.51
+ $X2=0 $Y2=0
cc_830 N_A_865_255#_c_1135_n N_A_1445_69#_c_1336_n 0.00119574f $X=10.8 $Y=1.51
+ $X2=0 $Y2=0
cc_831 N_A_865_255#_c_1137_n N_A_1445_69#_c_1336_n 0.0268345f $X=11.465 $Y=1.08
+ $X2=0 $Y2=0
cc_832 N_A_865_255#_c_1131_n N_A_1445_69#_c_1339_n 0.0054896f $X=9.8 $Y=1.64
+ $X2=0 $Y2=0
cc_833 N_A_865_255#_c_1131_n N_A_1445_69#_c_1340_n 0.0470246f $X=9.8 $Y=1.64
+ $X2=0 $Y2=0
cc_834 N_A_865_255#_c_1132_n N_A_1445_69#_c_1340_n 2.57398e-19 $X=8.205 $Y=1.65
+ $X2=0 $Y2=0
cc_835 N_A_865_255#_c_1133_n N_A_1445_69#_c_1340_n 0.00302141f $X=8.37 $Y=1.65
+ $X2=0 $Y2=0
cc_836 N_A_865_255#_c_1131_n N_A_1445_69#_c_1341_n 0.0400225f $X=9.8 $Y=1.64
+ $X2=0 $Y2=0
cc_837 N_A_865_255#_c_1137_n N_A_1445_69#_c_1342_n 0.0161073f $X=11.465 $Y=1.08
+ $X2=0 $Y2=0
cc_838 N_A_865_255#_c_1137_n N_A_1445_69#_c_1343_n 3.77762e-19 $X=11.465 $Y=1.08
+ $X2=0 $Y2=0
cc_839 N_A_865_255#_M1012_g N_A_1641_21#_M1020_g 0.0493683f $X=7.92 $Y=0.775
+ $X2=0 $Y2=0
cc_840 N_A_865_255#_c_1131_n N_A_1641_21#_c_1531_n 0.0012061f $X=9.8 $Y=1.64
+ $X2=0 $Y2=0
cc_841 N_A_865_255#_c_1132_n N_A_1641_21#_c_1532_n 0.00871161f $X=8.205 $Y=1.65
+ $X2=0 $Y2=0
cc_842 N_A_865_255#_M1012_g N_A_1641_21#_c_1533_n 0.00311257f $X=7.92 $Y=0.775
+ $X2=0 $Y2=0
cc_843 N_A_865_255#_c_1131_n N_A_1641_21#_c_1533_n 0.00989616f $X=9.8 $Y=1.64
+ $X2=0 $Y2=0
cc_844 N_A_865_255#_c_1132_n N_A_1641_21#_c_1533_n 0.0205906f $X=8.205 $Y=1.65
+ $X2=0 $Y2=0
cc_845 N_A_865_255#_c_1133_n N_A_1641_21#_c_1533_n 0.00106005f $X=8.37 $Y=1.65
+ $X2=0 $Y2=0
cc_846 N_A_865_255#_c_1131_n N_A_1641_21#_c_1540_n 0.0621052f $X=9.8 $Y=1.64
+ $X2=0 $Y2=0
cc_847 N_A_865_255#_c_1147_n N_A_1641_21#_c_1540_n 0.0133575f $X=9.922 $Y=2.37
+ $X2=0 $Y2=0
cc_848 N_A_865_255#_M1010_g N_A_1641_21#_c_1536_n 8.44356e-19 $X=10.625 $Y=0.785
+ $X2=0 $Y2=0
cc_849 N_A_865_255#_c_1131_n N_A_1641_21#_c_1541_n 0.0187519f $X=9.8 $Y=1.64
+ $X2=0 $Y2=0
cc_850 N_A_865_255#_c_1147_n N_A_1641_21#_c_1542_n 0.0207473f $X=9.922 $Y=2.37
+ $X2=0 $Y2=0
cc_851 N_A_865_255#_c_1149_n N_A_1641_21#_c_1542_n 0.0131377f $X=10.045 $Y=2.455
+ $X2=0 $Y2=0
cc_852 N_A_865_255#_c_1131_n N_A_1641_21#_c_1543_n 0.00210664f $X=9.8 $Y=1.64
+ $X2=0 $Y2=0
cc_853 N_A_865_255#_c_1132_n N_A_1641_21#_c_1543_n 0.00236994f $X=8.205 $Y=1.65
+ $X2=0 $Y2=0
cc_854 N_A_865_255#_c_1133_n N_A_1641_21#_c_1543_n 2.06019e-19 $X=8.37 $Y=1.65
+ $X2=0 $Y2=0
cc_855 N_A_865_255#_M1010_g N_A_1641_21#_c_1537_n 0.00818731f $X=10.625 $Y=0.785
+ $X2=0 $Y2=0
cc_856 N_A_865_255#_M1010_g N_CLK_M1007_g 0.0257363f $X=10.625 $Y=0.785 $X2=0
+ $Y2=0
cc_857 N_A_865_255#_c_1136_n N_CLK_M1007_g 0.00677384f $X=11.047 $Y=1.345 $X2=0
+ $Y2=0
cc_858 N_A_865_255#_c_1137_n N_CLK_M1007_g 0.00735731f $X=11.465 $Y=1.08 $X2=0
+ $Y2=0
cc_859 N_A_865_255#_M1035_g N_CLK_M1018_g 0.0329588f $X=10.665 $Y=2.465 $X2=0
+ $Y2=0
cc_860 N_A_865_255#_c_1150_n N_CLK_M1018_g 0.0313823f $X=11.047 $Y=2.37 $X2=0
+ $Y2=0
cc_861 N_A_865_255#_c_1134_n N_CLK_M1018_g 0.00475944f $X=10.8 $Y=1.51 $X2=0
+ $Y2=0
cc_862 N_A_865_255#_c_1154_n N_CLK_M1018_g 0.0191568f $X=11.21 $Y=2.455 $X2=0
+ $Y2=0
cc_863 N_A_865_255#_c_1134_n N_CLK_c_1643_n 0.0078678f $X=10.8 $Y=1.51 $X2=0
+ $Y2=0
cc_864 N_A_865_255#_c_1137_n N_CLK_c_1643_n 0.00786529f $X=11.465 $Y=1.08 $X2=0
+ $Y2=0
cc_865 N_A_865_255#_c_1134_n N_CLK_c_1644_n 0.00417528f $X=10.8 $Y=1.51 $X2=0
+ $Y2=0
cc_866 N_A_865_255#_c_1135_n N_CLK_c_1644_n 0.0213966f $X=10.8 $Y=1.51 $X2=0
+ $Y2=0
cc_867 N_A_865_255#_c_1134_n N_CLK_c_1645_n 0.0011306f $X=10.8 $Y=1.51 $X2=0
+ $Y2=0
cc_868 N_A_865_255#_M1018_d N_CLK_c_1648_n 0.00760995f $X=11.325 $Y=1.835 $X2=0
+ $Y2=0
cc_869 N_A_865_255#_c_1134_n N_CLK_c_1648_n 0.0560592f $X=10.8 $Y=1.51 $X2=0
+ $Y2=0
cc_870 N_A_865_255#_c_1154_n N_CLK_c_1648_n 0.00661425f $X=11.21 $Y=2.455 $X2=0
+ $Y2=0
cc_871 N_A_865_255#_c_1137_n N_CLK_c_1648_n 0.0048381f $X=11.465 $Y=1.08 $X2=0
+ $Y2=0
cc_872 N_A_865_255#_c_1150_n N_VPWR_M1035_d 0.00213375f $X=11.047 $Y=2.37 $X2=0
+ $Y2=0
cc_873 N_A_865_255#_c_1154_n N_VPWR_M1035_d 0.00513142f $X=11.21 $Y=2.455 $X2=0
+ $Y2=0
cc_874 N_A_865_255#_M1037_g N_VPWR_c_1745_n 0.00676916f $X=4.4 $Y=2.525 $X2=0
+ $Y2=0
cc_875 N_A_865_255#_c_1139_n N_VPWR_c_1745_n 0.0256837f $X=7.12 $Y=3.15 $X2=0
+ $Y2=0
cc_876 N_A_865_255#_c_1139_n N_VPWR_c_1746_n 0.0252913f $X=7.12 $Y=3.15 $X2=0
+ $Y2=0
cc_877 N_A_865_255#_M1017_g N_VPWR_c_1746_n 6.6829e-19 $X=7.195 $Y=2.315 $X2=0
+ $Y2=0
cc_878 N_A_865_255#_M1035_g N_VPWR_c_1748_n 0.00718041f $X=10.665 $Y=2.465 $X2=0
+ $Y2=0
cc_879 N_A_865_255#_c_1149_n N_VPWR_c_1748_n 0.0218849f $X=10.045 $Y=2.455 $X2=0
+ $Y2=0
cc_880 N_A_865_255#_M1035_g N_VPWR_c_1749_n 0.0133121f $X=10.665 $Y=2.465 $X2=0
+ $Y2=0
cc_881 N_A_865_255#_c_1154_n N_VPWR_c_1749_n 0.0414242f $X=11.21 $Y=2.455 $X2=0
+ $Y2=0
cc_882 N_A_865_255#_c_1140_n N_VPWR_c_1754_n 0.0192779f $X=4.475 $Y=3.15 $X2=0
+ $Y2=0
cc_883 N_A_865_255#_c_1139_n N_VPWR_c_1755_n 0.0351105f $X=7.12 $Y=3.15 $X2=0
+ $Y2=0
cc_884 N_A_865_255#_M1035_g N_VPWR_c_1756_n 0.00486043f $X=10.665 $Y=2.465 $X2=0
+ $Y2=0
cc_885 N_A_865_255#_c_1154_n N_VPWR_c_1757_n 0.0139486f $X=11.21 $Y=2.455 $X2=0
+ $Y2=0
cc_886 N_A_865_255#_M1018_d N_VPWR_c_1742_n 0.0023243f $X=11.325 $Y=1.835 $X2=0
+ $Y2=0
cc_887 N_A_865_255#_c_1139_n N_VPWR_c_1742_n 0.0713545f $X=7.12 $Y=3.15 $X2=0
+ $Y2=0
cc_888 N_A_865_255#_c_1140_n N_VPWR_c_1742_n 0.00962546f $X=4.475 $Y=3.15 $X2=0
+ $Y2=0
cc_889 N_A_865_255#_M1035_g N_VPWR_c_1742_n 0.00589841f $X=10.665 $Y=2.465 $X2=0
+ $Y2=0
cc_890 N_A_865_255#_c_1148_n N_VPWR_c_1742_n 0.0231335f $X=10.715 $Y=2.455 $X2=0
+ $Y2=0
cc_891 N_A_865_255#_c_1149_n N_VPWR_c_1742_n 9.61647e-19 $X=10.045 $Y=2.455
+ $X2=0 $Y2=0
cc_892 N_A_865_255#_c_1154_n N_VPWR_c_1742_n 0.022291f $X=11.21 $Y=2.455 $X2=0
+ $Y2=0
cc_893 N_A_865_255#_c_1139_n N_VPWR_c_1763_n 0.0169195f $X=7.12 $Y=3.15 $X2=0
+ $Y2=0
cc_894 N_A_865_255#_M1037_g N_A_380_50#_c_1893_n 4.84158e-19 $X=4.4 $Y=2.525
+ $X2=0 $Y2=0
cc_895 N_A_865_255#_M1032_g N_A_380_50#_c_1893_n 9.22186e-19 $X=4.45 $Y=0.805
+ $X2=0 $Y2=0
cc_896 N_A_865_255#_M1037_g N_A_380_50#_c_1898_n 0.0028431f $X=4.4 $Y=2.525
+ $X2=0 $Y2=0
cc_897 N_A_865_255#_M1032_g N_A_380_50#_c_1936_n 0.0045374f $X=4.45 $Y=0.805
+ $X2=0 $Y2=0
cc_898 N_A_865_255#_M1010_g N_VGND_c_2009_n 0.00302439f $X=10.625 $Y=0.785 $X2=0
+ $Y2=0
cc_899 N_A_865_255#_M1012_g N_VGND_c_2013_n 0.00352658f $X=7.92 $Y=0.775 $X2=0
+ $Y2=0
cc_900 N_A_865_255#_M1010_g N_VGND_c_2017_n 0.00330473f $X=10.625 $Y=0.785 $X2=0
+ $Y2=0
cc_901 N_A_865_255#_M1032_g N_VGND_c_2020_n 9.39239e-19 $X=4.45 $Y=0.805 $X2=0
+ $Y2=0
cc_902 N_A_865_255#_M1012_g N_VGND_c_2020_n 0.00486331f $X=7.92 $Y=0.775 $X2=0
+ $Y2=0
cc_903 N_A_865_255#_M1010_g N_VGND_c_2020_n 0.00428598f $X=10.625 $Y=0.785 $X2=0
+ $Y2=0
cc_904 N_A_1445_69#_c_1331_n N_A_1641_21#_M1020_g 0.00276775f $X=7.365 $Y=0.49
+ $X2=0 $Y2=0
cc_905 N_A_1445_69#_c_1363_n N_A_1641_21#_M1020_g 0.00729768f $X=8.11 $Y=0.83
+ $X2=0 $Y2=0
cc_906 N_A_1445_69#_c_1333_n N_A_1641_21#_M1020_g 0.00553937f $X=8.215 $Y=1.135
+ $X2=0 $Y2=0
cc_907 N_A_1445_69#_c_1324_n N_A_1641_21#_c_1529_n 0.0103024f $X=9.375 $Y=1.125
+ $X2=0 $Y2=0
cc_908 N_A_1445_69#_c_1340_n N_A_1641_21#_c_1531_n 0.0145012f $X=9.48 $Y=1.26
+ $X2=0 $Y2=0
cc_909 N_A_1445_69#_c_1333_n N_A_1641_21#_c_1532_n 0.00135109f $X=8.215 $Y=1.135
+ $X2=0 $Y2=0
cc_910 N_A_1445_69#_c_1334_n N_A_1641_21#_c_1532_n 0.00210503f $X=8.32 $Y=1.22
+ $X2=0 $Y2=0
cc_911 N_A_1445_69#_c_1340_n N_A_1641_21#_c_1532_n 0.00198519f $X=9.48 $Y=1.26
+ $X2=0 $Y2=0
cc_912 N_A_1445_69#_c_1340_n N_A_1641_21#_c_1533_n 0.00299173f $X=9.48 $Y=1.26
+ $X2=0 $Y2=0
cc_913 N_A_1445_69#_M1014_g N_A_1641_21#_c_1540_n 0.00525337f $X=9.67 $Y=2.875
+ $X2=0 $Y2=0
cc_914 N_A_1445_69#_c_1324_n N_A_1641_21#_c_1534_n 0.0114379f $X=9.375 $Y=1.125
+ $X2=0 $Y2=0
cc_915 N_A_1445_69#_c_1335_n N_A_1641_21#_c_1534_n 0.0114797f $X=9.96 $Y=1.135
+ $X2=0 $Y2=0
cc_916 N_A_1445_69#_c_1337_n N_A_1641_21#_c_1534_n 0.0146126f $X=10.045 $Y=0.73
+ $X2=0 $Y2=0
cc_917 N_A_1445_69#_c_1339_n N_A_1641_21#_c_1534_n 0.00614302f $X=9.645 $Y=1.29
+ $X2=0 $Y2=0
cc_918 N_A_1445_69#_c_1340_n N_A_1641_21#_c_1534_n 0.0182692f $X=9.48 $Y=1.26
+ $X2=0 $Y2=0
cc_919 N_A_1445_69#_c_1324_n N_A_1641_21#_c_1535_n 5.59345e-19 $X=9.375 $Y=1.125
+ $X2=0 $Y2=0
cc_920 N_A_1445_69#_c_1336_n N_A_1641_21#_c_1536_n 0.00756892f $X=11.81 $Y=0.73
+ $X2=0 $Y2=0
cc_921 N_A_1445_69#_c_1337_n N_A_1641_21#_c_1536_n 0.0128231f $X=10.045 $Y=0.73
+ $X2=0 $Y2=0
cc_922 N_A_1445_69#_c_1339_n N_A_1641_21#_c_1536_n 0.00173763f $X=9.645 $Y=1.29
+ $X2=0 $Y2=0
cc_923 N_A_1445_69#_c_1341_n N_A_1641_21#_c_1536_n 0.0046284f $X=9.96 $Y=1.26
+ $X2=0 $Y2=0
cc_924 N_A_1445_69#_M1014_g N_A_1641_21#_c_1613_n 0.00370709f $X=9.67 $Y=2.875
+ $X2=0 $Y2=0
cc_925 N_A_1445_69#_M1014_g N_A_1641_21#_c_1542_n 0.0173909f $X=9.67 $Y=2.875
+ $X2=0 $Y2=0
cc_926 N_A_1445_69#_c_1324_n N_A_1641_21#_c_1537_n 0.00144479f $X=9.375 $Y=1.125
+ $X2=0 $Y2=0
cc_927 N_A_1445_69#_c_1336_n N_A_1641_21#_c_1537_n 0.00270068f $X=11.81 $Y=0.73
+ $X2=0 $Y2=0
cc_928 N_A_1445_69#_c_1337_n N_A_1641_21#_c_1537_n 0.00429217f $X=10.045 $Y=0.73
+ $X2=0 $Y2=0
cc_929 N_A_1445_69#_c_1341_n N_A_1641_21#_c_1537_n 8.55445e-19 $X=9.96 $Y=1.26
+ $X2=0 $Y2=0
cc_930 N_A_1445_69#_c_1336_n N_CLK_M1007_g 0.0148232f $X=11.81 $Y=0.73 $X2=0
+ $Y2=0
cc_931 N_A_1445_69#_c_1338_n N_CLK_M1007_g 0.00295477f $X=11.895 $Y=0.985 $X2=0
+ $Y2=0
cc_932 N_A_1445_69#_M1003_g N_CLK_c_1645_n 0.00278229f $X=12.38 $Y=2.155 $X2=0
+ $Y2=0
cc_933 N_A_1445_69#_c_1336_n N_CLK_c_1645_n 0.00341726f $X=11.81 $Y=0.73 $X2=0
+ $Y2=0
cc_934 N_A_1445_69#_c_1342_n N_CLK_c_1645_n 0.00257508f $X=12.29 $Y=1.08 $X2=0
+ $Y2=0
cc_935 N_A_1445_69#_c_1343_n N_CLK_c_1645_n 0.0136709f $X=12.29 $Y=1.08 $X2=0
+ $Y2=0
cc_936 N_A_1445_69#_M1003_g N_CLK_c_1648_n 0.0023112f $X=12.38 $Y=2.155 $X2=0
+ $Y2=0
cc_937 N_A_1445_69#_c_1329_n N_CLK_c_1648_n 8.53337e-19 $X=12.29 $Y=1.585 $X2=0
+ $Y2=0
cc_938 N_A_1445_69#_c_1336_n N_CLK_c_1648_n 0.00539271f $X=11.81 $Y=0.73 $X2=0
+ $Y2=0
cc_939 N_A_1445_69#_c_1342_n N_CLK_c_1648_n 0.00850251f $X=12.29 $Y=1.08 $X2=0
+ $Y2=0
cc_940 N_A_1445_69#_M1039_g N_A_2408_367#_M1016_g 0.0242603f $X=12.455 $Y=0.445
+ $X2=0 $Y2=0
cc_941 N_A_1445_69#_c_1343_n N_A_2408_367#_M1016_g 0.00562601f $X=12.29 $Y=1.08
+ $X2=0 $Y2=0
cc_942 N_A_1445_69#_M1003_g N_A_2408_367#_M1024_g 0.0152106f $X=12.38 $Y=2.155
+ $X2=0 $Y2=0
cc_943 N_A_1445_69#_M1003_g N_A_2408_367#_c_1692_n 4.43964e-19 $X=12.38 $Y=2.155
+ $X2=0 $Y2=0
cc_944 N_A_1445_69#_M1039_g N_A_2408_367#_c_1699_n 0.00563611f $X=12.455
+ $Y=0.445 $X2=0 $Y2=0
cc_945 N_A_1445_69#_M1003_g N_A_2408_367#_c_1693_n 0.0160408f $X=12.38 $Y=2.155
+ $X2=0 $Y2=0
cc_946 N_A_1445_69#_c_1328_n N_A_2408_367#_c_1693_n 0.00197252f $X=12.327
+ $Y=1.065 $X2=0 $Y2=0
cc_947 N_A_1445_69#_c_1329_n N_A_2408_367#_c_1693_n 0.00128002f $X=12.29
+ $Y=1.585 $X2=0 $Y2=0
cc_948 N_A_1445_69#_c_1342_n N_A_2408_367#_c_1693_n 0.0140901f $X=12.29 $Y=1.08
+ $X2=0 $Y2=0
cc_949 N_A_1445_69#_c_1329_n N_A_2408_367#_c_1694_n 0.00399224f $X=12.29
+ $Y=1.585 $X2=0 $Y2=0
cc_950 N_A_1445_69#_c_1342_n N_A_2408_367#_c_1694_n 0.0143779f $X=12.29 $Y=1.08
+ $X2=0 $Y2=0
cc_951 N_A_1445_69#_M1039_g N_A_2408_367#_c_1687_n 0.0108423f $X=12.455 $Y=0.445
+ $X2=0 $Y2=0
cc_952 N_A_1445_69#_c_1342_n N_A_2408_367#_c_1687_n 0.0033701f $X=12.29 $Y=1.08
+ $X2=0 $Y2=0
cc_953 N_A_1445_69#_M1039_g N_A_2408_367#_c_1688_n 0.00396576f $X=12.455
+ $Y=0.445 $X2=0 $Y2=0
cc_954 N_A_1445_69#_c_1328_n N_A_2408_367#_c_1688_n 0.00669514f $X=12.327
+ $Y=1.065 $X2=0 $Y2=0
cc_955 N_A_1445_69#_c_1336_n N_A_2408_367#_c_1688_n 0.0159105f $X=11.81 $Y=0.73
+ $X2=0 $Y2=0
cc_956 N_A_1445_69#_c_1342_n N_A_2408_367#_c_1688_n 0.0201379f $X=12.29 $Y=1.08
+ $X2=0 $Y2=0
cc_957 N_A_1445_69#_M1003_g N_A_2408_367#_c_1689_n 8.8953e-19 $X=12.38 $Y=2.155
+ $X2=0 $Y2=0
cc_958 N_A_1445_69#_M1039_g N_A_2408_367#_c_1689_n 0.00487214f $X=12.455
+ $Y=0.445 $X2=0 $Y2=0
cc_959 N_A_1445_69#_c_1342_n N_A_2408_367#_c_1689_n 0.0338837f $X=12.29 $Y=1.08
+ $X2=0 $Y2=0
cc_960 N_A_1445_69#_c_1343_n N_A_2408_367#_c_1689_n 0.0031447f $X=12.29 $Y=1.08
+ $X2=0 $Y2=0
cc_961 N_A_1445_69#_c_1342_n N_A_2408_367#_c_1690_n 7.12795e-19 $X=12.29 $Y=1.08
+ $X2=0 $Y2=0
cc_962 N_A_1445_69#_c_1343_n N_A_2408_367#_c_1690_n 0.0209636f $X=12.29 $Y=1.08
+ $X2=0 $Y2=0
cc_963 N_A_1445_69#_M1014_g N_VPWR_c_1747_n 0.00539298f $X=9.67 $Y=2.875 $X2=0
+ $Y2=0
cc_964 N_A_1445_69#_M1014_g N_VPWR_c_1748_n 0.00343734f $X=9.67 $Y=2.875 $X2=0
+ $Y2=0
cc_965 N_A_1445_69#_M1003_g N_VPWR_c_1750_n 0.0159393f $X=12.38 $Y=2.155 $X2=0
+ $Y2=0
cc_966 N_A_1445_69#_M1003_g N_VPWR_c_1757_n 0.00259749f $X=12.38 $Y=2.155 $X2=0
+ $Y2=0
cc_967 N_A_1445_69#_M1017_d N_VPWR_c_1742_n 0.00289524f $X=7.27 $Y=1.895 $X2=0
+ $Y2=0
cc_968 N_A_1445_69#_M1014_g N_VPWR_c_1742_n 0.0111498f $X=9.67 $Y=2.875 $X2=0
+ $Y2=0
cc_969 N_A_1445_69#_M1003_g N_VPWR_c_1742_n 0.00344639f $X=12.38 $Y=2.155 $X2=0
+ $Y2=0
cc_970 N_A_1445_69#_M1014_g N_VPWR_c_1764_n 4.78216e-19 $X=9.67 $Y=2.875 $X2=0
+ $Y2=0
cc_971 N_A_1445_69#_c_1336_n N_VGND_M1010_d 0.0111351f $X=11.81 $Y=0.73 $X2=0
+ $Y2=0
cc_972 N_A_1445_69#_c_1363_n N_VGND_c_2008_n 0.0140087f $X=8.11 $Y=0.83 $X2=0
+ $Y2=0
cc_973 N_A_1445_69#_c_1333_n N_VGND_c_2008_n 0.00372063f $X=8.215 $Y=1.135 $X2=0
+ $Y2=0
cc_974 N_A_1445_69#_c_1340_n N_VGND_c_2008_n 0.0239502f $X=9.48 $Y=1.26 $X2=0
+ $Y2=0
cc_975 N_A_1445_69#_c_1336_n N_VGND_c_2009_n 0.0250071f $X=11.81 $Y=0.73 $X2=0
+ $Y2=0
cc_976 N_A_1445_69#_M1039_g N_VGND_c_2010_n 0.00436793f $X=12.455 $Y=0.445 $X2=0
+ $Y2=0
cc_977 N_A_1445_69#_c_1331_n N_VGND_c_2013_n 0.0123538f $X=7.365 $Y=0.49 $X2=0
+ $Y2=0
cc_978 N_A_1445_69#_c_1363_n N_VGND_c_2013_n 0.0025998f $X=8.11 $Y=0.83 $X2=0
+ $Y2=0
cc_979 N_A_1445_69#_c_1365_n N_VGND_c_2013_n 0.00907103f $X=7.53 $Y=0.83 $X2=0
+ $Y2=0
cc_980 N_A_1445_69#_c_1336_n N_VGND_c_2017_n 0.00931085f $X=11.81 $Y=0.73 $X2=0
+ $Y2=0
cc_981 N_A_1445_69#_M1039_g N_VGND_c_2018_n 0.00417265f $X=12.455 $Y=0.445 $X2=0
+ $Y2=0
cc_982 N_A_1445_69#_c_1336_n N_VGND_c_2018_n 0.0146939f $X=11.81 $Y=0.73 $X2=0
+ $Y2=0
cc_983 N_A_1445_69#_c_1324_n N_VGND_c_2020_n 7.82699e-19 $X=9.375 $Y=1.125 $X2=0
+ $Y2=0
cc_984 N_A_1445_69#_M1039_g N_VGND_c_2020_n 0.00740088f $X=12.455 $Y=0.445 $X2=0
+ $Y2=0
cc_985 N_A_1445_69#_c_1331_n N_VGND_c_2020_n 0.00952535f $X=7.365 $Y=0.49 $X2=0
+ $Y2=0
cc_986 N_A_1445_69#_c_1363_n N_VGND_c_2020_n 0.00522755f $X=8.11 $Y=0.83 $X2=0
+ $Y2=0
cc_987 N_A_1445_69#_c_1365_n N_VGND_c_2020_n 0.0190506f $X=7.53 $Y=0.83 $X2=0
+ $Y2=0
cc_988 N_A_1445_69#_c_1336_n N_VGND_c_2020_n 0.0427601f $X=11.81 $Y=0.73 $X2=0
+ $Y2=0
cc_989 N_A_1445_69#_c_1363_n A_1599_113# 0.00225709f $X=8.11 $Y=0.83 $X2=-0.19
+ $Y2=-0.245
cc_990 N_A_1445_69#_c_1333_n A_1599_113# 7.95246e-19 $X=8.215 $Y=1.135 $X2=-0.19
+ $Y2=-0.245
cc_991 N_A_1641_21#_c_1613_n N_VPWR_c_1747_n 0.0154118f $X=9.455 $Y=2.91 $X2=0
+ $Y2=0
cc_992 N_A_1641_21#_M1023_d N_VPWR_c_1742_n 0.00380103f $X=9.315 $Y=2.665 $X2=0
+ $Y2=0
cc_993 N_A_1641_21#_M1031_g N_VPWR_c_1742_n 0.00458965f $X=8.405 $Y=2.875 $X2=0
+ $Y2=0
cc_994 N_A_1641_21#_c_1613_n N_VPWR_c_1742_n 0.00978578f $X=9.455 $Y=2.91 $X2=0
+ $Y2=0
cc_995 N_A_1641_21#_M1031_g N_VPWR_c_1763_n 0.00352442f $X=8.405 $Y=2.875 $X2=0
+ $Y2=0
cc_996 N_A_1641_21#_M1031_g N_VPWR_c_1764_n 0.00877798f $X=8.405 $Y=2.875 $X2=0
+ $Y2=0
cc_997 N_A_1641_21#_M1020_g N_VGND_c_2008_n 0.0144241f $X=8.28 $Y=0.775 $X2=0
+ $Y2=0
cc_998 N_A_1641_21#_c_1529_n N_VGND_c_2008_n 0.0256764f $X=9.825 $Y=0.18 $X2=0
+ $Y2=0
cc_999 N_A_1641_21#_c_1531_n N_VGND_c_2008_n 0.00613368f $X=8.58 $Y=1.17 $X2=0
+ $Y2=0
cc_1000 N_A_1641_21#_c_1534_n N_VGND_c_2008_n 0.0139807f $X=9.59 $Y=0.8 $X2=0
+ $Y2=0
cc_1001 N_A_1641_21#_c_1535_n N_VGND_c_2008_n 0.00797755f $X=9.705 $Y=0.365
+ $X2=0 $Y2=0
cc_1002 N_A_1641_21#_c_1536_n N_VGND_c_2009_n 0.00506563f $X=9.99 $Y=0.35 $X2=0
+ $Y2=0
cc_1003 N_A_1641_21#_c_1537_n N_VGND_c_2009_n 0.0019451f $X=9.99 $Y=0.18 $X2=0
+ $Y2=0
cc_1004 N_A_1641_21#_c_1530_n N_VGND_c_2013_n 0.00980412f $X=8.355 $Y=0.18 $X2=0
+ $Y2=0
cc_1005 N_A_1641_21#_c_1529_n N_VGND_c_2017_n 0.0371052f $X=9.825 $Y=0.18 $X2=0
+ $Y2=0
cc_1006 N_A_1641_21#_c_1535_n N_VGND_c_2017_n 0.0191482f $X=9.705 $Y=0.365 $X2=0
+ $Y2=0
cc_1007 N_A_1641_21#_c_1536_n N_VGND_c_2017_n 0.0284865f $X=9.99 $Y=0.35 $X2=0
+ $Y2=0
cc_1008 N_A_1641_21#_c_1529_n N_VGND_c_2020_n 0.0439255f $X=9.825 $Y=0.18 $X2=0
+ $Y2=0
cc_1009 N_A_1641_21#_c_1530_n N_VGND_c_2020_n 0.00801046f $X=8.355 $Y=0.18 $X2=0
+ $Y2=0
cc_1010 N_A_1641_21#_c_1535_n N_VGND_c_2020_n 0.00961688f $X=9.705 $Y=0.365
+ $X2=0 $Y2=0
cc_1011 N_A_1641_21#_c_1536_n N_VGND_c_2020_n 0.0149973f $X=9.99 $Y=0.35 $X2=0
+ $Y2=0
cc_1012 N_A_1641_21#_c_1537_n N_VGND_c_2020_n 0.0100269f $X=9.99 $Y=0.18 $X2=0
+ $Y2=0
cc_1013 N_CLK_c_1648_n N_A_2408_367#_c_1692_n 0.0514176f $X=11.715 $Y=1.51 $X2=0
+ $Y2=0
cc_1014 N_CLK_c_1648_n N_A_2408_367#_c_1694_n 0.0150205f $X=11.715 $Y=1.51 $X2=0
+ $Y2=0
cc_1015 N_CLK_M1018_g N_VPWR_c_1749_n 0.00841898f $X=11.25 $Y=2.465 $X2=0 $Y2=0
cc_1016 N_CLK_M1018_g N_VPWR_c_1757_n 0.00431225f $X=11.25 $Y=2.465 $X2=0 $Y2=0
cc_1017 N_CLK_M1018_g N_VPWR_c_1742_n 0.00751203f $X=11.25 $Y=2.465 $X2=0 $Y2=0
cc_1018 N_CLK_c_1648_n N_VPWR_c_1742_n 0.0100517f $X=11.715 $Y=1.51 $X2=0 $Y2=0
cc_1019 N_CLK_M1007_g N_VGND_c_2009_n 0.00670283f $X=11.25 $Y=0.785 $X2=0 $Y2=0
cc_1020 N_CLK_M1007_g N_VGND_c_2018_n 0.00330473f $X=11.25 $Y=0.785 $X2=0 $Y2=0
cc_1021 N_CLK_M1007_g N_VGND_c_2020_n 0.0043803f $X=11.25 $Y=0.785 $X2=0 $Y2=0
cc_1022 N_A_2408_367#_c_1693_n N_VPWR_M1003_d 0.00351427f $X=12.665 $Y=1.76
+ $X2=0 $Y2=0
cc_1023 N_A_2408_367#_M1024_g N_VPWR_c_1750_n 0.0244185f $X=12.965 $Y=2.465
+ $X2=0 $Y2=0
cc_1024 N_A_2408_367#_c_1692_n N_VPWR_c_1750_n 0.0198415f $X=12.165 $Y=1.98
+ $X2=0 $Y2=0
cc_1025 N_A_2408_367#_c_1693_n N_VPWR_c_1750_n 0.0313762f $X=12.665 $Y=1.76
+ $X2=0 $Y2=0
cc_1026 N_A_2408_367#_c_1690_n N_VPWR_c_1750_n 9.80275e-19 $X=12.83 $Y=1.47
+ $X2=0 $Y2=0
cc_1027 N_A_2408_367#_M1024_g N_VPWR_c_1758_n 0.00486043f $X=12.965 $Y=2.465
+ $X2=0 $Y2=0
cc_1028 N_A_2408_367#_M1024_g N_VPWR_c_1742_n 0.00917987f $X=12.965 $Y=2.465
+ $X2=0 $Y2=0
cc_1029 N_A_2408_367#_c_1692_n N_VPWR_c_1742_n 0.00823744f $X=12.165 $Y=1.98
+ $X2=0 $Y2=0
cc_1030 N_A_2408_367#_M1016_g N_Q_c_1994_n 0.0237858f $X=12.965 $Y=0.655 $X2=0
+ $Y2=0
cc_1031 N_A_2408_367#_c_1693_n N_Q_c_1994_n 0.0136053f $X=12.665 $Y=1.76 $X2=0
+ $Y2=0
cc_1032 N_A_2408_367#_c_1689_n N_Q_c_1994_n 0.0549572f $X=12.83 $Y=1.47 $X2=0
+ $Y2=0
cc_1033 N_A_2408_367#_c_1687_n N_VGND_M1039_d 0.00349403f $X=12.665 $Y=0.73
+ $X2=0 $Y2=0
cc_1034 N_A_2408_367#_c_1689_n N_VGND_M1039_d 0.00302927f $X=12.83 $Y=1.47 $X2=0
+ $Y2=0
cc_1035 N_A_2408_367#_M1016_g N_VGND_c_2010_n 0.00815466f $X=12.965 $Y=0.655
+ $X2=0 $Y2=0
cc_1036 N_A_2408_367#_c_1687_n N_VGND_c_2010_n 0.0219838f $X=12.665 $Y=0.73
+ $X2=0 $Y2=0
cc_1037 N_A_2408_367#_c_1699_n N_VGND_c_2018_n 0.0137411f $X=12.24 $Y=0.44 $X2=0
+ $Y2=0
cc_1038 N_A_2408_367#_c_1687_n N_VGND_c_2018_n 0.00240763f $X=12.665 $Y=0.73
+ $X2=0 $Y2=0
cc_1039 N_A_2408_367#_M1016_g N_VGND_c_2019_n 0.00486043f $X=12.965 $Y=0.655
+ $X2=0 $Y2=0
cc_1040 N_A_2408_367#_M1039_s N_VGND_c_2020_n 0.00340962f $X=12.115 $Y=0.235
+ $X2=0 $Y2=0
cc_1041 N_A_2408_367#_M1016_g N_VGND_c_2020_n 0.00917987f $X=12.965 $Y=0.655
+ $X2=0 $Y2=0
cc_1042 N_A_2408_367#_c_1699_n N_VGND_c_2020_n 0.00949595f $X=12.24 $Y=0.44
+ $X2=0 $Y2=0
cc_1043 N_A_2408_367#_c_1687_n N_VGND_c_2020_n 0.00580796f $X=12.665 $Y=0.73
+ $X2=0 $Y2=0
cc_1044 N_VPWR_M1008_d N_A_380_50#_c_1899_n 0.00446845f $X=3.035 $Y=2.315 $X2=0
+ $Y2=0
cc_1045 N_VPWR_c_1744_n N_A_380_50#_c_1899_n 0.0175938f $X=3.205 $Y=2.77 $X2=0
+ $Y2=0
cc_1046 N_VPWR_c_1742_n N_A_380_50#_c_1899_n 0.0227422f $X=13.2 $Y=3.33 $X2=0
+ $Y2=0
cc_1047 N_VPWR_c_1743_n N_A_380_50#_c_1897_n 0.0230792f $X=1.485 $Y=2.46 $X2=0
+ $Y2=0
cc_1048 N_VPWR_c_1744_n N_A_380_50#_c_1897_n 0.00515726f $X=3.205 $Y=2.77 $X2=0
+ $Y2=0
cc_1049 N_VPWR_c_1753_n N_A_380_50#_c_1897_n 0.0154243f $X=3.04 $Y=3.33 $X2=0
+ $Y2=0
cc_1050 N_VPWR_c_1742_n N_A_380_50#_c_1897_n 0.0119923f $X=13.2 $Y=3.33 $X2=0
+ $Y2=0
cc_1051 N_VPWR_c_1744_n N_A_380_50#_c_1898_n 0.0132219f $X=3.205 $Y=2.77 $X2=0
+ $Y2=0
cc_1052 N_VPWR_c_1754_n N_A_380_50#_c_1898_n 0.0119038f $X=4.865 $Y=3.33 $X2=0
+ $Y2=0
cc_1053 N_VPWR_c_1742_n N_A_380_50#_c_1898_n 0.0123859f $X=13.2 $Y=3.33 $X2=0
+ $Y2=0
cc_1054 N_VPWR_c_1742_n A_1578_533# 0.00373269f $X=13.2 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_1055 N_VPWR_c_1742_n N_Q_M1024_d 0.00371702f $X=13.2 $Y=3.33 $X2=0 $Y2=0
cc_1056 N_VPWR_c_1758_n N_Q_c_1994_n 0.018528f $X=13.2 $Y=3.33 $X2=0 $Y2=0
cc_1057 N_VPWR_c_1742_n N_Q_c_1994_n 0.0104192f $X=13.2 $Y=3.33 $X2=0 $Y2=0
cc_1058 N_A_380_50#_c_1899_n A_513_463# 0.0104694f $X=3.48 $Y=2.4 $X2=-0.19
+ $Y2=-0.245
cc_1059 N_A_380_50#_c_1892_n N_VGND_M1027_d 2.89266e-19 $X=3.48 $Y=0.9 $X2=0
+ $Y2=0
cc_1060 N_A_380_50#_c_1949_n N_VGND_M1027_d 0.00207681f $X=3.582 $Y=0.9 $X2=0
+ $Y2=0
cc_1061 N_A_380_50#_c_1892_n N_VGND_c_2006_n 0.0020984f $X=3.48 $Y=0.9 $X2=0
+ $Y2=0
cc_1062 N_A_380_50#_c_1894_n N_VGND_c_2006_n 0.00381712f $X=4.015 $Y=0.9 $X2=0
+ $Y2=0
cc_1063 N_A_380_50#_c_1949_n N_VGND_c_2006_n 0.0172277f $X=3.582 $Y=0.9 $X2=0
+ $Y2=0
cc_1064 N_A_380_50#_c_1936_n N_VGND_c_2011_n 0.00347046f $X=4.13 $Y=0.82 $X2=0
+ $Y2=0
cc_1065 N_A_380_50#_c_1892_n N_VGND_c_2020_n 0.00764367f $X=3.48 $Y=0.9 $X2=0
+ $Y2=0
cc_1066 N_A_380_50#_c_1894_n N_VGND_c_2020_n 0.00847965f $X=4.015 $Y=0.9 $X2=0
+ $Y2=0
cc_1067 N_A_380_50#_c_1949_n N_VGND_c_2020_n 7.96362e-19 $X=3.582 $Y=0.9 $X2=0
+ $Y2=0
cc_1068 N_A_380_50#_c_1936_n N_VGND_c_2020_n 0.00495356f $X=4.13 $Y=0.82 $X2=0
+ $Y2=0
cc_1069 N_A_380_50#_c_1892_n N_noxref_24_M1000_d 0.00226056f $X=3.48 $Y=0.9
+ $X2=0 $Y2=0
cc_1070 N_A_380_50#_M1033_d N_noxref_24_c_2144_n 0.00996163f $X=1.9 $Y=0.25
+ $X2=0 $Y2=0
cc_1071 N_A_380_50#_c_1892_n N_noxref_24_c_2144_n 0.0129281f $X=3.48 $Y=0.9
+ $X2=0 $Y2=0
cc_1072 N_A_380_50#_c_1895_n N_noxref_24_c_2144_n 0.0227549f $X=2.155 $Y=0.7
+ $X2=0 $Y2=0
cc_1073 N_A_380_50#_c_1892_n N_noxref_24_c_2145_n 0.0167737f $X=3.48 $Y=0.9
+ $X2=0 $Y2=0
cc_1074 N_A_380_50#_c_1895_n N_noxref_24_c_2145_n 5.95629e-19 $X=2.155 $Y=0.7
+ $X2=0 $Y2=0
cc_1075 N_A_380_50#_c_1892_n noxref_26 0.00145645f $X=3.48 $Y=0.9 $X2=-0.19
+ $Y2=-0.245
cc_1076 N_Q_c_1994_n N_VGND_c_2019_n 0.018528f $X=13.18 $Y=0.42 $X2=0 $Y2=0
cc_1077 N_Q_M1016_d N_VGND_c_2020_n 0.00371702f $X=13.04 $Y=0.235 $X2=0 $Y2=0
cc_1078 N_Q_c_1994_n N_VGND_c_2020_n 0.0104192f $X=13.18 $Y=0.42 $X2=0 $Y2=0
cc_1079 N_VGND_c_2016_n N_noxref_24_c_2144_n 0.0864158f $X=3.405 $Y=0 $X2=0
+ $Y2=0
cc_1080 N_VGND_c_2020_n N_noxref_24_c_2144_n 0.0561734f $X=13.2 $Y=0 $X2=0 $Y2=0
cc_1081 N_VGND_c_2005_n N_noxref_24_c_2148_n 0.0196347f $X=0.73 $Y=0.525 $X2=0
+ $Y2=0
cc_1082 N_VGND_c_2016_n N_noxref_24_c_2148_n 0.0124385f $X=3.405 $Y=0 $X2=0
+ $Y2=0
cc_1083 N_VGND_c_2020_n N_noxref_24_c_2148_n 0.00789949f $X=13.2 $Y=0 $X2=0
+ $Y2=0
cc_1084 N_VGND_c_2006_n N_noxref_24_c_2145_n 0.0111082f $X=3.57 $Y=0.55 $X2=0
+ $Y2=0
cc_1085 N_VGND_c_2016_n N_noxref_24_c_2145_n 0.0211423f $X=3.405 $Y=0 $X2=0
+ $Y2=0
cc_1086 N_VGND_c_2020_n N_noxref_24_c_2145_n 0.0124918f $X=13.2 $Y=0 $X2=0 $Y2=0
cc_1087 N_noxref_24_c_2144_n noxref_25 0.00458445f $X=2.895 $Y=0.35 $X2=-0.19
+ $Y2=-0.245
cc_1088 N_noxref_24_c_2144_n noxref_26 0.0014993f $X=2.895 $Y=0.35 $X2=-0.19
+ $Y2=-0.245
