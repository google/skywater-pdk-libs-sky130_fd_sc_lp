* NGSPICE file created from sky130_fd_sc_lp__dfxbp_lp.ext - technology: sky130A

.subckt sky130_fd_sc_lp__dfxbp_lp CLK D VGND VNB VPB VPWR Q Q_N
M1000 a_297_85# D VGND VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=8.391e+11p ps=9.11e+06u
M1001 Q_N a_2062_367# VPWR VPB phighvt w=1e+06u l=250000u
+  ad=2.85e+11p pd=2.57e+06u as=1.99e+12p ps=1.598e+07u
M1002 a_239_403# D a_297_85# VNB nshort w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=0p ps=0u
M1003 a_2168_127# a_1507_321# VGND VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1004 VPWR a_615_93# a_349_323# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=5.6e+11p ps=5.12e+06u
M1005 a_1445_419# a_511_218# a_1339_153# VPB phighvt w=1e+06u l=250000u
+  ad=3.1e+11p pd=2.62e+06u as=2.8e+11p ps=2.56e+06u
M1006 VGND CLK a_125_85# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1007 VPWR a_1507_321# Q VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=2.85e+11p ps=2.57e+06u
M1008 a_239_403# a_511_218# a_455_85# VPB phighvt w=1e+06u l=250000u
+  ad=5.65e+11p pd=5.13e+06u as=2.8e+11p ps=2.56e+06u
M1009 VGND a_27_403# a_1049_125# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1010 VGND a_1507_321# a_1232_153# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=2.814e+11p ps=3.02e+06u
M1011 a_2010_127# a_1507_321# Q VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=1.176e+11p ps=1.4e+06u
M1012 a_2062_367# a_1507_321# a_2168_127# VNB nshort w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=0p ps=0u
M1013 VPWR CLK a_27_403# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=2.8e+11p ps=2.56e+06u
M1014 a_2062_367# a_1507_321# VPWR VPB phighvt w=1e+06u l=250000u
+  ad=2.85e+11p pd=2.57e+06u as=0p ps=0u
M1015 a_1507_321# a_1339_153# a_1742_57# VNB nshort w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=8.82e+10p ps=1.26e+06u
M1016 a_455_85# a_27_403# a_239_403# VNB nshort w=420000u l=150000u
+  ad=2.341e+11p pd=2.06e+06u as=0p ps=0u
M1017 VGND a_1507_321# a_2010_127# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_125_85# CLK a_27_403# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1019 VGND a_615_93# a_573_119# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1020 a_615_93# a_455_85# a_763_119# VNB nshort w=420000u l=150000u
+  ad=2.373e+11p pd=2.81e+06u as=8.82e+10p ps=1.26e+06u
M1021 VPWR a_1507_321# a_1445_419# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_1339_153# a_27_403# a_1232_153# VNB nshort w=420000u l=150000u
+  ad=1.9665e+11p pd=1.92e+06u as=0p ps=0u
M1023 a_1339_153# a_27_403# a_615_93# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=5.7e+11p ps=5.14e+06u
M1024 a_1742_57# a_1339_153# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 Q_N a_2062_367# a_2436_57# VNB nshort w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=8.82e+10p ps=1.26e+06u
M1026 a_455_85# a_27_403# a_349_323# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_615_93# a_455_85# VPWR VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_239_403# D VPWR VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1029 a_573_119# a_511_218# a_455_85# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 a_763_119# a_455_85# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_615_93# a_511_218# a_1339_153# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 a_2436_57# a_2062_367# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 VPWR a_27_403# a_511_218# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=2.85e+11p ps=2.57e+06u
M1034 a_1049_125# a_27_403# a_511_218# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.736e+11p ps=1.71e+06u
M1035 a_1507_321# a_1339_153# VPWR VPB phighvt w=1e+06u l=250000u
+  ad=2.85e+11p pd=2.57e+06u as=0p ps=0u
.ends

