* File: sky130_fd_sc_lp__ha_4.pex.spice
* Created: Fri Aug 28 10:36:35 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__HA_4%A_110_263# 1 2 3 4 15 19 23 27 31 35 39 43 45
+ 53 56 60 61 62 64 65 69 77 78 79 81 82 83 86 89 102 107
c239 102 0 1.0594e-19 $X=1.95 $Y=1.48
c240 81 0 2.95893e-20 $X=9.425 $Y=1.84
c241 56 0 3.13091e-20 $X=6.82 $Y=2.355
r242 101 102 6.12014 $w=3.3e-07 $l=3.5e-08 $layer=POLY_cond $X=1.915 $Y=1.48
+ $X2=1.95 $Y2=1.48
r243 98 99 6.12014 $w=3.3e-07 $l=3.5e-08 $layer=POLY_cond $X=1.485 $Y=1.48
+ $X2=1.52 $Y2=1.48
r244 97 98 69.0702 $w=3.3e-07 $l=3.95e-07 $layer=POLY_cond $X=1.09 $Y=1.48
+ $X2=1.485 $Y2=1.48
r245 96 97 6.12014 $w=3.3e-07 $l=3.5e-08 $layer=POLY_cond $X=1.055 $Y=1.48
+ $X2=1.09 $Y2=1.48
r246 92 94 6.12014 $w=3.3e-07 $l=3.5e-08 $layer=POLY_cond $X=0.625 $Y=1.48
+ $X2=0.66 $Y2=1.48
r247 90 110 10.7517 $w=4.73e-07 $l=2.2e-07 $layer=LI1_cond $X=9.272 $Y=0.925
+ $X2=9.272 $Y2=1.145
r248 90 107 5.66563 $w=4.73e-07 $l=2.25e-07 $layer=LI1_cond $X=9.272 $Y=0.925
+ $X2=9.272 $Y2=0.7
r249 89 90 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=0.925
+ $X2=9.36 $Y2=0.925
r250 85 86 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0.925
+ $X2=2.16 $Y2=0.925
r251 83 85 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.305 $Y=0.925
+ $X2=2.16 $Y2=0.925
r252 82 89 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=9.215 $Y=0.925
+ $X2=9.36 $Y2=0.925
r253 82 83 8.55196 $w=1.4e-07 $l=6.91e-06 $layer=MET1_cond $X=9.215 $Y=0.925
+ $X2=2.305 $Y2=0.925
r254 77 79 26.1869 $w=1.78e-07 $l=4.25e-07 $layer=LI1_cond $X=8.615 $Y=2.36
+ $X2=9.04 $Y2=2.36
r255 77 78 10.2135 $w=1.78e-07 $l=1.65e-07 $layer=LI1_cond $X=8.615 $Y=2.36
+ $X2=8.45 $Y2=2.36
r256 73 86 30.6631 $w=1.68e-07 $l=4.7e-07 $layer=LI1_cond $X=2.16 $Y=1.395
+ $X2=2.16 $Y2=0.925
r257 69 71 36.3313 $w=2.93e-07 $l=9.3e-07 $layer=LI1_cond $X=9.837 $Y=1.98
+ $X2=9.837 $Y2=2.91
r258 67 69 2.14862 $w=2.93e-07 $l=5.5e-08 $layer=LI1_cond $X=9.837 $Y=1.925
+ $X2=9.837 $Y2=1.98
r259 66 81 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.51 $Y=1.84
+ $X2=9.425 $Y2=1.84
r260 65 67 7.47753 $w=1.7e-07 $l=1.84673e-07 $layer=LI1_cond $X=9.69 $Y=1.84
+ $X2=9.837 $Y2=1.925
r261 65 66 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=9.69 $Y=1.84
+ $X2=9.51 $Y2=1.84
r262 64 81 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.425 $Y=1.755
+ $X2=9.425 $Y2=1.84
r263 64 110 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=9.425 $Y=1.755
+ $X2=9.425 $Y2=1.145
r264 61 81 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.34 $Y=1.84
+ $X2=9.425 $Y2=1.84
r265 61 62 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=9.34 $Y=1.84
+ $X2=9.125 $Y2=1.84
r266 60 79 1.06262 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=9.04 $Y=2.27 $X2=9.04
+ $Y2=2.36
r267 59 62 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.04 $Y=1.925
+ $X2=9.125 $Y2=1.84
r268 59 60 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=9.04 $Y=1.925
+ $X2=9.04 $Y2=2.27
r269 56 78 106.342 $w=1.68e-07 $l=1.63e-06 $layer=LI1_cond $X=6.82 $Y=2.355
+ $X2=8.45 $Y2=2.355
r270 53 56 17.9729 $w=2.18e-07 $l=3.39588e-07 $layer=LI1_cond $X=6.51 $Y=2.417
+ $X2=6.82 $Y2=2.355
r271 52 101 9.61737 $w=3.3e-07 $l=5.5e-08 $layer=POLY_cond $X=1.86 $Y=1.48
+ $X2=1.915 $Y2=1.48
r272 52 99 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.86 $Y=1.48
+ $X2=1.52 $Y2=1.48
r273 51 52 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.86
+ $Y=1.48 $X2=1.86 $Y2=1.48
r274 48 96 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=0.84 $Y=1.48
+ $X2=1.055 $Y2=1.48
r275 48 94 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=0.84 $Y=1.48
+ $X2=0.66 $Y2=1.48
r276 47 51 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=0.84 $Y=1.48
+ $X2=1.86 $Y2=1.48
r277 47 48 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.84
+ $Y=1.48 $X2=0.84 $Y2=1.48
r278 45 73 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.075 $Y=1.48
+ $X2=2.16 $Y2=1.395
r279 45 51 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=2.075 $Y=1.48
+ $X2=1.86 $Y2=1.48
r280 41 102 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.95 $Y=1.315
+ $X2=1.95 $Y2=1.48
r281 41 43 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.95 $Y=1.315
+ $X2=1.95 $Y2=0.655
r282 37 101 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.915 $Y=1.645
+ $X2=1.915 $Y2=1.48
r283 37 39 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=1.915 $Y=1.645
+ $X2=1.915 $Y2=2.465
r284 33 99 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.52 $Y=1.315
+ $X2=1.52 $Y2=1.48
r285 33 35 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.52 $Y=1.315
+ $X2=1.52 $Y2=0.655
r286 29 98 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.485 $Y=1.645
+ $X2=1.485 $Y2=1.48
r287 29 31 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=1.485 $Y=1.645
+ $X2=1.485 $Y2=2.465
r288 25 97 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.09 $Y=1.315
+ $X2=1.09 $Y2=1.48
r289 25 27 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.09 $Y=1.315
+ $X2=1.09 $Y2=0.655
r290 21 96 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.055 $Y=1.645
+ $X2=1.055 $Y2=1.48
r291 21 23 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=1.055 $Y=1.645
+ $X2=1.055 $Y2=2.465
r292 17 94 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.66 $Y=1.315
+ $X2=0.66 $Y2=1.48
r293 17 19 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.66 $Y=1.315
+ $X2=0.66 $Y2=0.655
r294 13 92 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.625 $Y=1.645
+ $X2=0.625 $Y2=1.48
r295 13 15 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=0.625 $Y=1.645
+ $X2=0.625 $Y2=2.465
r296 4 71 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=9.68
+ $Y=1.835 $X2=9.82 $Y2=2.91
r297 4 69 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=9.68
+ $Y=1.835 $X2=9.82 $Y2=1.98
r298 3 77 300 $w=1.7e-07 $l=6.71044e-07 $layer=licon1_PDIFF $count=2 $X=8.395
+ $Y=1.835 $X2=8.615 $Y2=2.405
r299 2 53 300 $w=1.7e-07 $l=7.85016e-07 $layer=licon1_PDIFF $count=2 $X=6.42
+ $Y=1.835 $X2=6.545 $Y2=2.56
r300 1 107 91 $w=1.7e-07 $l=4.3946e-07 $layer=licon1_NDIFF $count=2 $X=9.06
+ $Y=0.325 $X2=9.2 $Y2=0.7
.ends

.subckt PM_SKY130_FD_SC_LP__HA_4%A_454_263# 1 2 3 12 16 22 26 30 34 38 42 46 50
+ 52 56 60 62 64 66 75 77 78 79 80 81 82 84 86 90 94 96 98 101 102 104 107 113
+ 114 119 126 128
c267 126 0 1.60386e-19 $X=3.67 $Y=1.48
c268 86 0 1.61867e-19 $X=5.18 $Y=2.13
c269 75 0 2.54181e-20 $X=3.805 $Y=1.395
r270 128 129 30.474 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=9.005 $Y=1.4
+ $X2=9.005 $Y2=1.325
r271 125 126 6.12014 $w=3.3e-07 $l=3.5e-08 $layer=POLY_cond $X=3.635 $Y=1.48
+ $X2=3.67 $Y2=1.48
r272 122 123 6.12014 $w=3.3e-07 $l=3.5e-08 $layer=POLY_cond $X=3.205 $Y=1.48
+ $X2=3.24 $Y2=1.48
r273 118 120 6.12014 $w=3.3e-07 $l=3.5e-08 $layer=POLY_cond $X=2.775 $Y=1.48
+ $X2=2.81 $Y2=1.48
r274 118 119 30.474 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=2.775 $Y=1.48
+ $X2=2.7 $Y2=1.48
r275 114 116 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=6.385 $Y=2.015
+ $X2=6.385 $Y2=2.13
r276 109 111 4.10084 $w=2.38e-07 $l=8e-08 $layer=LI1_cond $X=4.352 $Y=2.13
+ $X2=4.352 $Y2=2.21
r277 108 109 9.7395 $w=2.38e-07 $l=1.9e-07 $layer=LI1_cond $X=4.352 $Y=1.94
+ $X2=4.352 $Y2=2.13
r278 105 131 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=9.005 $Y=1.49
+ $X2=9.005 $Y2=1.655
r279 105 128 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=9.005 $Y=1.49
+ $X2=9.005 $Y2=1.4
r280 104 105 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.005
+ $Y=1.49 $X2=9.005 $Y2=1.49
r281 102 104 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=8.775 $Y=1.49
+ $X2=9.005 $Y2=1.49
r282 100 102 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.69 $Y=1.575
+ $X2=8.775 $Y2=1.49
r283 100 101 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=8.69 $Y=1.575
+ $X2=8.69 $Y2=1.93
r284 99 114 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.47 $Y=2.015
+ $X2=6.385 $Y2=2.015
r285 98 101 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.605 $Y=2.015
+ $X2=8.69 $Y2=1.93
r286 98 99 139.289 $w=1.68e-07 $l=2.135e-06 $layer=LI1_cond $X=8.605 $Y=2.015
+ $X2=6.47 $Y2=2.015
r287 97 113 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=5.39 $Y=2.13
+ $X2=5.285 $Y2=2.13
r288 96 116 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.3 $Y=2.13
+ $X2=6.385 $Y2=2.13
r289 96 97 59.369 $w=1.68e-07 $l=9.1e-07 $layer=LI1_cond $X=6.3 $Y=2.13 $X2=5.39
+ $Y2=2.13
r290 92 113 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=5.285 $Y=2.215
+ $X2=5.285 $Y2=2.13
r291 92 94 36.7056 $w=2.08e-07 $l=6.95e-07 $layer=LI1_cond $X=5.285 $Y=2.215
+ $X2=5.285 $Y2=2.91
r292 88 90 13.134 $w=1.88e-07 $l=2.25e-07 $layer=LI1_cond $X=4.825 $Y=0.995
+ $X2=4.825 $Y2=0.77
r293 87 109 2.70854 $w=1.7e-07 $l=1.58e-07 $layer=LI1_cond $X=4.51 $Y=2.13
+ $X2=4.352 $Y2=2.13
r294 86 113 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=5.18 $Y=2.13
+ $X2=5.285 $Y2=2.13
r295 86 87 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.18 $Y=2.13
+ $X2=4.51 $Y2=2.13
r296 82 111 0.951208 $w=3.15e-07 $l=5e-09 $layer=LI1_cond $X=4.352 $Y=2.215
+ $X2=4.352 $Y2=2.21
r297 82 84 24.6952 $w=3.13e-07 $l=6.75e-07 $layer=LI1_cond $X=4.352 $Y=2.215
+ $X2=4.352 $Y2=2.89
r298 80 108 2.70854 $w=1.7e-07 $l=1.57e-07 $layer=LI1_cond $X=4.195 $Y=1.94
+ $X2=4.352 $Y2=1.94
r299 80 81 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=4.195 $Y=1.94
+ $X2=3.89 $Y2=1.94
r300 78 88 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=4.73 $Y=1.08
+ $X2=4.825 $Y2=0.995
r301 78 79 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=4.73 $Y=1.08
+ $X2=3.89 $Y2=1.08
r302 77 81 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.805 $Y=1.855
+ $X2=3.89 $Y2=1.94
r303 76 107 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.805 $Y=1.565
+ $X2=3.805 $Y2=1.48
r304 76 77 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=3.805 $Y=1.565
+ $X2=3.805 $Y2=1.855
r305 75 107 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.805 $Y=1.395
+ $X2=3.805 $Y2=1.48
r306 74 79 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.805 $Y=1.165
+ $X2=3.89 $Y2=1.08
r307 74 75 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=3.805 $Y=1.165
+ $X2=3.805 $Y2=1.395
r308 73 125 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=3.62 $Y=1.48
+ $X2=3.635 $Y2=1.48
r309 73 123 66.4473 $w=3.3e-07 $l=3.8e-07 $layer=POLY_cond $X=3.62 $Y=1.48
+ $X2=3.24 $Y2=1.48
r310 72 73 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=3.62
+ $Y=1.48 $X2=3.62 $Y2=1.48
r311 69 122 46.3382 $w=3.3e-07 $l=2.65e-07 $layer=POLY_cond $X=2.94 $Y=1.48
+ $X2=3.205 $Y2=1.48
r312 69 120 22.732 $w=3.3e-07 $l=1.3e-07 $layer=POLY_cond $X=2.94 $Y=1.48
+ $X2=2.81 $Y2=1.48
r313 68 72 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=2.94 $Y=1.48
+ $X2=3.62 $Y2=1.48
r314 68 69 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.94
+ $Y=1.48 $X2=2.94 $Y2=1.48
r315 66 107 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.72 $Y=1.48
+ $X2=3.805 $Y2=1.48
r316 66 72 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=3.72 $Y=1.48 $X2=3.62
+ $Y2=1.48
r317 63 64 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=9.415 $Y=1.4
+ $X2=9.605 $Y2=1.4
r318 58 64 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.605 $Y=1.475
+ $X2=9.605 $Y2=1.4
r319 58 60 507.638 $w=1.5e-07 $l=9.9e-07 $layer=POLY_cond $X=9.605 $Y=1.475
+ $X2=9.605 $Y2=2.465
r320 54 63 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.415 $Y=1.325
+ $X2=9.415 $Y2=1.4
r321 54 56 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=9.415 $Y=1.325
+ $X2=9.415 $Y2=0.745
r322 53 128 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.17 $Y=1.4
+ $X2=9.005 $Y2=1.4
r323 52 63 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.34 $Y=1.4
+ $X2=9.415 $Y2=1.4
r324 52 53 87.1702 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=9.34 $Y=1.4
+ $X2=9.17 $Y2=1.4
r325 50 129 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=8.985 $Y=0.745
+ $X2=8.985 $Y2=1.325
r326 46 131 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=8.915 $Y=2.465
+ $X2=8.915 $Y2=1.655
r327 40 126 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.67 $Y=1.315
+ $X2=3.67 $Y2=1.48
r328 40 42 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.67 $Y=1.315
+ $X2=3.67 $Y2=0.655
r329 36 125 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.635 $Y=1.645
+ $X2=3.635 $Y2=1.48
r330 36 38 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=3.635 $Y=1.645
+ $X2=3.635 $Y2=2.465
r331 32 123 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.24 $Y=1.315
+ $X2=3.24 $Y2=1.48
r332 32 34 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.24 $Y=1.315
+ $X2=3.24 $Y2=0.655
r333 28 122 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.205 $Y=1.645
+ $X2=3.205 $Y2=1.48
r334 28 30 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=3.205 $Y=1.645
+ $X2=3.205 $Y2=2.465
r335 24 120 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.81 $Y=1.315
+ $X2=2.81 $Y2=1.48
r336 24 26 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.81 $Y=1.315
+ $X2=2.81 $Y2=0.655
r337 20 118 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.775 $Y=1.645
+ $X2=2.775 $Y2=1.48
r338 20 22 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=2.775 $Y=1.645
+ $X2=2.775 $Y2=2.465
r339 19 62 5.30422 $w=1.5e-07 $l=9.3e-08 $layer=POLY_cond $X=2.455 $Y=1.39
+ $X2=2.362 $Y2=1.39
r340 19 119 125.628 $w=1.5e-07 $l=2.45e-07 $layer=POLY_cond $X=2.455 $Y=1.39
+ $X2=2.7 $Y2=1.39
r341 14 62 20.4101 $w=1.5e-07 $l=8.35165e-08 $layer=POLY_cond $X=2.38 $Y=1.315
+ $X2=2.362 $Y2=1.39
r342 14 16 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.38 $Y=1.315
+ $X2=2.38 $Y2=0.655
r343 10 62 20.4101 $w=1.5e-07 $l=8.30662e-08 $layer=POLY_cond $X=2.345 $Y=1.465
+ $X2=2.362 $Y2=1.39
r344 10 12 512.766 $w=1.5e-07 $l=1e-06 $layer=POLY_cond $X=2.345 $Y=1.465
+ $X2=2.345 $Y2=2.465
r345 3 113 400 $w=1.7e-07 $l=4.3946e-07 $layer=licon1_PDIFF $count=1 $X=5.155
+ $Y=1.835 $X2=5.295 $Y2=2.21
r346 3 94 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=5.155
+ $Y=1.835 $X2=5.295 $Y2=2.91
r347 2 111 400 $w=1.7e-07 $l=4.3946e-07 $layer=licon1_PDIFF $count=1 $X=4.255
+ $Y=1.835 $X2=4.395 $Y2=2.21
r348 2 84 400 $w=1.7e-07 $l=1.12282e-06 $layer=licon1_PDIFF $count=1 $X=4.255
+ $Y=1.835 $X2=4.395 $Y2=2.89
r349 1 90 182 $w=1.7e-07 $l=6.00937e-07 $layer=licon1_NDIFF $count=1 $X=4.685
+ $Y=0.235 $X2=4.825 $Y2=0.77
.ends

.subckt PM_SKY130_FD_SC_LP__HA_4%A 3 7 11 15 19 23 27 31 33 36 38 45 46 52 53 54
+ 70 72 74 80 85 87 91
c170 72 0 1.26425e-19 $X=7.78 $Y=1.51
c171 70 0 5.91746e-20 $X=7.21 $Y=1.51
c172 54 0 3.13091e-20 $X=6.875 $Y=1.58
c173 33 0 2.54181e-20 $X=4.545 $Y=1.51
c174 19 0 7.37997e-20 $X=7.19 $Y=2.465
r175 80 91 2.7304 $w=3.23e-07 $l=7.7e-08 $layer=LI1_cond $X=7.037 $Y=1.587
+ $X2=6.96 $Y2=1.587
r176 74 85 1.05478 $w=2.93e-07 $l=2.7e-08 $layer=LI1_cond $X=5.973 $Y=1.727
+ $X2=6 $Y2=1.727
r177 71 72 67.2922 $w=3.08e-07 $l=4.3e-07 $layer=POLY_cond $X=7.35 $Y=1.51
+ $X2=7.78 $Y2=1.51
r178 69 71 21.9091 $w=3.08e-07 $l=1.4e-07 $layer=POLY_cond $X=7.21 $Y=1.51
+ $X2=7.35 $Y2=1.51
r179 69 70 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.21
+ $Y=1.51 $X2=7.21 $Y2=1.51
r180 67 69 3.12987 $w=3.08e-07 $l=2e-08 $layer=POLY_cond $X=7.19 $Y=1.51
+ $X2=7.21 $Y2=1.51
r181 54 91 0.141839 $w=3.23e-07 $l=4e-09 $layer=LI1_cond $X=6.956 $Y=1.587
+ $X2=6.96 $Y2=1.587
r182 54 70 5.9927 $w=3.23e-07 $l=1.69e-07 $layer=LI1_cond $X=7.041 $Y=1.587
+ $X2=7.21 $Y2=1.587
r183 54 80 0.141839 $w=3.23e-07 $l=4e-09 $layer=LI1_cond $X=7.041 $Y=1.587
+ $X2=7.037 $Y2=1.587
r184 53 54 16.2679 $w=3.38e-07 $l=3.95e-07 $layer=LI1_cond $X=6.48 $Y=1.665
+ $X2=6.875 $Y2=1.665
r185 53 87 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=6.48 $Y=1.665
+ $X2=6.12 $Y2=1.665
r186 52 87 5.60678 $w=2.93e-07 $l=9.1e-08 $layer=LI1_cond $X=6.029 $Y=1.727
+ $X2=6.12 $Y2=1.727
r187 52 85 1.13291 $w=2.93e-07 $l=2.9e-08 $layer=LI1_cond $X=6.029 $Y=1.727
+ $X2=6 $Y2=1.727
r188 52 74 1.13291 $w=2.93e-07 $l=2.9e-08 $layer=LI1_cond $X=5.944 $Y=1.727
+ $X2=5.973 $Y2=1.727
r189 49 52 6.79746 $w=2.93e-07 $l=1.74e-07 $layer=LI1_cond $X=5.77 $Y=1.727
+ $X2=5.944 $Y2=1.727
r190 48 50 2.02551 $w=3.28e-07 $l=5.8e-08 $layer=LI1_cond $X=5.605 $Y=1.727
+ $X2=5.605 $Y2=1.785
r191 48 49 1.40979 $w=2.95e-07 $l=1.65e-07 $layer=LI1_cond $X=5.605 $Y=1.727
+ $X2=5.77 $Y2=1.727
r192 46 66 46.255 $w=3.35e-07 $l=1.65e-07 $layer=POLY_cond $X=5.602 $Y=1.51
+ $X2=5.602 $Y2=1.675
r193 46 65 46.255 $w=3.35e-07 $l=1.65e-07 $layer=POLY_cond $X=5.602 $Y=1.51
+ $X2=5.602 $Y2=1.345
r194 45 48 7.57819 $w=3.28e-07 $l=2.17e-07 $layer=LI1_cond $X=5.605 $Y=1.51
+ $X2=5.605 $Y2=1.727
r195 45 46 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.605
+ $Y=1.51 $X2=5.605 $Y2=1.51
r196 39 42 0.364908 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=4.715 $Y=1.785
+ $X2=4.63 $Y2=1.785
r197 38 50 4.28565 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=5.44 $Y=1.785
+ $X2=5.605 $Y2=1.785
r198 38 39 44.6717 $w=1.78e-07 $l=7.25e-07 $layer=LI1_cond $X=5.44 $Y=1.785
+ $X2=4.715 $Y2=1.785
r199 36 63 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.16 $Y=1.51
+ $X2=4.16 $Y2=1.675
r200 36 62 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.16 $Y=1.51
+ $X2=4.16 $Y2=1.345
r201 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.16
+ $Y=1.51 $X2=4.16 $Y2=1.51
r202 33 42 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=4.63 $Y=1.51
+ $X2=4.63 $Y2=1.785
r203 33 35 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=4.545 $Y=1.51
+ $X2=4.16 $Y2=1.51
r204 29 72 17.2143 $w=3.08e-07 $l=2.13014e-07 $layer=POLY_cond $X=7.89 $Y=1.675
+ $X2=7.78 $Y2=1.51
r205 29 31 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=7.89 $Y=1.675
+ $X2=7.89 $Y2=2.465
r206 25 72 19.5884 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.78 $Y=1.345
+ $X2=7.78 $Y2=1.51
r207 25 27 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=7.78 $Y=1.345 $X2=7.78
+ $Y2=0.745
r208 21 71 19.5884 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.35 $Y=1.345
+ $X2=7.35 $Y2=1.51
r209 21 23 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=7.35 $Y=1.345 $X2=7.35
+ $Y2=0.745
r210 17 67 19.5884 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.19 $Y=1.675
+ $X2=7.19 $Y2=1.51
r211 17 19 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=7.19 $Y=1.675
+ $X2=7.19 $Y2=2.465
r212 15 66 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=5.51 $Y=2.465
+ $X2=5.51 $Y2=1.675
r213 11 65 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=5.51 $Y=0.655
+ $X2=5.51 $Y2=1.345
r214 7 63 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=4.18 $Y=2.465
+ $X2=4.18 $Y2=1.675
r215 3 62 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=4.18 $Y=0.655
+ $X2=4.18 $Y2=1.345
.ends

.subckt PM_SKY130_FD_SC_LP__HA_4%B 3 7 9 13 17 19 21 23 26 30 34 36 37 40 42 48
+ 49 50 51 53 63 67
c165 67 0 7.37997e-20 $X=7.92 $Y=1.665
c166 42 0 1.36401e-19 $X=5.09 $Y=1.17
c167 9 0 1.61867e-19 $X=4.895 $Y=1.34
r168 64 67 13.4842 $w=3.8e-07 $l=4.2e-07 $layer=LI1_cond $X=8.34 $Y=1.417
+ $X2=7.92 $Y2=1.417
r169 63 64 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.34
+ $Y=1.51 $X2=8.34 $Y2=1.51
r170 61 63 3.44286 $w=2.8e-07 $l=2e-08 $layer=POLY_cond $X=8.32 $Y=1.51 $X2=8.34
+ $Y2=1.51
r171 53 54 30.474 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=5.06 $Y=1.34
+ $X2=5.06 $Y2=1.265
r172 51 67 5.46774 $w=1.7e-07 $l=2.48e-07 $layer=LI1_cond $X=7.92 $Y=1.665
+ $X2=7.92 $Y2=1.417
r173 48 59 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=6.145 $Y=1.26
+ $X2=6.145 $Y2=1.35
r174 47 50 8.69362 $w=2.58e-07 $l=1.65e-07 $layer=LI1_cond $X=6.145 $Y=1.215
+ $X2=6.31 $Y2=1.215
r175 47 49 8.69362 $w=2.58e-07 $l=1.65e-07 $layer=LI1_cond $X=6.145 $Y=1.215
+ $X2=5.98 $Y2=1.215
r176 47 48 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.145
+ $Y=1.26 $X2=6.145 $Y2=1.26
r177 45 56 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.06 $Y=1.43
+ $X2=5.06 $Y2=1.595
r178 45 53 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=5.06 $Y=1.43 $X2=5.06
+ $Y2=1.34
r179 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.06
+ $Y=1.43 $X2=5.06 $Y2=1.43
r180 42 44 12.8421 $w=2.47e-07 $l=2.6e-07 $layer=LI1_cond $X=5.09 $Y=1.17
+ $X2=5.09 $Y2=1.43
r181 40 67 15.4947 $w=3.8e-07 $l=4.72631e-07 $layer=LI1_cond $X=7.555 $Y=1.17
+ $X2=7.92 $Y2=1.417
r182 40 50 81.2246 $w=1.68e-07 $l=1.245e-06 $layer=LI1_cond $X=7.555 $Y=1.17
+ $X2=6.31 $Y2=1.17
r183 39 42 2.92482 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=5.26 $Y=1.17
+ $X2=5.09 $Y2=1.17
r184 39 49 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=5.26 $Y=1.17
+ $X2=5.98 $Y2=1.17
r185 32 63 37.0107 $w=2.8e-07 $l=2.85832e-07 $layer=POLY_cond $X=8.555 $Y=1.345
+ $X2=8.34 $Y2=1.51
r186 32 34 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=8.555 $Y=1.345
+ $X2=8.555 $Y2=0.745
r187 28 61 17.3521 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.32 $Y=1.675
+ $X2=8.32 $Y2=1.51
r188 28 30 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=8.32 $Y=1.675
+ $X2=8.32 $Y2=2.465
r189 24 37 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.76 $Y=1.425
+ $X2=6.76 $Y2=1.35
r190 24 26 533.277 $w=1.5e-07 $l=1.04e-06 $layer=POLY_cond $X=6.76 $Y=1.425
+ $X2=6.76 $Y2=2.465
r191 21 37 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.76 $Y=1.275
+ $X2=6.76 $Y2=1.35
r192 21 23 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=6.76 $Y=1.275
+ $X2=6.76 $Y2=0.745
r193 20 59 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.31 $Y=1.35
+ $X2=6.145 $Y2=1.35
r194 19 37 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.685 $Y=1.35
+ $X2=6.76 $Y2=1.35
r195 19 20 192.287 $w=1.5e-07 $l=3.75e-07 $layer=POLY_cond $X=6.685 $Y=1.35
+ $X2=6.31 $Y2=1.35
r196 17 56 446.106 $w=1.5e-07 $l=8.7e-07 $layer=POLY_cond $X=5.08 $Y=2.465
+ $X2=5.08 $Y2=1.595
r197 13 54 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=5.04 $Y=0.655
+ $X2=5.04 $Y2=1.265
r198 10 36 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.685 $Y=1.34
+ $X2=4.61 $Y2=1.34
r199 9 53 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.895 $Y=1.34
+ $X2=5.06 $Y2=1.34
r200 9 10 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=4.895 $Y=1.34
+ $X2=4.685 $Y2=1.34
r201 5 36 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.61 $Y=1.415
+ $X2=4.61 $Y2=1.34
r202 5 7 538.404 $w=1.5e-07 $l=1.05e-06 $layer=POLY_cond $X=4.61 $Y=1.415
+ $X2=4.61 $Y2=2.465
r203 1 36 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.61 $Y=1.265
+ $X2=4.61 $Y2=1.34
r204 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.61 $Y=1.265
+ $X2=4.61 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__HA_4%VPWR 1 2 3 4 5 6 7 8 9 28 30 36 42 48 54 60 64
+ 66 69 72 75 76 78 79 81 82 84 85 87 89 94 112 119 129 130 136 139 142 149
c174 54 0 1.60386e-19 $X=3.85 $Y=2.28
r175 149 150 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r176 139 140 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r177 136 137 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r178 133 134 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r179 130 150 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.84 $Y=3.33
+ $X2=9.36 $Y2=3.33
r180 129 130 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r181 127 149 12.1981 $w=1.7e-07 $l=2.85e-07 $layer=LI1_cond $X=9.52 $Y=3.33
+ $X2=9.235 $Y2=3.33
r182 127 129 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=9.52 $Y=3.33
+ $X2=9.84 $Y2=3.33
r183 126 150 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=9.36 $Y2=3.33
r184 125 126 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r185 123 126 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=8.88 $Y2=3.33
r186 123 146 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=7.44 $Y2=3.33
r187 122 125 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=7.92 $Y=3.33
+ $X2=8.88 $Y2=3.33
r188 122 123 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r189 120 122 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=7.685 $Y=3.33
+ $X2=7.92 $Y2=3.33
r190 119 149 12.1981 $w=1.7e-07 $l=2.85e-07 $layer=LI1_cond $X=8.95 $Y=3.33
+ $X2=9.235 $Y2=3.33
r191 119 125 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=8.95 $Y=3.33
+ $X2=8.88 $Y2=3.33
r192 118 146 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=7.44 $Y2=3.33
r193 117 118 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r194 115 118 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=3.33
+ $X2=6.96 $Y2=3.33
r195 114 117 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=6 $Y=3.33 $X2=6.96
+ $Y2=3.33
r196 114 115 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r197 112 120 4.88813 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=7.512 $Y=3.33
+ $X2=7.685 $Y2=3.33
r198 112 146 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r199 112 142 8.8521 $w=3.43e-07 $l=2.65e-07 $layer=LI1_cond $X=7.512 $Y=3.33
+ $X2=7.512 $Y2=3.065
r200 112 117 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=7.34 $Y=3.33
+ $X2=6.96 $Y2=3.33
r201 111 115 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=6 $Y2=3.33
r202 110 111 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r203 107 108 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r204 105 108 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.56 $Y2=3.33
r205 104 105 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r206 102 105 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r207 102 140 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r208 101 102 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r209 99 139 7.13466 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=2.255 $Y=3.33
+ $X2=2.127 $Y2=3.33
r210 99 101 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=2.255 $Y=3.33
+ $X2=2.64 $Y2=3.33
r211 98 140 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r212 98 137 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r213 97 98 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r214 95 136 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.435 $Y=3.33
+ $X2=1.27 $Y2=3.33
r215 95 97 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=1.435 $Y=3.33
+ $X2=1.68 $Y2=3.33
r216 94 139 7.13466 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=2 $Y=3.33
+ $X2=2.127 $Y2=3.33
r217 94 97 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=2 $Y=3.33 $X2=1.68
+ $Y2=3.33
r218 93 137 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r219 93 134 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r220 92 93 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r221 90 133 4.50939 $w=1.7e-07 $l=2.88e-07 $layer=LI1_cond $X=0.575 $Y=3.33
+ $X2=0.287 $Y2=3.33
r222 90 92 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=0.575 $Y=3.33
+ $X2=0.72 $Y2=3.33
r223 89 136 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.105 $Y=3.33
+ $X2=1.27 $Y2=3.33
r224 89 92 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=1.105 $Y=3.33
+ $X2=0.72 $Y2=3.33
r225 87 111 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=5.52 $Y2=3.33
r226 87 108 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=4.56 $Y2=3.33
r227 84 110 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=5.56 $Y=3.33
+ $X2=5.52 $Y2=3.33
r228 84 85 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.56 $Y=3.33
+ $X2=5.725 $Y2=3.33
r229 83 114 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=5.89 $Y=3.33 $X2=6
+ $Y2=3.33
r230 83 85 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.89 $Y=3.33
+ $X2=5.725 $Y2=3.33
r231 81 107 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=4.68 $Y=3.33
+ $X2=4.56 $Y2=3.33
r232 81 82 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.68 $Y=3.33
+ $X2=4.845 $Y2=3.33
r233 80 110 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=5.01 $Y=3.33
+ $X2=5.52 $Y2=3.33
r234 80 82 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.01 $Y=3.33
+ $X2=4.845 $Y2=3.33
r235 78 104 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=3.685 $Y=3.33
+ $X2=3.6 $Y2=3.33
r236 78 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.685 $Y=3.33
+ $X2=3.85 $Y2=3.33
r237 77 107 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=4.015 $Y=3.33
+ $X2=4.56 $Y2=3.33
r238 77 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.015 $Y=3.33
+ $X2=3.85 $Y2=3.33
r239 75 101 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=2.895 $Y=3.33
+ $X2=2.64 $Y2=3.33
r240 75 76 6.25164 $w=1.7e-07 $l=1.07e-07 $layer=LI1_cond $X=2.895 $Y=3.33
+ $X2=3.002 $Y2=3.33
r241 74 104 31.9679 $w=1.68e-07 $l=4.9e-07 $layer=LI1_cond $X=3.11 $Y=3.33
+ $X2=3.6 $Y2=3.33
r242 74 76 6.25164 $w=1.7e-07 $l=1.08e-07 $layer=LI1_cond $X=3.11 $Y=3.33
+ $X2=3.002 $Y2=3.33
r243 72 86 18.4391 $w=2.23e-07 $l=3.6e-07 $layer=LI1_cond $X=9.407 $Y=2.27
+ $X2=9.407 $Y2=2.63
r244 67 149 2.39972 $w=5.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.235 $Y=3.245
+ $X2=9.235 $Y2=3.33
r245 67 69 6.19023 $w=5.68e-07 $l=2.95e-07 $layer=LI1_cond $X=9.235 $Y=3.245
+ $X2=9.235 $Y2=2.95
r246 66 86 10.5188 $w=5.68e-07 $l=2.85e-07 $layer=LI1_cond $X=9.235 $Y=2.915
+ $X2=9.235 $Y2=2.63
r247 66 69 0.734434 $w=5.68e-07 $l=3.5e-08 $layer=LI1_cond $X=9.235 $Y=2.915
+ $X2=9.235 $Y2=2.95
r248 62 85 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.725 $Y=3.245
+ $X2=5.725 $Y2=3.33
r249 62 64 26.1919 $w=3.28e-07 $l=7.5e-07 $layer=LI1_cond $X=5.725 $Y=3.245
+ $X2=5.725 $Y2=2.495
r250 58 82 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.845 $Y=3.245
+ $X2=4.845 $Y2=3.33
r251 58 60 26.1919 $w=3.28e-07 $l=7.5e-07 $layer=LI1_cond $X=4.845 $Y=3.245
+ $X2=4.845 $Y2=2.495
r252 54 57 24.0965 $w=3.28e-07 $l=6.9e-07 $layer=LI1_cond $X=3.85 $Y=2.28
+ $X2=3.85 $Y2=2.97
r253 52 79 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.85 $Y=3.245
+ $X2=3.85 $Y2=3.33
r254 52 57 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=3.85 $Y=3.245
+ $X2=3.85 $Y2=2.97
r255 48 51 36.9854 $w=2.13e-07 $l=6.9e-07 $layer=LI1_cond $X=3.002 $Y=2.26
+ $X2=3.002 $Y2=2.95
r256 46 76 0.512231 $w=2.15e-07 $l=8.5e-08 $layer=LI1_cond $X=3.002 $Y=3.245
+ $X2=3.002 $Y2=3.33
r257 46 51 15.8126 $w=2.13e-07 $l=2.95e-07 $layer=LI1_cond $X=3.002 $Y=3.245
+ $X2=3.002 $Y2=2.95
r258 42 45 44.064 $w=2.53e-07 $l=9.75e-07 $layer=LI1_cond $X=2.127 $Y=1.975
+ $X2=2.127 $Y2=2.95
r259 40 139 0.067832 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=2.127 $Y=3.245
+ $X2=2.127 $Y2=3.33
r260 40 45 13.3322 $w=2.53e-07 $l=2.95e-07 $layer=LI1_cond $X=2.127 $Y=3.245
+ $X2=2.127 $Y2=2.95
r261 36 39 26.8903 $w=3.28e-07 $l=7.7e-07 $layer=LI1_cond $X=1.27 $Y=2.18
+ $X2=1.27 $Y2=2.95
r262 34 136 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.27 $Y=3.245
+ $X2=1.27 $Y2=3.33
r263 34 39 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.27 $Y=3.245
+ $X2=1.27 $Y2=2.95
r264 30 33 26.8903 $w=3.28e-07 $l=7.7e-07 $layer=LI1_cond $X=0.41 $Y=2.18
+ $X2=0.41 $Y2=2.95
r265 28 133 3.25678 $w=3.3e-07 $l=1.5995e-07 $layer=LI1_cond $X=0.41 $Y=3.245
+ $X2=0.287 $Y2=3.33
r266 28 33 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.41 $Y=3.245
+ $X2=0.41 $Y2=2.95
r267 9 72 300 $w=1.7e-07 $l=6.02682e-07 $layer=licon1_PDIFF $count=2 $X=8.99
+ $Y=1.835 $X2=9.39 $Y2=2.27
r268 9 69 600 $w=1.7e-07 $l=1.19931e-06 $layer=licon1_PDIFF $count=1 $X=8.99
+ $Y=1.835 $X2=9.165 $Y2=2.95
r269 8 142 600 $w=1.7e-07 $l=1.3515e-06 $layer=licon1_PDIFF $count=1 $X=7.265
+ $Y=1.835 $X2=7.52 $Y2=3.065
r270 7 64 300 $w=1.7e-07 $l=7.26636e-07 $layer=licon1_PDIFF $count=2 $X=5.585
+ $Y=1.835 $X2=5.725 $Y2=2.495
r271 6 60 300 $w=1.7e-07 $l=7.35663e-07 $layer=licon1_PDIFF $count=2 $X=4.685
+ $Y=1.835 $X2=4.845 $Y2=2.495
r272 5 57 400 $w=1.7e-07 $l=1.20297e-06 $layer=licon1_PDIFF $count=1 $X=3.71
+ $Y=1.835 $X2=3.85 $Y2=2.97
r273 5 54 400 $w=1.7e-07 $l=5.10221e-07 $layer=licon1_PDIFF $count=1 $X=3.71
+ $Y=1.835 $X2=3.85 $Y2=2.28
r274 4 51 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=2.85
+ $Y=1.835 $X2=2.99 $Y2=2.95
r275 4 48 400 $w=1.7e-07 $l=4.90026e-07 $layer=licon1_PDIFF $count=1 $X=2.85
+ $Y=1.835 $X2=2.99 $Y2=2.26
r276 3 45 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=1.99
+ $Y=1.835 $X2=2.13 $Y2=2.95
r277 3 42 400 $w=1.7e-07 $l=1.9799e-07 $layer=licon1_PDIFF $count=1 $X=1.99
+ $Y=1.835 $X2=2.13 $Y2=1.975
r278 2 39 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=1.13
+ $Y=1.835 $X2=1.27 $Y2=2.95
r279 2 36 400 $w=1.7e-07 $l=4.09054e-07 $layer=licon1_PDIFF $count=1 $X=1.13
+ $Y=1.835 $X2=1.27 $Y2=2.18
r280 1 33 400 $w=1.7e-07 $l=1.17584e-06 $layer=licon1_PDIFF $count=1 $X=0.285
+ $Y=1.835 $X2=0.41 $Y2=2.95
r281 1 30 400 $w=1.7e-07 $l=4.02679e-07 $layer=licon1_PDIFF $count=1 $X=0.285
+ $Y=1.835 $X2=0.41 $Y2=2.18
.ends

.subckt PM_SKY130_FD_SC_LP__HA_4%SUM 1 2 3 4 13 15 16 19 25 27 29 33 39 42 43 44
+ 45 49 51
r60 49 51 2.92684 $w=3.13e-07 $l=8e-08 $layer=LI1_cond $X=0.247 $Y=1.215
+ $X2=0.247 $Y2=1.295
r61 44 49 2.6726 $w=3.15e-07 $l=8.5e-08 $layer=LI1_cond $X=0.247 $Y=1.13
+ $X2=0.247 $Y2=1.215
r62 44 45 13.4635 $w=3.13e-07 $l=3.68e-07 $layer=LI1_cond $X=0.247 $Y=1.297
+ $X2=0.247 $Y2=1.665
r63 44 51 0.073171 $w=3.13e-07 $l=2e-09 $layer=LI1_cond $X=0.247 $Y=1.297
+ $X2=0.247 $Y2=1.295
r64 41 45 3.29269 $w=3.13e-07 $l=9e-08 $layer=LI1_cond $X=0.247 $Y=1.755
+ $X2=0.247 $Y2=1.665
r65 37 39 36.4833 $w=1.88e-07 $l=6.25e-07 $layer=LI1_cond $X=1.735 $Y=1.045
+ $X2=1.735 $Y2=0.42
r66 33 35 47.6343 $w=2.23e-07 $l=9.3e-07 $layer=LI1_cond $X=1.717 $Y=1.98
+ $X2=1.717 $Y2=2.91
r67 31 33 2.81708 $w=2.23e-07 $l=5.5e-08 $layer=LI1_cond $X=1.717 $Y=1.925
+ $X2=1.717 $Y2=1.98
r68 30 43 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=0.97 $Y=1.13
+ $X2=0.875 $Y2=1.13
r69 29 37 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=1.64 $Y=1.13
+ $X2=1.735 $Y2=1.045
r70 29 30 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.64 $Y=1.13
+ $X2=0.97 $Y2=1.13
r71 28 42 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=0.935 $Y=1.84
+ $X2=0.84 $Y2=1.84
r72 27 31 6.9898 $w=1.7e-07 $l=1.4854e-07 $layer=LI1_cond $X=1.605 $Y=1.84
+ $X2=1.717 $Y2=1.925
r73 27 28 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.605 $Y=1.84
+ $X2=0.935 $Y2=1.84
r74 23 43 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=0.875 $Y=1.045
+ $X2=0.875 $Y2=1.13
r75 23 25 36.4833 $w=1.88e-07 $l=6.25e-07 $layer=LI1_cond $X=0.875 $Y=1.045
+ $X2=0.875 $Y2=0.42
r76 19 21 54.2871 $w=1.88e-07 $l=9.3e-07 $layer=LI1_cond $X=0.84 $Y=1.98
+ $X2=0.84 $Y2=2.91
r77 17 42 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=0.84 $Y=1.925
+ $X2=0.84 $Y2=1.84
r78 17 19 3.21053 $w=1.88e-07 $l=5.5e-08 $layer=LI1_cond $X=0.84 $Y=1.925
+ $X2=0.84 $Y2=1.98
r79 16 41 7.64049 $w=1.7e-07 $l=1.95944e-07 $layer=LI1_cond $X=0.405 $Y=1.84
+ $X2=0.247 $Y2=1.755
r80 15 42 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=0.745 $Y=1.84
+ $X2=0.84 $Y2=1.84
r81 15 16 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=0.745 $Y=1.84
+ $X2=0.405 $Y2=1.84
r82 14 44 4.96789 $w=1.7e-07 $l=1.58e-07 $layer=LI1_cond $X=0.405 $Y=1.13
+ $X2=0.247 $Y2=1.13
r83 13 43 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=0.78 $Y=1.13
+ $X2=0.875 $Y2=1.13
r84 13 14 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.78 $Y=1.13
+ $X2=0.405 $Y2=1.13
r85 4 35 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=1.56
+ $Y=1.835 $X2=1.7 $Y2=2.91
r86 4 33 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.56
+ $Y=1.835 $X2=1.7 $Y2=1.98
r87 3 21 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=0.7
+ $Y=1.835 $X2=0.84 $Y2=2.91
r88 3 19 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.7
+ $Y=1.835 $X2=0.84 $Y2=1.98
r89 2 39 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=1.595
+ $Y=0.235 $X2=1.735 $Y2=0.42
r90 1 25 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=0.735
+ $Y=0.235 $X2=0.875 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__HA_4%COUT 1 2 3 4 14 17 19 21 25 31 33 35 36 37 38
c68 14 0 1.0594e-19 $X=2.51 $Y=1.755
r69 38 50 5.18599 $w=2.98e-07 $l=1.35e-07 $layer=LI1_cond $X=2.575 $Y=2.775
+ $X2=2.575 $Y2=2.91
r70 37 38 14.2135 $w=2.98e-07 $l=3.7e-07 $layer=LI1_cond $X=2.575 $Y=2.405
+ $X2=2.575 $Y2=2.775
r71 36 37 16.3263 $w=2.98e-07 $l=4.25e-07 $layer=LI1_cond $X=2.575 $Y=1.98
+ $X2=2.575 $Y2=2.405
r72 34 36 2.11281 $w=2.98e-07 $l=5.5e-08 $layer=LI1_cond $X=2.575 $Y=1.925
+ $X2=2.575 $Y2=1.98
r73 34 35 3.91525 $w=2.35e-07 $l=8.5e-08 $layer=LI1_cond $X=2.575 $Y=1.925
+ $X2=2.575 $Y2=1.84
r74 29 31 36.4833 $w=1.88e-07 $l=6.25e-07 $layer=LI1_cond $X=3.455 $Y=1.045
+ $X2=3.455 $Y2=0.42
r75 25 27 45.6073 $w=2.33e-07 $l=9.3e-07 $layer=LI1_cond $X=3.397 $Y=1.98
+ $X2=3.397 $Y2=2.91
r76 23 25 2.69721 $w=2.33e-07 $l=5.5e-08 $layer=LI1_cond $X=3.397 $Y=1.925
+ $X2=3.397 $Y2=1.98
r77 22 35 2.53056 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=2.725 $Y=1.84
+ $X2=2.575 $Y2=1.84
r78 21 23 7.04737 $w=1.7e-07 $l=1.53734e-07 $layer=LI1_cond $X=3.28 $Y=1.84
+ $X2=3.397 $Y2=1.925
r79 21 22 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=3.28 $Y=1.84
+ $X2=2.725 $Y2=1.84
r80 20 33 1.54918 $w=1.7e-07 $l=1.33e-07 $layer=LI1_cond $X=2.69 $Y=1.13
+ $X2=2.557 $Y2=1.13
r81 19 29 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=3.36 $Y=1.13
+ $X2=3.455 $Y2=1.045
r82 19 20 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.36 $Y=1.13
+ $X2=2.69 $Y2=1.13
r83 15 33 4.92476 $w=1.8e-07 $l=1.0225e-07 $layer=LI1_cond $X=2.595 $Y=1.045
+ $X2=2.557 $Y2=1.13
r84 15 17 36.4833 $w=1.88e-07 $l=6.25e-07 $layer=LI1_cond $X=2.595 $Y=1.045
+ $X2=2.595 $Y2=0.42
r85 14 35 3.91525 $w=2.35e-07 $l=1.12916e-07 $layer=LI1_cond $X=2.51 $Y=1.755
+ $X2=2.575 $Y2=1.84
r86 13 33 4.92476 $w=1.8e-07 $l=1.05924e-07 $layer=LI1_cond $X=2.51 $Y=1.215
+ $X2=2.557 $Y2=1.13
r87 13 14 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=2.51 $Y=1.215
+ $X2=2.51 $Y2=1.755
r88 4 27 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=3.28
+ $Y=1.835 $X2=3.42 $Y2=2.91
r89 4 25 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=3.28
+ $Y=1.835 $X2=3.42 $Y2=1.98
r90 3 50 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=2.42
+ $Y=1.835 $X2=2.56 $Y2=2.91
r91 3 36 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.42
+ $Y=1.835 $X2=2.56 $Y2=1.98
r92 2 31 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=3.315
+ $Y=0.235 $X2=3.455 $Y2=0.42
r93 1 17 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=2.455
+ $Y=0.235 $X2=2.595 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__HA_4%A_1367_367# 1 2 7 8 12
r29 12 15 3.49225 $w=3.28e-07 $l=1e-07 $layer=LI1_cond $X=8.105 $Y=2.695
+ $X2=8.105 $Y2=2.795
r30 8 11 6.63509 $w=2.85e-07 $l=2.45561e-07 $layer=LI1_cond $X=7.17 $Y=2.695
+ $X2=6.99 $Y2=2.85
r31 7 12 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.94 $Y=2.695
+ $X2=8.105 $Y2=2.695
r32 7 8 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=7.94 $Y=2.695 $X2=7.17
+ $Y2=2.695
r33 2 15 600 $w=1.7e-07 $l=1.02762e-06 $layer=licon1_PDIFF $count=1 $X=7.965
+ $Y=1.835 $X2=8.105 $Y2=2.795
r34 1 11 600 $w=1.7e-07 $l=1.08274e-06 $layer=licon1_PDIFF $count=1 $X=6.835
+ $Y=1.835 $X2=6.975 $Y2=2.85
.ends

.subckt PM_SKY130_FD_SC_LP__HA_4%VGND 1 2 3 4 5 6 7 8 27 29 33 37 41 45 49 53 55
+ 56 58 59 61 62 64 65 66 71 89 93 100 101 104 107 110 118
r163 118 120 3.27831 $w=5.21e-07 $l=2.63873e-07 $layer=LI1_cond $X=8.137 $Y=0.45
+ $X2=8.34 $Y2=0.59
r164 114 116 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0
+ $X2=8.4 $Y2=0
r165 113 118 10.5374 $w=5.21e-07 $l=4.5e-07 $layer=LI1_cond $X=8.137 $Y=0
+ $X2=8.137 $Y2=0.45
r166 113 116 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r167 113 114 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=0
+ $X2=7.92 $Y2=0
r168 110 111 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.96 $Y=0
+ $X2=6.96 $Y2=0
r169 107 108 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0
+ $X2=2.16 $Y2=0
r170 104 105 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r171 101 116 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=9.84 $Y=0
+ $X2=8.4 $Y2=0
r172 100 101 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.84 $Y=0
+ $X2=9.84 $Y2=0
r173 98 113 7.41575 $w=1.7e-07 $l=3.08e-07 $layer=LI1_cond $X=8.445 $Y=0
+ $X2=8.137 $Y2=0
r174 98 100 91.0107 $w=1.68e-07 $l=1.395e-06 $layer=LI1_cond $X=8.445 $Y=0
+ $X2=9.84 $Y2=0
r175 97 114 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0
+ $X2=7.92 $Y2=0
r176 97 111 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0
+ $X2=6.96 $Y2=0
r177 96 97 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r178 94 110 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.22 $Y=0
+ $X2=7.055 $Y2=0
r179 94 96 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=7.22 $Y=0 $X2=7.44
+ $Y2=0
r180 93 113 7.41575 $w=1.7e-07 $l=3.07e-07 $layer=LI1_cond $X=7.83 $Y=0
+ $X2=8.137 $Y2=0
r181 93 96 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=7.83 $Y=0 $X2=7.44
+ $Y2=0
r182 92 111 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.96
+ $Y2=0
r183 91 92 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6 $Y2=0
r184 89 110 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.89 $Y=0
+ $X2=7.055 $Y2=0
r185 89 91 58.0642 $w=1.68e-07 $l=8.9e-07 $layer=LI1_cond $X=6.89 $Y=0 $X2=6
+ $Y2=0
r186 88 92 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=6
+ $Y2=0
r187 87 88 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r188 84 87 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=4.08 $Y=0 $X2=5.52
+ $Y2=0
r189 84 85 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r190 82 85 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r191 81 82 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r192 79 82 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r193 79 108 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0
+ $X2=2.16 $Y2=0
r194 78 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r195 76 107 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.33 $Y=0
+ $X2=2.165 $Y2=0
r196 76 78 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=2.33 $Y=0 $X2=2.64
+ $Y2=0
r197 75 108 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0
+ $X2=2.16 $Y2=0
r198 75 105 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r199 74 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r200 72 104 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.47 $Y=0
+ $X2=1.305 $Y2=0
r201 72 74 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=1.47 $Y=0 $X2=1.68
+ $Y2=0
r202 71 107 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2 $Y=0 $X2=2.165
+ $Y2=0
r203 71 74 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=2 $Y=0 $X2=1.68
+ $Y2=0
r204 70 105 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r205 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r206 66 88 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=5.52
+ $Y2=0
r207 66 85 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=4.08
+ $Y2=0
r208 64 87 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=5.605 $Y=0 $X2=5.52
+ $Y2=0
r209 64 65 7.75133 $w=1.7e-07 $l=1.42e-07 $layer=LI1_cond $X=5.605 $Y=0
+ $X2=5.747 $Y2=0
r210 63 91 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=5.89 $Y=0 $X2=6
+ $Y2=0
r211 63 65 7.75133 $w=1.7e-07 $l=1.43e-07 $layer=LI1_cond $X=5.89 $Y=0 $X2=5.747
+ $Y2=0
r212 61 81 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=3.72 $Y=0 $X2=3.6
+ $Y2=0
r213 61 62 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=3.72 $Y=0 $X2=3.89
+ $Y2=0
r214 60 84 1.30481 $w=1.68e-07 $l=2e-08 $layer=LI1_cond $X=4.06 $Y=0 $X2=4.08
+ $Y2=0
r215 60 62 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=4.06 $Y=0 $X2=3.89
+ $Y2=0
r216 58 78 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=2.86 $Y=0 $X2=2.64
+ $Y2=0
r217 58 59 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.86 $Y=0 $X2=3.025
+ $Y2=0
r218 57 81 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=3.19 $Y=0 $X2=3.6
+ $Y2=0
r219 57 59 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.19 $Y=0 $X2=3.025
+ $Y2=0
r220 55 69 2.87059 $w=1.7e-07 $l=4e-08 $layer=LI1_cond $X=0.28 $Y=0 $X2=0.24
+ $Y2=0
r221 55 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.28 $Y=0 $X2=0.445
+ $Y2=0
r222 51 110 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.055 $Y=0.085
+ $X2=7.055 $Y2=0
r223 51 53 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=7.055 $Y=0.085
+ $X2=7.055 $Y2=0.45
r224 47 65 0.432977 $w=2.85e-07 $l=8.5e-08 $layer=LI1_cond $X=5.747 $Y=0.085
+ $X2=5.747 $Y2=0
r225 47 49 11.9288 $w=2.83e-07 $l=2.95e-07 $layer=LI1_cond $X=5.747 $Y=0.085
+ $X2=5.747 $Y2=0.38
r226 43 62 0.987631 $w=3.4e-07 $l=8.5e-08 $layer=LI1_cond $X=3.89 $Y=0.085
+ $X2=3.89 $Y2=0
r227 43 45 9.32123 $w=3.38e-07 $l=2.75e-07 $layer=LI1_cond $X=3.89 $Y=0.085
+ $X2=3.89 $Y2=0.36
r228 39 59 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.025 $Y=0.085
+ $X2=3.025 $Y2=0
r229 39 41 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=3.025 $Y=0.085
+ $X2=3.025 $Y2=0.36
r230 35 107 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.165 $Y=0.085
+ $X2=2.165 $Y2=0
r231 35 37 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=2.165 $Y=0.085
+ $X2=2.165 $Y2=0.55
r232 31 104 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.305 $Y=0.085
+ $X2=1.305 $Y2=0
r233 31 33 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=1.305 $Y=0.085
+ $X2=1.305 $Y2=0.36
r234 30 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.61 $Y=0 $X2=0.445
+ $Y2=0
r235 29 104 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.14 $Y=0
+ $X2=1.305 $Y2=0
r236 29 30 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=1.14 $Y=0 $X2=0.61
+ $Y2=0
r237 25 56 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.445 $Y=0.085
+ $X2=0.445 $Y2=0
r238 25 27 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=0.445 $Y=0.085
+ $X2=0.445 $Y2=0.36
r239 8 120 182 $w=1.7e-07 $l=6.03117e-07 $layer=licon1_NDIFF $count=1 $X=7.855
+ $Y=0.325 $X2=8.34 $Y2=0.59
r240 8 118 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=7.855
+ $Y=0.325 $X2=7.995 $Y2=0.45
r241 7 53 182 $w=1.7e-07 $l=2.755e-07 $layer=licon1_NDIFF $count=1 $X=6.835
+ $Y=0.325 $X2=7.055 $Y2=0.45
r242 6 49 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.585
+ $Y=0.235 $X2=5.725 $Y2=0.38
r243 5 45 91 $w=1.7e-07 $l=2.03101e-07 $layer=licon1_NDIFF $count=2 $X=3.745
+ $Y=0.235 $X2=3.895 $Y2=0.36
r244 4 41 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=2.885
+ $Y=0.235 $X2=3.025 $Y2=0.36
r245 3 37 182 $w=1.7e-07 $l=3.78583e-07 $layer=licon1_NDIFF $count=1 $X=2.025
+ $Y=0.235 $X2=2.165 $Y2=0.55
r246 2 33 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=1.165
+ $Y=0.235 $X2=1.305 $Y2=0.36
r247 1 27 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.3
+ $Y=0.235 $X2=0.445 $Y2=0.36
.ends

.subckt PM_SKY130_FD_SC_LP__HA_4%A_851_47# 1 2 9 14 16
c28 9 0 1.36401e-19 $X=5.105 $Y=0.35
r29 10 14 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.56 $Y=0.35
+ $X2=4.395 $Y2=0.35
r30 9 16 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.105 $Y=0.35
+ $X2=5.27 $Y2=0.35
r31 9 10 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=5.105 $Y=0.35
+ $X2=4.56 $Y2=0.35
r32 2 16 91 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_NDIFF $count=2 $X=5.115
+ $Y=0.235 $X2=5.27 $Y2=0.38
r33 1 14 91 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_NDIFF $count=2 $X=4.255
+ $Y=0.235 $X2=4.395 $Y2=0.37
.ends

.subckt PM_SKY130_FD_SC_LP__HA_4%A_1284_65# 1 2 3 4 15 17 18 21 23 25 30 31 32
+ 35 38 39
c87 23 0 1.26425e-19 $X=7.905 $Y=0.825
r88 39 41 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=7.99 $Y=0.825
+ $X2=7.99 $Y2=1.01
r89 33 35 1.61342 $w=2.48e-07 $l=3.5e-08 $layer=LI1_cond $X=9.805 $Y=0.435
+ $X2=9.805 $Y2=0.47
r90 31 33 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=9.68 $Y=0.35
+ $X2=9.805 $Y2=0.435
r91 31 32 53.8235 $w=1.68e-07 $l=8.25e-07 $layer=LI1_cond $X=9.68 $Y=0.35
+ $X2=8.855 $Y2=0.35
r92 28 30 26.5598 $w=1.88e-07 $l=4.55e-07 $layer=LI1_cond $X=8.76 $Y=0.925
+ $X2=8.76 $Y2=0.47
r93 27 32 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=8.76 $Y=0.435
+ $X2=8.855 $Y2=0.35
r94 27 30 2.04306 $w=1.88e-07 $l=3.5e-08 $layer=LI1_cond $X=8.76 $Y=0.435
+ $X2=8.76 $Y2=0.47
r95 26 41 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.075 $Y=1.01
+ $X2=7.99 $Y2=1.01
r96 25 28 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=8.665 $Y=1.01
+ $X2=8.76 $Y2=0.925
r97 25 26 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=8.665 $Y=1.01
+ $X2=8.075 $Y2=1.01
r98 24 38 6.78838 $w=1.85e-07 $l=1.32476e-07 $layer=LI1_cond $X=7.66 $Y=0.825
+ $X2=7.53 $Y2=0.82
r99 23 39 0.364908 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=7.905 $Y=0.825
+ $X2=7.99 $Y2=0.825
r100 23 24 15.096 $w=1.78e-07 $l=2.45e-07 $layer=LI1_cond $X=7.905 $Y=0.825
+ $X2=7.66 $Y2=0.825
r101 19 38 0.150961 $w=2.6e-07 $l=9.5e-08 $layer=LI1_cond $X=7.53 $Y=0.725
+ $X2=7.53 $Y2=0.82
r102 19 21 12.1893 $w=2.58e-07 $l=2.75e-07 $layer=LI1_cond $X=7.53 $Y=0.725
+ $X2=7.53 $Y2=0.45
r103 17 38 6.78838 $w=1.85e-07 $l=1.3e-07 $layer=LI1_cond $X=7.4 $Y=0.82
+ $X2=7.53 $Y2=0.82
r104 17 18 40.2775 $w=1.88e-07 $l=6.9e-07 $layer=LI1_cond $X=7.4 $Y=0.82
+ $X2=6.71 $Y2=0.82
r105 13 18 7.47963 $w=1.9e-07 $l=2.07123e-07 $layer=LI1_cond $X=6.545 $Y=0.725
+ $X2=6.71 $Y2=0.82
r106 13 15 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=6.545 $Y=0.725
+ $X2=6.545 $Y2=0.47
r107 4 35 91 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=2 $X=9.49
+ $Y=0.325 $X2=9.765 $Y2=0.47
r108 3 30 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=8.63
+ $Y=0.325 $X2=8.77 $Y2=0.47
r109 2 38 182 $w=1.7e-07 $l=5.60647e-07 $layer=licon1_NDIFF $count=1 $X=7.425
+ $Y=0.325 $X2=7.565 $Y2=0.82
r110 2 21 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=7.425
+ $Y=0.325 $X2=7.565 $Y2=0.45
r111 1 15 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=6.42
+ $Y=0.325 $X2=6.545 $Y2=0.47
.ends

