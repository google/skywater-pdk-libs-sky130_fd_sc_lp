* File: sky130_fd_sc_lp__o41ai_0.pxi.spice
* Created: Wed Sep  2 10:28:03 2020
* 
x_PM_SKY130_FD_SC_LP__O41AI_0%B1 N_B1_c_78_n N_B1_M1000_g N_B1_M1006_g
+ N_B1_c_79_n N_B1_c_80_n N_B1_c_86_n B1 B1 B1 N_B1_c_82_n N_B1_c_83_n
+ PM_SKY130_FD_SC_LP__O41AI_0%B1
x_PM_SKY130_FD_SC_LP__O41AI_0%A4 N_A4_c_122_n N_A4_M1004_g N_A4_M1001_g A4 A4
+ N_A4_c_125_n PM_SKY130_FD_SC_LP__O41AI_0%A4
x_PM_SKY130_FD_SC_LP__O41AI_0%A3 N_A3_c_171_n N_A3_M1003_g N_A3_M1002_g
+ N_A3_c_168_n A3 A3 A3 A3 A3 N_A3_c_170_n A3 A3 PM_SKY130_FD_SC_LP__O41AI_0%A3
x_PM_SKY130_FD_SC_LP__O41AI_0%A2 N_A2_c_217_n N_A2_M1007_g N_A2_M1009_g
+ N_A2_c_219_n N_A2_c_220_n N_A2_c_225_n A2 A2 A2 N_A2_c_222_n
+ PM_SKY130_FD_SC_LP__O41AI_0%A2
x_PM_SKY130_FD_SC_LP__O41AI_0%A1 N_A1_M1008_g N_A1_M1005_g N_A1_c_265_n
+ N_A1_c_269_n N_A1_c_270_n N_A1_c_271_n A1 A1 A1 N_A1_c_267_n
+ PM_SKY130_FD_SC_LP__O41AI_0%A1
x_PM_SKY130_FD_SC_LP__O41AI_0%VPWR N_VPWR_M1000_s N_VPWR_M1008_d N_VPWR_c_298_n
+ N_VPWR_c_299_n N_VPWR_c_300_n N_VPWR_c_301_n N_VPWR_c_302_n VPWR
+ N_VPWR_c_303_n N_VPWR_c_297_n N_VPWR_c_305_n PM_SKY130_FD_SC_LP__O41AI_0%VPWR
x_PM_SKY130_FD_SC_LP__O41AI_0%Y N_Y_M1006_s N_Y_M1000_d N_Y_c_333_n N_Y_c_334_n
+ Y Y Y Y Y Y N_Y_c_332_n N_Y_c_336_n Y PM_SKY130_FD_SC_LP__O41AI_0%Y
x_PM_SKY130_FD_SC_LP__O41AI_0%A_218_57# N_A_218_57#_M1006_d N_A_218_57#_M1002_d
+ N_A_218_57#_M1005_d N_A_218_57#_c_366_n N_A_218_57#_c_367_n
+ N_A_218_57#_c_368_n N_A_218_57#_c_369_n N_A_218_57#_c_370_n
+ N_A_218_57#_c_371_n N_A_218_57#_c_372_n PM_SKY130_FD_SC_LP__O41AI_0%A_218_57#
x_PM_SKY130_FD_SC_LP__O41AI_0%VGND N_VGND_M1001_d N_VGND_M1009_d N_VGND_c_411_n
+ N_VGND_c_412_n VGND N_VGND_c_413_n N_VGND_c_414_n N_VGND_c_415_n
+ N_VGND_c_416_n N_VGND_c_417_n N_VGND_c_418_n PM_SKY130_FD_SC_LP__O41AI_0%VGND
cc_1 VNB N_B1_c_78_n 0.0247985f $X=-0.19 $Y=-0.245 $X2=0.74 $Y2=1.26
cc_2 VNB N_B1_c_79_n 0.0255479f $X=-0.19 $Y=-0.245 $X2=0.74 $Y2=1.485
cc_3 VNB N_B1_c_80_n 0.0124559f $X=-0.19 $Y=-0.245 $X2=0.86 $Y2=2.115
cc_4 VNB B1 0.00425423f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.84
cc_5 VNB N_B1_c_82_n 0.0371551f $X=-0.19 $Y=-0.245 $X2=0.68 $Y2=0.98
cc_6 VNB N_B1_c_83_n 0.0210229f $X=-0.19 $Y=-0.245 $X2=0.802 $Y2=0.815
cc_7 VNB N_A4_c_122_n 0.0175448f $X=-0.19 $Y=-0.245 $X2=0.74 $Y2=1.26
cc_8 VNB N_A4_M1001_g 0.0391164f $X=-0.19 $Y=-0.245 $X2=1.015 $Y2=0.815
cc_9 VNB A4 0.00605736f $X=-0.19 $Y=-0.245 $X2=1.015 $Y2=0.495
cc_10 VNB N_A4_c_125_n 0.0164897f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_11 VNB N_A3_M1002_g 0.0368711f $X=-0.19 $Y=-0.245 $X2=0.95 $Y2=2.735
cc_12 VNB N_A3_c_168_n 0.0172416f $X=-0.19 $Y=-0.245 $X2=1.015 $Y2=0.495
cc_13 VNB A3 0.00622815f $X=-0.19 $Y=-0.245 $X2=0.74 $Y2=1.485
cc_14 VNB N_A3_c_170_n 0.0153056f $X=-0.19 $Y=-0.245 $X2=0.802 $Y2=0.995
cc_15 VNB N_A2_c_217_n 0.00724219f $X=-0.19 $Y=-0.245 $X2=0.74 $Y2=0.995
cc_16 VNB N_A2_M1009_g 0.0243905f $X=-0.19 $Y=-0.245 $X2=1.015 $Y2=0.815
cc_17 VNB N_A2_c_219_n 0.00826315f $X=-0.19 $Y=-0.245 $X2=0.86 $Y2=2.115
cc_18 VNB N_A2_c_220_n 0.0172416f $X=-0.19 $Y=-0.245 $X2=0.86 $Y2=2.265
cc_19 VNB A2 0.0053889f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_20 VNB N_A2_c_222_n 0.0137646f $X=-0.19 $Y=-0.245 $X2=0.68 $Y2=0.98
cc_21 VNB N_A1_M1005_g 0.048676f $X=-0.19 $Y=-0.245 $X2=0.95 $Y2=2.735
cc_22 VNB N_A1_c_265_n 0.0205269f $X=-0.19 $Y=-0.245 $X2=1.015 $Y2=0.495
cc_23 VNB A1 0.021494f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A1_c_267_n 0.0289472f $X=-0.19 $Y=-0.245 $X2=0.802 $Y2=0.995
cc_25 VNB N_VPWR_c_297_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB Y 0.0553139f $X=-0.19 $Y=-0.245 $X2=0.86 $Y2=2.265
cc_27 VNB N_Y_c_332_n 0.0155701f $X=-0.19 $Y=-0.245 $X2=0.745 $Y2=0.925
cc_28 VNB N_A_218_57#_c_366_n 0.00259016f $X=-0.19 $Y=-0.245 $X2=0.74 $Y2=1.485
cc_29 VNB N_A_218_57#_c_367_n 0.00859778f $X=-0.19 $Y=-0.245 $X2=0.86 $Y2=2.265
cc_30 VNB N_A_218_57#_c_368_n 0.00365738f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.84
cc_31 VNB N_A_218_57#_c_369_n 0.00104496f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_218_57#_c_370_n 0.0174243f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_218_57#_c_371_n 0.0208209f $X=-0.19 $Y=-0.245 $X2=0.802 $Y2=0.815
cc_34 VNB N_A_218_57#_c_372_n 0.00866545f $X=-0.19 $Y=-0.245 $X2=0.745 $Y2=0.925
cc_35 VNB N_VGND_c_411_n 0.00652431f $X=-0.19 $Y=-0.245 $X2=1.015 $Y2=0.815
cc_36 VNB N_VGND_c_412_n 0.00648667f $X=-0.19 $Y=-0.245 $X2=0.86 $Y2=2.115
cc_37 VNB N_VGND_c_413_n 0.0420235f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_38 VNB N_VGND_c_414_n 0.0171006f $X=-0.19 $Y=-0.245 $X2=0.802 $Y2=0.995
cc_39 VNB N_VGND_c_415_n 0.0175832f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_416_n 0.202556f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_417_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_418_n 0.00615512f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VPB N_B1_M1000_g 0.0249964f $X=-0.19 $Y=1.655 $X2=0.95 $Y2=2.735
cc_44 VPB N_B1_c_80_n 0.0337128f $X=-0.19 $Y=1.655 $X2=0.86 $Y2=2.115
cc_45 VPB N_B1_c_86_n 0.0192538f $X=-0.19 $Y=1.655 $X2=0.86 $Y2=2.265
cc_46 VPB B1 0.00283768f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=0.84
cc_47 VPB N_A4_c_122_n 0.0442881f $X=-0.19 $Y=1.655 $X2=0.74 $Y2=1.26
cc_48 VPB N_A4_M1004_g 0.0187368f $X=-0.19 $Y=1.655 $X2=0.95 $Y2=2.265
cc_49 VPB A4 0.00329903f $X=-0.19 $Y=1.655 $X2=1.015 $Y2=0.495
cc_50 VPB N_A3_c_171_n 0.0153056f $X=-0.19 $Y=1.655 $X2=0.74 $Y2=0.995
cc_51 VPB N_A3_M1003_g 0.0358005f $X=-0.19 $Y=1.655 $X2=0.83 $Y2=1.485
cc_52 VPB N_A3_c_168_n 0.00364608f $X=-0.19 $Y=1.655 $X2=1.015 $Y2=0.495
cc_53 VPB A3 0.00413981f $X=-0.19 $Y=1.655 $X2=0.74 $Y2=1.485
cc_54 VPB A3 0.00667562f $X=-0.19 $Y=1.655 $X2=0.86 $Y2=2.265
cc_55 VPB A3 0.00195351f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_56 VPB N_A2_M1007_g 0.0380527f $X=-0.19 $Y=1.655 $X2=0.95 $Y2=2.265
cc_57 VPB N_A2_c_220_n 0.00364608f $X=-0.19 $Y=1.655 $X2=0.86 $Y2=2.265
cc_58 VPB N_A2_c_225_n 0.0153343f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=0.84
cc_59 VPB A2 0.0112976f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_60 VPB N_A1_M1008_g 0.0232289f $X=-0.19 $Y=1.655 $X2=0.83 $Y2=1.485
cc_61 VPB N_A1_c_269_n 0.0159432f $X=-0.19 $Y=1.655 $X2=0.74 $Y2=1.485
cc_62 VPB N_A1_c_270_n 0.0242572f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=0.84
cc_63 VPB N_A1_c_271_n 0.0289472f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_64 VPB A1 0.0297991f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_298_n 0.0345701f $X=-0.19 $Y=1.655 $X2=1.015 $Y2=0.815
cc_66 VPB N_VPWR_c_299_n 0.0331777f $X=-0.19 $Y=1.655 $X2=0.86 $Y2=2.115
cc_67 VPB N_VPWR_c_300_n 0.0108943f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=0.84
cc_68 VPB N_VPWR_c_301_n 0.0505137f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_69 VPB N_VPWR_c_302_n 0.00607754f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_70 VPB N_VPWR_c_303_n 0.0202818f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_71 VPB N_VPWR_c_297_n 0.0951425f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_72 VPB N_VPWR_c_305_n 0.00555219f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_73 VPB N_Y_c_333_n 0.0176528f $X=-0.19 $Y=1.655 $X2=0.95 $Y2=2.735
cc_74 VPB N_Y_c_334_n 0.00391851f $X=-0.19 $Y=1.655 $X2=1.015 $Y2=0.495
cc_75 VPB Y 0.0229668f $X=-0.19 $Y=1.655 $X2=0.86 $Y2=2.265
cc_76 VPB N_Y_c_336_n 0.021652f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_77 N_B1_c_79_n N_A4_c_122_n 0.0207252f $X=0.74 $Y=1.485 $X2=0 $Y2=0
cc_78 N_B1_c_80_n N_A4_c_122_n 0.0111169f $X=0.86 $Y=2.115 $X2=0 $Y2=0
cc_79 N_B1_c_86_n N_A4_c_122_n 0.0083288f $X=0.86 $Y=2.265 $X2=0 $Y2=0
cc_80 N_B1_M1000_g N_A4_M1004_g 0.0121152f $X=0.95 $Y=2.735 $X2=0 $Y2=0
cc_81 N_B1_c_78_n N_A4_M1001_g 0.00691819f $X=0.74 $Y=1.26 $X2=0 $Y2=0
cc_82 B1 N_A4_M1001_g 0.001145f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_83 N_B1_c_83_n N_A4_M1001_g 0.0192065f $X=0.802 $Y=0.815 $X2=0 $Y2=0
cc_84 N_B1_c_78_n A4 0.00455303f $X=0.74 $Y=1.26 $X2=0 $Y2=0
cc_85 B1 A4 0.0509709f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_86 N_B1_c_82_n A4 0.00110323f $X=0.68 $Y=0.98 $X2=0 $Y2=0
cc_87 N_B1_c_78_n N_A4_c_125_n 0.0207252f $X=0.74 $Y=1.26 $X2=0 $Y2=0
cc_88 B1 N_A4_c_125_n 5.80364e-19 $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_89 N_B1_M1000_g N_VPWR_c_298_n 0.00501097f $X=0.95 $Y=2.735 $X2=0 $Y2=0
cc_90 N_B1_c_86_n N_VPWR_c_298_n 0.00465828f $X=0.86 $Y=2.265 $X2=0 $Y2=0
cc_91 N_B1_M1000_g N_VPWR_c_301_n 0.00545548f $X=0.95 $Y=2.735 $X2=0 $Y2=0
cc_92 N_B1_M1000_g N_VPWR_c_297_n 0.0113288f $X=0.95 $Y=2.735 $X2=0 $Y2=0
cc_93 N_B1_c_79_n N_Y_c_333_n 0.00251706f $X=0.74 $Y=1.485 $X2=0 $Y2=0
cc_94 N_B1_c_80_n N_Y_c_333_n 0.00968235f $X=0.86 $Y=2.115 $X2=0 $Y2=0
cc_95 N_B1_c_86_n N_Y_c_333_n 0.0162199f $X=0.86 $Y=2.265 $X2=0 $Y2=0
cc_96 B1 N_Y_c_333_n 0.0203662f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_97 N_B1_c_86_n N_Y_c_334_n 0.00523734f $X=0.86 $Y=2.265 $X2=0 $Y2=0
cc_98 N_B1_c_80_n Y 0.00895329f $X=0.86 $Y=2.115 $X2=0 $Y2=0
cc_99 B1 Y 0.0790616f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_100 N_B1_c_82_n Y 0.0179485f $X=0.68 $Y=0.98 $X2=0 $Y2=0
cc_101 N_B1_c_83_n Y 0.00394996f $X=0.802 $Y=0.815 $X2=0 $Y2=0
cc_102 B1 Y 0.0234363f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_103 N_B1_c_82_n Y 0.0057145f $X=0.68 $Y=0.98 $X2=0 $Y2=0
cc_104 B1 N_A_218_57#_c_366_n 9.72828e-19 $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_105 N_B1_c_83_n N_A_218_57#_c_366_n 0.00322908f $X=0.802 $Y=0.815 $X2=0 $Y2=0
cc_106 B1 N_A_218_57#_c_368_n 0.0123431f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_107 N_B1_c_82_n N_A_218_57#_c_368_n 0.0018709f $X=0.68 $Y=0.98 $X2=0 $Y2=0
cc_108 N_B1_c_83_n N_VGND_c_413_n 0.0053602f $X=0.802 $Y=0.815 $X2=0 $Y2=0
cc_109 N_B1_c_82_n N_VGND_c_416_n 2.5959e-19 $X=0.68 $Y=0.98 $X2=0 $Y2=0
cc_110 N_B1_c_83_n N_VGND_c_416_n 0.0113452f $X=0.802 $Y=0.815 $X2=0 $Y2=0
cc_111 N_A4_c_122_n N_A3_M1003_g 0.0402723f $X=1.347 $Y=1.703 $X2=0 $Y2=0
cc_112 N_A4_M1001_g N_A3_M1002_g 0.0214173f $X=1.445 $Y=0.495 $X2=0 $Y2=0
cc_113 N_A4_c_122_n N_A3_c_168_n 0.0207106f $X=1.347 $Y=1.703 $X2=0 $Y2=0
cc_114 N_A4_M1001_g A3 0.0107184f $X=1.445 $Y=0.495 $X2=0 $Y2=0
cc_115 A4 A3 0.0547608f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_116 N_A4_c_122_n A3 0.00662155f $X=1.347 $Y=1.703 $X2=0 $Y2=0
cc_117 A4 N_A3_c_170_n 5.51855e-19 $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_118 N_A4_c_125_n N_A3_c_170_n 0.0207106f $X=1.34 $Y=1.37 $X2=0 $Y2=0
cc_119 N_A4_M1004_g A3 0.00300987f $X=1.38 $Y=2.735 $X2=0 $Y2=0
cc_120 N_A4_M1004_g N_VPWR_c_301_n 0.00511657f $X=1.38 $Y=2.735 $X2=0 $Y2=0
cc_121 N_A4_M1004_g N_VPWR_c_297_n 0.00983613f $X=1.38 $Y=2.735 $X2=0 $Y2=0
cc_122 N_A4_c_122_n N_Y_c_333_n 0.0063185f $X=1.347 $Y=1.703 $X2=0 $Y2=0
cc_123 A4 N_Y_c_333_n 0.0227154f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_124 N_A4_c_122_n N_Y_c_334_n 0.00198944f $X=1.347 $Y=1.703 $X2=0 $Y2=0
cc_125 N_A4_M1004_g N_Y_c_334_n 0.0102188f $X=1.38 $Y=2.735 $X2=0 $Y2=0
cc_126 A4 Y 8.07776e-19 $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_127 N_A4_M1001_g N_A_218_57#_c_366_n 0.0020031f $X=1.445 $Y=0.495 $X2=0 $Y2=0
cc_128 N_A4_M1001_g N_A_218_57#_c_367_n 0.0133093f $X=1.445 $Y=0.495 $X2=0 $Y2=0
cc_129 A4 N_A_218_57#_c_367_n 0.00350455f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_130 N_A4_M1001_g N_A_218_57#_c_368_n 0.00162415f $X=1.445 $Y=0.495 $X2=0
+ $Y2=0
cc_131 A4 N_A_218_57#_c_368_n 0.0211942f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_132 N_A4_c_125_n N_A_218_57#_c_368_n 0.00148112f $X=1.34 $Y=1.37 $X2=0 $Y2=0
cc_133 N_A4_M1001_g N_A_218_57#_c_369_n 5.15328e-19 $X=1.445 $Y=0.495 $X2=0
+ $Y2=0
cc_134 N_A4_M1001_g N_VGND_c_411_n 0.00344564f $X=1.445 $Y=0.495 $X2=0 $Y2=0
cc_135 N_A4_M1001_g N_VGND_c_413_n 0.0053602f $X=1.445 $Y=0.495 $X2=0 $Y2=0
cc_136 N_A4_M1001_g N_VGND_c_416_n 0.00592151f $X=1.445 $Y=0.495 $X2=0 $Y2=0
cc_137 N_A3_M1002_g N_A2_c_217_n 0.0149859f $X=1.97 $Y=0.495 $X2=-0.19
+ $Y2=-0.245
cc_138 N_A3_M1003_g N_A2_M1007_g 0.0501884f $X=1.895 $Y=2.735 $X2=0 $Y2=0
cc_139 A3 N_A2_M1007_g 0.0138504f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_140 N_A3_M1002_g N_A2_M1009_g 0.0184426f $X=1.97 $Y=0.495 $X2=0 $Y2=0
cc_141 A3 N_A2_c_219_n 2.30253e-19 $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_142 N_A3_c_168_n N_A2_c_220_n 0.0135694f $X=1.895 $Y=1.715 $X2=0 $Y2=0
cc_143 N_A3_c_171_n N_A2_c_225_n 0.0135694f $X=1.895 $Y=1.88 $X2=0 $Y2=0
cc_144 N_A3_M1003_g A2 3.97208e-19 $X=1.895 $Y=2.735 $X2=0 $Y2=0
cc_145 A3 A2 0.0729476f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_146 N_A3_c_170_n A2 0.00232271f $X=1.895 $Y=1.375 $X2=0 $Y2=0
cc_147 A3 N_A2_c_222_n 0.00232293f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_148 N_A3_c_170_n N_A2_c_222_n 0.0135694f $X=1.895 $Y=1.375 $X2=0 $Y2=0
cc_149 A3 N_VPWR_c_299_n 0.0175026f $X=1.68 $Y=2.405 $X2=0 $Y2=0
cc_150 N_A3_M1003_g N_VPWR_c_301_n 0.00341069f $X=1.895 $Y=2.735 $X2=0 $Y2=0
cc_151 A3 N_VPWR_c_301_n 0.0261455f $X=1.68 $Y=2.405 $X2=0 $Y2=0
cc_152 N_A3_M1003_g N_VPWR_c_297_n 0.00522128f $X=1.895 $Y=2.735 $X2=0 $Y2=0
cc_153 A3 N_VPWR_c_297_n 0.0204413f $X=1.68 $Y=2.405 $X2=0 $Y2=0
cc_154 A3 N_Y_c_333_n 0.0145697f $X=1.595 $Y=1.95 $X2=0 $Y2=0
cc_155 N_A3_M1003_g N_Y_c_334_n 7.43211e-19 $X=1.895 $Y=2.735 $X2=0 $Y2=0
cc_156 A3 N_Y_c_334_n 0.0379813f $X=1.595 $Y=1.95 $X2=0 $Y2=0
cc_157 A3 A_291_483# 0.00705077f $X=1.68 $Y=2.405 $X2=-0.19 $Y2=-0.245
cc_158 A3 A_394_483# 0.00980737f $X=1.68 $Y=2.405 $X2=-0.19 $Y2=-0.245
cc_159 N_A3_M1002_g N_A_218_57#_c_367_n 0.0100356f $X=1.97 $Y=0.495 $X2=0 $Y2=0
cc_160 A3 N_A_218_57#_c_367_n 0.036263f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_161 N_A3_c_170_n N_A_218_57#_c_367_n 0.00102716f $X=1.895 $Y=1.375 $X2=0
+ $Y2=0
cc_162 N_A3_M1002_g N_A_218_57#_c_369_n 0.00747368f $X=1.97 $Y=0.495 $X2=0 $Y2=0
cc_163 N_A3_M1002_g N_A_218_57#_c_372_n 0.00199038f $X=1.97 $Y=0.495 $X2=0 $Y2=0
cc_164 A3 N_A_218_57#_c_372_n 0.00173297f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_165 N_A3_M1002_g N_VGND_c_411_n 0.00190645f $X=1.97 $Y=0.495 $X2=0 $Y2=0
cc_166 N_A3_M1002_g N_VGND_c_414_n 0.00530767f $X=1.97 $Y=0.495 $X2=0 $Y2=0
cc_167 N_A3_M1002_g N_VGND_c_416_n 0.0058535f $X=1.97 $Y=0.495 $X2=0 $Y2=0
cc_168 N_A2_M1009_g N_A1_M1005_g 0.0246249f $X=2.4 $Y=0.495 $X2=0 $Y2=0
cc_169 A2 N_A1_M1005_g 0.00748444f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_170 N_A2_c_220_n N_A1_c_265_n 0.0140366f $X=2.435 $Y=1.715 $X2=0 $Y2=0
cc_171 N_A2_M1007_g N_A1_c_269_n 0.00597573f $X=2.345 $Y=2.735 $X2=0 $Y2=0
cc_172 N_A2_M1007_g N_A1_c_270_n 0.0650144f $X=2.345 $Y=2.735 $X2=0 $Y2=0
cc_173 A2 N_A1_c_270_n 0.0128115f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_174 N_A2_c_225_n N_A1_c_271_n 0.0140366f $X=2.435 $Y=1.88 $X2=0 $Y2=0
cc_175 N_A2_M1007_g A1 2.04672e-19 $X=2.345 $Y=2.735 $X2=0 $Y2=0
cc_176 A2 A1 0.0831356f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_177 N_A2_c_222_n A1 5.39125e-19 $X=2.435 $Y=1.375 $X2=0 $Y2=0
cc_178 N_A2_c_222_n N_A1_c_267_n 0.0140366f $X=2.435 $Y=1.375 $X2=0 $Y2=0
cc_179 N_A2_M1007_g N_VPWR_c_299_n 0.00331874f $X=2.345 $Y=2.735 $X2=0 $Y2=0
cc_180 A2 N_VPWR_c_299_n 0.00279348f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_181 N_A2_M1007_g N_VPWR_c_301_n 0.00545548f $X=2.345 $Y=2.735 $X2=0 $Y2=0
cc_182 N_A2_M1007_g N_VPWR_c_297_n 0.0104754f $X=2.345 $Y=2.735 $X2=0 $Y2=0
cc_183 N_A2_M1009_g N_A_218_57#_c_369_n 0.00192977f $X=2.4 $Y=0.495 $X2=0 $Y2=0
cc_184 N_A2_c_217_n N_A_218_57#_c_370_n 0.00346177f $X=2.372 $Y=1.067 $X2=0
+ $Y2=0
cc_185 N_A2_M1009_g N_A_218_57#_c_370_n 0.008695f $X=2.4 $Y=0.495 $X2=0 $Y2=0
cc_186 A2 N_A_218_57#_c_370_n 0.0352532f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_187 N_A2_c_222_n N_A_218_57#_c_370_n 7.78583e-19 $X=2.435 $Y=1.375 $X2=0
+ $Y2=0
cc_188 N_A2_c_217_n N_A_218_57#_c_372_n 0.00193317f $X=2.372 $Y=1.067 $X2=0
+ $Y2=0
cc_189 A2 N_A_218_57#_c_372_n 0.00329776f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_190 N_A2_M1009_g N_VGND_c_412_n 0.00192154f $X=2.4 $Y=0.495 $X2=0 $Y2=0
cc_191 N_A2_M1009_g N_VGND_c_414_n 0.0053602f $X=2.4 $Y=0.495 $X2=0 $Y2=0
cc_192 N_A2_M1009_g N_VGND_c_416_n 0.00582181f $X=2.4 $Y=0.495 $X2=0 $Y2=0
cc_193 N_A1_M1008_g N_VPWR_c_299_n 0.0235506f $X=2.705 $Y=2.735 $X2=0 $Y2=0
cc_194 N_A1_c_270_n N_VPWR_c_299_n 0.00789145f $X=2.885 $Y=2.195 $X2=0 $Y2=0
cc_195 N_A1_c_271_n N_VPWR_c_299_n 5.1063e-19 $X=3.032 $Y=1.88 $X2=0 $Y2=0
cc_196 A1 N_VPWR_c_299_n 0.0131227f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_197 N_A1_M1008_g N_VPWR_c_301_n 0.00289303f $X=2.705 $Y=2.735 $X2=0 $Y2=0
cc_198 N_A1_M1008_g N_VPWR_c_297_n 0.00528764f $X=2.705 $Y=2.735 $X2=0 $Y2=0
cc_199 N_A1_M1005_g N_A_218_57#_c_370_n 0.0167922f $X=2.885 $Y=0.495 $X2=0 $Y2=0
cc_200 A1 N_A_218_57#_c_370_n 0.0317644f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_201 N_A1_c_267_n N_A_218_57#_c_370_n 0.00204946f $X=3 $Y=1.375 $X2=0 $Y2=0
cc_202 N_A1_M1005_g N_A_218_57#_c_371_n 0.00414679f $X=2.885 $Y=0.495 $X2=0
+ $Y2=0
cc_203 N_A1_M1005_g N_VGND_c_412_n 0.00342029f $X=2.885 $Y=0.495 $X2=0 $Y2=0
cc_204 N_A1_M1005_g N_VGND_c_415_n 0.0053602f $X=2.885 $Y=0.495 $X2=0 $Y2=0
cc_205 N_A1_M1005_g N_VGND_c_416_n 0.00646358f $X=2.885 $Y=0.495 $X2=0 $Y2=0
cc_206 N_VPWR_c_298_n N_Y_c_333_n 0.0227326f $X=0.735 $Y=2.57 $X2=0 $Y2=0
cc_207 N_VPWR_c_298_n N_Y_c_334_n 0.00147252f $X=0.735 $Y=2.57 $X2=0 $Y2=0
cc_208 N_VPWR_c_301_n N_Y_c_334_n 0.0200094f $X=2.71 $Y=3.33 $X2=0 $Y2=0
cc_209 N_VPWR_c_297_n N_Y_c_334_n 0.01142f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_210 Y N_VGND_c_413_n 0.0236302f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_211 N_Y_c_332_n N_VGND_c_413_n 0.0160774f $X=0.257 $Y=0.645 $X2=0 $Y2=0
cc_212 Y N_VGND_c_416_n 0.0189764f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_213 N_Y_c_332_n N_VGND_c_416_n 0.011873f $X=0.257 $Y=0.645 $X2=0 $Y2=0
cc_214 N_A_218_57#_c_367_n N_VGND_c_411_n 0.0234856f $X=2.04 $Y=0.915 $X2=0
+ $Y2=0
cc_215 N_A_218_57#_c_370_n N_VGND_c_412_n 0.0213314f $X=2.97 $Y=0.915 $X2=0
+ $Y2=0
cc_216 N_A_218_57#_c_366_n N_VGND_c_413_n 0.0103639f $X=1.23 $Y=0.495 $X2=0
+ $Y2=0
cc_217 N_A_218_57#_c_369_n N_VGND_c_414_n 0.0104258f $X=2.185 $Y=0.495 $X2=0
+ $Y2=0
cc_218 N_A_218_57#_c_371_n N_VGND_c_415_n 0.0128504f $X=3.1 $Y=0.495 $X2=0 $Y2=0
cc_219 N_A_218_57#_c_366_n N_VGND_c_416_n 0.0100107f $X=1.23 $Y=0.495 $X2=0
+ $Y2=0
cc_220 N_A_218_57#_c_367_n N_VGND_c_416_n 0.0108458f $X=2.04 $Y=0.915 $X2=0
+ $Y2=0
cc_221 N_A_218_57#_c_369_n N_VGND_c_416_n 0.00997979f $X=2.185 $Y=0.495 $X2=0
+ $Y2=0
cc_222 N_A_218_57#_c_370_n N_VGND_c_416_n 0.0107705f $X=2.97 $Y=0.915 $X2=0
+ $Y2=0
cc_223 N_A_218_57#_c_371_n N_VGND_c_416_n 0.0109445f $X=3.1 $Y=0.495 $X2=0 $Y2=0
