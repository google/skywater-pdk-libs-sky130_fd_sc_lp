* NGSPICE file created from sky130_fd_sc_lp__iso1n_lp2.ext - technology: sky130A

.subckt sky130_fd_sc_lp__iso1n_lp2 A SLEEP_B KAGND VGND VNB VPB VPWR X
M1000 VPWR SLEEP_B a_27_109# VPB phighvt w=1e+06u l=250000u
+  ad=6.05e+11p pd=5.21e+06u as=2.85e+11p ps=2.57e+06u
M1001 a_114_109# SLEEP_B a_27_109# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=1.197e+11p ps=1.41e+06u
M1002 a_350_109# A a_300_409# VPB phighvt w=1e+06u l=250000u
+  ad=2.85e+11p pd=2.57e+06u as=2.4e+11p ps=2.48e+06u
M1003 X a_350_109# VPWR VPB phighvt w=1e+06u l=250000u
+  ad=2.85e+11p pd=2.57e+06u as=0p ps=0u
M1004 a_350_109# a_27_109# a_272_109# VNB nshort w=420000u l=150000u
+  ad=1.512e+11p pd=1.56e+06u as=1.008e+11p ps=1.32e+06u
M1005 X a_350_109# a_610_109# VNB nshort w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=8.82e+10p ps=1.26e+06u
M1006 KAGND SLEEP_B a_114_109# VNB nshort w=420000u l=150000u
+  ad=2.352e+11p pd=2.8e+06u as=0p ps=0u
M1007 a_300_409# a_27_109# VPWR VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_272_109# a_27_109# KAGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 KAGND A a_452_109# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1010 a_610_109# a_350_109# KAGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_452_109# A a_350_109# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

