* File: sky130_fd_sc_lp__a2bb2o_4.pxi.spice
* Created: Fri Aug 28 09:56:00 2020
* 
x_PM_SKY130_FD_SC_LP__A2BB2O_4%B1 N_B1_M1002_g N_B1_M1011_g N_B1_M1007_g
+ N_B1_M1017_g N_B1_c_130_n N_B1_c_131_n N_B1_c_138_n N_B1_c_132_n N_B1_c_133_n
+ N_B1_c_134_n N_B1_c_143_p B1 B1 PM_SKY130_FD_SC_LP__A2BB2O_4%B1
x_PM_SKY130_FD_SC_LP__A2BB2O_4%B2 N_B2_M1005_g N_B2_M1019_g N_B2_M1021_g
+ N_B2_M1026_g B2 N_B2_c_215_n N_B2_c_212_n PM_SKY130_FD_SC_LP__A2BB2O_4%B2
x_PM_SKY130_FD_SC_LP__A2BB2O_4%A_436_21# N_A_436_21#_M1024_s N_A_436_21#_M1027_d
+ N_A_436_21#_M1000_s N_A_436_21#_M1001_g N_A_436_21#_M1003_g
+ N_A_436_21#_c_262_n N_A_436_21#_M1013_g N_A_436_21#_M1020_g
+ N_A_436_21#_c_265_n N_A_436_21#_c_266_n N_A_436_21#_c_278_p
+ N_A_436_21#_c_352_p N_A_436_21#_c_270_n N_A_436_21#_c_319_p
+ N_A_436_21#_c_300_p N_A_436_21#_c_286_p N_A_436_21#_c_293_p
+ N_A_436_21#_c_299_p N_A_436_21#_c_294_p N_A_436_21#_c_271_n
+ PM_SKY130_FD_SC_LP__A2BB2O_4%A_436_21#
x_PM_SKY130_FD_SC_LP__A2BB2O_4%A1_N N_A1_N_c_377_n N_A1_N_M1024_g N_A1_N_c_378_n
+ N_A1_N_M1004_g N_A1_N_M1025_g N_A1_N_M1018_g N_A1_N_c_380_n A1_N
+ N_A1_N_c_382_n N_A1_N_c_383_n N_A1_N_c_384_n PM_SKY130_FD_SC_LP__A2BB2O_4%A1_N
x_PM_SKY130_FD_SC_LP__A2BB2O_4%A2_N N_A2_N_c_459_n N_A2_N_M1010_g N_A2_N_M1000_g
+ N_A2_N_c_460_n N_A2_N_M1027_g N_A2_N_M1012_g A2_N N_A2_N_c_464_n
+ N_A2_N_c_461_n PM_SKY130_FD_SC_LP__A2BB2O_4%A2_N
x_PM_SKY130_FD_SC_LP__A2BB2O_4%A_200_47# N_A_200_47#_M1005_d N_A_200_47#_M1001_d
+ N_A_200_47#_M1003_d N_A_200_47#_M1006_g N_A_200_47#_M1009_g
+ N_A_200_47#_M1008_g N_A_200_47#_M1016_g N_A_200_47#_M1014_g
+ N_A_200_47#_M1022_g N_A_200_47#_M1015_g N_A_200_47#_M1023_g
+ N_A_200_47#_c_665_p N_A_200_47#_c_516_n N_A_200_47#_c_517_n
+ N_A_200_47#_c_518_n N_A_200_47#_c_582_p N_A_200_47#_c_655_p
+ N_A_200_47#_c_528_n N_A_200_47#_c_555_n N_A_200_47#_c_519_n
+ N_A_200_47#_c_520_n N_A_200_47#_c_616_p N_A_200_47#_c_521_n
+ N_A_200_47#_c_530_n N_A_200_47#_c_522_n PM_SKY130_FD_SC_LP__A2BB2O_4%A_200_47#
x_PM_SKY130_FD_SC_LP__A2BB2O_4%A_27_367# N_A_27_367#_M1011_d N_A_27_367#_M1019_s
+ N_A_27_367#_M1017_d N_A_27_367#_M1020_s N_A_27_367#_c_669_n
+ N_A_27_367#_c_679_n N_A_27_367#_c_720_p N_A_27_367#_c_683_n
+ N_A_27_367#_c_670_n N_A_27_367#_c_671_n N_A_27_367#_c_718_p
+ N_A_27_367#_c_672_n N_A_27_367#_c_673_n N_A_27_367#_c_691_n
+ PM_SKY130_FD_SC_LP__A2BB2O_4%A_27_367#
x_PM_SKY130_FD_SC_LP__A2BB2O_4%VPWR N_VPWR_M1011_s N_VPWR_M1026_d N_VPWR_M1004_s
+ N_VPWR_M1018_s N_VPWR_M1016_d N_VPWR_M1023_d N_VPWR_c_730_n N_VPWR_c_731_n
+ N_VPWR_c_732_n N_VPWR_c_733_n N_VPWR_c_734_n N_VPWR_c_735_n N_VPWR_c_736_n
+ N_VPWR_c_737_n N_VPWR_c_738_n VPWR N_VPWR_c_739_n N_VPWR_c_740_n
+ N_VPWR_c_741_n N_VPWR_c_742_n N_VPWR_c_743_n N_VPWR_c_744_n N_VPWR_c_745_n
+ N_VPWR_c_746_n N_VPWR_c_747_n N_VPWR_c_729_n PM_SKY130_FD_SC_LP__A2BB2O_4%VPWR
x_PM_SKY130_FD_SC_LP__A2BB2O_4%A_742_367# N_A_742_367#_M1004_d
+ N_A_742_367#_M1012_d N_A_742_367#_c_844_n
+ PM_SKY130_FD_SC_LP__A2BB2O_4%A_742_367#
x_PM_SKY130_FD_SC_LP__A2BB2O_4%X N_X_M1006_d N_X_M1014_d N_X_M1009_s N_X_M1022_s
+ N_X_c_909_p N_X_c_895_n N_X_c_854_n N_X_c_855_n N_X_c_860_n N_X_c_861_n
+ N_X_c_910_p N_X_c_899_n N_X_c_862_n N_X_c_856_n N_X_c_863_n X X N_X_c_858_n X
+ PM_SKY130_FD_SC_LP__A2BB2O_4%X
x_PM_SKY130_FD_SC_LP__A2BB2O_4%VGND N_VGND_M1002_d N_VGND_M1007_d N_VGND_M1013_s
+ N_VGND_M1010_s N_VGND_M1025_d N_VGND_M1008_s N_VGND_M1015_s N_VGND_c_915_n
+ N_VGND_c_916_n N_VGND_c_917_n N_VGND_c_918_n N_VGND_c_919_n N_VGND_c_920_n
+ N_VGND_c_921_n N_VGND_c_922_n N_VGND_c_923_n N_VGND_c_924_n N_VGND_c_925_n
+ N_VGND_c_926_n VGND N_VGND_c_927_n N_VGND_c_928_n N_VGND_c_929_n
+ N_VGND_c_930_n N_VGND_c_931_n N_VGND_c_932_n N_VGND_c_933_n N_VGND_c_934_n
+ PM_SKY130_FD_SC_LP__A2BB2O_4%VGND
x_PM_SKY130_FD_SC_LP__A2BB2O_4%A_114_47# N_A_114_47#_M1002_s N_A_114_47#_M1021_s
+ N_A_114_47#_c_1038_n N_A_114_47#_c_1034_n N_A_114_47#_c_1037_n
+ PM_SKY130_FD_SC_LP__A2BB2O_4%A_114_47#
cc_1 VNB N_B1_M1002_g 0.0349147f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.655
cc_2 VNB N_B1_M1007_g 0.0240558f $X=-0.19 $Y=-0.245 $X2=1.785 $Y2=0.655
cc_3 VNB N_B1_c_130_n 0.0152673f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=1.495
cc_4 VNB N_B1_c_131_n 0.0291717f $X=-0.19 $Y=-0.245 $X2=0.405 $Y2=1.51
cc_5 VNB N_B1_c_132_n 0.00299491f $X=-0.19 $Y=-0.245 $X2=1.635 $Y2=1.525
cc_6 VNB N_B1_c_133_n 0.00195814f $X=-0.19 $Y=-0.245 $X2=1.805 $Y2=1.51
cc_7 VNB N_B1_c_134_n 0.0223882f $X=-0.19 $Y=-0.245 $X2=1.805 $Y2=1.51
cc_8 VNB N_B2_M1005_g 0.0247747f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.655
cc_9 VNB N_B2_M1021_g 0.0232219f $X=-0.19 $Y=-0.245 $X2=1.785 $Y2=0.655
cc_10 VNB N_B2_c_212_n 0.0327253f $X=-0.19 $Y=-0.245 $X2=1.635 $Y2=1.525
cc_11 VNB N_A_436_21#_M1001_g 0.0197753f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_436_21#_M1003_g 0.0112741f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_436_21#_c_262_n 0.0472035f $X=-0.19 $Y=-0.245 $X2=0.405 $Y2=1.495
cc_14 VNB N_A_436_21#_M1013_g 0.0225024f $X=-0.19 $Y=-0.245 $X2=1.55 $Y2=1.645
cc_15 VNB N_A_436_21#_M1020_g 0.00276207f $X=-0.19 $Y=-0.245 $X2=1.805 $Y2=1.51
cc_16 VNB N_A_436_21#_c_265_n 0.00526723f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_436_21#_c_266_n 0.00232864f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A1_N_c_377_n 0.0173944f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.345
cc_19 VNB N_A1_N_c_378_n 0.048482f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A1_N_M1018_g 0.00781993f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A1_N_c_380_n 0.00120674f $X=-0.19 $Y=-0.245 $X2=1.825 $Y2=2.465
cc_22 VNB A1_N 0.00447847f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A1_N_c_382_n 0.0350204f $X=-0.19 $Y=-0.245 $X2=1.805 $Y2=1.51
cc_24 VNB N_A1_N_c_383_n 0.00933661f $X=-0.19 $Y=-0.245 $X2=1.805 $Y2=1.51
cc_25 VNB N_A1_N_c_384_n 0.0159135f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A2_N_c_459_n 0.0166528f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.345
cc_27 VNB N_A2_N_c_460_n 0.0166049f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A2_N_c_461_n 0.0610616f $X=-0.19 $Y=-0.245 $X2=1.55 $Y2=1.645
cc_29 VNB N_A_200_47#_M1006_g 0.0238557f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_200_47#_M1008_g 0.0217542f $X=-0.19 $Y=-0.245 $X2=0.405 $Y2=1.51
cc_31 VNB N_A_200_47#_M1014_g 0.0217342f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_200_47#_M1015_g 0.0265185f $X=-0.19 $Y=-0.245 $X2=0.405 $Y2=1.345
cc_33 VNB N_A_200_47#_c_516_n 0.00813562f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.95
cc_34 VNB N_A_200_47#_c_517_n 0.00370848f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=2.035
cc_35 VNB N_A_200_47#_c_518_n 0.00414742f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_200_47#_c_519_n 6.81766e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_200_47#_c_520_n 0.00355088f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_200_47#_c_521_n 0.00101212f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_200_47#_c_522_n 0.0729434f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_VPWR_c_729_n 0.302998f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_X_c_854_n 0.00304538f $X=-0.19 $Y=-0.245 $X2=1.55 $Y2=1.95
cc_42 VNB N_X_c_855_n 0.00365065f $X=-0.19 $Y=-0.245 $X2=1.635 $Y2=1.525
cc_43 VNB N_X_c_856_n 0.00144145f $X=-0.19 $Y=-0.245 $X2=1.805 $Y2=1.675
cc_44 VNB X 0.00169133f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=2.035
cc_45 VNB N_X_c_858_n 0.00754504f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB X 0.0195569f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_915_n 0.0113512f $X=-0.19 $Y=-0.245 $X2=1.55 $Y2=1.645
cc_48 VNB N_VGND_c_916_n 0.044354f $X=-0.19 $Y=-0.245 $X2=1.635 $Y2=1.525
cc_49 VNB N_VGND_c_917_n 0.00252888f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_918_n 0.0144243f $X=-0.19 $Y=-0.245 $X2=1.465 $Y2=2.035
cc_51 VNB N_VGND_c_919_n 0.00501912f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_920_n 0.0175865f $X=-0.19 $Y=-0.245 $X2=0.405 $Y2=1.345
cc_53 VNB N_VGND_c_921_n 0.0046469f $X=-0.19 $Y=-0.245 $X2=1.805 $Y2=1.675
cc_54 VNB N_VGND_c_922_n 3.16049e-19 $X=-0.19 $Y=-0.245 $X2=0.76 $Y2=2.035
cc_55 VNB N_VGND_c_923_n 0.0116416f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.95
cc_56 VNB N_VGND_c_924_n 0.0283468f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_VGND_c_925_n 0.0364888f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_926_n 0.00428723f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_927_n 0.0148832f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_928_n 0.0129398f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_929_n 0.0134763f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_930_n 0.0122171f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_VGND_c_931_n 0.00631953f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_VGND_c_932_n 0.0053824f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_VGND_c_933_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_VGND_c_934_n 0.349497f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_A_114_47#_c_1034_n 0.0074378f $X=-0.19 $Y=-0.245 $X2=1.825 $Y2=2.465
cc_68 VPB N_B1_M1011_g 0.0247289f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=2.465
cc_69 VPB N_B1_M1017_g 0.0195082f $X=-0.19 $Y=1.655 $X2=1.825 $Y2=2.465
cc_70 VPB N_B1_c_131_n 0.00665934f $X=-0.19 $Y=1.655 $X2=0.405 $Y2=1.51
cc_71 VPB N_B1_c_138_n 0.00284273f $X=-0.19 $Y=1.655 $X2=1.55 $Y2=1.95
cc_72 VPB N_B1_c_134_n 0.00707107f $X=-0.19 $Y=1.655 $X2=1.805 $Y2=1.51
cc_73 VPB B1 0.00126936f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.95
cc_74 VPB N_B2_M1019_g 0.0183444f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=2.465
cc_75 VPB N_B2_M1026_g 0.0187559f $X=-0.19 $Y=1.655 $X2=1.825 $Y2=2.465
cc_76 VPB N_B2_c_215_n 0.00260271f $X=-0.19 $Y=1.655 $X2=1.55 $Y2=1.95
cc_77 VPB N_B2_c_212_n 0.00481806f $X=-0.19 $Y=1.655 $X2=1.635 $Y2=1.525
cc_78 VPB N_A_436_21#_M1003_g 0.0200488f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_79 VPB N_A_436_21#_M1020_g 0.0239855f $X=-0.19 $Y=1.655 $X2=1.805 $Y2=1.51
cc_80 VPB N_A_436_21#_c_266_n 0.00138787f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_81 VPB N_A_436_21#_c_270_n 0.0158223f $X=-0.19 $Y=1.655 $X2=0.405 $Y2=1.345
cc_82 VPB N_A_436_21#_c_271_n 0.00126554f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_83 VPB N_A1_N_c_378_n 0.0279526f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_84 VPB N_A1_N_M1018_g 0.021214f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_85 VPB N_A2_N_M1000_g 0.0187244f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=2.465
cc_86 VPB N_A2_N_M1012_g 0.0195707f $X=-0.19 $Y=1.655 $X2=1.825 $Y2=1.675
cc_87 VPB N_A2_N_c_464_n 0.00349012f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_88 VPB N_A2_N_c_461_n 0.00452845f $X=-0.19 $Y=1.655 $X2=1.55 $Y2=1.645
cc_89 VPB N_A_200_47#_M1009_g 0.0196748f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_90 VPB N_A_200_47#_M1016_g 0.0189821f $X=-0.19 $Y=1.655 $X2=1.635 $Y2=1.525
cc_91 VPB N_A_200_47#_M1022_g 0.0188421f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_92 VPB N_A_200_47#_M1023_g 0.0232806f $X=-0.19 $Y=1.655 $X2=1.805 $Y2=1.675
cc_93 VPB N_A_200_47#_c_518_n 0.00412335f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_94 VPB N_A_200_47#_c_528_n 0.00981593f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_95 VPB N_A_200_47#_c_519_n 0.00177852f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_96 VPB N_A_200_47#_c_530_n 0.00450654f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_97 VPB N_A_200_47#_c_522_n 0.00744666f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_98 VPB N_A_27_367#_c_669_n 0.0248654f $X=-0.19 $Y=1.655 $X2=1.825 $Y2=2.465
cc_99 VPB N_A_27_367#_c_670_n 0.00383515f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=1.645
cc_100 VPB N_A_27_367#_c_671_n 0.00182139f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_101 VPB N_A_27_367#_c_672_n 0.00557433f $X=-0.19 $Y=1.655 $X2=0.405 $Y2=1.675
cc_102 VPB N_A_27_367#_c_673_n 0.0307716f $X=-0.19 $Y=1.655 $X2=1.805 $Y2=1.675
cc_103 VPB N_VPWR_c_730_n 4.02668e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_104 VPB N_VPWR_c_731_n 4.02668e-19 $X=-0.19 $Y=1.655 $X2=1.805 $Y2=1.525
cc_105 VPB N_VPWR_c_732_n 0.00730073f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=1.645
cc_106 VPB N_VPWR_c_733_n 0.00285717f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_107 VPB N_VPWR_c_734_n 3.19622e-19 $X=-0.19 $Y=1.655 $X2=0.405 $Y2=1.675
cc_108 VPB N_VPWR_c_735_n 0.0111354f $X=-0.19 $Y=1.655 $X2=0.715 $Y2=2.035
cc_109 VPB N_VPWR_c_736_n 0.0444288f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=2.035
cc_110 VPB N_VPWR_c_737_n 0.0357104f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_111 VPB N_VPWR_c_738_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_112 VPB N_VPWR_c_739_n 0.0158241f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_113 VPB N_VPWR_c_740_n 0.0133881f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_114 VPB N_VPWR_c_741_n 0.0356756f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_115 VPB N_VPWR_c_742_n 0.0138945f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_116 VPB N_VPWR_c_743_n 0.0146078f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_117 VPB N_VPWR_c_744_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_118 VPB N_VPWR_c_745_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_119 VPB N_VPWR_c_746_n 0.00522677f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_120 VPB N_VPWR_c_747_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_121 VPB N_VPWR_c_729_n 0.052543f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_122 VPB N_X_c_860_n 0.00304705f $X=-0.19 $Y=1.655 $X2=1.805 $Y2=1.525
cc_123 VPB N_X_c_861_n 0.00199724f $X=-0.19 $Y=1.655 $X2=1.805 $Y2=1.51
cc_124 VPB N_X_c_862_n 0.00461479f $X=-0.19 $Y=1.655 $X2=0.405 $Y2=1.675
cc_125 VPB N_X_c_863_n 0.00172486f $X=-0.19 $Y=1.655 $X2=0.715 $Y2=2.035
cc_126 VPB X 0.00455971f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_127 N_B1_M1002_g N_B2_M1005_g 0.0296196f $X=0.495 $Y=0.655 $X2=0 $Y2=0
cc_128 N_B1_M1011_g N_B2_M1019_g 0.0296196f $X=0.495 $Y=2.465 $X2=0 $Y2=0
cc_129 N_B1_c_143_p N_B2_M1019_g 0.0118001f $X=1.465 $Y=2.035 $X2=0 $Y2=0
cc_130 N_B1_M1007_g N_B2_M1021_g 0.0243644f $X=1.785 $Y=0.655 $X2=0 $Y2=0
cc_131 N_B1_M1017_g N_B2_M1026_g 0.0409027f $X=1.825 $Y=2.465 $X2=0 $Y2=0
cc_132 N_B1_c_143_p N_B2_M1026_g 0.0141918f $X=1.465 $Y=2.035 $X2=0 $Y2=0
cc_133 N_B1_c_130_n N_B2_c_215_n 0.019082f $X=0.545 $Y=1.495 $X2=0 $Y2=0
cc_134 N_B1_c_131_n N_B2_c_215_n 3.51309e-19 $X=0.405 $Y=1.51 $X2=0 $Y2=0
cc_135 N_B1_c_138_n N_B2_c_215_n 0.0102197f $X=1.55 $Y=1.95 $X2=0 $Y2=0
cc_136 N_B1_c_132_n N_B2_c_215_n 0.0200216f $X=1.635 $Y=1.525 $X2=0 $Y2=0
cc_137 N_B1_c_143_p N_B2_c_215_n 0.0265579f $X=1.465 $Y=2.035 $X2=0 $Y2=0
cc_138 B1 N_B2_c_215_n 0.00978927f $X=0.635 $Y=1.95 $X2=0 $Y2=0
cc_139 N_B1_c_130_n N_B2_c_212_n 0.0035905f $X=0.545 $Y=1.495 $X2=0 $Y2=0
cc_140 N_B1_c_131_n N_B2_c_212_n 0.0296196f $X=0.405 $Y=1.51 $X2=0 $Y2=0
cc_141 N_B1_c_138_n N_B2_c_212_n 0.0029626f $X=1.55 $Y=1.95 $X2=0 $Y2=0
cc_142 N_B1_c_132_n N_B2_c_212_n 0.00200312f $X=1.635 $Y=1.525 $X2=0 $Y2=0
cc_143 N_B1_c_134_n N_B2_c_212_n 0.0219175f $X=1.805 $Y=1.51 $X2=0 $Y2=0
cc_144 N_B1_c_143_p N_B2_c_212_n 5.38132e-19 $X=1.465 $Y=2.035 $X2=0 $Y2=0
cc_145 B1 N_B2_c_212_n 0.00450268f $X=0.635 $Y=1.95 $X2=0 $Y2=0
cc_146 N_B1_M1007_g N_A_436_21#_M1001_g 0.0221733f $X=1.785 $Y=0.655 $X2=0 $Y2=0
cc_147 N_B1_M1017_g N_A_436_21#_M1003_g 0.0183316f $X=1.825 $Y=2.465 $X2=0 $Y2=0
cc_148 N_B1_c_133_n N_A_436_21#_c_265_n 8.35289e-19 $X=1.805 $Y=1.51 $X2=0 $Y2=0
cc_149 N_B1_c_134_n N_A_436_21#_c_265_n 0.0207332f $X=1.805 $Y=1.51 $X2=0 $Y2=0
cc_150 N_B1_M1007_g N_A_200_47#_c_516_n 0.0144718f $X=1.785 $Y=0.655 $X2=0 $Y2=0
cc_151 N_B1_c_132_n N_A_200_47#_c_516_n 0.0144183f $X=1.635 $Y=1.525 $X2=0 $Y2=0
cc_152 N_B1_c_133_n N_A_200_47#_c_516_n 0.0239961f $X=1.805 $Y=1.51 $X2=0 $Y2=0
cc_153 N_B1_c_134_n N_A_200_47#_c_516_n 0.00450001f $X=1.805 $Y=1.51 $X2=0 $Y2=0
cc_154 N_B1_M1007_g N_A_200_47#_c_518_n 3.1212e-19 $X=1.785 $Y=0.655 $X2=0 $Y2=0
cc_155 N_B1_c_133_n N_A_200_47#_c_518_n 0.010362f $X=1.805 $Y=1.51 $X2=0 $Y2=0
cc_156 N_B1_c_134_n N_A_200_47#_c_518_n 3.24407e-19 $X=1.805 $Y=1.51 $X2=0 $Y2=0
cc_157 N_B1_c_143_p N_A_27_367#_M1019_s 0.00333507f $X=1.465 $Y=2.035 $X2=0
+ $Y2=0
cc_158 N_B1_M1011_g N_A_27_367#_c_669_n 0.00199721f $X=0.495 $Y=2.465 $X2=0
+ $Y2=0
cc_159 N_B1_c_130_n N_A_27_367#_c_669_n 0.011227f $X=0.545 $Y=1.495 $X2=0 $Y2=0
cc_160 N_B1_c_131_n N_A_27_367#_c_669_n 0.00323663f $X=0.405 $Y=1.51 $X2=0 $Y2=0
cc_161 B1 N_A_27_367#_c_669_n 0.00531237f $X=0.635 $Y=1.95 $X2=0 $Y2=0
cc_162 N_B1_M1011_g N_A_27_367#_c_679_n 0.0140136f $X=0.495 $Y=2.465 $X2=0 $Y2=0
cc_163 N_B1_c_130_n N_A_27_367#_c_679_n 0.00344318f $X=0.545 $Y=1.495 $X2=0
+ $Y2=0
cc_164 N_B1_c_143_p N_A_27_367#_c_679_n 0.0157622f $X=1.465 $Y=2.035 $X2=0 $Y2=0
cc_165 B1 N_A_27_367#_c_679_n 0.00897693f $X=0.635 $Y=1.95 $X2=0 $Y2=0
cc_166 N_B1_M1017_g N_A_27_367#_c_683_n 0.0151765f $X=1.825 $Y=2.465 $X2=0 $Y2=0
cc_167 N_B1_c_133_n N_A_27_367#_c_683_n 0.00597237f $X=1.805 $Y=1.51 $X2=0 $Y2=0
cc_168 N_B1_c_134_n N_A_27_367#_c_683_n 0.00167524f $X=1.805 $Y=1.51 $X2=0 $Y2=0
cc_169 N_B1_c_143_p N_A_27_367#_c_683_n 0.0221786f $X=1.465 $Y=2.035 $X2=0 $Y2=0
cc_170 N_B1_M1017_g N_A_27_367#_c_670_n 5.37707e-19 $X=1.825 $Y=2.465 $X2=0
+ $Y2=0
cc_171 N_B1_c_138_n N_A_27_367#_c_670_n 0.00373893f $X=1.55 $Y=1.95 $X2=0 $Y2=0
cc_172 N_B1_c_133_n N_A_27_367#_c_670_n 0.00280614f $X=1.805 $Y=1.51 $X2=0 $Y2=0
cc_173 N_B1_c_134_n N_A_27_367#_c_670_n 8.21235e-19 $X=1.805 $Y=1.51 $X2=0 $Y2=0
cc_174 N_B1_c_143_p N_A_27_367#_c_691_n 0.0135055f $X=1.465 $Y=2.035 $X2=0 $Y2=0
cc_175 N_B1_c_143_p N_VPWR_M1011_s 0.0037585f $X=1.465 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_176 B1 N_VPWR_M1011_s 0.00225932f $X=0.635 $Y=1.95 $X2=-0.19 $Y2=-0.245
cc_177 N_B1_c_138_n N_VPWR_M1026_d 0.00133236f $X=1.55 $Y=1.95 $X2=0 $Y2=0
cc_178 N_B1_c_143_p N_VPWR_M1026_d 0.00369416f $X=1.465 $Y=2.035 $X2=0 $Y2=0
cc_179 N_B1_M1011_g N_VPWR_c_730_n 0.0121813f $X=0.495 $Y=2.465 $X2=0 $Y2=0
cc_180 N_B1_M1017_g N_VPWR_c_731_n 0.010521f $X=1.825 $Y=2.465 $X2=0 $Y2=0
cc_181 N_B1_M1017_g N_VPWR_c_737_n 0.00564095f $X=1.825 $Y=2.465 $X2=0 $Y2=0
cc_182 N_B1_M1011_g N_VPWR_c_739_n 0.00486043f $X=0.495 $Y=2.465 $X2=0 $Y2=0
cc_183 N_B1_M1011_g N_VPWR_c_729_n 0.00919827f $X=0.495 $Y=2.465 $X2=0 $Y2=0
cc_184 N_B1_M1017_g N_VPWR_c_729_n 0.00950825f $X=1.825 $Y=2.465 $X2=0 $Y2=0
cc_185 N_B1_M1002_g N_VGND_c_916_n 0.00847481f $X=0.495 $Y=0.655 $X2=0 $Y2=0
cc_186 N_B1_c_130_n N_VGND_c_916_n 0.00999271f $X=0.545 $Y=1.495 $X2=0 $Y2=0
cc_187 N_B1_c_131_n N_VGND_c_916_n 0.00354571f $X=0.405 $Y=1.51 $X2=0 $Y2=0
cc_188 N_B1_M1007_g N_VGND_c_917_n 0.00297689f $X=1.785 $Y=0.655 $X2=0 $Y2=0
cc_189 N_B1_M1002_g N_VGND_c_925_n 0.00585385f $X=0.495 $Y=0.655 $X2=0 $Y2=0
cc_190 N_B1_M1007_g N_VGND_c_925_n 0.00547432f $X=1.785 $Y=0.655 $X2=0 $Y2=0
cc_191 N_B1_M1002_g N_VGND_c_934_n 0.0115261f $X=0.495 $Y=0.655 $X2=0 $Y2=0
cc_192 N_B1_M1007_g N_VGND_c_934_n 0.009873f $X=1.785 $Y=0.655 $X2=0 $Y2=0
cc_193 N_B1_M1002_g N_A_114_47#_c_1034_n 7.23352e-19 $X=0.495 $Y=0.655 $X2=0
+ $Y2=0
cc_194 N_B1_c_130_n N_A_114_47#_c_1034_n 0.0102844f $X=0.545 $Y=1.495 $X2=0
+ $Y2=0
cc_195 N_B1_M1007_g N_A_114_47#_c_1037_n 0.00709582f $X=1.785 $Y=0.655 $X2=0
+ $Y2=0
cc_196 N_B2_M1021_g N_A_200_47#_c_516_n 0.0160282f $X=1.355 $Y=0.655 $X2=0 $Y2=0
cc_197 N_B2_c_215_n N_A_200_47#_c_516_n 0.00441038f $X=1.06 $Y=1.51 $X2=0 $Y2=0
cc_198 N_B2_M1005_g N_A_200_47#_c_517_n 0.00484133f $X=0.925 $Y=0.655 $X2=0
+ $Y2=0
cc_199 N_B2_c_215_n N_A_200_47#_c_517_n 0.0182913f $X=1.06 $Y=1.51 $X2=0 $Y2=0
cc_200 N_B2_c_212_n N_A_200_47#_c_517_n 0.00249434f $X=1.355 $Y=1.51 $X2=0 $Y2=0
cc_201 N_B2_M1019_g N_A_27_367#_c_679_n 0.0122129f $X=0.925 $Y=2.465 $X2=0 $Y2=0
cc_202 N_B2_M1026_g N_A_27_367#_c_683_n 0.0129951f $X=1.355 $Y=2.465 $X2=0 $Y2=0
cc_203 N_B2_M1019_g N_VPWR_c_730_n 0.0105405f $X=0.925 $Y=2.465 $X2=0 $Y2=0
cc_204 N_B2_M1026_g N_VPWR_c_730_n 5.8398e-19 $X=1.355 $Y=2.465 $X2=0 $Y2=0
cc_205 N_B2_M1019_g N_VPWR_c_731_n 5.5535e-19 $X=0.925 $Y=2.465 $X2=0 $Y2=0
cc_206 N_B2_M1026_g N_VPWR_c_731_n 0.0093124f $X=1.355 $Y=2.465 $X2=0 $Y2=0
cc_207 N_B2_M1019_g N_VPWR_c_740_n 0.00486043f $X=0.925 $Y=2.465 $X2=0 $Y2=0
cc_208 N_B2_M1026_g N_VPWR_c_740_n 0.00564095f $X=1.355 $Y=2.465 $X2=0 $Y2=0
cc_209 N_B2_M1019_g N_VPWR_c_729_n 0.00824727f $X=0.925 $Y=2.465 $X2=0 $Y2=0
cc_210 N_B2_M1026_g N_VPWR_c_729_n 0.00948291f $X=1.355 $Y=2.465 $X2=0 $Y2=0
cc_211 N_B2_M1005_g N_VGND_c_925_n 0.00357877f $X=0.925 $Y=0.655 $X2=0 $Y2=0
cc_212 N_B2_M1021_g N_VGND_c_925_n 0.00357842f $X=1.355 $Y=0.655 $X2=0 $Y2=0
cc_213 N_B2_M1005_g N_VGND_c_934_n 0.00537654f $X=0.925 $Y=0.655 $X2=0 $Y2=0
cc_214 N_B2_M1021_g N_VGND_c_934_n 0.00537652f $X=1.355 $Y=0.655 $X2=0 $Y2=0
cc_215 N_B2_M1005_g N_A_114_47#_c_1038_n 0.012237f $X=0.925 $Y=0.655 $X2=0 $Y2=0
cc_216 N_B2_M1021_g N_A_114_47#_c_1038_n 0.00848835f $X=1.355 $Y=0.655 $X2=0
+ $Y2=0
cc_217 N_B2_M1005_g N_A_114_47#_c_1034_n 7.22995e-19 $X=0.925 $Y=0.655 $X2=0
+ $Y2=0
cc_218 N_B2_M1005_g N_A_114_47#_c_1037_n 5.24903e-19 $X=0.925 $Y=0.655 $X2=0
+ $Y2=0
cc_219 N_B2_M1021_g N_A_114_47#_c_1037_n 0.00702123f $X=1.355 $Y=0.655 $X2=0
+ $Y2=0
cc_220 N_A_436_21#_M1013_g N_A1_N_c_377_n 0.00989062f $X=2.685 $Y=0.655
+ $X2=-0.19 $Y2=-0.245
cc_221 N_A_436_21#_c_266_n N_A1_N_c_377_n 0.00321725f $X=2.84 $Y=1.44 $X2=-0.19
+ $Y2=-0.245
cc_222 N_A_436_21#_c_278_p N_A1_N_c_377_n 0.0111658f $X=3.575 $Y=0.81 $X2=-0.19
+ $Y2=-0.245
cc_223 N_A_436_21#_c_262_n N_A1_N_c_378_n 0.0167346f $X=2.61 $Y=1.35 $X2=0 $Y2=0
cc_224 N_A_436_21#_M1013_g N_A1_N_c_378_n 0.0017845f $X=2.685 $Y=0.655 $X2=0
+ $Y2=0
cc_225 N_A_436_21#_M1020_g N_A1_N_c_378_n 0.0014393f $X=2.685 $Y=2.465 $X2=0
+ $Y2=0
cc_226 N_A_436_21#_c_266_n N_A1_N_c_378_n 0.00489186f $X=2.84 $Y=1.44 $X2=0
+ $Y2=0
cc_227 N_A_436_21#_c_278_p N_A1_N_c_378_n 5.9866e-19 $X=3.575 $Y=0.81 $X2=0
+ $Y2=0
cc_228 N_A_436_21#_c_270_n N_A1_N_c_378_n 0.013952f $X=3.575 $Y=1.845 $X2=0
+ $Y2=0
cc_229 N_A_436_21#_c_271_n N_A1_N_c_378_n 0.0177016f $X=3.66 $Y=1.845 $X2=0
+ $Y2=0
cc_230 N_A_436_21#_c_286_p N_A1_N_M1018_g 0.00100552f $X=4.28 $Y=2.035 $X2=0
+ $Y2=0
cc_231 N_A_436_21#_c_262_n N_A1_N_c_380_n 7.09263e-19 $X=2.61 $Y=1.35 $X2=0
+ $Y2=0
cc_232 N_A_436_21#_M1013_g N_A1_N_c_380_n 4.86476e-19 $X=2.685 $Y=0.655 $X2=0
+ $Y2=0
cc_233 N_A_436_21#_c_266_n N_A1_N_c_380_n 0.0172135f $X=2.84 $Y=1.44 $X2=0 $Y2=0
cc_234 N_A_436_21#_c_278_p N_A1_N_c_380_n 0.0167996f $X=3.575 $Y=0.81 $X2=0
+ $Y2=0
cc_235 N_A_436_21#_c_270_n N_A1_N_c_380_n 0.0153096f $X=3.575 $Y=1.845 $X2=0
+ $Y2=0
cc_236 N_A_436_21#_M1024_s A1_N 0.00181776f $X=3.53 $Y=0.235 $X2=0 $Y2=0
cc_237 N_A_436_21#_c_293_p A1_N 0.0407703f $X=4.525 $Y=0.81 $X2=0 $Y2=0
cc_238 N_A_436_21#_c_294_p A1_N 0.015318f $X=3.705 $Y=0.81 $X2=0 $Y2=0
cc_239 N_A_436_21#_c_271_n A1_N 0.00560381f $X=3.66 $Y=1.845 $X2=0 $Y2=0
cc_240 N_A_436_21#_M1027_d N_A1_N_c_383_n 0.00181822f $X=4.55 $Y=0.235 $X2=0
+ $Y2=0
cc_241 N_A_436_21#_c_293_p N_A1_N_c_383_n 0.0183678f $X=4.525 $Y=0.81 $X2=0
+ $Y2=0
cc_242 N_A_436_21#_c_293_p N_A1_N_c_384_n 0.00210681f $X=4.525 $Y=0.81 $X2=0
+ $Y2=0
cc_243 N_A_436_21#_c_299_p N_A1_N_c_384_n 0.00498229f $X=4.69 $Y=0.42 $X2=0
+ $Y2=0
cc_244 N_A_436_21#_c_300_p N_A2_N_c_459_n 0.00655392f $X=3.67 $Y=0.42 $X2=-0.19
+ $Y2=-0.245
cc_245 N_A_436_21#_c_293_p N_A2_N_c_459_n 0.0098613f $X=4.525 $Y=0.81 $X2=-0.19
+ $Y2=-0.245
cc_246 N_A_436_21#_c_299_p N_A2_N_c_459_n 8.28349e-19 $X=4.69 $Y=0.42 $X2=-0.19
+ $Y2=-0.245
cc_247 N_A_436_21#_c_294_p N_A2_N_c_459_n 5.64397e-19 $X=3.705 $Y=0.81 $X2=-0.19
+ $Y2=-0.245
cc_248 N_A_436_21#_c_286_p N_A2_N_M1000_g 0.0090575f $X=4.28 $Y=2.035 $X2=0
+ $Y2=0
cc_249 N_A_436_21#_c_271_n N_A2_N_M1000_g 0.00167837f $X=3.66 $Y=1.845 $X2=0
+ $Y2=0
cc_250 N_A_436_21#_c_300_p N_A2_N_c_460_n 8.23834e-19 $X=3.67 $Y=0.42 $X2=0
+ $Y2=0
cc_251 N_A_436_21#_c_293_p N_A2_N_c_460_n 0.0103039f $X=4.525 $Y=0.81 $X2=0
+ $Y2=0
cc_252 N_A_436_21#_c_299_p N_A2_N_c_460_n 0.00684735f $X=4.69 $Y=0.42 $X2=0
+ $Y2=0
cc_253 N_A_436_21#_c_286_p N_A2_N_M1012_g 0.00554425f $X=4.28 $Y=2.035 $X2=0
+ $Y2=0
cc_254 N_A_436_21#_c_286_p N_A2_N_c_464_n 0.0210909f $X=4.28 $Y=2.035 $X2=0
+ $Y2=0
cc_255 N_A_436_21#_c_286_p N_A2_N_c_461_n 0.00542252f $X=4.28 $Y=2.035 $X2=0
+ $Y2=0
cc_256 N_A_436_21#_c_293_p N_A2_N_c_461_n 0.00131493f $X=4.525 $Y=0.81 $X2=0
+ $Y2=0
cc_257 N_A_436_21#_M1001_g N_A_200_47#_c_516_n 0.0188923f $X=2.255 $Y=0.655
+ $X2=0 $Y2=0
cc_258 N_A_436_21#_M1001_g N_A_200_47#_c_518_n 0.00102875f $X=2.255 $Y=0.655
+ $X2=0 $Y2=0
cc_259 N_A_436_21#_M1003_g N_A_200_47#_c_518_n 0.00706582f $X=2.255 $Y=2.465
+ $X2=0 $Y2=0
cc_260 N_A_436_21#_c_262_n N_A_200_47#_c_518_n 0.0156941f $X=2.61 $Y=1.35 $X2=0
+ $Y2=0
cc_261 N_A_436_21#_M1013_g N_A_200_47#_c_518_n 2.97573e-19 $X=2.685 $Y=0.655
+ $X2=0 $Y2=0
cc_262 N_A_436_21#_c_266_n N_A_200_47#_c_518_n 0.0345503f $X=2.84 $Y=1.44 $X2=0
+ $Y2=0
cc_263 N_A_436_21#_c_319_p N_A_200_47#_c_518_n 0.00923414f $X=2.925 $Y=1.845
+ $X2=0 $Y2=0
cc_264 N_A_436_21#_c_262_n N_A_200_47#_c_528_n 6.16877e-19 $X=2.61 $Y=1.35 $X2=0
+ $Y2=0
cc_265 N_A_436_21#_M1020_g N_A_200_47#_c_528_n 0.0171888f $X=2.685 $Y=2.465
+ $X2=0 $Y2=0
cc_266 N_A_436_21#_c_270_n N_A_200_47#_c_528_n 0.0230402f $X=3.575 $Y=1.845
+ $X2=0 $Y2=0
cc_267 N_A_436_21#_c_319_p N_A_200_47#_c_528_n 0.00912547f $X=2.925 $Y=1.845
+ $X2=0 $Y2=0
cc_268 N_A_436_21#_M1000_s N_A_200_47#_c_555_n 0.0035168f $X=4.14 $Y=1.835 $X2=0
+ $Y2=0
cc_269 N_A_436_21#_c_270_n N_A_200_47#_c_555_n 0.00447181f $X=3.575 $Y=1.845
+ $X2=0 $Y2=0
cc_270 N_A_436_21#_c_286_p N_A_200_47#_c_555_n 0.0364898f $X=4.28 $Y=2.035 $X2=0
+ $Y2=0
cc_271 N_A_436_21#_c_271_n N_A_200_47#_c_555_n 0.00972913f $X=3.66 $Y=1.845
+ $X2=0 $Y2=0
cc_272 N_A_436_21#_M1013_g N_A_200_47#_c_521_n 0.00138311f $X=2.685 $Y=0.655
+ $X2=0 $Y2=0
cc_273 N_A_436_21#_c_266_n N_A_200_47#_c_521_n 0.0121426f $X=2.84 $Y=1.44 $X2=0
+ $Y2=0
cc_274 N_A_436_21#_M1020_g N_A_200_47#_c_530_n 0.00200817f $X=2.685 $Y=2.465
+ $X2=0 $Y2=0
cc_275 N_A_436_21#_c_270_n N_A_200_47#_c_530_n 0.0132161f $X=3.575 $Y=1.845
+ $X2=0 $Y2=0
cc_276 N_A_436_21#_c_271_n N_A_200_47#_c_530_n 0.0028082f $X=3.66 $Y=1.845 $X2=0
+ $Y2=0
cc_277 N_A_436_21#_c_270_n N_A_27_367#_M1020_s 0.0014972f $X=3.575 $Y=1.845
+ $X2=0 $Y2=0
cc_278 N_A_436_21#_c_319_p N_A_27_367#_M1020_s 0.00119809f $X=2.925 $Y=1.845
+ $X2=0 $Y2=0
cc_279 N_A_436_21#_M1003_g N_A_27_367#_c_670_n 5.31076e-19 $X=2.255 $Y=2.465
+ $X2=0 $Y2=0
cc_280 N_A_436_21#_M1003_g N_A_27_367#_c_671_n 0.012237f $X=2.255 $Y=2.465 $X2=0
+ $Y2=0
cc_281 N_A_436_21#_M1020_g N_A_27_367#_c_671_n 0.00902986f $X=2.685 $Y=2.465
+ $X2=0 $Y2=0
cc_282 N_A_436_21#_M1003_g N_A_27_367#_c_672_n 5.24515e-19 $X=2.255 $Y=2.465
+ $X2=0 $Y2=0
cc_283 N_A_436_21#_M1020_g N_A_27_367#_c_672_n 0.00679325f $X=2.685 $Y=2.465
+ $X2=0 $Y2=0
cc_284 N_A_436_21#_c_270_n N_VPWR_M1004_s 0.00313148f $X=3.575 $Y=1.845 $X2=0
+ $Y2=0
cc_285 N_A_436_21#_M1003_g N_VPWR_c_731_n 0.00105139f $X=2.255 $Y=2.465 $X2=0
+ $Y2=0
cc_286 N_A_436_21#_M1020_g N_VPWR_c_732_n 0.00301839f $X=2.685 $Y=2.465 $X2=0
+ $Y2=0
cc_287 N_A_436_21#_M1003_g N_VPWR_c_737_n 0.00357877f $X=2.255 $Y=2.465 $X2=0
+ $Y2=0
cc_288 N_A_436_21#_M1020_g N_VPWR_c_737_n 0.00357842f $X=2.685 $Y=2.465 $X2=0
+ $Y2=0
cc_289 N_A_436_21#_M1000_s N_VPWR_c_729_n 0.00231436f $X=4.14 $Y=1.835 $X2=0
+ $Y2=0
cc_290 N_A_436_21#_M1003_g N_VPWR_c_729_n 0.00537654f $X=2.255 $Y=2.465 $X2=0
+ $Y2=0
cc_291 N_A_436_21#_M1020_g N_VPWR_c_729_n 0.00665087f $X=2.685 $Y=2.465 $X2=0
+ $Y2=0
cc_292 N_A_436_21#_c_286_p N_A_742_367#_M1004_d 0.00568075f $X=4.28 $Y=2.035
+ $X2=-0.19 $Y2=-0.245
cc_293 N_A_436_21#_M1000_s N_A_742_367#_c_844_n 0.00374953f $X=4.14 $Y=1.835
+ $X2=0 $Y2=0
cc_294 N_A_436_21#_c_266_n N_VGND_M1013_s 0.0026111f $X=2.84 $Y=1.44 $X2=0 $Y2=0
cc_295 N_A_436_21#_c_278_p N_VGND_M1013_s 0.0175031f $X=3.575 $Y=0.81 $X2=0
+ $Y2=0
cc_296 N_A_436_21#_c_352_p N_VGND_M1013_s 0.00116809f $X=2.925 $Y=0.81 $X2=0
+ $Y2=0
cc_297 N_A_436_21#_c_293_p N_VGND_M1010_s 0.00696198f $X=4.525 $Y=0.81 $X2=0
+ $Y2=0
cc_298 N_A_436_21#_M1001_g N_VGND_c_917_n 0.00897214f $X=2.255 $Y=0.655 $X2=0
+ $Y2=0
cc_299 N_A_436_21#_M1013_g N_VGND_c_917_n 6.13778e-19 $X=2.685 $Y=0.655 $X2=0
+ $Y2=0
cc_300 N_A_436_21#_c_278_p N_VGND_c_918_n 0.00200585f $X=3.575 $Y=0.81 $X2=0
+ $Y2=0
cc_301 N_A_436_21#_c_300_p N_VGND_c_918_n 0.01564f $X=3.67 $Y=0.42 $X2=0 $Y2=0
cc_302 N_A_436_21#_c_293_p N_VGND_c_918_n 0.00211143f $X=4.525 $Y=0.81 $X2=0
+ $Y2=0
cc_303 N_A_436_21#_c_293_p N_VGND_c_919_n 0.0251099f $X=4.525 $Y=0.81 $X2=0
+ $Y2=0
cc_304 N_A_436_21#_c_293_p N_VGND_c_920_n 0.0020834f $X=4.525 $Y=0.81 $X2=0
+ $Y2=0
cc_305 N_A_436_21#_c_299_p N_VGND_c_920_n 0.0188581f $X=4.69 $Y=0.42 $X2=0 $Y2=0
cc_306 N_A_436_21#_M1001_g N_VGND_c_929_n 0.00564095f $X=2.255 $Y=0.655 $X2=0
+ $Y2=0
cc_307 N_A_436_21#_M1013_g N_VGND_c_929_n 0.00486043f $X=2.685 $Y=0.655 $X2=0
+ $Y2=0
cc_308 N_A_436_21#_M1001_g N_VGND_c_930_n 5.59252e-19 $X=2.255 $Y=0.655 $X2=0
+ $Y2=0
cc_309 N_A_436_21#_M1013_g N_VGND_c_930_n 0.00922837f $X=2.685 $Y=0.655 $X2=0
+ $Y2=0
cc_310 N_A_436_21#_c_278_p N_VGND_c_930_n 0.0327177f $X=3.575 $Y=0.81 $X2=0
+ $Y2=0
cc_311 N_A_436_21#_c_352_p N_VGND_c_930_n 0.00964607f $X=2.925 $Y=0.81 $X2=0
+ $Y2=0
cc_312 N_A_436_21#_M1024_s N_VGND_c_934_n 0.00248381f $X=3.53 $Y=0.235 $X2=0
+ $Y2=0
cc_313 N_A_436_21#_M1027_d N_VGND_c_934_n 0.00223559f $X=4.55 $Y=0.235 $X2=0
+ $Y2=0
cc_314 N_A_436_21#_M1001_g N_VGND_c_934_n 0.00948291f $X=2.255 $Y=0.655 $X2=0
+ $Y2=0
cc_315 N_A_436_21#_M1013_g N_VGND_c_934_n 0.00819843f $X=2.685 $Y=0.655 $X2=0
+ $Y2=0
cc_316 N_A_436_21#_c_278_p N_VGND_c_934_n 0.00568502f $X=3.575 $Y=0.81 $X2=0
+ $Y2=0
cc_317 N_A_436_21#_c_352_p N_VGND_c_934_n 7.40073e-19 $X=2.925 $Y=0.81 $X2=0
+ $Y2=0
cc_318 N_A_436_21#_c_300_p N_VGND_c_934_n 0.00985449f $X=3.67 $Y=0.42 $X2=0
+ $Y2=0
cc_319 N_A_436_21#_c_293_p N_VGND_c_934_n 0.00955876f $X=4.525 $Y=0.81 $X2=0
+ $Y2=0
cc_320 N_A_436_21#_c_299_p N_VGND_c_934_n 0.0123659f $X=4.69 $Y=0.42 $X2=0 $Y2=0
cc_321 N_A1_N_c_377_n N_A2_N_c_459_n 0.0161562f $X=3.455 $Y=1.185 $X2=-0.19
+ $Y2=-0.245
cc_322 A1_N N_A2_N_c_459_n 0.00679595f $X=4.475 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_323 N_A1_N_c_378_n N_A2_N_M1000_g 0.0539105f $X=3.635 $Y=1.725 $X2=0 $Y2=0
cc_324 A1_N N_A2_N_c_460_n 0.00379334f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_325 N_A1_N_c_383_n N_A2_N_c_460_n 0.00327998f $X=4.945 $Y=1.35 $X2=0 $Y2=0
cc_326 N_A1_N_c_384_n N_A2_N_c_460_n 0.0167308f $X=4.945 $Y=1.185 $X2=0 $Y2=0
cc_327 N_A1_N_c_378_n N_A2_N_c_464_n 0.00338589f $X=3.635 $Y=1.725 $X2=0 $Y2=0
cc_328 N_A1_N_M1018_g N_A2_N_c_464_n 5.60461e-19 $X=4.925 $Y=2.465 $X2=0 $Y2=0
cc_329 N_A1_N_c_380_n N_A2_N_c_464_n 7.69237e-19 $X=3.41 $Y=1.15 $X2=0 $Y2=0
cc_330 A1_N N_A2_N_c_464_n 0.022512f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_331 N_A1_N_c_383_n N_A2_N_c_464_n 0.00743582f $X=4.945 $Y=1.35 $X2=0 $Y2=0
cc_332 N_A1_N_c_378_n N_A2_N_c_461_n 0.0228462f $X=3.635 $Y=1.725 $X2=0 $Y2=0
cc_333 N_A1_N_M1018_g N_A2_N_c_461_n 0.0619725f $X=4.925 $Y=2.465 $X2=0 $Y2=0
cc_334 N_A1_N_c_380_n N_A2_N_c_461_n 0.00143916f $X=3.41 $Y=1.15 $X2=0 $Y2=0
cc_335 A1_N N_A2_N_c_461_n 0.0259371f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_336 N_A1_N_c_382_n N_A2_N_c_461_n 0.01921f $X=4.945 $Y=1.35 $X2=0 $Y2=0
cc_337 N_A1_N_c_383_n N_A2_N_c_461_n 0.02062f $X=4.945 $Y=1.35 $X2=0 $Y2=0
cc_338 N_A1_N_c_382_n N_A_200_47#_M1006_g 0.0189487f $X=4.945 $Y=1.35 $X2=0
+ $Y2=0
cc_339 N_A1_N_c_383_n N_A_200_47#_M1006_g 0.00223786f $X=4.945 $Y=1.35 $X2=0
+ $Y2=0
cc_340 N_A1_N_c_384_n N_A_200_47#_M1006_g 0.0147361f $X=4.945 $Y=1.185 $X2=0
+ $Y2=0
cc_341 N_A1_N_c_378_n N_A_200_47#_c_555_n 0.0127989f $X=3.635 $Y=1.725 $X2=0
+ $Y2=0
cc_342 N_A1_N_M1018_g N_A_200_47#_c_555_n 0.0169207f $X=4.925 $Y=2.465 $X2=0
+ $Y2=0
cc_343 N_A1_N_M1018_g N_A_200_47#_c_519_n 0.0147046f $X=4.925 $Y=2.465 $X2=0
+ $Y2=0
cc_344 N_A1_N_M1018_g N_A_200_47#_c_520_n 0.00187922f $X=4.925 $Y=2.465 $X2=0
+ $Y2=0
cc_345 N_A1_N_c_382_n N_A_200_47#_c_520_n 8.13042e-19 $X=4.945 $Y=1.35 $X2=0
+ $Y2=0
cc_346 N_A1_N_c_383_n N_A_200_47#_c_520_n 0.00958868f $X=4.945 $Y=1.35 $X2=0
+ $Y2=0
cc_347 N_A1_N_c_378_n N_A_200_47#_c_530_n 0.00760963f $X=3.635 $Y=1.725 $X2=0
+ $Y2=0
cc_348 N_A1_N_M1018_g N_A_200_47#_c_522_n 0.0426433f $X=4.925 $Y=2.465 $X2=0
+ $Y2=0
cc_349 N_A1_N_c_382_n N_A_200_47#_c_522_n 0.00215311f $X=4.945 $Y=1.35 $X2=0
+ $Y2=0
cc_350 N_A1_N_c_378_n N_A_27_367#_c_671_n 5.6196e-19 $X=3.635 $Y=1.725 $X2=0
+ $Y2=0
cc_351 N_A1_N_c_378_n N_A_27_367#_c_672_n 0.00365671f $X=3.635 $Y=1.725 $X2=0
+ $Y2=0
cc_352 N_A1_N_c_378_n N_VPWR_c_732_n 0.0141923f $X=3.635 $Y=1.725 $X2=0 $Y2=0
cc_353 N_A1_N_M1018_g N_VPWR_c_733_n 0.0038871f $X=4.925 $Y=2.465 $X2=0 $Y2=0
cc_354 N_A1_N_c_378_n N_VPWR_c_741_n 0.00486043f $X=3.635 $Y=1.725 $X2=0 $Y2=0
cc_355 N_A1_N_M1018_g N_VPWR_c_741_n 0.00585385f $X=4.925 $Y=2.465 $X2=0 $Y2=0
cc_356 N_A1_N_c_378_n N_VPWR_c_729_n 0.00466752f $X=3.635 $Y=1.725 $X2=0 $Y2=0
cc_357 N_A1_N_M1018_g N_VPWR_c_729_n 0.0065574f $X=4.925 $Y=2.465 $X2=0 $Y2=0
cc_358 N_A1_N_c_383_n N_X_c_855_n 0.00770034f $X=4.945 $Y=1.35 $X2=0 $Y2=0
cc_359 N_A1_N_c_380_n N_VGND_M1013_s 9.64592e-19 $X=3.41 $Y=1.15 $X2=0 $Y2=0
cc_360 A1_N N_VGND_M1010_s 0.00342061f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_361 N_A1_N_c_377_n N_VGND_c_918_n 0.00364083f $X=3.455 $Y=1.185 $X2=0 $Y2=0
cc_362 N_A1_N_c_384_n N_VGND_c_920_n 0.0054895f $X=4.945 $Y=1.185 $X2=0 $Y2=0
cc_363 N_A1_N_c_382_n N_VGND_c_921_n 0.00276251f $X=4.945 $Y=1.35 $X2=0 $Y2=0
cc_364 N_A1_N_c_383_n N_VGND_c_921_n 2.50277e-19 $X=4.945 $Y=1.35 $X2=0 $Y2=0
cc_365 N_A1_N_c_384_n N_VGND_c_921_n 0.00300596f $X=4.945 $Y=1.185 $X2=0 $Y2=0
cc_366 N_A1_N_c_377_n N_VGND_c_930_n 0.00868226f $X=3.455 $Y=1.185 $X2=0 $Y2=0
cc_367 N_A1_N_c_377_n N_VGND_c_934_n 0.0043218f $X=3.455 $Y=1.185 $X2=0 $Y2=0
cc_368 N_A1_N_c_384_n N_VGND_c_934_n 0.00995442f $X=4.945 $Y=1.185 $X2=0 $Y2=0
cc_369 N_A2_N_M1000_g N_A_200_47#_c_555_n 0.0105614f $X=4.065 $Y=2.465 $X2=0
+ $Y2=0
cc_370 N_A2_N_M1012_g N_A_200_47#_c_555_n 0.0143791f $X=4.495 $Y=2.465 $X2=0
+ $Y2=0
cc_371 N_A2_N_M1000_g N_VPWR_c_732_n 0.00143205f $X=4.065 $Y=2.465 $X2=0 $Y2=0
cc_372 N_A2_N_M1000_g N_VPWR_c_741_n 0.00373071f $X=4.065 $Y=2.465 $X2=0 $Y2=0
cc_373 N_A2_N_M1012_g N_VPWR_c_741_n 0.00373071f $X=4.495 $Y=2.465 $X2=0 $Y2=0
cc_374 N_A2_N_M1000_g N_VPWR_c_729_n 0.00548684f $X=4.065 $Y=2.465 $X2=0 $Y2=0
cc_375 N_A2_N_M1012_g N_VPWR_c_729_n 0.00548684f $X=4.495 $Y=2.465 $X2=0 $Y2=0
cc_376 N_A2_N_M1000_g N_A_742_367#_c_844_n 0.0124277f $X=4.065 $Y=2.465 $X2=0
+ $Y2=0
cc_377 N_A2_N_M1012_g N_A_742_367#_c_844_n 0.0124277f $X=4.495 $Y=2.465 $X2=0
+ $Y2=0
cc_378 N_A2_N_c_459_n N_VGND_c_918_n 0.00428679f $X=3.89 $Y=1.185 $X2=0 $Y2=0
cc_379 N_A2_N_c_459_n N_VGND_c_919_n 0.00369955f $X=3.89 $Y=1.185 $X2=0 $Y2=0
cc_380 N_A2_N_c_460_n N_VGND_c_919_n 0.00507717f $X=4.475 $Y=1.185 $X2=0 $Y2=0
cc_381 N_A2_N_c_460_n N_VGND_c_920_n 0.00426006f $X=4.475 $Y=1.185 $X2=0 $Y2=0
cc_382 N_A2_N_c_459_n N_VGND_c_930_n 4.98814e-19 $X=3.89 $Y=1.185 $X2=0 $Y2=0
cc_383 N_A2_N_c_459_n N_VGND_c_934_n 0.006337f $X=3.89 $Y=1.185 $X2=0 $Y2=0
cc_384 N_A2_N_c_460_n N_VGND_c_934_n 0.0063111f $X=4.475 $Y=1.185 $X2=0 $Y2=0
cc_385 N_A_200_47#_c_528_n N_A_27_367#_M1020_s 0.00498046f $X=3.235 $Y=2.185
+ $X2=0 $Y2=0
cc_386 N_A_200_47#_c_516_n N_A_27_367#_c_670_n 0.00732675f $X=2.345 $Y=1.15
+ $X2=0 $Y2=0
cc_387 N_A_200_47#_c_518_n N_A_27_367#_c_670_n 0.00149665f $X=2.47 $Y=1.98 $X2=0
+ $Y2=0
cc_388 N_A_200_47#_M1003_d N_A_27_367#_c_671_n 0.00332344f $X=2.33 $Y=1.835
+ $X2=0 $Y2=0
cc_389 N_A_200_47#_c_582_p N_A_27_367#_c_671_n 0.0126348f $X=2.47 $Y=2.57 $X2=0
+ $Y2=0
cc_390 N_A_200_47#_c_528_n N_A_27_367#_c_671_n 0.00282113f $X=3.235 $Y=2.185
+ $X2=0 $Y2=0
cc_391 N_A_200_47#_c_528_n N_A_27_367#_c_672_n 0.0218796f $X=3.235 $Y=2.185
+ $X2=0 $Y2=0
cc_392 N_A_200_47#_c_530_n N_A_27_367#_c_672_n 0.00317136f $X=3.32 $Y=2.185
+ $X2=0 $Y2=0
cc_393 N_A_200_47#_c_555_n N_VPWR_M1004_s 0.00288705f $X=5.21 $Y=2.395 $X2=0
+ $Y2=0
cc_394 N_A_200_47#_c_530_n N_VPWR_M1004_s 0.00675234f $X=3.32 $Y=2.185 $X2=0
+ $Y2=0
cc_395 N_A_200_47#_c_555_n N_VPWR_M1018_s 0.00823584f $X=5.21 $Y=2.395 $X2=0
+ $Y2=0
cc_396 N_A_200_47#_c_519_n N_VPWR_M1018_s 0.0056566f $X=5.295 $Y=2.31 $X2=0
+ $Y2=0
cc_397 N_A_200_47#_c_555_n N_VPWR_c_732_n 0.00955265f $X=5.21 $Y=2.395 $X2=0
+ $Y2=0
cc_398 N_A_200_47#_c_530_n N_VPWR_c_732_n 0.0126358f $X=3.32 $Y=2.185 $X2=0
+ $Y2=0
cc_399 N_A_200_47#_M1009_g N_VPWR_c_733_n 0.008998f $X=5.42 $Y=2.465 $X2=0 $Y2=0
cc_400 N_A_200_47#_M1016_g N_VPWR_c_733_n 5.64123e-19 $X=5.86 $Y=2.465 $X2=0
+ $Y2=0
cc_401 N_A_200_47#_c_555_n N_VPWR_c_733_n 0.0192656f $X=5.21 $Y=2.395 $X2=0
+ $Y2=0
cc_402 N_A_200_47#_M1009_g N_VPWR_c_734_n 7.26754e-19 $X=5.42 $Y=2.465 $X2=0
+ $Y2=0
cc_403 N_A_200_47#_M1016_g N_VPWR_c_734_n 0.0143056f $X=5.86 $Y=2.465 $X2=0
+ $Y2=0
cc_404 N_A_200_47#_M1022_g N_VPWR_c_734_n 0.0142882f $X=6.29 $Y=2.465 $X2=0
+ $Y2=0
cc_405 N_A_200_47#_M1023_g N_VPWR_c_734_n 7.39378e-19 $X=6.72 $Y=2.465 $X2=0
+ $Y2=0
cc_406 N_A_200_47#_M1023_g N_VPWR_c_736_n 0.00341818f $X=6.72 $Y=2.465 $X2=0
+ $Y2=0
cc_407 N_A_200_47#_M1009_g N_VPWR_c_742_n 0.00564095f $X=5.42 $Y=2.465 $X2=0
+ $Y2=0
cc_408 N_A_200_47#_M1016_g N_VPWR_c_742_n 0.00486043f $X=5.86 $Y=2.465 $X2=0
+ $Y2=0
cc_409 N_A_200_47#_M1022_g N_VPWR_c_743_n 0.00486043f $X=6.29 $Y=2.465 $X2=0
+ $Y2=0
cc_410 N_A_200_47#_M1023_g N_VPWR_c_743_n 0.00585385f $X=6.72 $Y=2.465 $X2=0
+ $Y2=0
cc_411 N_A_200_47#_M1003_d N_VPWR_c_729_n 0.00225186f $X=2.33 $Y=1.835 $X2=0
+ $Y2=0
cc_412 N_A_200_47#_M1009_g N_VPWR_c_729_n 0.00859431f $X=5.42 $Y=2.465 $X2=0
+ $Y2=0
cc_413 N_A_200_47#_M1016_g N_VPWR_c_729_n 0.00827314f $X=5.86 $Y=2.465 $X2=0
+ $Y2=0
cc_414 N_A_200_47#_M1022_g N_VPWR_c_729_n 0.00824727f $X=6.29 $Y=2.465 $X2=0
+ $Y2=0
cc_415 N_A_200_47#_M1023_g N_VPWR_c_729_n 0.011446f $X=6.72 $Y=2.465 $X2=0 $Y2=0
cc_416 N_A_200_47#_c_555_n N_VPWR_c_729_n 0.0138997f $X=5.21 $Y=2.395 $X2=0
+ $Y2=0
cc_417 N_A_200_47#_c_530_n N_VPWR_c_729_n 0.00124074f $X=3.32 $Y=2.185 $X2=0
+ $Y2=0
cc_418 N_A_200_47#_c_555_n N_A_742_367#_M1004_d 0.00359746f $X=5.21 $Y=2.395
+ $X2=-0.19 $Y2=-0.245
cc_419 N_A_200_47#_c_555_n N_A_742_367#_M1012_d 0.00816237f $X=5.21 $Y=2.395
+ $X2=0 $Y2=0
cc_420 N_A_200_47#_c_555_n N_A_742_367#_c_844_n 0.0528662f $X=5.21 $Y=2.395
+ $X2=0 $Y2=0
cc_421 N_A_200_47#_M1008_g N_X_c_854_n 0.0138955f $X=5.825 $Y=0.655 $X2=0 $Y2=0
cc_422 N_A_200_47#_M1014_g N_X_c_854_n 0.014114f $X=6.255 $Y=0.655 $X2=0 $Y2=0
cc_423 N_A_200_47#_c_616_p N_X_c_854_n 0.0469271f $X=6.53 $Y=1.49 $X2=0 $Y2=0
cc_424 N_A_200_47#_c_522_n N_X_c_854_n 0.00261515f $X=6.685 $Y=1.49 $X2=0 $Y2=0
cc_425 N_A_200_47#_M1006_g N_X_c_855_n 0.00229451f $X=5.395 $Y=0.655 $X2=0 $Y2=0
cc_426 N_A_200_47#_c_616_p N_X_c_855_n 0.0186281f $X=6.53 $Y=1.49 $X2=0 $Y2=0
cc_427 N_A_200_47#_c_522_n N_X_c_855_n 0.00267516f $X=6.685 $Y=1.49 $X2=0 $Y2=0
cc_428 N_A_200_47#_M1016_g N_X_c_860_n 0.0130217f $X=5.86 $Y=2.465 $X2=0 $Y2=0
cc_429 N_A_200_47#_M1022_g N_X_c_860_n 0.013144f $X=6.29 $Y=2.465 $X2=0 $Y2=0
cc_430 N_A_200_47#_c_616_p N_X_c_860_n 0.0469272f $X=6.53 $Y=1.49 $X2=0 $Y2=0
cc_431 N_A_200_47#_c_522_n N_X_c_860_n 0.00258422f $X=6.685 $Y=1.49 $X2=0 $Y2=0
cc_432 N_A_200_47#_M1009_g N_X_c_861_n 6.52891e-19 $X=5.42 $Y=2.465 $X2=0 $Y2=0
cc_433 N_A_200_47#_c_519_n N_X_c_861_n 0.00947169f $X=5.295 $Y=2.31 $X2=0 $Y2=0
cc_434 N_A_200_47#_c_616_p N_X_c_861_n 0.0153878f $X=6.53 $Y=1.49 $X2=0 $Y2=0
cc_435 N_A_200_47#_c_522_n N_X_c_861_n 0.00293877f $X=6.685 $Y=1.49 $X2=0 $Y2=0
cc_436 N_A_200_47#_M1023_g N_X_c_862_n 0.0161899f $X=6.72 $Y=2.465 $X2=0 $Y2=0
cc_437 N_A_200_47#_c_616_p N_X_c_862_n 0.00444395f $X=6.53 $Y=1.49 $X2=0 $Y2=0
cc_438 N_A_200_47#_c_616_p N_X_c_856_n 0.015388f $X=6.53 $Y=1.49 $X2=0 $Y2=0
cc_439 N_A_200_47#_c_522_n N_X_c_856_n 0.00271819f $X=6.685 $Y=1.49 $X2=0 $Y2=0
cc_440 N_A_200_47#_c_616_p N_X_c_863_n 0.0178182f $X=6.53 $Y=1.49 $X2=0 $Y2=0
cc_441 N_A_200_47#_c_522_n N_X_c_863_n 0.00268515f $X=6.685 $Y=1.49 $X2=0 $Y2=0
cc_442 N_A_200_47#_M1015_g X 0.0162151f $X=6.685 $Y=0.655 $X2=0 $Y2=0
cc_443 N_A_200_47#_c_616_p X 0.00898195f $X=6.53 $Y=1.49 $X2=0 $Y2=0
cc_444 N_A_200_47#_c_522_n X 0.00116067f $X=6.685 $Y=1.49 $X2=0 $Y2=0
cc_445 N_A_200_47#_M1015_g X 0.00323451f $X=6.685 $Y=0.655 $X2=0 $Y2=0
cc_446 N_A_200_47#_c_616_p X 0.0136179f $X=6.53 $Y=1.49 $X2=0 $Y2=0
cc_447 N_A_200_47#_c_522_n X 0.0159329f $X=6.685 $Y=1.49 $X2=0 $Y2=0
cc_448 N_A_200_47#_c_516_n N_VGND_M1007_d 0.00218982f $X=2.345 $Y=1.15 $X2=0
+ $Y2=0
cc_449 N_A_200_47#_c_516_n N_VGND_c_917_n 0.0170224f $X=2.345 $Y=1.15 $X2=0
+ $Y2=0
cc_450 N_A_200_47#_M1006_g N_VGND_c_921_n 0.00167704f $X=5.395 $Y=0.655 $X2=0
+ $Y2=0
cc_451 N_A_200_47#_c_520_n N_VGND_c_921_n 0.00305572f $X=5.38 $Y=1.495 $X2=0
+ $Y2=0
cc_452 N_A_200_47#_M1006_g N_VGND_c_922_n 6.3872e-19 $X=5.395 $Y=0.655 $X2=0
+ $Y2=0
cc_453 N_A_200_47#_M1008_g N_VGND_c_922_n 0.0109629f $X=5.825 $Y=0.655 $X2=0
+ $Y2=0
cc_454 N_A_200_47#_M1014_g N_VGND_c_922_n 0.010871f $X=6.255 $Y=0.655 $X2=0
+ $Y2=0
cc_455 N_A_200_47#_M1015_g N_VGND_c_922_n 6.22495e-19 $X=6.685 $Y=0.655 $X2=0
+ $Y2=0
cc_456 N_A_200_47#_M1014_g N_VGND_c_924_n 6.30983e-19 $X=6.255 $Y=0.655 $X2=0
+ $Y2=0
cc_457 N_A_200_47#_M1015_g N_VGND_c_924_n 0.0130637f $X=6.685 $Y=0.655 $X2=0
+ $Y2=0
cc_458 N_A_200_47#_M1006_g N_VGND_c_927_n 0.00585385f $X=5.395 $Y=0.655 $X2=0
+ $Y2=0
cc_459 N_A_200_47#_M1008_g N_VGND_c_927_n 0.00486043f $X=5.825 $Y=0.655 $X2=0
+ $Y2=0
cc_460 N_A_200_47#_M1014_g N_VGND_c_928_n 0.00486043f $X=6.255 $Y=0.655 $X2=0
+ $Y2=0
cc_461 N_A_200_47#_M1015_g N_VGND_c_928_n 0.00486043f $X=6.685 $Y=0.655 $X2=0
+ $Y2=0
cc_462 N_A_200_47#_c_655_p N_VGND_c_929_n 0.0128073f $X=2.47 $Y=0.42 $X2=0 $Y2=0
cc_463 N_A_200_47#_M1005_d N_VGND_c_934_n 0.00225186f $X=1 $Y=0.235 $X2=0 $Y2=0
cc_464 N_A_200_47#_M1001_d N_VGND_c_934_n 0.00501859f $X=2.33 $Y=0.235 $X2=0
+ $Y2=0
cc_465 N_A_200_47#_M1006_g N_VGND_c_934_n 0.0106995f $X=5.395 $Y=0.655 $X2=0
+ $Y2=0
cc_466 N_A_200_47#_M1008_g N_VGND_c_934_n 0.00824727f $X=5.825 $Y=0.655 $X2=0
+ $Y2=0
cc_467 N_A_200_47#_M1014_g N_VGND_c_934_n 0.00824727f $X=6.255 $Y=0.655 $X2=0
+ $Y2=0
cc_468 N_A_200_47#_M1015_g N_VGND_c_934_n 0.00824727f $X=6.685 $Y=0.655 $X2=0
+ $Y2=0
cc_469 N_A_200_47#_c_655_p N_VGND_c_934_n 0.00769778f $X=2.47 $Y=0.42 $X2=0
+ $Y2=0
cc_470 N_A_200_47#_c_516_n N_A_114_47#_M1021_s 0.00176461f $X=2.345 $Y=1.15
+ $X2=0 $Y2=0
cc_471 N_A_200_47#_M1005_d N_A_114_47#_c_1038_n 0.00332344f $X=1 $Y=0.235 $X2=0
+ $Y2=0
cc_472 N_A_200_47#_c_665_p N_A_114_47#_c_1038_n 0.0125759f $X=1.14 $Y=0.76 $X2=0
+ $Y2=0
cc_473 N_A_200_47#_c_516_n N_A_114_47#_c_1038_n 0.00280043f $X=2.345 $Y=1.15
+ $X2=0 $Y2=0
cc_474 N_A_200_47#_c_517_n N_A_114_47#_c_1034_n 0.00206756f $X=1.235 $Y=1.15
+ $X2=0 $Y2=0
cc_475 N_A_200_47#_c_516_n N_A_114_47#_c_1037_n 0.0169932f $X=2.345 $Y=1.15
+ $X2=0 $Y2=0
cc_476 N_A_27_367#_c_679_n N_VPWR_M1011_s 0.00352062f $X=1.045 $Y=2.375
+ $X2=-0.19 $Y2=1.655
cc_477 N_A_27_367#_c_683_n N_VPWR_M1026_d 0.00480022f $X=1.935 $Y=2.375 $X2=0
+ $Y2=0
cc_478 N_A_27_367#_c_679_n N_VPWR_c_730_n 0.0170777f $X=1.045 $Y=2.375 $X2=0
+ $Y2=0
cc_479 N_A_27_367#_c_683_n N_VPWR_c_731_n 0.017285f $X=1.935 $Y=2.375 $X2=0
+ $Y2=0
cc_480 N_A_27_367#_c_671_n N_VPWR_c_732_n 0.0139f $X=2.735 $Y=2.99 $X2=0 $Y2=0
cc_481 N_A_27_367#_c_672_n N_VPWR_c_732_n 0.0195971f $X=2.9 $Y=2.535 $X2=0 $Y2=0
cc_482 N_A_27_367#_c_671_n N_VPWR_c_737_n 0.0526725f $X=2.735 $Y=2.99 $X2=0
+ $Y2=0
cc_483 N_A_27_367#_c_718_p N_VPWR_c_737_n 0.0142975f $X=2.175 $Y=2.99 $X2=0
+ $Y2=0
cc_484 N_A_27_367#_c_673_n N_VPWR_c_739_n 0.0192173f $X=0.26 $Y=2.45 $X2=0 $Y2=0
cc_485 N_A_27_367#_c_720_p N_VPWR_c_740_n 0.0131621f $X=1.14 $Y=2.465 $X2=0
+ $Y2=0
cc_486 N_A_27_367#_M1011_d N_VPWR_c_729_n 0.00388458f $X=0.135 $Y=1.835 $X2=0
+ $Y2=0
cc_487 N_A_27_367#_M1019_s N_VPWR_c_729_n 0.00467071f $X=1 $Y=1.835 $X2=0 $Y2=0
cc_488 N_A_27_367#_M1017_d N_VPWR_c_729_n 0.0033862f $X=1.9 $Y=1.835 $X2=0 $Y2=0
cc_489 N_A_27_367#_M1020_s N_VPWR_c_729_n 0.00215158f $X=2.76 $Y=1.835 $X2=0
+ $Y2=0
cc_490 N_A_27_367#_c_720_p N_VPWR_c_729_n 0.00808656f $X=1.14 $Y=2.465 $X2=0
+ $Y2=0
cc_491 N_A_27_367#_c_671_n N_VPWR_c_729_n 0.0323445f $X=2.735 $Y=2.99 $X2=0
+ $Y2=0
cc_492 N_A_27_367#_c_718_p N_VPWR_c_729_n 0.00932008f $X=2.175 $Y=2.99 $X2=0
+ $Y2=0
cc_493 N_A_27_367#_c_673_n N_VPWR_c_729_n 0.010808f $X=0.26 $Y=2.45 $X2=0 $Y2=0
cc_494 N_VPWR_c_729_n N_A_742_367#_M1004_d 0.00260949f $X=6.96 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_495 N_VPWR_c_729_n N_A_742_367#_M1012_d 0.00231436f $X=6.96 $Y=3.33 $X2=0
+ $Y2=0
cc_496 N_VPWR_c_741_n N_A_742_367#_c_844_n 0.0424961f $X=5.02 $Y=3.33 $X2=0
+ $Y2=0
cc_497 N_VPWR_c_729_n N_A_742_367#_c_844_n 0.0385305f $X=6.96 $Y=3.33 $X2=0
+ $Y2=0
cc_498 N_VPWR_c_729_n N_X_M1009_s 0.00579476f $X=6.96 $Y=3.33 $X2=0 $Y2=0
cc_499 N_VPWR_c_729_n N_X_M1022_s 0.00432284f $X=6.96 $Y=3.33 $X2=0 $Y2=0
cc_500 N_VPWR_c_742_n N_X_c_895_n 0.0128008f $X=5.91 $Y=3.33 $X2=0 $Y2=0
cc_501 N_VPWR_c_729_n N_X_c_895_n 0.00730372f $X=6.96 $Y=3.33 $X2=0 $Y2=0
cc_502 N_VPWR_M1016_d N_X_c_860_n 0.00176461f $X=5.935 $Y=1.835 $X2=0 $Y2=0
cc_503 N_VPWR_c_734_n N_X_c_860_n 0.0170777f $X=6.075 $Y=2.26 $X2=0 $Y2=0
cc_504 N_VPWR_c_743_n N_X_c_899_n 0.0135169f $X=6.8 $Y=3.33 $X2=0 $Y2=0
cc_505 N_VPWR_c_729_n N_X_c_899_n 0.00847534f $X=6.96 $Y=3.33 $X2=0 $Y2=0
cc_506 N_VPWR_M1023_d N_X_c_862_n 0.00652378f $X=6.795 $Y=1.835 $X2=0 $Y2=0
cc_507 N_VPWR_c_736_n N_X_c_862_n 0.0171623f $X=6.935 $Y=2.26 $X2=0 $Y2=0
cc_508 N_X_c_854_n N_VGND_M1008_s 0.00189202f $X=6.375 $Y=1.15 $X2=0 $Y2=0
cc_509 X N_VGND_M1015_s 6.05921e-19 $X=6.875 $Y=1.21 $X2=0 $Y2=0
cc_510 N_X_c_858_n N_VGND_M1015_s 0.00239048f $X=6.96 $Y=1.235 $X2=0 $Y2=0
cc_511 N_X_c_854_n N_VGND_c_922_n 0.0150989f $X=6.375 $Y=1.15 $X2=0 $Y2=0
cc_512 X N_VGND_c_924_n 0.0064684f $X=6.875 $Y=1.21 $X2=0 $Y2=0
cc_513 N_X_c_858_n N_VGND_c_924_n 0.0153275f $X=6.96 $Y=1.235 $X2=0 $Y2=0
cc_514 N_X_c_909_p N_VGND_c_927_n 0.0138717f $X=5.61 $Y=0.42 $X2=0 $Y2=0
cc_515 N_X_c_910_p N_VGND_c_928_n 0.0124525f $X=6.47 $Y=0.42 $X2=0 $Y2=0
cc_516 N_X_M1006_d N_VGND_c_934_n 0.00397496f $X=5.47 $Y=0.235 $X2=0 $Y2=0
cc_517 N_X_M1014_d N_VGND_c_934_n 0.00536646f $X=6.33 $Y=0.235 $X2=0 $Y2=0
cc_518 N_X_c_909_p N_VGND_c_934_n 0.00886411f $X=5.61 $Y=0.42 $X2=0 $Y2=0
cc_519 N_X_c_910_p N_VGND_c_934_n 0.00730901f $X=6.47 $Y=0.42 $X2=0 $Y2=0
cc_520 N_VGND_c_934_n N_A_114_47#_M1002_s 0.00223559f $X=6.96 $Y=0 $X2=-0.19
+ $Y2=-0.245
cc_521 N_VGND_c_934_n N_A_114_47#_M1021_s 0.00223559f $X=6.96 $Y=0 $X2=0 $Y2=0
cc_522 N_VGND_c_925_n N_A_114_47#_c_1038_n 0.031405f $X=1.905 $Y=0 $X2=0 $Y2=0
cc_523 N_VGND_c_934_n N_A_114_47#_c_1038_n 0.0195789f $X=6.96 $Y=0 $X2=0 $Y2=0
cc_524 N_VGND_c_916_n N_A_114_47#_c_1034_n 0.0230122f $X=0.28 $Y=0.38 $X2=0
+ $Y2=0
cc_525 N_VGND_c_925_n N_A_114_47#_c_1034_n 0.0157167f $X=1.905 $Y=0 $X2=0 $Y2=0
cc_526 N_VGND_c_934_n N_A_114_47#_c_1034_n 0.010808f $X=6.96 $Y=0 $X2=0 $Y2=0
cc_527 N_VGND_c_925_n N_A_114_47#_c_1037_n 0.0189944f $X=1.905 $Y=0 $X2=0 $Y2=0
cc_528 N_VGND_c_934_n N_A_114_47#_c_1037_n 0.0124345f $X=6.96 $Y=0 $X2=0 $Y2=0
