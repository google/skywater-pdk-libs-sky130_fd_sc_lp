* NGSPICE file created from sky130_fd_sc_lp__a21boi_2.ext - technology: sky130A

.subckt sky130_fd_sc_lp__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
M1000 VPWR A1 a_231_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=1.0185e+12p pd=7.85e+06u as=1.3734e+12p ps=1.226e+07u
M1001 VPWR A2 a_231_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1002 Y a_119_500# VGND VNB nshort w=840000u l=150000u
+  ad=5.376e+11p pd=4.64e+06u as=7.938e+11p ps=7.04e+06u
M1003 Y A1 a_502_65# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=4.704e+11p ps=4.48e+06u
M1004 a_231_367# a_119_500# Y VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=3.528e+11p ps=3.08e+06u
M1005 a_502_65# A1 Y VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_231_367# A1 VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND a_119_500# Y VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_231_367# A2 VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_502_65# A2 VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 Y a_119_500# a_231_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_119_500# B1_N VPWR VPB phighvt w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1012 VGND B1_N a_119_500# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1013 VGND A2 a_502_65# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

