* NGSPICE file created from sky130_fd_sc_lp__a2111o_1.ext - technology: sky130A

.subckt sky130_fd_sc_lp__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
M1000 VGND C1 a_105_239# VNB nshort w=840000u l=150000u
+  ad=1.155e+12p pd=7.79e+06u as=7.896e+11p ps=5.24e+06u
M1001 a_403_367# C1 a_325_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=4.914e+11p pd=3.3e+06u as=3.024e+11p ps=3e+06u
M1002 a_511_367# A2 VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=1.1151e+12p pd=6.81e+06u as=6.867e+11p ps=6.13e+06u
M1003 a_105_239# B1 VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_511_367# B1 a_403_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_673_49# A1 a_105_239# VNB nshort w=840000u l=150000u
+  ad=1.764e+11p pd=2.1e+06u as=0p ps=0u
M1006 VGND A2 a_673_49# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR A1 a_511_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPWR a_105_239# X VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=3.339e+11p ps=3.05e+06u
M1009 a_325_367# D1 a_105_239# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=3.339e+11p ps=3.05e+06u
M1010 VGND a_105_239# X VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=2.226e+11p ps=2.21e+06u
M1011 a_105_239# D1 VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

