* File: sky130_fd_sc_lp__dfxtp_2.pex.spice
* Created: Fri Aug 28 10:24:21 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__DFXTP_2%CLK 2 5 8 10 11 12 13 14 15 22 24
r25 22 24 45.5639 $w=3.95e-07 $l=1.65e-07 $layer=POLY_cond $X=0.352 $Y=1.005
+ $X2=0.352 $Y2=0.84
r26 14 15 12.5413 $w=3.38e-07 $l=3.7e-07 $layer=LI1_cond $X=0.255 $Y=2.035
+ $X2=0.255 $Y2=2.405
r27 13 14 12.5413 $w=3.38e-07 $l=3.7e-07 $layer=LI1_cond $X=0.255 $Y=1.665
+ $X2=0.255 $Y2=2.035
r28 12 13 12.5413 $w=3.38e-07 $l=3.7e-07 $layer=LI1_cond $X=0.255 $Y=1.295
+ $X2=0.255 $Y2=1.665
r29 11 12 12.5413 $w=3.38e-07 $l=3.7e-07 $layer=LI1_cond $X=0.255 $Y=0.925
+ $X2=0.255 $Y2=1.295
r30 11 22 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.32
+ $Y=1.005 $X2=0.32 $Y2=1.005
r31 8 10 620.447 $w=1.5e-07 $l=1.21e-06 $layer=POLY_cond $X=0.475 $Y=2.72
+ $X2=0.475 $Y2=1.51
r32 5 24 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.475 $Y=0.52
+ $X2=0.475 $Y2=0.84
r33 2 10 50.0695 $w=3.95e-07 $l=1.97e-07 $layer=POLY_cond $X=0.352 $Y=1.313
+ $X2=0.352 $Y2=1.51
r34 1 22 4.50555 $w=3.95e-07 $l=3.2e-08 $layer=POLY_cond $X=0.352 $Y=1.037
+ $X2=0.352 $Y2=1.005
r35 1 2 38.8604 $w=3.95e-07 $l=2.76e-07 $layer=POLY_cond $X=0.352 $Y=1.037
+ $X2=0.352 $Y2=1.313
.ends

.subckt PM_SKY130_FD_SC_LP__DFXTP_2%D 3 6 8 9 13 15
c40 8 0 3.84473e-21 $X=2.16 $Y=1.295
r41 13 16 88.6355 $w=4.55e-07 $l=5.05e-07 $layer=POLY_cond $X=2.167 $Y=1.295
+ $X2=2.167 $Y2=1.8
r42 13 15 47.0767 $w=4.55e-07 $l=1.65e-07 $layer=POLY_cond $X=2.167 $Y=1.295
+ $X2=2.167 $Y2=1.13
r43 8 9 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=2.105 $Y=1.295
+ $X2=2.105 $Y2=1.665
r44 8 13 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.105
+ $Y=1.295 $X2=2.105 $Y2=1.295
r45 6 16 320.479 $w=1.5e-07 $l=6.25e-07 $layer=POLY_cond $X=2.32 $Y=2.425
+ $X2=2.32 $Y2=1.8
r46 3 15 104.433 $w=1.5e-07 $l=3.25e-07 $layer=POLY_cond $X=2.085 $Y=0.805
+ $X2=2.085 $Y2=1.13
.ends

.subckt PM_SKY130_FD_SC_LP__DFXTP_2%A_240_443# 1 2 9 13 17 19 21 23 26 28 31 35
+ 37 40 41 42 45 46 48 51 52 53 54 55 56 57 60
c162 54 0 6.46168e-20 $X=5.075 $Y=1.555
c163 48 0 4.80136e-20 $X=3.52 $Y=2.85
c164 26 0 9.35787e-20 $X=2.93 $Y=1.535
r165 59 60 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.14
+ $Y=1.39 $X2=5.14 $Y2=1.39
r166 54 59 8.60334 $w=3.26e-07 $l=1.94808e-07 $layer=LI1_cond $X=5.075 $Y=1.555
+ $X2=5.14 $Y2=1.39
r167 54 55 44.9798 $w=1.78e-07 $l=7.3e-07 $layer=LI1_cond $X=5.075 $Y=1.555
+ $X2=5.075 $Y2=2.285
r168 52 55 6.82373 $w=1.7e-07 $l=1.25499e-07 $layer=LI1_cond $X=4.985 $Y=2.37
+ $X2=5.075 $Y2=2.285
r169 52 53 84.4866 $w=1.68e-07 $l=1.295e-06 $layer=LI1_cond $X=4.985 $Y=2.37
+ $X2=3.69 $Y2=2.37
r170 50 53 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.605 $Y=2.455
+ $X2=3.69 $Y2=2.37
r171 50 51 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3.605 $Y=2.455
+ $X2=3.605 $Y2=2.76
r172 49 57 4.92476 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.97 $Y=2.85
+ $X2=2.885 $Y2=2.85
r173 48 51 6.82373 $w=1.8e-07 $l=1.25499e-07 $layer=LI1_cond $X=3.52 $Y=2.85
+ $X2=3.605 $Y2=2.76
r174 48 49 33.8889 $w=1.78e-07 $l=5.5e-07 $layer=LI1_cond $X=3.52 $Y=2.85
+ $X2=2.97 $Y2=2.85
r175 45 46 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.885
+ $Y=1.55 $X2=2.885 $Y2=1.55
r176 43 57 1.54918 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=2.885 $Y=2.76
+ $X2=2.885 $Y2=2.85
r177 43 45 78.9412 $w=1.68e-07 $l=1.21e-06 $layer=LI1_cond $X=2.885 $Y=2.76
+ $X2=2.885 $Y2=1.55
r178 41 57 4.92476 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.8 $Y=2.85
+ $X2=2.885 $Y2=2.85
r179 41 42 32.6566 $w=1.78e-07 $l=5.3e-07 $layer=LI1_cond $X=2.8 $Y=2.85
+ $X2=2.27 $Y2=2.85
r180 40 42 6.81649 $w=1.8e-07 $l=1.27279e-07 $layer=LI1_cond $X=2.18 $Y=2.76
+ $X2=2.27 $Y2=2.85
r181 39 40 40.3586 $w=1.78e-07 $l=6.55e-07 $layer=LI1_cond $X=2.18 $Y=2.105
+ $X2=2.18 $Y2=2.76
r182 38 56 3.35233 $w=1.7e-07 $l=1.88e-07 $layer=LI1_cond $X=1.585 $Y=2.02
+ $X2=1.397 $Y2=2.02
r183 37 39 6.82373 $w=1.7e-07 $l=1.25499e-07 $layer=LI1_cond $X=2.09 $Y=2.02
+ $X2=2.18 $Y2=2.105
r184 37 38 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=2.09 $Y=2.02
+ $X2=1.585 $Y2=2.02
r185 33 56 3.22182 $w=2.92e-07 $l=1.19143e-07 $layer=LI1_cond $X=1.315 $Y=2.105
+ $X2=1.397 $Y2=2.02
r186 33 35 13.4675 $w=2.08e-07 $l=2.55e-07 $layer=LI1_cond $X=1.315 $Y=2.105
+ $X2=1.315 $Y2=2.36
r187 29 56 3.22182 $w=2.92e-07 $l=8.5e-08 $layer=LI1_cond $X=1.397 $Y=1.935
+ $X2=1.397 $Y2=2.02
r188 29 31 34.7269 $w=3.73e-07 $l=1.13e-06 $layer=LI1_cond $X=1.397 $Y=1.935
+ $X2=1.397 $Y2=0.805
r189 27 46 47.1618 $w=3.75e-07 $l=3.18e-07 $layer=POLY_cond $X=2.862 $Y=1.868
+ $X2=2.862 $Y2=1.55
r190 27 28 48.4185 $w=3.75e-07 $l=1.87e-07 $layer=POLY_cond $X=2.862 $Y=1.868
+ $X2=2.862 $Y2=2.055
r191 26 46 2.22462 $w=3.75e-07 $l=1.5e-08 $layer=POLY_cond $X=2.862 $Y=1.535
+ $X2=2.862 $Y2=1.55
r192 25 26 42.9311 $w=3.75e-07 $l=1.5e-07 $layer=POLY_cond $X=2.93 $Y=1.385
+ $X2=2.93 $Y2=1.535
r193 21 23 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=5.74 $Y=1.785
+ $X2=5.74 $Y2=2.105
r194 20 60 51.2425 $w=3.01e-07 $l=4.20666e-07 $layer=POLY_cond $X=5.41 $Y=1.71
+ $X2=5.177 $Y2=1.39
r195 19 21 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.665 $Y=1.71
+ $X2=5.74 $Y2=1.785
r196 19 20 130.755 $w=1.5e-07 $l=2.55e-07 $layer=POLY_cond $X=5.665 $Y=1.71
+ $X2=5.41 $Y2=1.71
r197 15 60 38.5481 $w=3.01e-07 $l=2.30499e-07 $layer=POLY_cond $X=5.02 $Y=1.225
+ $X2=5.177 $Y2=1.39
r198 15 17 215.362 $w=1.5e-07 $l=4.2e-07 $layer=POLY_cond $X=5.02 $Y=1.225
+ $X2=5.02 $Y2=0.805
r199 13 25 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=3.11 $Y=0.805
+ $X2=3.11 $Y2=1.385
r200 9 28 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=2.75 $Y=2.425
+ $X2=2.75 $Y2=2.055
r201 2 35 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=1.2
+ $Y=2.215 $X2=1.325 $Y2=2.36
r202 1 31 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=1.295
+ $Y=0.595 $X2=1.42 $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_LP__DFXTP_2%A_679_93# 1 2 9 13 17 20 21 22 24 31
c64 17 0 9.35787e-20 $X=3.77 $Y=1.57
c65 13 0 4.80136e-20 $X=3.81 $Y=2.425
r66 22 27 3.33156 $w=2.1e-07 $l=1.0247e-07 $layer=LI1_cond $X=4.7 $Y=1.915
+ $X2=4.705 $Y2=2.015
r67 22 24 61.5281 $w=2.08e-07 $l=1.165e-06 $layer=LI1_cond $X=4.7 $Y=1.915
+ $X2=4.7 $Y2=0.75
r68 20 27 3.49021 $w=2e-07 $l=1.1e-07 $layer=LI1_cond $X=4.595 $Y=2.015
+ $X2=4.705 $Y2=2.015
r69 20 21 36.6 $w=1.98e-07 $l=6.6e-07 $layer=LI1_cond $X=4.595 $Y=2.015
+ $X2=3.935 $Y2=2.015
r70 18 31 6.99445 $w=3.3e-07 $l=4e-08 $layer=POLY_cond $X=3.77 $Y=1.57 $X2=3.81
+ $Y2=1.57
r71 18 28 52.4584 $w=3.3e-07 $l=3e-07 $layer=POLY_cond $X=3.77 $Y=1.57 $X2=3.47
+ $Y2=1.57
r72 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.77
+ $Y=1.57 $X2=3.77 $Y2=1.57
r73 15 21 7.36389 $w=2e-07 $l=2.09105e-07 $layer=LI1_cond $X=3.77 $Y=1.915
+ $X2=3.935 $Y2=2.015
r74 15 17 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=3.77 $Y=1.915
+ $X2=3.77 $Y2=1.57
r75 11 31 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.81 $Y=1.735
+ $X2=3.81 $Y2=1.57
r76 11 13 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.81 $Y=1.735
+ $X2=3.81 $Y2=2.425
r77 7 28 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.47 $Y=1.405
+ $X2=3.47 $Y2=1.57
r78 7 9 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=3.47 $Y=1.405 $X2=3.47
+ $Y2=0.805
r79 2 27 600 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=4.51
+ $Y=1.895 $X2=4.65 $Y2=2.02
r80 1 24 91 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=2 $X=4.57
+ $Y=0.595 $X2=4.71 $Y2=0.75
.ends

.subckt PM_SKY130_FD_SC_LP__DFXTP_2%A_551_119# 1 2 9 13 16 18 19 22 23 29
c65 22 0 1.61944e-19 $X=4.34 $Y=1.51
c66 19 0 1.7508e-19 $X=3.35 $Y=1.14
r67 26 27 12.341 $w=3.46e-07 $l=3.5e-07 $layer=LI1_cond $X=2.895 $Y=0.932
+ $X2=3.245 $Y2=0.932
r68 23 30 45.5639 $w=3.95e-07 $l=1.65e-07 $layer=POLY_cond $X=4.372 $Y=1.51
+ $X2=4.372 $Y2=1.675
r69 23 29 45.5639 $w=3.95e-07 $l=1.65e-07 $layer=POLY_cond $X=4.372 $Y=1.51
+ $X2=4.372 $Y2=1.345
r70 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.34
+ $Y=1.51 $X2=4.34 $Y2=1.51
r71 20 22 13.1378 $w=2.48e-07 $l=2.85e-07 $layer=LI1_cond $X=4.3 $Y=1.225
+ $X2=4.3 $Y2=1.51
r72 19 27 6.86265 $w=3.46e-07 $l=2.55155e-07 $layer=LI1_cond $X=3.35 $Y=1.14
+ $X2=3.245 $Y2=0.932
r73 18 20 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=4.175 $Y=1.14
+ $X2=4.3 $Y2=1.225
r74 18 19 53.8235 $w=1.68e-07 $l=8.25e-07 $layer=LI1_cond $X=4.175 $Y=1.14
+ $X2=3.35 $Y2=1.14
r75 14 27 3.65847 $w=2.1e-07 $l=2.93e-07 $layer=LI1_cond $X=3.245 $Y=1.225
+ $X2=3.245 $Y2=0.932
r76 14 16 63.3766 $w=2.08e-07 $l=1.2e-06 $layer=LI1_cond $X=3.245 $Y=1.225
+ $X2=3.245 $Y2=2.425
r77 13 29 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=4.495 $Y=0.915
+ $X2=4.495 $Y2=1.345
r78 9 30 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=4.435 $Y=2.315
+ $X2=4.435 $Y2=1.675
r79 2 16 600 $w=1.7e-07 $l=5.04182e-07 $layer=licon1_PDIFF $count=1 $X=2.825
+ $Y=2.215 $X2=3.235 $Y2=2.425
r80 1 26 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.755
+ $Y=0.595 $X2=2.895 $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_LP__DFXTP_2%A_110_62# 1 2 7 8 12 16 17 18 19 20 23 25 29
+ 31 35 39 43 45 46 48 52
c129 35 0 6.46168e-20 $X=4.945 $Y=2.315
c130 23 0 3.84473e-21 $X=2.68 $Y=0.805
r131 51 54 29.7822 $w=4.43e-07 $l=1.15e-06 $layer=LI1_cond $X=0.817 $Y=1.395
+ $X2=0.817 $Y2=2.545
r132 51 52 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.955
+ $Y=1.395 $X2=0.955 $Y2=1.395
r133 48 51 23.3078 $w=4.43e-07 $l=9e-07 $layer=LI1_cond $X=0.817 $Y=0.495
+ $X2=0.817 $Y2=1.395
r134 42 43 58.9681 $w=1.5e-07 $l=1.15e-07 $layer=POLY_cond $X=1.54 $Y=1.305
+ $X2=1.655 $Y2=1.305
r135 41 52 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=0.955 $Y=1.38
+ $X2=0.955 $Y2=1.395
r136 37 39 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=5.59 $Y=0.255
+ $X2=5.59 $Y2=0.805
r137 33 35 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=4.945 $Y=3.075
+ $X2=4.945 $Y2=2.315
r138 32 46 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.525 $Y=3.15
+ $X2=3.45 $Y2=3.15
r139 31 33 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.87 $Y=3.15
+ $X2=4.945 $Y2=3.075
r140 31 32 689.67 $w=1.5e-07 $l=1.345e-06 $layer=POLY_cond $X=4.87 $Y=3.15
+ $X2=3.525 $Y2=3.15
r141 27 46 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.45 $Y=3.075
+ $X2=3.45 $Y2=3.15
r142 27 29 333.298 $w=1.5e-07 $l=6.5e-07 $layer=POLY_cond $X=3.45 $Y=3.075
+ $X2=3.45 $Y2=2.425
r143 26 45 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.755 $Y=0.18
+ $X2=2.68 $Y2=0.18
r144 25 37 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.515 $Y=0.18
+ $X2=5.59 $Y2=0.255
r145 25 26 1415.23 $w=1.5e-07 $l=2.76e-06 $layer=POLY_cond $X=5.515 $Y=0.18
+ $X2=2.755 $Y2=0.18
r146 21 45 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.68 $Y=0.255
+ $X2=2.68 $Y2=0.18
r147 21 23 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=2.68 $Y=0.255
+ $X2=2.68 $Y2=0.805
r148 19 45 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.605 $Y=0.18
+ $X2=2.68 $Y2=0.18
r149 19 20 448.67 $w=1.5e-07 $l=8.75e-07 $layer=POLY_cond $X=2.605 $Y=0.18
+ $X2=1.73 $Y2=0.18
r150 17 46 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.375 $Y=3.15
+ $X2=3.45 $Y2=3.15
r151 17 18 902.468 $w=1.5e-07 $l=1.76e-06 $layer=POLY_cond $X=3.375 $Y=3.15
+ $X2=1.615 $Y2=3.15
r152 14 43 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.655 $Y=1.23
+ $X2=1.655 $Y2=1.305
r153 14 16 217.926 $w=1.5e-07 $l=4.25e-07 $layer=POLY_cond $X=1.655 $Y=1.23
+ $X2=1.655 $Y2=0.805
r154 13 20 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.655 $Y=0.255
+ $X2=1.73 $Y2=0.18
r155 13 16 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=1.655 $Y=0.255
+ $X2=1.655 $Y2=0.805
r156 10 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.54 $Y=3.075
+ $X2=1.615 $Y2=3.15
r157 10 12 276.894 $w=1.5e-07 $l=5.4e-07 $layer=POLY_cond $X=1.54 $Y=3.075
+ $X2=1.54 $Y2=2.535
r158 9 42 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.54 $Y=1.38
+ $X2=1.54 $Y2=1.305
r159 9 12 592.245 $w=1.5e-07 $l=1.155e-06 $layer=POLY_cond $X=1.54 $Y=1.38
+ $X2=1.54 $Y2=2.535
r160 8 41 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=1.12 $Y=1.305
+ $X2=0.955 $Y2=1.38
r161 7 42 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.465 $Y=1.305
+ $X2=1.54 $Y2=1.305
r162 7 8 176.904 $w=1.5e-07 $l=3.45e-07 $layer=POLY_cond $X=1.465 $Y=1.305
+ $X2=1.12 $Y2=1.305
r163 2 54 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=0.55
+ $Y=2.4 $X2=0.69 $Y2=2.545
r164 1 48 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.31 $X2=0.69 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__DFXTP_2%A_1175_93# 1 2 9 11 13 15 17 20 22 24 26 29
+ 31 32 33 34 38 41 43 49 53
c96 31 0 1.00884e-19 $X=7.63 $Y=1.51
c97 9 0 6.87636e-20 $X=5.95 $Y=0.805
r98 55 56 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.27
+ $Y=1.51 $X2=7.27 $Y2=1.51
r99 53 55 9.61826 $w=2.41e-07 $l=1.9e-07 $layer=LI1_cond $X=7.08 $Y=1.615
+ $X2=7.27 $Y2=1.615
r100 49 51 15.9138 $w=4.73e-07 $l=4.25e-07 $layer=LI1_cond $X=6.927 $Y=0.52
+ $X2=6.927 $Y2=0.945
r101 43 46 5.5876 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=6.19 $Y=1.56
+ $X2=6.19 $Y2=1.72
r102 43 44 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.19
+ $Y=1.56 $X2=6.19 $Y2=1.56
r103 41 53 2.78154 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=7.08 $Y=1.425
+ $X2=7.08 $Y2=1.615
r104 41 51 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=7.08 $Y=1.425
+ $X2=7.08 $Y2=0.945
r105 36 53 6.22656 $w=2.41e-07 $l=2.43865e-07 $layer=LI1_cond $X=6.957 $Y=1.805
+ $X2=7.08 $Y2=1.615
r106 36 38 6.52588 $w=4.13e-07 $l=2.35e-07 $layer=LI1_cond $X=6.957 $Y=1.805
+ $X2=6.957 $Y2=2.04
r107 35 46 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.355 $Y=1.72
+ $X2=6.19 $Y2=1.72
r108 34 36 11.5531 $w=2.41e-07 $l=2.45854e-07 $layer=LI1_cond $X=6.75 $Y=1.72
+ $X2=6.957 $Y2=1.805
r109 34 35 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=6.75 $Y=1.72
+ $X2=6.355 $Y2=1.72
r110 31 56 62.9501 $w=3.3e-07 $l=3.6e-07 $layer=POLY_cond $X=7.63 $Y=1.51
+ $X2=7.27 $Y2=1.51
r111 31 32 6.91837 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=7.63 $Y=1.51
+ $X2=7.705 $Y2=1.51
r112 27 33 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.135 $Y=1.495
+ $X2=8.135 $Y2=1.42
r113 27 29 497.383 $w=1.5e-07 $l=9.7e-07 $layer=POLY_cond $X=8.135 $Y=1.495
+ $X2=8.135 $Y2=2.465
r114 24 33 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.135 $Y=1.345
+ $X2=8.135 $Y2=1.42
r115 24 26 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=8.135 $Y=1.345
+ $X2=8.135 $Y2=0.815
r116 23 32 6.91837 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=7.78 $Y=1.42
+ $X2=7.705 $Y2=1.51
r117 22 33 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.06 $Y=1.42
+ $X2=8.135 $Y2=1.42
r118 22 23 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=8.06 $Y=1.42
+ $X2=7.78 $Y2=1.42
r119 18 32 18.1359 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.705 $Y=1.675
+ $X2=7.705 $Y2=1.51
r120 18 20 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=7.705 $Y=1.675
+ $X2=7.705 $Y2=2.465
r121 15 32 18.1359 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.705 $Y=1.345
+ $X2=7.705 $Y2=1.51
r122 15 17 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=7.705 $Y=1.345
+ $X2=7.705 $Y2=0.815
r123 11 44 39.1513 $w=3.76e-07 $l=1.72337e-07 $layer=POLY_cond $X=6.1 $Y=1.725
+ $X2=6.115 $Y2=1.56
r124 11 13 194.851 $w=1.5e-07 $l=3.8e-07 $layer=POLY_cond $X=6.1 $Y=1.725
+ $X2=6.1 $Y2=2.105
r125 7 44 58.38 $w=3.76e-07 $l=3.88844e-07 $layer=POLY_cond $X=5.95 $Y=1.245
+ $X2=6.115 $Y2=1.56
r126 7 9 225.617 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=5.95 $Y=1.245
+ $X2=5.95 $Y2=0.805
r127 2 38 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=6.715
+ $Y=1.895 $X2=6.855 $Y2=2.04
r128 1 49 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.715
+ $Y=0.375 $X2=6.855 $Y2=0.52
.ends

.subckt PM_SKY130_FD_SC_LP__DFXTP_2%A_1004_379# 1 2 9 12 14 16 20 22 27 28 32 35
c75 28 0 1.69648e-19 $X=6.695 $Y=1.21
r76 32 36 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.73 $Y=1.29
+ $X2=6.73 $Y2=1.455
r77 32 35 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.73 $Y=1.29
+ $X2=6.73 $Y2=1.125
r78 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.73
+ $Y=1.29 $X2=6.73 $Y2=1.29
r79 28 31 3.54598 $w=2.58e-07 $l=8e-08 $layer=LI1_cond $X=6.695 $Y=1.21
+ $X2=6.695 $Y2=1.29
r80 23 25 11.5914 $w=4.21e-07 $l=5.11859e-07 $layer=LI1_cond $X=5.655 $Y=1.21
+ $X2=5.4 $Y2=0.81
r81 22 28 3.22376 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=6.565 $Y=1.21
+ $X2=6.695 $Y2=1.21
r82 22 23 59.369 $w=1.68e-07 $l=9.1e-07 $layer=LI1_cond $X=6.565 $Y=1.21
+ $X2=5.655 $Y2=1.21
r83 20 23 6.93546 $w=4.21e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.57 $Y=1.295
+ $X2=5.655 $Y2=1.21
r84 20 27 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=5.57 $Y=1.295
+ $X2=5.57 $Y2=1.875
r85 16 18 19.8076 $w=3.18e-07 $l=5.5e-07 $layer=LI1_cond $X=5.495 $Y=2.04
+ $X2=5.495 $Y2=2.59
r86 14 27 8.28018 $w=3.18e-07 $l=1.6e-07 $layer=LI1_cond $X=5.495 $Y=2.035
+ $X2=5.495 $Y2=1.875
r87 14 16 0.180069 $w=3.18e-07 $l=5e-09 $layer=LI1_cond $X=5.495 $Y=2.035
+ $X2=5.495 $Y2=2.04
r88 12 36 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=6.64 $Y=2.315
+ $X2=6.64 $Y2=1.455
r89 9 35 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=6.64 $Y=0.695
+ $X2=6.64 $Y2=1.125
r90 2 18 600 $w=1.7e-07 $l=8.76342e-07 $layer=licon1_PDIFF $count=1 $X=5.02
+ $Y=1.895 $X2=5.43 $Y2=2.59
r91 2 16 600 $w=1.7e-07 $l=4.77022e-07 $layer=licon1_PDIFF $count=1 $X=5.02
+ $Y=1.895 $X2=5.43 $Y2=2.04
r92 1 25 182 $w=1.7e-07 $l=3.04056e-07 $layer=licon1_NDIFF $count=1 $X=5.095
+ $Y=0.595 $X2=5.31 $Y2=0.81
.ends

.subckt PM_SKY130_FD_SC_LP__DFXTP_2%VPWR 1 2 3 4 5 6 19 21 25 29 33 39 43 45 50
+ 51 52 54 59 74 78 87 90 93 97
r100 96 97 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=3.33 $X2=8.4
+ $Y2=3.33
r101 93 94 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r102 90 91 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r103 87 88 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r104 84 85 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r105 82 97 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=8.4 $Y2=3.33
r106 82 94 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=7.44 $Y2=3.33
r107 81 82 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r108 79 93 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=7.615 $Y=3.33
+ $X2=7.475 $Y2=3.33
r109 79 81 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=7.615 $Y=3.33
+ $X2=7.92 $Y2=3.33
r110 78 96 3.8143 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=8.22 $Y=3.33 $X2=8.43
+ $Y2=3.33
r111 78 81 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=8.22 $Y=3.33 $X2=7.92
+ $Y2=3.33
r112 77 94 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=7.44 $Y2=3.33
r113 76 77 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r114 74 93 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=7.335 $Y=3.33
+ $X2=7.475 $Y2=3.33
r115 74 76 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=7.335 $Y=3.33
+ $X2=6.96 $Y2=3.33
r116 73 77 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=6.96
+ $Y2=3.33
r117 72 73 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r118 70 73 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=6 $Y2=3.33
r119 69 72 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=4.56 $Y=3.33 $X2=6
+ $Y2=3.33
r120 69 70 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r121 67 90 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.305 $Y=3.33
+ $X2=4.14 $Y2=3.33
r122 67 69 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=4.305 $Y=3.33
+ $X2=4.56 $Y2=3.33
r123 66 91 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r124 65 66 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r125 63 66 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.6 $Y2=3.33
r126 63 88 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r127 62 65 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=2.16 $Y=3.33
+ $X2=3.6 $Y2=3.33
r128 62 63 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r129 60 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.92 $Y=3.33
+ $X2=1.755 $Y2=3.33
r130 60 62 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=1.92 $Y=3.33
+ $X2=2.16 $Y2=3.33
r131 59 90 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.975 $Y=3.33
+ $X2=4.14 $Y2=3.33
r132 59 65 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=3.975 $Y=3.33
+ $X2=3.6 $Y2=3.33
r133 58 88 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r134 58 85 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.24 $Y2=3.33
r135 57 58 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r136 55 84 4.78091 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=3.33
+ $X2=0.212 $Y2=3.33
r137 55 57 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=0.425 $Y=3.33
+ $X2=1.2 $Y2=3.33
r138 54 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.59 $Y=3.33
+ $X2=1.755 $Y2=3.33
r139 54 57 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=1.59 $Y=3.33
+ $X2=1.2 $Y2=3.33
r140 52 70 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.32 $Y=3.33
+ $X2=4.56 $Y2=3.33
r141 52 91 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.32 $Y=3.33
+ $X2=4.08 $Y2=3.33
r142 50 72 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=6.15 $Y=3.33 $X2=6
+ $Y2=3.33
r143 50 51 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=6.15 $Y=3.33
+ $X2=6.34 $Y2=3.33
r144 49 76 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=6.53 $Y=3.33
+ $X2=6.96 $Y2=3.33
r145 49 51 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=6.53 $Y=3.33
+ $X2=6.34 $Y2=3.33
r146 45 48 47.5689 $w=2.33e-07 $l=9.7e-07 $layer=LI1_cond $X=8.337 $Y=1.98
+ $X2=8.337 $Y2=2.95
r147 43 96 3.23307 $w=2.35e-07 $l=1.28662e-07 $layer=LI1_cond $X=8.337 $Y=3.245
+ $X2=8.43 $Y2=3.33
r148 43 48 14.4668 $w=2.33e-07 $l=2.95e-07 $layer=LI1_cond $X=8.337 $Y=3.245
+ $X2=8.337 $Y2=2.95
r149 39 42 39.9239 $w=2.78e-07 $l=9.7e-07 $layer=LI1_cond $X=7.475 $Y=1.98
+ $X2=7.475 $Y2=2.95
r150 37 93 0.375625 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=7.475 $Y=3.245
+ $X2=7.475 $Y2=3.33
r151 37 42 12.1418 $w=2.78e-07 $l=2.95e-07 $layer=LI1_cond $X=7.475 $Y=3.245
+ $X2=7.475 $Y2=2.95
r152 33 36 14.7088 $w=3.78e-07 $l=4.85e-07 $layer=LI1_cond $X=6.34 $Y=2.105
+ $X2=6.34 $Y2=2.59
r153 31 51 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=6.34 $Y=3.245
+ $X2=6.34 $Y2=3.33
r154 31 36 19.8645 $w=3.78e-07 $l=6.55e-07 $layer=LI1_cond $X=6.34 $Y=3.245
+ $X2=6.34 $Y2=2.59
r155 27 90 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.14 $Y=3.245
+ $X2=4.14 $Y2=3.33
r156 27 29 18.3343 $w=3.28e-07 $l=5.25e-07 $layer=LI1_cond $X=4.14 $Y=3.245
+ $X2=4.14 $Y2=2.72
r157 23 87 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.755 $Y=3.245
+ $X2=1.755 $Y2=3.33
r158 23 25 29.8588 $w=3.28e-07 $l=8.55e-07 $layer=LI1_cond $X=1.755 $Y=3.245
+ $X2=1.755 $Y2=2.39
r159 19 84 2.98526 $w=3.3e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.26 $Y=3.245
+ $X2=0.212 $Y2=3.33
r160 19 21 16.0644 $w=3.28e-07 $l=4.6e-07 $layer=LI1_cond $X=0.26 $Y=3.245
+ $X2=0.26 $Y2=2.785
r161 6 48 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=8.21
+ $Y=1.835 $X2=8.35 $Y2=2.95
r162 6 45 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=8.21
+ $Y=1.835 $X2=8.35 $Y2=1.98
r163 5 42 400 $w=1.7e-07 $l=1.17584e-06 $layer=licon1_PDIFF $count=1 $X=7.365
+ $Y=1.835 $X2=7.49 $Y2=2.95
r164 5 39 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=7.365
+ $Y=1.835 $X2=7.49 $Y2=1.98
r165 4 36 600 $w=1.7e-07 $l=8.10417e-07 $layer=licon1_PDIFF $count=1 $X=6.175
+ $Y=1.895 $X2=6.425 $Y2=2.59
r166 4 33 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=6.175
+ $Y=1.895 $X2=6.315 $Y2=2.105
r167 3 29 600 $w=1.7e-07 $l=6.19516e-07 $layer=licon1_PDIFF $count=1 $X=3.885
+ $Y=2.215 $X2=4.14 $Y2=2.72
r168 2 25 300 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_PDIFF $count=2 $X=1.615
+ $Y=2.215 $X2=1.755 $Y2=2.39
r169 1 21 600 $w=1.7e-07 $l=4.43114e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.4 $X2=0.26 $Y2=2.785
.ends

.subckt PM_SKY130_FD_SC_LP__DFXTP_2%A_432_119# 1 2 9 11 16 18
c27 9 0 1.7508e-19 $X=2.535 $Y=1.315
r28 14 16 4.88915 $w=3.28e-07 $l=1.4e-07 $layer=LI1_cond $X=2.39 $Y=0.805
+ $X2=2.53 $Y2=0.805
r29 9 18 5.58789 $w=1.88e-07 $l=9.5e-08 $layer=LI1_cond $X=2.535 $Y=1.315
+ $X2=2.535 $Y2=1.22
r30 9 11 64.7943 $w=1.88e-07 $l=1.11e-06 $layer=LI1_cond $X=2.535 $Y=1.315
+ $X2=2.535 $Y2=2.425
r31 7 16 4.28565 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=2.53 $Y=0.97 $X2=2.53
+ $Y2=0.805
r32 7 18 15.404 $w=1.78e-07 $l=2.5e-07 $layer=LI1_cond $X=2.53 $Y=0.97 $X2=2.53
+ $Y2=1.22
r33 2 11 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=2.395
+ $Y=2.215 $X2=2.535 $Y2=2.425
r34 1 14 182 $w=1.7e-07 $l=3.18119e-07 $layer=licon1_NDIFF $count=1 $X=2.16
+ $Y=0.595 $X2=2.39 $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_LP__DFXTP_2%Q 1 2 7 8 9 10 11 12 13
r19 13 39 5.87094 $w=2.63e-07 $l=1.35e-07 $layer=LI1_cond $X=7.917 $Y=2.775
+ $X2=7.917 $Y2=2.91
r20 12 13 16.0907 $w=2.63e-07 $l=3.7e-07 $layer=LI1_cond $X=7.917 $Y=2.405
+ $X2=7.917 $Y2=2.775
r21 11 12 16.9605 $w=2.63e-07 $l=3.9e-07 $layer=LI1_cond $X=7.917 $Y=2.015
+ $X2=7.917 $Y2=2.405
r22 10 11 15.2209 $w=2.63e-07 $l=3.5e-07 $layer=LI1_cond $X=7.917 $Y=1.665
+ $X2=7.917 $Y2=2.015
r23 9 10 16.0907 $w=2.63e-07 $l=3.7e-07 $layer=LI1_cond $X=7.917 $Y=1.295
+ $X2=7.917 $Y2=1.665
r24 8 9 16.0907 $w=2.63e-07 $l=3.7e-07 $layer=LI1_cond $X=7.917 $Y=0.925
+ $X2=7.917 $Y2=1.295
r25 7 8 16.743 $w=2.63e-07 $l=3.85e-07 $layer=LI1_cond $X=7.917 $Y=0.54
+ $X2=7.917 $Y2=0.925
r26 2 39 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=7.78
+ $Y=1.835 $X2=7.92 $Y2=2.91
r27 2 11 400 $w=1.7e-07 $l=2.4e-07 $layer=licon1_PDIFF $count=1 $X=7.78 $Y=1.835
+ $X2=7.92 $Y2=2.015
r28 1 7 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=7.78
+ $Y=0.395 $X2=7.92 $Y2=0.54
.ends

.subckt PM_SKY130_FD_SC_LP__DFXTP_2%VGND 1 2 3 4 5 6 19 21 25 29 33 35 37 40 41
+ 42 51 55 60 65 83 86 90
c91 3 0 1.61944e-19 $X=3.545 $Y=0.595
r92 89 90 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r93 86 87 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r94 83 84 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=0 $X2=6 $Y2=0
r95 76 78 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r96 71 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r97 69 90 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=8.4
+ $Y2=0
r98 69 87 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=7.44
+ $Y2=0
r99 68 69 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r100 66 86 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=7.615 $Y=0 $X2=7.475
+ $Y2=0
r101 66 68 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=7.615 $Y=0
+ $X2=7.92 $Y2=0
r102 65 89 3.8143 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=8.22 $Y=0 $X2=8.43
+ $Y2=0
r103 65 68 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=8.22 $Y=0 $X2=7.92
+ $Y2=0
r104 64 87 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=7.44
+ $Y2=0
r105 64 84 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=6
+ $Y2=0
r106 63 64 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r107 61 83 11.5608 $w=1.7e-07 $l=2.6e-07 $layer=LI1_cond $X=6.52 $Y=0 $X2=6.26
+ $Y2=0
r108 61 63 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=6.52 $Y=0 $X2=6.96
+ $Y2=0
r109 60 86 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=7.335 $Y=0 $X2=7.475
+ $Y2=0
r110 60 63 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=7.335 $Y=0
+ $X2=6.96 $Y2=0
r111 59 84 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=4.56 $Y=0 $X2=6
+ $Y2=0
r112 58 59 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r113 56 58 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=4.425 $Y=0
+ $X2=4.56 $Y2=0
r114 55 83 11.5608 $w=1.7e-07 $l=2.6e-07 $layer=LI1_cond $X=6 $Y=0 $X2=6.26
+ $Y2=0
r115 55 58 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=6 $Y=0 $X2=4.56
+ $Y2=0
r116 54 76 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.6
+ $Y2=0
r117 53 54 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r118 51 80 10.3801 $w=9.03e-07 $l=7.7e-07 $layer=LI1_cond $X=3.972 $Y=0
+ $X2=3.972 $Y2=0.77
r119 51 56 11.0417 $w=1.7e-07 $l=4.53e-07 $layer=LI1_cond $X=3.972 $Y=0
+ $X2=4.425 $Y2=0
r120 51 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r121 51 76 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r122 51 53 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=3.52 $Y=0 $X2=2.16
+ $Y2=0
r123 50 54 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r124 49 50 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r125 47 50 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r126 47 72 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r127 46 49 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r128 46 47 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r129 44 71 4.78091 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=0
+ $X2=0.212 $Y2=0
r130 44 46 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.425 $Y=0 $X2=0.72
+ $Y2=0
r131 42 59 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.32 $Y=0
+ $X2=4.56 $Y2=0
r132 42 78 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.32 $Y=0
+ $X2=4.08 $Y2=0
r133 40 49 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=1.755 $Y=0 $X2=1.68
+ $Y2=0
r134 40 41 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=1.755 $Y=0 $X2=1.895
+ $Y2=0
r135 39 53 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=2.035 $Y=0
+ $X2=2.16 $Y2=0
r136 39 41 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=2.035 $Y=0 $X2=1.895
+ $Y2=0
r137 35 89 3.23307 $w=2.35e-07 $l=1.28662e-07 $layer=LI1_cond $X=8.337 $Y=0.085
+ $X2=8.43 $Y2=0
r138 35 37 22.3133 $w=2.33e-07 $l=4.55e-07 $layer=LI1_cond $X=8.337 $Y=0.085
+ $X2=8.337 $Y2=0.54
r139 31 86 0.375625 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=7.475 $Y=0.085
+ $X2=7.475 $Y2=0
r140 31 33 18.7272 $w=2.78e-07 $l=4.55e-07 $layer=LI1_cond $X=7.475 $Y=0.085
+ $X2=7.475 $Y2=0.54
r141 27 83 2.17428 $w=5.2e-07 $l=8.5e-08 $layer=LI1_cond $X=6.26 $Y=0.085
+ $X2=6.26 $Y2=0
r142 27 29 9.54563 $w=5.18e-07 $l=4.15e-07 $layer=LI1_cond $X=6.26 $Y=0.085
+ $X2=6.26 $Y2=0.5
r143 23 41 0.375625 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=1.895 $Y=0.085
+ $X2=1.895 $Y2=0
r144 23 25 29.6342 $w=2.78e-07 $l=7.2e-07 $layer=LI1_cond $X=1.895 $Y=0.085
+ $X2=1.895 $Y2=0.805
r145 19 71 2.98526 $w=3.3e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.212 $Y2=0
r146 19 21 15.1913 $w=3.28e-07 $l=4.35e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.26 $Y2=0.52
r147 6 37 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=8.21
+ $Y=0.395 $X2=8.35 $Y2=0.54
r148 5 33 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=7.365
+ $Y=0.395 $X2=7.49 $Y2=0.54
r149 4 29 91 $w=1.7e-07 $l=4.44972e-07 $layer=licon1_NDIFF $count=2 $X=6.025
+ $Y=0.595 $X2=6.425 $Y2=0.5
r150 3 80 91 $w=1.7e-07 $l=7.97716e-07 $layer=licon1_NDIFF $count=2 $X=3.545
+ $Y=0.595 $X2=4.26 $Y2=0.77
r151 2 25 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.73
+ $Y=0.595 $X2=1.87 $Y2=0.805
r152 1 21 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.31 $X2=0.26 $Y2=0.52
.ends

