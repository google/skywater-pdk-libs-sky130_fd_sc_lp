* File: sky130_fd_sc_lp__nor4_2.pxi.spice
* Created: Wed Sep  2 10:10:25 2020
* 
x_PM_SKY130_FD_SC_LP__NOR4_2%B N_B_M1003_g N_B_M1007_g N_B_M1004_g N_B_M1015_g
+ N_B_c_86_n N_B_c_87_n N_B_c_88_n N_B_c_97_n N_B_c_89_n B B N_B_c_91_n
+ PM_SKY130_FD_SC_LP__NOR4_2%B
x_PM_SKY130_FD_SC_LP__NOR4_2%A N_A_c_164_n N_A_M1010_g N_A_M1000_g N_A_c_166_n
+ N_A_M1014_g N_A_M1005_g A N_A_c_169_n PM_SKY130_FD_SC_LP__NOR4_2%A
x_PM_SKY130_FD_SC_LP__NOR4_2%C N_C_M1011_g N_C_M1001_g N_C_M1012_g N_C_M1009_g
+ N_C_c_222_n N_C_c_216_n C C N_C_c_219_n N_C_c_227_n
+ PM_SKY130_FD_SC_LP__NOR4_2%C
x_PM_SKY130_FD_SC_LP__NOR4_2%D N_D_c_308_n N_D_M1002_g N_D_M1006_g N_D_c_310_n
+ N_D_M1013_g N_D_M1008_g D N_D_c_313_n PM_SKY130_FD_SC_LP__NOR4_2%D
x_PM_SKY130_FD_SC_LP__NOR4_2%A_74_367# N_A_74_367#_M1007_s N_A_74_367#_M1015_s
+ N_A_74_367#_M1009_d N_A_74_367#_c_362_n N_A_74_367#_c_363_n
+ N_A_74_367#_c_368_n N_A_74_367#_c_373_n N_A_74_367#_c_382_n
+ N_A_74_367#_c_364_n N_A_74_367#_c_365_n PM_SKY130_FD_SC_LP__NOR4_2%A_74_367#
x_PM_SKY130_FD_SC_LP__NOR4_2%A_157_367# N_A_157_367#_M1007_d
+ N_A_157_367#_M1005_s N_A_157_367#_c_412_n N_A_157_367#_c_417_n
+ N_A_157_367#_c_418_n PM_SKY130_FD_SC_LP__NOR4_2%A_157_367#
x_PM_SKY130_FD_SC_LP__NOR4_2%VPWR N_VPWR_M1000_d N_VPWR_c_428_n VPWR
+ N_VPWR_c_429_n N_VPWR_c_430_n N_VPWR_c_427_n N_VPWR_c_432_n
+ PM_SKY130_FD_SC_LP__NOR4_2%VPWR
x_PM_SKY130_FD_SC_LP__NOR4_2%A_553_367# N_A_553_367#_M1001_s
+ N_A_553_367#_M1008_s N_A_553_367#_c_476_n N_A_553_367#_c_478_n
+ N_A_553_367#_c_479_n PM_SKY130_FD_SC_LP__NOR4_2%A_553_367#
x_PM_SKY130_FD_SC_LP__NOR4_2%Y N_Y_M1003_s N_Y_M1014_s N_Y_M1011_s N_Y_M1013_d
+ N_Y_M1006_d N_Y_c_572_p N_Y_c_505_n N_Y_c_506_n N_Y_c_508_n N_Y_c_496_n
+ N_Y_c_530_n N_Y_c_531_n N_Y_c_502_n N_Y_c_582_p N_Y_c_497_n N_Y_c_498_n
+ N_Y_c_499_n N_Y_c_542_n N_Y_c_500_n Y Y Y PM_SKY130_FD_SC_LP__NOR4_2%Y
x_PM_SKY130_FD_SC_LP__NOR4_2%VGND N_VGND_M1003_d N_VGND_M1010_d N_VGND_M1004_d
+ N_VGND_M1002_s N_VGND_M1012_d N_VGND_c_593_n N_VGND_c_594_n N_VGND_c_595_n
+ N_VGND_c_596_n N_VGND_c_597_n N_VGND_c_598_n N_VGND_c_599_n N_VGND_c_600_n
+ N_VGND_c_601_n N_VGND_c_602_n VGND N_VGND_c_603_n N_VGND_c_604_n
+ N_VGND_c_605_n N_VGND_c_606_n N_VGND_c_607_n N_VGND_c_608_n N_VGND_c_609_n
+ PM_SKY130_FD_SC_LP__NOR4_2%VGND
cc_1 VNB N_B_M1003_g 0.0349222f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=0.655
cc_2 VNB N_B_M1004_g 0.0258008f $X=-0.19 $Y=-0.245 $X2=2 $Y2=0.655
cc_3 VNB N_B_c_86_n 0.0360695f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.51
cc_4 VNB N_B_c_87_n 0.009048f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=1.51
cc_5 VNB N_B_c_88_n 0.00815588f $X=-0.19 $Y=-0.245 $X2=1.855 $Y2=1.7
cc_6 VNB N_B_c_89_n 0.0251325f $X=-0.19 $Y=-0.245 $X2=2.02 $Y2=1.51
cc_7 VNB B 0.0177963f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_8 VNB N_B_c_91_n 0.00375608f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=1.565
cc_9 VNB N_A_c_164_n 0.0162354f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=1.345
cc_10 VNB N_A_M1000_g 0.00687258f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=2.465
cc_11 VNB N_A_c_166_n 0.0155954f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_M1005_g 0.00648038f $X=-0.19 $Y=-0.245 $X2=2 $Y2=1.675
cc_13 VNB A 0.00282816f $X=-0.19 $Y=-0.245 $X2=2 $Y2=2.465
cc_14 VNB N_A_c_169_n 0.0357054f $X=-0.19 $Y=-0.245 $X2=2.02 $Y2=1.51
cc_15 VNB N_C_M1011_g 0.0258152f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=0.655
cc_16 VNB N_C_M1012_g 0.0281753f $X=-0.19 $Y=-0.245 $X2=2 $Y2=0.655
cc_17 VNB N_C_c_216_n 0.0281896f $X=-0.19 $Y=-0.245 $X2=2.02 $Y2=1.51
cc_18 VNB C 0.00236701f $X=-0.19 $Y=-0.245 $X2=2.02 $Y2=1.7
cc_19 VNB C 0.00444264f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_C_c_219_n 0.0276181f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.51
cc_21 VNB N_D_c_308_n 0.0161919f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=1.345
cc_22 VNB N_D_M1006_g 0.00726469f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=2.465
cc_23 VNB N_D_c_310_n 0.0161882f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_D_M1008_g 0.00547738f $X=-0.19 $Y=-0.245 $X2=2 $Y2=1.675
cc_25 VNB D 0.00132852f $X=-0.19 $Y=-0.245 $X2=2 $Y2=2.465
cc_26 VNB N_D_c_313_n 0.042942f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_VPWR_c_427_n 0.203486f $X=-0.19 $Y=-0.245 $X2=2.02 $Y2=1.51
cc_28 VNB N_Y_c_496_n 0.0172492f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_Y_c_497_n 0.0354975f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.565
cc_30 VNB N_Y_c_498_n 0.00307439f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_Y_c_499_n 0.00292596f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_Y_c_500_n 0.00310024f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB Y 0.0277724f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_593_n 0.0398917f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=1.51
cc_35 VNB N_VGND_c_594_n 0.0149039f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=1.7
cc_36 VNB N_VGND_c_595_n 3.31577e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_596_n 0.0163828f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_597_n 0.00443255f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_598_n 0.0158731f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.51
cc_40 VNB N_VGND_c_599_n 3.23981e-19 $X=-0.19 $Y=-0.245 $X2=2.02 $Y2=1.51
cc_41 VNB N_VGND_c_600_n 0.0261048f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.565
cc_42 VNB N_VGND_c_601_n 0.0126445f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_602_n 0.00567425f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.565
cc_44 VNB N_VGND_c_603_n 0.0129398f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_604_n 0.0183725f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_605_n 0.274182f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_606_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_607_n 0.00634414f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_608_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_609_n 0.00513431f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VPB N_B_M1007_g 0.0238089f $X=-0.19 $Y=1.655 $X2=0.71 $Y2=2.465
cc_52 VPB N_B_M1015_g 0.0204069f $X=-0.19 $Y=1.655 $X2=2 $Y2=2.465
cc_53 VPB N_B_c_86_n 0.0132856f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.51
cc_54 VPB N_B_c_87_n 5.846e-19 $X=-0.19 $Y=1.655 $X2=0.71 $Y2=1.51
cc_55 VPB N_B_c_88_n 0.0066258f $X=-0.19 $Y=1.655 $X2=1.855 $Y2=1.7
cc_56 VPB N_B_c_97_n 0.00268974f $X=-0.19 $Y=1.655 $X2=2.02 $Y2=1.51
cc_57 VPB N_B_c_89_n 0.00632477f $X=-0.19 $Y=1.655 $X2=2.02 $Y2=1.51
cc_58 VPB B 0.0175453f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_59 VPB N_B_c_91_n 6.53693e-19 $X=-0.19 $Y=1.655 $X2=0.855 $Y2=1.565
cc_60 VPB N_A_M1000_g 0.0186876f $X=-0.19 $Y=1.655 $X2=0.71 $Y2=2.465
cc_61 VPB N_A_M1005_g 0.0186243f $X=-0.19 $Y=1.655 $X2=2 $Y2=1.675
cc_62 VPB N_C_M1001_g 0.0198823f $X=-0.19 $Y=1.655 $X2=0.71 $Y2=2.465
cc_63 VPB N_C_M1009_g 0.0225139f $X=-0.19 $Y=1.655 $X2=2 $Y2=2.465
cc_64 VPB N_C_c_222_n 0.00135562f $X=-0.19 $Y=1.655 $X2=0.855 $Y2=1.7
cc_65 VPB N_C_c_216_n 0.00776914f $X=-0.19 $Y=1.655 $X2=2.02 $Y2=1.51
cc_66 VPB C 4.91959e-19 $X=-0.19 $Y=1.655 $X2=2.02 $Y2=1.7
cc_67 VPB C 0.00169029f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_68 VPB N_C_c_219_n 0.00661822f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.51
cc_69 VPB N_C_c_227_n 0.0110482f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=1.565
cc_70 VPB N_D_M1006_g 0.0187149f $X=-0.19 $Y=1.655 $X2=0.71 $Y2=2.465
cc_71 VPB N_D_M1008_g 0.0182714f $X=-0.19 $Y=1.655 $X2=2 $Y2=1.675
cc_72 VPB N_A_74_367#_c_362_n 0.00743506f $X=-0.19 $Y=1.655 $X2=2 $Y2=0.655
cc_73 VPB N_A_74_367#_c_363_n 0.0365382f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_74 VPB N_A_74_367#_c_364_n 0.00745923f $X=-0.19 $Y=1.655 $X2=0.71 $Y2=1.51
cc_75 VPB N_A_74_367#_c_365_n 0.0202768f $X=-0.19 $Y=1.655 $X2=2.02 $Y2=1.51
cc_76 VPB N_VPWR_c_428_n 4.89148e-19 $X=-0.19 $Y=1.655 $X2=0.71 $Y2=2.465
cc_77 VPB N_VPWR_c_429_n 0.0341103f $X=-0.19 $Y=1.655 $X2=2 $Y2=0.655
cc_78 VPB N_VPWR_c_430_n 0.0814688f $X=-0.19 $Y=1.655 $X2=0.855 $Y2=1.7
cc_79 VPB N_VPWR_c_427_n 0.0692467f $X=-0.19 $Y=1.655 $X2=2.02 $Y2=1.51
cc_80 VPB N_VPWR_c_432_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_81 VPB N_Y_c_502_n 0.00493654f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.51
cc_82 VPB Y 0.0218529f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_83 VPB Y 0.021652f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_84 N_B_M1003_g N_A_c_164_n 0.0240083f $X=0.71 $Y=0.655 $X2=-0.19 $Y2=-0.245
cc_85 N_B_M1007_g N_A_M1000_g 0.0240083f $X=0.71 $Y=2.465 $X2=0 $Y2=0
cc_86 N_B_c_88_n N_A_M1000_g 0.0104608f $X=1.855 $Y=1.7 $X2=0 $Y2=0
cc_87 N_B_M1004_g N_A_c_166_n 0.0241009f $X=2 $Y=0.655 $X2=0 $Y2=0
cc_88 N_B_M1015_g N_A_M1005_g 0.0362988f $X=2 $Y=2.465 $X2=0 $Y2=0
cc_89 N_B_c_88_n N_A_M1005_g 0.011748f $X=1.855 $Y=1.7 $X2=0 $Y2=0
cc_90 N_B_M1003_g A 0.00307913f $X=0.71 $Y=0.655 $X2=0 $Y2=0
cc_91 N_B_M1004_g A 4.11007e-19 $X=2 $Y=0.655 $X2=0 $Y2=0
cc_92 N_B_c_87_n A 2.70096e-19 $X=0.71 $Y=1.51 $X2=0 $Y2=0
cc_93 N_B_c_88_n A 0.0293198f $X=1.855 $Y=1.7 $X2=0 $Y2=0
cc_94 N_B_c_97_n A 3.42831e-19 $X=2.02 $Y=1.51 $X2=0 $Y2=0
cc_95 N_B_c_89_n A 3.98597e-19 $X=2.02 $Y=1.51 $X2=0 $Y2=0
cc_96 N_B_c_91_n A 0.00796181f $X=0.855 $Y=1.565 $X2=0 $Y2=0
cc_97 N_B_c_87_n N_A_c_169_n 0.0240083f $X=0.71 $Y=1.51 $X2=0 $Y2=0
cc_98 N_B_c_88_n N_A_c_169_n 0.00244902f $X=1.855 $Y=1.7 $X2=0 $Y2=0
cc_99 N_B_c_97_n N_A_c_169_n 0.00131996f $X=2.02 $Y=1.51 $X2=0 $Y2=0
cc_100 N_B_c_89_n N_A_c_169_n 0.0224106f $X=2.02 $Y=1.51 $X2=0 $Y2=0
cc_101 N_B_c_91_n N_A_c_169_n 0.00516007f $X=0.855 $Y=1.565 $X2=0 $Y2=0
cc_102 N_B_M1004_g N_C_M1011_g 0.0246786f $X=2 $Y=0.655 $X2=0 $Y2=0
cc_103 N_B_M1015_g N_C_M1001_g 0.0239904f $X=2 $Y=2.465 $X2=0 $Y2=0
cc_104 N_B_c_97_n N_C_M1001_g 2.92862e-19 $X=2.02 $Y=1.51 $X2=0 $Y2=0
cc_105 N_B_M1015_g N_C_c_222_n 0.00210138f $X=2 $Y=2.465 $X2=0 $Y2=0
cc_106 N_B_c_97_n N_C_c_222_n 0.0237413f $X=2.02 $Y=1.51 $X2=0 $Y2=0
cc_107 N_B_c_89_n N_C_c_222_n 8.70727e-19 $X=2.02 $Y=1.51 $X2=0 $Y2=0
cc_108 N_B_c_97_n N_C_c_216_n 8.89548e-19 $X=2.02 $Y=1.51 $X2=0 $Y2=0
cc_109 N_B_c_89_n N_C_c_216_n 0.0213644f $X=2.02 $Y=1.51 $X2=0 $Y2=0
cc_110 N_B_c_86_n N_A_74_367#_c_362_n 0.00166261f $X=0.635 $Y=1.51 $X2=0 $Y2=0
cc_111 B N_A_74_367#_c_362_n 0.0240828f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_112 N_B_M1007_g N_A_74_367#_c_368_n 0.0129469f $X=0.71 $Y=2.465 $X2=0 $Y2=0
cc_113 N_B_M1015_g N_A_74_367#_c_368_n 0.015522f $X=2 $Y=2.465 $X2=0 $Y2=0
cc_114 N_B_c_97_n N_A_74_367#_c_368_n 0.0146306f $X=2.02 $Y=1.51 $X2=0 $Y2=0
cc_115 N_B_c_89_n N_A_74_367#_c_368_n 2.66669e-19 $X=2.02 $Y=1.51 $X2=0 $Y2=0
cc_116 B N_A_74_367#_c_368_n 0.0786319f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_117 N_B_c_97_n N_A_74_367#_c_373_n 0.00655924f $X=2.02 $Y=1.51 $X2=0 $Y2=0
cc_118 N_B_c_89_n N_A_74_367#_c_373_n 4.804e-19 $X=2.02 $Y=1.51 $X2=0 $Y2=0
cc_119 N_B_M1007_g N_VPWR_c_428_n 0.00121672f $X=0.71 $Y=2.465 $X2=0 $Y2=0
cc_120 N_B_M1015_g N_VPWR_c_428_n 0.00121672f $X=2 $Y=2.465 $X2=0 $Y2=0
cc_121 N_B_M1007_g N_VPWR_c_429_n 0.00585385f $X=0.71 $Y=2.465 $X2=0 $Y2=0
cc_122 N_B_M1015_g N_VPWR_c_430_n 0.00585385f $X=2 $Y=2.465 $X2=0 $Y2=0
cc_123 N_B_M1007_g N_VPWR_c_427_n 0.0118825f $X=0.71 $Y=2.465 $X2=0 $Y2=0
cc_124 N_B_M1015_g N_VPWR_c_427_n 0.0114676f $X=2 $Y=2.465 $X2=0 $Y2=0
cc_125 N_B_c_88_n N_Y_c_505_n 0.00407359f $X=1.855 $Y=1.7 $X2=0 $Y2=0
cc_126 N_B_c_88_n N_Y_c_506_n 0.00525113f $X=1.855 $Y=1.7 $X2=0 $Y2=0
cc_127 N_B_c_91_n N_Y_c_506_n 0.00212286f $X=0.855 $Y=1.565 $X2=0 $Y2=0
cc_128 N_B_M1004_g N_Y_c_508_n 0.00813322f $X=2 $Y=0.655 $X2=0 $Y2=0
cc_129 N_B_M1004_g N_Y_c_496_n 0.0125576f $X=2 $Y=0.655 $X2=0 $Y2=0
cc_130 N_B_c_97_n N_Y_c_496_n 0.0173226f $X=2.02 $Y=1.51 $X2=0 $Y2=0
cc_131 N_B_c_89_n N_Y_c_496_n 0.00272601f $X=2.02 $Y=1.51 $X2=0 $Y2=0
cc_132 N_B_M1004_g N_Y_c_498_n 0.00744736f $X=2 $Y=0.655 $X2=0 $Y2=0
cc_133 N_B_c_88_n N_Y_c_498_n 0.0113857f $X=1.855 $Y=1.7 $X2=0 $Y2=0
cc_134 N_B_c_97_n N_Y_c_498_n 0.00781954f $X=2.02 $Y=1.51 $X2=0 $Y2=0
cc_135 N_B_c_89_n N_Y_c_498_n 0.00181877f $X=2.02 $Y=1.51 $X2=0 $Y2=0
cc_136 N_B_M1004_g N_Y_c_499_n 7.92182e-19 $X=2 $Y=0.655 $X2=0 $Y2=0
cc_137 N_B_M1003_g N_VGND_c_593_n 0.00745762f $X=0.71 $Y=0.655 $X2=0 $Y2=0
cc_138 N_B_c_86_n N_VGND_c_593_n 0.00653393f $X=0.635 $Y=1.51 $X2=0 $Y2=0
cc_139 B N_VGND_c_593_n 0.0188963f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_140 N_B_M1003_g N_VGND_c_594_n 0.00585385f $X=0.71 $Y=0.655 $X2=0 $Y2=0
cc_141 N_B_M1003_g N_VGND_c_595_n 6.02213e-19 $X=0.71 $Y=0.655 $X2=0 $Y2=0
cc_142 N_B_M1004_g N_VGND_c_595_n 6.5421e-19 $X=2 $Y=0.655 $X2=0 $Y2=0
cc_143 N_B_M1004_g N_VGND_c_596_n 0.0054895f $X=2 $Y=0.655 $X2=0 $Y2=0
cc_144 N_B_M1004_g N_VGND_c_597_n 0.00845096f $X=2 $Y=0.655 $X2=0 $Y2=0
cc_145 N_B_M1003_g N_VGND_c_605_n 0.0116396f $X=0.71 $Y=0.655 $X2=0 $Y2=0
cc_146 N_B_M1004_g N_VGND_c_605_n 0.0104279f $X=2 $Y=0.655 $X2=0 $Y2=0
cc_147 N_A_M1000_g N_A_74_367#_c_368_n 0.010446f $X=1.14 $Y=2.465 $X2=0 $Y2=0
cc_148 N_A_M1005_g N_A_74_367#_c_368_n 0.010446f $X=1.57 $Y=2.465 $X2=0 $Y2=0
cc_149 N_A_M1000_g N_A_157_367#_c_412_n 0.0122129f $X=1.14 $Y=2.465 $X2=0 $Y2=0
cc_150 N_A_M1005_g N_A_157_367#_c_412_n 0.0122129f $X=1.57 $Y=2.465 $X2=0 $Y2=0
cc_151 N_A_M1000_g N_VPWR_c_428_n 0.0116523f $X=1.14 $Y=2.465 $X2=0 $Y2=0
cc_152 N_A_M1005_g N_VPWR_c_428_n 0.0116523f $X=1.57 $Y=2.465 $X2=0 $Y2=0
cc_153 N_A_M1000_g N_VPWR_c_429_n 0.00486043f $X=1.14 $Y=2.465 $X2=0 $Y2=0
cc_154 N_A_M1005_g N_VPWR_c_430_n 0.00486043f $X=1.57 $Y=2.465 $X2=0 $Y2=0
cc_155 N_A_M1000_g N_VPWR_c_427_n 0.0082726f $X=1.14 $Y=2.465 $X2=0 $Y2=0
cc_156 N_A_M1005_g N_VPWR_c_427_n 0.0082726f $X=1.57 $Y=2.465 $X2=0 $Y2=0
cc_157 N_A_c_164_n N_Y_c_505_n 0.0122595f $X=1.14 $Y=1.185 $X2=0 $Y2=0
cc_158 N_A_c_166_n N_Y_c_505_n 0.0125665f $X=1.57 $Y=1.185 $X2=0 $Y2=0
cc_159 A N_Y_c_505_n 0.0262719f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_160 N_A_c_169_n N_Y_c_505_n 0.00230884f $X=1.57 $Y=1.35 $X2=0 $Y2=0
cc_161 N_A_c_164_n N_Y_c_498_n 7.83637e-19 $X=1.14 $Y=1.185 $X2=0 $Y2=0
cc_162 N_A_c_166_n N_Y_c_498_n 0.00591119f $X=1.57 $Y=1.185 $X2=0 $Y2=0
cc_163 A N_Y_c_498_n 0.00338435f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_164 N_A_c_169_n N_Y_c_498_n 0.00329154f $X=1.57 $Y=1.35 $X2=0 $Y2=0
cc_165 N_A_c_164_n N_VGND_c_594_n 0.00486043f $X=1.14 $Y=1.185 $X2=0 $Y2=0
cc_166 N_A_c_164_n N_VGND_c_595_n 0.0108299f $X=1.14 $Y=1.185 $X2=0 $Y2=0
cc_167 N_A_c_166_n N_VGND_c_595_n 0.0107926f $X=1.57 $Y=1.185 $X2=0 $Y2=0
cc_168 N_A_c_166_n N_VGND_c_596_n 0.00486043f $X=1.57 $Y=1.185 $X2=0 $Y2=0
cc_169 N_A_c_164_n N_VGND_c_605_n 0.0082726f $X=1.14 $Y=1.185 $X2=0 $Y2=0
cc_170 N_A_c_166_n N_VGND_c_605_n 0.0082726f $X=1.57 $Y=1.185 $X2=0 $Y2=0
cc_171 N_C_M1011_g N_D_c_308_n 0.021496f $X=2.62 $Y=0.655 $X2=-0.19 $Y2=-0.245
cc_172 N_C_c_222_n N_D_M1006_g 0.00113391f $X=2.56 $Y=1.51 $X2=0 $Y2=0
cc_173 N_C_c_216_n N_D_M1006_g 0.0445624f $X=2.56 $Y=1.51 $X2=0 $Y2=0
cc_174 C N_D_M1006_g 0.00440708f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_175 N_C_c_227_n N_D_M1006_g 0.0123173f $X=3.465 $Y=1.645 $X2=0 $Y2=0
cc_176 N_C_M1012_g N_D_c_310_n 0.0152095f $X=3.91 $Y=0.655 $X2=0 $Y2=0
cc_177 N_C_M1009_g N_D_M1008_g 0.0544989f $X=3.98 $Y=2.465 $X2=0 $Y2=0
cc_178 C N_D_M1008_g 0.0132719f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_179 N_C_c_219_n N_D_M1008_g 0.0167908f $X=4 $Y=1.51 $X2=0 $Y2=0
cc_180 N_C_M1011_g D 6.1494e-19 $X=2.62 $Y=0.655 $X2=0 $Y2=0
cc_181 N_C_M1012_g D 8.49572e-19 $X=3.91 $Y=0.655 $X2=0 $Y2=0
cc_182 N_C_c_222_n D 0.00470873f $X=2.56 $Y=1.51 $X2=0 $Y2=0
cc_183 N_C_c_216_n D 8.78769e-19 $X=2.56 $Y=1.51 $X2=0 $Y2=0
cc_184 C D 0.00706416f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_185 N_C_c_227_n D 0.0213498f $X=3.465 $Y=1.645 $X2=0 $Y2=0
cc_186 N_C_M1012_g N_D_c_313_n 0.0167908f $X=3.91 $Y=0.655 $X2=0 $Y2=0
cc_187 N_C_c_222_n N_D_c_313_n 3.38093e-19 $X=2.56 $Y=1.51 $X2=0 $Y2=0
cc_188 N_C_c_216_n N_D_c_313_n 0.0116732f $X=2.56 $Y=1.51 $X2=0 $Y2=0
cc_189 C N_D_c_313_n 0.00654642f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_190 N_C_c_227_n N_D_c_313_n 0.00474533f $X=3.465 $Y=1.645 $X2=0 $Y2=0
cc_191 N_C_c_222_n N_A_74_367#_M1015_s 0.00310933f $X=2.56 $Y=1.51 $X2=0 $Y2=0
cc_192 C N_A_74_367#_M1009_d 0.00161645f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_193 N_C_M1001_g N_A_74_367#_c_373_n 0.00289696f $X=2.69 $Y=2.465 $X2=0 $Y2=0
cc_194 N_C_c_222_n N_A_74_367#_c_373_n 0.011704f $X=2.56 $Y=1.51 $X2=0 $Y2=0
cc_195 N_C_c_216_n N_A_74_367#_c_373_n 6.8197e-19 $X=2.56 $Y=1.51 $X2=0 $Y2=0
cc_196 N_C_M1001_g N_A_74_367#_c_382_n 0.0117681f $X=2.69 $Y=2.465 $X2=0 $Y2=0
cc_197 N_C_M1001_g N_A_74_367#_c_364_n 0.0144843f $X=2.69 $Y=2.465 $X2=0 $Y2=0
cc_198 N_C_M1009_g N_A_74_367#_c_364_n 0.0114269f $X=3.98 $Y=2.465 $X2=0 $Y2=0
cc_199 N_C_M1001_g N_VPWR_c_430_n 0.00357877f $X=2.69 $Y=2.465 $X2=0 $Y2=0
cc_200 N_C_M1009_g N_VPWR_c_430_n 0.00357877f $X=3.98 $Y=2.465 $X2=0 $Y2=0
cc_201 N_C_M1001_g N_VPWR_c_427_n 0.00601842f $X=2.69 $Y=2.465 $X2=0 $Y2=0
cc_202 N_C_M1009_g N_VPWR_c_427_n 0.00667818f $X=3.98 $Y=2.465 $X2=0 $Y2=0
cc_203 N_C_c_227_n N_A_553_367#_M1001_s 0.00176461f $X=3.465 $Y=1.645 $X2=-0.19
+ $Y2=-0.245
cc_204 C N_A_553_367#_M1008_s 0.00177752f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_205 N_C_M1001_g N_A_553_367#_c_476_n 0.0056797f $X=2.69 $Y=2.465 $X2=0 $Y2=0
cc_206 N_C_c_227_n N_A_553_367#_c_476_n 0.015328f $X=3.465 $Y=1.645 $X2=0 $Y2=0
cc_207 N_C_M1001_g N_A_553_367#_c_478_n 0.00296602f $X=2.69 $Y=2.465 $X2=0 $Y2=0
cc_208 N_C_M1009_g N_A_553_367#_c_479_n 0.00321923f $X=3.98 $Y=2.465 $X2=0 $Y2=0
cc_209 N_C_c_227_n N_A_553_367#_c_479_n 0.00286677f $X=3.465 $Y=1.645 $X2=0
+ $Y2=0
cc_210 N_C_c_227_n N_Y_M1006_d 0.00176891f $X=3.465 $Y=1.645 $X2=0 $Y2=0
cc_211 N_C_M1011_g N_Y_c_508_n 8.96285e-19 $X=2.62 $Y=0.655 $X2=0 $Y2=0
cc_212 N_C_M1011_g N_Y_c_496_n 0.010512f $X=2.62 $Y=0.655 $X2=0 $Y2=0
cc_213 N_C_c_222_n N_Y_c_496_n 0.0191849f $X=2.56 $Y=1.51 $X2=0 $Y2=0
cc_214 N_C_c_216_n N_Y_c_496_n 0.00371134f $X=2.56 $Y=1.51 $X2=0 $Y2=0
cc_215 N_C_M1011_g N_Y_c_530_n 0.00755622f $X=2.62 $Y=0.655 $X2=0 $Y2=0
cc_216 C N_Y_c_531_n 0.00389245f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_217 N_C_M1009_g N_Y_c_502_n 0.0163465f $X=3.98 $Y=2.465 $X2=0 $Y2=0
cc_218 C N_Y_c_502_n 0.0292122f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_219 N_C_c_219_n N_Y_c_502_n 6.32008e-19 $X=4 $Y=1.51 $X2=0 $Y2=0
cc_220 N_C_M1012_g N_Y_c_497_n 0.0152243f $X=3.91 $Y=0.655 $X2=0 $Y2=0
cc_221 C N_Y_c_497_n 0.0252407f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_222 N_C_c_219_n N_Y_c_497_n 0.00447774f $X=4 $Y=1.51 $X2=0 $Y2=0
cc_223 N_C_M1011_g N_Y_c_499_n 0.00761178f $X=2.62 $Y=0.655 $X2=0 $Y2=0
cc_224 N_C_c_222_n N_Y_c_499_n 0.00619374f $X=2.56 $Y=1.51 $X2=0 $Y2=0
cc_225 N_C_c_216_n N_Y_c_499_n 0.00230862f $X=2.56 $Y=1.51 $X2=0 $Y2=0
cc_226 N_C_c_227_n N_Y_c_499_n 0.00398931f $X=3.465 $Y=1.645 $X2=0 $Y2=0
cc_227 N_C_M1009_g N_Y_c_542_n 6.30161e-19 $X=3.98 $Y=2.465 $X2=0 $Y2=0
cc_228 N_C_c_227_n N_Y_c_542_n 0.0292122f $X=3.465 $Y=1.645 $X2=0 $Y2=0
cc_229 N_C_M1012_g N_Y_c_500_n 2.17608e-19 $X=3.91 $Y=0.655 $X2=0 $Y2=0
cc_230 C N_Y_c_500_n 0.0134317f $X=3.515 $Y=1.58 $X2=0 $Y2=0
cc_231 N_C_M1012_g Y 0.00481066f $X=3.91 $Y=0.655 $X2=0 $Y2=0
cc_232 N_C_M1009_g Y 0.00614721f $X=3.98 $Y=2.465 $X2=0 $Y2=0
cc_233 C Y 0.0385629f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_234 N_C_c_219_n Y 0.0045832f $X=4 $Y=1.51 $X2=0 $Y2=0
cc_235 N_C_M1011_g N_VGND_c_597_n 0.00828502f $X=2.62 $Y=0.655 $X2=0 $Y2=0
cc_236 N_C_M1011_g N_VGND_c_598_n 0.00518588f $X=2.62 $Y=0.655 $X2=0 $Y2=0
cc_237 N_C_M1011_g N_VGND_c_599_n 6.18296e-19 $X=2.62 $Y=0.655 $X2=0 $Y2=0
cc_238 N_C_M1012_g N_VGND_c_599_n 5.68743e-19 $X=3.91 $Y=0.655 $X2=0 $Y2=0
cc_239 N_C_M1012_g N_VGND_c_600_n 0.0112405f $X=3.91 $Y=0.655 $X2=0 $Y2=0
cc_240 N_C_M1012_g N_VGND_c_603_n 0.00486043f $X=3.91 $Y=0.655 $X2=0 $Y2=0
cc_241 N_C_M1011_g N_VGND_c_605_n 0.00965935f $X=2.62 $Y=0.655 $X2=0 $Y2=0
cc_242 N_C_M1012_g N_VGND_c_605_n 0.0082726f $X=3.91 $Y=0.655 $X2=0 $Y2=0
cc_243 N_D_M1006_g N_A_74_367#_c_364_n 0.00968453f $X=3.12 $Y=2.465 $X2=0 $Y2=0
cc_244 N_D_M1008_g N_A_74_367#_c_364_n 0.00968453f $X=3.55 $Y=2.465 $X2=0 $Y2=0
cc_245 N_D_M1006_g N_VPWR_c_430_n 0.00357877f $X=3.12 $Y=2.465 $X2=0 $Y2=0
cc_246 N_D_M1008_g N_VPWR_c_430_n 0.00357877f $X=3.55 $Y=2.465 $X2=0 $Y2=0
cc_247 N_D_M1006_g N_VPWR_c_427_n 0.00544922f $X=3.12 $Y=2.465 $X2=0 $Y2=0
cc_248 N_D_M1008_g N_VPWR_c_427_n 0.00544922f $X=3.55 $Y=2.465 $X2=0 $Y2=0
cc_249 N_D_M1006_g N_A_553_367#_c_479_n 0.0118527f $X=3.12 $Y=2.465 $X2=0 $Y2=0
cc_250 N_D_M1008_g N_A_553_367#_c_479_n 0.0106438f $X=3.55 $Y=2.465 $X2=0 $Y2=0
cc_251 N_D_c_308_n N_Y_c_531_n 0.010119f $X=3.05 $Y=1.185 $X2=0 $Y2=0
cc_252 N_D_c_310_n N_Y_c_531_n 0.0123392f $X=3.48 $Y=1.185 $X2=0 $Y2=0
cc_253 D N_Y_c_531_n 0.020082f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_254 N_D_c_313_n N_Y_c_531_n 0.00133921f $X=3.55 $Y=1.35 $X2=0 $Y2=0
cc_255 N_D_M1008_g N_Y_c_502_n 0.00792748f $X=3.55 $Y=2.465 $X2=0 $Y2=0
cc_256 N_D_c_308_n N_Y_c_499_n 0.00476752f $X=3.05 $Y=1.185 $X2=0 $Y2=0
cc_257 D N_Y_c_499_n 0.00587155f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_258 N_D_M1006_g N_Y_c_542_n 0.0036983f $X=3.12 $Y=2.465 $X2=0 $Y2=0
cc_259 N_D_M1008_g N_Y_c_542_n 0.00342325f $X=3.55 $Y=2.465 $X2=0 $Y2=0
cc_260 N_D_c_310_n N_Y_c_500_n 0.00250412f $X=3.48 $Y=1.185 $X2=0 $Y2=0
cc_261 N_D_c_313_n N_Y_c_500_n 0.00117584f $X=3.55 $Y=1.35 $X2=0 $Y2=0
cc_262 N_D_c_308_n N_VGND_c_598_n 0.00486043f $X=3.05 $Y=1.185 $X2=0 $Y2=0
cc_263 N_D_c_308_n N_VGND_c_599_n 0.0102179f $X=3.05 $Y=1.185 $X2=0 $Y2=0
cc_264 N_D_c_310_n N_VGND_c_599_n 0.0100168f $X=3.48 $Y=1.185 $X2=0 $Y2=0
cc_265 N_D_c_310_n N_VGND_c_600_n 6.14008e-19 $X=3.48 $Y=1.185 $X2=0 $Y2=0
cc_266 N_D_c_310_n N_VGND_c_603_n 0.00486043f $X=3.48 $Y=1.185 $X2=0 $Y2=0
cc_267 N_D_c_308_n N_VGND_c_605_n 0.0045769f $X=3.05 $Y=1.185 $X2=0 $Y2=0
cc_268 N_D_c_310_n N_VGND_c_605_n 0.0045769f $X=3.48 $Y=1.185 $X2=0 $Y2=0
cc_269 N_A_74_367#_c_368_n N_A_157_367#_M1007_d 0.00353353f $X=2.085 $Y=2.04
+ $X2=-0.19 $Y2=1.655
cc_270 N_A_74_367#_c_368_n N_A_157_367#_M1005_s 0.00349947f $X=2.085 $Y=2.04
+ $X2=0 $Y2=0
cc_271 N_A_74_367#_c_368_n N_A_157_367#_c_412_n 0.0323235f $X=2.085 $Y=2.04
+ $X2=0 $Y2=0
cc_272 N_A_74_367#_c_368_n N_A_157_367#_c_417_n 0.0135055f $X=2.085 $Y=2.04
+ $X2=0 $Y2=0
cc_273 N_A_74_367#_c_368_n N_A_157_367#_c_418_n 0.0135055f $X=2.085 $Y=2.04
+ $X2=0 $Y2=0
cc_274 N_A_74_367#_c_368_n N_VPWR_M1000_d 0.00340044f $X=2.085 $Y=2.04 $X2=-0.19
+ $Y2=1.655
cc_275 N_A_74_367#_c_363_n N_VPWR_c_429_n 0.0190529f $X=0.495 $Y=2.91 $X2=0
+ $Y2=0
cc_276 N_A_74_367#_c_382_n N_VPWR_c_430_n 0.029652f $X=2.307 $Y=2.905 $X2=0
+ $Y2=0
cc_277 N_A_74_367#_c_364_n N_VPWR_c_430_n 0.103807f $X=4.1 $Y=2.99 $X2=0 $Y2=0
cc_278 N_A_74_367#_M1007_s N_VPWR_c_427_n 0.00249946f $X=0.37 $Y=1.835 $X2=0
+ $Y2=0
cc_279 N_A_74_367#_M1015_s N_VPWR_c_427_n 0.00475096f $X=2.075 $Y=1.835 $X2=0
+ $Y2=0
cc_280 N_A_74_367#_M1009_d N_VPWR_c_427_n 0.00215161f $X=4.055 $Y=1.835 $X2=0
+ $Y2=0
cc_281 N_A_74_367#_c_363_n N_VPWR_c_427_n 0.0113912f $X=0.495 $Y=2.91 $X2=0
+ $Y2=0
cc_282 N_A_74_367#_c_382_n N_VPWR_c_427_n 0.0173006f $X=2.307 $Y=2.905 $X2=0
+ $Y2=0
cc_283 N_A_74_367#_c_364_n N_VPWR_c_427_n 0.0663354f $X=4.1 $Y=2.99 $X2=0 $Y2=0
cc_284 N_A_74_367#_c_364_n N_A_553_367#_M1001_s 0.00332344f $X=4.1 $Y=2.99
+ $X2=-0.19 $Y2=1.655
cc_285 N_A_74_367#_c_364_n N_A_553_367#_M1008_s 0.00332774f $X=4.1 $Y=2.99 $X2=0
+ $Y2=0
cc_286 N_A_74_367#_c_373_n N_A_553_367#_c_476_n 0.00621108f $X=2.307 $Y=2.125
+ $X2=0 $Y2=0
cc_287 N_A_74_367#_c_382_n N_A_553_367#_c_476_n 0.0251686f $X=2.307 $Y=2.905
+ $X2=0 $Y2=0
cc_288 N_A_74_367#_c_382_n N_A_553_367#_c_478_n 0.0164505f $X=2.307 $Y=2.905
+ $X2=0 $Y2=0
cc_289 N_A_74_367#_c_364_n N_A_553_367#_c_478_n 0.014411f $X=4.1 $Y=2.99 $X2=0
+ $Y2=0
cc_290 N_A_74_367#_c_364_n N_A_553_367#_c_479_n 0.044282f $X=4.1 $Y=2.99 $X2=0
+ $Y2=0
cc_291 N_A_74_367#_c_364_n N_Y_M1006_d 0.00332774f $X=4.1 $Y=2.99 $X2=0 $Y2=0
cc_292 N_A_74_367#_M1009_d N_Y_c_502_n 0.00760562f $X=4.055 $Y=1.835 $X2=0 $Y2=0
cc_293 N_A_74_367#_c_365_n N_Y_c_502_n 0.0202647f $X=4.195 $Y=2.54 $X2=0 $Y2=0
cc_294 N_A_157_367#_c_412_n N_VPWR_M1000_d 0.00353353f $X=1.69 $Y=2.38 $X2=1.14
+ $Y2=1.185
cc_295 N_A_157_367#_c_412_n N_VPWR_c_428_n 0.0170777f $X=1.69 $Y=2.38 $X2=1.14
+ $Y2=2.465
cc_296 N_A_157_367#_c_417_n N_VPWR_c_429_n 0.0136943f $X=0.925 $Y=2.46 $X2=1.57
+ $Y2=0.655
cc_297 N_A_157_367#_c_418_n N_VPWR_c_430_n 0.0136943f $X=1.785 $Y=2.46 $X2=1.285
+ $Y2=1.35
cc_298 N_A_157_367#_M1007_d N_VPWR_c_427_n 0.0041489f $X=0.785 $Y=1.835
+ $X2=1.285 $Y2=1.35
cc_299 N_A_157_367#_M1005_s N_VPWR_c_427_n 0.0041489f $X=1.645 $Y=1.835
+ $X2=1.285 $Y2=1.35
cc_300 N_A_157_367#_c_417_n N_VPWR_c_427_n 0.00866972f $X=0.925 $Y=2.46
+ $X2=1.285 $Y2=1.35
cc_301 N_A_157_367#_c_418_n N_VPWR_c_427_n 0.00866972f $X=1.785 $Y=2.46
+ $X2=1.285 $Y2=1.35
cc_302 N_VPWR_c_427_n N_A_553_367#_M1001_s 0.00225186f $X=4.56 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_303 N_VPWR_c_427_n N_A_553_367#_M1008_s 0.00225186f $X=4.56 $Y=3.33 $X2=0
+ $Y2=0
cc_304 N_VPWR_c_427_n N_Y_M1006_d 0.00225186f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_305 N_A_553_367#_c_479_n N_Y_M1006_d 0.00348729f $X=3.765 $Y=2.61 $X2=0.71
+ $Y2=1.675
cc_306 N_A_553_367#_M1008_s N_Y_c_502_n 0.00404431f $X=3.625 $Y=1.835 $X2=0.385
+ $Y2=1.51
cc_307 N_A_553_367#_c_479_n N_Y_c_502_n 0.0146677f $X=3.765 $Y=2.61 $X2=0.385
+ $Y2=1.51
cc_308 N_A_553_367#_c_479_n N_Y_c_542_n 0.0164214f $X=3.765 $Y=2.61 $X2=0 $Y2=0
cc_309 N_Y_c_505_n N_VGND_M1010_d 0.00329816f $X=1.62 $Y=0.955 $X2=0 $Y2=0
cc_310 N_Y_c_531_n N_VGND_M1002_s 0.00425454f $X=3.59 $Y=0.93 $X2=0 $Y2=0
cc_311 N_Y_c_497_n N_VGND_M1012_d 0.00253571f $X=4.4 $Y=1.09 $X2=0 $Y2=0
cc_312 N_Y_c_572_p N_VGND_c_594_n 0.0125413f $X=0.925 $Y=0.43 $X2=0 $Y2=0
cc_313 N_Y_c_505_n N_VGND_c_595_n 0.0170777f $X=1.62 $Y=0.955 $X2=0 $Y2=0
cc_314 N_Y_c_508_n N_VGND_c_596_n 0.015688f $X=1.785 $Y=0.42 $X2=0 $Y2=0
cc_315 N_Y_c_508_n N_VGND_c_597_n 0.0444483f $X=1.785 $Y=0.42 $X2=0 $Y2=0
cc_316 N_Y_c_496_n N_VGND_c_597_n 0.0271222f $X=2.65 $Y=1.17 $X2=0 $Y2=0
cc_317 N_Y_c_530_n N_VGND_c_597_n 0.0452116f $X=2.835 $Y=0.42 $X2=0 $Y2=0
cc_318 N_Y_c_499_n N_VGND_c_597_n 0.00576821f $X=2.79 $Y=0.93 $X2=0 $Y2=0
cc_319 N_Y_c_530_n N_VGND_c_598_n 0.0170515f $X=2.835 $Y=0.42 $X2=0 $Y2=0
cc_320 N_Y_c_531_n N_VGND_c_599_n 0.016709f $X=3.59 $Y=0.93 $X2=0 $Y2=0
cc_321 N_Y_c_497_n N_VGND_c_600_n 0.0220026f $X=4.4 $Y=1.09 $X2=0 $Y2=0
cc_322 N_Y_c_582_p N_VGND_c_603_n 0.0124525f $X=3.695 $Y=0.42 $X2=0 $Y2=0
cc_323 N_Y_M1003_s N_VGND_c_605_n 0.00449877f $X=0.785 $Y=0.235 $X2=0 $Y2=0
cc_324 N_Y_M1014_s N_VGND_c_605_n 0.00380103f $X=1.645 $Y=0.235 $X2=0 $Y2=0
cc_325 N_Y_M1011_s N_VGND_c_605_n 0.00252268f $X=2.695 $Y=0.235 $X2=0 $Y2=0
cc_326 N_Y_M1013_d N_VGND_c_605_n 0.00407324f $X=3.555 $Y=0.235 $X2=0 $Y2=0
cc_327 N_Y_c_572_p N_VGND_c_605_n 0.00823619f $X=0.925 $Y=0.43 $X2=0 $Y2=0
cc_328 N_Y_c_508_n N_VGND_c_605_n 0.00984745f $X=1.785 $Y=0.42 $X2=0 $Y2=0
cc_329 N_Y_c_530_n N_VGND_c_605_n 0.0105335f $X=2.835 $Y=0.42 $X2=0 $Y2=0
cc_330 N_Y_c_531_n N_VGND_c_605_n 0.0105096f $X=3.59 $Y=0.93 $X2=0 $Y2=0
cc_331 N_Y_c_582_p N_VGND_c_605_n 0.00730901f $X=3.695 $Y=0.42 $X2=0 $Y2=0
cc_332 N_Y_c_500_n N_VGND_c_605_n 3.11813e-19 $X=3.695 $Y=0.93 $X2=0 $Y2=0
