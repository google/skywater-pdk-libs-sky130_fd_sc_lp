* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__and4_lp2 A B C D VGND VNB VPB VPWR X
X0 a_114_47# a_84_21# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 X a_84_21# a_114_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 VGND D a_294_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 VPWR D a_84_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X4 a_372_47# B a_450_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 X a_84_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X6 a_84_21# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X7 a_450_47# A a_84_21# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 VPWR B a_84_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X9 a_294_47# C a_372_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 a_84_21# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
.ends
