* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__sdfxbp_lp CLK D SCD SCE VGND VNB VPB VPWR Q Q_N
X0 a_1859_155# a_2089_254# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 a_2751_127# a_2089_254# a_2714_401# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 a_1278_155# a_706_66# a_1482_347# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X3 a_2040_352# a_2089_254# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X4 a_1127_155# a_975_347# a_1278_155# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 VGND a_1902_347# a_2331_57# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 VPWR a_2714_401# Q_N VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X7 a_2331_57# a_1902_347# a_2089_254# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 a_1482_347# a_1530_231# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X9 a_706_66# CLK a_789_66# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 a_27_409# SCE VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X11 a_343_417# a_975_347# a_1278_155# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X12 a_27_409# SCE a_141_125# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X13 a_1674_125# a_1278_155# a_1530_231# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X14 a_1902_347# a_975_347# a_2040_352# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X15 a_2593_127# a_2089_254# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X16 VGND a_2714_401# a_3015_57# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X17 VGND a_1278_155# a_1674_125# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X18 VPWR SCD a_239_417# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X19 a_141_125# SCE VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X20 a_239_417# a_27_409# a_343_417# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X21 VPWR a_1278_155# a_1530_231# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X22 a_1530_231# a_706_66# a_1902_347# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X23 a_3015_57# a_2714_401# Q_N VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X24 VPWR a_706_66# a_975_347# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X25 a_789_66# CLK VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X26 Q a_2089_254# a_2593_127# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X27 a_337_125# D a_343_417# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X28 a_1859_155# a_706_66# a_1902_347# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X29 VPWR a_1902_347# a_2089_254# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X30 VPWR a_2089_254# a_2714_401# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X31 VGND a_2089_254# a_2751_127# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X32 a_523_125# SCD VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X33 a_706_66# CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X34 a_1902_347# a_975_347# a_1530_231# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X35 Q a_2089_254# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X36 VGND a_27_409# a_337_125# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X37 VGND a_706_66# a_947_66# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X38 a_343_417# SCE a_523_125# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X39 a_1127_155# a_1530_231# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X40 a_449_417# SCE VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X41 a_1278_155# a_706_66# a_343_417# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X42 a_947_66# a_706_66# a_975_347# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X43 a_343_417# D a_449_417# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
.ends
