* File: sky130_fd_sc_lp__xor2_2.spice
* Created: Wed Sep  2 10:41:15 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__xor2_2.pex.spice"
.subckt sky130_fd_sc_lp__xor2_2  VNB VPB A B VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1003 N_VGND_M1003_d N_A_M1003_g N_A_149_65#_M1003_s VNB NSHORT L=0.15 W=0.84
+ AD=0.3349 AS=0.1176 PD=2.66 PS=1.12 NRD=14.28 NRS=0 M=1 R=5.6 SA=75000.3
+ SB=75005.3 A=0.126 P=1.98 MULT=1
MM1009 N_VGND_M1009_d N_B_M1009_g N_A_149_65#_M1003_s VNB NSHORT L=0.15 W=0.84
+ AD=0.20075 AS=0.1176 PD=1.39 PS=1.12 NRD=12.132 NRS=0 M=1 R=5.6 SA=75000.7
+ SB=75004.8 A=0.126 P=1.98 MULT=1
MM1011 N_VGND_M1009_d N_B_M1011_g N_A_149_65#_M1011_s VNB NSHORT L=0.15 W=0.84
+ AD=0.20075 AS=0.2142 PD=1.39 PS=1.35 NRD=12.132 NRS=16.428 M=1 R=5.6
+ SA=75001.3 SB=75004.2 A=0.126 P=1.98 MULT=1
MM1004 N_VGND_M1004_d N_A_M1004_g N_A_149_65#_M1011_s VNB NSHORT L=0.15 W=0.84
+ AD=0.21545 AS=0.2142 PD=1.425 PS=1.35 NRD=12.132 NRS=16.428 M=1 R=5.6 SA=75002
+ SB=75003.6 A=0.126 P=1.98 MULT=1
MM1007 N_VGND_M1004_d N_A_149_65#_M1007_g N_X_M1007_s VNB NSHORT L=0.15 W=0.84
+ AD=0.21545 AS=0.1176 PD=1.425 PS=1.12 NRD=17.136 NRS=0 M=1 R=5.6 SA=75002.6
+ SB=75003 A=0.126 P=1.98 MULT=1
MM1019 N_VGND_M1019_d N_A_149_65#_M1019_g N_X_M1007_s VNB NSHORT L=0.15 W=0.84
+ AD=0.20075 AS=0.1176 PD=1.39 PS=1.12 NRD=12.132 NRS=0 M=1 R=5.6 SA=75003
+ SB=75002.5 A=0.126 P=1.98 MULT=1
MM1008 N_A_814_65#_M1008_d N_A_M1008_g N_VGND_M1019_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.20075 PD=1.12 PS=1.39 NRD=0 NRS=12.132 M=1 R=5.6 SA=75003.6
+ SB=75001.9 A=0.126 P=1.98 MULT=1
MM1012 N_A_814_65#_M1008_d N_B_M1012_g N_X_M1012_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1281 PD=1.12 PS=1.145 NRD=0 NRS=0 M=1 R=5.6 SA=75004 SB=75001.5
+ A=0.126 P=1.98 MULT=1
MM1018 N_A_814_65#_M1018_d N_B_M1018_g N_X_M1012_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2709 AS=0.1281 PD=1.485 PS=1.145 NRD=26.064 NRS=3.564 M=1 R=5.6
+ SA=75004.5 SB=75001.1 A=0.126 P=1.98 MULT=1
MM1010 N_A_814_65#_M1018_d N_A_M1010_g N_VGND_M1010_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2709 AS=0.2814 PD=1.485 PS=2.35 NRD=0 NRS=9.996 M=1 R=5.6 SA=75005.3
+ SB=75000.3 A=0.126 P=1.98 MULT=1
MM1001 N_A_149_367#_M1001_d N_A_M1001_g N_VPWR_M1001_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.378 PD=1.54 PS=3.12 NRD=0 NRS=1.8124 M=1 R=8.4 SA=75000.2
+ SB=75001.6 A=0.189 P=2.82 MULT=1
MM1000 N_A_149_367#_M1001_d N_B_M1000_g N_A_149_65#_M1000_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.7
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1014 N_A_149_367#_M1014_d N_B_M1014_g N_A_149_65#_M1000_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.2331 AS=0.1764 PD=1.63 PS=1.54 NRD=3.1126 NRS=0 M=1 R=8.4
+ SA=75001.1 SB=75000.7 A=0.189 P=2.82 MULT=1
MM1015 N_A_149_367#_M1014_d N_A_M1015_g N_VPWR_M1015_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.2331 AS=0.3339 PD=1.63 PS=3.05 NRD=10.9335 NRS=0 M=1 R=8.4 SA=75001.6
+ SB=75000.2 A=0.189 P=2.82 MULT=1
MM1002 N_X_M1002_d N_A_149_65#_M1002_g N_A_532_367#_M1002_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75002.7 A=0.189 P=2.82 MULT=1
MM1016 N_X_M1002_d N_A_149_65#_M1016_g N_A_532_367#_M1016_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75002.2 A=0.189 P=2.82 MULT=1
MM1006 N_VPWR_M1006_d N_A_M1006_g N_A_532_367#_M1016_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.290975 AS=0.1764 PD=1.795 PS=1.54 NRD=13.2778 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75001.8 A=0.189 P=2.82 MULT=1
MM1005 N_VPWR_M1006_d N_B_M1005_g N_A_532_367#_M1005_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.290975 AS=0.1764 PD=1.795 PS=1.54 NRD=13.2778 NRS=0 M=1 R=8.4 SA=75001.6
+ SB=75001.2 A=0.189 P=2.82 MULT=1
MM1017 N_VPWR_M1017_d N_B_M1017_g N_A_532_367#_M1005_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.290975 AS=0.1764 PD=1.795 PS=1.54 NRD=13.2778 NRS=0 M=1 R=8.4 SA=75002.1
+ SB=75000.8 A=0.189 P=2.82 MULT=1
MM1013 N_VPWR_M1017_d N_A_M1013_g N_A_532_367#_M1013_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.290975 AS=0.3339 PD=1.795 PS=3.05 NRD=13.2778 NRS=0 M=1 R=8.4 SA=75002.7
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX20_noxref VNB VPB NWDIODE A=12.3463 P=16.97
*
.include "sky130_fd_sc_lp__xor2_2.pxi.spice"
*
.ends
*
*
