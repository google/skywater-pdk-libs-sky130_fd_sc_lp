* File: sky130_fd_sc_lp__o311ai_2.pex.spice
* Created: Wed Sep  2 10:23:52 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O311AI_2%A1 1 3 6 8 10 13 15 16 24
r41 22 24 28.8521 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.78 $Y=1.35
+ $X2=0.945 $Y2=1.35
r42 19 22 46.3382 $w=3.3e-07 $l=2.65e-07 $layer=POLY_cond $X=0.515 $Y=1.35
+ $X2=0.78 $Y2=1.35
r43 16 22 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.78
+ $Y=1.35 $X2=0.78 $Y2=1.35
r44 15 16 22.1269 $w=2.48e-07 $l=4.8e-07 $layer=LI1_cond $X=0.24 $Y=1.31
+ $X2=0.72 $Y2=1.31
r45 11 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.945 $Y=1.515
+ $X2=0.945 $Y2=1.35
r46 11 13 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=0.945 $Y=1.515
+ $X2=0.945 $Y2=2.465
r47 8 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.945 $Y=1.185
+ $X2=0.945 $Y2=1.35
r48 8 10 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.945 $Y=1.185
+ $X2=0.945 $Y2=0.655
r49 4 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.515 $Y=1.515
+ $X2=0.515 $Y2=1.35
r50 4 6 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=0.515 $Y=1.515
+ $X2=0.515 $Y2=2.465
r51 1 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.515 $Y=1.185
+ $X2=0.515 $Y2=1.35
r52 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.515 $Y=1.185
+ $X2=0.515 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__O311AI_2%A2 1 3 6 8 10 13 15 16 24
c52 13 0 4.40372e-20 $X=1.805 $Y=2.465
r53 22 24 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=1.735 $Y=1.35
+ $X2=1.805 $Y2=1.35
r54 19 22 62.9501 $w=3.3e-07 $l=3.6e-07 $layer=POLY_cond $X=1.375 $Y=1.35
+ $X2=1.735 $Y2=1.35
r55 16 22 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.735
+ $Y=1.35 $X2=1.735 $Y2=1.35
r56 15 16 22.1269 $w=2.48e-07 $l=4.8e-07 $layer=LI1_cond $X=1.2 $Y=1.31 $X2=1.68
+ $Y2=1.31
r57 11 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.805 $Y=1.515
+ $X2=1.805 $Y2=1.35
r58 11 13 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=1.805 $Y=1.515
+ $X2=1.805 $Y2=2.465
r59 8 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.805 $Y=1.185
+ $X2=1.805 $Y2=1.35
r60 8 10 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.805 $Y=1.185
+ $X2=1.805 $Y2=0.655
r61 4 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.375 $Y=1.515
+ $X2=1.375 $Y2=1.35
r62 4 6 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=1.375 $Y=1.515
+ $X2=1.375 $Y2=2.465
r63 1 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.375 $Y=1.185
+ $X2=1.375 $Y2=1.35
r64 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.375 $Y=1.185
+ $X2=1.375 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__O311AI_2%A3 3 5 7 10 12 14 15 16 17 27 29 39
c53 29 0 4.40372e-20 $X=2.68 $Y=1.355
c54 27 0 1.98392e-19 $X=3.045 $Y=1.5
c55 10 0 1.49555e-19 $X=3.045 $Y=0.655
r56 29 39 1.63459 $w=3.4e-07 $l=4e-08 $layer=LI1_cond $X=2.68 $Y=1.355 $X2=2.64
+ $Y2=1.355
r57 25 27 12.1854 $w=3.56e-07 $l=9e-08 $layer=POLY_cond $X=2.955 $Y=1.5
+ $X2=3.045 $Y2=1.5
r58 25 26 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.955
+ $Y=1.44 $X2=2.955 $Y2=1.44
r59 23 25 27.0787 $w=3.56e-07 $l=2e-07 $layer=POLY_cond $X=2.755 $Y=1.5
+ $X2=2.955 $Y2=1.5
r60 22 23 64.9888 $w=3.56e-07 $l=4.8e-07 $layer=POLY_cond $X=2.275 $Y=1.5
+ $X2=2.755 $Y2=1.5
r61 17 26 5.59274 $w=3.38e-07 $l=1.65e-07 $layer=LI1_cond $X=3.12 $Y=1.355
+ $X2=2.955 $Y2=1.355
r62 16 39 0.935333 $w=3e-07 $l=2.3e-08 $layer=LI1_cond $X=2.617 $Y=1.355
+ $X2=2.64 $Y2=1.355
r63 16 26 8.57553 $w=3.38e-07 $l=2.53e-07 $layer=LI1_cond $X=2.702 $Y=1.355
+ $X2=2.955 $Y2=1.355
r64 16 29 0.745698 $w=3.38e-07 $l=2.2e-08 $layer=LI1_cond $X=2.702 $Y=1.355
+ $X2=2.68 $Y2=1.355
r65 15 16 18.5847 $w=3e-07 $l=4.57e-07 $layer=LI1_cond $X=2.16 $Y=1.355
+ $X2=2.617 $Y2=1.355
r66 12 27 18.9551 $w=3.56e-07 $l=2.86575e-07 $layer=POLY_cond $X=3.185 $Y=1.725
+ $X2=3.045 $Y2=1.5
r67 12 14 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=3.185 $Y=1.725
+ $X2=3.185 $Y2=2.465
r68 8 27 23.0368 $w=1.5e-07 $l=2.25e-07 $layer=POLY_cond $X=3.045 $Y=1.275
+ $X2=3.045 $Y2=1.5
r69 8 10 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=3.045 $Y=1.275
+ $X2=3.045 $Y2=0.655
r70 5 23 23.0368 $w=1.5e-07 $l=2.25e-07 $layer=POLY_cond $X=2.755 $Y=1.725
+ $X2=2.755 $Y2=1.5
r71 5 7 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=2.755 $Y=1.725
+ $X2=2.755 $Y2=2.465
r72 1 22 23.0368 $w=1.5e-07 $l=2.25e-07 $layer=POLY_cond $X=2.275 $Y=1.275
+ $X2=2.275 $Y2=1.5
r73 1 3 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=2.275 $Y=1.275
+ $X2=2.275 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__O311AI_2%B1 1 3 4 6 7 9 10 12 13 14 21
c49 14 0 3.47947e-19 $X=4.08 $Y=1.295
c50 1 0 6.04418e-20 $X=3.475 $Y=1.185
r51 21 23 44.1752 $w=4.91e-07 $l=4.5e-07 $layer=POLY_cond $X=3.975 $Y=1.455
+ $X2=4.425 $Y2=1.455
r52 21 22 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.975
+ $Y=1.35 $X2=3.975 $Y2=1.35
r53 19 21 6.87169 $w=4.91e-07 $l=7e-08 $layer=POLY_cond $X=3.905 $Y=1.455
+ $X2=3.975 $Y2=1.455
r54 18 19 28.4684 $w=4.91e-07 $l=2.9e-07 $layer=POLY_cond $X=3.615 $Y=1.455
+ $X2=3.905 $Y2=1.455
r55 17 18 13.7434 $w=4.91e-07 $l=1.4e-07 $layer=POLY_cond $X=3.475 $Y=1.455
+ $X2=3.615 $Y2=1.455
r56 14 22 3.66686 $w=3.28e-07 $l=1.05e-07 $layer=LI1_cond $X=4.08 $Y=1.35
+ $X2=3.975 $Y2=1.35
r57 13 22 13.0959 $w=3.28e-07 $l=3.75e-07 $layer=LI1_cond $X=3.6 $Y=1.35
+ $X2=3.975 $Y2=1.35
r58 10 23 30.9498 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=4.425 $Y=1.725
+ $X2=4.425 $Y2=1.455
r59 10 12 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=4.425 $Y=1.725
+ $X2=4.425 $Y2=2.465
r60 7 19 30.9498 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=3.905 $Y=1.185
+ $X2=3.905 $Y2=1.455
r61 7 9 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=3.905 $Y=1.185
+ $X2=3.905 $Y2=0.655
r62 4 18 30.9498 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=3.615 $Y=1.725
+ $X2=3.615 $Y2=1.455
r63 4 6 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=3.615 $Y=1.725
+ $X2=3.615 $Y2=2.465
r64 1 17 30.9498 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=3.475 $Y=1.185
+ $X2=3.475 $Y2=1.455
r65 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=3.475 $Y=1.185
+ $X2=3.475 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__O311AI_2%C1 1 3 6 8 10 13 15 21
r44 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.47
+ $Y=1.46 $X2=5.47 $Y2=1.46
r45 19 21 32.3493 $w=3.3e-07 $l=1.85e-07 $layer=POLY_cond $X=5.285 $Y=1.46
+ $X2=5.47 $Y2=1.46
r46 17 19 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=4.855 $Y=1.46
+ $X2=5.285 $Y2=1.46
r47 15 22 5.00403 $w=3.78e-07 $l=1.65e-07 $layer=LI1_cond $X=5.485 $Y=1.295
+ $X2=5.485 $Y2=1.46
r48 11 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.285 $Y=1.625
+ $X2=5.285 $Y2=1.46
r49 11 13 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=5.285 $Y=1.625
+ $X2=5.285 $Y2=2.465
r50 8 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.285 $Y=1.295
+ $X2=5.285 $Y2=1.46
r51 8 10 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=5.285 $Y=1.295
+ $X2=5.285 $Y2=0.765
r52 4 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.855 $Y=1.625
+ $X2=4.855 $Y2=1.46
r53 4 6 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=4.855 $Y=1.625
+ $X2=4.855 $Y2=2.465
r54 1 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.855 $Y=1.295
+ $X2=4.855 $Y2=1.46
r55 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=4.855 $Y=1.295
+ $X2=4.855 $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_LP__O311AI_2%A_35_367# 1 2 3 12 16 17 20 24 28 30
r47 26 28 9.08657 $w=2.58e-07 $l=2.05e-07 $layer=LI1_cond $X=2.055 $Y=1.775
+ $X2=2.055 $Y2=1.98
r48 25 30 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.255 $Y=1.69
+ $X2=1.16 $Y2=1.69
r49 24 26 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=1.925 $Y=1.69
+ $X2=2.055 $Y2=1.775
r50 24 25 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.925 $Y=1.69
+ $X2=1.255 $Y2=1.69
r51 20 22 54.2871 $w=1.88e-07 $l=9.3e-07 $layer=LI1_cond $X=1.16 $Y=1.98
+ $X2=1.16 $Y2=2.91
r52 18 30 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.16 $Y=1.775
+ $X2=1.16 $Y2=1.69
r53 18 20 11.9665 $w=1.88e-07 $l=2.05e-07 $layer=LI1_cond $X=1.16 $Y=1.775
+ $X2=1.16 $Y2=1.98
r54 16 30 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.065 $Y=1.69
+ $X2=1.16 $Y2=1.69
r55 16 17 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.065 $Y=1.69
+ $X2=0.395 $Y2=1.69
r56 12 14 41.222 $w=2.58e-07 $l=9.3e-07 $layer=LI1_cond $X=0.265 $Y=1.98
+ $X2=0.265 $Y2=2.91
r57 10 17 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=0.265 $Y=1.775
+ $X2=0.395 $Y2=1.69
r58 10 12 9.08657 $w=2.58e-07 $l=2.05e-07 $layer=LI1_cond $X=0.265 $Y=1.775
+ $X2=0.265 $Y2=1.98
r59 3 28 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=1.88
+ $Y=1.835 $X2=2.02 $Y2=1.98
r60 2 22 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=1.02
+ $Y=1.835 $X2=1.16 $Y2=2.91
r61 2 20 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.02
+ $Y=1.835 $X2=1.16 $Y2=1.98
r62 1 14 400 $w=1.7e-07 $l=1.13578e-06 $layer=licon1_PDIFF $count=1 $X=0.175
+ $Y=1.835 $X2=0.3 $Y2=2.91
r63 1 12 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.175
+ $Y=1.835 $X2=0.3 $Y2=1.98
.ends

.subckt PM_SKY130_FD_SC_LP__O311AI_2%VPWR 1 2 3 12 18 24 28 30 35 43 50 51 54 57
+ 60
r74 60 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r75 57 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r76 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r77 51 61 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=5.04 $Y2=3.33
r78 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r79 48 60 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.235 $Y=3.33
+ $X2=5.07 $Y2=3.33
r80 48 50 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=5.235 $Y=3.33
+ $X2=5.52 $Y2=3.33
r81 47 61 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.04 $Y2=3.33
r82 47 58 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=4.08 $Y2=3.33
r83 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r84 44 57 13.764 $w=1.7e-07 $l=3.55e-07 $layer=LI1_cond $X=4.375 $Y=3.33
+ $X2=4.02 $Y2=3.33
r85 44 46 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=4.375 $Y=3.33
+ $X2=4.56 $Y2=3.33
r86 43 60 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.905 $Y=3.33
+ $X2=5.07 $Y2=3.33
r87 43 46 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=4.905 $Y=3.33
+ $X2=4.56 $Y2=3.33
r88 42 58 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r89 41 42 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r90 39 55 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r91 38 41 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=1.2 $Y=3.33 $X2=3.6
+ $Y2=3.33
r92 38 39 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r93 36 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.895 $Y=3.33
+ $X2=0.73 $Y2=3.33
r94 36 38 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.895 $Y=3.33
+ $X2=1.2 $Y2=3.33
r95 35 57 13.764 $w=1.7e-07 $l=3.55e-07 $layer=LI1_cond $X=3.665 $Y=3.33
+ $X2=4.02 $Y2=3.33
r96 35 41 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=3.665 $Y=3.33
+ $X2=3.6 $Y2=3.33
r97 33 55 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r98 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r99 30 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.565 $Y=3.33
+ $X2=0.73 $Y2=3.33
r100 30 32 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.565 $Y=3.33
+ $X2=0.24 $Y2=3.33
r101 28 42 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.88 $Y=3.33
+ $X2=3.6 $Y2=3.33
r102 28 39 0.468274 $w=4.9e-07 $l=1.68e-06 $layer=MET1_cond $X=2.88 $Y=3.33
+ $X2=1.2 $Y2=3.33
r103 24 27 28.2872 $w=3.28e-07 $l=8.1e-07 $layer=LI1_cond $X=5.07 $Y=2.14
+ $X2=5.07 $Y2=2.95
r104 22 60 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.07 $Y=3.245
+ $X2=5.07 $Y2=3.33
r105 22 27 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=5.07 $Y=3.245
+ $X2=5.07 $Y2=2.95
r106 18 21 13.9823 $w=7.08e-07 $l=8.3e-07 $layer=LI1_cond $X=4.02 $Y=2.12
+ $X2=4.02 $Y2=2.95
r107 16 57 2.89202 $w=7.1e-07 $l=8.5e-08 $layer=LI1_cond $X=4.02 $Y=3.245
+ $X2=4.02 $Y2=3.33
r108 16 21 4.96962 $w=7.08e-07 $l=2.95e-07 $layer=LI1_cond $X=4.02 $Y=3.245
+ $X2=4.02 $Y2=2.95
r109 12 15 32.1287 $w=3.28e-07 $l=9.2e-07 $layer=LI1_cond $X=0.73 $Y=2.03
+ $X2=0.73 $Y2=2.95
r110 10 54 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=3.245
+ $X2=0.73 $Y2=3.33
r111 10 15 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.73 $Y=3.245
+ $X2=0.73 $Y2=2.95
r112 3 27 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=4.93
+ $Y=1.835 $X2=5.07 $Y2=2.95
r113 3 24 400 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_PDIFF $count=1 $X=4.93
+ $Y=1.835 $X2=5.07 $Y2=2.14
r114 2 21 200 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=3 $X=3.69
+ $Y=1.835 $X2=3.83 $Y2=2.95
r115 2 18 200 $w=1.7e-07 $l=3.4803e-07 $layer=licon1_PDIFF $count=3 $X=3.69
+ $Y=1.835 $X2=3.83 $Y2=2.12
r116 1 15 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=0.59
+ $Y=1.835 $X2=0.73 $Y2=2.95
r117 1 12 400 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_PDIFF $count=1 $X=0.59
+ $Y=1.835 $X2=0.73 $Y2=2.03
.ends

.subckt PM_SKY130_FD_SC_LP__O311AI_2%A_290_367# 1 2 9 13 14 17
r24 17 20 27.2396 $w=3.28e-07 $l=7.8e-07 $layer=LI1_cond $X=2.97 $Y=2.12
+ $X2=2.97 $Y2=2.9
r25 15 20 0.174613 $w=3.28e-07 $l=5e-09 $layer=LI1_cond $X=2.97 $Y=2.905
+ $X2=2.97 $Y2=2.9
r26 13 15 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.805 $Y=2.99
+ $X2=2.97 $Y2=2.905
r27 13 14 68.5027 $w=1.68e-07 $l=1.05e-06 $layer=LI1_cond $X=2.805 $Y=2.99
+ $X2=1.755 $Y2=2.99
r28 9 12 30.3826 $w=3.28e-07 $l=8.7e-07 $layer=LI1_cond $X=1.59 $Y=2.03 $X2=1.59
+ $Y2=2.9
r29 7 14 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.59 $Y=2.905
+ $X2=1.755 $Y2=2.99
r30 7 12 0.174613 $w=3.28e-07 $l=5e-09 $layer=LI1_cond $X=1.59 $Y=2.905 $X2=1.59
+ $Y2=2.9
r31 2 20 400 $w=1.7e-07 $l=1.13284e-06 $layer=licon1_PDIFF $count=1 $X=2.83
+ $Y=1.835 $X2=2.97 $Y2=2.9
r32 2 17 400 $w=1.7e-07 $l=3.4803e-07 $layer=licon1_PDIFF $count=1 $X=2.83
+ $Y=1.835 $X2=2.97 $Y2=2.12
r33 1 12 400 $w=1.7e-07 $l=1.13284e-06 $layer=licon1_PDIFF $count=1 $X=1.45
+ $Y=1.835 $X2=1.59 $Y2=2.9
r34 1 9 400 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_PDIFF $count=1 $X=1.45
+ $Y=1.835 $X2=1.59 $Y2=2.03
.ends

.subckt PM_SKY130_FD_SC_LP__O311AI_2%Y 1 2 3 4 5 6 21 23 24 27 31 35 39 41 43 47
+ 51 52 58 59 69
r81 66 69 0.535558 $w=6.68e-07 $l=3e-08 $layer=LI1_cond $X=4.79 $Y=1.695
+ $X2=4.79 $Y2=1.665
r82 59 66 0.769716 $w=6.7e-07 $l=3.35e-07 $layer=LI1_cond $X=4.455 $Y=1.695
+ $X2=4.79 $Y2=1.695
r83 59 69 0.499854 $w=6.68e-07 $l=2.8e-08 $layer=LI1_cond $X=4.79 $Y=1.637
+ $X2=4.79 $Y2=1.665
r84 58 59 15.5046 $w=2.03e-07 $l=2.8e-07 $layer=LI1_cond $X=5.405 $Y=1.8
+ $X2=5.125 $Y2=1.8
r85 54 55 7.10805 $w=4.72e-07 $l=2.75e-07 $layer=LI1_cond $X=4.79 $Y=0.68
+ $X2=4.79 $Y2=0.955
r86 52 59 10.6576 $w=6.68e-07 $l=5.97e-07 $layer=LI1_cond $X=4.79 $Y=1.04
+ $X2=4.79 $Y2=1.637
r87 52 55 2.62839 $w=6.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.79 $Y=1.04 $X2=4.79
+ $Y2=0.955
r88 47 49 41.222 $w=2.58e-07 $l=9.3e-07 $layer=LI1_cond $X=5.535 $Y=1.98
+ $X2=5.535 $Y2=2.91
r89 45 58 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=5.535 $Y=1.885
+ $X2=5.405 $Y2=1.8
r90 45 47 4.21085 $w=2.58e-07 $l=9.5e-08 $layer=LI1_cond $X=5.535 $Y=1.885
+ $X2=5.535 $Y2=1.98
r91 41 57 2.81454 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.53 $Y=0.87 $X2=5.53
+ $Y2=0.955
r92 41 43 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=5.53 $Y=0.87
+ $X2=5.53 $Y2=0.5
r93 40 55 6.79641 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=5.125 $Y=0.955
+ $X2=4.79 $Y2=0.955
r94 39 57 4.47015 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=5.395 $Y=0.955
+ $X2=5.53 $Y2=0.955
r95 39 40 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=5.395 $Y=0.955
+ $X2=5.125 $Y2=0.955
r96 35 37 54.2871 $w=1.88e-07 $l=9.3e-07 $layer=LI1_cond $X=4.64 $Y=1.98
+ $X2=4.64 $Y2=2.91
r97 33 59 0.769716 $w=1.9e-07 $l=2.66927e-07 $layer=LI1_cond $X=4.64 $Y=1.885
+ $X2=4.455 $Y2=1.695
r98 33 35 5.54545 $w=1.88e-07 $l=9.5e-08 $layer=LI1_cond $X=4.64 $Y=1.885
+ $X2=4.64 $Y2=1.98
r99 32 51 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=3.495 $Y=1.78 $X2=3.4
+ $Y2=1.78
r100 31 59 6.23798 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.455 $Y=1.78
+ $X2=4.455 $Y2=1.695
r101 31 32 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=4.455 $Y=1.78
+ $X2=3.495 $Y2=1.78
r102 27 29 54.2871 $w=1.88e-07 $l=9.3e-07 $layer=LI1_cond $X=3.4 $Y=1.98 $X2=3.4
+ $Y2=2.91
r103 25 51 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=3.4 $Y=1.865
+ $X2=3.4 $Y2=1.78
r104 25 27 6.71292 $w=1.88e-07 $l=1.15e-07 $layer=LI1_cond $X=3.4 $Y=1.865
+ $X2=3.4 $Y2=1.98
r105 23 51 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=3.305 $Y=1.78
+ $X2=3.4 $Y2=1.78
r106 23 24 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.305 $Y=1.78
+ $X2=2.635 $Y2=1.78
r107 19 24 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=2.505 $Y=1.865
+ $X2=2.635 $Y2=1.78
r108 19 21 5.09734 $w=2.58e-07 $l=1.15e-07 $layer=LI1_cond $X=2.505 $Y=1.865
+ $X2=2.505 $Y2=1.98
r109 6 49 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=5.36
+ $Y=1.835 $X2=5.5 $Y2=2.91
r110 6 47 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=5.36
+ $Y=1.835 $X2=5.5 $Y2=1.98
r111 5 37 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=4.5
+ $Y=1.835 $X2=4.64 $Y2=2.91
r112 5 35 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=4.5
+ $Y=1.835 $X2=4.64 $Y2=1.98
r113 4 29 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=3.26
+ $Y=1.835 $X2=3.4 $Y2=2.91
r114 4 27 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=3.26
+ $Y=1.835 $X2=3.4 $Y2=1.98
r115 3 21 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=2.415
+ $Y=1.835 $X2=2.54 $Y2=1.98
r116 2 57 182 $w=1.7e-07 $l=6.76387e-07 $layer=licon1_NDIFF $count=1 $X=5.36
+ $Y=0.345 $X2=5.5 $Y2=0.955
r117 2 43 182 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=1 $X=5.36
+ $Y=0.345 $X2=5.5 $Y2=0.5
r118 1 54 91 $w=1.7e-07 $l=3.92556e-07 $layer=licon1_NDIFF $count=2 $X=4.515
+ $Y=0.345 $X2=4.64 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_LP__O311AI_2%A_35_47# 1 2 3 4 5 16 18 20 24 26 30 32 36
+ 38 43 45 47 49
r63 49 51 7.5352 $w=2.58e-07 $l=1.7e-07 $layer=LI1_cond $X=4.155 $Y=0.76
+ $X2=4.155 $Y2=0.93
r64 39 47 5.53942 $w=1.7e-07 $l=9.3e-08 $layer=LI1_cond $X=3.355 $Y=0.93
+ $X2=3.262 $Y2=0.93
r65 38 51 3.22376 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=4.025 $Y=0.93
+ $X2=4.155 $Y2=0.93
r66 38 39 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.025 $Y=0.93
+ $X2=3.355 $Y2=0.93
r67 34 47 1.03991 $w=1.85e-07 $l=8.5e-08 $layer=LI1_cond $X=3.262 $Y=0.845
+ $X2=3.262 $Y2=0.93
r68 34 36 25.4791 $w=1.83e-07 $l=4.25e-07 $layer=LI1_cond $X=3.262 $Y=0.845
+ $X2=3.262 $Y2=0.42
r69 33 45 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=2.155 $Y=0.93
+ $X2=2.04 $Y2=0.93
r70 32 47 5.53942 $w=1.7e-07 $l=9.2e-08 $layer=LI1_cond $X=3.17 $Y=0.93
+ $X2=3.262 $Y2=0.93
r71 32 33 66.2193 $w=1.68e-07 $l=1.015e-06 $layer=LI1_cond $X=3.17 $Y=0.93
+ $X2=2.155 $Y2=0.93
r72 28 45 0.280307 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.04 $Y=0.845
+ $X2=2.04 $Y2=0.93
r73 28 30 21.2951 $w=2.28e-07 $l=4.25e-07 $layer=LI1_cond $X=2.04 $Y=0.845
+ $X2=2.04 $Y2=0.42
r74 27 43 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.255 $Y=0.93
+ $X2=1.16 $Y2=0.93
r75 26 45 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=1.925 $Y=0.93
+ $X2=2.04 $Y2=0.93
r76 26 27 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.925 $Y=0.93
+ $X2=1.255 $Y2=0.93
r77 22 43 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.16 $Y=0.845
+ $X2=1.16 $Y2=0.93
r78 22 24 24.8086 $w=1.88e-07 $l=4.25e-07 $layer=LI1_cond $X=1.16 $Y=0.845
+ $X2=1.16 $Y2=0.42
r79 21 41 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.395 $Y=0.93
+ $X2=0.265 $Y2=0.93
r80 20 43 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.065 $Y=0.93
+ $X2=1.16 $Y2=0.93
r81 20 21 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.065 $Y=0.93
+ $X2=0.395 $Y2=0.93
r82 16 41 2.85134 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=0.265 $Y=0.845
+ $X2=0.265 $Y2=0.93
r83 16 18 18.838 $w=2.58e-07 $l=4.25e-07 $layer=LI1_cond $X=0.265 $Y=0.845
+ $X2=0.265 $Y2=0.42
r84 5 49 182 $w=1.7e-07 $l=5.90868e-07 $layer=licon1_NDIFF $count=1 $X=3.98
+ $Y=0.235 $X2=4.12 $Y2=0.76
r85 4 47 182 $w=1.7e-07 $l=7.61791e-07 $layer=licon1_NDIFF $count=1 $X=3.12
+ $Y=0.235 $X2=3.26 $Y2=0.93
r86 4 36 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=3.12
+ $Y=0.235 $X2=3.26 $Y2=0.42
r87 3 45 182 $w=1.7e-07 $l=7.68603e-07 $layer=licon1_NDIFF $count=1 $X=1.88
+ $Y=0.235 $X2=2.035 $Y2=0.93
r88 3 30 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=1.88
+ $Y=0.235 $X2=2.035 $Y2=0.42
r89 2 43 182 $w=1.7e-07 $l=7.61791e-07 $layer=licon1_NDIFF $count=1 $X=1.02
+ $Y=0.235 $X2=1.16 $Y2=0.93
r90 2 24 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=1.02
+ $Y=0.235 $X2=1.16 $Y2=0.42
r91 1 41 182 $w=1.7e-07 $l=7.54917e-07 $layer=licon1_NDIFF $count=1 $X=0.175
+ $Y=0.235 $X2=0.3 $Y2=0.93
r92 1 18 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=0.175
+ $Y=0.235 $X2=0.3 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__O311AI_2%VGND 1 2 3 12 16 19 20 21 23 32 41 42 45
r68 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r69 41 42 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r70 39 42 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=3.12 $Y=0 $X2=5.52
+ $Y2=0
r71 38 41 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=3.12 $Y=0 $X2=5.52
+ $Y2=0
r72 38 39 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r73 36 38 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=3 $Y=0 $X2=3.12
+ $Y2=0
r74 35 50 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r75 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r76 32 52 9.74582 $w=6.73e-07 $l=5.5e-07 $layer=LI1_cond $X=2.662 $Y=0 $X2=2.662
+ $Y2=0.55
r77 32 36 9.08255 $w=1.7e-07 $l=3.38e-07 $layer=LI1_cond $X=2.662 $Y=0 $X2=3
+ $Y2=0
r78 32 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r79 32 34 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=2.325 $Y=0 $X2=2.16
+ $Y2=0
r80 31 35 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r81 31 46 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r82 30 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r83 28 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.895 $Y=0 $X2=0.73
+ $Y2=0
r84 28 30 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.895 $Y=0 $X2=1.2
+ $Y2=0
r85 26 46 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r86 25 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r87 23 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.565 $Y=0 $X2=0.73
+ $Y2=0
r88 23 25 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.565 $Y=0 $X2=0.24
+ $Y2=0
r89 21 39 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.88 $Y=0 $X2=3.12
+ $Y2=0
r90 21 50 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.88 $Y=0 $X2=2.64
+ $Y2=0
r91 19 30 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=1.425 $Y=0 $X2=1.2
+ $Y2=0
r92 19 20 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.425 $Y=0 $X2=1.59
+ $Y2=0
r93 18 34 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=1.755 $Y=0 $X2=2.16
+ $Y2=0
r94 18 20 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.755 $Y=0 $X2=1.59
+ $Y2=0
r95 14 20 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.59 $Y=0.085
+ $X2=1.59 $Y2=0
r96 14 16 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=1.59 $Y=0.085
+ $X2=1.59 $Y2=0.55
r97 10 45 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=0.085
+ $X2=0.73 $Y2=0
r98 10 12 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=0.73 $Y=0.085
+ $X2=0.73 $Y2=0.55
r99 3 52 91 $w=1.7e-07 $l=6.17738e-07 $layer=licon1_NDIFF $count=2 $X=2.35
+ $Y=0.235 $X2=2.83 $Y2=0.55
r100 2 16 182 $w=1.7e-07 $l=3.78583e-07 $layer=licon1_NDIFF $count=1 $X=1.45
+ $Y=0.235 $X2=1.59 $Y2=0.55
r101 1 12 182 $w=1.7e-07 $l=3.78583e-07 $layer=licon1_NDIFF $count=1 $X=0.59
+ $Y=0.235 $X2=0.73 $Y2=0.55
.ends

.subckt PM_SKY130_FD_SC_LP__O311AI_2%A_710_47# 1 2 7 11 13
c26 7 0 6.04418e-20 $X=4.975 $Y=0.34
r27 13 16 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=3.69 $Y=0.34
+ $X2=3.69 $Y2=0.55
r28 9 11 5.07075 $w=2.48e-07 $l=1.1e-07 $layer=LI1_cond $X=5.1 $Y=0.425 $X2=5.1
+ $Y2=0.535
r29 8 13 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.855 $Y=0.34
+ $X2=3.69 $Y2=0.34
r30 7 9 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=4.975 $Y=0.34
+ $X2=5.1 $Y2=0.425
r31 7 8 73.0695 $w=1.68e-07 $l=1.12e-06 $layer=LI1_cond $X=4.975 $Y=0.34
+ $X2=3.855 $Y2=0.34
r32 2 11 182 $w=1.7e-07 $l=2.504e-07 $layer=licon1_NDIFF $count=1 $X=4.93
+ $Y=0.345 $X2=5.07 $Y2=0.535
r33 1 16 182 $w=1.7e-07 $l=3.78583e-07 $layer=licon1_NDIFF $count=1 $X=3.55
+ $Y=0.235 $X2=3.69 $Y2=0.55
.ends

