* File: sky130_fd_sc_lp__o2bb2a_0.spice
* Created: Fri Aug 28 11:11:29 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__o2bb2a_0.pex.spice"
.subckt sky130_fd_sc_lp__o2bb2a_0  VNB VPB A1_N A2_N B2 B1 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* B1	B1
* B2	B2
* A2_N	A2_N
* A1_N	A1_N
* VPB	VPB
* VNB	VNB
MM1002 N_VGND_M1002_d N_A_80_176#_M1002_g N_X_M1002_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75001
+ A=0.063 P=1.14 MULT=1
MM1003 A_224_70# N_A1_N_M1003_g N_VGND_M1002_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.0588 PD=0.66 PS=0.7 NRD=18.564 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1004 N_A_229_483#_M1004_d N_A2_N_M1004_g A_224_70# VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.0504 PD=1.37 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75001
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1001 N_A_512_47#_M1001_d N_A_229_483#_M1001_g N_A_80_176#_M1001_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1010 N_VGND_M1010_d N_B2_M1010_g N_A_512_47#_M1001_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1000 N_A_512_47#_M1000_d N_B1_M1000_g N_VGND_M1010_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.1 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1005 N_VPWR_M1005_d N_A_80_176#_M1005_g N_X_M1005_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.148045 AS=0.1696 PD=1.31019 PS=1.81 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75002 A=0.096 P=1.58 MULT=1
MM1007 N_A_229_483#_M1007_d N_A1_N_M1007_g N_VPWR_M1005_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.08925 AS=0.0971547 PD=0.845 PS=0.859811 NRD=68.0044 NRS=79.7259
+ M=1 R=2.8 SA=75000.8 SB=75002.4 A=0.063 P=1.14 MULT=1
MM1009 N_VPWR_M1009_d N_A2_N_M1009_g N_A_229_483#_M1007_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1449 AS=0.08925 PD=1.11 PS=0.845 NRD=178.226 NRS=0 M=1 R=2.8
+ SA=75001.4 SB=75001.8 A=0.063 P=1.14 MULT=1
MM1011 N_A_80_176#_M1011_d N_A_229_483#_M1011_g N_VPWR_M1009_d VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.0588 AS=0.1449 PD=0.7 PS=1.11 NRD=0 NRS=14.0658 M=1 R=2.8
+ SA=75002.2 SB=75001 A=0.063 P=1.14 MULT=1
MM1008 A_598_483# N_B2_M1008_g N_A_80_176#_M1011_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=23.443 NRS=0 M=1 R=2.8 SA=75002.6
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1006 N_VPWR_M1006_d N_B1_M1006_g A_598_483# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.1113 AS=0.0441 PD=1.37 PS=0.63 NRD=0 NRS=23.443 M=1 R=2.8 SA=75003
+ SB=75000.2 A=0.063 P=1.14 MULT=1
DX12_noxref VNB VPB NWDIODE A=7.8703 P=12.17
c_95 VPB 0 1.4009e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_lp__o2bb2a_0.pxi.spice"
*
.ends
*
*
