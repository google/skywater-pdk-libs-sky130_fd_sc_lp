* NGSPICE file created from sky130_fd_sc_lp__and4_lp.ext - technology: sky130A

.subckt sky130_fd_sc_lp__and4_lp A B C D VGND VNB VPB VPWR X
M1000 a_230_55# D VGND VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=2.856e+11p ps=3.04e+06u
M1001 a_422_55# B a_308_55# VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=1.764e+11p ps=1.68e+06u
M1002 a_186_485# A a_422_55# VNB nshort w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=0p ps=0u
M1003 a_186_485# B a_430_485# VPB phighvt w=420000u l=150000u
+  ad=2.352e+11p pd=2.8e+06u as=8.82e+10p ps=1.26e+06u
M1004 a_186_485# D a_114_485# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1005 a_114_485# D VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=3.549e+11p ps=4.21e+06u
M1006 a_720_55# a_186_485# VGND VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1007 a_430_485# B VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_746_485# a_186_485# VPWR VPB phighvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1009 X a_186_485# a_746_485# VPB phighvt w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=0p ps=0u
M1010 X a_186_485# a_720_55# VNB nshort w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=0p ps=0u
M1011 a_272_485# C a_186_485# VPB phighvt w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1012 VPWR A a_588_485# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1013 a_588_485# A a_186_485# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_308_55# C a_230_55# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VPWR C a_272_485# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

