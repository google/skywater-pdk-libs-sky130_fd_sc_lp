* File: sky130_fd_sc_lp__o311a_1.pxi.spice
* Created: Wed Sep  2 10:22:53 2020
* 
x_PM_SKY130_FD_SC_LP__O311A_1%A_80_21# N_A_80_21#_M1008_d N_A_80_21#_M1000_d
+ N_A_80_21#_M1009_d N_A_80_21#_M1003_g N_A_80_21#_M1002_g N_A_80_21#_c_64_n
+ N_A_80_21#_c_70_n N_A_80_21#_c_71_n N_A_80_21#_c_134_p N_A_80_21#_c_72_n
+ N_A_80_21#_c_65_n N_A_80_21#_c_74_n N_A_80_21#_c_75_n N_A_80_21#_c_76_n
+ N_A_80_21#_c_66_n N_A_80_21#_c_67_n PM_SKY130_FD_SC_LP__O311A_1%A_80_21#
x_PM_SKY130_FD_SC_LP__O311A_1%A1 N_A1_M1011_g N_A1_M1006_g A1 A1 A1 N_A1_c_157_n
+ N_A1_c_158_n PM_SKY130_FD_SC_LP__O311A_1%A1
x_PM_SKY130_FD_SC_LP__O311A_1%A2 N_A2_M1010_g N_A2_M1001_g A2 N_A2_c_196_n
+ N_A2_c_197_n PM_SKY130_FD_SC_LP__O311A_1%A2
x_PM_SKY130_FD_SC_LP__O311A_1%A3 N_A3_M1000_g N_A3_M1005_g A3 N_A3_c_225_n
+ N_A3_c_226_n N_A3_c_227_n PM_SKY130_FD_SC_LP__O311A_1%A3
x_PM_SKY130_FD_SC_LP__O311A_1%B1 N_B1_M1004_g N_B1_M1007_g B1 N_B1_c_255_n
+ N_B1_c_256_n N_B1_c_257_n PM_SKY130_FD_SC_LP__O311A_1%B1
x_PM_SKY130_FD_SC_LP__O311A_1%C1 N_C1_c_284_n N_C1_M1008_g N_C1_M1009_g C1
+ N_C1_c_287_n PM_SKY130_FD_SC_LP__O311A_1%C1
x_PM_SKY130_FD_SC_LP__O311A_1%X N_X_M1003_s N_X_M1002_s X X X X X X X
+ N_X_c_309_n X X PM_SKY130_FD_SC_LP__O311A_1%X
x_PM_SKY130_FD_SC_LP__O311A_1%VPWR N_VPWR_M1002_d N_VPWR_M1004_d N_VPWR_c_330_n
+ N_VPWR_c_331_n N_VPWR_c_332_n N_VPWR_c_333_n N_VPWR_c_334_n N_VPWR_c_335_n
+ VPWR N_VPWR_c_336_n N_VPWR_c_329_n PM_SKY130_FD_SC_LP__O311A_1%VPWR
x_PM_SKY130_FD_SC_LP__O311A_1%VGND N_VGND_M1003_d N_VGND_M1001_d N_VGND_c_374_n
+ N_VGND_c_375_n VGND N_VGND_c_376_n N_VGND_c_377_n N_VGND_c_378_n
+ N_VGND_c_379_n N_VGND_c_380_n N_VGND_c_381_n PM_SKY130_FD_SC_LP__O311A_1%VGND
x_PM_SKY130_FD_SC_LP__O311A_1%A_267_47# N_A_267_47#_M1011_d N_A_267_47#_M1005_d
+ N_A_267_47#_c_423_n N_A_267_47#_c_427_n N_A_267_47#_c_425_n
+ N_A_267_47#_c_434_n N_A_267_47#_c_444_n PM_SKY130_FD_SC_LP__O311A_1%A_267_47#
cc_1 VNB N_A_80_21#_M1003_g 0.0318906f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.655
cc_2 VNB N_A_80_21#_c_64_n 0.00366302f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.51
cc_3 VNB N_A_80_21#_c_65_n 0.00455367f $X=-0.19 $Y=-0.245 $X2=3.16 $Y2=1.705
cc_4 VNB N_A_80_21#_c_66_n 0.0317416f $X=-0.19 $Y=-0.245 $X2=3.455 $Y2=0.38
cc_5 VNB N_A_80_21#_c_67_n 0.033389f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.51
cc_6 VNB N_A1_M1006_g 0.00813787f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB A1 0.00134793f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB A1 0.0037497f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.345
cc_9 VNB N_A1_c_157_n 0.0336228f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=2.465
cc_10 VNB N_A1_c_158_n 0.0189532f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A2_M1010_g 0.00775149f $X=-0.19 $Y=-0.245 $X2=3.315 $Y2=1.835
cc_12 VNB A2 0.00376427f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A2_c_196_n 0.0304839f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.655
cc_14 VNB N_A2_c_197_n 0.0185224f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A3_M1000_g 0.00821743f $X=-0.19 $Y=-0.245 $X2=3.315 $Y2=1.835
cc_16 VNB N_A3_c_225_n 0.0296729f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.655
cc_17 VNB N_A3_c_226_n 0.00307435f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.655
cc_18 VNB N_A3_c_227_n 0.0188983f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_B1_M1004_g 0.00858759f $X=-0.19 $Y=-0.245 $X2=3.315 $Y2=1.835
cc_20 VNB N_B1_c_255_n 0.0302847f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.655
cc_21 VNB N_B1_c_256_n 0.00420217f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.655
cc_22 VNB N_B1_c_257_n 0.0169089f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_C1_c_284_n 0.0216661f $X=-0.19 $Y=-0.245 $X2=3.315 $Y2=0.235
cc_24 VNB N_C1_M1009_g 0.0103577f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB C1 0.0178007f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_C1_c_287_n 0.0502813f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_X_c_309_n 0.0622952f $X=-0.19 $Y=-0.245 $X2=2.425 $Y2=1.875
cc_28 VNB N_VPWR_c_329_n 0.163682f $X=-0.19 $Y=-0.245 $X2=3.485 $Y2=2.91
cc_29 VNB N_VGND_c_374_n 0.00958724f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_375_n 0.00561756f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_376_n 0.0182379f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_377_n 0.0272945f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_378_n 0.0454905f $X=-0.19 $Y=-0.245 $X2=2.425 $Y2=2.91
cc_34 VNB N_VGND_c_379_n 0.213666f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_380_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=3.16 $Y2=1.015
cc_36 VNB N_VGND_c_381_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=3.515 $Y2=1.98
cc_37 VPB N_A_80_21#_M1002_g 0.0237876f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=2.465
cc_38 VPB N_A_80_21#_c_64_n 2.68374e-19 $X=-0.19 $Y=1.655 $X2=0.63 $Y2=1.51
cc_39 VPB N_A_80_21#_c_70_n 0.0205106f $X=-0.19 $Y=1.655 $X2=2.26 $Y2=1.79
cc_40 VPB N_A_80_21#_c_71_n 0.00122076f $X=-0.19 $Y=1.655 $X2=0.795 $Y2=1.79
cc_41 VPB N_A_80_21#_c_72_n 0.0059616f $X=-0.19 $Y=1.655 $X2=3.075 $Y2=1.79
cc_42 VPB N_A_80_21#_c_65_n 7.87286e-19 $X=-0.19 $Y=1.655 $X2=3.16 $Y2=1.705
cc_43 VPB N_A_80_21#_c_74_n 0.0104494f $X=-0.19 $Y=1.655 $X2=3.515 $Y2=1.875
cc_44 VPB N_A_80_21#_c_75_n 0.0457335f $X=-0.19 $Y=1.655 $X2=3.485 $Y2=1.98
cc_45 VPB N_A_80_21#_c_76_n 0.00604273f $X=-0.19 $Y=1.655 $X2=2.425 $Y2=1.79
cc_46 VPB N_A_80_21#_c_67_n 0.00899059f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=1.51
cc_47 VPB N_A1_M1006_g 0.0203593f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_48 VPB N_A2_M1010_g 0.0194782f $X=-0.19 $Y=1.655 $X2=3.315 $Y2=1.835
cc_49 VPB N_A3_M1000_g 0.0205113f $X=-0.19 $Y=1.655 $X2=3.315 $Y2=1.835
cc_50 VPB N_B1_M1004_g 0.0213866f $X=-0.19 $Y=1.655 $X2=3.315 $Y2=1.835
cc_51 VPB N_C1_M1009_g 0.0258702f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_52 VPB X 0.0150733f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.655
cc_53 VPB N_X_c_309_n 0.0212121f $X=-0.19 $Y=1.655 $X2=2.425 $Y2=1.875
cc_54 VPB X 0.039458f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_55 VPB N_VPWR_c_330_n 0.0055721f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_56 VPB N_VPWR_c_331_n 0.00561589f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=2.465
cc_57 VPB N_VPWR_c_332_n 0.023359f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=1.51
cc_58 VPB N_VPWR_c_333_n 0.00631825f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=1.51
cc_59 VPB N_VPWR_c_334_n 0.0487205f $X=-0.19 $Y=1.655 $X2=2.26 $Y2=1.79
cc_60 VPB N_VPWR_c_335_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0.795 $Y2=1.79
cc_61 VPB N_VPWR_c_336_n 0.0222157f $X=-0.19 $Y=1.655 $X2=3.515 $Y2=2.91
cc_62 VPB N_VPWR_c_329_n 0.0508749f $X=-0.19 $Y=1.655 $X2=3.485 $Y2=2.91
cc_63 N_A_80_21#_c_64_n N_A1_M1006_g 0.0010934f $X=0.63 $Y=1.51 $X2=0 $Y2=0
cc_64 N_A_80_21#_c_70_n N_A1_M1006_g 0.0157503f $X=2.26 $Y=1.79 $X2=0 $Y2=0
cc_65 N_A_80_21#_c_67_n N_A1_M1006_g 0.0318058f $X=0.72 $Y=1.51 $X2=0 $Y2=0
cc_66 N_A_80_21#_M1003_g A1 0.00224812f $X=0.475 $Y=0.655 $X2=0 $Y2=0
cc_67 N_A_80_21#_M1003_g A1 7.70814e-19 $X=0.475 $Y=0.655 $X2=0 $Y2=0
cc_68 N_A_80_21#_c_64_n A1 0.00802539f $X=0.63 $Y=1.51 $X2=0 $Y2=0
cc_69 N_A_80_21#_c_70_n A1 0.0181796f $X=2.26 $Y=1.79 $X2=0 $Y2=0
cc_70 N_A_80_21#_c_67_n A1 5.43409e-19 $X=0.72 $Y=1.51 $X2=0 $Y2=0
cc_71 N_A_80_21#_M1003_g N_A1_c_157_n 0.0038878f $X=0.475 $Y=0.655 $X2=0 $Y2=0
cc_72 N_A_80_21#_c_64_n N_A1_c_157_n 6.29449e-19 $X=0.63 $Y=1.51 $X2=0 $Y2=0
cc_73 N_A_80_21#_c_70_n N_A1_c_157_n 0.00365927f $X=2.26 $Y=1.79 $X2=0 $Y2=0
cc_74 N_A_80_21#_c_67_n N_A1_c_157_n 0.0106594f $X=0.72 $Y=1.51 $X2=0 $Y2=0
cc_75 N_A_80_21#_M1003_g N_A1_c_158_n 0.0126802f $X=0.475 $Y=0.655 $X2=0 $Y2=0
cc_76 N_A_80_21#_c_70_n N_A2_M1010_g 0.0157853f $X=2.26 $Y=1.79 $X2=0 $Y2=0
cc_77 N_A_80_21#_c_70_n A2 0.018261f $X=2.26 $Y=1.79 $X2=0 $Y2=0
cc_78 N_A_80_21#_c_70_n N_A2_c_196_n 0.00434588f $X=2.26 $Y=1.79 $X2=0 $Y2=0
cc_79 N_A_80_21#_c_70_n N_A3_M1000_g 0.0151631f $X=2.26 $Y=1.79 $X2=0 $Y2=0
cc_80 N_A_80_21#_c_70_n N_A3_c_225_n 5.5094e-19 $X=2.26 $Y=1.79 $X2=0 $Y2=0
cc_81 N_A_80_21#_c_76_n N_A3_c_225_n 0.00578812f $X=2.425 $Y=1.79 $X2=0 $Y2=0
cc_82 N_A_80_21#_c_70_n N_A3_c_226_n 0.0144248f $X=2.26 $Y=1.79 $X2=0 $Y2=0
cc_83 N_A_80_21#_c_76_n N_A3_c_226_n 0.00581771f $X=2.425 $Y=1.79 $X2=0 $Y2=0
cc_84 N_A_80_21#_c_72_n N_B1_M1004_g 0.0162358f $X=3.075 $Y=1.79 $X2=0 $Y2=0
cc_85 N_A_80_21#_c_65_n N_B1_M1004_g 0.00352951f $X=3.16 $Y=1.705 $X2=0 $Y2=0
cc_86 N_A_80_21#_c_72_n N_B1_c_255_n 0.00573264f $X=3.075 $Y=1.79 $X2=0 $Y2=0
cc_87 N_A_80_21#_c_65_n N_B1_c_255_n 0.00588567f $X=3.16 $Y=1.705 $X2=0 $Y2=0
cc_88 N_A_80_21#_c_72_n N_B1_c_256_n 0.0192425f $X=3.075 $Y=1.79 $X2=0 $Y2=0
cc_89 N_A_80_21#_c_65_n N_B1_c_256_n 0.0220977f $X=3.16 $Y=1.705 $X2=0 $Y2=0
cc_90 N_A_80_21#_c_76_n N_B1_c_256_n 0.00695016f $X=2.425 $Y=1.79 $X2=0 $Y2=0
cc_91 N_A_80_21#_c_66_n N_B1_c_257_n 0.00588567f $X=3.455 $Y=0.38 $X2=0 $Y2=0
cc_92 N_A_80_21#_c_65_n N_C1_c_284_n 0.00869829f $X=3.16 $Y=1.705 $X2=-0.19
+ $Y2=-0.245
cc_93 N_A_80_21#_c_66_n N_C1_c_284_n 0.0218292f $X=3.455 $Y=0.38 $X2=-0.19
+ $Y2=-0.245
cc_94 N_A_80_21#_c_65_n N_C1_M1009_g 0.00972202f $X=3.16 $Y=1.705 $X2=0 $Y2=0
cc_95 N_A_80_21#_c_74_n N_C1_M1009_g 0.0175181f $X=3.515 $Y=1.875 $X2=0 $Y2=0
cc_96 N_A_80_21#_c_75_n N_C1_M1009_g 0.0109329f $X=3.485 $Y=1.98 $X2=0 $Y2=0
cc_97 N_A_80_21#_c_65_n C1 0.0224575f $X=3.16 $Y=1.705 $X2=0 $Y2=0
cc_98 N_A_80_21#_c_74_n C1 0.0161974f $X=3.515 $Y=1.875 $X2=0 $Y2=0
cc_99 N_A_80_21#_c_66_n C1 0.0153959f $X=3.455 $Y=0.38 $X2=0 $Y2=0
cc_100 N_A_80_21#_c_65_n N_C1_c_287_n 0.0084316f $X=3.16 $Y=1.705 $X2=0 $Y2=0
cc_101 N_A_80_21#_c_74_n N_C1_c_287_n 0.00910015f $X=3.515 $Y=1.875 $X2=0 $Y2=0
cc_102 N_A_80_21#_c_66_n N_C1_c_287_n 0.00796894f $X=3.455 $Y=0.38 $X2=0 $Y2=0
cc_103 N_A_80_21#_c_71_n N_X_M1002_s 0.00101483f $X=0.795 $Y=1.79 $X2=0 $Y2=0
cc_104 N_A_80_21#_M1002_g X 0.00344243f $X=0.72 $Y=2.465 $X2=0 $Y2=0
cc_105 N_A_80_21#_c_71_n X 0.00664499f $X=0.795 $Y=1.79 $X2=0 $Y2=0
cc_106 N_A_80_21#_c_67_n X 0.00572893f $X=0.72 $Y=1.51 $X2=0 $Y2=0
cc_107 N_A_80_21#_M1003_g N_X_c_309_n 0.022407f $X=0.475 $Y=0.655 $X2=0 $Y2=0
cc_108 N_A_80_21#_M1002_g N_X_c_309_n 0.00492504f $X=0.72 $Y=2.465 $X2=0 $Y2=0
cc_109 N_A_80_21#_c_64_n N_X_c_309_n 0.0276331f $X=0.63 $Y=1.51 $X2=0 $Y2=0
cc_110 N_A_80_21#_c_71_n N_X_c_309_n 0.0147537f $X=0.795 $Y=1.79 $X2=0 $Y2=0
cc_111 N_A_80_21#_M1002_g X 0.00855753f $X=0.72 $Y=2.465 $X2=0 $Y2=0
cc_112 N_A_80_21#_c_70_n N_VPWR_M1002_d 0.00299869f $X=2.26 $Y=1.79 $X2=-0.19
+ $Y2=-0.245
cc_113 N_A_80_21#_c_72_n N_VPWR_M1004_d 0.00263727f $X=3.075 $Y=1.79 $X2=0 $Y2=0
cc_114 N_A_80_21#_c_74_n N_VPWR_M1004_d 3.50796e-19 $X=3.515 $Y=1.875 $X2=0
+ $Y2=0
cc_115 N_A_80_21#_M1002_g N_VPWR_c_330_n 0.00911554f $X=0.72 $Y=2.465 $X2=0
+ $Y2=0
cc_116 N_A_80_21#_c_70_n N_VPWR_c_330_n 0.022455f $X=2.26 $Y=1.79 $X2=0 $Y2=0
cc_117 N_A_80_21#_c_72_n N_VPWR_c_331_n 0.0224185f $X=3.075 $Y=1.79 $X2=0 $Y2=0
cc_118 N_A_80_21#_M1002_g N_VPWR_c_332_n 0.0054895f $X=0.72 $Y=2.465 $X2=0 $Y2=0
cc_119 N_A_80_21#_c_134_p N_VPWR_c_334_n 0.0212513f $X=2.425 $Y=1.98 $X2=0 $Y2=0
cc_120 N_A_80_21#_c_75_n N_VPWR_c_336_n 0.0188974f $X=3.485 $Y=1.98 $X2=0 $Y2=0
cc_121 N_A_80_21#_M1000_d N_VPWR_c_329_n 0.00526034f $X=2.235 $Y=1.835 $X2=0
+ $Y2=0
cc_122 N_A_80_21#_M1009_d N_VPWR_c_329_n 0.00466411f $X=3.315 $Y=1.835 $X2=0
+ $Y2=0
cc_123 N_A_80_21#_M1002_g N_VPWR_c_329_n 0.0112575f $X=0.72 $Y=2.465 $X2=0 $Y2=0
cc_124 N_A_80_21#_c_134_p N_VPWR_c_329_n 0.0127519f $X=2.425 $Y=1.98 $X2=0 $Y2=0
cc_125 N_A_80_21#_c_75_n N_VPWR_c_329_n 0.0104192f $X=3.485 $Y=1.98 $X2=0 $Y2=0
cc_126 N_A_80_21#_c_70_n A_267_367# 0.00690616f $X=2.26 $Y=1.79 $X2=-0.19
+ $Y2=-0.245
cc_127 N_A_80_21#_c_70_n A_356_367# 0.00728771f $X=2.26 $Y=1.79 $X2=-0.19
+ $Y2=-0.245
cc_128 N_A_80_21#_M1003_g N_VGND_c_374_n 0.0109356f $X=0.475 $Y=0.655 $X2=0
+ $Y2=0
cc_129 N_A_80_21#_c_64_n N_VGND_c_374_n 0.013632f $X=0.63 $Y=1.51 $X2=0 $Y2=0
cc_130 N_A_80_21#_c_70_n N_VGND_c_374_n 0.00410457f $X=2.26 $Y=1.79 $X2=0 $Y2=0
cc_131 N_A_80_21#_c_67_n N_VGND_c_374_n 0.00155971f $X=0.72 $Y=1.51 $X2=0 $Y2=0
cc_132 N_A_80_21#_M1003_g N_VGND_c_376_n 0.00585385f $X=0.475 $Y=0.655 $X2=0
+ $Y2=0
cc_133 N_A_80_21#_c_66_n N_VGND_c_378_n 0.0339088f $X=3.455 $Y=0.38 $X2=0 $Y2=0
cc_134 N_A_80_21#_M1008_d N_VGND_c_379_n 0.00215158f $X=3.315 $Y=0.235 $X2=0
+ $Y2=0
cc_135 N_A_80_21#_M1003_g N_VGND_c_379_n 0.012342f $X=0.475 $Y=0.655 $X2=0 $Y2=0
cc_136 N_A_80_21#_c_66_n N_VGND_c_379_n 0.0203511f $X=3.455 $Y=0.38 $X2=0 $Y2=0
cc_137 N_A_80_21#_c_65_n A_591_47# 6.64472e-19 $X=3.16 $Y=1.705 $X2=-0.19
+ $Y2=-0.245
cc_138 N_A_80_21#_c_66_n A_591_47# 0.00841383f $X=3.455 $Y=0.38 $X2=-0.19
+ $Y2=-0.245
cc_139 N_A1_M1006_g N_A2_M1010_g 0.0765723f $X=1.26 $Y=2.465 $X2=0 $Y2=0
cc_140 A1 A2 0.0205786f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_141 N_A1_c_157_n A2 8.16502e-19 $X=1.17 $Y=1.35 $X2=0 $Y2=0
cc_142 A1 N_A2_c_196_n 0.00244711f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_143 N_A1_c_157_n N_A2_c_196_n 0.0212463f $X=1.17 $Y=1.35 $X2=0 $Y2=0
cc_144 A1 N_A2_c_197_n 8.43385e-19 $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_145 N_A1_c_158_n N_A2_c_197_n 0.0216646f $X=1.17 $Y=1.185 $X2=0 $Y2=0
cc_146 N_A1_M1006_g N_VPWR_c_330_n 0.00355844f $X=1.26 $Y=2.465 $X2=0 $Y2=0
cc_147 N_A1_M1006_g N_VPWR_c_334_n 0.00585385f $X=1.26 $Y=2.465 $X2=0 $Y2=0
cc_148 N_A1_M1006_g N_VPWR_c_329_n 0.0109773f $X=1.26 $Y=2.465 $X2=0 $Y2=0
cc_149 A1 N_VGND_M1003_d 0.00721244f $X=1.115 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_150 A1 N_VGND_c_374_n 0.0553397f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_151 N_A1_c_158_n N_VGND_c_374_n 0.00645322f $X=1.17 $Y=1.185 $X2=0 $Y2=0
cc_152 A1 N_VGND_c_377_n 0.00645621f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_153 N_A1_c_158_n N_VGND_c_377_n 0.00451445f $X=1.17 $Y=1.185 $X2=0 $Y2=0
cc_154 A1 N_VGND_c_379_n 0.00669557f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_155 N_A1_c_158_n N_VGND_c_379_n 0.00827112f $X=1.17 $Y=1.185 $X2=0 $Y2=0
cc_156 A1 N_A_267_47#_c_423_n 0.0336717f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_157 N_A1_c_158_n N_A_267_47#_c_423_n 0.00468441f $X=1.17 $Y=1.185 $X2=0 $Y2=0
cc_158 A1 N_A_267_47#_c_425_n 0.0135647f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_159 N_A1_c_158_n N_A_267_47#_c_425_n 0.00132724f $X=1.17 $Y=1.185 $X2=0 $Y2=0
cc_160 N_A2_M1010_g N_A3_M1000_g 0.073321f $X=1.705 $Y=2.465 $X2=0 $Y2=0
cc_161 A2 N_A3_c_225_n 2.86248e-19 $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_162 N_A2_c_196_n N_A3_c_225_n 0.02065f $X=1.71 $Y=1.35 $X2=0 $Y2=0
cc_163 A2 N_A3_c_226_n 0.0197284f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_164 N_A2_c_196_n N_A3_c_226_n 0.00318179f $X=1.71 $Y=1.35 $X2=0 $Y2=0
cc_165 N_A2_c_197_n N_A3_c_227_n 0.0260435f $X=1.71 $Y=1.185 $X2=0 $Y2=0
cc_166 N_A2_M1010_g N_VPWR_c_334_n 0.00585385f $X=1.705 $Y=2.465 $X2=0 $Y2=0
cc_167 N_A2_M1010_g N_VPWR_c_329_n 0.011138f $X=1.705 $Y=2.465 $X2=0 $Y2=0
cc_168 N_A2_c_197_n N_VGND_c_375_n 0.00581236f $X=1.71 $Y=1.185 $X2=0 $Y2=0
cc_169 N_A2_c_197_n N_VGND_c_377_n 0.00585385f $X=1.71 $Y=1.185 $X2=0 $Y2=0
cc_170 N_A2_c_197_n N_VGND_c_379_n 0.00690231f $X=1.71 $Y=1.185 $X2=0 $Y2=0
cc_171 A2 N_A_267_47#_c_427_n 0.0122723f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_172 N_A2_c_197_n N_A_267_47#_c_427_n 0.0107057f $X=1.71 $Y=1.185 $X2=0 $Y2=0
cc_173 A2 N_A_267_47#_c_425_n 0.0107175f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_174 N_A2_c_196_n N_A_267_47#_c_425_n 8.67081e-19 $X=1.71 $Y=1.35 $X2=0 $Y2=0
cc_175 N_A3_M1000_g N_B1_M1004_g 0.0306341f $X=2.16 $Y=2.465 $X2=0 $Y2=0
cc_176 N_A3_c_225_n N_B1_c_255_n 0.0204451f $X=2.25 $Y=1.35 $X2=0 $Y2=0
cc_177 N_A3_c_226_n N_B1_c_255_n 2.86406e-19 $X=2.25 $Y=1.35 $X2=0 $Y2=0
cc_178 N_A3_c_225_n N_B1_c_256_n 0.00219472f $X=2.25 $Y=1.35 $X2=0 $Y2=0
cc_179 N_A3_c_226_n N_B1_c_256_n 0.0262082f $X=2.25 $Y=1.35 $X2=0 $Y2=0
cc_180 N_A3_c_227_n N_B1_c_257_n 0.019799f $X=2.25 $Y=1.185 $X2=0 $Y2=0
cc_181 N_A3_M1000_g N_VPWR_c_334_n 0.00585385f $X=2.16 $Y=2.465 $X2=0 $Y2=0
cc_182 N_A3_M1000_g N_VPWR_c_329_n 0.0112318f $X=2.16 $Y=2.465 $X2=0 $Y2=0
cc_183 N_A3_c_227_n N_VGND_c_375_n 0.0058704f $X=2.25 $Y=1.185 $X2=0 $Y2=0
cc_184 N_A3_c_227_n N_VGND_c_378_n 0.00585385f $X=2.25 $Y=1.185 $X2=0 $Y2=0
cc_185 N_A3_c_227_n N_VGND_c_379_n 0.00708071f $X=2.25 $Y=1.185 $X2=0 $Y2=0
cc_186 N_A3_c_225_n N_A_267_47#_c_427_n 0.00450164f $X=2.25 $Y=1.35 $X2=0 $Y2=0
cc_187 N_A3_c_226_n N_A_267_47#_c_427_n 0.0193377f $X=2.25 $Y=1.35 $X2=0 $Y2=0
cc_188 N_A3_c_227_n N_A_267_47#_c_427_n 0.0153085f $X=2.25 $Y=1.185 $X2=0 $Y2=0
cc_189 N_B1_c_256_n N_C1_c_284_n 3.05388e-19 $X=2.79 $Y=1.35 $X2=-0.19
+ $Y2=-0.245
cc_190 N_B1_c_257_n N_C1_c_284_n 0.042616f $X=2.79 $Y=1.185 $X2=-0.19 $Y2=-0.245
cc_191 N_B1_M1004_g N_C1_c_287_n 0.0292819f $X=2.7 $Y=2.465 $X2=0 $Y2=0
cc_192 N_B1_c_255_n N_C1_c_287_n 0.042616f $X=2.79 $Y=1.35 $X2=0 $Y2=0
cc_193 N_B1_M1004_g N_VPWR_c_331_n 0.00348909f $X=2.7 $Y=2.465 $X2=0 $Y2=0
cc_194 N_B1_M1004_g N_VPWR_c_334_n 0.00585385f $X=2.7 $Y=2.465 $X2=0 $Y2=0
cc_195 N_B1_M1004_g N_VPWR_c_329_n 0.0112268f $X=2.7 $Y=2.465 $X2=0 $Y2=0
cc_196 N_B1_c_257_n N_VGND_c_378_n 0.00585385f $X=2.79 $Y=1.185 $X2=0 $Y2=0
cc_197 N_B1_c_257_n N_VGND_c_379_n 0.0109726f $X=2.79 $Y=1.185 $X2=0 $Y2=0
cc_198 N_B1_c_255_n N_A_267_47#_c_434_n 0.00410495f $X=2.79 $Y=1.35 $X2=0 $Y2=0
cc_199 N_B1_c_256_n N_A_267_47#_c_434_n 0.0217667f $X=2.79 $Y=1.35 $X2=0 $Y2=0
cc_200 N_C1_M1009_g N_VPWR_c_331_n 0.00930086f $X=3.24 $Y=2.465 $X2=0 $Y2=0
cc_201 N_C1_M1009_g N_VPWR_c_336_n 0.00585385f $X=3.24 $Y=2.465 $X2=0 $Y2=0
cc_202 N_C1_M1009_g N_VPWR_c_329_n 0.0120174f $X=3.24 $Y=2.465 $X2=0 $Y2=0
cc_203 N_C1_c_284_n N_VGND_c_378_n 0.00357668f $X=3.24 $Y=1.195 $X2=0 $Y2=0
cc_204 N_C1_c_284_n N_VGND_c_379_n 0.0062144f $X=3.24 $Y=1.195 $X2=0 $Y2=0
cc_205 X N_VPWR_c_332_n 0.0386099f $X=0.24 $Y=2.405 $X2=0 $Y2=0
cc_206 N_X_M1002_s N_VPWR_c_329_n 0.00215158f $X=0.38 $Y=1.835 $X2=0 $Y2=0
cc_207 X N_VPWR_c_329_n 0.0220939f $X=0.24 $Y=2.405 $X2=0 $Y2=0
cc_208 N_X_c_309_n N_VGND_c_374_n 0.00129956f $X=0.26 $Y=0.42 $X2=0 $Y2=0
cc_209 N_X_c_309_n N_VGND_c_376_n 0.0181659f $X=0.26 $Y=0.42 $X2=0 $Y2=0
cc_210 N_X_M1003_s N_VGND_c_379_n 0.00336915f $X=0.135 $Y=0.235 $X2=0 $Y2=0
cc_211 N_X_c_309_n N_VGND_c_379_n 0.0104192f $X=0.26 $Y=0.42 $X2=0 $Y2=0
cc_212 N_VPWR_c_329_n A_267_367# 0.0126346f $X=3.6 $Y=3.33 $X2=-0.19 $Y2=-0.245
cc_213 N_VPWR_c_329_n A_356_367# 0.0130629f $X=3.6 $Y=3.33 $X2=-0.19 $Y2=-0.245
cc_214 N_VGND_c_379_n N_A_267_47#_M1011_d 0.00693542f $X=3.6 $Y=0 $X2=-0.19
+ $Y2=-0.245
cc_215 N_VGND_c_379_n N_A_267_47#_M1005_d 0.00423472f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_216 N_VGND_c_374_n N_A_267_47#_c_423_n 0.00410639f $X=0.75 $Y=0.38 $X2=0
+ $Y2=0
cc_217 N_VGND_c_377_n N_A_267_47#_c_423_n 0.0135517f $X=1.885 $Y=0 $X2=0 $Y2=0
cc_218 N_VGND_c_379_n N_A_267_47#_c_423_n 0.00847534f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_219 N_VGND_M1001_d N_A_267_47#_c_427_n 0.0115133f $X=1.83 $Y=0.235 $X2=0
+ $Y2=0
cc_220 N_VGND_c_375_n N_A_267_47#_c_427_n 0.0255547f $X=2.05 $Y=0.55 $X2=0 $Y2=0
cc_221 N_VGND_c_379_n N_A_267_47#_c_427_n 0.0141077f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_222 N_VGND_c_378_n N_A_267_47#_c_444_n 0.0212513f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_223 N_VGND_c_379_n N_A_267_47#_c_444_n 0.0127519f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_224 N_VGND_c_379_n A_591_47# 0.00589804f $X=3.6 $Y=0 $X2=-0.19 $Y2=-0.245
