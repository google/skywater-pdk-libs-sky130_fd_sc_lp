* File: sky130_fd_sc_lp__o2bb2a_4.pxi.spice
* Created: Wed Sep  2 10:21:35 2020
* 
x_PM_SKY130_FD_SC_LP__O2BB2A_4%B1 N_B1_M1006_g N_B1_M1011_g N_B1_M1026_g
+ N_B1_M1009_g N_B1_c_132_n N_B1_c_133_n N_B1_c_139_n N_B1_c_140_n N_B1_c_134_n
+ N_B1_c_135_n N_B1_c_144_p B1 B1 B1 PM_SKY130_FD_SC_LP__O2BB2A_4%B1
x_PM_SKY130_FD_SC_LP__O2BB2A_4%B2 N_B2_M1014_g N_B2_M1008_g N_B2_M1024_g
+ N_B2_M1021_g B2 N_B2_c_224_n N_B2_c_221_n PM_SKY130_FD_SC_LP__O2BB2A_4%B2
x_PM_SKY130_FD_SC_LP__O2BB2A_4%A_462_21# N_A_462_21#_M1016_d N_A_462_21#_M1000_s
+ N_A_462_21#_M1020_s N_A_462_21#_c_273_n N_A_462_21#_M1003_g
+ N_A_462_21#_M1001_g N_A_462_21#_c_275_n N_A_462_21#_M1015_g
+ N_A_462_21#_M1019_g N_A_462_21#_c_277_n N_A_462_21#_c_278_n
+ N_A_462_21#_c_279_n N_A_462_21#_c_280_n N_A_462_21#_c_281_n
+ N_A_462_21#_c_328_p N_A_462_21#_c_295_p N_A_462_21#_c_282_n
+ N_A_462_21#_c_297_p N_A_462_21#_c_303_p PM_SKY130_FD_SC_LP__O2BB2A_4%A_462_21#
x_PM_SKY130_FD_SC_LP__O2BB2A_4%A1_N N_A1_N_M1000_g N_A1_N_M1004_g N_A1_N_M1007_g
+ N_A1_N_M1022_g N_A1_N_c_391_n N_A1_N_c_392_n N_A1_N_c_393_n A1_N
+ N_A1_N_c_394_n N_A1_N_c_395_n N_A1_N_c_396_n N_A1_N_c_397_n
+ PM_SKY130_FD_SC_LP__O2BB2A_4%A1_N
x_PM_SKY130_FD_SC_LP__O2BB2A_4%A2_N N_A2_N_c_477_n N_A2_N_M1012_g N_A2_N_c_473_n
+ N_A2_N_M1016_g N_A2_N_c_474_n N_A2_N_M1025_g N_A2_N_c_478_n N_A2_N_M1020_g
+ A2_N N_A2_N_c_475_n N_A2_N_c_476_n PM_SKY130_FD_SC_LP__O2BB2A_4%A2_N
x_PM_SKY130_FD_SC_LP__O2BB2A_4%A_218_367# N_A_218_367#_M1003_s
+ N_A_218_367#_M1008_d N_A_218_367#_M1001_d N_A_218_367#_M1010_g
+ N_A_218_367#_M1002_g N_A_218_367#_M1018_g N_A_218_367#_M1005_g
+ N_A_218_367#_M1023_g N_A_218_367#_M1013_g N_A_218_367#_M1027_g
+ N_A_218_367#_M1017_g N_A_218_367#_c_546_n N_A_218_367#_c_529_n
+ N_A_218_367#_c_530_n N_A_218_367#_c_573_n N_A_218_367#_c_575_n
+ N_A_218_367#_c_541_n N_A_218_367#_c_580_n N_A_218_367#_c_583_n
+ N_A_218_367#_c_584_n N_A_218_367#_c_531_n N_A_218_367#_c_532_n
+ N_A_218_367#_c_656_p N_A_218_367#_c_533_n N_A_218_367#_c_534_n
+ N_A_218_367#_c_598_n N_A_218_367#_c_535_n
+ PM_SKY130_FD_SC_LP__O2BB2A_4%A_218_367#
x_PM_SKY130_FD_SC_LP__O2BB2A_4%VPWR N_VPWR_M1011_d N_VPWR_M1026_d N_VPWR_M1019_s
+ N_VPWR_M1012_d N_VPWR_M1022_d N_VPWR_M1018_s N_VPWR_M1027_s N_VPWR_c_712_n
+ N_VPWR_c_713_n N_VPWR_c_740_n N_VPWR_c_714_n N_VPWR_c_715_n N_VPWR_c_716_n
+ N_VPWR_c_717_n N_VPWR_c_718_n N_VPWR_c_719_n N_VPWR_c_720_n N_VPWR_c_721_n
+ N_VPWR_c_722_n N_VPWR_c_723_n N_VPWR_c_724_n N_VPWR_c_725_n N_VPWR_c_726_n
+ VPWR N_VPWR_c_727_n N_VPWR_c_728_n N_VPWR_c_711_n N_VPWR_c_730_n
+ N_VPWR_c_731_n N_VPWR_c_732_n N_VPWR_c_733_n PM_SKY130_FD_SC_LP__O2BB2A_4%VPWR
x_PM_SKY130_FD_SC_LP__O2BB2A_4%A_132_367# N_A_132_367#_M1011_s
+ N_A_132_367#_M1021_s N_A_132_367#_c_839_n
+ PM_SKY130_FD_SC_LP__O2BB2A_4%A_132_367#
x_PM_SKY130_FD_SC_LP__O2BB2A_4%X N_X_M1002_s N_X_M1013_s N_X_M1010_d N_X_M1023_d
+ N_X_c_894_n N_X_c_857_n N_X_c_858_n N_X_c_872_n N_X_c_851_n N_X_c_852_n
+ N_X_c_898_n N_X_c_859_n N_X_c_909_p N_X_c_853_n N_X_c_860_n N_X_c_854_n X X
+ N_X_c_855_n N_X_c_861_n X X PM_SKY130_FD_SC_LP__O2BB2A_4%X
x_PM_SKY130_FD_SC_LP__O2BB2A_4%A_49_47# N_A_49_47#_M1006_d N_A_49_47#_M1014_d
+ N_A_49_47#_M1009_d N_A_49_47#_M1015_d N_A_49_47#_c_914_n N_A_49_47#_c_915_n
+ N_A_49_47#_c_916_n N_A_49_47#_c_957_p N_A_49_47#_c_922_n N_A_49_47#_c_923_n
+ N_A_49_47#_c_924_n N_A_49_47#_c_935_n N_A_49_47#_c_937_n
+ PM_SKY130_FD_SC_LP__O2BB2A_4%A_49_47#
x_PM_SKY130_FD_SC_LP__O2BB2A_4%VGND N_VGND_M1006_s N_VGND_M1024_s N_VGND_M1004_d
+ N_VGND_M1007_d N_VGND_M1005_d N_VGND_M1017_d N_VGND_c_973_n N_VGND_c_974_n
+ N_VGND_c_975_n N_VGND_c_976_n N_VGND_c_977_n N_VGND_c_978_n N_VGND_c_979_n
+ VGND N_VGND_c_980_n N_VGND_c_981_n N_VGND_c_982_n N_VGND_c_983_n
+ N_VGND_c_984_n N_VGND_c_985_n N_VGND_c_986_n N_VGND_c_987_n N_VGND_c_988_n
+ N_VGND_c_989_n N_VGND_c_990_n N_VGND_c_991_n PM_SKY130_FD_SC_LP__O2BB2A_4%VGND
x_PM_SKY130_FD_SC_LP__O2BB2A_4%A_768_47# N_A_768_47#_M1004_s N_A_768_47#_M1025_s
+ N_A_768_47#_c_1094_n N_A_768_47#_c_1099_n N_A_768_47#_c_1100_n
+ PM_SKY130_FD_SC_LP__O2BB2A_4%A_768_47#
cc_1 VNB N_B1_M1006_g 0.0313103f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=0.655
cc_2 VNB N_B1_M1009_g 0.0252295f $X=-0.19 $Y=-0.245 $X2=1.955 $Y2=0.655
cc_3 VNB N_B1_c_132_n 0.0121847f $X=-0.19 $Y=-0.245 $X2=0.625 $Y2=1.525
cc_4 VNB N_B1_c_133_n 0.0300535f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.51
cc_5 VNB N_B1_c_134_n 9.12083e-19 $X=-0.19 $Y=-0.245 $X2=1.93 $Y2=1.51
cc_6 VNB N_B1_c_135_n 0.0273938f $X=-0.19 $Y=-0.245 $X2=1.93 $Y2=1.51
cc_7 VNB N_B2_M1014_g 0.0229706f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=0.655
cc_8 VNB N_B2_M1024_g 0.024141f $X=-0.19 $Y=-0.245 $X2=1.875 $Y2=2.465
cc_9 VNB N_B2_c_221_n 0.0311857f $X=-0.19 $Y=-0.245 $X2=1.935 $Y2=1.65
cc_10 VNB N_A_462_21#_c_273_n 0.015373f $X=-0.19 $Y=-0.245 $X2=1.875 $Y2=2.465
cc_11 VNB N_A_462_21#_M1001_g 0.00719562f $X=-0.19 $Y=-0.245 $X2=1.955 $Y2=0.655
cc_12 VNB N_A_462_21#_c_275_n 0.0193362f $X=-0.19 $Y=-0.245 $X2=0.625 $Y2=1.525
cc_13 VNB N_A_462_21#_M1019_g 0.00856736f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.645
cc_14 VNB N_A_462_21#_c_277_n 0.00849724f $X=-0.19 $Y=-0.245 $X2=1.935 $Y2=1.65
cc_15 VNB N_A_462_21#_c_278_n 0.0701814f $X=-0.19 $Y=-0.245 $X2=1.93 $Y2=1.51
cc_16 VNB N_A_462_21#_c_279_n 0.0041688f $X=-0.19 $Y=-0.245 $X2=1.97 $Y2=1.65
cc_17 VNB N_A_462_21#_c_280_n 0.0032246f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=2.32
cc_18 VNB N_A_462_21#_c_281_n 0.00390097f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=2.32
cc_19 VNB N_A_462_21#_c_282_n 0.00322666f $X=-0.19 $Y=-0.245 $X2=1.93 $Y2=1.51
cc_20 VNB N_A1_N_M1000_g 0.00884745f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=0.655
cc_21 VNB N_A1_N_M1022_g 0.00784026f $X=-0.19 $Y=-0.245 $X2=1.955 $Y2=1.345
cc_22 VNB N_A1_N_c_391_n 0.00823115f $X=-0.19 $Y=-0.245 $X2=1.955 $Y2=0.655
cc_23 VNB N_A1_N_c_392_n 0.00686402f $X=-0.19 $Y=-0.245 $X2=0.625 $Y2=1.525
cc_24 VNB N_A1_N_c_393_n 0.0357139f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A1_N_c_394_n 0.0327889f $X=-0.19 $Y=-0.245 $X2=1.97 $Y2=1.51
cc_26 VNB N_A1_N_c_395_n 0.0196769f $X=-0.19 $Y=-0.245 $X2=1.93 $Y2=1.51
cc_27 VNB N_A1_N_c_396_n 0.0178263f $X=-0.19 $Y=-0.245 $X2=1.845 $Y2=2.405
cc_28 VNB N_A1_N_c_397_n 0.00691783f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A2_N_c_473_n 0.0154647f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A2_N_c_474_n 0.0154648f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=2.465
cc_31 VNB N_A2_N_c_475_n 0.00239161f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.51
cc_32 VNB N_A2_N_c_476_n 0.0450571f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.51
cc_33 VNB N_A_218_367#_M1002_g 0.0265723f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_218_367#_M1005_g 0.0217542f $X=-0.19 $Y=-0.245 $X2=1.935 $Y2=1.65
cc_35 VNB N_A_218_367#_M1013_g 0.0217348f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=2.32
cc_36 VNB N_A_218_367#_M1017_g 0.026556f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.675
cc_37 VNB N_A_218_367#_c_529_n 0.00353491f $X=-0.19 $Y=-0.245 $X2=1.68 $Y2=2.405
cc_38 VNB N_A_218_367#_c_530_n 0.0116889f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_218_367#_c_531_n 7.60855e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_218_367#_c_532_n 0.0033928f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_218_367#_c_533_n 0.00217252f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_218_367#_c_534_n 0.00134096f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_218_367#_c_535_n 0.0900397f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VPWR_c_711_n 0.322901f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_X_c_851_n 0.00305125f $X=-0.19 $Y=-0.245 $X2=1.935 $Y2=2.31
cc_46 VNB N_X_c_852_n 0.00186402f $X=-0.19 $Y=-0.245 $X2=1.97 $Y2=1.51
cc_47 VNB N_X_c_853_n 0.00237025f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.345
cc_48 VNB N_X_c_854_n 0.00144145f $X=-0.19 $Y=-0.245 $X2=1.93 $Y2=1.345
cc_49 VNB N_X_c_855_n 0.0137041f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=2.405
cc_50 VNB X 0.0222072f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_49_47#_c_914_n 0.0307328f $X=-0.19 $Y=-0.245 $X2=1.955 $Y2=0.655
cc_52 VNB N_A_49_47#_c_915_n 0.0088442f $X=-0.19 $Y=-0.245 $X2=0.625 $Y2=1.525
cc_53 VNB N_A_49_47#_c_916_n 0.0104404f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.525
cc_54 VNB N_VGND_c_973_n 3.99129e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_974_n 0.00274299f $X=-0.19 $Y=-0.245 $X2=1.935 $Y2=2.31
cc_56 VNB N_VGND_c_975_n 0.00875184f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_VGND_c_976_n 0.00602402f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=2.32
cc_58 VNB N_VGND_c_977_n 3.20903e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_978_n 0.0132365f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.345
cc_60 VNB N_VGND_c_979_n 0.0276525f $X=-0.19 $Y=-0.245 $X2=1.93 $Y2=1.51
cc_61 VNB N_VGND_c_980_n 0.0188763f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=2.405
cc_62 VNB N_VGND_c_981_n 0.0122054f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_VGND_c_982_n 0.0375643f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_VGND_c_983_n 0.0363525f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_VGND_c_984_n 0.0154314f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_VGND_c_985_n 0.0129398f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_986_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_VGND_c_987_n 0.00510247f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_VGND_c_988_n 0.00497021f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_VGND_c_989_n 0.0101874f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_VGND_c_990_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_VGND_c_991_n 0.382849f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VPB N_B1_M1011_g 0.0249715f $X=-0.19 $Y=1.655 $X2=0.585 $Y2=2.465
cc_74 VPB N_B1_M1026_g 0.0203427f $X=-0.19 $Y=1.655 $X2=1.875 $Y2=2.465
cc_75 VPB N_B1_c_133_n 0.00779349f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=1.51
cc_76 VPB N_B1_c_139_n 0.00135025f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=2.31
cc_77 VPB N_B1_c_140_n 0.00159562f $X=-0.19 $Y=1.655 $X2=1.935 $Y2=2.31
cc_78 VPB N_B1_c_135_n 0.00845424f $X=-0.19 $Y=1.655 $X2=1.93 $Y2=1.51
cc_79 VPB N_B2_M1008_g 0.0186664f $X=-0.19 $Y=1.655 $X2=0.585 $Y2=2.465
cc_80 VPB N_B2_M1021_g 0.0181024f $X=-0.19 $Y=1.655 $X2=1.955 $Y2=0.655
cc_81 VPB N_B2_c_224_n 0.00257788f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=2.31
cc_82 VPB N_B2_c_221_n 0.00471835f $X=-0.19 $Y=1.655 $X2=1.935 $Y2=1.65
cc_83 VPB N_A_462_21#_M1001_g 0.0216684f $X=-0.19 $Y=1.655 $X2=1.955 $Y2=0.655
cc_84 VPB N_A_462_21#_M1019_g 0.0223584f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=1.645
cc_85 VPB N_A_462_21#_c_280_n 0.00441782f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=2.32
cc_86 VPB N_A1_N_M1000_g 0.0231615f $X=-0.19 $Y=1.655 $X2=0.585 $Y2=0.655
cc_87 VPB N_A1_N_M1022_g 0.0210551f $X=-0.19 $Y=1.655 $X2=1.955 $Y2=1.345
cc_88 VPB N_A2_N_c_477_n 0.0163781f $X=-0.19 $Y=1.655 $X2=0.585 $Y2=1.345
cc_89 VPB N_A2_N_c_478_n 0.0161343f $X=-0.19 $Y=1.655 $X2=1.875 $Y2=2.465
cc_90 VPB N_A2_N_c_475_n 0.00374811f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=1.51
cc_91 VPB N_A2_N_c_476_n 0.0100019f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=1.51
cc_92 VPB N_A_218_367#_M1010_g 0.0198983f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_93 VPB N_A_218_367#_M1018_g 0.018773f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=1.51
cc_94 VPB N_A_218_367#_M1023_g 0.0187796f $X=-0.19 $Y=1.655 $X2=1.93 $Y2=1.51
cc_95 VPB N_A_218_367#_M1027_g 0.02291f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_96 VPB N_A_218_367#_c_529_n 0.00108378f $X=-0.19 $Y=1.655 $X2=1.68 $Y2=2.405
cc_97 VPB N_A_218_367#_c_541_n 0.00431174f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_98 VPB N_A_218_367#_c_531_n 0.00175231f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_99 VPB N_A_218_367#_c_534_n 6.64243e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_100 VPB N_A_218_367#_c_535_n 0.0141506f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_101 VPB N_VPWR_c_712_n 0.013523f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=1.645
cc_102 VPB N_VPWR_c_713_n 0.0558008f $X=-0.19 $Y=1.655 $X2=1.935 $Y2=1.65
cc_103 VPB N_VPWR_c_714_n 0.00310059f $X=-0.19 $Y=1.655 $X2=1.845 $Y2=2.405
cc_104 VPB N_VPWR_c_715_n 0.00374296f $X=-0.19 $Y=1.655 $X2=1.595 $Y2=2.32
cc_105 VPB N_VPWR_c_716_n 3.11597e-19 $X=-0.19 $Y=1.655 $X2=0.495 $Y2=1.675
cc_106 VPB N_VPWR_c_717_n 0.00214221f $X=-0.19 $Y=1.655 $X2=0.815 $Y2=2.405
cc_107 VPB N_VPWR_c_718_n 3.21684e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_108 VPB N_VPWR_c_719_n 0.0130339f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_109 VPB N_VPWR_c_720_n 0.0415892f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_110 VPB N_VPWR_c_721_n 0.0127224f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_111 VPB N_VPWR_c_722_n 0.00436638f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_112 VPB N_VPWR_c_723_n 0.0131493f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_113 VPB N_VPWR_c_724_n 0.00510611f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_114 VPB N_VPWR_c_725_n 0.0160952f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_115 VPB N_VPWR_c_726_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_116 VPB N_VPWR_c_727_n 0.0367428f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_117 VPB N_VPWR_c_728_n 0.0164632f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_118 VPB N_VPWR_c_711_n 0.0634202f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_119 VPB N_VPWR_c_730_n 0.00814565f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_120 VPB N_VPWR_c_731_n 0.0149992f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_121 VPB N_VPWR_c_732_n 0.0122128f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_122 VPB N_VPWR_c_733_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_123 VPB N_X_c_857_n 0.00301161f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=1.51
cc_124 VPB N_X_c_858_n 0.00210491f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=1.51
cc_125 VPB N_X_c_859_n 0.00959411f $X=-0.19 $Y=1.655 $X2=1.115 $Y2=2.32
cc_126 VPB N_X_c_860_n 0.00134754f $X=-0.19 $Y=1.655 $X2=1.93 $Y2=1.51
cc_127 VPB N_X_c_861_n 0.0190924f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_128 VPB X 0.00510498f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_129 N_B1_M1006_g N_B2_M1014_g 0.0296913f $X=0.585 $Y=0.655 $X2=0 $Y2=0
cc_130 N_B1_M1011_g N_B2_M1008_g 0.0296913f $X=0.585 $Y=2.465 $X2=0 $Y2=0
cc_131 N_B1_c_144_p N_B2_M1008_g 0.0125979f $X=1.845 $Y=2.405 $X2=0 $Y2=0
cc_132 N_B1_M1009_g N_B2_M1024_g 0.0338702f $X=1.955 $Y=0.655 $X2=0 $Y2=0
cc_133 N_B1_M1026_g N_B2_M1021_g 0.0511566f $X=1.875 $Y=2.465 $X2=0 $Y2=0
cc_134 N_B1_c_140_n N_B2_M1021_g 0.00133763f $X=1.935 $Y=2.31 $X2=0 $Y2=0
cc_135 N_B1_c_144_p N_B2_M1021_g 0.0111993f $X=1.845 $Y=2.405 $X2=0 $Y2=0
cc_136 N_B1_c_132_n N_B2_c_224_n 0.0196889f $X=0.625 $Y=1.525 $X2=0 $Y2=0
cc_137 N_B1_c_133_n N_B2_c_224_n 3.26233e-19 $X=0.495 $Y=1.51 $X2=0 $Y2=0
cc_138 N_B1_c_139_n N_B2_c_224_n 0.00864051f $X=0.72 $Y=2.31 $X2=0 $Y2=0
cc_139 N_B1_c_132_n N_B2_c_221_n 0.00192742f $X=0.625 $Y=1.525 $X2=0 $Y2=0
cc_140 N_B1_c_133_n N_B2_c_221_n 0.0296913f $X=0.495 $Y=1.51 $X2=0 $Y2=0
cc_141 N_B1_c_139_n N_B2_c_221_n 0.00779709f $X=0.72 $Y=2.31 $X2=0 $Y2=0
cc_142 N_B1_c_134_n N_B2_c_221_n 3.63568e-19 $X=1.93 $Y=1.51 $X2=0 $Y2=0
cc_143 N_B1_c_135_n N_B2_c_221_n 0.0168093f $X=1.93 $Y=1.51 $X2=0 $Y2=0
cc_144 N_B1_M1009_g N_A_462_21#_c_273_n 0.0264884f $X=1.955 $Y=0.655 $X2=0 $Y2=0
cc_145 N_B1_M1026_g N_A_462_21#_M1001_g 0.0150834f $X=1.875 $Y=2.465 $X2=0 $Y2=0
cc_146 N_B1_c_140_n N_A_462_21#_M1001_g 0.00164293f $X=1.935 $Y=2.31 $X2=0 $Y2=0
cc_147 N_B1_c_134_n N_A_462_21#_M1001_g 5.05442e-19 $X=1.93 $Y=1.51 $X2=0 $Y2=0
cc_148 N_B1_c_135_n N_A_462_21#_M1001_g 0.0046216f $X=1.93 $Y=1.51 $X2=0 $Y2=0
cc_149 N_B1_c_134_n N_A_462_21#_c_278_n 8.11235e-19 $X=1.93 $Y=1.51 $X2=0 $Y2=0
cc_150 N_B1_c_135_n N_A_462_21#_c_278_n 0.011224f $X=1.93 $Y=1.51 $X2=0 $Y2=0
cc_151 N_B1_c_144_p N_A_218_367#_M1008_d 0.0034413f $X=1.845 $Y=2.405 $X2=0
+ $Y2=0
cc_152 N_B1_M1026_g N_A_218_367#_c_546_n 0.0014675f $X=1.875 $Y=2.465 $X2=0
+ $Y2=0
cc_153 N_B1_c_139_n N_A_218_367#_c_546_n 0.0164762f $X=0.72 $Y=2.31 $X2=0 $Y2=0
cc_154 N_B1_c_140_n N_A_218_367#_c_546_n 0.015919f $X=1.935 $Y=2.31 $X2=0 $Y2=0
cc_155 N_B1_c_144_p N_A_218_367#_c_546_n 0.0373125f $X=1.845 $Y=2.405 $X2=0
+ $Y2=0
cc_156 N_B1_M1026_g N_A_218_367#_c_529_n 0.00154737f $X=1.875 $Y=2.465 $X2=0
+ $Y2=0
cc_157 N_B1_M1009_g N_A_218_367#_c_529_n 0.00347515f $X=1.955 $Y=0.655 $X2=0
+ $Y2=0
cc_158 N_B1_c_139_n N_A_218_367#_c_529_n 0.0041491f $X=0.72 $Y=2.31 $X2=0 $Y2=0
cc_159 N_B1_c_134_n N_A_218_367#_c_529_n 0.040718f $X=1.93 $Y=1.51 $X2=0 $Y2=0
cc_160 N_B1_c_135_n N_A_218_367#_c_529_n 0.00223682f $X=1.93 $Y=1.51 $X2=0 $Y2=0
cc_161 N_B1_M1009_g N_A_218_367#_c_530_n 0.0112304f $X=1.955 $Y=0.655 $X2=0
+ $Y2=0
cc_162 N_B1_c_134_n N_A_218_367#_c_530_n 0.0190017f $X=1.93 $Y=1.51 $X2=0 $Y2=0
cc_163 N_B1_c_135_n N_A_218_367#_c_530_n 0.00393324f $X=1.93 $Y=1.51 $X2=0 $Y2=0
cc_164 N_B1_M1026_g N_A_218_367#_c_534_n 2.1261e-19 $X=1.875 $Y=2.465 $X2=0
+ $Y2=0
cc_165 N_B1_M1009_g N_A_218_367#_c_534_n 5.98563e-19 $X=1.955 $Y=0.655 $X2=0
+ $Y2=0
cc_166 N_B1_c_140_n N_A_218_367#_c_534_n 0.0041902f $X=1.935 $Y=2.31 $X2=0 $Y2=0
cc_167 N_B1_c_134_n N_A_218_367#_c_534_n 0.00889929f $X=1.93 $Y=1.51 $X2=0 $Y2=0
cc_168 N_B1_c_135_n N_A_218_367#_c_534_n 9.60763e-19 $X=1.93 $Y=1.51 $X2=0 $Y2=0
cc_169 N_B1_c_140_n N_VPWR_M1026_d 0.00442299f $X=1.935 $Y=2.31 $X2=0 $Y2=0
cc_170 N_B1_c_144_p N_VPWR_M1026_d 0.00202754f $X=1.845 $Y=2.405 $X2=0 $Y2=0
cc_171 N_B1_M1011_g N_VPWR_c_713_n 0.00858005f $X=0.585 $Y=2.465 $X2=0 $Y2=0
cc_172 N_B1_c_132_n N_VPWR_c_713_n 0.0102342f $X=0.625 $Y=1.525 $X2=0 $Y2=0
cc_173 N_B1_c_133_n N_VPWR_c_713_n 0.00299509f $X=0.495 $Y=1.51 $X2=0 $Y2=0
cc_174 N_B1_c_139_n N_VPWR_c_713_n 0.0177887f $X=0.72 $Y=2.31 $X2=0 $Y2=0
cc_175 N_B1_M1026_g N_VPWR_c_740_n 0.00418029f $X=1.875 $Y=2.465 $X2=0 $Y2=0
cc_176 N_B1_c_144_p N_VPWR_c_740_n 0.00269489f $X=1.845 $Y=2.405 $X2=0 $Y2=0
cc_177 N_B1_M1026_g N_VPWR_c_714_n 0.00774034f $X=1.875 $Y=2.465 $X2=0 $Y2=0
cc_178 N_B1_M1026_g N_VPWR_c_715_n 0.00604976f $X=1.875 $Y=2.465 $X2=0 $Y2=0
cc_179 N_B1_c_140_n N_VPWR_c_715_n 0.0384426f $X=1.935 $Y=2.31 $X2=0 $Y2=0
cc_180 N_B1_c_144_p N_VPWR_c_715_n 0.0157553f $X=1.845 $Y=2.405 $X2=0 $Y2=0
cc_181 N_B1_M1011_g N_VPWR_c_727_n 0.00535845f $X=0.585 $Y=2.465 $X2=0 $Y2=0
cc_182 N_B1_M1026_g N_VPWR_c_727_n 0.00525069f $X=1.875 $Y=2.465 $X2=0 $Y2=0
cc_183 N_B1_M1011_g N_VPWR_c_711_n 0.0105135f $X=0.585 $Y=2.465 $X2=0 $Y2=0
cc_184 N_B1_M1026_g N_VPWR_c_711_n 0.00494384f $X=1.875 $Y=2.465 $X2=0 $Y2=0
cc_185 N_B1_c_144_p N_VPWR_c_711_n 0.00699733f $X=1.845 $Y=2.405 $X2=0 $Y2=0
cc_186 N_B1_c_139_n N_A_132_367#_M1011_s 0.00611063f $X=0.72 $Y=2.31 $X2=-0.19
+ $Y2=-0.245
cc_187 N_B1_c_144_p N_A_132_367#_M1011_s 0.00329722f $X=1.845 $Y=2.405 $X2=-0.19
+ $Y2=-0.245
cc_188 N_B1_c_144_p N_A_132_367#_M1021_s 0.00569401f $X=1.845 $Y=2.405 $X2=0
+ $Y2=0
cc_189 N_B1_M1011_g N_A_132_367#_c_839_n 0.0045886f $X=0.585 $Y=2.465 $X2=0
+ $Y2=0
cc_190 N_B1_c_139_n N_A_132_367#_c_839_n 0.0106827f $X=0.72 $Y=2.31 $X2=0 $Y2=0
cc_191 N_B1_c_144_p N_A_132_367#_c_839_n 0.0510051f $X=1.845 $Y=2.405 $X2=0
+ $Y2=0
cc_192 N_B1_M1006_g N_A_49_47#_c_915_n 0.0154323f $X=0.585 $Y=0.655 $X2=0 $Y2=0
cc_193 N_B1_c_132_n N_A_49_47#_c_915_n 0.0269924f $X=0.625 $Y=1.525 $X2=0 $Y2=0
cc_194 N_B1_c_133_n N_A_49_47#_c_915_n 0.00108047f $X=0.495 $Y=1.51 $X2=0 $Y2=0
cc_195 N_B1_c_132_n N_A_49_47#_c_916_n 0.0111416f $X=0.625 $Y=1.525 $X2=0 $Y2=0
cc_196 N_B1_c_133_n N_A_49_47#_c_916_n 0.00338214f $X=0.495 $Y=1.51 $X2=0 $Y2=0
cc_197 N_B1_M1009_g N_A_49_47#_c_922_n 0.00968247f $X=1.955 $Y=0.655 $X2=0 $Y2=0
cc_198 N_B1_M1009_g N_A_49_47#_c_923_n 0.00209799f $X=1.955 $Y=0.655 $X2=0 $Y2=0
cc_199 N_B1_M1009_g N_A_49_47#_c_924_n 0.00380015f $X=1.955 $Y=0.655 $X2=0 $Y2=0
cc_200 N_B1_M1006_g N_VGND_c_973_n 0.0127767f $X=0.585 $Y=0.655 $X2=0 $Y2=0
cc_201 N_B1_M1009_g N_VGND_c_974_n 0.00432564f $X=1.955 $Y=0.655 $X2=0 $Y2=0
cc_202 N_B1_M1006_g N_VGND_c_980_n 0.00486043f $X=0.585 $Y=0.655 $X2=0 $Y2=0
cc_203 N_B1_M1009_g N_VGND_c_982_n 0.00416296f $X=1.955 $Y=0.655 $X2=0 $Y2=0
cc_204 N_B1_M1006_g N_VGND_c_991_n 0.00926856f $X=0.585 $Y=0.655 $X2=0 $Y2=0
cc_205 N_B1_M1009_g N_VGND_c_991_n 0.00602095f $X=1.955 $Y=0.655 $X2=0 $Y2=0
cc_206 N_B2_M1008_g N_A_218_367#_c_546_n 0.00605797f $X=1.015 $Y=2.465 $X2=0
+ $Y2=0
cc_207 N_B2_M1021_g N_A_218_367#_c_546_n 0.0116137f $X=1.445 $Y=2.465 $X2=0
+ $Y2=0
cc_208 N_B2_c_224_n N_A_218_367#_c_546_n 0.0233186f $X=1.15 $Y=1.51 $X2=0 $Y2=0
cc_209 N_B2_c_221_n N_A_218_367#_c_546_n 5.72878e-19 $X=1.445 $Y=1.51 $X2=0
+ $Y2=0
cc_210 N_B2_M1014_g N_A_218_367#_c_529_n 5.93281e-19 $X=1.015 $Y=0.655 $X2=0
+ $Y2=0
cc_211 N_B2_M1008_g N_A_218_367#_c_529_n 4.07015e-19 $X=1.015 $Y=2.465 $X2=0
+ $Y2=0
cc_212 N_B2_M1024_g N_A_218_367#_c_529_n 0.00410858f $X=1.445 $Y=0.655 $X2=0
+ $Y2=0
cc_213 N_B2_M1021_g N_A_218_367#_c_529_n 0.00618678f $X=1.445 $Y=2.465 $X2=0
+ $Y2=0
cc_214 N_B2_c_224_n N_A_218_367#_c_529_n 0.0257707f $X=1.15 $Y=1.51 $X2=0 $Y2=0
cc_215 N_B2_c_221_n N_A_218_367#_c_529_n 0.00942339f $X=1.445 $Y=1.51 $X2=0
+ $Y2=0
cc_216 N_B2_M1024_g N_A_218_367#_c_573_n 0.00502252f $X=1.445 $Y=0.655 $X2=0
+ $Y2=0
cc_217 N_B2_M1021_g N_VPWR_c_714_n 0.00143366f $X=1.445 $Y=2.465 $X2=0 $Y2=0
cc_218 N_B2_M1008_g N_VPWR_c_727_n 0.00373071f $X=1.015 $Y=2.465 $X2=0 $Y2=0
cc_219 N_B2_M1021_g N_VPWR_c_727_n 0.00373071f $X=1.445 $Y=2.465 $X2=0 $Y2=0
cc_220 N_B2_M1008_g N_VPWR_c_711_n 0.00548684f $X=1.015 $Y=2.465 $X2=0 $Y2=0
cc_221 N_B2_M1021_g N_VPWR_c_711_n 0.00548684f $X=1.445 $Y=2.465 $X2=0 $Y2=0
cc_222 N_B2_M1008_g N_A_132_367#_c_839_n 0.0122888f $X=1.015 $Y=2.465 $X2=0
+ $Y2=0
cc_223 N_B2_M1021_g N_A_132_367#_c_839_n 0.0123797f $X=1.445 $Y=2.465 $X2=0
+ $Y2=0
cc_224 N_B2_M1014_g N_A_49_47#_c_915_n 0.0150759f $X=1.015 $Y=0.655 $X2=0 $Y2=0
cc_225 N_B2_M1024_g N_A_49_47#_c_915_n 0.00128644f $X=1.445 $Y=0.655 $X2=0 $Y2=0
cc_226 N_B2_c_224_n N_A_49_47#_c_915_n 0.0261363f $X=1.15 $Y=1.51 $X2=0 $Y2=0
cc_227 N_B2_c_221_n N_A_49_47#_c_915_n 0.00250341f $X=1.445 $Y=1.51 $X2=0 $Y2=0
cc_228 N_B2_M1024_g N_A_49_47#_c_922_n 0.0142582f $X=1.445 $Y=0.655 $X2=0 $Y2=0
cc_229 N_B2_M1024_g N_A_49_47#_c_924_n 5.96354e-19 $X=1.445 $Y=0.655 $X2=0 $Y2=0
cc_230 N_B2_M1014_g N_VGND_c_973_n 0.010963f $X=1.015 $Y=0.655 $X2=0 $Y2=0
cc_231 N_B2_M1024_g N_VGND_c_973_n 6.48667e-19 $X=1.445 $Y=0.655 $X2=0 $Y2=0
cc_232 N_B2_M1014_g N_VGND_c_974_n 5.14991e-19 $X=1.015 $Y=0.655 $X2=0 $Y2=0
cc_233 N_B2_M1024_g N_VGND_c_974_n 0.00667144f $X=1.445 $Y=0.655 $X2=0 $Y2=0
cc_234 N_B2_M1014_g N_VGND_c_981_n 0.00486043f $X=1.015 $Y=0.655 $X2=0 $Y2=0
cc_235 N_B2_M1024_g N_VGND_c_981_n 0.00355956f $X=1.445 $Y=0.655 $X2=0 $Y2=0
cc_236 N_B2_M1014_g N_VGND_c_991_n 0.00824727f $X=1.015 $Y=0.655 $X2=0 $Y2=0
cc_237 N_B2_M1024_g N_VGND_c_991_n 0.00415754f $X=1.445 $Y=0.655 $X2=0 $Y2=0
cc_238 N_A_462_21#_M1019_g N_A1_N_M1000_g 0.0187034f $X=2.98 $Y=2.465 $X2=0
+ $Y2=0
cc_239 N_A_462_21#_c_280_n N_A1_N_M1000_g 0.00958101f $X=3.385 $Y=1.93 $X2=0
+ $Y2=0
cc_240 N_A_462_21#_c_295_p N_A1_N_M1000_g 0.015771f $X=4.84 $Y=2.095 $X2=0 $Y2=0
cc_241 N_A_462_21#_c_295_p N_A1_N_c_391_n 0.00797884f $X=4.84 $Y=2.095 $X2=0
+ $Y2=0
cc_242 N_A_462_21#_c_297_p N_A1_N_c_391_n 0.030203f $X=4.41 $Y=0.79 $X2=0 $Y2=0
cc_243 N_A_462_21#_c_295_p N_A1_N_c_392_n 4.99242e-19 $X=4.84 $Y=2.095 $X2=0
+ $Y2=0
cc_244 N_A_462_21#_c_295_p N_A1_N_c_393_n 3.12905e-19 $X=4.84 $Y=2.095 $X2=0
+ $Y2=0
cc_245 N_A_462_21#_c_278_n N_A1_N_c_394_n 0.00900566f $X=3.015 $Y=1.35 $X2=0
+ $Y2=0
cc_246 N_A_462_21#_c_295_p N_A1_N_c_394_n 0.00372901f $X=4.84 $Y=2.095 $X2=0
+ $Y2=0
cc_247 N_A_462_21#_c_282_n N_A1_N_c_394_n 0.00317062f $X=3.385 $Y=1.35 $X2=0
+ $Y2=0
cc_248 N_A_462_21#_c_303_p N_A1_N_c_394_n 0.00254059f $X=4.245 $Y=0.785 $X2=0
+ $Y2=0
cc_249 N_A_462_21#_c_279_n N_A1_N_c_395_n 0.00621905f $X=3.385 $Y=1.185 $X2=0
+ $Y2=0
cc_250 N_A_462_21#_c_297_p N_A1_N_c_395_n 3.37063e-19 $X=4.41 $Y=0.79 $X2=0
+ $Y2=0
cc_251 N_A_462_21#_c_303_p N_A1_N_c_395_n 0.0145161f $X=4.245 $Y=0.785 $X2=0
+ $Y2=0
cc_252 N_A_462_21#_c_278_n N_A1_N_c_397_n 2.41395e-19 $X=3.015 $Y=1.35 $X2=0
+ $Y2=0
cc_253 N_A_462_21#_c_279_n N_A1_N_c_397_n 0.00835496f $X=3.385 $Y=1.185 $X2=0
+ $Y2=0
cc_254 N_A_462_21#_c_295_p N_A1_N_c_397_n 0.0184918f $X=4.84 $Y=2.095 $X2=0
+ $Y2=0
cc_255 N_A_462_21#_c_282_n N_A1_N_c_397_n 0.0284182f $X=3.385 $Y=1.35 $X2=0
+ $Y2=0
cc_256 N_A_462_21#_c_303_p N_A1_N_c_397_n 0.030203f $X=4.245 $Y=0.785 $X2=0
+ $Y2=0
cc_257 N_A_462_21#_c_295_p N_A2_N_c_477_n 0.0146239f $X=4.84 $Y=2.095 $X2=-0.19
+ $Y2=-0.245
cc_258 N_A_462_21#_c_297_p N_A2_N_c_473_n 0.00235948f $X=4.41 $Y=0.79 $X2=0
+ $Y2=0
cc_259 N_A_462_21#_c_303_p N_A2_N_c_473_n 0.00812413f $X=4.245 $Y=0.785 $X2=0
+ $Y2=0
cc_260 N_A_462_21#_c_297_p N_A2_N_c_474_n 0.00328463f $X=4.41 $Y=0.79 $X2=0
+ $Y2=0
cc_261 N_A_462_21#_c_295_p N_A2_N_c_478_n 0.0128888f $X=4.84 $Y=2.095 $X2=0
+ $Y2=0
cc_262 N_A_462_21#_c_295_p N_A2_N_c_475_n 0.0278233f $X=4.84 $Y=2.095 $X2=0
+ $Y2=0
cc_263 N_A_462_21#_c_295_p N_A2_N_c_476_n 7.59994e-19 $X=4.84 $Y=2.095 $X2=0
+ $Y2=0
cc_264 N_A_462_21#_c_297_p N_A2_N_c_476_n 5.59397e-19 $X=4.41 $Y=0.79 $X2=0
+ $Y2=0
cc_265 N_A_462_21#_c_273_n N_A_218_367#_c_530_n 0.0145498f $X=2.385 $Y=1.185
+ $X2=0 $Y2=0
cc_266 N_A_462_21#_c_275_n N_A_218_367#_c_575_n 0.00453825f $X=2.815 $Y=1.185
+ $X2=0 $Y2=0
cc_267 N_A_462_21#_M1001_g N_A_218_367#_c_541_n 0.00370352f $X=2.55 $Y=2.465
+ $X2=0 $Y2=0
cc_268 N_A_462_21#_M1019_g N_A_218_367#_c_541_n 0.00509386f $X=2.98 $Y=2.465
+ $X2=0 $Y2=0
cc_269 N_A_462_21#_c_278_n N_A_218_367#_c_541_n 0.00253535f $X=3.015 $Y=1.35
+ $X2=0 $Y2=0
cc_270 N_A_462_21#_c_280_n N_A_218_367#_c_541_n 0.00836964f $X=3.385 $Y=1.93
+ $X2=0 $Y2=0
cc_271 N_A_462_21#_M1001_g N_A_218_367#_c_580_n 0.00664624f $X=2.55 $Y=2.465
+ $X2=0 $Y2=0
cc_272 N_A_462_21#_M1019_g N_A_218_367#_c_580_n 0.013745f $X=2.98 $Y=2.465 $X2=0
+ $Y2=0
cc_273 N_A_462_21#_c_328_p N_A_218_367#_c_580_n 0.0151697f $X=3.475 $Y=2.095
+ $X2=0 $Y2=0
cc_274 N_A_462_21#_M1001_g N_A_218_367#_c_583_n 0.00622983f $X=2.55 $Y=2.465
+ $X2=0 $Y2=0
cc_275 N_A_462_21#_M1000_s N_A_218_367#_c_584_n 0.00494544f $X=3.825 $Y=1.835
+ $X2=0 $Y2=0
cc_276 N_A_462_21#_M1020_s N_A_218_367#_c_584_n 0.00494544f $X=4.7 $Y=1.835
+ $X2=0 $Y2=0
cc_277 N_A_462_21#_M1019_g N_A_218_367#_c_584_n 0.0139257f $X=2.98 $Y=2.465
+ $X2=0 $Y2=0
cc_278 N_A_462_21#_c_328_p N_A_218_367#_c_584_n 0.0146113f $X=3.475 $Y=2.095
+ $X2=0 $Y2=0
cc_279 N_A_462_21#_c_295_p N_A_218_367#_c_584_n 0.0824557f $X=4.84 $Y=2.095
+ $X2=0 $Y2=0
cc_280 N_A_462_21#_c_275_n N_A_218_367#_c_533_n 0.00545999f $X=2.815 $Y=1.185
+ $X2=0 $Y2=0
cc_281 N_A_462_21#_c_278_n N_A_218_367#_c_533_n 0.00224606f $X=3.015 $Y=1.35
+ $X2=0 $Y2=0
cc_282 N_A_462_21#_c_279_n N_A_218_367#_c_533_n 0.00536954f $X=3.385 $Y=1.185
+ $X2=0 $Y2=0
cc_283 N_A_462_21#_M1001_g N_A_218_367#_c_534_n 0.00547084f $X=2.55 $Y=2.465
+ $X2=0 $Y2=0
cc_284 N_A_462_21#_M1019_g N_A_218_367#_c_534_n 0.00209036f $X=2.98 $Y=2.465
+ $X2=0 $Y2=0
cc_285 N_A_462_21#_c_277_n N_A_218_367#_c_534_n 0.0245279f $X=3.295 $Y=1.35
+ $X2=0 $Y2=0
cc_286 N_A_462_21#_c_278_n N_A_218_367#_c_534_n 0.0180751f $X=3.015 $Y=1.35
+ $X2=0 $Y2=0
cc_287 N_A_462_21#_c_279_n N_A_218_367#_c_534_n 2.60067e-19 $X=3.385 $Y=1.185
+ $X2=0 $Y2=0
cc_288 N_A_462_21#_c_280_n N_A_218_367#_c_534_n 0.00725285f $X=3.385 $Y=1.93
+ $X2=0 $Y2=0
cc_289 N_A_462_21#_M1001_g N_A_218_367#_c_598_n 0.00200683f $X=2.55 $Y=2.465
+ $X2=0 $Y2=0
cc_290 N_A_462_21#_M1019_g N_A_218_367#_c_598_n 0.00101089f $X=2.98 $Y=2.465
+ $X2=0 $Y2=0
cc_291 N_A_462_21#_c_280_n N_VPWR_M1019_s 0.00315926f $X=3.385 $Y=1.93 $X2=0
+ $Y2=0
cc_292 N_A_462_21#_c_328_p N_VPWR_M1019_s 0.00933358f $X=3.475 $Y=2.095 $X2=0
+ $Y2=0
cc_293 N_A_462_21#_c_295_p N_VPWR_M1019_s 0.00638808f $X=4.84 $Y=2.095 $X2=0
+ $Y2=0
cc_294 N_A_462_21#_c_295_p N_VPWR_M1012_d 0.00404813f $X=4.84 $Y=2.095 $X2=0
+ $Y2=0
cc_295 N_A_462_21#_M1001_g N_VPWR_c_715_n 0.00410982f $X=2.55 $Y=2.465 $X2=0
+ $Y2=0
cc_296 N_A_462_21#_c_278_n N_VPWR_c_715_n 0.00318056f $X=3.015 $Y=1.35 $X2=0
+ $Y2=0
cc_297 N_A_462_21#_M1000_s N_VPWR_c_711_n 0.00360572f $X=3.825 $Y=1.835 $X2=0
+ $Y2=0
cc_298 N_A_462_21#_M1020_s N_VPWR_c_711_n 0.00360572f $X=4.7 $Y=1.835 $X2=0
+ $Y2=0
cc_299 N_A_462_21#_M1001_g N_VPWR_c_711_n 0.0100742f $X=2.55 $Y=2.465 $X2=0
+ $Y2=0
cc_300 N_A_462_21#_M1019_g N_VPWR_c_711_n 0.00427368f $X=2.98 $Y=2.465 $X2=0
+ $Y2=0
cc_301 N_A_462_21#_M1001_g N_VPWR_c_731_n 0.00533769f $X=2.55 $Y=2.465 $X2=0
+ $Y2=0
cc_302 N_A_462_21#_M1019_g N_VPWR_c_731_n 0.00363497f $X=2.98 $Y=2.465 $X2=0
+ $Y2=0
cc_303 N_A_462_21#_M1001_g N_VPWR_c_732_n 5.01907e-19 $X=2.55 $Y=2.465 $X2=0
+ $Y2=0
cc_304 N_A_462_21#_M1019_g N_VPWR_c_732_n 0.00872706f $X=2.98 $Y=2.465 $X2=0
+ $Y2=0
cc_305 N_A_462_21#_c_273_n N_A_49_47#_c_922_n 0.00207083f $X=2.385 $Y=1.185
+ $X2=0 $Y2=0
cc_306 N_A_462_21#_c_273_n N_A_49_47#_c_923_n 6.12373e-19 $X=2.385 $Y=1.185
+ $X2=0 $Y2=0
cc_307 N_A_462_21#_c_273_n N_A_49_47#_c_924_n 0.00361715f $X=2.385 $Y=1.185
+ $X2=0 $Y2=0
cc_308 N_A_462_21#_c_275_n N_A_49_47#_c_924_n 4.48149e-19 $X=2.815 $Y=1.185
+ $X2=0 $Y2=0
cc_309 N_A_462_21#_c_273_n N_A_49_47#_c_935_n 0.00849527f $X=2.385 $Y=1.185
+ $X2=0 $Y2=0
cc_310 N_A_462_21#_c_275_n N_A_49_47#_c_935_n 0.0119546f $X=2.815 $Y=1.185 $X2=0
+ $Y2=0
cc_311 N_A_462_21#_c_277_n N_A_49_47#_c_937_n 0.01522f $X=3.295 $Y=1.35 $X2=0
+ $Y2=0
cc_312 N_A_462_21#_c_278_n N_A_49_47#_c_937_n 0.00493639f $X=3.015 $Y=1.35 $X2=0
+ $Y2=0
cc_313 N_A_462_21#_c_279_n N_A_49_47#_c_937_n 0.00746692f $X=3.385 $Y=1.185
+ $X2=0 $Y2=0
cc_314 N_A_462_21#_c_281_n N_A_49_47#_c_937_n 0.0159382f $X=3.475 $Y=0.82 $X2=0
+ $Y2=0
cc_315 N_A_462_21#_c_279_n N_VGND_M1004_d 0.00231432f $X=3.385 $Y=1.185 $X2=0
+ $Y2=0
cc_316 N_A_462_21#_c_281_n N_VGND_M1004_d 0.00106532f $X=3.475 $Y=0.82 $X2=0
+ $Y2=0
cc_317 N_A_462_21#_c_303_p N_VGND_M1004_d 0.00629215f $X=4.245 $Y=0.785 $X2=0
+ $Y2=0
cc_318 N_A_462_21#_c_275_n N_VGND_c_975_n 0.00226038f $X=2.815 $Y=1.185 $X2=0
+ $Y2=0
cc_319 N_A_462_21#_c_281_n N_VGND_c_975_n 0.00782331f $X=3.475 $Y=0.82 $X2=0
+ $Y2=0
cc_320 N_A_462_21#_c_303_p N_VGND_c_975_n 0.0124148f $X=4.245 $Y=0.785 $X2=0
+ $Y2=0
cc_321 N_A_462_21#_c_273_n N_VGND_c_982_n 0.00357842f $X=2.385 $Y=1.185 $X2=0
+ $Y2=0
cc_322 N_A_462_21#_c_275_n N_VGND_c_982_n 0.00357877f $X=2.815 $Y=1.185 $X2=0
+ $Y2=0
cc_323 N_A_462_21#_c_281_n N_VGND_c_982_n 0.00152037f $X=3.475 $Y=0.82 $X2=0
+ $Y2=0
cc_324 N_A_462_21#_c_303_p N_VGND_c_983_n 0.00202355f $X=4.245 $Y=0.785 $X2=0
+ $Y2=0
cc_325 N_A_462_21#_M1016_d N_VGND_c_991_n 0.00225186f $X=4.27 $Y=0.235 $X2=0
+ $Y2=0
cc_326 N_A_462_21#_c_273_n N_VGND_c_991_n 0.00537652f $X=2.385 $Y=1.185 $X2=0
+ $Y2=0
cc_327 N_A_462_21#_c_275_n N_VGND_c_991_n 0.00665089f $X=2.815 $Y=1.185 $X2=0
+ $Y2=0
cc_328 N_A_462_21#_c_281_n N_VGND_c_991_n 0.00298618f $X=3.475 $Y=0.82 $X2=0
+ $Y2=0
cc_329 N_A_462_21#_c_303_p N_VGND_c_991_n 0.00548584f $X=4.245 $Y=0.785 $X2=0
+ $Y2=0
cc_330 N_A_462_21#_c_303_p N_A_768_47#_M1004_s 0.00377994f $X=4.245 $Y=0.785
+ $X2=-0.19 $Y2=-0.245
cc_331 N_A_462_21#_M1016_d N_A_768_47#_c_1094_n 0.0033589f $X=4.27 $Y=0.235
+ $X2=0 $Y2=0
cc_332 N_A_462_21#_c_297_p N_A_768_47#_c_1094_n 0.0154524f $X=4.41 $Y=0.79 $X2=0
+ $Y2=0
cc_333 N_A_462_21#_c_303_p N_A_768_47#_c_1094_n 0.0161465f $X=4.245 $Y=0.785
+ $X2=0 $Y2=0
cc_334 N_A1_N_c_391_n N_A2_N_c_473_n 0.00329748f $X=4.92 $Y=1.17 $X2=0 $Y2=0
cc_335 N_A1_N_c_395_n N_A2_N_c_473_n 0.0349274f $X=3.73 $Y=1.185 $X2=0 $Y2=0
cc_336 N_A1_N_c_397_n N_A2_N_c_473_n 0.00243476f $X=4.175 $Y=1.3 $X2=0 $Y2=0
cc_337 N_A1_N_c_391_n N_A2_N_c_474_n 0.00718805f $X=4.92 $Y=1.17 $X2=0 $Y2=0
cc_338 N_A1_N_c_396_n N_A2_N_c_474_n 0.0181137f $X=5.075 $Y=1.185 $X2=0 $Y2=0
cc_339 N_A1_N_M1000_g N_A2_N_c_475_n 8.35631e-19 $X=3.75 $Y=2.465 $X2=0 $Y2=0
cc_340 N_A1_N_M1022_g N_A2_N_c_475_n 0.00245571f $X=5.055 $Y=2.465 $X2=0 $Y2=0
cc_341 N_A1_N_c_391_n N_A2_N_c_475_n 0.0293508f $X=4.92 $Y=1.17 $X2=0 $Y2=0
cc_342 N_A1_N_c_392_n N_A2_N_c_475_n 0.00709956f $X=5.045 $Y=1.17 $X2=0 $Y2=0
cc_343 N_A1_N_c_393_n N_A2_N_c_475_n 5.28628e-19 $X=5.075 $Y=1.35 $X2=0 $Y2=0
cc_344 N_A1_N_c_397_n N_A2_N_c_475_n 0.00707169f $X=4.175 $Y=1.3 $X2=0 $Y2=0
cc_345 N_A1_N_M1000_g N_A2_N_c_476_n 0.0613841f $X=3.75 $Y=2.465 $X2=0 $Y2=0
cc_346 N_A1_N_M1022_g N_A2_N_c_476_n 0.0595878f $X=5.055 $Y=2.465 $X2=0 $Y2=0
cc_347 N_A1_N_c_391_n N_A2_N_c_476_n 0.0154165f $X=4.92 $Y=1.17 $X2=0 $Y2=0
cc_348 N_A1_N_c_392_n N_A2_N_c_476_n 0.00140148f $X=5.045 $Y=1.17 $X2=0 $Y2=0
cc_349 N_A1_N_c_393_n N_A2_N_c_476_n 0.0221724f $X=5.075 $Y=1.35 $X2=0 $Y2=0
cc_350 N_A1_N_c_394_n N_A2_N_c_476_n 0.0197277f $X=3.73 $Y=1.35 $X2=0 $Y2=0
cc_351 N_A1_N_c_397_n N_A2_N_c_476_n 0.0161016f $X=4.175 $Y=1.3 $X2=0 $Y2=0
cc_352 N_A1_N_c_392_n N_A_218_367#_M1002_g 0.00222399f $X=5.045 $Y=1.17 $X2=0
+ $Y2=0
cc_353 N_A1_N_c_393_n N_A_218_367#_M1002_g 0.00339141f $X=5.075 $Y=1.35 $X2=0
+ $Y2=0
cc_354 N_A1_N_c_396_n N_A_218_367#_M1002_g 0.00713592f $X=5.075 $Y=1.185 $X2=0
+ $Y2=0
cc_355 N_A1_N_M1000_g N_A_218_367#_c_584_n 0.0136307f $X=3.75 $Y=2.465 $X2=0
+ $Y2=0
cc_356 N_A1_N_M1022_g N_A_218_367#_c_584_n 0.0172496f $X=5.055 $Y=2.465 $X2=0
+ $Y2=0
cc_357 N_A1_N_M1022_g N_A_218_367#_c_531_n 0.0114386f $X=5.055 $Y=2.465 $X2=0
+ $Y2=0
cc_358 N_A1_N_M1022_g N_A_218_367#_c_532_n 7.27247e-19 $X=5.055 $Y=2.465 $X2=0
+ $Y2=0
cc_359 N_A1_N_c_392_n N_A_218_367#_c_532_n 0.009103f $X=5.045 $Y=1.17 $X2=0
+ $Y2=0
cc_360 N_A1_N_c_393_n N_A_218_367#_c_532_n 8.35889e-19 $X=5.075 $Y=1.35 $X2=0
+ $Y2=0
cc_361 N_A1_N_M1022_g N_A_218_367#_c_535_n 0.0465226f $X=5.055 $Y=2.465 $X2=0
+ $Y2=0
cc_362 N_A1_N_c_392_n N_A_218_367#_c_535_n 6.16624e-19 $X=5.045 $Y=1.17 $X2=0
+ $Y2=0
cc_363 N_A1_N_c_393_n N_A_218_367#_c_535_n 0.0105346f $X=5.075 $Y=1.35 $X2=0
+ $Y2=0
cc_364 N_A1_N_M1000_g N_VPWR_c_716_n 0.0013557f $X=3.75 $Y=2.465 $X2=0 $Y2=0
cc_365 N_A1_N_M1022_g N_VPWR_c_716_n 0.00132283f $X=5.055 $Y=2.465 $X2=0 $Y2=0
cc_366 N_A1_N_M1022_g N_VPWR_c_717_n 0.00972443f $X=5.055 $Y=2.465 $X2=0 $Y2=0
cc_367 N_A1_N_M1000_g N_VPWR_c_721_n 0.0036352f $X=3.75 $Y=2.465 $X2=0 $Y2=0
cc_368 N_A1_N_M1022_g N_VPWR_c_723_n 0.0036352f $X=5.055 $Y=2.465 $X2=0 $Y2=0
cc_369 N_A1_N_M1000_g N_VPWR_c_711_n 0.0043775f $X=3.75 $Y=2.465 $X2=0 $Y2=0
cc_370 N_A1_N_M1022_g N_VPWR_c_711_n 0.00439469f $X=5.055 $Y=2.465 $X2=0 $Y2=0
cc_371 N_A1_N_M1000_g N_VPWR_c_732_n 0.0107073f $X=3.75 $Y=2.465 $X2=0 $Y2=0
cc_372 N_A1_N_c_393_n N_X_c_852_n 2.40499e-19 $X=5.075 $Y=1.35 $X2=0 $Y2=0
cc_373 N_A1_N_c_395_n N_A_49_47#_c_937_n 0.00451107f $X=3.73 $Y=1.185 $X2=0
+ $Y2=0
cc_374 N_A1_N_c_395_n N_VGND_c_975_n 0.00459147f $X=3.73 $Y=1.185 $X2=0 $Y2=0
cc_375 N_A1_N_c_393_n N_VGND_c_976_n 0.00231617f $X=5.075 $Y=1.35 $X2=0 $Y2=0
cc_376 N_A1_N_c_396_n N_VGND_c_976_n 0.00356229f $X=5.075 $Y=1.185 $X2=0 $Y2=0
cc_377 N_A1_N_c_395_n N_VGND_c_983_n 0.00424523f $X=3.73 $Y=1.185 $X2=0 $Y2=0
cc_378 N_A1_N_c_396_n N_VGND_c_983_n 0.00547432f $X=5.075 $Y=1.185 $X2=0 $Y2=0
cc_379 N_A1_N_c_395_n N_VGND_c_991_n 0.00713961f $X=3.73 $Y=1.185 $X2=0 $Y2=0
cc_380 N_A1_N_c_396_n N_VGND_c_991_n 0.0103951f $X=5.075 $Y=1.185 $X2=0 $Y2=0
cc_381 N_A1_N_c_391_n N_A_768_47#_c_1094_n 0.00374916f $X=4.92 $Y=1.17 $X2=0
+ $Y2=0
cc_382 N_A1_N_c_395_n N_A_768_47#_c_1094_n 0.00304519f $X=3.73 $Y=1.185 $X2=0
+ $Y2=0
cc_383 N_A1_N_c_396_n N_A_768_47#_c_1099_n 0.00265698f $X=5.075 $Y=1.185 $X2=0
+ $Y2=0
cc_384 N_A1_N_c_391_n N_A_768_47#_c_1100_n 0.013862f $X=4.92 $Y=1.17 $X2=0 $Y2=0
cc_385 N_A1_N_c_392_n N_A_768_47#_c_1100_n 0.00458624f $X=5.045 $Y=1.17 $X2=0
+ $Y2=0
cc_386 N_A1_N_c_393_n N_A_768_47#_c_1100_n 2.81739e-19 $X=5.075 $Y=1.35 $X2=0
+ $Y2=0
cc_387 N_A1_N_c_396_n N_A_768_47#_c_1100_n 0.00490196f $X=5.075 $Y=1.185 $X2=0
+ $Y2=0
cc_388 N_A2_N_c_477_n N_A_218_367#_c_584_n 0.012347f $X=4.18 $Y=1.725 $X2=0
+ $Y2=0
cc_389 N_A2_N_c_478_n N_A_218_367#_c_584_n 0.0125211f $X=4.625 $Y=1.725 $X2=0
+ $Y2=0
cc_390 N_A2_N_c_475_n N_A_218_367#_c_531_n 0.0062038f $X=4.51 $Y=1.51 $X2=0
+ $Y2=0
cc_391 N_A2_N_c_475_n N_A_218_367#_c_532_n 0.00224029f $X=4.51 $Y=1.51 $X2=0
+ $Y2=0
cc_392 N_A2_N_c_477_n N_VPWR_c_716_n 0.00964774f $X=4.18 $Y=1.725 $X2=0 $Y2=0
cc_393 N_A2_N_c_478_n N_VPWR_c_716_n 0.00882798f $X=4.625 $Y=1.725 $X2=0 $Y2=0
cc_394 N_A2_N_c_478_n N_VPWR_c_717_n 0.00136612f $X=4.625 $Y=1.725 $X2=0 $Y2=0
cc_395 N_A2_N_c_477_n N_VPWR_c_721_n 0.0036352f $X=4.18 $Y=1.725 $X2=0 $Y2=0
cc_396 N_A2_N_c_478_n N_VPWR_c_723_n 0.00407237f $X=4.625 $Y=1.725 $X2=0 $Y2=0
cc_397 N_A2_N_c_477_n N_VPWR_c_711_n 0.00439469f $X=4.18 $Y=1.725 $X2=0 $Y2=0
cc_398 N_A2_N_c_478_n N_VPWR_c_711_n 0.00484671f $X=4.625 $Y=1.725 $X2=0 $Y2=0
cc_399 N_A2_N_c_477_n N_VPWR_c_732_n 0.00136669f $X=4.18 $Y=1.725 $X2=0 $Y2=0
cc_400 N_A2_N_c_473_n N_VGND_c_983_n 0.00357877f $X=4.195 $Y=1.185 $X2=0 $Y2=0
cc_401 N_A2_N_c_474_n N_VGND_c_983_n 0.00357877f $X=4.625 $Y=1.185 $X2=0 $Y2=0
cc_402 N_A2_N_c_473_n N_VGND_c_991_n 0.00537654f $X=4.195 $Y=1.185 $X2=0 $Y2=0
cc_403 N_A2_N_c_474_n N_VGND_c_991_n 0.00537654f $X=4.625 $Y=1.185 $X2=0 $Y2=0
cc_404 N_A2_N_c_473_n N_A_768_47#_c_1094_n 0.00961843f $X=4.195 $Y=1.185 $X2=0
+ $Y2=0
cc_405 N_A2_N_c_474_n N_A_768_47#_c_1094_n 0.0109843f $X=4.625 $Y=1.185 $X2=0
+ $Y2=0
cc_406 N_A_218_367#_c_584_n N_VPWR_M1019_s 0.0182777f $X=5.34 $Y=2.52 $X2=0
+ $Y2=0
cc_407 N_A_218_367#_c_584_n N_VPWR_M1012_d 0.00381036f $X=5.34 $Y=2.52 $X2=0
+ $Y2=0
cc_408 N_A_218_367#_c_584_n N_VPWR_M1022_d 0.00835531f $X=5.34 $Y=2.52 $X2=0
+ $Y2=0
cc_409 N_A_218_367#_c_531_n N_VPWR_M1022_d 0.00712828f $X=5.425 $Y=2.43 $X2=0
+ $Y2=0
cc_410 N_A_218_367#_c_530_n N_VPWR_c_715_n 0.00723383f $X=2.505 $Y=1.085 $X2=0
+ $Y2=0
cc_411 N_A_218_367#_c_541_n N_VPWR_c_715_n 0.0253916f $X=2.76 $Y=1.9 $X2=0 $Y2=0
cc_412 N_A_218_367#_c_584_n N_VPWR_c_716_n 0.0165322f $X=5.34 $Y=2.52 $X2=0
+ $Y2=0
cc_413 N_A_218_367#_M1010_g N_VPWR_c_717_n 0.00325225f $X=5.56 $Y=2.465 $X2=0
+ $Y2=0
cc_414 N_A_218_367#_c_584_n N_VPWR_c_717_n 0.0212369f $X=5.34 $Y=2.52 $X2=0
+ $Y2=0
cc_415 N_A_218_367#_M1010_g N_VPWR_c_718_n 7.57256e-19 $X=5.56 $Y=2.465 $X2=0
+ $Y2=0
cc_416 N_A_218_367#_M1018_g N_VPWR_c_718_n 0.0144481f $X=5.99 $Y=2.465 $X2=0
+ $Y2=0
cc_417 N_A_218_367#_M1023_g N_VPWR_c_718_n 0.0142791f $X=6.42 $Y=2.465 $X2=0
+ $Y2=0
cc_418 N_A_218_367#_M1027_g N_VPWR_c_718_n 7.27171e-19 $X=6.85 $Y=2.465 $X2=0
+ $Y2=0
cc_419 N_A_218_367#_M1023_g N_VPWR_c_719_n 0.00486043f $X=6.42 $Y=2.465 $X2=0
+ $Y2=0
cc_420 N_A_218_367#_M1027_g N_VPWR_c_719_n 0.00486043f $X=6.85 $Y=2.465 $X2=0
+ $Y2=0
cc_421 N_A_218_367#_M1023_g N_VPWR_c_720_n 7.42371e-19 $X=6.42 $Y=2.465 $X2=0
+ $Y2=0
cc_422 N_A_218_367#_M1027_g N_VPWR_c_720_n 0.015609f $X=6.85 $Y=2.465 $X2=0
+ $Y2=0
cc_423 N_A_218_367#_c_584_n N_VPWR_c_721_n 0.00670101f $X=5.34 $Y=2.52 $X2=0
+ $Y2=0
cc_424 N_A_218_367#_c_584_n N_VPWR_c_723_n 0.00690435f $X=5.34 $Y=2.52 $X2=0
+ $Y2=0
cc_425 N_A_218_367#_M1010_g N_VPWR_c_725_n 0.0056066f $X=5.56 $Y=2.465 $X2=0
+ $Y2=0
cc_426 N_A_218_367#_M1018_g N_VPWR_c_725_n 0.00486043f $X=5.99 $Y=2.465 $X2=0
+ $Y2=0
cc_427 N_A_218_367#_c_584_n N_VPWR_c_725_n 7.50781e-19 $X=5.34 $Y=2.52 $X2=0
+ $Y2=0
cc_428 N_A_218_367#_M1008_d N_VPWR_c_711_n 0.00231436f $X=1.09 $Y=1.835 $X2=0
+ $Y2=0
cc_429 N_A_218_367#_M1001_d N_VPWR_c_711_n 0.00243967f $X=2.625 $Y=1.835 $X2=0
+ $Y2=0
cc_430 N_A_218_367#_M1010_g N_VPWR_c_711_n 0.0101581f $X=5.56 $Y=2.465 $X2=0
+ $Y2=0
cc_431 N_A_218_367#_M1018_g N_VPWR_c_711_n 0.00824727f $X=5.99 $Y=2.465 $X2=0
+ $Y2=0
cc_432 N_A_218_367#_M1023_g N_VPWR_c_711_n 0.00824727f $X=6.42 $Y=2.465 $X2=0
+ $Y2=0
cc_433 N_A_218_367#_M1027_g N_VPWR_c_711_n 0.00824727f $X=6.85 $Y=2.465 $X2=0
+ $Y2=0
cc_434 N_A_218_367#_c_583_n N_VPWR_c_711_n 0.0101905f $X=2.765 $Y=2.91 $X2=0
+ $Y2=0
cc_435 N_A_218_367#_c_584_n N_VPWR_c_711_n 0.035681f $X=5.34 $Y=2.52 $X2=0 $Y2=0
cc_436 N_A_218_367#_c_598_n N_VPWR_c_711_n 0.00181391f $X=2.76 $Y=2.52 $X2=0
+ $Y2=0
cc_437 N_A_218_367#_c_583_n N_VPWR_c_731_n 0.0163698f $X=2.765 $Y=2.91 $X2=0
+ $Y2=0
cc_438 N_A_218_367#_c_584_n N_VPWR_c_731_n 0.00134205f $X=5.34 $Y=2.52 $X2=0
+ $Y2=0
cc_439 N_A_218_367#_c_598_n N_VPWR_c_731_n 7.19283e-19 $X=2.76 $Y=2.52 $X2=0
+ $Y2=0
cc_440 N_A_218_367#_c_584_n N_VPWR_c_732_n 0.0430389f $X=5.34 $Y=2.52 $X2=0
+ $Y2=0
cc_441 N_A_218_367#_c_546_n N_A_132_367#_M1021_s 0.0027969f $X=1.485 $Y=2.035
+ $X2=0 $Y2=0
cc_442 N_A_218_367#_c_529_n N_A_132_367#_M1021_s 7.96451e-19 $X=1.575 $Y=1.93
+ $X2=0 $Y2=0
cc_443 N_A_218_367#_M1008_d N_A_132_367#_c_839_n 0.00366227f $X=1.09 $Y=1.835
+ $X2=0 $Y2=0
cc_444 N_A_218_367#_M1018_g N_X_c_857_n 0.0133996f $X=5.99 $Y=2.465 $X2=0 $Y2=0
cc_445 N_A_218_367#_M1023_g N_X_c_857_n 0.0135857f $X=6.42 $Y=2.465 $X2=0 $Y2=0
cc_446 N_A_218_367#_c_656_p N_X_c_857_n 0.0469373f $X=7.01 $Y=1.49 $X2=0 $Y2=0
cc_447 N_A_218_367#_c_535_n N_X_c_857_n 0.00289796f $X=7.115 $Y=1.49 $X2=0 $Y2=0
cc_448 N_A_218_367#_M1010_g N_X_c_858_n 7.38449e-19 $X=5.56 $Y=2.465 $X2=0 $Y2=0
cc_449 N_A_218_367#_c_531_n N_X_c_858_n 0.0102784f $X=5.425 $Y=2.43 $X2=0 $Y2=0
cc_450 N_A_218_367#_c_656_p N_X_c_858_n 0.0153308f $X=7.01 $Y=1.49 $X2=0 $Y2=0
cc_451 N_A_218_367#_c_535_n N_X_c_858_n 0.0028903f $X=7.115 $Y=1.49 $X2=0 $Y2=0
cc_452 N_A_218_367#_M1002_g N_X_c_872_n 0.0137938f $X=5.825 $Y=0.655 $X2=0 $Y2=0
cc_453 N_A_218_367#_M1005_g N_X_c_851_n 0.0147781f $X=6.255 $Y=0.655 $X2=0 $Y2=0
cc_454 N_A_218_367#_M1013_g N_X_c_851_n 0.0147781f $X=6.685 $Y=0.655 $X2=0 $Y2=0
cc_455 N_A_218_367#_c_656_p N_X_c_851_n 0.0471383f $X=7.01 $Y=1.49 $X2=0 $Y2=0
cc_456 N_A_218_367#_c_535_n N_X_c_851_n 0.00290124f $X=7.115 $Y=1.49 $X2=0 $Y2=0
cc_457 N_A_218_367#_M1002_g N_X_c_852_n 0.0100433f $X=5.825 $Y=0.655 $X2=0 $Y2=0
cc_458 N_A_218_367#_c_656_p N_X_c_852_n 0.0208668f $X=7.01 $Y=1.49 $X2=0 $Y2=0
cc_459 N_A_218_367#_c_535_n N_X_c_852_n 0.00299787f $X=7.115 $Y=1.49 $X2=0 $Y2=0
cc_460 N_A_218_367#_M1027_g N_X_c_859_n 0.0157201f $X=6.85 $Y=2.465 $X2=0 $Y2=0
cc_461 N_A_218_367#_c_656_p N_X_c_859_n 0.0320881f $X=7.01 $Y=1.49 $X2=0 $Y2=0
cc_462 N_A_218_367#_c_535_n N_X_c_859_n 0.00763465f $X=7.115 $Y=1.49 $X2=0 $Y2=0
cc_463 N_A_218_367#_M1017_g N_X_c_853_n 0.0167079f $X=7.115 $Y=0.655 $X2=0 $Y2=0
cc_464 N_A_218_367#_c_656_p N_X_c_853_n 0.0124393f $X=7.01 $Y=1.49 $X2=0 $Y2=0
cc_465 N_A_218_367#_c_656_p N_X_c_860_n 0.0145237f $X=7.01 $Y=1.49 $X2=0 $Y2=0
cc_466 N_A_218_367#_c_535_n N_X_c_860_n 0.00299787f $X=7.115 $Y=1.49 $X2=0 $Y2=0
cc_467 N_A_218_367#_c_656_p N_X_c_854_n 0.0153308f $X=7.01 $Y=1.49 $X2=0 $Y2=0
cc_468 N_A_218_367#_c_535_n N_X_c_854_n 0.0028903f $X=7.115 $Y=1.49 $X2=0 $Y2=0
cc_469 N_A_218_367#_M1027_g X 0.00244976f $X=6.85 $Y=2.465 $X2=0 $Y2=0
cc_470 N_A_218_367#_M1017_g X 0.0148812f $X=7.115 $Y=0.655 $X2=0 $Y2=0
cc_471 N_A_218_367#_c_656_p X 0.0138085f $X=7.01 $Y=1.49 $X2=0 $Y2=0
cc_472 N_A_218_367#_c_530_n N_A_49_47#_M1009_d 0.00176773f $X=2.505 $Y=1.085
+ $X2=0 $Y2=0
cc_473 N_A_218_367#_c_529_n N_A_49_47#_c_915_n 0.00482399f $X=1.575 $Y=1.93
+ $X2=0 $Y2=0
cc_474 N_A_218_367#_c_573_n N_A_49_47#_c_915_n 0.00929066f $X=1.665 $Y=1.085
+ $X2=0 $Y2=0
cc_475 N_A_218_367#_c_530_n N_A_49_47#_c_922_n 0.0370161f $X=2.505 $Y=1.085
+ $X2=0 $Y2=0
cc_476 N_A_218_367#_c_573_n N_A_49_47#_c_922_n 0.00982569f $X=1.665 $Y=1.085
+ $X2=0 $Y2=0
cc_477 N_A_218_367#_M1003_s N_A_49_47#_c_935_n 0.00332931f $X=2.46 $Y=0.235
+ $X2=0 $Y2=0
cc_478 N_A_218_367#_c_530_n N_A_49_47#_c_935_n 0.00319453f $X=2.505 $Y=1.085
+ $X2=0 $Y2=0
cc_479 N_A_218_367#_c_575_n N_A_49_47#_c_935_n 0.0139642f $X=2.6 $Y=0.77 $X2=0
+ $Y2=0
cc_480 N_A_218_367#_c_530_n N_VGND_M1024_s 0.00167596f $X=2.505 $Y=1.085 $X2=0
+ $Y2=0
cc_481 N_A_218_367#_c_573_n N_VGND_M1024_s 9.76226e-19 $X=1.665 $Y=1.085 $X2=0
+ $Y2=0
cc_482 N_A_218_367#_M1002_g N_VGND_c_976_n 0.00202686f $X=5.825 $Y=0.655 $X2=0
+ $Y2=0
cc_483 N_A_218_367#_c_532_n N_VGND_c_976_n 0.00717404f $X=5.51 $Y=1.49 $X2=0
+ $Y2=0
cc_484 N_A_218_367#_c_656_p N_VGND_c_976_n 0.0065067f $X=7.01 $Y=1.49 $X2=0
+ $Y2=0
cc_485 N_A_218_367#_c_535_n N_VGND_c_976_n 0.00515928f $X=7.115 $Y=1.49 $X2=0
+ $Y2=0
cc_486 N_A_218_367#_M1002_g N_VGND_c_977_n 7.07939e-19 $X=5.825 $Y=0.655 $X2=0
+ $Y2=0
cc_487 N_A_218_367#_M1005_g N_VGND_c_977_n 0.0110403f $X=6.255 $Y=0.655 $X2=0
+ $Y2=0
cc_488 N_A_218_367#_M1013_g N_VGND_c_977_n 0.0108821f $X=6.685 $Y=0.655 $X2=0
+ $Y2=0
cc_489 N_A_218_367#_M1017_g N_VGND_c_977_n 6.25324e-19 $X=7.115 $Y=0.655 $X2=0
+ $Y2=0
cc_490 N_A_218_367#_M1013_g N_VGND_c_979_n 6.25324e-19 $X=6.685 $Y=0.655 $X2=0
+ $Y2=0
cc_491 N_A_218_367#_M1017_g N_VGND_c_979_n 0.0117461f $X=7.115 $Y=0.655 $X2=0
+ $Y2=0
cc_492 N_A_218_367#_M1002_g N_VGND_c_984_n 0.0054895f $X=5.825 $Y=0.655 $X2=0
+ $Y2=0
cc_493 N_A_218_367#_M1005_g N_VGND_c_984_n 0.00486043f $X=6.255 $Y=0.655 $X2=0
+ $Y2=0
cc_494 N_A_218_367#_M1013_g N_VGND_c_985_n 0.00486043f $X=6.685 $Y=0.655 $X2=0
+ $Y2=0
cc_495 N_A_218_367#_M1017_g N_VGND_c_985_n 0.00486043f $X=7.115 $Y=0.655 $X2=0
+ $Y2=0
cc_496 N_A_218_367#_M1003_s N_VGND_c_991_n 0.00225186f $X=2.46 $Y=0.235 $X2=0
+ $Y2=0
cc_497 N_A_218_367#_M1002_g N_VGND_c_991_n 0.0104069f $X=5.825 $Y=0.655 $X2=0
+ $Y2=0
cc_498 N_A_218_367#_M1005_g N_VGND_c_991_n 0.00824727f $X=6.255 $Y=0.655 $X2=0
+ $Y2=0
cc_499 N_A_218_367#_M1013_g N_VGND_c_991_n 0.00824727f $X=6.685 $Y=0.655 $X2=0
+ $Y2=0
cc_500 N_A_218_367#_M1017_g N_VGND_c_991_n 0.00824727f $X=7.115 $Y=0.655 $X2=0
+ $Y2=0
cc_501 N_VPWR_c_711_n N_A_132_367#_M1011_s 0.00231436f $X=7.44 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_502 N_VPWR_c_711_n N_A_132_367#_M1021_s 0.00253344f $X=7.44 $Y=3.33 $X2=0
+ $Y2=0
cc_503 N_VPWR_c_727_n N_A_132_367#_c_839_n 0.0442127f $X=1.935 $Y=3.33 $X2=0
+ $Y2=0
cc_504 N_VPWR_c_711_n N_A_132_367#_c_839_n 0.0399976f $X=7.44 $Y=3.33 $X2=0
+ $Y2=0
cc_505 N_VPWR_c_711_n N_X_M1010_d 0.00536646f $X=7.44 $Y=3.33 $X2=0 $Y2=0
cc_506 N_VPWR_c_711_n N_X_M1023_d 0.00571434f $X=7.44 $Y=3.33 $X2=0 $Y2=0
cc_507 N_VPWR_c_725_n N_X_c_894_n 0.0124525f $X=6.04 $Y=3.33 $X2=0 $Y2=0
cc_508 N_VPWR_c_711_n N_X_c_894_n 0.00730901f $X=7.44 $Y=3.33 $X2=0 $Y2=0
cc_509 N_VPWR_M1018_s N_X_c_857_n 0.00176773f $X=6.065 $Y=1.835 $X2=0 $Y2=0
cc_510 N_VPWR_c_718_n N_X_c_857_n 0.0171443f $X=6.205 $Y=2.18 $X2=0 $Y2=0
cc_511 N_VPWR_c_719_n N_X_c_898_n 0.0120977f $X=6.9 $Y=3.33 $X2=0 $Y2=0
cc_512 N_VPWR_c_711_n N_X_c_898_n 0.00691495f $X=7.44 $Y=3.33 $X2=0 $Y2=0
cc_513 N_VPWR_M1027_s N_X_c_859_n 0.00263371f $X=6.925 $Y=1.835 $X2=0 $Y2=0
cc_514 N_VPWR_c_720_n N_X_c_859_n 0.022088f $X=7.065 $Y=2.18 $X2=0 $Y2=0
cc_515 N_VPWR_c_713_n N_A_49_47#_c_916_n 0.00492604f $X=0.37 $Y=1.98 $X2=0 $Y2=0
cc_516 N_X_c_851_n N_VGND_M1005_d 0.00177068f $X=6.805 $Y=1.14 $X2=0 $Y2=0
cc_517 N_X_c_853_n N_VGND_M1017_d 0.00103467f $X=7.345 $Y=1.14 $X2=0 $Y2=0
cc_518 N_X_c_855_n N_VGND_M1017_d 0.00135843f $X=7.47 $Y=1.235 $X2=0 $Y2=0
cc_519 N_X_c_851_n N_VGND_c_977_n 0.0172078f $X=6.805 $Y=1.14 $X2=0 $Y2=0
cc_520 N_X_c_853_n N_VGND_c_979_n 0.00979637f $X=7.345 $Y=1.14 $X2=0 $Y2=0
cc_521 N_X_c_855_n N_VGND_c_979_n 0.013572f $X=7.47 $Y=1.235 $X2=0 $Y2=0
cc_522 N_X_c_872_n N_VGND_c_984_n 0.015688f $X=6.04 $Y=0.42 $X2=0 $Y2=0
cc_523 N_X_c_909_p N_VGND_c_985_n 0.0124525f $X=6.9 $Y=0.42 $X2=0 $Y2=0
cc_524 N_X_M1002_s N_VGND_c_991_n 0.00380103f $X=5.9 $Y=0.235 $X2=0 $Y2=0
cc_525 N_X_M1013_s N_VGND_c_991_n 0.00536646f $X=6.76 $Y=0.235 $X2=0 $Y2=0
cc_526 N_X_c_872_n N_VGND_c_991_n 0.00984745f $X=6.04 $Y=0.42 $X2=0 $Y2=0
cc_527 N_X_c_909_p N_VGND_c_991_n 0.00730901f $X=6.9 $Y=0.42 $X2=0 $Y2=0
cc_528 N_A_49_47#_c_915_n N_VGND_M1006_s 0.00176461f $X=1.135 $Y=1.15 $X2=-0.19
+ $Y2=-0.245
cc_529 N_A_49_47#_c_922_n N_VGND_M1024_s 0.00507645f $X=2.005 $Y=0.74 $X2=0
+ $Y2=0
cc_530 N_A_49_47#_c_915_n N_VGND_c_973_n 0.0170777f $X=1.135 $Y=1.15 $X2=0 $Y2=0
cc_531 N_A_49_47#_c_922_n N_VGND_c_974_n 0.0205525f $X=2.005 $Y=0.74 $X2=0 $Y2=0
cc_532 N_A_49_47#_c_937_n N_VGND_c_975_n 0.0181025f $X=3.03 $Y=0.42 $X2=0 $Y2=0
cc_533 N_A_49_47#_c_914_n N_VGND_c_980_n 0.0178111f $X=0.37 $Y=0.42 $X2=0 $Y2=0
cc_534 N_A_49_47#_c_957_p N_VGND_c_981_n 0.0124525f $X=1.23 $Y=0.42 $X2=0 $Y2=0
cc_535 N_A_49_47#_c_922_n N_VGND_c_981_n 0.00235807f $X=2.005 $Y=0.74 $X2=0
+ $Y2=0
cc_536 N_A_49_47#_c_922_n N_VGND_c_982_n 0.00244463f $X=2.005 $Y=0.74 $X2=0
+ $Y2=0
cc_537 N_A_49_47#_c_923_n N_VGND_c_982_n 0.018869f $X=2.17 $Y=0.435 $X2=0 $Y2=0
cc_538 N_A_49_47#_c_935_n N_VGND_c_982_n 0.0329194f $X=2.93 $Y=0.345 $X2=0 $Y2=0
cc_539 N_A_49_47#_c_937_n N_VGND_c_982_n 0.0131188f $X=3.03 $Y=0.42 $X2=0 $Y2=0
cc_540 N_A_49_47#_M1006_d N_VGND_c_991_n 0.00371702f $X=0.245 $Y=0.235 $X2=0
+ $Y2=0
cc_541 N_A_49_47#_M1014_d N_VGND_c_991_n 0.00396356f $X=1.09 $Y=0.235 $X2=0
+ $Y2=0
cc_542 N_A_49_47#_M1009_d N_VGND_c_991_n 0.00223559f $X=2.03 $Y=0.235 $X2=0
+ $Y2=0
cc_543 N_A_49_47#_M1015_d N_VGND_c_991_n 0.00319523f $X=2.89 $Y=0.235 $X2=0
+ $Y2=0
cc_544 N_A_49_47#_c_914_n N_VGND_c_991_n 0.0100304f $X=0.37 $Y=0.42 $X2=0 $Y2=0
cc_545 N_A_49_47#_c_957_p N_VGND_c_991_n 0.0073074f $X=1.23 $Y=0.42 $X2=0 $Y2=0
cc_546 N_A_49_47#_c_922_n N_VGND_c_991_n 0.00998089f $X=2.005 $Y=0.74 $X2=0
+ $Y2=0
cc_547 N_A_49_47#_c_923_n N_VGND_c_991_n 0.0123965f $X=2.17 $Y=0.435 $X2=0 $Y2=0
cc_548 N_A_49_47#_c_935_n N_VGND_c_991_n 0.0210677f $X=2.93 $Y=0.345 $X2=0 $Y2=0
cc_549 N_A_49_47#_c_937_n N_VGND_c_991_n 0.00758115f $X=3.03 $Y=0.42 $X2=0 $Y2=0
cc_550 N_VGND_c_991_n N_A_768_47#_M1004_s 0.00223577f $X=7.44 $Y=0 $X2=-0.19
+ $Y2=-0.245
cc_551 N_VGND_c_991_n N_A_768_47#_M1025_s 0.00223562f $X=7.44 $Y=0 $X2=0 $Y2=0
cc_552 N_VGND_c_983_n N_A_768_47#_c_1094_n 0.0514187f $X=5.175 $Y=0 $X2=0 $Y2=0
cc_553 N_VGND_c_991_n N_A_768_47#_c_1094_n 0.0334963f $X=7.44 $Y=0 $X2=0 $Y2=0
cc_554 N_VGND_c_983_n N_A_768_47#_c_1099_n 0.0157627f $X=5.175 $Y=0 $X2=0 $Y2=0
cc_555 N_VGND_c_991_n N_A_768_47#_c_1099_n 0.00991281f $X=7.44 $Y=0 $X2=0 $Y2=0
