* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__buf_8 A VGND VNB VPB VPWR X
M1000 VPWR A a_27_47# VPB phighvt w=1.26e+06u l=150000u
+  ad=2.1231e+12p pd=1.849e+07u as=6.867e+11p ps=6.13e+06u
M1001 X a_27_47# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=1.4112e+12p pd=1.232e+07u as=0p ps=0u
M1002 VGND a_27_47# X VNB nshort w=840000u l=150000u
+  ad=1.4154e+12p pd=1.345e+07u as=9.408e+11p ps=8.96e+06u
M1003 VPWR a_27_47# X VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 X a_27_47# VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VPWR a_27_47# X VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND A a_27_47# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=4.578e+11p ps=4.45e+06u
M1007 a_27_47# A VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPWR a_27_47# X VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND a_27_47# X VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND a_27_47# X VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 X a_27_47# VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_27_47# A VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VPWR a_27_47# X VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 X a_27_47# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 X a_27_47# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 X a_27_47# VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 X a_27_47# VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 X a_27_47# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VGND a_27_47# X VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VPWR A a_27_47# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VGND A a_27_47# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
