* File: sky130_fd_sc_lp__a32oi_2.pxi.spice
* Created: Wed Sep  2 09:28:21 2020
* 
x_PM_SKY130_FD_SC_LP__A32OI_2%B2 N_B2_c_91_n N_B2_M1012_g N_B2_M1005_g
+ N_B2_c_93_n N_B2_M1013_g N_B2_M1011_g N_B2_c_95_n B2 B2 N_B2_c_97_n
+ PM_SKY130_FD_SC_LP__A32OI_2%B2
x_PM_SKY130_FD_SC_LP__A32OI_2%B1 N_B1_M1003_g N_B1_M1000_g N_B1_M1009_g
+ N_B1_M1008_g N_B1_c_142_n B1 N_B1_c_143_n N_B1_c_144_n N_B1_c_145_n
+ PM_SKY130_FD_SC_LP__A32OI_2%B1
x_PM_SKY130_FD_SC_LP__A32OI_2%A1 N_A1_M1016_g N_A1_M1007_g N_A1_M1015_g
+ N_A1_M1019_g A1 N_A1_c_200_n N_A1_c_197_n PM_SKY130_FD_SC_LP__A32OI_2%A1
x_PM_SKY130_FD_SC_LP__A32OI_2%A2 N_A2_M1004_g N_A2_M1002_g N_A2_M1010_g
+ N_A2_M1018_g A2 A2 A2 N_A2_c_252_n PM_SKY130_FD_SC_LP__A32OI_2%A2
x_PM_SKY130_FD_SC_LP__A32OI_2%A3 N_A3_M1001_g N_A3_c_300_n N_A3_M1006_g
+ N_A3_M1014_g N_A3_c_302_n N_A3_M1017_g A3 N_A3_c_304_n
+ PM_SKY130_FD_SC_LP__A32OI_2%A3
x_PM_SKY130_FD_SC_LP__A32OI_2%A_43_367# N_A_43_367#_M1005_s N_A_43_367#_M1011_s
+ N_A_43_367#_M1008_d N_A_43_367#_M1019_d N_A_43_367#_M1018_d
+ N_A_43_367#_M1014_d N_A_43_367#_c_337_n N_A_43_367#_c_338_n
+ N_A_43_367#_c_344_n N_A_43_367#_c_369_p N_A_43_367#_c_346_n
+ N_A_43_367#_c_348_n N_A_43_367#_c_349_n N_A_43_367#_c_352_n
+ N_A_43_367#_c_383_p N_A_43_367#_c_355_n N_A_43_367#_c_356_n
+ N_A_43_367#_c_339_n N_A_43_367#_c_382_p N_A_43_367#_c_340_n
+ N_A_43_367#_c_341_n N_A_43_367#_c_397_p PM_SKY130_FD_SC_LP__A32OI_2%A_43_367#
x_PM_SKY130_FD_SC_LP__A32OI_2%Y N_Y_M1003_d N_Y_M1007_d N_Y_M1005_d N_Y_M1000_s
+ N_Y_c_414_n N_Y_c_410_n N_Y_c_411_n N_Y_c_427_n N_Y_c_412_n N_Y_c_433_n
+ N_Y_c_408_n N_Y_c_409_n N_Y_c_441_n Y Y Y Y N_Y_c_453_n N_Y_c_455_n Y
+ PM_SKY130_FD_SC_LP__A32OI_2%Y
x_PM_SKY130_FD_SC_LP__A32OI_2%VPWR N_VPWR_M1016_s N_VPWR_M1002_s N_VPWR_M1001_s
+ N_VPWR_c_496_n N_VPWR_c_497_n N_VPWR_c_498_n N_VPWR_c_499_n VPWR
+ N_VPWR_c_500_n N_VPWR_c_501_n N_VPWR_c_495_n N_VPWR_c_503_n N_VPWR_c_504_n
+ N_VPWR_c_505_n PM_SKY130_FD_SC_LP__A32OI_2%VPWR
x_PM_SKY130_FD_SC_LP__A32OI_2%A_43_65# N_A_43_65#_M1012_s N_A_43_65#_M1013_s
+ N_A_43_65#_M1009_s N_A_43_65#_c_570_n N_A_43_65#_c_576_n N_A_43_65#_c_571_n
+ N_A_43_65#_c_572_n N_A_43_65#_c_573_n N_A_43_65#_c_574_n
+ PM_SKY130_FD_SC_LP__A32OI_2%A_43_65#
x_PM_SKY130_FD_SC_LP__A32OI_2%VGND N_VGND_M1012_d N_VGND_M1006_d N_VGND_M1017_d
+ N_VGND_c_605_n N_VGND_c_606_n N_VGND_c_607_n N_VGND_c_608_n VGND
+ N_VGND_c_609_n N_VGND_c_610_n N_VGND_c_611_n N_VGND_c_612_n N_VGND_c_613_n
+ N_VGND_c_614_n PM_SKY130_FD_SC_LP__A32OI_2%VGND
x_PM_SKY130_FD_SC_LP__A32OI_2%A_509_65# N_A_509_65#_M1007_s N_A_509_65#_M1015_s
+ N_A_509_65#_M1010_s N_A_509_65#_c_671_n N_A_509_65#_c_672_n
+ N_A_509_65#_c_673_n N_A_509_65#_c_674_n N_A_509_65#_c_675_n
+ N_A_509_65#_c_676_n N_A_509_65#_c_677_n PM_SKY130_FD_SC_LP__A32OI_2%A_509_65#
x_PM_SKY130_FD_SC_LP__A32OI_2%A_778_65# N_A_778_65#_M1004_d N_A_778_65#_M1006_s
+ N_A_778_65#_c_713_n N_A_778_65#_c_711_n N_A_778_65#_c_712_n
+ N_A_778_65#_c_733_n PM_SKY130_FD_SC_LP__A32OI_2%A_778_65#
cc_1 VNB N_B2_c_91_n 0.021507f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=1.275
cc_2 VNB N_B2_M1005_g 0.0026762f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=2.465
cc_3 VNB N_B2_c_93_n 0.0166401f $X=-0.19 $Y=-0.245 $X2=0.985 $Y2=1.275
cc_4 VNB N_B2_M1011_g 0.002573f $X=-0.19 $Y=-0.245 $X2=0.985 $Y2=2.465
cc_5 VNB N_B2_c_95_n 0.003077f $X=-0.19 $Y=-0.245 $X2=0.895 $Y2=1.44
cc_6 VNB B2 0.0244591f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_7 VNB N_B2_c_97_n 0.0630706f $X=-0.19 $Y=-0.245 $X2=0.985 $Y2=1.44
cc_8 VNB N_B1_M1003_g 0.0198589f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=0.745
cc_9 VNB N_B1_M1000_g 0.0083402f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_B1_M1009_g 0.0258596f $X=-0.19 $Y=-0.245 $X2=0.985 $Y2=2.465
cc_11 VNB N_B1_c_142_n 0.00536961f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_B1_c_143_n 0.00884974f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_B1_c_144_n 0.0285979f $X=-0.19 $Y=-0.245 $X2=0.4 $Y2=1.44
cc_14 VNB N_B1_c_145_n 0.0017692f $X=-0.19 $Y=-0.245 $X2=0.4 $Y2=1.44
cc_15 VNB N_A1_M1007_g 0.0254324f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A1_M1015_g 0.0194466f $X=-0.19 $Y=-0.245 $X2=0.985 $Y2=1.605
cc_17 VNB N_A1_c_197_n 0.0588454f $X=-0.19 $Y=-0.245 $X2=0.4 $Y2=1.44
cc_18 VNB N_A2_M1004_g 0.0198658f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=0.745
cc_19 VNB N_A2_M1010_g 0.0254946f $X=-0.19 $Y=-0.245 $X2=0.985 $Y2=1.605
cc_20 VNB A2 0.00529114f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A2_c_252_n 0.05824f $X=-0.19 $Y=-0.245 $X2=0.985 $Y2=1.44
cc_22 VNB N_A3_M1001_g 0.00676868f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=0.745
cc_23 VNB N_A3_c_300_n 0.0186908f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=2.465
cc_24 VNB N_A3_M1014_g 0.0103812f $X=-0.19 $Y=-0.245 $X2=0.985 $Y2=0.745
cc_25 VNB N_A3_c_302_n 0.0211802f $X=-0.19 $Y=-0.245 $X2=0.985 $Y2=2.465
cc_26 VNB A3 0.021492f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=1.4
cc_27 VNB N_A3_c_304_n 0.0802101f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_Y_c_408_n 0.0184568f $X=-0.19 $Y=-0.245 $X2=0.895 $Y2=1.44
cc_29 VNB N_Y_c_409_n 0.00297453f $X=-0.19 $Y=-0.245 $X2=0.985 $Y2=1.44
cc_30 VNB N_VPWR_c_495_n 0.263193f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_43_65#_c_570_n 0.0230663f $X=-0.19 $Y=-0.245 $X2=0.985 $Y2=2.465
cc_32 VNB N_A_43_65#_c_571_n 0.00755006f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=1.4
cc_33 VNB N_A_43_65#_c_572_n 0.00705819f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_34 VNB N_A_43_65#_c_573_n 0.00185825f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_35 VNB N_A_43_65#_c_574_n 0.00482896f $X=-0.19 $Y=-0.245 $X2=0.4 $Y2=1.44
cc_36 VNB N_VGND_c_605_n 0.00280617f $X=-0.19 $Y=-0.245 $X2=0.985 $Y2=2.465
cc_37 VNB N_VGND_c_606_n 0.00966991f $X=-0.19 $Y=-0.245 $X2=0.895 $Y2=1.4
cc_38 VNB N_VGND_c_607_n 0.0123554f $X=-0.19 $Y=-0.245 $X2=0.895 $Y2=1.44
cc_39 VNB N_VGND_c_608_n 0.0335597f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_40 VNB N_VGND_c_609_n 0.0187828f $X=-0.19 $Y=-0.245 $X2=0.4 $Y2=1.44
cc_41 VNB N_VGND_c_610_n 0.0943507f $X=-0.19 $Y=-0.245 $X2=0.895 $Y2=1.44
cc_42 VNB N_VGND_c_611_n 0.0130715f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_612_n 0.00549308f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_613_n 0.00521013f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_614_n 0.353991f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_509_65#_c_671_n 0.00473978f $X=-0.19 $Y=-0.245 $X2=0.985 $Y2=2.465
cc_47 VNB N_A_509_65#_c_672_n 0.00266623f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_509_65#_c_673_n 0.00439196f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=1.4
cc_49 VNB N_A_509_65#_c_674_n 0.00291322f $X=-0.19 $Y=-0.245 $X2=0.895 $Y2=1.44
cc_50 VNB N_A_509_65#_c_675_n 0.00700408f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_51 VNB N_A_509_65#_c_676_n 0.00454207f $X=-0.19 $Y=-0.245 $X2=0.4 $Y2=1.44
cc_52 VNB N_A_509_65#_c_677_n 0.00140772f $X=-0.19 $Y=-0.245 $X2=0.4 $Y2=1.44
cc_53 VNB N_A_778_65#_c_711_n 0.0179344f $X=-0.19 $Y=-0.245 $X2=0.985 $Y2=1.605
cc_54 VNB N_A_778_65#_c_712_n 0.0023296f $X=-0.19 $Y=-0.245 $X2=0.985 $Y2=2.465
cc_55 VPB N_B2_M1005_g 0.0244786f $X=-0.19 $Y=1.655 $X2=0.555 $Y2=2.465
cc_56 VPB N_B2_M1011_g 0.0187382f $X=-0.19 $Y=1.655 $X2=0.985 $Y2=2.465
cc_57 VPB B2 0.0107404f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_58 VPB N_B1_M1000_g 0.0187371f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_59 VPB N_B1_M1008_g 0.020766f $X=-0.19 $Y=1.655 $X2=0.895 $Y2=1.44
cc_60 VPB N_B1_c_144_n 0.010238f $X=-0.19 $Y=1.655 $X2=0.4 $Y2=1.44
cc_61 VPB N_B1_c_145_n 0.00376825f $X=-0.19 $Y=1.655 $X2=0.4 $Y2=1.44
cc_62 VPB N_A1_M1016_g 0.0246263f $X=-0.19 $Y=1.655 $X2=0.555 $Y2=0.745
cc_63 VPB N_A1_M1019_g 0.0234311f $X=-0.19 $Y=1.655 $X2=0.485 $Y2=1.4
cc_64 VPB N_A1_c_200_n 0.00228291f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_65 VPB N_A1_c_197_n 0.0179389f $X=-0.19 $Y=1.655 $X2=0.4 $Y2=1.44
cc_66 VPB N_A2_M1002_g 0.0220019f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_67 VPB N_A2_M1018_g 0.0215554f $X=-0.19 $Y=1.655 $X2=0.485 $Y2=1.4
cc_68 VPB A2 0.00958948f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_69 VPB N_A2_c_252_n 0.0185612f $X=-0.19 $Y=1.655 $X2=0.985 $Y2=1.44
cc_70 VPB N_A3_M1001_g 0.0191364f $X=-0.19 $Y=1.655 $X2=0.555 $Y2=0.745
cc_71 VPB N_A3_M1014_g 0.0257505f $X=-0.19 $Y=1.655 $X2=0.985 $Y2=0.745
cc_72 VPB N_A_43_367#_c_337_n 0.00746637f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_73 VPB N_A_43_367#_c_338_n 0.0370247f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_74 VPB N_A_43_367#_c_339_n 0.003563f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_75 VPB N_A_43_367#_c_340_n 0.0142718f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_76 VPB N_A_43_367#_c_341_n 0.0435297f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_77 VPB N_Y_c_410_n 0.00544527f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_78 VPB N_Y_c_411_n 0.00228659f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_79 VPB N_Y_c_412_n 0.00362291f $X=-0.19 $Y=1.655 $X2=0.4 $Y2=1.44
cc_80 VPB Y 0.00168346f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_81 VPB N_VPWR_c_496_n 0.00192049f $X=-0.19 $Y=1.655 $X2=0.985 $Y2=2.465
cc_82 VPB N_VPWR_c_497_n 3.99129e-19 $X=-0.19 $Y=1.655 $X2=0.895 $Y2=1.4
cc_83 VPB N_VPWR_c_498_n 0.0129398f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_84 VPB N_VPWR_c_499_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_85 VPB N_VPWR_c_500_n 0.0147271f $X=-0.19 $Y=1.655 $X2=0.985 $Y2=1.44
cc_86 VPB N_VPWR_c_501_n 0.0220585f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_87 VPB N_VPWR_c_495_n 0.0573441f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_88 VPB N_VPWR_c_503_n 0.0616335f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_89 VPB N_VPWR_c_504_n 0.0149125f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_90 VPB N_VPWR_c_505_n 0.0110121f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_91 N_B2_c_93_n N_B1_M1003_g 0.0186907f $X=0.985 $Y=1.275 $X2=0 $Y2=0
cc_92 N_B2_c_95_n N_B1_M1003_g 0.00171011f $X=0.895 $Y=1.44 $X2=0 $Y2=0
cc_93 N_B2_M1011_g N_B1_M1000_g 0.0186907f $X=0.985 $Y=2.465 $X2=0 $Y2=0
cc_94 N_B2_c_97_n N_B1_c_142_n 0.0186907f $X=0.985 $Y=1.44 $X2=0 $Y2=0
cc_95 B2 N_A_43_367#_c_338_n 0.0229113f $X=0.155 $Y=1.58 $X2=0 $Y2=0
cc_96 N_B2_c_97_n N_A_43_367#_c_338_n 0.00106234f $X=0.985 $Y=1.44 $X2=0 $Y2=0
cc_97 N_B2_M1005_g N_A_43_367#_c_344_n 0.0115031f $X=0.555 $Y=2.465 $X2=0 $Y2=0
cc_98 N_B2_M1011_g N_A_43_367#_c_344_n 0.0115031f $X=0.985 $Y=2.465 $X2=0 $Y2=0
cc_99 N_B2_M1005_g N_Y_c_414_n 0.0116775f $X=0.555 $Y=2.465 $X2=0 $Y2=0
cc_100 N_B2_M1011_g N_Y_c_414_n 0.0103476f $X=0.985 $Y=2.465 $X2=0 $Y2=0
cc_101 N_B2_M1011_g N_Y_c_410_n 0.0111034f $X=0.985 $Y=2.465 $X2=0 $Y2=0
cc_102 N_B2_c_95_n N_Y_c_410_n 0.00869731f $X=0.895 $Y=1.44 $X2=0 $Y2=0
cc_103 N_B2_M1005_g N_Y_c_411_n 0.00767224f $X=0.555 $Y=2.465 $X2=0 $Y2=0
cc_104 N_B2_M1011_g N_Y_c_411_n 0.00241999f $X=0.985 $Y=2.465 $X2=0 $Y2=0
cc_105 N_B2_c_95_n N_Y_c_411_n 0.027089f $X=0.895 $Y=1.44 $X2=0 $Y2=0
cc_106 B2 N_Y_c_411_n 0.005505f $X=0.155 $Y=1.58 $X2=0 $Y2=0
cc_107 N_B2_c_97_n N_Y_c_411_n 0.00256759f $X=0.985 $Y=1.44 $X2=0 $Y2=0
cc_108 N_B2_M1011_g N_Y_c_412_n 4.58312e-19 $X=0.985 $Y=2.465 $X2=0 $Y2=0
cc_109 N_B2_c_93_n N_Y_c_409_n 8.21499e-19 $X=0.985 $Y=1.275 $X2=0 $Y2=0
cc_110 N_B2_M1005_g N_VPWR_c_495_n 0.00635116f $X=0.555 $Y=2.465 $X2=0 $Y2=0
cc_111 N_B2_M1011_g N_VPWR_c_495_n 0.00537654f $X=0.985 $Y=2.465 $X2=0 $Y2=0
cc_112 N_B2_M1005_g N_VPWR_c_503_n 0.00357877f $X=0.555 $Y=2.465 $X2=0 $Y2=0
cc_113 N_B2_M1011_g N_VPWR_c_503_n 0.00357877f $X=0.985 $Y=2.465 $X2=0 $Y2=0
cc_114 N_B2_c_91_n N_A_43_65#_c_570_n 3.18679e-19 $X=0.555 $Y=1.275 $X2=0 $Y2=0
cc_115 N_B2_c_91_n N_A_43_65#_c_576_n 0.0123501f $X=0.555 $Y=1.275 $X2=0 $Y2=0
cc_116 N_B2_c_93_n N_A_43_65#_c_576_n 0.0124617f $X=0.985 $Y=1.275 $X2=0 $Y2=0
cc_117 N_B2_c_95_n N_A_43_65#_c_576_n 0.0283744f $X=0.895 $Y=1.44 $X2=0 $Y2=0
cc_118 B2 N_A_43_65#_c_576_n 0.00219355f $X=0.155 $Y=1.58 $X2=0 $Y2=0
cc_119 N_B2_c_97_n N_A_43_65#_c_576_n 0.00214617f $X=0.985 $Y=1.44 $X2=0 $Y2=0
cc_120 B2 N_A_43_65#_c_571_n 0.0230488f $X=0.155 $Y=1.58 $X2=0 $Y2=0
cc_121 N_B2_c_97_n N_A_43_65#_c_571_n 0.00130258f $X=0.985 $Y=1.44 $X2=0 $Y2=0
cc_122 N_B2_c_93_n N_A_43_65#_c_573_n 4.90985e-19 $X=0.985 $Y=1.275 $X2=0 $Y2=0
cc_123 N_B2_c_91_n N_VGND_c_605_n 0.0112436f $X=0.555 $Y=1.275 $X2=0 $Y2=0
cc_124 N_B2_c_93_n N_VGND_c_605_n 0.00884972f $X=0.985 $Y=1.275 $X2=0 $Y2=0
cc_125 N_B2_c_91_n N_VGND_c_609_n 0.00414769f $X=0.555 $Y=1.275 $X2=0 $Y2=0
cc_126 N_B2_c_93_n N_VGND_c_610_n 0.00414769f $X=0.985 $Y=1.275 $X2=0 $Y2=0
cc_127 N_B2_c_91_n N_VGND_c_614_n 0.00825965f $X=0.555 $Y=1.275 $X2=0 $Y2=0
cc_128 N_B2_c_93_n N_VGND_c_614_n 0.0078848f $X=0.985 $Y=1.275 $X2=0 $Y2=0
cc_129 N_B1_M1008_g N_A1_M1016_g 0.0291915f $X=1.845 $Y=2.465 $X2=0 $Y2=0
cc_130 N_B1_c_144_n N_A1_c_200_n 2.86633e-19 $X=2.06 $Y=1.51 $X2=0 $Y2=0
cc_131 N_B1_c_145_n N_A1_c_200_n 0.0259188f $X=2.06 $Y=1.51 $X2=0 $Y2=0
cc_132 N_B1_c_144_n N_A1_c_197_n 0.0232961f $X=2.06 $Y=1.51 $X2=0 $Y2=0
cc_133 N_B1_c_145_n N_A1_c_197_n 0.00218889f $X=2.06 $Y=1.51 $X2=0 $Y2=0
cc_134 N_B1_M1000_g N_A_43_367#_c_346_n 0.0115031f $X=1.415 $Y=2.465 $X2=0 $Y2=0
cc_135 N_B1_M1008_g N_A_43_367#_c_346_n 0.0143316f $X=1.845 $Y=2.465 $X2=0 $Y2=0
cc_136 N_B1_M1008_g N_A_43_367#_c_348_n 0.00186948f $X=1.845 $Y=2.465 $X2=0
+ $Y2=0
cc_137 N_B1_M1008_g N_A_43_367#_c_349_n 0.00762323f $X=1.845 $Y=2.465 $X2=0
+ $Y2=0
cc_138 N_B1_M1000_g N_Y_c_414_n 6.32676e-19 $X=1.415 $Y=2.465 $X2=0 $Y2=0
cc_139 N_B1_M1000_g N_Y_c_410_n 0.0148906f $X=1.415 $Y=2.465 $X2=0 $Y2=0
cc_140 N_B1_M1003_g N_Y_c_427_n 0.00532477f $X=1.415 $Y=0.745 $X2=0 $Y2=0
cc_141 N_B1_M1009_g N_Y_c_427_n 0.0108481f $X=1.845 $Y=0.745 $X2=0 $Y2=0
cc_142 N_B1_M1000_g N_Y_c_412_n 0.00608255f $X=1.415 $Y=2.465 $X2=0 $Y2=0
cc_143 N_B1_M1008_g N_Y_c_412_n 0.00428499f $X=1.845 $Y=2.465 $X2=0 $Y2=0
cc_144 N_B1_c_143_n N_Y_c_412_n 0.00231975f $X=1.77 $Y=1.51 $X2=0 $Y2=0
cc_145 N_B1_c_145_n N_Y_c_412_n 0.00467424f $X=2.06 $Y=1.51 $X2=0 $Y2=0
cc_146 N_B1_M1000_g N_Y_c_433_n 0.00653266f $X=1.415 $Y=2.465 $X2=0 $Y2=0
cc_147 N_B1_M1008_g N_Y_c_433_n 0.00916872f $X=1.845 $Y=2.465 $X2=0 $Y2=0
cc_148 N_B1_M1009_g N_Y_c_408_n 0.0126997f $X=1.845 $Y=0.745 $X2=0 $Y2=0
cc_149 N_B1_c_144_n N_Y_c_408_n 0.00746539f $X=2.06 $Y=1.51 $X2=0 $Y2=0
cc_150 N_B1_c_145_n N_Y_c_408_n 0.0266536f $X=2.06 $Y=1.51 $X2=0 $Y2=0
cc_151 N_B1_M1003_g N_Y_c_409_n 0.00484921f $X=1.415 $Y=0.745 $X2=0 $Y2=0
cc_152 N_B1_M1009_g N_Y_c_409_n 0.0020193f $X=1.845 $Y=0.745 $X2=0 $Y2=0
cc_153 N_B1_c_143_n N_Y_c_409_n 0.00262919f $X=1.77 $Y=1.51 $X2=0 $Y2=0
cc_154 N_B1_M1008_g N_Y_c_441_n 0.0146217f $X=1.845 $Y=2.465 $X2=0 $Y2=0
cc_155 N_B1_c_144_n N_Y_c_441_n 0.00167113f $X=2.06 $Y=1.51 $X2=0 $Y2=0
cc_156 N_B1_c_145_n N_Y_c_441_n 0.0268307f $X=2.06 $Y=1.51 $X2=0 $Y2=0
cc_157 N_B1_M1000_g N_VPWR_c_495_n 0.00537654f $X=1.415 $Y=2.465 $X2=0 $Y2=0
cc_158 N_B1_M1008_g N_VPWR_c_495_n 0.00594945f $X=1.845 $Y=2.465 $X2=0 $Y2=0
cc_159 N_B1_M1000_g N_VPWR_c_503_n 0.00357877f $X=1.415 $Y=2.465 $X2=0 $Y2=0
cc_160 N_B1_M1008_g N_VPWR_c_503_n 0.00357877f $X=1.845 $Y=2.465 $X2=0 $Y2=0
cc_161 N_B1_M1008_g N_VPWR_c_504_n 0.00103424f $X=1.845 $Y=2.465 $X2=0 $Y2=0
cc_162 N_B1_M1003_g N_A_43_65#_c_572_n 0.0117888f $X=1.415 $Y=0.745 $X2=0 $Y2=0
cc_163 N_B1_M1009_g N_A_43_65#_c_572_n 0.0127722f $X=1.845 $Y=0.745 $X2=0 $Y2=0
cc_164 N_B1_M1003_g N_VGND_c_605_n 5.59621e-19 $X=1.415 $Y=0.745 $X2=0 $Y2=0
cc_165 N_B1_M1003_g N_VGND_c_610_n 0.0030414f $X=1.415 $Y=0.745 $X2=0 $Y2=0
cc_166 N_B1_M1009_g N_VGND_c_610_n 0.0030414f $X=1.845 $Y=0.745 $X2=0 $Y2=0
cc_167 N_B1_M1003_g N_VGND_c_614_n 0.00435814f $X=1.415 $Y=0.745 $X2=0 $Y2=0
cc_168 N_B1_M1009_g N_VGND_c_614_n 0.00484828f $X=1.845 $Y=0.745 $X2=0 $Y2=0
cc_169 N_B1_M1009_g N_A_509_65#_c_673_n 6.31847e-19 $X=1.845 $Y=0.745 $X2=0
+ $Y2=0
cc_170 N_A1_M1015_g N_A2_M1004_g 0.0179726f $X=3.385 $Y=0.745 $X2=0 $Y2=0
cc_171 N_A1_M1019_g N_A2_M1002_g 0.0130324f $X=3.385 $Y=2.465 $X2=0 $Y2=0
cc_172 N_A1_c_197_n A2 0.00319856f $X=3.385 $Y=1.51 $X2=0 $Y2=0
cc_173 N_A1_c_197_n N_A2_c_252_n 0.0179726f $X=3.385 $Y=1.51 $X2=0 $Y2=0
cc_174 N_A1_M1016_g N_A_43_367#_c_346_n 0.00186905f $X=2.51 $Y=2.465 $X2=0 $Y2=0
cc_175 N_A1_M1016_g N_A_43_367#_c_349_n 0.00767499f $X=2.51 $Y=2.465 $X2=0 $Y2=0
cc_176 N_A1_M1016_g N_A_43_367#_c_352_n 0.0170366f $X=2.51 $Y=2.465 $X2=0 $Y2=0
cc_177 N_A1_M1019_g N_A_43_367#_c_352_n 0.0180292f $X=3.385 $Y=2.465 $X2=0 $Y2=0
cc_178 N_A1_c_197_n N_A_43_367#_c_352_n 8.6126e-19 $X=3.385 $Y=1.51 $X2=0 $Y2=0
cc_179 N_A1_M1016_g N_Y_c_433_n 9.05045e-19 $X=2.51 $Y=2.465 $X2=0 $Y2=0
cc_180 N_A1_M1007_g N_Y_c_408_n 0.012645f $X=2.955 $Y=0.745 $X2=0 $Y2=0
cc_181 N_A1_c_200_n N_Y_c_408_n 0.0236922f $X=2.6 $Y=1.51 $X2=0 $Y2=0
cc_182 N_A1_c_197_n N_Y_c_408_n 0.0125553f $X=3.385 $Y=1.51 $X2=0 $Y2=0
cc_183 N_A1_M1016_g N_Y_c_441_n 0.015205f $X=2.51 $Y=2.465 $X2=0 $Y2=0
cc_184 N_A1_c_200_n N_Y_c_441_n 0.0228449f $X=2.6 $Y=1.51 $X2=0 $Y2=0
cc_185 N_A1_c_197_n N_Y_c_441_n 0.00703103f $X=3.385 $Y=1.51 $X2=0 $Y2=0
cc_186 N_A1_M1007_g Y 0.0013353f $X=2.955 $Y=0.745 $X2=0 $Y2=0
cc_187 N_A1_M1015_g Y 0.00296996f $X=3.385 $Y=0.745 $X2=0 $Y2=0
cc_188 N_A1_M1007_g N_Y_c_453_n 0.0108489f $X=2.955 $Y=0.745 $X2=0 $Y2=0
cc_189 N_A1_M1015_g N_Y_c_453_n 0.00506777f $X=3.385 $Y=0.745 $X2=0 $Y2=0
cc_190 N_A1_M1019_g N_Y_c_455_n 0.00726696f $X=3.385 $Y=2.465 $X2=0 $Y2=0
cc_191 N_A1_M1016_g Y 0.00519078f $X=2.51 $Y=2.465 $X2=0 $Y2=0
cc_192 N_A1_M1007_g Y 0.00542709f $X=2.955 $Y=0.745 $X2=0 $Y2=0
cc_193 N_A1_M1015_g Y 0.00297013f $X=3.385 $Y=0.745 $X2=0 $Y2=0
cc_194 N_A1_M1019_g Y 0.00899772f $X=3.385 $Y=2.465 $X2=0 $Y2=0
cc_195 N_A1_c_200_n Y 0.0191526f $X=2.6 $Y=1.51 $X2=0 $Y2=0
cc_196 N_A1_c_197_n Y 0.0285648f $X=3.385 $Y=1.51 $X2=0 $Y2=0
cc_197 N_A1_M1019_g N_VPWR_c_496_n 5.91826e-19 $X=3.385 $Y=2.465 $X2=0 $Y2=0
cc_198 N_A1_M1019_g N_VPWR_c_500_n 0.00486043f $X=3.385 $Y=2.465 $X2=0 $Y2=0
cc_199 N_A1_M1016_g N_VPWR_c_495_n 0.00883374f $X=2.51 $Y=2.465 $X2=0 $Y2=0
cc_200 N_A1_M1019_g N_VPWR_c_495_n 0.00840461f $X=3.385 $Y=2.465 $X2=0 $Y2=0
cc_201 N_A1_M1016_g N_VPWR_c_503_n 0.00486043f $X=2.51 $Y=2.465 $X2=0 $Y2=0
cc_202 N_A1_M1016_g N_VPWR_c_504_n 0.0156966f $X=2.51 $Y=2.465 $X2=0 $Y2=0
cc_203 N_A1_M1019_g N_VPWR_c_504_n 0.0140679f $X=3.385 $Y=2.465 $X2=0 $Y2=0
cc_204 N_A1_M1007_g N_A_43_65#_c_572_n 6.31847e-19 $X=2.955 $Y=0.745 $X2=0 $Y2=0
cc_205 N_A1_M1007_g N_VGND_c_610_n 0.0030414f $X=2.955 $Y=0.745 $X2=0 $Y2=0
cc_206 N_A1_M1015_g N_VGND_c_610_n 0.0030414f $X=3.385 $Y=0.745 $X2=0 $Y2=0
cc_207 N_A1_M1007_g N_VGND_c_614_n 0.00484828f $X=2.955 $Y=0.745 $X2=0 $Y2=0
cc_208 N_A1_M1015_g N_VGND_c_614_n 0.00435814f $X=3.385 $Y=0.745 $X2=0 $Y2=0
cc_209 N_A1_M1007_g N_A_509_65#_c_672_n 0.0128187f $X=2.955 $Y=0.745 $X2=0 $Y2=0
cc_210 N_A1_M1015_g N_A_509_65#_c_672_n 0.0119279f $X=3.385 $Y=0.745 $X2=0 $Y2=0
cc_211 N_A1_M1015_g N_A_509_65#_c_674_n 0.00105828f $X=3.385 $Y=0.745 $X2=0
+ $Y2=0
cc_212 N_A2_M1018_g N_A3_M1001_g 0.01869f $X=4.695 $Y=2.465 $X2=0 $Y2=0
cc_213 A2 N_A3_c_304_n 0.00167934f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_214 N_A2_c_252_n N_A3_c_304_n 0.01869f $X=4.695 $Y=1.51 $X2=0 $Y2=0
cc_215 A2 N_A_43_367#_c_355_n 0.0218862f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_216 N_A2_M1002_g N_A_43_367#_c_356_n 0.0137046f $X=3.895 $Y=2.465 $X2=0 $Y2=0
cc_217 N_A2_M1018_g N_A_43_367#_c_356_n 0.0151769f $X=4.695 $Y=2.465 $X2=0 $Y2=0
cc_218 A2 N_A_43_367#_c_356_n 0.0614961f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_219 N_A2_c_252_n N_A_43_367#_c_356_n 0.00269998f $X=4.695 $Y=1.51 $X2=0 $Y2=0
cc_220 N_A2_M1018_g N_A_43_367#_c_339_n 0.00250406f $X=4.695 $Y=2.465 $X2=0
+ $Y2=0
cc_221 N_A2_M1004_g Y 9.50304e-19 $X=3.815 $Y=0.745 $X2=0 $Y2=0
cc_222 N_A2_M1002_g Y 7.82547e-19 $X=3.895 $Y=2.465 $X2=0 $Y2=0
cc_223 A2 Y 0.0260513f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_224 N_A2_M1002_g N_VPWR_c_496_n 0.0175399f $X=3.895 $Y=2.465 $X2=0 $Y2=0
cc_225 N_A2_M1018_g N_VPWR_c_496_n 0.0172734f $X=4.695 $Y=2.465 $X2=0 $Y2=0
cc_226 N_A2_M1018_g N_VPWR_c_497_n 7.27171e-19 $X=4.695 $Y=2.465 $X2=0 $Y2=0
cc_227 N_A2_M1018_g N_VPWR_c_498_n 0.00486043f $X=4.695 $Y=2.465 $X2=0 $Y2=0
cc_228 N_A2_M1002_g N_VPWR_c_500_n 0.00486043f $X=3.895 $Y=2.465 $X2=0 $Y2=0
cc_229 N_A2_M1002_g N_VPWR_c_495_n 0.00845345f $X=3.895 $Y=2.465 $X2=0 $Y2=0
cc_230 N_A2_M1018_g N_VPWR_c_495_n 0.0082726f $X=4.695 $Y=2.465 $X2=0 $Y2=0
cc_231 N_A2_M1002_g N_VPWR_c_504_n 5.54446e-19 $X=3.895 $Y=2.465 $X2=0 $Y2=0
cc_232 N_A2_M1010_g N_VGND_c_606_n 0.00245665f $X=4.245 $Y=0.745 $X2=0 $Y2=0
cc_233 N_A2_M1004_g N_VGND_c_610_n 0.0030414f $X=3.815 $Y=0.745 $X2=0 $Y2=0
cc_234 N_A2_M1010_g N_VGND_c_610_n 0.0030414f $X=4.245 $Y=0.745 $X2=0 $Y2=0
cc_235 N_A2_M1004_g N_VGND_c_614_n 0.00435814f $X=3.815 $Y=0.745 $X2=0 $Y2=0
cc_236 N_A2_M1010_g N_VGND_c_614_n 0.00484828f $X=4.245 $Y=0.745 $X2=0 $Y2=0
cc_237 N_A2_M1004_g N_A_509_65#_c_674_n 0.00105828f $X=3.815 $Y=0.745 $X2=0
+ $Y2=0
cc_238 A2 N_A_509_65#_c_674_n 0.0131937f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_239 N_A2_M1004_g N_A_509_65#_c_675_n 0.0119279f $X=3.815 $Y=0.745 $X2=0 $Y2=0
cc_240 N_A2_M1010_g N_A_509_65#_c_675_n 0.0128187f $X=4.245 $Y=0.745 $X2=0 $Y2=0
cc_241 N_A2_M1004_g N_A_778_65#_c_713_n 0.00506691f $X=3.815 $Y=0.745 $X2=0
+ $Y2=0
cc_242 N_A2_M1010_g N_A_778_65#_c_713_n 0.0108481f $X=4.245 $Y=0.745 $X2=0 $Y2=0
cc_243 N_A2_M1010_g N_A_778_65#_c_711_n 0.0112556f $X=4.245 $Y=0.745 $X2=0 $Y2=0
cc_244 A2 N_A_778_65#_c_711_n 0.0325691f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_245 N_A2_c_252_n N_A_778_65#_c_711_n 0.0126712f $X=4.695 $Y=1.51 $X2=0 $Y2=0
cc_246 N_A2_M1004_g N_A_778_65#_c_712_n 0.0033274f $X=3.815 $Y=0.745 $X2=0 $Y2=0
cc_247 N_A2_M1010_g N_A_778_65#_c_712_n 0.00169274f $X=4.245 $Y=0.745 $X2=0
+ $Y2=0
cc_248 A2 N_A_778_65#_c_712_n 0.0262733f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_249 N_A2_c_252_n N_A_778_65#_c_712_n 0.00288587f $X=4.695 $Y=1.51 $X2=0 $Y2=0
cc_250 N_A3_M1001_g N_A_43_367#_c_340_n 0.0146899f $X=5.125 $Y=2.465 $X2=0 $Y2=0
cc_251 N_A3_M1014_g N_A_43_367#_c_340_n 0.0163258f $X=5.555 $Y=2.465 $X2=0 $Y2=0
cc_252 A3 N_A_43_367#_c_340_n 0.01211f $X=5.915 $Y=1.21 $X2=0 $Y2=0
cc_253 N_A3_c_304_n N_A_43_367#_c_340_n 0.0122977f $X=5.84 $Y=1.36 $X2=0 $Y2=0
cc_254 N_A3_M1001_g N_VPWR_c_496_n 6.94228e-19 $X=5.125 $Y=2.465 $X2=0 $Y2=0
cc_255 N_A3_M1001_g N_VPWR_c_497_n 0.0142189f $X=5.125 $Y=2.465 $X2=0 $Y2=0
cc_256 N_A3_M1014_g N_VPWR_c_497_n 0.0161992f $X=5.555 $Y=2.465 $X2=0 $Y2=0
cc_257 N_A3_M1001_g N_VPWR_c_498_n 0.00486043f $X=5.125 $Y=2.465 $X2=0 $Y2=0
cc_258 N_A3_M1014_g N_VPWR_c_501_n 0.00486043f $X=5.555 $Y=2.465 $X2=0 $Y2=0
cc_259 N_A3_M1001_g N_VPWR_c_495_n 0.0082726f $X=5.125 $Y=2.465 $X2=0 $Y2=0
cc_260 N_A3_M1014_g N_VPWR_c_495_n 0.0093271f $X=5.555 $Y=2.465 $X2=0 $Y2=0
cc_261 N_A3_c_300_n N_VGND_c_606_n 0.0126339f $X=5.275 $Y=1.195 $X2=0 $Y2=0
cc_262 N_A3_c_302_n N_VGND_c_606_n 6.15775e-19 $X=5.705 $Y=1.195 $X2=0 $Y2=0
cc_263 N_A3_c_304_n N_VGND_c_606_n 7.36808e-19 $X=5.84 $Y=1.36 $X2=0 $Y2=0
cc_264 N_A3_c_300_n N_VGND_c_608_n 6.49724e-19 $X=5.275 $Y=1.195 $X2=0 $Y2=0
cc_265 N_A3_c_302_n N_VGND_c_608_n 0.0162804f $X=5.705 $Y=1.195 $X2=0 $Y2=0
cc_266 A3 N_VGND_c_608_n 0.0248138f $X=5.915 $Y=1.21 $X2=0 $Y2=0
cc_267 N_A3_c_304_n N_VGND_c_608_n 0.00506784f $X=5.84 $Y=1.36 $X2=0 $Y2=0
cc_268 N_A3_c_300_n N_VGND_c_611_n 0.00477554f $X=5.275 $Y=1.195 $X2=0 $Y2=0
cc_269 N_A3_c_302_n N_VGND_c_611_n 0.00477554f $X=5.705 $Y=1.195 $X2=0 $Y2=0
cc_270 N_A3_c_300_n N_VGND_c_614_n 0.00825815f $X=5.275 $Y=1.195 $X2=0 $Y2=0
cc_271 N_A3_c_302_n N_VGND_c_614_n 0.00825815f $X=5.705 $Y=1.195 $X2=0 $Y2=0
cc_272 N_A3_c_300_n N_A_509_65#_c_676_n 8.44365e-19 $X=5.275 $Y=1.195 $X2=0
+ $Y2=0
cc_273 N_A3_c_300_n N_A_778_65#_c_711_n 0.0113656f $X=5.275 $Y=1.195 $X2=0 $Y2=0
cc_274 N_A3_c_302_n N_A_778_65#_c_711_n 0.00349191f $X=5.705 $Y=1.195 $X2=0
+ $Y2=0
cc_275 A3 N_A_778_65#_c_711_n 0.00398701f $X=5.915 $Y=1.21 $X2=0 $Y2=0
cc_276 N_A3_c_304_n N_A_778_65#_c_711_n 0.0225105f $X=5.84 $Y=1.36 $X2=0 $Y2=0
cc_277 N_A_43_367#_c_344_n N_Y_M1005_d 0.00332344f $X=1.105 $Y=2.99 $X2=0 $Y2=0
cc_278 N_A_43_367#_c_346_n N_Y_M1000_s 0.00332344f $X=2.015 $Y=2.99 $X2=0 $Y2=0
cc_279 N_A_43_367#_c_344_n N_Y_c_414_n 0.0159805f $X=1.105 $Y=2.99 $X2=0 $Y2=0
cc_280 N_A_43_367#_M1011_s N_Y_c_410_n 0.00176461f $X=1.06 $Y=1.835 $X2=0 $Y2=0
cc_281 N_A_43_367#_c_369_p N_Y_c_410_n 0.0135055f $X=1.2 $Y=2.2 $X2=0 $Y2=0
cc_282 N_A_43_367#_c_346_n N_Y_c_433_n 0.0159805f $X=2.015 $Y=2.99 $X2=0 $Y2=0
cc_283 N_A_43_367#_c_348_n N_Y_c_433_n 0.0115078f $X=2.18 $Y=2.46 $X2=0 $Y2=0
cc_284 N_A_43_367#_c_349_n N_Y_c_433_n 0.017477f $X=2.18 $Y=2.905 $X2=0 $Y2=0
cc_285 N_A_43_367#_M1008_d N_Y_c_441_n 0.0119078f $X=1.92 $Y=1.835 $X2=0 $Y2=0
cc_286 N_A_43_367#_c_348_n N_Y_c_441_n 0.0271453f $X=2.18 $Y=2.46 $X2=0 $Y2=0
cc_287 N_A_43_367#_c_352_n N_Y_c_441_n 0.0392711f $X=3.505 $Y=2.375 $X2=0 $Y2=0
cc_288 N_A_43_367#_c_352_n N_Y_c_455_n 0.0219943f $X=3.505 $Y=2.375 $X2=0 $Y2=0
cc_289 N_A_43_367#_c_352_n N_VPWR_M1016_s 0.015923f $X=3.505 $Y=2.375 $X2=-0.19
+ $Y2=1.655
cc_290 N_A_43_367#_c_356_n N_VPWR_M1002_s 0.0131419f $X=4.815 $Y=2.005 $X2=0
+ $Y2=0
cc_291 N_A_43_367#_c_340_n N_VPWR_M1001_s 0.00176461f $X=5.675 $Y=1.84 $X2=0
+ $Y2=0
cc_292 N_A_43_367#_c_356_n N_VPWR_c_496_n 0.0471803f $X=4.815 $Y=2.005 $X2=0
+ $Y2=0
cc_293 N_A_43_367#_c_340_n N_VPWR_c_497_n 0.0170777f $X=5.675 $Y=1.84 $X2=0
+ $Y2=0
cc_294 N_A_43_367#_c_382_p N_VPWR_c_498_n 0.0124525f $X=4.91 $Y=2.445 $X2=0
+ $Y2=0
cc_295 N_A_43_367#_c_383_p N_VPWR_c_500_n 0.0180775f $X=3.64 $Y=2.485 $X2=0
+ $Y2=0
cc_296 N_A_43_367#_c_341_n N_VPWR_c_501_n 0.0178111f $X=5.77 $Y=1.98 $X2=0 $Y2=0
cc_297 N_A_43_367#_M1005_s N_VPWR_c_495_n 0.00215161f $X=0.215 $Y=1.835 $X2=0
+ $Y2=0
cc_298 N_A_43_367#_M1011_s N_VPWR_c_495_n 0.00223565f $X=1.06 $Y=1.835 $X2=0
+ $Y2=0
cc_299 N_A_43_367#_M1008_d N_VPWR_c_495_n 0.00732452f $X=1.92 $Y=1.835 $X2=0
+ $Y2=0
cc_300 N_A_43_367#_M1019_d N_VPWR_c_495_n 0.0060098f $X=3.46 $Y=1.835 $X2=0
+ $Y2=0
cc_301 N_A_43_367#_M1018_d N_VPWR_c_495_n 0.00536646f $X=4.77 $Y=1.835 $X2=0
+ $Y2=0
cc_302 N_A_43_367#_M1014_d N_VPWR_c_495_n 0.00371702f $X=5.63 $Y=1.835 $X2=0
+ $Y2=0
cc_303 N_A_43_367#_c_337_n N_VPWR_c_495_n 0.0101029f $X=0.305 $Y=2.905 $X2=0
+ $Y2=0
cc_304 N_A_43_367#_c_344_n N_VPWR_c_495_n 0.023676f $X=1.105 $Y=2.99 $X2=0 $Y2=0
cc_305 N_A_43_367#_c_346_n N_VPWR_c_495_n 0.0384562f $X=2.015 $Y=2.99 $X2=0
+ $Y2=0
cc_306 N_A_43_367#_c_383_p N_VPWR_c_495_n 0.0104192f $X=3.64 $Y=2.485 $X2=0
+ $Y2=0
cc_307 N_A_43_367#_c_382_p N_VPWR_c_495_n 0.00729844f $X=4.91 $Y=2.445 $X2=0
+ $Y2=0
cc_308 N_A_43_367#_c_341_n N_VPWR_c_495_n 0.0100304f $X=5.77 $Y=1.98 $X2=0 $Y2=0
cc_309 N_A_43_367#_c_397_p N_VPWR_c_495_n 0.00738676f $X=1.2 $Y=2.99 $X2=0 $Y2=0
cc_310 N_A_43_367#_c_337_n N_VPWR_c_503_n 0.0179183f $X=0.305 $Y=2.905 $X2=0
+ $Y2=0
cc_311 N_A_43_367#_c_344_n N_VPWR_c_503_n 0.0361172f $X=1.105 $Y=2.99 $X2=0
+ $Y2=0
cc_312 N_A_43_367#_c_346_n N_VPWR_c_503_n 0.0621503f $X=2.015 $Y=2.99 $X2=0
+ $Y2=0
cc_313 N_A_43_367#_c_397_p N_VPWR_c_503_n 0.0125234f $X=1.2 $Y=2.99 $X2=0 $Y2=0
cc_314 N_A_43_367#_c_346_n N_VPWR_c_504_n 0.0123794f $X=2.015 $Y=2.99 $X2=0
+ $Y2=0
cc_315 N_A_43_367#_c_349_n N_VPWR_c_504_n 0.0187893f $X=2.18 $Y=2.905 $X2=0
+ $Y2=0
cc_316 N_A_43_367#_c_352_n N_VPWR_c_504_n 0.0531571f $X=3.505 $Y=2.375 $X2=0
+ $Y2=0
cc_317 N_A_43_367#_c_356_n N_A_778_65#_c_711_n 0.00348361f $X=4.815 $Y=2.005
+ $X2=0 $Y2=0
cc_318 N_A_43_367#_c_339_n N_A_778_65#_c_711_n 0.00708768f $X=4.91 $Y=2.09 $X2=0
+ $Y2=0
cc_319 N_A_43_367#_c_340_n N_A_778_65#_c_711_n 0.0180213f $X=5.675 $Y=1.84 $X2=0
+ $Y2=0
cc_320 N_Y_c_441_n N_VPWR_M1016_s 0.0111123f $X=3.005 $Y=2.02 $X2=-0.19
+ $Y2=-0.245
cc_321 N_Y_c_455_n N_VPWR_M1016_s 0.00412384f $X=3.17 $Y=1.92 $X2=-0.19
+ $Y2=-0.245
cc_322 Y N_VPWR_M1016_s 0.00174419f $X=3.12 $Y=1.295 $X2=-0.19 $Y2=-0.245
cc_323 N_Y_M1005_d N_VPWR_c_495_n 0.00225186f $X=0.63 $Y=1.835 $X2=0 $Y2=0
cc_324 N_Y_M1000_s N_VPWR_c_495_n 0.00225186f $X=1.49 $Y=1.835 $X2=0 $Y2=0
cc_325 N_Y_c_408_n N_A_43_65#_M1009_s 0.00371875f $X=3.005 $Y=1.16 $X2=0 $Y2=0
cc_326 N_Y_c_410_n N_A_43_65#_c_576_n 0.00548784f $X=1.465 $Y=1.78 $X2=0 $Y2=0
cc_327 N_Y_M1003_d N_A_43_65#_c_572_n 0.00176461f $X=1.49 $Y=0.325 $X2=0 $Y2=0
cc_328 N_Y_c_427_n N_A_43_65#_c_572_n 0.0159398f $X=1.63 $Y=0.69 $X2=0 $Y2=0
cc_329 N_Y_c_408_n N_A_43_65#_c_572_n 0.00280043f $X=3.005 $Y=1.16 $X2=0 $Y2=0
cc_330 N_Y_c_408_n N_A_43_65#_c_574_n 0.0257834f $X=3.005 $Y=1.16 $X2=0 $Y2=0
cc_331 N_Y_c_408_n N_A_509_65#_M1007_s 0.00371875f $X=3.005 $Y=1.16 $X2=-0.19
+ $Y2=-0.245
cc_332 N_Y_c_408_n N_A_509_65#_c_671_n 0.0257834f $X=3.005 $Y=1.16 $X2=0 $Y2=0
cc_333 N_Y_M1007_d N_A_509_65#_c_672_n 0.00176461f $X=3.03 $Y=0.325 $X2=0 $Y2=0
cc_334 N_Y_c_408_n N_A_509_65#_c_672_n 0.00280043f $X=3.005 $Y=1.16 $X2=0 $Y2=0
cc_335 N_Y_c_453_n N_A_509_65#_c_672_n 0.0160148f $X=3.17 $Y=0.69 $X2=0 $Y2=0
cc_336 Y N_A_509_65#_c_674_n 0.00697473f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_337 Y N_A_778_65#_c_712_n 0.00132601f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_338 N_A_43_65#_c_576_n N_VGND_M1012_d 0.00355045f $X=1.105 $Y=0.955 $X2=-0.19
+ $Y2=-0.245
cc_339 N_A_43_65#_c_570_n N_VGND_c_605_n 0.0148073f $X=0.34 $Y=0.48 $X2=0 $Y2=0
cc_340 N_A_43_65#_c_576_n N_VGND_c_605_n 0.0170777f $X=1.105 $Y=0.955 $X2=0
+ $Y2=0
cc_341 N_A_43_65#_c_573_n N_VGND_c_605_n 0.00915965f $X=1.295 $Y=0.35 $X2=0
+ $Y2=0
cc_342 N_A_43_65#_c_570_n N_VGND_c_609_n 0.0133857f $X=0.34 $Y=0.48 $X2=0 $Y2=0
cc_343 N_A_43_65#_c_572_n N_VGND_c_610_n 0.0618603f $X=1.965 $Y=0.35 $X2=0 $Y2=0
cc_344 N_A_43_65#_c_573_n N_VGND_c_610_n 0.0128106f $X=1.295 $Y=0.35 $X2=0 $Y2=0
cc_345 N_A_43_65#_c_570_n N_VGND_c_614_n 0.00972454f $X=0.34 $Y=0.48 $X2=0 $Y2=0
cc_346 N_A_43_65#_c_572_n N_VGND_c_614_n 0.036406f $X=1.965 $Y=0.35 $X2=0 $Y2=0
cc_347 N_A_43_65#_c_573_n N_VGND_c_614_n 0.0073517f $X=1.295 $Y=0.35 $X2=0 $Y2=0
cc_348 N_A_43_65#_c_574_n N_A_509_65#_c_671_n 0.0336785f $X=2.13 $Y=0.47 $X2=0
+ $Y2=0
cc_349 N_A_43_65#_c_572_n N_A_509_65#_c_673_n 0.0137129f $X=1.965 $Y=0.35 $X2=0
+ $Y2=0
cc_350 N_VGND_c_610_n N_A_509_65#_c_672_n 0.0397112f $X=4.895 $Y=0 $X2=0 $Y2=0
cc_351 N_VGND_c_614_n N_A_509_65#_c_672_n 0.0236582f $X=6 $Y=0 $X2=0 $Y2=0
cc_352 N_VGND_c_610_n N_A_509_65#_c_673_n 0.0221491f $X=4.895 $Y=0 $X2=0 $Y2=0
cc_353 N_VGND_c_614_n N_A_509_65#_c_673_n 0.0127478f $X=6 $Y=0 $X2=0 $Y2=0
cc_354 N_VGND_c_606_n N_A_509_65#_c_675_n 0.0134079f $X=5.06 $Y=0.39 $X2=0 $Y2=0
cc_355 N_VGND_c_610_n N_A_509_65#_c_675_n 0.0618603f $X=4.895 $Y=0 $X2=0 $Y2=0
cc_356 N_VGND_c_614_n N_A_509_65#_c_675_n 0.036406f $X=6 $Y=0 $X2=0 $Y2=0
cc_357 N_VGND_c_606_n N_A_509_65#_c_676_n 0.0348796f $X=5.06 $Y=0.39 $X2=0 $Y2=0
cc_358 N_VGND_c_610_n N_A_509_65#_c_677_n 0.0128106f $X=4.895 $Y=0 $X2=0 $Y2=0
cc_359 N_VGND_c_614_n N_A_509_65#_c_677_n 0.0073517f $X=6 $Y=0 $X2=0 $Y2=0
cc_360 N_VGND_c_614_n N_A_778_65#_M1006_s 0.00536646f $X=6 $Y=0 $X2=0 $Y2=0
cc_361 N_VGND_M1006_d N_A_778_65#_c_711_n 0.00221108f $X=4.935 $Y=0.245 $X2=0
+ $Y2=0
cc_362 N_VGND_c_606_n N_A_778_65#_c_711_n 0.0220026f $X=5.06 $Y=0.39 $X2=0 $Y2=0
cc_363 N_VGND_c_611_n N_A_778_65#_c_733_n 0.0124525f $X=5.755 $Y=0 $X2=0 $Y2=0
cc_364 N_VGND_c_614_n N_A_778_65#_c_733_n 0.00730901f $X=6 $Y=0 $X2=0 $Y2=0
cc_365 N_A_509_65#_c_675_n N_A_778_65#_M1004_d 0.00176461f $X=4.365 $Y=0.35
+ $X2=-0.19 $Y2=-0.245
cc_366 N_A_509_65#_c_675_n N_A_778_65#_c_713_n 0.0159398f $X=4.365 $Y=0.35 $X2=0
+ $Y2=0
cc_367 N_A_509_65#_M1010_s N_A_778_65#_c_711_n 0.00371875f $X=4.32 $Y=0.325
+ $X2=0 $Y2=0
cc_368 N_A_509_65#_c_675_n N_A_778_65#_c_711_n 0.00280043f $X=4.365 $Y=0.35
+ $X2=0 $Y2=0
cc_369 N_A_509_65#_c_676_n N_A_778_65#_c_711_n 0.0257834f $X=4.53 $Y=0.47 $X2=0
+ $Y2=0
cc_370 N_A_509_65#_c_674_n N_A_778_65#_c_712_n 0.00697473f $X=3.6 $Y=0.47 $X2=0
+ $Y2=0
