* File: sky130_fd_sc_lp__or2_lp.pex.spice
* Created: Wed Sep  2 10:29:27 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__OR2_LP%A 3 7 11 17 20 21 22 23 34
c35 21 0 5.8403e-20 $X=0.72 $Y=1.295
r36 34 35 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.605
+ $Y=1.345 $X2=0.605 $Y2=1.345
r37 22 23 6.23308 $w=7.08e-07 $l=3.7e-07 $layer=LI1_cond $X=0.48 $Y=1.665
+ $X2=0.48 $Y2=2.035
r38 22 35 5.39078 $w=7.08e-07 $l=3.2e-07 $layer=LI1_cond $X=0.48 $Y=1.665
+ $X2=0.48 $Y2=1.345
r39 21 35 0.842309 $w=7.08e-07 $l=5e-08 $layer=LI1_cond $X=0.48 $Y=1.295
+ $X2=0.48 $Y2=1.345
r40 19 34 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.605 $Y=1.685
+ $X2=0.605 $Y2=1.345
r41 19 20 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.605 $Y=1.685
+ $X2=0.605 $Y2=1.85
r42 16 34 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=0.605 $Y=1.33
+ $X2=0.605 $Y2=1.345
r43 16 17 153.83 $w=1.5e-07 $l=3e-07 $layer=POLY_cond $X=0.605 $Y=1.255
+ $X2=0.905 $Y2=1.255
r44 13 16 46.1489 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=0.515 $Y=1.255
+ $X2=0.605 $Y2=1.255
r45 9 17 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.905 $Y=1.18
+ $X2=0.905 $Y2=1.255
r46 9 11 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=0.905 $Y=1.18 $X2=0.905
+ $Y2=0.78
r47 7 20 358.936 $w=1.5e-07 $l=7e-07 $layer=POLY_cond $X=0.695 $Y=2.55 $X2=0.695
+ $Y2=1.85
r48 1 13 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.515 $Y=1.18
+ $X2=0.515 $Y2=1.255
r49 1 3 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=0.515 $Y=1.18 $X2=0.515
+ $Y2=0.78
.ends

.subckt PM_SKY130_FD_SC_LP__OR2_LP%B 3 5 6 7 9 10 12 17 20 21 22 23 29
c51 17 0 5.8403e-20 $X=1.695 $Y=1.175
r52 22 23 13.5582 $w=3.38e-07 $l=4e-07 $layer=LI1_cond $X=1.625 $Y=1.265
+ $X2=1.625 $Y2=1.665
r53 22 29 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.62
+ $Y=1.265 $X2=1.62 $Y2=1.265
r54 21 22 11.5244 $w=3.38e-07 $l=3.4e-07 $layer=LI1_cond $X=1.625 $Y=0.925
+ $X2=1.625 $Y2=1.265
r55 20 21 12.5413 $w=3.38e-07 $l=3.7e-07 $layer=LI1_cond $X=1.625 $Y=0.555
+ $X2=1.625 $Y2=0.925
r56 19 29 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=1.62 $Y=1.62
+ $X2=1.62 $Y2=1.265
r57 16 29 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=1.62 $Y=1.25
+ $X2=1.62 $Y2=1.265
r58 16 17 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.62 $Y=1.175
+ $X2=1.695 $Y2=1.175
r59 13 16 146.138 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=1.335 $Y=1.175
+ $X2=1.62 $Y2=1.175
r60 10 17 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.695 $Y=1.1
+ $X2=1.695 $Y2=1.175
r61 10 12 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.695 $Y=1.1
+ $X2=1.695 $Y2=0.78
r62 7 13 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.335 $Y=1.1
+ $X2=1.335 $Y2=1.175
r63 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.335 $Y=1.1 $X2=1.335
+ $Y2=0.78
r64 5 19 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=1.455 $Y=1.695
+ $X2=1.62 $Y2=1.62
r65 5 6 151.266 $w=1.5e-07 $l=2.95e-07 $layer=POLY_cond $X=1.455 $Y=1.695
+ $X2=1.16 $Y2=1.695
r66 1 6 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.085 $Y=1.77
+ $X2=1.16 $Y2=1.695
r67 1 3 399.957 $w=1.5e-07 $l=7.8e-07 $layer=POLY_cond $X=1.085 $Y=1.77
+ $X2=1.085 $Y2=2.55
.ends

.subckt PM_SKY130_FD_SC_LP__OR2_LP%A_196_114# 1 2 9 13 17 21 24 27 29 33 37 40
+ 46
r79 45 46 21.9602 $w=6.7e-07 $l=2.75e-07 $layer=POLY_cond $X=2.46 $Y=1.925
+ $X2=2.735 $Y2=1.925
r80 44 45 9.18334 $w=6.7e-07 $l=1.15e-07 $layer=POLY_cond $X=2.345 $Y=1.925
+ $X2=2.46 $Y2=1.925
r81 37 39 10.7321 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=1.12 $Y=0.78
+ $X2=1.12 $Y2=1.01
r82 34 44 12.3775 $w=6.7e-07 $l=1.55e-07 $layer=POLY_cond $X=2.19 $Y=1.925
+ $X2=2.345 $Y2=1.925
r83 34 41 7.18696 $w=6.7e-07 $l=9e-08 $layer=POLY_cond $X=2.19 $Y=1.925 $X2=2.1
+ $Y2=1.925
r84 33 34 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.19
+ $Y=1.755 $X2=2.19 $Y2=1.755
r85 31 33 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=2.19 $Y=2.09
+ $X2=2.19 $Y2=1.755
r86 30 40 2.90867 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=1.465 $Y=2.175
+ $X2=1.29 $Y2=2.175
r87 29 31 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.025 $Y=2.175
+ $X2=2.19 $Y2=2.09
r88 29 30 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=2.025 $Y=2.175
+ $X2=1.465 $Y2=2.175
r89 25 40 3.58051 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=1.29 $Y=2.26 $X2=1.29
+ $Y2=2.175
r90 25 27 9.54881 $w=3.48e-07 $l=2.9e-07 $layer=LI1_cond $X=1.29 $Y=2.26
+ $X2=1.29 $Y2=2.55
r91 24 40 3.58051 $w=2.6e-07 $l=1.25499e-07 $layer=LI1_cond $X=1.2 $Y=2.09
+ $X2=1.29 $Y2=2.175
r92 24 39 70.4599 $w=1.68e-07 $l=1.08e-06 $layer=LI1_cond $X=1.2 $Y=2.09 $X2=1.2
+ $Y2=1.01
r93 19 46 38.9565 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=2.735 $Y=1.59
+ $X2=2.735 $Y2=1.925
r94 19 21 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=2.735 $Y=1.59
+ $X2=2.735 $Y2=0.78
r95 15 45 38.9565 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=2.46 $Y=2.26
+ $X2=2.46 $Y2=1.925
r96 15 17 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=2.46 $Y=2.26 $X2=2.46
+ $Y2=2.66
r97 11 44 38.9565 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=2.345 $Y=1.59
+ $X2=2.345 $Y2=1.925
r98 11 13 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=2.345 $Y=1.59
+ $X2=2.345 $Y2=0.78
r99 7 41 38.9565 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=2.1 $Y=2.26 $X2=2.1
+ $Y2=1.925
r100 7 9 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=2.1 $Y=2.26 $X2=2.1
+ $Y2=2.66
r101 2 27 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=1.16
+ $Y=2.34 $X2=1.3 $Y2=2.55
r102 1 37 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.98
+ $Y=0.57 $X2=1.12 $Y2=0.78
.ends

.subckt PM_SKY130_FD_SC_LP__OR2_LP%VPWR 1 2 9 13 16 17 19 20 21 37 38
r32 37 38 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r33 35 38 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r34 34 37 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.16 $Y=3.33 $X2=3.12
+ $Y2=3.33
r35 34 35 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r36 28 31 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.72 $Y=3.33 $X2=1.68
+ $Y2=3.33
r37 28 29 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r38 25 29 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r39 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r40 21 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r41 21 29 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.72 $Y2=3.33
r42 21 31 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r43 19 31 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=1.72 $Y=3.33 $X2=1.68
+ $Y2=3.33
r44 19 20 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.72 $Y=3.33
+ $X2=1.885 $Y2=3.33
r45 18 34 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=2.05 $Y=3.33
+ $X2=2.16 $Y2=3.33
r46 18 20 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.05 $Y=3.33
+ $X2=1.885 $Y2=3.33
r47 16 24 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=0.315 $Y=3.33
+ $X2=0.24 $Y2=3.33
r48 16 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.315 $Y=3.33
+ $X2=0.48 $Y2=3.33
r49 15 28 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=0.645 $Y=3.33
+ $X2=0.72 $Y2=3.33
r50 15 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.645 $Y=3.33
+ $X2=0.48 $Y2=3.33
r51 11 20 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.885 $Y=3.245
+ $X2=1.885 $Y2=3.33
r52 11 13 20.4297 $w=3.28e-07 $l=5.85e-07 $layer=LI1_cond $X=1.885 $Y=3.245
+ $X2=1.885 $Y2=2.66
r53 7 17 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.48 $Y=3.245 $X2=0.48
+ $Y2=3.33
r54 7 9 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=0.48 $Y=3.245
+ $X2=0.48 $Y2=2.55
r55 2 13 600 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=1 $X=1.74
+ $Y=2.45 $X2=1.885 $Y2=2.66
r56 1 9 600 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=1 $X=0.335
+ $Y=2.34 $X2=0.48 $Y2=2.55
.ends

.subckt PM_SKY130_FD_SC_LP__OR2_LP%X 1 2 10 13 14 15 16 17 45 48
r25 45 52 0.421154 $w=7.08e-07 $l=2.5e-08 $layer=LI1_cond $X=2.88 $Y=2.405
+ $X2=2.88 $Y2=2.43
r26 17 54 1.89723 $w=7.23e-07 $l=1.15e-07 $layer=LI1_cond $X=2.872 $Y=2.775
+ $X2=2.872 $Y2=2.66
r27 16 54 3.29953 $w=7.23e-07 $l=2e-07 $layer=LI1_cond $X=2.872 $Y=2.46
+ $X2=2.872 $Y2=2.66
r28 16 52 0.494929 $w=7.23e-07 $l=3e-08 $layer=LI1_cond $X=2.872 $Y=2.46
+ $X2=2.872 $Y2=2.43
r29 16 45 0.505385 $w=7.08e-07 $l=3e-08 $layer=LI1_cond $X=2.88 $Y=2.375
+ $X2=2.88 $Y2=2.405
r30 15 16 5.7277 $w=7.08e-07 $l=3.4e-07 $layer=LI1_cond $X=2.88 $Y=2.035
+ $X2=2.88 $Y2=2.375
r31 14 15 6.23308 $w=7.08e-07 $l=3.7e-07 $layer=LI1_cond $X=2.88 $Y=1.665
+ $X2=2.88 $Y2=2.035
r32 14 35 2.19 $w=7.08e-07 $l=1.3e-07 $layer=LI1_cond $X=2.88 $Y=1.665 $X2=2.88
+ $Y2=1.535
r33 13 35 4.04308 $w=7.08e-07 $l=2.4e-07 $layer=LI1_cond $X=2.88 $Y=1.295
+ $X2=2.88 $Y2=1.535
r34 13 48 10.0269 $w=7.08e-07 $l=1.15e-07 $layer=LI1_cond $X=2.88 $Y=1.295
+ $X2=2.88 $Y2=1.18
r35 12 48 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=2.87 $Y=1.01
+ $X2=2.87 $Y2=1.18
r36 10 12 10.7321 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=2.95 $Y=0.78
+ $X2=2.95 $Y2=1.01
r37 2 54 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=2.535
+ $Y=2.45 $X2=2.675 $Y2=2.66
r38 1 10 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.81
+ $Y=0.57 $X2=2.95 $Y2=0.78
.ends

.subckt PM_SKY130_FD_SC_LP__OR2_LP%VGND 1 2 7 9 13 15 17 27 28 34
r35 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r36 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r37 28 35 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.16
+ $Y2=0
r38 27 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r39 25 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.295 $Y=0 $X2=2.13
+ $Y2=0
r40 25 27 53.8235 $w=1.68e-07 $l=8.25e-07 $layer=LI1_cond $X=2.295 $Y=0 $X2=3.12
+ $Y2=0
r41 21 32 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r42 20 23 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r43 20 21 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r44 18 31 4.68787 $w=1.7e-07 $l=2.33e-07 $layer=LI1_cond $X=0.465 $Y=0 $X2=0.232
+ $Y2=0
r45 18 20 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.465 $Y=0 $X2=0.72
+ $Y2=0
r46 17 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.965 $Y=0 $X2=2.13
+ $Y2=0
r47 17 23 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.965 $Y=0 $X2=1.68
+ $Y2=0
r48 15 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r49 15 21 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=0.72
+ $Y2=0
r50 15 23 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r51 11 34 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.13 $Y=0.085
+ $X2=2.13 $Y2=0
r52 11 13 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=2.13 $Y=0.085
+ $X2=2.13 $Y2=0.78
r53 7 31 3.0783 $w=3.3e-07 $l=1.14039e-07 $layer=LI1_cond $X=0.3 $Y=0.085
+ $X2=0.232 $Y2=0
r54 7 9 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=0.3 $Y=0.085 $X2=0.3
+ $Y2=0.78
r55 2 13 182 $w=1.7e-07 $l=4.5299e-07 $layer=licon1_NDIFF $count=1 $X=1.77
+ $Y=0.57 $X2=2.13 $Y2=0.78
r56 1 9 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.155
+ $Y=0.57 $X2=0.3 $Y2=0.78
.ends

