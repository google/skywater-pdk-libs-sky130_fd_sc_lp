* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__a2bb2o_m A1_N A2_N B1 B2 VGND VNB VPB VPWR X
X0 VPWR B1 a_479_429# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X1 VGND A1_N a_210_125# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 VPWR A1_N a_223_535# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X3 a_223_535# A2_N a_210_125# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X4 X a_85_345# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X5 a_551_125# B1 VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 a_210_125# A2_N VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 a_85_345# a_210_125# a_479_429# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X8 X a_85_345# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 a_85_345# B2 a_551_125# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 VGND a_210_125# a_85_345# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X11 a_479_429# B2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
.ends
