* File: sky130_fd_sc_lp__and2b_m.pex.spice
* Created: Fri Aug 28 10:05:36 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__AND2B_M%A_N 1 3 4 6 8 10
r34 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.605
+ $Y=1.045 $X2=0.605 $Y2=1.045
r35 8 10 10.6318 $w=5.38e-07 $l=4.8e-07 $layer=LI1_cond $X=0.72 $Y=1.11 $X2=1.2
+ $Y2=1.11
r36 8 18 2.5472 $w=5.38e-07 $l=1.15e-07 $layer=LI1_cond $X=0.72 $Y=1.11
+ $X2=0.605 $Y2=1.11
r37 4 17 64.2376 $w=2.83e-07 $l=3.63731e-07 $layer=POLY_cond $X=0.725 $Y=1.36
+ $X2=0.62 $Y2=1.045
r38 4 6 428.16 $w=1.5e-07 $l=8.35e-07 $layer=POLY_cond $X=0.725 $Y=1.36
+ $X2=0.725 $Y2=2.195
r39 1 17 38.6899 $w=2.83e-07 $l=2.11069e-07 $layer=POLY_cond $X=0.515 $Y=0.88
+ $X2=0.62 $Y2=1.045
r40 1 3 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.515 $Y=0.88
+ $X2=0.515 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_LP__AND2B_M%A_35_70# 1 2 11 13 14 15 17 19 21 24 25 27
+ 29 32 35 37
c62 24 0 1.77961e-19 $X=1.175 $Y=1.66
c63 13 0 4.76071e-20 $X=1.54 $Y=0.84
r64 32 34 9.38152 $w=2.13e-07 $l=1.65e-07 $layer=LI1_cond $X=0.277 $Y=0.495
+ $X2=0.277 $Y2=0.66
r65 27 29 8.97835 $w=2.08e-07 $l=1.7e-07 $layer=LI1_cond $X=0.34 $Y=2.13
+ $X2=0.51 $Y2=2.13
r66 25 38 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.175 $Y=1.66
+ $X2=1.175 $Y2=1.825
r67 25 37 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.175 $Y=1.66
+ $X2=1.175 $Y2=1.495
r68 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.175
+ $Y=1.66 $X2=1.175 $Y2=1.66
r69 22 35 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.34 $Y=1.66
+ $X2=0.255 $Y2=1.66
r70 22 24 54.4759 $w=1.68e-07 $l=8.35e-07 $layer=LI1_cond $X=0.34 $Y=1.66
+ $X2=1.175 $Y2=1.66
r71 21 27 6.91519 $w=2.1e-07 $l=1.41244e-07 $layer=LI1_cond $X=0.255 $Y=2.025
+ $X2=0.34 $Y2=2.13
r72 20 35 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.255 $Y=1.745
+ $X2=0.255 $Y2=1.66
r73 20 21 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=0.255 $Y=1.745
+ $X2=0.255 $Y2=2.025
r74 19 35 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.255 $Y=1.575
+ $X2=0.255 $Y2=1.66
r75 19 34 59.6952 $w=1.68e-07 $l=9.15e-07 $layer=LI1_cond $X=0.255 $Y=1.575
+ $X2=0.255 $Y2=0.66
r76 15 17 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.615 $Y=0.765
+ $X2=1.615 $Y2=0.445
r77 13 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.54 $Y=0.84
+ $X2=1.615 $Y2=0.765
r78 13 14 102.553 $w=1.5e-07 $l=2e-07 $layer=POLY_cond $X=1.54 $Y=0.84 $X2=1.34
+ $Y2=0.84
r79 11 38 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=1.265 $Y=2.195
+ $X2=1.265 $Y2=1.825
r80 7 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.265 $Y=0.915
+ $X2=1.34 $Y2=0.84
r81 7 37 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=1.265 $Y=0.915
+ $X2=1.265 $Y2=1.495
r82 2 29 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.385
+ $Y=1.985 $X2=0.51 $Y2=2.13
r83 1 32 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.175
+ $Y=0.35 $X2=0.3 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__AND2B_M%B 3 7 9 10 11 16
c34 16 0 2.70404e-19 $X=1.955 $Y=1.32
r35 16 19 82.9202 $w=5e-07 $l=5.05e-07 $layer=POLY_cond $X=1.87 $Y=1.32 $X2=1.87
+ $Y2=1.825
r36 16 18 46.5382 $w=5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.87 $Y=1.32 $X2=1.87
+ $Y2=1.155
r37 16 17 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.955
+ $Y=1.32 $X2=1.955 $Y2=1.32
r38 11 17 10.6025 $w=3.73e-07 $l=3.45e-07 $layer=LI1_cond $X=2.057 $Y=1.665
+ $X2=2.057 $Y2=1.32
r39 10 17 0.768295 $w=3.73e-07 $l=2.5e-08 $layer=LI1_cond $X=2.057 $Y=1.295
+ $X2=2.057 $Y2=1.32
r40 9 10 11.3708 $w=3.73e-07 $l=3.7e-07 $layer=LI1_cond $X=2.057 $Y=0.925
+ $X2=2.057 $Y2=1.295
r41 7 18 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=1.975 $Y=0.445
+ $X2=1.975 $Y2=1.155
r42 3 19 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=1.695 $Y=2.195
+ $X2=1.695 $Y2=1.825
.ends

.subckt PM_SKY130_FD_SC_LP__AND2B_M%A_255_47# 1 2 7 11 14 15 20 22 27 34
r56 32 34 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=1.66 $Y=2.94 $X2=1.66
+ $Y2=2.85
r57 26 27 0.68658 $w=2.08e-07 $l=1.3e-08 $layer=LI1_cond $X=1.592 $Y=2.26
+ $X2=1.605 $Y2=2.26
r58 24 26 5.91515 $w=2.08e-07 $l=1.12e-07 $layer=LI1_cond $X=1.48 $Y=2.26
+ $X2=1.592 $Y2=2.26
r59 22 27 1.9771 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.605 $Y=2.155
+ $X2=1.605 $Y2=2.26
r60 21 22 100.471 $w=1.68e-07 $l=1.54e-06 $layer=LI1_cond $X=1.605 $Y=0.615
+ $X2=1.605 $Y2=2.155
r61 20 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.66
+ $Y=2.94 $X2=1.66 $Y2=2.94
r62 19 26 1.19342 $w=1.95e-07 $l=1.05e-07 $layer=LI1_cond $X=1.592 $Y=2.365
+ $X2=1.592 $Y2=2.26
r63 19 20 27.8695 $w=1.93e-07 $l=4.9e-07 $layer=LI1_cond $X=1.592 $Y=2.365
+ $X2=1.592 $Y2=2.855
r64 15 21 6.91519 $w=2.1e-07 $l=1.41244e-07 $layer=LI1_cond $X=1.52 $Y=0.51
+ $X2=1.605 $Y2=0.615
r65 15 17 6.33766 $w=2.08e-07 $l=1.2e-07 $layer=LI1_cond $X=1.52 $Y=0.51 $X2=1.4
+ $Y2=0.51
r66 11 14 897.34 $w=1.5e-07 $l=1.75e-06 $layer=POLY_cond $X=2.405 $Y=0.445
+ $X2=2.405 $Y2=2.195
r67 9 14 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=2.405 $Y=2.775
+ $X2=2.405 $Y2=2.195
r68 8 34 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.825 $Y=2.85
+ $X2=1.66 $Y2=2.85
r69 7 9 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.33 $Y=2.85
+ $X2=2.405 $Y2=2.775
r70 7 8 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=2.33 $Y=2.85
+ $X2=1.825 $Y2=2.85
r71 2 24 600 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=1 $X=1.34
+ $Y=1.985 $X2=1.48 $Y2=2.26
r72 1 17 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=1.275
+ $Y=0.235 $X2=1.4 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_LP__AND2B_M%VPWR 1 2 9 13 16 17 18 24 30 31 34
r37 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r38 31 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r39 30 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r40 28 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.335 $Y=3.33
+ $X2=2.17 $Y2=3.33
r41 28 30 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.335 $Y=3.33
+ $X2=2.64 $Y2=3.33
r42 27 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r43 26 27 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r44 24 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.005 $Y=3.33
+ $X2=2.17 $Y2=3.33
r45 24 26 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=2.005 $Y=3.33
+ $X2=1.68 $Y2=3.33
r46 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r47 18 27 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=1.68 $Y2=3.33
r48 18 22 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=0.72 $Y2=3.33
r49 16 21 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=0.855 $Y=3.33
+ $X2=0.72 $Y2=3.33
r50 16 17 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=0.855 $Y=3.33
+ $X2=0.96 $Y2=3.33
r51 15 26 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=1.065 $Y=3.33
+ $X2=1.68 $Y2=3.33
r52 15 17 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.065 $Y=3.33
+ $X2=0.96 $Y2=3.33
r53 11 34 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.17 $Y=3.245
+ $X2=2.17 $Y2=3.33
r54 11 13 34.3987 $w=3.28e-07 $l=9.85e-07 $layer=LI1_cond $X=2.17 $Y=3.245
+ $X2=2.17 $Y2=2.26
r55 7 17 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=0.96 $Y=3.245
+ $X2=0.96 $Y2=3.33
r56 7 9 52.0216 $w=2.08e-07 $l=9.85e-07 $layer=LI1_cond $X=0.96 $Y=3.245
+ $X2=0.96 $Y2=2.26
r57 2 13 600 $w=1.7e-07 $l=5.19615e-07 $layer=licon1_PDIFF $count=1 $X=1.77
+ $Y=1.985 $X2=2.17 $Y2=2.26
r58 1 9 600 $w=1.7e-07 $l=3.45868e-07 $layer=licon1_PDIFF $count=1 $X=0.8
+ $Y=1.985 $X2=0.96 $Y2=2.26
.ends

.subckt PM_SKY130_FD_SC_LP__AND2B_M%X 1 2 7 8 9 10 11 12 13
r10 12 13 19.5411 $w=2.08e-07 $l=3.7e-07 $layer=LI1_cond $X=2.62 $Y=2.405
+ $X2=2.62 $Y2=2.775
r11 12 34 14.5238 $w=2.08e-07 $l=2.75e-07 $layer=LI1_cond $X=2.62 $Y=2.405
+ $X2=2.62 $Y2=2.13
r12 11 34 5.01732 $w=2.08e-07 $l=9.5e-08 $layer=LI1_cond $X=2.62 $Y=2.035
+ $X2=2.62 $Y2=2.13
r13 10 11 19.5411 $w=2.08e-07 $l=3.7e-07 $layer=LI1_cond $X=2.62 $Y=1.665
+ $X2=2.62 $Y2=2.035
r14 9 10 19.5411 $w=2.08e-07 $l=3.7e-07 $layer=LI1_cond $X=2.62 $Y=1.295
+ $X2=2.62 $Y2=1.665
r15 8 9 19.5411 $w=2.08e-07 $l=3.7e-07 $layer=LI1_cond $X=2.62 $Y=0.925 $X2=2.62
+ $Y2=1.295
r16 7 8 21.9177 $w=2.08e-07 $l=4.15e-07 $layer=LI1_cond $X=2.62 $Y=0.51 $X2=2.62
+ $Y2=0.925
r17 2 34 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.48
+ $Y=1.985 $X2=2.62 $Y2=2.13
r18 1 7 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=2.48
+ $Y=0.235 $X2=2.62 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_LP__AND2B_M%VGND 1 2 9 13 15 17 22 29 30 33 36
c38 22 0 4.76071e-20 $X=2.085 $Y=0
c39 13 0 9.24432e-20 $X=2.19 $Y=0.38
r40 36 37 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r41 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r42 30 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=2.16
+ $Y2=0
r43 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r44 27 36 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.275 $Y=0 $X2=2.18
+ $Y2=0
r45 27 29 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=2.275 $Y=0 $X2=2.64
+ $Y2=0
r46 26 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r47 25 26 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r48 23 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.895 $Y=0 $X2=0.73
+ $Y2=0
r49 23 25 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.895 $Y=0 $X2=1.2
+ $Y2=0
r50 22 36 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.085 $Y=0 $X2=2.18
+ $Y2=0
r51 22 25 57.738 $w=1.68e-07 $l=8.85e-07 $layer=LI1_cond $X=2.085 $Y=0 $X2=1.2
+ $Y2=0
r52 20 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r53 19 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r54 17 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.565 $Y=0 $X2=0.73
+ $Y2=0
r55 17 19 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.565 $Y=0 $X2=0.24
+ $Y2=0
r56 15 37 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=2.16
+ $Y2=0
r57 15 26 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=1.2
+ $Y2=0
r58 11 36 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=2.18 $Y=0.085
+ $X2=2.18 $Y2=0
r59 11 13 17.2201 $w=1.88e-07 $l=2.95e-07 $layer=LI1_cond $X=2.18 $Y=0.085
+ $X2=2.18 $Y2=0.38
r60 7 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=0.085 $X2=0.73
+ $Y2=0
r61 7 9 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=0.73 $Y=0.085 $X2=0.73
+ $Y2=0.495
r62 2 13 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=2.05
+ $Y=0.235 $X2=2.19 $Y2=0.38
r63 1 9 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=0.59
+ $Y=0.35 $X2=0.73 $Y2=0.495
.ends

