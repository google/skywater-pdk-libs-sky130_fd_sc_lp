* File: sky130_fd_sc_lp__o31ai_2.pxi.spice
* Created: Wed Sep  2 10:25:21 2020
* 
x_PM_SKY130_FD_SC_LP__O31AI_2%A1 N_A1_M1002_g N_A1_c_74_n N_A1_M1000_g
+ N_A1_M1009_g N_A1_c_76_n N_A1_M1010_g A1 A1 A1 N_A1_c_78_n
+ PM_SKY130_FD_SC_LP__O31AI_2%A1
x_PM_SKY130_FD_SC_LP__O31AI_2%A2 N_A2_M1004_g N_A2_c_124_n N_A2_M1003_g
+ N_A2_M1015_g N_A2_c_126_n N_A2_M1014_g N_A2_c_127_n N_A2_c_128_n A2 A2
+ PM_SKY130_FD_SC_LP__O31AI_2%A2
x_PM_SKY130_FD_SC_LP__O31AI_2%A3 N_A3_M1008_g N_A3_M1005_g N_A3_M1013_g
+ N_A3_M1006_g A3 N_A3_c_181_n N_A3_c_185_n PM_SKY130_FD_SC_LP__O31AI_2%A3
x_PM_SKY130_FD_SC_LP__O31AI_2%B1 N_B1_c_235_n N_B1_M1001_g N_B1_M1007_g
+ N_B1_c_236_n N_B1_M1011_g N_B1_M1012_g B1 N_B1_c_238_n N_B1_c_248_n
+ PM_SKY130_FD_SC_LP__O31AI_2%B1
x_PM_SKY130_FD_SC_LP__O31AI_2%A_44_367# N_A_44_367#_M1002_s N_A_44_367#_M1009_s
+ N_A_44_367#_M1015_s N_A_44_367#_c_279_n N_A_44_367#_c_280_n
+ N_A_44_367#_c_281_n N_A_44_367#_c_294_n N_A_44_367#_c_282_n
+ N_A_44_367#_c_283_n N_A_44_367#_c_284_n PM_SKY130_FD_SC_LP__O31AI_2%A_44_367#
x_PM_SKY130_FD_SC_LP__O31AI_2%VPWR N_VPWR_M1002_d N_VPWR_M1007_s N_VPWR_c_331_n
+ N_VPWR_c_332_n VPWR N_VPWR_c_333_n N_VPWR_c_334_n N_VPWR_c_330_n
+ N_VPWR_c_336_n N_VPWR_c_337_n PM_SKY130_FD_SC_LP__O31AI_2%VPWR
x_PM_SKY130_FD_SC_LP__O31AI_2%A_299_367# N_A_299_367#_M1004_d
+ N_A_299_367#_M1005_d N_A_299_367#_c_392_n N_A_299_367#_c_387_n
+ N_A_299_367#_c_383_n N_A_299_367#_c_399_p
+ PM_SKY130_FD_SC_LP__O31AI_2%A_299_367#
x_PM_SKY130_FD_SC_LP__O31AI_2%Y N_Y_M1001_s N_Y_M1005_s N_Y_M1006_s N_Y_M1012_d
+ N_Y_c_400_n N_Y_c_401_n N_Y_c_419_n N_Y_c_403_n N_Y_c_404_n Y Y Y N_Y_c_423_n
+ N_Y_c_459_n N_Y_c_407_n N_Y_c_402_n PM_SKY130_FD_SC_LP__O31AI_2%Y
x_PM_SKY130_FD_SC_LP__O31AI_2%A_58_65# N_A_58_65#_M1000_d N_A_58_65#_M1010_d
+ N_A_58_65#_M1014_s N_A_58_65#_M1013_s N_A_58_65#_M1011_d N_A_58_65#_c_473_n
+ N_A_58_65#_c_474_n N_A_58_65#_c_483_n N_A_58_65#_c_475_n N_A_58_65#_c_490_n
+ N_A_58_65#_c_476_n N_A_58_65#_c_498_n N_A_58_65#_c_511_n N_A_58_65#_c_477_n
+ N_A_58_65#_c_478_n N_A_58_65#_c_479_n N_A_58_65#_c_488_n N_A_58_65#_c_496_n
+ PM_SKY130_FD_SC_LP__O31AI_2%A_58_65#
x_PM_SKY130_FD_SC_LP__O31AI_2%VGND N_VGND_M1000_s N_VGND_M1003_d N_VGND_M1008_d
+ N_VGND_c_540_n N_VGND_c_541_n N_VGND_c_542_n VGND N_VGND_c_543_n
+ N_VGND_c_544_n N_VGND_c_545_n N_VGND_c_546_n N_VGND_c_547_n N_VGND_c_548_n
+ N_VGND_c_549_n PM_SKY130_FD_SC_LP__O31AI_2%VGND
cc_1 VNB N_A1_M1002_g 0.00394324f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=2.465
cc_2 VNB N_A1_c_74_n 0.021262f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.275
cc_3 VNB N_A1_M1009_g 0.00257528f $X=-0.19 $Y=-0.245 $X2=0.99 $Y2=2.465
cc_4 VNB N_A1_c_76_n 0.0160346f $X=-0.19 $Y=-0.245 $X2=1.06 $Y2=1.275
cc_5 VNB A1 0.0295303f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.21
cc_6 VNB N_A1_c_78_n 0.0569008f $X=-0.19 $Y=-0.245 $X2=1.06 $Y2=1.44
cc_7 VNB N_A2_M1004_g 0.00257528f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=2.465
cc_8 VNB N_A2_c_124_n 0.0196555f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.275
cc_9 VNB N_A2_M1015_g 0.00394324f $X=-0.19 $Y=-0.245 $X2=0.99 $Y2=2.465
cc_10 VNB N_A2_c_126_n 0.0194178f $X=-0.19 $Y=-0.245 $X2=1.06 $Y2=1.275
cc_11 VNB N_A2_c_127_n 0.0379833f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_12 VNB N_A2_c_128_n 0.0482166f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB A2 0.00649944f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.44
cc_14 VNB N_A3_M1008_g 0.0184779f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=2.465
cc_15 VNB N_A3_M1013_g 0.0202442f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A3_c_181_n 0.0402093f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.44
cc_17 VNB N_B1_c_235_n 0.0162438f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=1.605
cc_18 VNB N_B1_c_236_n 0.0198728f $X=-0.19 $Y=-0.245 $X2=0.99 $Y2=1.605
cc_19 VNB B1 0.0268654f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_B1_c_238_n 0.0767573f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.44
cc_21 VNB N_VPWR_c_330_n 0.203486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_Y_c_400_n 0.0141385f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_23 VNB N_Y_c_401_n 8.5472e-19 $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_24 VNB N_Y_c_402_n 0.00598491f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_58_65#_c_473_n 0.0075508f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_26 VNB N_A_58_65#_c_474_n 0.0230663f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_58_65#_c_475_n 0.00202603f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_58_65#_c_476_n 0.00208925f $X=-0.19 $Y=-0.245 $X2=0.99 $Y2=1.44
cc_29 VNB N_A_58_65#_c_477_n 0.0119082f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_58_65#_c_478_n 0.00259911f $X=-0.19 $Y=-0.245 $X2=0.97 $Y2=1.367
cc_31 VNB N_A_58_65#_c_479_n 0.0233568f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_540_n 0.00232955f $X=-0.19 $Y=-0.245 $X2=1.06 $Y2=0.745
cc_33 VNB N_VGND_c_541_n 0.00915907f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_542_n 0.00239616f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.44
cc_35 VNB N_VGND_c_543_n 0.0157131f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.44
cc_36 VNB N_VGND_c_544_n 0.0166912f $X=-0.19 $Y=-0.245 $X2=1.06 $Y2=1.44
cc_37 VNB N_VGND_c_545_n 0.0421193f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_546_n 0.282962f $X=-0.19 $Y=-0.245 $X2=0.97 $Y2=1.367
cc_39 VNB N_VGND_c_547_n 0.0266626f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_548_n 0.0114447f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_549_n 0.00546567f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VPB N_A1_M1002_g 0.0245735f $X=-0.19 $Y=1.655 $X2=0.56 $Y2=2.465
cc_43 VPB N_A1_M1009_g 0.0187384f $X=-0.19 $Y=1.655 $X2=0.99 $Y2=2.465
cc_44 VPB N_A2_M1004_g 0.0187384f $X=-0.19 $Y=1.655 $X2=0.56 $Y2=2.465
cc_45 VPB N_A2_M1015_g 0.0245735f $X=-0.19 $Y=1.655 $X2=0.99 $Y2=2.465
cc_46 VPB N_A3_M1005_g 0.023966f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=0.745
cc_47 VPB N_A3_M1006_g 0.0206484f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_48 VPB N_A3_c_181_n 0.00817398f $X=-0.19 $Y=1.655 $X2=0.54 $Y2=1.44
cc_49 VPB N_A3_c_185_n 0.0036462f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_50 VPB N_B1_M1007_g 0.0200972f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=0.745
cc_51 VPB N_B1_M1012_g 0.0248653f $X=-0.19 $Y=1.655 $X2=1.06 $Y2=0.745
cc_52 VPB N_B1_c_238_n 0.00898331f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=1.44
cc_53 VPB N_A_44_367#_c_279_n 0.0470856f $X=-0.19 $Y=1.655 $X2=1.06 $Y2=1.275
cc_54 VPB N_A_44_367#_c_280_n 0.00223696f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_55 VPB N_A_44_367#_c_281_n 0.0100658f $X=-0.19 $Y=1.655 $X2=1.115 $Y2=1.21
cc_56 VPB N_A_44_367#_c_282_n 0.0063518f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_57 VPB N_A_44_367#_c_283_n 0.0080533f $X=-0.19 $Y=1.655 $X2=0.97 $Y2=1.44
cc_58 VPB N_A_44_367#_c_284_n 0.00285383f $X=-0.19 $Y=1.655 $X2=0.99 $Y2=1.44
cc_59 VPB N_VPWR_c_331_n 0.00474108f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_60 VPB N_VPWR_c_332_n 4.89148e-19 $X=-0.19 $Y=1.655 $X2=1.115 $Y2=1.21
cc_61 VPB N_VPWR_c_333_n 0.0743549f $X=-0.19 $Y=1.655 $X2=0.54 $Y2=1.44
cc_62 VPB N_VPWR_c_334_n 0.0153759f $X=-0.19 $Y=1.655 $X2=0.24 $Y2=1.367
cc_63 VPB N_VPWR_c_330_n 0.0510684f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_64 VPB N_VPWR_c_336_n 0.0241944f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=1.367
cc_65 VPB N_VPWR_c_337_n 0.00436868f $X=-0.19 $Y=1.655 $X2=1.2 $Y2=1.367
cc_66 VPB N_A_299_367#_c_383_n 0.0108867f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_67 VPB N_Y_c_403_n 0.0121034f $X=-0.19 $Y=1.655 $X2=0.54 $Y2=1.44
cc_68 VPB N_Y_c_404_n 0.0435297f $X=-0.19 $Y=1.655 $X2=0.56 $Y2=1.44
cc_69 VPB Y 0.00593029f $X=-0.19 $Y=1.655 $X2=0.97 $Y2=1.44
cc_70 VPB Y 0.00236249f $X=-0.19 $Y=1.655 $X2=1.06 $Y2=1.44
cc_71 VPB N_Y_c_407_n 0.0126606f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_72 VPB N_Y_c_402_n 0.00301911f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_73 N_A1_M1009_g N_A2_M1004_g 0.0241183f $X=0.99 $Y=2.465 $X2=0 $Y2=0
cc_74 N_A1_c_76_n N_A2_c_124_n 0.0143218f $X=1.06 $Y=1.275 $X2=0 $Y2=0
cc_75 A1 N_A2_c_124_n 4.38371e-19 $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_76 A1 N_A2_c_127_n 0.00209436f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_77 N_A1_c_78_n N_A2_c_127_n 0.0231268f $X=1.06 $Y=1.44 $X2=0 $Y2=0
cc_78 N_A1_c_76_n A2 2.52514e-19 $X=1.06 $Y=1.275 $X2=0 $Y2=0
cc_79 A1 A2 0.0278597f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_80 N_A1_M1002_g N_A_44_367#_c_279_n 0.0166971f $X=0.56 $Y=2.465 $X2=0 $Y2=0
cc_81 N_A1_M1009_g N_A_44_367#_c_279_n 7.29074e-19 $X=0.99 $Y=2.465 $X2=0 $Y2=0
cc_82 N_A1_M1002_g N_A_44_367#_c_280_n 0.01115f $X=0.56 $Y=2.465 $X2=0 $Y2=0
cc_83 N_A1_M1009_g N_A_44_367#_c_280_n 0.01115f $X=0.99 $Y=2.465 $X2=0 $Y2=0
cc_84 A1 N_A_44_367#_c_280_n 0.0386902f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_85 N_A1_c_78_n N_A_44_367#_c_280_n 0.00276559f $X=1.06 $Y=1.44 $X2=0 $Y2=0
cc_86 N_A1_M1002_g N_A_44_367#_c_281_n 0.00356805f $X=0.56 $Y=2.465 $X2=0 $Y2=0
cc_87 A1 N_A_44_367#_c_281_n 0.0284279f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_88 N_A1_c_78_n N_A_44_367#_c_281_n 0.00282435f $X=1.06 $Y=1.44 $X2=0 $Y2=0
cc_89 N_A1_M1002_g N_A_44_367#_c_294_n 7.29074e-19 $X=0.56 $Y=2.465 $X2=0 $Y2=0
cc_90 N_A1_M1009_g N_A_44_367#_c_294_n 0.0154189f $X=0.99 $Y=2.465 $X2=0 $Y2=0
cc_91 N_A1_M1009_g N_A_44_367#_c_284_n 0.00238146f $X=0.99 $Y=2.465 $X2=0 $Y2=0
cc_92 A1 N_A_44_367#_c_284_n 0.0210981f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_93 N_A1_c_78_n N_A_44_367#_c_284_n 0.00209851f $X=1.06 $Y=1.44 $X2=0 $Y2=0
cc_94 N_A1_M1002_g N_VPWR_c_331_n 0.00288887f $X=0.56 $Y=2.465 $X2=0 $Y2=0
cc_95 N_A1_M1009_g N_VPWR_c_331_n 0.00288887f $X=0.99 $Y=2.465 $X2=0 $Y2=0
cc_96 N_A1_M1009_g N_VPWR_c_333_n 0.0054895f $X=0.99 $Y=2.465 $X2=0 $Y2=0
cc_97 N_A1_M1002_g N_VPWR_c_330_n 0.0107693f $X=0.56 $Y=2.465 $X2=0 $Y2=0
cc_98 N_A1_M1009_g N_VPWR_c_330_n 0.00979102f $X=0.99 $Y=2.465 $X2=0 $Y2=0
cc_99 N_A1_M1002_g N_VPWR_c_336_n 0.0054895f $X=0.56 $Y=2.465 $X2=0 $Y2=0
cc_100 A1 N_A_58_65#_c_473_n 0.0219955f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_101 N_A1_c_78_n N_A_58_65#_c_473_n 8.68713e-19 $X=1.06 $Y=1.44 $X2=0 $Y2=0
cc_102 N_A1_c_74_n N_A_58_65#_c_474_n 0.00186805f $X=0.63 $Y=1.275 $X2=0 $Y2=0
cc_103 N_A1_c_74_n N_A_58_65#_c_483_n 0.0120955f $X=0.63 $Y=1.275 $X2=0 $Y2=0
cc_104 N_A1_c_76_n N_A_58_65#_c_483_n 0.0120955f $X=1.06 $Y=1.275 $X2=0 $Y2=0
cc_105 A1 N_A_58_65#_c_483_n 0.0426015f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_106 N_A1_c_78_n N_A_58_65#_c_483_n 5.87177e-19 $X=1.06 $Y=1.44 $X2=0 $Y2=0
cc_107 N_A1_c_76_n N_A_58_65#_c_475_n 4.35595e-19 $X=1.06 $Y=1.275 $X2=0 $Y2=0
cc_108 A1 N_A_58_65#_c_488_n 0.00853317f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_109 N_A1_c_74_n N_VGND_c_540_n 0.0112436f $X=0.63 $Y=1.275 $X2=0 $Y2=0
cc_110 N_A1_c_76_n N_VGND_c_540_n 0.00887263f $X=1.06 $Y=1.275 $X2=0 $Y2=0
cc_111 N_A1_c_76_n N_VGND_c_543_n 0.00414769f $X=1.06 $Y=1.275 $X2=0 $Y2=0
cc_112 N_A1_c_74_n N_VGND_c_546_n 0.00827884f $X=0.63 $Y=1.275 $X2=0 $Y2=0
cc_113 N_A1_c_76_n N_VGND_c_546_n 0.0078848f $X=1.06 $Y=1.275 $X2=0 $Y2=0
cc_114 N_A1_c_74_n N_VGND_c_547_n 0.00414769f $X=0.63 $Y=1.275 $X2=0 $Y2=0
cc_115 N_A2_c_126_n N_A3_M1008_g 0.0135452f $X=2.34 $Y=1.275 $X2=0 $Y2=0
cc_116 A2 N_A3_M1008_g 2.90819e-19 $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_117 N_A2_c_128_n N_A3_c_181_n 0.0180412f $X=2.265 $Y=1.44 $X2=0 $Y2=0
cc_118 N_A2_M1004_g N_A_44_367#_c_294_n 0.0153991f $X=1.42 $Y=2.465 $X2=0 $Y2=0
cc_119 N_A2_M1015_g N_A_44_367#_c_294_n 6.81261e-19 $X=1.85 $Y=2.465 $X2=0 $Y2=0
cc_120 N_A2_M1004_g N_A_44_367#_c_282_n 0.0122341f $X=1.42 $Y=2.465 $X2=0 $Y2=0
cc_121 N_A2_M1015_g N_A_44_367#_c_282_n 0.0147181f $X=1.85 $Y=2.465 $X2=0 $Y2=0
cc_122 N_A2_c_127_n N_A_44_367#_c_282_n 0.00276559f $X=1.925 $Y=1.44 $X2=0 $Y2=0
cc_123 N_A2_c_128_n N_A_44_367#_c_282_n 0.00804572f $X=2.265 $Y=1.44 $X2=0 $Y2=0
cc_124 A2 N_A_44_367#_c_282_n 0.0602653f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_125 N_A2_M1004_g N_A_44_367#_c_283_n 6.32885e-19 $X=1.42 $Y=2.465 $X2=0 $Y2=0
cc_126 N_A2_M1015_g N_A_44_367#_c_283_n 0.0152181f $X=1.85 $Y=2.465 $X2=0 $Y2=0
cc_127 N_A2_M1004_g N_A_44_367#_c_284_n 0.00263866f $X=1.42 $Y=2.465 $X2=0 $Y2=0
cc_128 N_A2_M1004_g N_VPWR_c_333_n 0.0054895f $X=1.42 $Y=2.465 $X2=0 $Y2=0
cc_129 N_A2_M1015_g N_VPWR_c_333_n 0.00357877f $X=1.85 $Y=2.465 $X2=0 $Y2=0
cc_130 N_A2_M1004_g N_VPWR_c_330_n 0.0099382f $X=1.42 $Y=2.465 $X2=0 $Y2=0
cc_131 N_A2_M1015_g N_VPWR_c_330_n 0.00675087f $X=1.85 $Y=2.465 $X2=0 $Y2=0
cc_132 N_A2_M1015_g N_A_299_367#_c_383_n 0.0135436f $X=1.85 $Y=2.465 $X2=0 $Y2=0
cc_133 N_A2_c_126_n N_Y_c_401_n 0.00163626f $X=2.34 $Y=1.275 $X2=0 $Y2=0
cc_134 A2 N_Y_c_401_n 0.00156421f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_135 N_A2_M1015_g Y 0.00151539f $X=1.85 $Y=2.465 $X2=0 $Y2=0
cc_136 N_A2_M1015_g N_Y_c_407_n 5.51873e-19 $X=1.85 $Y=2.465 $X2=0 $Y2=0
cc_137 N_A2_c_126_n N_Y_c_402_n 0.00379037f $X=2.34 $Y=1.275 $X2=0 $Y2=0
cc_138 A2 N_Y_c_402_n 0.0114342f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_139 N_A2_c_124_n N_A_58_65#_c_475_n 4.73912e-19 $X=1.49 $Y=1.275 $X2=0 $Y2=0
cc_140 N_A2_c_124_n N_A_58_65#_c_490_n 0.0149296f $X=1.49 $Y=1.275 $X2=0 $Y2=0
cc_141 N_A2_c_126_n N_A_58_65#_c_490_n 0.0112498f $X=2.34 $Y=1.275 $X2=0 $Y2=0
cc_142 N_A2_c_127_n N_A_58_65#_c_490_n 0.00305891f $X=1.925 $Y=1.44 $X2=0 $Y2=0
cc_143 A2 N_A_58_65#_c_490_n 0.0587587f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_144 N_A2_c_126_n N_A_58_65#_c_476_n 0.00816228f $X=2.34 $Y=1.275 $X2=0 $Y2=0
cc_145 N_A2_c_127_n N_A_58_65#_c_488_n 0.0015791f $X=1.925 $Y=1.44 $X2=0 $Y2=0
cc_146 N_A2_c_126_n N_A_58_65#_c_496_n 0.0115511f $X=2.34 $Y=1.275 $X2=0 $Y2=0
cc_147 N_A2_c_124_n N_VGND_c_540_n 4.87122e-19 $X=1.49 $Y=1.275 $X2=0 $Y2=0
cc_148 N_A2_c_124_n N_VGND_c_541_n 0.00258596f $X=1.49 $Y=1.275 $X2=0 $Y2=0
cc_149 N_A2_c_126_n N_VGND_c_541_n 0.00338144f $X=2.34 $Y=1.275 $X2=0 $Y2=0
cc_150 N_A2_c_126_n N_VGND_c_542_n 3.99488e-19 $X=2.34 $Y=1.275 $X2=0 $Y2=0
cc_151 N_A2_c_124_n N_VGND_c_543_n 0.00499542f $X=1.49 $Y=1.275 $X2=0 $Y2=0
cc_152 N_A2_c_126_n N_VGND_c_544_n 0.00411073f $X=2.34 $Y=1.275 $X2=0 $Y2=0
cc_153 N_A2_c_124_n N_VGND_c_546_n 0.0100168f $X=1.49 $Y=1.275 $X2=0 $Y2=0
cc_154 N_A2_c_126_n N_VGND_c_546_n 0.00763133f $X=2.34 $Y=1.275 $X2=0 $Y2=0
cc_155 N_A3_M1013_g N_B1_c_235_n 0.0267591f $X=3.2 $Y=0.745 $X2=-0.19 $Y2=-0.245
cc_156 N_A3_M1006_g N_B1_M1007_g 0.020306f $X=3.31 $Y=2.465 $X2=0 $Y2=0
cc_157 N_A3_c_181_n N_B1_M1007_g 3.38109e-19 $X=3.25 $Y=1.51 $X2=0 $Y2=0
cc_158 N_A3_c_185_n N_B1_M1007_g 0.00161173f $X=3.25 $Y=1.51 $X2=0 $Y2=0
cc_159 N_A3_c_181_n N_B1_c_238_n 0.0236844f $X=3.25 $Y=1.51 $X2=0 $Y2=0
cc_160 N_A3_c_185_n N_B1_c_238_n 0.00127153f $X=3.25 $Y=1.51 $X2=0 $Y2=0
cc_161 N_A3_c_181_n N_B1_c_248_n 6.8386e-19 $X=3.25 $Y=1.51 $X2=0 $Y2=0
cc_162 N_A3_c_185_n N_B1_c_248_n 0.0100581f $X=3.25 $Y=1.51 $X2=0 $Y2=0
cc_163 N_A3_M1005_g N_A_44_367#_c_282_n 9.23481e-19 $X=2.8 $Y=2.465 $X2=0 $Y2=0
cc_164 N_A3_M1005_g N_A_44_367#_c_283_n 0.00151145f $X=2.8 $Y=2.465 $X2=0 $Y2=0
cc_165 N_A3_M1006_g N_VPWR_c_332_n 0.00106288f $X=3.31 $Y=2.465 $X2=0 $Y2=0
cc_166 N_A3_M1005_g N_VPWR_c_333_n 0.00357877f $X=2.8 $Y=2.465 $X2=0 $Y2=0
cc_167 N_A3_M1006_g N_VPWR_c_333_n 0.00585385f $X=3.31 $Y=2.465 $X2=0 $Y2=0
cc_168 N_A3_M1005_g N_VPWR_c_330_n 0.00694461f $X=2.8 $Y=2.465 $X2=0 $Y2=0
cc_169 N_A3_M1006_g N_VPWR_c_330_n 0.0114351f $X=3.31 $Y=2.465 $X2=0 $Y2=0
cc_170 N_A3_M1005_g N_A_299_367#_c_383_n 0.0135141f $X=2.8 $Y=2.465 $X2=0 $Y2=0
cc_171 N_A3_M1013_g N_Y_c_400_n 0.0108338f $X=3.2 $Y=0.745 $X2=0 $Y2=0
cc_172 N_A3_c_181_n N_Y_c_400_n 0.00809154f $X=3.25 $Y=1.51 $X2=0 $Y2=0
cc_173 N_A3_c_185_n N_Y_c_400_n 0.026773f $X=3.25 $Y=1.51 $X2=0 $Y2=0
cc_174 N_A3_M1008_g N_Y_c_401_n 0.00714628f $X=2.77 $Y=0.745 $X2=0 $Y2=0
cc_175 N_A3_M1013_g N_Y_c_419_n 5.43466e-19 $X=3.2 $Y=0.745 $X2=0 $Y2=0
cc_176 N_A3_M1005_g Y 0.0132351f $X=2.8 $Y=2.465 $X2=0 $Y2=0
cc_177 N_A3_M1006_g Y 6.32592e-19 $X=3.31 $Y=2.465 $X2=0 $Y2=0
cc_178 N_A3_M1006_g Y 0.00430325f $X=3.31 $Y=2.465 $X2=0 $Y2=0
cc_179 N_A3_M1005_g N_Y_c_423_n 0.00558429f $X=2.8 $Y=2.465 $X2=0 $Y2=0
cc_180 N_A3_M1006_g N_Y_c_423_n 0.0142641f $X=3.31 $Y=2.465 $X2=0 $Y2=0
cc_181 N_A3_c_181_n N_Y_c_423_n 0.00310788f $X=3.25 $Y=1.51 $X2=0 $Y2=0
cc_182 N_A3_c_185_n N_Y_c_423_n 0.0256706f $X=3.25 $Y=1.51 $X2=0 $Y2=0
cc_183 N_A3_M1005_g N_Y_c_407_n 0.0118584f $X=2.8 $Y=2.465 $X2=0 $Y2=0
cc_184 N_A3_M1008_g N_Y_c_402_n 0.00199979f $X=2.77 $Y=0.745 $X2=0 $Y2=0
cc_185 N_A3_M1005_g N_Y_c_402_n 0.00495785f $X=2.8 $Y=2.465 $X2=0 $Y2=0
cc_186 N_A3_M1013_g N_Y_c_402_n 0.00181541f $X=3.2 $Y=0.745 $X2=0 $Y2=0
cc_187 N_A3_M1006_g N_Y_c_402_n 0.0010438f $X=3.31 $Y=2.465 $X2=0 $Y2=0
cc_188 N_A3_c_181_n N_Y_c_402_n 0.0140758f $X=3.25 $Y=1.51 $X2=0 $Y2=0
cc_189 N_A3_c_185_n N_Y_c_402_n 0.0230728f $X=3.25 $Y=1.51 $X2=0 $Y2=0
cc_190 N_A3_M1008_g N_A_58_65#_c_476_n 2.98511e-19 $X=2.77 $Y=0.745 $X2=0 $Y2=0
cc_191 N_A3_M1008_g N_A_58_65#_c_498_n 0.00981896f $X=2.77 $Y=0.745 $X2=0 $Y2=0
cc_192 N_A3_M1013_g N_A_58_65#_c_498_n 0.00982509f $X=3.2 $Y=0.745 $X2=0 $Y2=0
cc_193 N_A3_M1013_g N_A_58_65#_c_478_n 6.37722e-19 $X=3.2 $Y=0.745 $X2=0 $Y2=0
cc_194 N_A3_M1008_g N_A_58_65#_c_496_n 0.00331298f $X=2.77 $Y=0.745 $X2=0 $Y2=0
cc_195 N_A3_M1008_g N_VGND_c_542_n 0.00669238f $X=2.77 $Y=0.745 $X2=0 $Y2=0
cc_196 N_A3_M1013_g N_VGND_c_542_n 0.00677442f $X=3.2 $Y=0.745 $X2=0 $Y2=0
cc_197 N_A3_M1008_g N_VGND_c_544_n 0.00305694f $X=2.77 $Y=0.745 $X2=0 $Y2=0
cc_198 N_A3_M1013_g N_VGND_c_545_n 0.00305694f $X=3.2 $Y=0.745 $X2=0 $Y2=0
cc_199 N_A3_M1008_g N_VGND_c_546_n 0.00392857f $X=2.77 $Y=0.745 $X2=0 $Y2=0
cc_200 N_A3_M1013_g N_VGND_c_546_n 0.00398998f $X=3.2 $Y=0.745 $X2=0 $Y2=0
cc_201 N_B1_M1007_g N_VPWR_c_332_n 0.0156484f $X=3.895 $Y=2.465 $X2=0 $Y2=0
cc_202 N_B1_M1012_g N_VPWR_c_332_n 0.0161992f $X=4.325 $Y=2.465 $X2=0 $Y2=0
cc_203 N_B1_M1007_g N_VPWR_c_333_n 0.00486043f $X=3.895 $Y=2.465 $X2=0 $Y2=0
cc_204 N_B1_M1012_g N_VPWR_c_334_n 0.00486043f $X=4.325 $Y=2.465 $X2=0 $Y2=0
cc_205 N_B1_M1007_g N_VPWR_c_330_n 0.00873567f $X=3.895 $Y=2.465 $X2=0 $Y2=0
cc_206 N_B1_M1012_g N_VPWR_c_330_n 0.00917987f $X=4.325 $Y=2.465 $X2=0 $Y2=0
cc_207 N_B1_c_235_n N_Y_c_400_n 0.0113731f $X=3.7 $Y=1.275 $X2=0 $Y2=0
cc_208 N_B1_c_236_n N_Y_c_400_n 0.00807213f $X=4.13 $Y=1.275 $X2=0 $Y2=0
cc_209 B1 N_Y_c_400_n 0.00281226f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_210 N_B1_c_238_n N_Y_c_400_n 0.00321706f $X=4.325 $Y=1.47 $X2=0 $Y2=0
cc_211 N_B1_c_248_n N_Y_c_400_n 0.0333834f $X=4.26 $Y=1.397 $X2=0 $Y2=0
cc_212 N_B1_c_235_n N_Y_c_419_n 0.00673716f $X=3.7 $Y=1.275 $X2=0 $Y2=0
cc_213 N_B1_c_236_n N_Y_c_419_n 0.00654168f $X=4.13 $Y=1.275 $X2=0 $Y2=0
cc_214 N_B1_M1007_g N_Y_c_403_n 0.0143784f $X=3.895 $Y=2.465 $X2=0 $Y2=0
cc_215 N_B1_M1012_g N_Y_c_403_n 0.0138099f $X=4.325 $Y=2.465 $X2=0 $Y2=0
cc_216 B1 N_Y_c_403_n 0.0226029f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_217 N_B1_c_238_n N_Y_c_403_n 0.00868528f $X=4.325 $Y=1.47 $X2=0 $Y2=0
cc_218 N_B1_c_248_n N_Y_c_403_n 0.0474998f $X=4.26 $Y=1.397 $X2=0 $Y2=0
cc_219 N_B1_c_238_n Y 0.00461176f $X=4.325 $Y=1.47 $X2=0 $Y2=0
cc_220 N_B1_c_248_n Y 0.0104877f $X=4.26 $Y=1.397 $X2=0 $Y2=0
cc_221 N_B1_c_235_n N_A_58_65#_c_477_n 0.0112303f $X=3.7 $Y=1.275 $X2=0 $Y2=0
cc_222 N_B1_c_236_n N_A_58_65#_c_477_n 0.0125492f $X=4.13 $Y=1.275 $X2=0 $Y2=0
cc_223 B1 N_A_58_65#_c_479_n 0.0217678f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_224 N_B1_c_238_n N_A_58_65#_c_479_n 0.00164902f $X=4.325 $Y=1.47 $X2=0 $Y2=0
cc_225 N_B1_c_235_n N_VGND_c_542_n 5.53873e-19 $X=3.7 $Y=1.275 $X2=0 $Y2=0
cc_226 N_B1_c_235_n N_VGND_c_545_n 0.00302501f $X=3.7 $Y=1.275 $X2=0 $Y2=0
cc_227 N_B1_c_236_n N_VGND_c_545_n 0.00302501f $X=4.13 $Y=1.275 $X2=0 $Y2=0
cc_228 N_B1_c_235_n N_VGND_c_546_n 0.00441786f $X=3.7 $Y=1.275 $X2=0 $Y2=0
cc_229 N_B1_c_236_n N_VGND_c_546_n 0.00475908f $X=4.13 $Y=1.275 $X2=0 $Y2=0
cc_230 N_A_44_367#_c_280_n N_VPWR_M1002_d 0.00176461f $X=1.04 $Y=1.78 $X2=-0.19
+ $Y2=1.655
cc_231 N_A_44_367#_c_280_n N_VPWR_c_331_n 0.0135055f $X=1.04 $Y=1.78 $X2=0 $Y2=0
cc_232 N_A_44_367#_c_294_n N_VPWR_c_333_n 0.0189236f $X=1.205 $Y=1.98 $X2=0
+ $Y2=0
cc_233 N_A_44_367#_M1002_s N_VPWR_c_330_n 0.00215158f $X=0.22 $Y=1.835 $X2=0
+ $Y2=0
cc_234 N_A_44_367#_M1009_s N_VPWR_c_330_n 0.00223559f $X=1.065 $Y=1.835 $X2=0
+ $Y2=0
cc_235 N_A_44_367#_M1015_s N_VPWR_c_330_n 0.0021598f $X=1.925 $Y=1.835 $X2=0
+ $Y2=0
cc_236 N_A_44_367#_c_279_n N_VPWR_c_330_n 0.0125689f $X=0.345 $Y=1.98 $X2=0
+ $Y2=0
cc_237 N_A_44_367#_c_294_n N_VPWR_c_330_n 0.0123859f $X=1.205 $Y=1.98 $X2=0
+ $Y2=0
cc_238 N_A_44_367#_c_279_n N_VPWR_c_336_n 0.0210467f $X=0.345 $Y=1.98 $X2=0
+ $Y2=0
cc_239 N_A_44_367#_c_282_n N_A_299_367#_M1004_d 0.00176461f $X=1.9 $Y=1.78
+ $X2=-0.19 $Y2=1.655
cc_240 N_A_44_367#_c_282_n N_A_299_367#_c_387_n 0.0135055f $X=1.9 $Y=1.78 $X2=0
+ $Y2=0
cc_241 N_A_44_367#_M1015_s N_A_299_367#_c_383_n 0.00495471f $X=1.925 $Y=1.835
+ $X2=0 $Y2=0
cc_242 N_A_44_367#_c_283_n N_A_299_367#_c_383_n 0.0205857f $X=2.065 $Y=1.98
+ $X2=0 $Y2=0
cc_243 N_A_44_367#_c_283_n Y 0.0473989f $X=2.065 $Y=1.98 $X2=0 $Y2=0
cc_244 N_A_44_367#_c_282_n N_Y_c_407_n 0.00417062f $X=1.9 $Y=1.78 $X2=0 $Y2=0
cc_245 N_A_44_367#_c_283_n N_Y_c_407_n 0.0200157f $X=2.065 $Y=1.98 $X2=0 $Y2=0
cc_246 N_A_44_367#_c_282_n N_Y_c_402_n 0.00509857f $X=1.9 $Y=1.78 $X2=0 $Y2=0
cc_247 N_A_44_367#_c_282_n N_A_58_65#_c_490_n 9.24293e-19 $X=1.9 $Y=1.78 $X2=0
+ $Y2=0
cc_248 N_A_44_367#_c_284_n N_A_58_65#_c_488_n 0.00261601f $X=1.205 $Y=1.78 $X2=0
+ $Y2=0
cc_249 N_VPWR_c_330_n N_A_299_367#_M1004_d 0.00376627f $X=4.56 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_250 N_VPWR_c_330_n N_A_299_367#_M1005_d 0.00480031f $X=4.56 $Y=3.33 $X2=0
+ $Y2=0
cc_251 N_VPWR_c_333_n N_A_299_367#_c_392_n 0.0125234f $X=3.945 $Y=3.33 $X2=0
+ $Y2=0
cc_252 N_VPWR_c_330_n N_A_299_367#_c_392_n 0.00738676f $X=4.56 $Y=3.33 $X2=0
+ $Y2=0
cc_253 N_VPWR_c_333_n N_A_299_367#_c_383_n 0.0871502f $X=3.945 $Y=3.33 $X2=0
+ $Y2=0
cc_254 N_VPWR_c_330_n N_A_299_367#_c_383_n 0.0533245f $X=4.56 $Y=3.33 $X2=0
+ $Y2=0
cc_255 N_VPWR_c_330_n N_Y_M1005_s 0.0021598f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_256 N_VPWR_c_330_n N_Y_M1006_s 0.00615916f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_257 N_VPWR_c_330_n N_Y_M1012_d 0.00371702f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_258 N_VPWR_M1007_s N_Y_c_403_n 0.00176461f $X=3.97 $Y=1.835 $X2=0 $Y2=0
cc_259 N_VPWR_c_332_n N_Y_c_403_n 0.0170777f $X=4.11 $Y=2.18 $X2=0 $Y2=0
cc_260 N_VPWR_c_334_n N_Y_c_404_n 0.0178111f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_261 N_VPWR_c_330_n N_Y_c_404_n 0.0100304f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_262 N_VPWR_c_333_n N_Y_c_459_n 0.0238831f $X=3.945 $Y=3.33 $X2=0 $Y2=0
cc_263 N_VPWR_c_330_n N_Y_c_459_n 0.0139182f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_264 N_A_299_367#_c_383_n N_Y_M1005_s 0.0049601f $X=2.92 $Y=2.99 $X2=0 $Y2=0
cc_265 N_A_299_367#_c_383_n Y 0.0204673f $X=2.92 $Y=2.99 $X2=0 $Y2=0
cc_266 N_A_299_367#_M1005_d N_Y_c_423_n 0.0060896f $X=2.875 $Y=1.835 $X2=0 $Y2=0
cc_267 N_A_299_367#_c_399_p N_Y_c_423_n 0.0202007f $X=3.015 $Y=2.455 $X2=0 $Y2=0
cc_268 N_Y_c_400_n N_A_58_65#_M1013_s 0.00250873f $X=3.75 $Y=1.16 $X2=0 $Y2=0
cc_269 N_Y_c_400_n N_A_58_65#_c_498_n 0.0221903f $X=3.75 $Y=1.16 $X2=0 $Y2=0
cc_270 N_Y_c_401_n N_A_58_65#_c_498_n 0.0113922f $X=2.855 $Y=1.16 $X2=0 $Y2=0
cc_271 N_Y_c_400_n N_A_58_65#_c_511_n 0.01913f $X=3.75 $Y=1.16 $X2=0 $Y2=0
cc_272 N_Y_M1001_s N_A_58_65#_c_477_n 0.00176461f $X=3.775 $Y=0.325 $X2=0 $Y2=0
cc_273 N_Y_c_400_n N_A_58_65#_c_477_n 0.00275981f $X=3.75 $Y=1.16 $X2=0 $Y2=0
cc_274 N_Y_c_419_n N_A_58_65#_c_477_n 0.0159249f $X=3.915 $Y=0.68 $X2=0 $Y2=0
cc_275 N_Y_c_400_n N_VGND_M1008_d 0.00176891f $X=3.75 $Y=1.16 $X2=0 $Y2=0
cc_276 N_A_58_65#_c_483_n N_VGND_M1000_s 0.003325f $X=1.18 $Y=0.955 $X2=-0.19
+ $Y2=-0.245
cc_277 N_A_58_65#_c_490_n N_VGND_M1003_d 0.0154783f $X=2.345 $Y=0.955 $X2=0
+ $Y2=0
cc_278 N_A_58_65#_c_498_n N_VGND_M1008_d 0.00334372f $X=3.32 $Y=0.82 $X2=0 $Y2=0
cc_279 N_A_58_65#_c_474_n N_VGND_c_540_n 0.0148073f $X=0.415 $Y=0.48 $X2=0 $Y2=0
cc_280 N_A_58_65#_c_483_n N_VGND_c_540_n 0.0170777f $X=1.18 $Y=0.955 $X2=0 $Y2=0
cc_281 N_A_58_65#_c_475_n N_VGND_c_540_n 0.0148006f $X=1.275 $Y=0.48 $X2=0 $Y2=0
cc_282 N_A_58_65#_c_475_n N_VGND_c_541_n 7.63817e-19 $X=1.275 $Y=0.48 $X2=0
+ $Y2=0
cc_283 N_A_58_65#_c_490_n N_VGND_c_541_n 0.0449099f $X=2.345 $Y=0.955 $X2=0
+ $Y2=0
cc_284 N_A_58_65#_c_476_n N_VGND_c_541_n 0.0336233f $X=2.555 $Y=0.45 $X2=0 $Y2=0
cc_285 N_A_58_65#_c_476_n N_VGND_c_542_n 0.0121096f $X=2.555 $Y=0.45 $X2=0 $Y2=0
cc_286 N_A_58_65#_c_498_n N_VGND_c_542_n 0.016459f $X=3.32 $Y=0.82 $X2=0 $Y2=0
cc_287 N_A_58_65#_c_478_n N_VGND_c_542_n 0.00962585f $X=3.58 $Y=0.34 $X2=0 $Y2=0
cc_288 N_A_58_65#_c_475_n N_VGND_c_543_n 0.0118292f $X=1.275 $Y=0.48 $X2=0 $Y2=0
cc_289 N_A_58_65#_c_476_n N_VGND_c_544_n 0.0179638f $X=2.555 $Y=0.45 $X2=0 $Y2=0
cc_290 N_A_58_65#_c_498_n N_VGND_c_544_n 0.00196209f $X=3.32 $Y=0.82 $X2=0 $Y2=0
cc_291 N_A_58_65#_c_498_n N_VGND_c_545_n 0.00196209f $X=3.32 $Y=0.82 $X2=0 $Y2=0
cc_292 N_A_58_65#_c_477_n N_VGND_c_545_n 0.0608672f $X=4.25 $Y=0.34 $X2=0 $Y2=0
cc_293 N_A_58_65#_c_478_n N_VGND_c_545_n 0.0185749f $X=3.58 $Y=0.34 $X2=0 $Y2=0
cc_294 N_A_58_65#_c_474_n N_VGND_c_546_n 0.00972454f $X=0.415 $Y=0.48 $X2=0
+ $Y2=0
cc_295 N_A_58_65#_c_475_n N_VGND_c_546_n 0.00859378f $X=1.275 $Y=0.48 $X2=0
+ $Y2=0
cc_296 N_A_58_65#_c_476_n N_VGND_c_546_n 0.0112715f $X=2.555 $Y=0.45 $X2=0 $Y2=0
cc_297 N_A_58_65#_c_498_n N_VGND_c_546_n 0.00899218f $X=3.32 $Y=0.82 $X2=0 $Y2=0
cc_298 N_A_58_65#_c_477_n N_VGND_c_546_n 0.0339255f $X=4.25 $Y=0.34 $X2=0 $Y2=0
cc_299 N_A_58_65#_c_478_n N_VGND_c_546_n 0.0100962f $X=3.58 $Y=0.34 $X2=0 $Y2=0
cc_300 N_A_58_65#_c_474_n N_VGND_c_547_n 0.0133857f $X=0.415 $Y=0.48 $X2=0 $Y2=0
