* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__and4_m A B C D VGND VNB VPB VPWR X
X0 a_136_47# B a_208_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 a_53_47# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X2 a_53_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X3 VPWR a_53_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X4 VPWR A a_53_47# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X5 a_208_47# C a_316_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 a_316_47# D VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 VPWR C a_53_47# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X8 VGND a_53_47# X VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 a_53_47# A a_136_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
