* File: sky130_fd_sc_lp__clkinv_8.pxi.spice
* Created: Fri Aug 28 10:18:09 2020
* 
x_PM_SKY130_FD_SC_LP__CLKINV_8%A N_A_M1000_g N_A_M1003_g N_A_M1001_g N_A_M1005_g
+ N_A_M1002_g N_A_M1007_g N_A_M1004_g N_A_M1008_g N_A_M1006_g N_A_M1010_g
+ N_A_M1009_g N_A_M1012_g N_A_M1011_g N_A_M1014_g N_A_M1013_g N_A_M1015_g
+ N_A_M1018_g N_A_M1016_g N_A_M1017_g N_A_M1019_g A A A A A A A A A A
+ N_A_c_126_n PM_SKY130_FD_SC_LP__CLKINV_8%A
x_PM_SKY130_FD_SC_LP__CLKINV_8%VPWR N_VPWR_M1000_s N_VPWR_M1003_s N_VPWR_M1007_s
+ N_VPWR_M1010_s N_VPWR_M1014_s N_VPWR_M1016_s N_VPWR_M1019_s N_VPWR_c_274_n
+ N_VPWR_c_275_n N_VPWR_c_276_n N_VPWR_c_277_n N_VPWR_c_278_n N_VPWR_c_279_n
+ N_VPWR_c_280_n N_VPWR_c_281_n N_VPWR_c_282_n N_VPWR_c_283_n N_VPWR_c_284_n
+ N_VPWR_c_285_n N_VPWR_c_286_n N_VPWR_c_287_n N_VPWR_c_288_n N_VPWR_c_289_n
+ VPWR N_VPWR_c_290_n N_VPWR_c_291_n N_VPWR_c_292_n N_VPWR_c_293_n
+ N_VPWR_c_273_n PM_SKY130_FD_SC_LP__CLKINV_8%VPWR
x_PM_SKY130_FD_SC_LP__CLKINV_8%Y N_Y_M1001_s N_Y_M1004_s N_Y_M1009_s N_Y_M1013_s
+ N_Y_M1000_d N_Y_M1005_d N_Y_M1008_d N_Y_M1012_d N_Y_M1015_d N_Y_M1017_d
+ N_Y_c_365_n N_Y_c_366_n N_Y_c_367_n N_Y_c_383_n N_Y_c_384_n N_Y_c_482_n
+ N_Y_c_385_n N_Y_c_368_n N_Y_c_486_n N_Y_c_369_n N_Y_c_386_n N_Y_c_370_n
+ N_Y_c_490_n N_Y_c_371_n N_Y_c_387_n N_Y_c_372_n N_Y_c_494_n N_Y_c_373_n
+ N_Y_c_388_n N_Y_c_374_n N_Y_c_498_n N_Y_c_389_n N_Y_c_502_n N_Y_c_390_n
+ N_Y_c_391_n N_Y_c_375_n N_Y_c_392_n N_Y_c_376_n N_Y_c_393_n N_Y_c_377_n
+ N_Y_c_394_n N_Y_c_378_n N_Y_c_395_n N_Y_c_396_n Y Y N_Y_c_381_n
+ PM_SKY130_FD_SC_LP__CLKINV_8%Y
x_PM_SKY130_FD_SC_LP__CLKINV_8%VGND N_VGND_M1001_d N_VGND_M1002_d N_VGND_M1006_d
+ N_VGND_M1011_d N_VGND_M1018_d N_VGND_c_526_n N_VGND_c_527_n N_VGND_c_528_n
+ N_VGND_c_529_n N_VGND_c_530_n N_VGND_c_531_n N_VGND_c_532_n N_VGND_c_533_n
+ N_VGND_c_534_n N_VGND_c_535_n N_VGND_c_536_n N_VGND_c_537_n VGND
+ N_VGND_c_538_n N_VGND_c_539_n N_VGND_c_540_n N_VGND_c_541_n N_VGND_c_542_n
+ PM_SKY130_FD_SC_LP__CLKINV_8%VGND
cc_1 VNB N_A_M1000_g 0.00628988f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=2.465
cc_2 VNB N_A_M1003_g 0.00579465f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=2.465
cc_3 VNB N_A_M1001_g 0.0432088f $X=-0.19 $Y=-0.245 $X2=1.405 $Y2=0.56
cc_4 VNB N_A_M1005_g 0.00579762f $X=-0.19 $Y=-0.245 $X2=1.405 $Y2=2.465
cc_5 VNB N_A_M1002_g 0.0320798f $X=-0.19 $Y=-0.245 $X2=1.835 $Y2=0.56
cc_6 VNB N_A_M1007_g 0.00579762f $X=-0.19 $Y=-0.245 $X2=1.835 $Y2=2.465
cc_7 VNB N_A_M1004_g 0.0320798f $X=-0.19 $Y=-0.245 $X2=2.265 $Y2=0.56
cc_8 VNB N_A_M1008_g 0.00579762f $X=-0.19 $Y=-0.245 $X2=2.265 $Y2=2.465
cc_9 VNB N_A_M1006_g 0.0320798f $X=-0.19 $Y=-0.245 $X2=2.695 $Y2=0.56
cc_10 VNB N_A_M1010_g 0.00579762f $X=-0.19 $Y=-0.245 $X2=2.695 $Y2=2.465
cc_11 VNB N_A_M1009_g 0.0320798f $X=-0.19 $Y=-0.245 $X2=3.125 $Y2=0.56
cc_12 VNB N_A_M1012_g 0.00579762f $X=-0.19 $Y=-0.245 $X2=3.125 $Y2=2.465
cc_13 VNB N_A_M1011_g 0.0320798f $X=-0.19 $Y=-0.245 $X2=3.555 $Y2=0.56
cc_14 VNB N_A_M1014_g 0.00579762f $X=-0.19 $Y=-0.245 $X2=3.555 $Y2=2.465
cc_15 VNB N_A_M1013_g 0.0320798f $X=-0.19 $Y=-0.245 $X2=3.985 $Y2=0.56
cc_16 VNB N_A_M1015_g 0.00579762f $X=-0.19 $Y=-0.245 $X2=3.985 $Y2=2.465
cc_17 VNB N_A_M1018_g 0.0432088f $X=-0.19 $Y=-0.245 $X2=4.415 $Y2=0.56
cc_18 VNB N_A_M1016_g 0.00579762f $X=-0.19 $Y=-0.245 $X2=4.415 $Y2=2.465
cc_19 VNB N_A_M1017_g 0.00579365f $X=-0.19 $Y=-0.245 $X2=4.845 $Y2=2.465
cc_20 VNB N_A_M1019_g 0.00625137f $X=-0.19 $Y=-0.245 $X2=5.275 $Y2=2.465
cc_21 VNB N_A_c_126_n 0.275358f $X=-0.19 $Y=-0.245 $X2=5.275 $Y2=1.375
cc_22 VNB N_VPWR_c_273_n 0.243291f $X=-0.19 $Y=-0.245 $X2=1.405 $Y2=1.375
cc_23 VNB N_Y_c_365_n 0.0333088f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_Y_c_366_n 0.0278014f $X=-0.19 $Y=-0.245 $X2=2.695 $Y2=1.21
cc_25 VNB N_Y_c_367_n 0.0128703f $X=-0.19 $Y=-0.245 $X2=2.695 $Y2=0.56
cc_26 VNB N_Y_c_368_n 0.00119645f $X=-0.19 $Y=-0.245 $X2=3.125 $Y2=2.465
cc_27 VNB N_Y_c_369_n 0.00538522f $X=-0.19 $Y=-0.245 $X2=3.555 $Y2=2.465
cc_28 VNB N_Y_c_370_n 0.00110053f $X=-0.19 $Y=-0.245 $X2=3.985 $Y2=1.54
cc_29 VNB N_Y_c_371_n 0.00538522f $X=-0.19 $Y=-0.245 $X2=4.415 $Y2=1.54
cc_30 VNB N_Y_c_372_n 0.00110053f $X=-0.19 $Y=-0.245 $X2=4.845 $Y2=2.465
cc_31 VNB N_Y_c_373_n 0.00538522f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.21
cc_32 VNB N_Y_c_374_n 0.00119645f $X=-0.19 $Y=-0.245 $X2=4.475 $Y2=1.21
cc_33 VNB N_Y_c_375_n 0.00205825f $X=-0.19 $Y=-0.245 $X2=1.835 $Y2=1.375
cc_34 VNB N_Y_c_376_n 0.00205825f $X=-0.19 $Y=-0.245 $X2=2.695 $Y2=1.375
cc_35 VNB N_Y_c_377_n 0.00205825f $X=-0.19 $Y=-0.245 $X2=3.555 $Y2=1.375
cc_36 VNB N_Y_c_378_n 0.00205825f $X=-0.19 $Y=-0.245 $X2=4.845 $Y2=1.375
cc_37 VNB Y 0.0263263f $X=-0.19 $Y=-0.245 $X2=5.275 $Y2=1.375
cc_38 VNB Y 0.0337179f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_Y_c_381_n 0.0132875f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=1.375
cc_40 VNB N_VGND_c_526_n 0.0235135f $X=-0.19 $Y=-0.245 $X2=1.835 $Y2=0.56
cc_41 VNB N_VGND_c_527_n 0.00698312f $X=-0.19 $Y=-0.245 $X2=1.835 $Y2=2.465
cc_42 VNB N_VGND_c_528_n 0.00698312f $X=-0.19 $Y=-0.245 $X2=2.265 $Y2=0.56
cc_43 VNB N_VGND_c_529_n 0.00698312f $X=-0.19 $Y=-0.245 $X2=2.265 $Y2=2.465
cc_44 VNB N_VGND_c_530_n 0.0171844f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_531_n 0.0235135f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_532_n 0.0171844f $X=-0.19 $Y=-0.245 $X2=2.695 $Y2=2.465
cc_47 VNB N_VGND_c_533_n 0.00500104f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_534_n 0.0171844f $X=-0.19 $Y=-0.245 $X2=3.125 $Y2=0.56
cc_49 VNB N_VGND_c_535_n 0.00500104f $X=-0.19 $Y=-0.245 $X2=3.125 $Y2=0.56
cc_50 VNB N_VGND_c_536_n 0.0171844f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_537_n 0.00500104f $X=-0.19 $Y=-0.245 $X2=3.125 $Y2=1.54
cc_52 VNB N_VGND_c_538_n 0.0347608f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_539_n 0.0328515f $X=-0.19 $Y=-0.245 $X2=4.415 $Y2=1.21
cc_54 VNB N_VGND_c_540_n 0.326397f $X=-0.19 $Y=-0.245 $X2=4.415 $Y2=0.56
cc_55 VNB N_VGND_c_541_n 0.00567425f $X=-0.19 $Y=-0.245 $X2=4.415 $Y2=1.54
cc_56 VNB N_VGND_c_542_n 0.00567425f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VPB N_A_M1000_g 0.0234928f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=2.465
cc_58 VPB N_A_M1003_g 0.018718f $X=-0.19 $Y=1.655 $X2=0.975 $Y2=2.465
cc_59 VPB N_A_M1005_g 0.0187369f $X=-0.19 $Y=1.655 $X2=1.405 $Y2=2.465
cc_60 VPB N_A_M1007_g 0.0187369f $X=-0.19 $Y=1.655 $X2=1.835 $Y2=2.465
cc_61 VPB N_A_M1008_g 0.0187369f $X=-0.19 $Y=1.655 $X2=2.265 $Y2=2.465
cc_62 VPB N_A_M1010_g 0.0187369f $X=-0.19 $Y=1.655 $X2=2.695 $Y2=2.465
cc_63 VPB N_A_M1012_g 0.0187369f $X=-0.19 $Y=1.655 $X2=3.125 $Y2=2.465
cc_64 VPB N_A_M1014_g 0.0187369f $X=-0.19 $Y=1.655 $X2=3.555 $Y2=2.465
cc_65 VPB N_A_M1015_g 0.0187369f $X=-0.19 $Y=1.655 $X2=3.985 $Y2=2.465
cc_66 VPB N_A_M1016_g 0.0187369f $X=-0.19 $Y=1.655 $X2=4.415 $Y2=2.465
cc_67 VPB N_A_M1017_g 0.0187175f $X=-0.19 $Y=1.655 $X2=4.845 $Y2=2.465
cc_68 VPB N_A_M1019_g 0.0234742f $X=-0.19 $Y=1.655 $X2=5.275 $Y2=2.465
cc_69 VPB N_VPWR_c_274_n 0.0135558f $X=-0.19 $Y=1.655 $X2=1.835 $Y2=2.465
cc_70 VPB N_VPWR_c_275_n 0.0421937f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_71 VPB N_VPWR_c_276_n 0.00400996f $X=-0.19 $Y=1.655 $X2=2.265 $Y2=2.465
cc_72 VPB N_VPWR_c_277_n 0.00400996f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_73 VPB N_VPWR_c_278_n 0.00400996f $X=-0.19 $Y=1.655 $X2=3.125 $Y2=0.56
cc_74 VPB N_VPWR_c_279_n 0.00400996f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_75 VPB N_VPWR_c_280_n 0.0167849f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_76 VPB N_VPWR_c_281_n 0.00400996f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_77 VPB N_VPWR_c_282_n 0.0116028f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_78 VPB N_VPWR_c_283_n 0.00460237f $X=-0.19 $Y=1.655 $X2=3.985 $Y2=2.465
cc_79 VPB N_VPWR_c_284_n 0.0167849f $X=-0.19 $Y=1.655 $X2=4.415 $Y2=0.56
cc_80 VPB N_VPWR_c_285_n 0.00497514f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_81 VPB N_VPWR_c_286_n 0.0167849f $X=-0.19 $Y=1.655 $X2=4.415 $Y2=2.465
cc_82 VPB N_VPWR_c_287_n 0.00497514f $X=-0.19 $Y=1.655 $X2=4.415 $Y2=2.465
cc_83 VPB N_VPWR_c_288_n 0.0167849f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_84 VPB N_VPWR_c_289_n 0.00497514f $X=-0.19 $Y=1.655 $X2=4.845 $Y2=1.54
cc_85 VPB N_VPWR_c_290_n 0.0167849f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_86 VPB N_VPWR_c_291_n 0.0167406f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_87 VPB N_VPWR_c_292_n 0.00497514f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_88 VPB N_VPWR_c_293_n 0.00497514f $X=-0.19 $Y=1.655 $X2=0.68 $Y2=1.375
cc_89 VPB N_VPWR_c_273_n 0.0501806f $X=-0.19 $Y=1.655 $X2=1.405 $Y2=1.375
cc_90 VPB N_Y_c_365_n 0.0025871f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_91 VPB N_Y_c_383_n 0.00201395f $X=-0.19 $Y=1.655 $X2=2.695 $Y2=0.56
cc_92 VPB N_Y_c_384_n 0.00873266f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_93 VPB N_Y_c_385_n 0.00243013f $X=-0.19 $Y=1.655 $X2=3.125 $Y2=0.56
cc_94 VPB N_Y_c_386_n 0.00243013f $X=-0.19 $Y=1.655 $X2=3.985 $Y2=1.21
cc_95 VPB N_Y_c_387_n 0.00243013f $X=-0.19 $Y=1.655 $X2=4.415 $Y2=2.465
cc_96 VPB N_Y_c_388_n 0.00243013f $X=-0.19 $Y=1.655 $X2=2.555 $Y2=1.21
cc_97 VPB N_Y_c_389_n 0.00242094f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_98 VPB N_Y_c_390_n 0.0089125f $X=-0.19 $Y=1.655 $X2=0.68 $Y2=1.375
cc_99 VPB N_Y_c_391_n 0.00206951f $X=-0.19 $Y=1.655 $X2=1.405 $Y2=1.375
cc_100 VPB N_Y_c_392_n 0.00206951f $X=-0.19 $Y=1.655 $X2=2.265 $Y2=1.375
cc_101 VPB N_Y_c_393_n 0.00206951f $X=-0.19 $Y=1.655 $X2=3.125 $Y2=1.375
cc_102 VPB N_Y_c_394_n 0.00206951f $X=-0.19 $Y=1.655 $X2=3.985 $Y2=1.375
cc_103 VPB N_Y_c_395_n 0.00206951f $X=-0.19 $Y=1.655 $X2=5.1 $Y2=1.375
cc_104 VPB N_Y_c_396_n 0.00211646f $X=-0.19 $Y=1.655 $X2=5.1 $Y2=1.375
cc_105 VPB Y 0.00255258f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_106 N_A_M1000_g N_VPWR_c_275_n 0.00342038f $X=0.545 $Y=2.465 $X2=0 $Y2=0
cc_107 N_A_M1003_g N_VPWR_c_276_n 0.0016342f $X=0.975 $Y=2.465 $X2=0 $Y2=0
cc_108 N_A_M1005_g N_VPWR_c_276_n 0.0016342f $X=1.405 $Y=2.465 $X2=0 $Y2=0
cc_109 N_A_M1007_g N_VPWR_c_277_n 0.0016342f $X=1.835 $Y=2.465 $X2=0 $Y2=0
cc_110 N_A_M1008_g N_VPWR_c_277_n 0.0016342f $X=2.265 $Y=2.465 $X2=0 $Y2=0
cc_111 N_A_M1010_g N_VPWR_c_278_n 0.0016342f $X=2.695 $Y=2.465 $X2=0 $Y2=0
cc_112 N_A_M1012_g N_VPWR_c_278_n 0.0016342f $X=3.125 $Y=2.465 $X2=0 $Y2=0
cc_113 N_A_M1014_g N_VPWR_c_279_n 0.0016342f $X=3.555 $Y=2.465 $X2=0 $Y2=0
cc_114 N_A_M1015_g N_VPWR_c_279_n 0.0016342f $X=3.985 $Y=2.465 $X2=0 $Y2=0
cc_115 N_A_M1015_g N_VPWR_c_280_n 0.00585385f $X=3.985 $Y=2.465 $X2=0 $Y2=0
cc_116 N_A_M1016_g N_VPWR_c_280_n 0.00585385f $X=4.415 $Y=2.465 $X2=0 $Y2=0
cc_117 N_A_M1016_g N_VPWR_c_281_n 0.0016342f $X=4.415 $Y=2.465 $X2=0 $Y2=0
cc_118 N_A_M1017_g N_VPWR_c_281_n 0.0016342f $X=4.845 $Y=2.465 $X2=0 $Y2=0
cc_119 N_A_M1019_g N_VPWR_c_283_n 0.00341773f $X=5.275 $Y=2.465 $X2=0 $Y2=0
cc_120 N_A_M1005_g N_VPWR_c_284_n 0.00585385f $X=1.405 $Y=2.465 $X2=0 $Y2=0
cc_121 N_A_M1007_g N_VPWR_c_284_n 0.00585385f $X=1.835 $Y=2.465 $X2=0 $Y2=0
cc_122 N_A_M1008_g N_VPWR_c_286_n 0.00585385f $X=2.265 $Y=2.465 $X2=0 $Y2=0
cc_123 N_A_M1010_g N_VPWR_c_286_n 0.00585385f $X=2.695 $Y=2.465 $X2=0 $Y2=0
cc_124 N_A_M1012_g N_VPWR_c_288_n 0.00585385f $X=3.125 $Y=2.465 $X2=0 $Y2=0
cc_125 N_A_M1014_g N_VPWR_c_288_n 0.00585385f $X=3.555 $Y=2.465 $X2=0 $Y2=0
cc_126 N_A_M1000_g N_VPWR_c_290_n 0.00585385f $X=0.545 $Y=2.465 $X2=0 $Y2=0
cc_127 N_A_M1003_g N_VPWR_c_290_n 0.00585385f $X=0.975 $Y=2.465 $X2=0 $Y2=0
cc_128 N_A_M1017_g N_VPWR_c_291_n 0.00585385f $X=4.845 $Y=2.465 $X2=0 $Y2=0
cc_129 N_A_M1019_g N_VPWR_c_291_n 0.00585385f $X=5.275 $Y=2.465 $X2=0 $Y2=0
cc_130 N_A_M1000_g N_VPWR_c_273_n 0.0116226f $X=0.545 $Y=2.465 $X2=0 $Y2=0
cc_131 N_A_M1003_g N_VPWR_c_273_n 0.0106302f $X=0.975 $Y=2.465 $X2=0 $Y2=0
cc_132 N_A_M1005_g N_VPWR_c_273_n 0.0106302f $X=1.405 $Y=2.465 $X2=0 $Y2=0
cc_133 N_A_M1007_g N_VPWR_c_273_n 0.0106302f $X=1.835 $Y=2.465 $X2=0 $Y2=0
cc_134 N_A_M1008_g N_VPWR_c_273_n 0.0106302f $X=2.265 $Y=2.465 $X2=0 $Y2=0
cc_135 N_A_M1010_g N_VPWR_c_273_n 0.0106302f $X=2.695 $Y=2.465 $X2=0 $Y2=0
cc_136 N_A_M1012_g N_VPWR_c_273_n 0.0106302f $X=3.125 $Y=2.465 $X2=0 $Y2=0
cc_137 N_A_M1014_g N_VPWR_c_273_n 0.0106302f $X=3.555 $Y=2.465 $X2=0 $Y2=0
cc_138 N_A_M1015_g N_VPWR_c_273_n 0.0106302f $X=3.985 $Y=2.465 $X2=0 $Y2=0
cc_139 N_A_M1016_g N_VPWR_c_273_n 0.0106302f $X=4.415 $Y=2.465 $X2=0 $Y2=0
cc_140 N_A_M1017_g N_VPWR_c_273_n 0.0106302f $X=4.845 $Y=2.465 $X2=0 $Y2=0
cc_141 N_A_M1019_g N_VPWR_c_273_n 0.0115721f $X=5.275 $Y=2.465 $X2=0 $Y2=0
cc_142 A N_Y_c_365_n 0.0262109f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_143 N_A_c_126_n N_Y_c_365_n 0.0152693f $X=5.275 $Y=1.375 $X2=0 $Y2=0
cc_144 N_A_M1001_g N_Y_c_366_n 0.0155371f $X=1.405 $Y=0.56 $X2=0 $Y2=0
cc_145 A N_Y_c_366_n 0.073583f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_146 N_A_c_126_n N_Y_c_366_n 0.0221841f $X=5.275 $Y=1.375 $X2=0 $Y2=0
cc_147 N_A_M1000_g N_Y_c_383_n 0.0165938f $X=0.545 $Y=2.465 $X2=0 $Y2=0
cc_148 A N_Y_c_383_n 0.00860651f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_149 N_A_M1003_g N_Y_c_385_n 0.0146426f $X=0.975 $Y=2.465 $X2=0 $Y2=0
cc_150 N_A_M1005_g N_Y_c_385_n 0.0146426f $X=1.405 $Y=2.465 $X2=0 $Y2=0
cc_151 A N_Y_c_385_n 0.0443704f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_152 N_A_c_126_n N_Y_c_385_n 0.00224353f $X=5.275 $Y=1.375 $X2=0 $Y2=0
cc_153 N_A_M1001_g N_Y_c_368_n 0.00194229f $X=1.405 $Y=0.56 $X2=0 $Y2=0
cc_154 N_A_M1002_g N_Y_c_368_n 0.00105846f $X=1.835 $Y=0.56 $X2=0 $Y2=0
cc_155 N_A_M1002_g N_Y_c_369_n 0.0131322f $X=1.835 $Y=0.56 $X2=0 $Y2=0
cc_156 N_A_M1004_g N_Y_c_369_n 0.0131322f $X=2.265 $Y=0.56 $X2=0 $Y2=0
cc_157 A N_Y_c_369_n 0.0444367f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_158 N_A_c_126_n N_Y_c_369_n 0.00225043f $X=5.275 $Y=1.375 $X2=0 $Y2=0
cc_159 N_A_M1007_g N_Y_c_386_n 0.0146426f $X=1.835 $Y=2.465 $X2=0 $Y2=0
cc_160 N_A_M1008_g N_Y_c_386_n 0.0146426f $X=2.265 $Y=2.465 $X2=0 $Y2=0
cc_161 A N_Y_c_386_n 0.0443704f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_162 N_A_c_126_n N_Y_c_386_n 0.00224353f $X=5.275 $Y=1.375 $X2=0 $Y2=0
cc_163 N_A_M1004_g N_Y_c_370_n 0.00105846f $X=2.265 $Y=0.56 $X2=0 $Y2=0
cc_164 N_A_M1006_g N_Y_c_370_n 0.00105846f $X=2.695 $Y=0.56 $X2=0 $Y2=0
cc_165 N_A_M1006_g N_Y_c_371_n 0.0131322f $X=2.695 $Y=0.56 $X2=0 $Y2=0
cc_166 N_A_M1009_g N_Y_c_371_n 0.0131322f $X=3.125 $Y=0.56 $X2=0 $Y2=0
cc_167 A N_Y_c_371_n 0.0444367f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_168 N_A_c_126_n N_Y_c_371_n 0.00225043f $X=5.275 $Y=1.375 $X2=0 $Y2=0
cc_169 N_A_M1010_g N_Y_c_387_n 0.0146426f $X=2.695 $Y=2.465 $X2=0 $Y2=0
cc_170 N_A_M1012_g N_Y_c_387_n 0.0146426f $X=3.125 $Y=2.465 $X2=0 $Y2=0
cc_171 A N_Y_c_387_n 0.0443704f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_172 N_A_c_126_n N_Y_c_387_n 0.00224353f $X=5.275 $Y=1.375 $X2=0 $Y2=0
cc_173 N_A_M1009_g N_Y_c_372_n 0.00105846f $X=3.125 $Y=0.56 $X2=0 $Y2=0
cc_174 N_A_M1011_g N_Y_c_372_n 0.00105846f $X=3.555 $Y=0.56 $X2=0 $Y2=0
cc_175 N_A_M1011_g N_Y_c_373_n 0.0131322f $X=3.555 $Y=0.56 $X2=0 $Y2=0
cc_176 N_A_M1013_g N_Y_c_373_n 0.0131322f $X=3.985 $Y=0.56 $X2=0 $Y2=0
cc_177 A N_Y_c_373_n 0.0444367f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_178 N_A_c_126_n N_Y_c_373_n 0.00225043f $X=5.275 $Y=1.375 $X2=0 $Y2=0
cc_179 N_A_M1014_g N_Y_c_388_n 0.0146426f $X=3.555 $Y=2.465 $X2=0 $Y2=0
cc_180 N_A_M1015_g N_Y_c_388_n 0.0146426f $X=3.985 $Y=2.465 $X2=0 $Y2=0
cc_181 A N_Y_c_388_n 0.0443704f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_182 N_A_c_126_n N_Y_c_388_n 0.00224353f $X=5.275 $Y=1.375 $X2=0 $Y2=0
cc_183 N_A_M1013_g N_Y_c_374_n 0.00105846f $X=3.985 $Y=0.56 $X2=0 $Y2=0
cc_184 N_A_M1018_g N_Y_c_374_n 0.00194229f $X=4.415 $Y=0.56 $X2=0 $Y2=0
cc_185 N_A_M1016_g N_Y_c_389_n 0.0146426f $X=4.415 $Y=2.465 $X2=0 $Y2=0
cc_186 N_A_M1017_g N_Y_c_389_n 0.0146085f $X=4.845 $Y=2.465 $X2=0 $Y2=0
cc_187 A N_Y_c_389_n 0.0439938f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_188 N_A_c_126_n N_Y_c_389_n 0.00224353f $X=5.275 $Y=1.375 $X2=0 $Y2=0
cc_189 N_A_M1019_g N_Y_c_390_n 0.0170121f $X=5.275 $Y=2.465 $X2=0 $Y2=0
cc_190 A N_Y_c_390_n 0.00536724f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_191 A N_Y_c_391_n 0.0215081f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_192 N_A_c_126_n N_Y_c_391_n 0.00232957f $X=5.275 $Y=1.375 $X2=0 $Y2=0
cc_193 A N_Y_c_375_n 0.0218346f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_194 N_A_c_126_n N_Y_c_375_n 0.00232201f $X=5.275 $Y=1.375 $X2=0 $Y2=0
cc_195 A N_Y_c_392_n 0.0215081f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_196 N_A_c_126_n N_Y_c_392_n 0.00232957f $X=5.275 $Y=1.375 $X2=0 $Y2=0
cc_197 A N_Y_c_376_n 0.0218346f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_198 N_A_c_126_n N_Y_c_376_n 0.00232201f $X=5.275 $Y=1.375 $X2=0 $Y2=0
cc_199 A N_Y_c_393_n 0.0215081f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_200 N_A_c_126_n N_Y_c_393_n 0.00232957f $X=5.275 $Y=1.375 $X2=0 $Y2=0
cc_201 A N_Y_c_377_n 0.0218346f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_202 N_A_c_126_n N_Y_c_377_n 0.00232201f $X=5.275 $Y=1.375 $X2=0 $Y2=0
cc_203 A N_Y_c_394_n 0.0215081f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_204 N_A_c_126_n N_Y_c_394_n 0.00232957f $X=5.275 $Y=1.375 $X2=0 $Y2=0
cc_205 A N_Y_c_378_n 0.0218346f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_206 N_A_c_126_n N_Y_c_378_n 0.00232201f $X=5.275 $Y=1.375 $X2=0 $Y2=0
cc_207 A N_Y_c_395_n 0.0215081f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_208 N_A_c_126_n N_Y_c_395_n 0.00232957f $X=5.275 $Y=1.375 $X2=0 $Y2=0
cc_209 A N_Y_c_396_n 0.0219298f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_210 N_A_c_126_n N_Y_c_396_n 0.00232957f $X=5.275 $Y=1.375 $X2=0 $Y2=0
cc_211 N_A_M1018_g Y 0.0155371f $X=4.415 $Y=0.56 $X2=0 $Y2=0
cc_212 A Y 0.0705391f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_213 N_A_c_126_n Y 0.0223886f $X=5.275 $Y=1.375 $X2=0 $Y2=0
cc_214 A Y 0.0263702f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_215 N_A_c_126_n Y 0.0160643f $X=5.275 $Y=1.375 $X2=0 $Y2=0
cc_216 N_A_M1001_g N_VGND_c_526_n 0.0038152f $X=1.405 $Y=0.56 $X2=0 $Y2=0
cc_217 N_A_M1002_g N_VGND_c_527_n 0.00181038f $X=1.835 $Y=0.56 $X2=0 $Y2=0
cc_218 N_A_M1004_g N_VGND_c_527_n 0.00181038f $X=2.265 $Y=0.56 $X2=0 $Y2=0
cc_219 N_A_M1006_g N_VGND_c_528_n 0.00181038f $X=2.695 $Y=0.56 $X2=0 $Y2=0
cc_220 N_A_M1009_g N_VGND_c_528_n 0.00181038f $X=3.125 $Y=0.56 $X2=0 $Y2=0
cc_221 N_A_M1011_g N_VGND_c_529_n 0.00181038f $X=3.555 $Y=0.56 $X2=0 $Y2=0
cc_222 N_A_M1013_g N_VGND_c_529_n 0.00181038f $X=3.985 $Y=0.56 $X2=0 $Y2=0
cc_223 N_A_M1013_g N_VGND_c_530_n 0.00478016f $X=3.985 $Y=0.56 $X2=0 $Y2=0
cc_224 N_A_M1018_g N_VGND_c_530_n 0.00478016f $X=4.415 $Y=0.56 $X2=0 $Y2=0
cc_225 N_A_M1018_g N_VGND_c_531_n 0.0038152f $X=4.415 $Y=0.56 $X2=0 $Y2=0
cc_226 N_A_M1001_g N_VGND_c_532_n 0.00478016f $X=1.405 $Y=0.56 $X2=0 $Y2=0
cc_227 N_A_M1002_g N_VGND_c_532_n 0.00478016f $X=1.835 $Y=0.56 $X2=0 $Y2=0
cc_228 N_A_M1004_g N_VGND_c_534_n 0.00478016f $X=2.265 $Y=0.56 $X2=0 $Y2=0
cc_229 N_A_M1006_g N_VGND_c_534_n 0.00478016f $X=2.695 $Y=0.56 $X2=0 $Y2=0
cc_230 N_A_M1009_g N_VGND_c_536_n 0.00478016f $X=3.125 $Y=0.56 $X2=0 $Y2=0
cc_231 N_A_M1011_g N_VGND_c_536_n 0.00478016f $X=3.555 $Y=0.56 $X2=0 $Y2=0
cc_232 N_A_M1001_g N_VGND_c_540_n 0.0051579f $X=1.405 $Y=0.56 $X2=0 $Y2=0
cc_233 N_A_M1002_g N_VGND_c_540_n 0.00490796f $X=1.835 $Y=0.56 $X2=0 $Y2=0
cc_234 N_A_M1004_g N_VGND_c_540_n 0.00490796f $X=2.265 $Y=0.56 $X2=0 $Y2=0
cc_235 N_A_M1006_g N_VGND_c_540_n 0.00490796f $X=2.695 $Y=0.56 $X2=0 $Y2=0
cc_236 N_A_M1009_g N_VGND_c_540_n 0.00490796f $X=3.125 $Y=0.56 $X2=0 $Y2=0
cc_237 N_A_M1011_g N_VGND_c_540_n 0.00490796f $X=3.555 $Y=0.56 $X2=0 $Y2=0
cc_238 N_A_M1013_g N_VGND_c_540_n 0.00490796f $X=3.985 $Y=0.56 $X2=0 $Y2=0
cc_239 N_A_M1018_g N_VGND_c_540_n 0.0051579f $X=4.415 $Y=0.56 $X2=0 $Y2=0
cc_240 N_VPWR_c_273_n N_Y_M1000_d 0.00320275f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_241 N_VPWR_c_273_n N_Y_M1005_d 0.00320275f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_242 N_VPWR_c_273_n N_Y_M1008_d 0.00320275f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_243 N_VPWR_c_273_n N_Y_M1012_d 0.00320275f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_244 N_VPWR_c_273_n N_Y_M1015_d 0.00320275f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_245 N_VPWR_c_273_n N_Y_M1017_d 0.00302905f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_246 N_VPWR_M1000_s N_Y_c_383_n 7.1286e-19 $X=0.205 $Y=1.835 $X2=0 $Y2=0
cc_247 N_VPWR_c_275_n N_Y_c_383_n 0.00550656f $X=0.33 $Y=2.22 $X2=0 $Y2=0
cc_248 N_VPWR_M1000_s N_Y_c_384_n 0.00178451f $X=0.205 $Y=1.835 $X2=0 $Y2=0
cc_249 N_VPWR_c_275_n N_Y_c_384_n 0.0129974f $X=0.33 $Y=2.22 $X2=0 $Y2=0
cc_250 N_VPWR_c_290_n N_Y_c_482_n 0.0124051f $X=1.06 $Y=3.33 $X2=0 $Y2=0
cc_251 N_VPWR_c_273_n N_Y_c_482_n 0.00969167f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_252 N_VPWR_M1003_s N_Y_c_385_n 0.00176619f $X=1.05 $Y=1.835 $X2=0 $Y2=0
cc_253 N_VPWR_c_276_n N_Y_c_385_n 0.0135319f $X=1.19 $Y=2.22 $X2=0 $Y2=0
cc_254 N_VPWR_c_284_n N_Y_c_486_n 0.0124051f $X=1.92 $Y=3.33 $X2=0 $Y2=0
cc_255 N_VPWR_c_273_n N_Y_c_486_n 0.00969167f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_256 N_VPWR_M1007_s N_Y_c_386_n 0.00176619f $X=1.91 $Y=1.835 $X2=0 $Y2=0
cc_257 N_VPWR_c_277_n N_Y_c_386_n 0.0135319f $X=2.05 $Y=2.22 $X2=0 $Y2=0
cc_258 N_VPWR_c_286_n N_Y_c_490_n 0.0124051f $X=2.78 $Y=3.33 $X2=0 $Y2=0
cc_259 N_VPWR_c_273_n N_Y_c_490_n 0.00969167f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_260 N_VPWR_M1010_s N_Y_c_387_n 0.00176619f $X=2.77 $Y=1.835 $X2=0 $Y2=0
cc_261 N_VPWR_c_278_n N_Y_c_387_n 0.0135319f $X=2.91 $Y=2.22 $X2=0 $Y2=0
cc_262 N_VPWR_c_288_n N_Y_c_494_n 0.0124051f $X=3.64 $Y=3.33 $X2=0 $Y2=0
cc_263 N_VPWR_c_273_n N_Y_c_494_n 0.00969167f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_264 N_VPWR_M1014_s N_Y_c_388_n 0.00176619f $X=3.63 $Y=1.835 $X2=0 $Y2=0
cc_265 N_VPWR_c_279_n N_Y_c_388_n 0.0135319f $X=3.77 $Y=2.22 $X2=0 $Y2=0
cc_266 N_VPWR_c_280_n N_Y_c_498_n 0.0124051f $X=4.5 $Y=3.33 $X2=0 $Y2=0
cc_267 N_VPWR_c_273_n N_Y_c_498_n 0.00969167f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_268 N_VPWR_M1016_s N_Y_c_389_n 0.00176619f $X=4.49 $Y=1.835 $X2=0 $Y2=0
cc_269 N_VPWR_c_281_n N_Y_c_389_n 0.0135319f $X=4.63 $Y=2.22 $X2=0 $Y2=0
cc_270 N_VPWR_c_291_n N_Y_c_502_n 0.012556f $X=5.36 $Y=3.33 $X2=0 $Y2=0
cc_271 N_VPWR_c_273_n N_Y_c_502_n 0.00988321f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_272 N_VPWR_M1019_s N_Y_c_390_n 0.00250337f $X=5.35 $Y=1.835 $X2=0 $Y2=0
cc_273 N_VPWR_c_283_n N_Y_c_390_n 0.0183848f $X=5.49 $Y=2.22 $X2=0 $Y2=0
cc_274 N_Y_c_366_n N_VGND_c_526_n 0.0219547f $X=1.49 $Y=0.94 $X2=0 $Y2=0
cc_275 N_Y_c_369_n N_VGND_c_527_n 0.0169602f $X=2.35 $Y=0.94 $X2=0 $Y2=0
cc_276 N_Y_c_371_n N_VGND_c_528_n 0.0169602f $X=3.21 $Y=0.94 $X2=0 $Y2=0
cc_277 N_Y_c_373_n N_VGND_c_529_n 0.0169602f $X=4.07 $Y=0.94 $X2=0 $Y2=0
cc_278 N_Y_c_374_n N_VGND_c_530_n 0.00786011f $X=4.2 $Y=0.56 $X2=0 $Y2=0
cc_279 Y N_VGND_c_531_n 0.0219547f $X=5.435 $Y=0.84 $X2=0 $Y2=0
cc_280 N_Y_c_368_n N_VGND_c_532_n 0.00786011f $X=1.62 $Y=0.56 $X2=0 $Y2=0
cc_281 N_Y_c_370_n N_VGND_c_534_n 0.00786011f $X=2.48 $Y=0.56 $X2=0 $Y2=0
cc_282 N_Y_c_372_n N_VGND_c_536_n 0.00786011f $X=3.34 $Y=0.56 $X2=0 $Y2=0
cc_283 N_Y_c_366_n N_VGND_c_540_n 0.0297069f $X=1.49 $Y=0.94 $X2=0 $Y2=0
cc_284 N_Y_c_367_n N_VGND_c_540_n 0.00670311f $X=0.345 $Y=0.94 $X2=0 $Y2=0
cc_285 N_Y_c_368_n N_VGND_c_540_n 0.00924776f $X=1.62 $Y=0.56 $X2=0 $Y2=0
cc_286 N_Y_c_369_n N_VGND_c_540_n 0.0106287f $X=2.35 $Y=0.94 $X2=0 $Y2=0
cc_287 N_Y_c_370_n N_VGND_c_540_n 0.00924776f $X=2.48 $Y=0.56 $X2=0 $Y2=0
cc_288 N_Y_c_371_n N_VGND_c_540_n 0.0106287f $X=3.21 $Y=0.94 $X2=0 $Y2=0
cc_289 N_Y_c_372_n N_VGND_c_540_n 0.00924776f $X=3.34 $Y=0.56 $X2=0 $Y2=0
cc_290 N_Y_c_373_n N_VGND_c_540_n 0.0106287f $X=4.07 $Y=0.94 $X2=0 $Y2=0
cc_291 N_Y_c_374_n N_VGND_c_540_n 0.00924776f $X=4.2 $Y=0.56 $X2=0 $Y2=0
cc_292 Y N_VGND_c_540_n 0.0283045f $X=5.435 $Y=0.84 $X2=0 $Y2=0
cc_293 N_Y_c_381_n N_VGND_c_540_n 0.00729456f $X=5.527 $Y=1.04 $X2=0 $Y2=0
