* File: sky130_fd_sc_lp__o32ai_0.pxi.spice
* Created: Wed Sep  2 10:26:34 2020
* 
x_PM_SKY130_FD_SC_LP__O32AI_0%B1 N_B1_c_66_n N_B1_M1003_g N_B1_c_67_n
+ N_B1_M1006_g B1 B1 B1 B1 PM_SKY130_FD_SC_LP__O32AI_0%B1
x_PM_SKY130_FD_SC_LP__O32AI_0%B2 N_B2_M1007_g N_B2_M1000_g N_B2_c_99_n
+ N_B2_c_100_n B2 B2 N_B2_c_97_n PM_SKY130_FD_SC_LP__O32AI_0%B2
x_PM_SKY130_FD_SC_LP__O32AI_0%A3 N_A3_M1002_g N_A3_c_140_n N_A3_M1004_g
+ N_A3_c_145_n A3 A3 A3 A3 A3 N_A3_c_142_n PM_SKY130_FD_SC_LP__O32AI_0%A3
x_PM_SKY130_FD_SC_LP__O32AI_0%A2 N_A2_M1008_g N_A2_M1005_g N_A2_c_185_n
+ N_A2_c_190_n A2 A2 A2 A2 A2 N_A2_c_187_n PM_SKY130_FD_SC_LP__O32AI_0%A2
x_PM_SKY130_FD_SC_LP__O32AI_0%A1 N_A1_M1009_g N_A1_M1001_g N_A1_c_231_n
+ N_A1_c_232_n N_A1_c_227_n N_A1_c_234_n A1 A1 A1 N_A1_c_229_n
+ PM_SKY130_FD_SC_LP__O32AI_0%A1
x_PM_SKY130_FD_SC_LP__O32AI_0%VPWR N_VPWR_M1006_s N_VPWR_M1009_d N_VPWR_c_264_n
+ N_VPWR_c_265_n N_VPWR_c_266_n VPWR N_VPWR_c_267_n N_VPWR_c_268_n
+ N_VPWR_c_263_n N_VPWR_c_270_n PM_SKY130_FD_SC_LP__O32AI_0%VPWR
x_PM_SKY130_FD_SC_LP__O32AI_0%Y N_Y_M1003_d N_Y_M1007_d Y Y Y Y Y Y N_Y_c_302_n
+ Y Y PM_SKY130_FD_SC_LP__O32AI_0%Y
x_PM_SKY130_FD_SC_LP__O32AI_0%A_33_82# N_A_33_82#_M1003_s N_A_33_82#_M1000_d
+ N_A_33_82#_M1005_d N_A_33_82#_c_340_n N_A_33_82#_c_341_n N_A_33_82#_c_342_n
+ N_A_33_82#_c_343_n N_A_33_82#_c_344_n N_A_33_82#_c_345_n
+ PM_SKY130_FD_SC_LP__O32AI_0%A_33_82#
x_PM_SKY130_FD_SC_LP__O32AI_0%VGND N_VGND_M1002_d N_VGND_M1001_d N_VGND_c_380_n
+ N_VGND_c_381_n N_VGND_c_382_n N_VGND_c_383_n VGND N_VGND_c_384_n
+ N_VGND_c_385_n PM_SKY130_FD_SC_LP__O32AI_0%VGND
cc_1 VNB N_B1_c_66_n 0.0194136f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=0.94
cc_2 VNB N_B1_c_67_n 0.0799905f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.61
cc_3 VNB N_B1_M1006_g 0.0021491f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=2.775
cc_4 VNB B1 0.0345917f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_5 VNB N_B2_M1000_g 0.047337f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_6 VNB B2 0.00590685f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_B2_c_97_n 0.011193f $X=-0.19 $Y=-0.245 $X2=0.37 $Y2=1.105
cc_8 VNB N_A3_M1002_g 0.034294f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=0.62
cc_9 VNB N_A3_c_140_n 0.0180136f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=2.775
cc_10 VNB A3 0.00535933f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A3_c_142_n 0.0287989f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.295
cc_12 VNB N_A2_M1005_g 0.0343462f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A2_c_185_n 0.0179649f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.95
cc_14 VNB A2 0.00442373f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A2_c_187_n 0.015659f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A1_M1001_g 0.0423614f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A1_c_227_n 0.0209836f $X=-0.19 $Y=-0.245 $X2=0.37 $Y2=1.105
cc_18 VNB A1 0.0255889f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=0.925
cc_19 VNB N_A1_c_229_n 0.0175475f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_VPWR_c_263_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.665
cc_21 VNB Y 0.00168558f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_22 VNB N_Y_c_302_n 0.00189298f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.295
cc_23 VNB Y 0.00394974f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_33_82#_c_340_n 0.00747548f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_25 VNB N_A_33_82#_c_341_n 6.35322e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_33_82#_c_342_n 0.0294102f $X=-0.19 $Y=-0.245 $X2=0.435 $Y2=1.105
cc_27 VNB N_A_33_82#_c_343_n 0.00375536f $X=-0.19 $Y=-0.245 $X2=0.37 $Y2=1.105
cc_28 VNB N_A_33_82#_c_344_n 7.93408e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_33_82#_c_345_n 0.019351f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.105
cc_30 VNB N_VGND_c_380_n 0.029926f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_31 VNB N_VGND_c_381_n 0.0113717f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.95
cc_32 VNB N_VGND_c_382_n 0.0174847f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_383_n 0.00519339f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_384_n 0.0607781f $X=-0.19 $Y=-0.245 $X2=0.435 $Y2=1.105
cc_35 VNB N_VGND_c_385_n 0.220959f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VPB N_B1_M1006_g 0.058254f $X=-0.19 $Y=1.655 $X2=0.59 $Y2=2.775
cc_37 VPB B1 0.0367621f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_38 VPB N_B2_M1007_g 0.0237392f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=0.62
cc_39 VPB N_B2_c_99_n 0.021756f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.95
cc_40 VPB N_B2_c_100_n 0.0157583f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_41 VPB B2 0.00660172f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_42 VPB N_B2_c_97_n 0.00450569f $X=-0.19 $Y=1.655 $X2=0.37 $Y2=1.105
cc_43 VPB N_A3_c_140_n 0.00379865f $X=-0.19 $Y=1.655 $X2=0.59 $Y2=2.775
cc_44 VPB N_A3_M1004_g 0.0430376f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_45 VPB N_A3_c_145_n 0.0157612f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.95
cc_46 VPB A3 0.0053653f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_47 VPB N_A2_M1008_g 0.0389499f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=0.62
cc_48 VPB N_A2_c_185_n 0.00379902f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.95
cc_49 VPB N_A2_c_190_n 0.016786f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_50 VPB A2 0.00975002f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_51 VPB N_A1_M1009_g 0.027675f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=0.62
cc_52 VPB N_A1_c_231_n 0.0149304f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_53 VPB N_A1_c_232_n 0.0258865f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_54 VPB N_A1_c_227_n 0.0044374f $X=-0.19 $Y=1.655 $X2=0.37 $Y2=1.105
cc_55 VPB N_A1_c_234_n 0.0175475f $X=-0.19 $Y=1.655 $X2=0.37 $Y2=1.105
cc_56 VPB A1 0.03061f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=0.925
cc_57 VPB N_VPWR_c_264_n 0.013523f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_58 VPB N_VPWR_c_265_n 0.032559f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_59 VPB N_VPWR_c_266_n 0.00694267f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_60 VPB N_VPWR_c_267_n 0.0579169f $X=-0.19 $Y=1.655 $X2=0.37 $Y2=1.105
cc_61 VPB N_VPWR_c_268_n 0.0190089f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_62 VPB N_VPWR_c_263_n 0.06546f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.665
cc_63 VPB N_VPWR_c_270_n 0.00401341f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_64 VPB Y 0.00480454f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_65 VPB Y 0.0073994f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_66 N_B1_c_66_n N_B2_M1000_g 0.0197694f $X=0.505 $Y=0.94 $X2=0 $Y2=0
cc_67 N_B1_c_67_n N_B2_M1000_g 0.0221168f $X=0.59 $Y=1.61 $X2=0 $Y2=0
cc_68 B1 N_B2_M1000_g 4.85633e-19 $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_69 N_B1_M1006_g N_B2_c_100_n 0.0441339f $X=0.59 $Y=2.775 $X2=0 $Y2=0
cc_70 N_B1_c_67_n B2 5.75355e-19 $X=0.59 $Y=1.61 $X2=0 $Y2=0
cc_71 N_B1_c_67_n N_B2_c_97_n 0.0441339f $X=0.59 $Y=1.61 $X2=0 $Y2=0
cc_72 N_B1_M1006_g N_VPWR_c_265_n 0.00775271f $X=0.59 $Y=2.775 $X2=0 $Y2=0
cc_73 B1 N_VPWR_c_265_n 0.018491f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_74 N_B1_M1006_g N_VPWR_c_267_n 0.00531267f $X=0.59 $Y=2.775 $X2=0 $Y2=0
cc_75 N_B1_M1006_g N_VPWR_c_263_n 0.0102522f $X=0.59 $Y=2.775 $X2=0 $Y2=0
cc_76 N_B1_c_67_n Y 0.00557588f $X=0.59 $Y=1.61 $X2=0 $Y2=0
cc_77 N_B1_M1006_g Y 0.0225528f $X=0.59 $Y=2.775 $X2=0 $Y2=0
cc_78 N_B1_M1006_g Y 0.0122372f $X=0.59 $Y=2.775 $X2=0 $Y2=0
cc_79 N_B1_c_66_n N_Y_c_302_n 0.00379195f $X=0.505 $Y=0.94 $X2=0 $Y2=0
cc_80 N_B1_c_67_n N_Y_c_302_n 0.00477415f $X=0.59 $Y=1.61 $X2=0 $Y2=0
cc_81 B1 N_Y_c_302_n 0.104182f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_82 N_B1_c_67_n Y 0.00479922f $X=0.59 $Y=1.61 $X2=0 $Y2=0
cc_83 N_B1_c_66_n N_A_33_82#_c_340_n 0.0114775f $X=0.505 $Y=0.94 $X2=0 $Y2=0
cc_84 N_B1_c_66_n N_A_33_82#_c_345_n 0.00820247f $X=0.505 $Y=0.94 $X2=0 $Y2=0
cc_85 N_B1_c_67_n N_A_33_82#_c_345_n 0.0011777f $X=0.59 $Y=1.61 $X2=0 $Y2=0
cc_86 B1 N_A_33_82#_c_345_n 0.0258364f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_87 N_B1_c_66_n N_VGND_c_384_n 8.96016e-19 $X=0.505 $Y=0.94 $X2=0 $Y2=0
cc_88 B1 N_VGND_c_385_n 0.0021706f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_89 N_B2_M1000_g N_A3_M1002_g 0.0302789f $X=1.005 $Y=0.62 $X2=0 $Y2=0
cc_90 N_B2_M1000_g N_A3_c_140_n 0.0051987f $X=1.005 $Y=0.62 $X2=0 $Y2=0
cc_91 B2 N_A3_c_140_n 0.00460306f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_92 N_B2_c_97_n N_A3_c_140_n 0.0113192f $X=1.07 $Y=1.725 $X2=0 $Y2=0
cc_93 N_B2_M1007_g N_A3_M1004_g 0.0162519f $X=0.98 $Y=2.775 $X2=0 $Y2=0
cc_94 N_B2_c_100_n N_A3_M1004_g 0.0113192f $X=1.07 $Y=2.23 $X2=0 $Y2=0
cc_95 N_B2_c_99_n N_A3_c_145_n 0.0113192f $X=1.07 $Y=2.065 $X2=0 $Y2=0
cc_96 N_B2_M1007_g A3 0.00113245f $X=0.98 $Y=2.775 $X2=0 $Y2=0
cc_97 N_B2_M1000_g A3 0.00132143f $X=1.005 $Y=0.62 $X2=0 $Y2=0
cc_98 B2 A3 0.0467619f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_99 N_B2_c_97_n A3 6.10052e-19 $X=1.07 $Y=1.725 $X2=0 $Y2=0
cc_100 N_B2_M1007_g N_VPWR_c_267_n 0.00378316f $X=0.98 $Y=2.775 $X2=0 $Y2=0
cc_101 N_B2_M1007_g N_VPWR_c_263_n 0.00567148f $X=0.98 $Y=2.775 $X2=0 $Y2=0
cc_102 N_B2_M1000_g Y 0.00268811f $X=1.005 $Y=0.62 $X2=0 $Y2=0
cc_103 B2 Y 0.0511475f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_104 N_B2_c_97_n Y 0.00803772f $X=1.07 $Y=1.725 $X2=0 $Y2=0
cc_105 N_B2_M1007_g Y 0.0220924f $X=0.98 $Y=2.775 $X2=0 $Y2=0
cc_106 N_B2_c_100_n Y 0.0013615f $X=1.07 $Y=2.23 $X2=0 $Y2=0
cc_107 B2 Y 0.0284935f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_108 N_B2_M1000_g N_Y_c_302_n 0.0128078f $X=1.005 $Y=0.62 $X2=0 $Y2=0
cc_109 N_B2_M1000_g Y 0.00615799f $X=1.005 $Y=0.62 $X2=0 $Y2=0
cc_110 N_B2_c_97_n Y 0.00120964f $X=1.07 $Y=1.725 $X2=0 $Y2=0
cc_111 N_B2_M1000_g N_A_33_82#_c_340_n 0.0134278f $X=1.005 $Y=0.62 $X2=0 $Y2=0
cc_112 N_B2_M1000_g N_A_33_82#_c_341_n 3.46989e-19 $X=1.005 $Y=0.62 $X2=0 $Y2=0
cc_113 B2 N_A_33_82#_c_342_n 0.00149542f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_114 N_B2_M1000_g N_A_33_82#_c_343_n 0.0014023f $X=1.005 $Y=0.62 $X2=0 $Y2=0
cc_115 B2 N_A_33_82#_c_343_n 0.00764495f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_116 N_B2_c_97_n N_A_33_82#_c_343_n 7.2323e-19 $X=1.07 $Y=1.725 $X2=0 $Y2=0
cc_117 N_B2_M1000_g N_A_33_82#_c_345_n 4.06422e-19 $X=1.005 $Y=0.62 $X2=0 $Y2=0
cc_118 N_B2_M1000_g N_VGND_c_384_n 9.02242e-19 $X=1.005 $Y=0.62 $X2=0 $Y2=0
cc_119 N_A3_M1004_g N_A2_M1008_g 0.0360685f $X=1.55 $Y=2.775 $X2=0 $Y2=0
cc_120 N_A3_M1002_g N_A2_M1005_g 0.00921903f $X=1.435 $Y=0.62 $X2=0 $Y2=0
cc_121 N_A3_c_140_n N_A2_c_185_n 0.0122526f $X=1.64 $Y=1.715 $X2=0 $Y2=0
cc_122 N_A3_c_145_n N_A2_c_190_n 0.0122526f $X=1.64 $Y=1.88 $X2=0 $Y2=0
cc_123 N_A3_M1004_g A2 0.00173102f $X=1.55 $Y=2.775 $X2=0 $Y2=0
cc_124 A3 A2 0.121699f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_125 N_A3_c_142_n A2 0.00210709f $X=1.64 $Y=1.375 $X2=0 $Y2=0
cc_126 A3 N_A2_c_187_n 0.00570596f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_127 N_A3_c_142_n N_A2_c_187_n 0.0122526f $X=1.64 $Y=1.375 $X2=0 $Y2=0
cc_128 N_A3_M1004_g N_VPWR_c_267_n 0.00492032f $X=1.55 $Y=2.775 $X2=0 $Y2=0
cc_129 A3 N_VPWR_c_267_n 0.00960038f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_130 N_A3_M1004_g N_VPWR_c_263_n 0.00916689f $X=1.55 $Y=2.775 $X2=0 $Y2=0
cc_131 A3 N_VPWR_c_263_n 0.00974272f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_132 N_A3_M1004_g Y 0.00821442f $X=1.55 $Y=2.775 $X2=0 $Y2=0
cc_133 A3 Y 0.0420807f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_134 N_A3_M1002_g N_Y_c_302_n 9.45291e-19 $X=1.435 $Y=0.62 $X2=0 $Y2=0
cc_135 A3 N_Y_c_302_n 0.00468475f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_136 N_A3_c_142_n Y 7.41495e-19 $X=1.64 $Y=1.375 $X2=0 $Y2=0
cc_137 A3 A_325_491# 0.00696696f $X=1.595 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_138 N_A3_M1002_g N_A_33_82#_c_340_n 0.00113299f $X=1.435 $Y=0.62 $X2=0 $Y2=0
cc_139 N_A3_M1002_g N_A_33_82#_c_341_n 0.00101119f $X=1.435 $Y=0.62 $X2=0 $Y2=0
cc_140 N_A3_M1002_g N_A_33_82#_c_342_n 0.0192278f $X=1.435 $Y=0.62 $X2=0 $Y2=0
cc_141 A3 N_A_33_82#_c_342_n 0.0223484f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_142 N_A3_c_142_n N_A_33_82#_c_342_n 0.00364271f $X=1.64 $Y=1.375 $X2=0 $Y2=0
cc_143 N_A3_M1002_g N_VGND_c_384_n 0.0122821f $X=1.435 $Y=0.62 $X2=0 $Y2=0
cc_144 N_A3_M1002_g N_VGND_c_385_n 0.00447788f $X=1.435 $Y=0.62 $X2=0 $Y2=0
cc_145 N_A2_M1005_g N_A1_M1001_g 0.023243f $X=2.26 $Y=0.62 $X2=0 $Y2=0
cc_146 N_A2_M1008_g N_A1_c_231_n 0.00612201f $X=2.12 $Y=2.775 $X2=0 $Y2=0
cc_147 A2 N_A1_c_231_n 7.18226e-19 $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_148 N_A2_M1008_g N_A1_c_232_n 0.0568453f $X=2.12 $Y=2.775 $X2=0 $Y2=0
cc_149 A2 N_A1_c_232_n 0.0104378f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_150 N_A2_c_185_n N_A1_c_227_n 0.0116592f $X=2.21 $Y=1.715 $X2=0 $Y2=0
cc_151 N_A2_c_190_n N_A1_c_234_n 0.0116592f $X=2.21 $Y=1.88 $X2=0 $Y2=0
cc_152 N_A2_M1008_g A1 7.95332e-19 $X=2.12 $Y=2.775 $X2=0 $Y2=0
cc_153 A2 A1 0.0828401f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_154 N_A2_c_187_n A1 0.00450916f $X=2.21 $Y=1.375 $X2=0 $Y2=0
cc_155 A2 N_A1_c_229_n 6.45798e-19 $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_156 N_A2_c_187_n N_A1_c_229_n 0.0116592f $X=2.21 $Y=1.375 $X2=0 $Y2=0
cc_157 A2 N_VPWR_c_266_n 0.0141025f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_158 N_A2_M1008_g N_VPWR_c_267_n 0.00382445f $X=2.12 $Y=2.775 $X2=0 $Y2=0
cc_159 A2 N_VPWR_c_267_n 0.0106905f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_160 N_A2_M1008_g N_VPWR_c_263_n 0.00578247f $X=2.12 $Y=2.775 $X2=0 $Y2=0
cc_161 A2 N_VPWR_c_263_n 0.01116f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_162 A2 A_439_491# 0.00613245f $X=2.075 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_163 N_A2_M1005_g N_A_33_82#_c_342_n 0.0150846f $X=2.26 $Y=0.62 $X2=0 $Y2=0
cc_164 A2 N_A_33_82#_c_342_n 0.0258323f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_165 N_A2_c_187_n N_A_33_82#_c_342_n 0.00261825f $X=2.21 $Y=1.375 $X2=0 $Y2=0
cc_166 N_A2_M1005_g N_A_33_82#_c_344_n 0.0010204f $X=2.26 $Y=0.62 $X2=0 $Y2=0
cc_167 N_A2_M1005_g N_VGND_c_382_n 0.00457257f $X=2.26 $Y=0.62 $X2=0 $Y2=0
cc_168 N_A2_M1005_g N_VGND_c_384_n 0.00917212f $X=2.26 $Y=0.62 $X2=0 $Y2=0
cc_169 N_A2_M1005_g N_VGND_c_385_n 0.00447788f $X=2.26 $Y=0.62 $X2=0 $Y2=0
cc_170 N_A1_M1009_g N_VPWR_c_266_n 0.00484825f $X=2.51 $Y=2.775 $X2=0 $Y2=0
cc_171 N_A1_c_232_n N_VPWR_c_266_n 0.00402495f $X=2.69 $Y=2.195 $X2=0 $Y2=0
cc_172 N_A1_c_234_n N_VPWR_c_266_n 2.5158e-19 $X=2.78 $Y=1.88 $X2=0 $Y2=0
cc_173 A1 N_VPWR_c_266_n 0.0153079f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_174 N_A1_M1009_g N_VPWR_c_267_n 0.00585385f $X=2.51 $Y=2.775 $X2=0 $Y2=0
cc_175 N_A1_M1009_g N_VPWR_c_263_n 0.011917f $X=2.51 $Y=2.775 $X2=0 $Y2=0
cc_176 N_A1_M1001_g N_A_33_82#_c_342_n 0.00551383f $X=2.69 $Y=0.62 $X2=0 $Y2=0
cc_177 A1 N_A_33_82#_c_342_n 0.00685711f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_178 N_A1_M1001_g N_A_33_82#_c_344_n 0.00103408f $X=2.69 $Y=0.62 $X2=0 $Y2=0
cc_179 N_A1_M1001_g N_VGND_c_380_n 0.00403646f $X=2.69 $Y=0.62 $X2=0 $Y2=0
cc_180 A1 N_VGND_c_380_n 0.0061266f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_181 N_A1_c_229_n N_VGND_c_380_n 9.04298e-19 $X=2.78 $Y=1.375 $X2=0 $Y2=0
cc_182 N_A1_M1001_g N_VGND_c_382_n 0.00548708f $X=2.69 $Y=0.62 $X2=0 $Y2=0
cc_183 N_A1_M1001_g N_VGND_c_384_n 5.28126e-19 $X=2.69 $Y=0.62 $X2=0 $Y2=0
cc_184 N_A1_M1001_g N_VGND_c_385_n 0.00533081f $X=2.69 $Y=0.62 $X2=0 $Y2=0
cc_185 N_VPWR_c_263_n A_133_491# 0.00206003f $X=3.12 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_186 N_VPWR_c_263_n N_Y_M1007_d 0.00652051f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_187 N_VPWR_c_265_n Y 0.0452904f $X=0.37 $Y=2.6 $X2=0 $Y2=0
cc_188 N_VPWR_c_267_n Y 0.0359884f $X=2.62 $Y=3.33 $X2=0 $Y2=0
cc_189 N_VPWR_c_263_n Y 0.0273899f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_190 N_VPWR_c_263_n A_325_491# 0.0095155f $X=3.12 $Y=3.33 $X2=-0.19 $Y2=-0.245
cc_191 N_VPWR_c_263_n A_439_491# 0.00551885f $X=3.12 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_192 A_133_491# Y 0.00157559f $X=0.665 $Y=2.455 $X2=2.725 $Y2=2.61
cc_193 N_Y_M1003_d N_A_33_82#_c_340_n 0.00248745f $X=0.58 $Y=0.41 $X2=0 $Y2=0
cc_194 N_Y_c_302_n N_A_33_82#_c_340_n 0.0196355f $X=0.79 $Y=0.705 $X2=0 $Y2=0
cc_195 N_Y_c_302_n N_A_33_82#_c_341_n 0.0117727f $X=0.79 $Y=0.705 $X2=0 $Y2=0
cc_196 N_Y_c_302_n N_A_33_82#_c_343_n 0.0143344f $X=0.79 $Y=0.705 $X2=0 $Y2=0
cc_197 N_A_33_82#_c_344_n N_VGND_c_382_n 0.00548314f $X=2.475 $Y=0.62 $X2=0
+ $Y2=0
cc_198 N_A_33_82#_c_340_n N_VGND_c_384_n 0.0712062f $X=1.125 $Y=0.34 $X2=0 $Y2=0
cc_199 N_A_33_82#_c_342_n N_VGND_c_384_n 0.0542712f $X=2.38 $Y=0.955 $X2=0 $Y2=0
cc_200 N_A_33_82#_c_345_n N_VGND_c_384_n 0.0226635f $X=0.29 $Y=0.34 $X2=0 $Y2=0
cc_201 N_A_33_82#_c_340_n N_VGND_c_385_n 0.0325733f $X=1.125 $Y=0.34 $X2=0 $Y2=0
cc_202 N_A_33_82#_c_344_n N_VGND_c_385_n 0.00679302f $X=2.475 $Y=0.62 $X2=0
+ $Y2=0
cc_203 N_A_33_82#_c_345_n N_VGND_c_385_n 0.0125932f $X=0.29 $Y=0.34 $X2=0 $Y2=0
