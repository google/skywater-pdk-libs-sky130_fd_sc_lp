* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__xor3_lp A B C VGND VNB VPB VPWR X
X0 a_1245_89# B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 a_494_419# a_580_21# a_57_113# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X2 a_580_21# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X3 VGND a_1459_406# a_2046_141# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 a_494_419# C a_1459_406# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 a_388_419# a_580_21# a_494_419# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 a_1860_141# C VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 a_144_113# A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 a_855_66# a_580_21# a_388_419# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X9 a_1459_406# a_1393_300# a_855_66# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 a_1393_300# C a_1860_141# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X11 a_1459_406# C a_855_66# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X12 a_57_113# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X13 a_57_113# a_580_21# a_855_66# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X14 VGND a_57_113# a_430_113# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X15 a_388_419# B a_494_419# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X16 a_57_113# B a_855_66# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X17 a_494_419# a_1393_300# a_1459_406# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X18 a_855_66# B a_388_419# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X19 a_494_419# B a_57_113# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X20 a_1393_300# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X21 VPWR a_1459_406# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X22 a_430_113# a_57_113# a_388_419# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X23 a_2046_141# a_1459_406# X VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X24 VPWR a_57_113# a_388_419# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X25 a_57_113# A a_144_113# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X26 a_580_21# B a_1245_89# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
