* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__or4b_2 A B C D_N VGND VNB VPB VPWR X
X0 VPWR A a_436_385# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X1 X a_189_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X2 a_508_385# C a_616_385# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X3 a_616_385# a_31_131# a_189_21# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X4 a_436_385# B a_508_385# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X5 VGND C a_189_21# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 a_31_131# D_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X7 VGND a_189_21# X VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X8 VGND A a_189_21# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 X a_189_21# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X10 a_189_21# a_31_131# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X11 a_189_21# B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 a_31_131# D_N VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X13 VPWR a_189_21# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
.ends
