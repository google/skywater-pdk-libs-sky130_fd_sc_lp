* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__o21ba_2 A1 A2 B1_N VGND VNB VPB VPWR X
M1000 a_186_21# a_28_131# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=3.654e+11p pd=3.1e+06u as=1.3125e+12p ps=9.95e+06u
M1001 X a_186_21# VGND VNB nshort w=840000u l=150000u
+  ad=2.352e+11p pd=2.24e+06u as=7.938e+11p ps=7.04e+06u
M1002 VGND A2 a_492_47# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=4.746e+11p ps=4.49e+06u
M1003 a_492_47# A1 VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VPWR A1 a_564_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=5.355e+11p ps=3.37e+06u
M1005 VGND a_186_21# X VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_564_367# A2 a_186_21# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_492_47# a_28_131# a_186_21# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=2.226e+11p ps=2.21e+06u
M1008 VGND B1_N a_28_131# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1009 VPWR a_186_21# X VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=3.528e+11p ps=3.08e+06u
M1010 VPWR B1_N a_28_131# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1011 X a_186_21# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
