* NGSPICE file created from sky130_fd_sc_lp__dfxtp_4.ext - technology: sky130A

.subckt sky130_fd_sc_lp__dfxtp_4 CLK D VGND VNB VPB VPWR Q
M1000 a_526_413# a_110_70# a_431_119# VNB nshort w=420000u l=150000u
+  ad=1.575e+11p pd=1.59e+06u as=1.596e+11p ps=1.6e+06u
M1001 VGND a_684_93# a_642_119# VNB nshort w=420000u l=150000u
+  ad=1.5787e+12p pd=1.465e+07u as=8.82e+10p ps=1.26e+06u
M1002 VPWR a_1112_93# Q VPB phighvt w=1.26e+06u l=150000u
+  ad=2.2113e+12p pd=1.945e+07u as=7.056e+11p ps=6.16e+06u
M1003 a_684_93# a_526_413# VPWR VPB phighvt w=840000u l=150000u
+  ad=2.352e+11p pd=2.24e+06u as=0p ps=0u
M1004 a_110_70# CLK VGND VNB nshort w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1005 a_642_119# a_217_413# a_526_413# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_1116_441# a_217_413# a_941_379# VPB phighvt w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=5.06225e+11p ps=3.13e+06u
M1007 a_941_379# a_217_413# a_684_93# VNB nshort w=420000u l=150000u
+  ad=1.491e+11p pd=1.55e+06u as=2.239e+11p ps=2.07e+06u
M1008 a_526_413# a_217_413# a_431_119# VPB phighvt w=420000u l=150000u
+  ad=2.31e+11p pd=1.94e+06u as=1.176e+11p ps=1.4e+06u
M1009 Q a_1112_93# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND a_1112_93# a_1070_119# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1011 VGND a_110_70# a_217_413# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1012 VPWR a_1112_93# a_1116_441# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 Q a_1112_93# VGND VNB nshort w=840000u l=150000u
+  ad=4.704e+11p pd=4.48e+06u as=0p ps=0u
M1014 Q a_1112_93# VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VPWR a_110_70# a_217_413# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.696e+11p ps=1.81e+06u
M1016 a_684_93# a_526_413# VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_1070_119# a_110_70# a_941_379# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 Q a_1112_93# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_431_119# D VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VGND a_1112_93# Q VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_941_379# a_110_70# a_684_93# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_666_413# a_110_70# a_526_413# VPB phighvt w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1023 a_110_70# CLK VPWR VPB phighvt w=640000u l=150000u
+  ad=1.696e+11p pd=1.81e+06u as=0p ps=0u
M1024 VPWR a_684_93# a_666_413# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 VPWR a_1112_93# Q VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_1112_93# a_941_379# VGND VNB nshort w=840000u l=150000u
+  ad=2.394e+11p pd=2.25e+06u as=0p ps=0u
M1027 a_431_119# D VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_1112_93# a_941_379# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=3.339e+11p pd=3.05e+06u as=0p ps=0u
M1029 VGND a_1112_93# Q VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

