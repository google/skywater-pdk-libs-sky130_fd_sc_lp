* File: sky130_fd_sc_lp__o211a_m.pxi.spice
* Created: Wed Sep  2 10:14:14 2020
* 
x_PM_SKY130_FD_SC_LP__O211A_M%A_80_60# N_A_80_60#_M1006_d N_A_80_60#_M1009_d
+ N_A_80_60#_M1001_d N_A_80_60#_M1002_g N_A_80_60#_M1003_g N_A_80_60#_c_63_n
+ N_A_80_60#_c_64_n N_A_80_60#_c_68_n N_A_80_60#_c_69_n N_A_80_60#_c_93_p
+ N_A_80_60#_c_70_n N_A_80_60#_c_65_n N_A_80_60#_c_72_n N_A_80_60#_c_73_n
+ N_A_80_60#_c_103_p N_A_80_60#_c_74_n PM_SKY130_FD_SC_LP__O211A_M%A_80_60#
x_PM_SKY130_FD_SC_LP__O211A_M%A1 N_A1_M1000_g N_A1_M1007_g N_A1_c_140_n
+ N_A1_c_141_n A1 N_A1_c_142_n N_A1_c_152_n PM_SKY130_FD_SC_LP__O211A_M%A1
x_PM_SKY130_FD_SC_LP__O211A_M%A2 N_A2_M1009_g N_A2_M1005_g N_A2_c_180_n
+ N_A2_c_181_n A2 N_A2_c_182_n N_A2_c_183_n PM_SKY130_FD_SC_LP__O211A_M%A2
x_PM_SKY130_FD_SC_LP__O211A_M%B1 N_B1_M1004_g N_B1_M1008_g N_B1_c_215_n B1 B1
+ N_B1_c_218_n N_B1_c_219_n PM_SKY130_FD_SC_LP__O211A_M%B1
x_PM_SKY130_FD_SC_LP__O211A_M%C1 N_C1_M1006_g N_C1_c_250_n N_C1_M1001_g
+ N_C1_c_252_n C1 C1 N_C1_c_254_n PM_SKY130_FD_SC_LP__O211A_M%C1
x_PM_SKY130_FD_SC_LP__O211A_M%X N_X_M1002_s N_X_M1003_s X X X X X X X X
+ PM_SKY130_FD_SC_LP__O211A_M%X
x_PM_SKY130_FD_SC_LP__O211A_M%VPWR N_VPWR_M1003_d N_VPWR_M1004_d N_VPWR_c_293_n
+ N_VPWR_c_294_n N_VPWR_c_295_n N_VPWR_c_305_n VPWR N_VPWR_c_296_n
+ N_VPWR_c_297_n N_VPWR_c_292_n N_VPWR_c_299_n N_VPWR_c_300_n
+ PM_SKY130_FD_SC_LP__O211A_M%VPWR
x_PM_SKY130_FD_SC_LP__O211A_M%VGND N_VGND_M1002_d N_VGND_M1000_d N_VGND_c_321_n
+ N_VGND_c_322_n N_VGND_c_323_n N_VGND_c_324_n VGND N_VGND_c_325_n
+ N_VGND_c_326_n N_VGND_c_327_n N_VGND_c_328_n PM_SKY130_FD_SC_LP__O211A_M%VGND
x_PM_SKY130_FD_SC_LP__O211A_M%A_217_49# N_A_217_49#_M1000_s N_A_217_49#_M1005_d
+ N_A_217_49#_c_381_n N_A_217_49#_c_365_n N_A_217_49#_c_366_n
+ N_A_217_49#_c_390_n PM_SKY130_FD_SC_LP__O211A_M%A_217_49#
cc_1 VNB N_A_80_60#_M1002_g 0.0285645f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.64
cc_2 VNB N_A_80_60#_c_63_n 0.00192066f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=1.19
cc_3 VNB N_A_80_60#_c_64_n 0.0740293f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=1.19
cc_4 VNB N_A_80_60#_c_65_n 0.0189258f $X=-0.19 $Y=-0.245 $X2=2.54 $Y2=1.675
cc_5 VNB N_A1_M1000_g 0.0304128f $X=-0.19 $Y=-0.245 $X2=2.875 $Y2=1.855
cc_6 VNB N_A1_M1007_g 0.00457477f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_A1_c_140_n 0.0220408f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.64
cc_8 VNB N_A1_c_141_n 0.0200699f $X=-0.19 $Y=-0.245 $X2=0.8 $Y2=1.695
cc_9 VNB N_A1_c_142_n 0.0263365f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=1.675
cc_10 VNB N_A2_M1009_g 0.00439424f $X=-0.19 $Y=-0.245 $X2=2.875 $Y2=1.855
cc_11 VNB N_A2_M1005_g 0.0231562f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A2_c_180_n 0.0206201f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.64
cc_13 VNB N_A2_c_181_n 0.0150924f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.64
cc_14 VNB N_A2_c_182_n 0.0150937f $X=-0.19 $Y=-0.245 $X2=0.8 $Y2=2.065
cc_15 VNB N_A2_c_183_n 0.00975262f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_B1_M1008_g 0.0574094f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_B1_c_215_n 0.00596296f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.64
cc_18 VNB N_C1_M1006_g 0.0267476f $X=-0.19 $Y=-0.245 $X2=2.875 $Y2=1.855
cc_19 VNB N_C1_c_250_n 0.0232771f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_C1_M1001_g 0.0118126f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_C1_c_252_n 0.0249286f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.64
cc_22 VNB C1 0.0367574f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.64
cc_23 VNB N_C1_c_254_n 0.0250755f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB X 0.0488112f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_VPWR_c_292_n 0.143779f $X=-0.19 $Y=-0.245 $X2=2.105 $Y2=1.77
cc_26 VNB N_VGND_c_321_n 0.0117547f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_322_n 0.00313631f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_323_n 0.0193716f $X=-0.19 $Y=-0.245 $X2=0.8 $Y2=2.065
cc_29 VNB N_VGND_c_324_n 0.0036546f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_325_n 0.018332f $X=-0.19 $Y=-0.245 $X2=0.795 $Y2=1.76
cc_31 VNB N_VGND_c_326_n 0.0441542f $X=-0.19 $Y=-0.245 $X2=2.93 $Y2=1.78
cc_32 VNB N_VGND_c_327_n 0.211831f $X=-0.19 $Y=-0.245 $X2=2.625 $Y2=1.78
cc_33 VNB N_VGND_c_328_n 0.00517647f $X=-0.19 $Y=-0.245 $X2=3.015 $Y2=2
cc_34 VNB N_A_217_49#_c_365_n 0.014987f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.64
cc_35 VNB N_A_217_49#_c_366_n 0.00320514f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.64
cc_36 VPB N_A_80_60#_M1003_g 0.0268613f $X=-0.19 $Y=1.655 $X2=0.8 $Y2=2.065
cc_37 VPB N_A_80_60#_c_64_n 0.0134548f $X=-0.19 $Y=1.655 $X2=0.71 $Y2=1.19
cc_38 VPB N_A_80_60#_c_68_n 0.0279224f $X=-0.19 $Y=1.655 $X2=1.895 $Y2=1.76
cc_39 VPB N_A_80_60#_c_69_n 0.00244704f $X=-0.19 $Y=1.655 $X2=0.795 $Y2=1.76
cc_40 VPB N_A_80_60#_c_70_n 0.00550269f $X=-0.19 $Y=1.655 $X2=2.455 $Y2=1.77
cc_41 VPB N_A_80_60#_c_65_n 3.46711e-19 $X=-0.19 $Y=1.655 $X2=2.54 $Y2=1.675
cc_42 VPB N_A_80_60#_c_72_n 0.0101815f $X=-0.19 $Y=1.655 $X2=2.93 $Y2=1.78
cc_43 VPB N_A_80_60#_c_73_n 0.00367204f $X=-0.19 $Y=1.655 $X2=2 $Y2=1.77
cc_44 VPB N_A_80_60#_c_74_n 2.18656e-19 $X=-0.19 $Y=1.655 $X2=2.54 $Y2=1.77
cc_45 VPB N_A1_M1007_g 0.0252069f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_46 VPB N_A2_M1009_g 0.0200155f $X=-0.19 $Y=1.655 $X2=2.875 $Y2=1.855
cc_47 VPB N_B1_M1004_g 0.0154304f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_48 VPB N_B1_c_215_n 0.00595442f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.64
cc_49 VPB N_B1_c_218_n 0.0816439f $X=-0.19 $Y=1.655 $X2=0.71 $Y2=1.675
cc_50 VPB N_B1_c_219_n 0.0265204f $X=-0.19 $Y=1.655 $X2=0.71 $Y2=1.19
cc_51 VPB N_C1_M1001_g 0.0304814f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_52 VPB X 0.0196642f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_53 VPB X 0.0607658f $X=-0.19 $Y=1.655 $X2=3.025 $Y2=1.865
cc_54 VPB N_VPWR_c_293_n 0.0431984f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_55 VPB N_VPWR_c_294_n 0.0346096f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.64
cc_56 VPB N_VPWR_c_295_n 0.0375592f $X=-0.19 $Y=1.655 $X2=0.8 $Y2=1.695
cc_57 VPB N_VPWR_c_296_n 0.0281855f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_58 VPB N_VPWR_c_297_n 0.0215547f $X=-0.19 $Y=1.655 $X2=2.455 $Y2=1.77
cc_59 VPB N_VPWR_c_292_n 0.103787f $X=-0.19 $Y=1.655 $X2=2.105 $Y2=1.77
cc_60 VPB N_VPWR_c_299_n 0.00632158f $X=-0.19 $Y=1.655 $X2=2.93 $Y2=1.78
cc_61 VPB N_VPWR_c_300_n 0.00324402f $X=-0.19 $Y=1.655 $X2=3.025 $Y2=2
cc_62 N_A_80_60#_c_63_n N_A1_M1007_g 4.7509e-19 $X=0.71 $Y=1.19 $X2=0 $Y2=0
cc_63 N_A_80_60#_c_64_n N_A1_M1007_g 0.0181093f $X=0.71 $Y=1.19 $X2=0 $Y2=0
cc_64 N_A_80_60#_c_68_n N_A1_M1007_g 0.0155502f $X=1.895 $Y=1.76 $X2=0 $Y2=0
cc_65 N_A_80_60#_M1002_g N_A1_c_140_n 0.00278227f $X=0.475 $Y=0.64 $X2=0 $Y2=0
cc_66 N_A_80_60#_c_63_n N_A1_c_140_n 0.0019545f $X=0.71 $Y=1.19 $X2=0 $Y2=0
cc_67 N_A_80_60#_c_64_n N_A1_c_140_n 0.0356609f $X=0.71 $Y=1.19 $X2=0 $Y2=0
cc_68 N_A_80_60#_c_68_n N_A1_c_140_n 3.9729e-19 $X=1.895 $Y=1.76 $X2=0 $Y2=0
cc_69 N_A_80_60#_c_68_n N_A1_c_141_n 0.00751645f $X=1.895 $Y=1.76 $X2=0 $Y2=0
cc_70 N_A_80_60#_c_63_n N_A1_c_152_n 0.0218505f $X=0.71 $Y=1.19 $X2=0 $Y2=0
cc_71 N_A_80_60#_c_64_n N_A1_c_152_n 0.00185206f $X=0.71 $Y=1.19 $X2=0 $Y2=0
cc_72 N_A_80_60#_c_68_n N_A1_c_152_n 0.0242882f $X=1.895 $Y=1.76 $X2=0 $Y2=0
cc_73 N_A_80_60#_c_68_n N_A2_M1009_g 0.0124797f $X=1.895 $Y=1.76 $X2=0 $Y2=0
cc_74 N_A_80_60#_c_73_n N_A2_M1009_g 3.10746e-19 $X=2 $Y=1.77 $X2=0 $Y2=0
cc_75 N_A_80_60#_c_68_n N_A2_c_181_n 0.00100329f $X=1.895 $Y=1.76 $X2=0 $Y2=0
cc_76 N_A_80_60#_c_73_n N_A2_c_181_n 0.0042646f $X=2 $Y=1.77 $X2=0 $Y2=0
cc_77 N_A_80_60#_c_68_n N_A2_c_183_n 0.0222421f $X=1.895 $Y=1.76 $X2=0 $Y2=0
cc_78 N_A_80_60#_c_65_n N_A2_c_183_n 0.0199689f $X=2.54 $Y=1.675 $X2=0 $Y2=0
cc_79 N_A_80_60#_c_73_n N_A2_c_183_n 0.0117611f $X=2 $Y=1.77 $X2=0 $Y2=0
cc_80 N_A_80_60#_c_93_p N_B1_M1004_g 0.00527251f $X=2 $Y=2 $X2=0 $Y2=0
cc_81 N_A_80_60#_c_70_n N_B1_M1004_g 0.00925448f $X=2.455 $Y=1.77 $X2=0 $Y2=0
cc_82 N_A_80_60#_c_65_n N_B1_M1008_g 0.0150334f $X=2.54 $Y=1.675 $X2=0 $Y2=0
cc_83 N_A_80_60#_c_70_n N_B1_c_215_n 0.0119379f $X=2.455 $Y=1.77 $X2=0 $Y2=0
cc_84 N_A_80_60#_c_93_p N_B1_c_218_n 8.77563e-19 $X=2 $Y=2 $X2=0 $Y2=0
cc_85 N_A_80_60#_c_70_n N_B1_c_218_n 0.00258754f $X=2.455 $Y=1.77 $X2=0 $Y2=0
cc_86 N_A_80_60#_c_68_n N_B1_c_219_n 0.00883518f $X=1.895 $Y=1.76 $X2=0 $Y2=0
cc_87 N_A_80_60#_c_93_p N_B1_c_219_n 0.0101619f $X=2 $Y=2 $X2=0 $Y2=0
cc_88 N_A_80_60#_c_70_n N_B1_c_219_n 0.0067323f $X=2.455 $Y=1.77 $X2=0 $Y2=0
cc_89 N_A_80_60#_c_65_n N_C1_M1006_g 0.00915069f $X=2.54 $Y=1.675 $X2=0 $Y2=0
cc_90 N_A_80_60#_c_103_p N_C1_M1006_g 0.015655f $X=2.94 $Y=0.495 $X2=0 $Y2=0
cc_91 N_A_80_60#_c_65_n N_C1_M1001_g 0.0037079f $X=2.54 $Y=1.675 $X2=0 $Y2=0
cc_92 N_A_80_60#_c_72_n N_C1_M1001_g 0.0176756f $X=2.93 $Y=1.78 $X2=0 $Y2=0
cc_93 N_A_80_60#_c_74_n N_C1_M1001_g 6.00243e-19 $X=2.54 $Y=1.77 $X2=0 $Y2=0
cc_94 N_A_80_60#_c_72_n N_C1_c_252_n 0.00436867f $X=2.93 $Y=1.78 $X2=0 $Y2=0
cc_95 N_A_80_60#_c_65_n C1 0.0488668f $X=2.54 $Y=1.675 $X2=0 $Y2=0
cc_96 N_A_80_60#_c_72_n C1 0.0247047f $X=2.93 $Y=1.78 $X2=0 $Y2=0
cc_97 N_A_80_60#_c_103_p C1 0.0162922f $X=2.94 $Y=0.495 $X2=0 $Y2=0
cc_98 N_A_80_60#_c_103_p N_C1_c_254_n 0.00159853f $X=2.94 $Y=0.495 $X2=0 $Y2=0
cc_99 N_A_80_60#_M1002_g X 0.0181494f $X=0.475 $Y=0.64 $X2=0 $Y2=0
cc_100 N_A_80_60#_M1003_g X 0.00533094f $X=0.8 $Y=2.065 $X2=0 $Y2=0
cc_101 N_A_80_60#_c_63_n X 0.0407263f $X=0.71 $Y=1.19 $X2=0 $Y2=0
cc_102 N_A_80_60#_c_64_n X 0.0256666f $X=0.71 $Y=1.19 $X2=0 $Y2=0
cc_103 N_A_80_60#_c_69_n X 0.0132301f $X=0.795 $Y=1.76 $X2=0 $Y2=0
cc_104 N_A_80_60#_M1003_g X 0.00808288f $X=0.8 $Y=2.065 $X2=0 $Y2=0
cc_105 N_A_80_60#_c_64_n X 0.00854841f $X=0.71 $Y=1.19 $X2=0 $Y2=0
cc_106 N_A_80_60#_c_69_n X 0.0082536f $X=0.795 $Y=1.76 $X2=0 $Y2=0
cc_107 N_A_80_60#_c_72_n N_VPWR_M1004_d 4.58388e-19 $X=2.93 $Y=1.78 $X2=0 $Y2=0
cc_108 N_A_80_60#_c_74_n N_VPWR_M1004_d 0.00190923f $X=2.54 $Y=1.77 $X2=0 $Y2=0
cc_109 N_A_80_60#_M1003_g N_VPWR_c_293_n 0.00377781f $X=0.8 $Y=2.065 $X2=0 $Y2=0
cc_110 N_A_80_60#_c_68_n N_VPWR_c_293_n 0.0260134f $X=1.895 $Y=1.76 $X2=0 $Y2=0
cc_111 N_A_80_60#_c_72_n N_VPWR_c_305_n 0.00461854f $X=2.93 $Y=1.78 $X2=0 $Y2=0
cc_112 N_A_80_60#_c_74_n N_VPWR_c_305_n 0.0132852f $X=2.54 $Y=1.77 $X2=0 $Y2=0
cc_113 N_A_80_60#_M1002_g N_VGND_c_321_n 0.00509177f $X=0.475 $Y=0.64 $X2=0
+ $Y2=0
cc_114 N_A_80_60#_c_63_n N_VGND_c_321_n 0.00984623f $X=0.71 $Y=1.19 $X2=0 $Y2=0
cc_115 N_A_80_60#_c_64_n N_VGND_c_321_n 0.00206487f $X=0.71 $Y=1.19 $X2=0 $Y2=0
cc_116 N_A_80_60#_M1002_g N_VGND_c_323_n 0.00511809f $X=0.475 $Y=0.64 $X2=0
+ $Y2=0
cc_117 N_A_80_60#_c_103_p N_VGND_c_326_n 0.0229998f $X=2.94 $Y=0.495 $X2=0 $Y2=0
cc_118 N_A_80_60#_M1006_d N_VGND_c_327_n 0.00231826f $X=2.8 $Y=0.245 $X2=0 $Y2=0
cc_119 N_A_80_60#_M1002_g N_VGND_c_327_n 0.00526787f $X=0.475 $Y=0.64 $X2=0
+ $Y2=0
cc_120 N_A_80_60#_c_103_p N_VGND_c_327_n 0.0208199f $X=2.94 $Y=0.495 $X2=0 $Y2=0
cc_121 N_A_80_60#_c_65_n N_A_217_49#_c_365_n 0.0104563f $X=2.54 $Y=1.675 $X2=0
+ $Y2=0
cc_122 N_A_80_60#_M1002_g N_A_217_49#_c_366_n 0.0017257f $X=0.475 $Y=0.64 $X2=0
+ $Y2=0
cc_123 N_A_80_60#_c_65_n A_488_49# 2.78135e-19 $X=2.54 $Y=1.675 $X2=-0.19
+ $Y2=-0.245
cc_124 N_A_80_60#_c_103_p A_488_49# 0.00135771f $X=2.94 $Y=0.495 $X2=-0.19
+ $Y2=-0.245
cc_125 N_A1_M1007_g N_A2_M1009_g 0.0310901f $X=1.425 $Y=2.065 $X2=0 $Y2=0
cc_126 N_A1_M1000_g N_A2_M1005_g 0.0205019f $X=1.425 $Y=0.455 $X2=0 $Y2=0
cc_127 N_A1_c_141_n N_A2_c_181_n 0.0310901f $X=1.292 $Y=1.575 $X2=0 $Y2=0
cc_128 N_A1_c_140_n N_A2_c_182_n 0.0104693f $X=1.292 $Y=1.055 $X2=0 $Y2=0
cc_129 N_A1_c_142_n N_A2_c_182_n 0.0147982f $X=1.25 $Y=1.07 $X2=0 $Y2=0
cc_130 N_A1_c_152_n N_A2_c_182_n 5.07778e-19 $X=1.25 $Y=1.07 $X2=0 $Y2=0
cc_131 N_A1_c_140_n N_A2_c_183_n 4.92301e-19 $X=1.292 $Y=1.055 $X2=0 $Y2=0
cc_132 N_A1_c_141_n N_A2_c_183_n 4.92301e-19 $X=1.292 $Y=1.575 $X2=0 $Y2=0
cc_133 N_A1_c_142_n N_A2_c_183_n 0.00255877f $X=1.25 $Y=1.07 $X2=0 $Y2=0
cc_134 N_A1_c_152_n N_A2_c_183_n 0.039558f $X=1.25 $Y=1.07 $X2=0 $Y2=0
cc_135 N_A1_c_140_n X 6.41024e-19 $X=1.292 $Y=1.055 $X2=0 $Y2=0
cc_136 N_A1_c_152_n X 9.55227e-19 $X=1.25 $Y=1.07 $X2=0 $Y2=0
cc_137 N_A1_M1007_g N_VPWR_c_293_n 0.00908673f $X=1.425 $Y=2.065 $X2=0 $Y2=0
cc_138 N_A1_M1000_g N_VGND_c_321_n 0.00492171f $X=1.425 $Y=0.455 $X2=0 $Y2=0
cc_139 N_A1_M1000_g N_VGND_c_322_n 0.0110152f $X=1.425 $Y=0.455 $X2=0 $Y2=0
cc_140 N_A1_M1000_g N_VGND_c_325_n 0.0034661f $X=1.425 $Y=0.455 $X2=0 $Y2=0
cc_141 N_A1_M1000_g N_VGND_c_327_n 0.0054408f $X=1.425 $Y=0.455 $X2=0 $Y2=0
cc_142 N_A1_M1000_g N_A_217_49#_c_365_n 0.0130444f $X=1.425 $Y=0.455 $X2=0 $Y2=0
cc_143 N_A1_c_140_n N_A_217_49#_c_365_n 0.00155403f $X=1.292 $Y=1.055 $X2=0
+ $Y2=0
cc_144 N_A1_c_141_n N_A_217_49#_c_365_n 3.9729e-19 $X=1.292 $Y=1.575 $X2=0 $Y2=0
cc_145 N_A1_c_152_n N_A_217_49#_c_365_n 0.00862208f $X=1.25 $Y=1.07 $X2=0 $Y2=0
cc_146 N_A1_c_140_n N_A_217_49#_c_366_n 0.00550875f $X=1.292 $Y=1.055 $X2=0
+ $Y2=0
cc_147 N_A1_c_152_n N_A_217_49#_c_366_n 0.0153796f $X=1.25 $Y=1.07 $X2=0 $Y2=0
cc_148 N_A2_M1009_g N_B1_M1008_g 5.63706e-19 $X=1.785 $Y=2.065 $X2=0 $Y2=0
cc_149 N_A2_M1005_g N_B1_M1008_g 0.0204185f $X=1.935 $Y=0.455 $X2=0 $Y2=0
cc_150 N_A2_c_182_n N_B1_M1008_g 0.0331733f $X=1.875 $Y=1.07 $X2=0 $Y2=0
cc_151 N_A2_c_183_n N_B1_M1008_g 0.00182186f $X=1.875 $Y=1.07 $X2=0 $Y2=0
cc_152 N_A2_M1009_g N_B1_c_215_n 0.0194622f $X=1.785 $Y=2.065 $X2=0 $Y2=0
cc_153 N_A2_M1009_g N_B1_c_219_n 0.00540408f $X=1.785 $Y=2.065 $X2=0 $Y2=0
cc_154 N_A2_M1005_g N_VGND_c_322_n 0.00403298f $X=1.935 $Y=0.455 $X2=0 $Y2=0
cc_155 N_A2_M1005_g N_VGND_c_326_n 0.0041676f $X=1.935 $Y=0.455 $X2=0 $Y2=0
cc_156 N_A2_M1005_g N_VGND_c_327_n 0.006026f $X=1.935 $Y=0.455 $X2=0 $Y2=0
cc_157 N_A2_M1005_g N_A_217_49#_c_365_n 0.0115714f $X=1.935 $Y=0.455 $X2=0 $Y2=0
cc_158 N_A2_c_182_n N_A_217_49#_c_365_n 0.00516074f $X=1.875 $Y=1.07 $X2=0 $Y2=0
cc_159 N_A2_c_183_n N_A_217_49#_c_365_n 0.033073f $X=1.875 $Y=1.07 $X2=0 $Y2=0
cc_160 N_B1_M1008_g N_C1_M1006_g 0.0805832f $X=2.365 $Y=0.455 $X2=0 $Y2=0
cc_161 N_B1_M1004_g N_C1_M1001_g 0.0119951f $X=2.325 $Y=2.065 $X2=0 $Y2=0
cc_162 N_B1_M1008_g N_C1_M1001_g 0.00864948f $X=2.365 $Y=0.455 $X2=0 $Y2=0
cc_163 N_B1_c_219_n N_VPWR_c_293_n 0.0289419f $X=2.235 $Y=2.6 $X2=0 $Y2=0
cc_164 N_B1_c_218_n N_VPWR_c_294_n 0.00643118f $X=2.235 $Y=2.6 $X2=0 $Y2=0
cc_165 N_B1_c_219_n N_VPWR_c_294_n 0.0416352f $X=2.235 $Y=2.6 $X2=0 $Y2=0
cc_166 N_B1_M1004_g N_VPWR_c_295_n 0.00706853f $X=2.325 $Y=2.065 $X2=0 $Y2=0
cc_167 N_B1_c_218_n N_VPWR_c_295_n 0.00635852f $X=2.235 $Y=2.6 $X2=0 $Y2=0
cc_168 N_B1_c_219_n N_VPWR_c_295_n 0.0388295f $X=2.235 $Y=2.6 $X2=0 $Y2=0
cc_169 N_B1_c_218_n N_VPWR_c_292_n 0.00853149f $X=2.235 $Y=2.6 $X2=0 $Y2=0
cc_170 N_B1_c_219_n N_VPWR_c_292_n 0.0286705f $X=2.235 $Y=2.6 $X2=0 $Y2=0
cc_171 N_B1_M1008_g N_VGND_c_326_n 0.00575161f $X=2.365 $Y=0.455 $X2=0 $Y2=0
cc_172 N_B1_M1008_g N_VGND_c_327_n 0.0107404f $X=2.365 $Y=0.455 $X2=0 $Y2=0
cc_173 N_B1_M1008_g N_A_217_49#_c_365_n 0.00126505f $X=2.365 $Y=0.455 $X2=0
+ $Y2=0
cc_174 N_C1_M1001_g N_VPWR_c_295_n 0.00779611f $X=2.8 $Y=2.065 $X2=0 $Y2=0
cc_175 N_C1_M1001_g N_VPWR_c_305_n 0.00558458f $X=2.8 $Y=2.065 $X2=0 $Y2=0
cc_176 N_C1_M1006_g N_VGND_c_326_n 0.00366017f $X=2.725 $Y=0.455 $X2=0 $Y2=0
cc_177 N_C1_M1006_g N_VGND_c_327_n 0.00624653f $X=2.725 $Y=0.455 $X2=0 $Y2=0
cc_178 C1 N_VGND_c_327_n 0.00659571f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_179 X N_VPWR_c_293_n 0.0644344f $X=0.24 $Y=2.035 $X2=0 $Y2=0
cc_180 X N_VPWR_c_296_n 0.0195785f $X=0.24 $Y=2.035 $X2=0 $Y2=0
cc_181 X N_VPWR_c_292_n 0.0223074f $X=0.24 $Y=2.035 $X2=0 $Y2=0
cc_182 X N_VGND_c_323_n 0.00871478f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_183 X N_VGND_c_327_n 0.0111671f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_184 N_VGND_c_327_n N_A_217_49#_M1000_s 0.00311927f $X=3.12 $Y=0 $X2=-0.19
+ $Y2=-0.245
cc_185 N_VGND_c_327_n N_A_217_49#_M1005_d 0.00369724f $X=3.12 $Y=0 $X2=0 $Y2=0
cc_186 N_VGND_c_321_n N_A_217_49#_c_381_n 0.0133862f $X=0.69 $Y=0.575 $X2=0
+ $Y2=0
cc_187 N_VGND_c_325_n N_A_217_49#_c_381_n 0.00775693f $X=1.475 $Y=0 $X2=0 $Y2=0
cc_188 N_VGND_c_327_n N_A_217_49#_c_381_n 0.00682159f $X=3.12 $Y=0 $X2=0 $Y2=0
cc_189 N_VGND_M1000_d N_A_217_49#_c_365_n 0.00257168f $X=1.5 $Y=0.245 $X2=0
+ $Y2=0
cc_190 N_VGND_c_322_n N_A_217_49#_c_365_n 0.0194062f $X=1.64 $Y=0.37 $X2=0 $Y2=0
cc_191 N_VGND_c_325_n N_A_217_49#_c_365_n 0.00256318f $X=1.475 $Y=0 $X2=0 $Y2=0
cc_192 N_VGND_c_326_n N_A_217_49#_c_365_n 0.00331392f $X=3.12 $Y=0 $X2=0 $Y2=0
cc_193 N_VGND_c_327_n N_A_217_49#_c_365_n 0.0121173f $X=3.12 $Y=0 $X2=0 $Y2=0
cc_194 N_VGND_c_321_n N_A_217_49#_c_366_n 0.00566601f $X=0.69 $Y=0.575 $X2=0
+ $Y2=0
cc_195 N_VGND_c_326_n N_A_217_49#_c_390_n 0.00781074f $X=3.12 $Y=0 $X2=0 $Y2=0
cc_196 N_VGND_c_327_n N_A_217_49#_c_390_n 0.00755398f $X=3.12 $Y=0 $X2=0 $Y2=0
cc_197 N_VGND_c_327_n A_488_49# 0.00224596f $X=3.12 $Y=0 $X2=-0.19 $Y2=-0.245
