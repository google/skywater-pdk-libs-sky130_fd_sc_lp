* File: sky130_fd_sc_lp__dlxtn_2.spice
* Created: Wed Sep  2 09:48:31 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__dlxtn_2.pex.spice"
.subckt sky130_fd_sc_lp__dlxtn_2  VNB VPB D GATE_N VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* GATE_N	GATE_N
* D	D
* VPB	VPB
* VNB	VNB
MM1007 N_VGND_M1007_d N_D_M1007_g N_A_57_130#_M1007_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0756 AS=0.1113 PD=0.78 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1017 N_A_242_130#_M1017_d N_GATE_N_M1017_g N_VGND_M1007_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1113 AS=0.0756 PD=1.37 PS=0.78 NRD=0 NRS=22.848 M=1 R=2.8
+ SA=75000.7 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1006 N_VGND_M1006_d N_A_242_130#_M1006_g N_A_349_481#_M1006_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75002.6 A=0.063 P=1.14 MULT=1
MM1019 A_669_47# N_A_57_130#_M1019_g N_VGND_M1006_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75002.2 A=0.063 P=1.14 MULT=1
MM1014 N_A_663_481#_M1014_d N_A_242_130#_M1014_g A_669_47# VNB NSHORT L=0.15
+ W=0.42 AD=0.0819 AS=0.0441 PD=0.81 PS=0.63 NRD=31.428 NRS=14.28 M=1 R=2.8
+ SA=75001 SB=75001.8 A=0.063 P=1.14 MULT=1
MM1004 A_849_47# N_A_349_481#_M1004_g N_A_663_481#_M1014_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0819 AS=0.0819 PD=0.81 PS=0.81 NRD=39.996 NRS=0 M=1 R=2.8
+ SA=75001.5 SB=75001.3 A=0.063 P=1.14 MULT=1
MM1008 N_VGND_M1008_d N_A_849_419#_M1008_g A_849_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.0924 AS=0.0819 PD=0.823333 PS=0.81 NRD=32.856 NRS=39.996 M=1 R=2.8
+ SA=75002.1 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1005 N_A_849_419#_M1005_d N_A_663_481#_M1005_g N_VGND_M1008_d VNB NSHORT
+ L=0.15 W=0.84 AD=0.2226 AS=0.1848 PD=2.21 PS=1.64667 NRD=0 NRS=0 M=1 R=5.6
+ SA=75001.4 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1001 N_VGND_M1001_d N_A_849_419#_M1001_g N_Q_M1001_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1009 N_VGND_M1009_d N_A_849_419#_M1009_g N_Q_M1001_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1010 N_VPWR_M1010_d N_D_M1010_g N_A_57_130#_M1010_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0896 AS=0.1696 PD=0.92 PS=1.81 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75000.6 A=0.096 P=1.58 MULT=1
MM1002 N_A_242_130#_M1002_d N_GATE_N_M1002_g N_VPWR_M1010_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1696 AS=0.0896 PD=1.81 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.6 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1011 N_VPWR_M1011_d N_A_242_130#_M1011_g N_A_349_481#_M1011_s VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.2064 AS=0.1696 PD=1.285 PS=1.81 NRD=83.0946 NRS=0 M=1
+ R=4.26667 SA=75000.2 SB=75002.7 A=0.096 P=1.58 MULT=1
MM1015 A_591_481# N_A_57_130#_M1015_g N_VPWR_M1011_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0672 AS=0.2064 PD=0.85 PS=1.285 NRD=15.3857 NRS=29.2348 M=1 R=4.26667
+ SA=75001 SB=75001.9 A=0.096 P=1.58 MULT=1
MM1016 N_A_663_481#_M1016_d N_A_349_481#_M1016_g A_591_481# VPB PHIGHVT L=0.15
+ W=0.64 AD=0.134098 AS=0.0672 PD=1.24377 PS=0.85 NRD=0 NRS=15.3857 M=1
+ R=4.26667 SA=75001.3 SB=75001.6 A=0.096 P=1.58 MULT=1
MM1003 A_771_481# N_A_242_130#_M1003_g N_A_663_481#_M1016_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0819 AS=0.0880019 PD=0.81 PS=0.816226 NRD=65.6601 NRS=53.9386 M=1
+ R=2.8 SA=75001.9 SB=75001.7 A=0.063 P=1.14 MULT=1
MM1013 N_VPWR_M1013_d N_A_849_419#_M1013_g A_771_481# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.150675 AS=0.0819 PD=1.0625 PS=0.81 NRD=276.726 NRS=65.6601 M=1 R=2.8
+ SA=75002.4 SB=75001.2 A=0.063 P=1.14 MULT=1
MM1000 N_A_849_419#_M1000_d N_A_663_481#_M1000_g N_VPWR_M1013_d VPB PHIGHVT
+ L=0.15 W=1.26 AD=0.3339 AS=0.452025 PD=3.05 PS=3.1875 NRD=0 NRS=0 M=1 R=8.4
+ SA=75001.3 SB=75000.2 A=0.189 P=2.82 MULT=1
MM1012 N_VPWR_M1012_d N_A_849_419#_M1012_g N_Q_M1012_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1018 N_VPWR_M1018_d N_A_849_419#_M1018_g N_Q_M1012_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX20_noxref VNB VPB NWDIODE A=14.301 P=19.2
c_137 VPB 0 2.4855e-20 $X=0 $Y=3.085
*
.include "sky130_fd_sc_lp__dlxtn_2.pxi.spice"
*
.ends
*
*
