# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__invlp_4
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__invlp_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.320000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  2.520000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.385000 1.345000 4.095000 1.675000 ;
        RECT 1.565000 1.675000 2.755000 1.780000 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  1.411200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605000 1.180000 1.215000 1.410000 ;
        RECT 1.045000 1.005000 3.235000 1.175000 ;
        RECT 1.045000 1.175000 1.215000 1.180000 ;
        RECT 1.045000 1.410000 1.215000 1.950000 ;
        RECT 1.045000 1.950000 3.255000 2.120000 ;
        RECT 1.925000 2.120000 2.255000 2.735000 ;
        RECT 2.055000 0.595000 2.225000 1.005000 ;
        RECT 2.905000 0.595000 3.235000 1.005000 ;
        RECT 2.925000 1.845000 3.255000 1.950000 ;
        RECT 2.925000 2.120000 3.255000 2.735000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 4.320000 0.085000 ;
        RECT 0.115000  0.085000 0.365000 1.125000 ;
        RECT 1.045000  0.085000 1.375000 0.495000 ;
        RECT 3.915000  0.085000 4.165000 1.125000 ;
      LAYER mcon ;
        RECT 0.155000 -0.085000 0.325000 0.085000 ;
        RECT 0.635000 -0.085000 0.805000 0.085000 ;
        RECT 1.115000 -0.085000 1.285000 0.085000 ;
        RECT 1.595000 -0.085000 1.765000 0.085000 ;
        RECT 2.075000 -0.085000 2.245000 0.085000 ;
        RECT 2.555000 -0.085000 2.725000 0.085000 ;
        RECT 3.035000 -0.085000 3.205000 0.085000 ;
        RECT 3.515000 -0.085000 3.685000 0.085000 ;
        RECT 3.995000 -0.085000 4.165000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.320000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.245000 4.320000 3.415000 ;
        RECT 0.135000 1.815000 0.385000 3.245000 ;
        RECT 0.995000 2.630000 1.245000 3.245000 ;
        RECT 3.855000 1.845000 4.185000 3.245000 ;
      LAYER mcon ;
        RECT 0.155000 3.245000 0.325000 3.415000 ;
        RECT 0.635000 3.245000 0.805000 3.415000 ;
        RECT 1.115000 3.245000 1.285000 3.415000 ;
        RECT 1.595000 3.245000 1.765000 3.415000 ;
        RECT 2.075000 3.245000 2.245000 3.415000 ;
        RECT 2.555000 3.245000 2.725000 3.415000 ;
        RECT 3.035000 3.245000 3.205000 3.415000 ;
        RECT 3.515000 3.245000 3.685000 3.415000 ;
        RECT 3.995000 3.245000 4.165000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 4.320000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.545000 0.255000 0.875000 0.665000 ;
      RECT 0.545000 0.665000 1.875000 0.835000 ;
      RECT 0.545000 0.835000 0.875000 1.010000 ;
      RECT 0.565000 1.815000 0.815000 2.290000 ;
      RECT 0.565000 2.290000 1.755000 2.460000 ;
      RECT 0.565000 2.460000 0.815000 3.075000 ;
      RECT 1.425000 2.460000 1.755000 2.905000 ;
      RECT 1.425000 2.905000 3.685000 3.075000 ;
      RECT 1.545000 0.255000 3.735000 0.425000 ;
      RECT 1.545000 0.425000 1.875000 0.665000 ;
      RECT 2.405000 0.425000 2.735000 0.835000 ;
      RECT 2.425000 2.290000 2.755000 2.905000 ;
      RECT 3.405000 0.425000 3.735000 1.125000 ;
      RECT 3.435000 1.845000 3.685000 2.905000 ;
  END
END sky130_fd_sc_lp__invlp_4
