* File: sky130_fd_sc_lp__a311oi_lp.spice
* Created: Wed Sep  2 09:25:59 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__a311oi_lp.pex.spice"
.subckt sky130_fd_sc_lp__a311oi_lp  VNB VPB A1 A2 A3 B1 C1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* C1	C1
* B1	B1
* A3	A3
* A2	A2
* A1	A1
* VPB	VPB
* VNB	VNB
MM1006 A_116_47# N_A1_M1006_g N_Y_M1006_s VNB NSHORT L=0.15 W=0.42 AD=0.0504
+ AS=0.1197 PD=0.66 PS=1.41 NRD=18.564 NRS=0 M=1 R=2.8 SA=75000.2 SB=75002.6
+ A=0.063 P=1.14 MULT=1
MM1003 A_194_47# N_A2_M1003_g A_116_47# VNB NSHORT L=0.15 W=0.42 AD=0.0504
+ AS=0.0504 PD=0.66 PS=0.66 NRD=18.564 NRS=18.564 M=1 R=2.8 SA=75000.6
+ SB=75002.2 A=0.063 P=1.14 MULT=1
MM1002 N_VGND_M1002_d N_A3_M1002_g A_194_47# VNB NSHORT L=0.15 W=0.42 AD=0.0588
+ AS=0.0504 PD=0.7 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75001 SB=75001.8
+ A=0.063 P=1.14 MULT=1
MM1009 A_358_47# N_B1_M1009_g N_VGND_M1002_d VNB NSHORT L=0.15 W=0.42 AD=0.0441
+ AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75001.4 SB=75001.4
+ A=0.063 P=1.14 MULT=1
MM1007 N_Y_M1007_d N_B1_M1007_g A_358_47# VNB NSHORT L=0.15 W=0.42 AD=0.0588
+ AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.8 SB=75001 A=0.063
+ P=1.14 MULT=1
MM1010 A_516_47# N_C1_M1010_g N_Y_M1007_d VNB NSHORT L=0.15 W=0.42 AD=0.0441
+ AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75002.2 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1011 N_VGND_M1011_d N_C1_M1011_g A_516_47# VNB NSHORT L=0.15 W=0.42 AD=0.1197
+ AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75002.6 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1001 N_A_134_409#_M1001_d N_A1_M1001_g N_VPWR_M1001_s VPB PHIGHVT L=0.25 W=1
+ AD=0.14 AS=0.285 PD=1.28 PS=2.57 NRD=0 NRS=0 M=1 R=4 SA=125000 SB=125002
+ A=0.25 P=2.5 MULT=1
MM1005 N_VPWR_M1005_d N_A2_M1005_g N_A_134_409#_M1001_d VPB PHIGHVT L=0.25 W=1
+ AD=0.15 AS=0.14 PD=1.3 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125001 SB=125002 A=0.25
+ P=2.5 MULT=1
MM1000 N_A_134_409#_M1000_d N_A3_M1000_g N_VPWR_M1005_d VPB PHIGHVT L=0.25 W=1
+ AD=0.14 AS=0.15 PD=1.28 PS=1.3 NRD=0 NRS=3.9203 M=1 R=4 SA=125001 SB=125001
+ A=0.25 P=2.5 MULT=1
MM1008 A_456_409# N_B1_M1008_g N_A_134_409#_M1000_d VPB PHIGHVT L=0.25 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=16.7253 NRS=0 M=1 R=4 SA=125002 SB=125001
+ A=0.25 P=2.5 MULT=1
MM1004 N_Y_M1004_d N_C1_M1004_g A_456_409# VPB PHIGHVT L=0.25 W=1 AD=0.285
+ AS=0.14 PD=2.57 PS=1.28 NRD=0 NRS=16.7253 M=1 R=4 SA=125002 SB=125000 A=0.25
+ P=2.5 MULT=1
DX12_noxref VNB VPB NWDIODE A=6.9751 P=11.21
*
.include "sky130_fd_sc_lp__a311oi_lp.pxi.spice"
*
.ends
*
*
