* File: sky130_fd_sc_lp__o221ai_0.pex.spice
* Created: Fri Aug 28 11:08:13 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O221AI_0%C1 3 7 9 12 13
r34 12 15 45.3519 $w=3.85e-07 $l=1.65e-07 $layer=POLY_cond $X=0.447 $Y=2.015
+ $X2=0.447 $Y2=2.18
r35 12 14 45.3519 $w=3.85e-07 $l=1.65e-07 $layer=POLY_cond $X=0.447 $Y=2.015
+ $X2=0.447 $Y2=1.85
r36 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.42
+ $Y=2.015 $X2=0.42 $Y2=2.015
r37 9 13 9.01912 $w=2.28e-07 $l=1.8e-07 $layer=LI1_cond $X=0.24 $Y=2.035
+ $X2=0.42 $Y2=2.035
r38 7 15 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.565 $Y=2.66
+ $X2=0.565 $Y2=2.18
r39 3 14 720.436 $w=1.5e-07 $l=1.405e-06 $layer=POLY_cond $X=0.475 $Y=0.445
+ $X2=0.475 $Y2=1.85
.ends

.subckt PM_SKY130_FD_SC_LP__O221AI_0%B1 3 7 9 10 11 16 19 24
c50 24 0 1.72602e-19 $X=1.197 $Y=1.41
c51 16 0 1.31003e-19 $X=0.995 $Y=1.3
r52 17 19 6.1 $w=1.98e-07 $l=1.1e-07 $layer=LI1_cond $X=0.995 $Y=1.31 $X2=1.105
+ $Y2=1.31
r53 16 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.995 $Y=1.3
+ $X2=0.995 $Y2=1.135
r54 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.995
+ $Y=1.3 $X2=0.995 $Y2=1.3
r55 11 24 15.2875 $w=1.83e-07 $l=2.55e-07 $layer=LI1_cond $X=1.197 $Y=1.665
+ $X2=1.197 $Y2=1.41
r56 10 24 3.55727 $w=1.85e-07 $l=1e-07 $layer=LI1_cond $X=1.197 $Y=1.31
+ $X2=1.197 $Y2=1.41
r57 10 19 3.27269 $w=2e-07 $l=9.2e-08 $layer=LI1_cond $X=1.197 $Y=1.31 $X2=1.105
+ $Y2=1.31
r58 9 17 15.25 $w=1.98e-07 $l=2.75e-07 $layer=LI1_cond $X=0.72 $Y=1.31 $X2=0.995
+ $Y2=1.31
r59 5 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.995 $Y=1.465
+ $X2=0.995 $Y2=1.3
r60 5 7 612.755 $w=1.5e-07 $l=1.195e-06 $layer=POLY_cond $X=0.995 $Y=1.465
+ $X2=0.995 $Y2=2.66
r61 3 18 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=0.905 $Y=0.445
+ $X2=0.905 $Y2=1.135
.ends

.subckt PM_SKY130_FD_SC_LP__O221AI_0%B2 3 7 13 15 16 17 18 19 20 21 30 35 37 39
+ 50
r58 35 37 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.085 $Y=2.015
+ $X2=3.085 $Y2=1.85
r59 30 33 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.445 $Y=2.015
+ $X2=1.445 $Y2=2.18
r60 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.445
+ $Y=2.015 $X2=1.445 $Y2=2.015
r61 20 21 13.3251 $w=3.18e-07 $l=3.7e-07 $layer=LI1_cond $X=3.115 $Y=2.405
+ $X2=3.115 $Y2=2.775
r62 20 50 9.54367 $w=3.18e-07 $l=2.65e-07 $layer=LI1_cond $X=3.115 $Y=2.405
+ $X2=3.115 $Y2=2.14
r63 19 50 2.855 $w=3.2e-07 $l=1.05e-07 $layer=LI1_cond $X=3.115 $Y=2.035
+ $X2=3.115 $Y2=2.14
r64 19 39 4.35048 $w=2.1e-07 $l=1.6e-07 $layer=LI1_cond $X=3.115 $Y=2.035
+ $X2=2.955 $Y2=2.035
r65 19 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.085
+ $Y=2.015 $X2=3.085 $Y2=2.015
r66 18 39 16.6364 $w=2.08e-07 $l=3.15e-07 $layer=LI1_cond $X=2.64 $Y=2.035
+ $X2=2.955 $Y2=2.035
r67 17 18 25.3506 $w=2.08e-07 $l=4.8e-07 $layer=LI1_cond $X=2.16 $Y=2.035
+ $X2=2.64 $Y2=2.035
r68 16 17 25.3506 $w=2.08e-07 $l=4.8e-07 $layer=LI1_cond $X=1.68 $Y=2.035
+ $X2=2.16 $Y2=2.035
r69 16 31 12.4113 $w=2.08e-07 $l=2.35e-07 $layer=LI1_cond $X=1.68 $Y=2.035
+ $X2=1.445 $Y2=2.035
r70 15 31 12.9394 $w=2.08e-07 $l=2.45e-07 $layer=LI1_cond $X=1.2 $Y=2.035
+ $X2=1.445 $Y2=2.035
r71 11 13 153.83 $w=1.5e-07 $l=3e-07 $layer=POLY_cond $X=2.695 $Y=1.135
+ $X2=2.995 $Y2=1.135
r72 9 13 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.995 $Y=1.21
+ $X2=2.995 $Y2=1.135
r73 9 37 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=2.995 $Y=1.21
+ $X2=2.995 $Y2=1.85
r74 5 11 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.695 $Y=1.06
+ $X2=2.695 $Y2=1.135
r75 5 7 315.351 $w=1.5e-07 $l=6.15e-07 $layer=POLY_cond $X=2.695 $Y=1.06
+ $X2=2.695 $Y2=0.445
r76 3 33 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.355 $Y=2.66
+ $X2=1.355 $Y2=2.18
.ends

.subckt PM_SKY130_FD_SC_LP__O221AI_0%A2 1 3 5 8 12 14 15 23
c49 23 0 1.6655e-19 $X=1.895 $Y=1.475
c50 15 0 1.31003e-19 $X=2.16 $Y=1.665
c51 12 0 1.72602e-19 $X=1.445 $Y=0.85
c52 8 0 1.46389e-19 $X=1.895 $Y=2.66
r53 21 23 33.2236 $w=3.3e-07 $l=1.9e-07 $layer=POLY_cond $X=1.705 $Y=1.475
+ $X2=1.895 $Y2=1.475
r54 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.705
+ $Y=1.475 $X2=1.705 $Y2=1.475
r55 18 21 45.4639 $w=3.3e-07 $l=2.6e-07 $layer=POLY_cond $X=1.445 $Y=1.475
+ $X2=1.705 $Y2=1.475
r56 15 22 12.0937 $w=4.48e-07 $l=4.55e-07 $layer=LI1_cond $X=2.16 $Y=1.535
+ $X2=1.705 $Y2=1.535
r57 14 22 0.664488 $w=4.48e-07 $l=2.5e-08 $layer=LI1_cond $X=1.68 $Y=1.535
+ $X2=1.705 $Y2=1.535
r58 10 12 56.4043 $w=1.5e-07 $l=1.1e-07 $layer=POLY_cond $X=1.335 $Y=0.85
+ $X2=1.445 $Y2=0.85
r59 6 23 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.895 $Y=1.64
+ $X2=1.895 $Y2=1.475
r60 6 8 523.021 $w=1.5e-07 $l=1.02e-06 $layer=POLY_cond $X=1.895 $Y=1.64
+ $X2=1.895 $Y2=2.66
r61 5 18 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.445 $Y=1.31
+ $X2=1.445 $Y2=1.475
r62 4 12 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.445 $Y=0.925
+ $X2=1.445 $Y2=0.85
r63 4 5 197.415 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=1.445 $Y=0.925
+ $X2=1.445 $Y2=1.31
r64 1 10 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.335 $Y=0.775
+ $X2=1.335 $Y2=0.85
r65 1 3 106.04 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=1.335 $Y=0.775
+ $X2=1.335 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__O221AI_0%A1 1 2 5 9 12 13 20
c42 13 0 1.6655e-19 $X=3.12 $Y=1.665
r43 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.545
+ $Y=1.585 $X2=2.545 $Y2=1.585
r44 18 20 49.8355 $w=3.3e-07 $l=2.85e-07 $layer=POLY_cond $X=2.26 $Y=1.585
+ $X2=2.545 $Y2=1.585
r45 16 18 0.874306 $w=3.3e-07 $l=5e-09 $layer=POLY_cond $X=2.255 $Y=1.585
+ $X2=2.26 $Y2=1.585
r46 12 13 16.5126 $w=3.33e-07 $l=4.8e-07 $layer=LI1_cond $X=2.64 $Y=1.587
+ $X2=3.12 $Y2=1.587
r47 12 21 3.26812 $w=3.33e-07 $l=9.5e-08 $layer=LI1_cond $X=2.64 $Y=1.587
+ $X2=2.545 $Y2=1.587
r48 9 11 335.862 $w=1.5e-07 $l=6.55e-07 $layer=POLY_cond $X=2.265 $Y=0.445
+ $X2=2.265 $Y2=1.1
r49 3 16 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.255 $Y=1.75
+ $X2=2.255 $Y2=1.585
r50 3 5 466.617 $w=1.5e-07 $l=9.1e-07 $layer=POLY_cond $X=2.255 $Y=1.75
+ $X2=2.255 $Y2=2.66
r51 2 18 19.6935 $w=1.6e-07 $l=1.65e-07 $layer=POLY_cond $X=2.26 $Y=1.42
+ $X2=2.26 $Y2=1.585
r52 1 11 37.4638 $w=1.6e-07 $l=8e-08 $layer=POLY_cond $X=2.26 $Y=1.18 $X2=2.26
+ $Y2=1.1
r53 1 2 111.231 $w=1.6e-07 $l=2.4e-07 $layer=POLY_cond $X=2.26 $Y=1.18 $X2=2.26
+ $Y2=1.42
.ends

.subckt PM_SKY130_FD_SC_LP__O221AI_0%Y 1 2 3 12 16 17 18 21 23 25 26 27 28 33
c66 28 0 1.46389e-19 $X=1.68 $Y=2.775
r67 27 33 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.63 $Y=2.405
+ $X2=1.465 $Y2=2.405
r68 27 28 8.20134 $w=4.98e-07 $l=2.85e-07 $layer=LI1_cond $X=1.63 $Y=2.49
+ $X2=1.63 $Y2=2.775
r69 26 33 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=1.2 $Y=2.405
+ $X2=1.465 $Y2=2.405
r70 24 26 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.935 $Y=2.405
+ $X2=1.2 $Y2=2.405
r71 24 25 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.935 $Y=2.405
+ $X2=0.85 $Y2=2.405
r72 21 25 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.85 $Y=2.32 $X2=0.85
+ $Y2=2.405
r73 20 21 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=0.85 $Y=1.75
+ $X2=0.85 $Y2=2.32
r74 19 23 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.445 $Y=2.405
+ $X2=0.315 $Y2=2.405
r75 18 25 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.765 $Y=2.405
+ $X2=0.85 $Y2=2.405
r76 18 19 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=0.765 $Y=2.405
+ $X2=0.445 $Y2=2.405
r77 16 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.765 $Y=1.665
+ $X2=0.85 $Y2=1.75
r78 16 17 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=0.765 $Y=1.665
+ $X2=0.365 $Y2=1.665
r79 10 17 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=0.23 $Y=1.58
+ $X2=0.365 $Y2=1.665
r80 10 12 48.4453 $w=2.68e-07 $l=1.135e-06 $layer=LI1_cond $X=0.23 $Y=1.58
+ $X2=0.23 $Y2=0.445
r81 3 27 300 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_PDIFF $count=2 $X=1.43
+ $Y=2.34 $X2=1.63 $Y2=2.485
r82 2 23 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.225
+ $Y=2.34 $X2=0.35 $Y2=2.485
r83 1 12 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__O221AI_0%VPWR 1 2 9 13 16 17 18 20 33 34 37
r43 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r44 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r45 31 34 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r46 30 31 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r47 28 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r48 27 30 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=3.33 $X2=2.16
+ $Y2=3.33
r49 27 28 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r50 25 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.945 $Y=3.33
+ $X2=0.78 $Y2=3.33
r51 25 27 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.945 $Y=3.33
+ $X2=1.2 $Y2=3.33
r52 23 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r53 22 23 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r54 20 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.615 $Y=3.33
+ $X2=0.78 $Y2=3.33
r55 20 22 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.615 $Y=3.33
+ $X2=0.24 $Y2=3.33
r56 18 31 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r57 18 28 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r58 16 30 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=2.365 $Y=3.33
+ $X2=2.16 $Y2=3.33
r59 16 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.365 $Y=3.33
+ $X2=2.53 $Y2=3.33
r60 15 33 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=2.695 $Y=3.33
+ $X2=3.12 $Y2=3.33
r61 15 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.695 $Y=3.33
+ $X2=2.53 $Y2=3.33
r62 11 17 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.53 $Y=3.245
+ $X2=2.53 $Y2=3.33
r63 11 13 26.1919 $w=3.28e-07 $l=7.5e-07 $layer=LI1_cond $X=2.53 $Y=3.245
+ $X2=2.53 $Y2=2.495
r64 7 37 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.78 $Y=3.245 $X2=0.78
+ $Y2=3.33
r65 7 9 16.0644 $w=3.28e-07 $l=4.6e-07 $layer=LI1_cond $X=0.78 $Y=3.245 $X2=0.78
+ $Y2=2.785
r66 2 13 300 $w=1.7e-07 $l=2.66458e-07 $layer=licon1_PDIFF $count=2 $X=2.33
+ $Y=2.34 $X2=2.53 $Y2=2.495
r67 1 9 600 $w=1.7e-07 $l=5.10221e-07 $layer=licon1_PDIFF $count=1 $X=0.64
+ $Y=2.34 $X2=0.78 $Y2=2.785
.ends

.subckt PM_SKY130_FD_SC_LP__O221AI_0%A_110_47# 1 2 8 10 11 15 18 21 22
r44 21 22 10.774 $w=1.73e-07 $l=1.7e-07 $layer=LI1_cond $X=1.465 $Y=0.957
+ $X2=1.635 $Y2=0.957
r45 18 20 8.71257 $w=2.88e-07 $l=1.7e-07 $layer=LI1_cond $X=0.69 $Y=0.445
+ $X2=0.69 $Y2=0.615
r46 13 15 16.2476 $w=3.03e-07 $l=4.3e-07 $layer=LI1_cond $X=2.922 $Y=0.875
+ $X2=2.922 $Y2=0.445
r47 11 13 7.55824 $w=1.7e-07 $l=1.898e-07 $layer=LI1_cond $X=2.77 $Y=0.96
+ $X2=2.922 $Y2=0.875
r48 11 22 74.0481 $w=1.68e-07 $l=1.135e-06 $layer=LI1_cond $X=2.77 $Y=0.96
+ $X2=1.635 $Y2=0.96
r49 10 21 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=0.715 $Y=0.955
+ $X2=1.465 $Y2=0.955
r50 8 10 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.63 $Y=0.87
+ $X2=0.715 $Y2=0.955
r51 8 20 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.63 $Y=0.87
+ $X2=0.63 $Y2=0.615
r52 2 15 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.77
+ $Y=0.235 $X2=2.91 $Y2=0.445
r53 1 18 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.235 $X2=0.69 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__O221AI_0%A_196_47# 1 2 7 10 15
r27 10 12 6.99698 $w=2.78e-07 $l=1.7e-07 $layer=LI1_cond $X=1.145 $Y=0.445
+ $X2=1.145 $Y2=0.615
r28 8 12 3.65648 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=1.285 $Y=0.615
+ $X2=1.145 $Y2=0.615
r29 7 15 6.87422 $w=2.83e-07 $l=1.7e-07 $layer=LI1_cond $X=2.457 $Y=0.615
+ $X2=2.457 $Y2=0.445
r30 7 8 67.1979 $w=1.68e-07 $l=1.03e-06 $layer=LI1_cond $X=2.315 $Y=0.615
+ $X2=1.285 $Y2=0.615
r31 2 15 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.34
+ $Y=0.235 $X2=2.48 $Y2=0.445
r32 1 10 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.98
+ $Y=0.235 $X2=1.12 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__O221AI_0%VGND 1 4 19 20 25 28
r36 27 28 8.86124 $w=4.43e-07 $l=1.65e-07 $layer=LI1_cond $X=1.97 $Y=0.137
+ $X2=2.135 $Y2=0.137
r37 23 27 7.5103 $w=4.43e-07 $l=2.9e-07 $layer=LI1_cond $X=1.68 $Y=0.137
+ $X2=1.97 $Y2=0.137
r38 23 25 10.1561 $w=4.43e-07 $l=2.15e-07 $layer=LI1_cond $X=1.68 $Y=0.137
+ $X2=1.465 $Y2=0.137
r39 19 20 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r40 17 20 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r41 16 19 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r42 16 28 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=2.16 $Y=0 $X2=2.135
+ $Y2=0
r43 16 17 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r44 12 25 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=1.2 $Y=0 $X2=1.465
+ $Y2=0
r45 12 13 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r46 9 13 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r47 8 12 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r48 8 9 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r49 4 17 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r50 4 13 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r51 4 23 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r52 1 27 91 $w=1.7e-07 $l=5.79655e-07 $layer=licon1_NDIFF $count=2 $X=1.41
+ $Y=0.235 $X2=1.97 $Y2=0.275
.ends

