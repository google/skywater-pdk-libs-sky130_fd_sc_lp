* File: sky130_fd_sc_lp__srdlrtp_1.spice
* Created: Fri Aug 28 11:33:01 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__srdlrtp_1.pex.spice"
.subckt sky130_fd_sc_lp__srdlrtp_1  VNB VPB D RESET_B GATE SLEEP_B VPWR KAPWR Q
+ VGND
* 
* VGND	VGND
* Q	Q
* KAPWR	KAPWR
* VPWR	VPWR
* SLEEP_B	SLEEP_B
* GATE	GATE
* RESET_B	RESET_B
* D	D
* VPB	VPB
* VNB	VNB
MM1005 A_114_97# N_D_M1005_g N_A_27_97#_M1005_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1197 PD=0.63 PS=1.41 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75003.9 A=0.063 P=1.14 MULT=1
MM1030 N_VGND_M1030_d N_RESET_B_M1030_g A_114_97# VNB NSHORT L=0.15 W=0.42
+ AD=0.0672 AS=0.0441 PD=0.74 PS=0.63 NRD=11.424 NRS=14.28 M=1 R=2.8 SA=75000.6
+ SB=75003.5 A=0.063 P=1.14 MULT=1
MM1025 N_A_280_97#_M1025_d N_A_27_97#_M1025_g N_VGND_M1030_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0588 AS=0.0672 PD=0.7 PS=0.74 NRD=0 NRS=0 M=1 R=2.8 SA=75001
+ SB=75003 A=0.063 P=1.14 MULT=1
MM1002 A_366_97# N_A_336_71#_M1002_g N_A_280_97#_M1025_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75001.5
+ SB=75002.6 A=0.063 P=1.14 MULT=1
MM1010 N_A_438_97#_M1010_d N_A_336_71#_M1010_g A_366_97# VNB NSHORT L=0.15
+ W=0.42 AD=0.1071 AS=0.0441 PD=0.93 PS=0.63 NRD=32.856 NRS=14.28 M=1 R=2.8
+ SA=75001.8 SB=75002.2 A=0.063 P=1.14 MULT=1
MM1024 A_570_97# N_A_393_335#_M1024_g N_A_438_97#_M1010_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.1071 PD=0.63 PS=0.93 NRD=14.28 NRS=32.856 M=1 R=2.8
+ SA=75002.5 SB=75001.6 A=0.063 P=1.14 MULT=1
MM1026 A_642_97# N_A_612_71#_M1026_g A_570_97# VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0441 PD=0.63 PS=0.63 NRD=14.28 NRS=14.28 M=1 R=2.8 SA=75002.8
+ SB=75001.2 A=0.063 P=1.14 MULT=1
MM1015 N_VGND_M1015_d N_A_612_71#_M1015_g A_642_97# VNB NSHORT L=0.15 W=0.42
+ AD=0.15785 AS=0.0441 PD=1.28 PS=0.63 NRD=91.656 NRS=14.28 M=1 R=2.8 SA=75003.2
+ SB=75000.9 A=0.063 P=1.14 MULT=1
MM1006 N_A_336_71#_M1006_d N_A_393_335#_M1006_g N_VGND_M1015_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1197 AS=0.15785 PD=1.41 PS=1.28 NRD=0 NRS=91.656 M=1 R=2.8
+ SA=75003.9 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1019 A_1069_97# N_GATE_M1019_g N_A_393_335#_M1019_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.1197 PD=0.66 PS=1.41 NRD=18.564 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.1 A=0.063 P=1.14 MULT=1
MM1020 A_1147_97# N_SLEEP_B_M1020_g A_1069_97# VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0504 PD=0.63 PS=0.66 NRD=14.28 NRS=18.564 M=1 R=2.8 SA=75000.6
+ SB=75001.7 A=0.063 P=1.14 MULT=1
MM1001 N_VGND_M1001_d N_SLEEP_B_M1001_g A_1147_97# VNB NSHORT L=0.15 W=0.42
+ AD=0.123675 AS=0.0441 PD=1.06 PS=0.63 NRD=24.276 NRS=14.28 M=1 R=2.8 SA=75001
+ SB=75001.3 A=0.063 P=1.14 MULT=1
MM1003 A_1344_97# N_SLEEP_B_M1003_g N_VGND_M1001_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.123675 PD=0.63 PS=1.06 NRD=14.28 NRS=34.284 M=1 R=2.8
+ SA=75001.6 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1029 N_A_1324_394#_M1029_d N_SLEEP_B_M1029_g A_1344_97# VNB NSHORT L=0.15
+ W=0.42 AD=0.168 AS=0.0441 PD=1.64 PS=0.63 NRD=32.856 NRS=14.28 M=1 R=2.8
+ SA=75001.9 SB=75000.3 A=0.063 P=1.14 MULT=1
MM1007 N_VGND_M1007_d N_A_1324_394#_M1007_g N_A_1624_47#_M1007_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.1069 AS=0.1197 PD=0.96 PS=1.41 NRD=24.276 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.6 A=0.063 P=1.14 MULT=1
MM1022 N_A_1624_47#_M1022_d N_RESET_B_M1022_g N_VGND_M1007_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0609 AS=0.1069 PD=0.71 PS=0.96 NRD=1.428 NRS=24.276 M=1 R=2.8
+ SA=75000.8 SB=75001 A=0.063 P=1.14 MULT=1
MM1011 A_1917_47# N_A_438_97#_M1011_g N_A_1624_47#_M1022_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.0609 PD=0.63 PS=0.71 NRD=14.28 NRS=1.428 M=1 R=2.8
+ SA=75001.2 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1013 N_A_612_71#_M1013_d N_A_438_97#_M1013_g A_1917_47# VNB NSHORT L=0.15
+ W=0.42 AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8
+ SA=75001.6 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1017 N_VGND_M1017_d N_A_438_97#_M1017_g N_A_2120_55#_M1017_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0952 AS=0.1197 PD=0.823333 PS=1.41 NRD=32.856 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1016 N_Q_M1016_d N_A_2120_55#_M1016_g N_VGND_M1017_d VNB NSHORT L=0.15 W=0.84
+ AD=0.2394 AS=0.1904 PD=2.25 PS=1.64667 NRD=0 NRS=0 M=1 R=5.6 SA=75000.5
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1032 N_A_27_97#_M1032_d N_D_M1032_g N_VPWR_M1032_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.112 AS=0.1824 PD=0.99 PS=1.85 NRD=21.5321 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75002.1 A=0.096 P=1.58 MULT=1
MM1031 N_VPWR_M1031_d N_RESET_B_M1031_g N_A_27_97#_M1032_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1488 AS=0.112 PD=1.105 PS=0.99 NRD=35.3812 NRS=0 M=1 R=4.26667
+ SA=75000.7 SB=75001.6 A=0.096 P=1.58 MULT=1
MM1008 N_A_280_97#_M1008_d N_A_27_97#_M1008_g N_VPWR_M1031_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.0896 AS=0.1488 PD=0.92 PS=1.105 NRD=0 NRS=21.5321 M=1 R=4.26667
+ SA=75001.3 SB=75001 A=0.096 P=1.58 MULT=1
MM1018 A_423_487# N_A_393_335#_M1018_g N_A_280_97#_M1008_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.0672 AS=0.0896 PD=0.85 PS=0.92 NRD=15.3857 NRS=0 M=1 R=4.26667
+ SA=75001.8 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1021 N_A_438_97#_M1021_d N_A_393_335#_M1021_g A_423_487# VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1824 AS=0.0672 PD=1.85 PS=0.85 NRD=0 NRS=15.3857 M=1 R=4.26667
+ SA=75002.1 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1033 N_VPWR_M1033_d N_A_393_335#_M1033_g N_A_336_71#_M1033_s VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.4358 AS=0.26615 PD=3.32 PS=2.15 NRD=192.666 NRS=35.3812 M=1
+ R=4.26667 SA=75000.3 SB=75000.3 A=0.096 P=1.58 MULT=1
MM1000 N_A_393_335#_M1000_d N_GATE_M1000_g N_KAPWR_M1000_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.27195 AS=0.1824 PD=1.9 PS=1.85 NRD=113.866 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75001.6 A=0.096 P=1.58 MULT=1
MM1035 N_KAPWR_M1035_d N_SLEEP_B_M1035_g N_A_393_335#_M1000_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.138693 AS=0.27195 PD=1.08878 PS=1.9 NRD=35.3812 NRS=113.866 M=1
+ R=4.26667 SA=75000.9 SB=75001 A=0.096 P=1.58 MULT=1
MM1023 N_A_1324_394#_M1023_d N_SLEEP_B_M1023_g N_KAPWR_M1035_d VPB PHIGHVT
+ L=0.25 W=1 AD=0.5131 AS=0.216707 PD=3.58 PS=1.70122 NRD=90.226 NRS=0 M=1 R=4
+ SA=125001 SB=125000 A=0.25 P=2.5 MULT=1
MM1027 A_1565_419# N_A_336_71#_M1027_g N_A_438_97#_M1027_s VPB PHIGHVT L=0.25
+ W=1 AD=0.105 AS=0.285 PD=1.21 PS=2.57 NRD=9.8303 NRS=0 M=1 R=4 SA=125000
+ SB=125002 A=0.25 P=2.5 MULT=1
MM1028 N_KAPWR_M1028_d N_A_612_71#_M1028_g A_1565_419# VPB PHIGHVT L=0.25 W=1
+ AD=0.145 AS=0.105 PD=1.29 PS=1.21 NRD=1.9503 NRS=9.8303 M=1 R=4 SA=125001
+ SB=125002 A=0.25 P=2.5 MULT=1
MM1009 A_1765_419# N_A_1324_394#_M1009_g N_KAPWR_M1028_d VPB PHIGHVT L=0.25 W=1
+ AD=0.105 AS=0.145 PD=1.21 PS=1.29 NRD=9.8303 NRS=0 M=1 R=4 SA=125001 SB=125001
+ A=0.25 P=2.5 MULT=1
MM1014 N_A_612_71#_M1014_d N_RESET_B_M1014_g A_1765_419# VPB PHIGHVT L=0.25 W=1
+ AD=0.255 AS=0.105 PD=1.51 PS=1.21 NRD=22.6353 NRS=9.8303 M=1 R=4 SA=125002
+ SB=125001 A=0.25 P=2.5 MULT=1
MM1004 N_KAPWR_M1004_d N_A_438_97#_M1004_g N_A_612_71#_M1014_d VPB PHIGHVT
+ L=0.25 W=1 AD=0.285 AS=0.255 PD=2.57 PS=1.51 NRD=0 NRS=22.6353 M=1 R=4
+ SA=125002 SB=125000 A=0.25 P=2.5 MULT=1
MM1034 N_VPWR_M1034_d N_A_438_97#_M1034_g N_A_2120_55#_M1034_s VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.144674 AS=0.1824 PD=1.11495 PS=1.85 NRD=36.1495 NRS=0 M=1
+ R=4.26667 SA=75000.2 SB=75000.8 A=0.096 P=1.58 MULT=1
MM1012 N_Q_M1012_d N_A_2120_55#_M1012_g N_VPWR_M1034_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3591 AS=0.284826 PD=3.09 PS=2.19505 NRD=0 NRS=0 M=1 R=8.4 SA=75000.5
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX36_noxref VNB VPB NWDIODE A=23.6357 P=29
c_120 VNB 0 1.20584e-19 $X=0 $Y=0
*
.include "sky130_fd_sc_lp__srdlrtp_1.pxi.spice"
*
.ends
*
*
