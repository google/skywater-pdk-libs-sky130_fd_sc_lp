* File: sky130_fd_sc_lp__a2111o_1.pxi.spice
* Created: Wed Sep  2 09:16:13 2020
* 
x_PM_SKY130_FD_SC_LP__A2111O_1%A_105_239# N_A_105_239#_M1011_d
+ N_A_105_239#_M1003_d N_A_105_239#_M1009_s N_A_105_239#_M1008_g
+ N_A_105_239#_c_66_n N_A_105_239#_M1010_g N_A_105_239#_c_67_n
+ N_A_105_239#_c_68_n N_A_105_239#_c_69_n N_A_105_239#_c_114_p
+ N_A_105_239#_c_74_n N_A_105_239#_c_119_p N_A_105_239#_c_75_n
+ N_A_105_239#_c_136_p N_A_105_239#_c_70_n N_A_105_239#_c_94_p
+ N_A_105_239#_c_71_n PM_SKY130_FD_SC_LP__A2111O_1%A_105_239#
x_PM_SKY130_FD_SC_LP__A2111O_1%D1 N_D1_M1011_g N_D1_M1009_g D1 D1 N_D1_c_148_n
+ PM_SKY130_FD_SC_LP__A2111O_1%D1
x_PM_SKY130_FD_SC_LP__A2111O_1%C1 N_C1_M1000_g N_C1_M1001_g C1 C1 C1 C1
+ N_C1_c_183_n N_C1_c_184_n PM_SKY130_FD_SC_LP__A2111O_1%C1
x_PM_SKY130_FD_SC_LP__A2111O_1%B1 N_B1_M1003_g N_B1_M1004_g B1 N_B1_c_222_n
+ N_B1_c_223_n PM_SKY130_FD_SC_LP__A2111O_1%B1
x_PM_SKY130_FD_SC_LP__A2111O_1%A1 N_A1_M1007_g N_A1_M1005_g A1 A1 N_A1_c_259_n
+ N_A1_c_260_n PM_SKY130_FD_SC_LP__A2111O_1%A1
x_PM_SKY130_FD_SC_LP__A2111O_1%A2 N_A2_c_294_n N_A2_M1006_g N_A2_M1002_g A2 A2
+ N_A2_c_297_n PM_SKY130_FD_SC_LP__A2111O_1%A2
x_PM_SKY130_FD_SC_LP__A2111O_1%X N_X_M1010_s N_X_M1008_s X X X X X X X
+ N_X_c_319_n N_X_c_321_n PM_SKY130_FD_SC_LP__A2111O_1%X
x_PM_SKY130_FD_SC_LP__A2111O_1%VPWR N_VPWR_M1008_d N_VPWR_M1007_d N_VPWR_c_336_n
+ N_VPWR_c_337_n N_VPWR_c_338_n N_VPWR_c_339_n VPWR N_VPWR_c_340_n
+ N_VPWR_c_335_n N_VPWR_c_342_n PM_SKY130_FD_SC_LP__A2111O_1%VPWR
x_PM_SKY130_FD_SC_LP__A2111O_1%A_511_367# N_A_511_367#_M1004_d
+ N_A_511_367#_M1002_d N_A_511_367#_c_388_n N_A_511_367#_c_389_n
+ N_A_511_367#_c_397_n N_A_511_367#_c_386_n N_A_511_367#_c_387_n
+ PM_SKY130_FD_SC_LP__A2111O_1%A_511_367#
x_PM_SKY130_FD_SC_LP__A2111O_1%VGND N_VGND_M1010_d N_VGND_M1000_d N_VGND_M1006_d
+ N_VGND_c_410_n N_VGND_c_411_n N_VGND_c_412_n N_VGND_c_413_n N_VGND_c_414_n
+ VGND N_VGND_c_415_n N_VGND_c_416_n N_VGND_c_417_n N_VGND_c_418_n
+ PM_SKY130_FD_SC_LP__A2111O_1%VGND
cc_1 VNB N_A_105_239#_M1008_g 0.00838258f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=2.465
cc_2 VNB N_A_105_239#_c_66_n 0.0211217f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.195
cc_3 VNB N_A_105_239#_c_67_n 0.00202682f $X=-0.19 $Y=-0.245 $X2=0.795 $Y2=1.36
cc_4 VNB N_A_105_239#_c_68_n 0.0482582f $X=-0.19 $Y=-0.245 $X2=0.795 $Y2=1.36
cc_5 VNB N_A_105_239#_c_69_n 0.0080457f $X=-0.19 $Y=-0.245 $X2=1.63 $Y2=1.08
cc_6 VNB N_A_105_239#_c_70_n 0.00970604f $X=-0.19 $Y=-0.245 $X2=2.53 $Y2=1.08
cc_7 VNB N_A_105_239#_c_71_n 0.00482346f $X=-0.19 $Y=-0.245 $X2=1.745 $Y2=1.08
cc_8 VNB N_D1_M1011_g 0.0270466f $X=-0.19 $Y=-0.245 $X2=1.21 $Y2=1.835
cc_9 VNB D1 0.00943733f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.525
cc_10 VNB N_D1_c_148_n 0.0253069f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.195
cc_11 VNB N_C1_M1000_g 0.025331f $X=-0.19 $Y=-0.245 $X2=1.21 $Y2=1.835
cc_12 VNB N_C1_c_183_n 0.0246582f $X=-0.19 $Y=-0.245 $X2=0.797 $Y2=1.92
cc_13 VNB N_C1_c_184_n 0.00425744f $X=-0.19 $Y=-0.245 $X2=0.797 $Y2=1.36
cc_14 VNB N_B1_M1003_g 0.0287133f $X=-0.19 $Y=-0.245 $X2=1.21 $Y2=1.835
cc_15 VNB N_B1_c_222_n 0.0287806f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=2.465
cc_16 VNB N_B1_c_223_n 0.00448124f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A1_M1007_g 0.00527299f $X=-0.19 $Y=-0.245 $X2=1.21 $Y2=1.835
cc_18 VNB A1 0.0122521f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.525
cc_19 VNB N_A1_c_259_n 0.0316323f $X=-0.19 $Y=-0.245 $X2=0.797 $Y2=1.165
cc_20 VNB N_A1_c_260_n 0.0195118f $X=-0.19 $Y=-0.245 $X2=0.797 $Y2=1.36
cc_21 VNB N_A2_c_294_n 0.0219493f $X=-0.19 $Y=-0.245 $X2=1.585 $Y2=0.245
cc_22 VNB N_A2_M1002_g 0.00580554f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB A2 0.0271596f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A2_c_297_n 0.0533707f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=0.665
cc_25 VNB X 0.00583199f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.525
cc_26 VNB N_X_c_319_n 0.0684881f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=1.08
cc_27 VNB N_VPWR_c_335_n 0.183584f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_410_n 0.00525703f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.195
cc_29 VNB N_VGND_c_411_n 0.0341491f $X=-0.19 $Y=-0.245 $X2=0.797 $Y2=1.92
cc_30 VNB N_VGND_c_412_n 0.0113717f $X=-0.19 $Y=-0.245 $X2=0.795 $Y2=1.36
cc_31 VNB N_VGND_c_413_n 0.0346846f $X=-0.19 $Y=-0.245 $X2=0.795 $Y2=1.36
cc_32 VNB N_VGND_c_414_n 0.00521013f $X=-0.19 $Y=-0.245 $X2=1.63 $Y2=1.08
cc_33 VNB N_VGND_c_415_n 0.0149753f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=2.005
cc_34 VNB N_VGND_c_416_n 0.237465f $X=-0.19 $Y=-0.245 $X2=2.885 $Y2=0.42
cc_35 VNB N_VGND_c_417_n 0.034368f $X=-0.19 $Y=-0.245 $X2=1.745 $Y2=1.08
cc_36 VNB N_VGND_c_418_n 0.00634414f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VPB N_A_105_239#_M1008_g 0.025711f $X=-0.19 $Y=1.655 $X2=0.6 $Y2=2.465
cc_38 VPB N_A_105_239#_c_67_n 0.00397391f $X=-0.19 $Y=1.655 $X2=0.795 $Y2=1.36
cc_39 VPB N_A_105_239#_c_74_n 0.0139819f $X=-0.19 $Y=1.655 $X2=1.17 $Y2=2.005
cc_40 VPB N_A_105_239#_c_75_n 0.0101473f $X=-0.19 $Y=1.655 $X2=1.335 $Y2=2.095
cc_41 VPB N_D1_M1009_g 0.022669f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_42 VPB D1 0.0108122f $X=-0.19 $Y=1.655 $X2=0.6 $Y2=1.525
cc_43 VPB N_D1_c_148_n 0.00652754f $X=-0.19 $Y=1.655 $X2=0.64 $Y2=1.195
cc_44 VPB N_C1_M1001_g 0.0191011f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_45 VPB N_C1_c_183_n 0.00640484f $X=-0.19 $Y=1.655 $X2=0.797 $Y2=1.92
cc_46 VPB N_C1_c_184_n 0.00143494f $X=-0.19 $Y=1.655 $X2=0.797 $Y2=1.36
cc_47 VPB N_B1_M1004_g 0.0228712f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_48 VPB N_B1_c_222_n 0.00836056f $X=-0.19 $Y=1.655 $X2=0.6 $Y2=2.465
cc_49 VPB N_B1_c_223_n 0.00313968f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_50 VPB N_A1_M1007_g 0.0220182f $X=-0.19 $Y=1.655 $X2=1.21 $Y2=1.835
cc_51 VPB A1 0.00514175f $X=-0.19 $Y=1.655 $X2=0.6 $Y2=1.525
cc_52 VPB N_A2_M1002_g 0.0246361f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_53 VPB A2 0.0138149f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_54 VPB X 0.00882392f $X=-0.19 $Y=1.655 $X2=0.6 $Y2=1.525
cc_55 VPB N_X_c_321_n 0.0599565f $X=-0.19 $Y=1.655 $X2=1.745 $Y2=0.42
cc_56 VPB N_VPWR_c_336_n 0.0107864f $X=-0.19 $Y=1.655 $X2=0.6 $Y2=2.465
cc_57 VPB N_VPWR_c_337_n 4.89148e-19 $X=-0.19 $Y=1.655 $X2=0.64 $Y2=0.665
cc_58 VPB N_VPWR_c_338_n 0.0613615f $X=-0.19 $Y=1.655 $X2=0.797 $Y2=1.92
cc_59 VPB N_VPWR_c_339_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0.797 $Y2=1.36
cc_60 VPB N_VPWR_c_340_n 0.0206265f $X=-0.19 $Y=1.655 $X2=1.335 $Y2=2.91
cc_61 VPB N_VPWR_c_335_n 0.0610852f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_62 VPB N_VPWR_c_342_n 0.023192f $X=-0.19 $Y=1.655 $X2=1.725 $Y2=0.42
cc_63 VPB N_A_511_367#_c_386_n 0.00745115f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_64 VPB N_A_511_367#_c_387_n 0.0369431f $X=-0.19 $Y=1.655 $X2=0.64 $Y2=0.665
cc_65 N_A_105_239#_c_66_n N_D1_M1011_g 0.0049101f $X=0.64 $Y=1.195 $X2=0 $Y2=0
cc_66 N_A_105_239#_c_67_n N_D1_M1011_g 0.00119286f $X=0.795 $Y=1.36 $X2=0 $Y2=0
cc_67 N_A_105_239#_c_68_n N_D1_M1011_g 0.00423349f $X=0.795 $Y=1.36 $X2=0 $Y2=0
cc_68 N_A_105_239#_c_69_n N_D1_M1011_g 0.0146932f $X=1.63 $Y=1.08 $X2=0 $Y2=0
cc_69 N_A_105_239#_c_67_n N_D1_M1009_g 0.00396707f $X=0.795 $Y=1.36 $X2=0 $Y2=0
cc_70 N_A_105_239#_c_74_n N_D1_M1009_g 0.00304054f $X=1.17 $Y=2.005 $X2=0 $Y2=0
cc_71 N_A_105_239#_c_75_n N_D1_M1009_g 0.0166633f $X=1.335 $Y=2.095 $X2=0 $Y2=0
cc_72 N_A_105_239#_c_67_n D1 0.0347947f $X=0.795 $Y=1.36 $X2=0 $Y2=0
cc_73 N_A_105_239#_c_68_n D1 0.00170917f $X=0.795 $Y=1.36 $X2=0 $Y2=0
cc_74 N_A_105_239#_c_69_n D1 0.0435774f $X=1.63 $Y=1.08 $X2=0 $Y2=0
cc_75 N_A_105_239#_c_74_n D1 0.0340237f $X=1.17 $Y=2.005 $X2=0 $Y2=0
cc_76 N_A_105_239#_c_71_n D1 0.0130406f $X=1.745 $Y=1.08 $X2=0 $Y2=0
cc_77 N_A_105_239#_M1008_g N_D1_c_148_n 0.00169675f $X=0.6 $Y=2.465 $X2=0 $Y2=0
cc_78 N_A_105_239#_c_67_n N_D1_c_148_n 5.18034e-19 $X=0.795 $Y=1.36 $X2=0 $Y2=0
cc_79 N_A_105_239#_c_68_n N_D1_c_148_n 0.00611744f $X=0.795 $Y=1.36 $X2=0 $Y2=0
cc_80 N_A_105_239#_c_69_n N_D1_c_148_n 0.0012307f $X=1.63 $Y=1.08 $X2=0 $Y2=0
cc_81 N_A_105_239#_c_74_n N_D1_c_148_n 0.0010224f $X=1.17 $Y=2.005 $X2=0 $Y2=0
cc_82 N_A_105_239#_c_70_n N_C1_M1000_g 0.0169156f $X=2.53 $Y=1.08 $X2=0 $Y2=0
cc_83 N_A_105_239#_c_94_p N_C1_M1000_g 3.84467e-19 $X=3.075 $Y=0.42 $X2=0 $Y2=0
cc_84 N_A_105_239#_c_74_n N_C1_M1001_g 4.68513e-19 $X=1.17 $Y=2.005 $X2=0 $Y2=0
cc_85 N_A_105_239#_c_75_n N_C1_M1001_g 0.00297603f $X=1.335 $Y=2.095 $X2=0 $Y2=0
cc_86 N_A_105_239#_c_70_n N_C1_c_183_n 0.00123224f $X=2.53 $Y=1.08 $X2=0 $Y2=0
cc_87 N_A_105_239#_c_74_n N_C1_c_184_n 0.00619288f $X=1.17 $Y=2.005 $X2=0 $Y2=0
cc_88 N_A_105_239#_c_75_n N_C1_c_184_n 0.0298582f $X=1.335 $Y=2.095 $X2=0 $Y2=0
cc_89 N_A_105_239#_c_70_n N_C1_c_184_n 0.026284f $X=2.53 $Y=1.08 $X2=0 $Y2=0
cc_90 N_A_105_239#_c_70_n N_B1_M1003_g 0.0146248f $X=2.53 $Y=1.08 $X2=0 $Y2=0
cc_91 N_A_105_239#_c_94_p N_B1_M1003_g 0.0120962f $X=3.075 $Y=0.42 $X2=0 $Y2=0
cc_92 N_A_105_239#_c_70_n N_B1_c_222_n 0.00184634f $X=2.53 $Y=1.08 $X2=0 $Y2=0
cc_93 N_A_105_239#_c_70_n N_B1_c_223_n 0.0327261f $X=2.53 $Y=1.08 $X2=0 $Y2=0
cc_94 N_A_105_239#_c_70_n A1 0.0188077f $X=2.53 $Y=1.08 $X2=0 $Y2=0
cc_95 N_A_105_239#_c_70_n N_A1_c_259_n 0.00487617f $X=2.53 $Y=1.08 $X2=0 $Y2=0
cc_96 N_A_105_239#_c_70_n N_A1_c_260_n 0.00381905f $X=2.53 $Y=1.08 $X2=0 $Y2=0
cc_97 N_A_105_239#_c_94_p N_A1_c_260_n 0.0145895f $X=3.075 $Y=0.42 $X2=0 $Y2=0
cc_98 N_A_105_239#_c_94_p N_A2_c_294_n 0.00200143f $X=3.075 $Y=0.42 $X2=-0.19
+ $Y2=-0.245
cc_99 N_A_105_239#_M1008_g X 0.0078902f $X=0.6 $Y=2.465 $X2=0 $Y2=0
cc_100 N_A_105_239#_c_66_n N_X_c_319_n 0.00501121f $X=0.64 $Y=1.195 $X2=0 $Y2=0
cc_101 N_A_105_239#_c_67_n N_X_c_319_n 0.0487435f $X=0.795 $Y=1.36 $X2=0 $Y2=0
cc_102 N_A_105_239#_c_68_n N_X_c_319_n 0.0078902f $X=0.795 $Y=1.36 $X2=0 $Y2=0
cc_103 N_A_105_239#_c_114_p N_X_c_319_n 0.0106024f $X=0.905 $Y=1.08 $X2=0 $Y2=0
cc_104 N_A_105_239#_M1008_g N_X_c_321_n 0.00430917f $X=0.6 $Y=2.465 $X2=0 $Y2=0
cc_105 N_A_105_239#_c_67_n N_X_c_321_n 0.00412028f $X=0.795 $Y=1.36 $X2=0 $Y2=0
cc_106 N_A_105_239#_c_67_n N_VPWR_M1008_d 0.00221326f $X=0.795 $Y=1.36 $X2=-0.19
+ $Y2=-0.245
cc_107 N_A_105_239#_c_74_n N_VPWR_M1008_d 0.00115411f $X=1.17 $Y=2.005 $X2=-0.19
+ $Y2=-0.245
cc_108 N_A_105_239#_c_119_p N_VPWR_M1008_d 0.00346372f $X=0.905 $Y=2.005
+ $X2=-0.19 $Y2=-0.245
cc_109 N_A_105_239#_M1008_g N_VPWR_c_336_n 0.0203207f $X=0.6 $Y=2.465 $X2=0
+ $Y2=0
cc_110 N_A_105_239#_c_74_n N_VPWR_c_336_n 0.00610503f $X=1.17 $Y=2.005 $X2=0
+ $Y2=0
cc_111 N_A_105_239#_c_119_p N_VPWR_c_336_n 0.0155529f $X=0.905 $Y=2.005 $X2=0
+ $Y2=0
cc_112 N_A_105_239#_c_75_n N_VPWR_c_336_n 0.0627569f $X=1.335 $Y=2.095 $X2=0
+ $Y2=0
cc_113 N_A_105_239#_c_75_n N_VPWR_c_338_n 0.0210467f $X=1.335 $Y=2.095 $X2=0
+ $Y2=0
cc_114 N_A_105_239#_M1009_s N_VPWR_c_335_n 0.00215158f $X=1.21 $Y=1.835 $X2=0
+ $Y2=0
cc_115 N_A_105_239#_M1008_g N_VPWR_c_335_n 0.00927852f $X=0.6 $Y=2.465 $X2=0
+ $Y2=0
cc_116 N_A_105_239#_c_75_n N_VPWR_c_335_n 0.0125689f $X=1.335 $Y=2.095 $X2=0
+ $Y2=0
cc_117 N_A_105_239#_M1008_g N_VPWR_c_342_n 0.00486043f $X=0.6 $Y=2.465 $X2=0
+ $Y2=0
cc_118 N_A_105_239#_c_69_n N_VGND_M1010_d 0.00604702f $X=1.63 $Y=1.08 $X2=-0.19
+ $Y2=-0.245
cc_119 N_A_105_239#_c_114_p N_VGND_M1010_d 0.00147181f $X=0.905 $Y=1.08
+ $X2=-0.19 $Y2=-0.245
cc_120 N_A_105_239#_c_70_n N_VGND_M1000_d 0.00308172f $X=2.53 $Y=1.08 $X2=0
+ $Y2=0
cc_121 N_A_105_239#_c_70_n N_VGND_c_410_n 0.022455f $X=2.53 $Y=1.08 $X2=0 $Y2=0
cc_122 N_A_105_239#_c_70_n N_VGND_c_411_n 0.00159689f $X=2.53 $Y=1.08 $X2=0
+ $Y2=0
cc_123 N_A_105_239#_c_94_p N_VGND_c_411_n 0.0262773f $X=3.075 $Y=0.42 $X2=0
+ $Y2=0
cc_124 N_A_105_239#_c_94_p N_VGND_c_413_n 0.0456424f $X=3.075 $Y=0.42 $X2=0
+ $Y2=0
cc_125 N_A_105_239#_c_136_p N_VGND_c_415_n 0.0138717f $X=1.725 $Y=0.42 $X2=0
+ $Y2=0
cc_126 N_A_105_239#_M1011_d N_VGND_c_416_n 0.00397496f $X=1.585 $Y=0.245 $X2=0
+ $Y2=0
cc_127 N_A_105_239#_M1003_d N_VGND_c_416_n 0.00529143f $X=2.555 $Y=0.245 $X2=0
+ $Y2=0
cc_128 N_A_105_239#_c_66_n N_VGND_c_416_n 0.00931388f $X=0.64 $Y=1.195 $X2=0
+ $Y2=0
cc_129 N_A_105_239#_c_136_p N_VGND_c_416_n 0.00886411f $X=1.725 $Y=0.42 $X2=0
+ $Y2=0
cc_130 N_A_105_239#_c_94_p N_VGND_c_416_n 0.0271594f $X=3.075 $Y=0.42 $X2=0
+ $Y2=0
cc_131 N_A_105_239#_c_66_n N_VGND_c_417_n 0.0176064f $X=0.64 $Y=1.195 $X2=0
+ $Y2=0
cc_132 N_A_105_239#_c_68_n N_VGND_c_417_n 9.58071e-19 $X=0.795 $Y=1.36 $X2=0
+ $Y2=0
cc_133 N_A_105_239#_c_69_n N_VGND_c_417_n 0.0402322f $X=1.63 $Y=1.08 $X2=0 $Y2=0
cc_134 N_A_105_239#_c_114_p N_VGND_c_417_n 0.0139808f $X=0.905 $Y=1.08 $X2=0
+ $Y2=0
cc_135 N_D1_M1011_g N_C1_M1000_g 0.0236875f $X=1.51 $Y=0.665 $X2=0 $Y2=0
cc_136 D1 N_C1_M1000_g 0.00310374f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_137 N_D1_M1009_g N_C1_M1001_g 0.0474166f $X=1.55 $Y=2.465 $X2=0 $Y2=0
cc_138 N_D1_c_148_n N_C1_c_183_n 0.0474166f $X=1.46 $Y=1.51 $X2=0 $Y2=0
cc_139 N_D1_M1009_g N_C1_c_184_n 0.00409234f $X=1.55 $Y=2.465 $X2=0 $Y2=0
cc_140 D1 N_C1_c_184_n 0.0347616f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_141 N_D1_c_148_n N_C1_c_184_n 3.43721e-19 $X=1.46 $Y=1.51 $X2=0 $Y2=0
cc_142 N_D1_M1009_g N_VPWR_c_336_n 0.0036497f $X=1.55 $Y=2.465 $X2=0 $Y2=0
cc_143 N_D1_M1009_g N_VPWR_c_338_n 0.0054895f $X=1.55 $Y=2.465 $X2=0 $Y2=0
cc_144 N_D1_M1009_g N_VPWR_c_335_n 0.0112391f $X=1.55 $Y=2.465 $X2=0 $Y2=0
cc_145 N_D1_M1011_g N_VGND_c_415_n 0.00479301f $X=1.51 $Y=0.665 $X2=0 $Y2=0
cc_146 N_D1_M1011_g N_VGND_c_416_n 0.00828353f $X=1.51 $Y=0.665 $X2=0 $Y2=0
cc_147 N_D1_M1011_g N_VGND_c_417_n 0.0111902f $X=1.51 $Y=0.665 $X2=0 $Y2=0
cc_148 N_C1_M1000_g N_B1_M1003_g 0.0253716f $X=1.94 $Y=0.665 $X2=0 $Y2=0
cc_149 N_C1_c_184_n N_B1_M1003_g 0.0162326f $X=2.03 $Y=1.51 $X2=0 $Y2=0
cc_150 N_C1_M1001_g N_B1_M1004_g 0.0414535f $X=1.94 $Y=2.465 $X2=0 $Y2=0
cc_151 N_C1_c_183_n N_B1_c_222_n 0.0207938f $X=2.03 $Y=1.51 $X2=0 $Y2=0
cc_152 N_C1_c_183_n N_B1_c_223_n 3.40353e-19 $X=2.03 $Y=1.51 $X2=0 $Y2=0
cc_153 N_C1_c_184_n N_B1_c_223_n 0.0330561f $X=2.03 $Y=1.51 $X2=0 $Y2=0
cc_154 N_C1_M1001_g N_VPWR_c_338_n 0.00491168f $X=1.94 $Y=2.465 $X2=0 $Y2=0
cc_155 N_C1_c_184_n N_VPWR_c_338_n 0.0115705f $X=2.03 $Y=1.51 $X2=0 $Y2=0
cc_156 N_C1_M1001_g N_VPWR_c_335_n 0.00866672f $X=1.94 $Y=2.465 $X2=0 $Y2=0
cc_157 N_C1_c_184_n N_VPWR_c_335_n 0.0112666f $X=2.03 $Y=1.51 $X2=0 $Y2=0
cc_158 N_C1_c_184_n A_403_367# 0.0181179f $X=2.03 $Y=1.51 $X2=-0.19 $Y2=-0.245
cc_159 N_C1_c_184_n N_A_511_367#_c_388_n 0.00992069f $X=2.03 $Y=1.51 $X2=0 $Y2=0
cc_160 N_C1_M1001_g N_A_511_367#_c_389_n 0.00120141f $X=1.94 $Y=2.465 $X2=0
+ $Y2=0
cc_161 N_C1_c_184_n N_A_511_367#_c_389_n 0.0495232f $X=2.03 $Y=1.51 $X2=0 $Y2=0
cc_162 N_C1_M1000_g N_VGND_c_410_n 0.00173463f $X=1.94 $Y=0.665 $X2=0 $Y2=0
cc_163 N_C1_M1000_g N_VGND_c_415_n 0.00575161f $X=1.94 $Y=0.665 $X2=0 $Y2=0
cc_164 N_C1_M1000_g N_VGND_c_416_n 0.0108419f $X=1.94 $Y=0.665 $X2=0 $Y2=0
cc_165 N_C1_M1000_g N_VGND_c_417_n 6.23669e-19 $X=1.94 $Y=0.665 $X2=0 $Y2=0
cc_166 N_B1_M1004_g N_A1_M1007_g 0.006591f $X=2.48 $Y=2.465 $X2=0 $Y2=0
cc_167 N_B1_c_222_n N_A1_M1007_g 0.00403328f $X=2.6 $Y=1.51 $X2=0 $Y2=0
cc_168 N_B1_c_223_n N_A1_M1007_g 5.58179e-19 $X=2.6 $Y=1.51 $X2=0 $Y2=0
cc_169 N_B1_M1003_g A1 0.00267026f $X=2.48 $Y=0.665 $X2=0 $Y2=0
cc_170 N_B1_M1004_g A1 4.0152e-19 $X=2.48 $Y=2.465 $X2=0 $Y2=0
cc_171 N_B1_c_222_n A1 0.00123581f $X=2.6 $Y=1.51 $X2=0 $Y2=0
cc_172 N_B1_c_223_n A1 0.0372162f $X=2.6 $Y=1.51 $X2=0 $Y2=0
cc_173 N_B1_M1003_g N_A1_c_259_n 0.00300418f $X=2.48 $Y=0.665 $X2=0 $Y2=0
cc_174 N_B1_c_222_n N_A1_c_259_n 0.0126694f $X=2.6 $Y=1.51 $X2=0 $Y2=0
cc_175 N_B1_c_223_n N_A1_c_259_n 6.72924e-19 $X=2.6 $Y=1.51 $X2=0 $Y2=0
cc_176 N_B1_M1003_g N_A1_c_260_n 0.0054909f $X=2.48 $Y=0.665 $X2=0 $Y2=0
cc_177 N_B1_M1004_g N_VPWR_c_338_n 0.0054895f $X=2.48 $Y=2.465 $X2=0 $Y2=0
cc_178 N_B1_M1004_g N_VPWR_c_335_n 0.0109499f $X=2.48 $Y=2.465 $X2=0 $Y2=0
cc_179 N_B1_M1004_g N_A_511_367#_c_388_n 0.002494f $X=2.48 $Y=2.465 $X2=0 $Y2=0
cc_180 N_B1_c_222_n N_A_511_367#_c_388_n 0.00140711f $X=2.6 $Y=1.51 $X2=0 $Y2=0
cc_181 N_B1_c_223_n N_A_511_367#_c_388_n 0.0218695f $X=2.6 $Y=1.51 $X2=0 $Y2=0
cc_182 N_B1_M1004_g N_A_511_367#_c_389_n 0.0155982f $X=2.48 $Y=2.465 $X2=0 $Y2=0
cc_183 N_B1_M1003_g N_VGND_c_410_n 0.00634658f $X=2.48 $Y=0.665 $X2=0 $Y2=0
cc_184 N_B1_M1003_g N_VGND_c_413_n 0.00539298f $X=2.48 $Y=0.665 $X2=0 $Y2=0
cc_185 N_B1_M1003_g N_VGND_c_416_n 0.0107839f $X=2.48 $Y=0.665 $X2=0 $Y2=0
cc_186 N_A1_c_260_n N_A2_c_294_n 0.0433441f $X=3.185 $Y=1.21 $X2=-0.19
+ $Y2=-0.245
cc_187 N_A1_M1007_g N_A2_M1002_g 0.0445854f $X=3.25 $Y=2.465 $X2=0 $Y2=0
cc_188 A1 N_A2_M1002_g 0.0071336f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_189 A1 A2 0.045102f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_190 A1 N_A2_c_297_n 0.0181405f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_191 N_A1_c_259_n N_A2_c_297_n 0.0433441f $X=3.2 $Y=1.375 $X2=0 $Y2=0
cc_192 N_A1_M1007_g N_VPWR_c_337_n 0.0167102f $X=3.25 $Y=2.465 $X2=0 $Y2=0
cc_193 N_A1_M1007_g N_VPWR_c_338_n 0.00486043f $X=3.25 $Y=2.465 $X2=0 $Y2=0
cc_194 N_A1_M1007_g N_VPWR_c_335_n 0.00888845f $X=3.25 $Y=2.465 $X2=0 $Y2=0
cc_195 A1 N_A_511_367#_c_388_n 0.0120677f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_196 N_A1_c_259_n N_A_511_367#_c_388_n 5.77357e-19 $X=3.2 $Y=1.375 $X2=0 $Y2=0
cc_197 N_A1_M1007_g N_A_511_367#_c_397_n 0.0122129f $X=3.25 $Y=2.465 $X2=0 $Y2=0
cc_198 A1 N_A_511_367#_c_397_n 0.0384822f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_199 N_A1_c_260_n N_VGND_c_411_n 0.003284f $X=3.185 $Y=1.21 $X2=0 $Y2=0
cc_200 N_A1_c_260_n N_VGND_c_413_n 0.00539298f $X=3.185 $Y=1.21 $X2=0 $Y2=0
cc_201 N_A1_c_260_n N_VGND_c_416_n 0.0105081f $X=3.185 $Y=1.21 $X2=0 $Y2=0
cc_202 N_A2_M1002_g N_VPWR_c_337_n 0.0167102f $X=3.68 $Y=2.465 $X2=0 $Y2=0
cc_203 N_A2_M1002_g N_VPWR_c_340_n 0.00486043f $X=3.68 $Y=2.465 $X2=0 $Y2=0
cc_204 N_A2_M1002_g N_VPWR_c_335_n 0.00930295f $X=3.68 $Y=2.465 $X2=0 $Y2=0
cc_205 N_A2_M1002_g N_A_511_367#_c_397_n 0.0140148f $X=3.68 $Y=2.465 $X2=0 $Y2=0
cc_206 A2 N_A_511_367#_c_386_n 0.0176196f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_207 N_A2_c_297_n N_A_511_367#_c_386_n 0.00302448f $X=3.95 $Y=1.375 $X2=0
+ $Y2=0
cc_208 N_A2_c_294_n N_VGND_c_411_n 0.0229543f $X=3.65 $Y=1.21 $X2=0 $Y2=0
cc_209 A2 N_VGND_c_411_n 0.014096f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_210 N_A2_c_297_n N_VGND_c_411_n 0.00629566f $X=3.95 $Y=1.375 $X2=0 $Y2=0
cc_211 N_A2_c_294_n N_VGND_c_413_n 0.00477554f $X=3.65 $Y=1.21 $X2=0 $Y2=0
cc_212 N_A2_c_294_n N_VGND_c_416_n 0.00814835f $X=3.65 $Y=1.21 $X2=0 $Y2=0
cc_213 N_X_M1008_s N_VPWR_c_335_n 0.00371702f $X=0.26 $Y=1.835 $X2=0 $Y2=0
cc_214 N_X_c_321_n N_VPWR_c_335_n 0.0152789f $X=0.385 $Y=1.98 $X2=0 $Y2=0
cc_215 N_X_c_321_n N_VPWR_c_342_n 0.0274888f $X=0.385 $Y=1.98 $X2=0 $Y2=0
cc_216 N_X_M1010_s N_VGND_c_416_n 0.00368844f $X=0.3 $Y=0.245 $X2=0 $Y2=0
cc_217 N_X_c_319_n N_VGND_c_416_n 0.016834f $X=0.425 $Y=0.42 $X2=0 $Y2=0
cc_218 N_X_c_319_n N_VGND_c_417_n 0.0303563f $X=0.425 $Y=0.42 $X2=0 $Y2=0
cc_219 N_VPWR_c_335_n A_325_367# 0.010279f $X=4.08 $Y=3.33 $X2=-0.19 $Y2=-0.245
cc_220 N_VPWR_c_335_n A_403_367# 0.00816765f $X=4.08 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_221 N_VPWR_c_335_n N_A_511_367#_M1004_d 0.00662261f $X=4.08 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_222 N_VPWR_c_335_n N_A_511_367#_M1002_d 0.00371702f $X=4.08 $Y=3.33 $X2=0
+ $Y2=0
cc_223 N_VPWR_c_338_n N_A_511_367#_c_389_n 0.0395943f $X=3.3 $Y=3.33 $X2=0 $Y2=0
cc_224 N_VPWR_c_335_n N_A_511_367#_c_389_n 0.0230659f $X=4.08 $Y=3.33 $X2=0
+ $Y2=0
cc_225 N_VPWR_M1007_d N_A_511_367#_c_397_n 0.00353353f $X=3.325 $Y=1.835 $X2=0
+ $Y2=0
cc_226 N_VPWR_c_337_n N_A_511_367#_c_397_n 0.0170777f $X=3.465 $Y=2.375 $X2=0
+ $Y2=0
cc_227 N_VPWR_c_340_n N_A_511_367#_c_387_n 0.0178111f $X=4.08 $Y=3.33 $X2=0
+ $Y2=0
cc_228 N_VPWR_c_335_n N_A_511_367#_c_387_n 0.0100304f $X=4.08 $Y=3.33 $X2=0
+ $Y2=0
cc_229 N_VGND_c_416_n A_673_49# 0.00899413f $X=4.08 $Y=0 $X2=-0.19 $Y2=-0.245
