* File: sky130_fd_sc_lp__a2bb2oi_1.pex.spice
* Created: Fri Aug 28 09:56:38 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A2BB2OI_1%A1_N 3 6 8 10 17 19
r26 17 20 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.4 $Y=1.375
+ $X2=0.4 $Y2=1.54
r27 17 19 50.583 $w=3.3e-07 $l=1.9e-07 $layer=POLY_cond $X=0.4 $Y=1.375 $X2=0.4
+ $Y2=1.185
r28 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.4
+ $Y=1.375 $X2=0.4 $Y2=1.375
r29 10 18 7.08787 $w=5.38e-07 $l=3.2e-07 $layer=LI1_cond $X=0.72 $Y=1.48 $X2=0.4
+ $Y2=1.48
r30 8 18 3.54394 $w=5.38e-07 $l=1.6e-07 $layer=LI1_cond $X=0.24 $Y=1.48 $X2=0.4
+ $Y2=1.48
r31 6 20 474.309 $w=1.5e-07 $l=9.25e-07 $layer=POLY_cond $X=0.49 $Y=2.465
+ $X2=0.49 $Y2=1.54
r32 3 19 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.49 $Y=0.655
+ $X2=0.49 $Y2=1.185
.ends

.subckt PM_SKY130_FD_SC_LP__A2BB2OI_1%A2_N 1 3 4 6 7
r33 7 10 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.16
+ $Y=1.35 $X2=1.16 $Y2=1.35
r34 4 10 40.6804 $w=4.5e-07 $l=2.26164e-07 $layer=POLY_cond $X=0.92 $Y=1.185
+ $X2=1.065 $Y2=1.35
r35 4 6 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.92 $Y=1.185 $X2=0.92
+ $Y2=0.655
r36 1 10 63.1737 $w=4.5e-07 $l=4.58258e-07 $layer=POLY_cond $X=0.88 $Y=1.725
+ $X2=1.065 $Y2=1.35
r37 1 3 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=0.88 $Y=1.725 $X2=0.88
+ $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__A2BB2OI_1%A_113_47# 1 2 9 12 16 18 19 20 22 24 29 34
+ 35 36 39
c68 36 0 6.54081e-20 $X=1.725 $Y=1.2
c69 34 0 9.66306e-21 $X=1.73 $Y=1.35
r70 35 40 46.3065 $w=3.4e-07 $l=1.65e-07 $layer=POLY_cond $X=1.735 $Y=1.35
+ $X2=1.735 $Y2=1.515
r71 35 39 46.3065 $w=3.4e-07 $l=1.65e-07 $layer=POLY_cond $X=1.735 $Y=1.35
+ $X2=1.735 $Y2=1.185
r72 34 37 8.13106 $w=3.38e-07 $l=1.65e-07 $layer=LI1_cond $X=1.725 $Y=1.35
+ $X2=1.725 $Y2=1.515
r73 34 36 7.62263 $w=3.38e-07 $l=1.5e-07 $layer=LI1_cond $X=1.725 $Y=1.35
+ $X2=1.725 $Y2=1.2
r74 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.73
+ $Y=1.35 $X2=1.73 $Y2=1.35
r75 30 32 8.02632 $w=3.04e-07 $l=2e-07 $layer=LI1_cond $X=1.095 $Y=1.78
+ $X2=1.095 $Y2=1.98
r76 29 37 11.0909 $w=1.78e-07 $l=1.8e-07 $layer=LI1_cond $X=1.645 $Y=1.695
+ $X2=1.645 $Y2=1.515
r77 26 36 11.399 $w=1.78e-07 $l=1.85e-07 $layer=LI1_cond $X=1.645 $Y=1.015
+ $X2=1.645 $Y2=1.2
r78 25 30 4.13891 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.26 $Y=1.78
+ $X2=1.095 $Y2=1.78
r79 24 29 6.82373 $w=1.7e-07 $l=1.25499e-07 $layer=LI1_cond $X=1.555 $Y=1.78
+ $X2=1.645 $Y2=1.695
r80 24 25 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.555 $Y=1.78
+ $X2=1.26 $Y2=1.78
r81 20 32 3.97847 $w=3.3e-07 $l=1.05e-07 $layer=LI1_cond $X=1.095 $Y=2.085
+ $X2=1.095 $Y2=1.98
r82 20 22 30.208 $w=3.28e-07 $l=8.65e-07 $layer=LI1_cond $X=1.095 $Y=2.085
+ $X2=1.095 $Y2=2.95
r83 18 26 6.82373 $w=1.7e-07 $l=1.25499e-07 $layer=LI1_cond $X=1.555 $Y=0.93
+ $X2=1.645 $Y2=1.015
r84 18 19 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=1.555 $Y=0.93
+ $X2=0.8 $Y2=0.93
r85 14 19 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=0.705 $Y=0.845
+ $X2=0.8 $Y2=0.93
r86 14 16 24.8086 $w=1.88e-07 $l=4.25e-07 $layer=LI1_cond $X=0.705 $Y=0.845
+ $X2=0.705 $Y2=0.42
r87 12 40 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=1.83 $Y=2.465
+ $X2=1.83 $Y2=1.515
r88 9 39 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.83 $Y=0.655
+ $X2=1.83 $Y2=1.185
r89 2 32 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.955
+ $Y=1.835 $X2=1.095 $Y2=1.98
r90 2 22 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=0.955
+ $Y=1.835 $X2=1.095 $Y2=2.95
r91 1 16 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=0.565
+ $Y=0.235 $X2=0.705 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__A2BB2OI_1%B2 3 7 9 10 14
c41 9 0 2.66849e-20 $X=2.16 $Y=1.295
c42 3 0 7.50712e-20 $X=2.26 $Y=0.655
r43 14 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.31 $Y=1.375
+ $X2=2.31 $Y2=1.54
r44 14 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.31 $Y=1.375
+ $X2=2.31 $Y2=1.21
r45 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.31
+ $Y=1.375 $X2=2.31 $Y2=1.375
r46 10 15 9.82966 $w=3.38e-07 $l=2.9e-07 $layer=LI1_cond $X=2.235 $Y=1.665
+ $X2=2.235 $Y2=1.375
r47 9 15 2.71163 $w=3.38e-07 $l=8e-08 $layer=LI1_cond $X=2.235 $Y=1.295
+ $X2=2.235 $Y2=1.375
r48 7 17 474.309 $w=1.5e-07 $l=9.25e-07 $layer=POLY_cond $X=2.265 $Y=2.465
+ $X2=2.265 $Y2=1.54
r49 3 16 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=2.26 $Y=0.655
+ $X2=2.26 $Y2=1.21
.ends

.subckt PM_SKY130_FD_SC_LP__A2BB2OI_1%B1 3 7 9 10 17
c30 3 0 2.66849e-20 $X=2.79 $Y=0.655
r31 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.01
+ $Y=1.375 $X2=3.01 $Y2=1.375
r32 15 17 34.0979 $w=3.3e-07 $l=1.95e-07 $layer=POLY_cond $X=2.815 $Y=1.375
+ $X2=3.01 $Y2=1.375
r33 13 15 4.37153 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=2.79 $Y=1.375
+ $X2=2.815 $Y2=1.375
r34 10 18 9.28357 $w=3.58e-07 $l=2.9e-07 $layer=LI1_cond $X=3.095 $Y=1.665
+ $X2=3.095 $Y2=1.375
r35 9 18 2.56098 $w=3.58e-07 $l=8e-08 $layer=LI1_cond $X=3.095 $Y=1.295
+ $X2=3.095 $Y2=1.375
r36 5 15 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.815 $Y=1.54
+ $X2=2.815 $Y2=1.375
r37 5 7 474.309 $w=1.5e-07 $l=9.25e-07 $layer=POLY_cond $X=2.815 $Y=1.54
+ $X2=2.815 $Y2=2.465
r38 1 13 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.79 $Y=1.21
+ $X2=2.79 $Y2=1.375
r39 1 3 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=2.79 $Y=1.21 $X2=2.79
+ $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__A2BB2OI_1%VPWR 1 2 7 9 15 18 19 20 30 31
r44 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r45 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r46 28 31 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r47 27 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r48 25 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r49 24 27 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=0.72 $Y=3.33
+ $X2=2.16 $Y2=3.33
r50 24 25 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r51 22 34 4.746 $w=1.7e-07 $l=2.2e-07 $layer=LI1_cond $X=0.44 $Y=3.33 $X2=0.22
+ $Y2=3.33
r52 22 24 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=0.44 $Y=3.33
+ $X2=0.72 $Y2=3.33
r53 20 28 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r54 20 25 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.72 $Y2=3.33
r55 18 27 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=2.38 $Y=3.33
+ $X2=2.16 $Y2=3.33
r56 18 19 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.38 $Y=3.33
+ $X2=2.545 $Y2=3.33
r57 17 30 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=2.71 $Y=3.33
+ $X2=3.12 $Y2=3.33
r58 17 19 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.71 $Y=3.33
+ $X2=2.545 $Y2=3.33
r59 13 19 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.545 $Y=3.245
+ $X2=2.545 $Y2=3.33
r60 13 15 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=2.545 $Y=3.245
+ $X2=2.545 $Y2=2.83
r61 9 12 33.0018 $w=3.28e-07 $l=9.45e-07 $layer=LI1_cond $X=0.275 $Y=2.005
+ $X2=0.275 $Y2=2.95
r62 7 34 3.02018 $w=3.3e-07 $l=1.09087e-07 $layer=LI1_cond $X=0.275 $Y=3.245
+ $X2=0.22 $Y2=3.33
r63 7 12 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.275 $Y=3.245
+ $X2=0.275 $Y2=2.95
r64 2 15 600 $w=1.7e-07 $l=1.0927e-06 $layer=licon1_PDIFF $count=1 $X=2.34
+ $Y=1.835 $X2=2.545 $Y2=2.83
r65 1 12 400 $w=1.7e-07 $l=1.17584e-06 $layer=licon1_PDIFF $count=1 $X=0.15
+ $Y=1.835 $X2=0.275 $Y2=2.95
r66 1 9 400 $w=1.7e-07 $l=2.23942e-07 $layer=licon1_PDIFF $count=1 $X=0.15
+ $Y=1.835 $X2=0.275 $Y2=2.005
.ends

.subckt PM_SKY130_FD_SC_LP__A2BB2OI_1%Y 1 2 7 11 13 14 16 17 20 21
r51 21 29 4.78707 $w=3.23e-07 $l=1.35e-07 $layer=LI1_cond $X=1.612 $Y=2.775
+ $X2=1.612 $Y2=2.91
r52 20 21 13.1201 $w=3.23e-07 $l=3.7e-07 $layer=LI1_cond $X=1.612 $Y=2.405
+ $X2=1.612 $Y2=2.775
r53 17 20 7.09196 $w=3.23e-07 $l=2e-07 $layer=LI1_cond $X=1.612 $Y=2.205
+ $X2=1.612 $Y2=2.405
r54 17 19 2.64734 $w=3.25e-07 $l=8.5e-08 $layer=LI1_cond $X=1.612 $Y=2.205
+ $X2=1.612 $Y2=2.12
r55 15 16 65.5668 $w=1.68e-07 $l=1.005e-06 $layer=LI1_cond $X=2.66 $Y=1.03
+ $X2=2.66 $Y2=2.035
r56 13 15 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.575 $Y=0.945
+ $X2=2.66 $Y2=1.03
r57 13 14 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=2.575 $Y=0.945
+ $X2=2.15 $Y2=0.945
r58 9 14 6.87494 $w=1.7e-07 $l=1.36015e-07 $layer=LI1_cond $X=2.05 $Y=0.86
+ $X2=2.15 $Y2=0.945
r59 9 11 24.4 $w=1.98e-07 $l=4.4e-07 $layer=LI1_cond $X=2.05 $Y=0.86 $X2=2.05
+ $Y2=0.42
r60 8 19 5.07667 $w=1.7e-07 $l=1.63e-07 $layer=LI1_cond $X=1.775 $Y=2.12
+ $X2=1.612 $Y2=2.12
r61 7 16 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.575 $Y=2.12
+ $X2=2.66 $Y2=2.035
r62 7 8 52.1925 $w=1.68e-07 $l=8e-07 $layer=LI1_cond $X=2.575 $Y=2.12 $X2=1.775
+ $Y2=2.12
r63 2 29 400 $w=1.7e-07 $l=1.13578e-06 $layer=licon1_PDIFF $count=1 $X=1.49
+ $Y=1.835 $X2=1.615 $Y2=2.91
r64 2 19 400 $w=1.7e-07 $l=3.41833e-07 $layer=licon1_PDIFF $count=1 $X=1.49
+ $Y=1.835 $X2=1.615 $Y2=2.12
r65 1 11 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=1.905
+ $Y=0.235 $X2=2.045 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__A2BB2OI_1%A_381_367# 1 2 9 11 12 17 20
r23 15 20 3.17288 $w=2.97e-07 $l=9.35682e-08 $layer=LI1_cond $X=3.055 $Y=2.375
+ $X2=3.037 $Y2=2.46
r24 15 17 11.5244 $w=2.78e-07 $l=2.8e-07 $layer=LI1_cond $X=3.055 $Y=2.375
+ $X2=3.055 $Y2=2.095
r25 11 20 3.41642 $w=1.7e-07 $l=1.57e-07 $layer=LI1_cond $X=2.88 $Y=2.46
+ $X2=3.037 $Y2=2.46
r26 11 12 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.88 $Y=2.46
+ $X2=2.21 $Y2=2.46
r27 7 12 7.24806 $w=1.7e-07 $l=1.70276e-07 $layer=LI1_cond $X=2.077 $Y=2.545
+ $X2=2.21 $Y2=2.46
r28 7 9 0.217442 $w=2.63e-07 $l=5e-09 $layer=LI1_cond $X=2.077 $Y=2.545
+ $X2=2.077 $Y2=2.55
r29 2 20 300 $w=1.7e-07 $l=7.31659e-07 $layer=licon1_PDIFF $count=2 $X=2.89
+ $Y=1.835 $X2=3.03 $Y2=2.5
r30 2 17 600 $w=1.7e-07 $l=3.2249e-07 $layer=licon1_PDIFF $count=1 $X=2.89
+ $Y=1.835 $X2=3.03 $Y2=2.095
r31 1 9 300 $w=1.7e-07 $l=7.84156e-07 $layer=licon1_PDIFF $count=2 $X=1.905
+ $Y=1.835 $X2=2.05 $Y2=2.55
.ends

.subckt PM_SKY130_FD_SC_LP__A2BB2OI_1%VGND 1 2 3 10 12 14 16 18 25 36 42 45
r45 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r46 40 42 10.1628 $w=7.58e-07 $l=1e-07 $layer=LI1_cond $X=1.68 $Y=0.295 $X2=1.78
+ $Y2=0.295
r47 38 40 1.02296 $w=7.58e-07 $l=6.5e-08 $layer=LI1_cond $X=1.615 $Y=0.295
+ $X2=1.68 $Y2=0.295
r48 34 38 6.53122 $w=7.58e-07 $l=4.15e-07 $layer=LI1_cond $X=1.2 $Y=0.295
+ $X2=1.615 $Y2=0.295
r49 34 36 12.2087 $w=7.58e-07 $l=2.3e-07 $layer=LI1_cond $X=1.2 $Y=0.295
+ $X2=0.97 $Y2=0.295
r50 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r51 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r52 29 45 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r53 28 42 56.107 $w=1.68e-07 $l=8.6e-07 $layer=LI1_cond $X=2.64 $Y=0 $X2=1.78
+ $Y2=0
r54 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r55 25 44 4.11661 $w=1.7e-07 $l=2.17e-07 $layer=LI1_cond $X=2.925 $Y=0 $X2=3.142
+ $Y2=0
r56 25 28 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=2.925 $Y=0 $X2=2.64
+ $Y2=0
r57 24 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r58 24 32 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r59 23 36 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=0.72 $Y=0 $X2=0.97
+ $Y2=0
r60 23 24 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r61 21 31 4.746 $w=1.7e-07 $l=2.2e-07 $layer=LI1_cond $X=0.44 $Y=0 $X2=0.22
+ $Y2=0
r62 21 23 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=0.44 $Y=0 $X2=0.72
+ $Y2=0
r63 18 29 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r64 18 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r65 18 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r66 14 44 3.16808 $w=2.7e-07 $l=1.19143e-07 $layer=LI1_cond $X=3.06 $Y=0.085
+ $X2=3.142 $Y2=0
r67 14 16 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=3.06 $Y=0.085
+ $X2=3.06 $Y2=0.38
r68 10 31 3.02018 $w=3.3e-07 $l=1.09087e-07 $layer=LI1_cond $X=0.275 $Y=0.085
+ $X2=0.22 $Y2=0
r69 10 12 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.275 $Y=0.085
+ $X2=0.275 $Y2=0.38
r70 3 16 91 $w=1.7e-07 $l=2.26164e-07 $layer=licon1_NDIFF $count=2 $X=2.865
+ $Y=0.235 $X2=3.03 $Y2=0.38
r71 2 38 91 $w=1.7e-07 $l=7.6138e-07 $layer=licon1_NDIFF $count=2 $X=0.995
+ $Y=0.235 $X2=1.615 $Y2=0.55
r72 1 12 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.15
+ $Y=0.235 $X2=0.275 $Y2=0.38
.ends

