# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__or4bb_m
  CLASS CORE ;
  FOREIGN sky130_fd_sc_lp__or4bb_m ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.320000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.035000 2.015000 3.505000 2.320000 ;
        RECT 3.035000 2.320000 3.205000 2.910000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.555000 0.975000 3.015000 1.485000 ;
    END
  END B
  PIN C_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.455000 0.775000 0.805000 1.445000 ;
    END
  END C_N
  PIN D_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.585000 2.005000 1.160000 2.525000 ;
    END
  END D_N
  PIN X
    ANTENNADIFFAREA  0.222600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.935000 2.320000 4.225000 2.910000 ;
        RECT 3.955000 0.345000 4.225000 0.675000 ;
        RECT 4.055000 0.675000 4.225000 2.320000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.320000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.320000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.320000 0.085000 ;
      RECT 0.000000  3.245000 4.320000 3.415000 ;
      RECT 0.105000  0.265000 0.480000 0.595000 ;
      RECT 0.105000  0.595000 0.275000 1.625000 ;
      RECT 0.105000  1.625000 2.375000 1.795000 ;
      RECT 0.105000  1.795000 0.365000 2.960000 ;
      RECT 0.585000  2.760000 0.775000 3.245000 ;
      RECT 0.700000  0.085000 0.910000 0.555000 ;
      RECT 1.015000  2.695000 1.735000 3.025000 ;
      RECT 1.130000  0.355000 1.340000 0.735000 ;
      RECT 1.130000  0.735000 1.705000 0.905000 ;
      RECT 1.535000  0.905000 1.705000 1.445000 ;
      RECT 1.650000  0.085000 1.860000 0.545000 ;
      RECT 1.700000  2.175000 2.855000 2.505000 ;
      RECT 2.080000  0.365000 2.290000 0.625000 ;
      RECT 2.080000  0.625000 3.365000 0.795000 ;
      RECT 2.205000  1.365000 2.375000 1.625000 ;
      RECT 2.470000  0.085000 2.800000 0.445000 ;
      RECT 2.685000  1.665000 3.875000 1.835000 ;
      RECT 2.685000  1.835000 2.855000 2.175000 ;
      RECT 3.020000  0.345000 3.365000 0.625000 ;
      RECT 3.195000  0.795000 3.365000 1.665000 ;
      RECT 3.385000  2.595000 3.715000 3.245000 ;
      RECT 3.545000  0.085000 3.735000 0.545000 ;
      RECT 3.705000  1.025000 3.875000 1.665000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
  END
END sky130_fd_sc_lp__or4bb_m
END LIBRARY
