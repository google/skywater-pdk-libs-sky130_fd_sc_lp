* File: sky130_fd_sc_lp__o2bb2ai_0.pex.spice
* Created: Fri Aug 28 11:12:26 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O2BB2AI_0%A1_N 2 5 7 8 11 15 17 18 19 20 21 22 23 31
r42 22 23 13.9805 $w=3.03e-07 $l=3.7e-07 $layer=LI1_cond $X=0.237 $Y=2.405
+ $X2=0.237 $Y2=2.775
r43 21 22 13.9805 $w=3.03e-07 $l=3.7e-07 $layer=LI1_cond $X=0.237 $Y=2.035
+ $X2=0.237 $Y2=2.405
r44 20 21 13.9805 $w=3.03e-07 $l=3.7e-07 $layer=LI1_cond $X=0.237 $Y=1.665
+ $X2=0.237 $Y2=2.035
r45 19 20 13.9805 $w=3.03e-07 $l=3.7e-07 $layer=LI1_cond $X=0.237 $Y=1.295
+ $X2=0.237 $Y2=1.665
r46 18 19 13.9805 $w=3.03e-07 $l=3.7e-07 $layer=LI1_cond $X=0.237 $Y=0.925
+ $X2=0.237 $Y2=1.295
r47 18 31 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.27
+ $Y=1.005 $X2=0.27 $Y2=1.005
r48 16 31 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.27 $Y=1.345
+ $X2=0.27 $Y2=1.005
r49 16 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.27 $Y=1.345
+ $X2=0.27 $Y2=1.51
r50 15 31 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=0.27 $Y=0.99
+ $X2=0.27 $Y2=1.005
r51 14 15 43.5886 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=0.345 $Y=0.84
+ $X2=0.345 $Y2=0.99
r52 9 11 243.564 $w=1.5e-07 $l=4.75e-07 $layer=POLY_cond $X=1.065 $Y=2.26
+ $X2=1.065 $Y2=2.735
r53 7 9 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.99 $Y=2.185
+ $X2=1.065 $Y2=2.26
r54 7 8 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=0.99 $Y=2.185
+ $X2=0.435 $Y2=2.185
r55 5 14 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=0.51 $Y=0.49 $X2=0.51
+ $Y2=0.84
r56 2 8 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.36 $Y=2.11
+ $X2=0.435 $Y2=2.185
r57 2 17 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=0.36 $Y=2.11 $X2=0.36
+ $Y2=1.51
.ends

.subckt PM_SKY130_FD_SC_LP__O2BB2AI_0%A2_N 3 5 6 9 13 14 15 16 17 23
r52 23 24 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.84
+ $Y=1.395 $X2=0.84 $Y2=1.395
r53 16 17 9.91637 $w=4.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.79 $Y=1.665
+ $X2=0.79 $Y2=2.035
r54 16 24 7.23627 $w=4.28e-07 $l=2.7e-07 $layer=LI1_cond $X=0.79 $Y=1.665
+ $X2=0.79 $Y2=1.395
r55 15 24 2.6801 $w=4.28e-07 $l=1e-07 $layer=LI1_cond $X=0.79 $Y=1.295 $X2=0.79
+ $Y2=1.395
r56 14 15 9.91637 $w=4.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.79 $Y=0.925
+ $X2=0.79 $Y2=1.295
r57 13 23 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=0.84 $Y=1.75
+ $X2=0.84 $Y2=1.395
r58 12 23 41.8716 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.84 $Y=1.23
+ $X2=0.84 $Y2=1.395
r59 7 9 428.16 $w=1.5e-07 $l=8.35e-07 $layer=POLY_cond $X=1.495 $Y=1.9 $X2=1.495
+ $Y2=2.735
r60 6 13 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=1.005 $Y=1.825
+ $X2=0.84 $Y2=1.75
r61 5 7 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.42 $Y=1.825
+ $X2=1.495 $Y2=1.9
r62 5 6 212.798 $w=1.5e-07 $l=4.15e-07 $layer=POLY_cond $X=1.42 $Y=1.825
+ $X2=1.005 $Y2=1.825
r63 3 12 379.447 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=0.9 $Y=0.49 $X2=0.9
+ $Y2=1.23
.ends

.subckt PM_SKY130_FD_SC_LP__O2BB2AI_0%A_195_56# 1 2 7 8 11 15 18 19 21 26 32 34
+ 36 37 38 39
c74 8 0 2.57313e-20 $X=1.545 $Y=0.885
r75 36 38 8.48848 $w=3.48e-07 $l=1.65e-07 $layer=LI1_cond $X=1.37 $Y=0.975
+ $X2=1.37 $Y2=0.81
r76 36 37 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.38
+ $Y=0.975 $X2=1.38 $Y2=0.975
r77 34 39 58.0813 $w=1.88e-07 $l=9.95e-07 $layer=LI1_cond $X=1.29 $Y=2.395
+ $X2=1.29 $Y2=1.4
r78 30 32 5.76222 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=1.115 $Y=0.49
+ $X2=1.28 $Y2=0.49
r79 26 39 8.15412 $w=3.48e-07 $l=1.75e-07 $layer=LI1_cond $X=1.37 $Y=1.225
+ $X2=1.37 $Y2=1.4
r80 25 36 0.329269 $w=3.48e-07 $l=1e-08 $layer=LI1_cond $X=1.37 $Y=0.985
+ $X2=1.37 $Y2=0.975
r81 25 26 7.90247 $w=3.48e-07 $l=2.4e-07 $layer=LI1_cond $X=1.37 $Y=0.985
+ $X2=1.37 $Y2=1.225
r82 23 32 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.28 $Y=0.655
+ $X2=1.28 $Y2=0.49
r83 23 38 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=1.28 $Y=0.655
+ $X2=1.28 $Y2=0.81
r84 19 34 6.19398 $w=2.33e-07 $l=1.17e-07 $layer=LI1_cond $X=1.267 $Y=2.512
+ $X2=1.267 $Y2=2.395
r85 19 21 2.35393 $w=2.33e-07 $l=4.8e-08 $layer=LI1_cond $X=1.267 $Y=2.512
+ $X2=1.267 $Y2=2.56
r86 17 37 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=1.38 $Y=0.96
+ $X2=1.38 $Y2=0.975
r87 13 18 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.925 $Y=0.96
+ $X2=1.925 $Y2=0.885
r88 13 15 910.16 $w=1.5e-07 $l=1.775e-06 $layer=POLY_cond $X=1.925 $Y=0.96
+ $X2=1.925 $Y2=2.735
r89 9 18 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.925 $Y=0.81
+ $X2=1.925 $Y2=0.885
r90 9 11 187.16 $w=1.5e-07 $l=3.65e-07 $layer=POLY_cond $X=1.925 $Y=0.81
+ $X2=1.925 $Y2=0.445
r91 8 17 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=1.545 $Y=0.885
+ $X2=1.38 $Y2=0.96
r92 7 18 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.85 $Y=0.885
+ $X2=1.925 $Y2=0.885
r93 7 8 156.394 $w=1.5e-07 $l=3.05e-07 $layer=POLY_cond $X=1.85 $Y=0.885
+ $X2=1.545 $Y2=0.885
r94 2 21 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=1.14
+ $Y=2.415 $X2=1.28 $Y2=2.56
r95 1 30 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.975
+ $Y=0.28 $X2=1.115 $Y2=0.49
.ends

.subckt PM_SKY130_FD_SC_LP__O2BB2AI_0%B2 3 7 11 12 13 14 18
c42 18 0 1.77059e-19 $X=2.405 $Y=1.32
c43 12 0 1.77059e-19 $X=2.405 $Y=1.825
c44 11 0 3.17149e-19 $X=2.405 $Y=1.66
c45 7 0 8.03548e-20 $X=2.395 $Y=0.445
r46 18 19 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.405
+ $Y=1.32 $X2=2.405 $Y2=1.32
r47 14 19 9.35513 $w=4.23e-07 $l=3.45e-07 $layer=LI1_cond $X=2.277 $Y=1.665
+ $X2=2.277 $Y2=1.32
r48 13 19 0.677908 $w=4.23e-07 $l=2.5e-08 $layer=LI1_cond $X=2.277 $Y=1.295
+ $X2=2.277 $Y2=1.32
r49 11 18 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.405 $Y=1.66
+ $X2=2.405 $Y2=1.32
r50 11 12 40.8701 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.405 $Y=1.66
+ $X2=2.405 $Y2=1.825
r51 10 18 38.0424 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.405 $Y=1.155
+ $X2=2.405 $Y2=1.32
r52 7 10 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=2.395 $Y=0.445
+ $X2=2.395 $Y2=1.155
r53 3 12 466.617 $w=1.5e-07 $l=9.1e-07 $layer=POLY_cond $X=2.355 $Y=2.735
+ $X2=2.355 $Y2=1.825
.ends

.subckt PM_SKY130_FD_SC_LP__O2BB2AI_0%B1 3 7 11 14 16 17 19 20 21 22 23 24 29
c43 22 0 3.83247e-20 $X=3.12 $Y=1.295
c44 17 0 1.6034e-19 $X=2.855 $Y=0.915
c45 11 0 1.77746e-19 $X=2.885 $Y=2.065
r46 29 30 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.975
+ $Y=1.375 $X2=2.975 $Y2=1.375
r47 23 24 11.0754 $w=3.83e-07 $l=3.7e-07 $layer=LI1_cond $X=3.082 $Y=1.665
+ $X2=3.082 $Y2=2.035
r48 23 30 8.68074 $w=3.83e-07 $l=2.9e-07 $layer=LI1_cond $X=3.082 $Y=1.665
+ $X2=3.082 $Y2=1.375
r49 22 30 2.39469 $w=3.83e-07 $l=8e-08 $layer=LI1_cond $X=3.082 $Y=1.295
+ $X2=3.082 $Y2=1.375
r50 20 29 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.975 $Y=1.715
+ $X2=2.975 $Y2=1.375
r51 20 21 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.975 $Y=1.715
+ $X2=2.975 $Y2=1.88
r52 19 29 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.975 $Y=1.21
+ $X2=2.975 $Y2=1.375
r53 17 19 151.266 $w=1.5e-07 $l=2.95e-07 $layer=POLY_cond $X=2.885 $Y=0.915
+ $X2=2.885 $Y2=1.21
r54 16 17 47.3682 $w=2.1e-07 $l=1.5e-07 $layer=POLY_cond $X=2.855 $Y=0.765
+ $X2=2.855 $Y2=0.915
r55 12 14 71.7872 $w=1.5e-07 $l=1.4e-07 $layer=POLY_cond $X=2.745 $Y=2.14
+ $X2=2.885 $Y2=2.14
r56 11 14 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.885 $Y=2.065
+ $X2=2.885 $Y2=2.14
r57 11 21 94.8617 $w=1.5e-07 $l=1.85e-07 $layer=POLY_cond $X=2.885 $Y=2.065
+ $X2=2.885 $Y2=1.88
r58 7 16 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.825 $Y=0.445
+ $X2=2.825 $Y2=0.765
r59 1 12 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.745 $Y=2.215
+ $X2=2.745 $Y2=2.14
r60 1 3 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=2.745 $Y=2.215
+ $X2=2.745 $Y2=2.735
.ends

.subckt PM_SKY130_FD_SC_LP__O2BB2AI_0%VPWR 1 2 3 14 18 20 22 24 26 31 37 40 44
r44 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r45 37 38 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r46 35 44 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r47 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r48 32 40 8.23795 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=1.865 $Y=3.33
+ $X2=1.71 $Y2=3.33
r49 32 34 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=1.865 $Y=3.33
+ $X2=2.64 $Y2=3.33
r50 31 43 4.52492 $w=1.7e-07 $l=2.82e-07 $layer=LI1_cond $X=2.795 $Y=3.33
+ $X2=3.077 $Y2=3.33
r51 31 34 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=2.795 $Y=3.33
+ $X2=2.64 $Y2=3.33
r52 30 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r53 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r54 27 37 7.94884 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=0.98 $Y=3.33
+ $X2=0.832 $Y2=3.33
r55 27 29 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=0.98 $Y=3.33 $X2=1.2
+ $Y2=3.33
r56 26 40 8.23795 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=1.555 $Y=3.33
+ $X2=1.71 $Y2=3.33
r57 26 29 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=1.555 $Y=3.33
+ $X2=1.2 $Y2=3.33
r58 24 35 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r59 24 30 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r60 24 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r61 20 43 3.24126 $w=3.3e-07 $l=1.53734e-07 $layer=LI1_cond $X=2.96 $Y=3.245
+ $X2=3.077 $Y2=3.33
r62 20 22 23.9219 $w=3.28e-07 $l=6.85e-07 $layer=LI1_cond $X=2.96 $Y=3.245
+ $X2=2.96 $Y2=2.56
r63 16 40 0.701276 $w=3.1e-07 $l=8.5e-08 $layer=LI1_cond $X=1.71 $Y=3.245
+ $X2=1.71 $Y2=3.33
r64 16 18 25.4653 $w=3.08e-07 $l=6.85e-07 $layer=LI1_cond $X=1.71 $Y=3.245
+ $X2=1.71 $Y2=2.56
r65 12 37 0.543863 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=0.832 $Y=3.245
+ $X2=0.832 $Y2=3.33
r66 12 14 26.7601 $w=2.93e-07 $l=6.85e-07 $layer=LI1_cond $X=0.832 $Y=3.245
+ $X2=0.832 $Y2=2.56
r67 3 22 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=2.82
+ $Y=2.415 $X2=2.96 $Y2=2.56
r68 2 18 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=1.57
+ $Y=2.415 $X2=1.71 $Y2=2.56
r69 1 14 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.725
+ $Y=2.415 $X2=0.85 $Y2=2.56
.ends

.subckt PM_SKY130_FD_SC_LP__O2BB2AI_0%Y 1 2 9 11 16 18 19 29 31
c51 29 0 1.77059e-19 $X=1.725 $Y=1.57
c52 18 0 3.54117e-19 $X=1.595 $Y=1.58
c53 9 0 1.77746e-19 $X=2.17 $Y=2.175
r54 24 31 2.54215 $w=3.38e-07 $l=7.5e-08 $layer=LI1_cond $X=1.725 $Y=1.74
+ $X2=1.725 $Y2=1.665
r55 19 25 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=1.68 $Y=2.09
+ $X2=1.725 $Y2=2.09
r56 19 25 0.949071 $w=3.38e-07 $l=2.8e-08 $layer=LI1_cond $X=1.725 $Y=1.977
+ $X2=1.725 $Y2=2.005
r57 18 31 0.169477 $w=3.38e-07 $l=5e-09 $layer=LI1_cond $X=1.725 $Y=1.66
+ $X2=1.725 $Y2=1.665
r58 18 29 5.92976 $w=3.38e-07 $l=9e-08 $layer=LI1_cond $X=1.725 $Y=1.66
+ $X2=1.725 $Y2=1.57
r59 18 19 7.86373 $w=3.38e-07 $l=2.32e-07 $layer=LI1_cond $X=1.725 $Y=1.745
+ $X2=1.725 $Y2=1.977
r60 18 24 0.169477 $w=3.38e-07 $l=5e-09 $layer=LI1_cond $X=1.725 $Y=1.745
+ $X2=1.725 $Y2=1.74
r61 14 16 3.49225 $w=3.28e-07 $l=1e-07 $layer=LI1_cond $X=1.71 $Y=0.445 $X2=1.81
+ $Y2=0.445
r62 9 25 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=2.17 $Y=2.09
+ $X2=1.725 $Y2=2.09
r63 9 11 16.433 $w=2.68e-07 $l=3.85e-07 $layer=LI1_cond $X=2.17 $Y=2.175
+ $X2=2.17 $Y2=2.56
r64 7 16 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.81 $Y=0.61 $X2=1.81
+ $Y2=0.445
r65 7 29 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.81 $Y=0.61 $X2=1.81
+ $Y2=1.57
r66 2 11 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=2
+ $Y=2.415 $X2=2.14 $Y2=2.56
r67 1 14 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=1.585
+ $Y=0.235 $X2=1.71 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__O2BB2AI_0%VGND 1 2 7 9 13 15 17 27 28 34
c41 28 0 1.86071e-19 $X=3.12 $Y=0
r42 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r43 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r44 28 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.64
+ $Y2=0
r45 27 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r46 25 34 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.735 $Y=0 $X2=2.605
+ $Y2=0
r47 25 27 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=2.735 $Y=0 $X2=3.12
+ $Y2=0
r48 24 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r49 23 24 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r50 21 32 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r51 20 23 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=0.72 $Y=0 $X2=2.16
+ $Y2=0
r52 20 21 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r53 18 31 4.70058 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=0.46 $Y=0 $X2=0.23
+ $Y2=0
r54 18 20 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=0.46 $Y=0 $X2=0.72
+ $Y2=0
r55 17 34 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.475 $Y=0 $X2=2.605
+ $Y2=0
r56 17 23 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=2.475 $Y=0 $X2=2.16
+ $Y2=0
r57 15 24 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r58 15 21 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=0.72
+ $Y2=0
r59 11 34 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=2.605 $Y=0.085
+ $X2=2.605 $Y2=0
r60 11 13 15.9569 $w=2.58e-07 $l=3.6e-07 $layer=LI1_cond $X=2.605 $Y=0.085
+ $X2=2.605 $Y2=0.445
r61 7 31 3.0656 $w=3.3e-07 $l=1.12916e-07 $layer=LI1_cond $X=0.295 $Y=0.085
+ $X2=0.23 $Y2=0
r62 7 9 14.1436 $w=3.28e-07 $l=4.05e-07 $layer=LI1_cond $X=0.295 $Y=0.085
+ $X2=0.295 $Y2=0.49
r63 2 13 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.47
+ $Y=0.235 $X2=2.61 $Y2=0.445
r64 1 9 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.17
+ $Y=0.28 $X2=0.295 $Y2=0.49
.ends

.subckt PM_SKY130_FD_SC_LP__O2BB2AI_0%A_400_47# 1 2 9 11 12 15
c29 15 0 4.20301e-20 $X=3.04 $Y=0.445
r30 13 15 12.8689 $w=2.98e-07 $l=3.35e-07 $layer=LI1_cond $X=3.055 $Y=0.78
+ $X2=3.055 $Y2=0.445
r31 11 13 7.51767 $w=1.7e-07 $l=1.8775e-07 $layer=LI1_cond $X=2.905 $Y=0.865
+ $X2=3.055 $Y2=0.78
r32 11 12 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=2.905 $Y=0.865
+ $X2=2.305 $Y2=0.865
r33 7 12 7.07814 $w=1.7e-07 $l=1.56844e-07 $layer=LI1_cond $X=2.185 $Y=0.78
+ $X2=2.305 $Y2=0.865
r34 7 9 16.0862 $w=2.38e-07 $l=3.35e-07 $layer=LI1_cond $X=2.185 $Y=0.78
+ $X2=2.185 $Y2=0.445
r35 2 15 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.9
+ $Y=0.235 $X2=3.04 $Y2=0.445
r36 1 9 182 $w=1.7e-07 $l=2.86182e-07 $layer=licon1_NDIFF $count=1 $X=2 $Y=0.235
+ $X2=2.18 $Y2=0.445
.ends

