* File: sky130_fd_sc_lp__and4bb_1.pex.spice
* Created: Wed Sep  2 09:34:01 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__AND4BB_1%A_N 3 7 11 12 13 18 20 22
r42 20 22 0.785757 $w=4.38e-07 $l=3e-08 $layer=LI1_cond $X=0.66 $Y=2.005
+ $X2=0.66 $Y2=2.035
r43 18 19 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.525
+ $Y=1.835 $X2=0.525 $Y2=1.835
r44 12 20 1.08585 $w=4.4e-07 $l=2.8e-08 $layer=LI1_cond $X=0.66 $Y=1.977
+ $X2=0.66 $Y2=2.005
r45 12 19 4.63209 $w=3.74e-07 $l=1.42e-07 $layer=LI1_cond $X=0.66 $Y=1.977
+ $X2=0.66 $Y2=1.835
r46 12 13 8.98382 $w=4.38e-07 $l=3.43e-07 $layer=LI1_cond $X=0.66 $Y=2.062
+ $X2=0.66 $Y2=2.405
r47 12 22 0.707181 $w=4.38e-07 $l=2.7e-08 $layer=LI1_cond $X=0.66 $Y=2.062
+ $X2=0.66 $Y2=2.035
r48 11 18 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.525 $Y=2.175
+ $X2=0.525 $Y2=1.835
r49 10 18 40.8701 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.525 $Y=1.67
+ $X2=0.525 $Y2=1.835
r50 5 11 57.73 $w=2.63e-07 $l=3.3908e-07 $layer=POLY_cond $X=0.575 $Y=2.49
+ $X2=0.525 $Y2=2.175
r51 5 7 192.287 $w=1.5e-07 $l=3.75e-07 $layer=POLY_cond $X=0.575 $Y=2.49
+ $X2=0.575 $Y2=2.865
r52 3 10 617.883 $w=1.5e-07 $l=1.205e-06 $layer=POLY_cond $X=0.475 $Y=0.465
+ $X2=0.475 $Y2=1.67
.ends

.subckt PM_SKY130_FD_SC_LP__AND4BB_1%B_N 3 8 10 11 12 15 16 17
r47 15 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.995 $Y=0.95
+ $X2=0.995 $Y2=1.115
r48 15 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.995 $Y=0.95
+ $X2=0.995 $Y2=0.785
r49 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.995
+ $Y=0.95 $X2=0.995 $Y2=0.95
r50 12 16 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=0.72 $Y=0.95
+ $X2=0.995 $Y2=0.95
r51 10 11 58.3064 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=0.99 $Y=1.925
+ $X2=0.99 $Y2=2.075
r52 10 18 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=0.975 $Y=1.925
+ $X2=0.975 $Y2=1.115
r53 8 11 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.005 $Y=2.865
+ $X2=1.005 $Y2=2.075
r54 3 17 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.905 $Y=0.465
+ $X2=0.905 $Y2=0.785
.ends

.subckt PM_SKY130_FD_SC_LP__AND4BB_1%A_27_51# 1 2 7 11 15 17 20 23 28 31 35 37
+ 38 39
r78 37 38 10.0716 $w=1.88e-07 $l=1.7e-07 $layer=LI1_cond $X=0.925 $Y=1.472
+ $X2=1.095 $Y2=1.472
r79 32 35 6.46067 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=0.175 $Y=2.865
+ $X2=0.36 $Y2=2.865
r80 29 39 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=1.425 $Y=1.52
+ $X2=1.425 $Y2=1.43
r81 28 38 19.2632 $w=1.88e-07 $l=3.3e-07 $layer=LI1_cond $X=1.425 $Y=1.52
+ $X2=1.095 $Y2=1.52
r82 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.425
+ $Y=1.52 $X2=1.425 $Y2=1.52
r83 25 31 2.53056 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=0.39 $Y=1.415
+ $X2=0.24 $Y2=1.415
r84 25 37 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=0.39 $Y=1.415
+ $X2=0.925 $Y2=1.415
r85 23 32 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.175 $Y=2.7
+ $X2=0.175 $Y2=2.865
r86 22 31 3.91525 $w=2.35e-07 $l=1.12916e-07 $layer=LI1_cond $X=0.175 $Y=1.5
+ $X2=0.24 $Y2=1.415
r87 22 23 78.2888 $w=1.68e-07 $l=1.2e-06 $layer=LI1_cond $X=0.175 $Y=1.5
+ $X2=0.175 $Y2=2.7
r88 18 31 3.91525 $w=2.35e-07 $l=8.5e-08 $layer=LI1_cond $X=0.24 $Y=1.33
+ $X2=0.24 $Y2=1.415
r89 18 20 33.805 $w=2.98e-07 $l=8.8e-07 $layer=LI1_cond $X=0.24 $Y=1.33 $X2=0.24
+ $Y2=0.45
r90 13 17 20.4101 $w=1.5e-07 $l=9.08295e-08 $layer=POLY_cond $X=2.06 $Y=1.355
+ $X2=2.025 $Y2=1.43
r91 13 15 251.255 $w=1.5e-07 $l=4.9e-07 $layer=POLY_cond $X=2.06 $Y=1.355
+ $X2=2.06 $Y2=0.865
r92 9 17 20.4101 $w=1.5e-07 $l=9.08295e-08 $layer=POLY_cond $X=1.99 $Y=1.505
+ $X2=2.025 $Y2=1.43
r93 9 11 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=1.99 $Y=1.505
+ $X2=1.99 $Y2=2.175
r94 8 39 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.59 $Y=1.43
+ $X2=1.425 $Y2=1.43
r95 7 17 5.30422 $w=1.5e-07 $l=1.1e-07 $layer=POLY_cond $X=1.915 $Y=1.43
+ $X2=2.025 $Y2=1.43
r96 7 8 166.649 $w=1.5e-07 $l=3.25e-07 $layer=POLY_cond $X=1.915 $Y=1.43
+ $X2=1.59 $Y2=1.43
r97 2 35 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=0.235
+ $Y=2.655 $X2=0.36 $Y2=2.865
r98 1 20 182 $w=1.7e-07 $l=2.498e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.255 $X2=0.26 $Y2=0.45
.ends

.subckt PM_SKY130_FD_SC_LP__AND4BB_1%A_196_51# 1 2 9 11 15 18 19 20 23 24 26 27
+ 29 34
r82 33 34 3.80841 $w=3.58e-07 $l=8.5e-08 $layer=LI1_cond $X=1.415 $Y=0.435
+ $X2=1.5 $Y2=0.435
r83 31 33 9.44363 $w=3.58e-07 $l=2.95e-07 $layer=LI1_cond $X=1.12 $Y=0.435
+ $X2=1.415 $Y2=0.435
r84 28 29 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=1.855 $Y=1.255
+ $X2=1.855 $Y2=1.785
r85 26 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.77 $Y=1.17
+ $X2=1.855 $Y2=1.255
r86 26 27 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=1.77 $Y=1.17 $X2=1.5
+ $Y2=1.17
r87 24 37 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.51 $Y=0.38
+ $X2=2.51 $Y2=0.545
r88 23 34 46.5587 $w=2.48e-07 $l=1.01e-06 $layer=LI1_cond $X=2.51 $Y=0.38
+ $X2=1.5 $Y2=0.38
r89 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.51
+ $Y=0.38 $X2=2.51 $Y2=0.38
r90 19 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.77 $Y=1.87
+ $X2=1.855 $Y2=1.785
r91 19 20 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=1.77 $Y=1.87
+ $X2=1.385 $Y2=1.87
r92 18 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.415 $Y=1.085
+ $X2=1.5 $Y2=1.17
r93 17 33 5.14255 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=1.415 $Y=0.615
+ $X2=1.415 $Y2=0.435
r94 17 18 30.6631 $w=1.68e-07 $l=4.7e-07 $layer=LI1_cond $X=1.415 $Y=0.615
+ $X2=1.415 $Y2=1.085
r95 13 20 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=1.255 $Y=1.955
+ $X2=1.385 $Y2=1.87
r96 13 15 40.3355 $w=2.58e-07 $l=9.1e-07 $layer=LI1_cond $X=1.255 $Y=1.955
+ $X2=1.255 $Y2=2.865
r97 9 11 671.723 $w=1.5e-07 $l=1.31e-06 $layer=POLY_cond $X=2.42 $Y=0.865
+ $X2=2.42 $Y2=2.175
r98 9 37 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.42 $Y=0.865
+ $X2=2.42 $Y2=0.545
r99 2 15 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=1.08
+ $Y=2.655 $X2=1.22 $Y2=2.865
r100 1 31 182 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_NDIFF $count=1 $X=0.98
+ $Y=0.255 $X2=1.12 $Y2=0.45
.ends

.subckt PM_SKY130_FD_SC_LP__AND4BB_1%C 3 7 8 10 17 19
r35 17 20 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.87 $Y=1.35
+ $X2=2.87 $Y2=1.515
r36 17 19 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.87 $Y=1.35
+ $X2=2.87 $Y2=1.185
r37 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.87
+ $Y=1.35 $X2=2.87 $Y2=1.35
r38 10 18 3.90875 $w=7.63e-07 $l=2.5e-07 $layer=LI1_cond $X=3.12 $Y=1.132
+ $X2=2.87 $Y2=1.132
r39 8 18 3.59605 $w=7.63e-07 $l=2.3e-07 $layer=LI1_cond $X=2.64 $Y=1.132
+ $X2=2.87 $Y2=1.132
r40 7 19 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.96 $Y=0.865
+ $X2=2.96 $Y2=1.185
r41 3 20 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.89 $Y=2.175
+ $X2=2.89 $Y2=1.515
.ends

.subckt PM_SKY130_FD_SC_LP__AND4BB_1%D 3 6 7 13
r27 10 13 24.4806 $w=3.3e-07 $l=1.4e-07 $layer=POLY_cond $X=3.18 $Y=2.92
+ $X2=3.32 $Y2=2.92
r28 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.18
+ $Y=2.92 $X2=3.18 $Y2=2.92
r29 7 11 4.64178 $w=3.58e-07 $l=1.45e-07 $layer=LI1_cond $X=3.165 $Y=2.775
+ $X2=3.165 $Y2=2.92
r30 3 6 671.723 $w=1.5e-07 $l=1.31e-06 $layer=POLY_cond $X=3.32 $Y=0.865
+ $X2=3.32 $Y2=2.175
r31 1 13 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.32 $Y=2.755
+ $X2=3.32 $Y2=2.92
r32 1 6 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=3.32 $Y=2.755 $X2=3.32
+ $Y2=2.175
.ends

.subckt PM_SKY130_FD_SC_LP__AND4BB_1%A_344_131# 1 2 3 12 16 18 23 26 28 32 34 38
+ 39 41 42
r74 39 45 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.77 $Y=1.51
+ $X2=3.77 $Y2=1.675
r75 39 44 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.77 $Y=1.51
+ $X2=3.77 $Y2=1.345
r76 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.77
+ $Y=1.51 $X2=3.77 $Y2=1.51
r77 36 38 8.98906 $w=2.48e-07 $l=1.95e-07 $layer=LI1_cond $X=3.73 $Y=1.705
+ $X2=3.73 $Y2=1.51
r78 35 42 7.13466 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=3.24 $Y=1.79
+ $X2=3.112 $Y2=1.79
r79 34 36 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.605 $Y=1.79
+ $X2=3.73 $Y2=1.705
r80 34 35 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=3.605 $Y=1.79
+ $X2=3.24 $Y2=1.79
r81 30 42 0.067832 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=3.112 $Y=1.875
+ $X2=3.112 $Y2=1.79
r82 30 32 13.5582 $w=2.53e-07 $l=3e-07 $layer=LI1_cond $X=3.112 $Y=1.875
+ $X2=3.112 $Y2=2.175
r83 29 41 1.97946 $w=1.7e-07 $l=1.03e-07 $layer=LI1_cond $X=2.315 $Y=1.79
+ $X2=2.212 $Y2=1.79
r84 28 42 7.13466 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=2.985 $Y=1.79
+ $X2=3.112 $Y2=1.79
r85 28 29 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.985 $Y=1.79
+ $X2=2.315 $Y2=1.79
r86 24 41 4.45556 $w=2.02e-07 $l=8.5e-08 $layer=LI1_cond $X=2.212 $Y=1.875
+ $X2=2.212 $Y2=1.79
r87 24 26 16.2306 $w=2.03e-07 $l=3e-07 $layer=LI1_cond $X=2.212 $Y=1.875
+ $X2=2.212 $Y2=2.175
r88 23 41 4.45556 $w=2.02e-07 $l=8.59942e-08 $layer=LI1_cond $X=2.21 $Y=1.705
+ $X2=2.212 $Y2=1.79
r89 22 23 43.8091 $w=1.98e-07 $l=7.9e-07 $layer=LI1_cond $X=2.21 $Y=0.915
+ $X2=2.21 $Y2=1.705
r90 18 22 6.89002 $w=2.4e-07 $l=1.62481e-07 $layer=LI1_cond $X=2.11 $Y=0.795
+ $X2=2.21 $Y2=0.915
r91 18 20 12.7249 $w=2.38e-07 $l=2.65e-07 $layer=LI1_cond $X=2.11 $Y=0.795
+ $X2=1.845 $Y2=0.795
r92 16 45 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.845 $Y=2.465
+ $X2=3.845 $Y2=1.675
r93 12 44 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.845 $Y=0.655
+ $X2=3.845 $Y2=1.345
r94 3 32 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=2.965
+ $Y=1.965 $X2=3.105 $Y2=2.175
r95 2 26 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=2.065
+ $Y=1.965 $X2=2.205 $Y2=2.175
r96 1 20 182 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=1 $X=1.72
+ $Y=0.655 $X2=1.845 $Y2=0.82
.ends

.subckt PM_SKY130_FD_SC_LP__AND4BB_1%VPWR 1 2 3 4 15 17 21 25 30 32 35 37 42 47
+ 54 55 58 61 64 67
r58 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r59 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r60 61 62 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r61 59 62 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r62 58 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r63 55 68 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.6 $Y2=3.33
r64 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r65 52 67 6.81202 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=3.755 $Y=3.33
+ $X2=3.635 $Y2=3.33
r66 52 54 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=3.755 $Y=3.33
+ $X2=4.08 $Y2=3.33
r67 51 68 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r68 51 65 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.64 $Y2=3.33
r69 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r70 48 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.815 $Y=3.33
+ $X2=2.65 $Y2=3.33
r71 48 50 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.815 $Y=3.33
+ $X2=3.12 $Y2=3.33
r72 47 67 6.81202 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=3.515 $Y=3.33
+ $X2=3.635 $Y2=3.33
r73 47 50 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=3.515 $Y=3.33
+ $X2=3.12 $Y2=3.33
r74 43 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.94 $Y=3.33
+ $X2=1.775 $Y2=3.33
r75 43 45 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=1.94 $Y=3.33
+ $X2=2.16 $Y2=3.33
r76 42 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.485 $Y=3.33
+ $X2=2.65 $Y2=3.33
r77 42 45 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=2.485 $Y=3.33
+ $X2=2.16 $Y2=3.33
r78 40 59 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r79 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r80 37 58 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.625 $Y=3.33
+ $X2=0.79 $Y2=3.33
r81 37 39 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=0.625 $Y=3.33
+ $X2=0.24 $Y2=3.33
r82 35 65 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r83 35 62 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r84 35 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r85 32 34 6.59091 $w=3.43e-07 $l=1.65e-07 $layer=LI1_cond $X=3.582 $Y=2.21
+ $X2=3.582 $Y2=2.375
r86 30 34 11.2843 $w=2.38e-07 $l=2.35e-07 $layer=LI1_cond $X=3.635 $Y=2.61
+ $X2=3.635 $Y2=2.375
r87 28 67 0.135687 $w=2.4e-07 $l=8.5e-08 $layer=LI1_cond $X=3.635 $Y=3.245
+ $X2=3.635 $Y2=3.33
r88 28 30 30.4917 $w=2.38e-07 $l=6.35e-07 $layer=LI1_cond $X=3.635 $Y=3.245
+ $X2=3.635 $Y2=2.61
r89 23 64 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.65 $Y=3.245
+ $X2=2.65 $Y2=3.33
r90 23 25 37.3671 $w=3.28e-07 $l=1.07e-06 $layer=LI1_cond $X=2.65 $Y=3.245
+ $X2=2.65 $Y2=2.175
r91 19 61 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.775 $Y=3.245
+ $X2=1.775 $Y2=3.33
r92 19 21 35.4464 $w=3.28e-07 $l=1.015e-06 $layer=LI1_cond $X=1.775 $Y=3.245
+ $X2=1.775 $Y2=2.23
r93 18 58 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.955 $Y=3.33
+ $X2=0.79 $Y2=3.33
r94 17 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.61 $Y=3.33
+ $X2=1.775 $Y2=3.33
r95 17 18 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=1.61 $Y=3.33
+ $X2=0.955 $Y2=3.33
r96 13 58 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.79 $Y=3.245
+ $X2=0.79 $Y2=3.33
r97 13 15 13.2706 $w=3.28e-07 $l=3.8e-07 $layer=LI1_cond $X=0.79 $Y=3.245
+ $X2=0.79 $Y2=2.865
r98 4 32 600 $w=1.7e-07 $l=3.07124e-07 $layer=licon1_PDIFF $count=1 $X=3.395
+ $Y=1.965 $X2=3.535 $Y2=2.21
r99 4 30 300 $w=1.7e-07 $l=7.53392e-07 $layer=licon1_PDIFF $count=2 $X=3.395
+ $Y=1.965 $X2=3.63 $Y2=2.61
r100 3 25 600 $w=1.7e-07 $l=2.76857e-07 $layer=licon1_PDIFF $count=1 $X=2.495
+ $Y=1.965 $X2=2.65 $Y2=2.175
r101 2 21 600 $w=1.7e-07 $l=3.21481e-07 $layer=licon1_PDIFF $count=1 $X=1.65
+ $Y=1.965 $X2=1.775 $Y2=2.23
r102 1 15 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=0.65
+ $Y=2.655 $X2=0.79 $Y2=2.865
.ends

.subckt PM_SKY130_FD_SC_LP__AND4BB_1%X 1 2 7 9 15 16 17 23 29
r20 21 29 0.557634 $w=3.08e-07 $l=1.5e-08 $layer=LI1_cond $X=4.08 $Y=0.94
+ $X2=4.08 $Y2=0.925
r21 17 31 5.66655 $w=3.08e-07 $l=1.2e-07 $layer=LI1_cond $X=4.08 $Y=0.975
+ $X2=4.08 $Y2=1.095
r22 17 21 1.30115 $w=3.08e-07 $l=3.5e-08 $layer=LI1_cond $X=4.08 $Y=0.975
+ $X2=4.08 $Y2=0.94
r23 17 29 1.30115 $w=3.08e-07 $l=3.5e-08 $layer=LI1_cond $X=4.08 $Y=0.89
+ $X2=4.08 $Y2=0.925
r24 16 17 12.4538 $w=3.08e-07 $l=3.35e-07 $layer=LI1_cond $X=4.08 $Y=0.555
+ $X2=4.08 $Y2=0.89
r25 16 23 5.0187 $w=3.08e-07 $l=1.35e-07 $layer=LI1_cond $X=4.08 $Y=0.555
+ $X2=4.08 $Y2=0.42
r26 15 31 49.645 $w=2.08e-07 $l=9.4e-07 $layer=LI1_cond $X=4.13 $Y=2.035
+ $X2=4.13 $Y2=1.095
r27 9 11 26.3947 $w=3.08e-07 $l=7.1e-07 $layer=LI1_cond $X=4.08 $Y=2.2 $X2=4.08
+ $Y2=2.91
r28 7 15 6.96769 $w=3.08e-07 $l=1.55e-07 $layer=LI1_cond $X=4.08 $Y=2.19
+ $X2=4.08 $Y2=2.035
r29 7 9 0.371756 $w=3.08e-07 $l=1e-08 $layer=LI1_cond $X=4.08 $Y=2.19 $X2=4.08
+ $Y2=2.2
r30 2 11 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=3.92
+ $Y=1.835 $X2=4.06 $Y2=2.91
r31 2 9 400 $w=1.7e-07 $l=4.29331e-07 $layer=licon1_PDIFF $count=1 $X=3.92
+ $Y=1.835 $X2=4.06 $Y2=2.2
r32 1 23 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=3.92
+ $Y=0.235 $X2=4.06 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__AND4BB_1%VGND 1 2 9 13 17 19 24 34 35 38 41
r41 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r42 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r43 35 42 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.6
+ $Y2=0
r44 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r45 32 41 8.42608 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=3.755 $Y=0 $X2=3.595
+ $Y2=0
r46 32 34 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=3.755 $Y=0 $X2=4.08
+ $Y2=0
r47 31 42 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r48 30 31 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r49 28 39 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r50 27 30 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=3.12
+ $Y2=0
r51 27 28 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r52 25 38 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.82 $Y=0 $X2=0.69
+ $Y2=0
r53 25 27 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=0.82 $Y=0 $X2=1.2
+ $Y2=0
r54 24 41 8.42608 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=3.435 $Y=0 $X2=3.595
+ $Y2=0
r55 24 30 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=3.435 $Y=0 $X2=3.12
+ $Y2=0
r56 22 39 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r57 21 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r58 19 38 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.56 $Y=0 $X2=0.69
+ $Y2=0
r59 19 21 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=0.56 $Y=0 $X2=0.24
+ $Y2=0
r60 17 31 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r61 17 28 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.2
+ $Y2=0
r62 13 15 19.8076 $w=3.18e-07 $l=5.5e-07 $layer=LI1_cond $X=3.595 $Y=0.38
+ $X2=3.595 $Y2=0.93
r63 11 41 0.800721 $w=3.2e-07 $l=8.5e-08 $layer=LI1_cond $X=3.595 $Y=0.085
+ $X2=3.595 $Y2=0
r64 11 13 10.6241 $w=3.18e-07 $l=2.95e-07 $layer=LI1_cond $X=3.595 $Y=0.085
+ $X2=3.595 $Y2=0.38
r65 7 38 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=0.085
+ $X2=0.69 $Y2=0
r66 7 9 16.1785 $w=2.58e-07 $l=3.65e-07 $layer=LI1_cond $X=0.69 $Y=0.085
+ $X2=0.69 $Y2=0.45
r67 2 15 182 $w=1.7e-07 $l=3.51781e-07 $layer=licon1_NDIFF $count=1 $X=3.395
+ $Y=0.655 $X2=3.57 $Y2=0.93
r68 2 13 182 $w=1.7e-07 $l=3.745e-07 $layer=licon1_NDIFF $count=1 $X=3.395
+ $Y=0.655 $X2=3.63 $Y2=0.38
r69 1 9 182 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.255 $X2=0.69 $Y2=0.45
.ends

