* File: sky130_fd_sc_lp__dlygate4s15_1.spice
* Created: Wed Sep  2 09:49:58 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__dlygate4s15_1.pex.spice"
.subckt sky130_fd_sc_lp__dlygate4s15_1  VNB VPB A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* VPB	VPB
* VNB	VNB
MM1005 N_VGND_M1005_d N_A_M1005_g N_A_27_52#_M1005_s VNB NSHORT L=0.15 W=0.42
+ AD=0.1554 AS=0.1113 PD=1.16 PS=1.37 NRD=15.708 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1002 N_A_288_52#_M1002_d N_A_27_52#_M1002_g N_VGND_M1005_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1113 AS=0.1554 PD=1.37 PS=1.16 NRD=0 NRS=115.704 M=1 R=2.8
+ SA=75001.1 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1006 N_VGND_M1006_d N_A_288_52#_M1006_g N_A_405_136#_M1006_s VNB NSHORT L=0.15
+ W=0.42 AD=0.1337 AS=0.1113 PD=1.02 PS=1.37 NRD=118.56 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001 A=0.063 P=1.14 MULT=1
MM1001 N_X_M1001_d N_A_405_136#_M1001_g N_VGND_M1006_d VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.2674 PD=2.21 PS=2.04 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1004 N_VPWR_M1004_d N_A_M1004_g N_A_27_52#_M1004_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.1554 AS=0.1113 PD=1.16 PS=1.37 NRD=21.0987 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1000 N_A_288_52#_M1000_d N_A_27_52#_M1000_g N_VPWR_M1004_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1113 AS=0.1554 PD=1.37 PS=1.16 NRD=0 NRS=194.636 M=1 R=2.8
+ SA=75001.1 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1007 N_VPWR_M1007_d N_A_288_52#_M1007_g N_A_405_136#_M1007_s VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.1281 AS=0.1113 PD=0.975 PS=1.37 NRD=194.636 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001 A=0.063 P=1.14 MULT=1
MM1003 N_X_M1003_d N_A_405_136#_M1003_g N_VPWR_M1007_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.3843 PD=3.05 PS=2.925 NRD=0 NRS=0 M=1 R=8.4 SA=75000.5
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX8_noxref VNB VPB NWDIODE A=7.8703 P=12.17
c_36 VNB 0 1.65637e-19 $X=0 $Y=0
*
.include "sky130_fd_sc_lp__dlygate4s15_1.pxi.spice"
*
.ends
*
*
