* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__nand3b_4 A_N B C VGND VNB VPB VPWR Y
X0 VGND C a_652_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X1 Y a_35_74# a_225_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X2 a_225_47# B a_652_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X3 Y a_35_74# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X4 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X5 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X6 a_652_47# C VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X7 VGND C a_652_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X8 a_652_47# B a_225_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X9 a_35_74# A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X10 a_652_47# C VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X11 a_35_74# A_N VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X12 Y a_35_74# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X13 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X14 VPWR a_35_74# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X15 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X16 a_225_47# a_35_74# Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X17 Y a_35_74# a_225_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X18 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X19 a_225_47# a_35_74# Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X20 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X21 a_225_47# B a_652_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X22 VPWR a_35_74# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X23 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X24 a_652_47# B a_225_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X25 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
.ends
