* File: sky130_fd_sc_lp__o22ai_0.pex.spice
* Created: Fri Aug 28 11:10:22 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O22AI_0%B1 3 5 8 12 14 15 16 17 23 25
c37 25 0 3.52235e-20 $X=0.345 $Y=0.955
c38 14 0 2.97974e-20 $X=0.24 $Y=0.925
r39 23 26 88.3231 $w=4.6e-07 $l=5.05e-07 $layer=POLY_cond $X=0.345 $Y=1.12
+ $X2=0.345 $Y2=1.625
r40 23 25 47.2161 $w=4.6e-07 $l=1.65e-07 $layer=POLY_cond $X=0.345 $Y=1.12
+ $X2=0.345 $Y2=0.955
r41 23 24 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.28
+ $Y=1.12 $X2=0.28 $Y2=1.12
r42 16 17 14.2135 $w=2.98e-07 $l=3.7e-07 $layer=LI1_cond $X=0.235 $Y=1.665
+ $X2=0.235 $Y2=2.035
r43 15 16 14.2135 $w=2.98e-07 $l=3.7e-07 $layer=LI1_cond $X=0.235 $Y=1.295
+ $X2=0.235 $Y2=1.665
r44 15 24 6.72258 $w=2.98e-07 $l=1.75e-07 $layer=LI1_cond $X=0.235 $Y=1.295
+ $X2=0.235 $Y2=1.12
r45 14 24 7.49088 $w=2.98e-07 $l=1.95e-07 $layer=LI1_cond $X=0.235 $Y=0.925
+ $X2=0.235 $Y2=1.12
r46 10 12 71.7872 $w=1.5e-07 $l=1.4e-07 $layer=POLY_cond $X=0.5 $Y=2.195
+ $X2=0.64 $Y2=2.195
r47 6 12 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.64 $Y=2.27 $X2=0.64
+ $Y2=2.195
r48 6 8 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=0.64 $Y=2.27 $X2=0.64
+ $Y2=2.735
r49 5 10 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.5 $Y=2.12 $X2=0.5
+ $Y2=2.195
r50 5 26 253.819 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=0.5 $Y=2.12 $X2=0.5
+ $Y2=1.625
r51 3 25 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.5 $Y=0.635 $X2=0.5
+ $Y2=0.955
.ends

.subckt PM_SKY130_FD_SC_LP__O22AI_0%B2 3 7 11 12 13 14 15 20
c44 20 0 7.8289e-20 $X=0.98 $Y=1.375
c45 12 0 1.83811e-19 $X=0.98 $Y=1.88
c46 3 0 1.91902e-19 $X=1.005 $Y=0.635
r47 20 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.98
+ $Y=1.375 $X2=0.98 $Y2=1.375
r48 14 15 10.6601 $w=3.98e-07 $l=3.7e-07 $layer=LI1_cond $X=1.095 $Y=1.665
+ $X2=1.095 $Y2=2.035
r49 14 21 8.35521 $w=3.98e-07 $l=2.9e-07 $layer=LI1_cond $X=1.095 $Y=1.665
+ $X2=1.095 $Y2=1.375
r50 13 21 2.30489 $w=3.98e-07 $l=8e-08 $layer=LI1_cond $X=1.095 $Y=1.295
+ $X2=1.095 $Y2=1.375
r51 11 20 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.98 $Y=1.715
+ $X2=0.98 $Y2=1.375
r52 11 12 40.8701 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.98 $Y=1.715
+ $X2=0.98 $Y2=1.88
r53 10 20 38.9318 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.98 $Y=1.21
+ $X2=0.98 $Y2=1.375
r54 7 12 438.415 $w=1.5e-07 $l=8.55e-07 $layer=POLY_cond $X=1.03 $Y=2.735
+ $X2=1.03 $Y2=1.88
r55 3 10 294.84 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.005 $Y=0.635
+ $X2=1.005 $Y2=1.21
.ends

.subckt PM_SKY130_FD_SC_LP__O22AI_0%A2 3 7 9 10 11 16
c39 7 0 6.95905e-20 $X=1.46 $Y=2.735
c40 3 0 2.86929e-19 $X=1.46 $Y=0.635
r41 16 19 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.55 $Y=1.51
+ $X2=1.55 $Y2=1.675
r42 16 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.55 $Y=1.51
+ $X2=1.55 $Y2=1.345
r43 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.55
+ $Y=1.51 $X2=1.55 $Y2=1.51
r44 10 11 11.6823 $w=3.63e-07 $l=3.7e-07 $layer=LI1_cond $X=1.647 $Y=1.665
+ $X2=1.647 $Y2=2.035
r45 10 17 4.89394 $w=3.63e-07 $l=1.55e-07 $layer=LI1_cond $X=1.647 $Y=1.665
+ $X2=1.647 $Y2=1.51
r46 9 17 6.78836 $w=3.63e-07 $l=2.15e-07 $layer=LI1_cond $X=1.647 $Y=1.295
+ $X2=1.647 $Y2=1.51
r47 7 19 543.532 $w=1.5e-07 $l=1.06e-06 $layer=POLY_cond $X=1.46 $Y=2.735
+ $X2=1.46 $Y2=1.675
r48 3 18 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=1.46 $Y=0.635
+ $X2=1.46 $Y2=1.345
.ends

.subckt PM_SKY130_FD_SC_LP__O22AI_0%A1 3 5 7 8 9 12 14 15 16
c32 14 0 1.09219e-19 $X=2.16 $Y=1.295
r33 15 16 13.5366 $w=3.13e-07 $l=3.7e-07 $layer=LI1_cond $X=2.157 $Y=1.665
+ $X2=2.157 $Y2=2.035
r34 14 15 13.5366 $w=3.13e-07 $l=3.7e-07 $layer=LI1_cond $X=2.157 $Y=1.295
+ $X2=2.157 $Y2=1.665
r35 14 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.13
+ $Y=1.375 $X2=2.13 $Y2=1.375
r36 10 12 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=1.85 $Y=1.99
+ $X2=2.04 $Y2=1.99
r37 9 12 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.04 $Y=1.915
+ $X2=2.04 $Y2=1.99
r38 8 21 38.716 $w=2.81e-07 $l=1.80291e-07 $layer=POLY_cond $X=2.04 $Y=1.54
+ $X2=2.072 $Y2=1.375
r39 8 9 192.287 $w=1.5e-07 $l=3.75e-07 $layer=POLY_cond $X=2.04 $Y=1.54 $X2=2.04
+ $Y2=1.915
r40 5 21 82.4562 $w=2.81e-07 $l=4.87996e-07 $layer=POLY_cond $X=1.925 $Y=0.955
+ $X2=2.072 $Y2=1.375
r41 5 7 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.925 $Y=0.955
+ $X2=1.925 $Y2=0.635
r42 1 10 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.85 $Y=2.065
+ $X2=1.85 $Y2=1.99
r43 1 3 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=1.85 $Y=2.065 $X2=1.85
+ $Y2=2.735
.ends

.subckt PM_SKY130_FD_SC_LP__O22AI_0%VPWR 1 2 7 8 9 11 15 17 30
r31 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r32 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r33 24 30 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r34 23 24 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r35 21 27 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r36 20 23 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.72 $Y=3.33 $X2=1.68
+ $Y2=3.33
r37 20 21 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r38 18 26 5.96248 $w=1.7e-07 $l=2.95e-07 $layer=LI1_cond $X=0.59 $Y=3.33
+ $X2=0.295 $Y2=3.33
r39 18 20 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=0.59 $Y=3.33
+ $X2=0.72 $Y2=3.33
r40 17 29 4.31539 $w=1.7e-07 $l=2.32e-07 $layer=LI1_cond $X=1.935 $Y=3.33
+ $X2=2.167 $Y2=3.33
r41 17 23 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=1.935 $Y=3.33
+ $X2=1.68 $Y2=3.33
r42 15 24 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r43 15 21 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r44 9 29 3.16214 $w=2.95e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.082 $Y=3.245
+ $X2=2.167 $Y2=3.33
r45 9 11 26.7601 $w=2.93e-07 $l=6.85e-07 $layer=LI1_cond $X=2.082 $Y=3.245
+ $X2=2.082 $Y2=2.56
r46 8 26 2.97113 $w=4.65e-07 $l=1.11781e-07 $layer=LI1_cond $X=0.357 $Y=3.245
+ $X2=0.295 $Y2=3.33
r47 7 14 9.42339 $w=4.65e-07 $l=3.32e-07 $layer=LI1_cond $X=0.357 $Y=2.892
+ $X2=0.357 $Y2=2.56
r48 7 8 9.07991 $w=4.63e-07 $l=3.53e-07 $layer=LI1_cond $X=0.357 $Y=2.892
+ $X2=0.357 $Y2=3.245
r49 2 11 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=1.925
+ $Y=2.415 $X2=2.065 $Y2=2.56
r50 1 14 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.165
+ $Y=2.415 $X2=0.29 $Y2=2.56
.ends

.subckt PM_SKY130_FD_SC_LP__O22AI_0%Y 1 2 7 8 11 12 18
c39 18 0 3.59675e-19 $X=1.08 $Y=2.395
c40 7 0 1.77711e-19 $X=0.64 $Y=1.005
r41 12 29 2.70645 $w=6.83e-07 $l=1.55e-07 $layer=LI1_cond $X=1.422 $Y=2.405
+ $X2=1.422 $Y2=2.56
r42 12 18 0.17461 $w=6.83e-07 $l=1e-08 $layer=LI1_cond $X=1.422 $Y=2.405
+ $X2=1.422 $Y2=2.395
r43 11 19 3.23184 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=0.64 $Y=2.395
+ $X2=0.725 $Y2=2.395
r44 11 18 18.3876 $w=1.88e-07 $l=3.15e-07 $layer=LI1_cond $X=0.765 $Y=2.395
+ $X2=1.08 $Y2=2.395
r45 11 19 2.33493 $w=1.88e-07 $l=4e-08 $layer=LI1_cond $X=0.765 $Y=2.395
+ $X2=0.725 $Y2=2.395
r46 8 11 3.61205 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=0.64 $Y=2.3 $X2=0.64
+ $Y2=2.395
r47 7 10 13.765 $w=3.59e-07 $l=3.57911e-07 $layer=LI1_cond $X=0.64 $Y=1.005
+ $X2=0.755 $Y2=0.7
r48 7 8 84.4866 $w=1.68e-07 $l=1.295e-06 $layer=LI1_cond $X=0.64 $Y=1.005
+ $X2=0.64 $Y2=2.3
r49 2 29 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=1.105
+ $Y=2.415 $X2=1.245 $Y2=2.56
r50 1 10 182 $w=1.7e-07 $l=3.67083e-07 $layer=licon1_NDIFF $count=1 $X=0.575
+ $Y=0.425 $X2=0.79 $Y2=0.7
.ends

.subckt PM_SKY130_FD_SC_LP__O22AI_0%A_27_85# 1 2 3 10 15 16 17 20 22
c37 17 0 7.8289e-20 $X=1.355 $Y=0.955
r38 22 25 7.50834 $w=3.28e-07 $l=2.15e-07 $layer=LI1_cond $X=0.28 $Y=0.34
+ $X2=0.28 $Y2=0.555
r39 18 20 9.67229 $w=2.78e-07 $l=2.35e-07 $layer=LI1_cond $X=2.165 $Y=0.87
+ $X2=2.165 $Y2=0.635
r40 16 18 7.36005 $w=1.7e-07 $l=1.77482e-07 $layer=LI1_cond $X=2.025 $Y=0.955
+ $X2=2.165 $Y2=0.87
r41 16 17 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.025 $Y=0.955
+ $X2=1.355 $Y2=0.955
r42 13 17 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=1.245 $Y=0.87
+ $X2=1.355 $Y2=0.955
r43 13 15 12.3102 $w=2.18e-07 $l=2.35e-07 $layer=LI1_cond $X=1.245 $Y=0.87
+ $X2=1.245 $Y2=0.635
r44 12 15 11.0006 $w=2.18e-07 $l=2.1e-07 $layer=LI1_cond $X=1.245 $Y=0.425
+ $X2=1.245 $Y2=0.635
r45 11 22 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.445 $Y=0.34
+ $X2=0.28 $Y2=0.34
r46 10 12 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=1.135 $Y=0.34
+ $X2=1.245 $Y2=0.425
r47 10 11 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.135 $Y=0.34
+ $X2=0.445 $Y2=0.34
r48 3 20 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2
+ $Y=0.425 $X2=2.14 $Y2=0.635
r49 2 15 182 $w=1.7e-07 $l=2.78747e-07 $layer=licon1_NDIFF $count=1 $X=1.08
+ $Y=0.425 $X2=1.24 $Y2=0.635
r50 1 25 182 $w=1.7e-07 $l=1.99687e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.425 $X2=0.28 $Y2=0.555
.ends

.subckt PM_SKY130_FD_SC_LP__O22AI_0%VGND 1 6 8 10 20 21 24
c22 21 0 3.52235e-20 $X=2.16 $Y=0
c23 6 0 1.62105e-19 $X=1.69 $Y=0.59
r24 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r25 21 25 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.68
+ $Y2=0
r26 20 21 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r27 18 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.855 $Y=0 $X2=1.69
+ $Y2=0
r28 18 20 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.855 $Y=0 $X2=2.16
+ $Y2=0
r29 12 16 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r30 12 13 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r31 10 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.525 $Y=0 $X2=1.69
+ $Y2=0
r32 10 16 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=1.525 $Y=0 $X2=1.2
+ $Y2=0
r33 8 25 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r34 8 13 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.24
+ $Y2=0
r35 8 16 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r36 4 24 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.69 $Y=0.085 $X2=1.69
+ $Y2=0
r37 4 6 17.6359 $w=3.28e-07 $l=5.05e-07 $layer=LI1_cond $X=1.69 $Y=0.085
+ $X2=1.69 $Y2=0.59
r38 1 6 182 $w=1.7e-07 $l=2.29783e-07 $layer=licon1_NDIFF $count=1 $X=1.535
+ $Y=0.425 $X2=1.69 $Y2=0.59
.ends

