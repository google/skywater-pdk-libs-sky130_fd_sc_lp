* File: sky130_fd_sc_lp__a21oi_2.pxi.spice
* Created: Fri Aug 28 09:51:44 2020
* 
x_PM_SKY130_FD_SC_LP__A21OI_2%A2 N_A2_M1003_g N_A2_M1009_g N_A2_M1006_g
+ N_A2_M1010_g N_A2_c_62_n N_A2_c_63_n A2 N_A2_c_65_n N_A2_c_66_n
+ PM_SKY130_FD_SC_LP__A21OI_2%A2
x_PM_SKY130_FD_SC_LP__A21OI_2%A1 N_A1_c_129_n N_A1_M1007_g N_A1_M1000_g
+ N_A1_c_131_n N_A1_M1011_g N_A1_M1004_g A1 A1 N_A1_c_134_n
+ PM_SKY130_FD_SC_LP__A21OI_2%A1
x_PM_SKY130_FD_SC_LP__A21OI_2%B1 N_B1_M1002_g N_B1_M1001_g N_B1_M1008_g
+ N_B1_M1005_g B1 B1 N_B1_c_181_n PM_SKY130_FD_SC_LP__A21OI_2%B1
x_PM_SKY130_FD_SC_LP__A21OI_2%A_27_367# N_A_27_367#_M1009_d N_A_27_367#_M1000_s
+ N_A_27_367#_M1010_d N_A_27_367#_M1005_d N_A_27_367#_c_227_n
+ N_A_27_367#_c_228_n N_A_27_367#_c_233_n N_A_27_367#_c_252_p
+ N_A_27_367#_c_236_n N_A_27_367#_c_240_n N_A_27_367#_c_253_p
+ N_A_27_367#_c_229_n N_A_27_367#_c_230_n N_A_27_367#_c_241_n
+ PM_SKY130_FD_SC_LP__A21OI_2%A_27_367#
x_PM_SKY130_FD_SC_LP__A21OI_2%VPWR N_VPWR_M1009_s N_VPWR_M1004_d N_VPWR_c_269_n
+ N_VPWR_c_270_n VPWR N_VPWR_c_271_n N_VPWR_c_272_n N_VPWR_c_273_n
+ N_VPWR_c_268_n N_VPWR_c_275_n N_VPWR_c_276_n PM_SKY130_FD_SC_LP__A21OI_2%VPWR
x_PM_SKY130_FD_SC_LP__A21OI_2%Y N_Y_M1007_d N_Y_M1002_d N_Y_M1001_s N_Y_c_318_n
+ N_Y_c_353_p N_Y_c_313_n N_Y_c_316_n N_Y_c_324_n N_Y_c_332_n N_Y_c_314_n Y Y
+ PM_SKY130_FD_SC_LP__A21OI_2%Y
x_PM_SKY130_FD_SC_LP__A21OI_2%VGND N_VGND_M1003_s N_VGND_M1006_s N_VGND_M1008_s
+ N_VGND_c_361_n N_VGND_c_362_n N_VGND_c_363_n N_VGND_c_364_n N_VGND_c_365_n
+ N_VGND_c_366_n N_VGND_c_367_n N_VGND_c_368_n VGND N_VGND_c_369_n
+ N_VGND_c_370_n PM_SKY130_FD_SC_LP__A21OI_2%VGND
x_PM_SKY130_FD_SC_LP__A21OI_2%A_110_47# N_A_110_47#_M1003_d N_A_110_47#_M1011_s
+ N_A_110_47#_c_406_n N_A_110_47#_c_412_n N_A_110_47#_c_408_n
+ PM_SKY130_FD_SC_LP__A21OI_2%A_110_47#
cc_1 VNB N_A2_M1003_g 0.0308122f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.655
cc_2 VNB N_A2_M1009_g 0.00167964f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.465
cc_3 VNB N_A2_M1006_g 0.0256976f $X=-0.19 $Y=-0.245 $X2=1.765 $Y2=0.655
cc_4 VNB N_A2_c_62_n 0.00704248f $X=-0.19 $Y=-0.245 $X2=1.525 $Y2=1.695
cc_5 VNB N_A2_c_63_n 0.005168f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.46
cc_6 VNB A2 0.00455627f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.58
cc_7 VNB N_A2_c_65_n 0.0541816f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.46
cc_8 VNB N_A2_c_66_n 0.0241592f $X=-0.19 $Y=-0.245 $X2=1.785 $Y2=1.51
cc_9 VNB N_A1_c_129_n 0.0164428f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.295
cc_10 VNB N_A1_M1000_g 0.00678716f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.465
cc_11 VNB N_A1_c_131_n 0.0164438f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A1_M1004_g 0.0063761f $X=-0.19 $Y=-0.245 $X2=1.805 $Y2=1.675
cc_13 VNB A1 0.00569679f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A1_c_134_n 0.0361364f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_B1_M1002_g 0.0251759f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.655
cc_16 VNB N_B1_M1008_g 0.0277011f $X=-0.19 $Y=-0.245 $X2=1.765 $Y2=0.655
cc_17 VNB B1 0.00572042f $X=-0.19 $Y=-0.245 $X2=0.455 $Y2=1.695
cc_18 VNB N_B1_c_181_n 0.0338851f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_VPWR_c_268_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_Y_c_313_n 0.0256103f $X=-0.19 $Y=-0.245 $X2=0.455 $Y2=1.695
cc_21 VNB N_Y_c_314_n 0.00284176f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.46
cc_22 VNB Y 0.0271736f $X=-0.19 $Y=-0.245 $X2=1.785 $Y2=1.51
cc_23 VNB N_VGND_c_361_n 0.0102287f $X=-0.19 $Y=-0.245 $X2=1.765 $Y2=0.655
cc_24 VNB N_VGND_c_362_n 0.0403734f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_363_n 4.02668e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_364_n 0.0261076f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.46
cc_27 VNB N_VGND_c_365_n 0.0348843f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.695
cc_28 VNB N_VGND_c_366_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_367_n 0.0133881f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_368_n 0.00513431f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.46
cc_31 VNB N_VGND_c_369_n 0.0121672f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_370_n 0.196391f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VPB N_A2_M1009_g 0.0247639f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.465
cc_34 VPB N_A2_M1010_g 0.01894f $X=-0.19 $Y=1.655 $X2=1.805 $Y2=2.465
cc_35 VPB N_A2_c_62_n 0.00619409f $X=-0.19 $Y=1.655 $X2=1.525 $Y2=1.695
cc_36 VPB N_A2_c_63_n 0.00739931f $X=-0.19 $Y=1.655 $X2=0.29 $Y2=1.46
cc_37 VPB A2 0.00191077f $X=-0.19 $Y=1.655 $X2=1.595 $Y2=1.58
cc_38 VPB N_A2_c_66_n 0.0061965f $X=-0.19 $Y=1.655 $X2=1.785 $Y2=1.51
cc_39 VPB N_A1_M1000_g 0.0186439f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.465
cc_40 VPB N_A1_M1004_g 0.0190258f $X=-0.19 $Y=1.655 $X2=1.805 $Y2=1.675
cc_41 VPB N_B1_M1001_g 0.0182394f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.465
cc_42 VPB N_B1_M1005_g 0.0224081f $X=-0.19 $Y=1.655 $X2=1.805 $Y2=2.465
cc_43 VPB B1 0.00726268f $X=-0.19 $Y=1.655 $X2=0.455 $Y2=1.695
cc_44 VPB N_B1_c_181_n 0.00486419f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_45 VPB N_A_27_367#_c_227_n 0.00849777f $X=-0.19 $Y=1.655 $X2=1.805 $Y2=1.675
cc_46 VPB N_A_27_367#_c_228_n 0.0360021f $X=-0.19 $Y=1.655 $X2=1.805 $Y2=2.465
cc_47 VPB N_A_27_367#_c_229_n 0.00746637f $X=-0.19 $Y=1.655 $X2=0.29 $Y2=1.46
cc_48 VPB N_A_27_367#_c_230_n 0.0242278f $X=-0.19 $Y=1.655 $X2=1.785 $Y2=1.51
cc_49 VPB N_VPWR_c_269_n 4.02668e-19 $X=-0.19 $Y=1.655 $X2=1.765 $Y2=1.345
cc_50 VPB N_VPWR_c_270_n 4.02668e-19 $X=-0.19 $Y=1.655 $X2=1.805 $Y2=1.675
cc_51 VPB N_VPWR_c_271_n 0.0153759f $X=-0.19 $Y=1.655 $X2=1.525 $Y2=1.695
cc_52 VPB N_VPWR_c_272_n 0.0133881f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_53 VPB N_VPWR_c_273_n 0.0418173f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=1.46
cc_54 VPB N_VPWR_c_268_n 0.0537912f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_55 VPB N_VPWR_c_275_n 0.00436868f $X=-0.19 $Y=1.655 $X2=1.785 $Y2=1.51
cc_56 VPB N_VPWR_c_276_n 0.00436868f $X=-0.19 $Y=1.655 $X2=1.697 $Y2=1.51
cc_57 VPB N_Y_c_316_n 0.0183542f $X=-0.19 $Y=1.655 $X2=0.29 $Y2=1.46
cc_58 VPB Y 0.0145346f $X=-0.19 $Y=1.655 $X2=1.785 $Y2=1.51
cc_59 N_A2_M1003_g N_A1_c_129_n 0.0257724f $X=0.475 $Y=0.655 $X2=-0.19
+ $Y2=-0.245
cc_60 N_A2_M1009_g N_A1_M1000_g 0.0257724f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_61 N_A2_c_62_n N_A1_M1000_g 0.0108336f $X=1.525 $Y=1.695 $X2=0 $Y2=0
cc_62 N_A2_M1006_g N_A1_c_131_n 0.0405834f $X=1.765 $Y=0.655 $X2=0 $Y2=0
cc_63 N_A2_M1010_g N_A1_M1004_g 0.0320246f $X=1.805 $Y=2.465 $X2=0 $Y2=0
cc_64 N_A2_c_62_n N_A1_M1004_g 0.0114482f $X=1.525 $Y=1.695 $X2=0 $Y2=0
cc_65 N_A2_M1003_g A1 0.00397177f $X=0.475 $Y=0.655 $X2=0 $Y2=0
cc_66 N_A2_M1006_g A1 7.66902e-19 $X=1.765 $Y=0.655 $X2=0 $Y2=0
cc_67 N_A2_c_62_n A1 0.0535137f $X=1.525 $Y=1.695 $X2=0 $Y2=0
cc_68 N_A2_c_63_n A1 0.0117208f $X=0.29 $Y=1.46 $X2=0 $Y2=0
cc_69 A2 A1 0.00752997f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_70 N_A2_c_62_n N_A1_c_134_n 0.00246815f $X=1.525 $Y=1.695 $X2=0 $Y2=0
cc_71 N_A2_c_63_n N_A1_c_134_n 0.00106093f $X=0.29 $Y=1.46 $X2=0 $Y2=0
cc_72 A2 N_A1_c_134_n 0.00489027f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_73 N_A2_c_65_n N_A1_c_134_n 0.0257724f $X=0.475 $Y=1.46 $X2=0 $Y2=0
cc_74 N_A2_c_66_n N_A1_c_134_n 0.020778f $X=1.785 $Y=1.51 $X2=0 $Y2=0
cc_75 N_A2_M1006_g N_B1_M1002_g 0.0339979f $X=1.765 $Y=0.655 $X2=0 $Y2=0
cc_76 N_A2_M1010_g N_B1_M1001_g 0.0190708f $X=1.805 $Y=2.465 $X2=0 $Y2=0
cc_77 A2 N_B1_M1001_g 2.03567e-19 $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_78 N_A2_M1010_g B1 6.86664e-19 $X=1.805 $Y=2.465 $X2=0 $Y2=0
cc_79 A2 B1 0.0266409f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_80 N_A2_c_66_n B1 0.00179125f $X=1.785 $Y=1.51 $X2=0 $Y2=0
cc_81 A2 N_B1_c_181_n 7.22186e-19 $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_82 N_A2_c_66_n N_B1_c_181_n 0.0212337f $X=1.785 $Y=1.51 $X2=0 $Y2=0
cc_83 N_A2_c_63_n N_A_27_367#_c_227_n 0.020011f $X=0.29 $Y=1.46 $X2=0 $Y2=0
cc_84 N_A2_c_65_n N_A_27_367#_c_227_n 0.00121139f $X=0.475 $Y=1.46 $X2=0 $Y2=0
cc_85 N_A2_M1009_g N_A_27_367#_c_233_n 0.0121528f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_86 N_A2_c_62_n N_A_27_367#_c_233_n 0.0350175f $X=1.525 $Y=1.695 $X2=0 $Y2=0
cc_87 N_A2_c_63_n N_A_27_367#_c_233_n 0.00596721f $X=0.29 $Y=1.46 $X2=0 $Y2=0
cc_88 N_A2_M1010_g N_A_27_367#_c_236_n 0.0136928f $X=1.805 $Y=2.465 $X2=0 $Y2=0
cc_89 N_A2_c_62_n N_A_27_367#_c_236_n 0.0175636f $X=1.525 $Y=1.695 $X2=0 $Y2=0
cc_90 A2 N_A_27_367#_c_236_n 0.0219774f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_91 N_A2_c_66_n N_A_27_367#_c_236_n 4.82069e-19 $X=1.785 $Y=1.51 $X2=0 $Y2=0
cc_92 N_A2_c_66_n N_A_27_367#_c_240_n 0.00108953f $X=1.785 $Y=1.51 $X2=0 $Y2=0
cc_93 N_A2_c_62_n N_A_27_367#_c_241_n 0.0154593f $X=1.525 $Y=1.695 $X2=0 $Y2=0
cc_94 N_A2_M1009_g N_VPWR_c_269_n 0.0156794f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_95 N_A2_M1010_g N_VPWR_c_270_n 0.0132628f $X=1.805 $Y=2.465 $X2=0 $Y2=0
cc_96 N_A2_M1009_g N_VPWR_c_271_n 0.00486043f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_97 N_A2_M1010_g N_VPWR_c_273_n 0.00564095f $X=1.805 $Y=2.465 $X2=0 $Y2=0
cc_98 N_A2_M1009_g N_VPWR_c_268_n 0.00917987f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_99 N_A2_M1010_g N_VPWR_c_268_n 0.00950825f $X=1.805 $Y=2.465 $X2=0 $Y2=0
cc_100 N_A2_M1006_g N_Y_c_318_n 0.0157392f $X=1.765 $Y=0.655 $X2=0 $Y2=0
cc_101 N_A2_c_62_n N_Y_c_318_n 0.00410755f $X=1.525 $Y=1.695 $X2=0 $Y2=0
cc_102 A2 N_Y_c_318_n 0.0143846f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_103 N_A2_c_66_n N_Y_c_318_n 0.00248855f $X=1.785 $Y=1.51 $X2=0 $Y2=0
cc_104 N_A2_M1003_g N_VGND_c_362_n 0.00849399f $X=0.475 $Y=0.655 $X2=0 $Y2=0
cc_105 N_A2_c_63_n N_VGND_c_362_n 0.0175611f $X=0.29 $Y=1.46 $X2=0 $Y2=0
cc_106 N_A2_c_65_n N_VGND_c_362_n 0.00176788f $X=0.475 $Y=1.46 $X2=0 $Y2=0
cc_107 N_A2_M1006_g N_VGND_c_363_n 0.0100599f $X=1.765 $Y=0.655 $X2=0 $Y2=0
cc_108 N_A2_M1003_g N_VGND_c_365_n 0.00547432f $X=0.475 $Y=0.655 $X2=0 $Y2=0
cc_109 N_A2_M1006_g N_VGND_c_365_n 0.00564095f $X=1.765 $Y=0.655 $X2=0 $Y2=0
cc_110 N_A2_M1003_g N_VGND_c_370_n 0.0106866f $X=0.475 $Y=0.655 $X2=0 $Y2=0
cc_111 N_A2_M1006_g N_VGND_c_370_n 0.00961799f $X=1.765 $Y=0.655 $X2=0 $Y2=0
cc_112 N_A2_M1003_g N_A_110_47#_c_406_n 0.00843205f $X=0.475 $Y=0.655 $X2=0
+ $Y2=0
cc_113 N_A2_c_62_n N_A_110_47#_c_406_n 0.00221879f $X=1.525 $Y=1.695 $X2=0 $Y2=0
cc_114 N_A2_M1003_g N_A_110_47#_c_408_n 0.00202381f $X=0.475 $Y=0.655 $X2=0
+ $Y2=0
cc_115 N_A1_M1000_g N_A_27_367#_c_233_n 0.0122129f $X=0.905 $Y=2.465 $X2=0 $Y2=0
cc_116 N_A1_M1004_g N_A_27_367#_c_236_n 0.0129951f $X=1.335 $Y=2.465 $X2=0 $Y2=0
cc_117 N_A1_M1000_g N_VPWR_c_269_n 0.0138551f $X=0.905 $Y=2.465 $X2=0 $Y2=0
cc_118 N_A1_M1004_g N_VPWR_c_269_n 6.78754e-19 $X=1.335 $Y=2.465 $X2=0 $Y2=0
cc_119 N_A1_M1000_g N_VPWR_c_270_n 6.45189e-19 $X=0.905 $Y=2.465 $X2=0 $Y2=0
cc_120 N_A1_M1004_g N_VPWR_c_270_n 0.0121565f $X=1.335 $Y=2.465 $X2=0 $Y2=0
cc_121 N_A1_M1000_g N_VPWR_c_272_n 0.00486043f $X=0.905 $Y=2.465 $X2=0 $Y2=0
cc_122 N_A1_M1004_g N_VPWR_c_272_n 0.00564095f $X=1.335 $Y=2.465 $X2=0 $Y2=0
cc_123 N_A1_M1000_g N_VPWR_c_268_n 0.00824727f $X=0.905 $Y=2.465 $X2=0 $Y2=0
cc_124 N_A1_M1004_g N_VPWR_c_268_n 0.00948291f $X=1.335 $Y=2.465 $X2=0 $Y2=0
cc_125 N_A1_c_131_n N_Y_c_318_n 0.0105255f $X=1.335 $Y=1.185 $X2=0 $Y2=0
cc_126 A1 N_Y_c_318_n 0.00659228f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_127 A1 N_Y_c_324_n 0.0152957f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_128 N_A1_c_134_n N_Y_c_324_n 0.00235264f $X=1.335 $Y=1.35 $X2=0 $Y2=0
cc_129 N_A1_c_131_n N_VGND_c_363_n 0.0010882f $X=1.335 $Y=1.185 $X2=0 $Y2=0
cc_130 N_A1_c_129_n N_VGND_c_365_n 0.00357842f $X=0.905 $Y=1.185 $X2=0 $Y2=0
cc_131 N_A1_c_131_n N_VGND_c_365_n 0.00357877f $X=1.335 $Y=1.185 $X2=0 $Y2=0
cc_132 N_A1_c_129_n N_VGND_c_370_n 0.00537652f $X=0.905 $Y=1.185 $X2=0 $Y2=0
cc_133 N_A1_c_131_n N_VGND_c_370_n 0.00544922f $X=1.335 $Y=1.185 $X2=0 $Y2=0
cc_134 N_A1_c_129_n N_A_110_47#_c_406_n 0.00913566f $X=0.905 $Y=1.185 $X2=0
+ $Y2=0
cc_135 N_A1_c_131_n N_A_110_47#_c_406_n 5.20784e-19 $X=1.335 $Y=1.185 $X2=0
+ $Y2=0
cc_136 A1 N_A_110_47#_c_406_n 0.0165822f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_137 N_A1_c_129_n N_A_110_47#_c_412_n 0.010474f $X=0.905 $Y=1.185 $X2=0 $Y2=0
cc_138 N_A1_c_131_n N_A_110_47#_c_412_n 0.009382f $X=1.335 $Y=1.185 $X2=0 $Y2=0
cc_139 N_A1_c_129_n N_A_110_47#_c_408_n 5.89773e-19 $X=0.905 $Y=1.185 $X2=0
+ $Y2=0
cc_140 B1 N_A_27_367#_c_240_n 0.00540484f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_141 N_B1_M1001_g N_A_27_367#_c_229_n 0.0115031f $X=2.235 $Y=2.465 $X2=0 $Y2=0
cc_142 N_B1_M1005_g N_A_27_367#_c_229_n 0.0114565f $X=2.665 $Y=2.465 $X2=0 $Y2=0
cc_143 N_B1_M1001_g N_VPWR_c_270_n 0.00105138f $X=2.235 $Y=2.465 $X2=0 $Y2=0
cc_144 N_B1_M1001_g N_VPWR_c_273_n 0.00357877f $X=2.235 $Y=2.465 $X2=0 $Y2=0
cc_145 N_B1_M1005_g N_VPWR_c_273_n 0.00357877f $X=2.665 $Y=2.465 $X2=0 $Y2=0
cc_146 N_B1_M1001_g N_VPWR_c_268_n 0.00537654f $X=2.235 $Y=2.465 $X2=0 $Y2=0
cc_147 N_B1_M1005_g N_VPWR_c_268_n 0.00643596f $X=2.665 $Y=2.465 $X2=0 $Y2=0
cc_148 N_B1_M1002_g N_Y_c_318_n 0.0140845f $X=2.235 $Y=0.655 $X2=0 $Y2=0
cc_149 B1 N_Y_c_318_n 0.0100253f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_150 N_B1_M1008_g N_Y_c_313_n 0.0155045f $X=2.665 $Y=0.655 $X2=0 $Y2=0
cc_151 B1 N_Y_c_313_n 0.0140316f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_152 N_B1_M1005_g N_Y_c_316_n 0.0129759f $X=2.665 $Y=2.465 $X2=0 $Y2=0
cc_153 B1 N_Y_c_316_n 0.0115162f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_154 N_B1_M1001_g N_Y_c_332_n 0.0116173f $X=2.235 $Y=2.465 $X2=0 $Y2=0
cc_155 N_B1_M1005_g N_Y_c_332_n 0.0159266f $X=2.665 $Y=2.465 $X2=0 $Y2=0
cc_156 B1 N_Y_c_332_n 0.0230948f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_157 N_B1_c_181_n N_Y_c_332_n 6.37898e-19 $X=2.665 $Y=1.51 $X2=0 $Y2=0
cc_158 N_B1_M1002_g N_Y_c_314_n 0.00321539f $X=2.235 $Y=0.655 $X2=0 $Y2=0
cc_159 B1 N_Y_c_314_n 0.0126632f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_160 N_B1_c_181_n N_Y_c_314_n 0.00245863f $X=2.665 $Y=1.51 $X2=0 $Y2=0
cc_161 N_B1_M1008_g Y 0.00907351f $X=2.665 $Y=0.655 $X2=0 $Y2=0
cc_162 N_B1_M1005_g Y 0.0058705f $X=2.665 $Y=2.465 $X2=0 $Y2=0
cc_163 B1 Y 0.0292889f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_164 N_B1_c_181_n Y 0.00207593f $X=2.665 $Y=1.51 $X2=0 $Y2=0
cc_165 N_B1_M1002_g N_VGND_c_363_n 0.00894125f $X=2.235 $Y=0.655 $X2=0 $Y2=0
cc_166 N_B1_M1008_g N_VGND_c_363_n 5.54009e-19 $X=2.665 $Y=0.655 $X2=0 $Y2=0
cc_167 N_B1_M1002_g N_VGND_c_364_n 6.22172e-19 $X=2.235 $Y=0.655 $X2=0 $Y2=0
cc_168 N_B1_M1008_g N_VGND_c_364_n 0.0112869f $X=2.665 $Y=0.655 $X2=0 $Y2=0
cc_169 N_B1_M1002_g N_VGND_c_367_n 0.00564095f $X=2.235 $Y=0.655 $X2=0 $Y2=0
cc_170 N_B1_M1008_g N_VGND_c_367_n 0.00486043f $X=2.665 $Y=0.655 $X2=0 $Y2=0
cc_171 N_B1_M1002_g N_VGND_c_370_n 0.00948291f $X=2.235 $Y=0.655 $X2=0 $Y2=0
cc_172 N_B1_M1008_g N_VGND_c_370_n 0.00824727f $X=2.665 $Y=0.655 $X2=0 $Y2=0
cc_173 N_A_27_367#_c_233_n N_VPWR_M1009_s 0.00353353f $X=1.025 $Y=2.04 $X2=-0.19
+ $Y2=1.655
cc_174 N_A_27_367#_c_236_n N_VPWR_M1004_d 0.00427917f $X=1.905 $Y=2.04 $X2=0
+ $Y2=0
cc_175 N_A_27_367#_c_233_n N_VPWR_c_269_n 0.0170777f $X=1.025 $Y=2.04 $X2=0
+ $Y2=0
cc_176 N_A_27_367#_c_236_n N_VPWR_c_270_n 0.017285f $X=1.905 $Y=2.04 $X2=0 $Y2=0
cc_177 N_A_27_367#_c_228_n N_VPWR_c_271_n 0.0178111f $X=0.26 $Y=2.495 $X2=0
+ $Y2=0
cc_178 N_A_27_367#_c_252_p N_VPWR_c_272_n 0.0131621f $X=1.12 $Y=2.495 $X2=0
+ $Y2=0
cc_179 N_A_27_367#_c_253_p N_VPWR_c_273_n 0.0132331f $X=2.01 $Y=2.905 $X2=0
+ $Y2=0
cc_180 N_A_27_367#_c_229_n N_VPWR_c_273_n 0.0540354f $X=2.785 $Y=2.99 $X2=0
+ $Y2=0
cc_181 N_A_27_367#_M1009_d N_VPWR_c_268_n 0.00371702f $X=0.135 $Y=1.835 $X2=0
+ $Y2=0
cc_182 N_A_27_367#_M1000_s N_VPWR_c_268_n 0.00467071f $X=0.98 $Y=1.835 $X2=0
+ $Y2=0
cc_183 N_A_27_367#_M1010_d N_VPWR_c_268_n 0.00307052f $X=1.88 $Y=1.835 $X2=0
+ $Y2=0
cc_184 N_A_27_367#_M1005_d N_VPWR_c_268_n 0.00215161f $X=2.74 $Y=1.835 $X2=0
+ $Y2=0
cc_185 N_A_27_367#_c_228_n N_VPWR_c_268_n 0.0100304f $X=0.26 $Y=2.495 $X2=0
+ $Y2=0
cc_186 N_A_27_367#_c_252_p N_VPWR_c_268_n 0.00808656f $X=1.12 $Y=2.495 $X2=0
+ $Y2=0
cc_187 N_A_27_367#_c_253_p N_VPWR_c_268_n 0.00816431f $X=2.01 $Y=2.905 $X2=0
+ $Y2=0
cc_188 N_A_27_367#_c_229_n N_VPWR_c_268_n 0.0337842f $X=2.785 $Y=2.99 $X2=0
+ $Y2=0
cc_189 N_A_27_367#_c_229_n N_Y_M1001_s 0.00332344f $X=2.785 $Y=2.99 $X2=0 $Y2=0
cc_190 N_A_27_367#_M1005_d N_Y_c_316_n 0.00943791f $X=2.74 $Y=1.835 $X2=0 $Y2=0
cc_191 N_A_27_367#_c_230_n N_Y_c_316_n 0.0208033f $X=2.88 $Y=2.435 $X2=0 $Y2=0
cc_192 N_A_27_367#_c_229_n N_Y_c_332_n 0.0159805f $X=2.785 $Y=2.99 $X2=0 $Y2=0
cc_193 N_A_27_367#_M1005_d Y 0.00139965f $X=2.74 $Y=1.835 $X2=0 $Y2=0
cc_194 N_VPWR_c_268_n N_Y_M1001_s 0.00225186f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_195 N_Y_c_318_n N_VGND_M1006_s 0.00730886f $X=2.335 $Y=0.95 $X2=0 $Y2=0
cc_196 N_Y_c_313_n N_VGND_M1008_s 0.00253846f $X=2.97 $Y=1.09 $X2=0 $Y2=0
cc_197 N_Y_c_318_n N_VGND_c_363_n 0.017285f $X=2.335 $Y=0.95 $X2=0 $Y2=0
cc_198 N_Y_c_313_n N_VGND_c_364_n 0.0226345f $X=2.97 $Y=1.09 $X2=0 $Y2=0
cc_199 N_Y_c_353_p N_VGND_c_367_n 0.0131621f $X=2.45 $Y=0.42 $X2=0 $Y2=0
cc_200 N_Y_M1007_d N_VGND_c_370_n 0.00224381f $X=0.98 $Y=0.235 $X2=0 $Y2=0
cc_201 N_Y_M1002_d N_VGND_c_370_n 0.00467071f $X=2.31 $Y=0.235 $X2=0 $Y2=0
cc_202 N_Y_c_353_p N_VGND_c_370_n 0.00808656f $X=2.45 $Y=0.42 $X2=0 $Y2=0
cc_203 N_Y_c_318_n N_A_110_47#_M1011_s 0.00436932f $X=2.335 $Y=0.95 $X2=0 $Y2=0
cc_204 N_Y_M1007_d N_A_110_47#_c_412_n 0.00332344f $X=0.98 $Y=0.235 $X2=0 $Y2=0
cc_205 N_Y_c_318_n N_A_110_47#_c_412_n 0.0177178f $X=2.335 $Y=0.95 $X2=0 $Y2=0
cc_206 N_Y_c_324_n N_A_110_47#_c_412_n 0.0122234f $X=1.12 $Y=0.76 $X2=0 $Y2=0
cc_207 N_VGND_c_370_n N_A_110_47#_M1003_d 0.00223559f $X=3.12 $Y=0 $X2=-0.19
+ $Y2=-0.245
cc_208 N_VGND_c_370_n N_A_110_47#_M1011_s 0.00314812f $X=3.12 $Y=0 $X2=0 $Y2=0
cc_209 N_VGND_c_365_n N_A_110_47#_c_412_n 0.0458243f $X=1.835 $Y=0 $X2=0 $Y2=0
cc_210 N_VGND_c_370_n N_A_110_47#_c_412_n 0.0293225f $X=3.12 $Y=0 $X2=0 $Y2=0
cc_211 N_VGND_c_365_n N_A_110_47#_c_408_n 0.01906f $X=1.835 $Y=0 $X2=0 $Y2=0
cc_212 N_VGND_c_370_n N_A_110_47#_c_408_n 0.0124545f $X=3.12 $Y=0 $X2=0 $Y2=0
