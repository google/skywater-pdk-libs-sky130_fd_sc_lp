* File: sky130_fd_sc_lp__a32o_1.spice
* Created: Wed Sep  2 09:27:34 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__a32o_1.pex.spice"
.subckt sky130_fd_sc_lp__a32o_1  VNB VPB A3 A2 A1 B1 B2 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* B2	B2
* B1	B1
* A1	A1
* A2	A2
* A3	A3
* VPB	VPB
* VNB	VNB
MM1006 N_VGND_M1006_d N_A_80_21#_M1006_g N_X_M1006_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2583 AS=0.2226 PD=1.455 PS=2.21 NRD=23.928 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75003 A=0.126 P=1.98 MULT=1
MM1002 A_263_47# N_A3_M1002_g N_VGND_M1006_d VNB NSHORT L=0.15 W=0.84 AD=0.1323
+ AS=0.2583 PD=1.155 PS=1.455 NRD=14.64 NRS=23.928 M=1 R=5.6 SA=75001 SB=75002.3
+ A=0.126 P=1.98 MULT=1
MM1007 A_356_47# N_A2_M1007_g A_263_47# VNB NSHORT L=0.15 W=0.84 AD=0.1407
+ AS=0.1323 PD=1.175 PS=1.155 NRD=16.068 NRS=14.64 M=1 R=5.6 SA=75001.4
+ SB=75001.8 A=0.126 P=1.98 MULT=1
MM1004 N_A_80_21#_M1004_d N_A1_M1004_g A_356_47# VNB NSHORT L=0.15 W=0.84
+ AD=0.2646 AS=0.1407 PD=1.47 PS=1.175 NRD=0 NRS=16.068 M=1 R=5.6 SA=75001.9
+ SB=75001.3 A=0.126 P=1.98 MULT=1
MM1001 A_609_47# N_B1_M1001_g N_A_80_21#_M1004_d VNB NSHORT L=0.15 W=0.84
+ AD=0.0882 AS=0.2646 PD=1.05 PS=1.47 NRD=7.14 NRS=0 M=1 R=5.6 SA=75002.7
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1010 N_VGND_M1010_d N_B2_M1010_g A_609_47# VNB NSHORT L=0.15 W=0.84 AD=0.2226
+ AS=0.0882 PD=2.21 PS=1.05 NRD=0 NRS=7.14 M=1 R=5.6 SA=75003 SB=75000.2 A=0.126
+ P=1.98 MULT=1
MM1005 N_VPWR_M1005_d N_A_80_21#_M1005_g N_X_M1005_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.22365 AS=0.3339 PD=1.615 PS=3.05 NRD=0.7683 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75002.9 A=0.189 P=2.82 MULT=1
MM1008 N_A_249_367#_M1008_d N_A3_M1008_g N_VPWR_M1005_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.22365 PD=1.54 PS=1.615 NRD=0 NRS=10.9335 M=1 R=8.4
+ SA=75000.7 SB=75002.4 A=0.189 P=2.82 MULT=1
MM1000 N_VPWR_M1000_d N_A2_M1000_g N_A_249_367#_M1008_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.4284 AS=0.1764 PD=1.94 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75001.9 A=0.189 P=2.82 MULT=1
MM1009 N_A_249_367#_M1009_d N_A1_M1009_g N_VPWR_M1000_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.4284 PD=1.54 PS=1.94 NRD=0 NRS=0 M=1 R=8.4 SA=75002
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1003 N_A_80_21#_M1003_d N_B1_M1003_g N_A_249_367#_M1009_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.2016 AS=0.1764 PD=1.58 PS=1.54 NRD=1.5563 NRS=0 M=1 R=8.4
+ SA=75002.4 SB=75000.7 A=0.189 P=2.82 MULT=1
MM1011 N_A_249_367#_M1011_d N_B2_M1011_g N_A_80_21#_M1003_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.2016 PD=3.05 PS=1.58 NRD=0 NRS=4.6886 M=1 R=8.4
+ SA=75002.9 SB=75000.2 A=0.189 P=2.82 MULT=1
DX12_noxref VNB VPB NWDIODE A=7.8703 P=12.17
*
.include "sky130_fd_sc_lp__a32o_1.pxi.spice"
*
.ends
*
*
