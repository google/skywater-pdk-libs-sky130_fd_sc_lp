* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__ebufn_lp2 A TE_B VGND VNB VPB VPWR Z
X0 a_114_47# A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 a_27_47# A a_114_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 Z a_27_47# a_475_419# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X3 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X4 a_475_419# TE_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X5 VGND TE_B a_606_153# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 Z a_27_47# a_425_193# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 a_606_153# TE_B a_232_231# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 a_425_193# a_232_231# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 VPWR TE_B a_232_231# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
.ends
