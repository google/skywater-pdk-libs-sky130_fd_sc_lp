* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__o32ai_lp A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
M1000 Y B2 a_134_419# VPB phighvt w=1e+06u l=250000u
+  ad=2.8e+11p pd=2.56e+06u as=2.4e+11p ps=2.48e+06u
M1001 VPWR A1 a_463_419# VPB phighvt w=1e+06u l=250000u
+  ad=5.7e+11p pd=5.14e+06u as=3.2e+11p ps=2.64e+06u
M1002 a_338_419# A3 Y VPB phighvt w=1e+06u l=250000u
+  ad=3.75e+11p pd=2.75e+06u as=0p ps=0u
M1003 a_27_179# B2 Y VNB nshort w=420000u l=150000u
+  ad=4.934e+11p pd=4.95e+06u as=1.176e+11p ps=1.4e+06u
M1004 a_463_419# A2 a_338_419# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VGND A3 a_27_179# VNB nshort w=420000u l=150000u
+  ad=4.095e+11p pd=3.63e+06u as=0p ps=0u
M1006 a_27_179# A2 VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND A1 a_27_179# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_134_419# B1 VPWR VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1009 Y B1 a_27_179# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
