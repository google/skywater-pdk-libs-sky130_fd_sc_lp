* NGSPICE file created from sky130_fd_sc_lp__inv_m.ext - technology: sky130A

.subckt sky130_fd_sc_lp__inv_m A VGND VNB VPB VPWR Y
M1000 Y A VGND VNB nshort w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=1.113e+11p ps=1.37e+06u
M1001 Y A VPWR VPB phighvt w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=1.113e+11p ps=1.37e+06u
.ends

