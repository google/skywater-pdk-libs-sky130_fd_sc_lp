* File: sky130_fd_sc_lp__mux4_lp.pxi.spice
* Created: Fri Aug 28 10:46:30 2020
* 
x_PM_SKY130_FD_SC_LP__MUX4_LP%A_84_21# N_A_84_21#_M1016_d N_A_84_21#_M1013_d
+ N_A_84_21#_M1006_g N_A_84_21#_M1005_g N_A_84_21#_c_207_n N_A_84_21#_c_208_n
+ N_A_84_21#_M1026_g N_A_84_21#_c_209_n N_A_84_21#_c_210_n N_A_84_21#_c_211_n
+ N_A_84_21#_c_212_n N_A_84_21#_c_213_n N_A_84_21#_c_214_n
+ PM_SKY130_FD_SC_LP__MUX4_LP%A_84_21#
x_PM_SKY130_FD_SC_LP__MUX4_LP%S1 N_S1_c_285_n N_S1_c_286_n N_S1_c_287_n
+ N_S1_M1016_g N_S1_c_301_n N_S1_M1001_g N_S1_c_288_n N_S1_c_289_n N_S1_c_290_n
+ N_S1_M1017_g N_S1_c_291_n N_S1_c_292_n N_S1_c_293_n N_S1_M1022_g N_S1_c_295_n
+ N_S1_M1007_g N_S1_c_296_n N_S1_c_297_n N_S1_c_298_n N_S1_c_307_n N_S1_c_325_n
+ N_S1_c_335_p N_S1_c_308_n S1 N_S1_c_300_n PM_SKY130_FD_SC_LP__MUX4_LP%S1
x_PM_SKY130_FD_SC_LP__MUX4_LP%A_320_366# N_A_320_366#_M1017_s
+ N_A_320_366#_M1022_s N_A_320_366#_c_442_n N_A_320_366#_M1013_g
+ N_A_320_366#_c_435_n N_A_320_366#_M1025_g N_A_320_366#_c_444_n
+ N_A_320_366#_c_437_n N_A_320_366#_c_438_n N_A_320_366#_c_439_n
+ N_A_320_366#_c_440_n N_A_320_366#_c_446_n N_A_320_366#_c_441_n
+ PM_SKY130_FD_SC_LP__MUX4_LP%A_320_366#
x_PM_SKY130_FD_SC_LP__MUX4_LP%A3 N_A3_M1002_g N_A3_c_522_n N_A3_c_523_n
+ N_A3_M1027_g N_A3_c_524_n A3 A3 N_A3_c_526_n PM_SKY130_FD_SC_LP__MUX4_LP%A3
x_PM_SKY130_FD_SC_LP__MUX4_LP%S0 N_S0_M1003_g N_S0_M1008_g N_S0_M1019_g
+ N_S0_M1004_g N_S0_c_570_n N_S0_M1014_g N_S0_M1028_g N_S0_c_571_n N_S0_M1020_g
+ N_S0_c_572_n N_S0_c_573_n N_S0_c_574_n N_S0_c_575_n N_S0_c_576_n N_S0_c_577_n
+ N_S0_c_578_n N_S0_c_579_n N_S0_c_580_n N_S0_c_614_p N_S0_c_615_p N_S0_c_616_p
+ N_S0_c_596_n N_S0_c_651_p N_S0_c_581_n N_S0_c_582_n N_S0_c_583_n N_S0_c_584_n
+ N_S0_c_585_n S0 S0 S0 N_S0_c_586_n N_S0_c_587_n N_S0_c_588_n N_S0_c_589_n
+ N_S0_c_590_n S0 PM_SKY130_FD_SC_LP__MUX4_LP%S0
x_PM_SKY130_FD_SC_LP__MUX4_LP%A_946_317# N_A_946_317#_M1020_d
+ N_A_946_317#_M1028_d N_A_946_317#_M1015_g N_A_946_317#_c_779_n
+ N_A_946_317#_M1011_g N_A_946_317#_M1023_g N_A_946_317#_c_781_n
+ N_A_946_317#_c_782_n N_A_946_317#_c_783_n N_A_946_317#_c_784_n
+ N_A_946_317#_M1024_g N_A_946_317#_c_785_n N_A_946_317#_c_799_n
+ N_A_946_317#_c_800_n N_A_946_317#_c_841_n N_A_946_317#_c_843_n
+ N_A_946_317#_c_894_p N_A_946_317#_c_786_n N_A_946_317#_c_850_n
+ N_A_946_317#_c_854_n N_A_946_317#_c_856_n N_A_946_317#_c_787_n
+ N_A_946_317#_c_788_n N_A_946_317#_c_789_n N_A_946_317#_c_803_n
+ N_A_946_317#_c_790_n N_A_946_317#_c_791_n N_A_946_317#_c_804_n
+ N_A_946_317#_c_792_n N_A_946_317#_c_793_n
+ PM_SKY130_FD_SC_LP__MUX4_LP%A_946_317#
x_PM_SKY130_FD_SC_LP__MUX4_LP%A2 N_A2_M1012_g N_A2_c_972_n N_A2_c_973_n
+ N_A2_M1009_g N_A2_c_974_n A2 N_A2_c_976_n N_A2_c_977_n
+ PM_SKY130_FD_SC_LP__MUX4_LP%A2
x_PM_SKY130_FD_SC_LP__MUX4_LP%A1 N_A1_c_1026_n N_A1_M1010_g N_A1_M1018_g
+ N_A1_c_1028_n A1 N_A1_c_1030_n PM_SKY130_FD_SC_LP__MUX4_LP%A1
x_PM_SKY130_FD_SC_LP__MUX4_LP%A0 N_A0_M1000_g N_A0_M1021_g A0 A0 A0
+ N_A0_c_1072_n PM_SKY130_FD_SC_LP__MUX4_LP%A0
x_PM_SKY130_FD_SC_LP__MUX4_LP%X N_X_M1006_s N_X_M1005_s X X X X X X X
+ PM_SKY130_FD_SC_LP__MUX4_LP%X
x_PM_SKY130_FD_SC_LP__MUX4_LP%VPWR N_VPWR_M1005_d N_VPWR_M1022_d N_VPWR_M1009_d
+ N_VPWR_M1021_d N_VPWR_c_1127_n N_VPWR_c_1128_n N_VPWR_c_1129_n N_VPWR_c_1130_n
+ N_VPWR_c_1131_n N_VPWR_c_1132_n N_VPWR_c_1133_n N_VPWR_c_1134_n VPWR
+ N_VPWR_c_1135_n N_VPWR_c_1136_n N_VPWR_c_1126_n N_VPWR_c_1138_n
+ N_VPWR_c_1139_n PM_SKY130_FD_SC_LP__MUX4_LP%VPWR
x_PM_SKY130_FD_SC_LP__MUX4_LP%A_245_411# N_A_245_411#_M1016_s
+ N_A_245_411#_M1003_d N_A_245_411#_M1013_s N_A_245_411#_M1015_d
+ N_A_245_411#_c_1224_n N_A_245_411#_c_1225_n N_A_245_411#_c_1226_n
+ N_A_245_411#_c_1231_n N_A_245_411#_c_1253_n N_A_245_411#_c_1232_n
+ N_A_245_411#_c_1233_n N_A_245_411#_c_1234_n N_A_245_411#_c_1227_n
+ N_A_245_411#_c_1235_n N_A_245_411#_c_1276_n N_A_245_411#_c_1236_n
+ N_A_245_411#_c_1228_n N_A_245_411#_c_1291_n N_A_245_411#_c_1229_n
+ N_A_245_411#_c_1306_n N_A_245_411#_c_1238_n N_A_245_411#_c_1336_n
+ N_A_245_411#_c_1292_n PM_SKY130_FD_SC_LP__MUX4_LP%A_245_411#
x_PM_SKY130_FD_SC_LP__MUX4_LP%A_470_57# N_A_470_57#_M1025_d N_A_470_57#_M1019_d
+ N_A_470_57#_M1001_d N_A_470_57#_M1023_d N_A_470_57#_c_1370_n
+ N_A_470_57#_c_1385_n N_A_470_57#_c_1386_n N_A_470_57#_c_1387_n
+ N_A_470_57#_c_1371_n N_A_470_57#_c_1372_n N_A_470_57#_c_1373_n
+ N_A_470_57#_c_1374_n N_A_470_57#_c_1375_n N_A_470_57#_c_1376_n
+ N_A_470_57#_c_1377_n N_A_470_57#_c_1378_n N_A_470_57#_c_1379_n
+ N_A_470_57#_c_1380_n N_A_470_57#_c_1381_n N_A_470_57#_c_1382_n
+ N_A_470_57#_c_1383_n N_A_470_57#_c_1384_n
+ PM_SKY130_FD_SC_LP__MUX4_LP%A_470_57#
x_PM_SKY130_FD_SC_LP__MUX4_LP%VGND N_VGND_M1026_d N_VGND_M1007_d N_VGND_M1012_d
+ N_VGND_M1000_d N_VGND_c_1550_n N_VGND_c_1551_n N_VGND_c_1552_n N_VGND_c_1553_n
+ N_VGND_c_1554_n N_VGND_c_1555_n N_VGND_c_1556_n N_VGND_c_1557_n VGND
+ N_VGND_c_1558_n N_VGND_c_1559_n N_VGND_c_1560_n N_VGND_c_1561_n
+ N_VGND_c_1562_n N_VGND_c_1563_n PM_SKY130_FD_SC_LP__MUX4_LP%VGND
cc_1 VNB N_A_84_21#_M1006_g 0.0411935f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.445
cc_2 VNB N_A_84_21#_M1005_g 0.0307035f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=2.545
cc_3 VNB N_A_84_21#_c_207_n 0.0221231f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=1.185
cc_4 VNB N_A_84_21#_c_208_n 0.0160229f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=0.73
cc_5 VNB N_A_84_21#_c_209_n 0.00854607f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=1.185
cc_6 VNB N_A_84_21#_c_210_n 0.0105137f $X=-0.19 $Y=-0.245 $X2=1.975 $Y2=1.127
cc_7 VNB N_A_84_21#_c_211_n 0.052709f $X=-0.19 $Y=-0.245 $X2=1.14 $Y2=1.095
cc_8 VNB N_A_84_21#_c_212_n 0.00826795f $X=-0.19 $Y=-0.245 $X2=2.06 $Y2=0.495
cc_9 VNB N_A_84_21#_c_213_n 0.00862991f $X=-0.19 $Y=-0.245 $X2=2.07 $Y2=2.2
cc_10 VNB N_A_84_21#_c_214_n 0.00145736f $X=-0.19 $Y=-0.245 $X2=2.065 $Y2=1.127
cc_11 VNB N_S1_c_285_n 0.0189834f $X=-0.19 $Y=-0.245 $X2=1.92 $Y2=0.285
cc_12 VNB N_S1_c_286_n 0.0323947f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_S1_c_287_n 0.0177199f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_S1_c_288_n 0.00897638f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=1.26
cc_15 VNB N_S1_c_289_n 0.0188308f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=2.545
cc_16 VNB N_S1_c_290_n 0.015f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=2.545
cc_17 VNB N_S1_c_291_n 0.0156167f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=0.73
cc_18 VNB N_S1_c_292_n 0.0156867f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=0.445
cc_19 VNB N_S1_c_293_n 0.0142553f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=1.185
cc_20 VNB N_S1_M1022_g 0.0017411f $X=-0.19 $Y=-0.245 $X2=1.14 $Y2=1.127
cc_21 VNB N_S1_c_295_n 0.0153824f $X=-0.19 $Y=-0.245 $X2=1.14 $Y2=1.095
cc_22 VNB N_S1_c_296_n 0.02413f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_S1_c_297_n 0.00669963f $X=-0.19 $Y=-0.245 $X2=2.07 $Y2=2.2
cc_24 VNB N_S1_c_298_n 0.00340752f $X=-0.19 $Y=-0.245 $X2=1.042 $Y2=1.095
cc_25 VNB S1 0.00394494f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_S1_c_300_n 0.0161613f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_320_366#_c_435_n 0.0198286f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=1.26
cc_28 VNB N_A_320_366#_M1025_g 0.0321106f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_320_366#_c_437_n 0.00586716f $X=-0.19 $Y=-0.245 $X2=0.545
+ $Y2=1.185
cc_30 VNB N_A_320_366#_c_438_n 0.00621783f $X=-0.19 $Y=-0.245 $X2=2.06 $Y2=0.495
cc_31 VNB N_A_320_366#_c_439_n 0.00541714f $X=-0.19 $Y=-0.245 $X2=2.07 $Y2=1.26
cc_32 VNB N_A_320_366#_c_440_n 0.00720808f $X=-0.19 $Y=-0.245 $X2=2.07 $Y2=2.2
cc_33 VNB N_A_320_366#_c_441_n 0.06934f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A3_c_522_n 0.0264063f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A3_c_523_n 0.0164498f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.11
cc_36 VNB N_A3_c_524_n 0.0155512f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=2.545
cc_37 VNB A3 0.0047459f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A3_c_526_n 0.0175878f $X=-0.19 $Y=-0.245 $X2=1.14 $Y2=1.095
cc_39 VNB N_S0_M1019_g 0.0328162f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_S0_c_570_n 0.0135932f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.185
cc_41 VNB N_S0_c_571_n 0.0172354f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_S0_c_572_n 0.0265258f $X=-0.19 $Y=-0.245 $X2=2.07 $Y2=2.2
cc_43 VNB N_S0_c_573_n 0.0319973f $X=-0.19 $Y=-0.245 $X2=1.042 $Y2=1.185
cc_44 VNB N_S0_c_574_n 0.0107984f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_S0_c_575_n 0.00481757f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_S0_c_576_n 6.35056e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_S0_c_577_n 0.0162332f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_S0_c_578_n 2.87724e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_S0_c_579_n 0.00475759f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_S0_c_580_n 0.0334674f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_S0_c_581_n 0.00365003f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_S0_c_582_n 0.010833f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_S0_c_583_n 0.00294166f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_S0_c_584_n 0.0211165f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_S0_c_585_n 3.82079e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_S0_c_586_n 0.0181899f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_S0_c_587_n 0.0121582f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_S0_c_588_n 0.00968476f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_S0_c_589_n 0.00492178f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_S0_c_590_n 0.0447233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_A_946_317#_c_779_n 0.00822316f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=1.26
cc_62 VNB N_A_946_317#_M1011_g 0.0674944f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=1.185
cc_63 VNB N_A_946_317#_c_781_n 0.00740892f $X=-0.19 $Y=-0.245 $X2=1.975
+ $Y2=1.127
cc_64 VNB N_A_946_317#_c_782_n 0.00505016f $X=-0.19 $Y=-0.245 $X2=1.14 $Y2=1.127
cc_65 VNB N_A_946_317#_c_783_n 0.0379595f $X=-0.19 $Y=-0.245 $X2=1.14 $Y2=1.095
cc_66 VNB N_A_946_317#_c_784_n 0.0198709f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_A_946_317#_c_785_n 0.0136767f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_A_946_317#_c_786_n 0.0149807f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_946_317#_c_787_n 0.0236757f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_A_946_317#_c_788_n 0.0312005f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_A_946_317#_c_789_n 0.00221406f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_A_946_317#_c_790_n 0.0537963f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_A_946_317#_c_791_n 0.0010407f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_A_946_317#_c_792_n 0.0144611f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_A_946_317#_c_793_n 0.0164761f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_A2_c_972_n 0.0259223f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_A2_c_973_n 0.0031101f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.445
cc_78 VNB N_A2_c_974_n 0.0345801f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=2.545
cc_79 VNB A2 0.00308413f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=2.545
cc_80 VNB N_A2_c_976_n 0.0324613f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.185
cc_81 VNB N_A2_c_977_n 0.0194783f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=0.445
cc_82 VNB N_A1_c_1026_n 0.00303211f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_A1_M1018_g 0.0386106f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.445
cc_84 VNB N_A1_c_1028_n 0.014806f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=1.26
cc_85 VNB A1 0.00528493f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=2.545
cc_86 VNB N_A1_c_1030_n 0.0273411f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=1.185
cc_87 VNB N_A0_M1000_g 0.0422819f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_A0_M1021_g 0.0130205f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.11
cc_89 VNB A0 0.0188187f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=1.26
cc_90 VNB N_A0_c_1072_n 0.033684f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.185
cc_91 VNB X 0.0568045f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.11
cc_92 VNB N_VPWR_c_1126_n 0.422413f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_93 VNB N_A_245_411#_c_1224_n 0.0145754f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_94 VNB N_A_245_411#_c_1225_n 0.00645764f $X=-0.19 $Y=-0.245 $X2=0.975
+ $Y2=1.185
cc_95 VNB N_A_245_411#_c_1226_n 9.57196e-19 $X=-0.19 $Y=-0.245 $X2=0.67
+ $Y2=1.185
cc_96 VNB N_A_245_411#_c_1227_n 0.00675634f $X=-0.19 $Y=-0.245 $X2=2.06
+ $Y2=0.495
cc_97 VNB N_A_245_411#_c_1228_n 0.0165971f $X=-0.19 $Y=-0.245 $X2=2.065
+ $Y2=1.127
cc_98 VNB N_A_245_411#_c_1229_n 0.00231163f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_99 VNB N_A_470_57#_c_1370_n 0.0195704f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=2.545
cc_100 VNB N_A_470_57#_c_1371_n 9.89651e-19 $X=-0.19 $Y=-0.245 $X2=1.14
+ $Y2=1.127
cc_101 VNB N_A_470_57#_c_1372_n 0.00410658f $X=-0.19 $Y=-0.245 $X2=1.14
+ $Y2=1.095
cc_102 VNB N_A_470_57#_c_1373_n 0.0184279f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_103 VNB N_A_470_57#_c_1374_n 0.00199632f $X=-0.19 $Y=-0.245 $X2=2.06
+ $Y2=0.995
cc_104 VNB N_A_470_57#_c_1375_n 0.00361572f $X=-0.19 $Y=-0.245 $X2=2.06
+ $Y2=0.495
cc_105 VNB N_A_470_57#_c_1376_n 0.0105964f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_106 VNB N_A_470_57#_c_1377_n 0.00311572f $X=-0.19 $Y=-0.245 $X2=2.07 $Y2=1.26
cc_107 VNB N_A_470_57#_c_1378_n 0.00219628f $X=-0.19 $Y=-0.245 $X2=2.07 $Y2=2.2
cc_108 VNB N_A_470_57#_c_1379_n 0.0295711f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_109 VNB N_A_470_57#_c_1380_n 0.00367292f $X=-0.19 $Y=-0.245 $X2=2.065
+ $Y2=1.127
cc_110 VNB N_A_470_57#_c_1381_n 8.39137e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_111 VNB N_A_470_57#_c_1382_n 0.00623451f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_112 VNB N_A_470_57#_c_1383_n 0.00913583f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_113 VNB N_A_470_57#_c_1384_n 0.00774356f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_114 VNB N_VGND_c_1550_n 0.00519098f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=1.185
cc_115 VNB N_VGND_c_1551_n 0.0123039f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=0.445
cc_116 VNB N_VGND_c_1552_n 0.00518129f $X=-0.19 $Y=-0.245 $X2=1.14 $Y2=1.095
cc_117 VNB N_VGND_c_1553_n 0.00280619f $X=-0.19 $Y=-0.245 $X2=2.06 $Y2=0.495
cc_118 VNB N_VGND_c_1554_n 0.0631208f $X=-0.19 $Y=-0.245 $X2=2.07 $Y2=1.26
cc_119 VNB N_VGND_c_1555_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=2.07 $Y2=2.2
cc_120 VNB N_VGND_c_1556_n 0.0616104f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_121 VNB N_VGND_c_1557_n 0.00478105f $X=-0.19 $Y=-0.245 $X2=2.065 $Y2=1.127
cc_122 VNB N_VGND_c_1558_n 0.0256527f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_123 VNB N_VGND_c_1559_n 0.0555781f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_124 VNB N_VGND_c_1560_n 0.0268233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_125 VNB N_VGND_c_1561_n 0.511585f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_126 VNB N_VGND_c_1562_n 0.00510127f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_127 VNB N_VGND_c_1563_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_128 VPB N_A_84_21#_M1005_g 0.0508236f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=2.545
cc_129 VPB N_A_84_21#_c_213_n 0.00296293f $X=-0.19 $Y=1.655 $X2=2.07 $Y2=2.2
cc_130 VPB N_S1_c_301_n 0.0232596f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=0.445
cc_131 VPB N_S1_c_288_n 0.00927962f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=1.26
cc_132 VPB N_S1_c_289_n 0.056526f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=2.545
cc_133 VPB N_S1_c_293_n 0.0119211f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=1.185
cc_134 VPB N_S1_M1022_g 0.0547147f $X=-0.19 $Y=1.655 $X2=1.14 $Y2=1.127
cc_135 VPB N_S1_c_298_n 0.00861531f $X=-0.19 $Y=1.655 $X2=1.042 $Y2=1.095
cc_136 VPB N_S1_c_307_n 0.00117059f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_137 VPB N_S1_c_308_n 2.10075e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_138 VPB S1 0.00371825f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_139 VPB N_S1_c_300_n 0.0185764f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_140 VPB N_A_320_366#_c_442_n 0.0244856f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=1.11
cc_141 VPB N_A_320_366#_c_435_n 0.0100704f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=1.26
cc_142 VPB N_A_320_366#_c_444_n 0.0331632f $X=-0.19 $Y=1.655 $X2=0.855 $Y2=0.445
cc_143 VPB N_A_320_366#_c_439_n 0.00133644f $X=-0.19 $Y=1.655 $X2=2.07 $Y2=1.26
cc_144 VPB N_A_320_366#_c_446_n 0.00755464f $X=-0.19 $Y=1.655 $X2=1.042
+ $Y2=1.095
cc_145 VPB N_A3_M1002_g 0.0294588f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_146 VPB A3 0.00292819f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_147 VPB N_A3_c_526_n 0.0239275f $X=-0.19 $Y=1.655 $X2=1.14 $Y2=1.095
cc_148 VPB N_S0_M1008_g 0.0422461f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_149 VPB N_S0_M1004_g 0.026445f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_150 VPB N_S0_M1028_g 0.028845f $X=-0.19 $Y=1.655 $X2=1.14 $Y2=1.095
cc_151 VPB N_S0_c_577_n 0.00444402f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_152 VPB N_S0_c_578_n 7.50383e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_153 VPB N_S0_c_596_n 0.00335728f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_154 VPB N_S0_c_583_n 8.94876e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_155 VPB N_S0_c_584_n 0.0104043f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_156 VPB N_S0_c_585_n 0.00505021f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_157 VPB N_S0_c_587_n 0.0196171f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_158 VPB N_S0_c_588_n 0.0239444f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_159 VPB N_S0_c_589_n 0.00421325f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_160 VPB N_A_946_317#_M1015_g 0.0310702f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=0.445
cc_161 VPB N_A_946_317#_c_779_n 0.0121535f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=1.26
cc_162 VPB N_A_946_317#_M1023_g 0.0373428f $X=-0.19 $Y=1.655 $X2=0.855 $Y2=0.445
cc_163 VPB N_A_946_317#_c_781_n 0.0189938f $X=-0.19 $Y=1.655 $X2=1.975 $Y2=1.127
cc_164 VPB N_A_946_317#_c_782_n 0.00579409f $X=-0.19 $Y=1.655 $X2=1.14 $Y2=1.127
cc_165 VPB N_A_946_317#_c_799_n 0.00949946f $X=-0.19 $Y=1.655 $X2=2.07 $Y2=1.26
cc_166 VPB N_A_946_317#_c_800_n 0.0106346f $X=-0.19 $Y=1.655 $X2=2.07 $Y2=2.2
cc_167 VPB N_A_946_317#_c_788_n 0.0301851f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_168 VPB N_A_946_317#_c_789_n 0.00220869f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_169 VPB N_A_946_317#_c_803_n 0.00825803f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_170 VPB N_A_946_317#_c_804_n 0.0337683f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_171 VPB N_A_946_317#_c_793_n 0.0287572f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_172 VPB N_A2_c_973_n 0.00639951f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=0.445
cc_173 VPB N_A2_M1009_g 0.0352016f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_174 VPB N_A1_c_1026_n 0.00649733f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_175 VPB N_A1_M1010_g 0.0342362f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_176 VPB N_A0_M1021_g 0.038581f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=1.11
cc_177 VPB X 0.0573842f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=1.11
cc_178 VPB N_VPWR_c_1127_n 0.0110533f $X=-0.19 $Y=1.655 $X2=0.855 $Y2=0.73
cc_179 VPB N_VPWR_c_1128_n 0.00475965f $X=-0.19 $Y=1.655 $X2=1.975 $Y2=1.127
cc_180 VPB N_VPWR_c_1129_n 0.00283116f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_181 VPB N_VPWR_c_1130_n 4.89148e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_182 VPB N_VPWR_c_1131_n 0.0686967f $X=-0.19 $Y=1.655 $X2=2.07 $Y2=2.2
cc_183 VPB N_VPWR_c_1132_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_184 VPB N_VPWR_c_1133_n 0.0490717f $X=-0.19 $Y=1.655 $X2=1.042 $Y2=1.095
cc_185 VPB N_VPWR_c_1134_n 0.00436868f $X=-0.19 $Y=1.655 $X2=1.042 $Y2=1.185
cc_186 VPB N_VPWR_c_1135_n 0.069946f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_187 VPB N_VPWR_c_1136_n 0.0212611f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_188 VPB N_VPWR_c_1126_n 0.0720697f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_189 VPB N_VPWR_c_1138_n 0.0244124f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_190 VPB N_VPWR_c_1139_n 0.00631443f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_191 VPB N_A_245_411#_c_1224_n 0.00717313f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_192 VPB N_A_245_411#_c_1231_n 0.0218391f $X=-0.19 $Y=1.655 $X2=0.855 $Y2=0.73
cc_193 VPB N_A_245_411#_c_1232_n 0.00345005f $X=-0.19 $Y=1.655 $X2=0.545
+ $Y2=1.185
cc_194 VPB N_A_245_411#_c_1233_n 0.00757689f $X=-0.19 $Y=1.655 $X2=1.14
+ $Y2=1.127
cc_195 VPB N_A_245_411#_c_1234_n 0.0135978f $X=-0.19 $Y=1.655 $X2=1.14 $Y2=1.095
cc_196 VPB N_A_245_411#_c_1235_n 0.00312609f $X=-0.19 $Y=1.655 $X2=2.07 $Y2=1.26
cc_197 VPB N_A_245_411#_c_1236_n 0.0023998f $X=-0.19 $Y=1.655 $X2=2.07 $Y2=2.2
cc_198 VPB N_A_245_411#_c_1228_n 0.00847022f $X=-0.19 $Y=1.655 $X2=2.065
+ $Y2=1.127
cc_199 VPB N_A_245_411#_c_1238_n 0.00158626f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_200 VPB N_A_470_57#_c_1385_n 0.00461654f $X=-0.19 $Y=1.655 $X2=0.855 $Y2=0.73
cc_201 VPB N_A_470_57#_c_1386_n 0.00735968f $X=-0.19 $Y=1.655 $X2=0.855
+ $Y2=0.445
cc_202 VPB N_A_470_57#_c_1387_n 3.95783e-19 $X=-0.19 $Y=1.655 $X2=0.545
+ $Y2=1.185
cc_203 VPB N_A_470_57#_c_1382_n 0.00371478f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_204 N_A_84_21#_c_210_n N_S1_c_286_n 0.0146095f $X=1.975 $Y=1.127 $X2=0 $Y2=0
cc_205 N_A_84_21#_c_211_n N_S1_c_286_n 0.018572f $X=1.14 $Y=1.095 $X2=0 $Y2=0
cc_206 N_A_84_21#_c_212_n N_S1_c_286_n 0.00127618f $X=2.06 $Y=0.495 $X2=0 $Y2=0
cc_207 N_A_84_21#_c_213_n N_S1_c_286_n 0.00121768f $X=2.07 $Y=2.2 $X2=0 $Y2=0
cc_208 N_A_84_21#_c_211_n N_S1_c_287_n 5.77446e-19 $X=1.14 $Y=1.095 $X2=0 $Y2=0
cc_209 N_A_84_21#_c_212_n N_S1_c_287_n 0.00393355f $X=2.06 $Y=0.495 $X2=0 $Y2=0
cc_210 N_A_84_21#_c_213_n N_S1_c_289_n 0.00454584f $X=2.07 $Y=2.2 $X2=0 $Y2=0
cc_211 N_A_84_21#_c_210_n N_S1_c_296_n 0.00849309f $X=1.975 $Y=1.127 $X2=0 $Y2=0
cc_212 N_A_84_21#_c_211_n N_S1_c_296_n 0.00564489f $X=1.14 $Y=1.095 $X2=0 $Y2=0
cc_213 N_A_84_21#_M1005_g N_S1_c_298_n 3.48181e-19 $X=0.545 $Y=2.545 $X2=0 $Y2=0
cc_214 N_A_84_21#_c_210_n N_S1_c_298_n 0.0508228f $X=1.975 $Y=1.127 $X2=0 $Y2=0
cc_215 N_A_84_21#_c_211_n N_S1_c_298_n 9.88671e-19 $X=1.14 $Y=1.095 $X2=0 $Y2=0
cc_216 N_A_84_21#_c_213_n N_S1_c_298_n 0.0255053f $X=2.07 $Y=2.2 $X2=0 $Y2=0
cc_217 N_A_84_21#_c_213_n N_S1_c_307_n 0.037629f $X=2.07 $Y=2.2 $X2=0 $Y2=0
cc_218 N_A_84_21#_M1013_d N_S1_c_325_n 0.0121996f $X=1.85 $Y=2.055 $X2=0 $Y2=0
cc_219 N_A_84_21#_c_213_n N_S1_c_325_n 0.0130962f $X=2.07 $Y=2.2 $X2=0 $Y2=0
cc_220 N_A_84_21#_c_213_n N_S1_c_308_n 0.0320976f $X=2.07 $Y=2.2 $X2=0 $Y2=0
cc_221 N_A_84_21#_c_213_n S1 0.0263487f $X=2.07 $Y=2.2 $X2=0 $Y2=0
cc_222 N_A_84_21#_M1005_g N_S1_c_300_n 0.0107444f $X=0.545 $Y=2.545 $X2=0 $Y2=0
cc_223 N_A_84_21#_c_210_n N_S1_c_300_n 0.00564068f $X=1.975 $Y=1.127 $X2=0 $Y2=0
cc_224 N_A_84_21#_c_211_n N_S1_c_300_n 0.0169737f $X=1.14 $Y=1.095 $X2=0 $Y2=0
cc_225 N_A_84_21#_c_213_n N_A_320_366#_c_442_n 0.00338412f $X=2.07 $Y=2.2 $X2=0
+ $Y2=0
cc_226 N_A_84_21#_c_213_n N_A_320_366#_c_435_n 0.0143852f $X=2.07 $Y=2.2 $X2=0
+ $Y2=0
cc_227 N_A_84_21#_c_212_n N_A_320_366#_M1025_g 0.0070087f $X=2.06 $Y=0.495 $X2=0
+ $Y2=0
cc_228 N_A_84_21#_c_210_n N_A_320_366#_c_444_n 0.00373598f $X=1.975 $Y=1.127
+ $X2=0 $Y2=0
cc_229 N_A_84_21#_c_213_n N_A_320_366#_c_444_n 0.00638471f $X=2.07 $Y=2.2 $X2=0
+ $Y2=0
cc_230 N_A_84_21#_c_213_n N_A_320_366#_c_437_n 0.00425929f $X=2.07 $Y=2.2 $X2=0
+ $Y2=0
cc_231 N_A_84_21#_c_214_n N_A_320_366#_c_437_n 0.0222091f $X=2.065 $Y=1.127
+ $X2=0 $Y2=0
cc_232 N_A_84_21#_c_210_n N_A_320_366#_c_441_n 0.0037679f $X=1.975 $Y=1.127
+ $X2=0 $Y2=0
cc_233 N_A_84_21#_c_213_n N_A_320_366#_c_441_n 0.00418435f $X=2.07 $Y=2.2 $X2=0
+ $Y2=0
cc_234 N_A_84_21#_c_214_n N_A_320_366#_c_441_n 0.0100973f $X=2.065 $Y=1.127
+ $X2=0 $Y2=0
cc_235 N_A_84_21#_M1006_g X 0.0207681f $X=0.495 $Y=0.445 $X2=0 $Y2=0
cc_236 N_A_84_21#_M1005_g X 0.0519906f $X=0.545 $Y=2.545 $X2=0 $Y2=0
cc_237 N_A_84_21#_c_208_n X 0.00163211f $X=0.855 $Y=0.73 $X2=0 $Y2=0
cc_238 N_A_84_21#_c_209_n X 0.00552932f $X=0.545 $Y=1.185 $X2=0 $Y2=0
cc_239 N_A_84_21#_M1005_g N_VPWR_c_1127_n 0.0195419f $X=0.545 $Y=2.545 $X2=0
+ $Y2=0
cc_240 N_A_84_21#_M1005_g N_VPWR_c_1126_n 0.014085f $X=0.545 $Y=2.545 $X2=0
+ $Y2=0
cc_241 N_A_84_21#_M1005_g N_VPWR_c_1138_n 0.00769046f $X=0.545 $Y=2.545 $X2=0
+ $Y2=0
cc_242 N_A_84_21#_M1006_g N_A_245_411#_c_1224_n 0.00478961f $X=0.495 $Y=0.445
+ $X2=0 $Y2=0
cc_243 N_A_84_21#_M1005_g N_A_245_411#_c_1224_n 0.0223939f $X=0.545 $Y=2.545
+ $X2=0 $Y2=0
cc_244 N_A_84_21#_c_207_n N_A_245_411#_c_1224_n 0.00935388f $X=0.975 $Y=1.185
+ $X2=0 $Y2=0
cc_245 N_A_84_21#_c_209_n N_A_245_411#_c_1224_n 0.002958f $X=0.545 $Y=1.185
+ $X2=0 $Y2=0
cc_246 N_A_84_21#_c_210_n N_A_245_411#_c_1224_n 0.0195629f $X=1.975 $Y=1.127
+ $X2=0 $Y2=0
cc_247 N_A_84_21#_c_211_n N_A_245_411#_c_1224_n 0.00384531f $X=1.14 $Y=1.095
+ $X2=0 $Y2=0
cc_248 N_A_84_21#_c_207_n N_A_245_411#_c_1225_n 5.0882e-19 $X=0.975 $Y=1.185
+ $X2=0 $Y2=0
cc_249 N_A_84_21#_c_208_n N_A_245_411#_c_1225_n 0.00590357f $X=0.855 $Y=0.73
+ $X2=0 $Y2=0
cc_250 N_A_84_21#_c_210_n N_A_245_411#_c_1225_n 0.0601578f $X=1.975 $Y=1.127
+ $X2=0 $Y2=0
cc_251 N_A_84_21#_c_211_n N_A_245_411#_c_1225_n 0.0181987f $X=1.14 $Y=1.095
+ $X2=0 $Y2=0
cc_252 N_A_84_21#_c_212_n N_A_245_411#_c_1225_n 0.0107524f $X=2.06 $Y=0.495
+ $X2=0 $Y2=0
cc_253 N_A_84_21#_M1006_g N_A_245_411#_c_1226_n 0.00120086f $X=0.495 $Y=0.445
+ $X2=0 $Y2=0
cc_254 N_A_84_21#_c_208_n N_A_245_411#_c_1226_n 9.50782e-19 $X=0.855 $Y=0.73
+ $X2=0 $Y2=0
cc_255 N_A_84_21#_c_211_n N_A_245_411#_c_1226_n 6.11155e-19 $X=1.14 $Y=1.095
+ $X2=0 $Y2=0
cc_256 N_A_84_21#_M1005_g N_A_245_411#_c_1253_n 0.00880696f $X=0.545 $Y=2.545
+ $X2=0 $Y2=0
cc_257 N_A_84_21#_M1005_g N_A_245_411#_c_1232_n 3.95513e-19 $X=0.545 $Y=2.545
+ $X2=0 $Y2=0
cc_258 N_A_84_21#_M1005_g N_A_245_411#_c_1233_n 0.00521226f $X=0.545 $Y=2.545
+ $X2=0 $Y2=0
cc_259 N_A_84_21#_M1013_d N_A_245_411#_c_1234_n 0.00495203f $X=1.85 $Y=2.055
+ $X2=0 $Y2=0
cc_260 N_A_84_21#_c_208_n N_A_245_411#_c_1227_n 0.00327684f $X=0.855 $Y=0.73
+ $X2=0 $Y2=0
cc_261 N_A_84_21#_c_212_n N_A_245_411#_c_1227_n 0.0142704f $X=2.06 $Y=0.495
+ $X2=0 $Y2=0
cc_262 N_A_84_21#_c_212_n N_A_470_57#_c_1383_n 0.0178601f $X=2.06 $Y=0.495 $X2=0
+ $Y2=0
cc_263 N_A_84_21#_M1006_g N_VGND_c_1550_n 0.00182636f $X=0.495 $Y=0.445 $X2=0
+ $Y2=0
cc_264 N_A_84_21#_c_208_n N_VGND_c_1550_n 0.00992618f $X=0.855 $Y=0.73 $X2=0
+ $Y2=0
cc_265 N_A_84_21#_c_211_n N_VGND_c_1550_n 0.0010653f $X=1.14 $Y=1.095 $X2=0
+ $Y2=0
cc_266 N_A_84_21#_c_212_n N_VGND_c_1554_n 0.0113273f $X=2.06 $Y=0.495 $X2=0
+ $Y2=0
cc_267 N_A_84_21#_M1006_g N_VGND_c_1558_n 0.00549284f $X=0.495 $Y=0.445 $X2=0
+ $Y2=0
cc_268 N_A_84_21#_c_208_n N_VGND_c_1558_n 0.00354737f $X=0.855 $Y=0.73 $X2=0
+ $Y2=0
cc_269 N_A_84_21#_M1006_g N_VGND_c_1561_n 0.010905f $X=0.495 $Y=0.445 $X2=0
+ $Y2=0
cc_270 N_A_84_21#_c_208_n N_VGND_c_1561_n 0.00400114f $X=0.855 $Y=0.73 $X2=0
+ $Y2=0
cc_271 N_A_84_21#_c_212_n N_VGND_c_1561_n 0.00650045f $X=2.06 $Y=0.495 $X2=0
+ $Y2=0
cc_272 N_S1_c_289_n N_A_320_366#_c_442_n 0.0274325f $X=3.025 $Y=1.525 $X2=0
+ $Y2=0
cc_273 N_S1_c_307_n N_A_320_366#_c_442_n 0.0172452f $X=1.72 $Y=2.545 $X2=0 $Y2=0
cc_274 N_S1_c_325_n N_A_320_366#_c_442_n 0.006143f $X=2.335 $Y=2.63 $X2=0 $Y2=0
cc_275 N_S1_c_335_p N_A_320_366#_c_442_n 0.00623529f $X=1.805 $Y=2.63 $X2=0
+ $Y2=0
cc_276 N_S1_c_308_n N_A_320_366#_c_442_n 8.21354e-19 $X=2.42 $Y=2.545 $X2=0
+ $Y2=0
cc_277 N_S1_c_285_n N_A_320_366#_c_435_n 0.0119502f $X=1.545 $Y=1.545 $X2=0
+ $Y2=0
cc_278 N_S1_c_289_n N_A_320_366#_c_435_n 0.0115845f $X=3.025 $Y=1.525 $X2=0
+ $Y2=0
cc_279 N_S1_c_298_n N_A_320_366#_c_435_n 0.00281667f $X=1.635 $Y=1.635 $X2=0
+ $Y2=0
cc_280 N_S1_c_307_n N_A_320_366#_c_435_n 5.84409e-19 $X=1.72 $Y=2.545 $X2=0
+ $Y2=0
cc_281 S1 N_A_320_366#_c_435_n 0.0011383f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_282 N_S1_c_300_n N_A_320_366#_c_435_n 0.0023981f $X=1.195 $Y=1.545 $X2=0
+ $Y2=0
cc_283 N_S1_c_286_n N_A_320_366#_M1025_g 0.0040815f $X=1.62 $Y=1.47 $X2=0 $Y2=0
cc_284 N_S1_c_287_n N_A_320_366#_M1025_g 0.0155289f $X=1.845 $Y=0.78 $X2=0 $Y2=0
cc_285 N_S1_c_285_n N_A_320_366#_c_444_n 0.00623493f $X=1.545 $Y=1.545 $X2=0
+ $Y2=0
cc_286 N_S1_c_289_n N_A_320_366#_c_444_n 0.0046586f $X=3.025 $Y=1.525 $X2=0
+ $Y2=0
cc_287 N_S1_c_298_n N_A_320_366#_c_444_n 9.71934e-19 $X=1.635 $Y=1.635 $X2=0
+ $Y2=0
cc_288 N_S1_c_307_n N_A_320_366#_c_444_n 0.0127588f $X=1.72 $Y=2.545 $X2=0 $Y2=0
cc_289 N_S1_c_325_n N_A_320_366#_c_444_n 0.00298537f $X=2.335 $Y=2.63 $X2=0
+ $Y2=0
cc_290 N_S1_c_289_n N_A_320_366#_c_437_n 0.00543819f $X=3.025 $Y=1.525 $X2=0
+ $Y2=0
cc_291 S1 N_A_320_366#_c_437_n 0.0269724f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_292 N_S1_c_290_n N_A_320_366#_c_438_n 0.00739798f $X=3.345 $Y=1 $X2=0 $Y2=0
cc_293 N_S1_c_288_n N_A_320_366#_c_439_n 0.0169021f $X=3.27 $Y=1.525 $X2=0 $Y2=0
cc_294 N_S1_c_289_n N_A_320_366#_c_439_n 8.40573e-19 $X=3.025 $Y=1.525 $X2=0
+ $Y2=0
cc_295 N_S1_c_291_n N_A_320_366#_c_439_n 0.00393255f $X=3.345 $Y=1.45 $X2=0
+ $Y2=0
cc_296 N_S1_M1022_g N_A_320_366#_c_439_n 4.39693e-19 $X=3.675 $Y=2.595 $X2=0
+ $Y2=0
cc_297 S1 N_A_320_366#_c_439_n 0.00520614f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_298 N_S1_c_289_n N_A_320_366#_c_440_n 0.00716255f $X=3.025 $Y=1.525 $X2=0
+ $Y2=0
cc_299 N_S1_c_290_n N_A_320_366#_c_440_n 0.00478236f $X=3.345 $Y=1 $X2=0 $Y2=0
cc_300 N_S1_c_288_n N_A_320_366#_c_446_n 0.0108011f $X=3.27 $Y=1.525 $X2=0 $Y2=0
cc_301 N_S1_c_289_n N_A_320_366#_c_446_n 0.00380821f $X=3.025 $Y=1.525 $X2=0
+ $Y2=0
cc_302 N_S1_M1022_g N_A_320_366#_c_446_n 0.00675139f $X=3.675 $Y=2.595 $X2=0
+ $Y2=0
cc_303 N_S1_c_308_n N_A_320_366#_c_446_n 0.00302561f $X=2.42 $Y=2.545 $X2=0
+ $Y2=0
cc_304 S1 N_A_320_366#_c_446_n 0.0128001f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_305 N_S1_c_286_n N_A_320_366#_c_441_n 0.0119502f $X=1.62 $Y=1.47 $X2=0 $Y2=0
cc_306 N_S1_c_289_n N_A_320_366#_c_441_n 0.0145032f $X=3.025 $Y=1.525 $X2=0
+ $Y2=0
cc_307 N_S1_c_290_n N_A_320_366#_c_441_n 0.00423749f $X=3.345 $Y=1 $X2=0 $Y2=0
cc_308 S1 N_A_320_366#_c_441_n 0.00234775f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_309 N_S1_M1022_g N_A3_M1002_g 0.0371507f $X=3.675 $Y=2.595 $X2=0 $Y2=0
cc_310 N_S1_c_293_n N_A3_c_522_n 0.00263899f $X=3.675 $Y=1.6 $X2=0 $Y2=0
cc_311 N_S1_c_295_n N_A3_c_523_n 0.00435161f $X=3.705 $Y=1 $X2=0 $Y2=0
cc_312 N_S1_c_292_n N_A3_c_524_n 0.00249474f $X=3.63 $Y=1.075 $X2=0 $Y2=0
cc_313 N_S1_c_293_n A3 0.00442033f $X=3.675 $Y=1.6 $X2=0 $Y2=0
cc_314 N_S1_c_293_n N_A3_c_526_n 0.0192879f $X=3.675 $Y=1.6 $X2=0 $Y2=0
cc_315 N_S1_M1022_g N_VPWR_c_1128_n 0.00476179f $X=3.675 $Y=2.595 $X2=0 $Y2=0
cc_316 N_S1_c_301_n N_VPWR_c_1135_n 0.00556532f $X=2.45 $Y=2.015 $X2=0 $Y2=0
cc_317 N_S1_M1022_g N_VPWR_c_1135_n 0.00710941f $X=3.675 $Y=2.595 $X2=0 $Y2=0
cc_318 N_S1_c_301_n N_VPWR_c_1126_n 0.0088375f $X=2.45 $Y=2.015 $X2=0 $Y2=0
cc_319 N_S1_M1022_g N_VPWR_c_1126_n 0.0106422f $X=3.675 $Y=2.595 $X2=0 $Y2=0
cc_320 N_S1_c_298_n N_A_245_411#_c_1224_n 0.0205268f $X=1.635 $Y=1.635 $X2=0
+ $Y2=0
cc_321 N_S1_c_300_n N_A_245_411#_c_1224_n 0.00115317f $X=1.195 $Y=1.545 $X2=0
+ $Y2=0
cc_322 N_S1_c_287_n N_A_245_411#_c_1225_n 0.00334114f $X=1.845 $Y=0.78 $X2=0
+ $Y2=0
cc_323 N_S1_c_296_n N_A_245_411#_c_1225_n 0.0098201f $X=1.845 $Y=0.855 $X2=0
+ $Y2=0
cc_324 N_S1_c_285_n N_A_245_411#_c_1231_n 4.98296e-19 $X=1.545 $Y=1.545 $X2=0
+ $Y2=0
cc_325 N_S1_c_298_n N_A_245_411#_c_1231_n 0.0331524f $X=1.635 $Y=1.635 $X2=0
+ $Y2=0
cc_326 N_S1_c_307_n N_A_245_411#_c_1231_n 0.0129384f $X=1.72 $Y=2.545 $X2=0
+ $Y2=0
cc_327 N_S1_c_300_n N_A_245_411#_c_1231_n 0.00748916f $X=1.195 $Y=1.545 $X2=0
+ $Y2=0
cc_328 N_S1_c_307_n N_A_245_411#_c_1233_n 0.0272825f $X=1.72 $Y=2.545 $X2=0
+ $Y2=0
cc_329 N_S1_c_335_p N_A_245_411#_c_1233_n 0.0131328f $X=1.805 $Y=2.63 $X2=0
+ $Y2=0
cc_330 N_S1_c_301_n N_A_245_411#_c_1234_n 0.0184812f $X=2.45 $Y=2.015 $X2=0
+ $Y2=0
cc_331 N_S1_M1022_g N_A_245_411#_c_1234_n 0.00417077f $X=3.675 $Y=2.595 $X2=0
+ $Y2=0
cc_332 N_S1_c_325_n N_A_245_411#_c_1234_n 0.0382906f $X=2.335 $Y=2.63 $X2=0
+ $Y2=0
cc_333 N_S1_c_335_p N_A_245_411#_c_1234_n 0.0114486f $X=1.805 $Y=2.63 $X2=0
+ $Y2=0
cc_334 N_S1_c_287_n N_A_245_411#_c_1227_n 0.00481483f $X=1.845 $Y=0.78 $X2=0
+ $Y2=0
cc_335 N_S1_c_301_n N_A_245_411#_c_1235_n 0.00446511f $X=2.45 $Y=2.015 $X2=0
+ $Y2=0
cc_336 N_S1_M1022_g N_A_245_411#_c_1235_n 0.00655757f $X=3.675 $Y=2.595 $X2=0
+ $Y2=0
cc_337 N_S1_M1022_g N_A_245_411#_c_1276_n 0.020721f $X=3.675 $Y=2.595 $X2=0
+ $Y2=0
cc_338 N_S1_c_290_n N_A_470_57#_c_1370_n 0.0104769f $X=3.345 $Y=1 $X2=0 $Y2=0
cc_339 N_S1_c_295_n N_A_470_57#_c_1370_n 4.426e-19 $X=3.705 $Y=1 $X2=0 $Y2=0
cc_340 N_S1_c_301_n N_A_470_57#_c_1385_n 0.00269994f $X=2.45 $Y=2.015 $X2=0
+ $Y2=0
cc_341 N_S1_M1022_g N_A_470_57#_c_1385_n 0.00486181f $X=3.675 $Y=2.595 $X2=0
+ $Y2=0
cc_342 N_S1_c_325_n N_A_470_57#_c_1385_n 0.0131327f $X=2.335 $Y=2.63 $X2=0 $Y2=0
cc_343 N_S1_c_308_n N_A_470_57#_c_1385_n 0.0144721f $X=2.42 $Y=2.545 $X2=0 $Y2=0
cc_344 N_S1_c_288_n N_A_470_57#_c_1386_n 4.54873e-19 $X=3.27 $Y=1.525 $X2=0
+ $Y2=0
cc_345 N_S1_c_289_n N_A_470_57#_c_1386_n 0.00242009f $X=3.025 $Y=1.525 $X2=0
+ $Y2=0
cc_346 N_S1_c_293_n N_A_470_57#_c_1386_n 0.00265854f $X=3.675 $Y=1.6 $X2=0 $Y2=0
cc_347 N_S1_M1022_g N_A_470_57#_c_1386_n 0.0156705f $X=3.675 $Y=2.595 $X2=0
+ $Y2=0
cc_348 N_S1_c_301_n N_A_470_57#_c_1387_n 0.00223949f $X=2.45 $Y=2.015 $X2=0
+ $Y2=0
cc_349 N_S1_c_289_n N_A_470_57#_c_1387_n 0.00691129f $X=3.025 $Y=1.525 $X2=0
+ $Y2=0
cc_350 N_S1_c_308_n N_A_470_57#_c_1387_n 0.0128379f $X=2.42 $Y=2.545 $X2=0 $Y2=0
cc_351 S1 N_A_470_57#_c_1387_n 0.00393582f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_352 N_S1_c_290_n N_A_470_57#_c_1371_n 0.0145527f $X=3.345 $Y=1 $X2=0 $Y2=0
cc_353 N_S1_c_292_n N_A_470_57#_c_1371_n 0.00583894f $X=3.63 $Y=1.075 $X2=0
+ $Y2=0
cc_354 N_S1_c_295_n N_A_470_57#_c_1371_n 0.00377817f $X=3.705 $Y=1 $X2=0 $Y2=0
cc_355 N_S1_c_297_n N_A_470_57#_c_1371_n 0.00152064f $X=3.345 $Y=1.075 $X2=0
+ $Y2=0
cc_356 N_S1_c_291_n N_A_470_57#_c_1372_n 0.00138184f $X=3.345 $Y=1.45 $X2=0
+ $Y2=0
cc_357 N_S1_c_293_n N_A_470_57#_c_1372_n 0.0088796f $X=3.675 $Y=1.6 $X2=0 $Y2=0
cc_358 N_S1_M1022_g N_A_470_57#_c_1372_n 0.0218798f $X=3.675 $Y=2.595 $X2=0
+ $Y2=0
cc_359 N_S1_c_292_n N_A_470_57#_c_1373_n 7.93859e-19 $X=3.63 $Y=1.075 $X2=0
+ $Y2=0
cc_360 N_S1_c_291_n N_A_470_57#_c_1374_n 0.00341825f $X=3.345 $Y=1.45 $X2=0
+ $Y2=0
cc_361 N_S1_c_292_n N_A_470_57#_c_1374_n 0.0124443f $X=3.63 $Y=1.075 $X2=0 $Y2=0
cc_362 N_S1_c_293_n N_A_470_57#_c_1374_n 0.0051919f $X=3.675 $Y=1.6 $X2=0 $Y2=0
cc_363 N_S1_c_297_n N_A_470_57#_c_1374_n 3.40191e-19 $X=3.345 $Y=1.075 $X2=0
+ $Y2=0
cc_364 N_S1_c_295_n N_A_470_57#_c_1375_n 0.00255917f $X=3.705 $Y=1 $X2=0 $Y2=0
cc_365 N_S1_c_290_n N_A_470_57#_c_1383_n 0.00451449f $X=3.345 $Y=1 $X2=0 $Y2=0
cc_366 N_S1_c_287_n N_VGND_c_1550_n 0.00226784f $X=1.845 $Y=0.78 $X2=0 $Y2=0
cc_367 N_S1_c_290_n N_VGND_c_1551_n 4.62581e-19 $X=3.345 $Y=1 $X2=0 $Y2=0
cc_368 N_S1_c_295_n N_VGND_c_1551_n 0.0095274f $X=3.705 $Y=1 $X2=0 $Y2=0
cc_369 N_S1_c_287_n N_VGND_c_1554_n 0.00502664f $X=1.845 $Y=0.78 $X2=0 $Y2=0
cc_370 N_S1_c_290_n N_VGND_c_1554_n 7.27864e-19 $X=3.345 $Y=1 $X2=0 $Y2=0
cc_371 N_S1_c_295_n N_VGND_c_1554_n 0.00402651f $X=3.705 $Y=1 $X2=0 $Y2=0
cc_372 N_S1_c_296_n N_VGND_c_1554_n 4.81257e-19 $X=1.845 $Y=0.855 $X2=0 $Y2=0
cc_373 N_S1_c_287_n N_VGND_c_1561_n 0.010456f $X=1.845 $Y=0.78 $X2=0 $Y2=0
cc_374 N_S1_c_295_n N_VGND_c_1561_n 0.00423264f $X=3.705 $Y=1 $X2=0 $Y2=0
cc_375 N_A_320_366#_c_442_n N_VPWR_c_1127_n 0.00323237f $X=1.725 $Y=1.98 $X2=0
+ $Y2=0
cc_376 N_A_320_366#_c_442_n N_VPWR_c_1135_n 0.00556532f $X=1.725 $Y=1.98 $X2=0
+ $Y2=0
cc_377 N_A_320_366#_M1022_s N_VPWR_c_1126_n 0.00398722f $X=3.185 $Y=1.675 $X2=0
+ $Y2=0
cc_378 N_A_320_366#_c_442_n N_VPWR_c_1126_n 0.0088375f $X=1.725 $Y=1.98 $X2=0
+ $Y2=0
cc_379 N_A_320_366#_c_442_n N_A_245_411#_c_1231_n 0.0038744f $X=1.725 $Y=1.98
+ $X2=0 $Y2=0
cc_380 N_A_320_366#_c_442_n N_A_245_411#_c_1233_n 0.0195137f $X=1.725 $Y=1.98
+ $X2=0 $Y2=0
cc_381 N_A_320_366#_M1022_s N_A_245_411#_c_1234_n 0.00451394f $X=3.185 $Y=1.675
+ $X2=0 $Y2=0
cc_382 N_A_320_366#_c_442_n N_A_245_411#_c_1234_n 0.0170224f $X=1.725 $Y=1.98
+ $X2=0 $Y2=0
cc_383 N_A_320_366#_M1022_s N_A_245_411#_c_1235_n 0.00379262f $X=3.185 $Y=1.675
+ $X2=0 $Y2=0
cc_384 N_A_320_366#_M1022_s N_A_245_411#_c_1276_n 0.00668635f $X=3.185 $Y=1.675
+ $X2=0 $Y2=0
cc_385 N_A_320_366#_M1022_s N_A_245_411#_c_1236_n 0.00207005f $X=3.185 $Y=1.675
+ $X2=0 $Y2=0
cc_386 N_A_320_366#_c_437_n N_A_470_57#_c_1370_n 0.00796773f $X=2.885 $Y=1.155
+ $X2=0 $Y2=0
cc_387 N_A_320_366#_c_438_n N_A_470_57#_c_1370_n 0.0242908f $X=3.05 $Y=0.78
+ $X2=0 $Y2=0
cc_388 N_A_320_366#_M1022_s N_A_470_57#_c_1386_n 0.00862078f $X=3.185 $Y=1.675
+ $X2=0 $Y2=0
cc_389 N_A_320_366#_c_446_n N_A_470_57#_c_1386_n 0.0275074f $X=3.33 $Y=1.82
+ $X2=0 $Y2=0
cc_390 N_A_320_366#_c_438_n N_A_470_57#_c_1371_n 0.0146569f $X=3.05 $Y=0.78
+ $X2=0 $Y2=0
cc_391 N_A_320_366#_c_440_n N_A_470_57#_c_1371_n 0.0104004f $X=3.05 $Y=1.155
+ $X2=0 $Y2=0
cc_392 N_A_320_366#_c_439_n N_A_470_57#_c_1372_n 0.0130459f $X=3.13 $Y=1.655
+ $X2=0 $Y2=0
cc_393 N_A_320_366#_c_440_n N_A_470_57#_c_1372_n 0.00120313f $X=3.05 $Y=1.155
+ $X2=0 $Y2=0
cc_394 N_A_320_366#_c_446_n N_A_470_57#_c_1372_n 0.0235821f $X=3.33 $Y=1.82
+ $X2=0 $Y2=0
cc_395 N_A_320_366#_c_440_n N_A_470_57#_c_1374_n 0.0142981f $X=3.05 $Y=1.155
+ $X2=0 $Y2=0
cc_396 N_A_320_366#_c_446_n N_A_470_57#_c_1374_n 8.64673e-19 $X=3.33 $Y=1.82
+ $X2=0 $Y2=0
cc_397 N_A_320_366#_M1025_g N_A_470_57#_c_1383_n 0.0070399f $X=2.275 $Y=0.495
+ $X2=0 $Y2=0
cc_398 N_A_320_366#_c_437_n N_A_470_57#_c_1383_n 0.0186362f $X=2.885 $Y=1.155
+ $X2=0 $Y2=0
cc_399 N_A_320_366#_c_438_n N_A_470_57#_c_1383_n 0.0074161f $X=3.05 $Y=0.78
+ $X2=0 $Y2=0
cc_400 N_A_320_366#_c_441_n N_A_470_57#_c_1383_n 0.00660528f $X=2.275 $Y=1.155
+ $X2=0 $Y2=0
cc_401 N_A_320_366#_M1025_g N_VGND_c_1554_n 0.00502664f $X=2.275 $Y=0.495 $X2=0
+ $Y2=0
cc_402 N_A_320_366#_M1025_g N_VGND_c_1561_n 0.010456f $X=2.275 $Y=0.495 $X2=0
+ $Y2=0
cc_403 N_A3_c_522_n N_S0_c_573_n 0.00540522f $X=4.415 $Y=1.55 $X2=0 $Y2=0
cc_404 N_A3_c_524_n N_S0_c_573_n 0.00420284f $X=4.5 $Y=1.075 $X2=0 $Y2=0
cc_405 N_A3_c_523_n N_S0_c_586_n 0.0246693f $X=4.5 $Y=1 $X2=0 $Y2=0
cc_406 N_A3_M1002_g N_A_946_317#_M1015_g 0.042919f $X=4.365 $Y=2.595 $X2=0 $Y2=0
cc_407 N_A3_c_526_n N_A_946_317#_c_793_n 0.042919f $X=4.415 $Y=1.715 $X2=0 $Y2=0
cc_408 A3 N_VPWR_M1022_d 0.00424199f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_409 N_A3_M1002_g N_VPWR_c_1128_n 0.00476179f $X=4.365 $Y=2.595 $X2=0 $Y2=0
cc_410 N_A3_M1002_g N_VPWR_c_1131_n 0.00710941f $X=4.365 $Y=2.595 $X2=0 $Y2=0
cc_411 N_A3_M1002_g N_VPWR_c_1126_n 0.00913969f $X=4.365 $Y=2.595 $X2=0 $Y2=0
cc_412 N_A3_M1002_g N_A_245_411#_c_1276_n 0.0227229f $X=4.365 $Y=2.595 $X2=0
+ $Y2=0
cc_413 A3 N_A_245_411#_c_1276_n 0.0143783f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_414 N_A3_c_526_n N_A_245_411#_c_1276_n 7.15e-19 $X=4.415 $Y=1.715 $X2=0 $Y2=0
cc_415 N_A3_c_522_n N_A_245_411#_c_1228_n 0.016772f $X=4.415 $Y=1.55 $X2=0 $Y2=0
cc_416 N_A3_c_523_n N_A_245_411#_c_1228_n 0.00264951f $X=4.5 $Y=1 $X2=0 $Y2=0
cc_417 N_A3_c_524_n N_A_245_411#_c_1228_n 0.00475245f $X=4.5 $Y=1.075 $X2=0
+ $Y2=0
cc_418 A3 N_A_245_411#_c_1228_n 0.0407859f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_419 N_A3_c_523_n N_A_245_411#_c_1291_n 0.00689729f $X=4.5 $Y=1 $X2=0 $Y2=0
cc_420 N_A3_M1002_g N_A_245_411#_c_1292_n 0.00164029f $X=4.365 $Y=2.595 $X2=0
+ $Y2=0
cc_421 N_A3_M1002_g N_A_470_57#_c_1386_n 9.46887e-19 $X=4.365 $Y=2.595 $X2=0
+ $Y2=0
cc_422 N_A3_M1002_g N_A_470_57#_c_1372_n 3.08636e-19 $X=4.365 $Y=2.595 $X2=0
+ $Y2=0
cc_423 N_A3_c_522_n N_A_470_57#_c_1372_n 0.00397367f $X=4.415 $Y=1.55 $X2=0
+ $Y2=0
cc_424 A3 N_A_470_57#_c_1372_n 0.0405332f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_425 N_A3_c_526_n N_A_470_57#_c_1372_n 3.55881e-19 $X=4.415 $Y=1.715 $X2=0
+ $Y2=0
cc_426 N_A3_c_522_n N_A_470_57#_c_1373_n 0.0053754f $X=4.415 $Y=1.55 $X2=0 $Y2=0
cc_427 N_A3_c_524_n N_A_470_57#_c_1373_n 8.61822e-19 $X=4.5 $Y=1.075 $X2=0 $Y2=0
cc_428 A3 N_A_470_57#_c_1373_n 0.0236294f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_429 N_A3_c_526_n N_A_470_57#_c_1373_n 0.00222585f $X=4.415 $Y=1.715 $X2=0
+ $Y2=0
cc_430 N_A3_c_523_n N_A_470_57#_c_1375_n 0.00911956f $X=4.5 $Y=1 $X2=0 $Y2=0
cc_431 N_A3_c_524_n N_A_470_57#_c_1375_n 0.00372307f $X=4.5 $Y=1.075 $X2=0 $Y2=0
cc_432 N_A3_c_523_n N_A_470_57#_c_1376_n 0.0104098f $X=4.5 $Y=1 $X2=0 $Y2=0
cc_433 N_A3_c_524_n N_A_470_57#_c_1376_n 0.00191382f $X=4.5 $Y=1.075 $X2=0 $Y2=0
cc_434 N_A3_c_523_n N_VGND_c_1551_n 9.58275e-19 $X=4.5 $Y=1 $X2=0 $Y2=0
cc_435 N_A3_c_523_n N_VGND_c_1556_n 7.10185e-19 $X=4.5 $Y=1 $X2=0 $Y2=0
cc_436 N_S0_c_589_n N_A_946_317#_M1028_d 8.72743e-19 $X=9.455 $Y=1.77 $X2=0
+ $Y2=0
cc_437 N_S0_c_582_n N_A_946_317#_c_779_n 3.15372e-19 $X=5.565 $Y=1.245 $X2=0
+ $Y2=0
cc_438 N_S0_c_573_n N_A_946_317#_M1011_g 0.0213362f $X=5.035 $Y=1.21 $X2=0 $Y2=0
cc_439 N_S0_c_582_n N_A_946_317#_M1011_g 0.021801f $X=5.565 $Y=1.245 $X2=0 $Y2=0
cc_440 N_S0_c_583_n N_A_946_317#_M1011_g 0.00223814f $X=5.98 $Y=1.36 $X2=0 $Y2=0
cc_441 N_S0_c_584_n N_A_946_317#_M1011_g 0.0175302f $X=5.98 $Y=1.595 $X2=0 $Y2=0
cc_442 N_S0_c_586_n N_A_946_317#_M1011_g 0.017703f $X=5.035 $Y=1.045 $X2=0 $Y2=0
cc_443 N_S0_M1004_g N_A_946_317#_M1023_g 0.023725f $X=8.335 $Y=2.595 $X2=0 $Y2=0
cc_444 N_S0_c_614_p N_A_946_317#_M1023_g 0.0231149f $X=7.525 $Y=2.545 $X2=0
+ $Y2=0
cc_445 N_S0_c_615_p N_A_946_317#_M1023_g 0.00640239f $X=8.18 $Y=2.63 $X2=0 $Y2=0
cc_446 N_S0_c_616_p N_A_946_317#_M1023_g 0.00613589f $X=7.61 $Y=2.63 $X2=0 $Y2=0
cc_447 N_S0_c_587_n N_A_946_317#_M1023_g 0.00218291f $X=8.345 $Y=1.77 $X2=0
+ $Y2=0
cc_448 N_S0_c_580_n N_A_946_317#_c_782_n 0.0113388f $X=7.445 $Y=1.245 $X2=0
+ $Y2=0
cc_449 N_S0_c_614_p N_A_946_317#_c_782_n 0.0016482f $X=7.525 $Y=2.545 $X2=0
+ $Y2=0
cc_450 N_S0_c_585_n N_A_946_317#_c_782_n 0.00880328f $X=7.445 $Y=1.675 $X2=0
+ $Y2=0
cc_451 N_S0_c_579_n N_A_946_317#_c_783_n 0.00123283f $X=7.445 $Y=1.245 $X2=0
+ $Y2=0
cc_452 N_S0_c_596_n N_A_946_317#_c_783_n 6.0922e-19 $X=8.265 $Y=2.15 $X2=0 $Y2=0
cc_453 N_S0_c_585_n N_A_946_317#_c_783_n 4.3694e-19 $X=7.445 $Y=1.675 $X2=0
+ $Y2=0
cc_454 N_S0_c_587_n N_A_946_317#_c_783_n 0.0126146f $X=8.345 $Y=1.77 $X2=0 $Y2=0
cc_455 N_S0_M1019_g N_A_946_317#_c_784_n 0.0179217f $X=7.385 $Y=0.445 $X2=0
+ $Y2=0
cc_456 N_S0_M1019_g N_A_946_317#_c_785_n 0.00404858f $X=7.385 $Y=0.445 $X2=0
+ $Y2=0
cc_457 N_S0_c_579_n N_A_946_317#_c_785_n 3.93205e-19 $X=7.445 $Y=1.245 $X2=0
+ $Y2=0
cc_458 N_S0_c_580_n N_A_946_317#_c_785_n 0.0205496f $X=7.445 $Y=1.245 $X2=0
+ $Y2=0
cc_459 N_S0_c_581_n N_A_946_317#_c_799_n 0.00828215f $X=5.395 $Y=1.245 $X2=0
+ $Y2=0
cc_460 N_S0_c_582_n N_A_946_317#_c_799_n 0.00355478f $X=5.565 $Y=1.245 $X2=0
+ $Y2=0
cc_461 N_S0_M1008_g N_A_946_317#_c_800_n 0.0237439f $X=5.925 $Y=2.595 $X2=0
+ $Y2=0
cc_462 N_S0_c_574_n N_A_946_317#_c_800_n 0.00635776f $X=5.815 $Y=1.36 $X2=0
+ $Y2=0
cc_463 N_S0_c_575_n N_A_946_317#_c_800_n 0.00645348f $X=6.325 $Y=1.36 $X2=0
+ $Y2=0
cc_464 N_S0_c_577_n N_A_946_317#_c_800_n 0.0539694f $X=7.28 $Y=1.675 $X2=0 $Y2=0
cc_465 N_S0_c_578_n N_A_946_317#_c_800_n 0.0122682f $X=6.495 $Y=1.675 $X2=0
+ $Y2=0
cc_466 N_S0_c_614_p N_A_946_317#_c_800_n 0.0131128f $X=7.525 $Y=2.545 $X2=0
+ $Y2=0
cc_467 N_S0_c_583_n N_A_946_317#_c_800_n 0.0235528f $X=5.98 $Y=1.36 $X2=0 $Y2=0
cc_468 N_S0_c_584_n N_A_946_317#_c_800_n 6.54454e-19 $X=5.98 $Y=1.595 $X2=0
+ $Y2=0
cc_469 N_S0_c_614_p N_A_946_317#_c_841_n 0.0291541f $X=7.525 $Y=2.545 $X2=0
+ $Y2=0
cc_470 N_S0_c_616_p N_A_946_317#_c_841_n 0.0127795f $X=7.61 $Y=2.63 $X2=0 $Y2=0
cc_471 N_S0_M1004_g N_A_946_317#_c_843_n 0.0182381f $X=8.335 $Y=2.595 $X2=0
+ $Y2=0
cc_472 N_S0_c_615_p N_A_946_317#_c_843_n 0.0409707f $X=8.18 $Y=2.63 $X2=0 $Y2=0
cc_473 N_S0_c_616_p N_A_946_317#_c_843_n 0.0114161f $X=7.61 $Y=2.63 $X2=0 $Y2=0
cc_474 N_S0_c_572_n N_A_946_317#_c_786_n 0.0183754f $X=9.585 $Y=0.805 $X2=0
+ $Y2=0
cc_475 N_S0_c_588_n N_A_946_317#_c_786_n 0.00261212f $X=9.455 $Y=1.77 $X2=0
+ $Y2=0
cc_476 N_S0_c_589_n N_A_946_317#_c_786_n 0.00426014f $X=9.455 $Y=1.77 $X2=0
+ $Y2=0
cc_477 N_S0_c_590_n N_A_946_317#_c_786_n 0.00991423f $X=9.455 $Y=1.605 $X2=0
+ $Y2=0
cc_478 N_S0_M1004_g N_A_946_317#_c_850_n 0.00534229f $X=8.335 $Y=2.595 $X2=0
+ $Y2=0
cc_479 N_S0_M1028_g N_A_946_317#_c_850_n 8.79206e-19 $X=9.415 $Y=2.595 $X2=0
+ $Y2=0
cc_480 N_S0_c_615_p N_A_946_317#_c_850_n 0.00896052f $X=8.18 $Y=2.63 $X2=0 $Y2=0
cc_481 N_S0_c_651_p N_A_946_317#_c_850_n 0.002079f $X=8.265 $Y=2.545 $X2=0 $Y2=0
cc_482 N_S0_M1028_g N_A_946_317#_c_854_n 0.0138442f $X=9.415 $Y=2.595 $X2=0
+ $Y2=0
cc_483 N_S0_c_589_n N_A_946_317#_c_854_n 0.0429652f $X=9.455 $Y=1.77 $X2=0 $Y2=0
cc_484 N_S0_M1004_g N_A_946_317#_c_856_n 0.00147421f $X=8.335 $Y=2.595 $X2=0
+ $Y2=0
cc_485 N_S0_c_651_p N_A_946_317#_c_856_n 0.00902915f $X=8.265 $Y=2.545 $X2=0
+ $Y2=0
cc_486 N_S0_c_589_n N_A_946_317#_c_856_n 0.00921165f $X=9.455 $Y=1.77 $X2=0
+ $Y2=0
cc_487 N_S0_c_570_n N_A_946_317#_c_787_n 0.0013866f $X=9.225 $Y=0.73 $X2=0 $Y2=0
cc_488 N_S0_c_571_n N_A_946_317#_c_787_n 0.0093683f $X=9.585 $Y=0.73 $X2=0 $Y2=0
cc_489 N_S0_c_572_n N_A_946_317#_c_787_n 0.00870351f $X=9.585 $Y=0.805 $X2=0
+ $Y2=0
cc_490 N_S0_M1028_g N_A_946_317#_c_788_n 0.00553621f $X=9.415 $Y=2.595 $X2=0
+ $Y2=0
cc_491 N_S0_c_588_n N_A_946_317#_c_788_n 0.00338477f $X=9.455 $Y=1.77 $X2=0
+ $Y2=0
cc_492 N_S0_c_589_n N_A_946_317#_c_788_n 0.0396803f $X=9.455 $Y=1.77 $X2=0 $Y2=0
cc_493 N_S0_c_590_n N_A_946_317#_c_788_n 0.00917137f $X=9.455 $Y=1.605 $X2=0
+ $Y2=0
cc_494 N_S0_c_573_n N_A_946_317#_c_789_n 0.00117858f $X=5.035 $Y=1.21 $X2=0
+ $Y2=0
cc_495 N_S0_c_581_n N_A_946_317#_c_789_n 0.0209342f $X=5.395 $Y=1.245 $X2=0
+ $Y2=0
cc_496 N_S0_c_583_n N_A_946_317#_c_789_n 0.00422602f $X=5.98 $Y=1.36 $X2=0 $Y2=0
cc_497 N_S0_c_584_n N_A_946_317#_c_789_n 3.78332e-19 $X=5.98 $Y=1.595 $X2=0
+ $Y2=0
cc_498 N_S0_M1008_g N_A_946_317#_c_803_n 8.40163e-19 $X=5.925 $Y=2.595 $X2=0
+ $Y2=0
cc_499 N_S0_c_582_n N_A_946_317#_c_803_n 0.00898593f $X=5.565 $Y=1.245 $X2=0
+ $Y2=0
cc_500 N_S0_c_583_n N_A_946_317#_c_803_n 0.0010798f $X=5.98 $Y=1.36 $X2=0 $Y2=0
cc_501 N_S0_c_584_n N_A_946_317#_c_803_n 0.00488911f $X=5.98 $Y=1.595 $X2=0
+ $Y2=0
cc_502 N_S0_c_596_n N_A_946_317#_c_790_n 4.43735e-19 $X=8.265 $Y=2.15 $X2=0
+ $Y2=0
cc_503 N_S0_c_587_n N_A_946_317#_c_790_n 0.00550103f $X=8.345 $Y=1.77 $X2=0
+ $Y2=0
cc_504 N_S0_c_596_n N_A_946_317#_c_791_n 0.0028536f $X=8.265 $Y=2.15 $X2=0 $Y2=0
cc_505 N_S0_c_587_n N_A_946_317#_c_791_n 4.94591e-19 $X=8.345 $Y=1.77 $X2=0
+ $Y2=0
cc_506 N_S0_M1028_g N_A_946_317#_c_804_n 0.0115954f $X=9.415 $Y=2.595 $X2=0
+ $Y2=0
cc_507 N_S0_c_588_n N_A_946_317#_c_804_n 2.70301e-19 $X=9.455 $Y=1.77 $X2=0
+ $Y2=0
cc_508 N_S0_c_589_n N_A_946_317#_c_804_n 0.00386371f $X=9.455 $Y=1.77 $X2=0
+ $Y2=0
cc_509 N_S0_c_572_n N_A_946_317#_c_792_n 8.86742e-19 $X=9.585 $Y=0.805 $X2=0
+ $Y2=0
cc_510 N_S0_c_573_n N_A_946_317#_c_793_n 0.0216115f $X=5.035 $Y=1.21 $X2=0 $Y2=0
cc_511 N_S0_c_581_n N_A_946_317#_c_793_n 0.00428109f $X=5.395 $Y=1.245 $X2=0
+ $Y2=0
cc_512 N_S0_c_584_n N_A_946_317#_c_793_n 0.00248089f $X=5.98 $Y=1.595 $X2=0
+ $Y2=0
cc_513 N_S0_c_575_n N_A2_c_972_n 0.00597575f $X=6.325 $Y=1.36 $X2=0 $Y2=0
cc_514 N_S0_M1008_g N_A2_c_973_n 0.0683052f $X=5.925 $Y=2.595 $X2=0 $Y2=0
cc_515 N_S0_c_577_n N_A2_c_973_n 0.00557448f $X=7.28 $Y=1.675 $X2=0 $Y2=0
cc_516 N_S0_c_578_n N_A2_c_973_n 0.00374657f $X=6.495 $Y=1.675 $X2=0 $Y2=0
cc_517 N_S0_c_575_n N_A2_c_974_n 0.00906983f $X=6.325 $Y=1.36 $X2=0 $Y2=0
cc_518 N_S0_c_576_n N_A2_c_974_n 0.00424705f $X=6.41 $Y=1.59 $X2=0 $Y2=0
cc_519 N_S0_c_577_n N_A2_c_974_n 0.00133605f $X=7.28 $Y=1.675 $X2=0 $Y2=0
cc_520 N_S0_c_578_n N_A2_c_974_n 9.04512e-19 $X=6.495 $Y=1.675 $X2=0 $Y2=0
cc_521 N_S0_c_583_n N_A2_c_974_n 0.00107882f $X=5.98 $Y=1.36 $X2=0 $Y2=0
cc_522 N_S0_c_584_n N_A2_c_974_n 0.0206524f $X=5.98 $Y=1.595 $X2=0 $Y2=0
cc_523 N_S0_c_574_n A2 0.00323948f $X=5.815 $Y=1.36 $X2=0 $Y2=0
cc_524 N_S0_c_582_n A2 0.00352108f $X=5.565 $Y=1.245 $X2=0 $Y2=0
cc_525 N_S0_c_583_n A2 0.0211332f $X=5.98 $Y=1.36 $X2=0 $Y2=0
cc_526 N_S0_c_584_n A2 2.80518e-19 $X=5.98 $Y=1.595 $X2=0 $Y2=0
cc_527 N_S0_c_574_n N_A2_c_976_n 7.8466e-19 $X=5.815 $Y=1.36 $X2=0 $Y2=0
cc_528 N_S0_c_583_n N_A2_c_976_n 0.00365775f $X=5.98 $Y=1.36 $X2=0 $Y2=0
cc_529 N_S0_c_584_n N_A2_c_976_n 0.0119133f $X=5.98 $Y=1.595 $X2=0 $Y2=0
cc_530 N_S0_c_577_n N_A1_c_1026_n 0.010068f $X=7.28 $Y=1.675 $X2=0 $Y2=0
cc_531 N_S0_c_614_p N_A1_c_1026_n 0.00112992f $X=7.525 $Y=2.545 $X2=0 $Y2=0
cc_532 N_S0_c_614_p N_A1_M1010_g 6.16357e-19 $X=7.525 $Y=2.545 $X2=0 $Y2=0
cc_533 N_S0_M1019_g N_A1_M1018_g 0.0533184f $X=7.385 $Y=0.445 $X2=0 $Y2=0
cc_534 N_S0_c_576_n N_A1_c_1028_n 8.13086e-19 $X=6.41 $Y=1.59 $X2=0 $Y2=0
cc_535 N_S0_c_577_n N_A1_c_1028_n 0.00516357f $X=7.28 $Y=1.675 $X2=0 $Y2=0
cc_536 N_S0_c_579_n N_A1_c_1028_n 0.00632616f $X=7.445 $Y=1.245 $X2=0 $Y2=0
cc_537 N_S0_c_575_n A1 0.00761148f $X=6.325 $Y=1.36 $X2=0 $Y2=0
cc_538 N_S0_c_577_n A1 0.0235706f $X=7.28 $Y=1.675 $X2=0 $Y2=0
cc_539 N_S0_c_579_n A1 0.0226851f $X=7.445 $Y=1.245 $X2=0 $Y2=0
cc_540 N_S0_c_580_n A1 0.00187622f $X=7.445 $Y=1.245 $X2=0 $Y2=0
cc_541 N_S0_c_577_n N_A1_c_1030_n 0.00393012f $X=7.28 $Y=1.675 $X2=0 $Y2=0
cc_542 N_S0_c_579_n N_A1_c_1030_n 4.09747e-19 $X=7.445 $Y=1.245 $X2=0 $Y2=0
cc_543 N_S0_c_580_n N_A1_c_1030_n 0.0207636f $X=7.445 $Y=1.245 $X2=0 $Y2=0
cc_544 N_S0_c_570_n N_A0_M1000_g 0.0187334f $X=9.225 $Y=0.73 $X2=0 $Y2=0
cc_545 N_S0_c_590_n N_A0_M1000_g 0.00875429f $X=9.455 $Y=1.605 $X2=0 $Y2=0
cc_546 N_S0_M1004_g N_A0_M1021_g 0.0557853f $X=8.335 $Y=2.595 $X2=0 $Y2=0
cc_547 N_S0_c_651_p N_A0_M1021_g 0.00115747f $X=8.265 $Y=2.545 $X2=0 $Y2=0
cc_548 N_S0_c_587_n N_A0_M1021_g 0.0184684f $X=8.345 $Y=1.77 $X2=0 $Y2=0
cc_549 N_S0_c_589_n N_A0_M1021_g 0.0311122f $X=9.455 $Y=1.77 $X2=0 $Y2=0
cc_550 N_S0_c_590_n N_A0_M1021_g 0.0608138f $X=9.455 $Y=1.605 $X2=0 $Y2=0
cc_551 N_S0_c_572_n A0 8.69706e-19 $X=9.585 $Y=0.805 $X2=0 $Y2=0
cc_552 N_S0_c_596_n A0 0.00511548f $X=8.265 $Y=2.15 $X2=0 $Y2=0
cc_553 N_S0_c_587_n A0 0.00296311f $X=8.345 $Y=1.77 $X2=0 $Y2=0
cc_554 N_S0_c_588_n A0 9.62038e-19 $X=9.455 $Y=1.77 $X2=0 $Y2=0
cc_555 N_S0_c_589_n A0 0.0866049f $X=9.455 $Y=1.77 $X2=0 $Y2=0
cc_556 N_S0_c_590_n A0 0.0139602f $X=9.455 $Y=1.605 $X2=0 $Y2=0
cc_557 N_S0_c_589_n N_A0_c_1072_n 0.00204657f $X=9.455 $Y=1.77 $X2=0 $Y2=0
cc_558 N_S0_c_590_n N_A0_c_1072_n 0.0186787f $X=9.455 $Y=1.605 $X2=0 $Y2=0
cc_559 N_S0_c_589_n N_VPWR_M1021_d 0.00198707f $X=9.455 $Y=1.77 $X2=0 $Y2=0
cc_560 N_S0_M1008_g N_VPWR_c_1129_n 0.00427944f $X=5.925 $Y=2.595 $X2=0 $Y2=0
cc_561 N_S0_M1004_g N_VPWR_c_1130_n 0.00110534f $X=8.335 $Y=2.595 $X2=0 $Y2=0
cc_562 N_S0_M1028_g N_VPWR_c_1130_n 0.0135263f $X=9.415 $Y=2.595 $X2=0 $Y2=0
cc_563 N_S0_M1008_g N_VPWR_c_1131_n 0.00975641f $X=5.925 $Y=2.595 $X2=0 $Y2=0
cc_564 N_S0_M1004_g N_VPWR_c_1133_n 0.00599941f $X=8.335 $Y=2.595 $X2=0 $Y2=0
cc_565 N_S0_M1028_g N_VPWR_c_1136_n 0.00840199f $X=9.415 $Y=2.595 $X2=0 $Y2=0
cc_566 N_S0_M1008_g N_VPWR_c_1126_n 0.0186811f $X=5.925 $Y=2.595 $X2=0 $Y2=0
cc_567 N_S0_M1004_g N_VPWR_c_1126_n 0.00855775f $X=8.335 $Y=2.595 $X2=0 $Y2=0
cc_568 N_S0_M1028_g N_VPWR_c_1126_n 0.0085752f $X=9.415 $Y=2.595 $X2=0 $Y2=0
cc_569 N_S0_c_573_n N_A_245_411#_c_1228_n 0.00242817f $X=5.035 $Y=1.21 $X2=0
+ $Y2=0
cc_570 N_S0_c_581_n N_A_245_411#_c_1228_n 0.0250964f $X=5.395 $Y=1.245 $X2=0
+ $Y2=0
cc_571 N_S0_c_586_n N_A_245_411#_c_1228_n 0.00367136f $X=5.035 $Y=1.045 $X2=0
+ $Y2=0
cc_572 N_S0_c_573_n N_A_245_411#_c_1229_n 0.00323185f $X=5.035 $Y=1.21 $X2=0
+ $Y2=0
cc_573 N_S0_c_581_n N_A_245_411#_c_1229_n 0.0317809f $X=5.395 $Y=1.245 $X2=0
+ $Y2=0
cc_574 N_S0_c_586_n N_A_245_411#_c_1229_n 0.0109865f $X=5.035 $Y=1.045 $X2=0
+ $Y2=0
cc_575 N_S0_M1008_g N_A_245_411#_c_1238_n 0.011059f $X=5.925 $Y=2.595 $X2=0
+ $Y2=0
cc_576 N_S0_M1008_g N_A_245_411#_c_1292_n 0.0154787f $X=5.925 $Y=2.595 $X2=0
+ $Y2=0
cc_577 N_S0_c_615_p N_A_470_57#_M1023_d 0.0186609f $X=8.18 $Y=2.63 $X2=0 $Y2=0
cc_578 N_S0_c_581_n N_A_470_57#_c_1376_n 0.00479602f $X=5.395 $Y=1.245 $X2=0
+ $Y2=0
cc_579 N_S0_c_586_n N_A_470_57#_c_1376_n 0.00703101f $X=5.035 $Y=1.045 $X2=0
+ $Y2=0
cc_580 N_S0_M1019_g N_A_470_57#_c_1379_n 0.012536f $X=7.385 $Y=0.445 $X2=0 $Y2=0
cc_581 N_S0_c_575_n N_A_470_57#_c_1379_n 0.0025498f $X=6.325 $Y=1.36 $X2=0 $Y2=0
cc_582 N_S0_c_579_n N_A_470_57#_c_1379_n 0.0195978f $X=7.445 $Y=1.245 $X2=0
+ $Y2=0
cc_583 N_S0_c_580_n N_A_470_57#_c_1379_n 7.91444e-19 $X=7.445 $Y=1.245 $X2=0
+ $Y2=0
cc_584 N_S0_c_575_n N_A_470_57#_c_1380_n 0.00826197f $X=6.325 $Y=1.36 $X2=0
+ $Y2=0
cc_585 N_S0_M1019_g N_A_470_57#_c_1381_n 0.0132855f $X=7.385 $Y=0.445 $X2=0
+ $Y2=0
cc_586 N_S0_M1019_g N_A_470_57#_c_1382_n 0.00318133f $X=7.385 $Y=0.445 $X2=0
+ $Y2=0
cc_587 N_S0_M1004_g N_A_470_57#_c_1382_n 0.00157734f $X=8.335 $Y=2.595 $X2=0
+ $Y2=0
cc_588 N_S0_c_579_n N_A_470_57#_c_1382_n 0.0374213f $X=7.445 $Y=1.245 $X2=0
+ $Y2=0
cc_589 N_S0_c_580_n N_A_470_57#_c_1382_n 0.00174446f $X=7.445 $Y=1.245 $X2=0
+ $Y2=0
cc_590 N_S0_c_614_p N_A_470_57#_c_1382_n 0.0408204f $X=7.525 $Y=2.545 $X2=0
+ $Y2=0
cc_591 N_S0_c_615_p N_A_470_57#_c_1382_n 0.0130962f $X=8.18 $Y=2.63 $X2=0 $Y2=0
cc_592 N_S0_c_596_n N_A_470_57#_c_1382_n 0.0315869f $X=8.265 $Y=2.15 $X2=0 $Y2=0
cc_593 N_S0_c_585_n N_A_470_57#_c_1382_n 0.012867f $X=7.445 $Y=1.675 $X2=0 $Y2=0
cc_594 N_S0_c_587_n N_A_470_57#_c_1382_n 9.67698e-19 $X=8.345 $Y=1.77 $X2=0
+ $Y2=0
cc_595 N_S0_c_579_n N_A_470_57#_c_1384_n 0.00543421f $X=7.445 $Y=1.245 $X2=0
+ $Y2=0
cc_596 N_S0_c_580_n N_A_470_57#_c_1384_n 4.97199e-19 $X=7.445 $Y=1.245 $X2=0
+ $Y2=0
cc_597 N_S0_c_589_n A_1692_419# 0.00579363f $X=9.455 $Y=1.77 $X2=-0.19
+ $Y2=-0.245
cc_598 N_S0_c_570_n N_VGND_c_1553_n 0.0127929f $X=9.225 $Y=0.73 $X2=0 $Y2=0
cc_599 N_S0_c_571_n N_VGND_c_1553_n 0.00239794f $X=9.585 $Y=0.73 $X2=0 $Y2=0
cc_600 N_S0_c_586_n N_VGND_c_1556_n 7.10185e-19 $X=5.035 $Y=1.045 $X2=0 $Y2=0
cc_601 N_S0_M1019_g N_VGND_c_1559_n 0.00438531f $X=7.385 $Y=0.445 $X2=0 $Y2=0
cc_602 N_S0_c_570_n N_VGND_c_1560_n 0.00486043f $X=9.225 $Y=0.73 $X2=0 $Y2=0
cc_603 N_S0_c_571_n N_VGND_c_1560_n 0.00549284f $X=9.585 $Y=0.73 $X2=0 $Y2=0
cc_604 N_S0_c_572_n N_VGND_c_1560_n 6.21075e-19 $X=9.585 $Y=0.805 $X2=0 $Y2=0
cc_605 N_S0_M1019_g N_VGND_c_1561_n 0.00646541f $X=7.385 $Y=0.445 $X2=0 $Y2=0
cc_606 N_S0_c_570_n N_VGND_c_1561_n 0.00445031f $X=9.225 $Y=0.73 $X2=0 $Y2=0
cc_607 N_S0_c_571_n N_VGND_c_1561_n 0.00719421f $X=9.585 $Y=0.73 $X2=0 $Y2=0
cc_608 N_S0_c_572_n N_VGND_c_1561_n 8.18184e-19 $X=9.585 $Y=0.805 $X2=0 $Y2=0
cc_609 N_A_946_317#_c_800_n N_A2_M1009_g 0.0220755f $X=7.09 $Y=2.025 $X2=0 $Y2=0
cc_610 N_A_946_317#_c_841_n N_A2_M1009_g 9.65029e-19 $X=7.175 $Y=2.895 $X2=0
+ $Y2=0
cc_611 N_A_946_317#_M1011_g A2 0.00162537f $X=5.485 $Y=0.445 $X2=0 $Y2=0
cc_612 N_A_946_317#_M1011_g N_A2_c_976_n 0.0199393f $X=5.485 $Y=0.445 $X2=0
+ $Y2=0
cc_613 N_A_946_317#_M1011_g N_A2_c_977_n 0.0374235f $X=5.485 $Y=0.445 $X2=0
+ $Y2=0
cc_614 N_A_946_317#_c_782_n N_A1_c_1026_n 0.0422137f $X=7.655 $Y=1.725 $X2=0
+ $Y2=0
cc_615 N_A_946_317#_M1023_g N_A1_M1010_g 0.0422137f $X=7.53 $Y=2.595 $X2=0 $Y2=0
cc_616 N_A_946_317#_c_800_n N_A1_M1010_g 0.0182149f $X=7.09 $Y=2.025 $X2=0 $Y2=0
cc_617 N_A_946_317#_c_841_n N_A1_M1010_g 0.0179507f $X=7.175 $Y=2.895 $X2=0
+ $Y2=0
cc_618 N_A_946_317#_c_894_p N_A1_M1010_g 0.00521921f $X=7.26 $Y=2.98 $X2=0 $Y2=0
cc_619 N_A_946_317#_c_784_n N_A0_M1000_g 0.0129437f $X=7.925 $Y=0.765 $X2=0
+ $Y2=0
cc_620 N_A_946_317#_c_786_n N_A0_M1000_g 0.012262f $X=9.635 $Y=0.945 $X2=0 $Y2=0
cc_621 N_A_946_317#_c_790_n N_A0_M1000_g 0.0176003f $X=8.305 $Y=0.93 $X2=0 $Y2=0
cc_622 N_A_946_317#_c_791_n N_A0_M1000_g 6.05143e-19 $X=8.47 $Y=0.897 $X2=0
+ $Y2=0
cc_623 N_A_946_317#_c_843_n N_A0_M1021_g 0.00584552f $X=8.635 $Y=2.98 $X2=0
+ $Y2=0
cc_624 N_A_946_317#_c_850_n N_A0_M1021_g 0.0104295f $X=8.72 $Y=2.895 $X2=0 $Y2=0
cc_625 N_A_946_317#_c_854_n N_A0_M1021_g 0.0123294f $X=9.515 $Y=2.415 $X2=0
+ $Y2=0
cc_626 N_A_946_317#_c_856_n N_A0_M1021_g 0.00284897f $X=8.805 $Y=2.415 $X2=0
+ $Y2=0
cc_627 N_A_946_317#_c_804_n N_A0_M1021_g 8.69744e-19 $X=9.68 $Y=2.495 $X2=0
+ $Y2=0
cc_628 N_A_946_317#_c_783_n A0 0.00462818f $X=7.895 $Y=1.65 $X2=0 $Y2=0
cc_629 N_A_946_317#_c_788_n A0 0.0133435f $X=9.885 $Y=2.33 $X2=0 $Y2=0
cc_630 N_A_946_317#_c_790_n A0 0.00189482f $X=8.305 $Y=0.93 $X2=0 $Y2=0
cc_631 N_A_946_317#_c_791_n A0 0.0852851f $X=8.47 $Y=0.897 $X2=0 $Y2=0
cc_632 N_A_946_317#_c_786_n N_A0_c_1072_n 0.00473222f $X=9.635 $Y=0.945 $X2=0
+ $Y2=0
cc_633 N_A_946_317#_c_800_n N_VPWR_M1009_d 0.00213411f $X=7.09 $Y=2.025 $X2=0
+ $Y2=0
cc_634 N_A_946_317#_c_854_n N_VPWR_M1021_d 0.00380882f $X=9.515 $Y=2.415 $X2=0
+ $Y2=0
cc_635 N_A_946_317#_c_800_n N_VPWR_c_1129_n 0.0169845f $X=7.09 $Y=2.025 $X2=0
+ $Y2=0
cc_636 N_A_946_317#_c_843_n N_VPWR_c_1130_n 0.0129587f $X=8.635 $Y=2.98 $X2=0
+ $Y2=0
cc_637 N_A_946_317#_c_850_n N_VPWR_c_1130_n 0.0146335f $X=8.72 $Y=2.895 $X2=0
+ $Y2=0
cc_638 N_A_946_317#_c_854_n N_VPWR_c_1130_n 0.0160419f $X=9.515 $Y=2.415 $X2=0
+ $Y2=0
cc_639 N_A_946_317#_c_804_n N_VPWR_c_1130_n 0.0260067f $X=9.68 $Y=2.495 $X2=0
+ $Y2=0
cc_640 N_A_946_317#_M1015_g N_VPWR_c_1131_n 0.00701311f $X=4.855 $Y=2.595 $X2=0
+ $Y2=0
cc_641 N_A_946_317#_M1023_g N_VPWR_c_1133_n 0.00599941f $X=7.53 $Y=2.595 $X2=0
+ $Y2=0
cc_642 N_A_946_317#_c_843_n N_VPWR_c_1133_n 0.0842305f $X=8.635 $Y=2.98 $X2=0
+ $Y2=0
cc_643 N_A_946_317#_c_894_p N_VPWR_c_1133_n 0.00921717f $X=7.26 $Y=2.98 $X2=0
+ $Y2=0
cc_644 N_A_946_317#_c_804_n N_VPWR_c_1136_n 0.0281861f $X=9.68 $Y=2.495 $X2=0
+ $Y2=0
cc_645 N_A_946_317#_M1028_d N_VPWR_c_1126_n 0.0023218f $X=9.54 $Y=2.095 $X2=0
+ $Y2=0
cc_646 N_A_946_317#_M1015_g N_VPWR_c_1126_n 0.0100017f $X=4.855 $Y=2.595 $X2=0
+ $Y2=0
cc_647 N_A_946_317#_M1023_g N_VPWR_c_1126_n 0.00842247f $X=7.53 $Y=2.595 $X2=0
+ $Y2=0
cc_648 N_A_946_317#_c_843_n N_VPWR_c_1126_n 0.0554116f $X=8.635 $Y=2.98 $X2=0
+ $Y2=0
cc_649 N_A_946_317#_c_894_p N_VPWR_c_1126_n 0.00623238f $X=7.26 $Y=2.98 $X2=0
+ $Y2=0
cc_650 N_A_946_317#_c_854_n N_VPWR_c_1126_n 0.0116288f $X=9.515 $Y=2.415 $X2=0
+ $Y2=0
cc_651 N_A_946_317#_c_804_n N_VPWR_c_1126_n 0.0173447f $X=9.68 $Y=2.495 $X2=0
+ $Y2=0
cc_652 N_A_946_317#_c_800_n N_A_245_411#_M1015_d 0.00415987f $X=7.09 $Y=2.025
+ $X2=0 $Y2=0
cc_653 N_A_946_317#_c_803_n N_A_245_411#_M1015_d 0.00734059f $X=5.55 $Y=1.83
+ $X2=0 $Y2=0
cc_654 N_A_946_317#_c_789_n N_A_245_411#_c_1228_n 0.0237518f $X=5.05 $Y=1.75
+ $X2=0 $Y2=0
cc_655 N_A_946_317#_c_793_n N_A_245_411#_c_1228_n 0.00905561f $X=5.215 $Y=1.75
+ $X2=0 $Y2=0
cc_656 N_A_946_317#_M1011_g N_A_245_411#_c_1229_n 0.00514465f $X=5.485 $Y=0.445
+ $X2=0 $Y2=0
cc_657 N_A_946_317#_M1015_g N_A_245_411#_c_1306_n 0.0192072f $X=4.855 $Y=2.595
+ $X2=0 $Y2=0
cc_658 N_A_946_317#_c_789_n N_A_245_411#_c_1306_n 0.00172794f $X=5.05 $Y=1.75
+ $X2=0 $Y2=0
cc_659 N_A_946_317#_M1015_g N_A_245_411#_c_1238_n 0.00748675f $X=4.855 $Y=2.595
+ $X2=0 $Y2=0
cc_660 N_A_946_317#_c_799_n N_A_245_411#_c_1238_n 0.00547233f $X=5.465 $Y=1.83
+ $X2=0 $Y2=0
cc_661 N_A_946_317#_c_789_n N_A_245_411#_c_1238_n 0.0179112f $X=5.05 $Y=1.75
+ $X2=0 $Y2=0
cc_662 N_A_946_317#_c_803_n N_A_245_411#_c_1238_n 0.00109864f $X=5.55 $Y=1.83
+ $X2=0 $Y2=0
cc_663 N_A_946_317#_c_793_n N_A_245_411#_c_1238_n 0.00165966f $X=5.215 $Y=1.75
+ $X2=0 $Y2=0
cc_664 N_A_946_317#_M1015_g N_A_245_411#_c_1292_n 0.0118765f $X=4.855 $Y=2.595
+ $X2=0 $Y2=0
cc_665 N_A_946_317#_c_843_n N_A_470_57#_M1023_d 0.0108596f $X=8.635 $Y=2.98
+ $X2=0 $Y2=0
cc_666 N_A_946_317#_M1011_g N_A_470_57#_c_1376_n 0.0130367f $X=5.485 $Y=0.445
+ $X2=0 $Y2=0
cc_667 N_A_946_317#_c_784_n N_A_470_57#_c_1381_n 0.025843f $X=7.925 $Y=0.765
+ $X2=0 $Y2=0
cc_668 N_A_946_317#_M1023_g N_A_470_57#_c_1382_n 0.00540411f $X=7.53 $Y=2.595
+ $X2=0 $Y2=0
cc_669 N_A_946_317#_c_781_n N_A_470_57#_c_1382_n 0.00976008f $X=7.82 $Y=1.725
+ $X2=0 $Y2=0
cc_670 N_A_946_317#_c_783_n N_A_470_57#_c_1382_n 0.0236546f $X=7.895 $Y=1.65
+ $X2=0 $Y2=0
cc_671 N_A_946_317#_c_785_n N_A_470_57#_c_1382_n 0.00878829f $X=7.82 $Y=0.945
+ $X2=0 $Y2=0
cc_672 N_A_946_317#_c_791_n N_A_470_57#_c_1382_n 0.00935127f $X=8.47 $Y=0.897
+ $X2=0 $Y2=0
cc_673 N_A_946_317#_c_784_n N_A_470_57#_c_1384_n 0.00234501f $X=7.925 $Y=0.765
+ $X2=0 $Y2=0
cc_674 N_A_946_317#_c_785_n N_A_470_57#_c_1384_n 0.00547038f $X=7.82 $Y=0.945
+ $X2=0 $Y2=0
cc_675 N_A_946_317#_c_791_n N_A_470_57#_c_1384_n 0.0104333f $X=8.47 $Y=0.897
+ $X2=0 $Y2=0
cc_676 N_A_946_317#_c_800_n A_1210_419# 0.00728771f $X=7.09 $Y=2.025 $X2=-0.19
+ $Y2=-0.245
cc_677 N_A_946_317#_c_841_n A_1433_419# 0.00716453f $X=7.175 $Y=2.895 $X2=-0.19
+ $Y2=-0.245
cc_678 N_A_946_317#_c_843_n A_1433_419# 0.00415466f $X=8.635 $Y=2.98 $X2=-0.19
+ $Y2=-0.245
cc_679 N_A_946_317#_c_894_p A_1433_419# 3.79893e-19 $X=7.26 $Y=2.98 $X2=-0.19
+ $Y2=-0.245
cc_680 N_A_946_317#_c_843_n A_1692_419# 0.00616714f $X=8.635 $Y=2.98 $X2=-0.19
+ $Y2=-0.245
cc_681 N_A_946_317#_c_850_n A_1692_419# 0.00429116f $X=8.72 $Y=2.895 $X2=-0.19
+ $Y2=-0.245
cc_682 N_A_946_317#_c_856_n A_1692_419# 0.00249153f $X=8.805 $Y=2.415 $X2=-0.19
+ $Y2=-0.245
cc_683 N_A_946_317#_c_786_n N_VGND_c_1553_n 0.0250214f $X=9.635 $Y=0.945 $X2=0
+ $Y2=0
cc_684 N_A_946_317#_c_787_n N_VGND_c_1553_n 0.0137333f $X=9.8 $Y=0.47 $X2=0
+ $Y2=0
cc_685 N_A_946_317#_M1011_g N_VGND_c_1556_n 0.00359964f $X=5.485 $Y=0.445 $X2=0
+ $Y2=0
cc_686 N_A_946_317#_c_784_n N_VGND_c_1559_n 0.00421428f $X=7.925 $Y=0.765 $X2=0
+ $Y2=0
cc_687 N_A_946_317#_c_790_n N_VGND_c_1559_n 0.00822282f $X=8.305 $Y=0.93 $X2=0
+ $Y2=0
cc_688 N_A_946_317#_c_787_n N_VGND_c_1560_n 0.0201256f $X=9.8 $Y=0.47 $X2=0
+ $Y2=0
cc_689 N_A_946_317#_M1020_d N_VGND_c_1561_n 0.00232985f $X=9.66 $Y=0.235 $X2=0
+ $Y2=0
cc_690 N_A_946_317#_M1011_g N_VGND_c_1561_n 0.00674206f $X=5.485 $Y=0.445 $X2=0
+ $Y2=0
cc_691 N_A_946_317#_c_784_n N_VGND_c_1561_n 0.0080497f $X=7.925 $Y=0.765 $X2=0
+ $Y2=0
cc_692 N_A_946_317#_c_786_n N_VGND_c_1561_n 0.0260467f $X=9.635 $Y=0.945 $X2=0
+ $Y2=0
cc_693 N_A_946_317#_c_787_n N_VGND_c_1561_n 0.0127743f $X=9.8 $Y=0.47 $X2=0
+ $Y2=0
cc_694 N_A_946_317#_c_790_n N_VGND_c_1561_n 0.0111244f $X=8.305 $Y=0.93 $X2=0
+ $Y2=0
cc_695 N_A_946_317#_c_791_n N_VGND_c_1561_n 0.0114918f $X=8.47 $Y=0.897 $X2=0
+ $Y2=0
cc_696 N_A2_c_973_n N_A1_c_1026_n 0.0180877f $X=6.48 $Y=1.775 $X2=0 $Y2=0
cc_697 N_A2_M1009_g N_A1_M1010_g 0.0180877f $X=6.48 $Y=2.595 $X2=0 $Y2=0
cc_698 N_A2_c_972_n N_A1_M1018_g 0.00542612f $X=6.355 $Y=1.02 $X2=0 $Y2=0
cc_699 N_A2_c_974_n N_A1_c_1028_n 0.00696886f $X=6.48 $Y=1.65 $X2=0 $Y2=0
cc_700 N_A2_c_972_n A1 0.00167239f $X=6.355 $Y=1.02 $X2=0 $Y2=0
cc_701 A2 A1 3.16546e-19 $X=5.915 $Y=0.84 $X2=0 $Y2=0
cc_702 N_A2_c_972_n N_A1_c_1030_n 0.017187f $X=6.355 $Y=1.02 $X2=0 $Y2=0
cc_703 N_A2_M1009_g N_VPWR_c_1129_n 0.0230465f $X=6.48 $Y=2.595 $X2=0 $Y2=0
cc_704 N_A2_M1009_g N_VPWR_c_1131_n 0.008763f $X=6.48 $Y=2.595 $X2=0 $Y2=0
cc_705 N_A2_M1009_g N_VPWR_c_1126_n 0.0146299f $X=6.48 $Y=2.595 $X2=0 $Y2=0
cc_706 A2 N_A_245_411#_c_1229_n 0.00423536f $X=5.915 $Y=0.84 $X2=0 $Y2=0
cc_707 N_A2_c_972_n N_A_470_57#_c_1376_n 0.00393242f $X=6.355 $Y=1.02 $X2=0
+ $Y2=0
cc_708 A2 N_A_470_57#_c_1376_n 0.00997911f $X=5.915 $Y=0.84 $X2=0 $Y2=0
cc_709 N_A2_c_976_n N_A_470_57#_c_1376_n 0.00300828f $X=5.935 $Y=0.93 $X2=0
+ $Y2=0
cc_710 N_A2_c_977_n N_A_470_57#_c_1376_n 0.0121502f $X=5.935 $Y=0.765 $X2=0
+ $Y2=0
cc_711 N_A2_c_977_n N_A_470_57#_c_1378_n 0.00862241f $X=5.935 $Y=0.765 $X2=0
+ $Y2=0
cc_712 N_A2_c_972_n N_A_470_57#_c_1379_n 0.00247306f $X=6.355 $Y=1.02 $X2=0
+ $Y2=0
cc_713 N_A2_c_972_n N_A_470_57#_c_1380_n 0.00525342f $X=6.355 $Y=1.02 $X2=0
+ $Y2=0
cc_714 A2 N_A_470_57#_c_1380_n 0.01084f $X=5.915 $Y=0.84 $X2=0 $Y2=0
cc_715 N_A2_c_976_n N_A_470_57#_c_1380_n 0.0032053f $X=5.935 $Y=0.93 $X2=0 $Y2=0
cc_716 N_A2_c_977_n N_A_470_57#_c_1380_n 0.00121802f $X=5.935 $Y=0.765 $X2=0
+ $Y2=0
cc_717 N_A2_c_977_n N_VGND_c_1552_n 0.00267147f $X=5.935 $Y=0.765 $X2=0 $Y2=0
cc_718 N_A2_c_977_n N_VGND_c_1556_n 0.00359964f $X=5.935 $Y=0.765 $X2=0 $Y2=0
cc_719 N_A2_c_977_n N_VGND_c_1561_n 0.00674206f $X=5.935 $Y=0.765 $X2=0 $Y2=0
cc_720 N_A1_M1010_g N_VPWR_c_1129_n 0.00389552f $X=7.04 $Y=2.595 $X2=0 $Y2=0
cc_721 N_A1_M1010_g N_VPWR_c_1133_n 0.00862827f $X=7.04 $Y=2.595 $X2=0 $Y2=0
cc_722 N_A1_M1010_g N_VPWR_c_1126_n 0.0140404f $X=7.04 $Y=2.595 $X2=0 $Y2=0
cc_723 N_A1_M1018_g N_A_470_57#_c_1378_n 0.00456175f $X=6.995 $Y=0.445 $X2=0
+ $Y2=0
cc_724 N_A1_M1018_g N_A_470_57#_c_1379_n 0.0139773f $X=6.995 $Y=0.445 $X2=0
+ $Y2=0
cc_725 A1 N_A_470_57#_c_1379_n 0.0235707f $X=6.875 $Y=1.21 $X2=0 $Y2=0
cc_726 N_A1_c_1030_n N_A_470_57#_c_1379_n 0.00402927f $X=6.905 $Y=1.245 $X2=0
+ $Y2=0
cc_727 N_A1_M1018_g N_VGND_c_1552_n 0.0105069f $X=6.995 $Y=0.445 $X2=0 $Y2=0
cc_728 N_A1_M1018_g N_VGND_c_1559_n 0.00438531f $X=6.995 $Y=0.445 $X2=0 $Y2=0
cc_729 N_A1_M1018_g N_VGND_c_1561_n 0.00745669f $X=6.995 $Y=0.445 $X2=0 $Y2=0
cc_730 N_A0_M1021_g N_VPWR_c_1130_n 0.0116219f $X=8.875 $Y=2.595 $X2=0 $Y2=0
cc_731 N_A0_M1021_g N_VPWR_c_1133_n 0.00832595f $X=8.875 $Y=2.595 $X2=0 $Y2=0
cc_732 N_A0_M1021_g N_VPWR_c_1126_n 0.00777522f $X=8.875 $Y=2.595 $X2=0 $Y2=0
cc_733 A0 N_A_470_57#_c_1382_n 0.0123807f $X=9.275 $Y=1.21 $X2=0 $Y2=0
cc_734 N_A0_M1000_g N_VGND_c_1553_n 0.0245566f $X=8.795 $Y=0.445 $X2=0 $Y2=0
cc_735 N_A0_M1000_g N_VGND_c_1559_n 0.00486043f $X=8.795 $Y=0.445 $X2=0 $Y2=0
cc_736 N_A0_M1000_g N_VGND_c_1561_n 0.0054803f $X=8.795 $Y=0.445 $X2=0 $Y2=0
cc_737 X N_VPWR_c_1127_n 0.0484297f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_738 X N_VPWR_c_1126_n 0.0125808f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_739 X N_VPWR_c_1138_n 0.0220321f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_740 X N_A_245_411#_c_1224_n 0.0804059f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_741 X N_A_245_411#_c_1226_n 0.0132378f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_742 X N_A_245_411#_c_1253_n 0.0129587f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_743 X N_VGND_c_1550_n 0.00669147f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_744 X N_VGND_c_1558_n 0.0197885f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_745 N_X_M1006_s N_VGND_c_1561_n 0.00232985f $X=0.135 $Y=0.235 $X2=0 $Y2=0
cc_746 X N_VGND_c_1561_n 0.0125808f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_747 N_VPWR_c_1126_n N_A_245_411#_M1015_d 0.024694f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_748 N_VPWR_M1005_d N_A_245_411#_c_1231_n 0.00233567f $X=0.67 $Y=2.045 $X2=0
+ $Y2=0
cc_749 N_VPWR_c_1127_n N_A_245_411#_c_1231_n 0.0139786f $X=0.81 $Y=2.495 $X2=0
+ $Y2=0
cc_750 N_VPWR_M1005_d N_A_245_411#_c_1253_n 7.70949e-19 $X=0.67 $Y=2.045 $X2=0
+ $Y2=0
cc_751 N_VPWR_c_1127_n N_A_245_411#_c_1253_n 0.00777198f $X=0.81 $Y=2.495 $X2=0
+ $Y2=0
cc_752 N_VPWR_c_1127_n N_A_245_411#_c_1232_n 0.0121618f $X=0.81 $Y=2.495 $X2=0
+ $Y2=0
cc_753 N_VPWR_c_1135_n N_A_245_411#_c_1232_n 0.0168561f $X=3.855 $Y=3.33 $X2=0
+ $Y2=0
cc_754 N_VPWR_c_1126_n N_A_245_411#_c_1232_n 0.00967329f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_755 N_VPWR_c_1127_n N_A_245_411#_c_1233_n 0.0372755f $X=0.81 $Y=2.495 $X2=0
+ $Y2=0
cc_756 N_VPWR_c_1135_n N_A_245_411#_c_1234_n 0.110317f $X=3.855 $Y=3.33 $X2=0
+ $Y2=0
cc_757 N_VPWR_c_1126_n N_A_245_411#_c_1234_n 0.0662824f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_758 N_VPWR_M1022_d N_A_245_411#_c_1276_n 0.0113828f $X=3.8 $Y=2.095 $X2=0
+ $Y2=0
cc_759 N_VPWR_c_1128_n N_A_245_411#_c_1276_n 0.0236971f $X=4.02 $Y=3.03 $X2=0
+ $Y2=0
cc_760 N_VPWR_c_1131_n N_A_245_411#_c_1276_n 0.00493296f $X=6.58 $Y=3.33 $X2=0
+ $Y2=0
cc_761 N_VPWR_c_1135_n N_A_245_411#_c_1276_n 0.00859354f $X=3.855 $Y=3.33 $X2=0
+ $Y2=0
cc_762 N_VPWR_c_1126_n N_A_245_411#_c_1276_n 0.0250386f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_763 N_VPWR_c_1131_n N_A_245_411#_c_1306_n 0.00382225f $X=6.58 $Y=3.33 $X2=0
+ $Y2=0
cc_764 N_VPWR_c_1126_n N_A_245_411#_c_1306_n 0.00595176f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_765 N_VPWR_c_1131_n N_A_245_411#_c_1336_n 0.00279764f $X=6.58 $Y=3.33 $X2=0
+ $Y2=0
cc_766 N_VPWR_c_1126_n N_A_245_411#_c_1336_n 0.00510631f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_767 N_VPWR_c_1131_n N_A_245_411#_c_1292_n 0.0197322f $X=6.58 $Y=3.33 $X2=0
+ $Y2=0
cc_768 N_VPWR_c_1126_n N_A_245_411#_c_1292_n 0.012508f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_769 N_VPWR_c_1126_n N_A_470_57#_M1023_d 0.00453461f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_770 N_VPWR_c_1126_n A_898_419# 0.00282312f $X=9.84 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_771 N_VPWR_c_1126_n A_1210_419# 0.0130629f $X=9.84 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_772 N_VPWR_c_1126_n A_1433_419# 0.00193244f $X=9.84 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_773 N_VPWR_c_1126_n A_1692_419# 0.00233503f $X=9.84 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_774 N_A_245_411#_c_1234_n N_A_470_57#_M1001_d 0.00596193f $X=3.115 $Y=2.98
+ $X2=0 $Y2=0
cc_775 N_A_245_411#_c_1234_n N_A_470_57#_c_1385_n 0.0177763f $X=3.115 $Y=2.98
+ $X2=0 $Y2=0
cc_776 N_A_245_411#_c_1235_n N_A_470_57#_c_1385_n 0.00219908f $X=3.2 $Y=2.895
+ $X2=0 $Y2=0
cc_777 N_A_245_411#_c_1236_n N_A_470_57#_c_1385_n 0.01416f $X=3.285 $Y=2.6 $X2=0
+ $Y2=0
cc_778 N_A_245_411#_c_1234_n N_A_470_57#_c_1386_n 0.00589553f $X=3.115 $Y=2.98
+ $X2=0 $Y2=0
cc_779 N_A_245_411#_c_1276_n N_A_470_57#_c_1386_n 0.0296113f $X=4.535 $Y=2.6
+ $X2=0 $Y2=0
cc_780 N_A_245_411#_c_1236_n N_A_470_57#_c_1386_n 0.013241f $X=3.285 $Y=2.6
+ $X2=0 $Y2=0
cc_781 N_A_245_411#_c_1228_n N_A_470_57#_c_1373_n 0.0128712f $X=4.62 $Y=2.515
+ $X2=0 $Y2=0
cc_782 N_A_245_411#_c_1228_n N_A_470_57#_c_1375_n 0.0171644f $X=4.62 $Y=2.515
+ $X2=0 $Y2=0
cc_783 N_A_245_411#_c_1291_n N_A_470_57#_c_1375_n 0.0187932f $X=4.705 $Y=0.74
+ $X2=0 $Y2=0
cc_784 N_A_245_411#_M1003_d N_A_470_57#_c_1376_n 0.00392215f $X=5.05 $Y=0.505
+ $X2=0 $Y2=0
cc_785 N_A_245_411#_c_1291_n N_A_470_57#_c_1376_n 0.0101805f $X=4.705 $Y=0.74
+ $X2=0 $Y2=0
cc_786 N_A_245_411#_c_1229_n N_A_470_57#_c_1376_n 0.0394408f $X=5.19 $Y=0.78
+ $X2=0 $Y2=0
cc_787 N_A_245_411#_c_1228_n A_898_419# 0.00168077f $X=4.62 $Y=2.515 $X2=-0.19
+ $Y2=-0.245
cc_788 N_A_245_411#_c_1336_n A_898_419# 0.00232661f $X=4.62 $Y=2.6 $X2=-0.19
+ $Y2=-0.245
cc_789 N_A_245_411#_c_1226_n A_114_47# 0.00177266f $X=0.795 $Y=0.73 $X2=-0.19
+ $Y2=-0.245
cc_790 N_A_245_411#_c_1225_n N_VGND_M1026_d 0.00238807f $X=1.465 $Y=0.73
+ $X2=-0.19 $Y2=-0.245
cc_791 N_A_245_411#_c_1225_n N_VGND_c_1550_n 0.0195984f $X=1.465 $Y=0.73 $X2=0
+ $Y2=0
cc_792 N_A_245_411#_c_1227_n N_VGND_c_1550_n 0.0134837f $X=1.63 $Y=0.495 $X2=0
+ $Y2=0
cc_793 N_A_245_411#_c_1225_n N_VGND_c_1554_n 0.00408821f $X=1.465 $Y=0.73 $X2=0
+ $Y2=0
cc_794 N_A_245_411#_c_1227_n N_VGND_c_1554_n 0.0216851f $X=1.63 $Y=0.495 $X2=0
+ $Y2=0
cc_795 N_A_245_411#_c_1225_n N_VGND_c_1558_n 0.00173934f $X=1.465 $Y=0.73 $X2=0
+ $Y2=0
cc_796 N_A_245_411#_c_1226_n N_VGND_c_1558_n 0.0026378f $X=0.795 $Y=0.73 $X2=0
+ $Y2=0
cc_797 N_A_245_411#_M1003_d N_VGND_c_1561_n 0.00203662f $X=5.05 $Y=0.505 $X2=0
+ $Y2=0
cc_798 N_A_245_411#_c_1225_n N_VGND_c_1561_n 0.0106216f $X=1.465 $Y=0.73 $X2=0
+ $Y2=0
cc_799 N_A_245_411#_c_1226_n N_VGND_c_1561_n 0.00502909f $X=0.795 $Y=0.73 $X2=0
+ $Y2=0
cc_800 N_A_245_411#_c_1227_n N_VGND_c_1561_n 0.0125086f $X=1.63 $Y=0.495 $X2=0
+ $Y2=0
cc_801 N_A_245_411#_c_1228_n A_915_101# 6.96297e-19 $X=4.62 $Y=2.515 $X2=-0.19
+ $Y2=-0.245
cc_802 N_A_245_411#_c_1291_n A_915_101# 7.93133e-19 $X=4.705 $Y=0.74 $X2=-0.19
+ $Y2=-0.245
cc_803 N_A_245_411#_c_1229_n A_915_101# 0.00692367f $X=5.19 $Y=0.78 $X2=-0.19
+ $Y2=-0.245
cc_804 N_A_470_57#_c_1375_n N_VGND_M1007_d 0.00998235f $X=4.27 $Y=1.125 $X2=0
+ $Y2=0
cc_805 N_A_470_57#_c_1376_n N_VGND_M1012_d 0.0123776f $X=6.265 $Y=0.35 $X2=0
+ $Y2=0
cc_806 N_A_470_57#_c_1378_n N_VGND_M1012_d 0.00758552f $X=6.35 $Y=0.73 $X2=0
+ $Y2=0
cc_807 N_A_470_57#_c_1370_n N_VGND_c_1551_n 0.0133864f $X=3.395 $Y=0.35 $X2=0
+ $Y2=0
cc_808 N_A_470_57#_c_1371_n N_VGND_c_1551_n 0.0339147f $X=3.48 $Y=1.125 $X2=0
+ $Y2=0
cc_809 N_A_470_57#_c_1374_n N_VGND_c_1551_n 0.0198809f $X=3.765 $Y=1.21 $X2=0
+ $Y2=0
cc_810 N_A_470_57#_c_1375_n N_VGND_c_1551_n 0.0367753f $X=4.27 $Y=1.125 $X2=0
+ $Y2=0
cc_811 N_A_470_57#_c_1377_n N_VGND_c_1551_n 0.0141598f $X=4.355 $Y=0.35 $X2=0
+ $Y2=0
cc_812 N_A_470_57#_c_1376_n N_VGND_c_1552_n 0.0136054f $X=6.265 $Y=0.35 $X2=0
+ $Y2=0
cc_813 N_A_470_57#_c_1378_n N_VGND_c_1552_n 0.00820853f $X=6.35 $Y=0.73 $X2=0
+ $Y2=0
cc_814 N_A_470_57#_c_1379_n N_VGND_c_1552_n 0.0187531f $X=7.545 $Y=0.815 $X2=0
+ $Y2=0
cc_815 N_A_470_57#_c_1370_n N_VGND_c_1554_n 0.0563044f $X=3.395 $Y=0.35 $X2=0
+ $Y2=0
cc_816 N_A_470_57#_c_1383_n N_VGND_c_1554_n 0.0214013f $X=2.49 $Y=0.35 $X2=0
+ $Y2=0
cc_817 N_A_470_57#_c_1376_n N_VGND_c_1556_n 0.119254f $X=6.265 $Y=0.35 $X2=0
+ $Y2=0
cc_818 N_A_470_57#_c_1377_n N_VGND_c_1556_n 0.0114622f $X=4.355 $Y=0.35 $X2=0
+ $Y2=0
cc_819 N_A_470_57#_c_1379_n N_VGND_c_1556_n 0.00269575f $X=7.545 $Y=0.815 $X2=0
+ $Y2=0
cc_820 N_A_470_57#_c_1379_n N_VGND_c_1559_n 0.00967367f $X=7.545 $Y=0.815 $X2=0
+ $Y2=0
cc_821 N_A_470_57#_c_1381_n N_VGND_c_1559_n 0.0251191f $X=7.71 $Y=0.47 $X2=0
+ $Y2=0
cc_822 N_A_470_57#_M1019_d N_VGND_c_1561_n 0.00356488f $X=7.46 $Y=0.235 $X2=0
+ $Y2=0
cc_823 N_A_470_57#_c_1370_n N_VGND_c_1561_n 0.0342298f $X=3.395 $Y=0.35 $X2=0
+ $Y2=0
cc_824 N_A_470_57#_c_1376_n N_VGND_c_1561_n 0.0765665f $X=6.265 $Y=0.35 $X2=0
+ $Y2=0
cc_825 N_A_470_57#_c_1377_n N_VGND_c_1561_n 0.00657784f $X=4.355 $Y=0.35 $X2=0
+ $Y2=0
cc_826 N_A_470_57#_c_1379_n N_VGND_c_1561_n 0.0223173f $X=7.545 $Y=0.815 $X2=0
+ $Y2=0
cc_827 N_A_470_57#_c_1381_n N_VGND_c_1561_n 0.0154606f $X=7.71 $Y=0.47 $X2=0
+ $Y2=0
cc_828 N_A_470_57#_c_1383_n N_VGND_c_1561_n 0.0124501f $X=2.49 $Y=0.35 $X2=0
+ $Y2=0
cc_829 N_A_470_57#_c_1371_n A_684_101# 0.00356941f $X=3.48 $Y=1.125 $X2=-0.19
+ $Y2=-0.245
cc_830 N_A_470_57#_c_1376_n A_1112_47# 0.00601709f $X=6.265 $Y=0.35 $X2=-0.19
+ $Y2=-0.245
cc_831 A_114_47# N_VGND_c_1561_n 0.00417822f $X=0.57 $Y=0.235 $X2=0 $Y2=0
cc_832 N_VGND_c_1561_n A_1112_47# 0.00193256f $X=9.84 $Y=0 $X2=-0.19 $Y2=-0.245
cc_833 N_VGND_c_1561_n A_1414_47# 0.00312641f $X=9.84 $Y=0 $X2=-0.19 $Y2=-0.245
cc_834 N_VGND_c_1561_n A_1600_47# 0.0111053f $X=9.84 $Y=0 $X2=-0.19 $Y2=-0.245
cc_835 N_VGND_c_1561_n A_1860_47# 0.00314438f $X=9.84 $Y=0 $X2=-0.19 $Y2=-0.245
