* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__o21ba_2 A1 A2 B1_N VGND VNB VPB VPWR X
X0 a_186_21# a_28_131# a_492_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X1 VGND A1 a_492_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X2 a_28_131# B1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X3 a_492_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X4 VPWR a_28_131# a_186_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X5 a_28_131# B1_N VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 VGND a_186_21# X VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X7 X a_186_21# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X8 X a_186_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X9 a_186_21# A2 a_564_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X10 VPWR a_186_21# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X11 a_564_367# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
.ends
