* File: sky130_fd_sc_lp__and2b_m.pxi.spice
* Created: Fri Aug 28 10:05:36 2020
* 
x_PM_SKY130_FD_SC_LP__AND2B_M%A_N N_A_N_c_55_n N_A_N_M1007_g N_A_N_c_56_n
+ N_A_N_M1000_g A_N A_N PM_SKY130_FD_SC_LP__AND2B_M%A_N
x_PM_SKY130_FD_SC_LP__AND2B_M%A_35_70# N_A_35_70#_M1007_s N_A_35_70#_M1000_s
+ N_A_35_70#_M1006_g N_A_35_70#_c_89_n N_A_35_70#_c_90_n N_A_35_70#_c_91_n
+ N_A_35_70#_M1002_g N_A_35_70#_c_92_n N_A_35_70#_c_99_n N_A_35_70#_c_93_n
+ N_A_35_70#_c_94_n N_A_35_70#_c_102_n N_A_35_70#_c_103_n N_A_35_70#_c_95_n
+ N_A_35_70#_c_96_n N_A_35_70#_c_97_n PM_SKY130_FD_SC_LP__AND2B_M%A_35_70#
x_PM_SKY130_FD_SC_LP__AND2B_M%B N_B_M1003_g N_B_M1005_g B B B N_B_c_153_n
+ PM_SKY130_FD_SC_LP__AND2B_M%B
x_PM_SKY130_FD_SC_LP__AND2B_M%A_255_47# N_A_255_47#_M1002_s N_A_255_47#_M1006_d
+ N_A_255_47#_c_188_n N_A_255_47#_M1004_g N_A_255_47#_M1001_g
+ N_A_255_47#_c_186_n N_A_255_47#_c_190_n N_A_255_47#_c_187_n
+ N_A_255_47#_c_203_n N_A_255_47#_c_192_n PM_SKY130_FD_SC_LP__AND2B_M%A_255_47#
x_PM_SKY130_FD_SC_LP__AND2B_M%VPWR N_VPWR_M1000_d N_VPWR_M1003_d N_VPWR_c_242_n
+ N_VPWR_c_243_n N_VPWR_c_244_n N_VPWR_c_245_n VPWR N_VPWR_c_246_n
+ N_VPWR_c_247_n N_VPWR_c_241_n N_VPWR_c_249_n PM_SKY130_FD_SC_LP__AND2B_M%VPWR
x_PM_SKY130_FD_SC_LP__AND2B_M%X N_X_M1004_d N_X_M1001_d X X X X X X X
+ PM_SKY130_FD_SC_LP__AND2B_M%X
x_PM_SKY130_FD_SC_LP__AND2B_M%VGND N_VGND_M1007_d N_VGND_M1005_d N_VGND_c_288_n
+ N_VGND_c_289_n VGND N_VGND_c_290_n N_VGND_c_291_n N_VGND_c_292_n
+ N_VGND_c_293_n N_VGND_c_294_n N_VGND_c_295_n PM_SKY130_FD_SC_LP__AND2B_M%VGND
cc_1 VNB N_A_N_c_55_n 0.0229734f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=0.88
cc_2 VNB N_A_N_c_56_n 0.0471157f $X=-0.19 $Y=-0.245 $X2=0.725 $Y2=1.36
cc_3 VNB N_A_N_M1000_g 0.017386f $X=-0.19 $Y=-0.245 $X2=0.725 $Y2=2.195
cc_4 VNB A_N 0.01582f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=0.84
cc_5 VNB N_A_35_70#_c_89_n 0.0246039f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_6 VNB N_A_35_70#_c_90_n 0.0105814f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_A_35_70#_c_91_n 0.0195534f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_35_70#_c_92_n 0.042416f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.11
cc_9 VNB N_A_35_70#_c_93_n 0.00811682f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=1.11
cc_10 VNB N_A_35_70#_c_94_n 0.0145978f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_35_70#_c_95_n 0.0137458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_35_70#_c_96_n 0.00376122f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_35_70#_c_97_n 0.0329928f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_B_M1005_g 0.0349511f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB B 0.0109846f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_B_c_153_n 0.0518586f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=1.045
cc_17 VNB N_A_255_47#_M1004_g 0.0680429f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_255_47#_c_186_n 0.00310175f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_255_47#_c_187_n 0.0107282f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_VPWR_c_241_n 0.123877f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB X 0.0501493f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_VGND_c_288_n 0.0102033f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_VGND_c_289_n 0.00482866f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_VGND_c_290_n 0.0181026f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.045
cc_25 VNB N_VGND_c_291_n 0.0346119f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_292_n 0.0197547f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_293_n 0.181599f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_294_n 0.00598062f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_295_n 0.00362723f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VPB N_A_N_M1000_g 0.0370224f $X=-0.19 $Y=1.655 $X2=0.725 $Y2=2.195
cc_31 VPB N_A_35_70#_M1006_g 0.0229603f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_32 VPB N_A_35_70#_c_99_n 0.0142692f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=1.11
cc_33 VPB N_A_35_70#_c_93_n 0.00751706f $X=-0.19 $Y=1.655 $X2=1.2 $Y2=1.11
cc_34 VPB N_A_35_70#_c_94_n 0.0187745f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_35 VPB N_A_35_70#_c_102_n 0.0164141f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_36 VPB N_A_35_70#_c_103_n 0.00227427f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_37 VPB N_A_35_70#_c_96_n 0.00423137f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_38 VPB N_B_M1003_g 0.0187113f $X=-0.19 $Y=1.655 $X2=0.515 $Y2=0.56
cc_39 VPB B 0.00957038f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_40 VPB N_B_c_153_n 0.0256603f $X=-0.19 $Y=1.655 $X2=0.62 $Y2=1.045
cc_41 VPB N_A_255_47#_c_188_n 0.0517083f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_42 VPB N_A_255_47#_M1004_g 0.0427932f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_43 VPB N_A_255_47#_c_190_n 0.00982965f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_44 VPB N_A_255_47#_c_187_n 0.00287456f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_45 VPB N_A_255_47#_c_192_n 0.0461514f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_46 VPB N_VPWR_c_242_n 0.0386043f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_47 VPB N_VPWR_c_243_n 0.0178503f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_48 VPB N_VPWR_c_244_n 0.0293511f $X=-0.19 $Y=1.655 $X2=0.62 $Y2=1.045
cc_49 VPB N_VPWR_c_245_n 0.00401341f $X=-0.19 $Y=1.655 $X2=0.605 $Y2=1.045
cc_50 VPB N_VPWR_c_246_n 0.0270348f $X=-0.19 $Y=1.655 $X2=1.2 $Y2=1.11
cc_51 VPB N_VPWR_c_247_n 0.0182027f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_52 VPB N_VPWR_c_241_n 0.0972115f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_53 VPB N_VPWR_c_249_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_54 VPB X 0.0411867f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_55 N_A_N_M1000_g N_A_35_70#_M1006_g 0.0154002f $X=0.725 $Y=2.195 $X2=0 $Y2=0
cc_56 N_A_N_c_55_n N_A_35_70#_c_90_n 0.00263248f $X=0.515 $Y=0.88 $X2=0 $Y2=0
cc_57 N_A_N_c_56_n N_A_35_70#_c_90_n 0.00849795f $X=0.725 $Y=1.36 $X2=0 $Y2=0
cc_58 A_N N_A_35_70#_c_90_n 0.00470045f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_59 N_A_N_c_55_n N_A_35_70#_c_92_n 0.0149945f $X=0.515 $Y=0.88 $X2=0 $Y2=0
cc_60 N_A_N_c_56_n N_A_35_70#_c_92_n 8.20771e-19 $X=0.725 $Y=1.36 $X2=0 $Y2=0
cc_61 N_A_N_M1000_g N_A_35_70#_c_92_n 0.00585822f $X=0.725 $Y=2.195 $X2=0 $Y2=0
cc_62 A_N N_A_35_70#_c_92_n 0.0418963f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_63 N_A_N_M1000_g N_A_35_70#_c_99_n 0.00764363f $X=0.725 $Y=2.195 $X2=0 $Y2=0
cc_64 N_A_N_c_56_n N_A_35_70#_c_93_n 0.00335553f $X=0.725 $Y=1.36 $X2=0 $Y2=0
cc_65 N_A_N_M1000_g N_A_35_70#_c_93_n 0.0157762f $X=0.725 $Y=2.195 $X2=0 $Y2=0
cc_66 A_N N_A_35_70#_c_93_n 0.0545826f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_67 N_A_N_M1000_g N_A_35_70#_c_94_n 0.0218758f $X=0.725 $Y=2.195 $X2=0 $Y2=0
cc_68 A_N N_A_35_70#_c_94_n 0.00451733f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_69 N_A_N_M1000_g N_A_35_70#_c_103_n 0.00428852f $X=0.725 $Y=2.195 $X2=0 $Y2=0
cc_70 N_A_N_c_55_n N_A_35_70#_c_95_n 4.41817e-19 $X=0.515 $Y=0.88 $X2=0 $Y2=0
cc_71 N_A_N_c_56_n N_A_35_70#_c_97_n 0.00919109f $X=0.725 $Y=1.36 $X2=0 $Y2=0
cc_72 A_N N_A_35_70#_c_97_n 0.01635f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_73 A_N N_B_c_153_n 2.22503e-19 $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_74 A_N N_A_255_47#_c_186_n 0.00303235f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_75 A_N N_A_255_47#_c_187_n 0.0333477f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_76 N_A_N_M1000_g N_VPWR_c_242_n 0.00338988f $X=0.725 $Y=2.195 $X2=0 $Y2=0
cc_77 N_A_N_M1000_g N_VPWR_c_241_n 0.00393927f $X=0.725 $Y=2.195 $X2=0 $Y2=0
cc_78 N_A_N_c_55_n N_VGND_c_288_n 0.0106688f $X=0.515 $Y=0.88 $X2=0 $Y2=0
cc_79 N_A_N_c_56_n N_VGND_c_288_n 0.00115686f $X=0.725 $Y=1.36 $X2=0 $Y2=0
cc_80 A_N N_VGND_c_288_n 0.019543f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_81 N_A_N_c_55_n N_VGND_c_290_n 0.00396895f $X=0.515 $Y=0.88 $X2=0 $Y2=0
cc_82 N_A_N_c_55_n N_VGND_c_293_n 0.00653476f $X=0.515 $Y=0.88 $X2=0 $Y2=0
cc_83 A_N N_VGND_c_293_n 0.0158439f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_84 N_A_35_70#_c_94_n N_B_M1003_g 0.0217618f $X=1.175 $Y=1.66 $X2=0 $Y2=0
cc_85 N_A_35_70#_c_91_n N_B_M1005_g 0.0508176f $X=1.615 $Y=0.765 $X2=0 $Y2=0
cc_86 N_A_35_70#_c_97_n N_B_M1005_g 0.00335829f $X=1.175 $Y=1.495 $X2=0 $Y2=0
cc_87 N_A_35_70#_c_89_n B 4.52911e-19 $X=1.54 $Y=0.84 $X2=0 $Y2=0
cc_88 N_A_35_70#_c_89_n N_B_c_153_n 0.00389988f $X=1.54 $Y=0.84 $X2=0 $Y2=0
cc_89 N_A_35_70#_c_97_n N_B_c_153_n 0.0217618f $X=1.175 $Y=1.495 $X2=0 $Y2=0
cc_90 N_A_35_70#_c_90_n N_A_255_47#_c_186_n 0.00952216f $X=1.34 $Y=0.84 $X2=0
+ $Y2=0
cc_91 N_A_35_70#_c_91_n N_A_255_47#_c_186_n 0.00603715f $X=1.615 $Y=0.765 $X2=0
+ $Y2=0
cc_92 N_A_35_70#_M1006_g N_A_255_47#_c_190_n 0.00134899f $X=1.265 $Y=2.195 $X2=0
+ $Y2=0
cc_93 N_A_35_70#_c_89_n N_A_255_47#_c_187_n 0.011406f $X=1.54 $Y=0.84 $X2=0
+ $Y2=0
cc_94 N_A_35_70#_c_91_n N_A_255_47#_c_187_n 0.00539348f $X=1.615 $Y=0.765 $X2=0
+ $Y2=0
cc_95 N_A_35_70#_c_93_n N_A_255_47#_c_187_n 0.0128545f $X=1.175 $Y=1.66 $X2=0
+ $Y2=0
cc_96 N_A_35_70#_c_94_n N_A_255_47#_c_187_n 0.0079633f $X=1.175 $Y=1.66 $X2=0
+ $Y2=0
cc_97 N_A_35_70#_c_97_n N_A_255_47#_c_187_n 0.00755573f $X=1.175 $Y=1.495 $X2=0
+ $Y2=0
cc_98 N_A_35_70#_M1006_g N_A_255_47#_c_203_n 0.00402967f $X=1.265 $Y=2.195 $X2=0
+ $Y2=0
cc_99 N_A_35_70#_c_93_n N_A_255_47#_c_203_n 8.29608e-19 $X=1.175 $Y=1.66 $X2=0
+ $Y2=0
cc_100 N_A_35_70#_M1006_g N_VPWR_c_242_n 0.00425398f $X=1.265 $Y=2.195 $X2=0
+ $Y2=0
cc_101 N_A_35_70#_c_93_n N_VPWR_c_242_n 0.010005f $X=1.175 $Y=1.66 $X2=0 $Y2=0
cc_102 N_A_35_70#_c_94_n N_VPWR_c_242_n 0.00124349f $X=1.175 $Y=1.66 $X2=0 $Y2=0
cc_103 N_A_35_70#_M1006_g N_VPWR_c_241_n 0.00393927f $X=1.265 $Y=2.195 $X2=0
+ $Y2=0
cc_104 N_A_35_70#_c_91_n N_VGND_c_288_n 0.00441631f $X=1.615 $Y=0.765 $X2=0
+ $Y2=0
cc_105 N_A_35_70#_c_95_n N_VGND_c_288_n 0.0103887f $X=0.3 $Y=0.495 $X2=0 $Y2=0
cc_106 N_A_35_70#_c_95_n N_VGND_c_290_n 0.0102241f $X=0.3 $Y=0.495 $X2=0 $Y2=0
cc_107 N_A_35_70#_c_90_n N_VGND_c_291_n 0.00115038f $X=1.34 $Y=0.84 $X2=0 $Y2=0
cc_108 N_A_35_70#_c_91_n N_VGND_c_291_n 0.00387067f $X=1.615 $Y=0.765 $X2=0
+ $Y2=0
cc_109 N_A_35_70#_c_90_n N_VGND_c_293_n 0.00121127f $X=1.34 $Y=0.84 $X2=0 $Y2=0
cc_110 N_A_35_70#_c_91_n N_VGND_c_293_n 0.00677977f $X=1.615 $Y=0.765 $X2=0
+ $Y2=0
cc_111 N_A_35_70#_c_95_n N_VGND_c_293_n 0.00792374f $X=0.3 $Y=0.495 $X2=0 $Y2=0
cc_112 N_B_M1003_g N_A_255_47#_M1004_g 0.0099952f $X=1.695 $Y=2.195 $X2=0 $Y2=0
cc_113 N_B_M1005_g N_A_255_47#_M1004_g 0.0305376f $X=1.975 $Y=0.445 $X2=0 $Y2=0
cc_114 B N_A_255_47#_M1004_g 0.00796966f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_115 N_B_c_153_n N_A_255_47#_M1004_g 0.0393306f $X=1.955 $Y=1.32 $X2=0 $Y2=0
cc_116 N_B_M1005_g N_A_255_47#_c_186_n 9.538e-19 $X=1.975 $Y=0.445 $X2=0 $Y2=0
cc_117 N_B_M1003_g N_A_255_47#_c_190_n 0.00526027f $X=1.695 $Y=2.195 $X2=0 $Y2=0
cc_118 N_B_M1003_g N_A_255_47#_c_187_n 0.00967667f $X=1.695 $Y=2.195 $X2=0 $Y2=0
cc_119 N_B_M1005_g N_A_255_47#_c_187_n 0.00247195f $X=1.975 $Y=0.445 $X2=0 $Y2=0
cc_120 B N_A_255_47#_c_187_n 0.0701227f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_121 N_B_c_153_n N_A_255_47#_c_187_n 0.0183151f $X=1.955 $Y=1.32 $X2=0 $Y2=0
cc_122 N_B_M1003_g N_A_255_47#_c_203_n 0.0039653f $X=1.695 $Y=2.195 $X2=0 $Y2=0
cc_123 N_B_M1003_g N_A_255_47#_c_192_n 0.00891663f $X=1.695 $Y=2.195 $X2=0 $Y2=0
cc_124 N_B_M1003_g N_VPWR_c_243_n 0.00355358f $X=1.695 $Y=2.195 $X2=0 $Y2=0
cc_125 B N_VPWR_c_243_n 0.0130394f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_126 N_B_c_153_n N_VPWR_c_243_n 8.23511e-19 $X=1.955 $Y=1.32 $X2=0 $Y2=0
cc_127 B X 0.0579585f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_128 N_B_M1005_g N_VGND_c_289_n 0.00285763f $X=1.975 $Y=0.445 $X2=0 $Y2=0
cc_129 B N_VGND_c_289_n 0.00821139f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_130 N_B_M1005_g N_VGND_c_291_n 0.00585385f $X=1.975 $Y=0.445 $X2=0 $Y2=0
cc_131 N_B_M1005_g N_VGND_c_293_n 0.00613579f $X=1.975 $Y=0.445 $X2=0 $Y2=0
cc_132 B N_VGND_c_293_n 0.00802068f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_133 N_A_255_47#_c_190_n N_VPWR_c_242_n 0.0259151f $X=1.592 $Y=2.855 $X2=0
+ $Y2=0
cc_134 N_A_255_47#_c_187_n N_VPWR_c_242_n 0.00213552f $X=1.605 $Y=2.155 $X2=0
+ $Y2=0
cc_135 N_A_255_47#_c_203_n N_VPWR_c_242_n 0.0117555f $X=1.605 $Y=2.26 $X2=0
+ $Y2=0
cc_136 N_A_255_47#_c_192_n N_VPWR_c_242_n 0.00489234f $X=1.66 $Y=2.85 $X2=0
+ $Y2=0
cc_137 N_A_255_47#_c_188_n N_VPWR_c_243_n 0.0254733f $X=2.33 $Y=2.85 $X2=0 $Y2=0
cc_138 N_A_255_47#_M1004_g N_VPWR_c_243_n 0.0128556f $X=2.405 $Y=0.445 $X2=0
+ $Y2=0
cc_139 N_A_255_47#_c_190_n N_VPWR_c_243_n 0.0367073f $X=1.592 $Y=2.855 $X2=0
+ $Y2=0
cc_140 N_A_255_47#_c_203_n N_VPWR_c_243_n 0.0101868f $X=1.605 $Y=2.26 $X2=0
+ $Y2=0
cc_141 N_A_255_47#_c_192_n N_VPWR_c_243_n 0.00374798f $X=1.66 $Y=2.85 $X2=0
+ $Y2=0
cc_142 N_A_255_47#_c_188_n N_VPWR_c_246_n 0.00445258f $X=2.33 $Y=2.85 $X2=0
+ $Y2=0
cc_143 N_A_255_47#_c_190_n N_VPWR_c_246_n 0.0152941f $X=1.592 $Y=2.855 $X2=0
+ $Y2=0
cc_144 N_A_255_47#_c_192_n N_VPWR_c_246_n 0.00593936f $X=1.66 $Y=2.85 $X2=0
+ $Y2=0
cc_145 N_A_255_47#_c_188_n N_VPWR_c_247_n 0.00449461f $X=2.33 $Y=2.85 $X2=0
+ $Y2=0
cc_146 N_A_255_47#_c_188_n N_VPWR_c_241_n 0.009566f $X=2.33 $Y=2.85 $X2=0 $Y2=0
cc_147 N_A_255_47#_c_190_n N_VPWR_c_241_n 0.0104794f $X=1.592 $Y=2.855 $X2=0
+ $Y2=0
cc_148 N_A_255_47#_c_192_n N_VPWR_c_241_n 0.00814482f $X=1.66 $Y=2.85 $X2=0
+ $Y2=0
cc_149 N_A_255_47#_M1004_g X 0.0504487f $X=2.405 $Y=0.445 $X2=0 $Y2=0
cc_150 N_A_255_47#_c_186_n N_VGND_c_288_n 0.0102737f $X=1.52 $Y=0.51 $X2=0 $Y2=0
cc_151 N_A_255_47#_M1004_g N_VGND_c_289_n 0.00274937f $X=2.405 $Y=0.445 $X2=0
+ $Y2=0
cc_152 N_A_255_47#_c_186_n N_VGND_c_291_n 0.0142558f $X=1.52 $Y=0.51 $X2=0 $Y2=0
cc_153 N_A_255_47#_M1004_g N_VGND_c_292_n 0.00585385f $X=2.405 $Y=0.445 $X2=0
+ $Y2=0
cc_154 N_A_255_47#_M1002_s N_VGND_c_293_n 0.00236038f $X=1.275 $Y=0.235 $X2=0
+ $Y2=0
cc_155 N_A_255_47#_M1004_g N_VGND_c_293_n 0.0117829f $X=2.405 $Y=0.445 $X2=0
+ $Y2=0
cc_156 N_A_255_47#_c_186_n N_VGND_c_293_n 0.015066f $X=1.52 $Y=0.51 $X2=0 $Y2=0
cc_157 N_VPWR_c_243_n X 0.0421725f $X=2.17 $Y=2.26 $X2=0 $Y2=0
cc_158 N_VPWR_c_247_n X 0.00623633f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_159 N_VPWR_c_241_n X 0.00710559f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_160 X N_VGND_c_292_n 0.00877924f $X=2.555 $Y=0.47 $X2=0 $Y2=0
cc_161 N_X_M1004_d N_VGND_c_293_n 0.0042053f $X=2.48 $Y=0.235 $X2=0 $Y2=0
cc_162 X N_VGND_c_293_n 0.00770513f $X=2.555 $Y=0.47 $X2=0 $Y2=0
cc_163 N_VGND_c_293_n A_338_47# 0.00817721f $X=2.64 $Y=0 $X2=-0.19 $Y2=-0.245
