* File: sky130_fd_sc_lp__a22o_4.spice
* Created: Fri Aug 28 09:54:23 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__a22o_4.pex.spice"
.subckt sky130_fd_sc_lp__a22o_4  VNB VPB B2 B1 A2 A1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A1	A1
* A2	A2
* B1	B1
* B2	B2
* VPB	VPB
* VNB	VNB
MM1003 N_VGND_M1003_d N_A_103_263#_M1003_g N_X_M1003_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75005.1 A=0.126 P=1.98 MULT=1
MM1010 N_VGND_M1010_d N_A_103_263#_M1010_g N_X_M1003_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75004.7 A=0.126 P=1.98 MULT=1
MM1021 N_VGND_M1010_d N_A_103_263#_M1021_g N_X_M1021_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.1
+ SB=75004.3 A=0.126 P=1.98 MULT=1
MM1022 N_VGND_M1022_d N_A_103_263#_M1022_g N_X_M1021_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1491 AS=0.1176 PD=1.195 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.5
+ SB=75003.9 A=0.126 P=1.98 MULT=1
MM1015 N_VGND_M1022_d N_B2_M1015_g N_A_632_47#_M1015_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1491 AS=0.1176 PD=1.195 PS=1.12 NRD=10.704 NRS=0 M=1 R=5.6 SA=75002
+ SB=75003.3 A=0.126 P=1.98 MULT=1
MM1001 N_A_103_263#_M1001_d N_B1_M1001_g N_A_632_47#_M1015_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002.4
+ SB=75002.9 A=0.126 P=1.98 MULT=1
MM1006 N_A_103_263#_M1001_d N_B1_M1006_g N_A_632_47#_M1006_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002.8
+ SB=75002.5 A=0.126 P=1.98 MULT=1
MM1020 N_VGND_M1020_d N_B2_M1020_g N_A_632_47#_M1006_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1806 AS=0.1176 PD=1.27 PS=1.12 NRD=2.856 NRS=0 M=1 R=5.6 SA=75003.3
+ SB=75002.1 A=0.126 P=1.98 MULT=1
MM1013 N_A_1006_47#_M1013_d N_A2_M1013_g N_VGND_M1020_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1806 PD=1.12 PS=1.27 NRD=0 NRS=18.564 M=1 R=5.6 SA=75003.9
+ SB=75001.5 A=0.126 P=1.98 MULT=1
MM1007 N_A_1006_47#_M1013_d N_A1_M1007_g N_A_103_263#_M1007_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75004.3
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1018 N_A_1006_47#_M1018_d N_A1_M1018_g N_A_103_263#_M1007_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75004.7
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1016 N_A_1006_47#_M1018_d N_A2_M1016_g N_VGND_M1016_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75005.1
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1000 N_X_M1000_d N_A_103_263#_M1000_g N_VPWR_M1000_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75001.5 A=0.189 P=2.82 MULT=1
MM1008 N_X_M1000_d N_A_103_263#_M1008_g N_VPWR_M1008_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1011 N_X_M1011_d N_A_103_263#_M1011_g N_VPWR_M1008_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1014 N_X_M1011_d N_A_103_263#_M1014_g N_VPWR_M1014_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75001.5
+ SB=75000.2 A=0.189 P=2.82 MULT=1
MM1005 N_A_549_367#_M1005_d N_B2_M1005_g N_A_103_263#_M1005_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75003.3 A=0.189 P=2.82 MULT=1
MM1004 N_A_549_367#_M1004_d N_B1_M1004_g N_A_103_263#_M1005_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75002.9 A=0.189 P=2.82 MULT=1
MM1019 N_A_549_367#_M1004_d N_B1_M1019_g N_A_103_263#_M1019_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75002.5 A=0.189 P=2.82 MULT=1
MM1023 N_A_549_367#_M1023_d N_B2_M1023_g N_A_103_263#_M1019_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.2205 AS=0.1764 PD=1.61 PS=1.54 NRD=6.2449 NRS=0 M=1 R=8.4
+ SA=75001.5 SB=75002.1 A=0.189 P=2.82 MULT=1
MM1012 N_VPWR_M1012_d N_A2_M1012_g N_A_549_367#_M1023_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.2268 AS=0.2205 PD=1.62 PS=1.61 NRD=6.2449 NRS=4.6886 M=1 R=8.4
+ SA=75002 SB=75001.6 A=0.189 P=2.82 MULT=1
MM1002 N_VPWR_M1012_d N_A1_M1002_g N_A_549_367#_M1002_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.2268 AS=0.1764 PD=1.62 PS=1.54 NRD=6.2449 NRS=0 M=1 R=8.4
+ SA=75002.5 SB=75001.1 A=0.189 P=2.82 MULT=1
MM1009 N_VPWR_M1009_d N_A1_M1009_g N_A_549_367#_M1002_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.9
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1017 N_VPWR_M1009_d N_A2_M1017_g N_A_549_367#_M1017_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75003.3
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX24_noxref VNB VPB NWDIODE A=13.2415 P=17.93
*
.include "sky130_fd_sc_lp__a22o_4.pxi.spice"
*
.ends
*
*
