* File: sky130_fd_sc_lp__a21oi_m.pxi.spice
* Created: Wed Sep  2 09:20:57 2020
* 
x_PM_SKY130_FD_SC_LP__A21OI_M%A2 N_A2_c_49_n N_A2_M1001_g N_A2_M1005_g
+ N_A2_c_51_n N_A2_c_52_n N_A2_c_57_n A2 A2 A2 A2 N_A2_c_54_n
+ PM_SKY130_FD_SC_LP__A21OI_M%A2
x_PM_SKY130_FD_SC_LP__A21OI_M%A1 N_A1_M1002_g N_A1_M1004_g N_A1_c_89_n
+ N_A1_c_94_n A1 A1 A1 A1 N_A1_c_91_n PM_SKY130_FD_SC_LP__A21OI_M%A1
x_PM_SKY130_FD_SC_LP__A21OI_M%B1 N_B1_M1003_g N_B1_M1000_g N_B1_c_136_n
+ N_B1_c_137_n B1 B1 N_B1_c_138_n N_B1_c_139_n PM_SKY130_FD_SC_LP__A21OI_M%B1
x_PM_SKY130_FD_SC_LP__A21OI_M%A_27_504# N_A_27_504#_M1001_s N_A_27_504#_M1004_d
+ N_A_27_504#_c_173_n N_A_27_504#_c_174_n N_A_27_504#_c_175_n
+ N_A_27_504#_c_176_n PM_SKY130_FD_SC_LP__A21OI_M%A_27_504#
x_PM_SKY130_FD_SC_LP__A21OI_M%VPWR N_VPWR_M1001_d N_VPWR_c_198_n VPWR
+ N_VPWR_c_199_n N_VPWR_c_200_n N_VPWR_c_197_n N_VPWR_c_202_n
+ PM_SKY130_FD_SC_LP__A21OI_M%VPWR
x_PM_SKY130_FD_SC_LP__A21OI_M%Y N_Y_M1002_d N_Y_M1003_d N_Y_c_224_n N_Y_c_219_n
+ N_Y_c_220_n N_Y_c_221_n Y N_Y_c_223_n PM_SKY130_FD_SC_LP__A21OI_M%Y
x_PM_SKY130_FD_SC_LP__A21OI_M%VGND N_VGND_M1005_s N_VGND_M1000_d N_VGND_c_247_n
+ N_VGND_c_248_n N_VGND_c_249_n N_VGND_c_250_n VGND N_VGND_c_251_n
+ N_VGND_c_252_n PM_SKY130_FD_SC_LP__A21OI_M%VGND
cc_1 VNB N_A2_c_49_n 0.00892806f $X=-0.19 $Y=-0.245 $X2=0.335 $Y2=2.14
cc_2 VNB N_A2_M1005_g 0.0275084f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=0.445
cc_3 VNB N_A2_c_51_n 0.0369223f $X=-0.19 $Y=-0.245 $X2=0.35 $Y2=0.99
cc_4 VNB N_A2_c_52_n 0.0233012f $X=-0.19 $Y=-0.245 $X2=0.275 $Y2=1.51
cc_5 VNB A2 0.00769149f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_6 VNB N_A2_c_54_n 0.0375699f $X=-0.19 $Y=-0.245 $X2=0.275 $Y2=1.005
cc_7 VNB N_A1_M1002_g 0.040321f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.29
cc_8 VNB N_A1_c_89_n 0.0165156f $X=-0.19 $Y=-0.245 $X2=0.275 $Y2=0.99
cc_9 VNB A1 0.00916315f $X=-0.19 $Y=-0.245 $X2=0.35 $Y2=0.99
cc_10 VNB N_A1_c_91_n 0.0163297f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_11 VNB N_B1_M1000_g 0.0387192f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=0.84
cc_12 VNB N_B1_c_136_n 0.0236573f $X=-0.19 $Y=-0.245 $X2=0.275 $Y2=0.99
cc_13 VNB N_B1_c_137_n 0.00489944f $X=-0.19 $Y=-0.245 $X2=0.35 $Y2=0.84
cc_14 VNB N_B1_c_138_n 0.0167796f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.215
cc_15 VNB N_B1_c_139_n 0.00590315f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_VPWR_c_197_n 0.0840719f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.215
cc_17 VNB N_Y_c_219_n 0.0169098f $X=-0.19 $Y=-0.245 $X2=0.275 $Y2=0.99
cc_18 VNB N_Y_c_220_n 0.00485541f $X=-0.19 $Y=-0.245 $X2=0.35 $Y2=0.84
cc_19 VNB N_Y_c_221_n 0.0390303f $X=-0.19 $Y=-0.245 $X2=0.275 $Y2=1.345
cc_20 VNB N_VGND_c_247_n 0.012433f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=0.84
cc_21 VNB N_VGND_c_248_n 0.00495479f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=0.445
cc_22 VNB N_VGND_c_249_n 0.012155f $X=-0.19 $Y=-0.245 $X2=0.275 $Y2=0.99
cc_23 VNB N_VGND_c_250_n 0.0126513f $X=-0.19 $Y=-0.245 $X2=0.35 $Y2=0.99
cc_24 VNB N_VGND_c_251_n 0.0294198f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_252_n 0.129999f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VPB N_A2_c_49_n 0.0318286f $X=-0.19 $Y=1.655 $X2=0.335 $Y2=2.14
cc_27 VPB N_A2_M1001_g 0.0279535f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.73
cc_28 VPB N_A2_c_57_n 0.0255288f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.215
cc_29 VPB A2 0.0173406f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_30 VPB N_A1_M1004_g 0.0423944f $X=-0.19 $Y=1.655 $X2=0.515 $Y2=0.84
cc_31 VPB N_A1_c_89_n 0.00508708f $X=-0.19 $Y=1.655 $X2=0.275 $Y2=0.99
cc_32 VPB N_A1_c_94_n 0.0160361f $X=-0.19 $Y=1.655 $X2=0.35 $Y2=0.84
cc_33 VPB A1 0.00527014f $X=-0.19 $Y=1.655 $X2=0.35 $Y2=0.99
cc_34 VPB N_B1_M1003_g 0.0594057f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.29
cc_35 VPB N_B1_c_137_n 0.013919f $X=-0.19 $Y=1.655 $X2=0.35 $Y2=0.84
cc_36 VPB N_B1_c_139_n 0.00613967f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_37 VPB N_A_27_504#_c_173_n 0.00224906f $X=-0.19 $Y=1.655 $X2=0.515 $Y2=0.445
cc_38 VPB N_A_27_504#_c_174_n 0.0174607f $X=-0.19 $Y=1.655 $X2=0.275 $Y2=0.99
cc_39 VPB N_A_27_504#_c_175_n 0.00896362f $X=-0.19 $Y=1.655 $X2=0.35 $Y2=0.84
cc_40 VPB N_A_27_504#_c_176_n 9.04027e-19 $X=-0.19 $Y=1.655 $X2=0.275 $Y2=1.51
cc_41 VPB N_VPWR_c_198_n 0.00986829f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_42 VPB N_VPWR_c_199_n 0.0195493f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_43 VPB N_VPWR_c_200_n 0.0344639f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_44 VPB N_VPWR_c_197_n 0.0658703f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.215
cc_45 VPB N_VPWR_c_202_n 0.00401341f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_46 VPB N_Y_c_221_n 0.0438885f $X=-0.19 $Y=1.655 $X2=0.275 $Y2=1.345
cc_47 VPB N_Y_c_223_n 0.0160816f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_48 N_A2_M1005_g N_A1_M1002_g 0.0555919f $X=0.515 $Y=0.445 $X2=0 $Y2=0
cc_49 A2 N_A1_M1002_g 3.30198e-19 $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_50 N_A2_c_54_n N_A1_M1002_g 0.00727198f $X=0.275 $Y=1.005 $X2=0 $Y2=0
cc_51 N_A2_c_49_n N_A1_M1004_g 0.00574499f $X=0.335 $Y=2.14 $X2=0 $Y2=0
cc_52 N_A2_c_57_n N_A1_M1004_g 0.026932f $X=0.475 $Y=2.215 $X2=0 $Y2=0
cc_53 A2 N_A1_M1004_g 2.04016e-19 $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_54 N_A2_c_49_n N_A1_c_89_n 0.0195802f $X=0.335 $Y=2.14 $X2=0 $Y2=0
cc_55 N_A2_c_52_n N_A1_c_89_n 0.00875475f $X=0.275 $Y=1.51 $X2=0 $Y2=0
cc_56 N_A2_c_49_n A1 0.00402141f $X=0.335 $Y=2.14 $X2=0 $Y2=0
cc_57 N_A2_c_51_n A1 0.00137533f $X=0.35 $Y=0.99 $X2=0 $Y2=0
cc_58 A2 A1 0.0671896f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_59 N_A2_c_54_n A1 0.00381655f $X=0.275 $Y=1.005 $X2=0 $Y2=0
cc_60 A2 N_A1_c_91_n 7.59337e-19 $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_61 N_A2_c_54_n N_A1_c_91_n 0.00875475f $X=0.275 $Y=1.005 $X2=0 $Y2=0
cc_62 N_A2_M1001_g N_A_27_504#_c_173_n 0.00143084f $X=0.475 $Y=2.73 $X2=0 $Y2=0
cc_63 N_A2_M1001_g N_A_27_504#_c_174_n 0.0169197f $X=0.475 $Y=2.73 $X2=0 $Y2=0
cc_64 N_A2_c_57_n N_A_27_504#_c_174_n 0.00171009f $X=0.475 $Y=2.215 $X2=0 $Y2=0
cc_65 N_A2_c_57_n N_A_27_504#_c_175_n 0.0036012f $X=0.475 $Y=2.215 $X2=0 $Y2=0
cc_66 A2 N_A_27_504#_c_175_n 0.0174687f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_67 N_A2_M1001_g N_VPWR_c_198_n 0.00329204f $X=0.475 $Y=2.73 $X2=0 $Y2=0
cc_68 N_A2_M1001_g N_VPWR_c_199_n 0.00563421f $X=0.475 $Y=2.73 $X2=0 $Y2=0
cc_69 N_A2_M1001_g N_VPWR_c_197_n 0.00539454f $X=0.475 $Y=2.73 $X2=0 $Y2=0
cc_70 N_A2_M1005_g N_VGND_c_248_n 0.00460896f $X=0.515 $Y=0.445 $X2=0 $Y2=0
cc_71 N_A2_c_51_n N_VGND_c_248_n 0.00262124f $X=0.35 $Y=0.99 $X2=0 $Y2=0
cc_72 A2 N_VGND_c_248_n 0.00847718f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_73 N_A2_M1005_g N_VGND_c_251_n 0.00585385f $X=0.515 $Y=0.445 $X2=0 $Y2=0
cc_74 N_A2_M1005_g N_VGND_c_252_n 0.0114989f $X=0.515 $Y=0.445 $X2=0 $Y2=0
cc_75 N_A2_c_51_n N_VGND_c_252_n 0.0020393f $X=0.35 $Y=0.99 $X2=0 $Y2=0
cc_76 A2 N_VGND_c_252_n 0.00211986f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_77 N_A1_c_94_n N_B1_M1003_g 0.0436682f $X=0.815 $Y=1.9 $X2=0 $Y2=0
cc_78 A1 N_B1_M1003_g 0.00196704f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_79 N_A1_M1002_g N_B1_M1000_g 0.0260773f $X=0.875 $Y=0.445 $X2=0 $Y2=0
cc_80 A1 N_B1_M1000_g 0.00129508f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_81 N_A1_c_89_n N_B1_c_136_n 0.00904753f $X=0.815 $Y=1.735 $X2=0 $Y2=0
cc_82 N_A1_c_94_n N_B1_c_137_n 0.00904753f $X=0.815 $Y=1.9 $X2=0 $Y2=0
cc_83 N_A1_M1002_g N_B1_c_138_n 0.00639158f $X=0.875 $Y=0.445 $X2=0 $Y2=0
cc_84 A1 N_B1_c_138_n 6.378e-19 $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_85 N_A1_c_91_n N_B1_c_138_n 0.00904753f $X=0.815 $Y=1.395 $X2=0 $Y2=0
cc_86 N_A1_M1002_g N_B1_c_139_n 9.74622e-19 $X=0.875 $Y=0.445 $X2=0 $Y2=0
cc_87 A1 N_B1_c_139_n 0.0439645f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_88 N_A1_c_91_n N_B1_c_139_n 0.00372884f $X=0.815 $Y=1.395 $X2=0 $Y2=0
cc_89 N_A1_M1004_g N_A_27_504#_c_174_n 0.0139964f $X=0.905 $Y=2.73 $X2=0 $Y2=0
cc_90 N_A1_c_94_n N_A_27_504#_c_174_n 7.53204e-19 $X=0.815 $Y=1.9 $X2=0 $Y2=0
cc_91 A1 N_A_27_504#_c_174_n 0.0207532f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_92 N_A1_M1004_g N_A_27_504#_c_176_n 6.71115e-19 $X=0.905 $Y=2.73 $X2=0 $Y2=0
cc_93 N_A1_M1004_g N_VPWR_c_198_n 0.00329204f $X=0.905 $Y=2.73 $X2=0 $Y2=0
cc_94 N_A1_M1004_g N_VPWR_c_200_n 0.00563421f $X=0.905 $Y=2.73 $X2=0 $Y2=0
cc_95 N_A1_M1004_g N_VPWR_c_197_n 0.00539454f $X=0.905 $Y=2.73 $X2=0 $Y2=0
cc_96 N_A1_M1002_g N_Y_c_224_n 0.00511937f $X=0.875 $Y=0.445 $X2=0 $Y2=0
cc_97 N_A1_M1002_g N_Y_c_220_n 0.00505296f $X=0.875 $Y=0.445 $X2=0 $Y2=0
cc_98 N_A1_M1002_g N_VGND_c_250_n 0.00148212f $X=0.875 $Y=0.445 $X2=0 $Y2=0
cc_99 N_A1_M1002_g N_VGND_c_251_n 0.00585385f $X=0.875 $Y=0.445 $X2=0 $Y2=0
cc_100 N_A1_M1002_g N_VGND_c_252_n 0.00808671f $X=0.875 $Y=0.445 $X2=0 $Y2=0
cc_101 A1 N_VGND_c_252_n 0.00960739f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_102 N_B1_M1003_g N_A_27_504#_c_174_n 0.00227506f $X=1.335 $Y=2.73 $X2=0 $Y2=0
cc_103 N_B1_c_139_n N_A_27_504#_c_174_n 0.00437675f $X=1.385 $Y=1.245 $X2=0
+ $Y2=0
cc_104 N_B1_M1003_g N_A_27_504#_c_176_n 5.44271e-19 $X=1.335 $Y=2.73 $X2=0 $Y2=0
cc_105 N_B1_M1003_g N_VPWR_c_200_n 0.00563421f $X=1.335 $Y=2.73 $X2=0 $Y2=0
cc_106 N_B1_M1003_g N_VPWR_c_197_n 0.00539454f $X=1.335 $Y=2.73 $X2=0 $Y2=0
cc_107 N_B1_M1000_g N_Y_c_224_n 2.0895e-19 $X=1.38 $Y=0.445 $X2=0 $Y2=0
cc_108 N_B1_M1000_g N_Y_c_219_n 0.0134962f $X=1.38 $Y=0.445 $X2=0 $Y2=0
cc_109 N_B1_c_138_n N_Y_c_219_n 0.00351522f $X=1.385 $Y=1.245 $X2=0 $Y2=0
cc_110 N_B1_c_139_n N_Y_c_219_n 0.012661f $X=1.385 $Y=1.245 $X2=0 $Y2=0
cc_111 N_B1_c_138_n N_Y_c_220_n 2.16099e-19 $X=1.385 $Y=1.245 $X2=0 $Y2=0
cc_112 N_B1_c_139_n N_Y_c_220_n 0.00932176f $X=1.385 $Y=1.245 $X2=0 $Y2=0
cc_113 N_B1_M1003_g N_Y_c_221_n 0.021895f $X=1.335 $Y=2.73 $X2=0 $Y2=0
cc_114 N_B1_M1000_g N_Y_c_221_n 0.00813157f $X=1.38 $Y=0.445 $X2=0 $Y2=0
cc_115 N_B1_c_138_n N_Y_c_221_n 0.0163648f $X=1.385 $Y=1.245 $X2=0 $Y2=0
cc_116 N_B1_c_139_n N_Y_c_221_n 0.048424f $X=1.385 $Y=1.245 $X2=0 $Y2=0
cc_117 N_B1_M1000_g N_VGND_c_250_n 0.00979919f $X=1.38 $Y=0.445 $X2=0 $Y2=0
cc_118 N_B1_M1000_g N_VGND_c_251_n 0.0035715f $X=1.38 $Y=0.445 $X2=0 $Y2=0
cc_119 N_B1_M1000_g N_VGND_c_252_n 0.00446383f $X=1.38 $Y=0.445 $X2=0 $Y2=0
cc_120 N_A_27_504#_c_174_n N_VPWR_c_198_n 0.0142847f $X=1.015 $Y=2.385 $X2=0
+ $Y2=0
cc_121 N_A_27_504#_c_173_n N_VPWR_c_199_n 0.00519224f $X=0.26 $Y=2.665 $X2=0
+ $Y2=0
cc_122 N_A_27_504#_c_176_n N_VPWR_c_200_n 0.00467386f $X=1.12 $Y=2.645 $X2=0
+ $Y2=0
cc_123 N_A_27_504#_c_173_n N_VPWR_c_197_n 0.00688714f $X=0.26 $Y=2.665 $X2=0
+ $Y2=0
cc_124 N_A_27_504#_c_174_n N_VPWR_c_197_n 0.0146356f $X=1.015 $Y=2.385 $X2=0
+ $Y2=0
cc_125 N_A_27_504#_c_176_n N_VPWR_c_197_n 0.00677835f $X=1.12 $Y=2.645 $X2=0
+ $Y2=0
cc_126 N_A_27_504#_c_174_n N_Y_c_221_n 0.00756459f $X=1.015 $Y=2.385 $X2=0 $Y2=0
cc_127 N_A_27_504#_c_176_n N_Y_c_221_n 0.00216499f $X=1.12 $Y=2.645 $X2=0 $Y2=0
cc_128 N_VPWR_c_200_n N_Y_c_223_n 0.0101583f $X=1.68 $Y=3.33 $X2=0 $Y2=0
cc_129 N_VPWR_c_197_n N_Y_c_223_n 0.0124384f $X=1.68 $Y=3.33 $X2=0 $Y2=0
cc_130 N_Y_c_219_n N_VGND_c_249_n 0.00114637f $X=1.65 $Y=0.75 $X2=0 $Y2=0
cc_131 N_Y_c_219_n N_VGND_c_250_n 0.0227232f $X=1.65 $Y=0.75 $X2=0 $Y2=0
cc_132 N_Y_c_224_n N_VGND_c_251_n 0.00725952f $X=1.165 $Y=0.51 $X2=0 $Y2=0
cc_133 N_Y_c_219_n N_VGND_c_251_n 0.00283061f $X=1.65 $Y=0.75 $X2=0 $Y2=0
cc_134 N_Y_M1002_d N_VGND_c_252_n 0.00767588f $X=0.95 $Y=0.235 $X2=0 $Y2=0
cc_135 N_Y_c_224_n N_VGND_c_252_n 0.00615038f $X=1.165 $Y=0.51 $X2=0 $Y2=0
cc_136 N_Y_c_219_n N_VGND_c_252_n 0.0077335f $X=1.65 $Y=0.75 $X2=0 $Y2=0
cc_137 N_VGND_c_252_n A_118_47# 0.00437433f $X=1.68 $Y=0 $X2=-0.19 $Y2=-0.245
