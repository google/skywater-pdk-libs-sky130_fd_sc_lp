# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__o2bb2ai_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_lp__o2bb2ai_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.760000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1_N
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.375000 0.805000 1.920000 ;
        RECT 0.085000 1.920000 2.010000 2.090000 ;
        RECT 1.695000 1.295000 2.010000 1.920000 ;
    END
  END A1_N
  PIN A2_N
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.985000 1.210000 1.455000 1.750000 ;
    END
  END A2_N
  PIN B1
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.565000 1.345000 3.815000 1.920000 ;
        RECT 3.565000 1.920000 5.675000 2.090000 ;
        RECT 5.325000 1.295000 5.675000 1.920000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.995000 1.210000 5.155000 1.750000 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  0.991200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.900000 0.595000 3.230000 2.260000 ;
        RECT 2.900000 2.260000 4.550000 2.590000 ;
        RECT 2.900000 2.590000 3.230000 3.075000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 5.760000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 5.760000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.760000 0.085000 ;
      RECT 0.000000  3.245000 5.760000 3.415000 ;
      RECT 0.170000  0.085000 0.475000 1.205000 ;
      RECT 0.170000  2.270000 0.500000 3.245000 ;
      RECT 0.645000  0.305000 1.710000 0.660000 ;
      RECT 0.645000  0.660000 0.860000 1.090000 ;
      RECT 0.670000  2.260000 2.350000 2.430000 ;
      RECT 0.670000  2.430000 0.860000 3.075000 ;
      RECT 1.030000  0.830000 2.350000 1.040000 ;
      RECT 1.030000  2.600000 1.360000 3.245000 ;
      RECT 1.530000  2.430000 2.350000 2.450000 ;
      RECT 1.530000  2.450000 1.755000 3.075000 ;
      RECT 1.890000  0.085000 2.220000 0.660000 ;
      RECT 1.925000  2.620000 2.730000 3.245000 ;
      RECT 2.180000  1.040000 2.350000 1.375000 ;
      RECT 2.180000  1.375000 2.565000 1.625000 ;
      RECT 2.180000  1.625000 2.350000 2.260000 ;
      RECT 2.520000  0.255000 3.670000 0.425000 ;
      RECT 2.520000  0.425000 2.730000 1.205000 ;
      RECT 2.520000  1.815000 2.730000 2.620000 ;
      RECT 3.400000  2.760000 3.630000 3.245000 ;
      RECT 3.410000  0.425000 3.670000 0.870000 ;
      RECT 3.410000  0.870000 5.460000 1.040000 ;
      RECT 3.800000  2.760000 4.950000 3.075000 ;
      RECT 3.840000  0.085000 4.170000 0.700000 ;
      RECT 4.340000  0.325000 4.530000 0.870000 ;
      RECT 4.700000  0.085000 5.030000 0.700000 ;
      RECT 4.720000  2.260000 4.950000 2.760000 ;
      RECT 5.130000  2.260000 5.460000 3.245000 ;
      RECT 5.200000  0.325000 5.460000 0.870000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
  END
END sky130_fd_sc_lp__o2bb2ai_2
END LIBRARY
