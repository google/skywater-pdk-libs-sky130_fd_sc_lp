* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
M1000 a_302_367# a_27_508# Y VPB phighvt w=1.26e+06u l=150000u
+  ad=6.867e+11p pd=6.13e+06u as=3.339e+11p ps=3.05e+06u
M1001 VPWR B1_N a_27_508# VPB phighvt w=420000u l=150000u
+  ad=5.901e+11p pd=4.65e+06u as=1.113e+11p ps=1.37e+06u
M1002 VGND B1_N a_27_508# VNB nshort w=420000u l=150000u
+  ad=4.914e+11p pd=4.64e+06u as=1.113e+11p ps=1.37e+06u
M1003 a_302_367# A2 VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 Y a_27_508# VGND VNB nshort w=840000u l=150000u
+  ad=2.898e+11p pd=2.37e+06u as=0p ps=0u
M1005 a_380_47# A1 Y VNB nshort w=840000u l=150000u
+  ad=3.528e+11p pd=2.52e+06u as=0p ps=0u
M1006 VPWR A1 a_302_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND A2 a_380_47# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
