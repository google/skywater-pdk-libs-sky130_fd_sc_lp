# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__or3b_lp
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__or3b_lp ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.800000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.376000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.005000 1.035000 3.715000 1.410000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.376000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.810000 1.675000 3.715000 2.150000 ;
    END
  END B
  PIN C_N
    ANTENNAGATEAREA  0.376000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.445000 1.175000 0.835000 1.845000 ;
    END
  END C_N
  PIN X
    ANTENNADIFFAREA  0.404700 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.245000 2.075000 4.685000 2.890000 ;
        RECT 4.245000 2.890000 4.575000 3.065000 ;
        RECT 4.355000 0.440000 4.685000 0.945000 ;
        RECT 4.445000 0.945000 4.685000 2.075000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 4.800000 0.085000 ;
        RECT 0.905000  0.085000 1.235000 0.645000 ;
        RECT 1.875000  0.895000 2.405000 1.145000 ;
        RECT 2.235000  0.085000 2.405000 0.895000 ;
        RECT 3.565000  0.085000 3.895000 0.855000 ;
      LAYER mcon ;
        RECT 0.155000 -0.085000 0.325000 0.085000 ;
        RECT 0.635000 -0.085000 0.805000 0.085000 ;
        RECT 1.115000 -0.085000 1.285000 0.085000 ;
        RECT 1.595000 -0.085000 1.765000 0.085000 ;
        RECT 2.075000 -0.085000 2.245000 0.085000 ;
        RECT 2.555000 -0.085000 2.725000 0.085000 ;
        RECT 3.035000 -0.085000 3.205000 0.085000 ;
        RECT 3.515000 -0.085000 3.685000 0.085000 ;
        RECT 3.995000 -0.085000 4.165000 0.085000 ;
        RECT 4.475000 -0.085000 4.645000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.800000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.245000 4.800000 3.415000 ;
        RECT 0.645000 2.025000 0.975000 3.245000 ;
        RECT 3.605000 2.680000 3.935000 3.245000 ;
      LAYER mcon ;
        RECT 0.155000 3.245000 0.325000 3.415000 ;
        RECT 0.635000 3.245000 0.805000 3.415000 ;
        RECT 1.115000 3.245000 1.285000 3.415000 ;
        RECT 1.595000 3.245000 1.765000 3.415000 ;
        RECT 2.075000 3.245000 2.245000 3.415000 ;
        RECT 2.555000 3.245000 2.725000 3.415000 ;
        RECT 3.035000 3.245000 3.205000 3.415000 ;
        RECT 3.515000 3.245000 3.685000 3.415000 ;
        RECT 3.995000 3.245000 4.165000 3.415000 ;
        RECT 4.475000 3.245000 4.645000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 4.800000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.095000 0.265000 0.445000 0.825000 ;
      RECT 0.095000 0.825000 1.345000 0.995000 ;
      RECT 0.095000 0.995000 0.265000 2.025000 ;
      RECT 0.095000 2.025000 0.445000 3.065000 ;
      RECT 1.015000 0.995000 1.345000 1.450000 ;
      RECT 1.295000 1.845000 1.625000 2.895000 ;
      RECT 1.295000 2.895000 2.915000 3.065000 ;
      RECT 1.525000 0.265000 2.055000 0.675000 ;
      RECT 1.525000 0.675000 1.695000 1.325000 ;
      RECT 1.525000 1.325000 2.825000 1.495000 ;
      RECT 1.825000 1.495000 2.155000 2.715000 ;
      RECT 2.460000 1.495000 2.630000 2.330000 ;
      RECT 2.460000 2.330000 4.065000 2.500000 ;
      RECT 2.585000 2.680000 2.915000 2.895000 ;
      RECT 2.655000 0.485000 3.075000 0.855000 ;
      RECT 2.655000 0.855000 2.825000 1.325000 ;
      RECT 3.895000 1.225000 4.225000 1.895000 ;
      RECT 3.895000 1.895000 4.065000 2.330000 ;
  END
END sky130_fd_sc_lp__or3b_lp
