* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__mux2i_lp2 A0 A1 S VGND VNB VPB VPWR Y
X0 VPWR S a_148_419# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X1 a_148_419# A0 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X2 a_422_47# a_490_21# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 VGND S a_256_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 VGND S a_609_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 a_410_419# a_490_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X6 VPWR S a_490_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X7 Y A0 a_422_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 Y A1 a_410_419# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X9 a_609_47# S a_490_21# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 a_256_47# A1 Y VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
