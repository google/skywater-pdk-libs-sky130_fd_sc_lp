* File: sky130_fd_sc_lp__and3_m.pex.spice
* Created: Fri Aug 28 10:06:30 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__AND3_M%A 3 7 9 10 14
r24 14 17 83.3779 $w=4.9e-07 $l=5.05e-07 $layer=POLY_cond $X=0.425 $Y=1.005
+ $X2=0.425 $Y2=1.51
r25 14 16 46.2534 $w=4.9e-07 $l=1.65e-07 $layer=POLY_cond $X=0.425 $Y=1.005
+ $X2=0.425 $Y2=0.84
r26 14 15 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.345
+ $Y=1.005 $X2=0.345 $Y2=1.005
r27 10 15 12.153 $w=2.73e-07 $l=2.9e-07 $layer=LI1_cond $X=0.292 $Y=1.295
+ $X2=0.292 $Y2=1.005
r28 9 15 3.35256 $w=2.73e-07 $l=8e-08 $layer=LI1_cond $X=0.292 $Y=0.925
+ $X2=0.292 $Y2=1.005
r29 7 17 335.862 $w=1.5e-07 $l=6.55e-07 $layer=POLY_cond $X=0.595 $Y=2.165
+ $X2=0.595 $Y2=1.51
r30 3 16 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.595 $Y=0.445
+ $X2=0.595 $Y2=0.84
.ends

.subckt PM_SKY130_FD_SC_LP__AND3_M%B 3 6 9 10 11 12 13 14 19
r41 19 20 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.045
+ $Y=0.93 $X2=1.045 $Y2=0.93
r42 14 20 12.9428 $w=3.23e-07 $l=3.65e-07 $layer=LI1_cond $X=1.122 $Y=1.295
+ $X2=1.122 $Y2=0.93
r43 13 20 0.177299 $w=3.23e-07 $l=5e-09 $layer=LI1_cond $X=1.122 $Y=0.925
+ $X2=1.122 $Y2=0.93
r44 12 13 13.1201 $w=3.23e-07 $l=3.7e-07 $layer=LI1_cond $X=1.122 $Y=0.555
+ $X2=1.122 $Y2=0.925
r45 10 19 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.045 $Y=1.27
+ $X2=1.045 $Y2=0.93
r46 10 11 38.6168 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.045 $Y=1.27
+ $X2=1.045 $Y2=1.435
r47 9 19 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.045 $Y=0.765
+ $X2=1.045 $Y2=0.93
r48 6 11 374.319 $w=1.5e-07 $l=7.3e-07 $layer=POLY_cond $X=1.025 $Y=2.165
+ $X2=1.025 $Y2=1.435
r49 3 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.955 $Y=0.445
+ $X2=0.955 $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_LP__AND3_M%C 3 7 11 12 13 14 15 20
c46 3 0 2.49619e-19 $X=1.455 $Y=2.165
r47 20 23 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.585 $Y=1.32
+ $X2=1.585 $Y2=1.485
r48 20 22 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.585 $Y=1.32
+ $X2=1.585 $Y2=1.155
r49 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.585
+ $Y=1.32 $X2=1.585 $Y2=1.32
r50 15 21 15.0035 $w=2.63e-07 $l=3.45e-07 $layer=LI1_cond $X=1.632 $Y=1.665
+ $X2=1.632 $Y2=1.32
r51 14 21 1.08721 $w=2.63e-07 $l=2.5e-08 $layer=LI1_cond $X=1.632 $Y=1.295
+ $X2=1.632 $Y2=1.32
r52 13 14 16.0907 $w=2.63e-07 $l=3.7e-07 $layer=LI1_cond $X=1.632 $Y=0.925
+ $X2=1.632 $Y2=1.295
r53 11 12 53.9552 $w=1.9e-07 $l=1.5e-07 $layer=POLY_cond $X=1.475 $Y=1.675
+ $X2=1.475 $Y2=1.825
r54 11 23 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=1.495 $Y=1.675
+ $X2=1.495 $Y2=1.485
r55 7 22 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=1.495 $Y=0.445
+ $X2=1.495 $Y2=1.155
r56 3 12 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=1.455 $Y=2.165
+ $X2=1.455 $Y2=1.825
.ends

.subckt PM_SKY130_FD_SC_LP__AND3_M%A_51_47# 1 2 3 10 15 16 18 20 23 27 29 34 35
+ 36 37 38 40 50
r88 48 50 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=1.3 $Y=2.91 $X2=1.3
+ $Y2=2.82
r89 38 48 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.3
+ $Y=2.91 $X2=1.3 $Y2=2.91
r90 38 40 38.29 $w=2.08e-07 $l=7.25e-07 $layer=LI1_cond $X=1.24 $Y=2.825
+ $X2=1.24 $Y2=2.1
r91 37 44 14.1928 $w=2.1e-07 $l=2.4e-07 $layer=LI1_cond $X=1.24 $Y=2.04 $X2=1.24
+ $Y2=1.8
r92 37 40 3.16883 $w=2.08e-07 $l=6e-08 $layer=LI1_cond $X=1.24 $Y=2.04 $X2=1.24
+ $Y2=2.1
r93 35 44 1.129 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.135 $Y=1.8 $X2=1.24
+ $Y2=1.8
r94 35 36 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=1.135 $Y=1.8
+ $X2=0.78 $Y2=1.8
r95 34 36 6.25812 $w=3.56e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.695 $Y=1.715
+ $X2=0.78 $Y2=1.8
r96 34 42 10.7949 $w=3.56e-07 $l=4.2e-07 $layer=LI1_cond $X=0.695 $Y=1.715
+ $X2=0.38 $Y2=1.96
r97 33 34 68.8289 $w=1.68e-07 $l=1.055e-06 $layer=LI1_cond $X=0.695 $Y=0.66
+ $X2=0.695 $Y2=1.715
r98 29 33 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.61 $Y=0.495
+ $X2=0.695 $Y2=0.66
r99 29 31 8.03218 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=0.61 $Y=0.495
+ $X2=0.38 $Y2=0.495
r100 25 27 71.7872 $w=1.5e-07 $l=1.4e-07 $layer=POLY_cond $X=1.925 $Y=0.84
+ $X2=2.065 $Y2=0.84
r101 21 23 92.2979 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=1.885 $Y=1.77
+ $X2=2.065 $Y2=1.77
r102 20 23 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.065 $Y=1.695
+ $X2=2.065 $Y2=1.77
r103 19 27 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.065 $Y=0.915
+ $X2=2.065 $Y2=0.84
r104 19 20 399.957 $w=1.5e-07 $l=7.8e-07 $layer=POLY_cond $X=2.065 $Y=0.915
+ $X2=2.065 $Y2=1.695
r105 16 25 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.925 $Y=0.765
+ $X2=1.925 $Y2=0.84
r106 16 18 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.925 $Y=0.765
+ $X2=1.925 $Y2=0.445
r107 13 15 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=1.885 $Y=2.745
+ $X2=1.885 $Y2=2.165
r108 12 21 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.885 $Y=1.845
+ $X2=1.885 $Y2=1.77
r109 12 15 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.885 $Y=1.845
+ $X2=1.885 $Y2=2.165
r110 11 50 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.465 $Y=2.82
+ $X2=1.3 $Y2=2.82
r111 10 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.81 $Y=2.82
+ $X2=1.885 $Y2=2.745
r112 10 11 176.904 $w=1.5e-07 $l=3.45e-07 $layer=POLY_cond $X=1.81 $Y=2.82
+ $X2=1.465 $Y2=2.82
r113 3 40 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.1
+ $Y=1.955 $X2=1.24 $Y2=2.1
r114 2 42 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.255
+ $Y=1.955 $X2=0.38 $Y2=2.1
r115 1 31 182 $w=1.7e-07 $l=3.16386e-07 $layer=licon1_NDIFF $count=1 $X=0.255
+ $Y=0.235 $X2=0.38 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__AND3_M%VPWR 1 2 9 11 14 15 16 18 21 29 30 33
c40 18 0 1.63777e-19 $X=1.67 $Y=2.23
r41 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r42 30 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r43 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r44 27 33 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.815 $Y=3.33
+ $X2=1.73 $Y2=3.33
r45 27 29 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.815 $Y=3.33
+ $X2=2.16 $Y2=3.33
r46 24 25 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r47 21 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r48 21 25 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r49 18 20 8.79328 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=1.69 $Y=2.23
+ $X2=1.69 $Y2=2.395
r50 15 24 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=0.725 $Y=3.33
+ $X2=0.72 $Y2=3.33
r51 15 16 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=0.725 $Y=3.33
+ $X2=0.82 $Y2=3.33
r52 14 33 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.73 $Y=3.245
+ $X2=1.73 $Y2=3.33
r53 14 20 55.4545 $w=1.68e-07 $l=8.5e-07 $layer=LI1_cond $X=1.73 $Y=3.245
+ $X2=1.73 $Y2=2.395
r54 12 16 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=0.915 $Y=3.33
+ $X2=0.82 $Y2=3.33
r55 11 33 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.645 $Y=3.33
+ $X2=1.73 $Y2=3.33
r56 11 12 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=1.645 $Y=3.33
+ $X2=0.915 $Y2=3.33
r57 7 16 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=0.82 $Y=3.245
+ $X2=0.82 $Y2=3.33
r58 7 9 59.2488 $w=1.88e-07 $l=1.015e-06 $layer=LI1_cond $X=0.82 $Y=3.245
+ $X2=0.82 $Y2=2.23
r59 2 18 600 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=1 $X=1.53
+ $Y=1.955 $X2=1.67 $Y2=2.23
r60 1 9 600 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=1 $X=0.67
+ $Y=1.955 $X2=0.81 $Y2=2.23
.ends

.subckt PM_SKY130_FD_SC_LP__AND3_M%X 1 2 7 8 9 10 11 12 13
c19 7 0 8.58422e-20 $X=2.16 $Y=0.555
r20 12 13 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=2.12 $Y=2.405
+ $X2=2.12 $Y2=2.775
r21 11 12 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=2.12 $Y=2.035
+ $X2=2.12 $Y2=2.405
r22 10 11 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=2.12 $Y=1.665
+ $X2=2.12 $Y2=2.035
r23 9 10 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=2.12 $Y=1.295
+ $X2=2.12 $Y2=1.665
r24 8 9 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=2.12 $Y=0.925 $X2=2.12
+ $Y2=1.295
r25 7 8 19.1306 $w=2.48e-07 $l=4.15e-07 $layer=LI1_cond $X=2.12 $Y=0.51 $X2=2.12
+ $Y2=0.925
r26 2 11 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.96
+ $Y=1.955 $X2=2.1 $Y2=2.1
r27 1 7 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=2 $Y=0.235
+ $X2=2.14 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_LP__AND3_M%VGND 1 6 8 10 17 18 21
r31 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r32 18 22 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.68
+ $Y2=0
r33 17 18 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r34 15 21 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.815 $Y=0 $X2=1.71
+ $Y2=0
r35 15 17 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.815 $Y=0 $X2=2.16
+ $Y2=0
r36 12 13 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r37 10 21 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.605 $Y=0 $X2=1.71
+ $Y2=0
r38 10 12 89.0535 $w=1.68e-07 $l=1.365e-06 $layer=LI1_cond $X=1.605 $Y=0
+ $X2=0.24 $Y2=0
r39 8 22 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r40 8 13 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.24
+ $Y2=0
r41 4 21 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=1.71 $Y=0.085
+ $X2=1.71 $Y2=0
r42 4 6 15.5801 $w=2.08e-07 $l=2.95e-07 $layer=LI1_cond $X=1.71 $Y=0.085
+ $X2=1.71 $Y2=0.38
r43 1 6 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=1.57
+ $Y=0.235 $X2=1.71 $Y2=0.38
.ends

