* File: sky130_fd_sc_lp__a22oi_m.pxi.spice
* Created: Wed Sep  2 09:23:29 2020
* 
x_PM_SKY130_FD_SC_LP__A22OI_M%B2 N_B2_c_56_n N_B2_M1007_g N_B2_M1005_g
+ N_B2_c_58_n N_B2_c_59_n N_B2_c_64_n B2 B2 B2 B2 B2 N_B2_c_61_n
+ PM_SKY130_FD_SC_LP__A22OI_M%B2
x_PM_SKY130_FD_SC_LP__A22OI_M%B1 N_B1_M1003_g N_B1_c_94_n N_B1_M1006_g
+ N_B1_c_96_n B1 B1 B1 B1 N_B1_c_98_n PM_SKY130_FD_SC_LP__A22OI_M%B1
x_PM_SKY130_FD_SC_LP__A22OI_M%A1 N_A1_M1002_g N_A1_c_133_n N_A1_M1001_g
+ N_A1_c_138_n A1 A1 A1 A1 A1 N_A1_c_135_n PM_SKY130_FD_SC_LP__A22OI_M%A1
x_PM_SKY130_FD_SC_LP__A22OI_M%A2 N_A2_M1004_g N_A2_c_183_n N_A2_M1000_g
+ N_A2_c_178_n N_A2_c_179_n N_A2_c_185_n N_A2_c_180_n A2 A2 A2 A2 N_A2_c_182_n
+ PM_SKY130_FD_SC_LP__A22OI_M%A2
x_PM_SKY130_FD_SC_LP__A22OI_M%A_39_496# N_A_39_496#_M1005_s N_A_39_496#_M1006_d
+ N_A_39_496#_M1000_d N_A_39_496#_c_212_n N_A_39_496#_c_213_n
+ N_A_39_496#_c_214_n N_A_39_496#_c_238_p N_A_39_496#_c_215_n
+ PM_SKY130_FD_SC_LP__A22OI_M%A_39_496#
x_PM_SKY130_FD_SC_LP__A22OI_M%Y N_Y_M1003_d N_Y_M1005_d N_Y_c_246_n N_Y_c_243_n
+ Y PM_SKY130_FD_SC_LP__A22OI_M%Y
x_PM_SKY130_FD_SC_LP__A22OI_M%VPWR N_VPWR_M1001_d N_VPWR_c_273_n VPWR
+ N_VPWR_c_274_n N_VPWR_c_275_n N_VPWR_c_272_n N_VPWR_c_277_n
+ PM_SKY130_FD_SC_LP__A22OI_M%VPWR
x_PM_SKY130_FD_SC_LP__A22OI_M%VGND N_VGND_M1007_s N_VGND_M1004_d N_VGND_c_297_n
+ N_VGND_c_298_n N_VGND_c_299_n N_VGND_c_300_n VGND N_VGND_c_301_n
+ N_VGND_c_302_n PM_SKY130_FD_SC_LP__A22OI_M%VGND
cc_1 VNB N_B2_c_56_n 0.00457352f $X=-0.19 $Y=-0.245 $X2=0.36 $Y2=1.75
cc_2 VNB N_B2_M1007_g 0.0302642f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=0.445
cc_3 VNB N_B2_c_58_n 0.0399363f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=0.995
cc_4 VNB N_B2_c_59_n 0.0249762f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.59
cc_5 VNB B2 0.00859675f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_6 VNB N_B2_c_61_n 0.0372496f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.085
cc_7 VNB N_B1_M1003_g 0.0208857f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=0.92
cc_8 VNB N_B1_c_94_n 0.0228547f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_B1_M1006_g 0.0072981f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=2.69
cc_10 VNB N_B1_c_96_n 0.0193017f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=0.995
cc_11 VNB B1 0.00888916f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.07
cc_12 VNB N_B1_c_98_n 0.0156795f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A1_M1002_g 0.0414809f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=0.92
cc_14 VNB N_A1_c_133_n 0.0115169f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB A1 0.00781335f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.07
cc_16 VNB N_A1_c_135_n 0.0156833f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_17 VNB N_A2_M1004_g 0.0318009f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=0.92
cc_18 VNB N_A2_c_178_n 0.00396825f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=2.69
cc_19 VNB N_A2_c_179_n 0.0402198f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A2_c_180_n 0.0234333f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.825
cc_21 VNB A2 0.00797133f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A2_c_182_n 0.0378399f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_Y_c_243_n 0.00522729f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=2.69
cc_24 VNB Y 0.0128806f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.07
cc_25 VNB N_VPWR_c_272_n 0.103974f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_297_n 0.0134838f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.9
cc_27 VNB N_VGND_c_298_n 0.00485511f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=2.69
cc_28 VNB N_VGND_c_299_n 0.0125039f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=0.995
cc_29 VNB N_VGND_c_300_n 0.015566f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_301_n 0.0412005f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.59
cc_31 VNB N_VGND_c_302_n 0.15203f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VPB N_B2_c_56_n 0.00431409f $X=-0.19 $Y=1.655 $X2=0.36 $Y2=1.75
cc_33 VPB N_B2_M1005_g 0.0418541f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=2.69
cc_34 VPB N_B2_c_64_n 0.0332691f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.825
cc_35 VPB B2 0.0368417f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_36 VPB N_B1_M1006_g 0.0495099f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=2.69
cc_37 VPB B1 0.00970151f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.07
cc_38 VPB N_A1_c_133_n 0.0104351f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_39 VPB N_A1_M1001_g 0.0357933f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=2.69
cc_40 VPB N_A1_c_138_n 0.0163803f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=0.995
cc_41 VPB A1 0.00535083f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.07
cc_42 VPB N_A2_c_183_n 0.020215f $X=-0.19 $Y=1.655 $X2=0.59 $Y2=0.445
cc_43 VPB N_A2_c_178_n 0.038344f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=2.69
cc_44 VPB N_A2_c_185_n 0.0251077f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.59
cc_45 VPB A2 0.0172796f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_46 VPB N_A_39_496#_c_212_n 0.00808721f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_47 VPB N_A_39_496#_c_213_n 0.0136673f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.425
cc_48 VPB N_A_39_496#_c_214_n 0.00540395f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.59
cc_49 VPB N_A_39_496#_c_215_n 0.0188356f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_50 VPB Y 0.0130321f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.07
cc_51 VPB N_VPWR_c_273_n 0.00777104f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_52 VPB N_VPWR_c_274_n 0.0404542f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_53 VPB N_VPWR_c_275_n 0.0178394f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.825
cc_54 VPB N_VPWR_c_272_n 0.0660237f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_55 VPB N_VPWR_c_277_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_56 N_B2_M1007_g N_B1_M1003_g 0.0304551f $X=0.59 $Y=0.445 $X2=0 $Y2=0
cc_57 N_B2_c_61_n N_B1_c_94_n 0.00357325f $X=0.27 $Y=1.085 $X2=0 $Y2=0
cc_58 N_B2_c_59_n N_B1_M1006_g 0.00218954f $X=0.27 $Y=1.59 $X2=0 $Y2=0
cc_59 N_B2_c_64_n N_B1_M1006_g 0.0421312f $X=0.635 $Y=1.825 $X2=0 $Y2=0
cc_60 N_B2_c_59_n N_B1_c_96_n 0.00357325f $X=0.27 $Y=1.59 $X2=0 $Y2=0
cc_61 N_B2_M1007_g B1 2.01599e-19 $X=0.59 $Y=0.445 $X2=0 $Y2=0
cc_62 N_B2_c_64_n B1 0.00111375f $X=0.635 $Y=1.825 $X2=0 $Y2=0
cc_63 N_B2_c_58_n N_B1_c_98_n 0.0304551f $X=0.59 $Y=0.995 $X2=0 $Y2=0
cc_64 B2 N_A_39_496#_M1005_s 0.00196532f $X=0.155 $Y=0.84 $X2=-0.19 $Y2=-0.245
cc_65 N_B2_M1005_g N_A_39_496#_c_212_n 0.012045f $X=0.635 $Y=2.69 $X2=0 $Y2=0
cc_66 N_B2_M1005_g N_A_39_496#_c_215_n 0.00124499f $X=0.635 $Y=2.69 $X2=0 $Y2=0
cc_67 B2 N_A_39_496#_c_215_n 0.0143889f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_68 N_B2_M1007_g N_Y_c_246_n 0.0120061f $X=0.59 $Y=0.445 $X2=0 $Y2=0
cc_69 N_B2_M1007_g Y 0.0100684f $X=0.59 $Y=0.445 $X2=0 $Y2=0
cc_70 N_B2_M1005_g Y 0.024889f $X=0.635 $Y=2.69 $X2=0 $Y2=0
cc_71 N_B2_c_58_n Y 0.00515365f $X=0.59 $Y=0.995 $X2=0 $Y2=0
cc_72 N_B2_c_64_n Y 0.00698754f $X=0.635 $Y=1.825 $X2=0 $Y2=0
cc_73 B2 Y 0.0876116f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_74 N_B2_c_61_n Y 0.00459224f $X=0.27 $Y=1.085 $X2=0 $Y2=0
cc_75 N_B2_M1005_g N_VPWR_c_274_n 8.70008e-19 $X=0.635 $Y=2.69 $X2=0 $Y2=0
cc_76 B2 N_VPWR_c_272_n 0.0011335f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_77 N_B2_M1007_g N_VGND_c_298_n 0.00654365f $X=0.59 $Y=0.445 $X2=0 $Y2=0
cc_78 N_B2_c_58_n N_VGND_c_298_n 0.00357108f $X=0.59 $Y=0.995 $X2=0 $Y2=0
cc_79 B2 N_VGND_c_298_n 0.00631716f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_80 N_B2_M1007_g N_VGND_c_301_n 0.00507464f $X=0.59 $Y=0.445 $X2=0 $Y2=0
cc_81 N_B2_M1007_g N_VGND_c_302_n 0.00966711f $X=0.59 $Y=0.445 $X2=0 $Y2=0
cc_82 B2 N_VGND_c_302_n 0.00390326f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_83 N_B1_M1003_g N_A1_M1002_g 0.0159426f $X=0.95 $Y=0.445 $X2=0 $Y2=0
cc_84 B1 N_A1_M1002_g 0.00889198f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_85 N_B1_c_98_n N_A1_M1002_g 0.0133344f $X=1.045 $Y=1.005 $X2=0 $Y2=0
cc_86 N_B1_M1006_g N_A1_c_133_n 0.0502966f $X=1.065 $Y=2.69 $X2=0 $Y2=0
cc_87 N_B1_c_96_n N_A1_c_133_n 0.0133344f $X=1.042 $Y=1.51 $X2=0 $Y2=0
cc_88 N_B1_M1003_g A1 9.57474e-19 $X=0.95 $Y=0.445 $X2=0 $Y2=0
cc_89 N_B1_M1006_g A1 5.542e-19 $X=1.065 $Y=2.69 $X2=0 $Y2=0
cc_90 B1 A1 0.0819142f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_91 N_B1_c_98_n A1 6.46197e-19 $X=1.045 $Y=1.005 $X2=0 $Y2=0
cc_92 N_B1_c_94_n N_A1_c_135_n 0.0133344f $X=1.042 $Y=1.343 $X2=0 $Y2=0
cc_93 N_B1_M1006_g N_A_39_496#_c_212_n 0.0128998f $X=1.065 $Y=2.69 $X2=0 $Y2=0
cc_94 N_B1_M1006_g N_A_39_496#_c_214_n 0.0013183f $X=1.065 $Y=2.69 $X2=0 $Y2=0
cc_95 B1 N_A_39_496#_c_214_n 0.00742998f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_96 N_B1_M1003_g N_Y_c_243_n 0.0143212f $X=0.95 $Y=0.445 $X2=0 $Y2=0
cc_97 B1 N_Y_c_243_n 0.024105f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_98 N_B1_c_98_n N_Y_c_243_n 0.00134056f $X=1.045 $Y=1.005 $X2=0 $Y2=0
cc_99 N_B1_M1003_g Y 0.010907f $X=0.95 $Y=0.445 $X2=0 $Y2=0
cc_100 N_B1_M1006_g Y 0.0127807f $X=1.065 $Y=2.69 $X2=0 $Y2=0
cc_101 B1 Y 0.0985885f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_102 N_B1_M1006_g N_VPWR_c_274_n 8.70008e-19 $X=1.065 $Y=2.69 $X2=0 $Y2=0
cc_103 N_B1_M1003_g N_VGND_c_301_n 0.00373071f $X=0.95 $Y=0.445 $X2=0 $Y2=0
cc_104 N_B1_M1003_g N_VGND_c_302_n 0.00559034f $X=0.95 $Y=0.445 $X2=0 $Y2=0
cc_105 B1 N_VGND_c_302_n 0.00106056f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_106 N_A1_M1002_g N_A2_M1004_g 0.0587801f $X=1.495 $Y=0.445 $X2=0 $Y2=0
cc_107 A1 N_A2_M1004_g 0.00766094f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_108 N_A1_c_133_n N_A2_c_178_n 0.0196f $X=1.587 $Y=1.813 $X2=0 $Y2=0
cc_109 N_A1_M1001_g N_A2_c_178_n 0.00662288f $X=1.495 $Y=2.69 $X2=0 $Y2=0
cc_110 A1 N_A2_c_178_n 0.0034028f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_111 N_A1_M1001_g N_A2_c_185_n 0.0226309f $X=1.495 $Y=2.69 $X2=0 $Y2=0
cc_112 N_A1_c_133_n N_A2_c_180_n 0.00876259f $X=1.587 $Y=1.813 $X2=0 $Y2=0
cc_113 N_A1_M1002_g A2 3.14547e-19 $X=1.495 $Y=0.445 $X2=0 $Y2=0
cc_114 A1 A2 0.0663925f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_115 N_A1_c_135_n A2 7.66262e-19 $X=1.59 $Y=1.475 $X2=0 $Y2=0
cc_116 N_A1_M1002_g N_A2_c_182_n 0.0063482f $X=1.495 $Y=0.445 $X2=0 $Y2=0
cc_117 A1 N_A2_c_182_n 0.00389542f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_118 N_A1_c_135_n N_A2_c_182_n 0.00876259f $X=1.59 $Y=1.475 $X2=0 $Y2=0
cc_119 N_A1_M1001_g N_A_39_496#_c_212_n 0.00111521f $X=1.495 $Y=2.69 $X2=0 $Y2=0
cc_120 N_A1_M1001_g N_A_39_496#_c_213_n 0.013717f $X=1.495 $Y=2.69 $X2=0 $Y2=0
cc_121 N_A1_c_138_n N_A_39_496#_c_213_n 9.03173e-19 $X=1.587 $Y=1.98 $X2=0 $Y2=0
cc_122 A1 N_A_39_496#_c_213_n 0.0188853f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_123 N_A1_M1002_g N_Y_c_243_n 0.00374285f $X=1.495 $Y=0.445 $X2=0 $Y2=0
cc_124 A1 N_Y_c_243_n 0.0119446f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_125 N_A1_M1001_g N_VPWR_c_273_n 0.00608121f $X=1.495 $Y=2.69 $X2=0 $Y2=0
cc_126 N_A1_M1001_g N_VPWR_c_274_n 0.00444095f $X=1.495 $Y=2.69 $X2=0 $Y2=0
cc_127 N_A1_M1001_g N_VPWR_c_272_n 0.00442501f $X=1.495 $Y=2.69 $X2=0 $Y2=0
cc_128 N_A1_M1002_g N_VGND_c_301_n 0.00505689f $X=1.495 $Y=0.445 $X2=0 $Y2=0
cc_129 A1 N_VGND_c_301_n 0.00604823f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_130 N_A1_M1002_g N_VGND_c_302_n 0.00884089f $X=1.495 $Y=0.445 $X2=0 $Y2=0
cc_131 A1 N_VGND_c_302_n 0.00849221f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_132 A1 A_314_47# 0.00139886f $X=1.595 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_133 N_A2_c_183_n N_A_39_496#_c_213_n 0.00831432f $X=1.925 $Y=2.37 $X2=0 $Y2=0
cc_134 N_A2_c_185_n N_A_39_496#_c_213_n 0.0148221f $X=2.07 $Y=2.295 $X2=0 $Y2=0
cc_135 A2 N_A_39_496#_c_213_n 0.0151121f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_136 N_A2_c_183_n N_VPWR_c_273_n 0.0140831f $X=1.925 $Y=2.37 $X2=0 $Y2=0
cc_137 N_A2_c_183_n N_VPWR_c_275_n 0.00444095f $X=1.925 $Y=2.37 $X2=0 $Y2=0
cc_138 N_A2_c_183_n N_VPWR_c_272_n 0.00442501f $X=1.925 $Y=2.37 $X2=0 $Y2=0
cc_139 N_A2_M1004_g N_VGND_c_300_n 0.00491682f $X=1.855 $Y=0.445 $X2=0 $Y2=0
cc_140 N_A2_c_179_n N_VGND_c_300_n 0.0049813f $X=2.13 $Y=1.07 $X2=0 $Y2=0
cc_141 A2 N_VGND_c_300_n 0.00930502f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_142 N_A2_M1004_g N_VGND_c_301_n 0.00585385f $X=1.855 $Y=0.445 $X2=0 $Y2=0
cc_143 N_A2_M1004_g N_VGND_c_302_n 0.0114683f $X=1.855 $Y=0.445 $X2=0 $Y2=0
cc_144 A2 N_VGND_c_302_n 0.00107888f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_145 N_A_39_496#_c_212_n N_Y_M1005_d 0.00180746f $X=1.195 $Y=2.975 $X2=0 $Y2=0
cc_146 N_A_39_496#_c_212_n Y 0.0172718f $X=1.195 $Y=2.975 $X2=0 $Y2=0
cc_147 N_A_39_496#_c_214_n Y 0.013494f $X=1.365 $Y=2.405 $X2=0 $Y2=0
cc_148 N_A_39_496#_c_213_n N_VPWR_M1001_d 0.00178209f $X=2.055 $Y=2.405
+ $X2=-0.19 $Y2=1.655
cc_149 N_A_39_496#_c_212_n N_VPWR_c_273_n 0.0133632f $X=1.195 $Y=2.975 $X2=0
+ $Y2=0
cc_150 N_A_39_496#_c_213_n N_VPWR_c_273_n 0.0159264f $X=2.055 $Y=2.405 $X2=0
+ $Y2=0
cc_151 N_A_39_496#_c_212_n N_VPWR_c_274_n 0.0517471f $X=1.195 $Y=2.975 $X2=0
+ $Y2=0
cc_152 N_A_39_496#_c_215_n N_VPWR_c_274_n 0.0206108f $X=0.34 $Y=2.775 $X2=0
+ $Y2=0
cc_153 N_A_39_496#_c_238_p N_VPWR_c_275_n 0.00439013f $X=2.14 $Y=2.625 $X2=0
+ $Y2=0
cc_154 N_A_39_496#_c_212_n N_VPWR_c_272_n 0.0322666f $X=1.195 $Y=2.975 $X2=0
+ $Y2=0
cc_155 N_A_39_496#_c_213_n N_VPWR_c_272_n 0.0126337f $X=2.055 $Y=2.405 $X2=0
+ $Y2=0
cc_156 N_A_39_496#_c_238_p N_VPWR_c_272_n 0.00601105f $X=2.14 $Y=2.625 $X2=0
+ $Y2=0
cc_157 N_A_39_496#_c_215_n N_VPWR_c_272_n 0.0124745f $X=0.34 $Y=2.775 $X2=0
+ $Y2=0
cc_158 N_Y_c_246_n N_VGND_c_298_n 0.0162495f $X=0.78 $Y=0.495 $X2=0 $Y2=0
cc_159 N_Y_c_246_n N_VGND_c_301_n 0.00665067f $X=0.78 $Y=0.495 $X2=0 $Y2=0
cc_160 N_Y_c_243_n N_VGND_c_301_n 0.0193476f $X=1.165 $Y=0.495 $X2=0 $Y2=0
cc_161 N_Y_M1003_d N_VGND_c_302_n 0.00806684f $X=1.025 $Y=0.235 $X2=0 $Y2=0
cc_162 N_Y_c_246_n N_VGND_c_302_n 0.00609033f $X=0.78 $Y=0.495 $X2=0 $Y2=0
cc_163 N_Y_c_243_n N_VGND_c_302_n 0.0171629f $X=1.165 $Y=0.495 $X2=0 $Y2=0
cc_164 N_Y_c_246_n A_133_47# 6.6248e-19 $X=0.78 $Y=0.495 $X2=-0.19 $Y2=-0.245
cc_165 N_Y_c_243_n A_133_47# 4.13878e-19 $X=1.165 $Y=0.495 $X2=-0.19 $Y2=-0.245
cc_166 N_VGND_c_302_n A_133_47# 0.00173518f $X=2.16 $Y=0 $X2=-0.19 $Y2=-0.245
cc_167 N_VGND_c_302_n A_314_47# 0.00251844f $X=2.16 $Y=0 $X2=-0.19 $Y2=-0.245
