* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
X0 a_80_246# A1 a_480_56# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X1 VGND B2 a_294_56# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X2 X a_80_246# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X3 a_80_246# B1 a_217_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X4 a_480_56# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X5 VPWR A2 a_217_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X6 X a_80_246# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X7 a_217_367# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X8 a_217_367# B2 a_80_246# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X9 a_294_56# B1 a_80_246# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
.ends
