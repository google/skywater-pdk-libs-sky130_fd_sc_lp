* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__a2bb2oi_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
X0 a_459_39# A1_N VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X1 VGND A2_N a_459_39# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X2 a_30_367# a_459_39# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X3 VPWR B1 a_30_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X4 VPWR B2 a_30_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X5 a_113_65# B2 Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X6 Y B2 a_113_65# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X7 a_30_367# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X8 Y a_459_39# a_30_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X9 a_113_65# B1 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X10 VPWR A1_N a_699_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X11 a_30_367# B2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X12 a_699_367# A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X13 VGND a_459_39# Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X14 Y a_459_39# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X15 a_459_39# A2_N VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X16 VGND A1_N a_459_39# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X17 a_459_39# A2_N a_699_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X18 a_699_367# A2_N a_459_39# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X19 VGND B1 a_113_65# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
.ends
