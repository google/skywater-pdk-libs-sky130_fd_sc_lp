* File: sky130_fd_sc_lp__o32ai_4.spice
* Created: Fri Aug 28 11:18:33 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__o32ai_4.pex.spice"
.subckt sky130_fd_sc_lp__o32ai_4  VNB VPB B2 B1 A3 A2 A1 Y VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Y	Y
* A1	A1
* A2	A2
* A3	A3
* B1	B1
* B2	B2
* VPB	VPB
* VNB	VNB
MM1003 N_Y_M1003_d N_B2_M1003_g N_A_30_47#_M1003_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75009.5 A=0.126 P=1.98 MULT=1
MM1018 N_Y_M1003_d N_B2_M1018_g N_A_30_47#_M1018_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75009.1 A=0.126 P=1.98 MULT=1
MM1020 N_Y_M1020_d N_B2_M1020_g N_A_30_47#_M1018_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.1
+ SB=75008.6 A=0.126 P=1.98 MULT=1
MM1027 N_Y_M1020_d N_B2_M1027_g N_A_30_47#_M1027_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.5
+ SB=75008.2 A=0.126 P=1.98 MULT=1
MM1001 N_Y_M1001_d N_B1_M1001_g N_A_30_47#_M1027_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.9
+ SB=75007.8 A=0.126 P=1.98 MULT=1
MM1015 N_Y_M1001_d N_B1_M1015_g N_A_30_47#_M1015_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002.3
+ SB=75007.3 A=0.126 P=1.98 MULT=1
MM1024 N_Y_M1024_d N_B1_M1024_g N_A_30_47#_M1015_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002.8
+ SB=75006.9 A=0.126 P=1.98 MULT=1
MM1039 N_Y_M1024_d N_B1_M1039_g N_A_30_47#_M1039_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1638 PD=1.12 PS=1.23 NRD=0 NRS=0 M=1 R=5.6 SA=75003.2
+ SB=75006.5 A=0.126 P=1.98 MULT=1
MM1009 N_VGND_M1009_d N_A3_M1009_g N_A_30_47#_M1039_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1638 PD=1.12 PS=1.23 NRD=0 NRS=15.708 M=1 R=5.6 SA=75003.7
+ SB=75005.9 A=0.126 P=1.98 MULT=1
MM1021 N_VGND_M1009_d N_A3_M1021_g N_A_30_47#_M1021_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.147 PD=1.12 PS=1.19 NRD=0 NRS=4.992 M=1 R=5.6 SA=75004.2
+ SB=75005.5 A=0.126 P=1.98 MULT=1
MM1031 N_VGND_M1031_d N_A3_M1031_g N_A_30_47#_M1021_s VNB NSHORT L=0.15 W=0.84
+ AD=0.147 AS=0.147 PD=1.19 PS=1.19 NRD=9.996 NRS=4.992 M=1 R=5.6 SA=75004.7
+ SB=75005 A=0.126 P=1.98 MULT=1
MM1034 N_VGND_M1031_d N_A3_M1034_g N_A_30_47#_M1034_s VNB NSHORT L=0.15 W=0.84
+ AD=0.147 AS=0.3129 PD=1.19 PS=1.585 NRD=0 NRS=22.848 M=1 R=5.6 SA=75005.2
+ SB=75004.5 A=0.126 P=1.98 MULT=1
MM1004 N_VGND_M1004_d N_A2_M1004_g N_A_30_47#_M1034_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.3129 PD=1.12 PS=1.585 NRD=0 NRS=43.56 M=1 R=5.6 SA=75006.1
+ SB=75003.6 A=0.126 P=1.98 MULT=1
MM1010 N_VGND_M1004_d N_A2_M1010_g N_A_30_47#_M1010_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75006.5
+ SB=75003.2 A=0.126 P=1.98 MULT=1
MM1019 N_VGND_M1019_d N_A2_M1019_g N_A_30_47#_M1010_s VNB NSHORT L=0.15 W=0.84
+ AD=0.273 AS=0.1176 PD=1.49 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75006.9 SB=75002.8
+ A=0.126 P=1.98 MULT=1
MM1032 N_VGND_M1019_d N_A2_M1032_g N_A_30_47#_M1032_s VNB NSHORT L=0.15 W=0.84
+ AD=0.273 AS=0.1365 PD=1.49 PS=1.165 NRD=0 NRS=0 M=1 R=5.6 SA=75007.7 SB=75002
+ A=0.126 P=1.98 MULT=1
MM1007 N_A_30_47#_M1032_s N_A1_M1007_g N_VGND_M1007_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1365 AS=0.1176 PD=1.165 PS=1.12 NRD=6.42 NRS=0 M=1 R=5.6 SA=75008.2
+ SB=75001.5 A=0.126 P=1.98 MULT=1
MM1011 N_A_30_47#_M1011_d N_A1_M1011_g N_VGND_M1007_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75008.6
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1035 N_A_30_47#_M1011_d N_A1_M1035_g N_VGND_M1035_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75009.1
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1036 N_A_30_47#_M1036_d N_A1_M1036_g N_VGND_M1035_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75009.5
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1006 N_A_30_367#_M1006_d N_B2_M1006_g N_Y_M1006_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75003.2 A=0.189 P=2.82 MULT=1
MM1014 N_A_30_367#_M1014_d N_B2_M1014_g N_Y_M1006_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75002.8 A=0.189 P=2.82 MULT=1
MM1025 N_A_30_367#_M1014_d N_B2_M1025_g N_Y_M1025_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75002.4 A=0.189 P=2.82 MULT=1
MM1028 N_A_30_367#_M1028_d N_B2_M1028_g N_Y_M1025_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.19845 AS=0.1764 PD=1.575 PS=1.54 NRD=5.4569 NRS=0 M=1 R=8.4 SA=75001.5
+ SB=75001.9 A=0.189 P=2.82 MULT=1
MM1013 N_VPWR_M1013_d N_B1_M1013_g N_A_30_367#_M1028_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.19845 PD=1.54 PS=1.575 NRD=0 NRS=0 M=1 R=8.4 SA=75001.9
+ SB=75001.5 A=0.189 P=2.82 MULT=1
MM1023 N_VPWR_M1013_d N_B1_M1023_g N_A_30_367#_M1023_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.4
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1029 N_VPWR_M1029_d N_B1_M1029_g N_A_30_367#_M1023_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.8
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1037 N_VPWR_M1029_d N_B1_M1037_g N_A_30_367#_M1037_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75003.2
+ SB=75000.2 A=0.189 P=2.82 MULT=1
MM1002 N_Y_M1002_d N_A3_M1002_g N_A_829_349#_M1002_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75003.2 A=0.189 P=2.82 MULT=1
MM1008 N_Y_M1002_d N_A3_M1008_g N_A_829_349#_M1008_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75002.8 A=0.189 P=2.82 MULT=1
MM1030 N_Y_M1030_d N_A3_M1030_g N_A_829_349#_M1008_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75002.3 A=0.189 P=2.82 MULT=1
MM1033 N_Y_M1030_d N_A3_M1033_g N_A_829_349#_M1033_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.5
+ SB=75001.9 A=0.189 P=2.82 MULT=1
MM1005 N_A_829_349#_M1033_s N_A2_M1005_g N_A_1256_349#_M1005_s VPB PHIGHVT
+ L=0.15 W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75001.9 SB=75001.5 A=0.189 P=2.82 MULT=1
MM1016 N_A_829_349#_M1016_d N_A2_M1016_g N_A_1256_349#_M1005_s VPB PHIGHVT
+ L=0.15 W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75002.3 SB=75001.1 A=0.189 P=2.82 MULT=1
MM1022 N_A_829_349#_M1016_d N_A2_M1022_g N_A_1256_349#_M1022_s VPB PHIGHVT
+ L=0.15 W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75002.8 SB=75000.6 A=0.189 P=2.82 MULT=1
MM1038 N_A_829_349#_M1038_d N_A2_M1038_g N_A_1256_349#_M1022_s VPB PHIGHVT
+ L=0.15 W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75003.2 SB=75000.2 A=0.189 P=2.82 MULT=1
MM1000 N_VPWR_M1000_d N_A1_M1000_g N_A_1256_349#_M1000_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75001.5 A=0.189 P=2.82 MULT=1
MM1012 N_VPWR_M1012_d N_A1_M1012_g N_A_1256_349#_M1000_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1017 N_VPWR_M1012_d N_A1_M1017_g N_A_1256_349#_M1017_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1026 N_VPWR_M1026_d N_A1_M1026_g N_A_1256_349#_M1017_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.5
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX40_noxref VNB VPB NWDIODE A=20.7676 P=25.79
*
.include "sky130_fd_sc_lp__o32ai_4.pxi.spice"
*
.ends
*
*
