* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__o311a_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
X0 VGND A3 a_731_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X1 a_1196_367# A2 a_910_345# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X2 a_731_47# B1 a_476_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X3 VPWR C1 a_81_23# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X4 a_81_23# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X5 a_910_345# A2 a_1196_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X6 a_731_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X7 VGND A2 a_731_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X8 a_476_47# C1 a_81_23# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X9 a_731_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X10 a_81_23# C1 a_476_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X11 VPWR a_81_23# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X12 a_476_47# B1 a_731_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X13 X a_81_23# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X14 VPWR A1 a_1196_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X15 VGND a_81_23# X VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X16 a_1196_367# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X17 a_81_23# A3 a_910_345# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X18 a_81_23# C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X19 VGND A1 a_731_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X20 VPWR a_81_23# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X21 X a_81_23# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X22 a_731_47# A3 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X23 X a_81_23# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X24 a_910_345# A3 a_81_23# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X25 VGND a_81_23# X VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X26 X a_81_23# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X27 VPWR B1 a_81_23# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
.ends
