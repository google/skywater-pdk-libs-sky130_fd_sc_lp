# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_sc_lp__nor3b_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_lp__nor3b_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.720000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.995000 1.355000 2.685000 1.525000 ;
        RECT 1.115000 1.185000 1.955000 1.325000 ;
        RECT 1.115000 1.325000 2.685000 1.355000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.865000 1.210000 5.670000 1.335000 ;
        RECT 4.865000 1.335000 6.215000 1.505000 ;
    END
  END B
  PIN C_N
    ANTENNAGATEAREA  0.315000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.445000 1.185000 0.825000 1.515000 ;
    END
  END C_N
  PIN Y
    ANTENNADIFFAREA  2.116800 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.305000 0.255000 1.570000 0.845000 ;
        RECT 1.305000 0.845000 2.470000 0.985000 ;
        RECT 1.305000 0.985000 6.635000 1.015000 ;
        RECT 2.210000 1.015000 6.635000 1.040000 ;
        RECT 2.210000 1.040000 4.260000 1.155000 ;
        RECT 2.240000 0.255000 2.470000 0.845000 ;
        RECT 3.140000 0.255000 3.330000 0.985000 ;
        RECT 3.330000 1.675000 6.635000 1.855000 ;
        RECT 3.330000 1.855000 4.400000 2.145000 ;
        RECT 4.000000 0.255000 4.255000 0.870000 ;
        RECT 4.000000 0.870000 6.040000 0.985000 ;
        RECT 4.925000 0.255000 5.180000 0.870000 ;
        RECT 5.840000 1.040000 6.635000 1.155000 ;
        RECT 5.850000 0.255000 6.040000 0.870000 ;
        RECT 6.385000 1.155000 6.635000 1.675000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 6.720000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.000000 0.000000 6.720000 0.245000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.655000 6.910000 3.520000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 6.720000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.720000 0.085000 ;
      RECT 0.000000  3.245000 6.720000 3.415000 ;
      RECT 0.095000  0.255000 0.580000 1.015000 ;
      RECT 0.095000  1.015000 0.275000 1.705000 ;
      RECT 0.095000  1.705000 3.065000 1.875000 ;
      RECT 0.095000  1.875000 0.420000 3.075000 ;
      RECT 0.600000  2.105000 0.930000 3.245000 ;
      RECT 0.805000  0.085000 1.135000 1.015000 ;
      RECT 1.100000  2.045000 2.220000 2.225000 ;
      RECT 1.100000  2.225000 1.290000 3.065000 ;
      RECT 1.460000  2.395000 1.790000 3.245000 ;
      RECT 1.740000  0.085000 2.070000 0.675000 ;
      RECT 1.960000  2.225000 2.220000 2.325000 ;
      RECT 1.960000  2.325000 5.320000 2.495000 ;
      RECT 1.960000  2.495000 2.150000 3.065000 ;
      RECT 2.320000  2.665000 2.650000 3.245000 ;
      RECT 2.640000  0.085000 2.970000 0.815000 ;
      RECT 2.895000  1.325000 4.585000 1.505000 ;
      RECT 2.895000  1.505000 3.065000 1.705000 ;
      RECT 2.900000  2.665000 4.030000 2.875000 ;
      RECT 2.900000  2.875000 5.680000 2.885000 ;
      RECT 2.900000  2.885000 6.610000 3.075000 ;
      RECT 3.500000  0.085000 3.830000 0.815000 ;
      RECT 4.425000  0.085000 4.755000 0.700000 ;
      RECT 4.990000  2.025000 6.180000 2.205000 ;
      RECT 4.990000  2.205000 5.320000 2.325000 ;
      RECT 4.990000  2.495000 5.320000 2.705000 ;
      RECT 5.350000  0.085000 5.680000 0.700000 ;
      RECT 5.490000  2.375000 5.680000 2.875000 ;
      RECT 5.850000  2.205000 6.180000 2.705000 ;
      RECT 6.210000  0.085000 6.540000 0.815000 ;
      RECT 6.350000  2.025000 6.610000 2.885000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
  END
END sky130_fd_sc_lp__nor3b_4
END LIBRARY
