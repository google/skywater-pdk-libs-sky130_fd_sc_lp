* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__a2bb2o_lp A1_N A2_N B1 B2 VGND VNB VPB VPWR X
X0 X a_63_57# a_584_74# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 a_63_57# B2 a_150_57# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 a_314_57# a_284_31# a_63_57# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 a_43_408# B2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X4 a_150_57# B1 VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 VGND a_284_31# a_314_57# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 X a_63_57# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X7 a_900_74# A2_N VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 a_584_74# a_63_57# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 VPWR A1_N a_794_409# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X10 VGND A1_N a_742_74# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X11 VPWR B1 a_43_408# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X12 a_43_408# a_284_31# a_63_57# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X13 a_742_74# A1_N a_284_31# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X14 a_794_409# A2_N a_284_31# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X15 a_284_31# A2_N a_900_74# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
