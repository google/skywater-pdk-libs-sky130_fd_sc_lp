* File: sky130_fd_sc_lp__o21ai_m.pex.spice
* Created: Wed Sep  2 10:16:27 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O21AI_M%A1 2 5 9 11 12 13 14 19 20
r29 19 21 46.2775 $w=4.25e-07 $l=1.65e-07 $layer=POLY_cond $X=0.337 $Y=1.12
+ $X2=0.337 $Y2=0.955
r30 19 20 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.29
+ $Y=1.12 $X2=0.29 $Y2=1.12
r31 13 14 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.29 $Y=1.665
+ $X2=0.29 $Y2=2.035
r32 12 13 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.29 $Y=1.295
+ $X2=0.29 $Y2=1.665
r33 12 20 6.11144 $w=3.28e-07 $l=1.75e-07 $layer=LI1_cond $X=0.29 $Y=1.295
+ $X2=0.29 $Y2=1.12
r34 9 11 387.138 $w=1.5e-07 $l=7.55e-07 $layer=POLY_cond $X=0.475 $Y=2.38
+ $X2=0.475 $Y2=1.625
r35 5 21 251.255 $w=1.5e-07 $l=4.9e-07 $layer=POLY_cond $X=0.475 $Y=0.465
+ $X2=0.475 $Y2=0.955
r36 2 11 52.4279 $w=4.25e-07 $l=2.12e-07 $layer=POLY_cond $X=0.337 $Y=1.413
+ $X2=0.337 $Y2=1.625
r37 1 19 6.15041 $w=4.25e-07 $l=4.7e-08 $layer=POLY_cond $X=0.337 $Y=1.167
+ $X2=0.337 $Y2=1.12
r38 1 2 32.1915 $w=4.25e-07 $l=2.46e-07 $layer=POLY_cond $X=0.337 $Y=1.167
+ $X2=0.337 $Y2=1.413
.ends

.subckt PM_SKY130_FD_SC_LP__O21AI_M%A2 4 7 10 11 12 16
c35 4 0 1.09464e-19 $X=0.835 $Y=2.38
r36 16 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.925 $Y=2.915
+ $X2=0.925 $Y2=2.75
r37 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.925
+ $Y=2.915 $X2=0.925 $Y2=2.915
r38 12 17 10.2233 $w=3.08e-07 $l=2.75e-07 $layer=LI1_cond $X=1.2 $Y=2.845
+ $X2=0.925 $Y2=2.845
r39 11 17 7.62099 $w=3.08e-07 $l=2.05e-07 $layer=LI1_cond $X=0.72 $Y=2.845
+ $X2=0.925 $Y2=2.845
r40 9 10 43.7534 $w=2.2e-07 $l=1.5e-07 $layer=POLY_cond $X=0.87 $Y=1.91 $X2=0.87
+ $Y2=2.06
r41 7 9 740.947 $w=1.5e-07 $l=1.445e-06 $layer=POLY_cond $X=0.905 $Y=0.465
+ $X2=0.905 $Y2=1.91
r42 4 18 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=0.835 $Y=2.38
+ $X2=0.835 $Y2=2.75
r43 4 10 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.835 $Y=2.38
+ $X2=0.835 $Y2=2.06
.ends

.subckt PM_SKY130_FD_SC_LP__O21AI_M%B1 3 7 11 12 13 14 18 19
c35 18 0 3.66836e-20 $X=1.385 $Y=1.245
c36 3 0 9.67899e-20 $X=1.335 $Y=0.465
r37 18 19 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.385
+ $Y=1.245 $X2=1.385 $Y2=1.245
r38 13 14 12.0114 $w=3.53e-07 $l=3.7e-07 $layer=LI1_cond $X=1.292 $Y=1.295
+ $X2=1.292 $Y2=1.665
r39 13 19 1.62316 $w=3.53e-07 $l=5e-08 $layer=LI1_cond $X=1.292 $Y=1.295
+ $X2=1.292 $Y2=1.245
r40 11 18 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.385 $Y=1.585
+ $X2=1.385 $Y2=1.245
r41 11 12 38.0424 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.385 $Y=1.585
+ $X2=1.385 $Y2=1.75
r42 10 18 40.8701 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.385 $Y=1.08
+ $X2=1.385 $Y2=1.245
r43 7 12 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=1.375 $Y=2.38
+ $X2=1.375 $Y2=1.75
r44 3 10 315.351 $w=1.5e-07 $l=6.15e-07 $layer=POLY_cond $X=1.335 $Y=0.465
+ $X2=1.335 $Y2=1.08
.ends

.subckt PM_SKY130_FD_SC_LP__O21AI_M%VPWR 1 2 7 9 11 13 15 17 27
c25 13 0 1.09464e-19 $X=1.59 $Y=2.445
r26 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r27 23 24 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r28 21 27 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r29 20 21 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r30 18 23 4.78091 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=3.33
+ $X2=0.212 $Y2=3.33
r31 18 20 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=0.425 $Y=3.33
+ $X2=1.2 $Y2=3.33
r32 17 26 3.62463 $w=1.7e-07 $l=2.17e-07 $layer=LI1_cond $X=1.485 $Y=3.33
+ $X2=1.702 $Y2=3.33
r33 17 20 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.485 $Y=3.33
+ $X2=1.2 $Y2=3.33
r34 15 21 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=0.96 $Y=3.33
+ $X2=1.2 $Y2=3.33
r35 15 24 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=0.96 $Y=3.33
+ $X2=0.24 $Y2=3.33
r36 11 26 3.29056 $w=2.1e-07 $l=1.4854e-07 $layer=LI1_cond $X=1.59 $Y=3.245
+ $X2=1.702 $Y2=3.33
r37 11 13 42.2511 $w=2.08e-07 $l=8e-07 $layer=LI1_cond $X=1.59 $Y=3.245 $X2=1.59
+ $Y2=2.445
r38 7 23 2.98526 $w=3.3e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.26 $Y=3.245
+ $X2=0.212 $Y2=3.33
r39 7 9 27.938 $w=3.28e-07 $l=8e-07 $layer=LI1_cond $X=0.26 $Y=3.245 $X2=0.26
+ $Y2=2.445
r40 2 13 600 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=1 $X=1.45
+ $Y=2.17 $X2=1.59 $Y2=2.445
r41 1 9 600 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.17 $X2=0.26 $Y2=2.445
.ends

.subckt PM_SKY130_FD_SC_LP__O21AI_M%Y 1 2 8 12 14 15 16
r30 16 26 3.26203 $w=5.48e-07 $l=1.5e-07 $layer=LI1_cond $X=1.2 $Y=2.205
+ $X2=1.05 $Y2=2.205
r31 15 26 7.17647 $w=5.48e-07 $l=3.3e-07 $layer=LI1_cond $X=0.72 $Y=2.205
+ $X2=1.05 $Y2=2.205
r32 14 16 14.494 $w=3.18e-07 $l=3.65e-07 $layer=LI1_cond $X=1.65 $Y=2.015
+ $X2=1.285 $Y2=2.015
r33 10 12 8.71429 $w=2.08e-07 $l=1.65e-07 $layer=LI1_cond $X=1.57 $Y=0.53
+ $X2=1.735 $Y2=0.53
r34 8 14 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.735 $Y=1.93
+ $X2=1.65 $Y2=2.015
r35 7 12 1.9771 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.735 $Y=0.635
+ $X2=1.735 $Y2=0.53
r36 7 8 84.4866 $w=1.68e-07 $l=1.295e-06 $layer=LI1_cond $X=1.735 $Y=0.635
+ $X2=1.735 $Y2=1.93
r37 2 26 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.91
+ $Y=2.17 $X2=1.05 $Y2=2.315
r38 1 10 182 $w=1.7e-07 $l=3.45868e-07 $layer=licon1_NDIFF $count=1 $X=1.41
+ $Y=0.255 $X2=1.57 $Y2=0.53
.ends

.subckt PM_SKY130_FD_SC_LP__O21AI_M%A_27_51# 1 2 9 11 12 15
c23 15 0 2.54743e-19 $X=1.12 $Y=0.53
c24 11 0 3.66836e-20 $X=1.035 $Y=0.77
r25 13 15 9.04785 $w=1.88e-07 $l=1.55e-07 $layer=LI1_cond $X=1.13 $Y=0.685
+ $X2=1.13 $Y2=0.53
r26 11 13 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=1.035 $Y=0.77
+ $X2=1.13 $Y2=0.685
r27 11 12 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.035 $Y=0.77
+ $X2=0.345 $Y2=0.77
r28 7 12 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=0.25 $Y=0.685
+ $X2=0.345 $Y2=0.77
r29 7 9 9.04785 $w=1.88e-07 $l=1.55e-07 $layer=LI1_cond $X=0.25 $Y=0.685
+ $X2=0.25 $Y2=0.53
r30 2 15 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=0.98
+ $Y=0.255 $X2=1.12 $Y2=0.53
r31 1 9 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.255 $X2=0.26 $Y2=0.53
.ends

.subckt PM_SKY130_FD_SC_LP__O21AI_M%VGND 1 6 8 10 17 18 21
r24 21 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r25 17 18 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r26 15 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.855 $Y=0 $X2=0.69
+ $Y2=0
r27 15 17 53.8235 $w=1.68e-07 $l=8.25e-07 $layer=LI1_cond $X=0.855 $Y=0 $X2=1.68
+ $Y2=0
r28 13 22 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r29 12 13 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r30 10 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.525 $Y=0 $X2=0.69
+ $Y2=0
r31 10 12 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.525 $Y=0 $X2=0.24
+ $Y2=0
r32 8 18 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=0.96 $Y=0 $X2=1.68
+ $Y2=0
r33 8 22 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=0.96 $Y=0 $X2=0.72
+ $Y2=0
r34 4 21 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=0.085 $X2=0.69
+ $Y2=0
r35 4 6 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=0.69 $Y=0.085
+ $X2=0.69 $Y2=0.4
r36 1 6 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.255 $X2=0.69 $Y2=0.4
.ends

