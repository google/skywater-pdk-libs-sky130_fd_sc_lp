* File: sky130_fd_sc_lp__dlxtn_4.pex.spice
* Created: Wed Sep  2 09:48:37 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__DLXTN_4%D 3 7 8 9 13 15
r34 13 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.525 $Y=1.355
+ $X2=0.525 $Y2=1.52
r35 13 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.525 $Y=1.355
+ $X2=0.525 $Y2=1.19
r36 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.525
+ $Y=1.355 $X2=0.525 $Y2=1.355
r37 8 9 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=0.72 $Y=1.355 $X2=1.2
+ $Y2=1.355
r38 8 14 6.80989 $w=3.28e-07 $l=1.95e-07 $layer=LI1_cond $X=0.72 $Y=1.355
+ $X2=0.525 $Y2=1.355
r39 7 15 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.555 $Y=0.87
+ $X2=0.555 $Y2=1.19
r40 3 16 617.883 $w=1.5e-07 $l=1.205e-06 $layer=POLY_cond $X=0.495 $Y=2.725
+ $X2=0.495 $Y2=1.52
.ends

.subckt PM_SKY130_FD_SC_LP__DLXTN_4%GATE_N 3 5 7 9 10 13 16 18 19 20 24
c58 20 0 6.38949e-20 $X=1.68 $Y=0.555
r59 24 27 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.585 $Y=0.365
+ $X2=1.585 $Y2=0.53
r60 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.585
+ $Y=0.365 $X2=1.585 $Y2=0.365
r61 20 25 2.95898 $w=3.68e-07 $l=9.5e-08 $layer=LI1_cond $X=1.68 $Y=0.465
+ $X2=1.585 $Y2=0.465
r62 19 25 11.9916 $w=3.68e-07 $l=3.85e-07 $layer=LI1_cond $X=1.2 $Y=0.465
+ $X2=1.585 $Y2=0.465
r63 14 16 41.0213 $w=1.5e-07 $l=8e-08 $layer=POLY_cond $X=0.925 $Y=1.835
+ $X2=1.005 $Y2=1.835
r64 13 27 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.495 $Y=1.19
+ $X2=1.495 $Y2=0.53
r65 11 18 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.08 $Y=1.265
+ $X2=1.005 $Y2=1.265
r66 10 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.42 $Y=1.265
+ $X2=1.495 $Y2=1.19
r67 10 11 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=1.42 $Y=1.265
+ $X2=1.08 $Y2=1.265
r68 9 16 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.005 $Y=1.76
+ $X2=1.005 $Y2=1.835
r69 8 18 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.005 $Y=1.34
+ $X2=1.005 $Y2=1.265
r70 8 9 215.362 $w=1.5e-07 $l=4.2e-07 $layer=POLY_cond $X=1.005 $Y=1.34
+ $X2=1.005 $Y2=1.76
r71 5 18 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.005 $Y=1.19
+ $X2=1.005 $Y2=1.265
r72 5 7 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.005 $Y=1.19
+ $X2=1.005 $Y2=0.87
r73 1 14 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.925 $Y=1.91
+ $X2=0.925 $Y2=1.835
r74 1 3 417.904 $w=1.5e-07 $l=8.15e-07 $layer=POLY_cond $X=0.925 $Y=1.91
+ $X2=0.925 $Y2=2.725
.ends

.subckt PM_SKY130_FD_SC_LP__DLXTN_4%A_200_481# 1 2 9 11 13 16 20 25 28 31 33 37
+ 38 40 41 42 43 45 46 47 50 51 53 56 59
c168 47 0 8.67612e-20 $X=3.565 $Y=1.495
c169 11 0 6.38949e-20 $X=2.365 $Y=0.77
r170 59 66 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.245 $Y=1.06
+ $X2=3.245 $Y2=0.895
r171 58 59 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.245
+ $Y=1.06 $X2=3.245 $Y2=1.06
r172 55 56 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.975
+ $Y=1.06 $X2=1.975 $Y2=1.06
r173 53 55 0.157216 $w=3.88e-07 $l=5e-09 $layer=LI1_cond $X=1.917 $Y=1.055
+ $X2=1.917 $Y2=1.06
r174 51 70 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.6 $Y=2.045
+ $X2=3.6 $Y2=2.21
r175 50 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.6
+ $Y=2.045 $X2=3.6 $Y2=2.045
r176 48 50 15.7353 $w=2.58e-07 $l=3.55e-07 $layer=LI1_cond $X=3.565 $Y=2.4
+ $X2=3.565 $Y2=2.045
r177 47 50 24.3786 $w=2.58e-07 $l=5.5e-07 $layer=LI1_cond $X=3.565 $Y=1.495
+ $X2=3.565 $Y2=2.045
r178 46 47 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=3.245 $Y=1.41
+ $X2=3.565 $Y2=1.41
r179 45 58 2.68691 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=3.245 $Y=1.145
+ $X2=3.245 $Y2=1.055
r180 45 46 6.28605 $w=3.28e-07 $l=1.8e-07 $layer=LI1_cond $X=3.245 $Y=1.145
+ $X2=3.245 $Y2=1.325
r181 44 53 5.24902 $w=1.8e-07 $l=2.23e-07 $layer=LI1_cond $X=2.14 $Y=1.055
+ $X2=1.917 $Y2=1.055
r182 43 58 4.92601 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=3.08 $Y=1.055
+ $X2=3.245 $Y2=1.055
r183 43 44 57.9192 $w=1.78e-07 $l=9.4e-07 $layer=LI1_cond $X=3.08 $Y=1.055
+ $X2=2.14 $Y2=1.055
r184 41 48 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=3.435 $Y=2.485
+ $X2=3.565 $Y2=2.4
r185 41 42 85.139 $w=1.68e-07 $l=1.305e-06 $layer=LI1_cond $X=3.435 $Y=2.485
+ $X2=2.13 $Y2=2.485
r186 39 42 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.045 $Y=2.57
+ $X2=2.13 $Y2=2.485
r187 39 40 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=2.045 $Y=2.57
+ $X2=2.045 $Y2=2.905
r188 37 40 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.96 $Y=2.99
+ $X2=2.045 $Y2=2.905
r189 37 38 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=1.96 $Y=2.99
+ $X2=1.305 $Y2=2.99
r190 33 53 4.40206 $w=3.88e-07 $l=2.83485e-07 $layer=LI1_cond $X=1.695 $Y=0.915
+ $X2=1.917 $Y2=1.055
r191 33 35 27.7273 $w=1.88e-07 $l=4.75e-07 $layer=LI1_cond $X=1.695 $Y=0.915
+ $X2=1.22 $Y2=0.915
r192 29 38 7.51767 $w=1.7e-07 $l=1.8775e-07 $layer=LI1_cond $X=1.155 $Y=2.905
+ $X2=1.305 $Y2=2.99
r193 29 31 13.2531 $w=2.98e-07 $l=3.45e-07 $layer=LI1_cond $X=1.155 $Y=2.905
+ $X2=1.155 $Y2=2.56
r194 27 56 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.975 $Y=1.4
+ $X2=1.975 $Y2=1.06
r195 27 28 42.4377 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.975 $Y=1.4
+ $X2=1.975 $Y2=1.565
r196 23 56 24.4806 $w=3.3e-07 $l=1.4e-07 $layer=POLY_cond $X=1.975 $Y=0.92
+ $X2=1.975 $Y2=1.06
r197 23 25 199.979 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=1.975 $Y=0.845
+ $X2=2.365 $Y2=0.845
r198 20 70 217.926 $w=1.5e-07 $l=4.25e-07 $layer=POLY_cond $X=3.51 $Y=2.635
+ $X2=3.51 $Y2=2.21
r199 16 66 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=3.155 $Y=0.445
+ $X2=3.155 $Y2=0.895
r200 11 25 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.365 $Y=0.77
+ $X2=2.365 $Y2=0.845
r201 11 13 104.433 $w=1.5e-07 $l=3.25e-07 $layer=POLY_cond $X=2.365 $Y=0.77
+ $X2=2.365 $Y2=0.445
r202 9 28 605.064 $w=1.5e-07 $l=1.18e-06 $layer=POLY_cond $X=1.91 $Y=2.745
+ $X2=1.91 $Y2=1.565
r203 2 31 300 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_PDIFF $count=2 $X=1
+ $Y=2.405 $X2=1.14 $Y2=2.56
r204 1 35 182 $w=1.7e-07 $l=3.07124e-07 $layer=licon1_NDIFF $count=1 $X=1.08
+ $Y=0.66 $X2=1.22 $Y2=0.905
.ends

.subckt PM_SKY130_FD_SC_LP__DLXTN_4%A_27_481# 1 2 9 13 18 19 21 24 26 30 31 36
+ 38
r82 33 36 5.76222 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.175 $Y=0.845
+ $X2=0.34 $Y2=0.845
r83 30 31 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.52
+ $Y=1.445 $X2=2.52 $Y2=1.445
r84 28 30 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=2.52 $Y=1.7
+ $X2=2.52 $Y2=1.445
r85 27 38 2.47289 $w=1.8e-07 $l=1.6e-07 $layer=LI1_cond $X=0.41 $Y=1.79 $X2=0.25
+ $Y2=1.79
r86 26 28 7.61292 $w=1.8e-07 $l=2.05122e-07 $layer=LI1_cond $X=2.355 $Y=1.79
+ $X2=2.52 $Y2=1.7
r87 26 27 119.843 $w=1.78e-07 $l=1.945e-06 $layer=LI1_cond $X=2.355 $Y=1.79
+ $X2=0.41 $Y2=1.79
r88 22 38 3.96879 $w=2.45e-07 $l=9e-08 $layer=LI1_cond $X=0.25 $Y=1.88 $X2=0.25
+ $Y2=1.79
r89 22 24 24.1293 $w=3.18e-07 $l=6.7e-07 $layer=LI1_cond $X=0.25 $Y=1.88
+ $X2=0.25 $Y2=2.55
r90 21 38 3.96879 $w=2.45e-07 $l=1.21861e-07 $layer=LI1_cond $X=0.175 $Y=1.7
+ $X2=0.25 $Y2=1.79
r91 20 33 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.175 $Y=1.01
+ $X2=0.175 $Y2=0.845
r92 20 21 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=0.175 $Y=1.01
+ $X2=0.175 $Y2=1.7
r93 18 31 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.52 $Y=1.785
+ $X2=2.52 $Y2=1.445
r94 18 19 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.52 $Y=1.785
+ $X2=2.52 $Y2=1.95
r95 17 31 62.5236 $w=2.12e-07 $l=3.50999e-07 $layer=POLY_cond $X=2.795 $Y=1.272
+ $X2=2.52 $Y2=1.445
r96 11 17 10.9192 $w=1.5e-07 $l=1.72e-07 $layer=POLY_cond $X=2.795 $Y=1.1
+ $X2=2.795 $Y2=1.272
r97 11 13 335.862 $w=1.5e-07 $l=6.55e-07 $layer=POLY_cond $X=2.795 $Y=1.1
+ $X2=2.795 $Y2=0.445
r98 9 19 407.649 $w=1.5e-07 $l=7.95e-07 $layer=POLY_cond $X=2.61 $Y=2.745
+ $X2=2.61 $Y2=1.95
r99 2 24 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.405 $X2=0.26 $Y2=2.55
r100 1 36 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=0.215
+ $Y=0.66 $X2=0.34 $Y2=0.845
.ends

.subckt PM_SKY130_FD_SC_LP__DLXTN_4%A_310_485# 1 2 9 11 12 15 18 21 24 25 28 30
+ 31 34 36 37 40 41 43 47
r124 46 47 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.785
+ $Y=0.98 $X2=3.785 $Y2=0.98
r125 43 46 9.42908 $w=3.28e-07 $l=2.7e-07 $layer=LI1_cond $X=3.785 $Y=0.71
+ $X2=3.785 $Y2=0.98
r126 40 41 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.06
+ $Y=1.76 $X2=3.06 $Y2=1.76
r127 38 40 10.1275 $w=3.28e-07 $l=2.9e-07 $layer=LI1_cond $X=3.06 $Y=2.05
+ $X2=3.06 $Y2=1.76
r128 36 43 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.62 $Y=0.71
+ $X2=3.785 $Y2=0.71
r129 36 37 90.3583 $w=1.68e-07 $l=1.385e-06 $layer=LI1_cond $X=3.62 $Y=0.71
+ $X2=2.235 $Y2=0.71
r130 32 37 6.87494 $w=1.7e-07 $l=1.36015e-07 $layer=LI1_cond $X=2.135 $Y=0.625
+ $X2=2.235 $Y2=0.71
r131 32 34 10.5364 $w=1.98e-07 $l=1.9e-07 $layer=LI1_cond $X=2.135 $Y=0.625
+ $X2=2.135 $Y2=0.435
r132 30 38 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.895 $Y=2.135
+ $X2=3.06 $Y2=2.05
r133 30 31 72.7433 $w=1.68e-07 $l=1.115e-06 $layer=LI1_cond $X=2.895 $Y=2.135
+ $X2=1.78 $Y2=2.135
r134 26 31 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.655 $Y=2.22
+ $X2=1.78 $Y2=2.135
r135 26 28 16.1342 $w=2.48e-07 $l=3.5e-07 $layer=LI1_cond $X=1.655 $Y=2.22
+ $X2=1.655 $Y2=2.57
r136 24 47 34.0979 $w=3.3e-07 $l=1.95e-07 $layer=POLY_cond $X=3.785 $Y=1.175
+ $X2=3.785 $Y2=0.98
r137 24 25 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.785 $Y=1.175
+ $X2=3.785 $Y2=1.34
r138 23 47 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.785 $Y=0.815
+ $X2=3.785 $Y2=0.98
r139 20 41 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=3.06 $Y=2.1
+ $X2=3.06 $Y2=1.76
r140 20 21 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.06 $Y=2.1
+ $X2=3.06 $Y2=2.265
r141 19 41 20.9834 $w=3.3e-07 $l=1.2e-07 $layer=POLY_cond $X=3.06 $Y=1.64
+ $X2=3.06 $Y2=1.76
r142 18 25 76.9149 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=3.695 $Y=1.49
+ $X2=3.695 $Y2=1.34
r143 15 23 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=3.695 $Y=0.445
+ $X2=3.695 $Y2=0.815
r144 12 19 114.514 $w=6.7e-08 $l=1.98997e-07 $layer=POLY_cond $X=3.225 $Y=1.565
+ $X2=3.06 $Y2=1.64
r145 11 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.62 $Y=1.565
+ $X2=3.695 $Y2=1.49
r146 11 12 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=3.62 $Y=1.565
+ $X2=3.225 $Y2=1.565
r147 9 21 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.97 $Y=2.745
+ $X2=2.97 $Y2=2.265
r148 2 28 600 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=1.55
+ $Y=2.425 $X2=1.695 $Y2=2.57
r149 1 34 182 $w=1.7e-07 $l=2.54951e-07 $layer=licon1_NDIFF $count=1 $X=2.025
+ $Y=0.235 $X2=2.15 $Y2=0.435
.ends

.subckt PM_SKY130_FD_SC_LP__DLXTN_4%A_795_423# 1 2 9 13 15 19 23 27 31 35 39 43
+ 47 51 53 55 57 58 60 64 68 73 75 81 86 87 88 89 92 102
c164 15 0 2.36442e-20 $X=4.25 $Y=1.43
c165 13 0 6.3117e-20 $X=4.235 $Y=0.445
r166 102 103 4.43558 $w=3.26e-07 $l=3e-08 $layer=POLY_cond $X=7.175 $Y=1.43
+ $X2=7.205 $Y2=1.43
r167 101 102 59.1411 $w=3.26e-07 $l=4e-07 $layer=POLY_cond $X=6.775 $Y=1.43
+ $X2=7.175 $Y2=1.43
r168 100 101 4.43558 $w=3.26e-07 $l=3e-08 $layer=POLY_cond $X=6.745 $Y=1.43
+ $X2=6.775 $Y2=1.43
r169 97 98 4.43558 $w=3.26e-07 $l=3e-08 $layer=POLY_cond $X=6.315 $Y=1.43
+ $X2=6.345 $Y2=1.43
r170 96 97 59.1411 $w=3.26e-07 $l=4e-07 $layer=POLY_cond $X=5.915 $Y=1.43
+ $X2=6.315 $Y2=1.43
r171 95 96 4.43558 $w=3.26e-07 $l=3e-08 $layer=POLY_cond $X=5.885 $Y=1.43
+ $X2=5.915 $Y2=1.43
r172 92 95 10.9545 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=5.81 $Y=1.43
+ $X2=5.885 $Y2=1.43
r173 85 86 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.3
+ $Y=1.76 $X2=4.3 $Y2=1.76
r174 82 100 31.7883 $w=3.26e-07 $l=2.15e-07 $layer=POLY_cond $X=6.53 $Y=1.43
+ $X2=6.745 $Y2=1.43
r175 82 98 27.3528 $w=3.26e-07 $l=1.85e-07 $layer=POLY_cond $X=6.53 $Y=1.43
+ $X2=6.345 $Y2=1.43
r176 81 82 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.53
+ $Y=1.43 $X2=6.53 $Y2=1.43
r177 79 92 52.4584 $w=3.3e-07 $l=3e-07 $layer=POLY_cond $X=5.51 $Y=1.43 $X2=5.81
+ $Y2=1.43
r178 78 81 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=5.51 $Y=1.43
+ $X2=6.53 $Y2=1.43
r179 78 79 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.51
+ $Y=1.43 $X2=5.51 $Y2=1.43
r180 76 89 1.44715 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=5.385 $Y=1.43
+ $X2=5.295 $Y2=1.43
r181 76 78 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=5.385 $Y=1.43
+ $X2=5.51 $Y2=1.43
r182 75 88 3.98977 $w=2.3e-07 $l=1.11018e-07 $layer=LI1_cond $X=5.29 $Y=1.675
+ $X2=5.23 $Y2=1.76
r183 74 89 5.04255 $w=1.75e-07 $l=8.74643e-08 $layer=LI1_cond $X=5.29 $Y=1.515
+ $X2=5.295 $Y2=1.43
r184 74 75 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=5.29 $Y=1.515
+ $X2=5.29 $Y2=1.675
r185 73 89 5.04255 $w=1.75e-07 $l=8.5e-08 $layer=LI1_cond $X=5.295 $Y=1.345
+ $X2=5.295 $Y2=1.43
r186 73 87 16.6364 $w=1.78e-07 $l=2.7e-07 $layer=LI1_cond $X=5.295 $Y=1.345
+ $X2=5.295 $Y2=1.075
r187 68 70 38.5472 $w=2.88e-07 $l=9.7e-07 $layer=LI1_cond $X=5.23 $Y=1.9
+ $X2=5.23 $Y2=2.87
r188 66 88 3.98977 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.23 $Y=1.845
+ $X2=5.23 $Y2=1.76
r189 66 68 2.18567 $w=2.88e-07 $l=5.5e-08 $layer=LI1_cond $X=5.23 $Y=1.845
+ $X2=5.23 $Y2=1.9
r190 62 87 11.0699 $w=4.93e-07 $l=2.47e-07 $layer=LI1_cond $X=5.137 $Y=0.828
+ $X2=5.137 $Y2=1.075
r191 62 64 9.85859 $w=4.93e-07 $l=4.08e-07 $layer=LI1_cond $X=5.137 $Y=0.828
+ $X2=5.137 $Y2=0.42
r192 61 85 3.71371 $w=1.7e-07 $l=1.2339e-07 $layer=LI1_cond $X=4.415 $Y=1.76
+ $X2=4.31 $Y2=1.72
r193 60 88 2.45049 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=5.085 $Y=1.76
+ $X2=5.23 $Y2=1.76
r194 60 61 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.085 $Y=1.76
+ $X2=4.415 $Y2=1.76
r195 58 86 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=4.3 $Y=2.1 $X2=4.3
+ $Y2=1.76
r196 57 58 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.3
+ $Y=2.1 $X2=4.3 $Y2=2.1
r197 55 85 3.20148 $w=2.1e-07 $l=1.25e-07 $layer=LI1_cond $X=4.31 $Y=1.845
+ $X2=4.31 $Y2=1.72
r198 55 57 13.4675 $w=2.08e-07 $l=2.55e-07 $layer=LI1_cond $X=4.31 $Y=1.845
+ $X2=4.31 $Y2=2.1
r199 53 86 37.7308 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.3 $Y=1.595
+ $X2=4.3 $Y2=1.76
r200 50 58 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=4.3 $Y=2.115
+ $X2=4.3 $Y2=2.1
r201 50 51 43.5886 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=4.22 $Y=2.115
+ $X2=4.22 $Y2=2.265
r202 45 103 20.933 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.205 $Y=1.595
+ $X2=7.205 $Y2=1.43
r203 45 47 446.106 $w=1.5e-07 $l=8.7e-07 $layer=POLY_cond $X=7.205 $Y=1.595
+ $X2=7.205 $Y2=2.465
r204 41 102 20.933 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.175 $Y=1.265
+ $X2=7.175 $Y2=1.43
r205 41 43 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=7.175 $Y=1.265
+ $X2=7.175 $Y2=0.655
r206 37 101 20.933 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.775 $Y=1.595
+ $X2=6.775 $Y2=1.43
r207 37 39 446.106 $w=1.5e-07 $l=8.7e-07 $layer=POLY_cond $X=6.775 $Y=1.595
+ $X2=6.775 $Y2=2.465
r208 33 100 20.933 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.745 $Y=1.265
+ $X2=6.745 $Y2=1.43
r209 33 35 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=6.745 $Y=1.265
+ $X2=6.745 $Y2=0.655
r210 29 98 20.933 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.345 $Y=1.595
+ $X2=6.345 $Y2=1.43
r211 29 31 446.106 $w=1.5e-07 $l=8.7e-07 $layer=POLY_cond $X=6.345 $Y=1.595
+ $X2=6.345 $Y2=2.465
r212 25 97 20.933 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.315 $Y=1.265
+ $X2=6.315 $Y2=1.43
r213 25 27 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=6.315 $Y=1.265
+ $X2=6.315 $Y2=0.655
r214 21 96 20.933 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.915 $Y=1.595
+ $X2=5.915 $Y2=1.43
r215 21 23 446.106 $w=1.5e-07 $l=8.7e-07 $layer=POLY_cond $X=5.915 $Y=1.595
+ $X2=5.915 $Y2=2.465
r216 17 95 20.933 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.885 $Y=1.265
+ $X2=5.885 $Y2=1.43
r217 17 19 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=5.885 $Y=1.265
+ $X2=5.885 $Y2=0.655
r218 15 54 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=4.25 $Y=1.43 $X2=4.25
+ $Y2=1.34
r219 15 53 64.1371 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=4.25 $Y=1.43
+ $X2=4.25 $Y2=1.595
r220 13 54 458.926 $w=1.5e-07 $l=8.95e-07 $layer=POLY_cond $X=4.235 $Y=0.445
+ $X2=4.235 $Y2=1.34
r221 9 51 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=4.05 $Y=2.635
+ $X2=4.05 $Y2=2.265
r222 2 70 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=5.04
+ $Y=1.755 $X2=5.18 $Y2=2.87
r223 2 68 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=5.04
+ $Y=1.755 $X2=5.18 $Y2=1.9
r224 1 64 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=4.855
+ $Y=0.235 $X2=4.995 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__DLXTN_4%A_609_485# 1 2 7 9 12 14 18 23 25 27 32 34
+ 39
r100 33 39 16.6118 $w=3.3e-07 $l=9.5e-08 $layer=POLY_cond $X=4.87 $Y=1.35
+ $X2=4.965 $Y2=1.35
r101 33 36 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=4.87 $Y=1.35 $X2=4.78
+ $Y2=1.35
r102 32 34 8.69362 $w=2.58e-07 $l=1.65e-07 $layer=LI1_cond $X=4.87 $Y=1.375
+ $X2=4.705 $Y2=1.375
r103 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.87
+ $Y=1.35 $X2=4.87 $Y2=1.35
r104 28 30 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=3.95 $Y=1.33
+ $X2=4.215 $Y2=1.33
r105 27 30 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=4.3 $Y=1.33
+ $X2=4.215 $Y2=1.33
r106 27 34 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=4.3 $Y=1.33
+ $X2=4.705 $Y2=1.33
r107 25 30 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.215 $Y=1.245
+ $X2=4.215 $Y2=1.33
r108 24 25 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=4.215 $Y=0.455
+ $X2=4.215 $Y2=1.245
r109 22 28 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.95 $Y=1.415
+ $X2=3.95 $Y2=1.33
r110 22 23 86.4438 $w=1.68e-07 $l=1.325e-06 $layer=LI1_cond $X=3.95 $Y=1.415
+ $X2=3.95 $Y2=2.74
r111 18 24 6.87494 $w=2e-07 $l=1.36015e-07 $layer=LI1_cond $X=4.13 $Y=0.355
+ $X2=4.215 $Y2=0.455
r112 18 20 39.65 $w=1.98e-07 $l=7.15e-07 $layer=LI1_cond $X=4.13 $Y=0.355
+ $X2=3.415 $Y2=0.355
r113 14 23 7.36005 $w=2.8e-07 $l=1.77482e-07 $layer=LI1_cond $X=3.865 $Y=2.88
+ $X2=3.95 $Y2=2.74
r114 14 16 27.9879 $w=2.78e-07 $l=6.8e-07 $layer=LI1_cond $X=3.865 $Y=2.88
+ $X2=3.185 $Y2=2.88
r115 10 39 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.965 $Y=1.515
+ $X2=4.965 $Y2=1.35
r116 10 12 446.106 $w=1.5e-07 $l=8.7e-07 $layer=POLY_cond $X=4.965 $Y=1.515
+ $X2=4.965 $Y2=2.385
r117 7 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.78 $Y=1.185
+ $X2=4.78 $Y2=1.35
r118 7 9 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=4.78 $Y=1.185
+ $X2=4.78 $Y2=0.655
r119 2 16 600 $w=1.7e-07 $l=4.95076e-07 $layer=licon1_PDIFF $count=1 $X=3.045
+ $Y=2.425 $X2=3.185 $Y2=2.855
r120 1 20 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=3.23
+ $Y=0.235 $X2=3.415 $Y2=0.36
.ends

.subckt PM_SKY130_FD_SC_LP__DLXTN_4%VPWR 1 2 3 4 5 6 21 25 28 31 35 41 45 47 52
+ 53 55 58 59 60 62 74 85 89 95 98 101 105
r110 104 105 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r111 101 102 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r112 98 99 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r113 95 96 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r114 93 105 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=7.44 $Y2=3.33
r115 93 102 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=6.48 $Y2=3.33
r116 92 93 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r117 90 101 7.94884 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=6.69 $Y=3.33
+ $X2=6.542 $Y2=3.33
r118 90 92 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=6.69 $Y=3.33
+ $X2=6.96 $Y2=3.33
r119 89 104 4.69085 $w=1.7e-07 $l=2.07e-07 $layer=LI1_cond $X=7.265 $Y=3.33
+ $X2=7.472 $Y2=3.33
r120 89 92 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=7.265 $Y=3.33
+ $X2=6.96 $Y2=3.33
r121 88 102 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33
+ $X2=6.48 $Y2=3.33
r122 87 88 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r123 85 101 7.94884 $w=1.7e-07 $l=1.47e-07 $layer=LI1_cond $X=6.395 $Y=3.33
+ $X2=6.542 $Y2=3.33
r124 85 87 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=6.395 $Y=3.33
+ $X2=6 $Y2=3.33
r125 84 88 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33 $X2=6
+ $Y2=3.33
r126 84 99 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=4.56 $Y2=3.33
r127 83 84 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r128 81 98 13.764 $w=1.7e-07 $l=3.55e-07 $layer=LI1_cond $X=4.915 $Y=3.33
+ $X2=4.56 $Y2=3.33
r129 81 83 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=4.915 $Y=3.33
+ $X2=5.52 $Y2=3.33
r130 80 99 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r131 79 80 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r132 76 79 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=2.64 $Y=3.33
+ $X2=4.08 $Y2=3.33
r133 76 77 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r134 74 98 13.764 $w=1.7e-07 $l=3.55e-07 $layer=LI1_cond $X=4.205 $Y=3.33
+ $X2=4.56 $Y2=3.33
r135 74 79 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=4.205 $Y=3.33
+ $X2=4.08 $Y2=3.33
r136 73 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r137 72 73 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r138 70 73 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r139 70 96 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r140 69 72 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=3.33 $X2=2.16
+ $Y2=3.33
r141 69 70 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r142 67 95 7.13466 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=0.835 $Y=3.33
+ $X2=0.707 $Y2=3.33
r143 67 69 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.835 $Y=3.33
+ $X2=1.2 $Y2=3.33
r144 65 96 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r145 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r146 62 95 7.13466 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=0.58 $Y=3.33
+ $X2=0.707 $Y2=3.33
r147 62 64 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=0.58 $Y=3.33
+ $X2=0.24 $Y2=3.33
r148 60 80 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.84 $Y=3.33
+ $X2=4.08 $Y2=3.33
r149 60 77 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=3.84 $Y=3.33
+ $X2=2.64 $Y2=3.33
r150 58 83 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=5.545 $Y=3.33
+ $X2=5.52 $Y2=3.33
r151 58 59 7.75133 $w=1.7e-07 $l=1.42e-07 $layer=LI1_cond $X=5.545 $Y=3.33
+ $X2=5.687 $Y2=3.33
r152 57 87 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=5.83 $Y=3.33 $X2=6
+ $Y2=3.33
r153 57 59 7.75133 $w=1.7e-07 $l=1.43e-07 $layer=LI1_cond $X=5.83 $Y=3.33
+ $X2=5.687 $Y2=3.33
r154 55 56 6.82277 $w=7.08e-07 $l=2e-07 $layer=LI1_cond $X=4.56 $Y=2.635
+ $X2=4.56 $Y2=2.435
r155 52 72 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=2.3 $Y=3.33
+ $X2=2.16 $Y2=3.33
r156 52 53 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.3 $Y=3.33 $X2=2.43
+ $Y2=3.33
r157 51 76 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=2.56 $Y=3.33 $X2=2.64
+ $Y2=3.33
r158 51 53 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.56 $Y=3.33
+ $X2=2.43 $Y2=3.33
r159 47 50 34.9334 $w=3.18e-07 $l=9.7e-07 $layer=LI1_cond $X=7.425 $Y=1.98
+ $X2=7.425 $Y2=2.95
r160 45 104 2.99127 $w=3.2e-07 $l=1.05924e-07 $layer=LI1_cond $X=7.425 $Y=3.245
+ $X2=7.472 $Y2=3.33
r161 45 50 10.6241 $w=3.18e-07 $l=2.95e-07 $layer=LI1_cond $X=7.425 $Y=3.245
+ $X2=7.425 $Y2=2.95
r162 41 44 29.6901 $w=2.93e-07 $l=7.6e-07 $layer=LI1_cond $X=6.542 $Y=2.19
+ $X2=6.542 $Y2=2.95
r163 39 101 0.543863 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=6.542 $Y=3.245
+ $X2=6.542 $Y2=3.33
r164 39 44 11.5244 $w=2.93e-07 $l=2.95e-07 $layer=LI1_cond $X=6.542 $Y=3.245
+ $X2=6.542 $Y2=2.95
r165 35 38 39.2235 $w=2.83e-07 $l=9.7e-07 $layer=LI1_cond $X=5.687 $Y=1.98
+ $X2=5.687 $Y2=2.95
r166 33 59 0.432977 $w=2.85e-07 $l=8.5e-08 $layer=LI1_cond $X=5.687 $Y=3.245
+ $X2=5.687 $Y2=3.33
r167 33 38 11.9288 $w=2.83e-07 $l=2.95e-07 $layer=LI1_cond $X=5.687 $Y=3.245
+ $X2=5.687 $Y2=2.95
r168 31 56 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=4.75 $Y=2.1
+ $X2=4.75 $Y2=2.435
r169 28 98 2.89202 $w=7.1e-07 $l=8.5e-08 $layer=LI1_cond $X=4.56 $Y=3.245
+ $X2=4.56 $Y2=3.33
r170 27 55 2.61116 $w=7.08e-07 $l=1.55e-07 $layer=LI1_cond $X=4.56 $Y=2.79
+ $X2=4.56 $Y2=2.635
r171 27 28 7.66501 $w=7.08e-07 $l=4.55e-07 $layer=LI1_cond $X=4.56 $Y=2.79
+ $X2=4.56 $Y2=3.245
r172 23 53 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=2.43 $Y=3.245
+ $X2=2.43 $Y2=3.33
r173 23 25 15.0704 $w=2.58e-07 $l=3.4e-07 $layer=LI1_cond $X=2.43 $Y=3.245
+ $X2=2.43 $Y2=2.905
r174 19 95 0.067832 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=0.707 $Y=3.245
+ $X2=0.707 $Y2=3.33
r175 19 21 30.9578 $w=2.53e-07 $l=6.85e-07 $layer=LI1_cond $X=0.707 $Y=3.245
+ $X2=0.707 $Y2=2.56
r176 6 50 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=7.28
+ $Y=1.835 $X2=7.42 $Y2=2.95
r177 6 47 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=7.28
+ $Y=1.835 $X2=7.42 $Y2=1.98
r178 5 44 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=6.42
+ $Y=1.835 $X2=6.56 $Y2=2.95
r179 5 41 400 $w=1.7e-07 $l=4.19196e-07 $layer=licon1_PDIFF $count=1 $X=6.42
+ $Y=1.835 $X2=6.56 $Y2=2.19
r180 4 38 400 $w=1.7e-07 $l=1.17584e-06 $layer=licon1_PDIFF $count=1 $X=5.575
+ $Y=1.835 $X2=5.7 $Y2=2.95
r181 4 35 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=5.575
+ $Y=1.835 $X2=5.7 $Y2=1.98
r182 3 55 300 $w=1.7e-07 $l=2.80624e-07 $layer=licon1_PDIFF $count=2 $X=4.125
+ $Y=2.425 $X2=4.29 $Y2=2.635
r183 3 31 300 $w=1.7e-07 $l=7.70552e-07 $layer=licon1_PDIFF $count=2 $X=4.125
+ $Y=2.425 $X2=4.75 $Y2=2.1
r184 2 25 600 $w=1.7e-07 $l=6.53605e-07 $layer=licon1_PDIFF $count=1 $X=1.985
+ $Y=2.425 $X2=2.395 $Y2=2.905
r185 1 21 300 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_PDIFF $count=2 $X=0.57
+ $Y=2.405 $X2=0.71 $Y2=2.56
.ends

.subckt PM_SKY130_FD_SC_LP__DLXTN_4%Q 1 2 3 4 15 19 23 24 25 26 27 28 29 30 39
+ 43 50
r52 45 50 1.00212 $w=2.28e-07 $l=2e-08 $layer=LI1_cond $X=6.98 $Y=1.685 $X2=6.98
+ $Y2=1.665
r53 37 43 4.1907 $w=2.18e-07 $l=8e-08 $layer=LI1_cond $X=6.985 $Y=1.005
+ $X2=6.985 $Y2=0.925
r54 30 56 45.6073 $w=2.33e-07 $l=9.3e-07 $layer=LI1_cond $X=6.977 $Y=1.98
+ $X2=6.977 $Y2=2.91
r55 30 51 6.13002 $w=2.33e-07 $l=1.25e-07 $layer=LI1_cond $X=6.977 $Y=1.98
+ $X2=6.977 $Y2=1.855
r56 29 45 3.95216 $w=2.32e-07 $l=8.6487e-08 $layer=LI1_cond $X=6.977 $Y=1.77
+ $X2=6.98 $Y2=1.685
r57 29 51 3.95216 $w=2.32e-07 $l=8.5e-08 $layer=LI1_cond $X=6.977 $Y=1.77
+ $X2=6.977 $Y2=1.855
r58 29 50 1.65351 $w=2.28e-07 $l=3.3e-08 $layer=LI1_cond $X=6.98 $Y=1.632
+ $X2=6.98 $Y2=1.665
r59 28 29 16.8858 $w=2.28e-07 $l=3.37e-07 $layer=LI1_cond $X=6.98 $Y=1.295
+ $X2=6.98 $Y2=1.632
r60 28 44 6.01275 $w=2.28e-07 $l=1.2e-07 $layer=LI1_cond $X=6.98 $Y=1.295
+ $X2=6.98 $Y2=1.175
r61 27 37 4.06715 $w=2.25e-07 $l=8.74643e-08 $layer=LI1_cond $X=6.98 $Y=1.09
+ $X2=6.985 $Y2=1.005
r62 27 44 4.06715 $w=2.25e-07 $l=8.5e-08 $layer=LI1_cond $X=6.98 $Y=1.09
+ $X2=6.98 $Y2=1.175
r63 27 43 0.157151 $w=2.18e-07 $l=3e-09 $layer=LI1_cond $X=6.985 $Y=0.922
+ $X2=6.985 $Y2=0.925
r64 27 39 26.2967 $w=2.18e-07 $l=5.02e-07 $layer=LI1_cond $X=6.985 $Y=0.922
+ $X2=6.985 $Y2=0.42
r65 25 29 2.49072 $w=1.7e-07 $l=1.17e-07 $layer=LI1_cond $X=6.86 $Y=1.77
+ $X2=6.977 $Y2=1.77
r66 25 26 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=6.86 $Y=1.77
+ $X2=6.225 $Y2=1.77
r67 23 27 2.36881 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=6.865 $Y=1.09
+ $X2=6.98 $Y2=1.09
r68 23 24 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=6.865 $Y=1.09
+ $X2=6.195 $Y2=1.09
r69 19 21 47.6343 $w=2.23e-07 $l=9.3e-07 $layer=LI1_cond $X=6.112 $Y=1.98
+ $X2=6.112 $Y2=2.91
r70 17 26 6.9898 $w=1.7e-07 $l=1.49579e-07 $layer=LI1_cond $X=6.112 $Y=1.855
+ $X2=6.225 $Y2=1.77
r71 17 19 6.40246 $w=2.23e-07 $l=1.25e-07 $layer=LI1_cond $X=6.112 $Y=1.855
+ $X2=6.112 $Y2=1.98
r72 13 24 6.9898 $w=1.7e-07 $l=1.49579e-07 $layer=LI1_cond $X=6.082 $Y=1.005
+ $X2=6.195 $Y2=1.09
r73 13 15 29.9635 $w=2.23e-07 $l=5.85e-07 $layer=LI1_cond $X=6.082 $Y=1.005
+ $X2=6.082 $Y2=0.42
r74 4 56 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=6.85
+ $Y=1.835 $X2=6.99 $Y2=2.91
r75 4 30 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=6.85
+ $Y=1.835 $X2=6.99 $Y2=1.98
r76 3 21 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=5.99
+ $Y=1.835 $X2=6.13 $Y2=2.91
r77 3 19 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=5.99
+ $Y=1.835 $X2=6.13 $Y2=1.98
r78 2 39 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=6.82
+ $Y=0.235 $X2=6.96 $Y2=0.42
r79 1 15 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=5.96
+ $Y=0.235 $X2=6.1 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__DLXTN_4%VGND 1 2 3 4 5 6 23 27 31 35 39 41 43 46 47
+ 48 50 58 70 74 80 83 86 89 93
r102 92 93 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r103 89 90 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r104 86 87 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r105 83 84 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r106 80 81 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r107 78 93 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=7.44
+ $Y2=0
r108 78 90 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=6.48
+ $Y2=0
r109 77 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r110 75 89 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.695 $Y=0 $X2=6.53
+ $Y2=0
r111 75 77 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=6.695 $Y=0
+ $X2=6.96 $Y2=0
r112 74 92 3.78308 $w=1.7e-07 $l=2.07e-07 $layer=LI1_cond $X=7.265 $Y=0
+ $X2=7.472 $Y2=0
r113 74 77 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=7.265 $Y=0
+ $X2=6.96 $Y2=0
r114 73 90 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.48
+ $Y2=0
r115 72 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6 $Y2=0
r116 70 89 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.365 $Y=0 $X2=6.53
+ $Y2=0
r117 70 72 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=6.365 $Y=0 $X2=6
+ $Y2=0
r118 69 73 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=6
+ $Y2=0
r119 69 87 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=4.56
+ $Y2=0
r120 68 69 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r121 66 86 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.72 $Y=0 $X2=4.595
+ $Y2=0
r122 66 68 52.1925 $w=1.68e-07 $l=8e-07 $layer=LI1_cond $X=4.72 $Y=0 $X2=5.52
+ $Y2=0
r123 65 87 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=4.56
+ $Y2=0
r124 64 65 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r125 62 84 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.64
+ $Y2=0
r126 61 64 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=3.12 $Y=0 $X2=4.08
+ $Y2=0
r127 61 62 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r128 59 83 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.745 $Y=0 $X2=2.58
+ $Y2=0
r129 59 61 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=2.745 $Y=0
+ $X2=3.12 $Y2=0
r130 58 86 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.47 $Y=0 $X2=4.595
+ $Y2=0
r131 58 64 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=4.47 $Y=0 $X2=4.08
+ $Y2=0
r132 57 84 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r133 56 57 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r134 54 57 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r135 54 81 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r136 53 56 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r137 53 54 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r138 51 80 6.92067 $w=1.7e-07 $l=1.23e-07 $layer=LI1_cond $X=0.885 $Y=0
+ $X2=0.762 $Y2=0
r139 51 53 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.885 $Y=0 $X2=1.2
+ $Y2=0
r140 50 83 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.415 $Y=0 $X2=2.58
+ $Y2=0
r141 50 56 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=2.415 $Y=0
+ $X2=2.16 $Y2=0
r142 48 65 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.84 $Y=0
+ $X2=4.08 $Y2=0
r143 48 62 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=3.84 $Y=0 $X2=3.12
+ $Y2=0
r144 46 68 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=5.555 $Y=0 $X2=5.52
+ $Y2=0
r145 46 47 6.92067 $w=1.7e-07 $l=1.22e-07 $layer=LI1_cond $X=5.555 $Y=0
+ $X2=5.677 $Y2=0
r146 45 72 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=5.8 $Y=0 $X2=6 $Y2=0
r147 45 47 6.92067 $w=1.7e-07 $l=1.23e-07 $layer=LI1_cond $X=5.8 $Y=0 $X2=5.677
+ $Y2=0
r148 41 92 3.23481 $w=2.3e-07 $l=1.27609e-07 $layer=LI1_cond $X=7.38 $Y=0.085
+ $X2=7.472 $Y2=0
r149 41 43 14.7813 $w=2.28e-07 $l=2.95e-07 $layer=LI1_cond $X=7.38 $Y=0.085
+ $X2=7.38 $Y2=0.38
r150 37 89 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.53 $Y=0.085
+ $X2=6.53 $Y2=0
r151 37 39 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=6.53 $Y=0.085
+ $X2=6.53 $Y2=0.38
r152 33 47 0.066131 $w=2.45e-07 $l=8.5e-08 $layer=LI1_cond $X=5.677 $Y=0.085
+ $X2=5.677 $Y2=0
r153 33 35 13.8764 $w=2.43e-07 $l=2.95e-07 $layer=LI1_cond $X=5.677 $Y=0.085
+ $X2=5.677 $Y2=0.38
r154 29 86 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.595 $Y=0.085
+ $X2=4.595 $Y2=0
r155 29 31 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=4.595 $Y=0.085
+ $X2=4.595 $Y2=0.38
r156 25 83 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.58 $Y=0.085
+ $X2=2.58 $Y2=0
r157 25 27 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.58 $Y=0.085
+ $X2=2.58 $Y2=0.36
r158 21 80 0.066131 $w=2.45e-07 $l=8.5e-08 $layer=LI1_cond $X=0.762 $Y=0.085
+ $X2=0.762 $Y2=0
r159 21 23 36.2196 $w=2.43e-07 $l=7.7e-07 $layer=LI1_cond $X=0.762 $Y=0.085
+ $X2=0.762 $Y2=0.855
r160 6 43 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=7.25
+ $Y=0.235 $X2=7.39 $Y2=0.38
r161 5 39 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.39
+ $Y=0.235 $X2=6.53 $Y2=0.38
r162 4 35 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=5.545
+ $Y=0.235 $X2=5.67 $Y2=0.38
r163 3 31 91 $w=1.7e-07 $l=3.19374e-07 $layer=licon1_NDIFF $count=2 $X=4.31
+ $Y=0.235 $X2=4.565 $Y2=0.38
r164 2 27 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=2.44
+ $Y=0.235 $X2=2.58 $Y2=0.36
r165 1 23 182 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_NDIFF $count=1 $X=0.63
+ $Y=0.66 $X2=0.77 $Y2=0.855
.ends

