* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__nor4b_4 A B C D_N VGND VNB VPB VPWR Y
X0 a_1009_367# B a_644_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X1 VPWR A a_1009_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X2 VGND a_27_367# Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X3 Y a_27_367# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X4 VGND A Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X5 Y a_27_367# a_217_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X6 a_217_367# C a_644_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X7 a_217_367# a_27_367# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X8 VGND B Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X9 Y B VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X10 VPWR A a_1009_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X11 Y a_27_367# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X12 Y C VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X13 a_1009_367# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X14 VGND C Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X15 a_644_367# B a_1009_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X16 Y C VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X17 Y A VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X18 a_27_367# D_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X19 a_644_367# C a_217_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X20 a_217_367# C a_644_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X21 VGND A Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X22 VGND C Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X23 a_644_367# C a_217_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X24 a_27_367# D_N VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X25 Y A VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X26 a_644_367# B a_1009_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X27 a_1009_367# B a_644_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X28 VGND B Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X29 Y B VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X30 Y a_27_367# a_217_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X31 a_217_367# a_27_367# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X32 VGND a_27_367# Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X33 a_1009_367# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
.ends
