* File: sky130_fd_sc_lp__o31a_m.spice
* Created: Fri Aug 28 11:16:00 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__o31a_m.pex.spice"
.subckt sky130_fd_sc_lp__o31a_m  VNB VPB A1 A2 A3 B1 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* B1	B1
* A3	A3
* A2	A2
* A1	A1
* VPB	VPB
* VNB	VNB
MM1006 N_VGND_M1006_d N_A_95_153#_M1006_g N_X_M1006_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75002.3
+ A=0.063 P=1.14 MULT=1
MM1000 N_A_239_47#_M1000_d N_A1_M1000_g N_VGND_M1006_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6 SB=75001.9
+ A=0.063 P=1.14 MULT=1
MM1001 N_VGND_M1001_d N_A2_M1001_g N_A_239_47#_M1000_d VNB NSHORT L=0.15 W=0.42
+ AD=0.07875 AS=0.0588 PD=0.795 PS=0.7 NRD=5.712 NRS=0 M=1 R=2.8 SA=75001.1
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1007 N_A_239_47#_M1007_d N_A3_M1007_g N_VGND_M1001_d VNB NSHORT L=0.15 W=0.42
+ AD=0.07035 AS=0.07875 PD=0.755 PS=0.795 NRD=0 NRS=21.42 M=1 R=2.8 SA=75001.6
+ SB=75000.9 A=0.063 P=1.14 MULT=1
MM1005 N_A_95_153#_M1005_d N_B1_M1005_g N_A_239_47#_M1007_d VNB NSHORT L=0.15
+ W=0.42 AD=0.2058 AS=0.07035 PD=1.82 PS=0.755 NRD=64.284 NRS=15.708 M=1 R=2.8
+ SA=75002.1 SB=75000.4 A=0.063 P=1.14 MULT=1
MM1003 N_VPWR_M1003_d N_A_95_153#_M1003_g N_X_M1003_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0819 AS=0.1113 PD=0.81 PS=1.37 NRD=32.8202 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.2 A=0.063 P=1.14 MULT=1
MM1008 A_239_397# N_A1_M1008_g N_VPWR_M1003_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0441 AS=0.0819 PD=0.63 PS=0.81 NRD=23.443 NRS=18.7544 M=1 R=2.8
+ SA=75000.7 SB=75001.6 A=0.063 P=1.14 MULT=1
MM1004 A_311_397# N_A2_M1004_g A_239_397# VPB PHIGHVT L=0.15 W=0.42 AD=0.0819
+ AS=0.0441 PD=0.81 PS=0.63 NRD=65.6601 NRS=23.443 M=1 R=2.8 SA=75001.1
+ SB=75001.3 A=0.063 P=1.14 MULT=1
MM1009 N_A_95_153#_M1009_d N_A3_M1009_g A_311_397# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0819 AS=0.0819 PD=0.81 PS=0.81 NRD=0 NRS=65.6601 M=1 R=2.8 SA=75001.6
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1002 N_VPWR_M1002_d N_B1_M1002_g N_A_95_153#_M1009_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.1113 AS=0.0819 PD=1.37 PS=0.81 NRD=0 NRS=51.5943 M=1 R=2.8 SA=75002.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9751 P=11.21
c_41 VNB 0 3.11919e-19 $X=0 $Y=0
c_69 VPB 0 2.80181e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_lp__o31a_m.pxi.spice"
*
.ends
*
*
