* File: sky130_fd_sc_lp__o221ai_lp.spice
* Created: Wed Sep  2 10:19:26 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__o221ai_lp.pex.spice"
.subckt sky130_fd_sc_lp__o221ai_lp  VNB VPB C1 B1 B2 A2 A1 Y VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Y	Y
* A1	A1
* A2	A2
* B2	B2
* B1	B1
* C1	C1
* VPB	VPB
* VNB	VNB
MM1004 N_A_216_55#_M1004_d N_C1_M1004_g N_Y_M1004_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.1197 PD=0.7 PS=1.41 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75002.9
+ A=0.063 P=1.14 MULT=1
MM1006 N_A_302_55#_M1006_d N_B1_M1006_g N_A_216_55#_M1004_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0756 AS=0.0588 PD=0.78 PS=0.7 NRD=22.848 NRS=0 M=1 R=2.8
+ SA=75000.6 SB=75002.4 A=0.063 P=1.14 MULT=1
MM1000 N_VGND_M1000_d N_A2_M1000_g N_A_302_55#_M1006_d VNB NSHORT L=0.15 W=0.42
+ AD=0.22155 AS=0.0756 PD=1.475 PS=0.78 NRD=22.848 NRS=0 M=1 R=2.8 SA=75001.1
+ SB=75001.9 A=0.063 P=1.14 MULT=1
MM1009 N_A_302_55#_M1009_d N_A1_M1009_g N_VGND_M1000_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.22155 PD=0.7 PS=1.475 NRD=0 NRS=198.564 M=1 R=2.8 SA=75002.4
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1002 N_A_216_55#_M1002_d N_B2_M1002_g N_A_302_55#_M1009_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1533 AS=0.0588 PD=1.57 PS=0.7 NRD=22.848 NRS=0 M=1 R=2.8
+ SA=75002.8 SB=75000.3 A=0.063 P=1.14 MULT=1
MM1003 N_VPWR_M1003_d N_C1_M1003_g N_Y_M1003_s VPB PHIGHVT L=0.25 W=1 AD=0.1925
+ AS=0.285 PD=1.385 PS=2.57 NRD=0 NRS=0 M=1 R=4 SA=125000 SB=125002 A=0.25 P=2.5
+ MULT=1
MM1007 A_347_419# N_B1_M1007_g N_VPWR_M1003_d VPB PHIGHVT L=0.25 W=1 AD=0.12
+ AS=0.1925 PD=1.24 PS=1.385 NRD=12.7853 NRS=20.685 M=1 R=4 SA=125001 SB=125002
+ A=0.25 P=2.5 MULT=1
MM1001 N_Y_M1001_d N_B2_M1001_g A_347_419# VPB PHIGHVT L=0.25 W=1 AD=0.16
+ AS=0.12 PD=1.32 PS=1.24 NRD=0 NRS=12.7853 M=1 R=4 SA=125001 SB=125001 A=0.25
+ P=2.5 MULT=1
MM1005 A_559_419# N_A2_M1005_g N_Y_M1001_d VPB PHIGHVT L=0.25 W=1 AD=0.12
+ AS=0.16 PD=1.24 PS=1.32 NRD=12.7853 NRS=7.8603 M=1 R=4 SA=125002 SB=125001
+ A=0.25 P=2.5 MULT=1
MM1008 N_VPWR_M1008_d N_A1_M1008_g A_559_419# VPB PHIGHVT L=0.25 W=1 AD=0.285
+ AS=0.12 PD=2.57 PS=1.24 NRD=0 NRS=12.7853 M=1 R=4 SA=125002 SB=125000 A=0.25
+ P=2.5 MULT=1
DX10_noxref VNB VPB NWDIODE A=8.7655 P=13.13
*
.include "sky130_fd_sc_lp__o221ai_lp.pxi.spice"
*
.ends
*
*
