* File: sky130_fd_sc_lp__dfstp_4.spice
* Created: Wed Sep  2 09:44:34 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__dfstp_4.pex.spice"
.subckt sky130_fd_sc_lp__dfstp_4  VNB VPB CLK D SET_B VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* SET_B	SET_B
* D	D
* CLK	CLK
* VPB	VPB
* VNB	VNB
MM1013 N_VGND_M1013_d N_CLK_M1013_g N_A_30_99#_M1013_s VNB NSHORT L=0.15 W=0.42
+ AD=0.13545 AS=0.1113 PD=1.065 PS=1.37 NRD=104.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1001 N_A_230_465#_M1001_d N_A_30_99#_M1001_g N_VGND_M1013_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1113 AS=0.13545 PD=1.37 PS=1.065 NRD=0 NRS=0 M=1 R=2.8 SA=75001
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1037 N_A_476_119#_M1037_d N_D_M1037_g N_VGND_M1037_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75001.4
+ A=0.063 P=1.14 MULT=1
MM1002 N_A_562_119#_M1002_d N_A_30_99#_M1002_g N_A_476_119#_M1037_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.6 SB=75001 A=0.063 P=1.14 MULT=1
MM1027 A_648_119# N_A_230_465#_M1027_g N_A_562_119#_M1002_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75001.1
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1035 N_VGND_M1035_d N_A_690_93#_M1035_g A_648_119# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.4
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1007 A_914_47# N_A_562_119#_M1007_g N_A_690_93#_M1007_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.1113 PD=0.63 PS=1.37 NRD=14.28 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75002.8 A=0.063 P=1.14 MULT=1
MM1009 N_VGND_M1009_d N_SET_B_M1009_g A_914_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.1554 AS=0.0441 PD=1.13717 PS=0.63 NRD=148.56 NRS=14.28 M=1 R=2.8
+ SA=75000.6 SB=75002.5 A=0.063 P=1.14 MULT=1
MM1015 A_1175_47# N_A_562_119#_M1015_g N_VGND_M1009_d VNB NSHORT L=0.15 W=0.64
+ AD=0.0672 AS=0.2368 PD=0.85 PS=1.73283 NRD=9.372 NRS=0 M=1 R=4.26667 SA=75001
+ SB=75001.9 A=0.096 P=1.58 MULT=1
MM1018 N_A_1247_47#_M1018_d N_A_230_465#_M1018_g A_1175_47# VNB NSHORT L=0.15
+ W=0.64 AD=0.135366 AS=0.0672 PD=1.24981 PS=0.85 NRD=10.776 NRS=9.372 M=1
+ R=4.26667 SA=75001.4 SB=75001.5 A=0.096 P=1.58 MULT=1
MM1021 A_1356_91# N_A_30_99#_M1021_g N_A_1247_47#_M1018_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.088834 PD=0.63 PS=0.820189 NRD=14.28 NRS=17.136 M=1
+ R=2.8 SA=75001.7 SB=75001.7 A=0.063 P=1.14 MULT=1
MM1008 A_1428_91# N_A_1398_65#_M1008_g A_1356_91# VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0441 PD=0.63 PS=0.63 NRD=14.28 NRS=14.28 M=1 R=2.8 SA=75002.1
+ SB=75001.3 A=0.063 P=1.14 MULT=1
MM1034 N_VGND_M1034_d N_SET_B_M1034_g A_1428_91# VNB NSHORT L=0.15 W=0.42
+ AD=0.1302 AS=0.0441 PD=1.04 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75002.4
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1028 N_A_1398_65#_M1028_d N_A_1247_47#_M1028_g N_VGND_M1034_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.1113 AS=0.1302 PD=1.37 PS=1.04 NRD=0 NRS=0 M=1 R=2.8
+ SA=75003.2 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1012 N_VGND_M1012_d N_A_1247_47#_M1012_g N_A_1989_49#_M1012_s VNB NSHORT
+ L=0.15 W=0.84 AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6
+ SA=75000.2 SB=75001.9 A=0.126 P=1.98 MULT=1
MM1010 N_VGND_M1012_d N_A_1989_49#_M1010_g N_Q_M1010_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75001.5 A=0.126 P=1.98 MULT=1
MM1023 N_VGND_M1023_d N_A_1989_49#_M1023_g N_Q_M1010_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.1
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1029 N_VGND_M1023_d N_A_1989_49#_M1029_g N_Q_M1029_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.5
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1030 N_VGND_M1030_d N_A_1989_49#_M1030_g N_Q_M1029_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.9
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1005 N_VPWR_M1005_d N_CLK_M1005_g N_A_30_99#_M1005_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0896 AS=0.1824 PD=0.92 PS=1.85 NRD=0 NRS=6.1464 M=1 R=4.26667 SA=75000.2
+ SB=75000.6 A=0.096 P=1.58 MULT=1
MM1025 N_A_230_465#_M1025_d N_A_30_99#_M1025_g N_VPWR_M1005_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1696 AS=0.0896 PD=1.81 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.6 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1031 N_A_476_119#_M1031_d N_D_M1031_g N_VPWR_M1031_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0588 AS=0.10995 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75003.1 A=0.063 P=1.14 MULT=1
MM1019 N_A_562_119#_M1019_d N_A_230_465#_M1019_g N_A_476_119#_M1031_d VPB
+ PHIGHVT L=0.15 W=0.42 AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.6 SB=75002.6 A=0.063 P=1.14 MULT=1
MM1000 A_690_463# N_A_30_99#_M1000_g N_A_562_119#_M1019_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=23.443 NRS=0 M=1 R=2.8 SA=75001
+ SB=75002.2 A=0.063 P=1.14 MULT=1
MM1006 N_VPWR_M1006_d N_A_690_93#_M1006_g A_690_463# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.08295 AS=0.0441 PD=0.815 PS=0.63 NRD=9.3772 NRS=23.443 M=1 R=2.8
+ SA=75001.4 SB=75001.8 A=0.063 P=1.14 MULT=1
MM1016 N_A_690_93#_M1016_d N_A_562_119#_M1016_g N_VPWR_M1006_d VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.0588 AS=0.08295 PD=0.7 PS=0.815 NRD=0 NRS=44.5417 M=1 R=2.8
+ SA=75002 SB=75001.3 A=0.063 P=1.14 MULT=1
MM1003 N_VPWR_M1003_d N_SET_B_M1003_g N_A_690_93#_M1016_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.112 AS=0.0588 PD=0.916667 PS=0.7 NRD=120.761 NRS=0 M=1 R=2.8
+ SA=75002.4 SB=75000.9 A=0.063 P=1.14 MULT=1
MM1020 N_A_1094_379#_M1020_d N_A_562_119#_M1020_g N_VPWR_M1003_d VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.2226 AS=0.224 PD=2.21 PS=1.83333 NRD=0 NRS=0 M=1 R=5.6
+ SA=75001.6 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1036 N_A_1247_47#_M1036_d N_A_230_465#_M1036_g N_A_1201_407#_M1036_s VPB
+ PHIGHVT L=0.15 W=0.42 AD=0.0896 AS=0.1113 PD=0.81 PS=1.37 NRD=32.8202 NRS=0
+ M=1 R=2.8 SA=75000.2 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1026 N_A_1094_379#_M1026_d N_A_30_99#_M1026_g N_A_1247_47#_M1036_d VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.3599 AS=0.1792 PD=2.86 PS=1.62 NRD=87.5665 NRS=5.8509 M=1
+ R=5.6 SA=75000.5 SB=75000.3 A=0.126 P=1.98 MULT=1
MM1014 N_VPWR_M1014_d N_A_1398_65#_M1014_g N_A_1201_407#_M1014_s VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1032 N_A_1247_47#_M1032_d N_SET_B_M1032_g N_VPWR_M1014_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1024 N_A_1398_65#_M1024_d N_A_1247_47#_M1024_g N_VPWR_M1024_s VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.1113 AS=0.1113 PD=1.37 PS=1.37 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1011 N_VPWR_M1011_d N_A_1247_47#_M1011_g N_A_1989_49#_M1011_s VPB PHIGHVT
+ L=0.15 W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.2 SB=75001.9 A=0.189 P=2.82 MULT=1
MM1004 N_Q_M1004_d N_A_1989_49#_M1004_g N_VPWR_M1011_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75001.5 A=0.189 P=2.82 MULT=1
MM1017 N_Q_M1004_d N_A_1989_49#_M1017_g N_VPWR_M1017_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1022 N_Q_M1022_d N_A_1989_49#_M1022_g N_VPWR_M1017_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.5
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1033 N_Q_M1022_d N_A_1989_49#_M1033_g N_VPWR_M1033_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75001.9
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX38_noxref VNB VPB NWDIODE A=24.1503 P=29.77
c_129 VNB 0 1.22064e-19 $X=0 $Y=0
*
.include "sky130_fd_sc_lp__dfstp_4.pxi.spice"
*
.ends
*
*
