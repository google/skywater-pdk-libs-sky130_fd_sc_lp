# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__o22ai_4
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__o22ai_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.680000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 1.345000 1.455000 1.630000 ;
        RECT 1.025000 1.630000 1.455000 1.950000 ;
        RECT 1.025000 1.950000 3.555000 2.120000 ;
        RECT 3.385000 1.345000 3.715000 1.525000 ;
        RECT 3.385000 1.525000 3.555000 1.950000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.810000 1.345000 3.205000 1.750000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.955000 1.355000 5.125000 1.535000 ;
        RECT 3.995000 1.210000 5.125000 1.355000 ;
        RECT 4.885000 1.005000 7.195000 1.175000 ;
        RECT 4.885000 1.175000 5.125000 1.210000 ;
        RECT 6.930000 1.175000 7.195000 1.515000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.305000 1.345000 6.655000 1.535000 ;
        RECT 5.810000 1.535000 6.120000 1.760000 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  2.352000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.920000 2.290000 3.960000 2.470000 ;
        RECT 1.920000 2.470000 3.050000 2.620000 ;
        RECT 3.790000 1.705000 5.640000 1.875000 ;
        RECT 3.790000 1.875000 3.960000 2.290000 ;
        RECT 3.985000 0.645000 7.535000 0.835000 ;
        RECT 3.985000 0.835000 4.715000 1.040000 ;
        RECT 5.370000 1.875000 5.640000 1.930000 ;
        RECT 5.370000 1.930000 6.560000 2.100000 ;
        RECT 5.370000 2.100000 5.700000 2.735000 ;
        RECT 6.230000 2.100000 6.560000 2.735000 ;
        RECT 6.290000 1.705000 7.535000 1.875000 ;
        RECT 6.290000 1.875000 6.560000 1.930000 ;
        RECT 7.365000 0.835000 7.535000 1.705000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 7.680000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 7.680000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.680000 0.085000 ;
      RECT 0.000000  3.245000 7.680000 3.415000 ;
      RECT 0.125000  0.255000 0.385000 1.005000 ;
      RECT 0.125000  1.005000 3.815000 1.175000 ;
      RECT 0.140000  1.815000 0.430000 3.245000 ;
      RECT 0.555000  0.085000 0.885000 0.825000 ;
      RECT 0.600000  1.815000 0.855000 2.290000 ;
      RECT 0.600000  2.290000 1.700000 2.460000 ;
      RECT 0.600000  2.460000 0.830000 3.075000 ;
      RECT 1.000000  2.630000 1.330000 3.245000 ;
      RECT 1.055000  0.255000 1.245000 1.005000 ;
      RECT 1.415000  0.085000 1.745000 0.825000 ;
      RECT 1.500000  2.460000 1.700000 2.790000 ;
      RECT 1.500000  2.790000 3.480000 3.075000 ;
      RECT 1.915000  0.255000 2.105000 1.005000 ;
      RECT 2.275000  0.085000 2.605000 0.825000 ;
      RECT 2.775000  0.255000 2.965000 1.005000 ;
      RECT 3.135000  0.085000 3.465000 0.825000 ;
      RECT 3.635000  0.255000 7.390000 0.475000 ;
      RECT 3.635000  0.475000 3.815000 1.005000 ;
      RECT 3.650000  2.640000 3.960000 3.245000 ;
      RECT 4.130000  2.045000 5.200000 2.225000 ;
      RECT 4.130000  2.225000 4.340000 3.075000 ;
      RECT 4.510000  2.395000 4.840000 3.245000 ;
      RECT 5.010000  2.225000 5.200000 2.905000 ;
      RECT 5.010000  2.905000 6.920000 3.075000 ;
      RECT 5.870000  2.270000 6.060000 2.905000 ;
      RECT 6.730000  2.045000 6.920000 2.905000 ;
      RECT 7.090000  2.105000 7.420000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
  END
END sky130_fd_sc_lp__o22ai_4
END LIBRARY
