* File: sky130_fd_sc_lp__a2bb2o_1.spice
* Created: Wed Sep  2 09:23:43 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__a2bb2o_1.pex.spice"
.subckt sky130_fd_sc_lp__a2bb2o_1  VNB VPB A1_N A2_N B2 B1 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* B1	B1
* B2	B2
* A2_N	A2_N
* A1_N	A1_N
* VPB	VPB
* VNB	VNB
MM1011 N_VGND_M1011_d N_A_91_269#_M1011_g N_X_M1011_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2254 AS=0.2226 PD=1.84 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75001.5 A=0.126 P=1.98 MULT=1
MM1005 N_A_271_47#_M1005_d N_A1_N_M1005_g N_VGND_M1011_d VNB NSHORT L=0.15
+ W=0.42 AD=0.07035 AS=0.1127 PD=0.755 PS=0.92 NRD=15.708 NRS=74.28 M=1 R=2.8
+ SA=75000.9 SB=75002.2 A=0.063 P=1.14 MULT=1
MM1006 N_VGND_M1006_d N_A2_N_M1006_g N_A_271_47#_M1005_d VNB NSHORT L=0.15
+ W=0.42 AD=0.09135 AS=0.07035 PD=0.855 PS=0.755 NRD=21.42 NRS=0 M=1 R=2.8
+ SA=75001.4 SB=75001.7 A=0.063 P=1.14 MULT=1
MM1008 N_A_91_269#_M1008_d N_A_271_47#_M1008_g N_VGND_M1006_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0588 AS=0.09135 PD=0.7 PS=0.855 NRD=0 NRS=22.848 M=1 R=2.8
+ SA=75001.9 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1002 A_571_47# N_B2_M1002_g N_A_91_269#_M1008_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.0588 PD=0.66 PS=0.7 NRD=18.564 NRS=0 M=1 R=2.8 SA=75002.4
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1003 N_VGND_M1003_d N_B1_M1003_g A_571_47# VNB NSHORT L=0.15 W=0.42 AD=0.1554
+ AS=0.0504 PD=1.58 PS=0.66 NRD=30 NRS=18.564 M=1 R=2.8 SA=75002.8 SB=75000.3
+ A=0.063 P=1.14 MULT=1
MM1009 N_VPWR_M1009_d N_A_91_269#_M1009_g N_X_M1009_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.307125 AS=0.3339 PD=2.5575 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75000.5 A=0.189 P=2.82 MULT=1
MM1000 A_271_367# N_A1_N_M1000_g N_VPWR_M1009_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0504 AS=0.102375 PD=0.66 PS=0.8525 NRD=30.4759 NRS=88.5318 M=1 R=2.8
+ SA=75000.8 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1007 N_A_271_47#_M1007_d N_A2_N_M1007_g A_271_367# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.1113 AS=0.0504 PD=1.37 PS=0.66 NRD=0 NRS=30.4759 M=1 R=2.8 SA=75001.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1010 N_A_505_529#_M1010_d N_A_271_47#_M1010_g N_A_91_269#_M1010_s VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1004 N_VPWR_M1004_d N_B2_M1004_g N_A_505_529#_M1010_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1001 N_A_505_529#_M1001_d N_B1_M1001_g N_VPWR_M1004_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.1
+ SB=75000.2 A=0.063 P=1.14 MULT=1
DX12_noxref VNB VPB NWDIODE A=7.8703 P=12.17
c_50 VNB 0 6.51563e-20 $X=0 $Y=0
*
.include "sky130_fd_sc_lp__a2bb2o_1.pxi.spice"
*
.ends
*
*
