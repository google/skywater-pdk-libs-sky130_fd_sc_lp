* File: sky130_fd_sc_lp__mux2_m.pex.spice
* Created: Fri Aug 28 10:44:36 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__MUX2_M%A_123_269# 1 2 9 13 17 18 21 22 24 25 27 29
+ 34
c74 29 0 1.45779e-19 $X=1.805 $Y=0.9
c75 27 0 3.43691e-20 $X=2.03 $Y=2.525
r76 31 34 6.71292 $w=1.88e-07 $l=1.15e-07 $layer=LI1_cond $X=2.03 $Y=2.62
+ $X2=2.145 $Y2=2.62
r77 27 31 1.386 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.03 $Y=2.525 $X2=2.03
+ $Y2=2.62
r78 26 29 7.2619 $w=3.78e-07 $l=3.28786e-07 $layer=LI1_cond $X=2.03 $Y=1.265
+ $X2=1.805 $Y2=1.03
r79 26 27 82.2032 $w=1.68e-07 $l=1.26e-06 $layer=LI1_cond $X=2.03 $Y=1.265
+ $X2=2.03 $Y2=2.525
r80 24 29 9.06643 $w=3.78e-07 $l=2.2798e-07 $layer=LI1_cond $X=1.64 $Y=1.18
+ $X2=1.805 $Y2=1.03
r81 24 25 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=1.64 $Y=1.18
+ $X2=0.865 $Y2=1.18
r82 21 22 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.78
+ $Y=1.51 $X2=0.78 $Y2=1.51
r83 19 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.78 $Y=1.265
+ $X2=0.865 $Y2=1.18
r84 19 21 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=0.78 $Y=1.265
+ $X2=0.78 $Y2=1.51
r85 17 22 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.78 $Y=1.85
+ $X2=0.78 $Y2=1.51
r86 17 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.78 $Y=1.85
+ $X2=0.78 $Y2=2.015
r87 16 22 41.8716 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.78 $Y=1.345
+ $X2=0.78 $Y2=1.51
r88 13 18 358.936 $w=1.5e-07 $l=7e-07 $layer=POLY_cond $X=0.87 $Y=2.715 $X2=0.87
+ $Y2=2.015
r89 9 16 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=0.72 $Y=0.835
+ $X2=0.72 $Y2=1.345
r90 2 34 600 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=2.005
+ $Y=2.505 $X2=2.145 $Y2=2.63
r91 1 29 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=1.665
+ $Y=0.625 $X2=1.805 $Y2=0.9
.ends

.subckt PM_SKY130_FD_SC_LP__MUX2_M%S 3 7 11 15 19 20 22 23 24 26 28 29 32 33 34
+ 35 42 47
c106 32 0 4.59407e-20 $X=2.66 $Y=2.43
r107 42 43 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.28
+ $Y=1.745 $X2=3.28 $Y2=1.745
r108 35 47 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.2 $Y=2.43 $X2=3.2
+ $Y2=2.345
r109 35 47 0.453993 $w=3.28e-07 $l=1.3e-08 $layer=LI1_cond $X=3.2 $Y=2.332
+ $X2=3.2 $Y2=2.345
r110 34 35 10.372 $w=3.28e-07 $l=2.97e-07 $layer=LI1_cond $X=3.2 $Y=2.035
+ $X2=3.2 $Y2=2.332
r111 34 43 10.1275 $w=3.28e-07 $l=2.9e-07 $layer=LI1_cond $X=3.2 $Y=2.035
+ $X2=3.2 $Y2=1.745
r112 33 43 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=3.2 $Y=1.665 $X2=3.2
+ $Y2=1.745
r113 32 35 15.0571 $w=3.13e-07 $l=3.75e-07 $layer=LI1_cond $X=2.66 $Y=2.43
+ $X2=3.035 $Y2=2.43
r114 29 46 18.1887 $w=3.18e-07 $l=1.2e-07 $layer=POLY_cond $X=1.45 $Y=2.18
+ $X2=1.57 $Y2=2.18
r115 29 44 33.3459 $w=3.18e-07 $l=2.2e-07 $layer=POLY_cond $X=1.45 $Y=2.18
+ $X2=1.23 $Y2=2.18
r116 28 31 8.74048 $w=2.53e-07 $l=1.65e-07 $layer=LI1_cond $X=1.492 $Y=2.18
+ $X2=1.492 $Y2=2.345
r117 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.45
+ $Y=2.18 $X2=1.45 $Y2=2.18
r118 25 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.575 $Y=2.515
+ $X2=2.66 $Y2=2.43
r119 25 26 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=2.575 $Y=2.515
+ $X2=2.575 $Y2=2.895
r120 23 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.49 $Y=2.98
+ $X2=2.575 $Y2=2.895
r121 23 24 56.7594 $w=1.68e-07 $l=8.7e-07 $layer=LI1_cond $X=2.49 $Y=2.98
+ $X2=1.62 $Y2=2.98
r122 22 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.535 $Y=2.895
+ $X2=1.62 $Y2=2.98
r123 22 31 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=1.535 $Y=2.895
+ $X2=1.535 $Y2=2.345
r124 19 42 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=3.28 $Y=2.085
+ $X2=3.28 $Y2=1.745
r125 19 20 41.8716 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.28 $Y=2.085
+ $X2=3.28 $Y2=2.25
r126 18 42 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.28 $Y=1.58
+ $X2=3.28 $Y2=1.745
r127 15 20 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.34 $Y=2.715
+ $X2=3.34 $Y2=2.25
r128 11 18 382.011 $w=1.5e-07 $l=7.45e-07 $layer=POLY_cond $X=3.19 $Y=0.835
+ $X2=3.19 $Y2=1.58
r129 5 46 20.3436 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.57 $Y=2.345
+ $X2=1.57 $Y2=2.18
r130 5 7 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=1.57 $Y=2.345
+ $X2=1.57 $Y2=2.715
r131 1 44 20.3436 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.23 $Y=2.015
+ $X2=1.23 $Y2=2.18
r132 1 3 605.064 $w=1.5e-07 $l=1.18e-06 $layer=POLY_cond $X=1.23 $Y=2.015
+ $X2=1.23 $Y2=0.835
.ends

.subckt PM_SKY130_FD_SC_LP__MUX2_M%A1 3 6 8 11 14 15 19 21
c59 19 0 1.6437e-19 $X=1.68 $Y=0.515
c60 6 0 1.91956e-19 $X=2.36 $Y=2.715
r61 21 24 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.38 $Y=2 $X2=2.38
+ $Y2=2.165
r62 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.38 $Y=2
+ $X2=2.38 $Y2=2
r63 15 22 9.07985 $w=3.28e-07 $l=2.6e-07 $layer=LI1_cond $X=2.64 $Y=2 $X2=2.38
+ $Y2=2
r64 14 22 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.38 $Y=1.835
+ $X2=2.38 $Y2=2
r65 13 14 91.3369 $w=1.68e-07 $l=1.4e-06 $layer=LI1_cond $X=2.38 $Y=0.435
+ $X2=2.38 $Y2=1.835
r66 11 19 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.68 $Y=0.35
+ $X2=1.68 $Y2=0.515
r67 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.68
+ $Y=0.35 $X2=1.68 $Y2=0.35
r68 8 13 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.295 $Y=0.35
+ $X2=2.38 $Y2=0.435
r69 8 10 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=2.295 $Y=0.35
+ $X2=1.68 $Y2=0.35
r70 6 24 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=2.36 $Y=2.715
+ $X2=2.36 $Y2=2.165
r71 3 19 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.59 $Y=0.835
+ $X2=1.59 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LP__MUX2_M%A0 3 7 9 10 12 13
c43 13 0 1.6437e-19 $X=1.68 $Y=1.665
r44 13 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.68
+ $Y=1.61 $X2=1.68 $Y2=1.61
r45 12 13 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=1.2 $Y=1.61 $X2=1.68
+ $Y2=1.61
r46 10 11 42.467 $w=2.27e-07 $l=2e-07 $layer=POLY_cond $X=1.93 $Y=1.595 $X2=2.13
+ $Y2=1.595
r47 9 17 30.6007 $w=3.3e-07 $l=1.75e-07 $layer=POLY_cond $X=1.855 $Y=1.61
+ $X2=1.68 $Y2=1.61
r48 9 10 15.6896 $w=3.3e-07 $l=8.21584e-08 $layer=POLY_cond $X=1.855 $Y=1.61
+ $X2=1.93 $Y2=1.595
r49 5 11 12.4931 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=2.13 $Y=1.445
+ $X2=2.13 $Y2=1.595
r50 5 7 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.13 $Y=1.445 $X2=2.13
+ $Y2=0.835
r51 1 10 12.4931 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=1.93 $Y=1.775
+ $X2=1.93 $Y2=1.595
r52 1 3 482 $w=1.5e-07 $l=9.4e-07 $layer=POLY_cond $X=1.93 $Y=1.775 $X2=1.93
+ $Y2=2.715
.ends

.subckt PM_SKY130_FD_SC_LP__MUX2_M%A_483_99# 1 2 7 9 12 14 16 17 20 21 29
c57 21 0 3.43691e-20 $X=2.74 $Y=1.32
c58 7 0 1.45779e-19 $X=2.49 $Y=1.155
r59 27 29 4.22511 $w=2.08e-07 $l=8e-08 $layer=LI1_cond $X=3.555 $Y=2.775
+ $X2=3.635 $Y2=2.775
r60 24 25 10.9735 $w=3.78e-07 $l=3.4e-07 $layer=LI1_cond $X=3.48 $Y=0.9 $X2=3.48
+ $Y2=1.24
r61 21 33 16.0074 $w=2.71e-07 $l=9e-08 $layer=POLY_cond $X=2.74 $Y=1.32 $X2=2.83
+ $Y2=1.32
r62 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.74
+ $Y=1.32 $X2=2.74 $Y2=1.32
r63 17 29 1.9771 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=3.635 $Y=2.67
+ $X2=3.635 $Y2=2.775
r64 16 25 6.48442 $w=3.78e-07 $l=1.92873e-07 $layer=LI1_cond $X=3.635 $Y=1.325
+ $X2=3.48 $Y2=1.24
r65 16 17 87.7487 $w=1.68e-07 $l=1.345e-06 $layer=LI1_cond $X=3.635 $Y=1.325
+ $X2=3.635 $Y2=2.67
r66 15 20 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.825 $Y=1.24
+ $X2=2.74 $Y2=1.24
r67 14 25 5.4359 $w=1.7e-07 $l=2.4e-07 $layer=LI1_cond $X=3.24 $Y=1.24 $X2=3.48
+ $Y2=1.24
r68 14 15 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=3.24 $Y=1.24
+ $X2=2.825 $Y2=1.24
r69 10 33 16.5906 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.83 $Y=1.485
+ $X2=2.83 $Y2=1.32
r70 10 12 630.702 $w=1.5e-07 $l=1.23e-06 $layer=POLY_cond $X=2.83 $Y=1.485
+ $X2=2.83 $Y2=2.715
r71 7 21 44.4649 $w=2.71e-07 $l=3.22102e-07 $layer=POLY_cond $X=2.49 $Y=1.155
+ $X2=2.74 $Y2=1.32
r72 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.49 $Y=1.155 $X2=2.49
+ $Y2=0.835
r73 2 27 600 $w=1.7e-07 $l=3.32716e-07 $layer=licon1_PDIFF $count=1 $X=3.415
+ $Y=2.505 $X2=3.555 $Y2=2.775
r74 1 24 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=3.265
+ $Y=0.625 $X2=3.405 $Y2=0.9
.ends

.subckt PM_SKY130_FD_SC_LP__MUX2_M%X 1 2 11 13 14 15 16 17 36
r17 17 36 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=0.24 $Y=2.695
+ $X2=0.655 $Y2=2.695
r18 17 23 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.24 $Y=2.695
+ $X2=0.24 $Y2=2.53
r19 16 23 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=0.24 $Y=2.405
+ $X2=0.24 $Y2=2.53
r20 15 16 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.24 $Y=2.035
+ $X2=0.24 $Y2=2.405
r21 14 15 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.24 $Y=1.665
+ $X2=0.24 $Y2=2.035
r22 13 14 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.24 $Y=1.295
+ $X2=0.24 $Y2=1.665
r23 8 13 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=0.24 $Y=0.915
+ $X2=0.24 $Y2=1.295
r24 7 11 9.25447 $w=3.28e-07 $l=2.65e-07 $layer=LI1_cond $X=0.24 $Y=0.75
+ $X2=0.505 $Y2=0.75
r25 7 8 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.24 $Y=0.75 $X2=0.24
+ $Y2=0.915
r26 2 36 600 $w=1.7e-07 $l=2.44643e-07 $layer=licon1_PDIFF $count=1 $X=0.53
+ $Y=2.505 $X2=0.655 $Y2=2.695
r27 1 11 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.36
+ $Y=0.625 $X2=0.505 $Y2=0.75
.ends

.subckt PM_SKY130_FD_SC_LP__MUX2_M%VPWR 1 2 9 13 15 17 22 29 30 33 36
c41 13 0 1.91956e-19 $X=3.045 $Y=2.78
r42 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r43 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r44 30 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=3.12 $Y2=3.33
r45 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r46 27 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.21 $Y=3.33
+ $X2=3.045 $Y2=3.33
r47 27 29 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=3.21 $Y=3.33 $X2=3.6
+ $Y2=3.33
r48 26 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r49 25 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r50 23 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.27 $Y=3.33
+ $X2=1.105 $Y2=3.33
r51 23 25 89.3797 $w=1.68e-07 $l=1.37e-06 $layer=LI1_cond $X=1.27 $Y=3.33
+ $X2=2.64 $Y2=3.33
r52 22 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.88 $Y=3.33
+ $X2=3.045 $Y2=3.33
r53 22 25 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=2.88 $Y=3.33
+ $X2=2.64 $Y2=3.33
r54 20 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r55 19 20 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r56 17 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.94 $Y=3.33
+ $X2=1.105 $Y2=3.33
r57 17 19 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=0.94 $Y=3.33
+ $X2=0.72 $Y2=3.33
r58 15 26 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=2.64 $Y2=3.33
r59 15 34 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=1.2 $Y2=3.33
r60 11 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.045 $Y=3.245
+ $X2=3.045 $Y2=3.33
r61 11 13 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=3.045 $Y=3.245
+ $X2=3.045 $Y2=2.78
r62 7 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.105 $Y=3.245
+ $X2=1.105 $Y2=3.33
r63 7 9 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=1.105 $Y=3.245
+ $X2=1.105 $Y2=2.78
r64 2 13 600 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=1 $X=2.905
+ $Y=2.505 $X2=3.045 $Y2=2.78
r65 1 9 600 $w=1.7e-07 $l=3.45868e-07 $layer=licon1_PDIFF $count=1 $X=0.945
+ $Y=2.505 $X2=1.105 $Y2=2.78
.ends

.subckt PM_SKY130_FD_SC_LP__MUX2_M%VGND 1 2 9 13 16 17 19 20 21 34 35
r39 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r40 32 35 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r41 31 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r42 28 31 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.64
+ $Y2=0
r43 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r44 25 29 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r45 24 25 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r46 21 32 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=2.64
+ $Y2=0
r47 21 29 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=1.2
+ $Y2=0
r48 19 31 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=2.645 $Y=0 $X2=2.64
+ $Y2=0
r49 19 20 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.645 $Y=0 $X2=2.81
+ $Y2=0
r50 18 34 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=2.975 $Y=0 $X2=3.6
+ $Y2=0
r51 18 20 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.975 $Y=0 $X2=2.81
+ $Y2=0
r52 16 24 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=0.79 $Y=0 $X2=0.72
+ $Y2=0
r53 16 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.79 $Y=0 $X2=0.955
+ $Y2=0
r54 15 28 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=1.12 $Y=0 $X2=1.2
+ $Y2=0
r55 15 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.12 $Y=0 $X2=0.955
+ $Y2=0
r56 11 20 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.81 $Y=0.085
+ $X2=2.81 $Y2=0
r57 11 13 23.9219 $w=3.28e-07 $l=6.85e-07 $layer=LI1_cond $X=2.81 $Y=0.085
+ $X2=2.81 $Y2=0.77
r58 7 17 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.955 $Y=0.085
+ $X2=0.955 $Y2=0
r59 7 9 23.9219 $w=3.28e-07 $l=6.85e-07 $layer=LI1_cond $X=0.955 $Y=0.085
+ $X2=0.955 $Y2=0.77
r60 2 13 182 $w=1.7e-07 $l=3.09112e-07 $layer=licon1_NDIFF $count=1 $X=2.565
+ $Y=0.625 $X2=2.81 $Y2=0.77
r61 1 9 182 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_NDIFF $count=1 $X=0.795
+ $Y=0.625 $X2=0.955 $Y2=0.77
.ends

