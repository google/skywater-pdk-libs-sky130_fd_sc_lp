* File: sky130_fd_sc_lp__o2bb2ai_1.pex.spice
* Created: Fri Aug 28 11:12:34 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O2BB2AI_1%A1_N 3 6 8 9 13 15
r26 13 16 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=0.387 $Y=1.375
+ $X2=0.387 $Y2=1.54
r27 13 15 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=0.387 $Y=1.375
+ $X2=0.387 $Y2=1.21
r28 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.365
+ $Y=1.375 $X2=0.365 $Y2=1.375
r29 9 14 9.1564 $w=3.63e-07 $l=2.9e-07 $layer=LI1_cond $X=0.267 $Y=1.665
+ $X2=0.267 $Y2=1.375
r30 8 14 2.5259 $w=3.63e-07 $l=8e-08 $layer=LI1_cond $X=0.267 $Y=1.295 $X2=0.267
+ $Y2=1.375
r31 6 16 474.309 $w=1.5e-07 $l=9.25e-07 $layer=POLY_cond $X=0.5 $Y=2.465 $X2=0.5
+ $Y2=1.54
r32 3 15 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.5 $Y=0.68 $X2=0.5
+ $Y2=1.21
.ends

.subckt PM_SKY130_FD_SC_LP__O2BB2AI_1%A2_N 3 6 8 11 12 13
c34 12 0 3.78943e-20 $X=0.95 $Y=1.375
r35 11 14 46.5827 $w=3.6e-07 $l=1.65e-07 $layer=POLY_cond $X=0.965 $Y=1.375
+ $X2=0.965 $Y2=1.54
r36 11 13 46.5827 $w=3.6e-07 $l=1.65e-07 $layer=POLY_cond $X=0.965 $Y=1.375
+ $X2=0.965 $Y2=1.21
r37 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.95
+ $Y=1.375 $X2=0.95 $Y2=1.375
r38 8 12 8.03218 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=0.72 $Y=1.375
+ $X2=0.95 $Y2=1.375
r39 6 14 474.309 $w=1.5e-07 $l=9.25e-07 $layer=POLY_cond $X=0.93 $Y=2.465
+ $X2=0.93 $Y2=1.54
r40 3 13 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.86 $Y=0.68 $X2=0.86
+ $Y2=1.21
.ends

.subckt PM_SKY130_FD_SC_LP__O2BB2AI_1%A_115_367# 1 2 9 13 15 16 19 23 24 27 31
+ 33 37 39
c74 16 0 1.30365e-19 $X=1.83 $Y=1.285
c75 15 0 3.78943e-20 $X=1.83 $Y=1.48
r76 37 39 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=1.29 $Y=1.04
+ $X2=1.29 $Y2=1.405
r77 36 37 10.3829 $w=3.28e-07 $l=2.2e-07 $layer=LI1_cond $X=1.18 $Y=0.82
+ $X2=1.18 $Y2=1.04
r78 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.595
+ $Y=1.51 $X2=1.595 $Y2=1.51
r79 31 40 15.8442 $w=2.08e-07 $l=3e-07 $layer=LI1_cond $X=1.31 $Y=1.54 $X2=1.31
+ $Y2=1.84
r80 31 39 7.56475 $w=2.08e-07 $l=1.35e-07 $layer=LI1_cond $X=1.31 $Y=1.54
+ $X2=1.31 $Y2=1.405
r81 31 33 7.68295 $w=2.68e-07 $l=1.8e-07 $layer=LI1_cond $X=1.415 $Y=1.54
+ $X2=1.595 $Y2=1.54
r82 27 36 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=1.15 $Y=0.405
+ $X2=1.15 $Y2=0.82
r83 23 40 1.9771 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.205 $Y=1.84
+ $X2=1.31 $Y2=1.84
r84 23 24 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=1.205 $Y=1.84
+ $X2=0.81 $Y2=1.84
r85 19 21 54.2871 $w=1.88e-07 $l=9.3e-07 $layer=LI1_cond $X=0.715 $Y=1.98
+ $X2=0.715 $Y2=2.91
r86 17 24 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=0.715 $Y=1.925
+ $X2=0.81 $Y2=1.84
r87 17 19 3.21053 $w=1.88e-07 $l=5.5e-08 $layer=LI1_cond $X=0.715 $Y=1.925
+ $X2=0.715 $Y2=1.98
r88 15 34 33.5118 $w=3.9e-07 $l=2.35e-07 $layer=POLY_cond $X=1.83 $Y=1.48
+ $X2=1.595 $Y2=1.48
r89 15 16 6.9036 $w=3.9e-07 $l=1.95e-07 $layer=POLY_cond $X=1.83 $Y=1.48
+ $X2=1.83 $Y2=1.285
r90 11 16 41.3382 $w=1.5e-07 $l=4.39375e-07 $layer=POLY_cond $X=1.935 $Y=1.675
+ $X2=1.83 $Y2=1.285
r91 11 13 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.935 $Y=1.675
+ $X2=1.935 $Y2=2.465
r92 7 16 41.3382 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.905 $Y=1.285
+ $X2=1.83 $Y2=1.285
r93 7 9 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=1.905 $Y=1.285
+ $X2=1.905 $Y2=0.655
r94 2 21 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=0.575
+ $Y=1.835 $X2=0.715 $Y2=2.91
r95 2 19 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.575
+ $Y=1.835 $X2=0.715 $Y2=1.98
r96 1 27 91 $w=1.7e-07 $l=2.78209e-07 $layer=licon1_NDIFF $count=2 $X=0.935
+ $Y=0.26 $X2=1.15 $Y2=0.405
.ends

.subckt PM_SKY130_FD_SC_LP__O2BB2AI_1%B2 3 7 9 11 12 13 21 27
c44 21 0 1.9443e-19 $X=2.415 $Y=1.375
c45 7 0 1.58364e-19 $X=2.445 $Y=2.465
c46 3 0 1.60614e-20 $X=2.335 $Y=0.655
r47 25 38 3.97524 $w=2.3e-07 $l=2e-07 $layer=LI1_cond $X=2.62 $Y=1.585 $X2=2.62
+ $Y2=1.385
r48 25 27 4.0085 $w=2.28e-07 $l=8e-08 $layer=LI1_cond $X=2.62 $Y=1.585 $X2=2.62
+ $Y2=1.665
r49 22 38 5.90627 $w=3.98e-07 $l=2.05e-07 $layer=LI1_cond $X=2.415 $Y=1.385
+ $X2=2.62 $Y2=1.385
r50 21 24 46.5827 $w=3.6e-07 $l=1.65e-07 $layer=POLY_cond $X=2.4 $Y=1.375
+ $X2=2.4 $Y2=1.54
r51 21 23 46.5827 $w=3.6e-07 $l=1.65e-07 $layer=POLY_cond $X=2.4 $Y=1.375
+ $X2=2.4 $Y2=1.21
r52 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.415
+ $Y=1.375 $X2=2.415 $Y2=1.375
r53 12 13 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=2.62 $Y=2.405
+ $X2=2.62 $Y2=2.775
r54 11 12 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=2.62 $Y=2.035
+ $X2=2.62 $Y2=2.405
r55 9 38 0.576222 $w=3.98e-07 $l=2e-08 $layer=LI1_cond $X=2.64 $Y=1.385 $X2=2.62
+ $Y2=1.385
r56 9 11 18.4391 $w=2.28e-07 $l=3.68e-07 $layer=LI1_cond $X=2.62 $Y=1.667
+ $X2=2.62 $Y2=2.035
r57 9 27 0.100212 $w=2.28e-07 $l=2e-09 $layer=LI1_cond $X=2.62 $Y=1.667 $X2=2.62
+ $Y2=1.665
r58 7 24 474.309 $w=1.5e-07 $l=9.25e-07 $layer=POLY_cond $X=2.445 $Y=2.465
+ $X2=2.445 $Y2=1.54
r59 3 23 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=2.335 $Y=0.655
+ $X2=2.335 $Y2=1.21
.ends

.subckt PM_SKY130_FD_SC_LP__O2BB2AI_1%B1 3 7 9 10 14
c27 9 0 1.74426e-19 $X=3.12 $Y=1.295
r28 14 17 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=2.972 $Y=1.375
+ $X2=2.972 $Y2=1.54
r29 14 16 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=2.972 $Y=1.375
+ $X2=2.972 $Y2=1.21
r30 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.99
+ $Y=1.375 $X2=2.99 $Y2=1.375
r31 10 15 9.03266 $w=3.68e-07 $l=2.9e-07 $layer=LI1_cond $X=3.09 $Y=1.665
+ $X2=3.09 $Y2=1.375
r32 9 15 2.49177 $w=3.68e-07 $l=8e-08 $layer=LI1_cond $X=3.09 $Y=1.295 $X2=3.09
+ $Y2=1.375
r33 7 17 474.309 $w=1.5e-07 $l=9.25e-07 $layer=POLY_cond $X=2.865 $Y=2.465
+ $X2=2.865 $Y2=1.54
r34 3 16 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=2.865 $Y=0.655
+ $X2=2.865 $Y2=1.21
.ends

.subckt PM_SKY130_FD_SC_LP__O2BB2AI_1%VPWR 1 2 3 10 12 18 22 24 28 30 35 44 48
r46 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r47 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r48 39 48 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r49 38 39 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r50 36 44 14.9939 $w=1.7e-07 $l=4.2e-07 $layer=LI1_cond $X=1.82 $Y=3.33 $X2=1.4
+ $Y2=3.33
r51 36 38 53.4973 $w=1.68e-07 $l=8.2e-07 $layer=LI1_cond $X=1.82 $Y=3.33
+ $X2=2.64 $Y2=3.33
r52 35 47 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=2.915 $Y=3.33
+ $X2=3.137 $Y2=3.33
r53 35 38 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=2.915 $Y=3.33
+ $X2=2.64 $Y2=3.33
r54 34 42 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r55 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r56 31 41 4.72267 $w=1.7e-07 $l=2.25e-07 $layer=LI1_cond $X=0.45 $Y=3.33
+ $X2=0.225 $Y2=3.33
r57 31 33 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=0.45 $Y=3.33 $X2=0.72
+ $Y2=3.33
r58 30 44 14.9939 $w=1.7e-07 $l=4.2e-07 $layer=LI1_cond $X=0.98 $Y=3.33 $X2=1.4
+ $Y2=3.33
r59 30 33 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=0.98 $Y=3.33
+ $X2=0.72 $Y2=3.33
r60 28 39 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r61 28 34 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.72 $Y2=3.33
r62 28 44 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r63 24 27 33.0018 $w=3.28e-07 $l=9.45e-07 $layer=LI1_cond $X=3.08 $Y=2.005
+ $X2=3.08 $Y2=2.95
r64 22 47 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=3.08 $Y=3.245
+ $X2=3.137 $Y2=3.33
r65 22 27 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=3.08 $Y=3.245
+ $X2=3.08 $Y2=2.95
r66 18 21 10.9641 $w=8.38e-07 $l=7.7e-07 $layer=LI1_cond $X=1.4 $Y=2.18 $X2=1.4
+ $Y2=2.95
r67 16 44 3.22441 $w=8.4e-07 $l=8.5e-08 $layer=LI1_cond $X=1.4 $Y=3.245 $X2=1.4
+ $Y2=3.33
r68 16 21 4.20051 $w=8.38e-07 $l=2.95e-07 $layer=LI1_cond $X=1.4 $Y=3.245
+ $X2=1.4 $Y2=2.95
r69 12 15 33.0018 $w=3.28e-07 $l=9.45e-07 $layer=LI1_cond $X=0.285 $Y=2.005
+ $X2=0.285 $Y2=2.95
r70 10 41 3.0435 $w=3.3e-07 $l=1.11018e-07 $layer=LI1_cond $X=0.285 $Y=3.245
+ $X2=0.225 $Y2=3.33
r71 10 15 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.285 $Y=3.245
+ $X2=0.285 $Y2=2.95
r72 3 27 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=2.94
+ $Y=1.835 $X2=3.08 $Y2=2.95
r73 3 24 400 $w=1.7e-07 $l=2.29565e-07 $layer=licon1_PDIFF $count=1 $X=2.94
+ $Y=1.835 $X2=3.08 $Y2=2.005
r74 2 21 200 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=3 $X=1.005
+ $Y=1.835 $X2=1.145 $Y2=2.95
r75 2 18 200 $w=1.7e-07 $l=4.09054e-07 $layer=licon1_PDIFF $count=3 $X=1.005
+ $Y=1.835 $X2=1.145 $Y2=2.18
r76 1 15 400 $w=1.7e-07 $l=1.17584e-06 $layer=licon1_PDIFF $count=1 $X=0.16
+ $Y=1.835 $X2=0.285 $Y2=2.95
r77 1 12 400 $w=1.7e-07 $l=2.23942e-07 $layer=licon1_PDIFF $count=1 $X=0.16
+ $Y=1.835 $X2=0.285 $Y2=2.005
.ends

.subckt PM_SKY130_FD_SC_LP__O2BB2AI_1%Y 1 2 12 15 16 17 18 19 20 21 41
c39 12 0 3.24794e-19 $X=2.015 $Y=1.15
r40 21 38 4.50956 $w=3.43e-07 $l=1.35e-07 $layer=LI1_cond $X=2.162 $Y=2.775
+ $X2=2.162 $Y2=2.91
r41 20 21 12.3595 $w=3.43e-07 $l=3.7e-07 $layer=LI1_cond $X=2.162 $Y=2.405
+ $X2=2.162 $Y2=2.775
r42 19 20 14.1968 $w=3.43e-07 $l=4.25e-07 $layer=LI1_cond $X=2.162 $Y=1.98
+ $X2=2.162 $Y2=2.405
r43 18 45 13.2051 $w=2.38e-07 $l=2.75e-07 $layer=LI1_cond $X=1.665 $Y=0.925
+ $X2=1.665 $Y2=0.65
r44 17 45 4.29829 $w=2.58e-07 $l=9.5e-08 $layer=LI1_cond $X=1.655 $Y=0.555
+ $X2=1.655 $Y2=0.65
r45 17 41 5.98384 $w=2.58e-07 $l=1.35e-07 $layer=LI1_cond $X=1.655 $Y=0.555
+ $X2=1.655 $Y2=0.42
r46 16 19 1.83723 $w=3.43e-07 $l=5.5e-08 $layer=LI1_cond $X=2.162 $Y=1.925
+ $X2=2.162 $Y2=1.98
r47 15 16 8.64642 $w=3.43e-07 $l=1.7e-07 $layer=LI1_cond $X=2.132 $Y=1.755
+ $X2=2.132 $Y2=1.925
r48 10 18 6.72258 $w=2.38e-07 $l=1.4e-07 $layer=LI1_cond $X=1.665 $Y=1.065
+ $X2=1.665 $Y2=0.925
r49 10 12 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=1.665 $Y=1.15
+ $X2=2.015 $Y2=1.15
r50 7 12 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.015 $Y=1.235
+ $X2=2.015 $Y2=1.15
r51 7 15 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=2.015 $Y=1.235
+ $X2=2.015 $Y2=1.755
r52 2 38 400 $w=1.7e-07 $l=1.15223e-06 $layer=licon1_PDIFF $count=1 $X=2.01
+ $Y=1.835 $X2=2.17 $Y2=2.91
r53 2 19 400 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_PDIFF $count=1 $X=2.01
+ $Y=1.835 $X2=2.17 $Y2=1.98
r54 1 41 91 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=2 $X=1.565
+ $Y=0.235 $X2=1.69 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__O2BB2AI_1%VGND 1 2 7 9 13 15 17 27 28 34
r41 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r42 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r43 28 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.64
+ $Y2=0
r44 27 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r45 25 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.785 $Y=0 $X2=2.62
+ $Y2=0
r46 25 27 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=2.785 $Y=0 $X2=3.12
+ $Y2=0
r47 24 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r48 23 24 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r49 21 32 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r50 20 23 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=0.72 $Y=0 $X2=2.16
+ $Y2=0
r51 20 21 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r52 18 31 4.72267 $w=1.7e-07 $l=2.25e-07 $layer=LI1_cond $X=0.45 $Y=0 $X2=0.225
+ $Y2=0
r53 18 20 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=0.45 $Y=0 $X2=0.72
+ $Y2=0
r54 17 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.455 $Y=0 $X2=2.62
+ $Y2=0
r55 17 23 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=2.455 $Y=0 $X2=2.16
+ $Y2=0
r56 15 24 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r57 15 21 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=0.72
+ $Y2=0
r58 11 34 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.62 $Y=0.085
+ $X2=2.62 $Y2=0
r59 11 13 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=2.62 $Y=0.085
+ $X2=2.62 $Y2=0.43
r60 7 31 3.0435 $w=3.3e-07 $l=1.11018e-07 $layer=LI1_cond $X=0.285 $Y=0.085
+ $X2=0.225 $Y2=0
r61 7 9 11.1752 $w=3.28e-07 $l=3.2e-07 $layer=LI1_cond $X=0.285 $Y=0.085
+ $X2=0.285 $Y2=0.405
r62 2 13 182 $w=1.7e-07 $l=2.91633e-07 $layer=licon1_NDIFF $count=1 $X=2.41
+ $Y=0.235 $X2=2.62 $Y2=0.43
r63 1 9 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.16
+ $Y=0.26 $X2=0.285 $Y2=0.405
.ends

.subckt PM_SKY130_FD_SC_LP__O2BB2AI_1%A_396_47# 1 2 7 9 11 14
r25 14 15 21.0647 $w=2.78e-07 $l=4.8e-07 $layer=LI1_cond $X=2.12 $Y=0.39
+ $X2=2.12 $Y2=0.87
r26 9 17 3.53583 $w=2.7e-07 $l=1.45e-07 $layer=LI1_cond $X=3.11 $Y=0.725
+ $X2=3.11 $Y2=0.87
r27 9 11 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=3.11 $Y=0.725
+ $X2=3.11 $Y2=0.43
r28 8 15 0.45714 $w=2.9e-07 $l=1.65e-07 $layer=LI1_cond $X=2.285 $Y=0.87
+ $X2=2.12 $Y2=0.87
r29 7 17 3.29198 $w=2.9e-07 $l=1.35e-07 $layer=LI1_cond $X=2.975 $Y=0.87
+ $X2=3.11 $Y2=0.87
r30 7 8 27.4202 $w=2.88e-07 $l=6.9e-07 $layer=LI1_cond $X=2.975 $Y=0.87
+ $X2=2.285 $Y2=0.87
r31 2 17 182 $w=1.7e-07 $l=7.61791e-07 $layer=licon1_NDIFF $count=1 $X=2.94
+ $Y=0.235 $X2=3.08 $Y2=0.93
r32 2 11 182 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_NDIFF $count=1 $X=2.94
+ $Y=0.235 $X2=3.08 $Y2=0.43
r33 1 14 91 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=2 $X=1.98
+ $Y=0.235 $X2=2.12 $Y2=0.39
.ends

