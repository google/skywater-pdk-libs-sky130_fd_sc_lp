* File: sky130_fd_sc_lp__nor2_0.pxi.spice
* Created: Wed Sep  2 10:07:16 2020
* 
x_PM_SKY130_FD_SC_LP__NOR2_0%A N_A_c_29_n N_A_M1003_g N_A_M1001_g N_A_c_31_n A A
+ A A N_A_c_33_n N_A_c_34_n PM_SKY130_FD_SC_LP__NOR2_0%A
x_PM_SKY130_FD_SC_LP__NOR2_0%B N_B_M1002_g N_B_M1000_g B B B B N_B_c_56_n
+ N_B_c_57_n PM_SKY130_FD_SC_LP__NOR2_0%B
x_PM_SKY130_FD_SC_LP__NOR2_0%VPWR N_VPWR_M1001_s N_VPWR_c_82_n N_VPWR_c_83_n
+ VPWR N_VPWR_c_84_n N_VPWR_c_81_n PM_SKY130_FD_SC_LP__NOR2_0%VPWR
x_PM_SKY130_FD_SC_LP__NOR2_0%Y N_Y_M1003_d N_Y_M1002_d Y Y Y Y Y Y N_Y_c_97_n Y
+ PM_SKY130_FD_SC_LP__NOR2_0%Y
x_PM_SKY130_FD_SC_LP__NOR2_0%VGND N_VGND_M1003_s N_VGND_M1000_d N_VGND_c_114_n
+ N_VGND_c_115_n N_VGND_c_116_n N_VGND_c_117_n VGND N_VGND_c_118_n
+ N_VGND_c_119_n PM_SKY130_FD_SC_LP__NOR2_0%VGND
cc_1 VNB N_A_c_29_n 0.0241976f $X=-0.19 $Y=-0.245 $X2=0.402 $Y2=1.353
cc_2 VNB N_A_M1001_g 0.00643653f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=2.735
cc_3 VNB N_A_c_31_n 0.0243907f $X=-0.19 $Y=-0.245 $X2=0.402 $Y2=1.55
cc_4 VNB A 0.0347357f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_5 VNB N_A_c_33_n 0.0243907f $X=-0.19 $Y=-0.245 $X2=0.37 $Y2=1.045
cc_6 VNB N_A_c_34_n 0.0212472f $X=-0.19 $Y=-0.245 $X2=0.402 $Y2=0.88
cc_7 VNB N_B_M1002_g 0.00508241f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=0.88
cc_8 VNB B 0.0337542f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=2.735
cc_9 VNB N_B_c_56_n 0.0838807f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_B_c_57_n 0.0198904f $X=-0.19 $Y=-0.245 $X2=0.402 $Y2=1.045
cc_11 VNB N_VPWR_c_81_n 0.0641695f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_12 VNB N_Y_c_97_n 0.00624061f $X=-0.19 $Y=-0.245 $X2=0.402 $Y2=0.88
cc_13 VNB N_VGND_c_114_n 0.0124811f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=2.735
cc_14 VNB N_VGND_c_115_n 0.0209751f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_VGND_c_116_n 0.0109361f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_16 VNB N_VGND_c_117_n 0.0231779f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_17 VNB N_VGND_c_118_n 0.0168361f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_VGND_c_119_n 0.111065f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.295
cc_19 VPB N_A_M1001_g 0.0625786f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=2.735
cc_20 VPB A 0.0302042f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_21 VPB N_B_M1002_g 0.0547621f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=0.88
cc_22 VPB B 0.034279f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=2.735
cc_23 VPB N_VPWR_c_82_n 0.011942f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=0.56
cc_24 VPB N_VPWR_c_83_n 0.0330547f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=1.55
cc_25 VPB N_VPWR_c_84_n 0.0262504f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_26 VPB N_VPWR_c_81_n 0.0523568f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_27 VPB N_Y_c_97_n 0.00562949f $X=-0.19 $Y=1.655 $X2=0.402 $Y2=0.88
cc_28 VPB Y 0.0376919f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_29 N_A_c_31_n N_B_M1002_g 0.0581393f $X=0.402 $Y=1.55 $X2=0 $Y2=0
cc_30 A N_B_c_56_n 9.50952e-19 $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_31 N_A_c_33_n N_B_c_56_n 0.0581393f $X=0.37 $Y=1.045 $X2=0 $Y2=0
cc_32 N_A_c_34_n N_B_c_57_n 0.0111277f $X=0.402 $Y=0.88 $X2=0 $Y2=0
cc_33 N_A_M1001_g N_VPWR_c_83_n 0.0110354f $X=0.525 $Y=2.735 $X2=0 $Y2=0
cc_34 A N_VPWR_c_83_n 0.0288227f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_35 N_A_M1001_g N_VPWR_c_84_n 0.00525707f $X=0.525 $Y=2.735 $X2=0 $Y2=0
cc_36 N_A_M1001_g N_VPWR_c_81_n 0.00933422f $X=0.525 $Y=2.735 $X2=0 $Y2=0
cc_37 A N_Y_c_97_n 0.108313f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_38 N_A_c_34_n N_Y_c_97_n 0.00991295f $X=0.402 $Y=0.88 $X2=0 $Y2=0
cc_39 N_A_c_29_n Y 0.00991295f $X=0.402 $Y=1.353 $X2=0 $Y2=0
cc_40 A N_VGND_c_115_n 0.0250475f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_41 N_A_c_33_n N_VGND_c_115_n 0.00156152f $X=0.37 $Y=1.045 $X2=0 $Y2=0
cc_42 N_A_c_34_n N_VGND_c_115_n 0.00782401f $X=0.402 $Y=0.88 $X2=0 $Y2=0
cc_43 N_A_c_34_n N_VGND_c_118_n 0.00460631f $X=0.402 $Y=0.88 $X2=0 $Y2=0
cc_44 A N_VGND_c_119_n 0.00348537f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_45 N_A_c_34_n N_VGND_c_119_n 0.00893712f $X=0.402 $Y=0.88 $X2=0 $Y2=0
cc_46 N_B_M1002_g N_VPWR_c_83_n 0.00131201f $X=0.915 $Y=2.735 $X2=0 $Y2=0
cc_47 N_B_M1002_g N_VPWR_c_84_n 0.00331858f $X=0.915 $Y=2.735 $X2=0 $Y2=0
cc_48 N_B_M1002_g N_VPWR_c_81_n 0.00567338f $X=0.915 $Y=2.735 $X2=0 $Y2=0
cc_49 N_B_M1002_g N_Y_c_97_n 0.0222176f $X=0.915 $Y=2.735 $X2=0 $Y2=0
cc_50 B N_Y_c_97_n 0.10413f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_51 N_B_c_56_n N_Y_c_97_n 0.0182901f $X=1.17 $Y=1.045 $X2=0 $Y2=0
cc_52 N_B_c_57_n N_Y_c_97_n 0.0112028f $X=1.087 $Y=0.88 $X2=0 $Y2=0
cc_53 N_B_M1002_g Y 0.0222477f $X=0.915 $Y=2.735 $X2=0 $Y2=0
cc_54 B Y 0.0223f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_55 N_B_c_57_n N_VGND_c_115_n 4.27056e-19 $X=1.087 $Y=0.88 $X2=0 $Y2=0
cc_56 B N_VGND_c_117_n 0.0235994f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_57 N_B_c_56_n N_VGND_c_117_n 0.00186616f $X=1.17 $Y=1.045 $X2=0 $Y2=0
cc_58 N_B_c_57_n N_VGND_c_117_n 0.00371692f $X=1.087 $Y=0.88 $X2=0 $Y2=0
cc_59 N_B_c_57_n N_VGND_c_118_n 0.00473473f $X=1.087 $Y=0.88 $X2=0 $Y2=0
cc_60 B N_VGND_c_119_n 0.0018004f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_61 N_B_c_56_n N_VGND_c_119_n 6.42459e-19 $X=1.17 $Y=1.045 $X2=0 $Y2=0
cc_62 N_B_c_57_n N_VGND_c_119_n 0.00937348f $X=1.087 $Y=0.88 $X2=0 $Y2=0
cc_63 N_VPWR_c_83_n Y 0.0270315f $X=0.31 $Y=2.56 $X2=0 $Y2=0
cc_64 N_VPWR_c_84_n Y 0.0473596f $X=1.2 $Y=3.33 $X2=0 $Y2=0
cc_65 N_VPWR_c_81_n Y 0.025284f $X=1.2 $Y=3.33 $X2=0 $Y2=0
cc_66 N_Y_c_97_n N_VGND_c_118_n 0.00821198f $X=0.74 $Y=0.55 $X2=0 $Y2=0
cc_67 N_Y_c_97_n N_VGND_c_119_n 0.00929282f $X=0.74 $Y=0.55 $X2=0 $Y2=0
