* File: sky130_fd_sc_lp__dlclkp_2.spice
* Created: Fri Aug 28 10:25:05 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__dlclkp_2.pex.spice"
.subckt sky130_fd_sc_lp__dlclkp_2  VNB VPB GATE CLK VPWR GCLK VGND
* 
* VGND	VGND
* GCLK	GCLK
* VPWR	VPWR
* CLK	CLK
* GATE	GATE
* VPB	VPB
* VNB	VNB
MM1005 N_VGND_M1005_d N_A_78_269#_M1005_g N_A_33_47#_M1005_s VNB NSHORT L=0.15
+ W=0.84 AD=0.22485 AS=0.2394 PD=1.84 PS=2.25 NRD=0 NRS=2.856 M=1 R=5.6
+ SA=75000.2 SB=75001.4 A=0.126 P=1.98 MULT=1
MM1020 A_258_81# N_GATE_M1020_g N_VGND_M1005_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.112425 PD=0.63 PS=0.92 NRD=14.28 NRS=75.708 M=1 R=2.8
+ SA=75000.9 SB=75002 A=0.063 P=1.14 MULT=1
MM1015 N_A_78_269#_M1015_d N_A_300_55#_M1015_g A_258_81# VNB NSHORT L=0.15
+ W=0.42 AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.3
+ SB=75001.6 A=0.063 P=1.14 MULT=1
MM1021 A_416_81# N_A_284_367#_M1021_g N_A_78_269#_M1015_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0672 AS=0.0588 PD=0.74 PS=0.7 NRD=30 NRS=0 M=1 R=2.8 SA=75001.7
+ SB=75001.2 A=0.063 P=1.14 MULT=1
MM1013 N_VGND_M1013_d N_A_33_47#_M1013_g A_416_81# VNB NSHORT L=0.15 W=0.42
+ AD=0.08295 AS=0.0672 PD=0.815 PS=0.74 NRD=27.132 NRS=30 M=1 R=2.8 SA=75002.2
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1019 N_A_284_367#_M1019_d N_A_300_55#_M1019_g N_VGND_M1013_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1113 AS=0.08295 PD=1.37 PS=0.815 NRD=0 NRS=5.712 M=1 R=2.8
+ SA=75002.7 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1007 N_VGND_M1007_d N_CLK_M1007_g N_A_300_55#_M1007_s VNB NSHORT L=0.15 W=0.42
+ AD=0.1766 AS=0.168 PD=1.425 PS=1.64 NRD=104.412 NRS=32.856 M=1 R=2.8
+ SA=75000.3 SB=75001.2 A=0.063 P=1.14 MULT=1
MM1006 A_1002_133# N_CLK_M1006_g N_VGND_M1007_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1766 PD=0.63 PS=1.425 NRD=14.28 NRS=104.412 M=1 R=2.8
+ SA=75000.9 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1002 N_A_1039_367#_M1002_d N_A_33_47#_M1002_g A_1002_133# VNB NSHORT L=0.15
+ W=0.42 AD=0.1113 AS=0.0441 PD=1.37 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8
+ SA=75001.3 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1003 N_VGND_M1003_d N_A_1039_367#_M1003_g N_GCLK_M1003_s VNB NSHORT L=0.15
+ W=0.84 AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1017 N_VGND_M1017_d N_A_1039_367#_M1017_g N_GCLK_M1003_s VNB NSHORT L=0.15
+ W=0.84 AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1009 N_VPWR_M1009_d N_A_78_269#_M1009_g N_A_33_47#_M1009_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.369943 AS=0.3339 PD=2.42716 PS=3.05 NRD=13.2778 NRS=0 M=1 R=8.4
+ SA=75000.2 SB=75001.2 A=0.189 P=2.82 MULT=1
MM1011 A_242_465# N_GATE_M1011_g N_VPWR_M1009_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0672 AS=0.187907 PD=0.85 PS=1.23284 NRD=15.3857 NRS=73.4416 M=1 R=4.26667
+ SA=75000.8 SB=75001.4 A=0.096 P=1.58 MULT=1
MM1004 N_A_78_269#_M1004_d N_A_284_367#_M1004_g A_242_465# VPB PHIGHVT L=0.15
+ W=0.64 AD=0.134098 AS=0.0672 PD=1.24377 PS=0.85 NRD=0 NRS=15.3857 M=1
+ R=4.26667 SA=75001.2 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1012 A_422_465# N_A_300_55#_M1012_g N_A_78_269#_M1004_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0441 AS=0.0880019 PD=0.63 PS=0.816226 NRD=23.443 NRS=51.5943 M=1
+ R=2.8 SA=75001.7 SB=75001 A=0.063 P=1.14 MULT=1
MM1014 N_VPWR_M1014_d N_A_33_47#_M1014_g A_422_465# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.146029 AS=0.0441 PD=1.12925 PS=0.63 NRD=56.2829 NRS=23.443 M=1 R=2.8
+ SA=75002.1 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1001 N_A_284_367#_M1001_d N_A_300_55#_M1001_g N_VPWR_M1014_d VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.1824 AS=0.222521 PD=1.85 PS=1.72075 NRD=0 NRS=90.0881 M=1
+ R=4.26667 SA=75001.3 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1008 N_VPWR_M1008_d N_CLK_M1008_g N_A_300_55#_M1008_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.20315 AS=0.3227 PD=1.51 PS=2.54 NRD=80.77 NRS=138.274 M=1
+ R=4.26667 SA=75000.3 SB=75002.3 A=0.096 P=1.58 MULT=1
MM1000 N_A_1039_367#_M1000_d N_CLK_M1000_g N_VPWR_M1008_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.12 AS=0.20315 PD=1.015 PS=1.51 NRD=15.3857 NRS=80.77 M=1 R=4.26667
+ SA=75000.9 SB=75001.7 A=0.096 P=1.58 MULT=1
MM1016 N_VPWR_M1016_d N_A_33_47#_M1016_g N_A_1039_367#_M1000_d VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.152354 AS=0.12 PD=1.152 PS=1.015 NRD=95.4071 NRS=3.5854 M=1
+ R=4.26667 SA=75001.4 SB=75001.2 A=0.096 P=1.58 MULT=1
MM1010 N_VPWR_M1016_d N_A_1039_367#_M1010_g N_GCLK_M1010_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.299946 AS=0.1764 PD=2.268 PS=1.54 NRD=4.6886 NRS=0 M=1 R=8.4
+ SA=75001.1 SB=75000.6 A=0.189 P=2.82 MULT=1
MM1018 N_VPWR_M1018_d N_A_1039_367#_M1018_g N_GCLK_M1010_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.6
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX22_noxref VNB VPB NWDIODE A=14.3299 P=19.35
c_81 VNB 0 1.79399e-19 $X=0 $Y=0
*
.include "sky130_fd_sc_lp__dlclkp_2.pxi.spice"
*
.ends
*
*
