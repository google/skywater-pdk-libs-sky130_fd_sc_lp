# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__isobufsrc_2
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__isobufsrc_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.360000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.600000 1.185000 0.885000 1.515000 ;
    END
  END A
  PIN SLEEP
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.055000 1.075000 2.815000 1.245000 ;
        RECT 1.055000 1.245000 1.775000 1.435000 ;
        RECT 2.555000 1.245000 2.815000 1.515000 ;
    END
  END SLEEP
  PIN X
    ANTENNADIFFAREA  0.823200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.435000 0.255000 1.695000 0.735000 ;
        RECT 1.435000 0.735000 3.275000 0.905000 ;
        RECT 1.820000 2.025000 3.275000 2.195000 ;
        RECT 1.820000 2.195000 2.150000 2.715000 ;
        RECT 2.365000 0.255000 2.555000 0.735000 ;
        RECT 2.985000 0.905000 3.275000 2.025000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.360000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.360000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.360000 0.085000 ;
      RECT 0.000000  3.245000 3.360000 3.415000 ;
      RECT 0.160000  0.700000 0.430000 1.685000 ;
      RECT 0.160000  1.685000 2.275000 1.855000 ;
      RECT 0.160000  1.855000 0.695000 2.210000 ;
      RECT 0.620000  0.085000 1.265000 0.885000 ;
      RECT 0.620000  0.885000 0.895000 1.015000 ;
      RECT 0.865000  2.025000 1.250000 3.245000 ;
      RECT 1.420000  2.025000 1.650000 2.895000 ;
      RECT 1.420000  2.895000 2.510000 3.075000 ;
      RECT 1.865000  0.085000 2.195000 0.565000 ;
      RECT 1.945000  1.415000 2.275000 1.685000 ;
      RECT 2.320000  2.365000 2.510000 2.895000 ;
      RECT 2.680000  2.365000 3.010000 3.245000 ;
      RECT 2.725000  0.085000 3.055000 0.565000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
  END
END sky130_fd_sc_lp__isobufsrc_2
