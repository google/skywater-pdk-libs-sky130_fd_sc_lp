* File: sky130_fd_sc_lp__a32oi_m.pex.spice
* Created: Wed Sep  2 09:28:41 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A32OI_M%B2 2 3 4 7 11 15 18 20 21 22 23 24 31
c39 11 0 7.48172e-20 $X=0.685 $Y=0.445
c40 7 0 1.7865e-19 $X=0.62 $Y=2.71
c41 3 0 1.66284e-19 $X=0.61 $Y=0.915
r42 23 24 20.5182 $w=1.98e-07 $l=3.7e-07 $layer=LI1_cond $X=0.255 $Y=2.035
+ $X2=0.255 $Y2=2.405
r43 22 23 20.5182 $w=1.98e-07 $l=3.7e-07 $layer=LI1_cond $X=0.255 $Y=1.665
+ $X2=0.255 $Y2=2.035
r44 21 22 20.5182 $w=1.98e-07 $l=3.7e-07 $layer=LI1_cond $X=0.255 $Y=1.295
+ $X2=0.255 $Y2=1.665
r45 20 21 20.5182 $w=1.98e-07 $l=3.7e-07 $layer=LI1_cond $X=0.255 $Y=0.925
+ $X2=0.255 $Y2=1.295
r46 20 31 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.27
+ $Y=1.005 $X2=0.27 $Y2=1.005
r47 16 18 133.319 $w=1.5e-07 $l=2.6e-07 $layer=POLY_cond $X=0.36 $Y=2.215
+ $X2=0.62 $Y2=2.215
r48 14 31 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.27 $Y=1.345
+ $X2=0.27 $Y2=1.005
r49 14 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.27 $Y=1.345
+ $X2=0.27 $Y2=1.51
r50 13 31 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=0.27 $Y=0.99
+ $X2=0.27 $Y2=1.005
r51 9 11 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.685 $Y=0.84
+ $X2=0.685 $Y2=0.445
r52 5 18 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.62 $Y=2.29 $X2=0.62
+ $Y2=2.215
r53 5 7 215.362 $w=1.5e-07 $l=4.2e-07 $layer=POLY_cond $X=0.62 $Y=2.29 $X2=0.62
+ $Y2=2.71
r54 4 13 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=0.435 $Y=0.915
+ $X2=0.27 $Y2=0.99
r55 3 9 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.61 $Y=0.915
+ $X2=0.685 $Y2=0.84
r56 3 4 89.734 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=0.61 $Y=0.915
+ $X2=0.435 $Y2=0.915
r57 2 16 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.36 $Y=2.14 $X2=0.36
+ $Y2=2.215
r58 2 15 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=0.36 $Y=2.14 $X2=0.36
+ $Y2=1.51
.ends

.subckt PM_SKY130_FD_SC_LP__A32OI_M%B1 3 7 11 12 13 14 15 16 22
c47 13 0 1.66284e-19 $X=1.2 $Y=0.925
c48 7 0 1.87176e-19 $X=1.05 $Y=2.71
c49 3 0 1.13091e-20 $X=1.045 $Y=0.445
r50 22 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.07
+ $Y=1.395 $X2=1.07 $Y2=1.395
r51 15 16 14.2135 $w=2.98e-07 $l=3.7e-07 $layer=LI1_cond $X=1.135 $Y=1.665
+ $X2=1.135 $Y2=2.035
r52 15 23 10.372 $w=2.98e-07 $l=2.7e-07 $layer=LI1_cond $X=1.135 $Y=1.665
+ $X2=1.135 $Y2=1.395
r53 14 23 3.84148 $w=2.98e-07 $l=1e-07 $layer=LI1_cond $X=1.135 $Y=1.295
+ $X2=1.135 $Y2=1.395
r54 13 14 14.2135 $w=2.98e-07 $l=3.7e-07 $layer=LI1_cond $X=1.135 $Y=0.925
+ $X2=1.135 $Y2=1.295
r55 11 22 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.07 $Y=1.735
+ $X2=1.07 $Y2=1.395
r56 11 12 38.6168 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.07 $Y=1.735
+ $X2=1.07 $Y2=1.9
r57 10 22 38.9318 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.07 $Y=1.23
+ $X2=1.07 $Y2=1.395
r58 7 12 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=1.05 $Y=2.71 $X2=1.05
+ $Y2=1.9
r59 3 10 402.521 $w=1.5e-07 $l=7.85e-07 $layer=POLY_cond $X=1.045 $Y=0.445
+ $X2=1.045 $Y2=1.23
.ends

.subckt PM_SKY130_FD_SC_LP__A32OI_M%A1 3 6 9 10 11 12 13 14 15 16 23
r49 15 16 17.7668 $w=2.38e-07 $l=3.7e-07 $layer=LI1_cond $X=1.645 $Y=1.665
+ $X2=1.645 $Y2=2.035
r50 14 15 17.7668 $w=2.38e-07 $l=3.7e-07 $layer=LI1_cond $X=1.645 $Y=1.295
+ $X2=1.645 $Y2=1.665
r51 13 14 17.7668 $w=2.38e-07 $l=3.7e-07 $layer=LI1_cond $X=1.645 $Y=0.925
+ $X2=1.645 $Y2=1.295
r52 13 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.61
+ $Y=0.93 $X2=1.61 $Y2=0.93
r53 12 13 17.7668 $w=2.38e-07 $l=3.7e-07 $layer=LI1_cond $X=1.645 $Y=0.555
+ $X2=1.645 $Y2=0.925
r54 10 23 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.61 $Y=1.27
+ $X2=1.61 $Y2=0.93
r55 10 11 40.8701 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.61 $Y=1.27
+ $X2=1.61 $Y2=1.435
r56 9 23 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.61 $Y=0.765
+ $X2=1.61 $Y2=0.93
r57 6 11 653.777 $w=1.5e-07 $l=1.275e-06 $layer=POLY_cond $X=1.56 $Y=2.71
+ $X2=1.56 $Y2=1.435
r58 3 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.52 $Y=0.445 $X2=1.52
+ $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_LP__A32OI_M%A2 3 6 9 11 12 13 14 15 16 23
c49 9 0 1.9934e-19 $X=2.07 $Y=2.71
r50 23 25 46.3065 $w=3.4e-07 $l=1.65e-07 $layer=POLY_cond $X=2.155 $Y=1.32
+ $X2=2.155 $Y2=1.155
r51 15 16 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=2.16 $Y=1.665
+ $X2=2.16 $Y2=2.035
r52 14 15 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=2.16 $Y=1.295
+ $X2=2.16 $Y2=1.665
r53 14 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.16
+ $Y=1.32 $X2=2.16 $Y2=1.32
r54 13 14 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=2.16 $Y=0.925
+ $X2=2.16 $Y2=1.295
r55 12 13 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=2.16 $Y=0.555
+ $X2=2.16 $Y2=0.925
r56 9 11 453.798 $w=1.5e-07 $l=8.85e-07 $layer=POLY_cond $X=2.07 $Y=2.71
+ $X2=2.07 $Y2=1.825
r57 6 11 45.4119 $w=3.4e-07 $l=1.7e-07 $layer=POLY_cond $X=2.155 $Y=1.655
+ $X2=2.155 $Y2=1.825
r58 5 23 0.848592 $w=3.4e-07 $l=5e-09 $layer=POLY_cond $X=2.155 $Y=1.325
+ $X2=2.155 $Y2=1.32
r59 5 6 56.007 $w=3.4e-07 $l=3.3e-07 $layer=POLY_cond $X=2.155 $Y=1.325
+ $X2=2.155 $Y2=1.655
r60 3 25 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=2.06 $Y=0.445
+ $X2=2.06 $Y2=1.155
.ends

.subckt PM_SKY130_FD_SC_LP__A32OI_M%A3 1 3 6 12 15 16 18 19 20 21 22 23 30
c39 6 0 1.9934e-19 $X=2.5 $Y=2.71
r40 30 31 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.73
+ $Y=1.71 $X2=2.73 $Y2=1.71
r41 22 23 16.4002 $w=2.58e-07 $l=3.7e-07 $layer=LI1_cond $X=2.685 $Y=2.035
+ $X2=2.685 $Y2=2.405
r42 22 31 14.4055 $w=2.58e-07 $l=3.25e-07 $layer=LI1_cond $X=2.685 $Y=2.035
+ $X2=2.685 $Y2=1.71
r43 21 31 1.99461 $w=2.58e-07 $l=4.5e-08 $layer=LI1_cond $X=2.685 $Y=1.665
+ $X2=2.685 $Y2=1.71
r44 20 21 16.4002 $w=2.58e-07 $l=3.7e-07 $layer=LI1_cond $X=2.685 $Y=1.295
+ $X2=2.685 $Y2=1.665
r45 19 20 16.4002 $w=2.58e-07 $l=3.7e-07 $layer=LI1_cond $X=2.685 $Y=0.925
+ $X2=2.685 $Y2=1.295
r46 18 30 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.73 $Y=1.545
+ $X2=2.73 $Y2=1.71
r47 15 30 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=2.73 $Y=2.065
+ $X2=2.73 $Y2=1.71
r48 15 16 43.5886 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=2.66 $Y=2.065
+ $X2=2.66 $Y2=2.215
r49 10 12 112.809 $w=1.5e-07 $l=2.2e-07 $layer=POLY_cond $X=2.42 $Y=0.84
+ $X2=2.64 $Y2=0.84
r50 8 12 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.64 $Y=0.915
+ $X2=2.64 $Y2=0.84
r51 8 18 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=2.64 $Y=0.915
+ $X2=2.64 $Y2=1.545
r52 6 16 253.819 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=2.5 $Y=2.71 $X2=2.5
+ $Y2=2.215
r53 1 10 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.42 $Y=0.765
+ $X2=2.42 $Y2=0.84
r54 1 3 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.42 $Y=0.765 $X2=2.42
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__A32OI_M%A_40_500# 1 2 3 10 15 16 17 20 23
c36 20 0 5.58598e-19 $X=2.285 $Y=2.645
c37 15 0 1.73472e-19 $X=1.285 $Y=2.645
r38 23 25 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=0.325 $Y=2.775
+ $X2=0.325 $Y2=2.975
r39 18 20 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=2.285 $Y=2.49
+ $X2=2.285 $Y2=2.645
r40 16 18 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.2 $Y=2.405
+ $X2=2.285 $Y2=2.49
r41 16 17 52.8449 $w=1.68e-07 $l=8.1e-07 $layer=LI1_cond $X=2.2 $Y=2.405
+ $X2=1.39 $Y2=2.405
r42 13 15 12.9394 $w=2.08e-07 $l=2.45e-07 $layer=LI1_cond $X=1.285 $Y=2.89
+ $X2=1.285 $Y2=2.645
r43 12 17 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=1.285 $Y=2.49
+ $X2=1.39 $Y2=2.405
r44 12 15 8.18615 $w=2.08e-07 $l=1.55e-07 $layer=LI1_cond $X=1.285 $Y=2.49
+ $X2=1.285 $Y2=2.645
r45 11 25 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.49 $Y=2.975
+ $X2=0.325 $Y2=2.975
r46 10 13 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=1.18 $Y=2.975
+ $X2=1.285 $Y2=2.89
r47 10 11 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.18 $Y=2.975
+ $X2=0.49 $Y2=2.975
r48 3 20 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.145
+ $Y=2.5 $X2=2.285 $Y2=2.645
r49 2 15 600 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_PDIFF $count=1 $X=1.125
+ $Y=2.5 $X2=1.285 $Y2=2.645
r50 1 23 600 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_PDIFF $count=1 $X=0.2
+ $Y=2.5 $X2=0.325 $Y2=2.775
.ends

.subckt PM_SKY130_FD_SC_LP__A32OI_M%Y 1 2 7 8 10 14 18
c40 18 0 1.7865e-19 $X=0.72 $Y=0.925
c41 14 0 8.61263e-20 $X=1.26 $Y=0.495
r42 14 16 4.66986 $w=1.88e-07 $l=8e-08 $layer=LI1_cond $X=1.25 $Y=0.495 $X2=1.25
+ $Y2=0.575
r43 10 18 89.7059 $w=1.68e-07 $l=1.375e-06 $layer=LI1_cond $X=0.72 $Y=2.3
+ $X2=0.72 $Y2=0.925
r44 10 12 14.6492 $w=3.44e-07 $l=3.70338e-07 $layer=LI1_cond $X=0.72 $Y=2.3
+ $X2=0.817 $Y2=2.625
r45 9 18 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.72 $Y=0.66
+ $X2=0.72 $Y2=0.925
r46 8 9 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.805 $Y=0.575
+ $X2=0.72 $Y2=0.66
r47 7 16 1.386 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.155 $Y=0.575 $X2=1.25
+ $Y2=0.575
r48 7 8 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=1.155 $Y=0.575
+ $X2=0.805 $Y2=0.575
r49 2 12 600 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=0.695
+ $Y=2.5 $X2=0.835 $Y2=2.625
r50 1 14 182 $w=1.7e-07 $l=3.2249e-07 $layer=licon1_NDIFF $count=1 $X=1.12
+ $Y=0.235 $X2=1.26 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__A32OI_M%VPWR 1 2 9 13 15 17 22 29 30 33 36
c35 9 0 1.87176e-19 $X=1.775 $Y=2.775
r36 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r37 30 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.64 $Y2=3.33
r38 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r39 27 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.88 $Y=3.33
+ $X2=2.715 $Y2=3.33
r40 27 29 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=2.88 $Y=3.33
+ $X2=3.12 $Y2=3.33
r41 26 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r42 25 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r43 23 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.94 $Y=3.33
+ $X2=1.775 $Y2=3.33
r44 23 25 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=1.94 $Y=3.33
+ $X2=2.16 $Y2=3.33
r45 22 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.55 $Y=3.33
+ $X2=2.715 $Y2=3.33
r46 22 25 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=2.55 $Y=3.33
+ $X2=2.16 $Y2=3.33
r47 19 20 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r48 17 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.61 $Y=3.33
+ $X2=1.775 $Y2=3.33
r49 17 19 89.3797 $w=1.68e-07 $l=1.37e-06 $layer=LI1_cond $X=1.61 $Y=3.33
+ $X2=0.24 $Y2=3.33
r50 15 26 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r51 15 20 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.24 $Y2=3.33
r52 15 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r53 11 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.715 $Y=3.245
+ $X2=2.715 $Y2=3.33
r54 11 13 16.4136 $w=3.28e-07 $l=4.7e-07 $layer=LI1_cond $X=2.715 $Y=3.245
+ $X2=2.715 $Y2=2.775
r55 7 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.775 $Y=3.245
+ $X2=1.775 $Y2=3.33
r56 7 9 16.4136 $w=3.28e-07 $l=4.7e-07 $layer=LI1_cond $X=1.775 $Y=3.245
+ $X2=1.775 $Y2=2.775
r57 2 13 600 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=1 $X=2.575
+ $Y=2.5 $X2=2.715 $Y2=2.775
r58 1 9 600 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=1 $X=1.635
+ $Y=2.5 $X2=1.775 $Y2=2.775
.ends

.subckt PM_SKY130_FD_SC_LP__A32OI_M%VGND 1 2 7 9 13 15 17 27 28 34
r45 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r46 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r47 28 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.64
+ $Y2=0
r48 27 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r49 25 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.8 $Y=0 $X2=2.635
+ $Y2=0
r50 25 27 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=2.8 $Y=0 $X2=3.12
+ $Y2=0
r51 24 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r52 23 24 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r53 21 32 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r54 20 23 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=0.72 $Y=0 $X2=2.16
+ $Y2=0
r55 20 21 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r56 18 31 4.70928 $w=1.7e-07 $l=2.28e-07 $layer=LI1_cond $X=0.455 $Y=0 $X2=0.227
+ $Y2=0
r57 18 20 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.455 $Y=0 $X2=0.72
+ $Y2=0
r58 17 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.47 $Y=0 $X2=2.635
+ $Y2=0
r59 17 23 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=2.47 $Y=0 $X2=2.16
+ $Y2=0
r60 15 24 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r61 15 21 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=0.72
+ $Y2=0
r62 11 34 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.635 $Y=0.085
+ $X2=2.635 $Y2=0
r63 11 13 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.635 $Y=0.085
+ $X2=2.635 $Y2=0.38
r64 7 31 3.0569 $w=3.3e-07 $l=1.12161e-07 $layer=LI1_cond $X=0.29 $Y=0.085
+ $X2=0.227 $Y2=0
r65 7 9 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.29 $Y=0.085
+ $X2=0.29 $Y2=0.38
r66 2 13 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=2.495
+ $Y=0.235 $X2=2.635 $Y2=0.38
r67 1 9 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.165
+ $Y=0.235 $X2=0.29 $Y2=0.38
.ends

