# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_lp__nor4b_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.280000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.870000 1.210000 4.645000 1.445000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.400000 1.345000 3.660000 1.615000 ;
        RECT 3.400000 1.615000 5.195000 1.785000 ;
        RECT 4.815000 1.185000 5.195000 1.615000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.865000 1.085000 2.880000 1.255000 ;
        RECT 0.865000 1.255000 1.065000 1.515000 ;
        RECT 2.490000 1.255000 2.880000 1.515000 ;
    END
  END C
  PIN D_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.185000 0.355000 1.515000 ;
    END
  END D_N
  PIN Y
    ANTENNADIFFAREA  1.293600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.535000 0.255000 1.795000 0.745000 ;
        RECT 1.535000 0.745000 3.825000 0.870000 ;
        RECT 1.535000 0.870000 4.685000 0.915000 ;
        RECT 1.585000 1.805000 3.230000 1.975000 ;
        RECT 1.585000 1.975000 2.735000 2.145000 ;
        RECT 2.465000 0.255000 2.725000 0.745000 ;
        RECT 3.060000 0.915000 4.685000 1.040000 ;
        RECT 3.060000 1.040000 3.700000 1.175000 ;
        RECT 3.060000 1.175000 3.230000 1.805000 ;
        RECT 3.565000 0.255000 3.825000 0.745000 ;
        RECT 4.495000 0.265000 4.685000 0.870000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 5.280000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.500000 0.500000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.800000 0.500000 3.300000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 5.280000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.280000 0.085000 ;
      RECT 0.000000  3.245000 5.280000 3.415000 ;
      RECT 0.095000  1.695000 1.415000 1.865000 ;
      RECT 0.095000  1.865000 0.355000 3.050000 ;
      RECT 0.150000  0.795000 0.695000 1.005000 ;
      RECT 0.525000  1.005000 0.695000 1.695000 ;
      RECT 0.525000  2.720000 0.855000 3.245000 ;
      RECT 0.865000  0.085000 1.365000 0.915000 ;
      RECT 1.105000  2.035000 1.415000 2.315000 ;
      RECT 1.105000  2.315000 3.235000 2.485000 ;
      RECT 1.105000  2.485000 1.410000 3.075000 ;
      RECT 1.245000  1.425000 2.320000 1.635000 ;
      RECT 1.245000  1.635000 1.415000 1.695000 ;
      RECT 1.580000  2.655000 2.735000 3.010000 ;
      RECT 1.965000  0.085000 2.295000 0.575000 ;
      RECT 2.905000  2.145000 5.185000 2.285000 ;
      RECT 2.905000  2.285000 3.815000 2.315000 ;
      RECT 2.905000  2.485000 3.235000 3.075000 ;
      RECT 2.985000  0.085000 3.315000 0.575000 ;
      RECT 3.440000  2.485000 3.770000 2.835000 ;
      RECT 3.440000  2.835000 4.755000 3.075000 ;
      RECT 3.645000  2.005000 5.185000 2.145000 ;
      RECT 3.995000  0.085000 4.325000 0.700000 ;
      RECT 3.995000  2.455000 5.195000 2.665000 ;
      RECT 4.855000  0.085000 5.185000 1.015000 ;
      RECT 4.935000  2.665000 5.195000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
  END
END sky130_fd_sc_lp__nor4b_2
END LIBRARY
