* File: sky130_fd_sc_lp__a41o_2.spice
* Created: Fri Aug 28 10:02:38 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__a41o_2.pex.spice"
.subckt sky130_fd_sc_lp__a41o_2  VNB VPB B1 A4 A3 A2 A1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A1	A1
* A2	A2
* A3	A3
* A4	A4
* B1	B1
* VPB	VPB
* VNB	VNB
MM1008 N_X_M1008_d N_A_90_53#_M1008_g N_VGND_M1008_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1011 N_X_M1008_d N_A_90_53#_M1011_g N_VGND_M1011_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1002 N_VGND_M1002_d N_B1_M1002_g N_A_90_53#_M1002_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1638 AS=0.2226 PD=1.23 PS=2.21 NRD=7.848 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75002.2 A=0.126 P=1.98 MULT=1
MM1006 A_561_49# N_A4_M1006_g N_VGND_M1002_d VNB NSHORT L=0.15 W=0.84 AD=0.0882
+ AS=0.1638 PD=1.05 PS=1.23 NRD=7.14 NRS=7.848 M=1 R=5.6 SA=75000.7 SB=75001.6
+ A=0.126 P=1.98 MULT=1
MM1007 A_633_49# N_A3_M1007_g A_561_49# VNB NSHORT L=0.15 W=0.84 AD=0.1638
+ AS=0.0882 PD=1.23 PS=1.05 NRD=19.992 NRS=7.14 M=1 R=5.6 SA=75001.1 SB=75001.3
+ A=0.126 P=1.98 MULT=1
MM1009 A_741_49# N_A2_M1009_g A_633_49# VNB NSHORT L=0.15 W=0.84 AD=0.1638
+ AS=0.1638 PD=1.23 PS=1.23 NRD=19.992 NRS=19.992 M=1 R=5.6 SA=75001.6
+ SB=75000.7 A=0.126 P=1.98 MULT=1
MM1003 N_A_90_53#_M1003_d N_A1_M1003_g A_741_49# VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1638 PD=2.21 PS=1.23 NRD=0 NRS=19.992 M=1 R=5.6 SA=75002.2
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1004 N_VPWR_M1004_d N_A_90_53#_M1004_g N_X_M1004_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1013 N_VPWR_M1013_d N_A_90_53#_M1013_g N_X_M1004_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75000.2 A=0.189 P=2.82 MULT=1
MM1005 N_A_453_367#_M1005_d N_B1_M1005_g N_A_90_53#_M1005_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75002.2 A=0.189 P=2.82 MULT=1
MM1001 N_VPWR_M1001_d N_A4_M1001_g N_A_453_367#_M1005_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.2016 AS=0.1764 PD=1.58 PS=1.54 NRD=3.1126 NRS=0 M=1 R=8.4
+ SA=75000.6 SB=75001.7 A=0.189 P=2.82 MULT=1
MM1012 N_A_453_367#_M1012_d N_A3_M1012_g N_VPWR_M1001_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.315 AS=0.2016 PD=1.76 PS=1.58 NRD=18.7544 NRS=3.1126 M=1 R=8.4
+ SA=75001.1 SB=75001.3 A=0.189 P=2.82 MULT=1
MM1000 N_VPWR_M1000_d N_A2_M1000_g N_A_453_367#_M1012_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.315 PD=1.54 PS=1.76 NRD=0 NRS=15.6221 M=1 R=8.4
+ SA=75001.7 SB=75000.6 A=0.189 P=2.82 MULT=1
MM1010 N_A_453_367#_M1010_d N_A1_M1010_g N_VPWR_M1000_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.2
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX14_noxref VNB VPB NWDIODE A=9.6607 P=14.09
*
.include "sky130_fd_sc_lp__a41o_2.pxi.spice"
*
.ends
*
*
