* File: sky130_fd_sc_lp__nand4bb_2.pex.spice
* Created: Wed Sep  2 10:06:46 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__NAND4BB_2%B_N 3 7 9 10 11 12 13 17
r33 17 18 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.56
+ $Y=0.94 $X2=0.56 $Y2=0.94
r34 13 18 10.7662 $w=3.78e-07 $l=3.55e-07 $layer=LI1_cond $X=0.655 $Y=1.295
+ $X2=0.655 $Y2=0.94
r35 12 18 0.454912 $w=3.78e-07 $l=1.5e-08 $layer=LI1_cond $X=0.655 $Y=0.925
+ $X2=0.655 $Y2=0.94
r36 10 17 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.56 $Y=1.28
+ $X2=0.56 $Y2=0.94
r37 10 11 45.2978 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.56 $Y=1.28
+ $X2=0.56 $Y2=1.445
r38 9 17 40.8701 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.56 $Y=0.775
+ $X2=0.56 $Y2=0.94
r39 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.61 $Y=0.455 $X2=0.61
+ $Y2=0.775
r40 3 11 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=0.475 $Y=2.075
+ $X2=0.475 $Y2=1.445
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4BB_2%A_N 3 6 9 10 11 12 13 17
r38 12 13 14.7036 $w=2.88e-07 $l=3.7e-07 $layer=LI1_cond $X=1.16 $Y=0.925
+ $X2=1.16 $Y2=1.295
r39 12 17 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.13
+ $Y=0.94 $X2=1.13 $Y2=0.94
r40 10 17 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.13 $Y=1.28
+ $X2=1.13 $Y2=0.94
r41 10 11 40.425 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.13 $Y=1.28
+ $X2=1.13 $Y2=1.445
r42 9 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.13 $Y=0.775
+ $X2=1.13 $Y2=0.94
r43 6 11 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=1.175 $Y=2.075
+ $X2=1.175 $Y2=1.445
r44 3 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.04 $Y=0.455 $X2=1.04
+ $Y2=0.775
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4BB_2%A_223_49# 1 2 9 13 17 21 23 27 36 39 40 43
+ 45
c75 23 0 2.94344e-20 $X=2.05 $Y=1.49
c76 9 0 1.20189e-19 $X=2.125 $Y=0.655
r77 43 45 8.47192 $w=3.38e-07 $l=1.65e-07 $layer=LI1_cond $X=1.645 $Y=1.49
+ $X2=1.645 $Y2=1.325
r78 43 44 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.7
+ $Y=1.49 $X2=1.7 $Y2=1.49
r79 39 40 5.20176 $w=5.08e-07 $l=1.65e-07 $layer=LI1_cond $X=1.56 $Y=2.01
+ $X2=1.56 $Y2=1.845
r80 34 36 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=1.255 $Y=0.44
+ $X2=1.56 $Y2=0.44
r81 31 43 0.169477 $w=3.38e-07 $l=5e-09 $layer=LI1_cond $X=1.645 $Y=1.495
+ $X2=1.645 $Y2=1.49
r82 31 40 11.8634 $w=3.38e-07 $l=3.5e-07 $layer=LI1_cond $X=1.645 $Y=1.495
+ $X2=1.645 $Y2=1.845
r83 29 36 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.56 $Y=0.605
+ $X2=1.56 $Y2=0.44
r84 29 45 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=1.56 $Y=0.605
+ $X2=1.56 $Y2=1.325
r85 26 27 13.9889 $w=3.3e-07 $l=8e-08 $layer=POLY_cond $X=2.555 $Y=1.49
+ $X2=2.635 $Y2=1.49
r86 25 26 61.2015 $w=3.3e-07 $l=3.5e-07 $layer=POLY_cond $X=2.205 $Y=1.49
+ $X2=2.555 $Y2=1.49
r87 24 25 13.9889 $w=3.3e-07 $l=8e-08 $layer=POLY_cond $X=2.125 $Y=1.49
+ $X2=2.205 $Y2=1.49
r88 23 44 61.2015 $w=3.3e-07 $l=3.5e-07 $layer=POLY_cond $X=2.05 $Y=1.49 $X2=1.7
+ $Y2=1.49
r89 23 24 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=2.05 $Y=1.49
+ $X2=2.125 $Y2=1.49
r90 19 27 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.635 $Y=1.655
+ $X2=2.635 $Y2=1.49
r91 19 21 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=2.635 $Y=1.655
+ $X2=2.635 $Y2=2.465
r92 15 26 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.555 $Y=1.325
+ $X2=2.555 $Y2=1.49
r93 15 17 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=2.555 $Y=1.325
+ $X2=2.555 $Y2=0.655
r94 11 25 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.205 $Y=1.655
+ $X2=2.205 $Y2=1.49
r95 11 13 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=2.205 $Y=1.655
+ $X2=2.205 $Y2=2.465
r96 7 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.125 $Y=1.325
+ $X2=2.125 $Y2=1.49
r97 7 9 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=2.125 $Y=1.325
+ $X2=2.125 $Y2=0.655
r98 2 39 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.25
+ $Y=1.865 $X2=1.39 $Y2=2.01
r99 1 34 182 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_NDIFF $count=1 $X=1.115
+ $Y=0.245 $X2=1.255 $Y2=0.44
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4BB_2%A_27_373# 1 2 9 13 17 21 24 27 29 32 33 34
+ 36 37 39 45 47 52
c103 29 0 2.94344e-20 $X=0.965 $Y=1.71
c104 21 0 6.36774e-20 $X=3.495 $Y=2.465
c105 13 0 6.36774e-20 $X=3.065 $Y=2.465
r106 48 50 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=2.995 $Y=1.485
+ $X2=3.065 $Y2=1.485
r107 42 45 7.15912 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=0.19 $Y=0.44
+ $X2=0.395 $Y2=0.44
r108 40 52 71.6931 $w=3.3e-07 $l=4.1e-07 $layer=POLY_cond $X=3.085 $Y=1.485
+ $X2=3.495 $Y2=1.485
r109 40 50 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=3.085 $Y=1.485
+ $X2=3.065 $Y2=1.485
r110 39 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.085
+ $Y=1.485 $X2=3.085 $Y2=1.485
r111 37 39 52.8951 $w=1.93e-07 $l=9.3e-07 $layer=LI1_cond $X=2.155 $Y=1.472
+ $X2=3.085 $Y2=1.472
r112 35 37 6.85817 $w=1.95e-07 $l=1.33918e-07 $layer=LI1_cond $X=2.07 $Y=1.57
+ $X2=2.155 $Y2=1.472
r113 35 36 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=2.07 $Y=1.57
+ $X2=2.07 $Y2=2.345
r114 33 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.985 $Y=2.43
+ $X2=2.07 $Y2=2.345
r115 33 34 55.4545 $w=1.68e-07 $l=8.5e-07 $layer=LI1_cond $X=1.985 $Y=2.43
+ $X2=1.135 $Y2=2.43
r116 32 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.05 $Y=2.345
+ $X2=1.135 $Y2=2.43
r117 31 32 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=1.05 $Y=1.795
+ $X2=1.05 $Y2=2.345
r118 30 47 2.87242 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=0.39 $Y=1.71
+ $X2=0.237 $Y2=1.71
r119 29 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.965 $Y=1.71
+ $X2=1.05 $Y2=1.795
r120 29 30 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=0.965 $Y=1.71
+ $X2=0.39 $Y2=1.71
r121 25 47 3.6114 $w=2.57e-07 $l=8.5e-08 $layer=LI1_cond $X=0.237 $Y=1.795
+ $X2=0.237 $Y2=1.71
r122 25 27 10.5798 $w=3.03e-07 $l=2.8e-07 $layer=LI1_cond $X=0.237 $Y=1.795
+ $X2=0.237 $Y2=2.075
r123 24 47 3.6114 $w=2.57e-07 $l=1.05924e-07 $layer=LI1_cond $X=0.19 $Y=1.625
+ $X2=0.237 $Y2=1.71
r124 23 42 3.38185 $w=2.1e-07 $l=1.65e-07 $layer=LI1_cond $X=0.19 $Y=0.605
+ $X2=0.19 $Y2=0.44
r125 23 24 53.8701 $w=2.08e-07 $l=1.02e-06 $layer=LI1_cond $X=0.19 $Y=0.605
+ $X2=0.19 $Y2=1.625
r126 19 52 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.495 $Y=1.65
+ $X2=3.495 $Y2=1.485
r127 19 21 417.904 $w=1.5e-07 $l=8.15e-07 $layer=POLY_cond $X=3.495 $Y=1.65
+ $X2=3.495 $Y2=2.465
r128 15 52 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.495 $Y=1.32
+ $X2=3.495 $Y2=1.485
r129 15 17 340.989 $w=1.5e-07 $l=6.65e-07 $layer=POLY_cond $X=3.495 $Y=1.32
+ $X2=3.495 $Y2=0.655
r130 11 50 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.065 $Y=1.65
+ $X2=3.065 $Y2=1.485
r131 11 13 417.904 $w=1.5e-07 $l=8.15e-07 $layer=POLY_cond $X=3.065 $Y=1.65
+ $X2=3.065 $Y2=2.465
r132 7 48 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.995 $Y=1.32
+ $X2=2.995 $Y2=1.485
r133 7 9 340.989 $w=1.5e-07 $l=6.65e-07 $layer=POLY_cond $X=2.995 $Y=1.32
+ $X2=2.995 $Y2=0.655
r134 2 27 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.865 $X2=0.26 $Y2=2.075
r135 1 45 182 $w=1.7e-07 $l=2.498e-07 $layer=licon1_NDIFF $count=1 $X=0.27
+ $Y=0.245 $X2=0.395 $Y2=0.44
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4BB_2%C 3 7 9 11 12 13 14 16 17 18
c54 13 0 1.00365e-19 $X=4.525 $Y=1.26
r55 24 26 12.4529 $w=3.29e-07 $l=8.5e-08 $layer=POLY_cond $X=4.36 $Y=1.35
+ $X2=4.445 $Y2=1.35
r56 24 25 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.36
+ $Y=1.35 $X2=4.36 $Y2=1.35
r57 22 24 0.732523 $w=3.29e-07 $l=5e-09 $layer=POLY_cond $X=4.355 $Y=1.35
+ $X2=4.36 $Y2=1.35
r58 21 22 62.997 $w=3.29e-07 $l=4.3e-07 $layer=POLY_cond $X=3.925 $Y=1.35
+ $X2=4.355 $Y2=1.35
r59 18 25 10.2439 $w=2.23e-07 $l=2e-07 $layer=LI1_cond $X=4.56 $Y=1.322 $X2=4.36
+ $Y2=1.322
r60 17 25 14.3415 $w=2.23e-07 $l=2.8e-07 $layer=LI1_cond $X=4.08 $Y=1.322
+ $X2=4.36 $Y2=1.322
r61 14 16 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=4.875 $Y=1.185
+ $X2=4.875 $Y2=0.655
r62 13 26 26.1409 $w=3.29e-07 $l=1.23693e-07 $layer=POLY_cond $X=4.525 $Y=1.26
+ $X2=4.445 $Y2=1.35
r63 12 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.8 $Y=1.26
+ $X2=4.875 $Y2=1.185
r64 12 13 141.011 $w=1.5e-07 $l=2.75e-07 $layer=POLY_cond $X=4.8 $Y=1.26
+ $X2=4.525 $Y2=1.26
r65 9 26 21.1507 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.445 $Y=1.185
+ $X2=4.445 $Y2=1.35
r66 9 11 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=4.445 $Y=1.185
+ $X2=4.445 $Y2=0.655
r67 5 22 21.1507 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.355 $Y=1.515
+ $X2=4.355 $Y2=1.35
r68 5 7 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=4.355 $Y=1.515
+ $X2=4.355 $Y2=2.465
r69 1 21 21.1507 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.925 $Y=1.515
+ $X2=3.925 $Y2=1.35
r70 1 3 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=3.925 $Y=1.515
+ $X2=3.925 $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4BB_2%D 1 3 4 5 8 10 12 15 17 18 24
c46 8 0 1.00365e-19 $X=5.305 $Y=0.655
r47 24 26 6.5847 $w=3.66e-07 $l=5e-08 $layer=POLY_cond $X=5.685 $Y=1.535
+ $X2=5.735 $Y2=1.535
r48 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.685
+ $Y=1.51 $X2=5.685 $Y2=1.51
r49 22 24 11.8525 $w=3.66e-07 $l=9e-08 $layer=POLY_cond $X=5.595 $Y=1.535
+ $X2=5.685 $Y2=1.535
r50 21 22 38.1913 $w=3.66e-07 $l=2.9e-07 $layer=POLY_cond $X=5.305 $Y=1.535
+ $X2=5.595 $Y2=1.535
r51 18 25 11.1698 $w=3.23e-07 $l=3.15e-07 $layer=LI1_cond $X=6 $Y=1.587
+ $X2=5.685 $Y2=1.587
r52 17 25 5.85086 $w=3.23e-07 $l=1.65e-07 $layer=LI1_cond $X=5.52 $Y=1.587
+ $X2=5.685 $Y2=1.587
r53 13 26 23.7042 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=5.735 $Y=1.345
+ $X2=5.735 $Y2=1.535
r54 13 15 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=5.735 $Y=1.345
+ $X2=5.735 $Y2=0.655
r55 10 22 23.7042 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=5.595 $Y=1.725
+ $X2=5.595 $Y2=1.535
r56 10 12 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=5.595 $Y=1.725
+ $X2=5.595 $Y2=2.465
r57 6 21 23.7042 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=5.305 $Y=1.345
+ $X2=5.305 $Y2=1.535
r58 6 8 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=5.305 $Y=1.345
+ $X2=5.305 $Y2=0.655
r59 4 21 36.3615 $w=3.66e-07 $l=1.94165e-07 $layer=POLY_cond $X=5.16 $Y=1.65
+ $X2=5.305 $Y2=1.535
r60 4 5 153.83 $w=1.5e-07 $l=3e-07 $layer=POLY_cond $X=5.16 $Y=1.65 $X2=4.86
+ $Y2=1.65
r61 1 5 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.785 $Y=1.725
+ $X2=4.86 $Y2=1.65
r62 1 3 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=4.785 $Y=1.725
+ $X2=4.785 $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4BB_2%VPWR 1 2 3 4 5 6 21 25 29 33 37 43 47 49
+ 54 55 56 57 58 60 72 77 83 86 89 93
r82 92 93 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r83 89 90 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r84 86 87 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r85 83 84 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r86 81 93 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33 $X2=6
+ $Y2=3.33
r87 81 90 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=4.56 $Y2=3.33
r88 80 81 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r89 78 89 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.735 $Y=3.33
+ $X2=4.57 $Y2=3.33
r90 78 80 51.2139 $w=1.68e-07 $l=7.85e-07 $layer=LI1_cond $X=4.735 $Y=3.33
+ $X2=5.52 $Y2=3.33
r91 77 92 4.48746 $w=1.7e-07 $l=2.97e-07 $layer=LI1_cond $X=5.645 $Y=3.33
+ $X2=5.942 $Y2=3.33
r92 77 80 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=5.645 $Y=3.33
+ $X2=5.52 $Y2=3.33
r93 76 90 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r94 76 87 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.6 $Y2=3.33
r95 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r96 73 86 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.875 $Y=3.33
+ $X2=3.71 $Y2=3.33
r97 73 75 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=3.875 $Y=3.33
+ $X2=4.08 $Y2=3.33
r98 72 89 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.405 $Y=3.33
+ $X2=4.57 $Y2=3.33
r99 72 75 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=4.405 $Y=3.33
+ $X2=4.08 $Y2=3.33
r100 70 71 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r101 68 71 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r102 68 84 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.72 $Y2=3.33
r103 67 68 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r104 65 83 6.70225 $w=1.7e-07 $l=1.18e-07 $layer=LI1_cond $X=0.795 $Y=3.33
+ $X2=0.677 $Y2=3.33
r105 65 67 57.738 $w=1.68e-07 $l=8.85e-07 $layer=LI1_cond $X=0.795 $Y=3.33
+ $X2=1.68 $Y2=3.33
r106 63 84 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r107 62 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r108 60 83 6.70225 $w=1.7e-07 $l=1.17e-07 $layer=LI1_cond $X=0.56 $Y=3.33
+ $X2=0.677 $Y2=3.33
r109 60 62 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=0.56 $Y=3.33
+ $X2=0.24 $Y2=3.33
r110 58 87 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r111 58 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.64 $Y2=3.33
r112 56 70 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=2.685 $Y=3.33
+ $X2=2.64 $Y2=3.33
r113 56 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.685 $Y=3.33
+ $X2=2.85 $Y2=3.33
r114 54 67 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=1.825 $Y=3.33
+ $X2=1.68 $Y2=3.33
r115 54 55 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.825 $Y=3.33
+ $X2=1.99 $Y2=3.33
r116 53 70 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=2.155 $Y=3.33
+ $X2=2.64 $Y2=3.33
r117 53 55 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.155 $Y=3.33
+ $X2=1.99 $Y2=3.33
r118 49 52 33.0018 $w=3.28e-07 $l=9.45e-07 $layer=LI1_cond $X=5.81 $Y=2.005
+ $X2=5.81 $Y2=2.95
r119 47 92 3.27872 $w=3.3e-07 $l=1.69245e-07 $layer=LI1_cond $X=5.81 $Y=3.245
+ $X2=5.942 $Y2=3.33
r120 47 52 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=5.81 $Y=3.245
+ $X2=5.81 $Y2=2.95
r121 43 46 32.1287 $w=3.28e-07 $l=9.2e-07 $layer=LI1_cond $X=4.57 $Y=2.03
+ $X2=4.57 $Y2=2.95
r122 41 89 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.57 $Y=3.245
+ $X2=4.57 $Y2=3.33
r123 41 46 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=4.57 $Y=3.245
+ $X2=4.57 $Y2=2.95
r124 37 40 27.0649 $w=3.28e-07 $l=7.75e-07 $layer=LI1_cond $X=3.71 $Y=2.175
+ $X2=3.71 $Y2=2.95
r125 35 86 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.71 $Y=3.245
+ $X2=3.71 $Y2=3.33
r126 35 40 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=3.71 $Y=3.245
+ $X2=3.71 $Y2=2.95
r127 34 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.015 $Y=3.33
+ $X2=2.85 $Y2=3.33
r128 33 86 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.545 $Y=3.33
+ $X2=3.71 $Y2=3.33
r129 33 34 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=3.545 $Y=3.33
+ $X2=3.015 $Y2=3.33
r130 29 32 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=2.85 $Y=2.27
+ $X2=2.85 $Y2=2.95
r131 27 57 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.85 $Y=3.245
+ $X2=2.85 $Y2=3.33
r132 27 32 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.85 $Y=3.245
+ $X2=2.85 $Y2=2.95
r133 23 55 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.99 $Y=3.245
+ $X2=1.99 $Y2=3.33
r134 23 25 14.8421 $w=3.28e-07 $l=4.25e-07 $layer=LI1_cond $X=1.99 $Y=3.245
+ $X2=1.99 $Y2=2.82
r135 19 83 0.207053 $w=2.35e-07 $l=8.5e-08 $layer=LI1_cond $X=0.677 $Y=3.245
+ $X2=0.677 $Y2=3.33
r136 19 21 54.6797 $w=2.33e-07 $l=1.115e-06 $layer=LI1_cond $X=0.677 $Y=3.245
+ $X2=0.677 $Y2=2.13
r137 6 52 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=5.67
+ $Y=1.835 $X2=5.81 $Y2=2.95
r138 6 49 400 $w=1.7e-07 $l=2.29565e-07 $layer=licon1_PDIFF $count=1 $X=5.67
+ $Y=1.835 $X2=5.81 $Y2=2.005
r139 5 46 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=4.43
+ $Y=1.835 $X2=4.57 $Y2=2.95
r140 5 43 400 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_PDIFF $count=1 $X=4.43
+ $Y=1.835 $X2=4.57 $Y2=2.03
r141 4 40 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=3.57
+ $Y=1.835 $X2=3.71 $Y2=2.95
r142 4 37 400 $w=1.7e-07 $l=4.0398e-07 $layer=licon1_PDIFF $count=1 $X=3.57
+ $Y=1.835 $X2=3.71 $Y2=2.175
r143 3 32 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=2.71
+ $Y=1.835 $X2=2.85 $Y2=2.95
r144 3 29 400 $w=1.7e-07 $l=5.00125e-07 $layer=licon1_PDIFF $count=1 $X=2.71
+ $Y=1.835 $X2=2.85 $Y2=2.27
r145 2 25 600 $w=1.7e-07 $l=1.04563e-06 $layer=licon1_PDIFF $count=1 $X=1.865
+ $Y=1.835 $X2=1.99 $Y2=2.82
r146 1 21 600 $w=1.7e-07 $l=3.35596e-07 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=1.865 $X2=0.71 $Y2=2.13
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4BB_2%Y 1 2 3 4 5 18 22 26 27 28 29 32 38 42 44
+ 46 49 50 54 55
r92 66 67 13.2207 $w=2.51e-07 $l=2.72e-07 $layer=LI1_cond $X=3.28 $Y=1.762
+ $X2=3.552 $Y2=1.762
r93 60 67 0.407084 $w=2.65e-07 $l=1.57e-07 $layer=LI1_cond $X=3.552 $Y=1.605
+ $X2=3.552 $Y2=1.762
r94 55 67 2.33307 $w=2.51e-07 $l=4.8e-08 $layer=LI1_cond $X=3.6 $Y=1.762
+ $X2=3.552 $Y2=1.762
r95 55 60 0.565349 $w=2.63e-07 $l=1.3e-08 $layer=LI1_cond $X=3.552 $Y=1.592
+ $X2=3.552 $Y2=1.605
r96 54 55 12.9161 $w=2.63e-07 $l=2.97e-07 $layer=LI1_cond $X=3.552 $Y=1.295
+ $X2=3.552 $Y2=1.592
r97 51 53 7.70806 $w=4.59e-07 $l=2.9e-07 $layer=LI1_cond $X=5.19 $Y=1.69
+ $X2=5.19 $Y2=1.98
r98 49 55 10.5579 $w=4.58e-07 $l=3.6e-07 $layer=LI1_cond $X=4.045 $Y=1.762
+ $X2=3.685 $Y2=1.762
r99 49 50 4.19778 $w=2.42e-07 $l=9.5e-08 $layer=LI1_cond $X=4.045 $Y=1.762
+ $X2=4.14 $Y2=1.762
r100 48 54 3.91396 $w=2.63e-07 $l=9e-08 $layer=LI1_cond $X=3.552 $Y=1.205
+ $X2=3.552 $Y2=1.295
r101 44 53 5.31394 $w=5.7e-07 $l=2.25e-07 $layer=LI1_cond $X=5.19 $Y=2.205
+ $X2=5.19 $Y2=1.98
r102 44 46 5.77055 $w=5.68e-07 $l=2.75e-07 $layer=LI1_cond $X=5.19 $Y=2.205
+ $X2=5.19 $Y2=2.48
r103 43 50 4.19778 $w=2.42e-07 $l=1.25956e-07 $layer=LI1_cond $X=4.235 $Y=1.69
+ $X2=4.14 $Y2=1.762
r104 42 51 6.62291 $w=1.7e-07 $l=2.85e-07 $layer=LI1_cond $X=4.905 $Y=1.69
+ $X2=5.19 $Y2=1.69
r105 42 43 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.905 $Y=1.69
+ $X2=4.235 $Y2=1.69
r106 38 40 54.2871 $w=1.88e-07 $l=9.3e-07 $layer=LI1_cond $X=4.14 $Y=1.98
+ $X2=4.14 $Y2=2.91
r107 36 50 2.23415 $w=1.9e-07 $l=1.58e-07 $layer=LI1_cond $X=4.14 $Y=1.92
+ $X2=4.14 $Y2=1.762
r108 36 38 3.50239 $w=1.88e-07 $l=6e-08 $layer=LI1_cond $X=4.14 $Y=1.92 $X2=4.14
+ $Y2=1.98
r109 32 34 54.2871 $w=1.88e-07 $l=9.3e-07 $layer=LI1_cond $X=3.28 $Y=1.98
+ $X2=3.28 $Y2=2.91
r110 30 66 2.36997 $w=1.9e-07 $l=1.58e-07 $layer=LI1_cond $X=3.28 $Y=1.92
+ $X2=3.28 $Y2=1.762
r111 30 32 3.50239 $w=1.88e-07 $l=6e-08 $layer=LI1_cond $X=3.28 $Y=1.92 $X2=3.28
+ $Y2=1.98
r112 28 66 5.61262 $w=2.51e-07 $l=1.24439e-07 $layer=LI1_cond $X=3.185 $Y=1.83
+ $X2=3.28 $Y2=1.762
r113 28 29 41.2828 $w=1.78e-07 $l=6.7e-07 $layer=LI1_cond $X=3.185 $Y=1.83
+ $X2=2.515 $Y2=1.83
r114 26 48 7.24806 $w=1.7e-07 $l=1.69245e-07 $layer=LI1_cond $X=3.42 $Y=1.12
+ $X2=3.552 $Y2=1.205
r115 26 27 64.262 $w=1.68e-07 $l=9.85e-07 $layer=LI1_cond $X=3.42 $Y=1.12
+ $X2=2.435 $Y2=1.12
r116 22 24 54.2871 $w=1.88e-07 $l=9.3e-07 $layer=LI1_cond $X=2.42 $Y=1.98
+ $X2=2.42 $Y2=2.91
r117 20 29 6.82297 $w=1.8e-07 $l=1.32571e-07 $layer=LI1_cond $X=2.42 $Y=1.92
+ $X2=2.515 $Y2=1.83
r118 20 22 3.50239 $w=1.88e-07 $l=6e-08 $layer=LI1_cond $X=2.42 $Y=1.92 $X2=2.42
+ $Y2=1.98
r119 16 27 6.9898 $w=1.7e-07 $l=1.49579e-07 $layer=LI1_cond $X=2.322 $Y=1.035
+ $X2=2.435 $Y2=1.12
r120 16 18 14.0854 $w=2.23e-07 $l=2.75e-07 $layer=LI1_cond $X=2.322 $Y=1.035
+ $X2=2.322 $Y2=0.76
r121 5 53 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=4.86
+ $Y=1.835 $X2=5 $Y2=1.98
r122 5 46 150 $w=1.7e-07 $l=8.66848e-07 $layer=licon1_PDIFF $count=4 $X=4.86
+ $Y=1.835 $X2=5.38 $Y2=2.48
r123 4 40 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=4
+ $Y=1.835 $X2=4.14 $Y2=2.91
r124 4 38 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=4
+ $Y=1.835 $X2=4.14 $Y2=1.98
r125 3 34 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=3.14
+ $Y=1.835 $X2=3.28 $Y2=2.91
r126 3 32 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=3.14
+ $Y=1.835 $X2=3.28 $Y2=1.98
r127 2 24 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=2.28
+ $Y=1.835 $X2=2.42 $Y2=2.91
r128 2 22 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.28
+ $Y=1.835 $X2=2.42 $Y2=1.98
r129 1 18 182 $w=1.7e-07 $l=5.90868e-07 $layer=licon1_NDIFF $count=1 $X=2.2
+ $Y=0.235 $X2=2.34 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4BB_2%VGND 1 2 11 15 17 19 29 30 33 36
r70 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r71 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r72 30 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=5.52
+ $Y2=0
r73 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6 $Y2=0
r74 27 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.685 $Y=0 $X2=5.52
+ $Y2=0
r75 27 29 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=5.685 $Y=0 $X2=6
+ $Y2=0
r76 26 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=5.52
+ $Y2=0
r77 25 26 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=5.04 $Y=0
+ $X2=5.04 $Y2=0
r78 23 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r79 22 25 250.524 $w=1.68e-07 $l=3.84e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=5.04
+ $Y2=0
r80 22 23 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=1.2 $Y=0
+ $X2=1.2 $Y2=0
r81 20 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.99 $Y=0 $X2=0.825
+ $Y2=0
r82 20 22 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=0.99 $Y=0 $X2=1.2
+ $Y2=0
r83 19 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.355 $Y=0 $X2=5.52
+ $Y2=0
r84 19 25 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=5.355 $Y=0 $X2=5.04
+ $Y2=0
r85 17 26 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=3.12 $Y=0 $X2=5.04
+ $Y2=0
r86 17 23 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=3.12 $Y=0 $X2=1.2
+ $Y2=0
r87 13 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.52 $Y=0.085
+ $X2=5.52 $Y2=0
r88 13 15 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=5.52 $Y=0.085
+ $X2=5.52 $Y2=0.38
r89 9 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.825 $Y=0.085
+ $X2=0.825 $Y2=0
r90 9 11 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=0.825 $Y=0.085
+ $X2=0.825 $Y2=0.43
r91 2 15 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.38
+ $Y=0.235 $X2=5.52 $Y2=0.38
r92 1 11 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=0.685
+ $Y=0.245 $X2=0.825 $Y2=0.43
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4BB_2%A_357_47# 1 2 3 12 14 15 20 23
c39 23 0 1.20189e-19 $X=2.77 $Y=0.38
r40 18 23 7.95398 $w=1.9e-07 $l=1.65e-07 $layer=LI1_cond $X=2.935 $Y=0.36
+ $X2=2.77 $Y2=0.36
r41 18 20 40.9307 $w=2.08e-07 $l=7.75e-07 $layer=LI1_cond $X=2.935 $Y=0.36
+ $X2=3.71 $Y2=0.36
r42 14 23 7.95398 $w=1.9e-07 $l=1.74714e-07 $layer=LI1_cond $X=2.605 $Y=0.34
+ $X2=2.77 $Y2=0.36
r43 14 15 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=2.605 $Y=0.34
+ $X2=2.015 $Y2=0.34
r44 10 15 6.87494 $w=1.7e-07 $l=1.36015e-07 $layer=LI1_cond $X=1.915 $Y=0.425
+ $X2=2.015 $Y2=0.34
r45 10 12 0.831818 $w=1.98e-07 $l=1.5e-08 $layer=LI1_cond $X=1.915 $Y=0.425
+ $X2=1.915 $Y2=0.44
r46 3 20 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=3.57
+ $Y=0.235 $X2=3.71 $Y2=0.38
r47 2 23 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.63
+ $Y=0.235 $X2=2.77 $Y2=0.38
r48 1 12 91 $w=1.7e-07 $l=2.60096e-07 $layer=licon1_NDIFF $count=2 $X=1.785
+ $Y=0.235 $X2=1.91 $Y2=0.44
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4BB_2%A_614_47# 1 2 11
r19 8 11 69.1466 $w=2.28e-07 $l=1.38e-06 $layer=LI1_cond $X=3.28 $Y=0.75
+ $X2=4.66 $Y2=0.75
r20 2 11 182 $w=1.7e-07 $l=5.80797e-07 $layer=licon1_NDIFF $count=1 $X=4.52
+ $Y=0.235 $X2=4.66 $Y2=0.75
r21 1 8 182 $w=1.7e-07 $l=5.90741e-07 $layer=licon1_NDIFF $count=1 $X=3.07
+ $Y=0.235 $X2=3.28 $Y2=0.73
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4BB_2%A_821_47# 1 2 3 10 14 16 17 20
r31 18 20 28.5895 $w=2.58e-07 $l=6.45e-07 $layer=LI1_cond $X=5.985 $Y=1.065
+ $X2=5.985 $Y2=0.42
r32 16 18 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=5.855 $Y=1.15
+ $X2=5.985 $Y2=1.065
r33 16 17 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.855 $Y=1.15
+ $X2=5.185 $Y2=1.15
r34 15 17 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=5.09 $Y=1.065
+ $X2=5.185 $Y2=1.15
r35 14 23 3.59031 $w=1.9e-07 $l=1.05e-07 $layer=LI1_cond $X=5.09 $Y=0.465
+ $X2=5.09 $Y2=0.36
r36 14 15 35.0239 $w=1.88e-07 $l=6e-07 $layer=LI1_cond $X=5.09 $Y=0.465 $X2=5.09
+ $Y2=1.065
r37 10 23 3.24837 $w=2.1e-07 $l=9.5e-08 $layer=LI1_cond $X=4.995 $Y=0.36
+ $X2=5.09 $Y2=0.36
r38 10 12 40.4026 $w=2.08e-07 $l=7.65e-07 $layer=LI1_cond $X=4.995 $Y=0.36
+ $X2=4.23 $Y2=0.36
r39 3 20 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=5.81
+ $Y=0.235 $X2=5.95 $Y2=0.42
r40 2 23 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=4.95
+ $Y=0.235 $X2=5.09 $Y2=0.42
r41 1 12 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=4.105
+ $Y=0.235 $X2=4.23 $Y2=0.38
.ends

