* File: sky130_fd_sc_lp__and2_2.pxi.spice
* Created: Fri Aug 28 10:04:22 2020
* 
x_PM_SKY130_FD_SC_LP__AND2_2%A N_A_c_55_n N_A_M1006_g N_A_c_51_n N_A_M1003_g
+ N_A_c_52_n A A N_A_c_53_n N_A_c_54_n PM_SKY130_FD_SC_LP__AND2_2%A
x_PM_SKY130_FD_SC_LP__AND2_2%B N_B_M1007_g N_B_M1000_g B N_B_c_87_n N_B_c_88_n
+ PM_SKY130_FD_SC_LP__AND2_2%B
x_PM_SKY130_FD_SC_LP__AND2_2%A_46_47# N_A_46_47#_M1003_s N_A_46_47#_M1006_d
+ N_A_46_47#_M1002_g N_A_46_47#_M1001_g N_A_46_47#_c_125_n N_A_46_47#_M1005_g
+ N_A_46_47#_M1004_g N_A_46_47#_c_128_n N_A_46_47#_c_129_n N_A_46_47#_c_130_n
+ N_A_46_47#_c_131_n N_A_46_47#_c_138_n N_A_46_47#_c_132_n N_A_46_47#_c_133_n
+ N_A_46_47#_c_191_p N_A_46_47#_c_163_n N_A_46_47#_c_134_n N_A_46_47#_c_135_n
+ PM_SKY130_FD_SC_LP__AND2_2%A_46_47#
x_PM_SKY130_FD_SC_LP__AND2_2%VPWR N_VPWR_M1006_s N_VPWR_M1000_d N_VPWR_M1004_d
+ N_VPWR_c_210_n N_VPWR_c_211_n N_VPWR_c_212_n N_VPWR_c_213_n N_VPWR_c_214_n
+ VPWR N_VPWR_c_215_n N_VPWR_c_216_n N_VPWR_c_217_n N_VPWR_c_209_n
+ PM_SKY130_FD_SC_LP__AND2_2%VPWR
x_PM_SKY130_FD_SC_LP__AND2_2%X N_X_M1002_d N_X_M1001_s N_X_c_242_n N_X_c_239_n X
+ X X N_X_c_240_n X PM_SKY130_FD_SC_LP__AND2_2%X
x_PM_SKY130_FD_SC_LP__AND2_2%VGND N_VGND_M1007_d N_VGND_M1005_s N_VGND_c_268_n
+ N_VGND_c_269_n N_VGND_c_270_n VGND N_VGND_c_271_n N_VGND_c_272_n
+ N_VGND_c_273_n N_VGND_c_274_n PM_SKY130_FD_SC_LP__AND2_2%VGND
cc_1 VNB N_A_c_51_n 0.0191349f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=0.765
cc_2 VNB N_A_c_52_n 0.0605573f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.46
cc_3 VNB N_A_c_53_n 0.057775f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.12
cc_4 VNB N_A_c_54_n 0.00111806f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.12
cc_5 VNB N_B_M1007_g 0.037553f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=2.195
cc_6 VNB N_B_M1000_g 0.00917592f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.12
cc_7 VNB N_B_c_87_n 0.0295893f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_8 VNB N_B_c_88_n 0.00763228f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_46_47#_M1002_g 0.0208283f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=0.765
cc_10 VNB N_A_46_47#_M1001_g 0.00269534f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_46_47#_c_125_n 0.0147888f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.12
cc_12 VNB N_A_46_47#_M1005_g 0.0276947f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_46_47#_M1004_g 0.0177377f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_46_47#_c_128_n 0.0106787f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_46_47#_c_129_n 0.016165f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_46_47#_c_130_n 0.00937438f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_46_47#_c_131_n 0.00748178f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_46_47#_c_132_n 0.00743847f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_46_47#_c_133_n 0.00194371f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_46_47#_c_134_n 0.00148477f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_46_47#_c_135_n 0.0297718f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_VPWR_c_209_n 0.103974f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_X_c_239_n 0.00207055f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_X_c_240_n 0.00252246f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_268_n 0.00503582f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=0.765
cc_26 VNB N_VGND_c_269_n 0.0118897f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_27 VNB N_VGND_c_270_n 0.0484852f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_271_n 0.0299618f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.12
cc_29 VNB N_VGND_c_272_n 0.0172812f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.665
cc_30 VNB N_VGND_c_273_n 0.00631792f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_274_n 0.15351f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VPB N_A_c_55_n 0.0231414f $X=-0.19 $Y=1.655 $X2=0.5 $Y2=1.875
cc_33 VPB N_A_c_52_n 0.0282416f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.46
cc_34 VPB N_A_c_54_n 0.00978796f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.12
cc_35 VPB N_B_M1000_g 0.0316267f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.12
cc_36 VPB N_A_46_47#_M1001_g 0.0226644f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_37 VPB N_A_46_47#_M1004_g 0.0265103f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_38 VPB N_A_46_47#_c_138_n 0.00415393f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_39 VPB N_A_46_47#_c_132_n 0.00473426f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_40 VPB N_A_46_47#_c_133_n 9.50817e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_41 VPB N_VPWR_c_210_n 0.0123504f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.46
cc_42 VPB N_VPWR_c_211_n 0.0588443f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_43 VPB N_VPWR_c_212_n 0.0168895f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.12
cc_44 VPB N_VPWR_c_213_n 0.0118638f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.295
cc_45 VPB N_VPWR_c_214_n 0.0646935f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.665
cc_46 VPB N_VPWR_c_215_n 0.0179158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_47 VPB N_VPWR_c_216_n 0.0170188f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_48 VPB N_VPWR_c_217_n 0.0066101f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_49 VPB N_VPWR_c_209_n 0.0631045f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_50 VPB N_X_c_240_n 0.00127276f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_51 N_A_c_51_n N_B_M1007_g 0.0506064f $X=0.57 $Y=0.765 $X2=0 $Y2=0
cc_52 N_A_c_53_n N_B_M1007_g 0.00792171f $X=0.27 $Y=1.12 $X2=0 $Y2=0
cc_53 N_A_c_54_n N_B_M1007_g 5.38096e-19 $X=0.27 $Y=1.12 $X2=0 $Y2=0
cc_54 N_A_c_52_n N_B_M1000_g 0.0224632f $X=0.27 $Y=1.46 $X2=0 $Y2=0
cc_55 N_A_c_54_n N_B_M1000_g 8.26537e-19 $X=0.27 $Y=1.12 $X2=0 $Y2=0
cc_56 N_A_c_52_n N_B_c_87_n 0.0176934f $X=0.27 $Y=1.46 $X2=0 $Y2=0
cc_57 N_A_c_54_n N_B_c_87_n 6.89525e-19 $X=0.27 $Y=1.12 $X2=0 $Y2=0
cc_58 N_A_c_52_n N_B_c_88_n 0.00192792f $X=0.27 $Y=1.46 $X2=0 $Y2=0
cc_59 N_A_c_53_n N_B_c_88_n 0.00106262f $X=0.27 $Y=1.12 $X2=0 $Y2=0
cc_60 N_A_c_54_n N_B_c_88_n 0.0244695f $X=0.27 $Y=1.12 $X2=0 $Y2=0
cc_61 N_A_c_51_n N_A_46_47#_c_129_n 0.0083467f $X=0.57 $Y=0.765 $X2=0 $Y2=0
cc_62 N_A_c_51_n N_A_46_47#_c_130_n 0.00444617f $X=0.57 $Y=0.765 $X2=0 $Y2=0
cc_63 N_A_c_53_n N_A_46_47#_c_130_n 0.00552355f $X=0.27 $Y=1.12 $X2=0 $Y2=0
cc_64 N_A_c_51_n N_A_46_47#_c_131_n 0.00155647f $X=0.57 $Y=0.765 $X2=0 $Y2=0
cc_65 N_A_c_53_n N_A_46_47#_c_131_n 0.0170643f $X=0.27 $Y=1.12 $X2=0 $Y2=0
cc_66 N_A_c_54_n N_A_46_47#_c_131_n 0.0208405f $X=0.27 $Y=1.12 $X2=0 $Y2=0
cc_67 N_A_c_52_n N_A_46_47#_c_138_n 0.00397717f $X=0.27 $Y=1.46 $X2=0 $Y2=0
cc_68 N_A_c_54_n N_A_46_47#_c_138_n 0.00644746f $X=0.27 $Y=1.12 $X2=0 $Y2=0
cc_69 N_A_c_52_n N_A_46_47#_c_133_n 0.00141817f $X=0.27 $Y=1.46 $X2=0 $Y2=0
cc_70 N_A_c_54_n N_A_46_47#_c_133_n 0.0134523f $X=0.27 $Y=1.12 $X2=0 $Y2=0
cc_71 N_A_c_55_n N_VPWR_c_211_n 0.0108046f $X=0.5 $Y=1.875 $X2=0 $Y2=0
cc_72 N_A_c_52_n N_VPWR_c_211_n 0.00445894f $X=0.27 $Y=1.46 $X2=0 $Y2=0
cc_73 N_A_c_54_n N_VPWR_c_211_n 0.025532f $X=0.27 $Y=1.12 $X2=0 $Y2=0
cc_74 N_A_c_55_n N_VPWR_c_209_n 0.00330899f $X=0.5 $Y=1.875 $X2=0 $Y2=0
cc_75 N_A_c_51_n N_VGND_c_271_n 0.0042339f $X=0.57 $Y=0.765 $X2=0 $Y2=0
cc_76 N_A_c_53_n N_VGND_c_271_n 4.685e-19 $X=0.27 $Y=1.12 $X2=0 $Y2=0
cc_77 N_A_c_51_n N_VGND_c_274_n 0.00695911f $X=0.57 $Y=0.765 $X2=0 $Y2=0
cc_78 N_B_M1007_g N_A_46_47#_M1002_g 0.0248238f $X=0.93 $Y=0.445 $X2=0 $Y2=0
cc_79 N_B_M1000_g N_A_46_47#_M1001_g 0.0179911f $X=0.93 $Y=2.195 $X2=0 $Y2=0
cc_80 N_B_M1007_g N_A_46_47#_c_129_n 0.00153508f $X=0.93 $Y=0.445 $X2=0 $Y2=0
cc_81 N_B_M1007_g N_A_46_47#_c_130_n 0.0125956f $X=0.93 $Y=0.445 $X2=0 $Y2=0
cc_82 N_B_c_87_n N_A_46_47#_c_130_n 0.00108763f $X=0.84 $Y=1.32 $X2=0 $Y2=0
cc_83 N_B_c_88_n N_A_46_47#_c_130_n 0.0220777f $X=0.84 $Y=1.32 $X2=0 $Y2=0
cc_84 N_B_M1000_g N_A_46_47#_c_138_n 0.00502546f $X=0.93 $Y=2.195 $X2=0 $Y2=0
cc_85 N_B_M1000_g N_A_46_47#_c_132_n 0.0154289f $X=0.93 $Y=2.195 $X2=0 $Y2=0
cc_86 N_B_c_87_n N_A_46_47#_c_132_n 2.36777e-19 $X=0.84 $Y=1.32 $X2=0 $Y2=0
cc_87 N_B_c_88_n N_A_46_47#_c_132_n 0.0113538f $X=0.84 $Y=1.32 $X2=0 $Y2=0
cc_88 N_B_c_87_n N_A_46_47#_c_133_n 0.00423302f $X=0.84 $Y=1.32 $X2=0 $Y2=0
cc_89 N_B_c_88_n N_A_46_47#_c_133_n 0.0190968f $X=0.84 $Y=1.32 $X2=0 $Y2=0
cc_90 N_B_c_87_n N_A_46_47#_c_163_n 0.00110914f $X=0.84 $Y=1.32 $X2=0 $Y2=0
cc_91 N_B_M1007_g N_A_46_47#_c_134_n 0.00574f $X=0.93 $Y=0.445 $X2=0 $Y2=0
cc_92 N_B_c_88_n N_A_46_47#_c_134_n 0.0179949f $X=0.84 $Y=1.32 $X2=0 $Y2=0
cc_93 N_B_c_87_n N_A_46_47#_c_135_n 0.0217502f $X=0.84 $Y=1.32 $X2=0 $Y2=0
cc_94 N_B_c_88_n N_A_46_47#_c_135_n 6.46178e-19 $X=0.84 $Y=1.32 $X2=0 $Y2=0
cc_95 N_B_M1000_g N_VPWR_c_211_n 5.51198e-19 $X=0.93 $Y=2.195 $X2=0 $Y2=0
cc_96 N_B_M1000_g N_VPWR_c_212_n 0.00303159f $X=0.93 $Y=2.195 $X2=0 $Y2=0
cc_97 N_B_M1000_g N_VPWR_c_209_n 0.00393927f $X=0.93 $Y=2.195 $X2=0 $Y2=0
cc_98 N_B_M1007_g N_VGND_c_268_n 0.00322925f $X=0.93 $Y=0.445 $X2=0 $Y2=0
cc_99 N_B_M1007_g N_VGND_c_271_n 0.00433717f $X=0.93 $Y=0.445 $X2=0 $Y2=0
cc_100 N_B_M1007_g N_VGND_c_274_n 0.00596326f $X=0.93 $Y=0.445 $X2=0 $Y2=0
cc_101 N_A_46_47#_M1001_g N_VPWR_c_212_n 0.00607841f $X=1.455 $Y=2.465 $X2=0
+ $Y2=0
cc_102 N_A_46_47#_c_138_n N_VPWR_c_212_n 0.00316461f $X=0.715 $Y=2.195 $X2=0
+ $Y2=0
cc_103 N_A_46_47#_c_132_n N_VPWR_c_212_n 0.0274404f $X=1.235 $Y=1.685 $X2=0
+ $Y2=0
cc_104 N_A_46_47#_c_135_n N_VPWR_c_212_n 5.72192e-19 $X=1.38 $Y=1.345 $X2=0
+ $Y2=0
cc_105 N_A_46_47#_M1004_g N_VPWR_c_214_n 0.00758113f $X=1.885 $Y=2.465 $X2=0
+ $Y2=0
cc_106 N_A_46_47#_M1001_g N_VPWR_c_216_n 0.00585385f $X=1.455 $Y=2.465 $X2=0
+ $Y2=0
cc_107 N_A_46_47#_M1004_g N_VPWR_c_216_n 0.00579312f $X=1.885 $Y=2.465 $X2=0
+ $Y2=0
cc_108 N_A_46_47#_M1001_g N_VPWR_c_209_n 0.0118494f $X=1.455 $Y=2.465 $X2=0
+ $Y2=0
cc_109 N_A_46_47#_M1004_g N_VPWR_c_209_n 0.0113933f $X=1.885 $Y=2.465 $X2=0
+ $Y2=0
cc_110 N_A_46_47#_M1005_g N_X_c_242_n 0.00769181f $X=1.885 $Y=0.655 $X2=0 $Y2=0
cc_111 N_A_46_47#_M1002_g N_X_c_239_n 6.01622e-19 $X=1.455 $Y=0.655 $X2=0 $Y2=0
cc_112 N_A_46_47#_c_125_n N_X_c_239_n 6.09999e-19 $X=1.81 $Y=1.345 $X2=0 $Y2=0
cc_113 N_A_46_47#_M1005_g N_X_c_239_n 0.00124306f $X=1.885 $Y=0.655 $X2=0 $Y2=0
cc_114 N_A_46_47#_c_134_n N_X_c_239_n 0.00814645f $X=1.35 $Y=1.27 $X2=0 $Y2=0
cc_115 N_A_46_47#_c_125_n X 0.0022221f $X=1.81 $Y=1.345 $X2=0 $Y2=0
cc_116 N_A_46_47#_M1004_g X 0.0108144f $X=1.885 $Y=2.465 $X2=0 $Y2=0
cc_117 N_A_46_47#_M1002_g N_X_c_240_n 0.00127767f $X=1.455 $Y=0.655 $X2=0 $Y2=0
cc_118 N_A_46_47#_M1001_g N_X_c_240_n 0.00478948f $X=1.455 $Y=2.465 $X2=0 $Y2=0
cc_119 N_A_46_47#_c_125_n N_X_c_240_n 0.0107265f $X=1.81 $Y=1.345 $X2=0 $Y2=0
cc_120 N_A_46_47#_M1005_g N_X_c_240_n 0.00836085f $X=1.885 $Y=0.655 $X2=0 $Y2=0
cc_121 N_A_46_47#_M1004_g N_X_c_240_n 0.0203599f $X=1.885 $Y=2.465 $X2=0 $Y2=0
cc_122 N_A_46_47#_c_128_n N_X_c_240_n 0.0058471f $X=1.885 $Y=1.345 $X2=0 $Y2=0
cc_123 N_A_46_47#_c_132_n N_X_c_240_n 0.0135986f $X=1.235 $Y=1.685 $X2=0 $Y2=0
cc_124 N_A_46_47#_c_191_p N_X_c_240_n 0.0236051f $X=1.35 $Y=1.385 $X2=0 $Y2=0
cc_125 N_A_46_47#_c_134_n N_X_c_240_n 0.0102619f $X=1.35 $Y=1.27 $X2=0 $Y2=0
cc_126 N_A_46_47#_c_135_n N_X_c_240_n 0.0012746f $X=1.38 $Y=1.345 $X2=0 $Y2=0
cc_127 N_A_46_47#_c_130_n N_VGND_M1007_d 0.0063976f $X=1.235 $Y=0.78 $X2=-0.19
+ $Y2=-0.245
cc_128 N_A_46_47#_c_134_n N_VGND_M1007_d 0.00253326f $X=1.35 $Y=1.27 $X2=-0.19
+ $Y2=-0.245
cc_129 N_A_46_47#_M1002_g N_VGND_c_268_n 0.00180476f $X=1.455 $Y=0.655 $X2=0
+ $Y2=0
cc_130 N_A_46_47#_c_130_n N_VGND_c_268_n 0.0220744f $X=1.235 $Y=0.78 $X2=0 $Y2=0
cc_131 N_A_46_47#_M1005_g N_VGND_c_270_n 0.00677253f $X=1.885 $Y=0.655 $X2=0
+ $Y2=0
cc_132 N_A_46_47#_c_129_n N_VGND_c_271_n 0.0179718f $X=0.355 $Y=0.445 $X2=0
+ $Y2=0
cc_133 N_A_46_47#_c_130_n N_VGND_c_271_n 0.00769607f $X=1.235 $Y=0.78 $X2=0
+ $Y2=0
cc_134 N_A_46_47#_M1002_g N_VGND_c_272_n 0.00560083f $X=1.455 $Y=0.655 $X2=0
+ $Y2=0
cc_135 N_A_46_47#_M1005_g N_VGND_c_272_n 0.00579312f $X=1.885 $Y=0.655 $X2=0
+ $Y2=0
cc_136 N_A_46_47#_c_130_n N_VGND_c_272_n 5.51759e-19 $X=1.235 $Y=0.78 $X2=0
+ $Y2=0
cc_137 N_A_46_47#_M1003_s N_VGND_c_274_n 0.00216892f $X=0.23 $Y=0.235 $X2=0
+ $Y2=0
cc_138 N_A_46_47#_M1002_g N_VGND_c_274_n 0.0100171f $X=1.455 $Y=0.655 $X2=0
+ $Y2=0
cc_139 N_A_46_47#_M1005_g N_VGND_c_274_n 0.0113933f $X=1.885 $Y=0.655 $X2=0
+ $Y2=0
cc_140 N_A_46_47#_c_129_n N_VGND_c_274_n 0.0124213f $X=0.355 $Y=0.445 $X2=0
+ $Y2=0
cc_141 N_A_46_47#_c_130_n N_VGND_c_274_n 0.0150124f $X=1.235 $Y=0.78 $X2=0 $Y2=0
cc_142 N_VPWR_c_209_n N_X_M1001_s 0.00223559f $X=2.16 $Y=3.33 $X2=0 $Y2=0
cc_143 N_VPWR_c_216_n X 0.0159213f $X=1.985 $Y=3.33 $X2=0 $Y2=0
cc_144 N_VPWR_c_209_n X 0.0109109f $X=2.16 $Y=3.33 $X2=0 $Y2=0
cc_145 N_VPWR_c_214_n N_X_c_240_n 0.0466161f $X=2.1 $Y=1.98 $X2=0 $Y2=0
cc_146 N_X_c_242_n N_VGND_c_270_n 0.0303711f $X=1.67 $Y=0.42 $X2=0 $Y2=0
cc_147 N_X_c_242_n N_VGND_c_272_n 0.0143246f $X=1.67 $Y=0.42 $X2=0 $Y2=0
cc_148 N_X_M1002_d N_VGND_c_274_n 0.00380103f $X=1.53 $Y=0.235 $X2=0 $Y2=0
cc_149 N_X_c_242_n N_VGND_c_274_n 0.00916141f $X=1.67 $Y=0.42 $X2=0 $Y2=0
cc_150 A_129_47# N_VGND_c_274_n 0.0026263f $X=0.645 $Y=0.235 $X2=2.16 $Y2=0
