* File: sky130_fd_sc_lp__a22oi_4.pxi.spice
* Created: Wed Sep  2 09:23:17 2020
* 
x_PM_SKY130_FD_SC_LP__A22OI_4%B2 N_B2_c_114_n N_B2_M1009_g N_B2_M1006_g
+ N_B2_c_116_n N_B2_M1010_g N_B2_M1015_g N_B2_c_118_n N_B2_M1018_g N_B2_M1023_g
+ N_B2_c_120_n N_B2_M1028_g N_B2_M1027_g B2 B2 B2 B2 B2 N_B2_c_123_n
+ N_B2_c_124_n PM_SKY130_FD_SC_LP__A22OI_4%B2
x_PM_SKY130_FD_SC_LP__A22OI_4%B1 N_B1_c_201_n N_B1_M1001_g N_B1_M1000_g
+ N_B1_c_203_n N_B1_M1011_g N_B1_M1008_g N_B1_c_205_n N_B1_M1020_g N_B1_M1016_g
+ N_B1_c_207_n N_B1_M1024_g N_B1_M1019_g B1 B1 B1 B1 N_B1_c_210_n N_B1_c_211_n
+ B1 PM_SKY130_FD_SC_LP__A22OI_4%B1
x_PM_SKY130_FD_SC_LP__A22OI_4%A1 N_A1_M1013_g N_A1_c_297_n N_A1_M1004_g
+ N_A1_M1017_g N_A1_c_299_n N_A1_M1005_g N_A1_M1026_g N_A1_c_301_n N_A1_M1021_g
+ N_A1_M1030_g N_A1_c_303_n N_A1_M1022_g A1 A1 A1 A1 N_A1_c_305_n
+ PM_SKY130_FD_SC_LP__A22OI_4%A1
x_PM_SKY130_FD_SC_LP__A22OI_4%A2 N_A2_c_387_n N_A2_M1003_g N_A2_M1002_g
+ N_A2_c_388_n N_A2_M1007_g N_A2_M1012_g N_A2_c_389_n N_A2_M1025_g N_A2_M1014_g
+ N_A2_c_390_n N_A2_M1029_g N_A2_M1031_g A2 A2 A2 N_A2_c_386_n
+ PM_SKY130_FD_SC_LP__A22OI_4%A2
x_PM_SKY130_FD_SC_LP__A22OI_4%A_89_367# N_A_89_367#_M1006_s N_A_89_367#_M1015_s
+ N_A_89_367#_M1027_s N_A_89_367#_M1008_s N_A_89_367#_M1019_s
+ N_A_89_367#_M1017_d N_A_89_367#_M1030_d N_A_89_367#_M1007_s
+ N_A_89_367#_M1029_s N_A_89_367#_c_453_n N_A_89_367#_c_454_n
+ N_A_89_367#_c_465_n N_A_89_367#_c_509_p N_A_89_367#_c_467_n
+ N_A_89_367#_c_513_p N_A_89_367#_c_469_n N_A_89_367#_c_516_p
+ N_A_89_367#_c_471_n N_A_89_367#_c_534_p N_A_89_367#_c_455_n
+ N_A_89_367#_c_456_n N_A_89_367#_c_538_p N_A_89_367#_c_457_n
+ N_A_89_367#_c_458_n N_A_89_367#_c_527_p N_A_89_367#_c_488_n
+ N_A_89_367#_c_528_p N_A_89_367#_c_495_n N_A_89_367#_c_459_n
+ N_A_89_367#_c_460_n N_A_89_367#_c_535_p N_A_89_367#_c_536_p
+ N_A_89_367#_c_537_p N_A_89_367#_c_461_n N_A_89_367#_c_501_n
+ PM_SKY130_FD_SC_LP__A22OI_4%A_89_367#
x_PM_SKY130_FD_SC_LP__A22OI_4%Y N_Y_M1001_s N_Y_M1020_s N_Y_M1004_s N_Y_M1021_s
+ N_Y_M1006_d N_Y_M1023_d N_Y_M1000_d N_Y_M1016_d N_Y_c_571_n N_Y_c_564_n
+ N_Y_c_565_n N_Y_c_582_n N_Y_c_566_n N_Y_c_562_n N_Y_c_589_n N_Y_c_568_n
+ N_Y_c_612_n N_Y_c_569_n N_Y_c_570_n N_Y_c_631_n N_Y_c_563_n Y Y Y Y Y
+ N_Y_c_594_n PM_SKY130_FD_SC_LP__A22OI_4%Y
x_PM_SKY130_FD_SC_LP__A22OI_4%VPWR N_VPWR_M1013_s N_VPWR_M1026_s N_VPWR_M1003_d
+ N_VPWR_M1025_d N_VPWR_c_677_n N_VPWR_c_678_n N_VPWR_c_679_n N_VPWR_c_680_n
+ N_VPWR_c_681_n N_VPWR_c_682_n N_VPWR_c_683_n N_VPWR_c_684_n VPWR
+ N_VPWR_c_685_n N_VPWR_c_686_n N_VPWR_c_687_n N_VPWR_c_676_n N_VPWR_c_689_n
+ N_VPWR_c_690_n PM_SKY130_FD_SC_LP__A22OI_4%VPWR
x_PM_SKY130_FD_SC_LP__A22OI_4%A_63_65# N_A_63_65#_M1009_d N_A_63_65#_M1010_d
+ N_A_63_65#_M1028_d N_A_63_65#_M1011_d N_A_63_65#_M1024_d N_A_63_65#_c_784_n
+ N_A_63_65#_c_792_n N_A_63_65#_c_785_n N_A_63_65#_c_786_n N_A_63_65#_c_798_n
+ N_A_63_65#_c_806_n N_A_63_65#_c_787_n N_A_63_65#_c_788_n N_A_63_65#_c_789_n
+ N_A_63_65#_c_803_n N_A_63_65#_c_790_n PM_SKY130_FD_SC_LP__A22OI_4%A_63_65#
x_PM_SKY130_FD_SC_LP__A22OI_4%VGND N_VGND_M1009_s N_VGND_M1018_s N_VGND_M1002_d
+ N_VGND_M1014_d N_VGND_c_838_n N_VGND_c_839_n N_VGND_c_840_n N_VGND_c_841_n
+ VGND N_VGND_c_842_n N_VGND_c_843_n N_VGND_c_844_n N_VGND_c_845_n
+ N_VGND_c_846_n N_VGND_c_847_n N_VGND_c_848_n N_VGND_c_849_n N_VGND_c_850_n
+ PM_SKY130_FD_SC_LP__A22OI_4%VGND
x_PM_SKY130_FD_SC_LP__A22OI_4%A_867_47# N_A_867_47#_M1004_d N_A_867_47#_M1005_d
+ N_A_867_47#_M1022_d N_A_867_47#_M1012_s N_A_867_47#_M1031_s
+ N_A_867_47#_c_935_n N_A_867_47#_c_944_n N_A_867_47#_c_945_n
+ N_A_867_47#_c_948_n N_A_867_47#_c_982_n N_A_867_47#_c_936_n
+ N_A_867_47#_c_937_n N_A_867_47#_c_938_n PM_SKY130_FD_SC_LP__A22OI_4%A_867_47#
cc_1 VNB N_B2_c_114_n 0.021262f $X=-0.19 $Y=-0.245 $X2=0.655 $Y2=1.275
cc_2 VNB N_B2_M1006_g 0.00394324f $X=-0.19 $Y=-0.245 $X2=0.785 $Y2=2.465
cc_3 VNB N_B2_c_116_n 0.0157949f $X=-0.19 $Y=-0.245 $X2=1.085 $Y2=1.275
cc_4 VNB N_B2_M1015_g 0.00249196f $X=-0.19 $Y=-0.245 $X2=1.215 $Y2=2.465
cc_5 VNB N_B2_c_118_n 0.0157949f $X=-0.19 $Y=-0.245 $X2=1.515 $Y2=1.275
cc_6 VNB N_B2_M1023_g 0.00249196f $X=-0.19 $Y=-0.245 $X2=1.645 $Y2=2.465
cc_7 VNB N_B2_c_120_n 0.0165356f $X=-0.19 $Y=-0.245 $X2=1.945 $Y2=1.275
cc_8 VNB N_B2_M1027_g 0.00256697f $X=-0.19 $Y=-0.245 $X2=2.075 $Y2=2.465
cc_9 VNB B2 0.0340307f $X=-0.19 $Y=-0.245 $X2=2.075 $Y2=1.21
cc_10 VNB N_B2_c_123_n 0.059687f $X=-0.19 $Y=-0.245 $X2=0.625 $Y2=1.44
cc_11 VNB N_B2_c_124_n 0.0841063f $X=-0.19 $Y=-0.245 $X2=2.075 $Y2=1.44
cc_12 VNB N_B1_c_201_n 0.0164878f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_B1_M1000_g 0.00208578f $X=-0.19 $Y=-0.245 $X2=0.785 $Y2=1.605
cc_14 VNB N_B1_c_203_n 0.0161955f $X=-0.19 $Y=-0.245 $X2=0.785 $Y2=2.465
cc_15 VNB N_B1_M1008_g 0.00263785f $X=-0.19 $Y=-0.245 $X2=1.215 $Y2=1.605
cc_16 VNB N_B1_c_205_n 0.0157063f $X=-0.19 $Y=-0.245 $X2=1.215 $Y2=2.465
cc_17 VNB N_B1_M1016_g 0.0026458f $X=-0.19 $Y=-0.245 $X2=1.645 $Y2=1.605
cc_18 VNB N_B1_c_207_n 0.0194324f $X=-0.19 $Y=-0.245 $X2=1.645 $Y2=2.465
cc_19 VNB N_B1_M1019_g 0.00275923f $X=-0.19 $Y=-0.245 $X2=2.075 $Y2=1.605
cc_20 VNB B1 0.0122105f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_21 VNB N_B1_c_210_n 0.103551f $X=-0.19 $Y=-0.245 $X2=1.305 $Y2=1.44
cc_22 VNB N_B1_c_211_n 0.00196937f $X=-0.19 $Y=-0.245 $X2=1.645 $Y2=1.44
cc_23 VNB N_A1_M1013_g 0.00716081f $X=-0.19 $Y=-0.245 $X2=0.655 $Y2=1.275
cc_24 VNB N_A1_c_297_n 0.0220814f $X=-0.19 $Y=-0.245 $X2=0.655 $Y2=0.745
cc_25 VNB N_A1_M1017_g 0.00706679f $X=-0.19 $Y=-0.245 $X2=1.085 $Y2=1.275
cc_26 VNB N_A1_c_299_n 0.0162054f $X=-0.19 $Y=-0.245 $X2=1.085 $Y2=0.745
cc_27 VNB N_A1_M1026_g 0.00731999f $X=-0.19 $Y=-0.245 $X2=1.515 $Y2=1.275
cc_28 VNB N_A1_c_301_n 0.0162054f $X=-0.19 $Y=-0.245 $X2=1.515 $Y2=0.745
cc_29 VNB N_A1_M1030_g 0.00798824f $X=-0.19 $Y=-0.245 $X2=1.945 $Y2=1.275
cc_30 VNB N_A1_c_303_n 0.0164438f $X=-0.19 $Y=-0.245 $X2=1.945 $Y2=0.745
cc_31 VNB A1 0.00947848f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_32 VNB N_A1_c_305_n 0.0976891f $X=-0.19 $Y=-0.245 $X2=1.085 $Y2=1.44
cc_33 VNB N_A2_M1002_g 0.0233464f $X=-0.19 $Y=-0.245 $X2=0.785 $Y2=1.605
cc_34 VNB N_A2_M1012_g 0.0233271f $X=-0.19 $Y=-0.245 $X2=1.215 $Y2=1.605
cc_35 VNB N_A2_M1014_g 0.0226024f $X=-0.19 $Y=-0.245 $X2=1.645 $Y2=1.605
cc_36 VNB N_A2_M1031_g 0.0306499f $X=-0.19 $Y=-0.245 $X2=2.075 $Y2=1.605
cc_37 VNB A2 0.0121507f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_38 VNB N_A2_c_386_n 0.080808f $X=-0.19 $Y=-0.245 $X2=0.965 $Y2=1.44
cc_39 VNB N_Y_c_562_n 0.00318651f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_Y_c_563_n 0.00892211f $X=-0.19 $Y=-0.245 $X2=1.645 $Y2=1.44
cc_41 VNB N_VPWR_c_676_n 0.342803f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_63_65#_c_784_n 0.0230663f $X=-0.19 $Y=-0.245 $X2=1.515 $Y2=0.745
cc_43 VNB N_A_63_65#_c_785_n 0.00742876f $X=-0.19 $Y=-0.245 $X2=1.645 $Y2=2.465
cc_44 VNB N_A_63_65#_c_786_n 0.00168668f $X=-0.19 $Y=-0.245 $X2=1.945 $Y2=1.275
cc_45 VNB N_A_63_65#_c_787_n 0.00199231f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.21
cc_46 VNB N_A_63_65#_c_788_n 0.00166051f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.21
cc_47 VNB N_A_63_65#_c_789_n 0.00465116f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_63_65#_c_790_n 0.00318981f $X=-0.19 $Y=-0.245 $X2=0.625 $Y2=1.44
cc_49 VNB N_VGND_c_838_n 0.00228974f $X=-0.19 $Y=-0.245 $X2=1.515 $Y2=1.275
cc_50 VNB N_VGND_c_839_n 0.00228974f $X=-0.19 $Y=-0.245 $X2=1.645 $Y2=2.465
cc_51 VNB N_VGND_c_840_n 3.99129e-19 $X=-0.19 $Y=-0.245 $X2=1.945 $Y2=0.745
cc_52 VNB N_VGND_c_841_n 3.99129e-19 $X=-0.19 $Y=-0.245 $X2=2.075 $Y2=2.465
cc_53 VNB N_VGND_c_842_n 0.0143206f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.21
cc_54 VNB N_VGND_c_843_n 0.106216f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_844_n 0.0129398f $X=-0.19 $Y=-0.245 $X2=0.625 $Y2=1.44
cc_56 VNB N_VGND_c_845_n 0.0153759f $X=-0.19 $Y=-0.245 $X2=1.215 $Y2=1.44
cc_57 VNB N_VGND_c_846_n 0.419675f $X=-0.19 $Y=-0.245 $X2=1.305 $Y2=1.44
cc_58 VNB N_VGND_c_847_n 0.0274581f $X=-0.19 $Y=-0.245 $X2=1.515 $Y2=1.44
cc_59 VNB N_VGND_c_848_n 0.00549308f $X=-0.19 $Y=-0.245 $X2=1.645 $Y2=1.44
cc_60 VNB N_VGND_c_849_n 0.00436918f $X=-0.19 $Y=-0.245 $X2=1.985 $Y2=1.44
cc_61 VNB N_VGND_c_850_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_A_867_47#_c_935_n 0.00317776f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_A_867_47#_c_936_n 0.016323f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_A_867_47#_c_937_n 0.0307328f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.21
cc_65 VNB N_A_867_47#_c_938_n 0.00218452f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VPB N_B2_M1006_g 0.026977f $X=-0.19 $Y=1.655 $X2=0.785 $Y2=2.465
cc_67 VPB N_B2_M1015_g 0.0186909f $X=-0.19 $Y=1.655 $X2=1.215 $Y2=2.465
cc_68 VPB N_B2_M1023_g 0.0186909f $X=-0.19 $Y=1.655 $X2=1.645 $Y2=2.465
cc_69 VPB N_B2_M1027_g 0.0188123f $X=-0.19 $Y=1.655 $X2=2.075 $Y2=2.465
cc_70 VPB N_B1_M1000_g 0.018308f $X=-0.19 $Y=1.655 $X2=0.785 $Y2=1.605
cc_71 VPB N_B1_M1008_g 0.0196366f $X=-0.19 $Y=1.655 $X2=1.215 $Y2=1.605
cc_72 VPB N_B1_M1016_g 0.0196366f $X=-0.19 $Y=1.655 $X2=1.645 $Y2=1.605
cc_73 VPB N_B1_M1019_g 0.0207315f $X=-0.19 $Y=1.655 $X2=2.075 $Y2=1.605
cc_74 VPB N_A1_M1013_g 0.0203056f $X=-0.19 $Y=1.655 $X2=0.655 $Y2=1.275
cc_75 VPB N_A1_M1017_g 0.018914f $X=-0.19 $Y=1.655 $X2=1.085 $Y2=1.275
cc_76 VPB N_A1_M1026_g 0.0194643f $X=-0.19 $Y=1.655 $X2=1.515 $Y2=1.275
cc_77 VPB N_A1_M1030_g 0.0198783f $X=-0.19 $Y=1.655 $X2=1.945 $Y2=1.275
cc_78 VPB N_A2_c_387_n 0.0162157f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_79 VPB N_A2_c_388_n 0.0159926f $X=-0.19 $Y=1.655 $X2=0.785 $Y2=2.465
cc_80 VPB N_A2_c_389_n 0.0157304f $X=-0.19 $Y=1.655 $X2=1.215 $Y2=2.465
cc_81 VPB N_A2_c_390_n 0.0211356f $X=-0.19 $Y=1.655 $X2=1.645 $Y2=2.465
cc_82 VPB A2 0.0182088f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_83 VPB N_A2_c_386_n 0.0303932f $X=-0.19 $Y=1.655 $X2=0.965 $Y2=1.44
cc_84 VPB N_A_89_367#_c_453_n 0.00746637f $X=-0.19 $Y=1.655 $X2=2.075 $Y2=2.465
cc_85 VPB N_A_89_367#_c_454_n 0.0427103f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_86 VPB N_A_89_367#_c_455_n 0.00576419f $X=-0.19 $Y=1.655 $X2=1.985 $Y2=1.44
cc_87 VPB N_A_89_367#_c_456_n 0.0035115f $X=-0.19 $Y=1.655 $X2=1.985 $Y2=1.44
cc_88 VPB N_A_89_367#_c_457_n 0.00374959f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=1.367
cc_89 VPB N_A_89_367#_c_458_n 0.0027807f $X=-0.19 $Y=1.655 $X2=0.965 $Y2=1.367
cc_90 VPB N_A_89_367#_c_459_n 0.0075508f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_91 VPB N_A_89_367#_c_460_n 0.0369431f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_92 VPB N_A_89_367#_c_461_n 0.00187503f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_93 VPB N_Y_c_564_n 0.0022809f $X=-0.19 $Y=1.655 $X2=2.075 $Y2=2.465
cc_94 VPB N_Y_c_565_n 0.00233203f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_95 VPB N_Y_c_566_n 0.00551076f $X=-0.19 $Y=1.655 $X2=2.075 $Y2=1.21
cc_96 VPB N_Y_c_562_n 6.05819e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_97 VPB N_Y_c_568_n 0.00508701f $X=-0.19 $Y=1.655 $X2=0.625 $Y2=1.44
cc_98 VPB N_Y_c_569_n 0.00233203f $X=-0.19 $Y=1.655 $X2=1.085 $Y2=1.44
cc_99 VPB N_Y_c_570_n 0.00267664f $X=-0.19 $Y=1.655 $X2=1.215 $Y2=1.44
cc_100 VPB N_VPWR_c_677_n 3.99129e-19 $X=-0.19 $Y=1.655 $X2=1.215 $Y2=2.465
cc_101 VPB N_VPWR_c_678_n 0.002101f $X=-0.19 $Y=1.655 $X2=1.645 $Y2=2.465
cc_102 VPB N_VPWR_c_679_n 3.16879e-19 $X=-0.19 $Y=1.655 $X2=2.075 $Y2=1.605
cc_103 VPB N_VPWR_c_680_n 3.99129e-19 $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_104 VPB N_VPWR_c_681_n 0.0149824f $X=-0.19 $Y=1.655 $X2=1.595 $Y2=1.21
cc_105 VPB N_VPWR_c_682_n 0.00436868f $X=-0.19 $Y=1.655 $X2=2.075 $Y2=1.21
cc_106 VPB N_VPWR_c_683_n 0.0129398f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_107 VPB N_VPWR_c_684_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_108 VPB N_VPWR_c_685_n 0.105445f $X=-0.19 $Y=1.655 $X2=0.625 $Y2=1.44
cc_109 VPB N_VPWR_c_686_n 0.0129398f $X=-0.19 $Y=1.655 $X2=1.085 $Y2=1.44
cc_110 VPB N_VPWR_c_687_n 0.0223767f $X=-0.19 $Y=1.655 $X2=2.075 $Y2=1.44
cc_111 VPB N_VPWR_c_676_n 0.0674407f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_112 VPB N_VPWR_c_689_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_113 VPB N_VPWR_c_690_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_114 N_B2_c_120_n N_B1_c_201_n 0.0224946f $X=1.945 $Y=1.275 $X2=-0.19
+ $Y2=-0.245
cc_115 B2 N_B1_c_201_n 0.0016646f $X=2.075 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_116 N_B2_M1027_g N_B1_M1000_g 0.0161492f $X=2.075 $Y=2.465 $X2=0 $Y2=0
cc_117 B2 N_B1_c_210_n 3.96827e-19 $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_118 N_B2_c_124_n N_B1_c_210_n 0.0260522f $X=2.075 $Y=1.44 $X2=0 $Y2=0
cc_119 N_B2_M1006_g N_A_89_367#_c_454_n 0.0029331f $X=0.785 $Y=2.465 $X2=0 $Y2=0
cc_120 B2 N_A_89_367#_c_454_n 0.0141878f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_121 N_B2_c_123_n N_A_89_367#_c_454_n 0.00644127f $X=0.625 $Y=1.44 $X2=0 $Y2=0
cc_122 N_B2_M1006_g N_A_89_367#_c_465_n 0.0115031f $X=0.785 $Y=2.465 $X2=0 $Y2=0
cc_123 N_B2_M1015_g N_A_89_367#_c_465_n 0.0115031f $X=1.215 $Y=2.465 $X2=0 $Y2=0
cc_124 N_B2_M1023_g N_A_89_367#_c_467_n 0.0115031f $X=1.645 $Y=2.465 $X2=0 $Y2=0
cc_125 N_B2_M1027_g N_A_89_367#_c_467_n 0.0115031f $X=2.075 $Y=2.465 $X2=0 $Y2=0
cc_126 N_B2_M1006_g N_Y_c_571_n 0.0123079f $X=0.785 $Y=2.465 $X2=0 $Y2=0
cc_127 N_B2_M1015_g N_Y_c_571_n 0.0130783f $X=1.215 $Y=2.465 $X2=0 $Y2=0
cc_128 N_B2_M1023_g N_Y_c_571_n 6.30056e-19 $X=1.645 $Y=2.465 $X2=0 $Y2=0
cc_129 N_B2_M1015_g N_Y_c_564_n 0.0112007f $X=1.215 $Y=2.465 $X2=0 $Y2=0
cc_130 N_B2_M1023_g N_Y_c_564_n 0.0112007f $X=1.645 $Y=2.465 $X2=0 $Y2=0
cc_131 B2 N_Y_c_564_n 0.0370126f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_132 N_B2_c_124_n N_Y_c_564_n 0.00287416f $X=2.075 $Y=1.44 $X2=0 $Y2=0
cc_133 N_B2_M1006_g N_Y_c_565_n 0.00811014f $X=0.785 $Y=2.465 $X2=0 $Y2=0
cc_134 N_B2_M1015_g N_Y_c_565_n 0.00231052f $X=1.215 $Y=2.465 $X2=0 $Y2=0
cc_135 B2 N_Y_c_565_n 0.0263482f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_136 N_B2_c_124_n N_Y_c_565_n 0.00298081f $X=2.075 $Y=1.44 $X2=0 $Y2=0
cc_137 N_B2_M1015_g N_Y_c_582_n 6.30056e-19 $X=1.215 $Y=2.465 $X2=0 $Y2=0
cc_138 N_B2_M1023_g N_Y_c_582_n 0.0130783f $X=1.645 $Y=2.465 $X2=0 $Y2=0
cc_139 N_B2_M1027_g N_Y_c_582_n 0.0130783f $X=2.075 $Y=2.465 $X2=0 $Y2=0
cc_140 N_B2_M1027_g N_Y_c_566_n 0.0111542f $X=2.075 $Y=2.465 $X2=0 $Y2=0
cc_141 B2 N_Y_c_566_n 0.0156705f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_142 B2 N_Y_c_562_n 0.0245335f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_143 N_B2_c_124_n N_Y_c_562_n 0.00406488f $X=2.075 $Y=1.44 $X2=0 $Y2=0
cc_144 N_B2_M1027_g N_Y_c_589_n 6.30056e-19 $X=2.075 $Y=2.465 $X2=0 $Y2=0
cc_145 N_B2_M1023_g N_Y_c_569_n 0.00231052f $X=1.645 $Y=2.465 $X2=0 $Y2=0
cc_146 N_B2_M1027_g N_Y_c_569_n 0.00231052f $X=2.075 $Y=2.465 $X2=0 $Y2=0
cc_147 B2 N_Y_c_569_n 0.0263482f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_148 N_B2_c_124_n N_Y_c_569_n 0.00298081f $X=2.075 $Y=1.44 $X2=0 $Y2=0
cc_149 N_B2_c_120_n N_Y_c_594_n 8.47781e-19 $X=1.945 $Y=1.275 $X2=0 $Y2=0
cc_150 N_B2_M1006_g N_VPWR_c_685_n 0.00357877f $X=0.785 $Y=2.465 $X2=0 $Y2=0
cc_151 N_B2_M1015_g N_VPWR_c_685_n 0.00357877f $X=1.215 $Y=2.465 $X2=0 $Y2=0
cc_152 N_B2_M1023_g N_VPWR_c_685_n 0.00357877f $X=1.645 $Y=2.465 $X2=0 $Y2=0
cc_153 N_B2_M1027_g N_VPWR_c_685_n 0.00357877f $X=2.075 $Y=2.465 $X2=0 $Y2=0
cc_154 N_B2_M1006_g N_VPWR_c_676_n 0.00647412f $X=0.785 $Y=2.465 $X2=0 $Y2=0
cc_155 N_B2_M1015_g N_VPWR_c_676_n 0.0053512f $X=1.215 $Y=2.465 $X2=0 $Y2=0
cc_156 N_B2_M1023_g N_VPWR_c_676_n 0.0053512f $X=1.645 $Y=2.465 $X2=0 $Y2=0
cc_157 N_B2_M1027_g N_VPWR_c_676_n 0.00537654f $X=2.075 $Y=2.465 $X2=0 $Y2=0
cc_158 N_B2_c_114_n N_A_63_65#_c_784_n 3.18679e-19 $X=0.655 $Y=1.275 $X2=0 $Y2=0
cc_159 N_B2_c_114_n N_A_63_65#_c_792_n 0.0120408f $X=0.655 $Y=1.275 $X2=0 $Y2=0
cc_160 N_B2_c_116_n N_A_63_65#_c_792_n 0.0120955f $X=1.085 $Y=1.275 $X2=0 $Y2=0
cc_161 B2 N_A_63_65#_c_792_n 0.0426015f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_162 N_B2_c_124_n N_A_63_65#_c_792_n 5.84859e-19 $X=2.075 $Y=1.44 $X2=0 $Y2=0
cc_163 B2 N_A_63_65#_c_785_n 0.0219949f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_164 N_B2_c_123_n N_A_63_65#_c_785_n 0.00170661f $X=0.625 $Y=1.44 $X2=0 $Y2=0
cc_165 N_B2_c_118_n N_A_63_65#_c_798_n 0.0120489f $X=1.515 $Y=1.275 $X2=0 $Y2=0
cc_166 N_B2_c_120_n N_A_63_65#_c_798_n 0.0120955f $X=1.945 $Y=1.275 $X2=0 $Y2=0
cc_167 B2 N_A_63_65#_c_798_n 0.0576144f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_168 N_B2_c_124_n N_A_63_65#_c_798_n 0.00111454f $X=2.075 $Y=1.44 $X2=0 $Y2=0
cc_169 N_B2_c_120_n N_A_63_65#_c_787_n 6.28789e-19 $X=1.945 $Y=1.275 $X2=0 $Y2=0
cc_170 B2 N_A_63_65#_c_803_n 0.0153383f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_171 N_B2_c_124_n N_A_63_65#_c_803_n 6.61019e-19 $X=2.075 $Y=1.44 $X2=0 $Y2=0
cc_172 N_B2_c_114_n N_VGND_c_838_n 0.0112436f $X=0.655 $Y=1.275 $X2=0 $Y2=0
cc_173 N_B2_c_116_n N_VGND_c_838_n 0.00879717f $X=1.085 $Y=1.275 $X2=0 $Y2=0
cc_174 N_B2_c_118_n N_VGND_c_838_n 4.78085e-19 $X=1.515 $Y=1.275 $X2=0 $Y2=0
cc_175 N_B2_c_116_n N_VGND_c_839_n 4.78085e-19 $X=1.085 $Y=1.275 $X2=0 $Y2=0
cc_176 N_B2_c_118_n N_VGND_c_839_n 0.00879717f $X=1.515 $Y=1.275 $X2=0 $Y2=0
cc_177 N_B2_c_120_n N_VGND_c_839_n 0.00882039f $X=1.945 $Y=1.275 $X2=0 $Y2=0
cc_178 N_B2_c_116_n N_VGND_c_842_n 0.00414769f $X=1.085 $Y=1.275 $X2=0 $Y2=0
cc_179 N_B2_c_118_n N_VGND_c_842_n 0.00414769f $X=1.515 $Y=1.275 $X2=0 $Y2=0
cc_180 N_B2_c_120_n N_VGND_c_843_n 0.00414769f $X=1.945 $Y=1.275 $X2=0 $Y2=0
cc_181 N_B2_c_114_n N_VGND_c_846_n 0.00828433f $X=0.655 $Y=1.275 $X2=0 $Y2=0
cc_182 N_B2_c_116_n N_VGND_c_846_n 0.00787505f $X=1.085 $Y=1.275 $X2=0 $Y2=0
cc_183 N_B2_c_118_n N_VGND_c_846_n 0.00787505f $X=1.515 $Y=1.275 $X2=0 $Y2=0
cc_184 N_B2_c_120_n N_VGND_c_846_n 0.0079379f $X=1.945 $Y=1.275 $X2=0 $Y2=0
cc_185 N_B2_c_114_n N_VGND_c_847_n 0.00414769f $X=0.655 $Y=1.275 $X2=0 $Y2=0
cc_186 N_B1_M1019_g N_A1_M1013_g 0.0152896f $X=3.875 $Y=2.465 $X2=0 $Y2=0
cc_187 B1 N_A1_M1013_g 0.00272194f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_188 B1 N_A1_M1017_g 2.5943e-19 $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_189 B1 A1 0.0145345f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_190 N_B1_c_207_n N_A1_c_305_n 0.00191622f $X=3.725 $Y=1.275 $X2=0 $Y2=0
cc_191 B1 N_A1_c_305_n 0.0234084f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_192 N_B1_c_210_n N_A1_c_305_n 0.0223074f $X=3.875 $Y=1.44 $X2=0 $Y2=0
cc_193 N_B1_M1000_g N_A_89_367#_c_469_n 0.0115031f $X=2.505 $Y=2.465 $X2=0 $Y2=0
cc_194 N_B1_M1008_g N_A_89_367#_c_469_n 0.0115031f $X=2.935 $Y=2.465 $X2=0 $Y2=0
cc_195 N_B1_M1016_g N_A_89_367#_c_471_n 0.0115031f $X=3.445 $Y=2.465 $X2=0 $Y2=0
cc_196 N_B1_M1019_g N_A_89_367#_c_471_n 0.0115031f $X=3.875 $Y=2.465 $X2=0 $Y2=0
cc_197 B1 N_A_89_367#_c_455_n 0.0214612f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_198 N_B1_M1019_g N_A_89_367#_c_456_n 7.62722e-19 $X=3.875 $Y=2.465 $X2=0
+ $Y2=0
cc_199 B1 N_A_89_367#_c_456_n 0.0204821f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_200 N_B1_c_210_n N_A_89_367#_c_456_n 0.00323402f $X=3.875 $Y=1.44 $X2=0 $Y2=0
cc_201 N_B1_M1000_g N_Y_c_582_n 6.30056e-19 $X=2.505 $Y=2.465 $X2=0 $Y2=0
cc_202 N_B1_c_210_n N_Y_c_566_n 0.00238284f $X=3.875 $Y=1.44 $X2=0 $Y2=0
cc_203 N_B1_c_201_n N_Y_c_562_n 0.00329464f $X=2.435 $Y=1.275 $X2=0 $Y2=0
cc_204 N_B1_M1000_g N_Y_c_562_n 0.00242187f $X=2.505 $Y=2.465 $X2=0 $Y2=0
cc_205 N_B1_c_203_n N_Y_c_562_n 7.89004e-19 $X=2.865 $Y=1.275 $X2=0 $Y2=0
cc_206 N_B1_M1008_g N_Y_c_562_n 9.19529e-19 $X=2.935 $Y=2.465 $X2=0 $Y2=0
cc_207 N_B1_c_210_n N_Y_c_562_n 0.0142957f $X=3.875 $Y=1.44 $X2=0 $Y2=0
cc_208 N_B1_c_211_n N_Y_c_562_n 0.0185536f $X=3.142 $Y=1.367 $X2=0 $Y2=0
cc_209 N_B1_M1000_g N_Y_c_589_n 0.0130783f $X=2.505 $Y=2.465 $X2=0 $Y2=0
cc_210 N_B1_M1008_g N_Y_c_589_n 0.0134529f $X=2.935 $Y=2.465 $X2=0 $Y2=0
cc_211 N_B1_M1016_g N_Y_c_589_n 6.11257e-19 $X=3.445 $Y=2.465 $X2=0 $Y2=0
cc_212 N_B1_M1008_g N_Y_c_568_n 0.0116393f $X=2.935 $Y=2.465 $X2=0 $Y2=0
cc_213 N_B1_M1016_g N_Y_c_568_n 0.0139549f $X=3.445 $Y=2.465 $X2=0 $Y2=0
cc_214 N_B1_M1019_g N_Y_c_568_n 0.00422635f $X=3.875 $Y=2.465 $X2=0 $Y2=0
cc_215 B1 N_Y_c_568_n 0.0511308f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_216 N_B1_c_210_n N_Y_c_568_n 0.00802618f $X=3.875 $Y=1.44 $X2=0 $Y2=0
cc_217 N_B1_c_211_n N_Y_c_568_n 0.0176985f $X=3.142 $Y=1.367 $X2=0 $Y2=0
cc_218 N_B1_M1008_g N_Y_c_612_n 6.11257e-19 $X=2.935 $Y=2.465 $X2=0 $Y2=0
cc_219 N_B1_M1016_g N_Y_c_612_n 0.0134529f $X=3.445 $Y=2.465 $X2=0 $Y2=0
cc_220 N_B1_M1019_g N_Y_c_612_n 0.0119685f $X=3.875 $Y=2.465 $X2=0 $Y2=0
cc_221 N_B1_M1000_g N_Y_c_570_n 0.012411f $X=2.505 $Y=2.465 $X2=0 $Y2=0
cc_222 N_B1_M1008_g N_Y_c_570_n 0.00230943f $X=2.935 $Y=2.465 $X2=0 $Y2=0
cc_223 N_B1_c_210_n N_Y_c_570_n 0.0034671f $X=3.875 $Y=1.44 $X2=0 $Y2=0
cc_224 N_B1_c_211_n N_Y_c_570_n 0.00843256f $X=3.142 $Y=1.367 $X2=0 $Y2=0
cc_225 N_B1_c_203_n N_Y_c_563_n 0.0117042f $X=2.865 $Y=1.275 $X2=0 $Y2=0
cc_226 N_B1_c_205_n N_Y_c_563_n 0.00997563f $X=3.295 $Y=1.275 $X2=0 $Y2=0
cc_227 N_B1_c_207_n N_Y_c_563_n 0.0126842f $X=3.725 $Y=1.275 $X2=0 $Y2=0
cc_228 B1 N_Y_c_563_n 0.105185f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_229 N_B1_c_210_n N_Y_c_563_n 0.00303546f $X=3.875 $Y=1.44 $X2=0 $Y2=0
cc_230 N_B1_c_211_n N_Y_c_563_n 0.0182793f $X=3.142 $Y=1.367 $X2=0 $Y2=0
cc_231 N_B1_c_201_n N_Y_c_594_n 0.0101064f $X=2.435 $Y=1.275 $X2=0 $Y2=0
cc_232 N_B1_c_203_n N_Y_c_594_n 0.00760513f $X=2.865 $Y=1.275 $X2=0 $Y2=0
cc_233 N_B1_c_205_n N_Y_c_594_n 0.00143575f $X=3.295 $Y=1.275 $X2=0 $Y2=0
cc_234 N_B1_c_210_n N_Y_c_594_n 0.0032772f $X=3.875 $Y=1.44 $X2=0 $Y2=0
cc_235 N_B1_c_211_n N_Y_c_594_n 0.00192124f $X=3.142 $Y=1.367 $X2=0 $Y2=0
cc_236 N_B1_M1019_g N_VPWR_c_677_n 9.44406e-19 $X=3.875 $Y=2.465 $X2=0 $Y2=0
cc_237 N_B1_M1000_g N_VPWR_c_685_n 0.00357877f $X=2.505 $Y=2.465 $X2=0 $Y2=0
cc_238 N_B1_M1008_g N_VPWR_c_685_n 0.00357877f $X=2.935 $Y=2.465 $X2=0 $Y2=0
cc_239 N_B1_M1016_g N_VPWR_c_685_n 0.00357877f $X=3.445 $Y=2.465 $X2=0 $Y2=0
cc_240 N_B1_M1019_g N_VPWR_c_685_n 0.00357877f $X=3.875 $Y=2.465 $X2=0 $Y2=0
cc_241 N_B1_M1000_g N_VPWR_c_676_n 0.00537654f $X=2.505 $Y=2.465 $X2=0 $Y2=0
cc_242 N_B1_M1008_g N_VPWR_c_676_n 0.00554494f $X=2.935 $Y=2.465 $X2=0 $Y2=0
cc_243 N_B1_M1016_g N_VPWR_c_676_n 0.00554494f $X=3.445 $Y=2.465 $X2=0 $Y2=0
cc_244 N_B1_M1019_g N_VPWR_c_676_n 0.00560871f $X=3.875 $Y=2.465 $X2=0 $Y2=0
cc_245 N_B1_c_201_n N_A_63_65#_c_798_n 0.00136247f $X=2.435 $Y=1.275 $X2=0 $Y2=0
cc_246 N_B1_c_201_n N_A_63_65#_c_806_n 0.00583424f $X=2.435 $Y=1.275 $X2=0 $Y2=0
cc_247 N_B1_c_205_n N_A_63_65#_c_788_n 0.0136567f $X=3.295 $Y=1.275 $X2=0 $Y2=0
cc_248 N_B1_c_207_n N_A_63_65#_c_789_n 0.014198f $X=3.725 $Y=1.275 $X2=0 $Y2=0
cc_249 N_B1_c_201_n N_A_63_65#_c_790_n 0.0113519f $X=2.435 $Y=1.275 $X2=0 $Y2=0
cc_250 N_B1_c_203_n N_A_63_65#_c_790_n 0.00913467f $X=2.865 $Y=1.275 $X2=0 $Y2=0
cc_251 N_B1_c_201_n N_VGND_c_839_n 5.93272e-19 $X=2.435 $Y=1.275 $X2=0 $Y2=0
cc_252 N_B1_c_201_n N_VGND_c_843_n 0.00302501f $X=2.435 $Y=1.275 $X2=0 $Y2=0
cc_253 N_B1_c_203_n N_VGND_c_843_n 0.00302501f $X=2.865 $Y=1.275 $X2=0 $Y2=0
cc_254 N_B1_c_205_n N_VGND_c_843_n 0.00302501f $X=3.295 $Y=1.275 $X2=0 $Y2=0
cc_255 N_B1_c_207_n N_VGND_c_843_n 0.00302501f $X=3.725 $Y=1.275 $X2=0 $Y2=0
cc_256 N_B1_c_201_n N_VGND_c_846_n 0.00440956f $X=2.435 $Y=1.275 $X2=0 $Y2=0
cc_257 N_B1_c_203_n N_VGND_c_846_n 0.00433762f $X=2.865 $Y=1.275 $X2=0 $Y2=0
cc_258 N_B1_c_205_n N_VGND_c_846_n 0.00434671f $X=3.295 $Y=1.275 $X2=0 $Y2=0
cc_259 N_B1_c_207_n N_VGND_c_846_n 0.0048466f $X=3.725 $Y=1.275 $X2=0 $Y2=0
cc_260 N_B1_c_207_n N_A_867_47#_c_935_n 7.06902e-19 $X=3.725 $Y=1.275 $X2=0
+ $Y2=0
cc_261 N_A1_c_303_n N_A2_M1002_g 0.0217853f $X=5.965 $Y=1.185 $X2=0 $Y2=0
cc_262 A1 N_A2_M1002_g 0.00639041f $X=6.395 $Y=1.21 $X2=0 $Y2=0
cc_263 N_A1_c_305_n N_A2_M1002_g 0.00600972f $X=5.745 $Y=1.35 $X2=0 $Y2=0
cc_264 A1 N_A2_M1012_g 0.00283029f $X=6.395 $Y=1.21 $X2=0 $Y2=0
cc_265 A1 A2 6.77207e-19 $X=6.395 $Y=1.21 $X2=0 $Y2=0
cc_266 N_A1_M1030_g N_A2_c_386_n 0.0271293f $X=5.745 $Y=2.465 $X2=0 $Y2=0
cc_267 A1 N_A2_c_386_n 0.0211692f $X=6.395 $Y=1.21 $X2=0 $Y2=0
cc_268 N_A1_M1013_g N_A_89_367#_c_455_n 0.013669f $X=4.41 $Y=2.465 $X2=0 $Y2=0
cc_269 N_A1_M1017_g N_A_89_367#_c_455_n 0.0168426f $X=4.84 $Y=2.465 $X2=0 $Y2=0
cc_270 A1 N_A_89_367#_c_455_n 0.00349003f $X=6.395 $Y=1.21 $X2=0 $Y2=0
cc_271 N_A1_c_305_n N_A_89_367#_c_455_n 0.00160418f $X=5.745 $Y=1.35 $X2=0 $Y2=0
cc_272 N_A1_M1026_g N_A_89_367#_c_457_n 0.0142598f $X=5.27 $Y=2.465 $X2=0 $Y2=0
cc_273 N_A1_M1030_g N_A_89_367#_c_457_n 0.0140916f $X=5.745 $Y=2.465 $X2=0 $Y2=0
cc_274 A1 N_A_89_367#_c_457_n 0.0293559f $X=6.395 $Y=1.21 $X2=0 $Y2=0
cc_275 N_A1_c_305_n N_A_89_367#_c_457_n 0.00374251f $X=5.745 $Y=1.35 $X2=0 $Y2=0
cc_276 N_A1_M1030_g N_A_89_367#_c_458_n 7.07765e-19 $X=5.745 $Y=2.465 $X2=0
+ $Y2=0
cc_277 A1 N_A_89_367#_c_458_n 0.0121906f $X=6.395 $Y=1.21 $X2=0 $Y2=0
cc_278 N_A1_c_305_n N_A_89_367#_c_458_n 0.00280242f $X=5.745 $Y=1.35 $X2=0 $Y2=0
cc_279 A1 N_A_89_367#_c_488_n 0.0143391f $X=6.395 $Y=1.21 $X2=0 $Y2=0
cc_280 A1 N_A_89_367#_c_461_n 0.0097664f $X=6.395 $Y=1.21 $X2=0 $Y2=0
cc_281 N_A1_c_305_n N_A_89_367#_c_461_n 0.00271666f $X=5.745 $Y=1.35 $X2=0 $Y2=0
cc_282 N_A1_M1013_g N_Y_c_568_n 2.94909e-19 $X=4.41 $Y=2.465 $X2=0 $Y2=0
cc_283 A1 N_Y_c_631_n 0.0137759f $X=6.395 $Y=1.21 $X2=0 $Y2=0
cc_284 N_A1_c_305_n N_Y_c_631_n 0.00275656f $X=5.745 $Y=1.35 $X2=0 $Y2=0
cc_285 N_A1_c_297_n N_Y_c_563_n 0.0165301f $X=4.675 $Y=1.185 $X2=0 $Y2=0
cc_286 N_A1_c_299_n N_Y_c_563_n 0.0105327f $X=5.105 $Y=1.185 $X2=0 $Y2=0
cc_287 N_A1_c_301_n N_Y_c_563_n 0.0105945f $X=5.535 $Y=1.185 $X2=0 $Y2=0
cc_288 A1 N_Y_c_563_n 0.047421f $X=6.395 $Y=1.21 $X2=0 $Y2=0
cc_289 N_A1_c_305_n N_Y_c_563_n 0.0131103f $X=5.745 $Y=1.35 $X2=0 $Y2=0
cc_290 N_A1_M1013_g N_VPWR_c_677_n 0.0156274f $X=4.41 $Y=2.465 $X2=0 $Y2=0
cc_291 N_A1_M1017_g N_VPWR_c_677_n 0.0142791f $X=4.84 $Y=2.465 $X2=0 $Y2=0
cc_292 N_A1_M1026_g N_VPWR_c_677_n 7.27171e-19 $X=5.27 $Y=2.465 $X2=0 $Y2=0
cc_293 N_A1_M1017_g N_VPWR_c_678_n 7.27171e-19 $X=4.84 $Y=2.465 $X2=0 $Y2=0
cc_294 N_A1_M1026_g N_VPWR_c_678_n 0.0142171f $X=5.27 $Y=2.465 $X2=0 $Y2=0
cc_295 N_A1_M1030_g N_VPWR_c_678_n 0.0016858f $X=5.745 $Y=2.465 $X2=0 $Y2=0
cc_296 N_A1_M1030_g N_VPWR_c_679_n 6.95886e-19 $X=5.745 $Y=2.465 $X2=0 $Y2=0
cc_297 N_A1_M1030_g N_VPWR_c_681_n 0.00585385f $X=5.745 $Y=2.465 $X2=0 $Y2=0
cc_298 N_A1_M1013_g N_VPWR_c_685_n 0.00486043f $X=4.41 $Y=2.465 $X2=0 $Y2=0
cc_299 N_A1_M1017_g N_VPWR_c_686_n 0.00486043f $X=4.84 $Y=2.465 $X2=0 $Y2=0
cc_300 N_A1_M1026_g N_VPWR_c_686_n 0.00486043f $X=5.27 $Y=2.465 $X2=0 $Y2=0
cc_301 N_A1_M1013_g N_VPWR_c_676_n 0.00850478f $X=4.41 $Y=2.465 $X2=0 $Y2=0
cc_302 N_A1_M1017_g N_VPWR_c_676_n 0.00824727f $X=4.84 $Y=2.465 $X2=0 $Y2=0
cc_303 N_A1_M1026_g N_VPWR_c_676_n 0.00824727f $X=5.27 $Y=2.465 $X2=0 $Y2=0
cc_304 N_A1_M1030_g N_VPWR_c_676_n 0.0106877f $X=5.745 $Y=2.465 $X2=0 $Y2=0
cc_305 N_A1_c_297_n N_A_63_65#_c_789_n 0.00244901f $X=4.675 $Y=1.185 $X2=0 $Y2=0
cc_306 N_A1_c_303_n N_VGND_c_840_n 0.00116114f $X=5.965 $Y=1.185 $X2=0 $Y2=0
cc_307 N_A1_c_297_n N_VGND_c_843_n 0.00362032f $X=4.675 $Y=1.185 $X2=0 $Y2=0
cc_308 N_A1_c_299_n N_VGND_c_843_n 0.00362032f $X=5.105 $Y=1.185 $X2=0 $Y2=0
cc_309 N_A1_c_301_n N_VGND_c_843_n 0.00362032f $X=5.535 $Y=1.185 $X2=0 $Y2=0
cc_310 N_A1_c_303_n N_VGND_c_843_n 0.00361998f $X=5.965 $Y=1.185 $X2=0 $Y2=0
cc_311 N_A1_c_297_n N_VGND_c_846_n 0.00665528f $X=4.675 $Y=1.185 $X2=0 $Y2=0
cc_312 N_A1_c_299_n N_VGND_c_846_n 0.00535559f $X=5.105 $Y=1.185 $X2=0 $Y2=0
cc_313 N_A1_c_301_n N_VGND_c_846_n 0.00535559f $X=5.535 $Y=1.185 $X2=0 $Y2=0
cc_314 N_A1_c_303_n N_VGND_c_846_n 0.00544446f $X=5.965 $Y=1.185 $X2=0 $Y2=0
cc_315 N_A1_c_297_n N_A_867_47#_c_935_n 0.0106283f $X=4.675 $Y=1.185 $X2=0 $Y2=0
cc_316 N_A1_c_299_n N_A_867_47#_c_935_n 0.0106283f $X=5.105 $Y=1.185 $X2=0 $Y2=0
cc_317 N_A1_c_301_n N_A_867_47#_c_935_n 0.0105595f $X=5.535 $Y=1.185 $X2=0 $Y2=0
cc_318 N_A1_c_303_n N_A_867_47#_c_935_n 0.0127727f $X=5.965 $Y=1.185 $X2=0 $Y2=0
cc_319 N_A1_c_303_n N_A_867_47#_c_944_n 7.92301e-19 $X=5.965 $Y=1.185 $X2=0
+ $Y2=0
cc_320 N_A1_c_301_n N_A_867_47#_c_945_n 7.86683e-19 $X=5.535 $Y=1.185 $X2=0
+ $Y2=0
cc_321 N_A1_c_303_n N_A_867_47#_c_945_n 0.00726126f $X=5.965 $Y=1.185 $X2=0
+ $Y2=0
cc_322 A1 N_A_867_47#_c_945_n 0.0186215f $X=6.395 $Y=1.21 $X2=0 $Y2=0
cc_323 A1 N_A_867_47#_c_948_n 0.0188602f $X=6.395 $Y=1.21 $X2=0 $Y2=0
cc_324 A1 N_A_867_47#_c_938_n 0.00256446f $X=6.395 $Y=1.21 $X2=0 $Y2=0
cc_325 N_A2_c_387_n N_A_89_367#_c_458_n 0.00250406f $X=6.175 $Y=1.725 $X2=0
+ $Y2=0
cc_326 N_A2_c_387_n N_A_89_367#_c_488_n 0.0133278f $X=6.175 $Y=1.725 $X2=0 $Y2=0
cc_327 N_A2_c_388_n N_A_89_367#_c_488_n 0.0156345f $X=6.605 $Y=1.725 $X2=0 $Y2=0
cc_328 N_A2_c_386_n N_A_89_367#_c_488_n 0.00285278f $X=7.595 $Y=1.51 $X2=0 $Y2=0
cc_329 N_A2_c_389_n N_A_89_367#_c_495_n 0.0122595f $X=7.035 $Y=1.725 $X2=0 $Y2=0
cc_330 N_A2_c_390_n N_A_89_367#_c_495_n 0.0122595f $X=7.465 $Y=1.725 $X2=0 $Y2=0
cc_331 A2 N_A_89_367#_c_495_n 0.0428504f $X=7.835 $Y=1.58 $X2=0 $Y2=0
cc_332 N_A2_c_386_n N_A_89_367#_c_495_n 6.31497e-19 $X=7.595 $Y=1.51 $X2=0 $Y2=0
cc_333 A2 N_A_89_367#_c_459_n 0.0220964f $X=7.835 $Y=1.58 $X2=0 $Y2=0
cc_334 N_A2_c_386_n N_A_89_367#_c_459_n 0.00121256f $X=7.595 $Y=1.51 $X2=0 $Y2=0
cc_335 A2 N_A_89_367#_c_501_n 0.013781f $X=7.835 $Y=1.58 $X2=0 $Y2=0
cc_336 N_A2_c_386_n N_A_89_367#_c_501_n 7.1239e-19 $X=7.595 $Y=1.51 $X2=0 $Y2=0
cc_337 N_A2_c_387_n N_VPWR_c_679_n 0.0146603f $X=6.175 $Y=1.725 $X2=0 $Y2=0
cc_338 N_A2_c_388_n N_VPWR_c_679_n 0.0145573f $X=6.605 $Y=1.725 $X2=0 $Y2=0
cc_339 N_A2_c_389_n N_VPWR_c_679_n 6.77662e-19 $X=7.035 $Y=1.725 $X2=0 $Y2=0
cc_340 N_A2_c_388_n N_VPWR_c_680_n 6.77662e-19 $X=6.605 $Y=1.725 $X2=0 $Y2=0
cc_341 N_A2_c_389_n N_VPWR_c_680_n 0.0145573f $X=7.035 $Y=1.725 $X2=0 $Y2=0
cc_342 N_A2_c_390_n N_VPWR_c_680_n 0.0164416f $X=7.465 $Y=1.725 $X2=0 $Y2=0
cc_343 N_A2_c_387_n N_VPWR_c_681_n 0.00486043f $X=6.175 $Y=1.725 $X2=0 $Y2=0
cc_344 N_A2_c_388_n N_VPWR_c_683_n 0.00486043f $X=6.605 $Y=1.725 $X2=0 $Y2=0
cc_345 N_A2_c_389_n N_VPWR_c_683_n 0.00486043f $X=7.035 $Y=1.725 $X2=0 $Y2=0
cc_346 N_A2_c_390_n N_VPWR_c_687_n 0.00486043f $X=7.465 $Y=1.725 $X2=0 $Y2=0
cc_347 N_A2_c_387_n N_VPWR_c_676_n 0.0082726f $X=6.175 $Y=1.725 $X2=0 $Y2=0
cc_348 N_A2_c_388_n N_VPWR_c_676_n 0.00824727f $X=6.605 $Y=1.725 $X2=0 $Y2=0
cc_349 N_A2_c_389_n N_VPWR_c_676_n 0.00824727f $X=7.035 $Y=1.725 $X2=0 $Y2=0
cc_350 N_A2_c_390_n N_VPWR_c_676_n 0.00933203f $X=7.465 $Y=1.725 $X2=0 $Y2=0
cc_351 N_A2_M1002_g N_VGND_c_840_n 0.00981715f $X=6.395 $Y=0.655 $X2=0 $Y2=0
cc_352 N_A2_M1012_g N_VGND_c_840_n 0.00846696f $X=6.825 $Y=0.655 $X2=0 $Y2=0
cc_353 N_A2_M1014_g N_VGND_c_840_n 5.48939e-19 $X=7.255 $Y=0.655 $X2=0 $Y2=0
cc_354 N_A2_M1012_g N_VGND_c_841_n 5.97034e-19 $X=6.825 $Y=0.655 $X2=0 $Y2=0
cc_355 N_A2_M1014_g N_VGND_c_841_n 0.0110161f $X=7.255 $Y=0.655 $X2=0 $Y2=0
cc_356 N_A2_M1031_g N_VGND_c_841_n 0.012818f $X=7.685 $Y=0.655 $X2=0 $Y2=0
cc_357 N_A2_M1002_g N_VGND_c_843_n 0.00486043f $X=6.395 $Y=0.655 $X2=0 $Y2=0
cc_358 N_A2_M1012_g N_VGND_c_844_n 0.00486043f $X=6.825 $Y=0.655 $X2=0 $Y2=0
cc_359 N_A2_M1014_g N_VGND_c_844_n 0.00486043f $X=7.255 $Y=0.655 $X2=0 $Y2=0
cc_360 N_A2_M1031_g N_VGND_c_845_n 0.00486043f $X=7.685 $Y=0.655 $X2=0 $Y2=0
cc_361 N_A2_M1002_g N_VGND_c_846_n 0.00449474f $X=6.395 $Y=0.655 $X2=0 $Y2=0
cc_362 N_A2_M1012_g N_VGND_c_846_n 0.00438968f $X=6.825 $Y=0.655 $X2=0 $Y2=0
cc_363 N_A2_M1014_g N_VGND_c_846_n 0.00824727f $X=7.255 $Y=0.655 $X2=0 $Y2=0
cc_364 N_A2_M1031_g N_VGND_c_846_n 0.00917987f $X=7.685 $Y=0.655 $X2=0 $Y2=0
cc_365 N_A2_M1002_g N_A_867_47#_c_948_n 0.012136f $X=6.395 $Y=0.655 $X2=0 $Y2=0
cc_366 N_A2_M1012_g N_A_867_47#_c_948_n 0.011437f $X=6.825 $Y=0.655 $X2=0 $Y2=0
cc_367 A2 N_A_867_47#_c_948_n 0.00401948f $X=7.835 $Y=1.58 $X2=0 $Y2=0
cc_368 N_A2_c_386_n N_A_867_47#_c_948_n 0.0031072f $X=7.595 $Y=1.51 $X2=0 $Y2=0
cc_369 N_A2_M1014_g N_A_867_47#_c_936_n 0.0136772f $X=7.255 $Y=0.655 $X2=0 $Y2=0
cc_370 N_A2_M1031_g N_A_867_47#_c_936_n 0.0164369f $X=7.685 $Y=0.655 $X2=0 $Y2=0
cc_371 A2 N_A_867_47#_c_936_n 0.0675649f $X=7.835 $Y=1.58 $X2=0 $Y2=0
cc_372 N_A2_c_386_n N_A_867_47#_c_936_n 0.00290124f $X=7.595 $Y=1.51 $X2=0 $Y2=0
cc_373 N_A2_M1002_g N_A_867_47#_c_938_n 0.00104114f $X=6.395 $Y=0.655 $X2=0
+ $Y2=0
cc_374 N_A2_M1012_g N_A_867_47#_c_938_n 0.00917009f $X=6.825 $Y=0.655 $X2=0
+ $Y2=0
cc_375 N_A2_M1014_g N_A_867_47#_c_938_n 3.93732e-19 $X=7.255 $Y=0.655 $X2=0
+ $Y2=0
cc_376 A2 N_A_867_47#_c_938_n 0.0230694f $X=7.835 $Y=1.58 $X2=0 $Y2=0
cc_377 N_A2_c_386_n N_A_867_47#_c_938_n 0.00299787f $X=7.595 $Y=1.51 $X2=0 $Y2=0
cc_378 N_A_89_367#_c_465_n N_Y_M1006_d 0.00332344f $X=1.335 $Y=2.99 $X2=0 $Y2=0
cc_379 N_A_89_367#_c_467_n N_Y_M1023_d 0.00332344f $X=2.195 $Y=2.99 $X2=0 $Y2=0
cc_380 N_A_89_367#_c_469_n N_Y_M1000_d 0.00332344f $X=3.055 $Y=2.99 $X2=0 $Y2=0
cc_381 N_A_89_367#_c_471_n N_Y_M1016_d 0.00332344f $X=3.995 $Y=2.99 $X2=0 $Y2=0
cc_382 N_A_89_367#_c_465_n N_Y_c_571_n 0.0159805f $X=1.335 $Y=2.99 $X2=0 $Y2=0
cc_383 N_A_89_367#_M1015_s N_Y_c_564_n 0.00176461f $X=1.29 $Y=1.835 $X2=0 $Y2=0
cc_384 N_A_89_367#_c_509_p N_Y_c_564_n 0.0135055f $X=1.43 $Y=2.21 $X2=0 $Y2=0
cc_385 N_A_89_367#_c_454_n N_Y_c_565_n 0.00246889f $X=0.57 $Y=1.99 $X2=0 $Y2=0
cc_386 N_A_89_367#_c_467_n N_Y_c_582_n 0.0159805f $X=2.195 $Y=2.99 $X2=0 $Y2=0
cc_387 N_A_89_367#_M1027_s N_Y_c_566_n 0.00176461f $X=2.15 $Y=1.835 $X2=0 $Y2=0
cc_388 N_A_89_367#_c_513_p N_Y_c_566_n 0.0135055f $X=2.29 $Y=2.21 $X2=0 $Y2=0
cc_389 N_A_89_367#_c_469_n N_Y_c_589_n 0.0159805f $X=3.055 $Y=2.99 $X2=0 $Y2=0
cc_390 N_A_89_367#_M1008_s N_Y_c_568_n 0.00261503f $X=3.01 $Y=1.835 $X2=0 $Y2=0
cc_391 N_A_89_367#_c_516_p N_Y_c_568_n 0.0200142f $X=3.2 $Y=2.21 $X2=0 $Y2=0
cc_392 N_A_89_367#_c_456_n N_Y_c_568_n 0.00877753f $X=4.29 $Y=1.84 $X2=0 $Y2=0
cc_393 N_A_89_367#_c_471_n N_Y_c_612_n 0.0159805f $X=3.995 $Y=2.99 $X2=0 $Y2=0
cc_394 N_A_89_367#_c_455_n N_VPWR_M1013_s 0.00176461f $X=4.96 $Y=1.84 $X2=-0.19
+ $Y2=1.655
cc_395 N_A_89_367#_c_457_n N_VPWR_M1026_s 0.00224297f $X=5.82 $Y=1.84 $X2=0
+ $Y2=0
cc_396 N_A_89_367#_c_488_n N_VPWR_M1003_d 0.00427768f $X=6.725 $Y=2.015 $X2=0
+ $Y2=0
cc_397 N_A_89_367#_c_495_n N_VPWR_M1025_d 0.00331527f $X=7.585 $Y=2.015 $X2=0
+ $Y2=0
cc_398 N_A_89_367#_c_455_n N_VPWR_c_677_n 0.0170777f $X=4.96 $Y=1.84 $X2=0 $Y2=0
cc_399 N_A_89_367#_c_457_n N_VPWR_c_678_n 0.0189527f $X=5.82 $Y=1.84 $X2=0 $Y2=0
cc_400 N_A_89_367#_c_488_n N_VPWR_c_679_n 0.0170777f $X=6.725 $Y=2.015 $X2=0
+ $Y2=0
cc_401 N_A_89_367#_c_495_n N_VPWR_c_680_n 0.0170777f $X=7.585 $Y=2.015 $X2=0
+ $Y2=0
cc_402 N_A_89_367#_c_527_p N_VPWR_c_681_n 0.0140491f $X=5.96 $Y=2.46 $X2=0 $Y2=0
cc_403 N_A_89_367#_c_528_p N_VPWR_c_683_n 0.0124525f $X=6.82 $Y=2.91 $X2=0 $Y2=0
cc_404 N_A_89_367#_c_453_n N_VPWR_c_685_n 0.0179183f $X=0.535 $Y=2.905 $X2=0
+ $Y2=0
cc_405 N_A_89_367#_c_465_n N_VPWR_c_685_n 0.0361172f $X=1.335 $Y=2.99 $X2=0
+ $Y2=0
cc_406 N_A_89_367#_c_467_n N_VPWR_c_685_n 0.0361172f $X=2.195 $Y=2.99 $X2=0
+ $Y2=0
cc_407 N_A_89_367#_c_469_n N_VPWR_c_685_n 0.0361172f $X=3.055 $Y=2.99 $X2=0
+ $Y2=0
cc_408 N_A_89_367#_c_471_n N_VPWR_c_685_n 0.0361172f $X=3.995 $Y=2.99 $X2=0
+ $Y2=0
cc_409 N_A_89_367#_c_534_p N_VPWR_c_685_n 0.0199062f $X=4.142 $Y=2.905 $X2=0
+ $Y2=0
cc_410 N_A_89_367#_c_535_p N_VPWR_c_685_n 0.0125234f $X=1.43 $Y=2.91 $X2=0 $Y2=0
cc_411 N_A_89_367#_c_536_p N_VPWR_c_685_n 0.0125234f $X=2.29 $Y=2.99 $X2=0 $Y2=0
cc_412 N_A_89_367#_c_537_p N_VPWR_c_685_n 0.0181484f $X=3.19 $Y=2.99 $X2=0 $Y2=0
cc_413 N_A_89_367#_c_538_p N_VPWR_c_686_n 0.0124525f $X=5.055 $Y=1.98 $X2=0
+ $Y2=0
cc_414 N_A_89_367#_c_460_n N_VPWR_c_687_n 0.0178111f $X=7.68 $Y=2.91 $X2=0 $Y2=0
cc_415 N_A_89_367#_M1006_s N_VPWR_c_676_n 0.00215161f $X=0.445 $Y=1.835 $X2=0
+ $Y2=0
cc_416 N_A_89_367#_M1015_s N_VPWR_c_676_n 0.00223565f $X=1.29 $Y=1.835 $X2=0
+ $Y2=0
cc_417 N_A_89_367#_M1027_s N_VPWR_c_676_n 0.00223565f $X=2.15 $Y=1.835 $X2=0
+ $Y2=0
cc_418 N_A_89_367#_M1008_s N_VPWR_c_676_n 0.00287898f $X=3.01 $Y=1.835 $X2=0
+ $Y2=0
cc_419 N_A_89_367#_M1019_s N_VPWR_c_676_n 0.00461905f $X=3.95 $Y=1.835 $X2=0
+ $Y2=0
cc_420 N_A_89_367#_M1017_d N_VPWR_c_676_n 0.00536646f $X=4.915 $Y=1.835 $X2=0
+ $Y2=0
cc_421 N_A_89_367#_M1030_d N_VPWR_c_676_n 0.00380103f $X=5.82 $Y=1.835 $X2=0
+ $Y2=0
cc_422 N_A_89_367#_M1007_s N_VPWR_c_676_n 0.00536646f $X=6.68 $Y=1.835 $X2=0
+ $Y2=0
cc_423 N_A_89_367#_M1029_s N_VPWR_c_676_n 0.00371702f $X=7.54 $Y=1.835 $X2=0
+ $Y2=0
cc_424 N_A_89_367#_c_453_n N_VPWR_c_676_n 0.0101029f $X=0.535 $Y=2.905 $X2=0
+ $Y2=0
cc_425 N_A_89_367#_c_465_n N_VPWR_c_676_n 0.023676f $X=1.335 $Y=2.99 $X2=0 $Y2=0
cc_426 N_A_89_367#_c_467_n N_VPWR_c_676_n 0.023676f $X=2.195 $Y=2.99 $X2=0 $Y2=0
cc_427 N_A_89_367#_c_469_n N_VPWR_c_676_n 0.023676f $X=3.055 $Y=2.99 $X2=0 $Y2=0
cc_428 N_A_89_367#_c_471_n N_VPWR_c_676_n 0.023676f $X=3.995 $Y=2.99 $X2=0 $Y2=0
cc_429 N_A_89_367#_c_534_p N_VPWR_c_676_n 0.0114689f $X=4.142 $Y=2.905 $X2=0
+ $Y2=0
cc_430 N_A_89_367#_c_538_p N_VPWR_c_676_n 0.00730901f $X=5.055 $Y=1.98 $X2=0
+ $Y2=0
cc_431 N_A_89_367#_c_527_p N_VPWR_c_676_n 0.00904266f $X=5.96 $Y=2.46 $X2=0
+ $Y2=0
cc_432 N_A_89_367#_c_528_p N_VPWR_c_676_n 0.00730901f $X=6.82 $Y=2.91 $X2=0
+ $Y2=0
cc_433 N_A_89_367#_c_460_n N_VPWR_c_676_n 0.0100304f $X=7.68 $Y=2.91 $X2=0 $Y2=0
cc_434 N_A_89_367#_c_535_p N_VPWR_c_676_n 0.00738676f $X=1.43 $Y=2.91 $X2=0
+ $Y2=0
cc_435 N_A_89_367#_c_536_p N_VPWR_c_676_n 0.00738676f $X=2.29 $Y=2.99 $X2=0
+ $Y2=0
cc_436 N_A_89_367#_c_537_p N_VPWR_c_676_n 0.010497f $X=3.19 $Y=2.99 $X2=0 $Y2=0
cc_437 N_Y_M1006_d N_VPWR_c_676_n 0.00225186f $X=0.86 $Y=1.835 $X2=0 $Y2=0
cc_438 N_Y_M1023_d N_VPWR_c_676_n 0.00225186f $X=1.72 $Y=1.835 $X2=0 $Y2=0
cc_439 N_Y_M1000_d N_VPWR_c_676_n 0.00225186f $X=2.58 $Y=1.835 $X2=0 $Y2=0
cc_440 N_Y_M1016_d N_VPWR_c_676_n 0.00225186f $X=3.52 $Y=1.835 $X2=0 $Y2=0
cc_441 N_Y_c_563_n N_A_63_65#_M1011_d 0.00336891f $X=5.645 $Y=0.927 $X2=0 $Y2=0
cc_442 N_Y_c_563_n N_A_63_65#_M1024_d 0.00529081f $X=5.645 $Y=0.927 $X2=0 $Y2=0
cc_443 N_Y_c_594_n N_A_63_65#_c_798_n 0.0135888f $X=2.65 $Y=0.7 $X2=0 $Y2=0
cc_444 N_Y_c_594_n N_A_63_65#_c_806_n 0.0197298f $X=2.65 $Y=0.7 $X2=0 $Y2=0
cc_445 N_Y_c_563_n N_A_63_65#_c_788_n 0.0584168f $X=5.645 $Y=0.927 $X2=0 $Y2=0
cc_446 N_Y_M1020_s N_A_63_65#_c_789_n 0.00177018f $X=3.37 $Y=0.325 $X2=0 $Y2=0
cc_447 N_Y_M1001_s N_A_63_65#_c_790_n 0.00176461f $X=2.51 $Y=0.325 $X2=0 $Y2=0
cc_448 N_Y_c_563_n N_A_63_65#_c_790_n 0.00378766f $X=5.645 $Y=0.927 $X2=0 $Y2=0
cc_449 N_Y_c_594_n N_A_63_65#_c_790_n 0.0200589f $X=2.65 $Y=0.7 $X2=0 $Y2=0
cc_450 N_Y_M1004_s N_VGND_c_846_n 0.00225919f $X=4.75 $Y=0.235 $X2=0 $Y2=0
cc_451 N_Y_M1021_s N_VGND_c_846_n 0.00225112f $X=5.61 $Y=0.235 $X2=0 $Y2=0
cc_452 N_Y_c_563_n N_VGND_c_846_n 0.0143579f $X=5.645 $Y=0.927 $X2=0 $Y2=0
cc_453 N_Y_c_563_n N_A_867_47#_M1004_d 0.00554433f $X=5.645 $Y=0.927 $X2=-0.19
+ $Y2=-0.245
cc_454 N_Y_c_563_n N_A_867_47#_M1005_d 0.00377422f $X=5.645 $Y=0.927 $X2=0 $Y2=0
cc_455 N_Y_M1004_s N_A_867_47#_c_935_n 0.00381621f $X=4.75 $Y=0.235 $X2=0 $Y2=0
cc_456 N_Y_M1021_s N_A_867_47#_c_935_n 0.00335534f $X=5.61 $Y=0.235 $X2=0 $Y2=0
cc_457 N_Y_c_631_n N_A_867_47#_c_935_n 0.0125888f $X=5.75 $Y=0.86 $X2=0 $Y2=0
cc_458 N_Y_c_563_n N_A_867_47#_c_935_n 0.046282f $X=5.645 $Y=0.927 $X2=0 $Y2=0
cc_459 N_A_63_65#_c_792_n N_VGND_M1009_s 0.003325f $X=1.205 $Y=0.955 $X2=-0.19
+ $Y2=-0.245
cc_460 N_A_63_65#_c_798_n N_VGND_M1018_s 0.003325f $X=2.065 $Y=0.955 $X2=0 $Y2=0
cc_461 N_A_63_65#_c_784_n N_VGND_c_838_n 0.0148073f $X=0.44 $Y=0.48 $X2=0 $Y2=0
cc_462 N_A_63_65#_c_792_n N_VGND_c_838_n 0.0170777f $X=1.205 $Y=0.955 $X2=0
+ $Y2=0
cc_463 N_A_63_65#_c_786_n N_VGND_c_838_n 0.0147905f $X=1.3 $Y=0.48 $X2=0 $Y2=0
cc_464 N_A_63_65#_c_786_n N_VGND_c_839_n 0.0147905f $X=1.3 $Y=0.48 $X2=0 $Y2=0
cc_465 N_A_63_65#_c_798_n N_VGND_c_839_n 0.0170777f $X=2.065 $Y=0.955 $X2=0
+ $Y2=0
cc_466 N_A_63_65#_c_787_n N_VGND_c_839_n 0.00962585f $X=2.245 $Y=0.34 $X2=0
+ $Y2=0
cc_467 N_A_63_65#_c_786_n N_VGND_c_842_n 0.00975394f $X=1.3 $Y=0.48 $X2=0 $Y2=0
cc_468 N_A_63_65#_c_787_n N_VGND_c_843_n 0.0129036f $X=2.245 $Y=0.34 $X2=0 $Y2=0
cc_469 N_A_63_65#_c_790_n N_VGND_c_843_n 0.117984f $X=2.995 $Y=0.445 $X2=0 $Y2=0
cc_470 N_A_63_65#_c_784_n N_VGND_c_846_n 0.00972454f $X=0.44 $Y=0.48 $X2=0 $Y2=0
cc_471 N_A_63_65#_c_786_n N_VGND_c_846_n 0.0070861f $X=1.3 $Y=0.48 $X2=0 $Y2=0
cc_472 N_A_63_65#_c_787_n N_VGND_c_846_n 0.00699798f $X=2.245 $Y=0.34 $X2=0
+ $Y2=0
cc_473 N_A_63_65#_c_790_n N_VGND_c_846_n 0.0656511f $X=2.995 $Y=0.445 $X2=0
+ $Y2=0
cc_474 N_A_63_65#_c_784_n N_VGND_c_847_n 0.0133857f $X=0.44 $Y=0.48 $X2=0 $Y2=0
cc_475 N_A_63_65#_c_789_n N_A_867_47#_c_935_n 0.0173369f $X=3.94 $Y=0.47 $X2=0
+ $Y2=0
cc_476 N_VGND_c_846_n N_A_867_47#_M1004_d 0.00215867f $X=7.92 $Y=0 $X2=-0.19
+ $Y2=-0.245
cc_477 N_VGND_c_846_n N_A_867_47#_M1005_d 0.00224306f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_478 N_VGND_c_846_n N_A_867_47#_M1022_d 0.00249042f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_479 N_VGND_c_846_n N_A_867_47#_M1012_s 0.00404131f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_480 N_VGND_c_846_n N_A_867_47#_M1031_s 0.00371702f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_481 N_VGND_c_843_n N_A_867_47#_c_935_n 0.0877189f $X=6.445 $Y=0 $X2=0 $Y2=0
cc_482 N_VGND_c_846_n N_A_867_47#_c_935_n 0.0615994f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_483 N_VGND_c_843_n N_A_867_47#_c_944_n 0.0140077f $X=6.445 $Y=0 $X2=0 $Y2=0
cc_484 N_VGND_c_846_n N_A_867_47#_c_944_n 0.00982246f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_485 N_VGND_M1002_d N_A_867_47#_c_948_n 0.00470865f $X=6.47 $Y=0.235 $X2=0
+ $Y2=0
cc_486 N_VGND_c_840_n N_A_867_47#_c_948_n 0.0171165f $X=6.61 $Y=0.48 $X2=0 $Y2=0
cc_487 N_VGND_c_846_n N_A_867_47#_c_948_n 0.00916249f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_488 N_VGND_c_844_n N_A_867_47#_c_982_n 0.0124525f $X=7.305 $Y=0 $X2=0 $Y2=0
cc_489 N_VGND_c_846_n N_A_867_47#_c_982_n 0.00730901f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_490 N_VGND_M1014_d N_A_867_47#_c_936_n 0.00177068f $X=7.33 $Y=0.235 $X2=0
+ $Y2=0
cc_491 N_VGND_c_841_n N_A_867_47#_c_936_n 0.0172078f $X=7.47 $Y=0.38 $X2=0 $Y2=0
cc_492 N_VGND_c_845_n N_A_867_47#_c_937_n 0.0178111f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_493 N_VGND_c_846_n N_A_867_47#_c_937_n 0.0100304f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_494 N_VGND_c_846_n N_A_867_47#_c_938_n 0.00318091f $X=7.92 $Y=0 $X2=0 $Y2=0
