* File: sky130_fd_sc_lp__a311oi_0.spice
* Created: Fri Aug 28 09:58:07 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__a311oi_0.pex.spice"
.subckt sky130_fd_sc_lp__a311oi_0  VNB VPB A3 A2 A1 B1 C1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* C1	C1
* B1	B1
* A1	A1
* A2	A2
* A3	A3
* VPB	VPB
* VNB	VNB
MM1006 A_180_47# N_A3_M1006_g N_VGND_M1006_s VNB NSHORT L=0.15 W=0.42 AD=0.0441
+ AS=0.2541 PD=0.63 PS=2.05 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.5 SB=75002.1
+ A=0.063 P=1.14 MULT=1
MM1007 A_252_47# N_A2_M1007_g A_180_47# VNB NSHORT L=0.15 W=0.42 AD=0.0441
+ AS=0.0441 PD=0.63 PS=0.63 NRD=14.28 NRS=14.28 M=1 R=2.8 SA=75000.9 SB=75001.8
+ A=0.063 P=1.14 MULT=1
MM1003 N_Y_M1003_d N_A1_M1003_g A_252_47# VNB NSHORT L=0.15 W=0.42 AD=0.0651
+ AS=0.0441 PD=0.73 PS=0.63 NRD=4.284 NRS=14.28 M=1 R=2.8 SA=75001.2 SB=75001.4
+ A=0.063 P=1.14 MULT=1
MM1009 N_VGND_M1009_d N_B1_M1009_g N_Y_M1003_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1302 AS=0.0651 PD=1.04 PS=0.73 NRD=0 NRS=4.284 M=1 R=2.8 SA=75001.7
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1004 N_Y_M1004_d N_C1_M1004_g N_VGND_M1009_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.1302 PD=1.37 PS=1.04 NRD=0 NRS=0 M=1 R=2.8 SA=75002.5
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1000 N_A_158_473#_M1000_d N_A3_M1000_g N_VPWR_M1000_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.0896 AS=0.1696 PD=0.92 PS=1.81 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75001.9 A=0.096 P=1.58 MULT=1
MM1005 N_VPWR_M1005_d N_A2_M1005_g N_A_158_473#_M1000_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.6 SB=75001.5 A=0.096 P=1.58 MULT=1
MM1001 N_A_158_473#_M1001_d N_A1_M1001_g N_VPWR_M1005_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1152 AS=0.0896 PD=1 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667 SA=75001.1
+ SB=75001.1 A=0.096 P=1.58 MULT=1
MM1002 A_432_473# N_B1_M1002_g N_A_158_473#_M1001_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0672 AS=0.1152 PD=0.85 PS=1 NRD=15.3857 NRS=24.6053 M=1 R=4.26667
+ SA=75001.6 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1008 N_Y_M1008_d N_C1_M1008_g A_432_473# VPB PHIGHVT L=0.15 W=0.64 AD=0.1696
+ AS=0.0672 PD=1.81 PS=0.85 NRD=0 NRS=15.3857 M=1 R=4.26667 SA=75001.9
+ SB=75000.2 A=0.096 P=1.58 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9751 P=11.21
c_72 VPB 0 2.80181e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_lp__a311oi_0.pxi.spice"
*
.ends
*
*
