* NGSPICE file created from sky130_fd_sc_lp__nor3b_1.ext - technology: sky130A

.subckt sky130_fd_sc_lp__nor3b_1 A B C_N VGND VNB VPB VPWR Y
M1000 VGND C_N a_82_131# VNB nshort w=420000u l=150000u
+  ad=5.187e+11p pd=4.73e+06u as=1.113e+11p ps=1.37e+06u
M1001 Y a_82_131# a_347_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=3.528e+11p pd=3.08e+06u as=4.914e+11p ps=3.3e+06u
M1002 Y A VGND VNB nshort w=840000u l=150000u
+  ad=4.872e+11p pd=4.52e+06u as=0p ps=0u
M1003 VGND B Y VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VPWR C_N a_82_131# VPB phighvt w=420000u l=150000u
+  ad=3.906e+11p pd=3.32e+06u as=1.113e+11p ps=1.37e+06u
M1005 Y a_82_131# VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_275_367# A VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=2.646e+11p pd=2.94e+06u as=0p ps=0u
M1007 a_347_367# B a_275_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

