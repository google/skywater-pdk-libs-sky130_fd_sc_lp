* File: sky130_fd_sc_lp__einvp_lp.spice
* Created: Fri Aug 28 10:34:14 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__einvp_lp.pex.spice"
.subckt sky130_fd_sc_lp__einvp_lp  VNB VPB A TE Z VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Z	Z
* TE	TE
* A	A
* VPB	VPB
* VNB	VNB
MM1005 A_134_141# N_A_M1005_g N_Z_M1005_s VNB NSHORT L=0.15 W=0.42 AD=0.0504
+ AS=0.16345 PD=0.66 PS=1.64 NRD=18.564 NRS=22.848 M=1 R=2.8 SA=75000.3
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1004 N_VGND_M1004_d N_TE_M1004_g A_134_141# VNB NSHORT L=0.15 W=0.42 AD=0.0931
+ AS=0.0504 PD=0.98 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75000.7 SB=75000.7
+ A=0.063 P=1.14 MULT=1
MM1002 A_314_101# N_TE_M1002_g N_VGND_M1004_d VNB NSHORT L=0.15 W=0.42 AD=0.0441
+ AS=0.0931 PD=0.63 PS=0.98 NRD=14.28 NRS=24.276 M=1 R=2.8 SA=75000.7 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1000 N_A_182_321#_M1000_d N_TE_M1000_g A_314_101# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.1
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1006 A_134_419# N_A_M1006_g N_Z_M1006_s VPB PHIGHVT L=0.25 W=1 AD=0.12
+ AS=0.285 PD=1.24 PS=2.57 NRD=12.7853 NRS=0 M=1 R=4 SA=125000 SB=125001 A=0.25
+ P=2.5 MULT=1
MM1001 N_VPWR_M1001_d N_A_182_321#_M1001_g A_134_419# VPB PHIGHVT L=0.25 W=1
+ AD=0.2825 AS=0.12 PD=1.565 PS=1.24 NRD=56.145 NRS=12.7853 M=1 R=4 SA=125001
+ SB=125001 A=0.25 P=2.5 MULT=1
MM1003 N_A_182_321#_M1003_d N_TE_M1003_g N_VPWR_M1001_d VPB PHIGHVT L=0.25 W=1
+ AD=0.285 AS=0.2825 PD=2.57 PS=1.565 NRD=0 NRS=0 M=1 R=4 SA=125001 SB=125000
+ A=0.25 P=2.5 MULT=1
DX7_noxref VNB VPB NWDIODE A=5.1847 P=9.29
*
.include "sky130_fd_sc_lp__einvp_lp.pxi.spice"
*
.ends
*
*
