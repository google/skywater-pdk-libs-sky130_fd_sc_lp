* File: sky130_fd_sc_lp__nor3_lp.pex.spice
* Created: Wed Sep  2 10:09:19 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__NOR3_LP%C 3 5 6 9 11 13 15 16 17 18 22
c49 17 0 2.70706e-20 $X=1.2 $Y=1.295
r50 17 18 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.22 $Y=1.295
+ $X2=1.22 $Y2=1.665
r51 17 22 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.22
+ $Y=1.34 $X2=1.22 $Y2=1.34
r52 16 22 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.22 $Y=1.68
+ $X2=1.22 $Y2=1.34
r53 14 22 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=1.22 $Y=1.325
+ $X2=1.22 $Y2=1.34
r54 14 15 13.5877 $w=2.4e-07 $l=7.5e-08 $layer=POLY_cond $X=1.22 $Y=1.325
+ $X2=1.22 $Y2=1.25
r55 11 16 47.383 $w=2.95e-07 $l=3.53129e-07 $layer=POLY_cond $X=1.36 $Y=1.97
+ $X2=1.22 $Y2=1.68
r56 11 13 110.86 $w=2.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.36 $Y=1.97
+ $X2=1.36 $Y2=2.545
r57 7 15 13.5877 $w=2.4e-07 $l=1.04283e-07 $layer=POLY_cond $X=1.15 $Y=1.175
+ $X2=1.22 $Y2=1.25
r58 7 9 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=1.15 $Y=1.175 $X2=1.15
+ $Y2=0.495
r59 5 15 12.1617 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.055 $Y=1.25
+ $X2=1.22 $Y2=1.25
r60 5 6 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=1.055 $Y=1.25
+ $X2=0.865 $Y2=1.25
r61 1 6 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.79 $Y=1.175
+ $X2=0.865 $Y2=1.25
r62 1 3 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=0.79 $Y=1.175 $X2=0.79
+ $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__NOR3_LP%B 1 3 8 10 12 16 19 20 21 22 23 24 25 26 43
c58 19 0 2.70706e-20 $X=1.89 $Y=1.18
r59 43 44 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.89
+ $Y=1.345 $X2=1.89 $Y2=1.345
r60 25 26 6.23308 $w=7.08e-07 $l=3.7e-07 $layer=LI1_cond $X=1.92 $Y=2.405
+ $X2=1.92 $Y2=2.775
r61 24 25 6.23308 $w=7.08e-07 $l=3.7e-07 $layer=LI1_cond $X=1.92 $Y=2.035
+ $X2=1.92 $Y2=2.405
r62 23 24 6.23308 $w=7.08e-07 $l=3.7e-07 $layer=LI1_cond $X=1.92 $Y=1.665
+ $X2=1.92 $Y2=2.035
r63 23 44 5.39078 $w=7.08e-07 $l=3.2e-07 $layer=LI1_cond $X=1.92 $Y=1.665
+ $X2=1.92 $Y2=1.345
r64 22 44 0.842309 $w=7.08e-07 $l=5e-08 $layer=LI1_cond $X=1.92 $Y=1.295
+ $X2=1.92 $Y2=1.345
r65 20 43 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.89 $Y=1.685
+ $X2=1.89 $Y2=1.345
r66 20 21 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.89 $Y=1.685
+ $X2=1.89 $Y2=1.85
r67 19 43 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.89 $Y=1.18
+ $X2=1.89 $Y2=1.345
r68 15 16 71.7872 $w=1.5e-07 $l=1.4e-07 $layer=POLY_cond $X=1.8 $Y=0.855
+ $X2=1.94 $Y2=0.855
r69 13 15 112.809 $w=1.5e-07 $l=2.2e-07 $layer=POLY_cond $X=1.58 $Y=0.855
+ $X2=1.8 $Y2=0.855
r70 10 16 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.94 $Y=0.78
+ $X2=1.94 $Y2=0.855
r71 10 12 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=1.94 $Y=0.78 $X2=1.94
+ $Y2=0.495
r72 8 21 172.675 $w=2.5e-07 $l=6.95e-07 $layer=POLY_cond $X=1.85 $Y=2.545
+ $X2=1.85 $Y2=1.85
r73 4 15 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.8 $Y=0.93 $X2=1.8
+ $Y2=0.855
r74 4 19 128.191 $w=1.5e-07 $l=2.5e-07 $layer=POLY_cond $X=1.8 $Y=0.93 $X2=1.8
+ $Y2=1.18
r75 1 13 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.58 $Y=0.78 $X2=1.58
+ $Y2=0.855
r76 1 3 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=1.58 $Y=0.78 $X2=1.58
+ $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__NOR3_LP%A 3 7 9 12 14 15 17 24
r32 24 26 80.7798 $w=5.6e-07 $l=5.05e-07 $layer=POLY_cond $X=2.575 $Y=1.17
+ $X2=2.575 $Y2=1.675
r33 24 25 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.69
+ $Y=1.17 $X2=2.69 $Y2=1.17
r34 17 25 6.63631 $w=7.73e-07 $l=4.3e-07 $layer=LI1_cond $X=3.12 $Y=1.392
+ $X2=2.69 $Y2=1.392
r35 15 25 0.771663 $w=7.73e-07 $l=5e-08 $layer=LI1_cond $X=2.64 $Y=1.392
+ $X2=2.69 $Y2=1.392
r36 14 26 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=2.37 $Y=1.915
+ $X2=2.37 $Y2=1.675
r37 10 24 30.7275 $w=2.8e-07 $l=2.29783e-07 $layer=POLY_cond $X=2.73 $Y=1.005
+ $X2=2.575 $Y2=1.17
r38 10 12 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=2.73 $Y=1.005
+ $X2=2.73 $Y2=0.495
r39 7 14 40.9178 $w=2.5e-07 $l=1.25e-07 $layer=POLY_cond $X=2.42 $Y=2.04
+ $X2=2.42 $Y2=1.915
r40 7 9 97.364 $w=2.5e-07 $l=5.05e-07 $layer=POLY_cond $X=2.42 $Y=2.04 $X2=2.42
+ $Y2=2.545
r41 1 24 30.7275 $w=2.8e-07 $l=2.75409e-07 $layer=POLY_cond $X=2.37 $Y=1.005
+ $X2=2.575 $Y2=1.17
r42 1 3 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=2.37 $Y=1.005 $X2=2.37
+ $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__NOR3_LP%Y 1 2 3 12 14 17 19 20 21 22 27 41 61
r51 42 55 2.22521 $w=7.1e-07 $l=5.2e-07 $layer=LI1_cond $X=0.48 $Y=2.025
+ $X2=0.48 $Y2=2.545
r52 27 61 5 $w=9.15e-07 $l=3.75e-07 $layer=LI1_cond $X=0.72 $Y=2.545 $X2=1.095
+ $Y2=2.545
r53 27 55 3.2 $w=9.15e-07 $l=2.4e-07 $layer=LI1_cond $X=0.72 $Y=2.545 $X2=0.48
+ $Y2=2.545
r54 22 55 3.2 $w=9.15e-07 $l=2.4e-07 $layer=LI1_cond $X=0.24 $Y=2.545 $X2=0.48
+ $Y2=2.545
r55 21 27 11.1165 $w=1.7e-07 $l=4.73e-07 $layer=LI1_cond $X=0.72 $Y=2.072
+ $X2=0.72 $Y2=2.545
r56 21 22 11.1165 $w=1.7e-07 $l=4.73e-07 $layer=LI1_cond $X=0.24 $Y=2.072
+ $X2=0.24 $Y2=2.545
r57 21 42 0.640155 $w=7.08e-07 $l=3.8e-08 $layer=LI1_cond $X=0.48 $Y=1.987
+ $X2=0.48 $Y2=2.025
r58 20 21 5.42447 $w=7.08e-07 $l=3.22e-07 $layer=LI1_cond $X=0.48 $Y=1.665
+ $X2=0.48 $Y2=1.987
r59 20 41 2.19 $w=7.08e-07 $l=1.3e-07 $layer=LI1_cond $X=0.48 $Y=1.665 $X2=0.48
+ $Y2=1.535
r60 19 41 4.65384 $w=7.1e-07 $l=2.4e-07 $layer=LI1_cond $X=0.48 $Y=1.295
+ $X2=0.48 $Y2=1.535
r61 19 47 8.28395 $w=5.67e-07 $l=3.85e-07 $layer=LI1_cond $X=0.48 $Y=1.295
+ $X2=0.48 $Y2=0.91
r62 17 18 18.7519 $w=2.7e-07 $l=4.15e-07 $layer=LI1_cond $X=2.155 $Y=0.495
+ $X2=2.155 $Y2=0.91
r63 15 47 7.95352 $w=1.7e-07 $l=3.55e-07 $layer=LI1_cond $X=0.835 $Y=0.91
+ $X2=0.48 $Y2=0.91
r64 14 18 3.44395 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.99 $Y=0.91
+ $X2=2.155 $Y2=0.91
r65 14 15 75.3529 $w=1.68e-07 $l=1.155e-06 $layer=LI1_cond $X=1.99 $Y=0.91
+ $X2=0.835 $Y2=0.91
r66 10 47 3.94259 $w=5.67e-07 $l=1.30767e-07 $layer=LI1_cond $X=0.575 $Y=0.825
+ $X2=0.48 $Y2=0.91
r67 10 12 11.5244 $w=3.28e-07 $l=3.3e-07 $layer=LI1_cond $X=0.575 $Y=0.825
+ $X2=0.575 $Y2=0.495
r68 3 61 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.95
+ $Y=2.045 $X2=1.095 $Y2=2.9
r69 3 61 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.95
+ $Y=2.045 $X2=1.095 $Y2=2.19
r70 2 17 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.015
+ $Y=0.285 $X2=2.155 $Y2=0.495
r71 1 12 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.43
+ $Y=0.285 $X2=0.575 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__NOR3_LP%VPWR 1 6 10 12 22 23 26
r21 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r22 23 27 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.64 $Y2=3.33
r23 22 23 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r24 20 26 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.85 $Y=3.33
+ $X2=2.685 $Y2=3.33
r25 20 22 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=2.85 $Y=3.33 $X2=3.12
+ $Y2=3.33
r26 19 27 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r27 18 19 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r28 14 18 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=0.24 $Y=3.33
+ $X2=2.16 $Y2=3.33
r29 14 15 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r30 12 26 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.52 $Y=3.33
+ $X2=2.685 $Y2=3.33
r31 12 18 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=2.52 $Y=3.33
+ $X2=2.16 $Y2=3.33
r32 10 19 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r33 10 15 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.24 $Y2=3.33
r34 6 9 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=2.685 $Y=2.19 $X2=2.685
+ $Y2=2.9
r35 4 26 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.685 $Y=3.245
+ $X2=2.685 $Y2=3.33
r36 4 9 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=2.685 $Y=3.245
+ $X2=2.685 $Y2=2.9
r37 1 9 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=2.545
+ $Y=2.045 $X2=2.685 $Y2=2.9
r38 1 6 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.545
+ $Y=2.045 $X2=2.685 $Y2=2.19
.ends

.subckt PM_SKY130_FD_SC_LP__NOR3_LP%VGND 1 2 9 11 13 15 17 22 31 35
r39 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r40 31 32 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r41 29 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r42 28 29 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r43 25 28 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r44 23 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.53 $Y=0 $X2=1.365
+ $Y2=0
r45 23 25 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=1.53 $Y=0 $X2=1.68
+ $Y2=0
r46 22 34 4.50438 $w=1.7e-07 $l=2.9e-07 $layer=LI1_cond $X=2.78 $Y=0 $X2=3.07
+ $Y2=0
r47 22 28 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=2.78 $Y=0 $X2=2.64
+ $Y2=0
r48 20 32 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r49 19 20 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r50 17 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.2 $Y=0 $X2=1.365
+ $Y2=0
r51 17 19 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=0 $X2=0.24
+ $Y2=0
r52 15 29 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r53 15 32 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r54 15 25 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r55 11 34 3.26179 $w=3.3e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.945 $Y=0.085
+ $X2=3.07 $Y2=0
r56 11 13 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=2.945 $Y=0.085
+ $X2=2.945 $Y2=0.495
r57 7 31 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.365 $Y=0.085
+ $X2=1.365 $Y2=0
r58 7 9 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.365 $Y=0.085
+ $X2=1.365 $Y2=0.455
r59 2 13 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.805
+ $Y=0.285 $X2=2.945 $Y2=0.495
r60 1 9 182 $w=1.7e-07 $l=2.29565e-07 $layer=licon1_NDIFF $count=1 $X=1.225
+ $Y=0.285 $X2=1.365 $Y2=0.455
.ends

