* File: sky130_fd_sc_lp__o21ai_lp.spice
* Created: Fri Aug 28 11:05:08 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__o21ai_lp.pex.spice"
.subckt sky130_fd_sc_lp__o21ai_lp  VNB VPB A1 A2 B1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B1	B1
* A2	A2
* A1	A1
* VPB	VPB
* VNB	VNB
MM1001 N_VGND_M1001_d N_A1_M1001_g N_A_64_57#_M1001_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0924 AS=0.1197 PD=0.86 PS=1.41 NRD=22.848 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.3 A=0.063 P=1.14 MULT=1
MM1003 N_A_64_57#_M1003_d N_A2_M1003_g N_VGND_M1001_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0924 PD=0.7 PS=0.86 NRD=0 NRS=22.848 M=1 R=2.8 SA=75000.8
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1005 N_Y_M1005_d N_B1_M1005_g N_A_64_57#_M1003_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1533 AS=0.0588 PD=1.57 PS=0.7 NRD=22.848 NRS=0 M=1 R=2.8 SA=75001.2
+ SB=75000.3 A=0.063 P=1.14 MULT=1
MM1000 A_155_409# N_A1_M1000_g N_VPWR_M1000_s VPB PHIGHVT L=0.25 W=1 AD=0.12
+ AS=0.285 PD=1.24 PS=2.57 NRD=12.7853 NRS=0 M=1 R=4 SA=125000 SB=125001 A=0.25
+ P=2.5 MULT=1
MM1004 N_Y_M1004_d N_A2_M1004_g A_155_409# VPB PHIGHVT L=0.25 W=1 AD=0.16
+ AS=0.12 PD=1.32 PS=1.24 NRD=0 NRS=12.7853 M=1 R=4 SA=125001 SB=125001 A=0.25
+ P=2.5 MULT=1
MM1002 N_VPWR_M1002_d N_B1_M1002_g N_Y_M1004_d VPB PHIGHVT L=0.25 W=1 AD=0.285
+ AS=0.16 PD=2.57 PS=1.32 NRD=0 NRS=7.8603 M=1 R=4 SA=125001 SB=125000 A=0.25
+ P=2.5 MULT=1
DX6_noxref VNB VPB NWDIODE A=5.1847 P=9.29
*
.include "sky130_fd_sc_lp__o21ai_lp.pxi.spice"
*
.ends
*
*
