* File: sky130_fd_sc_lp__busdriver2_20.pxi.spice
* Created: Wed Sep  2 09:37:06 2020
* 
x_PM_SKY130_FD_SC_LP__BUSDRIVER2_20%TE_B N_TE_B_c_389_n N_TE_B_M1020_g
+ N_TE_B_M1004_g N_TE_B_c_391_n N_TE_B_c_392_n N_TE_B_M1024_g N_TE_B_M1007_g
+ N_TE_B_c_394_n TE_B N_TE_B_c_396_n PM_SKY130_FD_SC_LP__BUSDRIVER2_20%TE_B
x_PM_SKY130_FD_SC_LP__BUSDRIVER2_20%A_114_47# N_A_114_47#_M1020_s
+ N_A_114_47#_M1004_s N_A_114_47#_M1049_g N_A_114_47#_M1010_g
+ N_A_114_47#_M1054_g N_A_114_47#_c_432_n N_A_114_47#_c_433_n
+ N_A_114_47#_M1043_g N_A_114_47#_M1068_g N_A_114_47#_c_436_n
+ N_A_114_47#_M1071_g N_A_114_47#_c_438_n N_A_114_47#_M1003_g
+ N_A_114_47#_c_439_n N_A_114_47#_c_440_n N_A_114_47#_c_441_n
+ N_A_114_47#_M1011_g N_A_114_47#_c_442_n N_A_114_47#_M1015_g
+ N_A_114_47#_c_443_n N_A_114_47#_M1016_g N_A_114_47#_c_444_n
+ N_A_114_47#_M1035_g N_A_114_47#_c_445_n N_A_114_47#_c_446_n
+ N_A_114_47#_c_447_n N_A_114_47#_M1039_g N_A_114_47#_c_448_n
+ N_A_114_47#_M1044_g N_A_114_47#_c_449_n N_A_114_47#_c_450_n
+ N_A_114_47#_M1045_g N_A_114_47#_c_451_n N_A_114_47#_c_452_n
+ N_A_114_47#_M1047_g N_A_114_47#_c_453_n N_A_114_47#_c_454_n
+ N_A_114_47#_M1051_g N_A_114_47#_c_455_n N_A_114_47#_c_456_n
+ N_A_114_47#_M1057_g N_A_114_47#_c_457_n N_A_114_47#_c_458_n
+ N_A_114_47#_M1066_g N_A_114_47#_c_459_n N_A_114_47#_c_460_n
+ N_A_114_47#_M1070_g N_A_114_47#_c_461_n N_A_114_47#_c_462_n
+ N_A_114_47#_M1080_g N_A_114_47#_c_463_n N_A_114_47#_c_464_n
+ N_A_114_47#_c_465_n N_A_114_47#_c_466_n N_A_114_47#_c_467_n
+ N_A_114_47#_c_468_n N_A_114_47#_c_469_n N_A_114_47#_c_596_p
+ N_A_114_47#_c_470_n N_A_114_47#_c_486_n N_A_114_47#_c_508_p
+ N_A_114_47#_c_509_p N_A_114_47#_c_471_n N_A_114_47#_c_472_n
+ PM_SKY130_FD_SC_LP__BUSDRIVER2_20%A_114_47#
x_PM_SKY130_FD_SC_LP__BUSDRIVER2_20%A_286_367# N_A_286_367#_M1010_s
+ N_A_286_367#_M1049_d N_A_286_367#_M1068_d N_A_286_367#_c_731_n
+ N_A_286_367#_M1001_g N_A_286_367#_c_704_n N_A_286_367#_c_705_n
+ N_A_286_367#_c_734_n N_A_286_367#_M1005_g N_A_286_367#_c_706_n
+ N_A_286_367#_c_736_n N_A_286_367#_M1012_g N_A_286_367#_c_707_n
+ N_A_286_367#_c_738_n N_A_286_367#_M1018_g N_A_286_367#_c_708_n
+ N_A_286_367#_c_740_n N_A_286_367#_M1019_g N_A_286_367#_c_709_n
+ N_A_286_367#_c_742_n N_A_286_367#_M1022_g N_A_286_367#_c_710_n
+ N_A_286_367#_c_744_n N_A_286_367#_M1037_g N_A_286_367#_c_711_n
+ N_A_286_367#_c_746_n N_A_286_367#_M1040_g N_A_286_367#_c_712_n
+ N_A_286_367#_c_748_n N_A_286_367#_M1041_g N_A_286_367#_c_749_n
+ N_A_286_367#_M1055_g N_A_286_367#_c_750_n N_A_286_367#_M1058_g
+ N_A_286_367#_c_751_n N_A_286_367#_M1061_g N_A_286_367#_c_752_n
+ N_A_286_367#_M1064_g N_A_286_367#_c_753_n N_A_286_367#_M1065_g
+ N_A_286_367#_c_754_n N_A_286_367#_M1069_g N_A_286_367#_c_755_n
+ N_A_286_367#_M1074_g N_A_286_367#_c_756_n N_A_286_367#_M1077_g
+ N_A_286_367#_c_713_n N_A_286_367#_c_714_n N_A_286_367#_c_759_n
+ N_A_286_367#_M1084_g N_A_286_367#_c_715_n N_A_286_367#_c_761_n
+ N_A_286_367#_M1087_g N_A_286_367#_c_716_n N_A_286_367#_c_763_n
+ N_A_286_367#_M1089_g N_A_286_367#_c_717_n N_A_286_367#_c_718_n
+ N_A_286_367#_c_719_n N_A_286_367#_c_720_n N_A_286_367#_c_721_n
+ N_A_286_367#_c_722_n N_A_286_367#_c_723_n N_A_286_367#_c_724_n
+ N_A_286_367#_c_725_n N_A_286_367#_c_777_n N_A_286_367#_c_726_n
+ N_A_286_367#_c_774_n N_A_286_367#_c_775_n N_A_286_367#_c_808_n
+ N_A_286_367#_c_727_n N_A_286_367#_c_728_n N_A_286_367#_c_729_n
+ N_A_286_367#_c_730_n PM_SKY130_FD_SC_LP__BUSDRIVER2_20%A_286_367#
x_PM_SKY130_FD_SC_LP__BUSDRIVER2_20%A_1909_21# N_A_1909_21#_M1028_d
+ N_A_1909_21#_M1082_d N_A_1909_21#_M1009_s N_A_1909_21#_M1034_s
+ N_A_1909_21#_M1072_s N_A_1909_21#_M1079_s N_A_1909_21#_c_1033_n
+ N_A_1909_21#_M1017_g N_A_1909_21#_c_1034_n N_A_1909_21#_c_1035_n
+ N_A_1909_21#_c_1036_n N_A_1909_21#_M1021_g N_A_1909_21#_c_1037_n
+ N_A_1909_21#_c_1038_n N_A_1909_21#_M1027_g N_A_1909_21#_c_1039_n
+ N_A_1909_21#_c_1040_n N_A_1909_21#_M1031_g N_A_1909_21#_c_1041_n
+ N_A_1909_21#_c_1042_n N_A_1909_21#_M1033_g N_A_1909_21#_c_1043_n
+ N_A_1909_21#_c_1044_n N_A_1909_21#_M1036_g N_A_1909_21#_M1000_g
+ N_A_1909_21#_c_1046_n N_A_1909_21#_M1048_g N_A_1909_21#_M1002_g
+ N_A_1909_21#_c_1048_n N_A_1909_21#_M1053_g N_A_1909_21#_M1006_g
+ N_A_1909_21#_c_1050_n N_A_1909_21#_M1059_g N_A_1909_21#_M1008_g
+ N_A_1909_21#_c_1052_n N_A_1909_21#_M1060_g N_A_1909_21#_M1013_g
+ N_A_1909_21#_c_1054_n N_A_1909_21#_M1067_g N_A_1909_21#_M1023_g
+ N_A_1909_21#_c_1056_n N_A_1909_21#_M1073_g N_A_1909_21#_M1025_g
+ N_A_1909_21#_c_1058_n N_A_1909_21#_M1081_g N_A_1909_21#_M1026_g
+ N_A_1909_21#_c_1060_n N_A_1909_21#_M1086_g N_A_1909_21#_M1030_g
+ N_A_1909_21#_M1032_g N_A_1909_21#_M1038_g N_A_1909_21#_M1042_g
+ N_A_1909_21#_M1046_g N_A_1909_21#_M1050_g N_A_1909_21#_M1056_g
+ N_A_1909_21#_M1062_g N_A_1909_21#_M1063_g N_A_1909_21#_M1075_g
+ N_A_1909_21#_M1078_g N_A_1909_21#_M1088_g N_A_1909_21#_c_1073_n
+ N_A_1909_21#_c_1074_n N_A_1909_21#_c_1075_n N_A_1909_21#_c_1076_n
+ N_A_1909_21#_c_1077_n N_A_1909_21#_c_1078_n N_A_1909_21#_c_1079_n
+ N_A_1909_21#_c_1080_n N_A_1909_21#_c_1118_p N_A_1909_21#_c_1121_p
+ N_A_1909_21#_c_1103_n N_A_1909_21#_c_1139_p N_A_1909_21#_c_1129_p
+ N_A_1909_21#_c_1140_p N_A_1909_21#_c_1104_n N_A_1909_21#_c_1141_p
+ N_A_1909_21#_c_1145_p N_A_1909_21#_c_1105_n N_A_1909_21#_c_1158_p
+ N_A_1909_21#_c_1081_n N_A_1909_21#_c_1119_p N_A_1909_21#_c_1142_p
+ N_A_1909_21#_c_1106_n N_A_1909_21#_c_1107_n N_A_1909_21#_c_1082_n
+ PM_SKY130_FD_SC_LP__BUSDRIVER2_20%A_1909_21#
x_PM_SKY130_FD_SC_LP__BUSDRIVER2_20%A N_A_M1009_g N_A_c_1479_n N_A_c_1480_n
+ N_A_M1014_g N_A_c_1481_n N_A_M1028_g N_A_M1034_g N_A_c_1483_n N_A_M1029_g
+ N_A_M1052_g N_A_c_1485_n N_A_M1082_g N_A_M1072_g N_A_c_1487_n N_A_M1083_g
+ N_A_M1076_g N_A_M1079_g N_A_M1085_g A A A A A A N_A_c_1492_n
+ PM_SKY130_FD_SC_LP__BUSDRIVER2_20%A
x_PM_SKY130_FD_SC_LP__BUSDRIVER2_20%VPWR N_VPWR_M1004_d N_VPWR_M1007_d
+ N_VPWR_M1054_s N_VPWR_M1071_s N_VPWR_M1005_d N_VPWR_M1018_d N_VPWR_M1022_d
+ N_VPWR_M1040_d N_VPWR_M1055_d N_VPWR_M1061_d N_VPWR_M1065_d N_VPWR_M1074_d
+ N_VPWR_M1084_d N_VPWR_M1089_d N_VPWR_M1009_d N_VPWR_M1014_d N_VPWR_M1052_d
+ N_VPWR_M1076_d N_VPWR_M1085_d N_VPWR_c_1613_n N_VPWR_c_1614_n N_VPWR_c_1615_n
+ N_VPWR_c_1616_n N_VPWR_c_1617_n N_VPWR_c_1618_n N_VPWR_c_1619_n
+ N_VPWR_c_1620_n N_VPWR_c_1621_n N_VPWR_c_1622_n N_VPWR_c_1623_n
+ N_VPWR_c_1624_n N_VPWR_c_1625_n N_VPWR_c_1626_n N_VPWR_c_1627_n
+ N_VPWR_c_1628_n N_VPWR_c_1629_n N_VPWR_c_1630_n N_VPWR_c_1631_n
+ N_VPWR_c_1632_n N_VPWR_c_1633_n N_VPWR_c_1634_n N_VPWR_c_1635_n
+ N_VPWR_c_1636_n N_VPWR_c_1637_n N_VPWR_c_1638_n N_VPWR_c_1639_n
+ N_VPWR_c_1640_n N_VPWR_c_1641_n N_VPWR_c_1642_n N_VPWR_c_1643_n
+ N_VPWR_c_1644_n N_VPWR_c_1645_n N_VPWR_c_1646_n N_VPWR_c_1647_n
+ N_VPWR_c_1648_n N_VPWR_c_1649_n N_VPWR_c_1650_n N_VPWR_c_1651_n
+ N_VPWR_c_1652_n N_VPWR_c_1653_n N_VPWR_c_1654_n N_VPWR_c_1655_n
+ N_VPWR_c_1656_n N_VPWR_c_1657_n N_VPWR_c_1658_n N_VPWR_c_1659_n
+ N_VPWR_c_1660_n N_VPWR_c_1661_n N_VPWR_c_1662_n N_VPWR_c_1663_n
+ N_VPWR_c_1664_n VPWR N_VPWR_c_1665_n N_VPWR_c_1666_n N_VPWR_c_1667_n
+ N_VPWR_c_1668_n N_VPWR_c_1612_n PM_SKY130_FD_SC_LP__BUSDRIVER2_20%VPWR
x_PM_SKY130_FD_SC_LP__BUSDRIVER2_20%A_630_367# N_A_630_367#_M1001_s
+ N_A_630_367#_M1012_s N_A_630_367#_M1019_s N_A_630_367#_M1037_s
+ N_A_630_367#_M1041_s N_A_630_367#_M1058_s N_A_630_367#_M1064_s
+ N_A_630_367#_M1069_s N_A_630_367#_M1077_s N_A_630_367#_M1087_s
+ N_A_630_367#_M1000_s N_A_630_367#_M1006_s N_A_630_367#_M1013_s
+ N_A_630_367#_M1025_s N_A_630_367#_M1030_s N_A_630_367#_M1038_s
+ N_A_630_367#_M1046_s N_A_630_367#_M1056_s N_A_630_367#_M1063_s
+ N_A_630_367#_M1078_s N_A_630_367#_c_1959_n N_A_630_367#_c_1963_n
+ N_A_630_367#_c_1967_n N_A_630_367#_c_1971_n N_A_630_367#_c_1975_n
+ N_A_630_367#_c_1979_n N_A_630_367#_c_1983_n N_A_630_367#_c_1987_n
+ N_A_630_367#_c_1991_n N_A_630_367#_c_1999_n N_A_630_367#_c_1937_n
+ N_A_630_367#_c_1938_n N_A_630_367#_c_1939_n N_A_630_367#_c_2015_n
+ N_A_630_367#_c_1940_n N_A_630_367#_c_2072_n N_A_630_367#_c_2074_n
+ N_A_630_367#_c_1941_n N_A_630_367#_c_1942_n N_A_630_367#_c_2081_n
+ N_A_630_367#_c_1943_n N_A_630_367#_c_2087_n N_A_630_367#_c_1944_n
+ N_A_630_367#_c_2093_n N_A_630_367#_c_1945_n N_A_630_367#_c_2099_n
+ N_A_630_367#_c_1946_n N_A_630_367#_c_2105_n N_A_630_367#_c_1947_n
+ N_A_630_367#_c_2111_n N_A_630_367#_c_1948_n N_A_630_367#_c_2117_n
+ N_A_630_367#_c_1949_n N_A_630_367#_c_2123_n N_A_630_367#_c_1950_n
+ N_A_630_367#_c_2130_n N_A_630_367#_c_2017_n N_A_630_367#_c_2022_n
+ N_A_630_367#_c_2028_n N_A_630_367#_c_2034_n N_A_630_367#_c_2040_n
+ N_A_630_367#_c_2046_n N_A_630_367#_c_2052_n N_A_630_367#_c_2058_n
+ N_A_630_367#_c_2064_n N_A_630_367#_c_2066_n N_A_630_367#_c_1951_n
+ N_A_630_367#_c_1952_n N_A_630_367#_c_1953_n N_A_630_367#_c_1954_n
+ N_A_630_367#_c_1955_n N_A_630_367#_c_1956_n N_A_630_367#_c_1957_n
+ N_A_630_367#_c_1958_n PM_SKY130_FD_SC_LP__BUSDRIVER2_20%A_630_367#
x_PM_SKY130_FD_SC_LP__BUSDRIVER2_20%Z N_Z_M1017_s N_Z_M1027_s N_Z_M1033_s
+ N_Z_M1048_s N_Z_M1059_s N_Z_M1067_s N_Z_M1081_s N_Z_M1000_d N_Z_M1002_d
+ N_Z_M1008_d N_Z_M1023_d N_Z_M1026_d N_Z_M1032_d N_Z_M1042_d N_Z_M1050_d
+ N_Z_M1062_d N_Z_M1075_d N_Z_M1088_d N_Z_c_2279_n N_Z_c_2280_n N_Z_c_2283_n
+ N_Z_c_2421_n N_Z_c_2284_n N_Z_c_2424_n N_Z_c_2285_n N_Z_c_2427_n N_Z_c_2286_n
+ N_Z_c_2430_n N_Z_c_2287_n N_Z_c_2433_n N_Z_c_2288_n N_Z_c_2436_n N_Z_c_2289_n
+ N_Z_c_2439_n N_Z_c_2290_n N_Z_c_2442_n N_Z_c_2291_n N_Z_c_2445_n N_Z_c_2292_n
+ N_Z_c_2293_n N_Z_c_2294_n N_Z_c_2295_n N_Z_c_2296_n N_Z_c_2297_n N_Z_c_2298_n
+ N_Z_c_2299_n N_Z_c_2300_n N_Z_c_2301_n N_Z_c_2302_n N_Z_c_2303_n Z Z Z
+ N_Z_c_2281_n Z PM_SKY130_FD_SC_LP__BUSDRIVER2_20%Z
x_PM_SKY130_FD_SC_LP__BUSDRIVER2_20%VGND N_VGND_M1020_d N_VGND_M1024_d
+ N_VGND_M1043_d N_VGND_M1003_d N_VGND_M1015_d N_VGND_M1035_d N_VGND_M1044_d
+ N_VGND_M1047_d N_VGND_M1057_d N_VGND_M1070_d N_VGND_M1028_s N_VGND_M1029_s
+ N_VGND_M1083_s N_VGND_c_2479_n N_VGND_c_2480_n N_VGND_c_2481_n N_VGND_c_2482_n
+ N_VGND_c_2483_n N_VGND_c_2484_n N_VGND_c_2485_n N_VGND_c_2486_n
+ N_VGND_c_2487_n N_VGND_c_2488_n N_VGND_c_2489_n N_VGND_c_2490_n
+ N_VGND_c_2491_n N_VGND_c_2492_n N_VGND_c_2493_n N_VGND_c_2494_n
+ N_VGND_c_2495_n N_VGND_c_2496_n N_VGND_c_2497_n N_VGND_c_2498_n
+ N_VGND_c_2499_n N_VGND_c_2500_n N_VGND_c_2501_n N_VGND_c_2502_n
+ N_VGND_c_2503_n N_VGND_c_2504_n N_VGND_c_2505_n N_VGND_c_2506_n
+ N_VGND_c_2507_n N_VGND_c_2508_n N_VGND_c_2509_n N_VGND_c_2510_n VGND
+ N_VGND_c_2511_n N_VGND_c_2512_n N_VGND_c_2513_n N_VGND_c_2514_n
+ N_VGND_c_2515_n N_VGND_c_2516_n N_VGND_c_2517_n N_VGND_c_2518_n
+ PM_SKY130_FD_SC_LP__BUSDRIVER2_20%VGND
x_PM_SKY130_FD_SC_LP__BUSDRIVER2_20%A_584_47# N_A_584_47#_M1003_s
+ N_A_584_47#_M1011_s N_A_584_47#_M1016_s N_A_584_47#_M1039_s
+ N_A_584_47#_M1045_s N_A_584_47#_M1051_s N_A_584_47#_M1066_s
+ N_A_584_47#_M1080_s N_A_584_47#_M1021_d N_A_584_47#_M1031_d
+ N_A_584_47#_M1036_d N_A_584_47#_M1053_d N_A_584_47#_M1060_d
+ N_A_584_47#_M1073_d N_A_584_47#_M1086_d N_A_584_47#_c_2722_n
+ N_A_584_47#_c_2735_n N_A_584_47#_c_2723_n N_A_584_47#_c_2898_n
+ N_A_584_47#_c_2745_n N_A_584_47#_c_2905_n N_A_584_47#_c_2749_n
+ N_A_584_47#_c_2753_n N_A_584_47#_c_2757_n N_A_584_47#_c_2761_n
+ N_A_584_47#_c_2764_n N_A_584_47#_c_2724_n N_A_584_47#_c_2725_n
+ N_A_584_47#_c_2778_n N_A_584_47#_c_2726_n N_A_584_47#_c_2788_n
+ N_A_584_47#_c_2727_n N_A_584_47#_c_2797_n N_A_584_47#_c_2835_n
+ N_A_584_47#_c_2800_n N_A_584_47#_c_2801_n N_A_584_47#_c_2803_n
+ N_A_584_47#_c_2805_n N_A_584_47#_c_2809_n N_A_584_47#_c_2728_n
+ N_A_584_47#_c_2729_n N_A_584_47#_c_2730_n
+ PM_SKY130_FD_SC_LP__BUSDRIVER2_20%A_584_47#
cc_1 VNB N_TE_B_c_389_n 0.0209923f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.185
cc_2 VNB N_TE_B_M1004_g 0.011142f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.465
cc_3 VNB N_TE_B_c_391_n 0.0101534f $X=-0.19 $Y=-0.245 $X2=0.85 $Y2=1.26
cc_4 VNB N_TE_B_c_392_n 0.0176508f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.185
cc_5 VNB N_TE_B_M1007_g 0.0166613f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=2.465
cc_6 VNB N_TE_B_c_394_n 0.00626286f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.26
cc_7 VNB TE_B 0.00656339f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_8 VNB N_TE_B_c_396_n 0.0541886f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=1.35
cc_9 VNB N_A_114_47#_M1049_g 0.00884464f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=1.26
cc_10 VNB N_A_114_47#_M1010_g 0.0292988f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.335
cc_11 VNB N_A_114_47#_M1054_g 0.00718155f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=1.26
cc_12 VNB N_A_114_47#_c_432_n 0.0108772f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_114_47#_c_433_n 0.0257156f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=1.35
cc_14 VNB N_A_114_47#_M1043_g 0.0292403f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_114_47#_M1068_g 0.00795f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_114_47#_c_436_n 0.0133327f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_114_47#_M1071_g 0.00922759f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_114_47#_c_438_n 0.0228233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_114_47#_c_439_n 0.0240999f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_114_47#_c_440_n 0.0753264f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_114_47#_c_441_n 0.0167375f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_114_47#_c_442_n 0.0160063f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_114_47#_c_443_n 0.0160063f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_114_47#_c_444_n 0.0167375f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_114_47#_c_445_n 0.0240999f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_114_47#_c_446_n 0.0868403f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_114_47#_c_447_n 0.0169473f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_114_47#_c_448_n 0.0175844f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_114_47#_c_449_n 0.0201385f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_114_47#_c_450_n 0.0171229f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_114_47#_c_451_n 0.0101163f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_114_47#_c_452_n 0.0157257f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_114_47#_c_453_n 0.00948073f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_114_47#_c_454_n 0.0157257f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_114_47#_c_455_n 0.0101163f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_114_47#_c_456_n 0.0157257f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_114_47#_c_457_n 0.00948073f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_114_47#_c_458_n 0.0157257f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_114_47#_c_459_n 0.0101163f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_114_47#_c_460_n 0.0157257f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_114_47#_c_461_n 0.0153631f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_114_47#_c_462_n 0.0157866f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_114_47#_c_463_n 0.00416623f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_114_47#_c_464_n 0.00476283f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_114_47#_c_465_n 0.00390043f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_114_47#_c_466_n 0.00390043f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_114_47#_c_467_n 0.00390043f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_114_47#_c_468_n 0.00390043f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_114_47#_c_469_n 0.00390043f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_114_47#_c_470_n 0.0080712f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_114_47#_c_471_n 0.0122581f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_114_47#_c_472_n 0.0432044f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_286_367#_c_704_n 0.00558275f $X=-0.19 $Y=-0.245 $X2=0.925
+ $Y2=1.335
cc_54 VNB N_A_286_367#_c_705_n 0.00407356f $X=-0.19 $Y=-0.245 $X2=0.925
+ $Y2=2.465
cc_55 VNB N_A_286_367#_c_706_n 0.00558275f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_56 VNB N_A_286_367#_c_707_n 0.00558275f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_286_367#_c_708_n 0.00558275f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_286_367#_c_709_n 0.00558275f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_286_367#_c_710_n 0.00558275f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_286_367#_c_711_n 0.00558275f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_A_286_367#_c_712_n 0.00619686f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_A_286_367#_c_713_n 0.00747967f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_A_286_367#_c_714_n 0.193431f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_A_286_367#_c_715_n 0.0075543f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_A_286_367#_c_716_n 0.0151222f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_A_286_367#_c_717_n 0.00300943f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_A_286_367#_c_718_n 0.00300943f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_A_286_367#_c_719_n 0.00300943f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_286_367#_c_720_n 0.00300943f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_A_286_367#_c_721_n 0.00300943f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_A_286_367#_c_722_n 0.00300943f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_A_286_367#_c_723_n 0.00308029f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_A_286_367#_c_724_n 0.00405366f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_A_286_367#_c_725_n 0.00405366f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_A_286_367#_c_726_n 0.00716792f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_A_286_367#_c_727_n 0.00688294f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_A_286_367#_c_728_n 0.00602717f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_A_286_367#_c_729_n 0.00232232f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_A_286_367#_c_730_n 0.0238032f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_A_1909_21#_c_1033_n 0.0165263f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_A_1909_21#_c_1034_n 0.0178584f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=1.35
cc_82 VNB N_A_1909_21#_c_1035_n 0.00674478f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_A_1909_21#_c_1036_n 0.0174693f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.35
cc_84 VNB N_A_1909_21#_c_1037_n 0.0184839f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_A_1909_21#_c_1038_n 0.0174526f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_A_1909_21#_c_1039_n 0.0184838f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_A_1909_21#_c_1040_n 0.016696f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_A_1909_21#_c_1041_n 0.0146842f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_A_1909_21#_c_1042_n 0.0152249f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_A_1909_21#_c_1043_n 0.0152334f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_A_1909_21#_c_1044_n 0.0152249f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_A_1909_21#_M1000_g 0.00117852f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_93 VNB N_A_1909_21#_c_1046_n 0.0159623f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_94 VNB N_A_1909_21#_M1002_g 9.64739e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_95 VNB N_A_1909_21#_c_1048_n 0.0159844f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_96 VNB N_A_1909_21#_M1006_g 9.66271e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_97 VNB N_A_1909_21#_c_1050_n 0.0160041f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_98 VNB N_A_1909_21#_M1008_g 9.66271e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_99 VNB N_A_1909_21#_c_1052_n 0.0160041f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_100 VNB N_A_1909_21#_M1013_g 9.66271e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_101 VNB N_A_1909_21#_c_1054_n 0.0160041f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_102 VNB N_A_1909_21#_M1023_g 9.66271e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_103 VNB N_A_1909_21#_c_1056_n 0.0160041f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_104 VNB N_A_1909_21#_M1025_g 9.66271e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_105 VNB N_A_1909_21#_c_1058_n 0.0160041f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_106 VNB N_A_1909_21#_M1026_g 9.66271e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_107 VNB N_A_1909_21#_c_1060_n 0.0219859f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_108 VNB N_A_1909_21#_M1030_g 9.66271e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_109 VNB N_A_1909_21#_M1032_g 9.66271e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_110 VNB N_A_1909_21#_M1038_g 9.66271e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_111 VNB N_A_1909_21#_M1042_g 9.66271e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_112 VNB N_A_1909_21#_M1046_g 9.66271e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_113 VNB N_A_1909_21#_M1050_g 9.66271e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_114 VNB N_A_1909_21#_M1056_g 9.66271e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_115 VNB N_A_1909_21#_M1062_g 9.66271e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_116 VNB N_A_1909_21#_M1063_g 0.00147483f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_117 VNB N_A_1909_21#_M1075_g 0.00147483f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_118 VNB N_A_1909_21#_M1078_g 0.00147483f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_119 VNB N_A_1909_21#_M1088_g 0.00233375f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_120 VNB N_A_1909_21#_c_1073_n 0.00621252f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_121 VNB N_A_1909_21#_c_1074_n 0.00621279f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_122 VNB N_A_1909_21#_c_1075_n 0.00624721f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_123 VNB N_A_1909_21#_c_1076_n 0.00666874f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_124 VNB N_A_1909_21#_c_1077_n 0.00165135f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_125 VNB N_A_1909_21#_c_1078_n 0.00236419f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_126 VNB N_A_1909_21#_c_1079_n 0.115373f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_127 VNB N_A_1909_21#_c_1080_n 0.00880557f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_128 VNB N_A_1909_21#_c_1081_n 0.00972274f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_129 VNB N_A_1909_21#_c_1082_n 0.650059f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_130 VNB N_A_c_1479_n 0.011419f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.465
cc_131 VNB N_A_c_1480_n 0.00833265f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.465
cc_132 VNB N_A_c_1481_n 0.0191729f $X=-0.19 $Y=-0.245 $X2=0.925 $Y2=0.655
cc_133 VNB N_A_M1034_g 0.00706566f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_134 VNB N_A_c_1483_n 0.0181593f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_135 VNB N_A_M1052_g 0.00706903f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_136 VNB N_A_c_1485_n 0.017472f $X=-0.19 $Y=-0.245 $X2=0.57 $Y2=1.35
cc_137 VNB N_A_M1072_g 0.00706903f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_138 VNB N_A_c_1487_n 0.0218877f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_139 VNB N_A_M1076_g 0.00721043f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_140 VNB N_A_M1079_g 0.00721043f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_141 VNB N_A_M1085_g 0.0111859f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_142 VNB A 0.0719111f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_143 VNB N_A_c_1492_n 0.18018f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_144 VNB N_VPWR_c_1612_n 1.03939f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_145 VNB N_A_630_367#_c_1937_n 0.00905481f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_146 VNB N_A_630_367#_c_1938_n 0.00426187f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_147 VNB N_Z_c_2279_n 0.0126176f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_148 VNB N_Z_c_2280_n 0.0176881f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_149 VNB N_Z_c_2281_n 0.00182111f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_150 VNB Z 0.0194829f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_151 VNB N_VGND_c_2479_n 0.0110036f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_152 VNB N_VGND_c_2480_n 0.0316927f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_153 VNB N_VGND_c_2481_n 0.00480599f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_154 VNB N_VGND_c_2482_n 0.0068991f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_155 VNB N_VGND_c_2483_n 0.00274299f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_156 VNB N_VGND_c_2484_n 3.0911e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_157 VNB N_VGND_c_2485_n 0.00274299f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_158 VNB N_VGND_c_2486_n 0.00561774f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_159 VNB N_VGND_c_2487_n 0.0047158f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_160 VNB N_VGND_c_2488_n 0.0047158f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_161 VNB N_VGND_c_2489_n 0.0047158f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_162 VNB N_VGND_c_2490_n 0.0185692f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_163 VNB N_VGND_c_2491_n 0.00561774f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_164 VNB N_VGND_c_2492_n 0.0345543f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_165 VNB N_VGND_c_2493_n 0.0260059f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_166 VNB N_VGND_c_2494_n 0.00631318f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_167 VNB N_VGND_c_2495_n 0.0116044f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_168 VNB N_VGND_c_2496_n 0.00436214f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_169 VNB N_VGND_c_2497_n 0.0116044f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_170 VNB N_VGND_c_2498_n 0.00510188f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_171 VNB N_VGND_c_2499_n 0.0173134f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_172 VNB N_VGND_c_2500_n 0.00631504f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_173 VNB N_VGND_c_2501_n 0.0180904f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_174 VNB N_VGND_c_2502_n 0.00326991f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_175 VNB N_VGND_c_2503_n 0.0188675f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_176 VNB N_VGND_c_2504_n 0.00326991f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_177 VNB N_VGND_c_2505_n 0.0188675f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_178 VNB N_VGND_c_2506_n 0.00326991f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_179 VNB N_VGND_c_2507_n 0.335017f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_180 VNB N_VGND_c_2508_n 0.0051639f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_181 VNB N_VGND_c_2509_n 0.0179931f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_182 VNB N_VGND_c_2510_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_183 VNB N_VGND_c_2511_n 0.0155644f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_184 VNB N_VGND_c_2512_n 0.0196816f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_185 VNB N_VGND_c_2513_n 0.0188675f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_186 VNB N_VGND_c_2514_n 0.0361928f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_187 VNB N_VGND_c_2515_n 1.37015f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_188 VNB N_VGND_c_2516_n 0.00631318f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_189 VNB N_VGND_c_2517_n 0.00510188f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_190 VNB N_VGND_c_2518_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_191 VNB N_A_584_47#_c_2722_n 0.00515289f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_192 VNB N_A_584_47#_c_2723_n 0.00232859f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_193 VNB N_A_584_47#_c_2724_n 0.00324175f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_194 VNB N_A_584_47#_c_2725_n 0.00240609f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_195 VNB N_A_584_47#_c_2726_n 0.00324175f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_196 VNB N_A_584_47#_c_2727_n 0.00653461f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_197 VNB N_A_584_47#_c_2728_n 0.00207104f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_198 VNB N_A_584_47#_c_2729_n 0.00207104f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_199 VNB N_A_584_47#_c_2730_n 0.0207635f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_200 VPB N_TE_B_M1004_g 0.0264715f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=2.465
cc_201 VPB N_TE_B_M1007_g 0.0197283f $X=-0.19 $Y=1.655 $X2=0.925 $Y2=2.465
cc_202 VPB N_A_114_47#_M1049_g 0.02002f $X=-0.19 $Y=1.655 $X2=0.57 $Y2=1.26
cc_203 VPB N_A_114_47#_M1054_g 0.018242f $X=-0.19 $Y=1.655 $X2=0.925 $Y2=1.26
cc_204 VPB N_A_114_47#_M1068_g 0.0188806f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_205 VPB N_A_114_47#_M1071_g 0.019225f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_206 VPB N_A_114_47#_c_470_n 0.00424242f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_207 VPB N_A_286_367#_c_731_n 0.016435f $X=-0.19 $Y=1.655 $X2=0.925 $Y2=1.185
cc_208 VPB N_A_286_367#_c_704_n 0.0042584f $X=-0.19 $Y=1.655 $X2=0.925 $Y2=1.335
cc_209 VPB N_A_286_367#_c_705_n 0.00231877f $X=-0.19 $Y=1.655 $X2=0.925
+ $Y2=2.465
cc_210 VPB N_A_286_367#_c_734_n 0.0162054f $X=-0.19 $Y=1.655 $X2=0.925 $Y2=2.465
cc_211 VPB N_A_286_367#_c_706_n 0.00425948f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_212 VPB N_A_286_367#_c_736_n 0.0162054f $X=-0.19 $Y=1.655 $X2=0.28 $Y2=1.35
cc_213 VPB N_A_286_367#_c_707_n 0.0042584f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_214 VPB N_A_286_367#_c_738_n 0.0162054f $X=-0.19 $Y=1.655 $X2=0.57 $Y2=1.35
cc_215 VPB N_A_286_367#_c_708_n 0.00425948f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_216 VPB N_A_286_367#_c_740_n 0.0162054f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_217 VPB N_A_286_367#_c_709_n 0.0042584f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_218 VPB N_A_286_367#_c_742_n 0.0162054f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_219 VPB N_A_286_367#_c_710_n 0.00425948f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_220 VPB N_A_286_367#_c_744_n 0.0162054f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_221 VPB N_A_286_367#_c_711_n 0.0042584f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_222 VPB N_A_286_367#_c_746_n 0.0162054f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_223 VPB N_A_286_367#_c_712_n 0.00388803f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_224 VPB N_A_286_367#_c_748_n 0.0162054f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_225 VPB N_A_286_367#_c_749_n 0.0162054f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_226 VPB N_A_286_367#_c_750_n 0.0162054f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_227 VPB N_A_286_367#_c_751_n 0.0164005f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_228 VPB N_A_286_367#_c_752_n 0.0164005f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_229 VPB N_A_286_367#_c_753_n 0.0162054f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_230 VPB N_A_286_367#_c_754_n 0.0162054f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_231 VPB N_A_286_367#_c_755_n 0.0161974f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_232 VPB N_A_286_367#_c_756_n 0.0157337f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_233 VPB N_A_286_367#_c_713_n 0.0049292f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_234 VPB N_A_286_367#_c_714_n 0.0469051f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_235 VPB N_A_286_367#_c_759_n 0.0157208f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_236 VPB N_A_286_367#_c_715_n 0.00421299f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_237 VPB N_A_286_367#_c_761_n 0.0157208f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_238 VPB N_A_286_367#_c_716_n 0.00804128f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_239 VPB N_A_286_367#_c_763_n 0.0201845f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_240 VPB N_A_286_367#_c_717_n 0.00111435f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_241 VPB N_A_286_367#_c_718_n 0.00111435f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_242 VPB N_A_286_367#_c_719_n 0.00111435f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_243 VPB N_A_286_367#_c_720_n 0.00111435f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_244 VPB N_A_286_367#_c_721_n 0.00111435f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_245 VPB N_A_286_367#_c_722_n 0.00111435f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_246 VPB N_A_286_367#_c_723_n 0.00111435f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_247 VPB N_A_286_367#_c_724_n 0.00111435f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_248 VPB N_A_286_367#_c_725_n 0.00111435f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_249 VPB N_A_286_367#_c_726_n 0.00311423f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_250 VPB N_A_286_367#_c_774_n 0.00351925f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_251 VPB N_A_286_367#_c_775_n 0.00674711f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_252 VPB N_A_286_367#_c_730_n 0.00538792f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_253 VPB N_A_1909_21#_M1000_g 0.0229316f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_254 VPB N_A_1909_21#_M1002_g 0.0190671f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_255 VPB N_A_1909_21#_M1006_g 0.0190975f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_256 VPB N_A_1909_21#_M1008_g 0.0190975f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_257 VPB N_A_1909_21#_M1013_g 0.0190975f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_258 VPB N_A_1909_21#_M1023_g 0.0190975f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_259 VPB N_A_1909_21#_M1025_g 0.0190975f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_260 VPB N_A_1909_21#_M1026_g 0.0190975f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_261 VPB N_A_1909_21#_M1030_g 0.0190796f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_262 VPB N_A_1909_21#_M1032_g 0.0190769f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_263 VPB N_A_1909_21#_M1038_g 0.0190139f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_264 VPB N_A_1909_21#_M1042_g 0.0190139f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_265 VPB N_A_1909_21#_M1046_g 0.0190139f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_266 VPB N_A_1909_21#_M1050_g 0.0190139f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_267 VPB N_A_1909_21#_M1056_g 0.0190139f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_268 VPB N_A_1909_21#_M1062_g 0.0190139f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_269 VPB N_A_1909_21#_M1063_g 0.0190139f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_270 VPB N_A_1909_21#_M1075_g 0.0190139f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_271 VPB N_A_1909_21#_M1078_g 0.0190139f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_272 VPB N_A_1909_21#_M1088_g 0.0255127f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_273 VPB N_A_1909_21#_c_1103_n 0.00229974f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_274 VPB N_A_1909_21#_c_1104_n 0.00229974f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_275 VPB N_A_1909_21#_c_1105_n 0.00480442f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_276 VPB N_A_1909_21#_c_1106_n 0.00235119f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_277 VPB N_A_1909_21#_c_1107_n 0.00235119f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_278 VPB N_A_M1009_g 0.0206394f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=0.655
cc_279 VPB N_A_c_1479_n 0.00433912f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=2.465
cc_280 VPB N_A_c_1480_n 0.00245547f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=2.465
cc_281 VPB N_A_M1014_g 0.0161014f $X=-0.19 $Y=1.655 $X2=0.57 $Y2=1.26
cc_282 VPB N_A_M1034_g 0.0185888f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_283 VPB N_A_M1052_g 0.0186072f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_284 VPB N_A_M1072_g 0.0186072f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_285 VPB N_A_M1076_g 0.0189208f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_286 VPB N_A_M1079_g 0.0189208f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_287 VPB N_A_M1085_g 0.0266775f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_288 VPB N_A_c_1492_n 0.00163176f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_289 VPB N_VPWR_c_1613_n 0.0109777f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_290 VPB N_VPWR_c_1614_n 0.0536171f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_291 VPB N_VPWR_c_1615_n 0.0115599f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_292 VPB N_VPWR_c_1616_n 0.0047158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_293 VPB N_VPWR_c_1617_n 0.0047158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_294 VPB N_VPWR_c_1618_n 0.00430763f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_295 VPB N_VPWR_c_1619_n 0.0195793f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_296 VPB N_VPWR_c_1620_n 0.00378659f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_297 VPB N_VPWR_c_1621_n 0.00378659f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_298 VPB N_VPWR_c_1622_n 0.00378659f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_299 VPB N_VPWR_c_1623_n 0.00378659f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_300 VPB N_VPWR_c_1624_n 0.00432085f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_301 VPB N_VPWR_c_1625_n 0.0202158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_302 VPB N_VPWR_c_1626_n 0.00430763f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_303 VPB N_VPWR_c_1627_n 0.00426383f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_304 VPB N_VPWR_c_1628_n 0.00563092f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_305 VPB N_VPWR_c_1629_n 0.0138665f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_306 VPB N_VPWR_c_1630_n 0.0218485f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_307 VPB N_VPWR_c_1631_n 0.0047158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_308 VPB N_VPWR_c_1632_n 0.0047158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_309 VPB N_VPWR_c_1633_n 0.0188675f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_310 VPB N_VPWR_c_1634_n 0.00472864f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_311 VPB N_VPWR_c_1635_n 0.0106521f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_312 VPB N_VPWR_c_1636_n 0.055403f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_313 VPB N_VPWR_c_1637_n 0.0131585f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_314 VPB N_VPWR_c_1638_n 0.00356964f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_315 VPB N_VPWR_c_1639_n 0.0188675f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_316 VPB N_VPWR_c_1640_n 0.00324402f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_317 VPB N_VPWR_c_1641_n 0.0188675f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_318 VPB N_VPWR_c_1642_n 0.00324402f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_319 VPB N_VPWR_c_1643_n 0.0198976f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_320 VPB N_VPWR_c_1644_n 0.00362871f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_321 VPB N_VPWR_c_1645_n 0.0195793f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_322 VPB N_VPWR_c_1646_n 0.00362871f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_323 VPB N_VPWR_c_1647_n 0.0195793f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_324 VPB N_VPWR_c_1648_n 0.00362871f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_325 VPB N_VPWR_c_1649_n 0.0195793f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_326 VPB N_VPWR_c_1650_n 0.00362871f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_327 VPB N_VPWR_c_1651_n 0.0195793f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_328 VPB N_VPWR_c_1652_n 0.00362871f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_329 VPB N_VPWR_c_1653_n 0.0195793f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_330 VPB N_VPWR_c_1654_n 0.00362871f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_331 VPB N_VPWR_c_1655_n 0.0185493f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_332 VPB N_VPWR_c_1656_n 0.00324402f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_333 VPB N_VPWR_c_1657_n 0.016013f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_334 VPB N_VPWR_c_1658_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_335 VPB N_VPWR_c_1659_n 0.223484f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_336 VPB N_VPWR_c_1660_n 0.0047828f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_337 VPB N_VPWR_c_1661_n 0.0188675f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_338 VPB N_VPWR_c_1662_n 0.00324402f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_339 VPB N_VPWR_c_1663_n 0.0188675f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_340 VPB N_VPWR_c_1664_n 0.00324402f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_341 VPB N_VPWR_c_1665_n 0.0196631f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_342 VPB N_VPWR_c_1666_n 0.00362871f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_343 VPB N_VPWR_c_1667_n 0.00362871f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_344 VPB N_VPWR_c_1668_n 0.00324402f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_345 VPB N_VPWR_c_1612_n 0.159044f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_346 VPB N_A_630_367#_c_1939_n 8.34152e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_347 VPB N_A_630_367#_c_1940_n 0.0146648f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_348 VPB N_A_630_367#_c_1941_n 0.00873754f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_349 VPB N_A_630_367#_c_1942_n 0.00505735f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_350 VPB N_A_630_367#_c_1943_n 0.00873754f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_351 VPB N_A_630_367#_c_1944_n 0.00873754f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_352 VPB N_A_630_367#_c_1945_n 0.00873754f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_353 VPB N_A_630_367#_c_1946_n 0.00873754f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_354 VPB N_A_630_367#_c_1947_n 0.00873754f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_355 VPB N_A_630_367#_c_1948_n 0.00873754f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_356 VPB N_A_630_367#_c_1949_n 0.00873754f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_357 VPB N_A_630_367#_c_1950_n 0.0137644f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_358 VPB N_A_630_367#_c_1951_n 0.00244498f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_359 VPB N_A_630_367#_c_1952_n 0.00244498f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_360 VPB N_A_630_367#_c_1953_n 0.00244498f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_361 VPB N_A_630_367#_c_1954_n 0.00244498f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_362 VPB N_A_630_367#_c_1955_n 0.00244498f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_363 VPB N_A_630_367#_c_1956_n 0.00244498f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_364 VPB N_A_630_367#_c_1957_n 0.00244498f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_365 VPB N_A_630_367#_c_1958_n 0.00244498f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_366 VPB N_Z_c_2283_n 0.00302716f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_367 VPB N_Z_c_2284_n 0.00313797f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_368 VPB N_Z_c_2285_n 0.00313797f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_369 VPB N_Z_c_2286_n 0.00313718f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_370 VPB N_Z_c_2287_n 0.00319476f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_371 VPB N_Z_c_2288_n 0.00313758f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_372 VPB N_Z_c_2289_n 0.00313758f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_373 VPB N_Z_c_2290_n 0.00313758f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_374 VPB N_Z_c_2291_n 0.0031404f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_375 VPB N_Z_c_2292_n 0.00305943f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_376 VPB N_Z_c_2293_n 0.00503673f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_377 VPB N_Z_c_2294_n 0.0129834f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_378 VPB N_Z_c_2295_n 0.00148939f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_379 VPB N_Z_c_2296_n 0.00148939f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_380 VPB N_Z_c_2297_n 0.00148939f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_381 VPB N_Z_c_2298_n 0.00150456f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_382 VPB N_Z_c_2299_n 0.00159601f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_383 VPB N_Z_c_2300_n 0.00148653f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_384 VPB N_Z_c_2301_n 0.00148653f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_385 VPB N_Z_c_2302_n 0.00148939f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_386 VPB N_Z_c_2303_n 0.00148939f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_387 VPB N_Z_c_2281_n 0.00833748f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_388 N_TE_B_c_392_n N_A_114_47#_M1010_g 0.0317687f $X=0.925 $Y=1.185 $X2=0
+ $Y2=0
cc_389 N_TE_B_M1007_g N_A_114_47#_c_433_n 0.0362432f $X=0.925 $Y=2.465 $X2=0
+ $Y2=0
cc_390 N_TE_B_c_389_n N_A_114_47#_c_470_n 0.00251768f $X=0.495 $Y=1.185 $X2=0
+ $Y2=0
cc_391 N_TE_B_c_391_n N_A_114_47#_c_470_n 0.012108f $X=0.85 $Y=1.26 $X2=0 $Y2=0
cc_392 N_TE_B_c_392_n N_A_114_47#_c_470_n 0.00260132f $X=0.925 $Y=1.185 $X2=0
+ $Y2=0
cc_393 N_TE_B_M1007_g N_A_114_47#_c_470_n 0.0121802f $X=0.925 $Y=2.465 $X2=0
+ $Y2=0
cc_394 TE_B N_A_114_47#_c_470_n 0.0235118f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_395 N_TE_B_c_396_n N_A_114_47#_c_470_n 0.00938712f $X=0.57 $Y=1.35 $X2=0
+ $Y2=0
cc_396 N_TE_B_c_392_n N_A_114_47#_c_486_n 0.0160662f $X=0.925 $Y=1.185 $X2=0
+ $Y2=0
cc_397 N_TE_B_M1007_g N_A_286_367#_c_777_n 4.08568e-19 $X=0.925 $Y=2.465 $X2=0
+ $Y2=0
cc_398 N_TE_B_M1007_g N_A_286_367#_c_726_n 4.58855e-19 $X=0.925 $Y=2.465 $X2=0
+ $Y2=0
cc_399 N_TE_B_M1004_g N_VPWR_c_1614_n 0.0228515f $X=0.495 $Y=2.465 $X2=0 $Y2=0
cc_400 N_TE_B_M1007_g N_VPWR_c_1614_n 8.30776e-19 $X=0.925 $Y=2.465 $X2=0 $Y2=0
cc_401 TE_B N_VPWR_c_1614_n 0.0180868f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_402 N_TE_B_c_396_n N_VPWR_c_1614_n 0.00224381f $X=0.57 $Y=1.35 $X2=0 $Y2=0
cc_403 N_TE_B_M1004_g N_VPWR_c_1615_n 8.27214e-19 $X=0.495 $Y=2.465 $X2=0 $Y2=0
cc_404 N_TE_B_M1007_g N_VPWR_c_1615_n 0.0198517f $X=0.925 $Y=2.465 $X2=0 $Y2=0
cc_405 N_TE_B_M1004_g N_VPWR_c_1637_n 0.00486043f $X=0.495 $Y=2.465 $X2=0 $Y2=0
cc_406 N_TE_B_M1007_g N_VPWR_c_1637_n 0.00486043f $X=0.925 $Y=2.465 $X2=0 $Y2=0
cc_407 N_TE_B_M1004_g N_VPWR_c_1612_n 0.00824727f $X=0.495 $Y=2.465 $X2=0 $Y2=0
cc_408 N_TE_B_M1007_g N_VPWR_c_1612_n 0.00824727f $X=0.925 $Y=2.465 $X2=0 $Y2=0
cc_409 N_TE_B_c_389_n N_VGND_c_2480_n 0.0146496f $X=0.495 $Y=1.185 $X2=0 $Y2=0
cc_410 N_TE_B_c_392_n N_VGND_c_2480_n 7.00016e-19 $X=0.925 $Y=1.185 $X2=0 $Y2=0
cc_411 TE_B N_VGND_c_2480_n 0.0247917f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_412 N_TE_B_c_396_n N_VGND_c_2480_n 0.00217868f $X=0.57 $Y=1.35 $X2=0 $Y2=0
cc_413 N_TE_B_c_392_n N_VGND_c_2481_n 0.00300298f $X=0.925 $Y=1.185 $X2=0 $Y2=0
cc_414 N_TE_B_c_389_n N_VGND_c_2511_n 0.00486043f $X=0.495 $Y=1.185 $X2=0 $Y2=0
cc_415 N_TE_B_c_392_n N_VGND_c_2511_n 0.0042361f $X=0.925 $Y=1.185 $X2=0 $Y2=0
cc_416 N_TE_B_c_389_n N_VGND_c_2515_n 0.00824727f $X=0.495 $Y=1.185 $X2=0 $Y2=0
cc_417 N_TE_B_c_392_n N_VGND_c_2515_n 0.00619616f $X=0.925 $Y=1.185 $X2=0 $Y2=0
cc_418 N_A_114_47#_c_486_n N_A_286_367#_M1010_s 0.0140131f $X=2.19 $Y=0.71
+ $X2=-0.19 $Y2=-0.245
cc_419 N_A_114_47#_M1071_g N_A_286_367#_c_705_n 0.023821f $X=2.645 $Y=2.465
+ $X2=0 $Y2=0
cc_420 N_A_114_47#_c_440_n N_A_286_367#_c_705_n 0.034655f $X=3.355 $Y=1.16 $X2=0
+ $Y2=0
cc_421 N_A_114_47#_c_471_n N_A_286_367#_c_705_n 0.00353499f $X=5.985 $Y=1.17
+ $X2=0 $Y2=0
cc_422 N_A_114_47#_c_439_n N_A_286_367#_c_706_n 0.034655f $X=3.715 $Y=1.16 $X2=0
+ $Y2=0
cc_423 N_A_114_47#_c_445_n N_A_286_367#_c_709_n 0.034655f $X=5.515 $Y=1.16 $X2=0
+ $Y2=0
cc_424 N_A_114_47#_c_449_n N_A_286_367#_c_714_n 0.190078f $X=6.535 $Y=1.06 $X2=0
+ $Y2=0
cc_425 N_A_114_47#_c_446_n N_A_286_367#_c_719_n 0.034655f $X=5.155 $Y=1.16 $X2=0
+ $Y2=0
cc_426 N_A_114_47#_c_472_n N_A_286_367#_c_722_n 0.034655f $X=6.15 $Y=1.16 $X2=0
+ $Y2=0
cc_427 N_A_114_47#_c_449_n N_A_286_367#_c_723_n 0.00548024f $X=6.535 $Y=1.06
+ $X2=0 $Y2=0
cc_428 N_A_114_47#_M1049_g N_A_286_367#_c_777_n 0.0131962f $X=1.355 $Y=2.465
+ $X2=0 $Y2=0
cc_429 N_A_114_47#_M1054_g N_A_286_367#_c_777_n 0.0144071f $X=1.785 $Y=2.465
+ $X2=0 $Y2=0
cc_430 N_A_114_47#_M1068_g N_A_286_367#_c_777_n 7.33648e-19 $X=2.215 $Y=2.465
+ $X2=0 $Y2=0
cc_431 N_A_114_47#_M1049_g N_A_286_367#_c_726_n 0.00705968f $X=1.355 $Y=2.465
+ $X2=0 $Y2=0
cc_432 N_A_114_47#_M1010_g N_A_286_367#_c_726_n 0.0102673f $X=1.515 $Y=0.655
+ $X2=0 $Y2=0
cc_433 N_A_114_47#_M1054_g N_A_286_367#_c_726_n 0.00882374f $X=1.785 $Y=2.465
+ $X2=0 $Y2=0
cc_434 N_A_114_47#_c_432_n N_A_286_367#_c_726_n 0.0135737f $X=2.1 $Y=1.41 $X2=0
+ $Y2=0
cc_435 N_A_114_47#_c_433_n N_A_286_367#_c_726_n 0.00953885f $X=1.86 $Y=1.41
+ $X2=0 $Y2=0
cc_436 N_A_114_47#_M1043_g N_A_286_367#_c_726_n 0.00347031f $X=2.175 $Y=0.655
+ $X2=0 $Y2=0
cc_437 N_A_114_47#_M1068_g N_A_286_367#_c_726_n 0.00302226f $X=2.215 $Y=2.465
+ $X2=0 $Y2=0
cc_438 N_A_114_47#_c_486_n N_A_286_367#_c_726_n 0.0255687f $X=2.19 $Y=0.71 $X2=0
+ $Y2=0
cc_439 N_A_114_47#_c_508_p N_A_286_367#_c_726_n 0.00209179f $X=2.275 $Y=1.005
+ $X2=0 $Y2=0
cc_440 N_A_114_47#_c_509_p N_A_286_367#_c_726_n 0.0263669f $X=2.36 $Y=1.17 $X2=0
+ $Y2=0
cc_441 N_A_114_47#_c_432_n N_A_286_367#_c_774_n 0.00139964f $X=2.1 $Y=1.41 $X2=0
+ $Y2=0
cc_442 N_A_114_47#_M1068_g N_A_286_367#_c_774_n 0.0145139f $X=2.215 $Y=2.465
+ $X2=0 $Y2=0
cc_443 N_A_114_47#_c_509_p N_A_286_367#_c_774_n 0.00245801f $X=2.36 $Y=1.17
+ $X2=0 $Y2=0
cc_444 N_A_114_47#_M1049_g N_A_286_367#_c_775_n 0.00307365f $X=1.355 $Y=2.465
+ $X2=0 $Y2=0
cc_445 N_A_114_47#_M1054_g N_A_286_367#_c_775_n 0.0106988f $X=1.785 $Y=2.465
+ $X2=0 $Y2=0
cc_446 N_A_114_47#_c_433_n N_A_286_367#_c_775_n 0.00350003f $X=1.86 $Y=1.41
+ $X2=0 $Y2=0
cc_447 N_A_114_47#_M1068_g N_A_286_367#_c_808_n 0.0143171f $X=2.215 $Y=2.465
+ $X2=0 $Y2=0
cc_448 N_A_114_47#_M1071_g N_A_286_367#_c_808_n 0.0130438f $X=2.645 $Y=2.465
+ $X2=0 $Y2=0
cc_449 N_A_114_47#_c_449_n N_A_286_367#_c_727_n 6.17508e-19 $X=6.535 $Y=1.06
+ $X2=0 $Y2=0
cc_450 N_A_114_47#_c_464_n N_A_286_367#_c_728_n 0.00368497f $X=6.61 $Y=1.06
+ $X2=0 $Y2=0
cc_451 N_A_114_47#_M1054_g N_A_286_367#_c_729_n 0.00107404f $X=1.785 $Y=2.465
+ $X2=0 $Y2=0
cc_452 N_A_114_47#_M1068_g N_A_286_367#_c_729_n 0.00867585f $X=2.215 $Y=2.465
+ $X2=0 $Y2=0
cc_453 N_A_114_47#_c_436_n N_A_286_367#_c_729_n 0.00240029f $X=2.57 $Y=1.41
+ $X2=0 $Y2=0
cc_454 N_A_114_47#_M1071_g N_A_286_367#_c_729_n 0.0095353f $X=2.645 $Y=2.465
+ $X2=0 $Y2=0
cc_455 N_A_114_47#_c_509_p N_A_286_367#_c_729_n 0.00790072f $X=2.36 $Y=1.17
+ $X2=0 $Y2=0
cc_456 N_A_114_47#_c_471_n N_A_286_367#_c_729_n 0.0196176f $X=5.985 $Y=1.17
+ $X2=0 $Y2=0
cc_457 N_A_114_47#_M1071_g N_A_286_367#_c_730_n 0.0129368f $X=2.645 $Y=2.465
+ $X2=0 $Y2=0
cc_458 N_A_114_47#_c_440_n N_A_286_367#_c_730_n 0.0255384f $X=3.355 $Y=1.16
+ $X2=0 $Y2=0
cc_459 N_A_114_47#_c_449_n N_A_286_367#_c_730_n 0.00417271f $X=6.535 $Y=1.06
+ $X2=0 $Y2=0
cc_460 N_A_114_47#_c_471_n N_A_286_367#_c_730_n 0.255303f $X=5.985 $Y=1.17 $X2=0
+ $Y2=0
cc_461 N_A_114_47#_c_462_n N_A_1909_21#_c_1033_n 0.014832f $X=9.19 $Y=0.985
+ $X2=0 $Y2=0
cc_462 N_A_114_47#_c_461_n N_A_1909_21#_c_1035_n 0.014832f $X=9.115 $Y=1.06
+ $X2=0 $Y2=0
cc_463 N_A_114_47#_c_470_n N_VPWR_c_1614_n 0.0454882f $X=0.71 $Y=0.93 $X2=0
+ $Y2=0
cc_464 N_A_114_47#_M1049_g N_VPWR_c_1615_n 0.00379088f $X=1.355 $Y=2.465 $X2=0
+ $Y2=0
cc_465 N_A_114_47#_c_470_n N_VPWR_c_1615_n 0.0436221f $X=0.71 $Y=0.93 $X2=0
+ $Y2=0
cc_466 N_A_114_47#_M1054_g N_VPWR_c_1616_n 0.00368607f $X=1.785 $Y=2.465 $X2=0
+ $Y2=0
cc_467 N_A_114_47#_M1068_g N_VPWR_c_1616_n 0.00368607f $X=2.215 $Y=2.465 $X2=0
+ $Y2=0
cc_468 N_A_114_47#_M1071_g N_VPWR_c_1617_n 0.00334938f $X=2.645 $Y=2.465 $X2=0
+ $Y2=0
cc_469 N_A_114_47#_c_470_n N_VPWR_c_1637_n 0.0110337f $X=0.71 $Y=0.93 $X2=0
+ $Y2=0
cc_470 N_A_114_47#_M1049_g N_VPWR_c_1639_n 0.00549284f $X=1.355 $Y=2.465 $X2=0
+ $Y2=0
cc_471 N_A_114_47#_M1054_g N_VPWR_c_1639_n 0.00549284f $X=1.785 $Y=2.465 $X2=0
+ $Y2=0
cc_472 N_A_114_47#_M1068_g N_VPWR_c_1641_n 0.00549284f $X=2.215 $Y=2.465 $X2=0
+ $Y2=0
cc_473 N_A_114_47#_M1071_g N_VPWR_c_1641_n 0.00549284f $X=2.645 $Y=2.465 $X2=0
+ $Y2=0
cc_474 N_A_114_47#_M1004_s N_VPWR_c_1612_n 0.00606379f $X=0.57 $Y=1.835 $X2=0
+ $Y2=0
cc_475 N_A_114_47#_M1049_g N_VPWR_c_1612_n 0.00981859f $X=1.355 $Y=2.465 $X2=0
+ $Y2=0
cc_476 N_A_114_47#_M1054_g N_VPWR_c_1612_n 0.00979325f $X=1.785 $Y=2.465 $X2=0
+ $Y2=0
cc_477 N_A_114_47#_M1068_g N_VPWR_c_1612_n 0.00979325f $X=2.215 $Y=2.465 $X2=0
+ $Y2=0
cc_478 N_A_114_47#_M1071_g N_VPWR_c_1612_n 0.00981859f $X=2.645 $Y=2.465 $X2=0
+ $Y2=0
cc_479 N_A_114_47#_c_470_n N_VPWR_c_1612_n 0.00648955f $X=0.71 $Y=0.93 $X2=0
+ $Y2=0
cc_480 N_A_114_47#_c_486_n N_VGND_M1024_d 0.0142964f $X=2.19 $Y=0.71 $X2=0 $Y2=0
cc_481 N_A_114_47#_c_486_n N_VGND_M1043_d 0.00415361f $X=2.19 $Y=0.71 $X2=0
+ $Y2=0
cc_482 N_A_114_47#_c_508_p N_VGND_M1043_d 0.00691765f $X=2.275 $Y=1.005 $X2=0
+ $Y2=0
cc_483 N_A_114_47#_c_471_n N_VGND_M1043_d 0.00567015f $X=5.985 $Y=1.17 $X2=0
+ $Y2=0
cc_484 N_A_114_47#_M1010_g N_VGND_c_2481_n 0.00442169f $X=1.515 $Y=0.655 $X2=0
+ $Y2=0
cc_485 N_A_114_47#_c_486_n N_VGND_c_2481_n 0.0235397f $X=2.19 $Y=0.71 $X2=0
+ $Y2=0
cc_486 N_A_114_47#_M1043_g N_VGND_c_2482_n 0.0126505f $X=2.175 $Y=0.655 $X2=0
+ $Y2=0
cc_487 N_A_114_47#_c_438_n N_VGND_c_2482_n 0.00308556f $X=3.28 $Y=0.985 $X2=0
+ $Y2=0
cc_488 N_A_114_47#_c_486_n N_VGND_c_2482_n 0.00151842f $X=2.19 $Y=0.71 $X2=0
+ $Y2=0
cc_489 N_A_114_47#_c_471_n N_VGND_c_2482_n 0.0106449f $X=5.985 $Y=1.17 $X2=0
+ $Y2=0
cc_490 N_A_114_47#_c_438_n N_VGND_c_2483_n 0.00427332f $X=3.28 $Y=0.985 $X2=0
+ $Y2=0
cc_491 N_A_114_47#_c_441_n N_VGND_c_2483_n 0.00670177f $X=3.79 $Y=0.985 $X2=0
+ $Y2=0
cc_492 N_A_114_47#_c_442_n N_VGND_c_2483_n 5.78217e-19 $X=4.22 $Y=0.985 $X2=0
+ $Y2=0
cc_493 N_A_114_47#_c_441_n N_VGND_c_2484_n 5.78217e-19 $X=3.79 $Y=0.985 $X2=0
+ $Y2=0
cc_494 N_A_114_47#_c_442_n N_VGND_c_2484_n 0.00666812f $X=4.22 $Y=0.985 $X2=0
+ $Y2=0
cc_495 N_A_114_47#_c_443_n N_VGND_c_2484_n 0.00666812f $X=4.65 $Y=0.985 $X2=0
+ $Y2=0
cc_496 N_A_114_47#_c_444_n N_VGND_c_2484_n 5.78217e-19 $X=5.08 $Y=0.985 $X2=0
+ $Y2=0
cc_497 N_A_114_47#_c_443_n N_VGND_c_2485_n 5.78217e-19 $X=4.65 $Y=0.985 $X2=0
+ $Y2=0
cc_498 N_A_114_47#_c_444_n N_VGND_c_2485_n 0.00670177f $X=5.08 $Y=0.985 $X2=0
+ $Y2=0
cc_499 N_A_114_47#_c_447_n N_VGND_c_2485_n 0.00427332f $X=5.59 $Y=0.985 $X2=0
+ $Y2=0
cc_500 N_A_114_47#_c_448_n N_VGND_c_2486_n 0.00460722f $X=6.02 $Y=0.985 $X2=0
+ $Y2=0
cc_501 N_A_114_47#_c_450_n N_VGND_c_2486_n 0.00460722f $X=6.61 $Y=0.985 $X2=0
+ $Y2=0
cc_502 N_A_114_47#_c_452_n N_VGND_c_2487_n 0.00351184f $X=7.04 $Y=0.985 $X2=0
+ $Y2=0
cc_503 N_A_114_47#_c_453_n N_VGND_c_2487_n 0.00201283f $X=7.395 $Y=1.06 $X2=0
+ $Y2=0
cc_504 N_A_114_47#_c_454_n N_VGND_c_2487_n 0.00351184f $X=7.47 $Y=0.985 $X2=0
+ $Y2=0
cc_505 N_A_114_47#_c_456_n N_VGND_c_2488_n 0.00351184f $X=7.9 $Y=0.985 $X2=0
+ $Y2=0
cc_506 N_A_114_47#_c_457_n N_VGND_c_2488_n 0.00201283f $X=8.255 $Y=1.06 $X2=0
+ $Y2=0
cc_507 N_A_114_47#_c_458_n N_VGND_c_2488_n 0.00351184f $X=8.33 $Y=0.985 $X2=0
+ $Y2=0
cc_508 N_A_114_47#_c_460_n N_VGND_c_2489_n 0.00351184f $X=8.76 $Y=0.985 $X2=0
+ $Y2=0
cc_509 N_A_114_47#_c_461_n N_VGND_c_2489_n 0.00201283f $X=9.115 $Y=1.06 $X2=0
+ $Y2=0
cc_510 N_A_114_47#_c_462_n N_VGND_c_2489_n 0.00351184f $X=9.19 $Y=0.985 $X2=0
+ $Y2=0
cc_511 N_A_114_47#_M1010_g N_VGND_c_2493_n 0.0042361f $X=1.515 $Y=0.655 $X2=0
+ $Y2=0
cc_512 N_A_114_47#_M1043_g N_VGND_c_2493_n 0.00423551f $X=2.175 $Y=0.655 $X2=0
+ $Y2=0
cc_513 N_A_114_47#_c_486_n N_VGND_c_2493_n 0.0150846f $X=2.19 $Y=0.71 $X2=0
+ $Y2=0
cc_514 N_A_114_47#_c_441_n N_VGND_c_2495_n 0.00355956f $X=3.79 $Y=0.985 $X2=0
+ $Y2=0
cc_515 N_A_114_47#_c_442_n N_VGND_c_2495_n 0.00355956f $X=4.22 $Y=0.985 $X2=0
+ $Y2=0
cc_516 N_A_114_47#_c_443_n N_VGND_c_2497_n 0.00355956f $X=4.65 $Y=0.985 $X2=0
+ $Y2=0
cc_517 N_A_114_47#_c_444_n N_VGND_c_2497_n 0.00355956f $X=5.08 $Y=0.985 $X2=0
+ $Y2=0
cc_518 N_A_114_47#_c_447_n N_VGND_c_2499_n 0.00418148f $X=5.59 $Y=0.985 $X2=0
+ $Y2=0
cc_519 N_A_114_47#_c_448_n N_VGND_c_2499_n 0.00418148f $X=6.02 $Y=0.985 $X2=0
+ $Y2=0
cc_520 N_A_114_47#_c_450_n N_VGND_c_2501_n 0.00418148f $X=6.61 $Y=0.985 $X2=0
+ $Y2=0
cc_521 N_A_114_47#_c_452_n N_VGND_c_2501_n 0.00549284f $X=7.04 $Y=0.985 $X2=0
+ $Y2=0
cc_522 N_A_114_47#_c_454_n N_VGND_c_2503_n 0.00549284f $X=7.47 $Y=0.985 $X2=0
+ $Y2=0
cc_523 N_A_114_47#_c_456_n N_VGND_c_2503_n 0.00549284f $X=7.9 $Y=0.985 $X2=0
+ $Y2=0
cc_524 N_A_114_47#_c_458_n N_VGND_c_2505_n 0.00549284f $X=8.33 $Y=0.985 $X2=0
+ $Y2=0
cc_525 N_A_114_47#_c_460_n N_VGND_c_2505_n 0.00549284f $X=8.76 $Y=0.985 $X2=0
+ $Y2=0
cc_526 N_A_114_47#_c_462_n N_VGND_c_2507_n 0.0054778f $X=9.19 $Y=0.985 $X2=0
+ $Y2=0
cc_527 N_A_114_47#_c_596_p N_VGND_c_2511_n 0.0110337f $X=0.71 $Y=0.43 $X2=0
+ $Y2=0
cc_528 N_A_114_47#_c_486_n N_VGND_c_2511_n 0.00360256f $X=2.19 $Y=0.71 $X2=0
+ $Y2=0
cc_529 N_A_114_47#_c_438_n N_VGND_c_2512_n 0.00418148f $X=3.28 $Y=0.985 $X2=0
+ $Y2=0
cc_530 N_A_114_47#_M1020_s N_VGND_c_2515_n 0.0043284f $X=0.57 $Y=0.235 $X2=0
+ $Y2=0
cc_531 N_A_114_47#_M1010_g N_VGND_c_2515_n 0.00679384f $X=1.515 $Y=0.655 $X2=0
+ $Y2=0
cc_532 N_A_114_47#_M1043_g N_VGND_c_2515_n 0.00789778f $X=2.175 $Y=0.655 $X2=0
+ $Y2=0
cc_533 N_A_114_47#_c_438_n N_VGND_c_2515_n 0.00744378f $X=3.28 $Y=0.985 $X2=0
+ $Y2=0
cc_534 N_A_114_47#_c_441_n N_VGND_c_2515_n 0.00423262f $X=3.79 $Y=0.985 $X2=0
+ $Y2=0
cc_535 N_A_114_47#_c_442_n N_VGND_c_2515_n 0.00423262f $X=4.22 $Y=0.985 $X2=0
+ $Y2=0
cc_536 N_A_114_47#_c_443_n N_VGND_c_2515_n 0.00423262f $X=4.65 $Y=0.985 $X2=0
+ $Y2=0
cc_537 N_A_114_47#_c_444_n N_VGND_c_2515_n 0.00423262f $X=5.08 $Y=0.985 $X2=0
+ $Y2=0
cc_538 N_A_114_47#_c_447_n N_VGND_c_2515_n 0.00604412f $X=5.59 $Y=0.985 $X2=0
+ $Y2=0
cc_539 N_A_114_47#_c_448_n N_VGND_c_2515_n 0.00622304f $X=6.02 $Y=0.985 $X2=0
+ $Y2=0
cc_540 N_A_114_47#_c_450_n N_VGND_c_2515_n 0.00622304f $X=6.61 $Y=0.985 $X2=0
+ $Y2=0
cc_541 N_A_114_47#_c_452_n N_VGND_c_2515_n 0.00997134f $X=7.04 $Y=0.985 $X2=0
+ $Y2=0
cc_542 N_A_114_47#_c_454_n N_VGND_c_2515_n 0.00997134f $X=7.47 $Y=0.985 $X2=0
+ $Y2=0
cc_543 N_A_114_47#_c_456_n N_VGND_c_2515_n 0.00997134f $X=7.9 $Y=0.985 $X2=0
+ $Y2=0
cc_544 N_A_114_47#_c_458_n N_VGND_c_2515_n 0.00997134f $X=8.33 $Y=0.985 $X2=0
+ $Y2=0
cc_545 N_A_114_47#_c_460_n N_VGND_c_2515_n 0.00997134f $X=8.76 $Y=0.985 $X2=0
+ $Y2=0
cc_546 N_A_114_47#_c_462_n N_VGND_c_2515_n 0.00996158f $X=9.19 $Y=0.985 $X2=0
+ $Y2=0
cc_547 N_A_114_47#_c_596_p N_VGND_c_2515_n 0.00648955f $X=0.71 $Y=0.43 $X2=0
+ $Y2=0
cc_548 N_A_114_47#_c_486_n N_VGND_c_2515_n 0.0346221f $X=2.19 $Y=0.71 $X2=0
+ $Y2=0
cc_549 N_A_114_47#_M1043_g N_A_584_47#_c_2722_n 0.00447047f $X=2.175 $Y=0.655
+ $X2=0 $Y2=0
cc_550 N_A_114_47#_c_438_n N_A_584_47#_c_2722_n 0.0076206f $X=3.28 $Y=0.985
+ $X2=0 $Y2=0
cc_551 N_A_114_47#_c_441_n N_A_584_47#_c_2722_n 5.96129e-19 $X=3.79 $Y=0.985
+ $X2=0 $Y2=0
cc_552 N_A_114_47#_c_486_n N_A_584_47#_c_2722_n 0.00111126f $X=2.19 $Y=0.71
+ $X2=0 $Y2=0
cc_553 N_A_114_47#_c_438_n N_A_584_47#_c_2735_n 0.00906605f $X=3.28 $Y=0.985
+ $X2=0 $Y2=0
cc_554 N_A_114_47#_c_439_n N_A_584_47#_c_2735_n 0.00415476f $X=3.715 $Y=1.16
+ $X2=0 $Y2=0
cc_555 N_A_114_47#_c_441_n N_A_584_47#_c_2735_n 0.011173f $X=3.79 $Y=0.985 $X2=0
+ $Y2=0
cc_556 N_A_114_47#_c_471_n N_A_584_47#_c_2735_n 0.0420906f $X=5.985 $Y=1.17
+ $X2=0 $Y2=0
cc_557 N_A_114_47#_M1043_g N_A_584_47#_c_2723_n 9.47371e-19 $X=2.175 $Y=0.655
+ $X2=0 $Y2=0
cc_558 N_A_114_47#_c_438_n N_A_584_47#_c_2723_n 0.00246487f $X=3.28 $Y=0.985
+ $X2=0 $Y2=0
cc_559 N_A_114_47#_c_440_n N_A_584_47#_c_2723_n 0.00709509f $X=3.355 $Y=1.16
+ $X2=0 $Y2=0
cc_560 N_A_114_47#_c_486_n N_A_584_47#_c_2723_n 0.00558438f $X=2.19 $Y=0.71
+ $X2=0 $Y2=0
cc_561 N_A_114_47#_c_508_p N_A_584_47#_c_2723_n 0.00107308f $X=2.275 $Y=1.005
+ $X2=0 $Y2=0
cc_562 N_A_114_47#_c_471_n N_A_584_47#_c_2723_n 0.0232551f $X=5.985 $Y=1.17
+ $X2=0 $Y2=0
cc_563 N_A_114_47#_c_442_n N_A_584_47#_c_2745_n 0.0107293f $X=4.22 $Y=0.985
+ $X2=0 $Y2=0
cc_564 N_A_114_47#_c_443_n N_A_584_47#_c_2745_n 0.0107293f $X=4.65 $Y=0.985
+ $X2=0 $Y2=0
cc_565 N_A_114_47#_c_446_n N_A_584_47#_c_2745_n 0.0023082f $X=5.155 $Y=1.16
+ $X2=0 $Y2=0
cc_566 N_A_114_47#_c_471_n N_A_584_47#_c_2745_n 0.0402196f $X=5.985 $Y=1.17
+ $X2=0 $Y2=0
cc_567 N_A_114_47#_c_444_n N_A_584_47#_c_2749_n 0.011173f $X=5.08 $Y=0.985 $X2=0
+ $Y2=0
cc_568 N_A_114_47#_c_445_n N_A_584_47#_c_2749_n 0.00415476f $X=5.515 $Y=1.16
+ $X2=0 $Y2=0
cc_569 N_A_114_47#_c_447_n N_A_584_47#_c_2749_n 0.00906605f $X=5.59 $Y=0.985
+ $X2=0 $Y2=0
cc_570 N_A_114_47#_c_471_n N_A_584_47#_c_2749_n 0.0420906f $X=5.985 $Y=1.17
+ $X2=0 $Y2=0
cc_571 N_A_114_47#_c_444_n N_A_584_47#_c_2753_n 5.96129e-19 $X=5.08 $Y=0.985
+ $X2=0 $Y2=0
cc_572 N_A_114_47#_c_447_n N_A_584_47#_c_2753_n 0.00691985f $X=5.59 $Y=0.985
+ $X2=0 $Y2=0
cc_573 N_A_114_47#_c_448_n N_A_584_47#_c_2753_n 0.00715928f $X=6.02 $Y=0.985
+ $X2=0 $Y2=0
cc_574 N_A_114_47#_c_450_n N_A_584_47#_c_2753_n 8.52731e-19 $X=6.61 $Y=0.985
+ $X2=0 $Y2=0
cc_575 N_A_114_47#_c_448_n N_A_584_47#_c_2757_n 0.00942392f $X=6.02 $Y=0.985
+ $X2=0 $Y2=0
cc_576 N_A_114_47#_c_449_n N_A_584_47#_c_2757_n 0.00836146f $X=6.535 $Y=1.06
+ $X2=0 $Y2=0
cc_577 N_A_114_47#_c_450_n N_A_584_47#_c_2757_n 0.0100267f $X=6.61 $Y=0.985
+ $X2=0 $Y2=0
cc_578 N_A_114_47#_c_471_n N_A_584_47#_c_2757_n 0.0104655f $X=5.985 $Y=1.17
+ $X2=0 $Y2=0
cc_579 N_A_114_47#_c_448_n N_A_584_47#_c_2761_n 8.52731e-19 $X=6.02 $Y=0.985
+ $X2=0 $Y2=0
cc_580 N_A_114_47#_c_450_n N_A_584_47#_c_2761_n 0.00758062f $X=6.61 $Y=0.985
+ $X2=0 $Y2=0
cc_581 N_A_114_47#_c_452_n N_A_584_47#_c_2761_n 0.00568122f $X=7.04 $Y=0.985
+ $X2=0 $Y2=0
cc_582 N_A_114_47#_c_448_n N_A_584_47#_c_2764_n 7.15856e-19 $X=6.02 $Y=0.985
+ $X2=0 $Y2=0
cc_583 N_A_114_47#_c_450_n N_A_584_47#_c_2764_n 0.00516629f $X=6.61 $Y=0.985
+ $X2=0 $Y2=0
cc_584 N_A_114_47#_c_451_n N_A_584_47#_c_2764_n 0.00264461f $X=6.965 $Y=1.06
+ $X2=0 $Y2=0
cc_585 N_A_114_47#_c_452_n N_A_584_47#_c_2764_n 0.00465882f $X=7.04 $Y=0.985
+ $X2=0 $Y2=0
cc_586 N_A_114_47#_c_454_n N_A_584_47#_c_2764_n 4.67286e-19 $X=7.47 $Y=0.985
+ $X2=0 $Y2=0
cc_587 N_A_114_47#_c_464_n N_A_584_47#_c_2764_n 4.29786e-19 $X=6.61 $Y=1.06
+ $X2=0 $Y2=0
cc_588 N_A_114_47#_c_465_n N_A_584_47#_c_2764_n 2.2335e-19 $X=7.04 $Y=1.06 $X2=0
+ $Y2=0
cc_589 N_A_114_47#_c_453_n N_A_584_47#_c_2724_n 0.0105811f $X=7.395 $Y=1.06
+ $X2=0 $Y2=0
cc_590 N_A_114_47#_c_465_n N_A_584_47#_c_2724_n 0.00736947f $X=7.04 $Y=1.06
+ $X2=0 $Y2=0
cc_591 N_A_114_47#_c_466_n N_A_584_47#_c_2724_n 0.00736947f $X=7.47 $Y=1.06
+ $X2=0 $Y2=0
cc_592 N_A_114_47#_c_451_n N_A_584_47#_c_2725_n 0.00426194f $X=6.965 $Y=1.06
+ $X2=0 $Y2=0
cc_593 N_A_114_47#_c_464_n N_A_584_47#_c_2725_n 0.00438771f $X=6.61 $Y=1.06
+ $X2=0 $Y2=0
cc_594 N_A_114_47#_c_465_n N_A_584_47#_c_2725_n 3.83268e-19 $X=7.04 $Y=1.06
+ $X2=0 $Y2=0
cc_595 N_A_114_47#_c_471_n N_A_584_47#_c_2725_n 0.00559377f $X=5.985 $Y=1.17
+ $X2=0 $Y2=0
cc_596 N_A_114_47#_c_452_n N_A_584_47#_c_2778_n 6.61624e-19 $X=7.04 $Y=0.985
+ $X2=0 $Y2=0
cc_597 N_A_114_47#_c_454_n N_A_584_47#_c_2778_n 0.0128096f $X=7.47 $Y=0.985
+ $X2=0 $Y2=0
cc_598 N_A_114_47#_c_455_n N_A_584_47#_c_2778_n 0.00264461f $X=7.825 $Y=1.06
+ $X2=0 $Y2=0
cc_599 N_A_114_47#_c_456_n N_A_584_47#_c_2778_n 0.0128098f $X=7.9 $Y=0.985 $X2=0
+ $Y2=0
cc_600 N_A_114_47#_c_458_n N_A_584_47#_c_2778_n 6.61637e-19 $X=8.33 $Y=0.985
+ $X2=0 $Y2=0
cc_601 N_A_114_47#_c_466_n N_A_584_47#_c_2778_n 2.2335e-19 $X=7.47 $Y=1.06 $X2=0
+ $Y2=0
cc_602 N_A_114_47#_c_467_n N_A_584_47#_c_2778_n 2.2335e-19 $X=7.9 $Y=1.06 $X2=0
+ $Y2=0
cc_603 N_A_114_47#_c_457_n N_A_584_47#_c_2726_n 0.0105811f $X=8.255 $Y=1.06
+ $X2=0 $Y2=0
cc_604 N_A_114_47#_c_467_n N_A_584_47#_c_2726_n 0.00736947f $X=7.9 $Y=1.06 $X2=0
+ $Y2=0
cc_605 N_A_114_47#_c_468_n N_A_584_47#_c_2726_n 0.00736947f $X=8.33 $Y=1.06
+ $X2=0 $Y2=0
cc_606 N_A_114_47#_c_456_n N_A_584_47#_c_2788_n 6.61637e-19 $X=7.9 $Y=0.985
+ $X2=0 $Y2=0
cc_607 N_A_114_47#_c_458_n N_A_584_47#_c_2788_n 0.0128098f $X=8.33 $Y=0.985
+ $X2=0 $Y2=0
cc_608 N_A_114_47#_c_459_n N_A_584_47#_c_2788_n 0.00264461f $X=8.685 $Y=1.06
+ $X2=0 $Y2=0
cc_609 N_A_114_47#_c_460_n N_A_584_47#_c_2788_n 0.0128098f $X=8.76 $Y=0.985
+ $X2=0 $Y2=0
cc_610 N_A_114_47#_c_462_n N_A_584_47#_c_2788_n 6.61637e-19 $X=9.19 $Y=0.985
+ $X2=0 $Y2=0
cc_611 N_A_114_47#_c_468_n N_A_584_47#_c_2788_n 2.2335e-19 $X=8.33 $Y=1.06 $X2=0
+ $Y2=0
cc_612 N_A_114_47#_c_469_n N_A_584_47#_c_2788_n 2.2335e-19 $X=8.76 $Y=1.06 $X2=0
+ $Y2=0
cc_613 N_A_114_47#_c_461_n N_A_584_47#_c_2727_n 0.020008f $X=9.115 $Y=1.06 $X2=0
+ $Y2=0
cc_614 N_A_114_47#_c_469_n N_A_584_47#_c_2727_n 0.00736947f $X=8.76 $Y=1.06
+ $X2=0 $Y2=0
cc_615 N_A_114_47#_c_460_n N_A_584_47#_c_2797_n 5.98671e-19 $X=8.76 $Y=0.985
+ $X2=0 $Y2=0
cc_616 N_A_114_47#_c_461_n N_A_584_47#_c_2797_n 3.30973e-19 $X=9.115 $Y=1.06
+ $X2=0 $Y2=0
cc_617 N_A_114_47#_c_462_n N_A_584_47#_c_2797_n 0.00891018f $X=9.19 $Y=0.985
+ $X2=0 $Y2=0
cc_618 N_A_114_47#_c_462_n N_A_584_47#_c_2800_n 0.00381664f $X=9.19 $Y=0.985
+ $X2=0 $Y2=0
cc_619 N_A_114_47#_c_446_n N_A_584_47#_c_2801_n 0.00238404f $X=5.155 $Y=1.16
+ $X2=0 $Y2=0
cc_620 N_A_114_47#_c_471_n N_A_584_47#_c_2801_n 0.013056f $X=5.985 $Y=1.17 $X2=0
+ $Y2=0
cc_621 N_A_114_47#_c_446_n N_A_584_47#_c_2803_n 0.00238404f $X=5.155 $Y=1.16
+ $X2=0 $Y2=0
cc_622 N_A_114_47#_c_471_n N_A_584_47#_c_2803_n 0.013056f $X=5.985 $Y=1.17 $X2=0
+ $Y2=0
cc_623 N_A_114_47#_c_447_n N_A_584_47#_c_2805_n 0.00176282f $X=5.59 $Y=0.985
+ $X2=0 $Y2=0
cc_624 N_A_114_47#_c_448_n N_A_584_47#_c_2805_n 0.00176282f $X=6.02 $Y=0.985
+ $X2=0 $Y2=0
cc_625 N_A_114_47#_c_471_n N_A_584_47#_c_2805_n 0.0207713f $X=5.985 $Y=1.17
+ $X2=0 $Y2=0
cc_626 N_A_114_47#_c_472_n N_A_584_47#_c_2805_n 0.00238404f $X=6.15 $Y=1.16
+ $X2=0 $Y2=0
cc_627 N_A_114_47#_c_450_n N_A_584_47#_c_2809_n 9.861e-19 $X=6.61 $Y=0.985 $X2=0
+ $Y2=0
cc_628 N_A_114_47#_c_452_n N_A_584_47#_c_2809_n 0.0024377f $X=7.04 $Y=0.985
+ $X2=0 $Y2=0
cc_629 N_A_114_47#_c_455_n N_A_584_47#_c_2728_n 0.00426194f $X=7.825 $Y=1.06
+ $X2=0 $Y2=0
cc_630 N_A_114_47#_c_466_n N_A_584_47#_c_2728_n 3.83268e-19 $X=7.47 $Y=1.06
+ $X2=0 $Y2=0
cc_631 N_A_114_47#_c_467_n N_A_584_47#_c_2728_n 3.83268e-19 $X=7.9 $Y=1.06 $X2=0
+ $Y2=0
cc_632 N_A_114_47#_c_459_n N_A_584_47#_c_2729_n 0.00426194f $X=8.685 $Y=1.06
+ $X2=0 $Y2=0
cc_633 N_A_114_47#_c_468_n N_A_584_47#_c_2729_n 3.83268e-19 $X=8.33 $Y=1.06
+ $X2=0 $Y2=0
cc_634 N_A_114_47#_c_469_n N_A_584_47#_c_2729_n 3.83268e-19 $X=8.76 $Y=1.06
+ $X2=0 $Y2=0
cc_635 N_A_286_367#_c_714_n N_A_1909_21#_c_1034_n 0.00700401f $X=10.05 $Y=1.65
+ $X2=0 $Y2=0
cc_636 N_A_286_367#_c_714_n N_A_1909_21#_c_1035_n 0.0172189f $X=10.05 $Y=1.65
+ $X2=0 $Y2=0
cc_637 N_A_286_367#_c_728_n N_A_1909_21#_c_1035_n 0.0015487f $X=9.615 $Y=1.51
+ $X2=0 $Y2=0
cc_638 N_A_286_367#_c_724_n N_A_1909_21#_c_1037_n 0.00700401f $X=10.405 $Y=1.65
+ $X2=0 $Y2=0
cc_639 N_A_286_367#_c_725_n N_A_1909_21#_c_1039_n 0.00700401f $X=10.835 $Y=1.65
+ $X2=0 $Y2=0
cc_640 N_A_286_367#_c_713_n N_A_1909_21#_c_1073_n 0.00700401f $X=10.33 $Y=1.65
+ $X2=0 $Y2=0
cc_641 N_A_286_367#_c_715_n N_A_1909_21#_c_1074_n 0.00700401f $X=10.76 $Y=1.65
+ $X2=0 $Y2=0
cc_642 N_A_286_367#_c_716_n N_A_1909_21#_c_1075_n 0.00700401f $X=11.19 $Y=1.65
+ $X2=0 $Y2=0
cc_643 N_A_286_367#_c_774_n N_VPWR_M1054_s 7.83958e-19 $X=2.265 $Y=1.9 $X2=0
+ $Y2=0
cc_644 N_A_286_367#_c_775_n N_VPWR_M1054_s 0.00101261f $X=2.01 $Y=1.9 $X2=0
+ $Y2=0
cc_645 N_A_286_367#_c_775_n N_VPWR_c_1615_n 0.00745032f $X=2.01 $Y=1.9 $X2=0
+ $Y2=0
cc_646 N_A_286_367#_c_775_n N_VPWR_c_1616_n 0.0129053f $X=2.01 $Y=1.9 $X2=0
+ $Y2=0
cc_647 N_A_286_367#_c_731_n N_VPWR_c_1617_n 0.00334938f $X=3.075 $Y=1.725 $X2=0
+ $Y2=0
cc_648 N_A_286_367#_c_730_n N_VPWR_c_1617_n 0.0138021f $X=6.39 $Y=1.515 $X2=0
+ $Y2=0
cc_649 N_A_286_367#_c_734_n N_VPWR_c_1618_n 0.00370529f $X=3.505 $Y=1.725 $X2=0
+ $Y2=0
cc_650 N_A_286_367#_c_736_n N_VPWR_c_1618_n 0.00243509f $X=3.935 $Y=1.725 $X2=0
+ $Y2=0
cc_651 N_A_286_367#_c_736_n N_VPWR_c_1619_n 0.00558004f $X=3.935 $Y=1.725 $X2=0
+ $Y2=0
cc_652 N_A_286_367#_c_738_n N_VPWR_c_1619_n 0.00558004f $X=4.365 $Y=1.725 $X2=0
+ $Y2=0
cc_653 N_A_286_367#_c_738_n N_VPWR_c_1620_n 0.00243509f $X=4.365 $Y=1.725 $X2=0
+ $Y2=0
cc_654 N_A_286_367#_c_740_n N_VPWR_c_1620_n 0.00243509f $X=4.795 $Y=1.725 $X2=0
+ $Y2=0
cc_655 N_A_286_367#_c_742_n N_VPWR_c_1621_n 0.00243509f $X=5.225 $Y=1.725 $X2=0
+ $Y2=0
cc_656 N_A_286_367#_c_744_n N_VPWR_c_1621_n 0.00243509f $X=5.655 $Y=1.725 $X2=0
+ $Y2=0
cc_657 N_A_286_367#_c_746_n N_VPWR_c_1622_n 0.00243509f $X=6.085 $Y=1.725 $X2=0
+ $Y2=0
cc_658 N_A_286_367#_c_748_n N_VPWR_c_1622_n 0.00243509f $X=6.515 $Y=1.725 $X2=0
+ $Y2=0
cc_659 N_A_286_367#_c_749_n N_VPWR_c_1623_n 0.00243509f $X=6.945 $Y=1.725 $X2=0
+ $Y2=0
cc_660 N_A_286_367#_c_750_n N_VPWR_c_1623_n 0.00243509f $X=7.375 $Y=1.725 $X2=0
+ $Y2=0
cc_661 N_A_286_367#_c_751_n N_VPWR_c_1624_n 0.00252142f $X=7.805 $Y=1.725 $X2=0
+ $Y2=0
cc_662 N_A_286_367#_c_752_n N_VPWR_c_1624_n 0.0118499f $X=8.255 $Y=1.725 $X2=0
+ $Y2=0
cc_663 N_A_286_367#_c_752_n N_VPWR_c_1625_n 0.00558004f $X=8.255 $Y=1.725 $X2=0
+ $Y2=0
cc_664 N_A_286_367#_c_753_n N_VPWR_c_1625_n 0.00558004f $X=8.685 $Y=1.725 $X2=0
+ $Y2=0
cc_665 N_A_286_367#_c_753_n N_VPWR_c_1626_n 0.00370529f $X=8.685 $Y=1.725 $X2=0
+ $Y2=0
cc_666 N_A_286_367#_c_754_n N_VPWR_c_1626_n 0.00243509f $X=9.115 $Y=1.725 $X2=0
+ $Y2=0
cc_667 N_A_286_367#_c_755_n N_VPWR_c_1627_n 0.00243509f $X=9.545 $Y=1.725 $X2=0
+ $Y2=0
cc_668 N_A_286_367#_c_756_n N_VPWR_c_1627_n 0.00370529f $X=9.975 $Y=1.725 $X2=0
+ $Y2=0
cc_669 N_A_286_367#_c_759_n N_VPWR_c_1628_n 0.00365752f $X=10.405 $Y=1.725 $X2=0
+ $Y2=0
cc_670 N_A_286_367#_c_715_n N_VPWR_c_1628_n 0.00222336f $X=10.76 $Y=1.65 $X2=0
+ $Y2=0
cc_671 N_A_286_367#_c_761_n N_VPWR_c_1628_n 0.0023508f $X=10.835 $Y=1.725 $X2=0
+ $Y2=0
cc_672 N_A_286_367#_c_761_n N_VPWR_c_1629_n 7.31436e-19 $X=10.835 $Y=1.725 $X2=0
+ $Y2=0
cc_673 N_A_286_367#_c_763_n N_VPWR_c_1629_n 0.0135992f $X=11.265 $Y=1.725 $X2=0
+ $Y2=0
cc_674 N_A_286_367#_c_777_n N_VPWR_c_1639_n 0.0177952f $X=1.57 $Y=2.9 $X2=0
+ $Y2=0
cc_675 N_A_286_367#_c_808_n N_VPWR_c_1641_n 0.0177952f $X=2.43 $Y=2.9 $X2=0
+ $Y2=0
cc_676 N_A_286_367#_c_731_n N_VPWR_c_1643_n 0.00558004f $X=3.075 $Y=1.725 $X2=0
+ $Y2=0
cc_677 N_A_286_367#_c_734_n N_VPWR_c_1643_n 0.00558004f $X=3.505 $Y=1.725 $X2=0
+ $Y2=0
cc_678 N_A_286_367#_c_740_n N_VPWR_c_1645_n 0.00558004f $X=4.795 $Y=1.725 $X2=0
+ $Y2=0
cc_679 N_A_286_367#_c_742_n N_VPWR_c_1645_n 0.00558004f $X=5.225 $Y=1.725 $X2=0
+ $Y2=0
cc_680 N_A_286_367#_c_744_n N_VPWR_c_1647_n 0.00558004f $X=5.655 $Y=1.725 $X2=0
+ $Y2=0
cc_681 N_A_286_367#_c_746_n N_VPWR_c_1647_n 0.00558004f $X=6.085 $Y=1.725 $X2=0
+ $Y2=0
cc_682 N_A_286_367#_c_748_n N_VPWR_c_1649_n 0.00558004f $X=6.515 $Y=1.725 $X2=0
+ $Y2=0
cc_683 N_A_286_367#_c_749_n N_VPWR_c_1649_n 0.00558004f $X=6.945 $Y=1.725 $X2=0
+ $Y2=0
cc_684 N_A_286_367#_c_750_n N_VPWR_c_1651_n 0.00558004f $X=7.375 $Y=1.725 $X2=0
+ $Y2=0
cc_685 N_A_286_367#_c_751_n N_VPWR_c_1651_n 0.00558004f $X=7.805 $Y=1.725 $X2=0
+ $Y2=0
cc_686 N_A_286_367#_c_754_n N_VPWR_c_1653_n 0.00558004f $X=9.115 $Y=1.725 $X2=0
+ $Y2=0
cc_687 N_A_286_367#_c_755_n N_VPWR_c_1653_n 0.00558004f $X=9.545 $Y=1.725 $X2=0
+ $Y2=0
cc_688 N_A_286_367#_c_756_n N_VPWR_c_1655_n 0.00549284f $X=9.975 $Y=1.725 $X2=0
+ $Y2=0
cc_689 N_A_286_367#_c_759_n N_VPWR_c_1655_n 0.00549284f $X=10.405 $Y=1.725 $X2=0
+ $Y2=0
cc_690 N_A_286_367#_c_761_n N_VPWR_c_1657_n 0.00549284f $X=10.835 $Y=1.725 $X2=0
+ $Y2=0
cc_691 N_A_286_367#_c_763_n N_VPWR_c_1657_n 0.00486043f $X=11.265 $Y=1.725 $X2=0
+ $Y2=0
cc_692 N_A_286_367#_M1049_d N_VPWR_c_1612_n 0.00223819f $X=1.43 $Y=1.835 $X2=0
+ $Y2=0
cc_693 N_A_286_367#_M1068_d N_VPWR_c_1612_n 0.00223819f $X=2.29 $Y=1.835 $X2=0
+ $Y2=0
cc_694 N_A_286_367#_c_731_n N_VPWR_c_1612_n 0.00995889f $X=3.075 $Y=1.725 $X2=0
+ $Y2=0
cc_695 N_A_286_367#_c_734_n N_VPWR_c_1612_n 0.00990622f $X=3.505 $Y=1.725 $X2=0
+ $Y2=0
cc_696 N_A_286_367#_c_736_n N_VPWR_c_1612_n 0.00990622f $X=3.935 $Y=1.725 $X2=0
+ $Y2=0
cc_697 N_A_286_367#_c_738_n N_VPWR_c_1612_n 0.00990622f $X=4.365 $Y=1.725 $X2=0
+ $Y2=0
cc_698 N_A_286_367#_c_740_n N_VPWR_c_1612_n 0.00990622f $X=4.795 $Y=1.725 $X2=0
+ $Y2=0
cc_699 N_A_286_367#_c_742_n N_VPWR_c_1612_n 0.00990622f $X=5.225 $Y=1.725 $X2=0
+ $Y2=0
cc_700 N_A_286_367#_c_744_n N_VPWR_c_1612_n 0.00990622f $X=5.655 $Y=1.725 $X2=0
+ $Y2=0
cc_701 N_A_286_367#_c_746_n N_VPWR_c_1612_n 0.00990622f $X=6.085 $Y=1.725 $X2=0
+ $Y2=0
cc_702 N_A_286_367#_c_748_n N_VPWR_c_1612_n 0.00990622f $X=6.515 $Y=1.725 $X2=0
+ $Y2=0
cc_703 N_A_286_367#_c_749_n N_VPWR_c_1612_n 0.00990622f $X=6.945 $Y=1.725 $X2=0
+ $Y2=0
cc_704 N_A_286_367#_c_750_n N_VPWR_c_1612_n 0.00990622f $X=7.375 $Y=1.725 $X2=0
+ $Y2=0
cc_705 N_A_286_367#_c_751_n N_VPWR_c_1612_n 0.00995748f $X=7.805 $Y=1.725 $X2=0
+ $Y2=0
cc_706 N_A_286_367#_c_752_n N_VPWR_c_1612_n 0.0100121f $X=8.255 $Y=1.725 $X2=0
+ $Y2=0
cc_707 N_A_286_367#_c_753_n N_VPWR_c_1612_n 0.00990622f $X=8.685 $Y=1.725 $X2=0
+ $Y2=0
cc_708 N_A_286_367#_c_754_n N_VPWR_c_1612_n 0.00990622f $X=9.115 $Y=1.725 $X2=0
+ $Y2=0
cc_709 N_A_286_367#_c_755_n N_VPWR_c_1612_n 0.00990622f $X=9.545 $Y=1.725 $X2=0
+ $Y2=0
cc_710 N_A_286_367#_c_756_n N_VPWR_c_1612_n 0.00976592f $X=9.975 $Y=1.725 $X2=0
+ $Y2=0
cc_711 N_A_286_367#_c_759_n N_VPWR_c_1612_n 0.00979325f $X=10.405 $Y=1.725 $X2=0
+ $Y2=0
cc_712 N_A_286_367#_c_761_n N_VPWR_c_1612_n 0.00979325f $X=10.835 $Y=1.725 $X2=0
+ $Y2=0
cc_713 N_A_286_367#_c_763_n N_VPWR_c_1612_n 0.00824727f $X=11.265 $Y=1.725 $X2=0
+ $Y2=0
cc_714 N_A_286_367#_c_777_n N_VPWR_c_1612_n 0.0123247f $X=1.57 $Y=2.9 $X2=0
+ $Y2=0
cc_715 N_A_286_367#_c_808_n N_VPWR_c_1612_n 0.0123247f $X=2.43 $Y=2.9 $X2=0
+ $Y2=0
cc_716 N_A_286_367#_c_734_n N_A_630_367#_c_1959_n 0.0111252f $X=3.505 $Y=1.725
+ $X2=0 $Y2=0
cc_717 N_A_286_367#_c_706_n N_A_630_367#_c_1959_n 0.00199111f $X=3.86 $Y=1.65
+ $X2=0 $Y2=0
cc_718 N_A_286_367#_c_736_n N_A_630_367#_c_1959_n 0.0111252f $X=3.935 $Y=1.725
+ $X2=0 $Y2=0
cc_719 N_A_286_367#_c_730_n N_A_630_367#_c_1959_n 0.0308981f $X=6.39 $Y=1.515
+ $X2=0 $Y2=0
cc_720 N_A_286_367#_c_738_n N_A_630_367#_c_1963_n 0.0111252f $X=4.365 $Y=1.725
+ $X2=0 $Y2=0
cc_721 N_A_286_367#_c_708_n N_A_630_367#_c_1963_n 0.00199111f $X=4.72 $Y=1.65
+ $X2=0 $Y2=0
cc_722 N_A_286_367#_c_740_n N_A_630_367#_c_1963_n 0.0111252f $X=4.795 $Y=1.725
+ $X2=0 $Y2=0
cc_723 N_A_286_367#_c_730_n N_A_630_367#_c_1963_n 0.0308981f $X=6.39 $Y=1.515
+ $X2=0 $Y2=0
cc_724 N_A_286_367#_c_742_n N_A_630_367#_c_1967_n 0.0111252f $X=5.225 $Y=1.725
+ $X2=0 $Y2=0
cc_725 N_A_286_367#_c_710_n N_A_630_367#_c_1967_n 0.00199111f $X=5.58 $Y=1.65
+ $X2=0 $Y2=0
cc_726 N_A_286_367#_c_744_n N_A_630_367#_c_1967_n 0.0111252f $X=5.655 $Y=1.725
+ $X2=0 $Y2=0
cc_727 N_A_286_367#_c_730_n N_A_630_367#_c_1967_n 0.0308981f $X=6.39 $Y=1.515
+ $X2=0 $Y2=0
cc_728 N_A_286_367#_c_746_n N_A_630_367#_c_1971_n 0.0111313f $X=6.085 $Y=1.725
+ $X2=0 $Y2=0
cc_729 N_A_286_367#_c_712_n N_A_630_367#_c_1971_n 0.00199111f $X=6.39 $Y=1.65
+ $X2=0 $Y2=0
cc_730 N_A_286_367#_c_748_n N_A_630_367#_c_1971_n 0.0112007f $X=6.515 $Y=1.725
+ $X2=0 $Y2=0
cc_731 N_A_286_367#_c_730_n N_A_630_367#_c_1971_n 0.031498f $X=6.39 $Y=1.515
+ $X2=0 $Y2=0
cc_732 N_A_286_367#_c_749_n N_A_630_367#_c_1975_n 0.0112007f $X=6.945 $Y=1.725
+ $X2=0 $Y2=0
cc_733 N_A_286_367#_c_750_n N_A_630_367#_c_1975_n 0.0112007f $X=7.375 $Y=1.725
+ $X2=0 $Y2=0
cc_734 N_A_286_367#_c_714_n N_A_630_367#_c_1975_n 0.0024034f $X=10.05 $Y=1.65
+ $X2=0 $Y2=0
cc_735 N_A_286_367#_c_728_n N_A_630_367#_c_1975_n 0.0328887f $X=9.615 $Y=1.51
+ $X2=0 $Y2=0
cc_736 N_A_286_367#_c_751_n N_A_630_367#_c_1979_n 0.0113207f $X=7.805 $Y=1.725
+ $X2=0 $Y2=0
cc_737 N_A_286_367#_c_752_n N_A_630_367#_c_1979_n 0.0113207f $X=8.255 $Y=1.725
+ $X2=0 $Y2=0
cc_738 N_A_286_367#_c_714_n N_A_630_367#_c_1979_n 0.00288408f $X=10.05 $Y=1.65
+ $X2=0 $Y2=0
cc_739 N_A_286_367#_c_728_n N_A_630_367#_c_1979_n 0.0343048f $X=9.615 $Y=1.51
+ $X2=0 $Y2=0
cc_740 N_A_286_367#_c_753_n N_A_630_367#_c_1983_n 0.0112007f $X=8.685 $Y=1.725
+ $X2=0 $Y2=0
cc_741 N_A_286_367#_c_754_n N_A_630_367#_c_1983_n 0.0112007f $X=9.115 $Y=1.725
+ $X2=0 $Y2=0
cc_742 N_A_286_367#_c_714_n N_A_630_367#_c_1983_n 0.0024034f $X=10.05 $Y=1.65
+ $X2=0 $Y2=0
cc_743 N_A_286_367#_c_728_n N_A_630_367#_c_1983_n 0.0328887f $X=9.615 $Y=1.51
+ $X2=0 $Y2=0
cc_744 N_A_286_367#_c_755_n N_A_630_367#_c_1987_n 0.0112007f $X=9.545 $Y=1.725
+ $X2=0 $Y2=0
cc_745 N_A_286_367#_c_756_n N_A_630_367#_c_1987_n 0.0144061f $X=9.975 $Y=1.725
+ $X2=0 $Y2=0
cc_746 N_A_286_367#_c_714_n N_A_630_367#_c_1987_n 0.00274341f $X=10.05 $Y=1.65
+ $X2=0 $Y2=0
cc_747 N_A_286_367#_c_728_n N_A_630_367#_c_1987_n 0.0178605f $X=9.615 $Y=1.51
+ $X2=0 $Y2=0
cc_748 N_A_286_367#_c_755_n N_A_630_367#_c_1991_n 6.75085e-19 $X=9.545 $Y=1.725
+ $X2=0 $Y2=0
cc_749 N_A_286_367#_c_756_n N_A_630_367#_c_1991_n 0.00382137f $X=9.975 $Y=1.725
+ $X2=0 $Y2=0
cc_750 N_A_286_367#_c_713_n N_A_630_367#_c_1991_n 0.00473883f $X=10.33 $Y=1.65
+ $X2=0 $Y2=0
cc_751 N_A_286_367#_c_714_n N_A_630_367#_c_1991_n 0.00297916f $X=10.05 $Y=1.65
+ $X2=0 $Y2=0
cc_752 N_A_286_367#_c_759_n N_A_630_367#_c_1991_n 0.00335948f $X=10.405 $Y=1.725
+ $X2=0 $Y2=0
cc_753 N_A_286_367#_c_761_n N_A_630_367#_c_1991_n 2.76623e-19 $X=10.835 $Y=1.725
+ $X2=0 $Y2=0
cc_754 N_A_286_367#_c_724_n N_A_630_367#_c_1991_n 0.00240982f $X=10.405 $Y=1.65
+ $X2=0 $Y2=0
cc_755 N_A_286_367#_c_728_n N_A_630_367#_c_1991_n 0.00288855f $X=9.615 $Y=1.51
+ $X2=0 $Y2=0
cc_756 N_A_286_367#_c_755_n N_A_630_367#_c_1999_n 6.78151e-19 $X=9.545 $Y=1.725
+ $X2=0 $Y2=0
cc_757 N_A_286_367#_c_756_n N_A_630_367#_c_1999_n 0.0135317f $X=9.975 $Y=1.725
+ $X2=0 $Y2=0
cc_758 N_A_286_367#_c_759_n N_A_630_367#_c_1999_n 0.0125271f $X=10.405 $Y=1.725
+ $X2=0 $Y2=0
cc_759 N_A_286_367#_c_715_n N_A_630_367#_c_1937_n 0.0107968f $X=10.76 $Y=1.65
+ $X2=0 $Y2=0
cc_760 N_A_286_367#_c_716_n N_A_630_367#_c_1937_n 0.00427623f $X=11.19 $Y=1.65
+ $X2=0 $Y2=0
cc_761 N_A_286_367#_c_724_n N_A_630_367#_c_1937_n 0.00735656f $X=10.405 $Y=1.65
+ $X2=0 $Y2=0
cc_762 N_A_286_367#_c_725_n N_A_630_367#_c_1937_n 0.00773704f $X=10.835 $Y=1.65
+ $X2=0 $Y2=0
cc_763 N_A_286_367#_c_713_n N_A_630_367#_c_1938_n 0.00419267f $X=10.33 $Y=1.65
+ $X2=0 $Y2=0
cc_764 N_A_286_367#_c_714_n N_A_630_367#_c_1938_n 0.0022608f $X=10.05 $Y=1.65
+ $X2=0 $Y2=0
cc_765 N_A_286_367#_c_724_n N_A_630_367#_c_1938_n 3.80481e-19 $X=10.405 $Y=1.65
+ $X2=0 $Y2=0
cc_766 N_A_286_367#_c_728_n N_A_630_367#_c_1938_n 0.0112293f $X=9.615 $Y=1.51
+ $X2=0 $Y2=0
cc_767 N_A_286_367#_c_759_n N_A_630_367#_c_1939_n 3.05764e-19 $X=10.405 $Y=1.725
+ $X2=0 $Y2=0
cc_768 N_A_286_367#_c_761_n N_A_630_367#_c_1939_n 0.00402916f $X=10.835 $Y=1.725
+ $X2=0 $Y2=0
cc_769 N_A_286_367#_c_716_n N_A_630_367#_c_1939_n 0.00551306f $X=11.19 $Y=1.65
+ $X2=0 $Y2=0
cc_770 N_A_286_367#_c_763_n N_A_630_367#_c_1939_n 0.00178495f $X=11.265 $Y=1.725
+ $X2=0 $Y2=0
cc_771 N_A_286_367#_c_725_n N_A_630_367#_c_1939_n 0.00240982f $X=10.835 $Y=1.65
+ $X2=0 $Y2=0
cc_772 N_A_286_367#_c_761_n N_A_630_367#_c_2015_n 0.0104717f $X=10.835 $Y=1.725
+ $X2=0 $Y2=0
cc_773 N_A_286_367#_c_763_n N_A_630_367#_c_1940_n 0.0200111f $X=11.265 $Y=1.725
+ $X2=0 $Y2=0
cc_774 N_A_286_367#_c_731_n N_A_630_367#_c_2017_n 0.0122836f $X=3.075 $Y=1.725
+ $X2=0 $Y2=0
cc_775 N_A_286_367#_c_704_n N_A_630_367#_c_2017_n 0.00208864f $X=3.43 $Y=1.65
+ $X2=0 $Y2=0
cc_776 N_A_286_367#_c_734_n N_A_630_367#_c_2017_n 0.0119767f $X=3.505 $Y=1.725
+ $X2=0 $Y2=0
cc_777 N_A_286_367#_c_736_n N_A_630_367#_c_2017_n 5.93278e-19 $X=3.935 $Y=1.725
+ $X2=0 $Y2=0
cc_778 N_A_286_367#_c_730_n N_A_630_367#_c_2017_n 0.0197346f $X=6.39 $Y=1.515
+ $X2=0 $Y2=0
cc_779 N_A_286_367#_c_734_n N_A_630_367#_c_2022_n 5.93278e-19 $X=3.505 $Y=1.725
+ $X2=0 $Y2=0
cc_780 N_A_286_367#_c_736_n N_A_630_367#_c_2022_n 0.0119767f $X=3.935 $Y=1.725
+ $X2=0 $Y2=0
cc_781 N_A_286_367#_c_707_n N_A_630_367#_c_2022_n 0.00208864f $X=4.29 $Y=1.65
+ $X2=0 $Y2=0
cc_782 N_A_286_367#_c_738_n N_A_630_367#_c_2022_n 0.0119767f $X=4.365 $Y=1.725
+ $X2=0 $Y2=0
cc_783 N_A_286_367#_c_740_n N_A_630_367#_c_2022_n 5.93278e-19 $X=4.795 $Y=1.725
+ $X2=0 $Y2=0
cc_784 N_A_286_367#_c_730_n N_A_630_367#_c_2022_n 0.0197346f $X=6.39 $Y=1.515
+ $X2=0 $Y2=0
cc_785 N_A_286_367#_c_738_n N_A_630_367#_c_2028_n 5.93278e-19 $X=4.365 $Y=1.725
+ $X2=0 $Y2=0
cc_786 N_A_286_367#_c_740_n N_A_630_367#_c_2028_n 0.0119767f $X=4.795 $Y=1.725
+ $X2=0 $Y2=0
cc_787 N_A_286_367#_c_709_n N_A_630_367#_c_2028_n 0.00208864f $X=5.15 $Y=1.65
+ $X2=0 $Y2=0
cc_788 N_A_286_367#_c_742_n N_A_630_367#_c_2028_n 0.0119767f $X=5.225 $Y=1.725
+ $X2=0 $Y2=0
cc_789 N_A_286_367#_c_744_n N_A_630_367#_c_2028_n 5.93278e-19 $X=5.655 $Y=1.725
+ $X2=0 $Y2=0
cc_790 N_A_286_367#_c_730_n N_A_630_367#_c_2028_n 0.0197346f $X=6.39 $Y=1.515
+ $X2=0 $Y2=0
cc_791 N_A_286_367#_c_742_n N_A_630_367#_c_2034_n 5.93278e-19 $X=5.225 $Y=1.725
+ $X2=0 $Y2=0
cc_792 N_A_286_367#_c_744_n N_A_630_367#_c_2034_n 0.0119767f $X=5.655 $Y=1.725
+ $X2=0 $Y2=0
cc_793 N_A_286_367#_c_711_n N_A_630_367#_c_2034_n 0.00208864f $X=6.01 $Y=1.65
+ $X2=0 $Y2=0
cc_794 N_A_286_367#_c_746_n N_A_630_367#_c_2034_n 0.0119767f $X=6.085 $Y=1.725
+ $X2=0 $Y2=0
cc_795 N_A_286_367#_c_748_n N_A_630_367#_c_2034_n 5.93278e-19 $X=6.515 $Y=1.725
+ $X2=0 $Y2=0
cc_796 N_A_286_367#_c_730_n N_A_630_367#_c_2034_n 0.0197346f $X=6.39 $Y=1.515
+ $X2=0 $Y2=0
cc_797 N_A_286_367#_c_746_n N_A_630_367#_c_2040_n 5.93278e-19 $X=6.085 $Y=1.725
+ $X2=0 $Y2=0
cc_798 N_A_286_367#_c_748_n N_A_630_367#_c_2040_n 0.0119922f $X=6.515 $Y=1.725
+ $X2=0 $Y2=0
cc_799 N_A_286_367#_c_749_n N_A_630_367#_c_2040_n 0.0119922f $X=6.945 $Y=1.725
+ $X2=0 $Y2=0
cc_800 N_A_286_367#_c_750_n N_A_630_367#_c_2040_n 5.93278e-19 $X=7.375 $Y=1.725
+ $X2=0 $Y2=0
cc_801 N_A_286_367#_c_714_n N_A_630_367#_c_2040_n 0.00250138f $X=10.05 $Y=1.65
+ $X2=0 $Y2=0
cc_802 N_A_286_367#_c_728_n N_A_630_367#_c_2040_n 0.0210041f $X=9.615 $Y=1.51
+ $X2=0 $Y2=0
cc_803 N_A_286_367#_c_749_n N_A_630_367#_c_2046_n 5.93278e-19 $X=6.945 $Y=1.725
+ $X2=0 $Y2=0
cc_804 N_A_286_367#_c_750_n N_A_630_367#_c_2046_n 0.0119922f $X=7.375 $Y=1.725
+ $X2=0 $Y2=0
cc_805 N_A_286_367#_c_751_n N_A_630_367#_c_2046_n 0.0120839f $X=7.805 $Y=1.725
+ $X2=0 $Y2=0
cc_806 N_A_286_367#_c_752_n N_A_630_367#_c_2046_n 5.90833e-19 $X=8.255 $Y=1.725
+ $X2=0 $Y2=0
cc_807 N_A_286_367#_c_714_n N_A_630_367#_c_2046_n 0.00250138f $X=10.05 $Y=1.65
+ $X2=0 $Y2=0
cc_808 N_A_286_367#_c_728_n N_A_630_367#_c_2046_n 0.0210041f $X=9.615 $Y=1.51
+ $X2=0 $Y2=0
cc_809 N_A_286_367#_c_751_n N_A_630_367#_c_2052_n 6.07264e-19 $X=7.805 $Y=1.725
+ $X2=0 $Y2=0
cc_810 N_A_286_367#_c_752_n N_A_630_367#_c_2052_n 0.0123432f $X=8.255 $Y=1.725
+ $X2=0 $Y2=0
cc_811 N_A_286_367#_c_753_n N_A_630_367#_c_2052_n 0.0119922f $X=8.685 $Y=1.725
+ $X2=0 $Y2=0
cc_812 N_A_286_367#_c_754_n N_A_630_367#_c_2052_n 5.93278e-19 $X=9.115 $Y=1.725
+ $X2=0 $Y2=0
cc_813 N_A_286_367#_c_714_n N_A_630_367#_c_2052_n 0.00250138f $X=10.05 $Y=1.65
+ $X2=0 $Y2=0
cc_814 N_A_286_367#_c_728_n N_A_630_367#_c_2052_n 0.0210041f $X=9.615 $Y=1.51
+ $X2=0 $Y2=0
cc_815 N_A_286_367#_c_753_n N_A_630_367#_c_2058_n 5.93278e-19 $X=8.685 $Y=1.725
+ $X2=0 $Y2=0
cc_816 N_A_286_367#_c_754_n N_A_630_367#_c_2058_n 0.0119922f $X=9.115 $Y=1.725
+ $X2=0 $Y2=0
cc_817 N_A_286_367#_c_755_n N_A_630_367#_c_2058_n 0.0119922f $X=9.545 $Y=1.725
+ $X2=0 $Y2=0
cc_818 N_A_286_367#_c_756_n N_A_630_367#_c_2058_n 5.93278e-19 $X=9.975 $Y=1.725
+ $X2=0 $Y2=0
cc_819 N_A_286_367#_c_714_n N_A_630_367#_c_2058_n 0.00250138f $X=10.05 $Y=1.65
+ $X2=0 $Y2=0
cc_820 N_A_286_367#_c_728_n N_A_630_367#_c_2058_n 0.0210041f $X=9.615 $Y=1.51
+ $X2=0 $Y2=0
cc_821 N_A_286_367#_c_756_n N_A_630_367#_c_2064_n 3.84191e-19 $X=9.975 $Y=1.725
+ $X2=0 $Y2=0
cc_822 N_A_286_367#_c_759_n N_A_630_367#_c_2064_n 0.0017646f $X=10.405 $Y=1.725
+ $X2=0 $Y2=0
cc_823 N_A_286_367#_c_761_n N_A_630_367#_c_2066_n 0.00245588f $X=10.835 $Y=1.725
+ $X2=0 $Y2=0
cc_824 N_A_286_367#_c_713_n N_Z_c_2279_n 7.6834e-19 $X=10.33 $Y=1.65 $X2=0 $Y2=0
cc_825 N_A_286_367#_c_714_n N_Z_c_2279_n 0.0016813f $X=10.05 $Y=1.65 $X2=0 $Y2=0
cc_826 N_A_286_367#_c_715_n N_Z_c_2279_n 7.69474e-19 $X=10.76 $Y=1.65 $X2=0
+ $Y2=0
cc_827 N_A_286_367#_c_716_n N_Z_c_2279_n 0.00158576f $X=11.19 $Y=1.65 $X2=0
+ $Y2=0
cc_828 N_A_286_367#_c_728_n N_Z_c_2279_n 0.00112414f $X=9.615 $Y=1.51 $X2=0
+ $Y2=0
cc_829 N_A_286_367#_c_716_n N_Z_c_2281_n 0.00702114f $X=11.19 $Y=1.65 $X2=0
+ $Y2=0
cc_830 N_A_286_367#_c_763_n N_Z_c_2281_n 0.00241354f $X=11.265 $Y=1.725 $X2=0
+ $Y2=0
cc_831 N_A_286_367#_M1010_s N_VGND_c_2515_n 0.00590798f $X=1.59 $Y=0.235 $X2=0
+ $Y2=0
cc_832 N_A_286_367#_c_714_n N_A_584_47#_c_2757_n 7.01567e-19 $X=10.05 $Y=1.65
+ $X2=0 $Y2=0
cc_833 N_A_286_367#_c_727_n N_A_584_47#_c_2757_n 0.00713351f $X=6.56 $Y=1.515
+ $X2=0 $Y2=0
cc_834 N_A_286_367#_c_714_n N_A_584_47#_c_2724_n 0.00305992f $X=10.05 $Y=1.65
+ $X2=0 $Y2=0
cc_835 N_A_286_367#_c_728_n N_A_584_47#_c_2724_n 0.0381685f $X=9.615 $Y=1.51
+ $X2=0 $Y2=0
cc_836 N_A_286_367#_c_714_n N_A_584_47#_c_2725_n 0.00218312f $X=10.05 $Y=1.65
+ $X2=0 $Y2=0
cc_837 N_A_286_367#_c_728_n N_A_584_47#_c_2725_n 0.0267119f $X=9.615 $Y=1.51
+ $X2=0 $Y2=0
cc_838 N_A_286_367#_c_714_n N_A_584_47#_c_2726_n 0.00305014f $X=10.05 $Y=1.65
+ $X2=0 $Y2=0
cc_839 N_A_286_367#_c_728_n N_A_584_47#_c_2726_n 0.0381685f $X=9.615 $Y=1.51
+ $X2=0 $Y2=0
cc_840 N_A_286_367#_c_714_n N_A_584_47#_c_2727_n 0.0106566f $X=10.05 $Y=1.65
+ $X2=0 $Y2=0
cc_841 N_A_286_367#_c_728_n N_A_584_47#_c_2727_n 0.0648805f $X=9.615 $Y=1.51
+ $X2=0 $Y2=0
cc_842 N_A_286_367#_c_714_n N_A_584_47#_c_2728_n 0.00218312f $X=10.05 $Y=1.65
+ $X2=0 $Y2=0
cc_843 N_A_286_367#_c_728_n N_A_584_47#_c_2728_n 0.0267119f $X=9.615 $Y=1.51
+ $X2=0 $Y2=0
cc_844 N_A_286_367#_c_714_n N_A_584_47#_c_2729_n 0.00218312f $X=10.05 $Y=1.65
+ $X2=0 $Y2=0
cc_845 N_A_286_367#_c_728_n N_A_584_47#_c_2729_n 0.0267119f $X=9.615 $Y=1.51
+ $X2=0 $Y2=0
cc_846 N_A_1909_21#_c_1118_p N_A_M1009_g 0.0149753f $X=21.645 $Y=1.98 $X2=0
+ $Y2=0
cc_847 N_A_1909_21#_c_1119_p N_A_M1009_g 0.00450851f $X=21.645 $Y=1.78 $X2=0
+ $Y2=0
cc_848 N_A_1909_21#_c_1080_n N_A_c_1479_n 0.0079007f $X=21.565 $Y=1.695 $X2=0
+ $Y2=0
cc_849 N_A_1909_21#_c_1121_p N_A_c_1479_n 0.00336446f $X=22.03 $Y=0.915 $X2=0
+ $Y2=0
cc_850 N_A_1909_21#_c_1119_p N_A_c_1479_n 0.00870347f $X=21.645 $Y=1.78 $X2=0
+ $Y2=0
cc_851 N_A_1909_21#_c_1078_n N_A_c_1480_n 0.00260673f $X=21.48 $Y=1.15 $X2=0
+ $Y2=0
cc_852 N_A_1909_21#_c_1079_n N_A_c_1480_n 0.00465205f $X=21.265 $Y=1.15 $X2=0
+ $Y2=0
cc_853 N_A_1909_21#_c_1080_n N_A_c_1480_n 0.00369289f $X=21.565 $Y=1.695 $X2=0
+ $Y2=0
cc_854 N_A_1909_21#_c_1119_p N_A_c_1480_n 2.22784e-19 $X=21.645 $Y=1.78 $X2=0
+ $Y2=0
cc_855 N_A_1909_21#_c_1118_p N_A_M1014_g 0.0164109f $X=21.645 $Y=1.98 $X2=0
+ $Y2=0
cc_856 N_A_1909_21#_c_1103_n N_A_M1014_g 0.00921648f $X=22.34 $Y=1.78 $X2=0
+ $Y2=0
cc_857 N_A_1909_21#_c_1129_p N_A_M1014_g 0.00108612f $X=22.505 $Y=1.98 $X2=0
+ $Y2=0
cc_858 N_A_1909_21#_c_1119_p N_A_M1014_g 0.00190031f $X=21.645 $Y=1.78 $X2=0
+ $Y2=0
cc_859 N_A_1909_21#_c_1079_n N_A_c_1481_n 0.00867997f $X=21.265 $Y=1.15 $X2=0
+ $Y2=0
cc_860 N_A_1909_21#_c_1121_p N_A_c_1481_n 0.0137301f $X=22.03 $Y=0.915 $X2=0
+ $Y2=0
cc_861 N_A_1909_21#_c_1081_n N_A_c_1481_n 0.00572835f $X=21.565 $Y=1.072 $X2=0
+ $Y2=0
cc_862 N_A_1909_21#_c_1080_n N_A_M1034_g 5.18796e-19 $X=21.565 $Y=1.695 $X2=0
+ $Y2=0
cc_863 N_A_1909_21#_c_1118_p N_A_M1034_g 0.00108612f $X=21.645 $Y=1.98 $X2=0
+ $Y2=0
cc_864 N_A_1909_21#_c_1103_n N_A_M1034_g 0.0112007f $X=22.34 $Y=1.78 $X2=0 $Y2=0
cc_865 N_A_1909_21#_c_1129_p N_A_M1034_g 0.0164109f $X=22.505 $Y=1.98 $X2=0
+ $Y2=0
cc_866 N_A_1909_21#_c_1106_n N_A_M1034_g 0.0024309f $X=22.505 $Y=1.78 $X2=0
+ $Y2=0
cc_867 N_A_1909_21#_c_1139_p N_A_c_1483_n 0.00848459f $X=22.195 $Y=0.38 $X2=0
+ $Y2=0
cc_868 N_A_1909_21#_c_1140_p N_A_c_1483_n 0.00947623f $X=23.05 $Y=0.915 $X2=0
+ $Y2=0
cc_869 N_A_1909_21#_c_1141_p N_A_c_1483_n 8.8778e-19 $X=23.215 $Y=0.43 $X2=0
+ $Y2=0
cc_870 N_A_1909_21#_c_1142_p N_A_c_1483_n 7.2817e-19 $X=22.195 $Y=0.915 $X2=0
+ $Y2=0
cc_871 N_A_1909_21#_c_1129_p N_A_M1052_g 0.0155573f $X=22.505 $Y=1.98 $X2=0
+ $Y2=0
cc_872 N_A_1909_21#_c_1104_n N_A_M1052_g 0.0112007f $X=23.2 $Y=1.78 $X2=0 $Y2=0
cc_873 N_A_1909_21#_c_1145_p N_A_M1052_g 7.68674e-19 $X=23.365 $Y=1.98 $X2=0
+ $Y2=0
cc_874 N_A_1909_21#_c_1106_n N_A_M1052_g 0.0024309f $X=22.505 $Y=1.78 $X2=0
+ $Y2=0
cc_875 N_A_1909_21#_c_1139_p N_A_c_1485_n 8.81771e-19 $X=22.195 $Y=0.38 $X2=0
+ $Y2=0
cc_876 N_A_1909_21#_c_1140_p N_A_c_1485_n 0.0102188f $X=23.05 $Y=0.915 $X2=0
+ $Y2=0
cc_877 N_A_1909_21#_c_1141_p N_A_c_1485_n 0.00815878f $X=23.215 $Y=0.43 $X2=0
+ $Y2=0
cc_878 N_A_1909_21#_c_1129_p N_A_M1072_g 7.68674e-19 $X=22.505 $Y=1.98 $X2=0
+ $Y2=0
cc_879 N_A_1909_21#_c_1104_n N_A_M1072_g 0.0112007f $X=23.2 $Y=1.78 $X2=0 $Y2=0
cc_880 N_A_1909_21#_c_1145_p N_A_M1072_g 0.0155573f $X=23.365 $Y=1.98 $X2=0
+ $Y2=0
cc_881 N_A_1909_21#_c_1107_n N_A_M1072_g 0.0024309f $X=23.365 $Y=1.78 $X2=0
+ $Y2=0
cc_882 N_A_1909_21#_c_1140_p N_A_c_1487_n 0.00222052f $X=23.05 $Y=0.915 $X2=0
+ $Y2=0
cc_883 N_A_1909_21#_c_1141_p N_A_c_1487_n 0.00654194f $X=23.215 $Y=0.43 $X2=0
+ $Y2=0
cc_884 N_A_1909_21#_c_1145_p N_A_M1076_g 0.0156985f $X=23.365 $Y=1.98 $X2=0
+ $Y2=0
cc_885 N_A_1909_21#_c_1105_n N_A_M1076_g 0.0113497f $X=24.085 $Y=1.78 $X2=0
+ $Y2=0
cc_886 N_A_1909_21#_c_1158_p N_A_M1076_g 7.93352e-19 $X=24.25 $Y=1.98 $X2=0
+ $Y2=0
cc_887 N_A_1909_21#_c_1107_n N_A_M1076_g 0.0024309f $X=23.365 $Y=1.78 $X2=0
+ $Y2=0
cc_888 N_A_1909_21#_c_1145_p N_A_M1079_g 7.56713e-19 $X=23.365 $Y=1.98 $X2=0
+ $Y2=0
cc_889 N_A_1909_21#_c_1105_n N_A_M1079_g 0.0137806f $X=24.085 $Y=1.78 $X2=0
+ $Y2=0
cc_890 N_A_1909_21#_c_1158_p N_A_M1079_g 0.0162907f $X=24.25 $Y=1.98 $X2=0 $Y2=0
cc_891 N_A_1909_21#_c_1105_n N_A_M1085_g 0.00824344f $X=24.085 $Y=1.78 $X2=0
+ $Y2=0
cc_892 N_A_1909_21#_c_1158_p N_A_M1085_g 0.0149753f $X=24.25 $Y=1.98 $X2=0 $Y2=0
cc_893 N_A_1909_21#_c_1080_n A 0.0151895f $X=21.565 $Y=1.695 $X2=0 $Y2=0
cc_894 N_A_1909_21#_c_1121_p A 0.0122485f $X=22.03 $Y=0.915 $X2=0 $Y2=0
cc_895 N_A_1909_21#_c_1103_n A 0.0358586f $X=22.34 $Y=1.78 $X2=0 $Y2=0
cc_896 N_A_1909_21#_c_1140_p A 0.0681321f $X=23.05 $Y=0.915 $X2=0 $Y2=0
cc_897 N_A_1909_21#_c_1104_n A 0.0371921f $X=23.2 $Y=1.78 $X2=0 $Y2=0
cc_898 N_A_1909_21#_c_1105_n A 0.0654549f $X=24.085 $Y=1.78 $X2=0 $Y2=0
cc_899 N_A_1909_21#_c_1081_n A 0.0113982f $X=21.565 $Y=1.072 $X2=0 $Y2=0
cc_900 N_A_1909_21#_c_1142_p A 0.0245648f $X=22.195 $Y=0.915 $X2=0 $Y2=0
cc_901 N_A_1909_21#_c_1106_n A 0.026461f $X=22.505 $Y=1.78 $X2=0 $Y2=0
cc_902 N_A_1909_21#_c_1107_n A 0.026461f $X=23.365 $Y=1.78 $X2=0 $Y2=0
cc_903 N_A_1909_21#_c_1080_n N_A_c_1492_n 0.0059146f $X=21.565 $Y=1.695 $X2=0
+ $Y2=0
cc_904 N_A_1909_21#_c_1103_n N_A_c_1492_n 0.00486222f $X=22.34 $Y=1.78 $X2=0
+ $Y2=0
cc_905 N_A_1909_21#_c_1140_p N_A_c_1492_n 0.00253182f $X=23.05 $Y=0.915 $X2=0
+ $Y2=0
cc_906 N_A_1909_21#_c_1104_n N_A_c_1492_n 0.00261742f $X=23.2 $Y=1.78 $X2=0
+ $Y2=0
cc_907 N_A_1909_21#_c_1105_n N_A_c_1492_n 0.00510265f $X=24.085 $Y=1.78 $X2=0
+ $Y2=0
cc_908 N_A_1909_21#_c_1119_p N_A_c_1492_n 0.00120528f $X=21.645 $Y=1.78 $X2=0
+ $Y2=0
cc_909 N_A_1909_21#_c_1142_p N_A_c_1492_n 0.00134539f $X=22.195 $Y=0.915 $X2=0
+ $Y2=0
cc_910 N_A_1909_21#_c_1106_n N_A_c_1492_n 0.00270827f $X=22.505 $Y=1.78 $X2=0
+ $Y2=0
cc_911 N_A_1909_21#_c_1107_n N_A_c_1492_n 0.00270827f $X=23.365 $Y=1.78 $X2=0
+ $Y2=0
cc_912 N_A_1909_21#_c_1103_n N_VPWR_M1014_d 0.00229297f $X=22.34 $Y=1.78 $X2=0
+ $Y2=0
cc_913 N_A_1909_21#_c_1104_n N_VPWR_M1052_d 0.00180746f $X=23.2 $Y=1.78 $X2=0
+ $Y2=0
cc_914 N_A_1909_21#_c_1105_n N_VPWR_M1076_d 0.00273408f $X=24.085 $Y=1.78 $X2=0
+ $Y2=0
cc_915 N_A_1909_21#_M1000_g N_VPWR_c_1629_n 0.00865603f $X=12.27 $Y=2.155 $X2=0
+ $Y2=0
cc_916 N_A_1909_21#_M1088_g N_VPWR_c_1630_n 0.00333514f $X=20.44 $Y=2.155 $X2=0
+ $Y2=0
cc_917 N_A_1909_21#_c_1078_n N_VPWR_c_1630_n 0.00933279f $X=21.48 $Y=1.15 $X2=0
+ $Y2=0
cc_918 N_A_1909_21#_c_1079_n N_VPWR_c_1630_n 0.0046469f $X=21.265 $Y=1.15 $X2=0
+ $Y2=0
cc_919 N_A_1909_21#_c_1119_p N_VPWR_c_1630_n 0.00274213f $X=21.645 $Y=1.78 $X2=0
+ $Y2=0
cc_920 N_A_1909_21#_c_1103_n N_VPWR_c_1631_n 0.00887783f $X=22.34 $Y=1.78 $X2=0
+ $Y2=0
cc_921 N_A_1909_21#_c_1104_n N_VPWR_c_1632_n 0.0129403f $X=23.2 $Y=1.78 $X2=0
+ $Y2=0
cc_922 N_A_1909_21#_c_1145_p N_VPWR_c_1633_n 0.0177952f $X=23.365 $Y=1.98 $X2=0
+ $Y2=0
cc_923 N_A_1909_21#_c_1105_n N_VPWR_c_1634_n 0.0130182f $X=24.085 $Y=1.78 $X2=0
+ $Y2=0
cc_924 N_A_1909_21#_c_1158_p N_VPWR_c_1634_n 0.0651913f $X=24.25 $Y=1.98 $X2=0
+ $Y2=0
cc_925 N_A_1909_21#_c_1105_n N_VPWR_c_1636_n 0.00274213f $X=24.085 $Y=1.78 $X2=0
+ $Y2=0
cc_926 N_A_1909_21#_M1000_g N_VPWR_c_1659_n 0.00394144f $X=12.27 $Y=2.155 $X2=0
+ $Y2=0
cc_927 N_A_1909_21#_M1002_g N_VPWR_c_1659_n 6.63248e-19 $X=12.7 $Y=2.155 $X2=0
+ $Y2=0
cc_928 N_A_1909_21#_M1006_g N_VPWR_c_1659_n 6.63248e-19 $X=13.13 $Y=2.155 $X2=0
+ $Y2=0
cc_929 N_A_1909_21#_M1008_g N_VPWR_c_1659_n 6.63248e-19 $X=13.56 $Y=2.155 $X2=0
+ $Y2=0
cc_930 N_A_1909_21#_M1013_g N_VPWR_c_1659_n 6.63248e-19 $X=13.99 $Y=2.155 $X2=0
+ $Y2=0
cc_931 N_A_1909_21#_M1023_g N_VPWR_c_1659_n 6.63248e-19 $X=14.42 $Y=2.155 $X2=0
+ $Y2=0
cc_932 N_A_1909_21#_M1025_g N_VPWR_c_1659_n 6.63248e-19 $X=14.85 $Y=2.155 $X2=0
+ $Y2=0
cc_933 N_A_1909_21#_M1026_g N_VPWR_c_1659_n 6.63248e-19 $X=15.28 $Y=2.155 $X2=0
+ $Y2=0
cc_934 N_A_1909_21#_M1030_g N_VPWR_c_1659_n 6.63248e-19 $X=15.71 $Y=2.155 $X2=0
+ $Y2=0
cc_935 N_A_1909_21#_M1032_g N_VPWR_c_1659_n 6.63248e-19 $X=16.14 $Y=2.155 $X2=0
+ $Y2=0
cc_936 N_A_1909_21#_M1038_g N_VPWR_c_1659_n 6.63248e-19 $X=16.57 $Y=2.155 $X2=0
+ $Y2=0
cc_937 N_A_1909_21#_M1042_g N_VPWR_c_1659_n 6.63248e-19 $X=17 $Y=2.155 $X2=0
+ $Y2=0
cc_938 N_A_1909_21#_M1046_g N_VPWR_c_1659_n 6.63248e-19 $X=17.43 $Y=2.155 $X2=0
+ $Y2=0
cc_939 N_A_1909_21#_M1050_g N_VPWR_c_1659_n 6.63248e-19 $X=17.86 $Y=2.155 $X2=0
+ $Y2=0
cc_940 N_A_1909_21#_M1056_g N_VPWR_c_1659_n 6.63248e-19 $X=18.29 $Y=2.155 $X2=0
+ $Y2=0
cc_941 N_A_1909_21#_M1062_g N_VPWR_c_1659_n 6.63248e-19 $X=18.72 $Y=2.155 $X2=0
+ $Y2=0
cc_942 N_A_1909_21#_M1063_g N_VPWR_c_1659_n 6.63248e-19 $X=19.15 $Y=2.155 $X2=0
+ $Y2=0
cc_943 N_A_1909_21#_M1075_g N_VPWR_c_1659_n 6.63248e-19 $X=19.58 $Y=2.155 $X2=0
+ $Y2=0
cc_944 N_A_1909_21#_M1078_g N_VPWR_c_1659_n 6.63248e-19 $X=20.01 $Y=2.155 $X2=0
+ $Y2=0
cc_945 N_A_1909_21#_M1088_g N_VPWR_c_1659_n 0.00394144f $X=20.44 $Y=2.155 $X2=0
+ $Y2=0
cc_946 N_A_1909_21#_c_1118_p N_VPWR_c_1661_n 0.0177952f $X=21.645 $Y=1.98 $X2=0
+ $Y2=0
cc_947 N_A_1909_21#_c_1129_p N_VPWR_c_1663_n 0.0177952f $X=22.505 $Y=1.98 $X2=0
+ $Y2=0
cc_948 N_A_1909_21#_c_1158_p N_VPWR_c_1665_n 0.0177952f $X=24.25 $Y=1.98 $X2=0
+ $Y2=0
cc_949 N_A_1909_21#_M1009_s N_VPWR_c_1612_n 0.00223819f $X=21.505 $Y=1.835 $X2=0
+ $Y2=0
cc_950 N_A_1909_21#_M1034_s N_VPWR_c_1612_n 0.00223819f $X=22.365 $Y=1.835 $X2=0
+ $Y2=0
cc_951 N_A_1909_21#_M1072_s N_VPWR_c_1612_n 0.00223819f $X=23.225 $Y=1.835 $X2=0
+ $Y2=0
cc_952 N_A_1909_21#_M1079_s N_VPWR_c_1612_n 0.00223819f $X=24.11 $Y=1.835 $X2=0
+ $Y2=0
cc_953 N_A_1909_21#_M1000_g N_VPWR_c_1612_n 0.00410091f $X=12.27 $Y=2.155 $X2=0
+ $Y2=0
cc_954 N_A_1909_21#_M1088_g N_VPWR_c_1612_n 0.00410091f $X=20.44 $Y=2.155 $X2=0
+ $Y2=0
cc_955 N_A_1909_21#_c_1118_p N_VPWR_c_1612_n 0.0123247f $X=21.645 $Y=1.98 $X2=0
+ $Y2=0
cc_956 N_A_1909_21#_c_1129_p N_VPWR_c_1612_n 0.0123247f $X=22.505 $Y=1.98 $X2=0
+ $Y2=0
cc_957 N_A_1909_21#_c_1145_p N_VPWR_c_1612_n 0.0123247f $X=23.365 $Y=1.98 $X2=0
+ $Y2=0
cc_958 N_A_1909_21#_c_1158_p N_VPWR_c_1612_n 0.0123247f $X=24.25 $Y=1.98 $X2=0
+ $Y2=0
cc_959 N_A_1909_21#_c_1037_n N_A_630_367#_c_1937_n 0.00495394f $X=10.565 $Y=1.06
+ $X2=0 $Y2=0
cc_960 N_A_1909_21#_c_1039_n N_A_630_367#_c_1937_n 0.00279834f $X=11.075 $Y=1.06
+ $X2=0 $Y2=0
cc_961 N_A_1909_21#_c_1034_n N_A_630_367#_c_1938_n 0.00380458f $X=10.055 $Y=1.06
+ $X2=0 $Y2=0
cc_962 N_A_1909_21#_M1000_g N_A_630_367#_c_1940_n 0.015395f $X=12.27 $Y=2.155
+ $X2=0 $Y2=0
cc_963 N_A_1909_21#_c_1082_n N_A_630_367#_c_1940_n 6.82908e-19 $X=20.515 $Y=1.15
+ $X2=0 $Y2=0
cc_964 N_A_1909_21#_M1000_g N_A_630_367#_c_2072_n 8.66862e-19 $X=12.27 $Y=2.155
+ $X2=0 $Y2=0
cc_965 N_A_1909_21#_M1002_g N_A_630_367#_c_2072_n 0.00264221f $X=12.7 $Y=2.155
+ $X2=0 $Y2=0
cc_966 N_A_1909_21#_M1000_g N_A_630_367#_c_2074_n 0.0220898f $X=12.27 $Y=2.155
+ $X2=0 $Y2=0
cc_967 N_A_1909_21#_M1002_g N_A_630_367#_c_2074_n 0.0109788f $X=12.7 $Y=2.155
+ $X2=0 $Y2=0
cc_968 N_A_1909_21#_M1006_g N_A_630_367#_c_2074_n 5.84508e-19 $X=13.13 $Y=2.155
+ $X2=0 $Y2=0
cc_969 N_A_1909_21#_M1002_g N_A_630_367#_c_1941_n 0.00835624f $X=12.7 $Y=2.155
+ $X2=0 $Y2=0
cc_970 N_A_1909_21#_M1006_g N_A_630_367#_c_1941_n 0.00835624f $X=13.13 $Y=2.155
+ $X2=0 $Y2=0
cc_971 N_A_1909_21#_M1000_g N_A_630_367#_c_1942_n 0.00147002f $X=12.27 $Y=2.155
+ $X2=0 $Y2=0
cc_972 N_A_1909_21#_M1002_g N_A_630_367#_c_1942_n 8.63014e-19 $X=12.7 $Y=2.155
+ $X2=0 $Y2=0
cc_973 N_A_1909_21#_M1002_g N_A_630_367#_c_2081_n 6.66834e-19 $X=12.7 $Y=2.155
+ $X2=0 $Y2=0
cc_974 N_A_1909_21#_M1006_g N_A_630_367#_c_2081_n 0.0127479f $X=13.13 $Y=2.155
+ $X2=0 $Y2=0
cc_975 N_A_1909_21#_M1008_g N_A_630_367#_c_2081_n 0.0127479f $X=13.56 $Y=2.155
+ $X2=0 $Y2=0
cc_976 N_A_1909_21#_M1013_g N_A_630_367#_c_2081_n 6.66834e-19 $X=13.99 $Y=2.155
+ $X2=0 $Y2=0
cc_977 N_A_1909_21#_M1008_g N_A_630_367#_c_1943_n 0.00835624f $X=13.56 $Y=2.155
+ $X2=0 $Y2=0
cc_978 N_A_1909_21#_M1013_g N_A_630_367#_c_1943_n 0.00835624f $X=13.99 $Y=2.155
+ $X2=0 $Y2=0
cc_979 N_A_1909_21#_M1008_g N_A_630_367#_c_2087_n 6.66834e-19 $X=13.56 $Y=2.155
+ $X2=0 $Y2=0
cc_980 N_A_1909_21#_M1013_g N_A_630_367#_c_2087_n 0.0127479f $X=13.99 $Y=2.155
+ $X2=0 $Y2=0
cc_981 N_A_1909_21#_M1023_g N_A_630_367#_c_2087_n 0.0127479f $X=14.42 $Y=2.155
+ $X2=0 $Y2=0
cc_982 N_A_1909_21#_M1025_g N_A_630_367#_c_2087_n 6.66834e-19 $X=14.85 $Y=2.155
+ $X2=0 $Y2=0
cc_983 N_A_1909_21#_M1023_g N_A_630_367#_c_1944_n 0.00835624f $X=14.42 $Y=2.155
+ $X2=0 $Y2=0
cc_984 N_A_1909_21#_M1025_g N_A_630_367#_c_1944_n 0.00835624f $X=14.85 $Y=2.155
+ $X2=0 $Y2=0
cc_985 N_A_1909_21#_M1023_g N_A_630_367#_c_2093_n 6.66834e-19 $X=14.42 $Y=2.155
+ $X2=0 $Y2=0
cc_986 N_A_1909_21#_M1025_g N_A_630_367#_c_2093_n 0.0127479f $X=14.85 $Y=2.155
+ $X2=0 $Y2=0
cc_987 N_A_1909_21#_M1026_g N_A_630_367#_c_2093_n 0.0127479f $X=15.28 $Y=2.155
+ $X2=0 $Y2=0
cc_988 N_A_1909_21#_M1030_g N_A_630_367#_c_2093_n 6.66834e-19 $X=15.71 $Y=2.155
+ $X2=0 $Y2=0
cc_989 N_A_1909_21#_M1026_g N_A_630_367#_c_1945_n 0.00835624f $X=15.28 $Y=2.155
+ $X2=0 $Y2=0
cc_990 N_A_1909_21#_M1030_g N_A_630_367#_c_1945_n 0.00835624f $X=15.71 $Y=2.155
+ $X2=0 $Y2=0
cc_991 N_A_1909_21#_M1026_g N_A_630_367#_c_2099_n 6.66834e-19 $X=15.28 $Y=2.155
+ $X2=0 $Y2=0
cc_992 N_A_1909_21#_M1030_g N_A_630_367#_c_2099_n 0.0127479f $X=15.71 $Y=2.155
+ $X2=0 $Y2=0
cc_993 N_A_1909_21#_M1032_g N_A_630_367#_c_2099_n 0.0127479f $X=16.14 $Y=2.155
+ $X2=0 $Y2=0
cc_994 N_A_1909_21#_M1038_g N_A_630_367#_c_2099_n 6.66834e-19 $X=16.57 $Y=2.155
+ $X2=0 $Y2=0
cc_995 N_A_1909_21#_M1032_g N_A_630_367#_c_1946_n 0.00835624f $X=16.14 $Y=2.155
+ $X2=0 $Y2=0
cc_996 N_A_1909_21#_M1038_g N_A_630_367#_c_1946_n 0.00835624f $X=16.57 $Y=2.155
+ $X2=0 $Y2=0
cc_997 N_A_1909_21#_M1032_g N_A_630_367#_c_2105_n 6.66834e-19 $X=16.14 $Y=2.155
+ $X2=0 $Y2=0
cc_998 N_A_1909_21#_M1038_g N_A_630_367#_c_2105_n 0.0127479f $X=16.57 $Y=2.155
+ $X2=0 $Y2=0
cc_999 N_A_1909_21#_M1042_g N_A_630_367#_c_2105_n 0.0127479f $X=17 $Y=2.155
+ $X2=0 $Y2=0
cc_1000 N_A_1909_21#_M1046_g N_A_630_367#_c_2105_n 6.66834e-19 $X=17.43 $Y=2.155
+ $X2=0 $Y2=0
cc_1001 N_A_1909_21#_M1042_g N_A_630_367#_c_1947_n 0.00835624f $X=17 $Y=2.155
+ $X2=0 $Y2=0
cc_1002 N_A_1909_21#_M1046_g N_A_630_367#_c_1947_n 0.00835624f $X=17.43 $Y=2.155
+ $X2=0 $Y2=0
cc_1003 N_A_1909_21#_M1042_g N_A_630_367#_c_2111_n 6.66834e-19 $X=17 $Y=2.155
+ $X2=0 $Y2=0
cc_1004 N_A_1909_21#_M1046_g N_A_630_367#_c_2111_n 0.0127479f $X=17.43 $Y=2.155
+ $X2=0 $Y2=0
cc_1005 N_A_1909_21#_M1050_g N_A_630_367#_c_2111_n 0.0127479f $X=17.86 $Y=2.155
+ $X2=0 $Y2=0
cc_1006 N_A_1909_21#_M1056_g N_A_630_367#_c_2111_n 6.66834e-19 $X=18.29 $Y=2.155
+ $X2=0 $Y2=0
cc_1007 N_A_1909_21#_M1050_g N_A_630_367#_c_1948_n 0.00835624f $X=17.86 $Y=2.155
+ $X2=0 $Y2=0
cc_1008 N_A_1909_21#_M1056_g N_A_630_367#_c_1948_n 0.00835624f $X=18.29 $Y=2.155
+ $X2=0 $Y2=0
cc_1009 N_A_1909_21#_M1050_g N_A_630_367#_c_2117_n 6.66834e-19 $X=17.86 $Y=2.155
+ $X2=0 $Y2=0
cc_1010 N_A_1909_21#_M1056_g N_A_630_367#_c_2117_n 0.0127479f $X=18.29 $Y=2.155
+ $X2=0 $Y2=0
cc_1011 N_A_1909_21#_M1062_g N_A_630_367#_c_2117_n 0.0127479f $X=18.72 $Y=2.155
+ $X2=0 $Y2=0
cc_1012 N_A_1909_21#_M1063_g N_A_630_367#_c_2117_n 6.66834e-19 $X=19.15 $Y=2.155
+ $X2=0 $Y2=0
cc_1013 N_A_1909_21#_M1062_g N_A_630_367#_c_1949_n 0.00835624f $X=18.72 $Y=2.155
+ $X2=0 $Y2=0
cc_1014 N_A_1909_21#_M1063_g N_A_630_367#_c_1949_n 0.00835624f $X=19.15 $Y=2.155
+ $X2=0 $Y2=0
cc_1015 N_A_1909_21#_M1062_g N_A_630_367#_c_2123_n 6.66834e-19 $X=18.72 $Y=2.155
+ $X2=0 $Y2=0
cc_1016 N_A_1909_21#_M1063_g N_A_630_367#_c_2123_n 0.0127479f $X=19.15 $Y=2.155
+ $X2=0 $Y2=0
cc_1017 N_A_1909_21#_M1075_g N_A_630_367#_c_2123_n 0.0127479f $X=19.58 $Y=2.155
+ $X2=0 $Y2=0
cc_1018 N_A_1909_21#_M1078_g N_A_630_367#_c_2123_n 6.66834e-19 $X=20.01 $Y=2.155
+ $X2=0 $Y2=0
cc_1019 N_A_1909_21#_M1075_g N_A_630_367#_c_1950_n 0.00835624f $X=19.58 $Y=2.155
+ $X2=0 $Y2=0
cc_1020 N_A_1909_21#_M1078_g N_A_630_367#_c_1950_n 0.00921926f $X=20.01 $Y=2.155
+ $X2=0 $Y2=0
cc_1021 N_A_1909_21#_M1088_g N_A_630_367#_c_1950_n 0.00146133f $X=20.44 $Y=2.155
+ $X2=0 $Y2=0
cc_1022 N_A_1909_21#_M1075_g N_A_630_367#_c_2130_n 6.66834e-19 $X=19.58 $Y=2.155
+ $X2=0 $Y2=0
cc_1023 N_A_1909_21#_M1078_g N_A_630_367#_c_2130_n 0.0127479f $X=20.01 $Y=2.155
+ $X2=0 $Y2=0
cc_1024 N_A_1909_21#_M1088_g N_A_630_367#_c_2130_n 0.0131924f $X=20.44 $Y=2.155
+ $X2=0 $Y2=0
cc_1025 N_A_1909_21#_M1006_g N_A_630_367#_c_1951_n 8.63014e-19 $X=13.13 $Y=2.155
+ $X2=0 $Y2=0
cc_1026 N_A_1909_21#_M1008_g N_A_630_367#_c_1951_n 8.63014e-19 $X=13.56 $Y=2.155
+ $X2=0 $Y2=0
cc_1027 N_A_1909_21#_M1013_g N_A_630_367#_c_1952_n 8.63014e-19 $X=13.99 $Y=2.155
+ $X2=0 $Y2=0
cc_1028 N_A_1909_21#_M1023_g N_A_630_367#_c_1952_n 8.63014e-19 $X=14.42 $Y=2.155
+ $X2=0 $Y2=0
cc_1029 N_A_1909_21#_M1025_g N_A_630_367#_c_1953_n 8.63014e-19 $X=14.85 $Y=2.155
+ $X2=0 $Y2=0
cc_1030 N_A_1909_21#_M1026_g N_A_630_367#_c_1953_n 8.63014e-19 $X=15.28 $Y=2.155
+ $X2=0 $Y2=0
cc_1031 N_A_1909_21#_M1030_g N_A_630_367#_c_1954_n 8.63014e-19 $X=15.71 $Y=2.155
+ $X2=0 $Y2=0
cc_1032 N_A_1909_21#_M1032_g N_A_630_367#_c_1954_n 8.63014e-19 $X=16.14 $Y=2.155
+ $X2=0 $Y2=0
cc_1033 N_A_1909_21#_M1038_g N_A_630_367#_c_1955_n 8.63014e-19 $X=16.57 $Y=2.155
+ $X2=0 $Y2=0
cc_1034 N_A_1909_21#_M1042_g N_A_630_367#_c_1955_n 8.63014e-19 $X=17 $Y=2.155
+ $X2=0 $Y2=0
cc_1035 N_A_1909_21#_M1046_g N_A_630_367#_c_1956_n 8.63014e-19 $X=17.43 $Y=2.155
+ $X2=0 $Y2=0
cc_1036 N_A_1909_21#_M1050_g N_A_630_367#_c_1956_n 8.63014e-19 $X=17.86 $Y=2.155
+ $X2=0 $Y2=0
cc_1037 N_A_1909_21#_M1056_g N_A_630_367#_c_1957_n 8.63014e-19 $X=18.29 $Y=2.155
+ $X2=0 $Y2=0
cc_1038 N_A_1909_21#_M1062_g N_A_630_367#_c_1957_n 8.63014e-19 $X=18.72 $Y=2.155
+ $X2=0 $Y2=0
cc_1039 N_A_1909_21#_M1063_g N_A_630_367#_c_1958_n 8.63014e-19 $X=19.15 $Y=2.155
+ $X2=0 $Y2=0
cc_1040 N_A_1909_21#_M1075_g N_A_630_367#_c_1958_n 8.63014e-19 $X=19.58 $Y=2.155
+ $X2=0 $Y2=0
cc_1041 N_A_1909_21#_c_1033_n N_Z_c_2279_n 0.00137326f $X=9.62 $Y=0.985 $X2=0
+ $Y2=0
cc_1042 N_A_1909_21#_c_1034_n N_Z_c_2279_n 0.00703917f $X=10.055 $Y=1.06 $X2=0
+ $Y2=0
cc_1043 N_A_1909_21#_c_1036_n N_Z_c_2279_n 0.0122752f $X=10.13 $Y=0.985 $X2=0
+ $Y2=0
cc_1044 N_A_1909_21#_c_1037_n N_Z_c_2279_n 0.00475429f $X=10.565 $Y=1.06 $X2=0
+ $Y2=0
cc_1045 N_A_1909_21#_c_1038_n N_Z_c_2279_n 0.0157102f $X=10.64 $Y=0.985 $X2=0
+ $Y2=0
cc_1046 N_A_1909_21#_c_1039_n N_Z_c_2279_n 0.00475386f $X=11.075 $Y=1.06 $X2=0
+ $Y2=0
cc_1047 N_A_1909_21#_c_1040_n N_Z_c_2279_n 0.0117416f $X=11.15 $Y=0.985 $X2=0
+ $Y2=0
cc_1048 N_A_1909_21#_c_1046_n N_Z_c_2280_n 0.0113651f $X=12.44 $Y=0.985 $X2=0
+ $Y2=0
cc_1049 N_A_1909_21#_c_1048_n N_Z_c_2280_n 0.01086f $X=12.87 $Y=0.985 $X2=0
+ $Y2=0
cc_1050 N_A_1909_21#_c_1050_n N_Z_c_2280_n 0.01086f $X=13.3 $Y=0.985 $X2=0 $Y2=0
cc_1051 N_A_1909_21#_c_1052_n N_Z_c_2280_n 0.01086f $X=13.73 $Y=0.985 $X2=0
+ $Y2=0
cc_1052 N_A_1909_21#_c_1054_n N_Z_c_2280_n 0.01086f $X=14.16 $Y=0.985 $X2=0
+ $Y2=0
cc_1053 N_A_1909_21#_c_1056_n N_Z_c_2280_n 0.01086f $X=14.59 $Y=0.985 $X2=0
+ $Y2=0
cc_1054 N_A_1909_21#_c_1058_n N_Z_c_2280_n 0.01086f $X=15.02 $Y=0.985 $X2=0
+ $Y2=0
cc_1055 N_A_1909_21#_c_1060_n N_Z_c_2280_n 0.0068359f $X=15.45 $Y=0.985 $X2=0
+ $Y2=0
cc_1056 N_A_1909_21#_c_1077_n N_Z_c_2280_n 0.21355f $X=15.33 $Y=1.2 $X2=0 $Y2=0
cc_1057 N_A_1909_21#_c_1082_n N_Z_c_2280_n 0.0217737f $X=20.515 $Y=1.15 $X2=0
+ $Y2=0
cc_1058 N_A_1909_21#_M1000_g N_Z_c_2283_n 0.0104764f $X=12.27 $Y=2.155 $X2=0
+ $Y2=0
cc_1059 N_A_1909_21#_M1002_g N_Z_c_2283_n 0.0156244f $X=12.7 $Y=2.155 $X2=0
+ $Y2=0
cc_1060 N_A_1909_21#_c_1077_n N_Z_c_2283_n 0.0297512f $X=15.33 $Y=1.2 $X2=0
+ $Y2=0
cc_1061 N_A_1909_21#_c_1082_n N_Z_c_2283_n 0.00264397f $X=20.515 $Y=1.15 $X2=0
+ $Y2=0
cc_1062 N_A_1909_21#_M1006_g N_Z_c_2284_n 0.0140452f $X=13.13 $Y=2.155 $X2=0
+ $Y2=0
cc_1063 N_A_1909_21#_M1008_g N_Z_c_2284_n 0.0140452f $X=13.56 $Y=2.155 $X2=0
+ $Y2=0
cc_1064 N_A_1909_21#_c_1077_n N_Z_c_2284_n 0.046956f $X=15.33 $Y=1.2 $X2=0 $Y2=0
cc_1065 N_A_1909_21#_c_1082_n N_Z_c_2284_n 0.0026313f $X=20.515 $Y=1.15 $X2=0
+ $Y2=0
cc_1066 N_A_1909_21#_M1013_g N_Z_c_2285_n 0.0140452f $X=13.99 $Y=2.155 $X2=0
+ $Y2=0
cc_1067 N_A_1909_21#_M1023_g N_Z_c_2285_n 0.0140452f $X=14.42 $Y=2.155 $X2=0
+ $Y2=0
cc_1068 N_A_1909_21#_c_1077_n N_Z_c_2285_n 0.046956f $X=15.33 $Y=1.2 $X2=0 $Y2=0
cc_1069 N_A_1909_21#_c_1082_n N_Z_c_2285_n 0.0026313f $X=20.515 $Y=1.15 $X2=0
+ $Y2=0
cc_1070 N_A_1909_21#_M1025_g N_Z_c_2286_n 0.0140452f $X=14.85 $Y=2.155 $X2=0
+ $Y2=0
cc_1071 N_A_1909_21#_M1026_g N_Z_c_2286_n 0.0140442f $X=15.28 $Y=2.155 $X2=0
+ $Y2=0
cc_1072 N_A_1909_21#_c_1077_n N_Z_c_2286_n 0.0469456f $X=15.33 $Y=1.2 $X2=0
+ $Y2=0
cc_1073 N_A_1909_21#_c_1082_n N_Z_c_2286_n 0.0026313f $X=20.515 $Y=1.15 $X2=0
+ $Y2=0
cc_1074 N_A_1909_21#_M1030_g N_Z_c_2287_n 0.0141004f $X=15.71 $Y=2.155 $X2=0
+ $Y2=0
cc_1075 N_A_1909_21#_M1032_g N_Z_c_2287_n 0.0141065f $X=16.14 $Y=2.155 $X2=0
+ $Y2=0
cc_1076 N_A_1909_21#_c_1077_n N_Z_c_2287_n 0.0159049f $X=15.33 $Y=1.2 $X2=0
+ $Y2=0
cc_1077 N_A_1909_21#_c_1078_n N_Z_c_2287_n 0.0300159f $X=21.48 $Y=1.15 $X2=0
+ $Y2=0
cc_1078 N_A_1909_21#_c_1082_n N_Z_c_2287_n 0.00226747f $X=20.515 $Y=1.15 $X2=0
+ $Y2=0
cc_1079 N_A_1909_21#_M1038_g N_Z_c_2288_n 0.0144336f $X=16.57 $Y=2.155 $X2=0
+ $Y2=0
cc_1080 N_A_1909_21#_M1042_g N_Z_c_2288_n 0.014457f $X=17 $Y=2.155 $X2=0 $Y2=0
cc_1081 N_A_1909_21#_c_1078_n N_Z_c_2288_n 0.0481189f $X=21.48 $Y=1.15 $X2=0
+ $Y2=0
cc_1082 N_A_1909_21#_c_1082_n N_Z_c_2288_n 0.00228443f $X=20.515 $Y=1.15 $X2=0
+ $Y2=0
cc_1083 N_A_1909_21#_M1046_g N_Z_c_2289_n 0.0144595f $X=17.43 $Y=2.155 $X2=0
+ $Y2=0
cc_1084 N_A_1909_21#_M1050_g N_Z_c_2289_n 0.0144595f $X=17.86 $Y=2.155 $X2=0
+ $Y2=0
cc_1085 N_A_1909_21#_c_1078_n N_Z_c_2289_n 0.0481189f $X=21.48 $Y=1.15 $X2=0
+ $Y2=0
cc_1086 N_A_1909_21#_c_1082_n N_Z_c_2289_n 0.00228443f $X=20.515 $Y=1.15 $X2=0
+ $Y2=0
cc_1087 N_A_1909_21#_M1056_g N_Z_c_2290_n 0.0144595f $X=18.29 $Y=2.155 $X2=0
+ $Y2=0
cc_1088 N_A_1909_21#_M1062_g N_Z_c_2290_n 0.0144595f $X=18.72 $Y=2.155 $X2=0
+ $Y2=0
cc_1089 N_A_1909_21#_c_1078_n N_Z_c_2290_n 0.0481189f $X=21.48 $Y=1.15 $X2=0
+ $Y2=0
cc_1090 N_A_1909_21#_c_1082_n N_Z_c_2290_n 0.00228443f $X=20.515 $Y=1.15 $X2=0
+ $Y2=0
cc_1091 N_A_1909_21#_M1063_g N_Z_c_2291_n 0.0144595f $X=19.15 $Y=2.155 $X2=0
+ $Y2=0
cc_1092 N_A_1909_21#_M1075_g N_Z_c_2291_n 0.0144595f $X=19.58 $Y=2.155 $X2=0
+ $Y2=0
cc_1093 N_A_1909_21#_c_1078_n N_Z_c_2291_n 0.048119f $X=21.48 $Y=1.15 $X2=0
+ $Y2=0
cc_1094 N_A_1909_21#_c_1082_n N_Z_c_2291_n 0.00224401f $X=20.515 $Y=1.15 $X2=0
+ $Y2=0
cc_1095 N_A_1909_21#_M1078_g N_Z_c_2292_n 0.0144595f $X=20.01 $Y=2.155 $X2=0
+ $Y2=0
cc_1096 N_A_1909_21#_M1088_g N_Z_c_2292_n 0.0146907f $X=20.44 $Y=2.155 $X2=0
+ $Y2=0
cc_1097 N_A_1909_21#_c_1078_n N_Z_c_2292_n 0.0488193f $X=21.48 $Y=1.15 $X2=0
+ $Y2=0
cc_1098 N_A_1909_21#_c_1079_n N_Z_c_2292_n 0.00121177f $X=21.265 $Y=1.15 $X2=0
+ $Y2=0
cc_1099 N_A_1909_21#_c_1082_n N_Z_c_2292_n 0.00224401f $X=20.515 $Y=1.15 $X2=0
+ $Y2=0
cc_1100 N_A_1909_21#_c_1078_n N_Z_c_2293_n 0.0201951f $X=21.48 $Y=1.15 $X2=0
+ $Y2=0
cc_1101 N_A_1909_21#_c_1079_n N_Z_c_2293_n 0.00579521f $X=21.265 $Y=1.15 $X2=0
+ $Y2=0
cc_1102 N_A_1909_21#_c_1080_n N_Z_c_2293_n 0.00600164f $X=21.565 $Y=1.695 $X2=0
+ $Y2=0
cc_1103 N_A_1909_21#_c_1119_p N_Z_c_2293_n 9.33846e-19 $X=21.645 $Y=1.78 $X2=0
+ $Y2=0
cc_1104 N_A_1909_21#_M1088_g N_Z_c_2294_n 0.00408335f $X=20.44 $Y=2.155 $X2=0
+ $Y2=0
cc_1105 N_A_1909_21#_c_1119_p N_Z_c_2294_n 0.0025951f $X=21.645 $Y=1.78 $X2=0
+ $Y2=0
cc_1106 N_A_1909_21#_c_1077_n N_Z_c_2295_n 0.0150652f $X=15.33 $Y=1.2 $X2=0
+ $Y2=0
cc_1107 N_A_1909_21#_c_1082_n N_Z_c_2295_n 0.00270827f $X=20.515 $Y=1.15 $X2=0
+ $Y2=0
cc_1108 N_A_1909_21#_c_1077_n N_Z_c_2296_n 0.0150652f $X=15.33 $Y=1.2 $X2=0
+ $Y2=0
cc_1109 N_A_1909_21#_c_1082_n N_Z_c_2296_n 0.00270827f $X=20.515 $Y=1.15 $X2=0
+ $Y2=0
cc_1110 N_A_1909_21#_c_1077_n N_Z_c_2297_n 0.0150652f $X=15.33 $Y=1.2 $X2=0
+ $Y2=0
cc_1111 N_A_1909_21#_c_1082_n N_Z_c_2297_n 0.00270827f $X=20.515 $Y=1.15 $X2=0
+ $Y2=0
cc_1112 N_A_1909_21#_c_1077_n N_Z_c_2298_n 0.0146792f $X=15.33 $Y=1.2 $X2=0
+ $Y2=0
cc_1113 N_A_1909_21#_c_1082_n N_Z_c_2298_n 0.00245286f $X=20.515 $Y=1.15 $X2=0
+ $Y2=0
cc_1114 N_A_1909_21#_M1032_g N_Z_c_2299_n 3.16435e-19 $X=16.14 $Y=2.155 $X2=0
+ $Y2=0
cc_1115 N_A_1909_21#_c_1078_n N_Z_c_2299_n 0.0153179f $X=21.48 $Y=1.15 $X2=0
+ $Y2=0
cc_1116 N_A_1909_21#_c_1082_n N_Z_c_2299_n 0.00235998f $X=20.515 $Y=1.15 $X2=0
+ $Y2=0
cc_1117 N_A_1909_21#_c_1078_n N_Z_c_2300_n 0.01535f $X=21.48 $Y=1.15 $X2=0 $Y2=0
cc_1118 N_A_1909_21#_c_1082_n N_Z_c_2300_n 0.00235998f $X=20.515 $Y=1.15 $X2=0
+ $Y2=0
cc_1119 N_A_1909_21#_c_1078_n N_Z_c_2301_n 0.01535f $X=21.48 $Y=1.15 $X2=0 $Y2=0
cc_1120 N_A_1909_21#_c_1082_n N_Z_c_2301_n 0.00235998f $X=20.515 $Y=1.15 $X2=0
+ $Y2=0
cc_1121 N_A_1909_21#_c_1078_n N_Z_c_2302_n 0.0153501f $X=21.48 $Y=1.15 $X2=0
+ $Y2=0
cc_1122 N_A_1909_21#_c_1082_n N_Z_c_2302_n 0.00231808f $X=20.515 $Y=1.15 $X2=0
+ $Y2=0
cc_1123 N_A_1909_21#_c_1078_n N_Z_c_2303_n 0.0153501f $X=21.48 $Y=1.15 $X2=0
+ $Y2=0
cc_1124 N_A_1909_21#_c_1082_n N_Z_c_2303_n 0.00231808f $X=20.515 $Y=1.15 $X2=0
+ $Y2=0
cc_1125 N_A_1909_21#_c_1042_n Z 0.00885835f $X=11.58 $Y=0.985 $X2=0 $Y2=0
cc_1126 N_A_1909_21#_c_1044_n Z 0.00885835f $X=12.01 $Y=0.985 $X2=0 $Y2=0
cc_1127 N_A_1909_21#_M1000_g N_Z_c_2281_n 0.00203693f $X=12.27 $Y=2.155 $X2=0
+ $Y2=0
cc_1128 N_A_1909_21#_c_1040_n Z 0.00272799f $X=11.15 $Y=0.985 $X2=0 $Y2=0
cc_1129 N_A_1909_21#_c_1041_n Z 0.0170718f $X=11.505 $Y=1.06 $X2=0 $Y2=0
cc_1130 N_A_1909_21#_c_1042_n Z 0.00302133f $X=11.58 $Y=0.985 $X2=0 $Y2=0
cc_1131 N_A_1909_21#_c_1043_n Z 0.0125397f $X=11.935 $Y=1.06 $X2=0 $Y2=0
cc_1132 N_A_1909_21#_c_1044_n Z 0.0029206f $X=12.01 $Y=0.985 $X2=0 $Y2=0
cc_1133 N_A_1909_21#_M1000_g Z 0.00800649f $X=12.27 $Y=2.155 $X2=0 $Y2=0
cc_1134 N_A_1909_21#_c_1046_n Z 0.0025678f $X=12.44 $Y=0.985 $X2=0 $Y2=0
cc_1135 N_A_1909_21#_M1002_g Z 8.85336e-19 $X=12.7 $Y=2.155 $X2=0 $Y2=0
cc_1136 N_A_1909_21#_c_1076_n Z 0.00564825f $X=11.58 $Y=1.06 $X2=0 $Y2=0
cc_1137 N_A_1909_21#_c_1077_n Z 0.0213392f $X=15.33 $Y=1.2 $X2=0 $Y2=0
cc_1138 N_A_1909_21#_c_1082_n Z 0.0255682f $X=20.515 $Y=1.15 $X2=0 $Y2=0
cc_1139 N_A_1909_21#_c_1121_p N_VGND_M1028_s 0.00327924f $X=22.03 $Y=0.915 $X2=0
+ $Y2=0
cc_1140 N_A_1909_21#_c_1081_n N_VGND_M1028_s 0.00280575f $X=21.565 $Y=1.072
+ $X2=0 $Y2=0
cc_1141 N_A_1909_21#_c_1140_p N_VGND_M1029_s 0.00719624f $X=23.05 $Y=0.915 $X2=0
+ $Y2=0
cc_1142 N_A_1909_21#_c_1121_p N_VGND_c_2490_n 0.0106432f $X=22.03 $Y=0.915 $X2=0
+ $Y2=0
cc_1143 N_A_1909_21#_c_1081_n N_VGND_c_2490_n 0.0108778f $X=21.565 $Y=1.072
+ $X2=0 $Y2=0
cc_1144 N_A_1909_21#_c_1140_p N_VGND_c_2491_n 0.0247309f $X=23.05 $Y=0.915 $X2=0
+ $Y2=0
cc_1145 N_A_1909_21#_c_1033_n N_VGND_c_2507_n 0.0035993f $X=9.62 $Y=0.985 $X2=0
+ $Y2=0
cc_1146 N_A_1909_21#_c_1036_n N_VGND_c_2507_n 0.00359964f $X=10.13 $Y=0.985
+ $X2=0 $Y2=0
cc_1147 N_A_1909_21#_c_1038_n N_VGND_c_2507_n 0.00359964f $X=10.64 $Y=0.985
+ $X2=0 $Y2=0
cc_1148 N_A_1909_21#_c_1040_n N_VGND_c_2507_n 0.00359964f $X=11.15 $Y=0.985
+ $X2=0 $Y2=0
cc_1149 N_A_1909_21#_c_1042_n N_VGND_c_2507_n 0.00359964f $X=11.58 $Y=0.985
+ $X2=0 $Y2=0
cc_1150 N_A_1909_21#_c_1044_n N_VGND_c_2507_n 0.00359964f $X=12.01 $Y=0.985
+ $X2=0 $Y2=0
cc_1151 N_A_1909_21#_c_1046_n N_VGND_c_2507_n 0.00359964f $X=12.44 $Y=0.985
+ $X2=0 $Y2=0
cc_1152 N_A_1909_21#_c_1048_n N_VGND_c_2507_n 0.00359964f $X=12.87 $Y=0.985
+ $X2=0 $Y2=0
cc_1153 N_A_1909_21#_c_1050_n N_VGND_c_2507_n 0.00359964f $X=13.3 $Y=0.985 $X2=0
+ $Y2=0
cc_1154 N_A_1909_21#_c_1052_n N_VGND_c_2507_n 0.00359964f $X=13.73 $Y=0.985
+ $X2=0 $Y2=0
cc_1155 N_A_1909_21#_c_1054_n N_VGND_c_2507_n 0.00359964f $X=14.16 $Y=0.985
+ $X2=0 $Y2=0
cc_1156 N_A_1909_21#_c_1056_n N_VGND_c_2507_n 0.00359964f $X=14.59 $Y=0.985
+ $X2=0 $Y2=0
cc_1157 N_A_1909_21#_c_1058_n N_VGND_c_2507_n 0.00359964f $X=15.02 $Y=0.985
+ $X2=0 $Y2=0
cc_1158 N_A_1909_21#_c_1060_n N_VGND_c_2507_n 0.00359964f $X=15.45 $Y=0.985
+ $X2=0 $Y2=0
cc_1159 N_A_1909_21#_c_1139_p N_VGND_c_2509_n 0.0165835f $X=22.195 $Y=0.38 $X2=0
+ $Y2=0
cc_1160 N_A_1909_21#_c_1141_p N_VGND_c_2513_n 0.0177952f $X=23.215 $Y=0.43 $X2=0
+ $Y2=0
cc_1161 N_A_1909_21#_M1028_d N_VGND_c_2515_n 0.00318548f $X=21.98 $Y=0.235 $X2=0
+ $Y2=0
cc_1162 N_A_1909_21#_M1082_d N_VGND_c_2515_n 0.00223819f $X=23.075 $Y=0.235
+ $X2=0 $Y2=0
cc_1163 N_A_1909_21#_c_1033_n N_VGND_c_2515_n 0.00565951f $X=9.62 $Y=0.985 $X2=0
+ $Y2=0
cc_1164 N_A_1909_21#_c_1036_n N_VGND_c_2515_n 0.00584091f $X=10.13 $Y=0.985
+ $X2=0 $Y2=0
cc_1165 N_A_1909_21#_c_1038_n N_VGND_c_2515_n 0.00575526f $X=10.64 $Y=0.985
+ $X2=0 $Y2=0
cc_1166 N_A_1909_21#_c_1040_n N_VGND_c_2515_n 0.00556152f $X=11.15 $Y=0.985
+ $X2=0 $Y2=0
cc_1167 N_A_1909_21#_c_1042_n N_VGND_c_2515_n 0.00535287f $X=11.58 $Y=0.985
+ $X2=0 $Y2=0
cc_1168 N_A_1909_21#_c_1044_n N_VGND_c_2515_n 0.00535287f $X=12.01 $Y=0.985
+ $X2=0 $Y2=0
cc_1169 N_A_1909_21#_c_1046_n N_VGND_c_2515_n 0.00535287f $X=12.44 $Y=0.985
+ $X2=0 $Y2=0
cc_1170 N_A_1909_21#_c_1048_n N_VGND_c_2515_n 0.00535287f $X=12.87 $Y=0.985
+ $X2=0 $Y2=0
cc_1171 N_A_1909_21#_c_1050_n N_VGND_c_2515_n 0.00535287f $X=13.3 $Y=0.985 $X2=0
+ $Y2=0
cc_1172 N_A_1909_21#_c_1052_n N_VGND_c_2515_n 0.00535287f $X=13.73 $Y=0.985
+ $X2=0 $Y2=0
cc_1173 N_A_1909_21#_c_1054_n N_VGND_c_2515_n 0.00535287f $X=14.16 $Y=0.985
+ $X2=0 $Y2=0
cc_1174 N_A_1909_21#_c_1056_n N_VGND_c_2515_n 0.00535287f $X=14.59 $Y=0.985
+ $X2=0 $Y2=0
cc_1175 N_A_1909_21#_c_1058_n N_VGND_c_2515_n 0.00535287f $X=15.02 $Y=0.985
+ $X2=0 $Y2=0
cc_1176 N_A_1909_21#_c_1060_n N_VGND_c_2515_n 0.00682329f $X=15.45 $Y=0.985
+ $X2=0 $Y2=0
cc_1177 N_A_1909_21#_c_1121_p N_VGND_c_2515_n 0.00600857f $X=22.03 $Y=0.915
+ $X2=0 $Y2=0
cc_1178 N_A_1909_21#_c_1139_p N_VGND_c_2515_n 0.0123283f $X=22.195 $Y=0.38 $X2=0
+ $Y2=0
cc_1179 N_A_1909_21#_c_1140_p N_VGND_c_2515_n 0.0118153f $X=23.05 $Y=0.915 $X2=0
+ $Y2=0
cc_1180 N_A_1909_21#_c_1141_p N_VGND_c_2515_n 0.0123247f $X=23.215 $Y=0.43 $X2=0
+ $Y2=0
cc_1181 N_A_1909_21#_c_1081_n N_VGND_c_2515_n 0.00212083f $X=21.565 $Y=1.072
+ $X2=0 $Y2=0
cc_1182 N_A_1909_21#_c_1035_n N_A_584_47#_c_2727_n 0.00932555f $X=9.695 $Y=1.06
+ $X2=0 $Y2=0
cc_1183 N_A_1909_21#_c_1033_n N_A_584_47#_c_2797_n 0.0101056f $X=9.62 $Y=0.985
+ $X2=0 $Y2=0
cc_1184 N_A_1909_21#_c_1035_n N_A_584_47#_c_2797_n 5.37409e-19 $X=9.695 $Y=1.06
+ $X2=0 $Y2=0
cc_1185 N_A_1909_21#_c_1036_n N_A_584_47#_c_2797_n 0.00107885f $X=10.13 $Y=0.985
+ $X2=0 $Y2=0
cc_1186 N_A_1909_21#_c_1033_n N_A_584_47#_c_2835_n 0.0120219f $X=9.62 $Y=0.985
+ $X2=0 $Y2=0
cc_1187 N_A_1909_21#_c_1036_n N_A_584_47#_c_2835_n 0.0124373f $X=10.13 $Y=0.985
+ $X2=0 $Y2=0
cc_1188 N_A_1909_21#_c_1038_n N_A_584_47#_c_2835_n 0.00936123f $X=10.64 $Y=0.985
+ $X2=0 $Y2=0
cc_1189 N_A_1909_21#_c_1040_n N_A_584_47#_c_2835_n 0.00936123f $X=11.15 $Y=0.985
+ $X2=0 $Y2=0
cc_1190 N_A_1909_21#_c_1041_n N_A_584_47#_c_2835_n 3.5085e-19 $X=11.505 $Y=1.06
+ $X2=0 $Y2=0
cc_1191 N_A_1909_21#_c_1042_n N_A_584_47#_c_2835_n 0.00880578f $X=11.58 $Y=0.985
+ $X2=0 $Y2=0
cc_1192 N_A_1909_21#_c_1043_n N_A_584_47#_c_2835_n 3.5085e-19 $X=11.935 $Y=1.06
+ $X2=0 $Y2=0
cc_1193 N_A_1909_21#_c_1044_n N_A_584_47#_c_2835_n 0.00880578f $X=12.01 $Y=0.985
+ $X2=0 $Y2=0
cc_1194 N_A_1909_21#_c_1046_n N_A_584_47#_c_2835_n 0.00881197f $X=12.44 $Y=0.985
+ $X2=0 $Y2=0
cc_1195 N_A_1909_21#_c_1048_n N_A_584_47#_c_2835_n 0.00881197f $X=12.87 $Y=0.985
+ $X2=0 $Y2=0
cc_1196 N_A_1909_21#_c_1050_n N_A_584_47#_c_2835_n 0.00881197f $X=13.3 $Y=0.985
+ $X2=0 $Y2=0
cc_1197 N_A_1909_21#_c_1052_n N_A_584_47#_c_2835_n 0.00881197f $X=13.73 $Y=0.985
+ $X2=0 $Y2=0
cc_1198 N_A_1909_21#_c_1054_n N_A_584_47#_c_2835_n 0.00881197f $X=14.16 $Y=0.985
+ $X2=0 $Y2=0
cc_1199 N_A_1909_21#_c_1056_n N_A_584_47#_c_2835_n 0.00881197f $X=14.59 $Y=0.985
+ $X2=0 $Y2=0
cc_1200 N_A_1909_21#_c_1058_n N_A_584_47#_c_2835_n 0.00875432f $X=15.02 $Y=0.985
+ $X2=0 $Y2=0
cc_1201 N_A_1909_21#_c_1060_n N_A_584_47#_c_2835_n 0.0137217f $X=15.45 $Y=0.985
+ $X2=0 $Y2=0
cc_1202 N_A_1909_21#_c_1077_n N_A_584_47#_c_2835_n 0.00382187f $X=15.33 $Y=1.2
+ $X2=0 $Y2=0
cc_1203 N_A_1909_21#_c_1033_n N_A_584_47#_c_2800_n 0.00211143f $X=9.62 $Y=0.985
+ $X2=0 $Y2=0
cc_1204 N_A_1909_21#_c_1077_n N_A_584_47#_c_2730_n 0.0172313f $X=15.33 $Y=1.2
+ $X2=0 $Y2=0
cc_1205 N_A_1909_21#_c_1078_n N_A_584_47#_c_2730_n 0.00651109f $X=21.48 $Y=1.15
+ $X2=0 $Y2=0
cc_1206 N_A_1909_21#_c_1082_n N_A_584_47#_c_2730_n 0.00560097f $X=20.515 $Y=1.15
+ $X2=0 $Y2=0
cc_1207 N_A_M1009_g N_VPWR_c_1630_n 0.00858283f $X=21.43 $Y=2.465 $X2=0 $Y2=0
cc_1208 N_A_M1014_g N_VPWR_c_1631_n 0.00368607f $X=21.86 $Y=2.465 $X2=0 $Y2=0
cc_1209 N_A_M1034_g N_VPWR_c_1631_n 0.00368607f $X=22.29 $Y=2.465 $X2=0 $Y2=0
cc_1210 N_A_M1052_g N_VPWR_c_1632_n 0.00271808f $X=22.72 $Y=2.465 $X2=0 $Y2=0
cc_1211 N_A_M1072_g N_VPWR_c_1632_n 0.00271808f $X=23.15 $Y=2.465 $X2=0 $Y2=0
cc_1212 N_A_M1072_g N_VPWR_c_1633_n 0.00549284f $X=23.15 $Y=2.465 $X2=0 $Y2=0
cc_1213 N_A_M1076_g N_VPWR_c_1633_n 0.00549284f $X=23.58 $Y=2.465 $X2=0 $Y2=0
cc_1214 N_A_M1076_g N_VPWR_c_1634_n 0.0027547f $X=23.58 $Y=2.465 $X2=0 $Y2=0
cc_1215 N_A_M1079_g N_VPWR_c_1634_n 0.00628394f $X=24.035 $Y=2.465 $X2=0 $Y2=0
cc_1216 N_A_M1085_g N_VPWR_c_1636_n 0.00858283f $X=24.465 $Y=2.465 $X2=0 $Y2=0
cc_1217 A N_VPWR_c_1636_n 0.0142489f $X=24.635 $Y=1.21 $X2=0 $Y2=0
cc_1218 N_A_M1009_g N_VPWR_c_1661_n 0.00549284f $X=21.43 $Y=2.465 $X2=0 $Y2=0
cc_1219 N_A_M1014_g N_VPWR_c_1661_n 0.00549284f $X=21.86 $Y=2.465 $X2=0 $Y2=0
cc_1220 N_A_M1034_g N_VPWR_c_1663_n 0.00549284f $X=22.29 $Y=2.465 $X2=0 $Y2=0
cc_1221 N_A_M1052_g N_VPWR_c_1663_n 0.00549284f $X=22.72 $Y=2.465 $X2=0 $Y2=0
cc_1222 N_A_M1079_g N_VPWR_c_1665_n 0.00549284f $X=24.035 $Y=2.465 $X2=0 $Y2=0
cc_1223 N_A_M1085_g N_VPWR_c_1665_n 0.00549284f $X=24.465 $Y=2.465 $X2=0 $Y2=0
cc_1224 N_A_M1009_g N_VPWR_c_1612_n 0.0110929f $X=21.43 $Y=2.465 $X2=0 $Y2=0
cc_1225 N_A_M1014_g N_VPWR_c_1612_n 0.00979325f $X=21.86 $Y=2.465 $X2=0 $Y2=0
cc_1226 N_A_M1034_g N_VPWR_c_1612_n 0.00979325f $X=22.29 $Y=2.465 $X2=0 $Y2=0
cc_1227 N_A_M1052_g N_VPWR_c_1612_n 0.00979325f $X=22.72 $Y=2.465 $X2=0 $Y2=0
cc_1228 N_A_M1072_g N_VPWR_c_1612_n 0.00979325f $X=23.15 $Y=2.465 $X2=0 $Y2=0
cc_1229 N_A_M1076_g N_VPWR_c_1612_n 0.00985703f $X=23.58 $Y=2.465 $X2=0 $Y2=0
cc_1230 N_A_M1079_g N_VPWR_c_1612_n 0.00992535f $X=24.035 $Y=2.465 $X2=0 $Y2=0
cc_1231 N_A_M1085_g N_VPWR_c_1612_n 0.0107443f $X=24.465 $Y=2.465 $X2=0 $Y2=0
cc_1232 N_A_c_1480_n N_Z_c_2293_n 0.00347253f $X=21.505 $Y=1.63 $X2=0 $Y2=0
cc_1233 N_A_M1009_g N_Z_c_2294_n 0.00301743f $X=21.43 $Y=2.465 $X2=0 $Y2=0
cc_1234 N_A_c_1481_n N_VGND_c_2490_n 0.0112564f $X=21.905 $Y=1.185 $X2=0 $Y2=0
cc_1235 N_A_c_1483_n N_VGND_c_2490_n 0.00118513f $X=22.41 $Y=1.185 $X2=0 $Y2=0
cc_1236 N_A_c_1483_n N_VGND_c_2491_n 0.00568946f $X=22.41 $Y=1.185 $X2=0 $Y2=0
cc_1237 N_A_c_1485_n N_VGND_c_2491_n 0.00568946f $X=23 $Y=1.185 $X2=0 $Y2=0
cc_1238 N_A_c_1487_n N_VGND_c_2492_n 0.0192091f $X=23.43 $Y=1.185 $X2=0 $Y2=0
cc_1239 A N_VGND_c_2492_n 0.0272938f $X=24.635 $Y=1.21 $X2=0 $Y2=0
cc_1240 N_A_c_1492_n N_VGND_c_2492_n 0.0025254f $X=24.375 $Y=1.35 $X2=0 $Y2=0
cc_1241 N_A_c_1481_n N_VGND_c_2509_n 0.00505556f $X=21.905 $Y=1.185 $X2=0 $Y2=0
cc_1242 N_A_c_1483_n N_VGND_c_2509_n 0.00550269f $X=22.41 $Y=1.185 $X2=0 $Y2=0
cc_1243 N_A_c_1485_n N_VGND_c_2513_n 0.00549284f $X=23 $Y=1.185 $X2=0 $Y2=0
cc_1244 N_A_c_1487_n N_VGND_c_2513_n 0.00549284f $X=23.43 $Y=1.185 $X2=0 $Y2=0
cc_1245 N_A_c_1481_n N_VGND_c_2515_n 0.00495475f $X=21.905 $Y=1.185 $X2=0 $Y2=0
cc_1246 N_A_c_1483_n N_VGND_c_2515_n 0.00669934f $X=22.41 $Y=1.185 $X2=0 $Y2=0
cc_1247 N_A_c_1485_n N_VGND_c_2515_n 0.00651517f $X=23 $Y=1.185 $X2=0 $Y2=0
cc_1248 N_A_c_1487_n N_VGND_c_2515_n 0.0113003f $X=23.43 $Y=1.185 $X2=0 $Y2=0
cc_1249 N_VPWR_c_1612_n N_A_630_367#_M1001_s 0.00297803f $X=24.72 $Y=3.33
+ $X2=-0.19 $Y2=-0.245
cc_1250 N_VPWR_c_1612_n N_A_630_367#_M1012_s 0.00297803f $X=24.72 $Y=3.33 $X2=0
+ $Y2=0
cc_1251 N_VPWR_c_1612_n N_A_630_367#_M1019_s 0.00297803f $X=24.72 $Y=3.33 $X2=0
+ $Y2=0
cc_1252 N_VPWR_c_1612_n N_A_630_367#_M1037_s 0.00297803f $X=24.72 $Y=3.33 $X2=0
+ $Y2=0
cc_1253 N_VPWR_c_1612_n N_A_630_367#_M1041_s 0.00297803f $X=24.72 $Y=3.33 $X2=0
+ $Y2=0
cc_1254 N_VPWR_c_1612_n N_A_630_367#_M1058_s 0.00297803f $X=24.72 $Y=3.33 $X2=0
+ $Y2=0
cc_1255 N_VPWR_c_1612_n N_A_630_367#_M1064_s 0.00297803f $X=24.72 $Y=3.33 $X2=0
+ $Y2=0
cc_1256 N_VPWR_c_1612_n N_A_630_367#_M1069_s 0.00297803f $X=24.72 $Y=3.33 $X2=0
+ $Y2=0
cc_1257 N_VPWR_c_1612_n N_A_630_367#_M1077_s 0.00223819f $X=24.72 $Y=3.33 $X2=0
+ $Y2=0
cc_1258 N_VPWR_c_1612_n N_A_630_367#_M1087_s 0.00415099f $X=24.72 $Y=3.33 $X2=0
+ $Y2=0
cc_1259 N_VPWR_M1005_d N_A_630_367#_c_1959_n 0.00325679f $X=3.58 $Y=1.835 $X2=0
+ $Y2=0
cc_1260 N_VPWR_c_1618_n N_A_630_367#_c_1959_n 0.0135055f $X=3.72 $Y=2.37 $X2=0
+ $Y2=0
cc_1261 N_VPWR_M1018_d N_A_630_367#_c_1963_n 0.00325679f $X=4.44 $Y=1.835 $X2=0
+ $Y2=0
cc_1262 N_VPWR_c_1620_n N_A_630_367#_c_1963_n 0.0135055f $X=4.58 $Y=2.37 $X2=0
+ $Y2=0
cc_1263 N_VPWR_M1022_d N_A_630_367#_c_1967_n 0.00325679f $X=5.3 $Y=1.835 $X2=0
+ $Y2=0
cc_1264 N_VPWR_c_1621_n N_A_630_367#_c_1967_n 0.0135055f $X=5.44 $Y=2.37 $X2=0
+ $Y2=0
cc_1265 N_VPWR_M1040_d N_A_630_367#_c_1971_n 0.00333197f $X=6.16 $Y=1.835 $X2=0
+ $Y2=0
cc_1266 N_VPWR_c_1622_n N_A_630_367#_c_1971_n 0.0135055f $X=6.3 $Y=2.37 $X2=0
+ $Y2=0
cc_1267 N_VPWR_M1055_d N_A_630_367#_c_1975_n 0.00333197f $X=7.02 $Y=1.835 $X2=0
+ $Y2=0
cc_1268 N_VPWR_c_1623_n N_A_630_367#_c_1975_n 0.0135055f $X=7.16 $Y=2.37 $X2=0
+ $Y2=0
cc_1269 N_VPWR_M1061_d N_A_630_367#_c_1979_n 0.00396171f $X=7.88 $Y=1.835 $X2=0
+ $Y2=0
cc_1270 N_VPWR_c_1624_n N_A_630_367#_c_1979_n 0.0144005f $X=8.02 $Y=2.37 $X2=0
+ $Y2=0
cc_1271 N_VPWR_M1065_d N_A_630_367#_c_1983_n 0.00333197f $X=8.76 $Y=1.835 $X2=0
+ $Y2=0
cc_1272 N_VPWR_c_1626_n N_A_630_367#_c_1983_n 0.0135055f $X=8.9 $Y=2.37 $X2=0
+ $Y2=0
cc_1273 N_VPWR_M1074_d N_A_630_367#_c_1987_n 0.00431837f $X=9.62 $Y=1.835 $X2=0
+ $Y2=0
cc_1274 N_VPWR_c_1627_n N_A_630_367#_c_1987_n 0.0135055f $X=9.76 $Y=2.37 $X2=0
+ $Y2=0
cc_1275 N_VPWR_c_1628_n N_A_630_367#_c_1991_n 0.00244279f $X=10.62 $Y=1.98 $X2=0
+ $Y2=0
cc_1276 N_VPWR_c_1655_n N_A_630_367#_c_1999_n 0.0177952f $X=10.535 $Y=3.33 $X2=0
+ $Y2=0
cc_1277 N_VPWR_c_1612_n N_A_630_367#_c_1999_n 0.0123247f $X=24.72 $Y=3.33 $X2=0
+ $Y2=0
cc_1278 N_VPWR_c_1628_n N_A_630_367#_c_1937_n 0.0129859f $X=10.62 $Y=1.98 $X2=0
+ $Y2=0
cc_1279 N_VPWR_c_1628_n N_A_630_367#_c_1939_n 0.00563274f $X=10.62 $Y=1.98 $X2=0
+ $Y2=0
cc_1280 N_VPWR_c_1657_n N_A_630_367#_c_2015_n 0.0144144f $X=11.315 $Y=3.33 $X2=0
+ $Y2=0
cc_1281 N_VPWR_c_1612_n N_A_630_367#_c_2015_n 0.00940713f $X=24.72 $Y=3.33 $X2=0
+ $Y2=0
cc_1282 N_VPWR_M1089_d N_A_630_367#_c_1940_n 0.00630433f $X=11.34 $Y=1.835 $X2=0
+ $Y2=0
cc_1283 N_VPWR_c_1629_n N_A_630_367#_c_1940_n 0.0214262f $X=11.48 $Y=2.53 $X2=0
+ $Y2=0
cc_1284 N_VPWR_c_1629_n N_A_630_367#_c_2074_n 0.014387f $X=11.48 $Y=2.53 $X2=0
+ $Y2=0
cc_1285 N_VPWR_c_1659_n N_A_630_367#_c_1941_n 0.0322076f $X=21.05 $Y=3.33 $X2=0
+ $Y2=0
cc_1286 N_VPWR_c_1612_n N_A_630_367#_c_1941_n 0.0198243f $X=24.72 $Y=3.33 $X2=0
+ $Y2=0
cc_1287 N_VPWR_c_1629_n N_A_630_367#_c_1942_n 0.00592055f $X=11.48 $Y=2.53 $X2=0
+ $Y2=0
cc_1288 N_VPWR_c_1659_n N_A_630_367#_c_1942_n 0.0222501f $X=21.05 $Y=3.33 $X2=0
+ $Y2=0
cc_1289 N_VPWR_c_1612_n N_A_630_367#_c_1942_n 0.0127687f $X=24.72 $Y=3.33 $X2=0
+ $Y2=0
cc_1290 N_VPWR_c_1659_n N_A_630_367#_c_1943_n 0.0322076f $X=21.05 $Y=3.33 $X2=0
+ $Y2=0
cc_1291 N_VPWR_c_1612_n N_A_630_367#_c_1943_n 0.0198243f $X=24.72 $Y=3.33 $X2=0
+ $Y2=0
cc_1292 N_VPWR_c_1659_n N_A_630_367#_c_1944_n 0.0322076f $X=21.05 $Y=3.33 $X2=0
+ $Y2=0
cc_1293 N_VPWR_c_1612_n N_A_630_367#_c_1944_n 0.0198243f $X=24.72 $Y=3.33 $X2=0
+ $Y2=0
cc_1294 N_VPWR_c_1659_n N_A_630_367#_c_1945_n 0.0322076f $X=21.05 $Y=3.33 $X2=0
+ $Y2=0
cc_1295 N_VPWR_c_1612_n N_A_630_367#_c_1945_n 0.0198243f $X=24.72 $Y=3.33 $X2=0
+ $Y2=0
cc_1296 N_VPWR_c_1659_n N_A_630_367#_c_1946_n 0.0322076f $X=21.05 $Y=3.33 $X2=0
+ $Y2=0
cc_1297 N_VPWR_c_1612_n N_A_630_367#_c_1946_n 0.0198243f $X=24.72 $Y=3.33 $X2=0
+ $Y2=0
cc_1298 N_VPWR_c_1659_n N_A_630_367#_c_1947_n 0.0322076f $X=21.05 $Y=3.33 $X2=0
+ $Y2=0
cc_1299 N_VPWR_c_1612_n N_A_630_367#_c_1947_n 0.0198243f $X=24.72 $Y=3.33 $X2=0
+ $Y2=0
cc_1300 N_VPWR_c_1659_n N_A_630_367#_c_1948_n 0.0322076f $X=21.05 $Y=3.33 $X2=0
+ $Y2=0
cc_1301 N_VPWR_c_1612_n N_A_630_367#_c_1948_n 0.0198243f $X=24.72 $Y=3.33 $X2=0
+ $Y2=0
cc_1302 N_VPWR_c_1659_n N_A_630_367#_c_1949_n 0.0322076f $X=21.05 $Y=3.33 $X2=0
+ $Y2=0
cc_1303 N_VPWR_c_1612_n N_A_630_367#_c_1949_n 0.0198243f $X=24.72 $Y=3.33 $X2=0
+ $Y2=0
cc_1304 N_VPWR_c_1630_n N_A_630_367#_c_1950_n 0.00590277f $X=21.215 $Y=1.98
+ $X2=0 $Y2=0
cc_1305 N_VPWR_c_1659_n N_A_630_367#_c_1950_n 0.0544577f $X=21.05 $Y=3.33 $X2=0
+ $Y2=0
cc_1306 N_VPWR_c_1612_n N_A_630_367#_c_1950_n 0.032593f $X=24.72 $Y=3.33 $X2=0
+ $Y2=0
cc_1307 N_VPWR_c_1630_n N_A_630_367#_c_2130_n 0.00219191f $X=21.215 $Y=1.98
+ $X2=0 $Y2=0
cc_1308 N_VPWR_c_1643_n N_A_630_367#_c_2017_n 0.00609757f $X=3.625 $Y=3.33 $X2=0
+ $Y2=0
cc_1309 N_VPWR_c_1612_n N_A_630_367#_c_2017_n 0.0102035f $X=24.72 $Y=3.33 $X2=0
+ $Y2=0
cc_1310 N_VPWR_c_1619_n N_A_630_367#_c_2022_n 0.00609757f $X=4.485 $Y=3.33 $X2=0
+ $Y2=0
cc_1311 N_VPWR_c_1612_n N_A_630_367#_c_2022_n 0.0102035f $X=24.72 $Y=3.33 $X2=0
+ $Y2=0
cc_1312 N_VPWR_c_1645_n N_A_630_367#_c_2028_n 0.00609757f $X=5.345 $Y=3.33 $X2=0
+ $Y2=0
cc_1313 N_VPWR_c_1612_n N_A_630_367#_c_2028_n 0.0102035f $X=24.72 $Y=3.33 $X2=0
+ $Y2=0
cc_1314 N_VPWR_c_1647_n N_A_630_367#_c_2034_n 0.00609757f $X=6.205 $Y=3.33 $X2=0
+ $Y2=0
cc_1315 N_VPWR_c_1612_n N_A_630_367#_c_2034_n 0.0102035f $X=24.72 $Y=3.33 $X2=0
+ $Y2=0
cc_1316 N_VPWR_c_1649_n N_A_630_367#_c_2040_n 0.00609757f $X=7.065 $Y=3.33 $X2=0
+ $Y2=0
cc_1317 N_VPWR_c_1612_n N_A_630_367#_c_2040_n 0.0102035f $X=24.72 $Y=3.33 $X2=0
+ $Y2=0
cc_1318 N_VPWR_c_1651_n N_A_630_367#_c_2046_n 0.00609757f $X=7.925 $Y=3.33 $X2=0
+ $Y2=0
cc_1319 N_VPWR_c_1612_n N_A_630_367#_c_2046_n 0.0102035f $X=24.72 $Y=3.33 $X2=0
+ $Y2=0
cc_1320 N_VPWR_c_1624_n N_A_630_367#_c_2052_n 0.03826f $X=8.02 $Y=2.37 $X2=0
+ $Y2=0
cc_1321 N_VPWR_c_1625_n N_A_630_367#_c_2052_n 0.00609757f $X=8.805 $Y=3.33 $X2=0
+ $Y2=0
cc_1322 N_VPWR_c_1612_n N_A_630_367#_c_2052_n 0.0102035f $X=24.72 $Y=3.33 $X2=0
+ $Y2=0
cc_1323 N_VPWR_c_1653_n N_A_630_367#_c_2058_n 0.00609757f $X=9.665 $Y=3.33 $X2=0
+ $Y2=0
cc_1324 N_VPWR_c_1612_n N_A_630_367#_c_2058_n 0.0102035f $X=24.72 $Y=3.33 $X2=0
+ $Y2=0
cc_1325 N_VPWR_c_1659_n N_A_630_367#_c_1951_n 0.0222501f $X=21.05 $Y=3.33 $X2=0
+ $Y2=0
cc_1326 N_VPWR_c_1612_n N_A_630_367#_c_1951_n 0.0127687f $X=24.72 $Y=3.33 $X2=0
+ $Y2=0
cc_1327 N_VPWR_c_1659_n N_A_630_367#_c_1952_n 0.0222501f $X=21.05 $Y=3.33 $X2=0
+ $Y2=0
cc_1328 N_VPWR_c_1612_n N_A_630_367#_c_1952_n 0.0127687f $X=24.72 $Y=3.33 $X2=0
+ $Y2=0
cc_1329 N_VPWR_c_1659_n N_A_630_367#_c_1953_n 0.0222501f $X=21.05 $Y=3.33 $X2=0
+ $Y2=0
cc_1330 N_VPWR_c_1612_n N_A_630_367#_c_1953_n 0.0127687f $X=24.72 $Y=3.33 $X2=0
+ $Y2=0
cc_1331 N_VPWR_c_1659_n N_A_630_367#_c_1954_n 0.0222501f $X=21.05 $Y=3.33 $X2=0
+ $Y2=0
cc_1332 N_VPWR_c_1612_n N_A_630_367#_c_1954_n 0.0127687f $X=24.72 $Y=3.33 $X2=0
+ $Y2=0
cc_1333 N_VPWR_c_1659_n N_A_630_367#_c_1955_n 0.0222501f $X=21.05 $Y=3.33 $X2=0
+ $Y2=0
cc_1334 N_VPWR_c_1612_n N_A_630_367#_c_1955_n 0.0127687f $X=24.72 $Y=3.33 $X2=0
+ $Y2=0
cc_1335 N_VPWR_c_1659_n N_A_630_367#_c_1956_n 0.0222501f $X=21.05 $Y=3.33 $X2=0
+ $Y2=0
cc_1336 N_VPWR_c_1612_n N_A_630_367#_c_1956_n 0.0127687f $X=24.72 $Y=3.33 $X2=0
+ $Y2=0
cc_1337 N_VPWR_c_1659_n N_A_630_367#_c_1957_n 0.0222501f $X=21.05 $Y=3.33 $X2=0
+ $Y2=0
cc_1338 N_VPWR_c_1612_n N_A_630_367#_c_1957_n 0.0127687f $X=24.72 $Y=3.33 $X2=0
+ $Y2=0
cc_1339 N_VPWR_c_1659_n N_A_630_367#_c_1958_n 0.0222501f $X=21.05 $Y=3.33 $X2=0
+ $Y2=0
cc_1340 N_VPWR_c_1612_n N_A_630_367#_c_1958_n 0.0127687f $X=24.72 $Y=3.33 $X2=0
+ $Y2=0
cc_1341 N_VPWR_c_1630_n N_Z_c_2294_n 0.0639967f $X=21.215 $Y=1.98 $X2=0 $Y2=0
cc_1342 N_VPWR_c_1659_n N_Z_c_2294_n 0.00643696f $X=21.05 $Y=3.33 $X2=0 $Y2=0
cc_1343 N_VPWR_c_1612_n N_Z_c_2294_n 0.00815161f $X=24.72 $Y=3.33 $X2=0 $Y2=0
cc_1344 N_A_630_367#_c_1940_n N_Z_M1000_d 0.0126241f $X=12.32 $Y=2.072 $X2=0
+ $Y2=0
cc_1345 N_A_630_367#_c_1937_n N_Z_c_2279_n 0.0260886f $X=10.885 $Y=1.55 $X2=0
+ $Y2=0
cc_1346 N_A_630_367#_c_1938_n N_Z_c_2279_n 0.0116838f $X=10.355 $Y=1.55 $X2=0
+ $Y2=0
cc_1347 N_A_630_367#_M1000_s N_Z_c_2283_n 0.00183453f $X=12.345 $Y=1.525 $X2=0
+ $Y2=0
cc_1348 N_A_630_367#_c_1940_n N_Z_c_2283_n 0.00576673f $X=12.32 $Y=2.072 $X2=0
+ $Y2=0
cc_1349 N_A_630_367#_c_2072_n N_Z_c_2283_n 0.0170548f $X=12.485 $Y=2.185 $X2=0
+ $Y2=0
cc_1350 N_A_630_367#_c_1941_n N_Z_c_2421_n 0.0138035f $X=13.18 $Y=2.975 $X2=0
+ $Y2=0
cc_1351 N_A_630_367#_M1006_s N_Z_c_2284_n 0.00177869f $X=13.205 $Y=1.525 $X2=0
+ $Y2=0
cc_1352 N_A_630_367#_c_2081_n N_Z_c_2284_n 0.0173823f $X=13.345 $Y=1.98 $X2=0
+ $Y2=0
cc_1353 N_A_630_367#_c_1943_n N_Z_c_2424_n 0.0138035f $X=14.04 $Y=2.975 $X2=0
+ $Y2=0
cc_1354 N_A_630_367#_M1013_s N_Z_c_2285_n 0.00177869f $X=14.065 $Y=1.525 $X2=0
+ $Y2=0
cc_1355 N_A_630_367#_c_2087_n N_Z_c_2285_n 0.0173823f $X=14.205 $Y=1.98 $X2=0
+ $Y2=0
cc_1356 N_A_630_367#_c_1944_n N_Z_c_2427_n 0.0138035f $X=14.9 $Y=2.975 $X2=0
+ $Y2=0
cc_1357 N_A_630_367#_M1025_s N_Z_c_2286_n 0.00177869f $X=14.925 $Y=1.525 $X2=0
+ $Y2=0
cc_1358 N_A_630_367#_c_2093_n N_Z_c_2286_n 0.0173823f $X=15.065 $Y=1.98 $X2=0
+ $Y2=0
cc_1359 N_A_630_367#_c_1945_n N_Z_c_2430_n 0.0138035f $X=15.76 $Y=2.975 $X2=0
+ $Y2=0
cc_1360 N_A_630_367#_M1030_s N_Z_c_2287_n 0.00177869f $X=15.785 $Y=1.525 $X2=0
+ $Y2=0
cc_1361 N_A_630_367#_c_2099_n N_Z_c_2287_n 0.0173823f $X=15.925 $Y=1.98 $X2=0
+ $Y2=0
cc_1362 N_A_630_367#_c_1946_n N_Z_c_2433_n 0.0138035f $X=16.62 $Y=2.975 $X2=0
+ $Y2=0
cc_1363 N_A_630_367#_M1038_s N_Z_c_2288_n 0.00178113f $X=16.645 $Y=1.525 $X2=0
+ $Y2=0
cc_1364 N_A_630_367#_c_2105_n N_Z_c_2288_n 0.017436f $X=16.785 $Y=1.98 $X2=0
+ $Y2=0
cc_1365 N_A_630_367#_c_1947_n N_Z_c_2436_n 0.0138035f $X=17.48 $Y=2.975 $X2=0
+ $Y2=0
cc_1366 N_A_630_367#_M1046_s N_Z_c_2289_n 0.00178113f $X=17.505 $Y=1.525 $X2=0
+ $Y2=0
cc_1367 N_A_630_367#_c_2111_n N_Z_c_2289_n 0.017436f $X=17.645 $Y=1.98 $X2=0
+ $Y2=0
cc_1368 N_A_630_367#_c_1948_n N_Z_c_2439_n 0.0138035f $X=18.34 $Y=2.975 $X2=0
+ $Y2=0
cc_1369 N_A_630_367#_M1056_s N_Z_c_2290_n 0.00178113f $X=18.365 $Y=1.525 $X2=0
+ $Y2=0
cc_1370 N_A_630_367#_c_2117_n N_Z_c_2290_n 0.017436f $X=18.505 $Y=1.98 $X2=0
+ $Y2=0
cc_1371 N_A_630_367#_c_1949_n N_Z_c_2442_n 0.0138035f $X=19.2 $Y=2.975 $X2=0
+ $Y2=0
cc_1372 N_A_630_367#_M1063_s N_Z_c_2291_n 0.00178113f $X=19.225 $Y=1.525 $X2=0
+ $Y2=0
cc_1373 N_A_630_367#_c_2123_n N_Z_c_2291_n 0.017436f $X=19.365 $Y=1.98 $X2=0
+ $Y2=0
cc_1374 N_A_630_367#_c_1950_n N_Z_c_2445_n 0.0138035f $X=20.06 $Y=2.975 $X2=0
+ $Y2=0
cc_1375 N_A_630_367#_M1078_s N_Z_c_2292_n 0.00178113f $X=20.085 $Y=1.525 $X2=0
+ $Y2=0
cc_1376 N_A_630_367#_c_2130_n N_Z_c_2292_n 0.017436f $X=20.225 $Y=1.98 $X2=0
+ $Y2=0
cc_1377 N_A_630_367#_c_2130_n N_Z_c_2294_n 0.0333436f $X=20.225 $Y=1.98 $X2=0
+ $Y2=0
cc_1378 N_A_630_367#_c_1937_n N_Z_c_2281_n 0.0116379f $X=10.885 $Y=1.55 $X2=0
+ $Y2=0
cc_1379 N_A_630_367#_c_1939_n N_Z_c_2281_n 0.0114848f $X=11.01 $Y=1.96 $X2=0
+ $Y2=0
cc_1380 N_A_630_367#_c_1940_n N_Z_c_2281_n 0.0682412f $X=12.32 $Y=2.072 $X2=0
+ $Y2=0
cc_1381 N_A_630_367#_c_1937_n Z 0.00368556f $X=10.885 $Y=1.55 $X2=0 $Y2=0
cc_1382 N_Z_M1017_s N_VGND_c_2515_n 0.00289884f $X=9.695 $Y=0.235 $X2=0 $Y2=0
cc_1383 N_Z_M1027_s N_VGND_c_2515_n 0.00289884f $X=10.715 $Y=0.235 $X2=0 $Y2=0
cc_1384 N_Z_M1033_s N_VGND_c_2515_n 0.00225465f $X=11.655 $Y=0.235 $X2=0 $Y2=0
cc_1385 N_Z_M1048_s N_VGND_c_2515_n 0.00225465f $X=12.515 $Y=0.235 $X2=0 $Y2=0
cc_1386 N_Z_M1059_s N_VGND_c_2515_n 0.00225465f $X=13.375 $Y=0.235 $X2=0 $Y2=0
cc_1387 N_Z_M1067_s N_VGND_c_2515_n 0.00225465f $X=14.235 $Y=0.235 $X2=0 $Y2=0
cc_1388 N_Z_M1081_s N_VGND_c_2515_n 0.00225465f $X=15.095 $Y=0.235 $X2=0 $Y2=0
cc_1389 N_Z_c_2279_n N_A_584_47#_M1021_d 0.0025542f $X=11.305 $Y=0.77 $X2=0
+ $Y2=0
cc_1390 N_Z_c_2279_n N_A_584_47#_M1031_d 2.28424e-19 $X=11.305 $Y=0.77 $X2=0
+ $Y2=0
cc_1391 Z N_A_584_47#_M1031_d 0.00152731f $X=11.675 $Y=0.84 $X2=0 $Y2=0
cc_1392 N_Z_c_2280_n N_A_584_47#_M1036_d 7.47571e-19 $X=15.235 $Y=0.73 $X2=0
+ $Y2=0
cc_1393 Z N_A_584_47#_M1036_d 9.93285e-19 $X=11.675 $Y=0.84 $X2=0 $Y2=0
cc_1394 N_Z_c_2280_n N_A_584_47#_M1053_d 0.00172357f $X=15.235 $Y=0.73 $X2=0
+ $Y2=0
cc_1395 N_Z_c_2280_n N_A_584_47#_M1060_d 0.00172357f $X=15.235 $Y=0.73 $X2=0
+ $Y2=0
cc_1396 N_Z_c_2280_n N_A_584_47#_M1073_d 0.00172357f $X=15.235 $Y=0.73 $X2=0
+ $Y2=0
cc_1397 N_Z_c_2279_n N_A_584_47#_c_2797_n 0.00973416f $X=11.305 $Y=0.77 $X2=0
+ $Y2=0
cc_1398 N_Z_M1017_s N_A_584_47#_c_2835_n 0.00480599f $X=9.695 $Y=0.235 $X2=0
+ $Y2=0
cc_1399 N_Z_M1027_s N_A_584_47#_c_2835_n 0.00480599f $X=10.715 $Y=0.235 $X2=0
+ $Y2=0
cc_1400 N_Z_M1033_s N_A_584_47#_c_2835_n 0.00326414f $X=11.655 $Y=0.235 $X2=0
+ $Y2=0
cc_1401 N_Z_M1048_s N_A_584_47#_c_2835_n 0.00326804f $X=12.515 $Y=0.235 $X2=0
+ $Y2=0
cc_1402 N_Z_M1059_s N_A_584_47#_c_2835_n 0.00326804f $X=13.375 $Y=0.235 $X2=0
+ $Y2=0
cc_1403 N_Z_M1067_s N_A_584_47#_c_2835_n 0.00326804f $X=14.235 $Y=0.235 $X2=0
+ $Y2=0
cc_1404 N_Z_M1081_s N_A_584_47#_c_2835_n 0.00326804f $X=15.095 $Y=0.235 $X2=0
+ $Y2=0
cc_1405 N_Z_c_2279_n N_A_584_47#_c_2835_n 0.085013f $X=11.305 $Y=0.77 $X2=0
+ $Y2=0
cc_1406 N_Z_c_2280_n N_A_584_47#_c_2835_n 0.160921f $X=15.235 $Y=0.73 $X2=0
+ $Y2=0
cc_1407 Z N_A_584_47#_c_2835_n 0.0531751f $X=11.675 $Y=0.84 $X2=0 $Y2=0
cc_1408 N_VGND_c_2515_n N_A_584_47#_M1003_s 0.00232985f $X=24.72 $Y=0 $X2=-0.19
+ $Y2=-0.245
cc_1409 N_VGND_c_2515_n N_A_584_47#_M1011_s 0.00266361f $X=24.72 $Y=0 $X2=0
+ $Y2=0
cc_1410 N_VGND_c_2515_n N_A_584_47#_M1016_s 0.00266361f $X=24.72 $Y=0 $X2=0
+ $Y2=0
cc_1411 N_VGND_c_2515_n N_A_584_47#_M1039_s 0.0022543f $X=24.72 $Y=0 $X2=0 $Y2=0
cc_1412 N_VGND_c_2515_n N_A_584_47#_M1045_s 0.0022543f $X=24.72 $Y=0 $X2=0 $Y2=0
cc_1413 N_VGND_c_2515_n N_A_584_47#_M1051_s 0.0022543f $X=24.72 $Y=0 $X2=0 $Y2=0
cc_1414 N_VGND_c_2515_n N_A_584_47#_M1066_s 0.0022543f $X=24.72 $Y=0 $X2=0 $Y2=0
cc_1415 N_VGND_c_2515_n N_A_584_47#_M1080_s 0.0022543f $X=24.72 $Y=0 $X2=0 $Y2=0
cc_1416 N_VGND_c_2515_n N_A_584_47#_M1021_d 0.00289079f $X=24.72 $Y=0 $X2=0
+ $Y2=0
cc_1417 N_VGND_c_2515_n N_A_584_47#_M1031_d 0.00223855f $X=24.72 $Y=0 $X2=0
+ $Y2=0
cc_1418 N_VGND_c_2515_n N_A_584_47#_M1036_d 0.00223855f $X=24.72 $Y=0 $X2=0
+ $Y2=0
cc_1419 N_VGND_c_2515_n N_A_584_47#_M1053_d 0.00223855f $X=24.72 $Y=0 $X2=0
+ $Y2=0
cc_1420 N_VGND_c_2515_n N_A_584_47#_M1060_d 0.00223855f $X=24.72 $Y=0 $X2=0
+ $Y2=0
cc_1421 N_VGND_c_2515_n N_A_584_47#_M1073_d 0.00223855f $X=24.72 $Y=0 $X2=0
+ $Y2=0
cc_1422 N_VGND_c_2515_n N_A_584_47#_M1086_d 0.00299285f $X=24.72 $Y=0 $X2=0
+ $Y2=0
cc_1423 N_VGND_c_2482_n N_A_584_47#_c_2722_n 0.0121355f $X=2.505 $Y=0.28 $X2=0
+ $Y2=0
cc_1424 N_VGND_c_2512_n N_A_584_47#_c_2722_n 0.0195379f $X=3.41 $Y=0 $X2=0 $Y2=0
cc_1425 N_VGND_c_2515_n N_A_584_47#_c_2722_n 0.0125146f $X=24.72 $Y=0 $X2=0
+ $Y2=0
cc_1426 N_VGND_M1003_d N_A_584_47#_c_2735_n 0.00483587f $X=3.355 $Y=0.235 $X2=0
+ $Y2=0
cc_1427 N_VGND_c_2483_n N_A_584_47#_c_2735_n 0.0195333f $X=3.575 $Y=0.385 $X2=0
+ $Y2=0
cc_1428 N_VGND_c_2495_n N_A_584_47#_c_2735_n 0.00244463f $X=4.27 $Y=0 $X2=0
+ $Y2=0
cc_1429 N_VGND_c_2512_n N_A_584_47#_c_2735_n 0.00244463f $X=3.41 $Y=0 $X2=0
+ $Y2=0
cc_1430 N_VGND_c_2515_n N_A_584_47#_c_2735_n 0.010327f $X=24.72 $Y=0 $X2=0 $Y2=0
cc_1431 N_VGND_c_2495_n N_A_584_47#_c_2898_n 0.0108803f $X=4.27 $Y=0 $X2=0 $Y2=0
cc_1432 N_VGND_c_2515_n N_A_584_47#_c_2898_n 0.00645603f $X=24.72 $Y=0 $X2=0
+ $Y2=0
cc_1433 N_VGND_M1015_d N_A_584_47#_c_2745_n 0.00331454f $X=4.295 $Y=0.235 $X2=0
+ $Y2=0
cc_1434 N_VGND_c_2484_n N_A_584_47#_c_2745_n 0.0152929f $X=4.435 $Y=0.385 $X2=0
+ $Y2=0
cc_1435 N_VGND_c_2495_n N_A_584_47#_c_2745_n 0.00244463f $X=4.27 $Y=0 $X2=0
+ $Y2=0
cc_1436 N_VGND_c_2497_n N_A_584_47#_c_2745_n 0.00244463f $X=5.13 $Y=0 $X2=0
+ $Y2=0
cc_1437 N_VGND_c_2515_n N_A_584_47#_c_2745_n 0.0103441f $X=24.72 $Y=0 $X2=0
+ $Y2=0
cc_1438 N_VGND_c_2497_n N_A_584_47#_c_2905_n 0.0108803f $X=5.13 $Y=0 $X2=0 $Y2=0
cc_1439 N_VGND_c_2515_n N_A_584_47#_c_2905_n 0.00645603f $X=24.72 $Y=0 $X2=0
+ $Y2=0
cc_1440 N_VGND_M1035_d N_A_584_47#_c_2749_n 0.00483587f $X=5.155 $Y=0.235 $X2=0
+ $Y2=0
cc_1441 N_VGND_c_2485_n N_A_584_47#_c_2749_n 0.0195333f $X=5.295 $Y=0.385 $X2=0
+ $Y2=0
cc_1442 N_VGND_c_2497_n N_A_584_47#_c_2749_n 0.00244463f $X=5.13 $Y=0 $X2=0
+ $Y2=0
cc_1443 N_VGND_c_2499_n N_A_584_47#_c_2749_n 0.00244463f $X=6.15 $Y=0 $X2=0
+ $Y2=0
cc_1444 N_VGND_c_2515_n N_A_584_47#_c_2749_n 0.010327f $X=24.72 $Y=0 $X2=0 $Y2=0
cc_1445 N_VGND_c_2499_n N_A_584_47#_c_2753_n 0.0176601f $X=6.15 $Y=0 $X2=0 $Y2=0
cc_1446 N_VGND_c_2515_n N_A_584_47#_c_2753_n 0.0124041f $X=24.72 $Y=0 $X2=0
+ $Y2=0
cc_1447 N_VGND_M1044_d N_A_584_47#_c_2757_n 0.00903372f $X=6.095 $Y=0.235 $X2=0
+ $Y2=0
cc_1448 N_VGND_c_2486_n N_A_584_47#_c_2757_n 0.0237737f $X=6.315 $Y=0.385 $X2=0
+ $Y2=0
cc_1449 N_VGND_c_2499_n N_A_584_47#_c_2757_n 0.00244463f $X=6.15 $Y=0 $X2=0
+ $Y2=0
cc_1450 N_VGND_c_2501_n N_A_584_47#_c_2757_n 0.00244463f $X=7.17 $Y=0 $X2=0
+ $Y2=0
cc_1451 N_VGND_c_2515_n N_A_584_47#_c_2757_n 0.0103098f $X=24.72 $Y=0 $X2=0
+ $Y2=0
cc_1452 N_VGND_c_2501_n N_A_584_47#_c_2761_n 0.0178561f $X=7.17 $Y=0 $X2=0 $Y2=0
cc_1453 N_VGND_c_2515_n N_A_584_47#_c_2761_n 0.0124703f $X=24.72 $Y=0 $X2=0
+ $Y2=0
cc_1454 N_VGND_c_2487_n N_A_584_47#_c_2724_n 0.0126012f $X=7.255 $Y=0.515 $X2=0
+ $Y2=0
cc_1455 N_VGND_c_2503_n N_A_584_47#_c_2778_n 0.0178561f $X=8.03 $Y=0 $X2=0 $Y2=0
cc_1456 N_VGND_c_2515_n N_A_584_47#_c_2778_n 0.0124703f $X=24.72 $Y=0 $X2=0
+ $Y2=0
cc_1457 N_VGND_c_2488_n N_A_584_47#_c_2726_n 0.0126012f $X=8.115 $Y=0.515 $X2=0
+ $Y2=0
cc_1458 N_VGND_c_2505_n N_A_584_47#_c_2788_n 0.0178561f $X=8.89 $Y=0 $X2=0 $Y2=0
cc_1459 N_VGND_c_2515_n N_A_584_47#_c_2788_n 0.0124703f $X=24.72 $Y=0 $X2=0
+ $Y2=0
cc_1460 N_VGND_c_2489_n N_A_584_47#_c_2727_n 0.0126012f $X=8.975 $Y=0.515 $X2=0
+ $Y2=0
cc_1461 N_VGND_c_2507_n N_A_584_47#_c_2835_n 0.317426f $X=21.52 $Y=0 $X2=0 $Y2=0
cc_1462 N_VGND_c_2515_n N_A_584_47#_c_2835_n 0.215381f $X=24.72 $Y=0 $X2=0 $Y2=0
cc_1463 N_VGND_c_2507_n N_A_584_47#_c_2800_n 0.017984f $X=21.52 $Y=0 $X2=0 $Y2=0
cc_1464 N_VGND_c_2515_n N_A_584_47#_c_2800_n 0.0125384f $X=24.72 $Y=0 $X2=0
+ $Y2=0
cc_1465 N_VGND_c_2507_n N_A_584_47#_c_2730_n 0.0213034f $X=21.52 $Y=0 $X2=0
+ $Y2=0
cc_1466 N_VGND_c_2515_n N_A_584_47#_c_2730_n 0.0126078f $X=24.72 $Y=0 $X2=0
+ $Y2=0
