* File: sky130_fd_sc_lp__o21bai_0.pex.spice
* Created: Wed Sep  2 10:17:20 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O21BAI_0%B1_N 2 3 4 5 7 10 15 16 17 18 19 24 25
c42 24 0 1.29656e-19 $X=0.27 $Y=1.12
r43 24 25 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.27
+ $Y=1.12 $X2=0.27 $Y2=1.12
r44 18 19 12.183 $w=3.48e-07 $l=3.7e-07 $layer=LI1_cond $X=0.26 $Y=1.665
+ $X2=0.26 $Y2=2.035
r45 17 18 12.183 $w=3.48e-07 $l=3.7e-07 $layer=LI1_cond $X=0.26 $Y=1.295
+ $X2=0.26 $Y2=1.665
r46 17 25 5.76222 $w=3.48e-07 $l=1.75e-07 $layer=LI1_cond $X=0.26 $Y=1.295
+ $X2=0.26 $Y2=1.12
r47 15 24 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.27 $Y=1.46
+ $X2=0.27 $Y2=1.12
r48 15 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.27 $Y=1.46
+ $X2=0.27 $Y2=1.625
r49 8 10 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=0.995 $Y=2.235
+ $X2=0.995 $Y2=2.575
r50 5 24 60.8238 $w=2.1e-07 $l=4.4833e-07 $layer=POLY_cond $X=0.535 $Y=0.785
+ $X2=0.27 $Y2=1.12
r51 5 7 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.535 $Y=0.785
+ $X2=0.535 $Y2=0.465
r52 3 8 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.92 $Y=2.16
+ $X2=0.995 $Y2=2.235
r53 3 4 248.691 $w=1.5e-07 $l=4.85e-07 $layer=POLY_cond $X=0.92 $Y=2.16
+ $X2=0.435 $Y2=2.16
r54 2 4 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.36 $Y=2.085
+ $X2=0.435 $Y2=2.16
r55 2 16 235.872 $w=1.5e-07 $l=4.6e-07 $layer=POLY_cond $X=0.36 $Y=2.085
+ $X2=0.36 $Y2=1.625
.ends

.subckt PM_SKY130_FD_SC_LP__O21BAI_0%A_39_51# 1 2 7 8 10 12 13 15 18 23 25 28 32
+ 34 35 39 40 42
c87 34 0 1.71295e-19 $X=0.675 $Y=0.78
r88 42 43 6.59928 $w=3.08e-07 $l=1.65e-07 $layer=LI1_cond $X=0.77 $Y=2.575
+ $X2=0.77 $Y2=2.41
r89 39 43 49.3246 $w=2.48e-07 $l=1.07e-06 $layer=LI1_cond $X=0.8 $Y=1.34 $X2=0.8
+ $Y2=2.41
r90 39 40 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.84
+ $Y=1.34 $X2=0.84 $Y2=1.34
r91 36 39 21.8964 $w=2.48e-07 $l=4.75e-07 $layer=LI1_cond $X=0.8 $Y=0.865
+ $X2=0.8 $Y2=1.34
r92 34 36 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.675 $Y=0.78
+ $X2=0.8 $Y2=0.865
r93 34 35 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=0.675 $Y=0.78
+ $X2=0.415 $Y2=0.78
r94 30 35 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=0.285 $Y=0.695
+ $X2=0.415 $Y2=0.78
r95 30 32 10.1947 $w=2.58e-07 $l=2.3e-07 $layer=LI1_cond $X=0.285 $Y=0.695
+ $X2=0.285 $Y2=0.465
r96 26 28 71.7872 $w=1.5e-07 $l=1.4e-07 $layer=POLY_cond $X=1.385 $Y=2.14
+ $X2=1.525 $Y2=2.14
r97 21 23 71.7872 $w=1.5e-07 $l=1.4e-07 $layer=POLY_cond $X=1.385 $Y=0.84
+ $X2=1.525 $Y2=0.84
r98 20 40 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=0.84 $Y=1.325
+ $X2=0.84 $Y2=1.34
r99 16 28 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.525 $Y=2.215
+ $X2=1.525 $Y2=2.14
r100 16 18 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=1.525 $Y=2.215
+ $X2=1.525 $Y2=2.685
r101 13 23 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.525 $Y=0.765
+ $X2=1.525 $Y2=0.84
r102 13 15 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.525 $Y=0.765
+ $X2=1.525 $Y2=0.445
r103 12 26 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.385 $Y=2.065
+ $X2=1.385 $Y2=2.14
r104 11 25 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.385 $Y=1.325
+ $X2=1.385 $Y2=1.25
r105 11 12 379.447 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=1.385 $Y=1.325
+ $X2=1.385 $Y2=2.065
r106 10 25 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.385 $Y=1.175
+ $X2=1.385 $Y2=1.25
r107 9 21 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.385 $Y=0.915
+ $X2=1.385 $Y2=0.84
r108 9 10 133.319 $w=1.5e-07 $l=2.6e-07 $layer=POLY_cond $X=1.385 $Y=0.915
+ $X2=1.385 $Y2=1.175
r109 8 20 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=1.005 $Y=1.25
+ $X2=0.84 $Y2=1.325
r110 7 25 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.31 $Y=1.25
+ $X2=1.385 $Y2=1.25
r111 7 8 156.394 $w=1.5e-07 $l=3.05e-07 $layer=POLY_cond $X=1.31 $Y=1.25
+ $X2=1.005 $Y2=1.25
r112 2 42 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=0.655
+ $Y=2.365 $X2=0.78 $Y2=2.575
r113 1 32 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.195
+ $Y=0.255 $X2=0.32 $Y2=0.465
.ends

.subckt PM_SKY130_FD_SC_LP__O21BAI_0%A2 3 7 11 12 13 14 18
c44 18 0 6.20788e-20 $X=1.865 $Y=1.32
c45 11 0 1.4009e-19 $X=1.865 $Y=1.66
r46 18 19 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.865
+ $Y=1.32 $X2=1.865 $Y2=1.32
r47 14 19 8.68731 $w=4.73e-07 $l=3.45e-07 $layer=LI1_cond $X=1.792 $Y=1.665
+ $X2=1.792 $Y2=1.32
r48 13 19 0.629515 $w=4.73e-07 $l=2.5e-08 $layer=LI1_cond $X=1.792 $Y=1.295
+ $X2=1.792 $Y2=1.32
r49 11 18 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.865 $Y=1.66
+ $X2=1.865 $Y2=1.32
r50 11 12 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.865 $Y=1.66
+ $X2=1.865 $Y2=1.825
r51 10 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.865 $Y=1.155
+ $X2=1.865 $Y2=1.32
r52 7 12 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=1.955 $Y=2.685
+ $X2=1.955 $Y2=1.825
r53 3 10 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=1.955 $Y=0.445
+ $X2=1.955 $Y2=1.155
.ends

.subckt PM_SKY130_FD_SC_LP__O21BAI_0%A1 3 7 11 12 13 14 15 20
r32 20 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.435
+ $Y=1.375 $X2=2.435 $Y2=1.375
r33 14 15 9.58211 $w=4.43e-07 $l=3.7e-07 $layer=LI1_cond $X=2.572 $Y=1.665
+ $X2=2.572 $Y2=2.035
r34 14 21 7.5103 $w=4.43e-07 $l=2.9e-07 $layer=LI1_cond $X=2.572 $Y=1.665
+ $X2=2.572 $Y2=1.375
r35 13 21 2.07181 $w=4.43e-07 $l=8e-08 $layer=LI1_cond $X=2.572 $Y=1.295
+ $X2=2.572 $Y2=1.375
r36 11 20 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.435 $Y=1.715
+ $X2=2.435 $Y2=1.375
r37 11 12 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.435 $Y=1.715
+ $X2=2.435 $Y2=1.88
r38 10 20 40.8701 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.435 $Y=1.21
+ $X2=2.435 $Y2=1.375
r39 7 10 392.266 $w=1.5e-07 $l=7.65e-07 $layer=POLY_cond $X=2.385 $Y=0.445
+ $X2=2.385 $Y2=1.21
r40 3 12 412.777 $w=1.5e-07 $l=8.05e-07 $layer=POLY_cond $X=2.345 $Y=2.685
+ $X2=2.345 $Y2=1.88
.ends

.subckt PM_SKY130_FD_SC_LP__O21BAI_0%VPWR 1 2 9 11 13 15 17 22 28 32
r31 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r32 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r33 26 32 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r34 25 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r35 23 28 8.88104 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=1.44 $Y=3.33
+ $X2=1.267 $Y2=3.33
r36 23 25 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=1.44 $Y=3.33
+ $X2=2.16 $Y2=3.33
r37 22 31 4.12929 $w=1.7e-07 $l=2.12e-07 $layer=LI1_cond $X=2.455 $Y=3.33
+ $X2=2.667 $Y2=3.33
r38 22 25 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=2.455 $Y=3.33
+ $X2=2.16 $Y2=3.33
r39 20 29 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r40 19 20 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r41 17 28 8.88104 $w=1.7e-07 $l=1.72e-07 $layer=LI1_cond $X=1.095 $Y=3.33
+ $X2=1.267 $Y2=3.33
r42 17 19 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.095 $Y=3.33
+ $X2=0.72 $Y2=3.33
r43 15 26 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=2.16 $Y2=3.33
r44 15 29 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=1.2 $Y2=3.33
r45 11 31 3.1554 $w=2.7e-07 $l=1.17346e-07 $layer=LI1_cond $X=2.59 $Y=3.245
+ $X2=2.667 $Y2=3.33
r46 11 13 31.3721 $w=2.68e-07 $l=7.35e-07 $layer=LI1_cond $X=2.59 $Y=3.245
+ $X2=2.59 $Y2=2.51
r47 7 28 1.03204 $w=3.45e-07 $l=8.5e-08 $layer=LI1_cond $X=1.267 $Y=3.245
+ $X2=1.267 $Y2=3.33
r48 7 9 24.552 $w=3.43e-07 $l=7.35e-07 $layer=LI1_cond $X=1.267 $Y=3.245
+ $X2=1.267 $Y2=2.51
r49 2 13 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=2.42
+ $Y=2.365 $X2=2.56 $Y2=2.51
r50 1 9 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=1.07
+ $Y=2.365 $X2=1.21 $Y2=2.51
.ends

.subckt PM_SKY130_FD_SC_LP__O21BAI_0%Y 1 2 7 11 13 14 15 16 17 26 36 40
c49 13 0 1.03241e-19 $X=1.115 $Y=0.47
r50 40 41 2.2834 $w=3.68e-07 $l=5.5e-08 $layer=LI1_cond $X=1.28 $Y=0.555
+ $X2=1.28 $Y2=0.61
r51 17 26 2.74877 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.24 $Y=2.09 $X2=1.24
+ $Y2=2.005
r52 17 26 1.1127 $w=2.88e-07 $l=2.8e-08 $layer=LI1_cond $X=1.24 $Y=1.977
+ $X2=1.24 $Y2=2.005
r53 16 17 12.3987 $w=2.88e-07 $l=3.12e-07 $layer=LI1_cond $X=1.24 $Y=1.665
+ $X2=1.24 $Y2=1.977
r54 15 16 14.7036 $w=2.88e-07 $l=3.7e-07 $layer=LI1_cond $X=1.24 $Y=1.295
+ $X2=1.24 $Y2=1.665
r55 14 15 14.7036 $w=2.88e-07 $l=3.7e-07 $layer=LI1_cond $X=1.24 $Y=0.925
+ $X2=1.24 $Y2=1.295
r56 13 40 0.467207 $w=3.68e-07 $l=1.5e-08 $layer=LI1_cond $X=1.28 $Y=0.54
+ $X2=1.28 $Y2=0.555
r57 13 36 2.95898 $w=3.68e-07 $l=9.5e-08 $layer=LI1_cond $X=1.28 $Y=0.54
+ $X2=1.28 $Y2=0.445
r58 13 14 11.9218 $w=2.88e-07 $l=3e-07 $layer=LI1_cond $X=1.24 $Y=0.625 $X2=1.24
+ $Y2=0.925
r59 13 41 0.596091 $w=2.88e-07 $l=1.5e-08 $layer=LI1_cond $X=1.24 $Y=0.625
+ $X2=1.24 $Y2=0.61
r60 9 11 12.3057 $w=2.93e-07 $l=3.15e-07 $layer=LI1_cond $X=1.757 $Y=2.175
+ $X2=1.757 $Y2=2.49
r61 8 17 4.68908 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=1.385 $Y=2.09
+ $X2=1.24 $Y2=2.09
r62 7 9 7.47753 $w=1.7e-07 $l=1.84673e-07 $layer=LI1_cond $X=1.61 $Y=2.09
+ $X2=1.757 $Y2=2.175
r63 7 8 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=1.61 $Y=2.09
+ $X2=1.385 $Y2=2.09
r64 2 11 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=1.6
+ $Y=2.365 $X2=1.74 $Y2=2.49
r65 1 36 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=1.185
+ $Y=0.235 $X2=1.31 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__O21BAI_0%VGND 1 2 9 13 15 17 22 29 30 33 36
c39 30 0 2.64147e-20 $X=2.64 $Y=0
c40 22 0 1.71295e-19 $X=2.04 $Y=0
r41 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r42 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r43 30 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=2.16
+ $Y2=0
r44 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r45 27 36 7.34436 $w=1.7e-07 $l=1.33e-07 $layer=LI1_cond $X=2.305 $Y=0 $X2=2.172
+ $Y2=0
r46 27 29 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=2.305 $Y=0 $X2=2.64
+ $Y2=0
r47 26 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r48 25 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r49 23 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.915 $Y=0 $X2=0.75
+ $Y2=0
r50 23 25 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=0.915 $Y=0 $X2=1.68
+ $Y2=0
r51 22 36 7.34436 $w=1.7e-07 $l=1.32e-07 $layer=LI1_cond $X=2.04 $Y=0 $X2=2.172
+ $Y2=0
r52 22 25 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=2.04 $Y=0 $X2=1.68
+ $Y2=0
r53 20 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r54 19 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r55 17 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.585 $Y=0 $X2=0.75
+ $Y2=0
r56 17 19 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.585 $Y=0 $X2=0.24
+ $Y2=0
r57 15 26 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=1.68
+ $Y2=0
r58 15 34 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=0.72
+ $Y2=0
r59 11 36 0.195364 $w=2.65e-07 $l=8.5e-08 $layer=LI1_cond $X=2.172 $Y=0.085
+ $X2=2.172 $Y2=0
r60 11 13 15.6558 $w=2.63e-07 $l=3.6e-07 $layer=LI1_cond $X=2.172 $Y=0.085
+ $X2=2.172 $Y2=0.445
r61 7 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.75 $Y=0.085 $X2=0.75
+ $Y2=0
r62 7 9 11.5244 $w=3.28e-07 $l=3.3e-07 $layer=LI1_cond $X=0.75 $Y=0.085 $X2=0.75
+ $Y2=0.415
r63 2 13 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.03
+ $Y=0.235 $X2=2.17 $Y2=0.445
r64 1 9 182 $w=1.7e-07 $l=2.19089e-07 $layer=licon1_NDIFF $count=1 $X=0.61
+ $Y=0.255 $X2=0.75 $Y2=0.415
.ends

.subckt PM_SKY130_FD_SC_LP__O21BAI_0%A_320_47# 1 2 9 11 12 15
c26 11 0 6.20788e-20 $X=2.475 $Y=0.865
r27 13 15 13.3127 $w=2.88e-07 $l=3.35e-07 $layer=LI1_cond $X=2.62 $Y=0.78
+ $X2=2.62 $Y2=0.445
r28 11 13 7.43784 $w=1.7e-07 $l=1.8262e-07 $layer=LI1_cond $X=2.475 $Y=0.865
+ $X2=2.62 $Y2=0.78
r29 11 12 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=2.475 $Y=0.865
+ $X2=1.87 $Y2=0.865
r30 7 12 7.04737 $w=1.7e-07 $l=1.54771e-07 $layer=LI1_cond $X=1.752 $Y=0.78
+ $X2=1.87 $Y2=0.865
r31 7 9 16.4284 $w=2.33e-07 $l=3.35e-07 $layer=LI1_cond $X=1.752 $Y=0.78
+ $X2=1.752 $Y2=0.445
r32 2 15 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.46
+ $Y=0.235 $X2=2.6 $Y2=0.445
r33 1 9 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.6
+ $Y=0.235 $X2=1.74 $Y2=0.445
.ends

