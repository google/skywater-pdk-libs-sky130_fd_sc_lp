* File: sky130_fd_sc_lp__dfbbn_1.pex.spice
* Created: Fri Aug 28 10:21:09 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__DFBBN_1%CLK_N 3 7 9 10 11 16 17
r24 16 19 88.6355 $w=4.55e-07 $l=5.05e-07 $layer=POLY_cond $X=0.342 $Y=1.12
+ $X2=0.342 $Y2=1.625
r25 16 18 47.0767 $w=4.55e-07 $l=1.65e-07 $layer=POLY_cond $X=0.342 $Y=1.12
+ $X2=0.342 $Y2=0.955
r26 16 17 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.28
+ $Y=1.12 $X2=0.28 $Y2=1.12
r27 10 11 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.28 $Y=1.665
+ $X2=0.28 $Y2=2.035
r28 9 10 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.28 $Y=1.295
+ $X2=0.28 $Y2=1.665
r29 9 17 6.11144 $w=3.28e-07 $l=1.75e-07 $layer=LI1_cond $X=0.28 $Y=1.295
+ $X2=0.28 $Y2=1.12
r30 7 19 564.043 $w=1.5e-07 $l=1.1e-06 $layer=POLY_cond $X=0.495 $Y=2.725
+ $X2=0.495 $Y2=1.625
r31 3 18 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=0.49 $Y=0.545
+ $X2=0.49 $Y2=0.955
.ends

.subckt PM_SKY130_FD_SC_LP__DFBBN_1%D 1 2 3 5 7 8 10 13 15 20
c53 20 0 1.12147e-19 $X=1.915 $Y=1.345
c54 5 0 3.3931e-19 $X=2.225 $Y=2.17
c55 1 0 1.77166e-19 $X=1.975 $Y=1.51
r56 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.915
+ $Y=1.345 $X2=1.915 $Y2=1.345
r57 15 20 8.20679 $w=3.28e-07 $l=2.35e-07 $layer=LI1_cond $X=1.68 $Y=1.345
+ $X2=1.915 $Y2=1.345
r58 11 13 128.191 $w=1.5e-07 $l=2.5e-07 $layer=POLY_cond $X=1.975 $Y=2.095
+ $X2=2.225 $Y2=2.095
r59 8 10 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.36 $Y=1.09 $X2=2.36
+ $Y2=0.805
r60 5 13 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.225 $Y=2.17
+ $X2=2.225 $Y2=2.095
r61 5 7 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.225 $Y=2.17 $X2=2.225
+ $Y2=2.455
r62 4 19 29.8144 $w=2.91e-07 $l=2.49199e-07 $layer=POLY_cond $X=2.08 $Y=1.165
+ $X2=1.915 $Y2=1.345
r63 3 8 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.285 $Y=1.165
+ $X2=2.36 $Y2=1.09
r64 3 4 105.117 $w=1.5e-07 $l=2.05e-07 $layer=POLY_cond $X=2.285 $Y=1.165
+ $X2=2.08 $Y2=1.165
r65 2 11 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.975 $Y=2.02
+ $X2=1.975 $Y2=2.095
r66 1 19 38.6072 $w=2.91e-07 $l=1.92678e-07 $layer=POLY_cond $X=1.975 $Y=1.51
+ $X2=1.915 $Y2=1.345
r67 1 2 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=1.975 $Y=1.51
+ $X2=1.975 $Y2=2.02
.ends

.subckt PM_SKY130_FD_SC_LP__DFBBN_1%A_113_67# 1 2 10 14 15 16 17 18 21 26 29 30
+ 32 38 43 46 50 51 53 54 56 57 58 60 61 62 63 64 65 66 69 70 73 77 79 80 84 90
+ 93
c251 93 0 1.6887e-19 $X=7.585 $Y=1.345
c252 80 0 5.9858e-20 $X=0.845 $Y=1.865
c253 50 0 8.05743e-20 $X=3.525 $Y=1.245
r254 84 93 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.585 $Y=1.51
+ $X2=7.585 $Y2=1.345
r255 83 84 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.585
+ $Y=1.51 $X2=7.585 $Y2=1.51
r256 78 90 39.8474 $w=6.29e-07 $l=5.2e-07 $layer=POLY_cond $X=0.945 $Y=1.547
+ $X2=1.465 $Y2=1.547
r257 77 79 6.56744 $w=4.38e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=1.36
+ $X2=0.845 $Y2=1.195
r258 77 78 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.945
+ $Y=1.36 $X2=0.945 $Y2=1.36
r259 75 79 19.7562 $w=2.43e-07 $l=4.2e-07 $layer=LI1_cond $X=0.747 $Y=0.775
+ $X2=0.747 $Y2=1.195
r260 73 75 8.82097 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=0.705 $Y=0.545
+ $X2=0.705 $Y2=0.775
r261 69 70 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=8.485
+ $Y=1.895 $X2=8.485 $Y2=1.895
r262 67 69 39.0659 $w=2.93e-07 $l=1e-06 $layer=LI1_cond $X=8.467 $Y=2.895
+ $X2=8.467 $Y2=1.895
r263 65 67 7.47753 $w=1.7e-07 $l=1.84673e-07 $layer=LI1_cond $X=8.32 $Y=2.98
+ $X2=8.467 $Y2=2.895
r264 65 66 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=8.32 $Y=2.98
+ $X2=7.53 $Y2=2.98
r265 64 66 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.445 $Y=2.895
+ $X2=7.53 $Y2=2.98
r266 63 83 9.00224 $w=2.93e-07 $l=2.13014e-07 $layer=LI1_cond $X=7.445 $Y=1.675
+ $X2=7.555 $Y2=1.51
r267 63 64 79.5936 $w=1.68e-07 $l=1.22e-06 $layer=LI1_cond $X=7.445 $Y=1.675
+ $X2=7.445 $Y2=2.895
r268 61 83 14.157 $w=2.93e-07 $l=4.26497e-07 $layer=LI1_cond $X=7.36 $Y=1.17
+ $X2=7.555 $Y2=1.51
r269 61 62 45.9947 $w=1.68e-07 $l=7.05e-07 $layer=LI1_cond $X=7.36 $Y=1.17
+ $X2=6.655 $Y2=1.17
r270 60 62 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.57 $Y=1.085
+ $X2=6.655 $Y2=1.17
r271 59 60 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=6.57 $Y=0.435
+ $X2=6.57 $Y2=1.085
r272 57 59 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.485 $Y=0.35
+ $X2=6.57 $Y2=0.435
r273 57 58 106.016 $w=1.68e-07 $l=1.625e-06 $layer=LI1_cond $X=6.485 $Y=0.35
+ $X2=4.86 $Y2=0.35
r274 55 58 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.775 $Y=0.435
+ $X2=4.86 $Y2=0.35
r275 55 56 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=4.775 $Y=0.435
+ $X2=4.775 $Y2=1.055
r276 53 56 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.69 $Y=1.14
+ $X2=4.775 $Y2=1.055
r277 53 54 69.8075 $w=1.68e-07 $l=1.07e-06 $layer=LI1_cond $X=4.69 $Y=1.14
+ $X2=3.62 $Y2=1.14
r278 50 51 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.525
+ $Y=1.245 $X2=3.525 $Y2=1.245
r279 48 54 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=3.525 $Y=1.225
+ $X2=3.62 $Y2=1.14
r280 48 50 1.16746 $w=1.88e-07 $l=2e-08 $layer=LI1_cond $X=3.525 $Y=1.225
+ $X2=3.525 $Y2=1.245
r281 46 80 23.9219 $w=3.28e-07 $l=6.85e-07 $layer=LI1_cond $X=0.79 $Y=2.55
+ $X2=0.79 $Y2=1.865
r282 43 80 6.50835 $w=4.38e-07 $l=2.2e-07 $layer=LI1_cond $X=0.845 $Y=1.645
+ $X2=0.845 $Y2=1.865
r283 42 77 1.44055 $w=4.38e-07 $l=5.5e-08 $layer=LI1_cond $X=0.845 $Y=1.415
+ $X2=0.845 $Y2=1.36
r284 42 43 6.02413 $w=4.38e-07 $l=2.3e-07 $layer=LI1_cond $X=0.845 $Y=1.415
+ $X2=0.845 $Y2=1.645
r285 38 70 71.6931 $w=3.3e-07 $l=4.1e-07 $layer=POLY_cond $X=8.485 $Y=2.305
+ $X2=8.485 $Y2=1.895
r286 35 38 161.521 $w=1.5e-07 $l=3.15e-07 $layer=POLY_cond $X=8.17 $Y=2.38
+ $X2=8.485 $Y2=2.38
r287 34 51 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.525 $Y=1.08
+ $X2=3.525 $Y2=1.245
r288 30 35 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.17 $Y=2.455
+ $X2=8.17 $Y2=2.38
r289 30 32 101.22 $w=1.5e-07 $l=3.15e-07 $layer=POLY_cond $X=8.17 $Y=2.455
+ $X2=8.17 $Y2=2.77
r290 29 93 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=7.645 $Y=0.915
+ $X2=7.645 $Y2=1.345
r291 26 34 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=3.435 $Y=0.76
+ $X2=3.435 $Y2=1.08
r292 23 26 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=3.435 $Y=0.255
+ $X2=3.435 $Y2=0.76
r293 19 21 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=2.655 $Y=3.005
+ $X2=2.655 $Y2=2.455
r294 17 19 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.58 $Y=3.08
+ $X2=2.655 $Y2=3.005
r295 17 18 471.745 $w=1.5e-07 $l=9.2e-07 $layer=POLY_cond $X=2.58 $Y=3.08
+ $X2=1.66 $Y2=3.08
r296 15 23 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.36 $Y=0.18
+ $X2=3.435 $Y2=0.255
r297 15 16 933.234 $w=1.5e-07 $l=1.82e-06 $layer=POLY_cond $X=3.36 $Y=0.18
+ $X2=1.54 $Y2=0.18
r298 12 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.585 $Y=3.005
+ $X2=1.66 $Y2=3.08
r299 12 14 225.617 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=1.585 $Y=3.005
+ $X2=1.585 $Y2=2.565
r300 11 90 9.19555 $w=6.29e-07 $l=4.08618e-07 $layer=POLY_cond $X=1.585 $Y=1.9
+ $X2=1.465 $Y2=1.547
r301 11 14 340.989 $w=1.5e-07 $l=6.65e-07 $layer=POLY_cond $X=1.585 $Y=1.9
+ $X2=1.585 $Y2=2.565
r302 8 90 37.3022 $w=1.5e-07 $l=3.52e-07 $layer=POLY_cond $X=1.465 $Y=1.195
+ $X2=1.465 $Y2=1.547
r303 8 10 199.979 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=1.465 $Y=1.195
+ $X2=1.465 $Y2=0.805
r304 7 16 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.465 $Y=0.255
+ $X2=1.54 $Y2=0.18
r305 7 10 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=1.465 $Y=0.255
+ $X2=1.465 $Y2=0.805
r306 2 46 300 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_PDIFF $count=2 $X=0.57
+ $Y=2.405 $X2=0.79 $Y2=2.55
r307 1 73 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.565
+ $Y=0.335 $X2=0.705 $Y2=0.545
.ends

.subckt PM_SKY130_FD_SC_LP__DFBBN_1%A_755_398# 1 2 7 9 12 14 16 20 24 27 28 29
+ 30 31 33 36 38 39 41 45 51 59
c152 45 0 1.99763e-19 $X=5.715 $Y=1.13
r153 55 57 10.6379 $w=2.58e-07 $l=2.4e-07 $layer=LI1_cond $X=6.22 $Y=1.565
+ $X2=6.46 $Y2=1.565
r154 51 53 6.80989 $w=3.28e-07 $l=1.95e-07 $layer=LI1_cond $X=5.85 $Y=2.395
+ $X2=5.85 $Y2=2.59
r155 45 47 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=5.715 $Y=1.13
+ $X2=5.715 $Y2=1.21
r156 41 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.015
+ $Y=1.565 $X2=7.015 $Y2=1.565
r157 39 57 3.7676 $w=2.58e-07 $l=8.5e-08 $layer=LI1_cond $X=6.545 $Y=1.565
+ $X2=6.46 $Y2=1.565
r158 39 41 20.8326 $w=2.58e-07 $l=4.7e-07 $layer=LI1_cond $X=6.545 $Y=1.565
+ $X2=7.015 $Y2=1.565
r159 37 57 3.22376 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=6.46 $Y=1.695
+ $X2=6.46 $Y2=1.565
r160 37 38 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=6.46 $Y=1.695
+ $X2=6.46 $Y2=1.915
r161 36 55 3.22376 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=6.22 $Y=1.435
+ $X2=6.22 $Y2=1.565
r162 35 36 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=6.22 $Y=1.295
+ $X2=6.22 $Y2=1.435
r163 34 50 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.015 $Y=2 $X2=5.85
+ $Y2=2
r164 33 38 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.375 $Y=2
+ $X2=6.46 $Y2=1.915
r165 33 34 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=6.375 $Y=2
+ $X2=6.015 $Y2=2
r166 32 47 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.88 $Y=1.21
+ $X2=5.715 $Y2=1.21
r167 31 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.135 $Y=1.21
+ $X2=6.22 $Y2=1.295
r168 31 32 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=6.135 $Y=1.21
+ $X2=5.88 $Y2=1.21
r169 30 51 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=5.85 $Y=2.31
+ $X2=5.85 $Y2=2.395
r170 29 50 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.85 $Y=2.085
+ $X2=5.85 $Y2=2
r171 29 30 7.85757 $w=3.28e-07 $l=2.25e-07 $layer=LI1_cond $X=5.85 $Y=2.085
+ $X2=5.85 $Y2=2.31
r172 27 51 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.685 $Y=2.395
+ $X2=5.85 $Y2=2.395
r173 27 28 87.4225 $w=1.68e-07 $l=1.34e-06 $layer=LI1_cond $X=5.685 $Y=2.395
+ $X2=4.345 $Y2=2.395
r174 25 59 35.3761 $w=3.27e-07 $l=2.4e-07 $layer=POLY_cond $X=4.245 $Y=1.947
+ $X2=4.005 $Y2=1.947
r175 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.245
+ $Y=1.92 $X2=4.245 $Y2=1.92
r176 22 28 6.85817 $w=1.7e-07 $l=1.33918e-07 $layer=LI1_cond $X=4.247 $Y=2.31
+ $X2=4.345 $Y2=2.395
r177 22 24 22.1818 $w=1.93e-07 $l=3.9e-07 $layer=LI1_cond $X=4.247 $Y=2.31
+ $X2=4.247 $Y2=1.92
r178 18 42 38.7084 $w=3.43e-07 $l=2.11069e-07 $layer=POLY_cond $X=7.135 $Y=1.4
+ $X2=7.03 $Y2=1.565
r179 18 20 248.691 $w=1.5e-07 $l=4.85e-07 $layer=POLY_cond $X=7.135 $Y=1.4
+ $X2=7.135 $Y2=0.915
r180 14 42 38.7084 $w=3.43e-07 $l=1.98997e-07 $layer=POLY_cond $X=7.105 $Y=1.73
+ $X2=7.03 $Y2=1.565
r181 14 16 299.968 $w=1.5e-07 $l=5.85e-07 $layer=POLY_cond $X=7.105 $Y=1.73
+ $X2=7.105 $Y2=2.315
r182 10 59 21.0057 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=4.005 $Y=1.755
+ $X2=4.005 $Y2=1.947
r183 10 12 510.202 $w=1.5e-07 $l=9.95e-07 $layer=POLY_cond $X=4.005 $Y=1.755
+ $X2=4.005 $Y2=0.76
r184 7 59 22.8471 $w=3.27e-07 $l=2.5916e-07 $layer=POLY_cond $X=3.85 $Y=2.14
+ $X2=4.005 $Y2=1.947
r185 7 9 101.22 $w=1.5e-07 $l=3.15e-07 $layer=POLY_cond $X=3.85 $Y=2.14 $X2=3.85
+ $Y2=2.455
r186 2 53 600 $w=1.7e-07 $l=9.98774e-07 $layer=licon1_PDIFF $count=1 $X=5.14
+ $Y=1.895 $X2=5.85 $Y2=2.59
r187 2 50 600 $w=1.7e-07 $l=7.97151e-07 $layer=licon1_PDIFF $count=1 $X=5.14
+ $Y=1.895 $X2=5.85 $Y2=2.08
r188 1 45 182 $w=1.7e-07 $l=9.0111e-07 $layer=licon1_NDIFF $count=1 $X=5.5
+ $Y=0.33 $X2=5.715 $Y2=1.13
.ends

.subckt PM_SKY130_FD_SC_LP__DFBBN_1%SET_B 3 7 11 14 15 17 20 22 24 25 31 35 36
+ 40
c141 11 0 8.77366e-20 $X=9.405 $Y=0.915
r142 40 43 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=9.415 $Y=1.665
+ $X2=9.415 $Y2=1.83
r143 40 42 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=9.415 $Y=1.665
+ $X2=9.415 $Y2=1.5
r144 35 38 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.975 $Y=1.57
+ $X2=4.975 $Y2=1.735
r145 35 37 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.975 $Y=1.57
+ $X2=4.975 $Y2=1.405
r146 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.975
+ $Y=1.57 $X2=4.975 $Y2=1.57
r147 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=1.665
+ $X2=8.88 $Y2=1.665
r148 27 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=1.665
+ $X2=5.04 $Y2=1.665
r149 25 27 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.185 $Y=1.665
+ $X2=5.04 $Y2=1.665
r150 24 31 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.735 $Y=1.665
+ $X2=8.88 $Y2=1.665
r151 24 25 4.39356 $w=1.4e-07 $l=3.55e-06 $layer=MET1_cond $X=8.735 $Y=1.665
+ $X2=5.185 $Y2=1.665
r152 22 32 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=9.36 $Y=1.665
+ $X2=8.88 $Y2=1.665
r153 22 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.415
+ $Y=1.665 $X2=9.415 $Y2=1.665
r154 18 20 87.1702 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=9.505 $Y=2.105
+ $X2=9.675 $Y2=2.105
r155 15 20 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.675 $Y=2.18
+ $X2=9.675 $Y2=2.105
r156 15 17 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=9.675 $Y=2.18
+ $X2=9.675 $Y2=2.675
r157 14 18 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.505 $Y=2.03
+ $X2=9.505 $Y2=2.105
r158 14 43 102.553 $w=1.5e-07 $l=2e-07 $layer=POLY_cond $X=9.505 $Y=2.03
+ $X2=9.505 $Y2=1.83
r159 11 42 299.968 $w=1.5e-07 $l=5.85e-07 $layer=POLY_cond $X=9.405 $Y=0.915
+ $X2=9.405 $Y2=1.5
r160 7 38 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=5.065 $Y=2.315
+ $X2=5.065 $Y2=1.735
r161 3 37 387.138 $w=1.5e-07 $l=7.55e-07 $layer=POLY_cond $X=4.99 $Y=0.65
+ $X2=4.99 $Y2=1.405
.ends

.subckt PM_SKY130_FD_SC_LP__DFBBN_1%A_546_449# 1 2 9 13 16 17 20 21 22 24 25 26
+ 28 29 31 32 35 42
c146 31 0 2.29376e-20 $X=5.79 $Y=1.57
c147 20 0 2.7703e-20 $X=3.885 $Y=2.225
r148 41 42 9.2801 $w=4.58e-07 $l=1.65e-07 $layer=LI1_cond $X=3.245 $Y=2.455
+ $X2=3.41 $Y2=2.455
r149 38 41 2.08014 $w=4.58e-07 $l=8e-08 $layer=LI1_cond $X=3.165 $Y=2.455
+ $X2=3.245 $Y2=2.455
r150 35 37 10.0337 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=3.085 $Y=0.74
+ $X2=3.085 $Y2=0.95
r151 32 45 49.6442 $w=2.67e-07 $l=2.75e-07 $layer=POLY_cond $X=5.79 $Y=1.57
+ $X2=6.065 $Y2=1.57
r152 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.79
+ $Y=1.57 $X2=5.79 $Y2=1.57
r153 29 31 12.6325 $w=2.58e-07 $l=2.85e-07 $layer=LI1_cond $X=5.505 $Y=1.605
+ $X2=5.79 $Y2=1.605
r154 27 29 7.21222 $w=2.6e-07 $l=1.67183e-07 $layer=LI1_cond $X=5.42 $Y=1.735
+ $X2=5.505 $Y2=1.605
r155 27 28 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=5.42 $Y=1.735
+ $X2=5.42 $Y2=1.96
r156 25 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.335 $Y=2.045
+ $X2=5.42 $Y2=1.96
r157 25 26 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=5.335 $Y=2.045
+ $X2=4.695 $Y2=2.045
r158 24 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.61 $Y=1.96
+ $X2=4.695 $Y2=2.045
r159 23 24 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=4.61 $Y=1.575
+ $X2=4.61 $Y2=1.96
r160 21 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.525 $Y=1.49
+ $X2=4.61 $Y2=1.575
r161 21 22 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=4.525 $Y=1.49
+ $X2=3.97 $Y2=1.49
r162 19 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.885 $Y=1.575
+ $X2=3.97 $Y2=1.49
r163 19 20 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=3.885 $Y=1.575
+ $X2=3.885 $Y2=2.225
r164 17 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.8 $Y=2.31
+ $X2=3.885 $Y2=2.225
r165 17 42 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=3.8 $Y=2.31
+ $X2=3.41 $Y2=2.31
r166 16 38 6.6364 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=3.165 $Y=2.225
+ $X2=3.165 $Y2=2.455
r167 16 37 83.1818 $w=1.68e-07 $l=1.275e-06 $layer=LI1_cond $X=3.165 $Y=2.225
+ $X2=3.165 $Y2=0.95
r168 11 45 16.2448 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.065 $Y=1.735
+ $X2=6.065 $Y2=1.57
r169 11 13 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=6.065 $Y=1.735
+ $X2=6.065 $Y2=2.315
r170 7 32 65.8914 $w=2.67e-07 $l=4.39829e-07 $layer=POLY_cond $X=5.425 $Y=1.405
+ $X2=5.79 $Y2=1.57
r171 7 9 387.138 $w=1.5e-07 $l=7.55e-07 $layer=POLY_cond $X=5.425 $Y=1.405
+ $X2=5.425 $Y2=0.65
r172 2 41 600 $w=1.7e-07 $l=6.11044e-07 $layer=licon1_PDIFF $count=1 $X=2.73
+ $Y=2.245 $X2=3.245 $Y2=2.455
r173 1 35 182 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_NDIFF $count=1 $X=2.865
+ $Y=0.595 $X2=3.085 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LP__DFBBN_1%A_223_119# 1 2 9 12 13 14 18 19 20 24 25 26
+ 28 29 30 31 33 34 35 37 39 42 43 47 51
c166 47 0 3.67402e-20 $X=2.455 $Y=1.645
c167 39 0 1.65878e-19 $X=1.37 $Y=2.39
c168 37 0 1.73432e-19 $X=1.37 $Y=2.21
c169 35 0 8.05743e-20 $X=2.79 $Y=1.66
c170 34 0 1.12147e-19 $X=2.715 $Y=1.645
c171 12 0 2.7703e-20 $X=3.045 $Y=2.02
r172 51 53 10.3829 $w=3.28e-07 $l=2.2e-07 $layer=LI1_cond $X=1.25 $Y=0.795
+ $X2=1.25 $Y2=1.015
r173 47 48 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.455
+ $Y=1.645 $X2=2.455 $Y2=1.645
r174 45 47 10.1947 $w=2.58e-07 $l=2.3e-07 $layer=LI1_cond $X=2.42 $Y=1.875
+ $X2=2.42 $Y2=1.645
r175 44 54 4.23499 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.535 $Y=1.96
+ $X2=1.37 $Y2=1.96
r176 43 45 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=2.29 $Y=1.96
+ $X2=2.42 $Y2=1.875
r177 43 44 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=2.29 $Y=1.96
+ $X2=1.535 $Y2=1.96
r178 42 54 5.80639 $w=3.09e-07 $l=1.03078e-07 $layer=LI1_cond $X=1.33 $Y=1.875
+ $X2=1.37 $Y2=1.96
r179 42 53 56.107 $w=1.68e-07 $l=8.6e-07 $layer=LI1_cond $X=1.33 $Y=1.875
+ $X2=1.33 $Y2=1.015
r180 37 54 9.30818 $w=3.3e-07 $l=2.5e-07 $layer=LI1_cond $X=1.37 $Y=2.21
+ $X2=1.37 $Y2=1.96
r181 37 39 6.28605 $w=3.28e-07 $l=1.8e-07 $layer=LI1_cond $X=1.37 $Y=2.21
+ $X2=1.37 $Y2=2.39
r182 35 36 56.9028 $w=2.16e-07 $l=2.55e-07 $layer=POLY_cond $X=2.79 $Y=1.66
+ $X2=3.045 $Y2=1.66
r183 34 48 45.4639 $w=3.3e-07 $l=2.6e-07 $layer=POLY_cond $X=2.715 $Y=1.645
+ $X2=2.455 $Y2=1.645
r184 34 35 16.704 $w=3.3e-07 $l=8.21584e-08 $layer=POLY_cond $X=2.715 $Y=1.645
+ $X2=2.79 $Y2=1.66
r185 31 33 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=8.39 $Y=1.31
+ $X2=8.39 $Y2=1.025
r186 29 31 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.315 $Y=1.385
+ $X2=8.39 $Y2=1.31
r187 29 30 105.117 $w=1.5e-07 $l=2.05e-07 $layer=POLY_cond $X=8.315 $Y=1.385
+ $X2=8.11 $Y2=1.385
r188 27 30 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.035 $Y=1.46
+ $X2=8.11 $Y2=1.385
r189 27 28 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=8.035 $Y=1.46
+ $X2=8.035 $Y2=1.915
r190 25 28 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.96 $Y=1.99
+ $X2=8.035 $Y2=1.915
r191 25 26 156.394 $w=1.5e-07 $l=3.05e-07 $layer=POLY_cond $X=7.96 $Y=1.99
+ $X2=7.655 $Y2=1.99
r192 22 24 264.074 $w=1.5e-07 $l=5.15e-07 $layer=POLY_cond $X=7.58 $Y=3.075
+ $X2=7.58 $Y2=2.56
r193 21 26 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.58 $Y=2.065
+ $X2=7.655 $Y2=1.99
r194 21 24 253.819 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=7.58 $Y=2.065
+ $X2=7.58 $Y2=2.56
r195 19 22 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.505 $Y=3.15
+ $X2=7.58 $Y2=3.075
r196 19 20 2035.68 $w=1.5e-07 $l=3.97e-06 $layer=POLY_cond $X=7.505 $Y=3.15
+ $X2=3.535 $Y2=3.15
r197 16 20 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.46 $Y=3.075
+ $X2=3.535 $Y2=3.15
r198 16 18 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=3.46 $Y=3.075
+ $X2=3.46 $Y2=2.455
r199 15 18 146.138 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.46 $Y=2.17
+ $X2=3.46 $Y2=2.455
r200 13 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.385 $Y=2.095
+ $X2=3.46 $Y2=2.17
r201 13 14 135.883 $w=1.5e-07 $l=2.65e-07 $layer=POLY_cond $X=3.385 $Y=2.095
+ $X2=3.12 $Y2=2.095
r202 12 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.045 $Y=2.02
+ $X2=3.12 $Y2=2.095
r203 11 36 11.3495 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=3.045 $Y=1.81
+ $X2=3.045 $Y2=1.66
r204 11 12 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=3.045 $Y=1.81
+ $X2=3.045 $Y2=2.02
r205 7 35 11.3495 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=2.79 $Y=1.48
+ $X2=2.79 $Y2=1.66
r206 7 9 346.117 $w=1.5e-07 $l=6.75e-07 $layer=POLY_cond $X=2.79 $Y=1.48
+ $X2=2.79 $Y2=0.805
r207 2 39 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=1.225
+ $Y=2.245 $X2=1.37 $Y2=2.39
r208 1 51 182 $w=1.7e-07 $l=2.58844e-07 $layer=licon1_NDIFF $count=1 $X=1.115
+ $Y=0.595 $X2=1.25 $Y2=0.795
.ends

.subckt PM_SKY130_FD_SC_LP__DFBBN_1%A_1741_137# 1 2 7 9 14 18 21 23 25 27 30 34
+ 36 37 40 44 46 49 50 53 54 56 58 62 66 68 69
c168 56 0 8.77366e-20 $X=10.13 $Y=0.79
c169 54 0 2.45307e-19 $X=9.89 $Y=2.235
c170 36 0 7.06233e-20 $X=12.915 $Y=1.26
r171 68 69 30.474 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=11.92 $Y=1.26
+ $X2=11.92 $Y2=1.185
r172 63 71 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=11.92 $Y=1.35
+ $X2=11.92 $Y2=1.515
r173 63 68 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=11.92 $Y=1.35
+ $X2=11.92 $Y2=1.26
r174 62 63 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.92
+ $Y=1.35 $X2=11.92 $Y2=1.35
r175 59 62 3.84148 $w=3.28e-07 $l=1.1e-07 $layer=LI1_cond $X=11.81 $Y=1.35
+ $X2=11.92 $Y2=1.35
r176 52 59 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.81 $Y=1.515
+ $X2=11.81 $Y2=1.35
r177 52 53 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=11.81 $Y=1.515
+ $X2=11.81 $Y2=2.205
r178 51 58 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.47 $Y=2.29
+ $X2=10.385 $Y2=2.29
r179 50 53 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=11.725 $Y=2.29
+ $X2=11.81 $Y2=2.205
r180 50 51 81.877 $w=1.68e-07 $l=1.255e-06 $layer=LI1_cond $X=11.725 $Y=2.29
+ $X2=10.47 $Y2=2.29
r181 49 58 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.385 $Y=2.205
+ $X2=10.385 $Y2=2.29
r182 48 56 10.37 $w=3e-07 $l=3.37994e-07 $layer=LI1_cond $X=10.385 $Y=1
+ $X2=10.13 $Y2=0.807
r183 48 49 78.615 $w=1.68e-07 $l=1.205e-06 $layer=LI1_cond $X=10.385 $Y=1
+ $X2=10.385 $Y2=2.205
r184 47 54 6.46576 $w=2.5e-07 $l=1.90526e-07 $layer=LI1_cond $X=10.055 $Y=2.29
+ $X2=9.89 $Y2=2.235
r185 46 58 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.3 $Y=2.29
+ $X2=10.385 $Y2=2.29
r186 46 47 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=10.3 $Y=2.29
+ $X2=10.055 $Y2=2.29
r187 44 54 0.364692 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=9.89 $Y=2.4
+ $X2=9.89 $Y2=2.235
r188 40 67 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=9.025 $Y=2.235
+ $X2=9.025 $Y2=2.4
r189 40 66 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=9.025 $Y=2.235
+ $X2=9.025 $Y2=2.07
r190 39 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.025
+ $Y=2.235 $X2=9.025 $Y2=2.235
r191 37 54 6.46576 $w=2.5e-07 $l=1.65e-07 $layer=LI1_cond $X=9.725 $Y=2.235
+ $X2=9.89 $Y2=2.235
r192 37 39 24.4458 $w=3.28e-07 $l=7e-07 $layer=LI1_cond $X=9.725 $Y=2.235
+ $X2=9.025 $Y2=2.235
r193 32 34 79.4787 $w=1.5e-07 $l=1.55e-07 $layer=POLY_cond $X=8.78 $Y=1.385
+ $X2=8.935 $Y2=1.385
r194 28 36 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=12.915 $Y=1.335
+ $X2=12.915 $Y2=1.26
r195 28 30 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=12.915 $Y=1.335
+ $X2=12.915 $Y2=2.155
r196 25 36 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=12.915 $Y=1.185
+ $X2=12.915 $Y2=1.26
r197 25 27 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=12.915 $Y=1.185
+ $X2=12.915 $Y2=0.895
r198 24 68 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=12.085 $Y=1.26
+ $X2=11.92 $Y2=1.26
r199 23 36 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=12.84 $Y=1.26
+ $X2=12.915 $Y2=1.26
r200 23 24 387.138 $w=1.5e-07 $l=7.55e-07 $layer=POLY_cond $X=12.84 $Y=1.26
+ $X2=12.085 $Y2=1.26
r201 21 71 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=11.945 $Y=2.345
+ $X2=11.945 $Y2=1.515
r202 18 69 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=11.925 $Y=0.655
+ $X2=11.925 $Y2=1.185
r203 14 67 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=8.965 $Y=2.77
+ $X2=8.965 $Y2=2.4
r204 10 34 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.935 $Y=1.46
+ $X2=8.935 $Y2=1.385
r205 10 66 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=8.935 $Y=1.46
+ $X2=8.935 $Y2=2.07
r206 7 32 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.78 $Y=1.31
+ $X2=8.78 $Y2=1.385
r207 7 9 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=8.78 $Y=1.31 $X2=8.78
+ $Y2=1.025
r208 2 44 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=9.75
+ $Y=2.255 $X2=9.89 $Y2=2.4
r209 1 56 182 $w=1.7e-07 $l=2.63106e-07 $layer=licon1_NDIFF $count=1 $X=9.97
+ $Y=0.595 $X2=10.13 $Y2=0.79
.ends

.subckt PM_SKY130_FD_SC_LP__DFBBN_1%A_1531_428# 1 2 9 13 15 20 26 29 30 31 35 41
c96 30 0 1.6887e-19 $X=7.905 $Y=2.12
r97 36 41 26.2292 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=9.955 $Y=1.625
+ $X2=10.105 $Y2=1.625
r98 36 38 10.4917 $w=3.3e-07 $l=6e-08 $layer=POLY_cond $X=9.955 $Y=1.625
+ $X2=9.895 $Y2=1.625
r99 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.955
+ $Y=1.625 $X2=9.955 $Y2=1.625
r100 32 35 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=9.86 $Y=1.625
+ $X2=9.955 $Y2=1.625
r101 29 32 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.86 $Y=1.46
+ $X2=9.86 $Y2=1.625
r102 28 29 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=9.86 $Y=1.32
+ $X2=9.86 $Y2=1.46
r103 27 31 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.26 $Y=1.235
+ $X2=8.095 $Y2=1.235
r104 26 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.775 $Y=1.235
+ $X2=9.86 $Y2=1.32
r105 26 27 98.8396 $w=1.68e-07 $l=1.515e-06 $layer=LI1_cond $X=9.775 $Y=1.235
+ $X2=8.26 $Y2=1.235
r106 24 31 3.70735 $w=2.5e-07 $l=1.18427e-07 $layer=LI1_cond $X=8.015 $Y=1.32
+ $X2=8.095 $Y2=1.235
r107 24 30 52.1925 $w=1.68e-07 $l=8e-07 $layer=LI1_cond $X=8.015 $Y=1.32
+ $X2=8.015 $Y2=2.12
r108 20 23 12.2229 $w=3.28e-07 $l=3.5e-07 $layer=LI1_cond $X=8.095 $Y=0.74
+ $X2=8.095 $Y2=1.09
r109 18 31 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=8.095 $Y=1.15
+ $X2=8.095 $Y2=1.235
r110 18 23 2.09535 $w=3.28e-07 $l=6e-08 $layer=LI1_cond $X=8.095 $Y=1.15
+ $X2=8.095 $Y2=1.09
r111 15 30 9.49412 $w=3.88e-07 $l=1.95e-07 $layer=LI1_cond $X=7.905 $Y=2.315
+ $X2=7.905 $Y2=2.12
r112 15 17 3.12821 $w=3.9e-07 $l=1e-07 $layer=LI1_cond $X=7.905 $Y=2.315
+ $X2=7.905 $Y2=2.415
r113 11 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.105 $Y=1.79
+ $X2=10.105 $Y2=1.625
r114 11 13 453.798 $w=1.5e-07 $l=8.85e-07 $layer=POLY_cond $X=10.105 $Y=1.79
+ $X2=10.105 $Y2=2.675
r115 7 38 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.895 $Y=1.46
+ $X2=9.895 $Y2=1.625
r116 7 9 279.457 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=9.895 $Y=1.46
+ $X2=9.895 $Y2=0.915
r117 2 17 600 $w=1.7e-07 $l=3.68951e-07 $layer=licon1_PDIFF $count=1 $X=7.655
+ $Y=2.14 $X2=7.875 $Y2=2.415
r118 1 23 182 $w=1.7e-07 $l=6.56239e-07 $layer=licon1_NDIFF $count=1 $X=7.72
+ $Y=0.595 $X2=8.095 $Y2=1.09
r119 1 20 182 $w=1.7e-07 $l=4.41588e-07 $layer=licon1_NDIFF $count=1 $X=7.72
+ $Y=0.595 $X2=8.095 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LP__DFBBN_1%A_1186_21# 1 2 10 11 12 13 14 17 22 23 25 26
+ 27 29 32 34 37 39 41 46
c120 32 0 1.21191e-19 $X=10.725 $Y=2.105
c121 23 0 1.24116e-19 $X=10.465 $Y=2.18
c122 14 0 2.227e-19 $X=6.08 $Y=1.12
r123 39 41 8.55602 $w=3.28e-07 $l=2.45e-07 $layer=LI1_cond $X=10.98 $Y=1.86
+ $X2=11.225 $Y2=1.86
r124 38 49 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=10.815 $Y=1.35
+ $X2=10.815 $Y2=1.515
r125 38 46 30.6007 $w=3.3e-07 $l=1.75e-07 $layer=POLY_cond $X=10.815 $Y=1.35
+ $X2=10.815 $Y2=1.175
r126 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.815
+ $Y=1.35 $X2=10.815 $Y2=1.35
r127 35 39 6.81649 $w=3.3e-07 $l=2.33345e-07 $layer=LI1_cond $X=10.815 $Y=1.695
+ $X2=10.98 $Y2=1.86
r128 35 37 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=10.815 $Y=1.695
+ $X2=10.815 $Y2=1.35
r129 34 45 18.0654 $w=2.6e-07 $l=3.85e-07 $layer=LI1_cond $X=10.815 $Y=0.83
+ $X2=11.2 $Y2=0.83
r130 34 37 12.2229 $w=3.28e-07 $l=3.5e-07 $layer=LI1_cond $X=10.815 $Y=1
+ $X2=10.815 $Y2=1.35
r131 30 32 133.319 $w=1.5e-07 $l=2.6e-07 $layer=POLY_cond $X=10.465 $Y=2.105
+ $X2=10.725 $Y2=2.105
r132 29 32 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=10.725 $Y=2.03
+ $X2=10.725 $Y2=2.105
r133 29 49 264.074 $w=1.5e-07 $l=5.15e-07 $layer=POLY_cond $X=10.725 $Y=2.03
+ $X2=10.725 $Y2=1.515
r134 26 46 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.65 $Y=1.175
+ $X2=10.815 $Y2=1.175
r135 26 27 105.117 $w=1.5e-07 $l=2.05e-07 $layer=POLY_cond $X=10.65 $Y=1.175
+ $X2=10.445 $Y2=1.175
r136 23 30 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=10.465 $Y=2.18
+ $X2=10.465 $Y2=2.105
r137 23 25 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=10.465 $Y=2.18
+ $X2=10.465 $Y2=2.675
r138 20 27 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=10.37 $Y=1.1
+ $X2=10.445 $Y2=1.175
r139 20 22 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=10.37 $Y=1.1
+ $X2=10.37 $Y2=0.705
r140 19 22 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=10.37 $Y=0.255
+ $X2=10.37 $Y2=0.705
r141 15 17 574.298 $w=1.5e-07 $l=1.12e-06 $layer=POLY_cond $X=6.455 $Y=1.195
+ $X2=6.455 $Y2=2.315
r142 13 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.38 $Y=1.12
+ $X2=6.455 $Y2=1.195
r143 13 14 153.83 $w=1.5e-07 $l=3e-07 $layer=POLY_cond $X=6.38 $Y=1.12 $X2=6.08
+ $Y2=1.12
r144 11 19 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=10.295 $Y=0.18
+ $X2=10.37 $Y2=0.255
r145 11 12 2161.31 $w=1.5e-07 $l=4.215e-06 $layer=POLY_cond $X=10.295 $Y=0.18
+ $X2=6.08 $Y2=0.18
r146 8 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.005 $Y=1.045
+ $X2=6.08 $Y2=1.12
r147 8 10 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=6.005 $Y=1.045
+ $X2=6.005 $Y2=0.65
r148 7 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.005 $Y=0.255
+ $X2=6.08 $Y2=0.18
r149 7 10 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=6.005 $Y=0.255
+ $X2=6.005 $Y2=0.65
r150 2 41 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=11.09
+ $Y=1.715 $X2=11.225 $Y2=1.86
r151 1 45 182 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_NDIFF $count=1 $X=11.055
+ $Y=0.655 $X2=11.2 $Y2=0.815
.ends

.subckt PM_SKY130_FD_SC_LP__DFBBN_1%RESET_B 3 6 8 11 13
c32 13 0 1.37465e-19 $X=11.355 $Y=1.185
r33 11 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=11.355 $Y=1.35
+ $X2=11.355 $Y2=1.515
r34 11 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=11.355 $Y=1.35
+ $X2=11.355 $Y2=1.185
r35 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.355
+ $Y=1.35 $X2=11.355 $Y2=1.35
r36 6 14 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=11.44 $Y=2.035
+ $X2=11.44 $Y2=1.515
r37 3 13 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=11.415 $Y=0.865
+ $X2=11.415 $Y2=1.185
.ends

.subckt PM_SKY130_FD_SC_LP__DFBBN_1%A_2511_137# 1 2 9 13 17 21 25 26 28
c49 28 0 7.06233e-20 $X=12.74 $Y=1.47
c50 21 0 1.76649e-19 $X=12.7 $Y=1.98
r51 26 31 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=13.365 $Y=1.47
+ $X2=13.365 $Y2=1.635
r52 26 30 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=13.365 $Y=1.47
+ $X2=13.365 $Y2=1.305
r53 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=13.365
+ $Y=1.47 $X2=13.365 $Y2=1.47
r54 23 28 0.364692 $w=3.3e-07 $l=1.25e-07 $layer=LI1_cond $X=12.865 $Y=1.47
+ $X2=12.74 $Y2=1.47
r55 23 25 17.4613 $w=3.28e-07 $l=5e-07 $layer=LI1_cond $X=12.865 $Y=1.47
+ $X2=13.365 $Y2=1.47
r56 19 28 6.46576 $w=2.5e-07 $l=1.65e-07 $layer=LI1_cond $X=12.74 $Y=1.635
+ $X2=12.74 $Y2=1.47
r57 19 21 15.9037 $w=2.48e-07 $l=3.45e-07 $layer=LI1_cond $X=12.74 $Y=1.635
+ $X2=12.74 $Y2=1.98
r58 15 28 6.46576 $w=2.5e-07 $l=1.65e-07 $layer=LI1_cond $X=12.74 $Y=1.305
+ $X2=12.74 $Y2=1.47
r59 15 17 18.9001 $w=2.48e-07 $l=4.1e-07 $layer=LI1_cond $X=12.74 $Y=1.305
+ $X2=12.74 $Y2=0.895
r60 13 31 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=13.425 $Y=2.465
+ $X2=13.425 $Y2=1.635
r61 9 30 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=13.425 $Y=0.685
+ $X2=13.425 $Y2=1.305
r62 2 21 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=12.565
+ $Y=1.835 $X2=12.7 $Y2=1.98
r63 1 17 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=12.555
+ $Y=0.685 $X2=12.7 $Y2=0.895
.ends

.subckt PM_SKY130_FD_SC_LP__DFBBN_1%VPWR 1 2 3 4 5 6 7 8 25 27 31 35 39 43 47 51
+ 55 60 61 63 64 66 67 68 83 90 102 106 113 114 120 123 126 129
r143 129 130 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.2 $Y=3.33
+ $X2=13.2 $Y2=3.33
r144 126 127 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.76 $Y=3.33
+ $X2=11.76 $Y2=3.33
r145 123 124 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r146 117 118 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r147 114 130 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.68 $Y=3.33
+ $X2=13.2 $Y2=3.33
r148 113 114 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.68 $Y=3.33
+ $X2=13.68 $Y2=3.33
r149 111 129 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=13.295 $Y=3.33
+ $X2=13.17 $Y2=3.33
r150 111 113 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=13.295 $Y=3.33
+ $X2=13.68 $Y2=3.33
r151 110 130 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.72 $Y=3.33
+ $X2=13.2 $Y2=3.33
r152 110 127 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=12.72 $Y=3.33
+ $X2=11.76 $Y2=3.33
r153 109 110 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=12.72 $Y=3.33
+ $X2=12.72 $Y2=3.33
r154 107 126 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.895 $Y=3.33
+ $X2=11.73 $Y2=3.33
r155 107 109 53.8235 $w=1.68e-07 $l=8.25e-07 $layer=LI1_cond $X=11.895 $Y=3.33
+ $X2=12.72 $Y2=3.33
r156 106 129 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=13.045 $Y=3.33
+ $X2=13.17 $Y2=3.33
r157 106 109 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=13.045 $Y=3.33
+ $X2=12.72 $Y2=3.33
r158 105 127 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=3.33
+ $X2=11.76 $Y2=3.33
r159 104 105 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.28 $Y=3.33
+ $X2=11.28 $Y2=3.33
r160 102 126 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.565 $Y=3.33
+ $X2=11.73 $Y2=3.33
r161 102 104 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=11.565 $Y=3.33
+ $X2=11.28 $Y2=3.33
r162 101 105 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=10.32 $Y=3.33
+ $X2=11.28 $Y2=3.33
r163 101 124 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=10.32 $Y=3.33
+ $X2=9.36 $Y2=3.33
r164 100 101 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.32 $Y=3.33
+ $X2=10.32 $Y2=3.33
r165 98 123 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.545 $Y=3.33
+ $X2=9.38 $Y2=3.33
r166 98 100 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=9.545 $Y=3.33
+ $X2=10.32 $Y2=3.33
r167 97 124 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=9.36 $Y2=3.33
r168 96 97 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r169 94 97 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=8.88 $Y2=3.33
r170 93 96 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=7.44 $Y=3.33
+ $X2=8.88 $Y2=3.33
r171 93 94 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r172 91 120 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.055 $Y=3.33
+ $X2=6.89 $Y2=3.33
r173 91 93 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=7.055 $Y=3.33
+ $X2=7.44 $Y2=3.33
r174 90 123 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.215 $Y=3.33
+ $X2=9.38 $Y2=3.33
r175 90 96 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=9.215 $Y=3.33
+ $X2=8.88 $Y2=3.33
r176 88 89 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r177 86 89 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=6.48 $Y2=3.33
r178 85 88 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=5.04 $Y=3.33
+ $X2=6.48 $Y2=3.33
r179 85 86 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r180 83 120 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.725 $Y=3.33
+ $X2=6.89 $Y2=3.33
r181 83 88 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=6.725 $Y=3.33
+ $X2=6.48 $Y2=3.33
r182 82 86 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.04 $Y2=3.33
r183 81 82 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r184 79 82 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=4.56 $Y2=3.33
r185 78 81 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=2.16 $Y=3.33
+ $X2=4.56 $Y2=3.33
r186 78 79 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r187 76 79 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r188 75 76 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r189 73 76 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r190 73 118 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r191 72 75 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r192 72 73 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r193 70 117 4.73185 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=3.33
+ $X2=0.222 $Y2=3.33
r194 70 72 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.445 $Y=3.33
+ $X2=0.72 $Y2=3.33
r195 68 94 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=7.44 $Y2=3.33
r196 68 89 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=6.48 $Y2=3.33
r197 68 120 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r198 66 100 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=10.515 $Y=3.33
+ $X2=10.32 $Y2=3.33
r199 66 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.515 $Y=3.33
+ $X2=10.68 $Y2=3.33
r200 65 104 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=10.845 $Y=3.33
+ $X2=11.28 $Y2=3.33
r201 65 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.845 $Y=3.33
+ $X2=10.68 $Y2=3.33
r202 63 81 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=4.605 $Y=3.33
+ $X2=4.56 $Y2=3.33
r203 63 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.605 $Y=3.33
+ $X2=4.77 $Y2=3.33
r204 62 85 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=4.935 $Y=3.33
+ $X2=5.04 $Y2=3.33
r205 62 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.935 $Y=3.33
+ $X2=4.77 $Y2=3.33
r206 60 75 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=1.715 $Y=3.33
+ $X2=1.68 $Y2=3.33
r207 60 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.715 $Y=3.33
+ $X2=1.88 $Y2=3.33
r208 59 78 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=2.045 $Y=3.33
+ $X2=2.16 $Y2=3.33
r209 59 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.045 $Y=3.33
+ $X2=1.88 $Y2=3.33
r210 55 58 22.3574 $w=2.48e-07 $l=4.85e-07 $layer=LI1_cond $X=13.17 $Y=1.98
+ $X2=13.17 $Y2=2.465
r211 53 129 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=13.17 $Y=3.245
+ $X2=13.17 $Y2=3.33
r212 53 58 35.9562 $w=2.48e-07 $l=7.8e-07 $layer=LI1_cond $X=13.17 $Y=3.245
+ $X2=13.17 $Y2=2.465
r213 49 126 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=11.73 $Y=3.245
+ $X2=11.73 $Y2=3.33
r214 49 51 16.4136 $w=3.28e-07 $l=4.7e-07 $layer=LI1_cond $X=11.73 $Y=3.245
+ $X2=11.73 $Y2=2.775
r215 45 67 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.68 $Y=3.245
+ $X2=10.68 $Y2=3.33
r216 45 47 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=10.68 $Y=3.245
+ $X2=10.68 $Y2=2.835
r217 41 123 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.38 $Y=3.245
+ $X2=9.38 $Y2=3.33
r218 41 43 13.969 $w=3.28e-07 $l=4e-07 $layer=LI1_cond $X=9.38 $Y=3.245 $X2=9.38
+ $Y2=2.845
r219 37 120 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.89 $Y=3.245
+ $X2=6.89 $Y2=3.33
r220 37 39 42.0816 $w=3.28e-07 $l=1.205e-06 $layer=LI1_cond $X=6.89 $Y=3.245
+ $X2=6.89 $Y2=2.04
r221 33 64 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.77 $Y=3.245
+ $X2=4.77 $Y2=3.33
r222 33 35 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=4.77 $Y=3.245
+ $X2=4.77 $Y2=2.825
r223 29 61 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.88 $Y=3.245
+ $X2=1.88 $Y2=3.33
r224 29 31 29.8588 $w=3.28e-07 $l=8.55e-07 $layer=LI1_cond $X=1.88 $Y=3.245
+ $X2=1.88 $Y2=2.39
r225 25 117 3.03433 $w=3.3e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.222 $Y2=3.33
r226 25 27 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.28 $Y2=2.55
r227 8 58 300 $w=1.7e-07 $l=7.31779e-07 $layer=licon1_PDIFF $count=2 $X=12.99
+ $Y=1.835 $X2=13.21 $Y2=2.465
r228 8 55 600 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_PDIFF $count=1 $X=12.99
+ $Y=1.835 $X2=13.21 $Y2=1.98
r229 7 51 600 $w=1.7e-07 $l=1.16254e-06 $layer=licon1_PDIFF $count=1 $X=11.515
+ $Y=1.715 $X2=11.73 $Y2=2.775
r230 6 47 600 $w=1.7e-07 $l=6.4622e-07 $layer=licon1_PDIFF $count=1 $X=10.54
+ $Y=2.255 $X2=10.68 $Y2=2.835
r231 5 43 600 $w=1.7e-07 $l=4.60977e-07 $layer=licon1_PDIFF $count=1 $X=9.04
+ $Y=2.56 $X2=9.38 $Y2=2.845
r232 4 39 300 $w=1.7e-07 $l=4.2638e-07 $layer=licon1_PDIFF $count=2 $X=6.53
+ $Y=1.895 $X2=6.89 $Y2=2.04
r233 3 35 600 $w=1.7e-07 $l=1.09733e-06 $layer=licon1_PDIFF $count=1 $X=3.925
+ $Y=2.245 $X2=4.77 $Y2=2.825
r234 2 31 300 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_PDIFF $count=2 $X=1.66
+ $Y=2.245 $X2=1.88 $Y2=2.39
r235 1 27 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.405 $X2=0.28 $Y2=2.55
.ends

.subckt PM_SKY130_FD_SC_LP__DFBBN_1%A_460_449# 1 2 9 12 14 17
c43 12 0 1.40426e-19 $X=2.815 $Y=2.305
r44 16 17 8.63679 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=2.655 $Y=1.13
+ $X2=2.655 $Y2=1.3
r45 12 14 16.3393 $w=2.8e-07 $l=4.60299e-07 $layer=LI1_cond $X=2.815 $Y=2.305
+ $X2=2.44 $Y2=2.495
r46 12 17 65.5668 $w=1.68e-07 $l=1.005e-06 $layer=LI1_cond $X=2.815 $Y=2.305
+ $X2=2.815 $Y2=1.3
r47 9 16 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=2.575 $Y=0.805
+ $X2=2.575 $Y2=1.13
r48 2 14 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=2.3
+ $Y=2.245 $X2=2.44 $Y2=2.455
r49 1 9 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.435
+ $Y=0.595 $X2=2.575 $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_LP__DFBBN_1%Q_N 1 2 9 13 16 17 18 19 20
c35 9 0 1.37465e-19 $X=12.14 $Y=0.43
r36 19 20 11.8446 $w=3.58e-07 $l=3.7e-07 $layer=LI1_cond $X=12.255 $Y=2.405
+ $X2=12.255 $Y2=2.775
r37 18 19 11.8446 $w=3.58e-07 $l=3.7e-07 $layer=LI1_cond $X=12.255 $Y=2.035
+ $X2=12.255 $Y2=2.405
r38 16 17 8.51103 $w=3.58e-07 $l=1.65e-07 $layer=LI1_cond $X=12.255 $Y=1.86
+ $X2=12.255 $Y2=1.695
r39 14 18 5.12197 $w=3.58e-07 $l=1.6e-07 $layer=LI1_cond $X=12.255 $Y=1.875
+ $X2=12.255 $Y2=2.035
r40 14 16 0.480185 $w=3.58e-07 $l=1.5e-08 $layer=LI1_cond $X=12.255 $Y=1.875
+ $X2=12.255 $Y2=1.86
r41 13 17 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=12.35 $Y=1.005
+ $X2=12.35 $Y2=1.695
r42 7 13 10.9702 $w=4.58e-07 $l=2.3e-07 $layer=LI1_cond $X=12.205 $Y=0.775
+ $X2=12.205 $Y2=1.005
r43 7 9 8.97059 $w=4.58e-07 $l=3.45e-07 $layer=LI1_cond $X=12.205 $Y=0.775
+ $X2=12.205 $Y2=0.43
r44 2 20 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=12.02
+ $Y=1.715 $X2=12.16 $Y2=2.83
r45 2 16 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=12.02
+ $Y=1.715 $X2=12.16 $Y2=1.86
r46 1 9 91 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_NDIFF $count=2 $X=12 $Y=0.235
+ $X2=12.14 $Y2=0.43
.ends

.subckt PM_SKY130_FD_SC_LP__DFBBN_1%Q 1 2 9 14 15 16 17 23 29
r23 21 29 0.746653 $w=3.53e-07 $l=2.3e-08 $layer=LI1_cond $X=13.652 $Y=0.948
+ $X2=13.652 $Y2=0.925
r24 17 31 7.88226 $w=3.53e-07 $l=1.46e-07 $layer=LI1_cond $X=13.652 $Y=0.979
+ $X2=13.652 $Y2=1.125
r25 17 21 1.00636 $w=3.53e-07 $l=3.1e-08 $layer=LI1_cond $X=13.652 $Y=0.979
+ $X2=13.652 $Y2=0.948
r26 17 29 1.00636 $w=3.53e-07 $l=3.1e-08 $layer=LI1_cond $X=13.652 $Y=0.894
+ $X2=13.652 $Y2=0.925
r27 16 17 11.005 $w=3.53e-07 $l=3.39e-07 $layer=LI1_cond $X=13.652 $Y=0.555
+ $X2=13.652 $Y2=0.894
r28 16 23 4.0579 $w=3.53e-07 $l=1.25e-07 $layer=LI1_cond $X=13.652 $Y=0.555
+ $X2=13.652 $Y2=0.43
r29 15 31 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=13.745 $Y=1.815
+ $X2=13.745 $Y2=1.125
r30 14 15 8.49906 $w=3.53e-07 $l=1.65e-07 $layer=LI1_cond $X=13.652 $Y=1.98
+ $X2=13.652 $Y2=1.815
r31 7 14 0.389558 $w=3.53e-07 $l=1.2e-08 $layer=LI1_cond $X=13.652 $Y=1.992
+ $X2=13.652 $Y2=1.98
r32 7 9 29.4766 $w=3.53e-07 $l=9.08e-07 $layer=LI1_cond $X=13.652 $Y=1.992
+ $X2=13.652 $Y2=2.9
r33 2 14 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=13.5
+ $Y=1.835 $X2=13.64 $Y2=1.98
r34 2 9 400 $w=1.7e-07 $l=1.13284e-06 $layer=licon1_PDIFF $count=1 $X=13.5
+ $Y=1.835 $X2=13.64 $Y2=2.9
r35 1 23 91 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=2 $X=13.5
+ $Y=0.265 $X2=13.64 $Y2=0.43
.ends

.subckt PM_SKY130_FD_SC_LP__DFBBN_1%VGND 1 2 3 4 5 6 7 22 24 28 32 36 40 44 50
+ 55 56 58 59 60 62 74 88 95 102 103 109 112 115 118
r129 118 119 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.2 $Y=0
+ $X2=13.2 $Y2=0
r130 115 116 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=11.76 $Y=0
+ $X2=11.76 $Y2=0
r131 109 110 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0
+ $X2=1.68 $Y2=0
r132 106 107 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0
+ $X2=0.24 $Y2=0
r133 103 119 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.68 $Y=0
+ $X2=13.2 $Y2=0
r134 102 103 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.68 $Y=0
+ $X2=13.68 $Y2=0
r135 100 118 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=13.295 $Y=0
+ $X2=13.17 $Y2=0
r136 100 102 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=13.295 $Y=0
+ $X2=13.68 $Y2=0
r137 99 119 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.72 $Y=0
+ $X2=13.2 $Y2=0
r138 99 116 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=12.72 $Y=0
+ $X2=11.76 $Y2=0
r139 98 99 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=12.72 $Y=0
+ $X2=12.72 $Y2=0
r140 96 115 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=11.795 $Y=0
+ $X2=11.67 $Y2=0
r141 96 98 60.3476 $w=1.68e-07 $l=9.25e-07 $layer=LI1_cond $X=11.795 $Y=0
+ $X2=12.72 $Y2=0
r142 95 118 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=13.045 $Y=0
+ $X2=13.17 $Y2=0
r143 95 98 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=13.045 $Y=0
+ $X2=12.72 $Y2=0
r144 94 116 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=0
+ $X2=11.76 $Y2=0
r145 93 94 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=11.28 $Y=0
+ $X2=11.28 $Y2=0
r146 91 94 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=9.36 $Y=0
+ $X2=11.28 $Y2=0
r147 90 93 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=9.36 $Y=0
+ $X2=11.28 $Y2=0
r148 90 91 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=9.36 $Y=0
+ $X2=9.36 $Y2=0
r149 88 115 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=11.545 $Y=0
+ $X2=11.67 $Y2=0
r150 88 93 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=11.545 $Y=0
+ $X2=11.28 $Y2=0
r151 87 91 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=0 $X2=9.36
+ $Y2=0
r152 86 87 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.88 $Y=0 $X2=8.88
+ $Y2=0
r153 84 87 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=7.44 $Y=0
+ $X2=8.88 $Y2=0
r154 83 86 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=7.44 $Y=0 $X2=8.88
+ $Y2=0
r155 83 84 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r156 81 112 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.085 $Y=0
+ $X2=6.96 $Y2=0
r157 81 83 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=7.085 $Y=0
+ $X2=7.44 $Y2=0
r158 79 80 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.48 $Y=0
+ $X2=6.48 $Y2=0
r159 77 80 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=4.56 $Y=0
+ $X2=6.48 $Y2=0
r160 76 79 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=4.56 $Y=0 $X2=6.48
+ $Y2=0
r161 76 77 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.56 $Y=0
+ $X2=4.56 $Y2=0
r162 74 112 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.835 $Y=0
+ $X2=6.96 $Y2=0
r163 74 79 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=6.835 $Y=0
+ $X2=6.48 $Y2=0
r164 73 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=4.56
+ $Y2=0
r165 72 73 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.08 $Y=0
+ $X2=4.08 $Y2=0
r166 70 73 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=2.16 $Y=0
+ $X2=4.08 $Y2=0
r167 70 110 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0
+ $X2=1.68 $Y2=0
r168 69 72 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=2.16 $Y=0 $X2=4.08
+ $Y2=0
r169 69 70 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.16 $Y=0
+ $X2=2.16 $Y2=0
r170 67 109 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.925 $Y=0
+ $X2=1.76 $Y2=0
r171 67 69 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=1.925 $Y=0
+ $X2=2.16 $Y2=0
r172 66 110 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r173 66 107 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.24
+ $Y2=0
r174 65 66 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r175 63 106 4.01803 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=0.36 $Y=0 $X2=0.18
+ $Y2=0
r176 63 65 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=0.36 $Y=0 $X2=1.2
+ $Y2=0
r177 62 109 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.595 $Y=0
+ $X2=1.76 $Y2=0
r178 62 65 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=1.595 $Y=0 $X2=1.2
+ $Y2=0
r179 60 84 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=7.44
+ $Y2=0
r180 60 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=6.48
+ $Y2=0
r181 60 112 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r182 58 86 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=8.945 $Y=0 $X2=8.88
+ $Y2=0
r183 58 59 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.945 $Y=0 $X2=9.11
+ $Y2=0
r184 57 90 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=9.275 $Y=0 $X2=9.36
+ $Y2=0
r185 57 59 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.275 $Y=0 $X2=9.11
+ $Y2=0
r186 55 72 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=4.18 $Y=0 $X2=4.08
+ $Y2=0
r187 55 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.18 $Y=0 $X2=4.345
+ $Y2=0
r188 54 76 3.26203 $w=1.68e-07 $l=5e-08 $layer=LI1_cond $X=4.51 $Y=0 $X2=4.56
+ $Y2=0
r189 54 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.51 $Y=0 $X2=4.345
+ $Y2=0
r190 50 52 25.3537 $w=2.48e-07 $l=5.5e-07 $layer=LI1_cond $X=13.17 $Y=0.41
+ $X2=13.17 $Y2=0.96
r191 48 118 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=13.17 $Y=0.085
+ $X2=13.17 $Y2=0
r192 48 50 14.9818 $w=2.48e-07 $l=3.25e-07 $layer=LI1_cond $X=13.17 $Y=0.085
+ $X2=13.17 $Y2=0.41
r193 44 46 20.9745 $w=2.48e-07 $l=4.55e-07 $layer=LI1_cond $X=11.67 $Y=0.38
+ $X2=11.67 $Y2=0.835
r194 42 115 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=11.67 $Y=0.085
+ $X2=11.67 $Y2=0
r195 42 44 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=11.67 $Y=0.085
+ $X2=11.67 $Y2=0.38
r196 38 59 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.11 $Y=0.085
+ $X2=9.11 $Y2=0
r197 38 40 23.9219 $w=3.28e-07 $l=6.85e-07 $layer=LI1_cond $X=9.11 $Y=0.085
+ $X2=9.11 $Y2=0.77
r198 34 112 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.96 $Y=0.085
+ $X2=6.96 $Y2=0
r199 34 36 30.194 $w=2.48e-07 $l=6.55e-07 $layer=LI1_cond $X=6.96 $Y=0.085
+ $X2=6.96 $Y2=0.74
r200 30 56 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.345 $Y=0.085
+ $X2=4.345 $Y2=0
r201 30 32 17.6359 $w=3.28e-07 $l=5.05e-07 $layer=LI1_cond $X=4.345 $Y=0.085
+ $X2=4.345 $Y2=0.59
r202 26 109 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.76 $Y=0.085
+ $X2=1.76 $Y2=0
r203 26 28 24.4458 $w=3.28e-07 $l=7e-07 $layer=LI1_cond $X=1.76 $Y=0.085
+ $X2=1.76 $Y2=0.785
r204 22 106 3.12513 $w=2.5e-07 $l=1.09087e-07 $layer=LI1_cond $X=0.235 $Y=0.085
+ $X2=0.18 $Y2=0
r205 22 24 21.205 $w=2.48e-07 $l=4.6e-07 $layer=LI1_cond $X=0.235 $Y=0.085
+ $X2=0.235 $Y2=0.545
r206 7 52 182 $w=1.7e-07 $l=3.68951e-07 $layer=licon1_NDIFF $count=1 $X=12.99
+ $Y=0.685 $X2=13.21 $Y2=0.96
r207 7 50 182 $w=1.7e-07 $l=3.68951e-07 $layer=licon1_NDIFF $count=1 $X=12.99
+ $Y=0.685 $X2=13.21 $Y2=0.41
r208 6 46 182 $w=1.7e-07 $l=2.96648e-07 $layer=licon1_NDIFF $count=1 $X=11.49
+ $Y=0.655 $X2=11.71 $Y2=0.835
r209 6 44 182 $w=1.7e-07 $l=3.68951e-07 $layer=licon1_NDIFF $count=1 $X=11.49
+ $Y=0.655 $X2=11.71 $Y2=0.38
r210 5 40 182 $w=1.7e-07 $l=2.76586e-07 $layer=licon1_NDIFF $count=1 $X=8.855
+ $Y=0.815 $X2=9.11 $Y2=0.77
r211 4 36 182 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=1 $X=6.775
+ $Y=0.595 $X2=6.92 $Y2=0.74
r212 3 32 182 $w=1.7e-07 $l=2.84297e-07 $layer=licon1_NDIFF $count=1 $X=4.08
+ $Y=0.55 $X2=4.345 $Y2=0.59
r213 2 28 182 $w=1.7e-07 $l=3.00333e-07 $layer=licon1_NDIFF $count=1 $X=1.54
+ $Y=0.595 $X2=1.76 $Y2=0.785
r214 1 24 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.335 $X2=0.275 $Y2=0.545
.ends

.subckt PM_SKY130_FD_SC_LP__DFBBN_1%A_1013_66# 1 2 7 12 15
r24 10 12 8.55446 $w=3.73e-07 $l=1.65e-07 $layer=LI1_cond $X=5.205 $Y=0.802
+ $X2=5.37 $Y2=0.802
r25 7 15 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.135 $Y=0.7 $X2=6.22
+ $Y2=0.7
r26 7 12 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=6.135 $Y=0.7
+ $X2=5.37 $Y2=0.7
r27 2 15 182 $w=1.7e-07 $l=5.15267e-07 $layer=licon1_NDIFF $count=1 $X=6.08
+ $Y=0.33 $X2=6.22 $Y2=0.78
r28 1 10 182 $w=1.7e-07 $l=4.95076e-07 $layer=licon1_NDIFF $count=1 $X=5.065
+ $Y=0.33 $X2=5.205 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_LP__DFBBN_1%A_1896_119# 1 2 9 11 12 13
r30 13 16 6.80989 $w=3.28e-07 $l=1.95e-07 $layer=LI1_cond $X=10.64 $Y=0.35
+ $X2=10.64 $Y2=0.545
r31 11 13 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.475 $Y=0.35
+ $X2=10.64 $Y2=0.35
r32 11 12 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=10.475 $Y=0.35
+ $X2=9.785 $Y2=0.35
r33 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=9.62 $Y=0.435
+ $X2=9.785 $Y2=0.35
r34 7 9 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=9.62 $Y=0.435 $X2=9.62
+ $Y2=0.77
r35 2 16 182 $w=1.7e-07 $l=2.63106e-07 $layer=licon1_NDIFF $count=1 $X=10.445
+ $Y=0.385 $X2=10.64 $Y2=0.545
r36 1 9 182 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=1 $X=9.48
+ $Y=0.595 $X2=9.62 $Y2=0.77
.ends

