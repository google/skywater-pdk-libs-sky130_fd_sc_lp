* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__maj3_lp A B C VGND VNB VPB VPWR X
M1000 a_154_125# B a_29_419# VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=3.20775e+11p ps=3.54e+06u
M1001 VGND C a_530_68# VNB nshort w=420000u l=150000u
+  ad=3.8505e+11p pd=3.69e+06u as=1.302e+11p ps=1.46e+06u
M1002 a_548_419# B a_29_419# VPB phighvt w=1e+06u l=250000u
+  ad=2.5e+11p pd=2.5e+06u as=6.45e+11p ps=5.29e+06u
M1003 X a_29_419# VPWR VPB phighvt w=1e+06u l=250000u
+  ad=2.85e+11p pd=2.57e+06u as=5.7e+11p ps=5.14e+06u
M1004 a_152_419# B a_29_419# VPB phighvt w=1e+06u l=250000u
+  ad=2.1e+11p pd=2.42e+06u as=0p ps=0u
M1005 VPWR C a_548_419# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_29_419# C a_350_125# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1007 X a_29_419# a_708_68# VNB nshort w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=8.82e+10p ps=1.26e+06u
M1008 a_29_419# C a_350_419# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=2.1e+11p ps=2.42e+06u
M1009 a_708_68# a_29_419# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND A a_154_125# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_530_68# B a_29_419# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_350_419# A VPWR VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VPWR A a_152_419# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_350_125# A VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
