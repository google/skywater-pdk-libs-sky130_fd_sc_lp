# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__and2_4
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__and2_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.360000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.315000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.325000 0.455000 1.750000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.315000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.635000 1.325000 1.020000 1.750000 ;
    END
  END B
  PIN X
    ANTENNADIFFAREA  1.176000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.530000 0.255000 1.720000 1.065000 ;
        RECT 1.530000 1.065000 3.260000 1.235000 ;
        RECT 1.530000 1.775000 3.260000 1.945000 ;
        RECT 1.530000 1.945000 1.720000 3.075000 ;
        RECT 2.390000 0.255000 2.580000 1.065000 ;
        RECT 2.390000 1.945000 2.580000 3.075000 ;
        RECT 2.855000 1.235000 3.260000 1.775000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.360000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.360000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.360000 0.085000 ;
      RECT 0.000000  3.245000 3.360000 3.415000 ;
      RECT 0.095000  0.255000 0.425000 0.985000 ;
      RECT 0.095000  0.985000 1.360000 1.155000 ;
      RECT 0.095000  1.920000 0.425000 3.245000 ;
      RECT 0.595000  1.930000 1.360000 2.100000 ;
      RECT 0.595000  2.100000 0.785000 3.075000 ;
      RECT 0.955000  0.085000 1.285000 0.815000 ;
      RECT 0.990000  2.270000 1.320000 3.245000 ;
      RECT 1.190000  1.155000 1.360000 1.405000 ;
      RECT 1.190000  1.405000 2.685000 1.605000 ;
      RECT 1.190000  1.605000 1.360000 1.930000 ;
      RECT 1.890000  0.085000 2.220000 0.885000 ;
      RECT 1.890000  2.115000 2.220000 3.245000 ;
      RECT 2.750000  0.085000 3.080000 0.885000 ;
      RECT 2.750000  2.115000 3.080000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
  END
END sky130_fd_sc_lp__and2_4
END LIBRARY
