* File: sky130_fd_sc_lp__a22oi_1.spice
* Created: Wed Sep  2 09:23:05 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__a22oi_1.pex.spice"
.subckt sky130_fd_sc_lp__a22oi_1  VNB VPB B2 B1 A1 A2 Y VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Y	Y
* A2	A2
* A1	A1
* B1	B1
* B2	B2
* VPB	VPB
* VNB	VNB
MM1004 A_148_69# N_B2_M1004_g N_VGND_M1004_s VNB NSHORT L=0.15 W=0.84 AD=0.0882
+ AS=0.2226 PD=1.05 PS=2.21 NRD=7.14 NRS=0 M=1 R=5.6 SA=75000.2 SB=75001.6
+ A=0.126 P=1.98 MULT=1
MM1007 N_Y_M1007_d N_B1_M1007_g A_148_69# VNB NSHORT L=0.15 W=0.84 AD=0.1701
+ AS=0.0882 PD=1.245 PS=1.05 NRD=12.852 NRS=7.14 M=1 R=5.6 SA=75000.6 SB=75001.3
+ A=0.126 P=1.98 MULT=1
MM1005 A_331_69# N_A1_M1005_g N_Y_M1007_d VNB NSHORT L=0.15 W=0.84 AD=0.1638
+ AS=0.1701 PD=1.23 PS=1.245 NRD=19.992 NRS=4.992 M=1 R=5.6 SA=75001.1
+ SB=75000.7 A=0.126 P=1.98 MULT=1
MM1001 N_VGND_M1001_d N_A2_M1001_g A_331_69# VNB NSHORT L=0.15 W=0.84 AD=0.2226
+ AS=0.1638 PD=2.21 PS=1.23 NRD=0 NRS=19.992 M=1 R=5.6 SA=75001.6 SB=75000.2
+ A=0.126 P=1.98 MULT=1
MM1002 N_Y_M1002_d N_B2_M1002_g N_A_65_367#_M1002_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75001.9 A=0.189 P=2.82 MULT=1
MM1006 N_A_65_367#_M1006_d N_B1_M1006_g N_Y_M1002_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.21105 AS=0.1764 PD=1.595 PS=1.54 NRD=4.6886 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75001.4 A=0.189 P=2.82 MULT=1
MM1003 N_VPWR_M1003_d N_A1_M1003_g N_A_65_367#_M1006_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3906 AS=0.21105 PD=1.88 PS=1.595 NRD=0 NRS=3.9006 M=1 R=8.4 SA=75001.1
+ SB=75001 A=0.189 P=2.82 MULT=1
MM1000 N_A_65_367#_M1000_d N_A2_M1000_g N_VPWR_M1003_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.3906 PD=3.05 PS=1.88 NRD=0 NRS=0 M=1 R=8.4 SA=75001.9
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX8_noxref VNB VPB NWDIODE A=6.0799 P=10.25
*
.include "sky130_fd_sc_lp__a22oi_1.pxi.spice"
*
.ends
*
*
