* File: sky130_fd_sc_lp__buflp_0.pex.spice
* Created: Fri Aug 28 10:12:08 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__BUFLP_0%A 3 7 11 15 17 18 19 20 26
r40 26 27 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.77
+ $Y=1.765 $X2=0.77 $Y2=1.765
r41 19 20 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.77 $Y=2.405
+ $X2=0.77 $Y2=2.775
r42 18 19 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.77 $Y=2.035
+ $X2=0.77 $Y2=2.405
r43 18 27 9.42908 $w=3.28e-07 $l=2.7e-07 $layer=LI1_cond $X=0.77 $Y=2.035
+ $X2=0.77 $Y2=1.765
r44 17 27 3.49225 $w=3.28e-07 $l=1e-07 $layer=LI1_cond $X=0.77 $Y=1.665 $X2=0.77
+ $Y2=1.765
r45 13 26 91.6154 $w=2.72e-07 $l=6.00054e-07 $layer=POLY_cond $X=0.955 $Y=2.27
+ $X2=0.747 $Y2=1.765
r46 13 15 199.979 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=0.955 $Y=2.27
+ $X2=0.955 $Y2=2.66
r47 9 26 31.3654 $w=2.72e-07 $l=2.52357e-07 $layer=POLY_cond $X=0.93 $Y=1.6
+ $X2=0.747 $Y2=1.765
r48 9 11 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=0.93 $Y=1.6 $X2=0.93
+ $Y2=0.81
r49 5 26 91.6154 $w=2.72e-07 $l=5.89012e-07 $layer=POLY_cond $X=0.565 $Y=2.27
+ $X2=0.747 $Y2=1.765
r50 5 7 199.979 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=0.565 $Y=2.27
+ $X2=0.565 $Y2=2.66
r51 1 26 31.3654 $w=2.72e-07 $l=2.77496e-07 $layer=POLY_cond $X=0.54 $Y=1.6
+ $X2=0.747 $Y2=1.765
r52 1 3 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=0.54 $Y=1.6 $X2=0.54
+ $Y2=0.81
.ends

.subckt PM_SKY130_FD_SC_LP__BUFLP_0%A_36_120# 1 2 9 13 17 21 28 31 34 38 40 44
+ 46 47
r62 46 47 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.41
+ $Y=1.375 $X2=1.41 $Y2=1.375
r63 41 44 3.47949 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.49 $Y=1.295
+ $X2=0.325 $Y2=1.295
r64 40 46 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.245 $Y=1.295
+ $X2=1.41 $Y2=1.295
r65 40 41 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=1.245 $Y=1.295
+ $X2=0.49 $Y2=1.295
r66 36 44 3.12539 $w=3.02e-07 $l=9.80051e-08 $layer=LI1_cond $X=0.297 $Y=1.38
+ $X2=0.325 $Y2=1.295
r67 36 38 53.641 $w=2.73e-07 $l=1.28e-06 $layer=LI1_cond $X=0.297 $Y=1.38
+ $X2=0.297 $Y2=2.66
r68 32 44 3.12539 $w=3.02e-07 $l=8.5e-08 $layer=LI1_cond $X=0.325 $Y=1.21
+ $X2=0.325 $Y2=1.295
r69 32 34 13.969 $w=3.28e-07 $l=4e-07 $layer=LI1_cond $X=0.325 $Y=1.21 $X2=0.325
+ $Y2=0.81
r70 30 47 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.41 $Y=1.715
+ $X2=1.41 $Y2=1.375
r71 30 31 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.41 $Y=1.715
+ $X2=1.41 $Y2=1.88
r72 27 28 71.7872 $w=1.5e-07 $l=1.4e-07 $layer=POLY_cond $X=1.75 $Y=1.285
+ $X2=1.89 $Y2=1.285
r73 26 47 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=1.41 $Y=1.36
+ $X2=1.41 $Y2=1.375
r74 26 27 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=1.41 $Y=1.285
+ $X2=1.75 $Y2=1.285
r75 23 26 25.6383 $w=1.5e-07 $l=5e-08 $layer=POLY_cond $X=1.36 $Y=1.285 $X2=1.41
+ $Y2=1.285
r76 19 28 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.89 $Y=1.36
+ $X2=1.89 $Y2=1.285
r77 19 21 610.191 $w=1.5e-07 $l=1.19e-06 $layer=POLY_cond $X=1.89 $Y=1.36
+ $X2=1.89 $Y2=2.55
r78 15 27 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.75 $Y=1.21
+ $X2=1.75 $Y2=1.285
r79 15 17 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=1.75 $Y=1.21 $X2=1.75
+ $Y2=0.81
r80 13 31 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=1.5 $Y=2.55 $X2=1.5
+ $Y2=1.88
r81 7 23 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.36 $Y=1.21 $X2=1.36
+ $Y2=1.285
r82 7 9 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=1.36 $Y=1.21 $X2=1.36
+ $Y2=0.81
r83 2 38 600 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=1 $X=0.205
+ $Y=2.45 $X2=0.35 $Y2=2.66
r84 1 34 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.18
+ $Y=0.6 $X2=0.325 $Y2=0.81
.ends

.subckt PM_SKY130_FD_SC_LP__BUFLP_0%VPWR 1 6 8 10 17 18 21
r27 17 18 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r28 15 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.45 $Y=3.33
+ $X2=1.285 $Y2=3.33
r29 15 17 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=1.45 $Y=3.33
+ $X2=2.16 $Y2=3.33
r30 12 13 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r31 10 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.12 $Y=3.33
+ $X2=1.285 $Y2=3.33
r32 10 12 57.4118 $w=1.68e-07 $l=8.8e-07 $layer=LI1_cond $X=1.12 $Y=3.33
+ $X2=0.24 $Y2=3.33
r33 8 18 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33 $X2=2.16
+ $Y2=3.33
r34 8 13 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33 $X2=0.24
+ $Y2=3.33
r35 8 21 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r36 4 21 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.285 $Y=3.245
+ $X2=1.285 $Y2=3.33
r37 4 6 30.3826 $w=3.28e-07 $l=8.7e-07 $layer=LI1_cond $X=1.285 $Y=3.245
+ $X2=1.285 $Y2=2.375
r38 1 6 300 $w=1.7e-07 $l=2.90086e-07 $layer=licon1_PDIFF $count=2 $X=1.03
+ $Y=2.45 $X2=1.285 $Y2=2.375
.ends

.subckt PM_SKY130_FD_SC_LP__BUFLP_0%X 1 2 7 8 9 10 11 12 13
r14 12 13 10.0722 $w=4.73e-07 $l=4e-07 $layer=LI1_cond $X=2.037 $Y=2.375
+ $X2=2.037 $Y2=2.775
r15 11 12 8.5614 $w=4.73e-07 $l=3.4e-07 $layer=LI1_cond $X=2.037 $Y=2.035
+ $X2=2.037 $Y2=2.375
r16 10 11 9.31682 $w=4.73e-07 $l=3.7e-07 $layer=LI1_cond $X=2.037 $Y=1.665
+ $X2=2.037 $Y2=2.035
r17 9 10 9.31682 $w=4.73e-07 $l=3.7e-07 $layer=LI1_cond $X=2.037 $Y=1.295
+ $X2=2.037 $Y2=1.665
r18 8 9 9.31682 $w=4.73e-07 $l=3.7e-07 $layer=LI1_cond $X=2.037 $Y=0.925
+ $X2=2.037 $Y2=1.295
r19 8 25 2.89577 $w=4.73e-07 $l=1.15e-07 $layer=LI1_cond $X=2.037 $Y=0.925
+ $X2=2.037 $Y2=0.81
r20 7 25 6.42105 $w=4.73e-07 $l=2.55e-07 $layer=LI1_cond $X=2.037 $Y=0.555
+ $X2=2.037 $Y2=0.81
r21 2 12 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=1.965
+ $Y=2.23 $X2=2.105 $Y2=2.375
r22 1 25 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.825
+ $Y=0.6 $X2=1.965 $Y2=0.81
.ends

.subckt PM_SKY130_FD_SC_LP__BUFLP_0%VGND 1 6 8 10 17 18 21
r26 17 18 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r27 15 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.31 $Y=0 $X2=1.145
+ $Y2=0
r28 15 17 55.4545 $w=1.68e-07 $l=8.5e-07 $layer=LI1_cond $X=1.31 $Y=0 $X2=2.16
+ $Y2=0
r29 12 13 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r30 10 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.98 $Y=0 $X2=1.145
+ $Y2=0
r31 10 12 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=0.98 $Y=0 $X2=0.72
+ $Y2=0
r32 8 18 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r33 8 13 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r34 8 21 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r35 4 21 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.145 $Y=0.085
+ $X2=1.145 $Y2=0
r36 4 6 25.3188 $w=3.28e-07 $l=7.25e-07 $layer=LI1_cond $X=1.145 $Y=0.085
+ $X2=1.145 $Y2=0.81
r37 1 6 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.005
+ $Y=0.6 $X2=1.145 $Y2=0.81
.ends

