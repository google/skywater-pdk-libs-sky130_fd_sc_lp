* File: sky130_fd_sc_lp__clkbuf_8.pex.spice
* Created: Wed Sep  2 09:38:39 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__CLKBUF_8%A 3 7 11 15 17 18 26
r39 25 26 34.3377 $w=6.7e-07 $l=4.3e-07 $layer=POLY_cond $X=0.475 $Y=1.235
+ $X2=0.905 $Y2=1.235
r40 22 25 16.3703 $w=6.7e-07 $l=2.05e-07 $layer=POLY_cond $X=0.27 $Y=1.235
+ $X2=0.475 $Y2=1.235
r41 22 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.27
+ $Y=1.065 $X2=0.27 $Y2=1.065
r42 18 23 8.41466 $w=3.13e-07 $l=2.3e-07 $layer=LI1_cond $X=0.242 $Y=1.295
+ $X2=0.242 $Y2=1.065
r43 17 23 5.12197 $w=3.13e-07 $l=1.4e-07 $layer=LI1_cond $X=0.242 $Y=0.925
+ $X2=0.242 $Y2=1.065
r44 13 26 38.9565 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=0.905 $Y=1.57
+ $X2=0.905 $Y2=1.235
r45 13 15 458.926 $w=1.5e-07 $l=8.95e-07 $layer=POLY_cond $X=0.905 $Y=1.57
+ $X2=0.905 $Y2=2.465
r46 9 26 38.9565 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=0.905 $Y=0.9
+ $X2=0.905 $Y2=1.235
r47 9 11 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=0.905 $Y=0.9
+ $X2=0.905 $Y2=0.445
r48 5 25 38.9565 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=0.475 $Y=1.57
+ $X2=0.475 $Y2=1.235
r49 5 7 458.926 $w=1.5e-07 $l=8.95e-07 $layer=POLY_cond $X=0.475 $Y=1.57
+ $X2=0.475 $Y2=2.465
r50 1 25 38.9565 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=0.475 $Y=0.9
+ $X2=0.475 $Y2=1.235
r51 1 3 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=0.475 $Y=0.9
+ $X2=0.475 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__CLKBUF_8%A_110_47# 1 2 9 13 17 21 25 29 33 37 41 45
+ 49 53 57 61 65 69 73 77 86 89 100
r156 99 100 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=3.915 $Y=1.32
+ $X2=4.345 $Y2=1.32
r157 98 99 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=3.485 $Y=1.32
+ $X2=3.915 $Y2=1.32
r158 95 96 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=2.625 $Y=1.32
+ $X2=3.055 $Y2=1.32
r159 94 95 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=2.195 $Y=1.32
+ $X2=2.625 $Y2=1.32
r160 93 94 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=1.765 $Y=1.32
+ $X2=2.195 $Y2=1.32
r161 87 98 41.9667 $w=3.3e-07 $l=2.4e-07 $layer=POLY_cond $X=3.245 $Y=1.32
+ $X2=3.485 $Y2=1.32
r162 87 96 33.2236 $w=3.3e-07 $l=1.9e-07 $layer=POLY_cond $X=3.245 $Y=1.32
+ $X2=3.055 $Y2=1.32
r163 86 87 48.4267 $w=1.7e-07 $l=5.1e-07 $layer=licon1_POLY $count=3 $X=3.245
+ $Y=1.32 $X2=3.245 $Y2=1.32
r164 84 93 38.4695 $w=3.3e-07 $l=2.2e-07 $layer=POLY_cond $X=1.545 $Y=1.32
+ $X2=1.765 $Y2=1.32
r165 84 90 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=1.545 $Y=1.32
+ $X2=1.335 $Y2=1.32
r166 83 86 59.3683 $w=3.28e-07 $l=1.7e-06 $layer=LI1_cond $X=1.545 $Y=1.32
+ $X2=3.245 $Y2=1.32
r167 83 84 48.4267 $w=1.7e-07 $l=5.1e-07 $layer=licon1_POLY $count=3 $X=1.545
+ $Y=1.32 $X2=1.545 $Y2=1.32
r168 81 89 0.364692 $w=3.3e-07 $l=1.25e-07 $layer=LI1_cond $X=0.82 $Y=1.32
+ $X2=0.695 $Y2=1.32
r169 81 83 25.3188 $w=3.28e-07 $l=7.25e-07 $layer=LI1_cond $X=0.82 $Y=1.32
+ $X2=1.545 $Y2=1.32
r170 77 79 39.1831 $w=2.48e-07 $l=8.5e-07 $layer=LI1_cond $X=0.695 $Y=2.04
+ $X2=0.695 $Y2=2.89
r171 75 89 6.46576 $w=2.5e-07 $l=1.65e-07 $layer=LI1_cond $X=0.695 $Y=1.485
+ $X2=0.695 $Y2=1.32
r172 75 77 25.5842 $w=2.48e-07 $l=5.55e-07 $layer=LI1_cond $X=0.695 $Y=1.485
+ $X2=0.695 $Y2=2.04
r173 71 89 6.46576 $w=2.5e-07 $l=1.65e-07 $layer=LI1_cond $X=0.695 $Y=1.155
+ $X2=0.695 $Y2=1.32
r174 71 73 32.7294 $w=2.48e-07 $l=7.1e-07 $layer=LI1_cond $X=0.695 $Y=1.155
+ $X2=0.695 $Y2=0.445
r175 67 100 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.345 $Y=1.485
+ $X2=4.345 $Y2=1.32
r176 67 69 502.511 $w=1.5e-07 $l=9.8e-07 $layer=POLY_cond $X=4.345 $Y=1.485
+ $X2=4.345 $Y2=2.465
r177 63 100 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.345 $Y=1.155
+ $X2=4.345 $Y2=1.32
r178 63 65 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=4.345 $Y=1.155
+ $X2=4.345 $Y2=0.445
r179 59 99 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.915 $Y=1.485
+ $X2=3.915 $Y2=1.32
r180 59 61 502.511 $w=1.5e-07 $l=9.8e-07 $layer=POLY_cond $X=3.915 $Y=1.485
+ $X2=3.915 $Y2=2.465
r181 55 99 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.915 $Y=1.155
+ $X2=3.915 $Y2=1.32
r182 55 57 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=3.915 $Y=1.155
+ $X2=3.915 $Y2=0.445
r183 51 98 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.485 $Y=1.485
+ $X2=3.485 $Y2=1.32
r184 51 53 502.511 $w=1.5e-07 $l=9.8e-07 $layer=POLY_cond $X=3.485 $Y=1.485
+ $X2=3.485 $Y2=2.465
r185 47 98 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.485 $Y=1.155
+ $X2=3.485 $Y2=1.32
r186 47 49 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=3.485 $Y=1.155
+ $X2=3.485 $Y2=0.445
r187 43 96 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.055 $Y=1.485
+ $X2=3.055 $Y2=1.32
r188 43 45 502.511 $w=1.5e-07 $l=9.8e-07 $layer=POLY_cond $X=3.055 $Y=1.485
+ $X2=3.055 $Y2=2.465
r189 39 96 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.055 $Y=1.155
+ $X2=3.055 $Y2=1.32
r190 39 41 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=3.055 $Y=1.155
+ $X2=3.055 $Y2=0.445
r191 35 95 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.625 $Y=1.485
+ $X2=2.625 $Y2=1.32
r192 35 37 502.511 $w=1.5e-07 $l=9.8e-07 $layer=POLY_cond $X=2.625 $Y=1.485
+ $X2=2.625 $Y2=2.465
r193 31 95 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.625 $Y=1.155
+ $X2=2.625 $Y2=1.32
r194 31 33 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=2.625 $Y=1.155
+ $X2=2.625 $Y2=0.445
r195 27 94 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.195 $Y=1.485
+ $X2=2.195 $Y2=1.32
r196 27 29 502.511 $w=1.5e-07 $l=9.8e-07 $layer=POLY_cond $X=2.195 $Y=1.485
+ $X2=2.195 $Y2=2.465
r197 23 94 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.195 $Y=1.155
+ $X2=2.195 $Y2=1.32
r198 23 25 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=2.195 $Y=1.155
+ $X2=2.195 $Y2=0.445
r199 19 93 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.765 $Y=1.485
+ $X2=1.765 $Y2=1.32
r200 19 21 502.511 $w=1.5e-07 $l=9.8e-07 $layer=POLY_cond $X=1.765 $Y=1.485
+ $X2=1.765 $Y2=2.465
r201 15 93 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.765 $Y=1.155
+ $X2=1.765 $Y2=1.32
r202 15 17 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=1.765 $Y=1.155
+ $X2=1.765 $Y2=0.445
r203 11 90 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.335 $Y=1.485
+ $X2=1.335 $Y2=1.32
r204 11 13 502.511 $w=1.5e-07 $l=9.8e-07 $layer=POLY_cond $X=1.335 $Y=1.485
+ $X2=1.335 $Y2=2.465
r205 7 90 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.335 $Y=1.155
+ $X2=1.335 $Y2=1.32
r206 7 9 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=1.335 $Y=1.155
+ $X2=1.335 $Y2=0.445
r207 2 79 400 $w=1.7e-07 $l=1.12282e-06 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=1.835 $X2=0.69 $Y2=2.89
r208 2 77 400 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=1.835 $X2=0.69 $Y2=2.04
r209 1 73 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.235 $X2=0.69 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__CLKBUF_8%VPWR 1 2 3 4 5 6 19 21 27 33 39 43 47 53 58
+ 59 61 62 63 64 65 77 84 85 91 94
r78 94 95 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r79 91 92 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r80 88 89 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r81 85 95 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=4.56 $Y2=3.33
r82 84 85 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r83 82 94 7.94884 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=4.725 $Y=3.33
+ $X2=4.577 $Y2=3.33
r84 82 84 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=4.725 $Y=3.33
+ $X2=5.04 $Y2=3.33
r85 81 95 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r86 81 92 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.6 $Y2=3.33
r87 80 81 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r88 78 91 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.83 $Y=3.33 $X2=3.7
+ $Y2=3.33
r89 78 80 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=3.83 $Y=3.33
+ $X2=4.08 $Y2=3.33
r90 77 94 7.94884 $w=1.7e-07 $l=1.47e-07 $layer=LI1_cond $X=4.43 $Y=3.33
+ $X2=4.577 $Y2=3.33
r91 77 80 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=4.43 $Y=3.33
+ $X2=4.08 $Y2=3.33
r92 72 73 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r93 70 73 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r94 70 89 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r95 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r96 67 88 4.45907 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=0.39 $Y=3.33
+ $X2=0.195 $Y2=3.33
r97 67 69 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=0.39 $Y=3.33
+ $X2=0.72 $Y2=3.33
r98 65 92 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r99 65 73 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=1.68 $Y2=3.33
r100 65 75 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r101 63 75 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=2.71 $Y=3.33 $X2=2.64
+ $Y2=3.33
r102 63 64 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.71 $Y=3.33
+ $X2=2.84 $Y2=3.33
r103 61 72 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.85 $Y=3.33
+ $X2=1.68 $Y2=3.33
r104 61 62 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.85 $Y=3.33
+ $X2=1.98 $Y2=3.33
r105 60 75 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=2.11 $Y=3.33
+ $X2=2.64 $Y2=3.33
r106 60 62 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.11 $Y=3.33
+ $X2=1.98 $Y2=3.33
r107 58 69 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=0.99 $Y=3.33
+ $X2=0.72 $Y2=3.33
r108 58 59 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.99 $Y=3.33
+ $X2=1.12 $Y2=3.33
r109 57 72 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=1.25 $Y=3.33
+ $X2=1.68 $Y2=3.33
r110 57 59 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.25 $Y=3.33
+ $X2=1.12 $Y2=3.33
r111 53 56 27.3461 $w=2.93e-07 $l=7e-07 $layer=LI1_cond $X=4.577 $Y=2.23
+ $X2=4.577 $Y2=2.93
r112 51 94 0.543863 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=4.577 $Y=3.245
+ $X2=4.577 $Y2=3.33
r113 51 56 12.3057 $w=2.93e-07 $l=3.15e-07 $layer=LI1_cond $X=4.577 $Y=3.245
+ $X2=4.577 $Y2=2.93
r114 47 50 31.0273 $w=2.58e-07 $l=7e-07 $layer=LI1_cond $X=3.7 $Y=2.23 $X2=3.7
+ $Y2=2.93
r115 45 91 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=3.7 $Y=3.245
+ $X2=3.7 $Y2=3.33
r116 45 50 13.9623 $w=2.58e-07 $l=3.15e-07 $layer=LI1_cond $X=3.7 $Y=3.245
+ $X2=3.7 $Y2=2.93
r117 44 64 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.97 $Y=3.33
+ $X2=2.84 $Y2=3.33
r118 43 91 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.57 $Y=3.33 $X2=3.7
+ $Y2=3.33
r119 43 44 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=3.57 $Y=3.33 $X2=2.97
+ $Y2=3.33
r120 39 42 31.0273 $w=2.58e-07 $l=7e-07 $layer=LI1_cond $X=2.84 $Y=2.23 $X2=2.84
+ $Y2=2.93
r121 37 64 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=2.84 $Y=3.245
+ $X2=2.84 $Y2=3.33
r122 37 42 13.9623 $w=2.58e-07 $l=3.15e-07 $layer=LI1_cond $X=2.84 $Y=3.245
+ $X2=2.84 $Y2=2.93
r123 33 36 31.0273 $w=2.58e-07 $l=7e-07 $layer=LI1_cond $X=1.98 $Y=2.23 $X2=1.98
+ $Y2=2.93
r124 31 62 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=1.98 $Y=3.245
+ $X2=1.98 $Y2=3.33
r125 31 36 13.9623 $w=2.58e-07 $l=3.15e-07 $layer=LI1_cond $X=1.98 $Y=3.245
+ $X2=1.98 $Y2=2.93
r126 27 30 37.676 $w=2.58e-07 $l=8.5e-07 $layer=LI1_cond $X=1.12 $Y=2.04
+ $X2=1.12 $Y2=2.89
r127 25 59 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=1.12 $Y=3.245
+ $X2=1.12 $Y2=3.33
r128 25 30 15.7353 $w=2.58e-07 $l=3.55e-07 $layer=LI1_cond $X=1.12 $Y=3.245
+ $X2=1.12 $Y2=2.89
r129 21 24 33.206 $w=2.93e-07 $l=8.5e-07 $layer=LI1_cond $X=0.242 $Y=2.04
+ $X2=0.242 $Y2=2.89
r130 19 88 3.01845 $w=2.95e-07 $l=1.05924e-07 $layer=LI1_cond $X=0.242 $Y=3.245
+ $X2=0.195 $Y2=3.33
r131 19 24 13.8684 $w=2.93e-07 $l=3.55e-07 $layer=LI1_cond $X=0.242 $Y=3.245
+ $X2=0.242 $Y2=2.89
r132 6 56 400 $w=1.7e-07 $l=1.1629e-06 $layer=licon1_PDIFF $count=1 $X=4.42
+ $Y=1.835 $X2=4.56 $Y2=2.93
r133 6 53 400 $w=1.7e-07 $l=4.59701e-07 $layer=licon1_PDIFF $count=1 $X=4.42
+ $Y=1.835 $X2=4.56 $Y2=2.23
r134 5 50 400 $w=1.7e-07 $l=1.1629e-06 $layer=licon1_PDIFF $count=1 $X=3.56
+ $Y=1.835 $X2=3.7 $Y2=2.93
r135 5 47 400 $w=1.7e-07 $l=4.59701e-07 $layer=licon1_PDIFF $count=1 $X=3.56
+ $Y=1.835 $X2=3.7 $Y2=2.23
r136 4 42 400 $w=1.7e-07 $l=1.1629e-06 $layer=licon1_PDIFF $count=1 $X=2.7
+ $Y=1.835 $X2=2.84 $Y2=2.93
r137 4 39 400 $w=1.7e-07 $l=4.59701e-07 $layer=licon1_PDIFF $count=1 $X=2.7
+ $Y=1.835 $X2=2.84 $Y2=2.23
r138 3 36 400 $w=1.7e-07 $l=1.1629e-06 $layer=licon1_PDIFF $count=1 $X=1.84
+ $Y=1.835 $X2=1.98 $Y2=2.93
r139 3 33 400 $w=1.7e-07 $l=4.59701e-07 $layer=licon1_PDIFF $count=1 $X=1.84
+ $Y=1.835 $X2=1.98 $Y2=2.23
r140 2 30 400 $w=1.7e-07 $l=1.12282e-06 $layer=licon1_PDIFF $count=1 $X=0.98
+ $Y=1.835 $X2=1.12 $Y2=2.89
r141 2 27 400 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=1 $X=0.98
+ $Y=1.835 $X2=1.12 $Y2=2.04
r142 1 24 400 $w=1.7e-07 $l=1.11575e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.835 $X2=0.26 $Y2=2.89
r143 1 21 400 $w=1.7e-07 $l=2.60096e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.835 $X2=0.26 $Y2=2.04
.ends

.subckt PM_SKY130_FD_SC_LP__CLKBUF_8%X 1 2 3 4 5 6 7 8 27 31 35 36 37 38 41 45
+ 49 51 55 59 63 65 69 73 77 78 79 80 81 82 83
r127 83 98 2.23356 $w=6.15e-07 $l=1.2e-07 $layer=LI1_cond $X=4.245 $Y=1.775
+ $X2=4.245 $Y2=1.655
r128 83 98 0.477938 $w=9.68e-07 $l=3.8e-08 $layer=LI1_cond $X=4.245 $Y=1.617
+ $X2=4.245 $Y2=1.655
r129 82 83 4.0499 $w=9.68e-07 $l=3.22e-07 $layer=LI1_cond $X=4.245 $Y=1.295
+ $X2=4.245 $Y2=1.617
r130 81 97 2.23356 $w=6.15e-07 $l=1.2e-07 $layer=LI1_cond $X=4.245 $Y=0.855
+ $X2=4.245 $Y2=0.975
r131 81 82 3.81093 $w=9.68e-07 $l=3.03e-07 $layer=LI1_cond $X=4.245 $Y=0.992
+ $X2=4.245 $Y2=1.295
r132 81 97 0.213814 $w=9.68e-07 $l=1.7e-08 $layer=LI1_cond $X=4.245 $Y=0.992
+ $X2=4.245 $Y2=0.975
r133 73 75 37.676 $w=2.58e-07 $l=8.5e-07 $layer=LI1_cond $X=4.13 $Y=2.04
+ $X2=4.13 $Y2=2.89
r134 71 83 2.23356 $w=6.15e-07 $l=1.67929e-07 $layer=LI1_cond $X=4.13 $Y=1.895
+ $X2=4.245 $Y2=1.775
r135 71 73 6.42709 $w=2.58e-07 $l=1.45e-07 $layer=LI1_cond $X=4.13 $Y=1.895
+ $X2=4.13 $Y2=2.04
r136 67 81 2.23356 $w=6.15e-07 $l=1.67929e-07 $layer=LI1_cond $X=4.13 $Y=0.735
+ $X2=4.245 $Y2=0.855
r137 67 69 12.8542 $w=2.58e-07 $l=2.9e-07 $layer=LI1_cond $X=4.13 $Y=0.735
+ $X2=4.13 $Y2=0.445
r138 66 80 5.51899 $w=2.4e-07 $l=1.3e-07 $layer=LI1_cond $X=3.4 $Y=1.775
+ $X2=3.27 $Y2=1.775
r139 65 83 4.87019 $w=2.4e-07 $l=4.85e-07 $layer=LI1_cond $X=3.76 $Y=1.775
+ $X2=4.245 $Y2=1.775
r140 65 66 17.2866 $w=2.38e-07 $l=3.6e-07 $layer=LI1_cond $X=3.76 $Y=1.775
+ $X2=3.4 $Y2=1.775
r141 64 79 5.51899 $w=2.4e-07 $l=1.3e-07 $layer=LI1_cond $X=3.4 $Y=0.855
+ $X2=3.27 $Y2=0.855
r142 63 81 4.87019 $w=2.4e-07 $l=4.85e-07 $layer=LI1_cond $X=3.76 $Y=0.855
+ $X2=4.245 $Y2=0.855
r143 63 64 17.2866 $w=2.38e-07 $l=3.6e-07 $layer=LI1_cond $X=3.76 $Y=0.855
+ $X2=3.4 $Y2=0.855
r144 59 61 37.676 $w=2.58e-07 $l=8.5e-07 $layer=LI1_cond $X=3.27 $Y=2.04
+ $X2=3.27 $Y2=2.89
r145 57 80 1.05597 $w=2.6e-07 $l=1.2e-07 $layer=LI1_cond $X=3.27 $Y=1.895
+ $X2=3.27 $Y2=1.775
r146 57 59 6.42709 $w=2.58e-07 $l=1.45e-07 $layer=LI1_cond $X=3.27 $Y=1.895
+ $X2=3.27 $Y2=2.04
r147 53 79 1.05597 $w=2.6e-07 $l=1.2e-07 $layer=LI1_cond $X=3.27 $Y=0.735
+ $X2=3.27 $Y2=0.855
r148 53 55 12.8542 $w=2.58e-07 $l=2.9e-07 $layer=LI1_cond $X=3.27 $Y=0.735
+ $X2=3.27 $Y2=0.445
r149 52 78 5.51899 $w=2.4e-07 $l=1.3e-07 $layer=LI1_cond $X=2.54 $Y=1.775
+ $X2=2.41 $Y2=1.775
r150 51 80 5.51899 $w=2.4e-07 $l=1.3e-07 $layer=LI1_cond $X=3.14 $Y=1.775
+ $X2=3.27 $Y2=1.775
r151 51 52 28.8111 $w=2.38e-07 $l=6e-07 $layer=LI1_cond $X=3.14 $Y=1.775
+ $X2=2.54 $Y2=1.775
r152 50 77 5.51899 $w=2.4e-07 $l=1.3e-07 $layer=LI1_cond $X=2.54 $Y=0.855
+ $X2=2.41 $Y2=0.855
r153 49 79 5.51899 $w=2.4e-07 $l=1.3e-07 $layer=LI1_cond $X=3.14 $Y=0.855
+ $X2=3.27 $Y2=0.855
r154 49 50 28.8111 $w=2.38e-07 $l=6e-07 $layer=LI1_cond $X=3.14 $Y=0.855
+ $X2=2.54 $Y2=0.855
r155 45 47 37.676 $w=2.58e-07 $l=8.5e-07 $layer=LI1_cond $X=2.41 $Y=2.04
+ $X2=2.41 $Y2=2.89
r156 43 78 1.05597 $w=2.6e-07 $l=1.2e-07 $layer=LI1_cond $X=2.41 $Y=1.895
+ $X2=2.41 $Y2=1.775
r157 43 45 6.42709 $w=2.58e-07 $l=1.45e-07 $layer=LI1_cond $X=2.41 $Y=1.895
+ $X2=2.41 $Y2=2.04
r158 39 77 1.05597 $w=2.6e-07 $l=1.2e-07 $layer=LI1_cond $X=2.41 $Y=0.735
+ $X2=2.41 $Y2=0.855
r159 39 41 12.8542 $w=2.58e-07 $l=2.9e-07 $layer=LI1_cond $X=2.41 $Y=0.735
+ $X2=2.41 $Y2=0.445
r160 37 78 5.51899 $w=2.4e-07 $l=1.3e-07 $layer=LI1_cond $X=2.28 $Y=1.775
+ $X2=2.41 $Y2=1.775
r161 37 38 28.8111 $w=2.38e-07 $l=6e-07 $layer=LI1_cond $X=2.28 $Y=1.775
+ $X2=1.68 $Y2=1.775
r162 35 77 5.51899 $w=2.4e-07 $l=1.3e-07 $layer=LI1_cond $X=2.28 $Y=0.855
+ $X2=2.41 $Y2=0.855
r163 35 36 28.8111 $w=2.38e-07 $l=6e-07 $layer=LI1_cond $X=2.28 $Y=0.855
+ $X2=1.68 $Y2=0.855
r164 31 33 37.676 $w=2.58e-07 $l=8.5e-07 $layer=LI1_cond $X=1.55 $Y=2.04
+ $X2=1.55 $Y2=2.89
r165 29 38 6.83069 $w=2.4e-07 $l=1.80278e-07 $layer=LI1_cond $X=1.55 $Y=1.895
+ $X2=1.68 $Y2=1.775
r166 29 31 6.42709 $w=2.58e-07 $l=1.45e-07 $layer=LI1_cond $X=1.55 $Y=1.895
+ $X2=1.55 $Y2=2.04
r167 25 36 6.83069 $w=2.4e-07 $l=1.80278e-07 $layer=LI1_cond $X=1.55 $Y=0.735
+ $X2=1.68 $Y2=0.855
r168 25 27 12.8542 $w=2.58e-07 $l=2.9e-07 $layer=LI1_cond $X=1.55 $Y=0.735
+ $X2=1.55 $Y2=0.445
r169 8 75 400 $w=1.7e-07 $l=1.12282e-06 $layer=licon1_PDIFF $count=1 $X=3.99
+ $Y=1.835 $X2=4.13 $Y2=2.89
r170 8 73 400 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=1 $X=3.99
+ $Y=1.835 $X2=4.13 $Y2=2.04
r171 7 61 400 $w=1.7e-07 $l=1.12282e-06 $layer=licon1_PDIFF $count=1 $X=3.13
+ $Y=1.835 $X2=3.27 $Y2=2.89
r172 7 59 400 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=1 $X=3.13
+ $Y=1.835 $X2=3.27 $Y2=2.04
r173 6 47 400 $w=1.7e-07 $l=1.12282e-06 $layer=licon1_PDIFF $count=1 $X=2.27
+ $Y=1.835 $X2=2.41 $Y2=2.89
r174 6 45 400 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=1 $X=2.27
+ $Y=1.835 $X2=2.41 $Y2=2.04
r175 5 33 400 $w=1.7e-07 $l=1.12282e-06 $layer=licon1_PDIFF $count=1 $X=1.41
+ $Y=1.835 $X2=1.55 $Y2=2.89
r176 5 31 400 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=1 $X=1.41
+ $Y=1.835 $X2=1.55 $Y2=2.04
r177 4 69 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=3.99
+ $Y=0.235 $X2=4.13 $Y2=0.445
r178 3 55 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=3.13
+ $Y=0.235 $X2=3.27 $Y2=0.445
r179 2 41 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.27
+ $Y=0.235 $X2=2.41 $Y2=0.445
r180 1 27 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.41
+ $Y=0.235 $X2=1.55 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__CLKBUF_8%VGND 1 2 3 4 5 6 19 21 25 29 33 35 39 43 46
+ 47 49 50 51 52 53 65 72 73 79 82
r83 82 83 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r84 79 80 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r85 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r86 73 83 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=4.56
+ $Y2=0
r87 72 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r88 70 82 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=4.73 $Y=0 $X2=4.58
+ $Y2=0
r89 70 72 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=4.73 $Y=0 $X2=5.04
+ $Y2=0
r90 69 83 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=4.56
+ $Y2=0
r91 69 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.6
+ $Y2=0
r92 68 69 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r93 66 79 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.83 $Y=0 $X2=3.7
+ $Y2=0
r94 66 68 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=3.83 $Y=0 $X2=4.08
+ $Y2=0
r95 65 82 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=4.43 $Y=0 $X2=4.58
+ $Y2=0
r96 65 68 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=4.43 $Y=0 $X2=4.08
+ $Y2=0
r97 60 61 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r98 58 61 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r99 58 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r100 57 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r101 55 76 3.93884 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=0.39 $Y=0 $X2=0.195
+ $Y2=0
r102 55 57 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=0.39 $Y=0 $X2=0.72
+ $Y2=0
r103 53 80 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r104 53 61 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=1.68
+ $Y2=0
r105 53 63 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r106 51 63 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=2.71 $Y=0 $X2=2.64
+ $Y2=0
r107 51 52 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.71 $Y=0 $X2=2.84
+ $Y2=0
r108 49 60 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.85 $Y=0 $X2=1.68
+ $Y2=0
r109 49 50 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.85 $Y=0 $X2=1.98
+ $Y2=0
r110 48 63 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=2.11 $Y=0 $X2=2.64
+ $Y2=0
r111 48 50 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.11 $Y=0 $X2=1.98
+ $Y2=0
r112 46 57 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=0.99 $Y=0 $X2=0.72
+ $Y2=0
r113 46 47 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.99 $Y=0 $X2=1.12
+ $Y2=0
r114 45 60 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=1.25 $Y=0 $X2=1.68
+ $Y2=0
r115 45 47 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.25 $Y=0 $X2=1.12
+ $Y2=0
r116 41 82 0.597483 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.58 $Y=0.085
+ $X2=4.58 $Y2=0
r117 41 43 12.1007 $w=2.98e-07 $l=3.15e-07 $layer=LI1_cond $X=4.58 $Y=0.085
+ $X2=4.58 $Y2=0.4
r118 37 79 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=3.7 $Y=0.085
+ $X2=3.7 $Y2=0
r119 37 39 13.9623 $w=2.58e-07 $l=3.15e-07 $layer=LI1_cond $X=3.7 $Y=0.085
+ $X2=3.7 $Y2=0.4
r120 36 52 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.97 $Y=0 $X2=2.84
+ $Y2=0
r121 35 79 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.57 $Y=0 $X2=3.7
+ $Y2=0
r122 35 36 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=3.57 $Y=0 $X2=2.97
+ $Y2=0
r123 31 52 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=2.84 $Y=0.085
+ $X2=2.84 $Y2=0
r124 31 33 13.9623 $w=2.58e-07 $l=3.15e-07 $layer=LI1_cond $X=2.84 $Y=0.085
+ $X2=2.84 $Y2=0.4
r125 27 50 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=1.98 $Y=0.085
+ $X2=1.98 $Y2=0
r126 27 29 13.9623 $w=2.58e-07 $l=3.15e-07 $layer=LI1_cond $X=1.98 $Y=0.085
+ $X2=1.98 $Y2=0.4
r127 23 47 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=1.12 $Y=0.085
+ $X2=1.12 $Y2=0
r128 23 25 15.9569 $w=2.58e-07 $l=3.6e-07 $layer=LI1_cond $X=1.12 $Y=0.085
+ $X2=1.12 $Y2=0.445
r129 19 76 3.17127 $w=2.45e-07 $l=1.15521e-07 $layer=LI1_cond $X=0.267 $Y=0.085
+ $X2=0.195 $Y2=0
r130 19 21 16.9339 $w=2.43e-07 $l=3.6e-07 $layer=LI1_cond $X=0.267 $Y=0.085
+ $X2=0.267 $Y2=0.445
r131 6 43 182 $w=1.7e-07 $l=2.26164e-07 $layer=licon1_NDIFF $count=1 $X=4.42
+ $Y=0.235 $X2=4.565 $Y2=0.4
r132 5 39 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=3.56
+ $Y=0.235 $X2=3.7 $Y2=0.4
r133 4 33 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=2.7
+ $Y=0.235 $X2=2.84 $Y2=0.4
r134 3 29 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=1.84
+ $Y=0.235 $X2=1.98 $Y2=0.4
r135 2 25 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.98
+ $Y=0.235 $X2=1.12 $Y2=0.445
r136 1 21 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.445
.ends

