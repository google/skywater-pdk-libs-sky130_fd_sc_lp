# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_lp__dfxtp_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.120000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.580000 1.125000 2.075000 1.795000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  1.176000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.420000 0.255000 7.650000 1.055000 ;
        RECT 7.420000 1.055000 9.035000 1.225000 ;
        RECT 7.425000 1.735000 9.035000 1.905000 ;
        RECT 7.425000 1.905000 7.650000 3.075000 ;
        RECT 8.320000 0.255000 8.510000 0.840000 ;
        RECT 8.320000 0.840000 9.035000 1.055000 ;
        RECT 8.320000 1.905000 9.035000 1.945000 ;
        RECT 8.320000 1.945000 8.510000 3.075000 ;
        RECT 8.795000 1.225000 9.035000 1.735000 ;
        RECT 8.795000 1.945000 9.035000 2.490000 ;
    END
  END Q
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.840000 0.425000 2.490000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 9.120000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.500000 0.500000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.800000 0.500000 3.300000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 9.120000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 9.120000 0.085000 ;
      RECT 0.000000  3.245000 9.120000 3.415000 ;
      RECT 0.095000  0.085000 0.425000 0.670000 ;
      RECT 0.095000  2.665000 0.425000 3.245000 ;
      RECT 0.595000  0.395000 0.855000 1.195000 ;
      RECT 0.595000  1.195000 1.030000 1.865000 ;
      RECT 0.595000  1.865000 0.855000 2.990000 ;
      RECT 1.045000  2.045000 2.075000 2.215000 ;
      RECT 1.045000  2.215000 1.315000 2.715000 ;
      RECT 1.200000  0.640000 1.480000 0.960000 ;
      RECT 1.200000  0.960000 1.410000 2.045000 ;
      RECT 1.535000  2.395000 1.725000 3.245000 ;
      RECT 1.650000  0.085000 1.980000 0.955000 ;
      RECT 1.905000  2.215000 2.075000 2.535000 ;
      RECT 1.905000  2.535000 3.495000 2.705000 ;
      RECT 2.220000  0.625000 2.550000 0.955000 ;
      RECT 2.245000  0.955000 2.415000 1.930000 ;
      RECT 2.245000  1.930000 2.425000 2.355000 ;
      RECT 2.595000  1.545000 2.775000 2.535000 ;
      RECT 2.720000  0.640000 3.050000 1.105000 ;
      RECT 2.720000  1.105000 4.220000 1.275000 ;
      RECT 2.720000  1.275000 3.145000 1.350000 ;
      RECT 2.945000  1.350000 3.145000 2.355000 ;
      RECT 3.325000  2.285000 4.930000 2.455000 ;
      RECT 3.325000  2.455000 3.495000 2.535000 ;
      RECT 3.420000  1.445000 3.750000 1.855000 ;
      RECT 3.420000  1.855000 4.560000 1.915000 ;
      RECT 3.420000  1.915000 4.580000 2.115000 ;
      RECT 3.705000  0.085000 4.035000 0.935000 ;
      RECT 3.760000  2.625000 4.090000 3.245000 ;
      RECT 3.960000  1.275000 4.220000 1.675000 ;
      RECT 4.290000  0.585000 4.560000 0.935000 ;
      RECT 4.390000  0.935000 4.560000 1.855000 ;
      RECT 4.730000  1.225000 4.930000 1.555000 ;
      RECT 4.760000  1.555000 4.930000 2.285000 ;
      RECT 4.895000  0.640000 5.280000 0.995000 ;
      RECT 5.110000  0.995000 5.280000 1.015000 ;
      RECT 5.110000  1.015000 6.410000 1.185000 ;
      RECT 5.110000  1.185000 5.360000 2.700000 ;
      RECT 5.560000  1.355000 5.890000 1.695000 ;
      RECT 5.560000  1.695000 6.750000 1.865000 ;
      RECT 5.785000  0.085000 6.115000 0.845000 ;
      RECT 6.010000  2.035000 6.340000 3.245000 ;
      RECT 6.150000  1.185000 6.410000 1.515000 ;
      RECT 6.295000  0.285000 6.750000 0.845000 ;
      RECT 6.510000  1.865000 6.750000 3.005000 ;
      RECT 6.580000  0.845000 6.750000 1.395000 ;
      RECT 6.580000  1.395000 8.615000 1.565000 ;
      RECT 6.580000  1.565000 6.750000 1.695000 ;
      RECT 6.960000  0.085000 7.250000 1.095000 ;
      RECT 6.960000  1.815000 7.255000 3.245000 ;
      RECT 7.820000  0.085000 8.150000 0.885000 ;
      RECT 7.820000  2.075000 8.150000 3.245000 ;
      RECT 8.680000  0.085000 9.010000 0.670000 ;
      RECT 8.680000  2.660000 9.010000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
      RECT 8.315000 -0.085000 8.485000 0.085000 ;
      RECT 8.315000  3.245000 8.485000 3.415000 ;
      RECT 8.795000 -0.085000 8.965000 0.085000 ;
      RECT 8.795000  3.245000 8.965000 3.415000 ;
  END
END sky130_fd_sc_lp__dfxtp_4
