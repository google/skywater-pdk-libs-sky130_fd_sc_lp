* File: sky130_fd_sc_lp__dfsbp_1.spice
* Created: Wed Sep  2 09:44:01 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__dfsbp_1.pex.spice"
.subckt sky130_fd_sc_lp__dfsbp_1  VNB VPB CLK D SET_B VPWR Q Q_N VGND
* 
* VGND	VGND
* Q_N	Q_N
* Q	Q
* VPWR	VPWR
* SET_B	SET_B
* D	D
* CLK	CLK
* VPB	VPB
* VNB	VNB
MM1025 N_A_111_156#_M1025_d N_CLK_M1025_g N_VGND_M1025_s VNB NSHORT L=0.15
+ W=0.42 AD=0.1281 AS=0.1113 PD=1.45 PS=1.37 NRD=11.424 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1011 N_VGND_M1011_d N_A_111_156#_M1011_g N_A_161_21#_M1011_s VNB NSHORT L=0.15
+ W=0.42 AD=0.1386 AS=0.1113 PD=1.08 PS=1.37 NRD=2.856 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75002.2 A=0.063 P=1.14 MULT=1
MM1008 N_A_494_119#_M1008_d N_D_M1008_g N_VGND_M1011_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.1386 PD=0.7 PS=1.08 NRD=0 NRS=105.708 M=1 R=2.8 SA=75001
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1010 N_A_580_119#_M1010_d N_A_111_156#_M1010_g N_A_494_119#_M1008_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8
+ SA=75001.4 SB=75001 A=0.063 P=1.14 MULT=1
MM1000 A_666_119# N_A_161_21#_M1000_g N_A_580_119#_M1010_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75001.9
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1023 N_VGND_M1023_d N_A_708_93#_M1023_g A_666_119# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75002.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1012 A_964_169# N_A_580_119#_M1012_g N_A_708_93#_M1012_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.1113 PD=0.63 PS=1.37 NRD=14.28 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1009 N_VGND_M1009_d N_SET_B_M1009_g A_964_169# VNB NSHORT L=0.15 W=0.42
+ AD=0.0855057 AS=0.0441 PD=0.80434 PS=0.63 NRD=28.56 NRS=14.28 M=1 R=2.8
+ SA=75000.6 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1026 N_A_1141_125#_M1026_d N_A_580_119#_M1026_g N_VGND_M1009_d VNB NSHORT
+ L=0.15 W=0.64 AD=0.1696 AS=0.130294 PD=1.81 PS=1.22566 NRD=0 NRS=0 M=1
+ R=4.26667 SA=75000.8 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1019 N_A_1331_151#_M1019_d N_A_111_156#_M1019_g N_A_1248_151#_M1019_s VNB
+ NSHORT L=0.15 W=0.42 AD=0.0905774 AS=0.1113 PD=0.820189 PS=1.37 NRD=19.992
+ NRS=0 M=1 R=2.8 SA=75000.2 SB=75000.9 A=0.063 P=1.14 MULT=1
MM1020 N_A_1141_125#_M1020_d N_A_161_21#_M1020_g N_A_1331_151#_M1019_d VNB
+ NSHORT L=0.15 W=0.64 AD=0.3459 AS=0.138023 PD=2.7 PS=1.24981 NRD=91.02
+ NRS=8.436 M=1 R=4.26667 SA=75000.6 SB=75000.3 A=0.096 P=1.58 MULT=1
MM1016 A_1657_71# N_A_1535_177#_M1016_g N_A_1248_151#_M1016_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.1113 PD=0.63 PS=1.37 NRD=14.28 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1005 N_VGND_M1005_d N_SET_B_M1005_g A_1657_71# VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.0441 PD=1.37 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1024 N_VGND_M1024_d N_A_1331_151#_M1024_g N_A_1535_177#_M1024_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1027 N_A_2005_119#_M1027_d N_A_1331_151#_M1027_g N_VGND_M1024_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.6 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1022 N_VGND_M1022_d N_A_2005_119#_M1022_g N_Q_M1022_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1827 AS=0.2226 PD=1.275 PS=2.21 NRD=15.708 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75000.8 A=0.126 P=1.98 MULT=1
MM1001 N_Q_N_M1001_d N_A_1331_151#_M1001_g N_VGND_M1022_d VNB NSHORT L=0.15
+ W=0.84 AD=0.2226 AS=0.1827 PD=2.21 PS=1.275 NRD=0 NRS=6.42 M=1 R=5.6
+ SA=75000.8 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1021 N_A_111_156#_M1021_d N_CLK_M1021_g N_VPWR_M1021_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1696 AS=0.1696 PD=1.81 PS=1.81 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1002 N_VPWR_M1002_d N_A_111_156#_M1002_g N_A_161_21#_M1002_s VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.171411 AS=0.1696 PD=1.56377 PS=1.81 NRD=41.5473 NRS=0 M=1
+ R=4.26667 SA=75000.2 SB=75002.5 A=0.096 P=1.58 MULT=1
MM1018 N_A_494_119#_M1018_d N_D_M1018_g N_VPWR_M1002_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0588 AS=0.112489 PD=0.7 PS=1.02623 NRD=0 NRS=56.2829 M=1 R=2.8 SA=75000.7
+ SB=75004.4 A=0.063 P=1.14 MULT=1
MM1003 N_A_580_119#_M1003_d N_A_161_21#_M1003_g N_A_494_119#_M1018_d VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8
+ SA=75001.1 SB=75004 A=0.063 P=1.14 MULT=1
MM1028 A_687_533# N_A_111_156#_M1028_g N_A_580_119#_M1003_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=23.443 NRS=0 M=1 R=2.8
+ SA=75001.6 SB=75003.6 A=0.063 P=1.14 MULT=1
MM1031 N_VPWR_M1031_d N_A_708_93#_M1031_g A_687_533# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.28875 AS=0.0441 PD=1.795 PS=0.63 NRD=0 NRS=23.443 M=1 R=2.8 SA=75001.9
+ SB=75003.2 A=0.063 P=1.14 MULT=1
MM1029 N_A_708_93#_M1029_d N_A_580_119#_M1029_g N_VPWR_M1031_d VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.0588 AS=0.28875 PD=0.7 PS=1.795 NRD=0 NRS=513.599 M=1 R=2.8
+ SA=75003.4 SB=75001.7 A=0.063 P=1.14 MULT=1
MM1013 N_VPWR_M1013_d N_SET_B_M1013_g N_A_708_93#_M1029_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0952 AS=0.0588 PD=0.823333 PS=0.7 NRD=44.5417 NRS=0 M=1 R=2.8
+ SA=75003.9 SB=75001.3 A=0.063 P=1.14 MULT=1
MM1032 A_1259_449# N_A_580_119#_M1032_g N_VPWR_M1013_d VPB PHIGHVT L=0.15 W=0.84
+ AD=0.1638 AS=0.1904 PD=1.23 PS=1.64667 NRD=32.8202 NRS=4.6886 M=1 R=5.6
+ SA=75002.3 SB=75001.4 A=0.126 P=1.98 MULT=1
MM1007 N_A_1331_151#_M1007_d N_A_111_156#_M1007_g A_1259_449# VPB PHIGHVT L=0.15
+ W=0.84 AD=0.1792 AS=0.1638 PD=1.62 PS=1.23 NRD=0 NRS=32.8202 M=1 R=5.6
+ SA=75002.9 SB=75000.9 A=0.126 P=1.98 MULT=1
MM1033 A_1472_449# N_A_161_21#_M1033_g N_A_1331_151#_M1007_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.06615 AS=0.0896 PD=0.735 PS=0.81 NRD=48.068 NRS=44.5417 M=1 R=2.8
+ SA=75001.3 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1030 N_VPWR_M1030_d N_A_1535_177#_M1030_g A_1472_449# VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0588 AS=0.06615 PD=0.7 PS=0.735 NRD=0 NRS=48.068 M=1 R=2.8
+ SA=75001.7 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1015 N_A_1331_151#_M1015_d N_SET_B_M1015_g N_VPWR_M1030_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75002.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1006 N_VPWR_M1006_d N_A_1331_151#_M1006_g N_A_1535_177#_M1006_s VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.0905774 AS=0.1113 PD=0.820189 PS=1.37 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1017 N_A_2005_119#_M1017_d N_A_1331_151#_M1017_g N_VPWR_M1006_d VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.1696 AS=0.138023 PD=1.81 PS=1.24981 NRD=0 NRS=17.6906 M=1
+ R=4.26667 SA=75000.6 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1014 N_VPWR_M1014_d N_A_2005_119#_M1014_g N_Q_M1014_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1004 N_Q_N_M1004_d N_A_1331_151#_M1004_g N_VPWR_M1014_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX34_noxref VNB VPB NWDIODE A=23.9839 P=29.45
c_133 VNB 0 1.05346e-19 $X=0 $Y=0
c_258 VPB 0 5.82661e-20 $X=0 $Y=3.085
*
.include "sky130_fd_sc_lp__dfsbp_1.pxi.spice"
*
.ends
*
*
