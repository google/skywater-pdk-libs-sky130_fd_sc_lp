* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__and2b_4 A_N B VGND VNB VPB VPWR X
X0 a_43_367# A_N VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 X a_213_23# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X2 VGND a_213_23# X VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X3 X a_213_23# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X4 VGND B a_616_49# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X5 VPWR a_213_23# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X6 VGND a_213_23# X VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X7 a_43_367# A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X8 VPWR a_213_23# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X9 X a_213_23# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X10 a_213_23# a_43_367# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X11 VPWR B a_213_23# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X12 a_616_49# a_43_367# a_213_23# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X13 X a_213_23# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
.ends
