* File: sky130_fd_sc_lp__or4_0.pxi.spice
* Created: Wed Sep  2 10:31:42 2020
* 
x_PM_SKY130_FD_SC_LP__OR4_0%D N_D_M1000_g N_D_c_70_n N_D_M1005_g D D D D
+ PM_SKY130_FD_SC_LP__OR4_0%D
x_PM_SKY130_FD_SC_LP__OR4_0%C N_C_M1009_g N_C_c_101_n N_C_M1003_g N_C_c_103_n C
+ C N_C_c_100_n PM_SKY130_FD_SC_LP__OR4_0%C
x_PM_SKY130_FD_SC_LP__OR4_0%B N_B_c_132_n N_B_M1006_g N_B_M1007_g N_B_c_134_n B
+ B N_B_c_136_n N_B_c_137_n PM_SKY130_FD_SC_LP__OR4_0%B
x_PM_SKY130_FD_SC_LP__OR4_0%A N_A_M1008_g N_A_M1002_g N_A_c_179_n A A
+ N_A_c_181_n PM_SKY130_FD_SC_LP__OR4_0%A
x_PM_SKY130_FD_SC_LP__OR4_0%A_54_482# N_A_54_482#_M1000_d N_A_54_482#_M1007_d
+ N_A_54_482#_M1005_s N_A_54_482#_M1001_g N_A_54_482#_M1004_g
+ N_A_54_482#_c_229_n N_A_54_482#_c_230_n N_A_54_482#_c_243_n
+ N_A_54_482#_c_231_n N_A_54_482#_c_232_n N_A_54_482#_c_263_n
+ N_A_54_482#_c_245_n N_A_54_482#_c_246_n N_A_54_482#_c_247_n
+ N_A_54_482#_c_233_n N_A_54_482#_c_234_n N_A_54_482#_c_235_n
+ N_A_54_482#_c_236_n N_A_54_482#_c_237_n N_A_54_482#_c_238_n
+ N_A_54_482#_c_239_n N_A_54_482#_c_257_n N_A_54_482#_c_305_n
+ N_A_54_482#_c_240_n N_A_54_482#_c_241_n PM_SKY130_FD_SC_LP__OR4_0%A_54_482#
x_PM_SKY130_FD_SC_LP__OR4_0%VPWR N_VPWR_M1008_d N_VPWR_c_345_n VPWR
+ N_VPWR_c_346_n N_VPWR_c_347_n N_VPWR_c_344_n N_VPWR_c_349_n
+ PM_SKY130_FD_SC_LP__OR4_0%VPWR
x_PM_SKY130_FD_SC_LP__OR4_0%X N_X_M1001_d N_X_M1004_d X X X X X X X N_X_c_375_n
+ X PM_SKY130_FD_SC_LP__OR4_0%X
x_PM_SKY130_FD_SC_LP__OR4_0%VGND N_VGND_M1000_s N_VGND_M1009_d N_VGND_M1002_d
+ N_VGND_c_393_n N_VGND_c_394_n N_VGND_c_395_n N_VGND_c_396_n N_VGND_c_397_n
+ VGND N_VGND_c_398_n N_VGND_c_399_n N_VGND_c_400_n
+ PM_SKY130_FD_SC_LP__OR4_0%VGND
cc_1 VNB N_D_M1000_g 0.0253963f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=0.47
cc_2 VNB N_D_c_70_n 0.0976963f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.51
cc_3 VNB N_D_M1005_g 0.00697166f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=2.62
cc_4 VNB D 0.0355568f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_5 VNB N_C_M1009_g 0.0594188f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=0.47
cc_6 VNB C 0.00368393f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.95
cc_7 VNB N_C_c_100_n 0.0199443f $X=-0.19 $Y=-0.245 $X2=0.395 $Y2=1.005
cc_8 VNB N_B_c_132_n 0.0223654f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=0.47
cc_9 VNB N_B_M1006_g 0.0111615f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.51
cc_10 VNB N_B_c_134_n 0.0209878f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_11 VNB B 0.00646799f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.95
cc_12 VNB N_B_c_136_n 0.0227888f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_B_c_137_n 0.0192272f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.005
cc_14 VNB N_A_M1002_g 0.0380708f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=2.62
cc_15 VNB N_A_c_179_n 0.0193963f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.95
cc_16 VNB A 0.00521233f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_c_181_n 0.015329f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_54_482#_M1001_g 0.0249562f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.95
cc_19 VNB N_A_54_482#_M1004_g 0.00645341f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_54_482#_c_229_n 0.0243393f $X=-0.19 $Y=-0.245 $X2=0.225 $Y2=0.925
cc_21 VNB N_A_54_482#_c_230_n 0.0188048f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_54_482#_c_231_n 0.00218526f $X=-0.19 $Y=-0.245 $X2=0.225 $Y2=2.035
cc_23 VNB N_A_54_482#_c_232_n 0.0129979f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_54_482#_c_233_n 0.0015054f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_54_482#_c_234_n 0.00685346f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_54_482#_c_235_n 0.0021482f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_54_482#_c_236_n 0.0025859f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_54_482#_c_237_n 0.00253179f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_54_482#_c_238_n 7.45068e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_54_482#_c_239_n 0.00963399f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_54_482#_c_240_n 0.0172591f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_54_482#_c_241_n 0.00418577f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VPWR_c_344_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB X 0.0530748f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=2.62
cc_35 VNB N_X_c_375_n 0.0177078f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_393_n 0.01337f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_37 VNB N_VGND_c_394_n 0.0206306f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.95
cc_38 VNB N_VGND_c_395_n 0.00547034f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_396_n 0.0180086f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.005
cc_40 VNB N_VGND_c_397_n 0.00526527f $X=-0.19 $Y=-0.245 $X2=0.225 $Y2=0.925
cc_41 VNB N_VGND_c_398_n 0.0352253f $X=-0.19 $Y=-0.245 $X2=0.225 $Y2=1.295
cc_42 VNB N_VGND_c_399_n 0.0222567f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_400_n 0.19926f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VPB N_D_M1005_g 0.0593877f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=2.62
cc_45 VPB D 0.0312547f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_46 VPB N_C_c_101_n 0.0153036f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=1.51
cc_47 VPB N_C_M1003_g 0.0241877f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=2.62
cc_48 VPB N_C_c_103_n 0.0208837f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_49 VPB C 0.00797178f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.95
cc_50 VPB N_C_c_100_n 6.17862e-19 $X=-0.19 $Y=1.655 $X2=0.395 $Y2=1.005
cc_51 VPB N_B_M1006_g 0.0468687f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=1.51
cc_52 VPB N_A_M1008_g 0.0423861f $X=-0.19 $Y=1.655 $X2=0.55 $Y2=0.47
cc_53 VPB N_A_c_179_n 0.0415803f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.95
cc_54 VPB A 0.00360562f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_55 VPB N_A_54_482#_M1004_g 0.0619946f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_56 VPB N_A_54_482#_c_243_n 0.0158541f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_57 VPB N_A_54_482#_c_231_n 0.00553896f $X=-0.19 $Y=1.655 $X2=0.225 $Y2=2.035
cc_58 VPB N_A_54_482#_c_245_n 0.00174618f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_59 VPB N_A_54_482#_c_246_n 0.0227741f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_60 VPB N_A_54_482#_c_247_n 6.08079e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_61 VPB N_A_54_482#_c_238_n 0.00371389f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_62 VPB N_VPWR_c_345_n 0.0209794f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=2.62
cc_63 VPB N_VPWR_c_346_n 0.055609f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_64 VPB N_VPWR_c_347_n 0.0213525f $X=-0.19 $Y=1.655 $X2=0.225 $Y2=0.925
cc_65 VPB N_VPWR_c_344_n 0.0766085f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_349_n 0.0131466f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_67 VPB X 0.0390621f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=2.62
cc_68 VPB X 0.0463799f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_69 N_D_M1000_g N_C_M1009_g 0.0188563f $X=0.55 $Y=0.47 $X2=0 $Y2=0
cc_70 N_D_c_70_n N_C_M1009_g 0.0234202f $X=0.61 $Y=1.51 $X2=0 $Y2=0
cc_71 N_D_M1005_g N_C_M1003_g 0.0329913f $X=0.61 $Y=2.62 $X2=0 $Y2=0
cc_72 N_D_M1005_g N_C_c_103_n 0.0208752f $X=0.61 $Y=2.62 $X2=0 $Y2=0
cc_73 N_D_M1005_g C 9.11948e-19 $X=0.61 $Y=2.62 $X2=0 $Y2=0
cc_74 N_D_c_70_n N_C_c_100_n 0.0208752f $X=0.61 $Y=1.51 $X2=0 $Y2=0
cc_75 D N_A_54_482#_c_243_n 0.00908703f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_76 N_D_c_70_n N_A_54_482#_c_231_n 0.00323924f $X=0.61 $Y=1.51 $X2=0 $Y2=0
cc_77 N_D_M1005_g N_A_54_482#_c_231_n 0.0287639f $X=0.61 $Y=2.62 $X2=0 $Y2=0
cc_78 N_D_M1000_g N_A_54_482#_c_232_n 0.00546619f $X=0.55 $Y=0.47 $X2=0 $Y2=0
cc_79 N_D_c_70_n N_A_54_482#_c_232_n 0.00270982f $X=0.61 $Y=1.51 $X2=0 $Y2=0
cc_80 D N_A_54_482#_c_232_n 0.0228946f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_81 N_D_c_70_n N_A_54_482#_c_239_n 0.012195f $X=0.61 $Y=1.51 $X2=0 $Y2=0
cc_82 D N_A_54_482#_c_239_n 0.066564f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_83 N_D_M1005_g N_A_54_482#_c_257_n 0.011747f $X=0.61 $Y=2.62 $X2=0 $Y2=0
cc_84 N_D_M1005_g N_VPWR_c_346_n 0.00367021f $X=0.61 $Y=2.62 $X2=0 $Y2=0
cc_85 N_D_M1005_g N_VPWR_c_344_n 0.00505379f $X=0.61 $Y=2.62 $X2=0 $Y2=0
cc_86 N_D_M1000_g N_VGND_c_394_n 0.00380474f $X=0.55 $Y=0.47 $X2=0 $Y2=0
cc_87 N_D_c_70_n N_VGND_c_394_n 0.00503784f $X=0.61 $Y=1.51 $X2=0 $Y2=0
cc_88 D N_VGND_c_394_n 0.0173875f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_89 N_D_M1000_g N_VGND_c_398_n 0.00560159f $X=0.55 $Y=0.47 $X2=0 $Y2=0
cc_90 N_D_M1000_g N_VGND_c_400_n 0.0113522f $X=0.55 $Y=0.47 $X2=0 $Y2=0
cc_91 D N_VGND_c_400_n 0.00419678f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_92 N_C_M1003_g N_B_M1006_g 0.0335549f $X=1.06 $Y=2.62 $X2=0 $Y2=0
cc_93 C N_B_M1006_g 0.012774f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_94 N_C_c_100_n N_B_M1006_g 0.0401838f $X=1.06 $Y=1.665 $X2=0 $Y2=0
cc_95 N_C_M1009_g B 0.00262889f $X=0.98 $Y=0.47 $X2=0 $Y2=0
cc_96 N_C_M1009_g N_B_c_136_n 0.0217701f $X=0.98 $Y=0.47 $X2=0 $Y2=0
cc_97 N_C_M1009_g N_B_c_137_n 0.00544163f $X=0.98 $Y=0.47 $X2=0 $Y2=0
cc_98 N_C_M1009_g N_A_54_482#_c_231_n 0.0019126f $X=0.98 $Y=0.47 $X2=0 $Y2=0
cc_99 N_C_M1003_g N_A_54_482#_c_231_n 0.00365078f $X=1.06 $Y=2.62 $X2=0 $Y2=0
cc_100 C N_A_54_482#_c_231_n 0.0457402f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_101 N_C_c_100_n N_A_54_482#_c_231_n 0.00456707f $X=1.06 $Y=1.665 $X2=0 $Y2=0
cc_102 N_C_M1009_g N_A_54_482#_c_232_n 0.0118925f $X=0.98 $Y=0.47 $X2=0 $Y2=0
cc_103 N_C_c_101_n N_A_54_482#_c_263_n 8.28639e-19 $X=1.06 $Y=2.17 $X2=0 $Y2=0
cc_104 N_C_M1003_g N_A_54_482#_c_263_n 0.0184741f $X=1.06 $Y=2.62 $X2=0 $Y2=0
cc_105 C N_A_54_482#_c_263_n 0.0246838f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_106 N_C_M1003_g N_A_54_482#_c_245_n 0.00122298f $X=1.06 $Y=2.62 $X2=0 $Y2=0
cc_107 C N_A_54_482#_c_247_n 0.0144747f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_108 N_C_M1003_g N_VPWR_c_346_n 0.00367106f $X=1.06 $Y=2.62 $X2=0 $Y2=0
cc_109 N_C_M1003_g N_VPWR_c_344_n 0.00505379f $X=1.06 $Y=2.62 $X2=0 $Y2=0
cc_110 N_C_M1009_g N_VGND_c_398_n 0.00790038f $X=0.98 $Y=0.47 $X2=0 $Y2=0
cc_111 N_C_M1009_g N_VGND_c_400_n 0.0110928f $X=0.98 $Y=0.47 $X2=0 $Y2=0
cc_112 B N_A_M1002_g 0.00136138f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_113 N_B_c_137_n N_A_M1002_g 0.0302217f $X=1.63 $Y=0.79 $X2=0 $Y2=0
cc_114 N_B_M1006_g N_A_c_179_n 0.0813327f $X=1.51 $Y=2.62 $X2=0 $Y2=0
cc_115 N_B_c_134_n N_A_c_179_n 0.00955055f $X=1.63 $Y=1.46 $X2=0 $Y2=0
cc_116 B N_A_c_179_n 4.69121e-19 $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_117 N_B_c_132_n A 8.21872e-19 $X=1.63 $Y=1.265 $X2=0 $Y2=0
cc_118 N_B_M1006_g A 0.0051867f $X=1.51 $Y=2.62 $X2=0 $Y2=0
cc_119 B A 0.0237542f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_120 N_B_c_132_n N_A_c_181_n 0.0080853f $X=1.63 $Y=1.265 $X2=0 $Y2=0
cc_121 B N_A_c_181_n 8.61885e-19 $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_122 B N_A_54_482#_c_232_n 0.0187631f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_123 N_B_M1006_g N_A_54_482#_c_263_n 0.0141168f $X=1.51 $Y=2.62 $X2=0 $Y2=0
cc_124 N_B_M1006_g N_A_54_482#_c_245_n 0.00571441f $X=1.51 $Y=2.62 $X2=0 $Y2=0
cc_125 N_B_c_134_n N_A_54_482#_c_246_n 8.14082e-19 $X=1.63 $Y=1.46 $X2=0 $Y2=0
cc_126 B N_A_54_482#_c_246_n 0.00693738f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_127 N_B_M1006_g N_A_54_482#_c_247_n 0.00769728f $X=1.51 $Y=2.62 $X2=0 $Y2=0
cc_128 N_B_c_134_n N_A_54_482#_c_247_n 3.07792e-19 $X=1.63 $Y=1.46 $X2=0 $Y2=0
cc_129 B N_A_54_482#_c_247_n 0.00578106f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_130 B N_A_54_482#_c_233_n 0.00412554f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_131 N_B_c_137_n N_A_54_482#_c_233_n 0.00386796f $X=1.63 $Y=0.79 $X2=0 $Y2=0
cc_132 B N_A_54_482#_c_235_n 0.0143975f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_133 N_B_c_136_n N_A_54_482#_c_235_n 0.00126769f $X=1.63 $Y=0.955 $X2=0 $Y2=0
cc_134 B N_A_54_482#_c_237_n 0.00523733f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_135 N_B_M1006_g N_VPWR_c_345_n 0.00125097f $X=1.51 $Y=2.62 $X2=0 $Y2=0
cc_136 N_B_M1006_g N_VPWR_c_346_n 0.00367038f $X=1.51 $Y=2.62 $X2=0 $Y2=0
cc_137 N_B_M1006_g N_VPWR_c_344_n 0.00505379f $X=1.51 $Y=2.62 $X2=0 $Y2=0
cc_138 N_B_c_137_n N_VGND_c_396_n 0.00560159f $X=1.63 $Y=0.79 $X2=0 $Y2=0
cc_139 B N_VGND_c_398_n 0.0149147f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_140 N_B_c_136_n N_VGND_c_398_n 0.00681461f $X=1.63 $Y=0.955 $X2=0 $Y2=0
cc_141 N_B_c_137_n N_VGND_c_398_n 0.00244456f $X=1.63 $Y=0.79 $X2=0 $Y2=0
cc_142 B N_VGND_c_400_n 0.00537277f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_143 N_B_c_136_n N_VGND_c_400_n 2.86346e-19 $X=1.63 $Y=0.955 $X2=0 $Y2=0
cc_144 N_B_c_137_n N_VGND_c_400_n 0.00711963f $X=1.63 $Y=0.79 $X2=0 $Y2=0
cc_145 N_A_M1002_g N_A_54_482#_M1001_g 0.0234827f $X=2.18 $Y=0.47 $X2=0 $Y2=0
cc_146 N_A_M1008_g N_A_54_482#_M1004_g 0.00834747f $X=1.87 $Y=2.62 $X2=0 $Y2=0
cc_147 N_A_c_179_n N_A_54_482#_M1004_g 0.0161972f $X=2.2 $Y=1.73 $X2=0 $Y2=0
cc_148 A N_A_54_482#_M1004_g 3.01831e-19 $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_149 A N_A_54_482#_c_229_n 3.07359e-19 $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_150 N_A_c_181_n N_A_54_482#_c_229_n 0.0083195f $X=2.2 $Y=1.375 $X2=0 $Y2=0
cc_151 N_A_c_179_n N_A_54_482#_c_230_n 0.0083195f $X=2.2 $Y=1.73 $X2=0 $Y2=0
cc_152 N_A_M1008_g N_A_54_482#_c_245_n 0.00358118f $X=1.87 $Y=2.62 $X2=0 $Y2=0
cc_153 N_A_M1008_g N_A_54_482#_c_246_n 0.0185601f $X=1.87 $Y=2.62 $X2=0 $Y2=0
cc_154 N_A_c_179_n N_A_54_482#_c_246_n 0.00722309f $X=2.2 $Y=1.73 $X2=0 $Y2=0
cc_155 A N_A_54_482#_c_246_n 0.0226162f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_156 N_A_M1002_g N_A_54_482#_c_233_n 0.00587321f $X=2.18 $Y=0.47 $X2=0 $Y2=0
cc_157 N_A_M1002_g N_A_54_482#_c_234_n 0.00821698f $X=2.18 $Y=0.47 $X2=0 $Y2=0
cc_158 A N_A_54_482#_c_234_n 0.0107941f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_159 N_A_c_181_n N_A_54_482#_c_234_n 0.0034905f $X=2.2 $Y=1.375 $X2=0 $Y2=0
cc_160 N_A_M1002_g N_A_54_482#_c_235_n 0.00236668f $X=2.18 $Y=0.47 $X2=0 $Y2=0
cc_161 N_A_c_179_n N_A_54_482#_c_235_n 6.67588e-19 $X=2.2 $Y=1.73 $X2=0 $Y2=0
cc_162 A N_A_54_482#_c_235_n 0.0126163f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_163 N_A_c_181_n N_A_54_482#_c_235_n 5.0609e-19 $X=2.2 $Y=1.375 $X2=0 $Y2=0
cc_164 N_A_M1002_g N_A_54_482#_c_237_n 0.00199412f $X=2.18 $Y=0.47 $X2=0 $Y2=0
cc_165 A N_A_54_482#_c_237_n 0.0509983f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_166 N_A_c_181_n N_A_54_482#_c_237_n 0.0016586f $X=2.2 $Y=1.375 $X2=0 $Y2=0
cc_167 N_A_M1008_g N_A_54_482#_c_238_n 0.00296117f $X=1.87 $Y=2.62 $X2=0 $Y2=0
cc_168 N_A_c_179_n N_A_54_482#_c_238_n 0.0016586f $X=2.2 $Y=1.73 $X2=0 $Y2=0
cc_169 N_A_M1002_g N_A_54_482#_c_305_n 0.00422327f $X=2.18 $Y=0.47 $X2=0 $Y2=0
cc_170 N_A_c_179_n N_A_54_482#_c_241_n 0.0016586f $X=2.2 $Y=1.73 $X2=0 $Y2=0
cc_171 N_A_M1008_g N_VPWR_c_345_n 0.0127476f $X=1.87 $Y=2.62 $X2=0 $Y2=0
cc_172 N_A_M1008_g N_VPWR_c_346_n 0.00405273f $X=1.87 $Y=2.62 $X2=0 $Y2=0
cc_173 N_A_M1008_g N_VPWR_c_344_n 0.00424518f $X=1.87 $Y=2.62 $X2=0 $Y2=0
cc_174 N_A_M1002_g N_VGND_c_395_n 0.00312753f $X=2.18 $Y=0.47 $X2=0 $Y2=0
cc_175 N_A_M1002_g N_VGND_c_396_n 0.00504402f $X=2.18 $Y=0.47 $X2=0 $Y2=0
cc_176 N_A_M1002_g N_VGND_c_400_n 0.00607344f $X=2.18 $Y=0.47 $X2=0 $Y2=0
cc_177 N_A_54_482#_c_263_n A_137_482# 0.00969419f $X=1.465 $Y=2.607 $X2=-0.19
+ $Y2=-0.245
cc_178 N_A_54_482#_c_263_n A_227_482# 0.00760697f $X=1.465 $Y=2.607 $X2=-0.19
+ $Y2=-0.245
cc_179 N_A_54_482#_M1004_g N_VPWR_c_345_n 0.00497163f $X=2.705 $Y=2.73 $X2=0
+ $Y2=0
cc_180 N_A_54_482#_c_245_n N_VPWR_c_345_n 0.00160929f $X=1.55 $Y=2.43 $X2=0
+ $Y2=0
cc_181 N_A_54_482#_c_246_n N_VPWR_c_345_n 0.0586867f $X=2.465 $Y=2.135 $X2=0
+ $Y2=0
cc_182 N_A_54_482#_c_243_n N_VPWR_c_346_n 0.00703076f $X=0.535 $Y=2.62 $X2=0
+ $Y2=0
cc_183 N_A_54_482#_c_263_n N_VPWR_c_346_n 0.0181337f $X=1.465 $Y=2.607 $X2=0
+ $Y2=0
cc_184 N_A_54_482#_c_257_n N_VPWR_c_346_n 0.00358385f $X=0.62 $Y=2.607 $X2=0
+ $Y2=0
cc_185 N_A_54_482#_M1004_g N_VPWR_c_347_n 0.0053511f $X=2.705 $Y=2.73 $X2=0
+ $Y2=0
cc_186 N_A_54_482#_M1004_g N_VPWR_c_344_n 0.0118241f $X=2.705 $Y=2.73 $X2=0
+ $Y2=0
cc_187 N_A_54_482#_c_243_n N_VPWR_c_344_n 0.0105152f $X=0.535 $Y=2.62 $X2=0
+ $Y2=0
cc_188 N_A_54_482#_c_263_n N_VPWR_c_344_n 0.029102f $X=1.465 $Y=2.607 $X2=0
+ $Y2=0
cc_189 N_A_54_482#_c_257_n N_VPWR_c_344_n 0.00532688f $X=0.62 $Y=2.607 $X2=0
+ $Y2=0
cc_190 N_A_54_482#_M1001_g X 0.00677575f $X=2.68 $Y=0.47 $X2=0 $Y2=0
cc_191 N_A_54_482#_M1004_g X 0.0184886f $X=2.705 $Y=2.73 $X2=0 $Y2=0
cc_192 N_A_54_482#_c_246_n X 0.010007f $X=2.465 $Y=2.135 $X2=0 $Y2=0
cc_193 N_A_54_482#_c_236_n X 0.0139296f $X=2.66 $Y=1.03 $X2=0 $Y2=0
cc_194 N_A_54_482#_c_237_n X 0.0390794f $X=2.66 $Y=1.335 $X2=0 $Y2=0
cc_195 N_A_54_482#_c_238_n X 0.028633f $X=2.612 $Y=2.05 $X2=0 $Y2=0
cc_196 N_A_54_482#_c_240_n X 0.0166276f $X=2.77 $Y=1.025 $X2=0 $Y2=0
cc_197 N_A_54_482#_c_236_n N_X_c_375_n 0.00428675f $X=2.66 $Y=1.03 $X2=0 $Y2=0
cc_198 N_A_54_482#_c_240_n N_X_c_375_n 0.0038259f $X=2.77 $Y=1.025 $X2=0 $Y2=0
cc_199 N_A_54_482#_M1004_g X 0.00731895f $X=2.705 $Y=2.73 $X2=0 $Y2=0
cc_200 N_A_54_482#_M1001_g N_VGND_c_395_n 0.00323971f $X=2.68 $Y=0.47 $X2=0
+ $Y2=0
cc_201 N_A_54_482#_c_234_n N_VGND_c_395_n 0.00963001f $X=2.465 $Y=0.945 $X2=0
+ $Y2=0
cc_202 N_A_54_482#_c_236_n N_VGND_c_395_n 0.0073714f $X=2.66 $Y=1.03 $X2=0 $Y2=0
cc_203 N_A_54_482#_c_305_n N_VGND_c_395_n 0.0251167f $X=2.06 $Y=0.47 $X2=0 $Y2=0
cc_204 N_A_54_482#_c_305_n N_VGND_c_396_n 0.013105f $X=2.06 $Y=0.47 $X2=0 $Y2=0
cc_205 N_A_54_482#_c_232_n N_VGND_c_398_n 0.0113476f $X=0.765 $Y=0.47 $X2=0
+ $Y2=0
cc_206 N_A_54_482#_M1001_g N_VGND_c_399_n 0.00560159f $X=2.68 $Y=0.47 $X2=0
+ $Y2=0
cc_207 N_A_54_482#_M1001_g N_VGND_c_400_n 0.00719246f $X=2.68 $Y=0.47 $X2=0
+ $Y2=0
cc_208 N_A_54_482#_c_232_n N_VGND_c_400_n 0.00977851f $X=0.765 $Y=0.47 $X2=0
+ $Y2=0
cc_209 N_A_54_482#_c_234_n N_VGND_c_400_n 0.00553439f $X=2.465 $Y=0.945 $X2=0
+ $Y2=0
cc_210 N_A_54_482#_c_236_n N_VGND_c_400_n 0.00613862f $X=2.66 $Y=1.03 $X2=0
+ $Y2=0
cc_211 N_A_54_482#_c_305_n N_VGND_c_400_n 0.0112979f $X=2.06 $Y=0.47 $X2=0 $Y2=0
cc_212 N_VPWR_c_345_n X 0.0293867f $X=2.47 $Y=2.555 $X2=0 $Y2=0
cc_213 N_VPWR_c_347_n X 0.0356959f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_214 N_VPWR_c_344_n X 0.0193447f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_215 N_X_c_375_n N_VGND_c_399_n 0.0249217f $X=3.15 $Y=0.47 $X2=0 $Y2=0
cc_216 N_X_c_375_n N_VGND_c_400_n 0.0190978f $X=3.15 $Y=0.47 $X2=0 $Y2=0
