* File: sky130_fd_sc_lp__sdlclkp_4.pex.spice
* Created: Fri Aug 28 11:31:38 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__SDLCLKP_4%SCE 3 7 11 14 15 16 17 18 19 26
r34 26 27 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.27
+ $Y=1.12 $X2=0.27 $Y2=1.12
r35 18 19 12.183 $w=3.48e-07 $l=3.7e-07 $layer=LI1_cond $X=0.26 $Y=2.035
+ $X2=0.26 $Y2=2.405
r36 17 18 12.183 $w=3.48e-07 $l=3.7e-07 $layer=LI1_cond $X=0.26 $Y=1.665
+ $X2=0.26 $Y2=2.035
r37 16 17 12.183 $w=3.48e-07 $l=3.7e-07 $layer=LI1_cond $X=0.26 $Y=1.295
+ $X2=0.26 $Y2=1.665
r38 16 27 5.76222 $w=3.48e-07 $l=1.75e-07 $layer=LI1_cond $X=0.26 $Y=1.295
+ $X2=0.26 $Y2=1.12
r39 15 27 6.42075 $w=3.48e-07 $l=1.95e-07 $layer=LI1_cond $X=0.26 $Y=0.925
+ $X2=0.26 $Y2=1.12
r40 13 26 47.5746 $w=4.15e-07 $l=3.55e-07 $layer=POLY_cond $X=0.312 $Y=1.475
+ $X2=0.312 $Y2=1.12
r41 13 14 44.0182 $w=4.15e-07 $l=1.5e-07 $layer=POLY_cond $X=0.327 $Y=1.475
+ $X2=0.327 $Y2=1.625
r42 11 26 2.01019 $w=4.15e-07 $l=1.5e-08 $layer=POLY_cond $X=0.312 $Y=1.105
+ $X2=0.312 $Y2=1.12
r43 10 11 44.0182 $w=4.15e-07 $l=1.5e-07 $layer=POLY_cond $X=0.387 $Y=0.955
+ $X2=0.387 $Y2=1.105
r44 7 10 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.595 $Y=0.56
+ $X2=0.595 $Y2=0.955
r45 3 14 530.713 $w=1.5e-07 $l=1.035e-06 $layer=POLY_cond $X=0.475 $Y=2.66
+ $X2=0.475 $Y2=1.625
.ends

.subckt PM_SKY130_FD_SC_LP__SDLCLKP_4%GATE 3 7 12 16 18 20 29 44
r58 29 30 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.15
+ $Y=1.09 $X2=1.15 $Y2=1.09
r59 18 20 7.70628 $w=7.43e-07 $l=4.8e-07 $layer=LI1_cond $X=1.68 $Y=1.417
+ $X2=2.16 $Y2=1.417
r60 18 44 5.85998 $w=7.43e-07 $l=3.65e-07 $layer=LI1_cond $X=1.68 $Y=1.417
+ $X2=1.315 $Y2=1.417
r61 16 44 1.89055 $w=8.63e-07 $l=1.15e-07 $layer=LI1_cond $X=1.2 $Y=1.357
+ $X2=1.315 $Y2=1.357
r62 16 30 0.705202 $w=8.63e-07 $l=5e-08 $layer=LI1_cond $X=1.2 $Y=1.357 $X2=1.15
+ $Y2=1.357
r63 15 29 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.15 $Y=0.925
+ $X2=1.15 $Y2=1.09
r64 12 29 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=1.15 $Y=1.445
+ $X2=1.15 $Y2=1.09
r65 9 12 161.521 $w=1.5e-07 $l=3.15e-07 $layer=POLY_cond $X=0.835 $Y=1.52
+ $X2=1.15 $Y2=1.52
r66 7 15 187.16 $w=1.5e-07 $l=3.65e-07 $layer=POLY_cond $X=1.06 $Y=0.56 $X2=1.06
+ $Y2=0.925
r67 1 9 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.835 $Y=1.595
+ $X2=0.835 $Y2=1.52
r68 1 3 546.096 $w=1.5e-07 $l=1.065e-06 $layer=POLY_cond $X=0.835 $Y=1.595
+ $X2=0.835 $Y2=2.66
.ends

.subckt PM_SKY130_FD_SC_LP__SDLCLKP_4%A_252_361# 1 2 8 9 10 11 12 15 17 18 20 21
+ 23 24 26 28 30 33 35 36 38 39 42 44 47 48 50 52 57
c148 57 0 1.62725e-19 $X=5.265 $Y=0.445
c149 50 0 1.28129e-19 $X=5.56 $Y=2.035
c150 44 0 1.81312e-19 $X=5.085 $Y=0.61
c151 18 0 1.54235e-19 $X=1.675 $Y=1.27
c152 17 0 1.43117e-19 $X=1.955 $Y=1.27
c153 15 0 3.58312e-20 $X=1.6 $Y=0.56
r154 52 54 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=3.785 $Y=0.35
+ $X2=3.785 $Y2=0.61
r155 48 50 16.1082 $w=2.08e-07 $l=3.05e-07 $layer=LI1_cond $X=5.255 $Y=2.035
+ $X2=5.56 $Y2=2.035
r156 47 48 6.91519 $w=2.1e-07 $l=1.41244e-07 $layer=LI1_cond $X=5.17 $Y=1.93
+ $X2=5.255 $Y2=2.035
r157 47 60 80.5722 $w=1.68e-07 $l=1.235e-06 $layer=LI1_cond $X=5.17 $Y=1.93
+ $X2=5.17 $Y2=0.695
r158 45 54 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.87 $Y=0.61
+ $X2=3.785 $Y2=0.61
r159 44 60 5.80707 $w=3.43e-07 $l=8.5e-08 $layer=LI1_cond $X=5.257 $Y=0.61
+ $X2=5.257 $Y2=0.695
r160 44 57 5.51168 $w=3.43e-07 $l=1.65e-07 $layer=LI1_cond $X=5.257 $Y=0.61
+ $X2=5.257 $Y2=0.445
r161 44 45 79.2674 $w=1.68e-07 $l=1.215e-06 $layer=LI1_cond $X=5.085 $Y=0.61
+ $X2=3.87 $Y2=0.61
r162 41 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.43
+ $Y=0.35 $X2=2.43 $Y2=0.35
r163 39 52 0.0262452 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=3.7 $Y=0.35
+ $X2=3.785 $Y2=0.35
r164 39 41 74.134 $w=1.88e-07 $l=1.27e-06 $layer=LI1_cond $X=3.7 $Y=0.35
+ $X2=2.43 $Y2=0.35
r165 37 42 147.758 $w=3.3e-07 $l=8.45e-07 $layer=POLY_cond $X=2.43 $Y=1.195
+ $X2=2.43 $Y2=0.35
r166 37 38 5.03009 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=2.43 $Y=1.195
+ $X2=2.43 $Y2=1.27
r167 31 33 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=3.525 $Y=3.075
+ $X2=3.525 $Y2=2.525
r168 28 30 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=3.095 $Y=1.195
+ $X2=3.095 $Y2=0.875
r169 27 38 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.595 $Y=1.27
+ $X2=2.43 $Y2=1.27
r170 26 28 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.02 $Y=1.27
+ $X2=3.095 $Y2=1.195
r171 26 27 217.926 $w=1.5e-07 $l=4.25e-07 $layer=POLY_cond $X=3.02 $Y=1.27
+ $X2=2.595 $Y2=1.27
r172 25 35 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.105 $Y=1.27
+ $X2=2.03 $Y2=1.27
r173 24 38 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.265 $Y=1.27
+ $X2=2.43 $Y2=1.27
r174 24 25 82.0426 $w=1.5e-07 $l=1.6e-07 $layer=POLY_cond $X=2.265 $Y=1.27
+ $X2=2.105 $Y2=1.27
r175 21 36 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.03 $Y=1.955
+ $X2=2.03 $Y2=1.88
r176 21 23 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=2.03 $Y=1.955
+ $X2=2.03 $Y2=2.385
r177 20 36 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.03 $Y=1.805
+ $X2=2.03 $Y2=1.88
r178 19 35 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.03 $Y=1.345
+ $X2=2.03 $Y2=1.27
r179 19 20 235.872 $w=1.5e-07 $l=4.6e-07 $layer=POLY_cond $X=2.03 $Y=1.345
+ $X2=2.03 $Y2=1.805
r180 17 35 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.955 $Y=1.27
+ $X2=2.03 $Y2=1.27
r181 17 18 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=1.955 $Y=1.27
+ $X2=1.675 $Y2=1.27
r182 13 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.6 $Y=1.195
+ $X2=1.675 $Y2=1.27
r183 13 15 325.606 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.6 $Y=1.195
+ $X2=1.6 $Y2=0.56
r184 11 31 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.45 $Y=3.15
+ $X2=3.525 $Y2=3.075
r185 11 12 1046.04 $w=1.5e-07 $l=2.04e-06 $layer=POLY_cond $X=3.45 $Y=3.15
+ $X2=1.41 $Y2=3.15
r186 9 36 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.955 $Y=1.88
+ $X2=2.03 $Y2=1.88
r187 9 10 279.457 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=1.955 $Y=1.88
+ $X2=1.41 $Y2=1.88
r188 8 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.335 $Y=3.075
+ $X2=1.41 $Y2=3.15
r189 7 10 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.335 $Y=1.955
+ $X2=1.41 $Y2=1.88
r190 7 8 574.298 $w=1.5e-07 $l=1.12e-06 $layer=POLY_cond $X=1.335 $Y=1.955
+ $X2=1.335 $Y2=3.075
r191 2 50 600 $w=1.7e-07 $l=2.54951e-07 $layer=licon1_PDIFF $count=1 $X=5.435
+ $Y=1.835 $X2=5.56 $Y2=2.035
r192 1 57 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=5.14
+ $Y=0.235 $X2=5.265 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__SDLCLKP_4%A_335_70# 1 2 7 11 13 15 17 19 21 28 31 36
+ 40
c75 21 0 3.58312e-20 $X=2.425 $Y=0.7
r76 36 37 8.2139 $w=3.78e-07 $l=1.65e-07 $layer=LI1_cond $X=2.415 $Y=2.21
+ $X2=2.415 $Y2=2.045
r77 31 33 4.88915 $w=3.28e-07 $l=1.4e-07 $layer=LI1_cond $X=1.815 $Y=0.56
+ $X2=1.815 $Y2=0.7
r78 29 40 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.51 $Y=1.74
+ $X2=2.675 $Y2=1.74
r79 28 37 18.7929 $w=1.78e-07 $l=3.05e-07 $layer=LI1_cond $X=2.515 $Y=1.74
+ $X2=2.515 $Y2=2.045
r80 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.51
+ $Y=1.74 $X2=2.51 $Y2=1.74
r81 25 28 58.8434 $w=1.78e-07 $l=9.55e-07 $layer=LI1_cond $X=2.515 $Y=0.785
+ $X2=2.515 $Y2=1.74
r82 22 33 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.98 $Y=0.7
+ $X2=1.815 $Y2=0.7
r83 21 25 6.82373 $w=1.7e-07 $l=1.25499e-07 $layer=LI1_cond $X=2.425 $Y=0.7
+ $X2=2.515 $Y2=0.785
r84 21 22 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=2.425 $Y=0.7
+ $X2=1.98 $Y2=0.7
r85 15 20 83.3023 $w=1.66e-07 $l=2.9483e-07 $layer=POLY_cond $X=3.525 $Y=1.375
+ $X2=3.505 $Y2=1.66
r86 15 17 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=3.525 $Y=1.375
+ $X2=3.525 $Y2=0.875
r87 14 19 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.17 $Y=1.66
+ $X2=3.095 $Y2=1.66
r88 13 20 5.24352 $w=1.5e-07 $l=9.5e-08 $layer=POLY_cond $X=3.41 $Y=1.66
+ $X2=3.505 $Y2=1.66
r89 13 14 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=3.41 $Y=1.66
+ $X2=3.17 $Y2=1.66
r90 9 19 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.095 $Y=1.735
+ $X2=3.095 $Y2=1.66
r91 9 11 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.095 $Y=1.735
+ $X2=3.095 $Y2=2.525
r92 7 19 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.02 $Y=1.66
+ $X2=3.095 $Y2=1.66
r93 7 40 176.904 $w=1.5e-07 $l=3.45e-07 $layer=POLY_cond $X=3.02 $Y=1.66
+ $X2=2.675 $Y2=1.66
r94 2 36 300 $w=1.7e-07 $l=2.67862e-07 $layer=licon1_PDIFF $count=2 $X=2.105
+ $Y=2.065 $X2=2.31 $Y2=2.21
r95 1 31 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.675
+ $Y=0.35 $X2=1.815 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_LP__SDLCLKP_4%A_762_107# 1 2 9 13 15 17 18 22 28 31 35
+ 36 39 40 41 43 44 48 53 55 57 61 62 68
c141 68 0 4.9125e-20 $X=6.75 $Y=1.675
c142 61 0 2.97134e-19 $X=6.75 $Y=1.51
c143 9 0 3.05678e-20 $X=3.885 $Y=0.875
r144 62 68 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.75 $Y=1.51
+ $X2=6.75 $Y2=1.675
r145 61 62 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.75
+ $Y=1.51 $X2=6.75 $Y2=1.51
r146 58 61 13.969 $w=3.28e-07 $l=4e-07 $layer=LI1_cond $X=6.35 $Y=1.51 $X2=6.75
+ $Y2=1.51
r147 51 53 4.93138 $w=2.13e-07 $l=9.2e-08 $layer=LI1_cond $X=4.725 $Y=0.972
+ $X2=4.817 $Y2=0.972
r148 48 66 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.975 $Y=1.93
+ $X2=3.975 $Y2=2.095
r149 48 65 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.975 $Y=1.93
+ $X2=3.975 $Y2=1.765
r150 47 48 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.975
+ $Y=1.93 $X2=3.975 $Y2=1.93
r151 44 47 7.22427 $w=3.33e-07 $l=2.1e-07 $layer=LI1_cond $X=3.972 $Y=1.72
+ $X2=3.972 $Y2=1.93
r152 42 58 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.35 $Y=1.675
+ $X2=6.35 $Y2=1.51
r153 42 43 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=6.35 $Y=1.675
+ $X2=6.35 $Y2=1.93
r154 40 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.265 $Y=2.015
+ $X2=6.35 $Y2=1.93
r155 40 41 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=6.265 $Y=2.015
+ $X2=6.075 $Y2=2.015
r156 38 41 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.99 $Y=2.1
+ $X2=6.075 $Y2=2.015
r157 38 39 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=5.99 $Y=2.1
+ $X2=5.99 $Y2=2.31
r158 37 57 2.80098 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=5.04 $Y=2.4
+ $X2=4.875 $Y2=2.4
r159 36 39 6.82373 $w=1.8e-07 $l=1.25499e-07 $layer=LI1_cond $X=5.905 $Y=2.4
+ $X2=5.99 $Y2=2.31
r160 36 37 53.298 $w=1.78e-07 $l=8.65e-07 $layer=LI1_cond $X=5.905 $Y=2.4
+ $X2=5.04 $Y2=2.4
r161 35 55 4.50329 $w=2e-07 $l=8.74643e-08 $layer=LI1_cond $X=4.817 $Y=1.635
+ $X2=4.812 $Y2=1.72
r162 34 53 1.33342 $w=1.95e-07 $l=1.08e-07 $layer=LI1_cond $X=4.817 $Y=1.08
+ $X2=4.817 $Y2=0.972
r163 34 35 31.5664 $w=1.93e-07 $l=5.55e-07 $layer=LI1_cond $X=4.817 $Y=1.08
+ $X2=4.817 $Y2=1.635
r164 31 57 3.67302 $w=2.67e-07 $l=1.17346e-07 $layer=LI1_cond $X=4.812 $Y=2.31
+ $X2=4.875 $Y2=2.4
r165 30 55 4.50329 $w=2e-07 $l=8.5e-08 $layer=LI1_cond $X=4.812 $Y=1.805
+ $X2=4.812 $Y2=1.72
r166 30 31 27.3215 $w=2.03e-07 $l=5.05e-07 $layer=LI1_cond $X=4.812 $Y=1.805
+ $X2=4.812 $Y2=2.31
r167 29 44 4.71304 $w=1.7e-07 $l=1.68e-07 $layer=LI1_cond $X=4.14 $Y=1.72
+ $X2=3.972 $Y2=1.72
r168 28 55 1.93381 $w=1.7e-07 $l=1.02e-07 $layer=LI1_cond $X=4.71 $Y=1.72
+ $X2=4.812 $Y2=1.72
r169 28 29 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=4.71 $Y=1.72
+ $X2=4.14 $Y2=1.72
r170 22 68 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=6.73 $Y=2.465
+ $X2=6.73 $Y2=1.675
r171 18 24 197.415 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=6.75 $Y=1.26
+ $X2=6.365 $Y2=1.26
r172 18 62 30.6007 $w=3.3e-07 $l=1.75e-07 $layer=POLY_cond $X=6.75 $Y=1.335
+ $X2=6.75 $Y2=1.51
r173 15 24 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.365 $Y=1.185
+ $X2=6.365 $Y2=1.26
r174 15 17 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=6.365 $Y=1.185
+ $X2=6.365 $Y2=0.655
r175 13 66 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=3.885 $Y=2.525
+ $X2=3.885 $Y2=2.095
r176 9 65 456.362 $w=1.5e-07 $l=8.9e-07 $layer=POLY_cond $X=3.885 $Y=0.875
+ $X2=3.885 $Y2=1.765
r177 2 57 300 $w=1.7e-07 $l=7.96932e-07 $layer=licon1_PDIFF $count=2 $X=4.735
+ $Y=1.695 $X2=4.875 $Y2=2.425
r178 1 51 182 $w=1.7e-07 $l=7.81873e-07 $layer=licon1_NDIFF $count=1 $X=4.585
+ $Y=0.245 $X2=4.725 $Y2=0.96
.ends

.subckt PM_SKY130_FD_SC_LP__SDLCLKP_4%A_634_133# 1 2 7 9 12 16 20 24 27 29
r67 25 29 23.4065 $w=2.78e-07 $l=1.35e-07 $layer=POLY_cond $X=4.375 $Y=1.36
+ $X2=4.51 $Y2=1.36
r68 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.375
+ $Y=1.36 $X2=4.375 $Y2=1.36
r69 22 27 2.50281 $w=2.15e-07 $l=1.48e-07 $layer=LI1_cond $X=3.475 $Y=1.357
+ $X2=3.327 $Y2=1.357
r70 22 24 48.2418 $w=2.13e-07 $l=9e-07 $layer=LI1_cond $X=3.475 $Y=1.357
+ $X2=4.375 $Y2=1.357
r71 18 27 3.94093 $w=2.95e-07 $l=1.08e-07 $layer=LI1_cond $X=3.327 $Y=1.465
+ $X2=3.327 $Y2=1.357
r72 18 20 41.6051 $w=2.93e-07 $l=1.065e-06 $layer=LI1_cond $X=3.327 $Y=1.465
+ $X2=3.327 $Y2=2.53
r73 14 27 3.94093 $w=2.95e-07 $l=1.07e-07 $layer=LI1_cond $X=3.327 $Y=1.25
+ $X2=3.327 $Y2=1.357
r74 14 16 14.6497 $w=2.93e-07 $l=3.75e-07 $layer=LI1_cond $X=3.327 $Y=1.25
+ $X2=3.327 $Y2=0.875
r75 10 29 26.0072 $w=2.78e-07 $l=2.2798e-07 $layer=POLY_cond $X=4.66 $Y=1.525
+ $X2=4.51 $Y2=1.36
r76 10 12 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=4.66 $Y=1.525 $X2=4.66
+ $Y2=2.325
r77 7 29 17.1848 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.51 $Y=1.195
+ $X2=4.51 $Y2=1.36
r78 7 9 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=4.51 $Y=1.195 $X2=4.51
+ $Y2=0.665
r79 2 20 600 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_PDIFF $count=1 $X=3.17
+ $Y=2.315 $X2=3.31 $Y2=2.53
r80 1 16 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=3.17
+ $Y=0.665 $X2=3.31 $Y2=0.875
.ends

.subckt PM_SKY130_FD_SC_LP__SDLCLKP_4%CLK 3 5 7 10 12 14 15 17 28
c55 17 0 4.9125e-20 $X=6 $Y=1.665
c56 12 0 1.28129e-19 $X=6.3 $Y=1.725
c57 10 0 1.62725e-19 $X=6.005 $Y=0.655
c58 3 0 1.81312e-19 $X=5.48 $Y=0.445
r59 27 28 37.7075 $w=2.94e-07 $l=2.3e-07 $layer=POLY_cond $X=5.775 $Y=1.535
+ $X2=6.005 $Y2=1.535
r60 25 27 33.6088 $w=2.94e-07 $l=2.05e-07 $layer=POLY_cond $X=5.57 $Y=1.535
+ $X2=5.775 $Y2=1.535
r61 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.57
+ $Y=1.51 $X2=5.57 $Y2=1.51
r62 23 25 14.7551 $w=2.94e-07 $l=9e-08 $layer=POLY_cond $X=5.48 $Y=1.535
+ $X2=5.57 $Y2=1.535
r63 17 26 9.35116 $w=5.48e-07 $l=4.3e-07 $layer=LI1_cond $X=6 $Y=1.485 $X2=5.57
+ $Y2=1.485
r64 15 26 1.08734 $w=5.48e-07 $l=5e-08 $layer=LI1_cond $X=5.52 $Y=1.485 $X2=5.57
+ $Y2=1.485
r65 12 28 48.3639 $w=2.94e-07 $l=3.78253e-07 $layer=POLY_cond $X=6.3 $Y=1.725
+ $X2=6.005 $Y2=1.535
r66 12 14 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=6.3 $Y=1.725 $X2=6.3
+ $Y2=2.465
r67 8 28 18.4939 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=6.005 $Y=1.345
+ $X2=6.005 $Y2=1.535
r68 8 10 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=6.005 $Y=1.345
+ $X2=6.005 $Y2=0.655
r69 5 27 18.4939 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=5.775 $Y=1.725
+ $X2=5.775 $Y2=1.535
r70 5 7 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=5.775 $Y=1.725
+ $X2=5.775 $Y2=2.155
r71 1 23 18.4939 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=5.48 $Y=1.345
+ $X2=5.48 $Y2=1.535
r72 1 3 461.489 $w=1.5e-07 $l=9e-07 $layer=POLY_cond $X=5.48 $Y=1.345 $X2=5.48
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__SDLCLKP_4%A_1275_367# 1 2 9 11 13 16 18 20 23 25 27
+ 30 32 34 39 43 44 45 46 48 54 58 59 60 73
c122 73 0 2.79516e-19 $X=8.615 $Y=1.35
c123 48 0 1.29324e-19 $X=7.11 $Y=1.845
c124 9 0 1.40035e-19 $X=7.265 $Y=2.465
r125 72 73 10.4917 $w=3.3e-07 $l=6e-08 $layer=POLY_cond $X=8.555 $Y=1.35
+ $X2=8.615 $Y2=1.35
r126 71 72 64.6987 $w=3.3e-07 $l=3.7e-07 $layer=POLY_cond $X=8.185 $Y=1.35
+ $X2=8.555 $Y2=1.35
r127 70 71 10.4917 $w=3.3e-07 $l=6e-08 $layer=POLY_cond $X=8.125 $Y=1.35
+ $X2=8.185 $Y2=1.35
r128 67 68 10.4917 $w=3.3e-07 $l=6e-08 $layer=POLY_cond $X=7.695 $Y=1.35
+ $X2=7.755 $Y2=1.35
r129 66 67 64.6987 $w=3.3e-07 $l=3.7e-07 $layer=POLY_cond $X=7.325 $Y=1.35
+ $X2=7.695 $Y2=1.35
r130 58 59 8.55446 $w=3.73e-07 $l=1.65e-07 $layer=LI1_cond $X=6.597 $Y=2.445
+ $X2=6.597 $Y2=2.28
r131 55 70 27.1035 $w=3.3e-07 $l=1.55e-07 $layer=POLY_cond $X=7.97 $Y=1.35
+ $X2=8.125 $Y2=1.35
r132 55 68 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=7.97 $Y=1.35
+ $X2=7.755 $Y2=1.35
r133 54 55 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=7.97
+ $Y=1.35 $X2=7.97 $Y2=1.35
r134 52 66 6.12014 $w=3.3e-07 $l=3.5e-08 $layer=POLY_cond $X=7.29 $Y=1.35
+ $X2=7.325 $Y2=1.35
r135 52 63 4.37153 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=7.29 $Y=1.35
+ $X2=7.265 $Y2=1.35
r136 51 54 31.3464 $w=2.48e-07 $l=6.8e-07 $layer=LI1_cond $X=7.29 $Y=1.31
+ $X2=7.97 $Y2=1.31
r137 51 52 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=7.29
+ $Y=1.35 $X2=7.29 $Y2=1.35
r138 49 60 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=7.11 $Y=1.31
+ $X2=7.11 $Y2=1.085
r139 49 51 4.37928 $w=2.48e-07 $l=9.5e-08 $layer=LI1_cond $X=7.195 $Y=1.31
+ $X2=7.29 $Y2=1.31
r140 47 49 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=7.11 $Y=1.435
+ $X2=7.11 $Y2=1.31
r141 47 48 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=7.11 $Y=1.435
+ $X2=7.11 $Y2=1.845
r142 45 48 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.025 $Y=1.93
+ $X2=7.11 $Y2=1.845
r143 45 46 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=7.025 $Y=1.93
+ $X2=6.785 $Y2=1.93
r144 43 60 0.364908 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=7.025 $Y=1.085
+ $X2=7.11 $Y2=1.085
r145 43 44 20.9495 $w=1.78e-07 $l=3.4e-07 $layer=LI1_cond $X=7.025 $Y=1.085
+ $X2=6.685 $Y2=1.085
r146 41 46 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.7 $Y=2.015
+ $X2=6.785 $Y2=1.93
r147 41 59 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=6.7 $Y=2.015
+ $X2=6.7 $Y2=2.28
r148 37 44 7.17723 $w=1.8e-07 $l=1.74284e-07 $layer=LI1_cond $X=6.55 $Y=0.995
+ $X2=6.685 $Y2=1.085
r149 37 39 24.5428 $w=2.68e-07 $l=5.75e-07 $layer=LI1_cond $X=6.55 $Y=0.995
+ $X2=6.55 $Y2=0.42
r150 32 73 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.615 $Y=1.185
+ $X2=8.615 $Y2=1.35
r151 32 34 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=8.615 $Y=1.185
+ $X2=8.615 $Y2=0.655
r152 28 72 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.555 $Y=1.515
+ $X2=8.555 $Y2=1.35
r153 28 30 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=8.555 $Y=1.515
+ $X2=8.555 $Y2=2.465
r154 25 71 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.185 $Y=1.185
+ $X2=8.185 $Y2=1.35
r155 25 27 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=8.185 $Y=1.185
+ $X2=8.185 $Y2=0.655
r156 21 70 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.125 $Y=1.515
+ $X2=8.125 $Y2=1.35
r157 21 23 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=8.125 $Y=1.515
+ $X2=8.125 $Y2=2.465
r158 18 68 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.755 $Y=1.185
+ $X2=7.755 $Y2=1.35
r159 18 20 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=7.755 $Y=1.185
+ $X2=7.755 $Y2=0.655
r160 14 67 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.695 $Y=1.515
+ $X2=7.695 $Y2=1.35
r161 14 16 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=7.695 $Y=1.515
+ $X2=7.695 $Y2=2.465
r162 11 66 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.325 $Y=1.185
+ $X2=7.325 $Y2=1.35
r163 11 13 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=7.325 $Y=1.185
+ $X2=7.325 $Y2=0.655
r164 7 63 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.265 $Y=1.515
+ $X2=7.265 $Y2=1.35
r165 7 9 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=7.265 $Y=1.515
+ $X2=7.265 $Y2=2.465
r166 2 58 300 $w=1.7e-07 $l=6.76387e-07 $layer=licon1_PDIFF $count=2 $X=6.375
+ $Y=1.835 $X2=6.515 $Y2=2.445
r167 1 39 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=6.44
+ $Y=0.235 $X2=6.58 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__SDLCLKP_4%VPWR 1 2 3 4 5 6 7 22 24 28 31 34 38 40 44
+ 48 52 54 59 61 63 68 73 78 83 92 95 98 101 104 108
c116 44 0 1.22416e-19 $X=7.05 $Y=2.35
c117 5 0 1.29324e-19 $X=6.805 $Y=1.835
r118 107 108 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r119 104 105 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r120 101 102 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r121 99 102 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=3.33
+ $X2=6.96 $Y2=3.33
r122 98 99 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r123 95 96 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r124 92 93 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r125 89 90 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r126 87 108 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=8.88 $Y2=3.33
r127 87 105 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=7.92 $Y2=3.33
r128 86 87 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=3.33 $X2=8.4
+ $Y2=3.33
r129 84 104 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=8.04 $Y=3.33
+ $X2=7.91 $Y2=3.33
r130 84 86 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=8.04 $Y=3.33
+ $X2=8.4 $Y2=3.33
r131 83 107 4.01281 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=8.675 $Y=3.33
+ $X2=8.897 $Y2=3.33
r132 83 86 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=8.675 $Y=3.33
+ $X2=8.4 $Y2=3.33
r133 82 105 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=7.92 $Y2=3.33
r134 82 102 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=6.96 $Y2=3.33
r135 81 82 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r136 79 101 6.81202 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=7.195 $Y=3.33
+ $X2=7.075 $Y2=3.33
r137 79 81 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=7.195 $Y=3.33
+ $X2=7.44 $Y2=3.33
r138 78 104 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=7.78 $Y=3.33
+ $X2=7.91 $Y2=3.33
r139 78 81 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=7.78 $Y=3.33
+ $X2=7.44 $Y2=3.33
r140 74 95 12.4999 $w=1.7e-07 $l=2.98e-07 $layer=LI1_cond $X=4.53 $Y=3.33
+ $X2=4.232 $Y2=3.33
r141 74 76 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=4.53 $Y=3.33 $X2=4.56
+ $Y2=3.33
r142 73 98 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=5.98 $Y=3.33
+ $X2=6.085 $Y2=3.33
r143 73 76 92.6417 $w=1.68e-07 $l=1.42e-06 $layer=LI1_cond $X=5.98 $Y=3.33
+ $X2=4.56 $Y2=3.33
r144 72 96 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r145 72 93 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=1.68 $Y2=3.33
r146 71 72 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r147 69 92 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.705 $Y=3.33
+ $X2=1.575 $Y2=3.33
r148 69 71 123.631 $w=1.68e-07 $l=1.895e-06 $layer=LI1_cond $X=1.705 $Y=3.33
+ $X2=3.6 $Y2=3.33
r149 68 95 12.4999 $w=1.7e-07 $l=2.97e-07 $layer=LI1_cond $X=3.935 $Y=3.33
+ $X2=4.232 $Y2=3.33
r150 68 71 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=3.935 $Y=3.33
+ $X2=3.6 $Y2=3.33
r151 67 93 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r152 67 90 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.24 $Y2=3.33
r153 66 67 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r154 64 89 4.21867 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=0.365 $Y=3.33
+ $X2=0.182 $Y2=3.33
r155 64 66 54.4759 $w=1.68e-07 $l=8.35e-07 $layer=LI1_cond $X=0.365 $Y=3.33
+ $X2=1.2 $Y2=3.33
r156 63 92 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.445 $Y=3.33
+ $X2=1.575 $Y2=3.33
r157 63 66 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=1.445 $Y=3.33
+ $X2=1.2 $Y2=3.33
r158 61 99 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=6 $Y2=3.33
r159 61 96 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=4.08 $Y2=3.33
r160 61 76 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r161 59 60 8.62559 $w=5.93e-07 $l=1.3e-07 $layer=LI1_cond $X=4.232 $Y=2.49
+ $X2=4.232 $Y2=2.36
r162 54 57 41.222 $w=2.58e-07 $l=9.3e-07 $layer=LI1_cond $X=8.805 $Y=1.98
+ $X2=8.805 $Y2=2.91
r163 52 107 3.19941 $w=2.6e-07 $l=1.27609e-07 $layer=LI1_cond $X=8.805 $Y=3.245
+ $X2=8.897 $Y2=3.33
r164 52 57 14.8488 $w=2.58e-07 $l=3.35e-07 $layer=LI1_cond $X=8.805 $Y=3.245
+ $X2=8.805 $Y2=2.91
r165 48 51 37.2328 $w=2.58e-07 $l=8.4e-07 $layer=LI1_cond $X=7.91 $Y=2.11
+ $X2=7.91 $Y2=2.95
r166 46 104 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=7.91 $Y=3.245
+ $X2=7.91 $Y2=3.33
r167 46 51 13.0758 $w=2.58e-07 $l=2.95e-07 $layer=LI1_cond $X=7.91 $Y=3.245
+ $X2=7.91 $Y2=2.95
r168 42 101 0.135687 $w=2.4e-07 $l=8.5e-08 $layer=LI1_cond $X=7.075 $Y=3.245
+ $X2=7.075 $Y2=3.33
r169 42 44 42.9765 $w=2.38e-07 $l=8.95e-07 $layer=LI1_cond $X=7.075 $Y=3.245
+ $X2=7.075 $Y2=2.35
r170 41 98 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=6.19 $Y=3.33
+ $X2=6.085 $Y2=3.33
r171 40 101 6.81202 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=6.955 $Y=3.33
+ $X2=7.075 $Y2=3.33
r172 40 41 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=6.955 $Y=3.33
+ $X2=6.19 $Y2=3.33
r173 36 98 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=6.085 $Y=3.245
+ $X2=6.085 $Y2=3.33
r174 36 38 15.5801 $w=2.08e-07 $l=2.95e-07 $layer=LI1_cond $X=6.085 $Y=3.245
+ $X2=6.085 $Y2=2.95
r175 34 60 12.2584 $w=1.88e-07 $l=2.1e-07 $layer=LI1_cond $X=4.435 $Y=2.15
+ $X2=4.435 $Y2=2.36
r176 31 95 2.50116 $w=5.95e-07 $l=8.5e-08 $layer=LI1_cond $X=4.232 $Y=3.245
+ $X2=4.232 $Y2=3.33
r177 30 59 3.35706 $w=5.93e-07 $l=1.67e-07 $layer=LI1_cond $X=4.232 $Y=2.657
+ $X2=4.232 $Y2=2.49
r178 30 31 11.8201 $w=5.93e-07 $l=5.88e-07 $layer=LI1_cond $X=4.232 $Y=2.657
+ $X2=4.232 $Y2=3.245
r179 26 92 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=1.575 $Y=3.245
+ $X2=1.575 $Y2=3.33
r180 26 28 34.5733 $w=2.58e-07 $l=7.8e-07 $layer=LI1_cond $X=1.575 $Y=3.245
+ $X2=1.575 $Y2=2.465
r181 22 89 3.06603 $w=2.7e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.23 $Y=3.245
+ $X2=0.182 $Y2=3.33
r182 22 24 17.9269 $w=2.68e-07 $l=4.2e-07 $layer=LI1_cond $X=0.23 $Y=3.245
+ $X2=0.23 $Y2=2.825
r183 7 57 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=8.63
+ $Y=1.835 $X2=8.77 $Y2=2.91
r184 7 54 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=8.63
+ $Y=1.835 $X2=8.77 $Y2=1.98
r185 6 51 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=7.77
+ $Y=1.835 $X2=7.91 $Y2=2.95
r186 6 48 400 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=1 $X=7.77
+ $Y=1.835 $X2=7.91 $Y2=2.11
r187 5 44 300 $w=1.7e-07 $l=6.2562e-07 $layer=licon1_PDIFF $count=2 $X=6.805
+ $Y=1.835 $X2=7.05 $Y2=2.35
r188 4 38 600 $w=1.7e-07 $l=1.22689e-06 $layer=licon1_PDIFF $count=1 $X=5.85
+ $Y=1.835 $X2=6.085 $Y2=2.95
r189 3 59 200 $w=1.7e-07 $l=5.65774e-07 $layer=licon1_PDIFF $count=3 $X=3.96
+ $Y=2.315 $X2=4.445 $Y2=2.49
r190 3 34 600 $w=1.7e-07 $l=5.61471e-07 $layer=licon1_PDIFF $count=1 $X=3.96
+ $Y=2.315 $X2=4.445 $Y2=2.15
r191 2 28 600 $w=1.7e-07 $l=4.58258e-07 $layer=licon1_PDIFF $count=1 $X=1.485
+ $Y=2.065 $X2=1.61 $Y2=2.465
r192 1 24 600 $w=1.7e-07 $l=5.43921e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.34 $X2=0.26 $Y2=2.825
.ends

.subckt PM_SKY130_FD_SC_LP__SDLCLKP_4%A_134_70# 1 2 3 4 14 17 19 22 23 24 27 32
+ 35
c75 19 0 2.97352e-19 $X=1.875 $Y=2.045
r76 32 34 8.06855 $w=2.68e-07 $l=1.65e-07 $layer=LI1_cond $X=0.84 $Y=0.56
+ $X2=0.84 $Y2=0.725
r77 27 30 81.1614 $w=2.33e-07 $l=1.655e-06 $layer=LI1_cond $X=2.892 $Y=0.875
+ $X2=2.892 $Y2=2.53
r78 25 30 17.4092 $w=2.33e-07 $l=3.55e-07 $layer=LI1_cond $X=2.892 $Y=2.885
+ $X2=2.892 $Y2=2.53
r79 23 25 6.91636 $w=1.9e-07 $l=1.57493e-07 $layer=LI1_cond $X=2.775 $Y=2.98
+ $X2=2.892 $Y2=2.885
r80 23 24 42.6124 $w=1.88e-07 $l=7.3e-07 $layer=LI1_cond $X=2.775 $Y=2.98
+ $X2=2.045 $Y2=2.98
r81 22 24 6.84389 $w=1.9e-07 $l=1.30767e-07 $layer=LI1_cond $X=1.96 $Y=2.885
+ $X2=2.045 $Y2=2.98
r82 21 22 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=1.96 $Y=2.13
+ $X2=1.96 $Y2=2.885
r83 20 35 4.03347 $w=1.7e-07 $l=2.55e-07 $layer=LI1_cond $X=1.215 $Y=2.045
+ $X2=0.96 $Y2=2.045
r84 19 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.875 $Y=2.045
+ $X2=1.96 $Y2=2.13
r85 19 20 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=1.875 $Y=2.045
+ $X2=1.215 $Y2=2.045
r86 15 35 2.73602 $w=3.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.96 $Y=2.13 $X2=0.96
+ $Y2=2.045
r87 15 17 8.32564 $w=5.08e-07 $l=3.55e-07 $layer=LI1_cond $X=0.96 $Y=2.13
+ $X2=0.96 $Y2=2.485
r88 14 35 2.73602 $w=3.5e-07 $l=1.9799e-07 $layer=LI1_cond $X=0.8 $Y=1.96
+ $X2=0.96 $Y2=2.045
r89 14 34 72.0909 $w=1.88e-07 $l=1.235e-06 $layer=LI1_cond $X=0.8 $Y=1.96
+ $X2=0.8 $Y2=0.725
r90 4 30 600 $w=1.7e-07 $l=2.7037e-07 $layer=licon1_PDIFF $count=1 $X=2.755
+ $Y=2.315 $X2=2.88 $Y2=2.53
r91 3 17 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=0.91
+ $Y=2.34 $X2=1.05 $Y2=2.485
r92 2 27 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=2.755
+ $Y=0.665 $X2=2.88 $Y2=0.875
r93 1 32 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.67
+ $Y=0.35 $X2=0.81 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_LP__SDLCLKP_4%GCLK 1 2 3 4 15 21 23 24 25 26 31 33 34 35
+ 36 37
r54 37 56 8.0085 $w=2.93e-07 $l=2.05e-07 $layer=LI1_cond $X=8.357 $Y=1.98
+ $X2=8.357 $Y2=1.775
r55 36 52 3.74047 $w=2.47e-07 $l=1.06325e-07 $layer=LI1_cond $X=8.357 $Y=1.69
+ $X2=8.405 $Y2=1.605
r56 36 56 3.74047 $w=2.47e-07 $l=8.5e-08 $layer=LI1_cond $X=8.357 $Y=1.69
+ $X2=8.357 $Y2=1.775
r57 36 52 0.720909 $w=1.98e-07 $l=1.3e-08 $layer=LI1_cond $X=8.405 $Y=1.592
+ $X2=8.405 $Y2=1.605
r58 35 36 16.47 $w=1.98e-07 $l=2.97e-07 $layer=LI1_cond $X=8.405 $Y=1.295
+ $X2=8.405 $Y2=1.592
r59 35 51 15.5273 $w=1.98e-07 $l=2.8e-07 $layer=LI1_cond $X=8.405 $Y=1.295
+ $X2=8.405 $Y2=1.015
r60 34 45 4.50329 $w=2e-07 $l=8.5e-08 $layer=LI1_cond $X=8.405 $Y=0.93 $X2=8.405
+ $Y2=0.845
r61 34 51 4.50329 $w=2e-07 $l=8.5e-08 $layer=LI1_cond $X=8.405 $Y=0.93 $X2=8.405
+ $Y2=1.015
r62 34 45 0.166364 $w=1.98e-07 $l=3e-09 $layer=LI1_cond $X=8.405 $Y=0.842
+ $X2=8.405 $Y2=0.845
r63 33 34 15.9155 $w=1.98e-07 $l=2.87e-07 $layer=LI1_cond $X=8.405 $Y=0.555
+ $X2=8.405 $Y2=0.842
r64 29 37 13.3996 $w=2.93e-07 $l=3.43e-07 $layer=LI1_cond $X=8.357 $Y=2.323
+ $X2=8.357 $Y2=1.98
r65 29 31 4.37538 $w=2.93e-07 $l=1.12e-07 $layer=LI1_cond $X=8.357 $Y=2.323
+ $X2=8.357 $Y2=2.435
r66 25 34 1.93381 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=8.305 $Y=0.93 $X2=8.405
+ $Y2=0.93
r67 25 26 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=8.305 $Y=0.93
+ $X2=7.635 $Y2=0.93
r68 23 36 2.72405 $w=1.7e-07 $l=1.47e-07 $layer=LI1_cond $X=8.21 $Y=1.69
+ $X2=8.357 $Y2=1.69
r69 23 24 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=8.21 $Y=1.69 $X2=7.61
+ $Y2=1.69
r70 19 26 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=7.54 $Y=0.845
+ $X2=7.635 $Y2=0.93
r71 19 21 24.8086 $w=1.88e-07 $l=4.25e-07 $layer=LI1_cond $X=7.54 $Y=0.845
+ $X2=7.54 $Y2=0.42
r72 15 17 43.7458 $w=2.43e-07 $l=9.3e-07 $layer=LI1_cond $X=7.487 $Y=1.98
+ $X2=7.487 $Y2=2.91
r73 13 24 7.11011 $w=1.7e-07 $l=1.5995e-07 $layer=LI1_cond $X=7.487 $Y=1.775
+ $X2=7.61 $Y2=1.69
r74 13 15 9.64289 $w=2.43e-07 $l=2.05e-07 $layer=LI1_cond $X=7.487 $Y=1.775
+ $X2=7.487 $Y2=1.98
r75 4 37 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=8.2
+ $Y=1.835 $X2=8.34 $Y2=1.98
r76 4 31 300 $w=1.7e-07 $l=6.66333e-07 $layer=licon1_PDIFF $count=2 $X=8.2
+ $Y=1.835 $X2=8.34 $Y2=2.435
r77 3 17 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=7.34
+ $Y=1.835 $X2=7.48 $Y2=2.91
r78 3 15 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=7.34
+ $Y=1.835 $X2=7.48 $Y2=1.98
r79 2 34 182 $w=1.7e-07 $l=7.61791e-07 $layer=licon1_NDIFF $count=1 $X=8.26
+ $Y=0.235 $X2=8.4 $Y2=0.93
r80 2 33 182 $w=1.7e-07 $l=4.19196e-07 $layer=licon1_NDIFF $count=1 $X=8.26
+ $Y=0.235 $X2=8.4 $Y2=0.59
r81 1 21 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=7.4
+ $Y=0.235 $X2=7.54 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__SDLCLKP_4%VGND 1 2 3 4 5 6 7 22 24 26 30 34 40 44 46
+ 48 51 52 53 55 67 71 76 85 89 95 98 102
c115 102 0 3.05678e-20 $X=8.88 $Y=0
r116 101 102 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=0
+ $X2=8.88 $Y2=0
r117 98 99 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r118 95 96 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r119 89 92 9.07985 $w=3.28e-07 $l=2.6e-07 $layer=LI1_cond $X=4.215 $Y=0
+ $X2=4.215 $Y2=0.26
r120 89 90 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r121 85 86 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r122 83 86 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r123 82 83 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r124 80 102 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=0 $X2=8.88
+ $Y2=0
r125 80 99 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=0 $X2=7.92
+ $Y2=0
r126 79 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r127 77 98 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.135 $Y=0 $X2=7.97
+ $Y2=0
r128 77 79 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=8.135 $Y=0 $X2=8.4
+ $Y2=0
r129 76 101 4.62176 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=8.675 $Y=0
+ $X2=8.897 $Y2=0
r130 76 79 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=8.675 $Y=0 $X2=8.4
+ $Y2=0
r131 75 99 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0 $X2=7.92
+ $Y2=0
r132 75 96 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0 $X2=6.96
+ $Y2=0
r133 74 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r134 72 95 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.275 $Y=0 $X2=7.11
+ $Y2=0
r135 72 74 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=7.275 $Y=0
+ $X2=7.44 $Y2=0
r136 71 98 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.805 $Y=0 $X2=7.97
+ $Y2=0
r137 71 74 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=7.805 $Y=0
+ $X2=7.44 $Y2=0
r138 70 96 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.96
+ $Y2=0
r139 69 70 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6 $Y2=0
r140 67 95 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.945 $Y=0 $X2=7.11
+ $Y2=0
r141 67 69 61.6524 $w=1.68e-07 $l=9.45e-07 $layer=LI1_cond $X=6.945 $Y=0 $X2=6
+ $Y2=0
r142 66 70 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=6
+ $Y2=0
r143 65 66 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r144 62 65 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=4.56 $Y=0 $X2=5.52
+ $Y2=0
r145 60 89 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.38 $Y=0 $X2=4.215
+ $Y2=0
r146 60 62 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=4.38 $Y=0 $X2=4.56
+ $Y2=0
r147 59 90 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=1.68 $Y=0 $X2=4.08
+ $Y2=0
r148 59 86 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r149 58 59 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r150 56 85 8.23795 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=1.48 $Y=0 $X2=1.325
+ $Y2=0
r151 56 58 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=1.48 $Y=0 $X2=1.68
+ $Y2=0
r152 55 89 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.05 $Y=0 $X2=4.215
+ $Y2=0
r153 55 58 154.62 $w=1.68e-07 $l=2.37e-06 $layer=LI1_cond $X=4.05 $Y=0 $X2=1.68
+ $Y2=0
r154 53 66 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.52
+ $Y2=0
r155 53 90 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=4.08
+ $Y2=0
r156 53 62 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r157 51 65 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=5.625 $Y=0
+ $X2=5.52 $Y2=0
r158 51 52 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.625 $Y=0 $X2=5.79
+ $Y2=0
r159 50 69 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=5.955 $Y=0 $X2=6
+ $Y2=0
r160 50 52 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.955 $Y=0 $X2=5.79
+ $Y2=0
r161 46 101 3.06035 $w=3.2e-07 $l=1.11781e-07 $layer=LI1_cond $X=8.835 $Y=0.085
+ $X2=8.897 $Y2=0
r162 46 48 10.6241 $w=3.18e-07 $l=2.95e-07 $layer=LI1_cond $X=8.835 $Y=0.085
+ $X2=8.835 $Y2=0.38
r163 42 98 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.97 $Y=0.085
+ $X2=7.97 $Y2=0
r164 42 44 15.8897 $w=3.28e-07 $l=4.55e-07 $layer=LI1_cond $X=7.97 $Y=0.085
+ $X2=7.97 $Y2=0.54
r165 38 95 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.11 $Y=0.085
+ $X2=7.11 $Y2=0
r166 38 40 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=7.11 $Y=0.085
+ $X2=7.11 $Y2=0.38
r167 34 36 19.2074 $w=3.28e-07 $l=5.5e-07 $layer=LI1_cond $X=5.79 $Y=0.38
+ $X2=5.79 $Y2=0.93
r168 32 52 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.79 $Y=0.085
+ $X2=5.79 $Y2=0
r169 32 34 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=5.79 $Y=0.085
+ $X2=5.79 $Y2=0.38
r170 28 85 0.701276 $w=3.1e-07 $l=8.5e-08 $layer=LI1_cond $X=1.325 $Y=0.085
+ $X2=1.325 $Y2=0
r171 28 30 17.6584 $w=3.08e-07 $l=4.75e-07 $layer=LI1_cond $X=1.325 $Y=0.085
+ $X2=1.325 $Y2=0.56
r172 27 82 4.56433 $w=1.7e-07 $l=2.68e-07 $layer=LI1_cond $X=0.535 $Y=0
+ $X2=0.267 $Y2=0
r173 26 85 8.23795 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=1.17 $Y=0 $X2=1.325
+ $Y2=0
r174 26 27 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=1.17 $Y=0
+ $X2=0.535 $Y2=0
r175 22 82 3.20184 $w=3.3e-07 $l=1.39155e-07 $layer=LI1_cond $X=0.37 $Y=0.085
+ $X2=0.267 $Y2=0
r176 22 24 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=0.37 $Y=0.085
+ $X2=0.37 $Y2=0.535
r177 7 48 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=8.69
+ $Y=0.235 $X2=8.83 $Y2=0.38
r178 6 44 182 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_NDIFF $count=1 $X=7.83
+ $Y=0.235 $X2=7.97 $Y2=0.54
r179 5 40 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=6.985
+ $Y=0.235 $X2=7.11 $Y2=0.38
r180 4 36 182 $w=1.7e-07 $l=8.03959e-07 $layer=licon1_NDIFF $count=1 $X=5.555
+ $Y=0.235 $X2=5.79 $Y2=0.93
r181 4 34 182 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_NDIFF $count=1 $X=5.555
+ $Y=0.235 $X2=5.79 $Y2=0.38
r182 3 92 182 $w=1.7e-07 $l=5.17011e-07 $layer=licon1_NDIFF $count=1 $X=3.96
+ $Y=0.665 $X2=4.215 $Y2=0.26
r183 2 30 182 $w=1.7e-07 $l=2.93428e-07 $layer=licon1_NDIFF $count=1 $X=1.135
+ $Y=0.35 $X2=1.335 $Y2=0.56
r184 1 24 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=0.245
+ $Y=0.35 $X2=0.37 $Y2=0.535
.ends

