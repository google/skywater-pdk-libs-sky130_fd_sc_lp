* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__mux4_2 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
M1000 a_196_125# S0 a_1223_119# VNB nshort w=420000u l=150000u
+  ad=2.289e+11p pd=2.77e+06u as=8.82e+10p ps=1.26e+06u
M1001 a_1381_119# a_859_351# a_196_125# VNB nshort w=420000u l=150000u
+  ad=1.344e+11p pd=1.48e+06u as=0p ps=0u
M1002 X a_110_125# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=3.528e+11p pd=3.08e+06u as=1.7686e+12p ps=1.21e+07u
M1003 a_196_125# a_80_293# a_110_125# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.176e+11p ps=1.4e+06u
M1004 VGND A0 a_1381_119# VNB nshort w=420000u l=150000u
+  ad=1.0748e+12p pd=8.96e+06u as=0p ps=0u
M1005 a_110_125# a_80_293# a_27_125# VPB phighvt w=640000u l=150000u
+  ad=1.792e+11p pd=1.84e+06u as=3.488e+11p ps=3.65e+06u
M1006 a_859_351# S0 VGND VNB nshort w=420000u l=150000u
+  ad=1.617e+11p pd=1.61e+06u as=0p ps=0u
M1007 a_1223_119# A1 VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_859_351# S0 VPWR VPB phighvt w=640000u l=150000u
+  ad=1.696e+11p pd=1.81e+06u as=0p ps=0u
M1009 a_27_125# S0 a_825_119# VNB nshort w=420000u l=150000u
+  ad=2.289e+11p pd=2.77e+06u as=8.82e+10p ps=1.26e+06u
M1010 VPWR A2 a_975_419# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.344e+11p ps=1.7e+06u
M1011 a_983_119# a_859_351# a_27_125# VNB nshort w=420000u l=150000u
+  ad=1.344e+11p pd=1.48e+06u as=0p ps=0u
M1012 a_975_419# S0 a_27_125# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_110_125# S1 a_27_125# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_1400_419# S0 a_196_125# VPB phighvt w=640000u l=150000u
+  ad=2.304e+11p pd=2e+06u as=4.096e+11p ps=3.84e+06u
M1015 X a_110_125# VGND VNB nshort w=840000u l=150000u
+  ad=2.352e+11p pd=2.24e+06u as=0p ps=0u
M1016 VPWR A0 a_1400_419# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_196_125# S1 a_110_125# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_825_119# A3 VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VPWR a_110_125# X VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VGND A2 a_983_119# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_817_419# A3 VPWR VPB phighvt w=640000u l=150000u
+  ad=1.344e+11p pd=1.7e+06u as=0p ps=0u
M1022 a_1223_419# A1 VPWR VPB phighvt w=640000u l=150000u
+  ad=1.344e+11p pd=1.7e+06u as=0p ps=0u
M1023 VGND S1 a_80_293# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.709e+11p ps=1.66e+06u
M1024 VGND a_110_125# X VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 VPWR S1 a_80_293# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=2.029e+11p ps=2e+06u
M1026 a_27_125# a_859_351# a_817_419# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_196_125# a_859_351# a_1223_419# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
