* NGSPICE file created from sky130_fd_sc_lp__a21bo_1.ext - technology: sky130A

.subckt sky130_fd_sc_lp__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
M1000 a_436_367# A2 VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=6.867e+11p pd=6.13e+06u as=8.589e+11p ps=6.55e+06u
M1001 a_436_367# a_237_367# a_80_43# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=3.339e+11p ps=3.05e+06u
M1002 a_237_367# B1_N VGND VNB nshort w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=8.651e+11p ps=7.38e+06u
M1003 a_556_47# A1 a_80_43# VNB nshort w=840000u l=150000u
+  ad=1.764e+11p pd=2.1e+06u as=3.78e+11p ps=2.58e+06u
M1004 VPWR A1 a_436_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VGND a_80_43# X VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=2.226e+11p ps=2.21e+06u
M1006 a_237_367# B1_N VPWR VPB phighvt w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1007 a_80_43# a_237_367# VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND A2 a_556_47# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR a_80_43# X VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=3.339e+11p ps=3.05e+06u
.ends

