* File: sky130_fd_sc_lp__ebufn_2.pex.spice
* Created: Wed Sep  2 09:50:45 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__EBUFN_2%A_96_21# 1 2 9 13 17 21 23 29 30 31 32 34 38
+ 39 43 45 52
c112 43 0 2.1839e-19 $X=4.035 $Y=2.525
c113 34 0 1.5751e-19 $X=4.035 $Y=2.615
c114 13 0 5.23685e-20 $X=0.555 $Y=2.465
r115 51 52 1.74861 $w=3.3e-07 $l=1e-08 $layer=POLY_cond $X=0.985 $Y=1.46
+ $X2=0.995 $Y2=1.46
r116 45 47 10.5766 $w=3.63e-07 $l=2.3e-07 $layer=LI1_cond $X=4.052 $Y=0.905
+ $X2=4.052 $Y2=1.135
r117 39 41 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=3.08 $Y=2.53
+ $X2=3.08 $Y2=2.7
r118 38 43 3.29812 $w=2.85e-07 $l=1.53542e-07 $layer=LI1_cond $X=4.15 $Y=2.435
+ $X2=4.035 $Y2=2.525
r119 38 47 84.8128 $w=1.68e-07 $l=1.3e-06 $layer=LI1_cond $X=4.15 $Y=2.435
+ $X2=4.15 $Y2=1.135
r120 34 43 3.29812 $w=2.85e-07 $l=9e-08 $layer=LI1_cond $X=4.035 $Y=2.615
+ $X2=4.035 $Y2=2.525
r121 34 36 4.27 $w=4e-07 $l=1.4e-07 $layer=LI1_cond $X=4.035 $Y=2.615 $X2=4.035
+ $Y2=2.755
r122 33 39 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.165 $Y=2.53
+ $X2=3.08 $Y2=2.53
r123 32 43 3.25423 $w=1.7e-07 $l=2.02485e-07 $layer=LI1_cond $X=3.835 $Y=2.53
+ $X2=4.035 $Y2=2.525
r124 32 33 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.835 $Y=2.53
+ $X2=3.165 $Y2=2.53
r125 30 41 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.995 $Y=2.7
+ $X2=3.08 $Y2=2.7
r126 30 31 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=2.995 $Y=2.7
+ $X2=2.485 $Y2=2.7
r127 29 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.4 $Y=2.615
+ $X2=2.485 $Y2=2.7
r128 28 29 64.5882 $w=1.68e-07 $l=9.9e-07 $layer=LI1_cond $X=2.4 $Y=1.625
+ $X2=2.4 $Y2=2.615
r129 26 51 13.9889 $w=3.3e-07 $l=8e-08 $layer=POLY_cond $X=0.905 $Y=1.46
+ $X2=0.985 $Y2=1.46
r130 26 48 61.2015 $w=3.3e-07 $l=3.5e-07 $layer=POLY_cond $X=0.905 $Y=1.46
+ $X2=0.555 $Y2=1.46
r131 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.905
+ $Y=1.46 $X2=0.905 $Y2=1.46
r132 23 28 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.315 $Y=1.46
+ $X2=2.4 $Y2=1.625
r133 23 25 49.2407 $w=3.28e-07 $l=1.41e-06 $layer=LI1_cond $X=2.315 $Y=1.46
+ $X2=0.905 $Y2=1.46
r134 19 52 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.995 $Y=1.295
+ $X2=0.995 $Y2=1.46
r135 19 21 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=0.995 $Y=1.295
+ $X2=0.995 $Y2=0.655
r136 15 51 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.985 $Y=1.625
+ $X2=0.985 $Y2=1.46
r137 15 17 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=0.985 $Y=1.625
+ $X2=0.985 $Y2=2.465
r138 11 48 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.555 $Y=1.625
+ $X2=0.555 $Y2=1.46
r139 11 13 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=0.555 $Y=1.625
+ $X2=0.555 $Y2=2.465
r140 7 48 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.555 $Y=1.295
+ $X2=0.555 $Y2=1.46
r141 7 9 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=0.555 $Y=1.295
+ $X2=0.555 $Y2=0.655
r142 2 36 600 $w=1.7e-07 $l=3.63318e-07 $layer=licon1_PDIFF $count=1 $X=3.86
+ $Y=2.455 $X2=4 $Y2=2.755
r143 1 45 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=3.895
+ $Y=0.695 $X2=4.035 $Y2=0.905
.ends

.subckt PM_SKY130_FD_SC_LP__EBUFN_2%A_284_21# 1 2 7 9 10 11 12 14 15 18 19 21 24
+ 27 28 32
c67 28 0 3.60707e-20 $X=2.77 $Y=0.42
c68 15 0 3.28377e-20 $X=2.605 $Y=1.26
c69 10 0 8.61933e-20 $X=1.92 $Y=1.26
c70 7 0 2.02596e-19 $X=1.495 $Y=1.185
r71 32 33 10.3486 $w=5.43e-07 $l=1.9e-07 $layer=LI1_cond $X=2.927 $Y=0.945
+ $X2=2.927 $Y2=1.135
r72 28 36 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.77 $Y=0.42
+ $X2=2.77 $Y2=0.585
r73 27 30 3.31686 $w=5.93e-07 $l=1.65e-07 $layer=LI1_cond $X=2.902 $Y=0.42
+ $X2=2.902 $Y2=0.585
r74 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.77
+ $Y=0.42 $X2=2.77 $Y2=0.42
r75 24 33 74.7005 $w=1.68e-07 $l=1.145e-06 $layer=LI1_cond $X=2.74 $Y=2.28
+ $X2=2.74 $Y2=1.135
r76 21 32 1.7996 $w=5.43e-07 $l=8.2e-08 $layer=LI1_cond $X=2.927 $Y=0.863
+ $X2=2.927 $Y2=0.945
r77 21 30 6.1011 $w=5.43e-07 $l=2.78e-07 $layer=LI1_cond $X=2.927 $Y=0.863
+ $X2=2.927 $Y2=0.585
r78 18 36 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=2.68 $Y=1.185 $X2=2.68
+ $Y2=0.585
r79 16 19 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.07 $Y=1.26
+ $X2=1.995 $Y2=1.26
r80 15 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.605 $Y=1.26
+ $X2=2.68 $Y2=1.185
r81 15 16 274.33 $w=1.5e-07 $l=5.35e-07 $layer=POLY_cond $X=2.605 $Y=1.26
+ $X2=2.07 $Y2=1.26
r82 12 19 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.995 $Y=1.185
+ $X2=1.995 $Y2=1.26
r83 12 14 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.995 $Y=1.185
+ $X2=1.995 $Y2=0.655
r84 10 19 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.92 $Y=1.26
+ $X2=1.995 $Y2=1.26
r85 10 11 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=1.92 $Y=1.26
+ $X2=1.57 $Y2=1.26
r86 7 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.495 $Y=1.185
+ $X2=1.57 $Y2=1.26
r87 7 9 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.495 $Y=1.185
+ $X2=1.495 $Y2=0.655
r88 2 24 600 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=2.595
+ $Y=2.135 $X2=2.74 $Y2=2.28
r89 1 32 182 $w=1.7e-07 $l=3.14245e-07 $layer=licon1_NDIFF $count=1 $X=2.89
+ $Y=0.695 $X2=3.035 $Y2=0.945
.ends

.subckt PM_SKY130_FD_SC_LP__EBUFN_2%TE_B 1 3 4 5 6 8 9 13 17 19 20 21 25 26
c82 26 0 3.28377e-20 $X=3.16 $Y=1.47
c83 13 0 1.99516e-19 $X=3.07 $Y=2.455
c84 5 0 7.3439e-20 $X=1.49 $Y=1.65
r85 28 29 74.1893 $w=3.3e-07 $l=3.25e-07 $layer=POLY_cond $X=3.16 $Y=1.65
+ $X2=3.16 $Y2=1.975
r86 25 28 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=3.16 $Y=1.47 $X2=3.16
+ $Y2=1.65
r87 25 27 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.16 $Y=1.47
+ $X2=3.16 $Y2=1.305
r88 25 26 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.16
+ $Y=1.47 $X2=3.16 $Y2=1.47
r89 20 21 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=3.16 $Y=1.665
+ $X2=3.16 $Y2=2.035
r90 20 26 6.80989 $w=3.28e-07 $l=1.95e-07 $layer=LI1_cond $X=3.16 $Y=1.665
+ $X2=3.16 $Y2=1.47
r91 17 27 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=3.25 $Y=0.905 $X2=3.25
+ $Y2=1.305
r92 13 29 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=3.07 $Y=2.455
+ $X2=3.07 $Y2=1.975
r93 10 19 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.92 $Y=1.65
+ $X2=1.845 $Y2=1.65
r94 9 28 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.995 $Y=1.65
+ $X2=3.16 $Y2=1.65
r95 9 10 551.223 $w=1.5e-07 $l=1.075e-06 $layer=POLY_cond $X=2.995 $Y=1.65
+ $X2=1.92 $Y2=1.65
r96 6 19 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.845 $Y=1.725
+ $X2=1.845 $Y2=1.65
r97 6 8 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=1.845 $Y=1.725
+ $X2=1.845 $Y2=2.465
r98 4 19 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.77 $Y=1.65
+ $X2=1.845 $Y2=1.65
r99 4 5 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=1.77 $Y=1.65 $X2=1.49
+ $Y2=1.65
r100 1 5 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.415 $Y=1.725
+ $X2=1.49 $Y2=1.65
r101 1 3 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=1.415 $Y=1.725
+ $X2=1.415 $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__EBUFN_2%A 3 7 11 12 13 14 18 19
c36 12 0 1.76383e-19 $X=3.73 $Y=1.975
r37 18 19 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.73
+ $Y=1.47 $X2=3.73 $Y2=1.47
r38 13 14 10.9334 $w=3.88e-07 $l=3.7e-07 $layer=LI1_cond $X=3.7 $Y=1.665 $X2=3.7
+ $Y2=2.035
r39 13 19 5.76222 $w=3.88e-07 $l=1.95e-07 $layer=LI1_cond $X=3.7 $Y=1.665
+ $X2=3.7 $Y2=1.47
r40 11 18 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=3.73 $Y=1.81
+ $X2=3.73 $Y2=1.47
r41 11 12 41.3509 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.73 $Y=1.81
+ $X2=3.73 $Y2=1.975
r42 10 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.73 $Y=1.305
+ $X2=3.73 $Y2=1.47
r43 7 10 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=3.82 $Y=0.905 $X2=3.82
+ $Y2=1.305
r44 3 12 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=3.785 $Y=2.775
+ $X2=3.785 $Y2=1.975
.ends

.subckt PM_SKY130_FD_SC_LP__EBUFN_2%A_39_367# 1 2 3 10 12 14 16 17 18 20 22
c52 20 0 1.38309e-20 $X=2.02 $Y=1.985
c53 18 0 7.23624e-20 $X=1.895 $Y=1.9
c54 16 0 5.23685e-20 $X=1.2 $Y=1.985
r55 20 31 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.02 $Y=1.985
+ $X2=2.02 $Y2=1.9
r56 20 22 42.6404 $w=2.48e-07 $l=9.25e-07 $layer=LI1_cond $X=2.02 $Y=1.985
+ $X2=2.02 $Y2=2.91
r57 19 27 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.365 $Y=1.9 $X2=1.2
+ $Y2=1.9
r58 18 31 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.895 $Y=1.9
+ $X2=2.02 $Y2=1.9
r59 18 19 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=1.895 $Y=1.9
+ $X2=1.365 $Y2=1.9
r60 17 29 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.2 $Y=2.905 $X2=1.2
+ $Y2=2.99
r61 16 27 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.2 $Y=1.985 $X2=1.2
+ $Y2=1.9
r62 16 17 32.1287 $w=3.28e-07 $l=9.2e-07 $layer=LI1_cond $X=1.2 $Y=1.985 $X2=1.2
+ $Y2=2.905
r63 15 25 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.505 $Y=2.99
+ $X2=0.34 $Y2=2.99
r64 14 29 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.035 $Y=2.99
+ $X2=1.2 $Y2=2.99
r65 14 15 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=1.035 $Y=2.99
+ $X2=0.505 $Y2=2.99
r66 10 25 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.34 $Y=2.905 $X2=0.34
+ $Y2=2.99
r67 10 12 23.9219 $w=3.28e-07 $l=6.85e-07 $layer=LI1_cond $X=0.34 $Y=2.905
+ $X2=0.34 $Y2=2.22
r68 3 31 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.92
+ $Y=1.835 $X2=2.06 $Y2=1.98
r69 3 22 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=1.92
+ $Y=1.835 $X2=2.06 $Y2=2.91
r70 2 29 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=1.06
+ $Y=1.835 $X2=1.2 $Y2=2.91
r71 2 27 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.06
+ $Y=1.835 $X2=1.2 $Y2=1.98
r72 1 25 400 $w=1.7e-07 $l=1.18528e-06 $layer=licon1_PDIFF $count=1 $X=0.195
+ $Y=1.835 $X2=0.34 $Y2=2.95
r73 1 12 400 $w=1.7e-07 $l=4.51719e-07 $layer=licon1_PDIFF $count=1 $X=0.195
+ $Y=1.835 $X2=0.34 $Y2=2.22
.ends

.subckt PM_SKY130_FD_SC_LP__EBUFN_2%Z 1 2 7 8 9 10 13 17 21 22
c35 13 0 1.40359e-19 $X=0.78 $Y=0.805
c36 7 0 6.22368e-20 $X=0.615 $Y=1.04
r37 21 22 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.24 $Y=1.295
+ $X2=0.24 $Y2=1.665
r38 20 22 6.51381 $w=2.28e-07 $l=1.3e-07 $layer=LI1_cond $X=0.24 $Y=1.795
+ $X2=0.24 $Y2=1.665
r39 19 21 8.51806 $w=2.28e-07 $l=1.7e-07 $layer=LI1_cond $X=0.24 $Y=1.125
+ $X2=0.24 $Y2=1.295
r40 15 17 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=0.77 $Y=1.965
+ $X2=0.77 $Y2=1.98
r41 11 13 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=0.78 $Y=0.955
+ $X2=0.78 $Y2=0.805
r42 10 20 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=0.355 $Y=1.88
+ $X2=0.24 $Y2=1.795
r43 9 15 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.685 $Y=1.88
+ $X2=0.77 $Y2=1.965
r44 9 10 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=0.685 $Y=1.88
+ $X2=0.355 $Y2=1.88
r45 8 19 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=0.355 $Y=1.04
+ $X2=0.24 $Y2=1.125
r46 7 11 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.615 $Y=1.04
+ $X2=0.78 $Y2=0.955
r47 7 8 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=0.615 $Y=1.04
+ $X2=0.355 $Y2=1.04
r48 2 17 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=0.63
+ $Y=1.835 $X2=0.77 $Y2=1.98
r49 1 13 182 $w=1.7e-07 $l=6.40625e-07 $layer=licon1_NDIFF $count=1 $X=0.63
+ $Y=0.235 $X2=0.78 $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_LP__EBUFN_2%VPWR 1 2 9 13 16 17 18 20 33 34 37
r54 37 38 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r55 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r56 31 34 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=4.08 $Y2=3.33
r57 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r58 28 37 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.715 $Y=3.33
+ $X2=1.63 $Y2=3.33
r59 28 30 91.6631 $w=1.68e-07 $l=1.405e-06 $layer=LI1_cond $X=1.715 $Y=3.33
+ $X2=3.12 $Y2=3.33
r60 27 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r61 26 27 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r62 23 27 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.2 $Y2=3.33
r63 22 26 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.24 $Y=3.33 $X2=1.2
+ $Y2=3.33
r64 22 23 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r65 20 37 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.545 $Y=3.33
+ $X2=1.63 $Y2=3.33
r66 20 26 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.545 $Y=3.33
+ $X2=1.2 $Y2=3.33
r67 18 31 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r68 18 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r69 16 30 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=3.335 $Y=3.33
+ $X2=3.12 $Y2=3.33
r70 16 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.335 $Y=3.33
+ $X2=3.5 $Y2=3.33
r71 15 33 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=3.665 $Y=3.33
+ $X2=4.08 $Y2=3.33
r72 15 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.665 $Y=3.33
+ $X2=3.5 $Y2=3.33
r73 11 17 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.5 $Y=3.245 $X2=3.5
+ $Y2=3.33
r74 11 13 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=3.5 $Y=3.245
+ $X2=3.5 $Y2=2.95
r75 7 37 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.63 $Y=3.245 $X2=1.63
+ $Y2=3.33
r76 7 9 60.3476 $w=1.68e-07 $l=9.25e-07 $layer=LI1_cond $X=1.63 $Y=3.245
+ $X2=1.63 $Y2=2.32
r77 2 13 600 $w=1.7e-07 $l=9.76499e-07 $layer=licon1_PDIFF $count=1 $X=3.145
+ $Y=2.135 $X2=3.5 $Y2=2.95
r78 1 9 300 $w=1.7e-07 $l=5.50568e-07 $layer=licon1_PDIFF $count=2 $X=1.49
+ $Y=1.835 $X2=1.63 $Y2=2.32
.ends

.subckt PM_SKY130_FD_SC_LP__EBUFN_2%A_27_47# 1 2 3 12 14 15 16 17 18 19 22
c49 18 0 7.3439e-20 $X=2.045 $Y=1.04
r50 20 22 18.6835 $w=3.28e-07 $l=5.35e-07 $layer=LI1_cond $X=2.21 $Y=0.955
+ $X2=2.21 $Y2=0.42
r51 18 20 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.045 $Y=1.04
+ $X2=2.21 $Y2=0.955
r52 18 19 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=2.045 $Y=1.04
+ $X2=1.445 $Y2=1.04
r53 17 19 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.28 $Y=0.955
+ $X2=1.445 $Y2=1.04
r54 16 25 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.28 $Y=0.425 $X2=1.28
+ $Y2=0.34
r55 16 17 18.5089 $w=3.28e-07 $l=5.3e-07 $layer=LI1_cond $X=1.28 $Y=0.425
+ $X2=1.28 $Y2=0.955
r56 14 25 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.115 $Y=0.34
+ $X2=1.28 $Y2=0.34
r57 14 15 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.115 $Y=0.34
+ $X2=0.445 $Y2=0.34
r58 10 15 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.28 $Y=0.425
+ $X2=0.445 $Y2=0.34
r59 10 12 4.01609 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=0.28 $Y=0.425
+ $X2=0.28 $Y2=0.54
r60 3 22 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=2.07
+ $Y=0.235 $X2=2.21 $Y2=0.42
r61 2 25 91 $w=1.7e-07 $l=2.8801e-07 $layer=licon1_NDIFF $count=2 $X=1.07
+ $Y=0.235 $X2=1.28 $Y2=0.42
r62 1 12 182 $w=1.7e-07 $l=3.70473e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.28 $Y2=0.54
.ends

.subckt PM_SKY130_FD_SC_LP__EBUFN_2%VGND 1 2 9 13 15 17 22 32 33 36 39
c48 33 0 3.60707e-20 $X=4.08 $Y=0
r49 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r50 36 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r51 33 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.6
+ $Y2=0
r52 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r53 30 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.7 $Y=0 $X2=3.535
+ $Y2=0
r54 30 32 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=3.7 $Y=0 $X2=4.08
+ $Y2=0
r55 29 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r56 28 29 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r57 25 28 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r58 23 36 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.875 $Y=0 $X2=1.75
+ $Y2=0
r59 23 25 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.875 $Y=0 $X2=2.16
+ $Y2=0
r60 22 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.37 $Y=0 $X2=3.535
+ $Y2=0
r61 22 28 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=3.37 $Y=0 $X2=3.12
+ $Y2=0
r62 20 37 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=0.24 $Y=0 $X2=1.68
+ $Y2=0
r63 19 20 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r64 17 36 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.625 $Y=0 $X2=1.75
+ $Y2=0
r65 17 19 90.3583 $w=1.68e-07 $l=1.385e-06 $layer=LI1_cond $X=1.625 $Y=0
+ $X2=0.24 $Y2=0
r66 15 29 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r67 15 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.68
+ $Y2=0
r68 15 25 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r69 11 39 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.535 $Y=0.085
+ $X2=3.535 $Y2=0
r70 11 13 28.6365 $w=3.28e-07 $l=8.2e-07 $layer=LI1_cond $X=3.535 $Y=0.085
+ $X2=3.535 $Y2=0.905
r71 7 36 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.75 $Y=0.085
+ $X2=1.75 $Y2=0
r72 7 9 19.1306 $w=2.48e-07 $l=4.15e-07 $layer=LI1_cond $X=1.75 $Y=0.085
+ $X2=1.75 $Y2=0.5
r73 2 13 182 $w=1.7e-07 $l=2.96985e-07 $layer=licon1_NDIFF $count=1 $X=3.325
+ $Y=0.695 $X2=3.535 $Y2=0.905
r74 1 9 182 $w=1.7e-07 $l=3.27605e-07 $layer=licon1_NDIFF $count=1 $X=1.57
+ $Y=0.235 $X2=1.71 $Y2=0.5
.ends

