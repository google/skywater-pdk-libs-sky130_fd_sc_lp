* File: sky130_fd_sc_lp__a21boi_2.pex.spice
* Created: Fri Aug 28 09:50:08 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A21BOI_2%B1_N 3 5 6 7 9 12 13 14 15 16 17 18 26
r35 26 27 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.385
+ $Y=1.02 $X2=0.385 $Y2=1.02
r36 17 18 11.0754 $w=3.83e-07 $l=3.7e-07 $layer=LI1_cond $X=0.277 $Y=2.035
+ $X2=0.277 $Y2=2.405
r37 16 17 11.0754 $w=3.83e-07 $l=3.7e-07 $layer=LI1_cond $X=0.277 $Y=1.665
+ $X2=0.277 $Y2=2.035
r38 15 16 11.0754 $w=3.83e-07 $l=3.7e-07 $layer=LI1_cond $X=0.277 $Y=1.295
+ $X2=0.277 $Y2=1.665
r39 15 27 8.23174 $w=3.83e-07 $l=2.75e-07 $layer=LI1_cond $X=0.277 $Y=1.295
+ $X2=0.277 $Y2=1.02
r40 14 27 2.84369 $w=3.83e-07 $l=9.5e-08 $layer=LI1_cond $X=0.277 $Y=0.925
+ $X2=0.277 $Y2=1.02
r41 13 14 11.0754 $w=3.83e-07 $l=3.7e-07 $layer=LI1_cond $X=0.277 $Y=0.555
+ $X2=0.277 $Y2=0.925
r42 11 26 47.1618 $w=3.75e-07 $l=3.18e-07 $layer=POLY_cond $X=0.407 $Y=1.338
+ $X2=0.407 $Y2=1.02
r43 11 12 48.4185 $w=3.75e-07 $l=1.87e-07 $layer=POLY_cond $X=0.407 $Y=1.338
+ $X2=0.407 $Y2=1.525
r44 10 26 2.22462 $w=3.75e-07 $l=1.5e-08 $layer=POLY_cond $X=0.407 $Y=1.005
+ $X2=0.407 $Y2=1.02
r45 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.97 $Y=0.855 $X2=0.97
+ $Y2=0.535
r46 6 10 33.9315 $w=1.5e-07 $l=2.2236e-07 $layer=POLY_cond $X=0.595 $Y=0.93
+ $X2=0.407 $Y2=1.005
r47 5 7 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.895 $Y=0.93
+ $X2=0.97 $Y2=0.855
r48 5 6 153.83 $w=1.5e-07 $l=3e-07 $layer=POLY_cond $X=0.895 $Y=0.93 $X2=0.595
+ $Y2=0.93
r49 3 12 607.628 $w=1.5e-07 $l=1.185e-06 $layer=POLY_cond $X=0.52 $Y=2.71
+ $X2=0.52 $Y2=1.525
.ends

.subckt PM_SKY130_FD_SC_LP__A21BOI_2%A_119_500# 1 2 7 9 11 14 16 18 20 23 25 26
+ 29 33 39 42
c77 42 0 1.90917e-19 $X=1 $Y=1.35
c78 18 0 6.82747e-20 $X=1.925 $Y=1.275
r79 40 42 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=1 $Y=1.44 $X2=1
+ $Y2=1.35
r80 39 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1 $Y=1.44
+ $X2=1 $Y2=1.44
r81 31 35 0.83239 $w=2.6e-07 $l=1.33e-07 $layer=LI1_cond $X=0.77 $Y=1.605
+ $X2=0.77 $Y2=1.472
r82 31 33 48.9788 $w=2.58e-07 $l=1.105e-06 $layer=LI1_cond $X=0.77 $Y=1.605
+ $X2=0.77 $Y2=2.71
r83 27 39 9.56745 $w=2.63e-07 $l=2.2e-07 $layer=LI1_cond $X=0.78 $Y=1.472 $X2=1
+ $Y2=1.472
r84 27 35 0.434884 $w=2.63e-07 $l=1e-08 $layer=LI1_cond $X=0.78 $Y=1.472
+ $X2=0.77 $Y2=1.472
r85 27 29 33.1327 $w=2.78e-07 $l=8.05e-07 $layer=LI1_cond $X=0.78 $Y=1.34
+ $X2=0.78 $Y2=0.535
r86 21 26 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.925 $Y=1.425
+ $X2=1.925 $Y2=1.35
r87 21 23 533.277 $w=1.5e-07 $l=1.04e-06 $layer=POLY_cond $X=1.925 $Y=1.425
+ $X2=1.925 $Y2=2.465
r88 18 26 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.925 $Y=1.275
+ $X2=1.925 $Y2=1.35
r89 18 20 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.925 $Y=1.275
+ $X2=1.925 $Y2=0.745
r90 17 25 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.57 $Y=1.35 $X2=1.495
+ $Y2=1.35
r91 16 26 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.85 $Y=1.35
+ $X2=1.925 $Y2=1.35
r92 16 17 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=1.85 $Y=1.35
+ $X2=1.57 $Y2=1.35
r93 12 25 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.495 $Y=1.425
+ $X2=1.495 $Y2=1.35
r94 12 14 533.277 $w=1.5e-07 $l=1.04e-06 $layer=POLY_cond $X=1.495 $Y=1.425
+ $X2=1.495 $Y2=2.465
r95 9 25 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.495 $Y=1.275 $X2=1.495
+ $Y2=1.35
r96 9 11 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.495 $Y=1.275
+ $X2=1.495 $Y2=0.745
r97 8 42 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.165 $Y=1.35 $X2=1
+ $Y2=1.35
r98 7 25 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.42 $Y=1.35 $X2=1.495
+ $Y2=1.35
r99 7 8 130.755 $w=1.5e-07 $l=2.55e-07 $layer=POLY_cond $X=1.42 $Y=1.35
+ $X2=1.165 $Y2=1.35
r100 2 33 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=0.595
+ $Y=2.5 $X2=0.735 $Y2=2.71
r101 1 29 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.63
+ $Y=0.325 $X2=0.755 $Y2=0.535
.ends

.subckt PM_SKY130_FD_SC_LP__A21BOI_2%A2 3 7 11 15 18 20 23 25 30 31 33 34 35 50
c93 3 0 3.15539e-19 $X=2.355 $Y=2.465
r94 48 50 2.55944 $w=1.93e-07 $l=4.5e-08 $layer=LI1_cond $X=2.595 $Y=2.022
+ $X2=2.64 $Y2=2.022
r95 34 35 14.9567 $w=3.63e-07 $l=3.95e-07 $layer=LI1_cond $X=3.12 $Y=2.022
+ $X2=3.515 $Y2=2.022
r96 33 48 3.20299 $w=1.95e-07 $l=8.5e-08 $layer=LI1_cond $X=2.51 $Y=2.022
+ $X2=2.595 $Y2=2.022
r97 33 34 26.1632 $w=1.93e-07 $l=4.6e-07 $layer=LI1_cond $X=2.66 $Y=2.022
+ $X2=3.12 $Y2=2.022
r98 33 50 1.13753 $w=1.93e-07 $l=2e-08 $layer=LI1_cond $X=2.66 $Y=2.022 $X2=2.64
+ $Y2=2.022
r99 31 46 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.895 $Y=1.51
+ $X2=3.895 $Y2=1.675
r100 31 45 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.895 $Y=1.51
+ $X2=3.895 $Y2=1.345
r101 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.895
+ $Y=1.51 $X2=3.895 $Y2=1.51
r102 27 30 10.5309 $w=2.88e-07 $l=2.65e-07 $layer=LI1_cond $X=3.63 $Y=1.5
+ $X2=3.895 $Y2=1.5
r103 23 43 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.415 $Y=1.51
+ $X2=2.415 $Y2=1.675
r104 23 42 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.415 $Y=1.51
+ $X2=2.415 $Y2=1.345
r105 22 25 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=2.415 $Y=1.51
+ $X2=2.51 $Y2=1.51
r106 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.415
+ $Y=1.51 $X2=2.415 $Y2=1.51
r107 20 35 3.14646 $w=2.3e-07 $l=9.7e-08 $layer=LI1_cond $X=3.63 $Y=1.925
+ $X2=3.63 $Y2=2.022
r108 19 27 2.09727 $w=2.3e-07 $l=1.45e-07 $layer=LI1_cond $X=3.63 $Y=1.645
+ $X2=3.63 $Y2=1.5
r109 19 20 14.0297 $w=2.28e-07 $l=2.8e-07 $layer=LI1_cond $X=3.63 $Y=1.645
+ $X2=3.63 $Y2=1.925
r110 18 33 3.65518 $w=1.7e-07 $l=9.7e-08 $layer=LI1_cond $X=2.51 $Y=1.925
+ $X2=2.51 $Y2=2.022
r111 17 25 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.51 $Y=1.595
+ $X2=2.51 $Y2=1.51
r112 17 18 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=2.51 $Y=1.595
+ $X2=2.51 $Y2=1.925
r113 15 46 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.805 $Y=2.465
+ $X2=3.805 $Y2=1.675
r114 11 45 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=3.805 $Y=0.745
+ $X2=3.805 $Y2=1.345
r115 7 42 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=2.435 $Y=0.745
+ $X2=2.435 $Y2=1.345
r116 3 43 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.355 $Y=2.465
+ $X2=2.355 $Y2=1.675
.ends

.subckt PM_SKY130_FD_SC_LP__A21BOI_2%A1 3 7 11 15 17 25
r57 23 25 73.4417 $w=3.3e-07 $l=4.2e-07 $layer=POLY_cond $X=2.955 $Y=1.51
+ $X2=3.375 $Y2=1.51
r58 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.955
+ $Y=1.51 $X2=2.955 $Y2=1.51
r59 21 23 1.74861 $w=3.3e-07 $l=1e-08 $layer=POLY_cond $X=2.945 $Y=1.51
+ $X2=2.955 $Y2=1.51
r60 19 21 13.9889 $w=3.3e-07 $l=8e-08 $layer=POLY_cond $X=2.865 $Y=1.51
+ $X2=2.945 $Y2=1.51
r61 17 24 5.85086 $w=3.23e-07 $l=1.65e-07 $layer=LI1_cond $X=3.12 $Y=1.587
+ $X2=2.955 $Y2=1.587
r62 13 25 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.375 $Y=1.675
+ $X2=3.375 $Y2=1.51
r63 13 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.375 $Y=1.675
+ $X2=3.375 $Y2=2.465
r64 9 25 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.375 $Y=1.345
+ $X2=3.375 $Y2=1.51
r65 9 11 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=3.375 $Y=1.345 $X2=3.375
+ $Y2=0.745
r66 5 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.945 $Y=1.675
+ $X2=2.945 $Y2=1.51
r67 5 7 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.945 $Y=1.675
+ $X2=2.945 $Y2=2.465
r68 1 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.865 $Y=1.345
+ $X2=2.865 $Y2=1.51
r69 1 3 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=2.865 $Y=1.345 $X2=2.865
+ $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_LP__A21BOI_2%VPWR 1 2 3 10 12 16 20 22 24 32 39 40 46 49
r58 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r59 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r60 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r61 40 50 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.6 $Y2=3.33
r62 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r63 37 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.755 $Y=3.33
+ $X2=3.59 $Y2=3.33
r64 37 39 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=3.755 $Y=3.33
+ $X2=4.08 $Y2=3.33
r65 36 50 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r66 36 47 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.64 $Y2=3.33
r67 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r68 33 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.815 $Y=3.33
+ $X2=2.65 $Y2=3.33
r69 33 35 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.815 $Y=3.33
+ $X2=3.12 $Y2=3.33
r70 32 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.425 $Y=3.33
+ $X2=3.59 $Y2=3.33
r71 32 35 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3.425 $Y=3.33
+ $X2=3.12 $Y2=3.33
r72 28 44 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r73 27 30 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=0.72 $Y=3.33
+ $X2=2.16 $Y2=3.33
r74 27 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r75 25 43 4.67962 $w=1.7e-07 $l=2.35e-07 $layer=LI1_cond $X=0.47 $Y=3.33
+ $X2=0.235 $Y2=3.33
r76 25 27 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=0.47 $Y=3.33
+ $X2=0.72 $Y2=3.33
r77 24 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.485 $Y=3.33
+ $X2=2.65 $Y2=3.33
r78 24 30 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=2.485 $Y=3.33
+ $X2=2.16 $Y2=3.33
r79 22 47 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r80 22 28 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=0.72 $Y2=3.33
r81 22 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r82 18 49 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.59 $Y=3.245
+ $X2=3.59 $Y2=3.33
r83 18 20 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=3.59 $Y=3.245
+ $X2=3.59 $Y2=2.765
r84 14 46 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.65 $Y=3.245
+ $X2=2.65 $Y2=3.33
r85 14 16 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=2.65 $Y=3.245
+ $X2=2.65 $Y2=2.78
r86 10 43 3.08656 $w=3.3e-07 $l=1.14782e-07 $layer=LI1_cond $X=0.305 $Y=3.245
+ $X2=0.235 $Y2=3.33
r87 10 12 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=0.305 $Y=3.245
+ $X2=0.305 $Y2=2.765
r88 3 20 600 $w=1.7e-07 $l=9.97547e-07 $layer=licon1_PDIFF $count=1 $X=3.45
+ $Y=1.835 $X2=3.59 $Y2=2.765
r89 2 16 600 $w=1.7e-07 $l=1.04925e-06 $layer=licon1_PDIFF $count=1 $X=2.43
+ $Y=1.835 $X2=2.65 $Y2=2.78
r90 1 12 600 $w=1.7e-07 $l=3.21481e-07 $layer=licon1_PDIFF $count=1 $X=0.18
+ $Y=2.5 $X2=0.305 $Y2=2.765
.ends

.subckt PM_SKY130_FD_SC_LP__A21BOI_2%A_231_367# 1 2 3 4 13 15 17 21 24 25 29 31
+ 35 42 44 46
r64 33 46 3.52026 $w=2.65e-07 $l=8.5e-08 $layer=LI1_cond $X=4.05 $Y=2.29
+ $X2=4.05 $Y2=2.375
r65 33 35 13.2318 $w=2.68e-07 $l=3.1e-07 $layer=LI1_cond $X=4.05 $Y=2.29
+ $X2=4.05 $Y2=1.98
r66 32 44 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=3.255 $Y=2.375
+ $X2=3.12 $Y2=2.375
r67 31 46 2.98021 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=3.915 $Y=2.375
+ $X2=4.05 $Y2=2.375
r68 31 32 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=3.915 $Y=2.375
+ $X2=3.255 $Y2=2.375
r69 27 44 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.12 $Y=2.46
+ $X2=3.12 $Y2=2.375
r70 27 29 14.7257 $w=2.68e-07 $l=3.45e-07 $layer=LI1_cond $X=3.12 $Y=2.46
+ $X2=3.12 $Y2=2.805
r71 26 42 2.53056 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=2.315 $Y=2.375
+ $X2=2.18 $Y2=2.375
r72 25 44 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=2.985 $Y=2.375
+ $X2=3.12 $Y2=2.375
r73 25 26 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.985 $Y=2.375
+ $X2=2.315 $Y2=2.375
r74 23 42 3.91525 $w=2.35e-07 $l=8.5e-08 $layer=LI1_cond $X=2.18 $Y=2.46
+ $X2=2.18 $Y2=2.375
r75 23 24 18.994 $w=2.68e-07 $l=4.45e-07 $layer=LI1_cond $X=2.18 $Y=2.46
+ $X2=2.18 $Y2=2.905
r76 19 42 3.91525 $w=2.35e-07 $l=1.00995e-07 $layer=LI1_cond $X=2.145 $Y=2.29
+ $X2=2.18 $Y2=2.375
r77 19 21 16.3591 $w=1.98e-07 $l=2.95e-07 $layer=LI1_cond $X=2.145 $Y=2.29
+ $X2=2.145 $Y2=1.995
r78 18 40 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.375 $Y=2.99
+ $X2=1.245 $Y2=2.99
r79 17 24 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=2.045 $Y=2.99
+ $X2=2.18 $Y2=2.905
r80 17 18 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.045 $Y=2.99
+ $X2=1.375 $Y2=2.99
r81 13 40 2.85134 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=1.245 $Y=2.905
+ $X2=1.245 $Y2=2.99
r82 13 15 40.3355 $w=2.58e-07 $l=9.1e-07 $layer=LI1_cond $X=1.245 $Y=2.905
+ $X2=1.245 $Y2=1.995
r83 4 46 300 $w=1.7e-07 $l=6.81414e-07 $layer=licon1_PDIFF $count=2 $X=3.88
+ $Y=1.835 $X2=4.02 $Y2=2.45
r84 4 35 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=3.88
+ $Y=1.835 $X2=4.02 $Y2=1.98
r85 3 44 600 $w=1.7e-07 $l=6.0597e-07 $layer=licon1_PDIFF $count=1 $X=3.02
+ $Y=1.835 $X2=3.16 $Y2=2.375
r86 3 29 600 $w=1.7e-07 $l=1.03764e-06 $layer=licon1_PDIFF $count=1 $X=3.02
+ $Y=1.835 $X2=3.16 $Y2=2.805
r87 2 42 300 $w=1.7e-07 $l=6.81414e-07 $layer=licon1_PDIFF $count=2 $X=2
+ $Y=1.835 $X2=2.14 $Y2=2.45
r88 2 21 600 $w=1.7e-07 $l=2.19089e-07 $layer=licon1_PDIFF $count=1 $X=2
+ $Y=1.835 $X2=2.14 $Y2=1.995
r89 1 40 400 $w=1.7e-07 $l=1.13578e-06 $layer=licon1_PDIFF $count=1 $X=1.155
+ $Y=1.835 $X2=1.28 $Y2=2.91
r90 1 15 400 $w=1.7e-07 $l=2.13542e-07 $layer=licon1_PDIFF $count=1 $X=1.155
+ $Y=1.835 $X2=1.28 $Y2=1.995
.ends

.subckt PM_SKY130_FD_SC_LP__A21BOI_2%Y 1 2 3 10 14 16 17 18 19 20 21 32 41 47
c56 47 0 1.56001e-19 $X=1.68 $Y=2.035
c57 41 0 1.90917e-19 $X=1.68 $Y=1.295
c58 20 0 1.59538e-19 $X=1.595 $Y=1.95
c59 18 0 1.37558e-19 $X=1.595 $Y=1.21
r60 45 47 1.74613 $w=3.28e-07 $l=5e-08 $layer=LI1_cond $X=1.71 $Y=1.985 $X2=1.71
+ $Y2=2.035
r61 38 41 2.30489 $w=2.48e-07 $l=5e-08 $layer=LI1_cond $X=1.67 $Y=1.245 $X2=1.67
+ $Y2=1.295
r62 21 52 8.3814 $w=3.28e-07 $l=2.4e-07 $layer=LI1_cond $X=1.71 $Y=2.405
+ $X2=1.71 $Y2=2.645
r63 20 45 0.873063 $w=3.28e-07 $l=2.5e-08 $layer=LI1_cond $X=1.71 $Y=1.96
+ $X2=1.71 $Y2=1.985
r64 20 57 5.59382 $w=3.28e-07 $l=1.4e-07 $layer=LI1_cond $X=1.71 $Y=1.96
+ $X2=1.71 $Y2=1.82
r65 20 21 12.3276 $w=3.28e-07 $l=3.53e-07 $layer=LI1_cond $X=1.71 $Y=2.052
+ $X2=1.71 $Y2=2.405
r66 20 47 0.593683 $w=3.28e-07 $l=1.7e-08 $layer=LI1_cond $X=1.71 $Y=2.052
+ $X2=1.71 $Y2=2.035
r67 19 57 7.14515 $w=2.48e-07 $l=1.55e-07 $layer=LI1_cond $X=1.67 $Y=1.665
+ $X2=1.67 $Y2=1.82
r68 18 30 3.64284 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=1.675 $Y=1.16
+ $X2=1.675 $Y2=1.075
r69 18 38 3.64284 $w=2.55e-07 $l=8.74643e-08 $layer=LI1_cond $X=1.675 $Y=1.16
+ $X2=1.67 $Y2=1.245
r70 18 19 16.2725 $w=2.48e-07 $l=3.53e-07 $layer=LI1_cond $X=1.67 $Y=1.312
+ $X2=1.67 $Y2=1.665
r71 18 41 0.783661 $w=2.48e-07 $l=1.7e-08 $layer=LI1_cond $X=1.67 $Y=1.312
+ $X2=1.67 $Y2=1.295
r72 17 30 6.64871 $w=2.58e-07 $l=1.5e-07 $layer=LI1_cond $X=1.675 $Y=0.925
+ $X2=1.675 $Y2=1.075
r73 16 17 16.4002 $w=2.58e-07 $l=3.7e-07 $layer=LI1_cond $X=1.675 $Y=0.555
+ $X2=1.675 $Y2=0.925
r74 16 32 4.6541 $w=2.58e-07 $l=1.05e-07 $layer=LI1_cond $X=1.675 $Y=0.555
+ $X2=1.675 $Y2=0.45
r75 12 14 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=3.16 $Y=1.075
+ $X2=3.16 $Y2=0.69
r76 11 18 2.83584 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.805 $Y=1.16
+ $X2=1.675 $Y2=1.16
r77 10 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.995 $Y=1.16
+ $X2=3.16 $Y2=1.075
r78 10 11 77.6364 $w=1.68e-07 $l=1.19e-06 $layer=LI1_cond $X=2.995 $Y=1.16
+ $X2=1.805 $Y2=1.16
r79 3 20 400 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=1.57
+ $Y=1.835 $X2=1.71 $Y2=1.96
r80 3 52 400 $w=1.7e-07 $l=8.77211e-07 $layer=licon1_PDIFF $count=1 $X=1.57
+ $Y=1.835 $X2=1.71 $Y2=2.645
r81 2 14 91 $w=1.7e-07 $l=4.62088e-07 $layer=licon1_NDIFF $count=2 $X=2.94
+ $Y=0.325 $X2=3.16 $Y2=0.69
r82 1 32 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=1.57
+ $Y=0.325 $X2=1.71 $Y2=0.45
.ends

.subckt PM_SKY130_FD_SC_LP__A21BOI_2%VGND 1 2 3 12 18 20 22 24 26 31 36 45 48 52
r57 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r58 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r59 43 52 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r60 42 43 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r61 40 43 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r62 39 42 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r63 39 40 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r64 37 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.305 $Y=0 $X2=2.14
+ $Y2=0
r65 37 39 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=2.305 $Y=0 $X2=2.64
+ $Y2=0
r66 36 51 4.36866 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=3.89 $Y=0 $X2=4.105
+ $Y2=0
r67 36 42 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=3.89 $Y=0 $X2=3.6
+ $Y2=0
r68 35 46 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r69 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r70 32 45 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.375 $Y=0 $X2=1.245
+ $Y2=0
r71 32 34 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.375 $Y=0 $X2=1.68
+ $Y2=0
r72 31 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.975 $Y=0 $X2=2.14
+ $Y2=0
r73 31 34 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.975 $Y=0 $X2=1.68
+ $Y2=0
r74 29 46 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r75 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r76 26 45 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.115 $Y=0 $X2=1.245
+ $Y2=0
r77 26 28 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=1.115 $Y=0 $X2=0.72
+ $Y2=0
r78 24 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r79 24 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.68
+ $Y2=0
r80 24 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r81 20 51 3.10886 $w=2.95e-07 $l=1.14039e-07 $layer=LI1_cond $X=4.037 $Y=0.085
+ $X2=4.105 $Y2=0
r82 20 22 15.0404 $w=2.93e-07 $l=3.85e-07 $layer=LI1_cond $X=4.037 $Y=0.085
+ $X2=4.037 $Y2=0.47
r83 16 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.14 $Y=0.085
+ $X2=2.14 $Y2=0
r84 16 18 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=2.14 $Y=0.085
+ $X2=2.14 $Y2=0.45
r85 12 14 23.7137 $w=2.58e-07 $l=5.35e-07 $layer=LI1_cond $X=1.245 $Y=0.47
+ $X2=1.245 $Y2=1.005
r86 10 45 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=1.245 $Y=0.085
+ $X2=1.245 $Y2=0
r87 10 12 17.065 $w=2.58e-07 $l=3.85e-07 $layer=LI1_cond $X=1.245 $Y=0.085
+ $X2=1.245 $Y2=0.47
r88 3 22 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.88
+ $Y=0.325 $X2=4.02 $Y2=0.47
r89 2 18 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=2 $Y=0.325
+ $X2=2.14 $Y2=0.45
r90 1 14 182 $w=1.7e-07 $l=7.88797e-07 $layer=licon1_NDIFF $count=1 $X=1.045
+ $Y=0.325 $X2=1.28 $Y2=1.005
r91 1 12 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=1.045
+ $Y=0.325 $X2=1.23 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_LP__A21BOI_2%A_502_65# 1 2 9 11 12 15
c27 12 0 6.82747e-20 $X=2.815 $Y=0.35
r28 13 15 1.79269 $w=2.23e-07 $l=3.5e-08 $layer=LI1_cond $X=3.607 $Y=0.435
+ $X2=3.607 $Y2=0.47
r29 11 13 6.9898 $w=1.7e-07 $l=1.4854e-07 $layer=LI1_cond $X=3.495 $Y=0.35
+ $X2=3.607 $Y2=0.435
r30 11 12 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=3.495 $Y=0.35
+ $X2=2.815 $Y2=0.35
r31 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.65 $Y=0.435
+ $X2=2.815 $Y2=0.35
r32 7 9 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=2.65 $Y=0.435
+ $X2=2.65 $Y2=0.45
r33 2 15 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.45
+ $Y=0.325 $X2=3.59 $Y2=0.47
r34 1 9 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=2.51
+ $Y=0.325 $X2=2.65 $Y2=0.45
.ends

