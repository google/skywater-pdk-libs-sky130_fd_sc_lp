# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__nor4bb_lp
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__nor4bb_lp ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.760000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.376000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.965000 0.825000 4.675000 1.495000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.376000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.385000 1.165000 3.715000 1.495000 ;
    END
  END B
  PIN C_N
    ANTENNAGATEAREA  0.376000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.465000 1.175000 0.835000 1.845000 ;
    END
  END C_N
  PIN D_N
    ANTENNAGATEAREA  0.376000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.855000 0.825000 5.185000 1.495000 ;
    END
  END D_N
  PIN Y
    ANTENNADIFFAREA  0.520200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.565000 0.265000 2.175000 0.815000 ;
        RECT 1.565000 0.815000 3.785000 0.985000 ;
        RECT 1.565000 0.985000 2.275000 1.675000 ;
        RECT 1.565000 1.675000 2.625000 1.780000 ;
        RECT 2.105000 1.780000 2.625000 2.005000 ;
        RECT 3.455000 0.265000 3.785000 0.815000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 5.760000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 5.760000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.760000 0.085000 ;
      RECT 0.000000  3.245000 5.760000 3.415000 ;
      RECT 0.115000  0.265000 0.595000 0.825000 ;
      RECT 0.115000  0.825000 1.385000 0.995000 ;
      RECT 0.115000  0.995000 0.285000 2.025000 ;
      RECT 0.115000  2.025000 0.365000 3.065000 ;
      RECT 0.645000  2.025000 0.975000 3.245000 ;
      RECT 1.055000  0.085000 1.385000 0.645000 ;
      RECT 1.055000  0.995000 1.385000 1.790000 ;
      RECT 1.205000  2.025000 1.535000 2.185000 ;
      RECT 1.205000  2.185000 3.155000 2.355000 ;
      RECT 1.205000  2.355000 1.535000 3.065000 ;
      RECT 1.735000  2.535000 2.065000 2.895000 ;
      RECT 1.735000  2.895000 3.715000 3.065000 ;
      RECT 2.520000  1.165000 2.975000 1.495000 ;
      RECT 2.635000  0.085000 2.965000 0.635000 ;
      RECT 2.805000  1.495000 2.975000 1.675000 ;
      RECT 2.805000  1.675000 5.595000 1.845000 ;
      RECT 2.825000  2.025000 3.155000 2.185000 ;
      RECT 2.825000  2.355000 3.155000 2.715000 ;
      RECT 3.385000  2.025000 3.715000 2.895000 ;
      RECT 4.305000  0.085000 4.635000 0.645000 ;
      RECT 4.405000  2.025000 4.735000 3.245000 ;
      RECT 4.975000  1.845000 5.595000 3.065000 ;
      RECT 5.265000  0.265000 5.595000 0.645000 ;
      RECT 5.425000  0.645000 5.595000 1.675000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
  END
END sky130_fd_sc_lp__nor4bb_lp
END LIBRARY
