# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__nor3b_2
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__nor3b_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.800000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.385000 1.335000 4.715000 1.750000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.440000 1.335000 3.215000 1.665000 ;
        RECT 2.860000 1.665000 3.215000 1.750000 ;
    END
  END B
  PIN C_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.450000 0.470000 2.130000 ;
    END
  END C_N
  PIN Y
    ANTENNADIFFAREA  1.146600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.475000 1.845000 1.805000 2.735000 ;
        RECT 1.595000 0.255000 1.925000 0.985000 ;
        RECT 1.595000 0.985000 2.850000 0.995000 ;
        RECT 1.595000 0.995000 3.750000 1.165000 ;
        RECT 1.595000 1.165000 1.805000 1.845000 ;
        RECT 2.620000 0.255000 2.850000 0.985000 ;
        RECT 3.520000 0.255000 3.750000 0.995000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.800000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.800000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.800000 0.085000 ;
      RECT 0.000000  3.245000 4.800000 3.415000 ;
      RECT 0.095000  0.700000 0.355000 1.110000 ;
      RECT 0.095000  1.110000 0.925000 1.185000 ;
      RECT 0.095000  1.185000 1.425000 1.280000 ;
      RECT 0.095000  2.300000 0.925000 2.470000 ;
      RECT 0.095000  2.470000 0.355000 2.915000 ;
      RECT 0.525000  0.085000 1.425000 0.940000 ;
      RECT 0.525000  2.640000 0.855000 3.245000 ;
      RECT 0.755000  1.280000 1.425000 1.515000 ;
      RECT 0.755000  1.515000 0.925000 2.300000 ;
      RECT 1.095000  1.805000 1.305000 2.905000 ;
      RECT 1.095000  2.905000 3.095000 3.075000 ;
      RECT 1.975000  1.805000 2.165000 2.905000 ;
      RECT 2.120000  0.085000 2.450000 0.815000 ;
      RECT 2.335000  1.845000 2.665000 1.920000 ;
      RECT 2.335000  1.920000 4.190000 2.090000 ;
      RECT 2.335000  2.090000 2.665000 2.735000 ;
      RECT 2.835000  2.260000 3.095000 2.905000 ;
      RECT 3.020000  0.085000 3.350000 0.825000 ;
      RECT 3.510000  2.260000 3.840000 3.245000 ;
      RECT 3.920000  0.085000 4.210000 1.095000 ;
      RECT 4.010000  2.090000 4.190000 3.075000 ;
      RECT 4.370000  1.920000 4.700000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
  END
END sky130_fd_sc_lp__nor3b_2
