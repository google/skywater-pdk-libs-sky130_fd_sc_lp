* File: sky130_fd_sc_lp__ebufn_2.spice
* Created: Fri Aug 28 10:31:41 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__ebufn_2.pex.spice"
.subckt sky130_fd_sc_lp__ebufn_2  VNB VPB TE_B A Z VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Z	Z
* A	A
* TE_B	TE_B
* VPB	VPB
* VNB	VNB
MM1001 N_Z_M1001_d N_A_96_21#_M1001_g N_A_27_47#_M1001_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1218 AS=0.2898 PD=1.13 PS=2.37 NRD=1.428 NRS=8.568 M=1 R=5.6
+ SA=75000.3 SB=75001.6 A=0.126 P=1.98 MULT=1
MM1009 N_Z_M1001_d N_A_96_21#_M1009_g N_A_27_47#_M1009_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1218 AS=0.147 PD=1.13 PS=1.19 NRD=0 NRS=9.996 M=1 R=5.6 SA=75000.7
+ SB=75001.2 A=0.126 P=1.98 MULT=1
MM1004 N_A_27_47#_M1009_s N_A_284_21#_M1004_g N_VGND_M1004_s VNB NSHORT L=0.15
+ W=0.84 AD=0.147 AS=0.147 PD=1.19 PS=1.19 NRD=0 NRS=0 M=1 R=5.6 SA=75001.2
+ SB=75000.7 A=0.126 P=1.98 MULT=1
MM1007 N_A_27_47#_M1007_d N_A_284_21#_M1007_g N_VGND_M1004_s VNB NSHORT L=0.15
+ W=0.84 AD=0.2394 AS=0.147 PD=2.25 PS=1.19 NRD=0 NRS=9.996 M=1 R=5.6 SA=75001.7
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1008 N_VGND_M1008_d N_TE_B_M1008_g N_A_284_21#_M1008_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0882 AS=0.1197 PD=0.84 PS=1.41 NRD=19.992 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1005 N_A_96_21#_M1005_d N_A_M1005_g N_VGND_M1008_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0882 PD=1.41 PS=0.84 NRD=0 NRS=19.992 M=1 R=2.8 SA=75000.8
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1002 N_Z_M1002_d N_A_96_21#_M1002_g N_A_39_367#_M1002_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.3591 PD=1.54 PS=3.09 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75001.5 A=0.189 P=2.82 MULT=1
MM1010 N_Z_M1002_d N_A_96_21#_M1010_g N_A_39_367#_M1010_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1000 N_A_39_367#_M1010_s N_TE_B_M1000_g N_VPWR_M1000_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1003 N_A_39_367#_M1003_d N_TE_B_M1003_g N_VPWR_M1000_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3591 AS=0.1764 PD=3.09 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.5
+ SB=75000.2 A=0.189 P=2.82 MULT=1
MM1006 N_VPWR_M1006_d N_TE_B_M1006_g N_A_284_21#_M1006_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1872 AS=0.256 PD=1.525 PS=2.08 NRD=73.087 NRS=35.3812 M=1
+ R=4.26667 SA=75000.3 SB=75000.5 A=0.096 P=1.58 MULT=1
MM1011 N_A_96_21#_M1011_d N_A_M1011_g N_VPWR_M1006_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1824 AS=0.1872 PD=1.85 PS=1.525 NRD=0 NRS=21.5321 M=1 R=4.26667
+ SA=75000.7 SB=75000.2 A=0.096 P=1.58 MULT=1
DX12_noxref VNB VPB NWDIODE A=8.7655 P=13.13
*
.include "sky130_fd_sc_lp__ebufn_2.pxi.spice"
*
.ends
*
*
