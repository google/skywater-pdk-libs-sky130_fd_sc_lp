* File: sky130_fd_sc_lp__fa_1.pxi.spice
* Created: Fri Aug 28 10:34:45 2020
* 
x_PM_SKY130_FD_SC_LP__FA_1%A_80_27# N_A_80_27#_M1026_d N_A_80_27#_M1008_d
+ N_A_80_27#_M1016_g N_A_80_27#_M1017_g N_A_80_27#_M1018_g N_A_80_27#_M1025_g
+ N_A_80_27#_c_163_n N_A_80_27#_c_177_p N_A_80_27#_c_269_p N_A_80_27#_c_164_n
+ N_A_80_27#_c_165_n N_A_80_27#_c_166_n N_A_80_27#_c_167_n N_A_80_27#_c_168_n
+ N_A_80_27#_c_178_p N_A_80_27#_c_175_n N_A_80_27#_c_176_n N_A_80_27#_c_169_n
+ PM_SKY130_FD_SC_LP__FA_1%A_80_27#
x_PM_SKY130_FD_SC_LP__FA_1%A N_A_M1004_g N_A_M1006_g N_A_M1005_g N_A_M1020_g
+ N_A_M1007_g N_A_c_307_n N_A_c_308_n N_A_M1010_g N_A_M1009_g N_A_M1019_g
+ N_A_c_311_n N_A_c_312_n N_A_c_323_n N_A_c_324_n N_A_c_325_n N_A_c_326_n
+ N_A_c_327_n N_A_c_328_n A N_A_c_313_n N_A_c_314_n N_A_c_315_n N_A_c_316_n
+ N_A_c_331_n N_A_c_332_n PM_SKY130_FD_SC_LP__FA_1%A
x_PM_SKY130_FD_SC_LP__FA_1%B N_B_M1008_g N_B_M1026_g N_B_c_515_n N_B_c_516_n
+ N_B_M1021_g N_B_M1012_g N_B_c_519_n N_B_c_520_n N_B_c_521_n N_B_M1022_g
+ N_B_c_523_n N_B_c_537_n N_B_M1002_g N_B_M1014_g N_B_M1000_g N_B_c_539_n
+ N_B_c_524_n N_B_c_525_n N_B_c_540_n N_B_c_526_n N_B_c_527_n N_B_c_541_n
+ N_B_c_528_n N_B_c_529_n B B N_B_c_532_n N_B_c_533_n PM_SKY130_FD_SC_LP__FA_1%B
x_PM_SKY130_FD_SC_LP__FA_1%CIN N_CIN_M1015_g N_CIN_M1001_g N_CIN_c_688_n
+ N_CIN_c_689_n N_CIN_c_690_n N_CIN_c_691_n N_CIN_M1024_g N_CIN_M1003_g
+ N_CIN_c_693_n N_CIN_M1027_g N_CIN_M1011_g N_CIN_c_695_n N_CIN_c_696_n
+ N_CIN_c_685_n N_CIN_c_697_n N_CIN_c_698_n N_CIN_c_699_n CIN CIN
+ PM_SKY130_FD_SC_LP__FA_1%CIN
x_PM_SKY130_FD_SC_LP__FA_1%A_1118_411# N_A_1118_411#_M1025_d
+ N_A_1118_411#_M1018_d N_A_1118_411#_M1023_g N_A_1118_411#_M1013_g
+ N_A_1118_411#_c_827_n N_A_1118_411#_c_828_n N_A_1118_411#_c_833_n
+ N_A_1118_411#_c_814_n N_A_1118_411#_c_821_n N_A_1118_411#_c_839_n
+ N_A_1118_411#_c_815_n N_A_1118_411#_c_816_n N_A_1118_411#_c_817_n
+ N_A_1118_411#_c_818_n PM_SKY130_FD_SC_LP__FA_1%A_1118_411#
x_PM_SKY130_FD_SC_LP__FA_1%COUT N_COUT_M1016_s N_COUT_M1017_s COUT COUT COUT
+ COUT COUT COUT N_COUT_c_890_n COUT PM_SKY130_FD_SC_LP__FA_1%COUT
x_PM_SKY130_FD_SC_LP__FA_1%VPWR N_VPWR_M1017_d N_VPWR_M1005_d N_VPWR_M1002_s
+ N_VPWR_M1003_d N_VPWR_M1019_d N_VPWR_c_907_n N_VPWR_c_908_n N_VPWR_c_909_n
+ N_VPWR_c_910_n N_VPWR_c_911_n N_VPWR_c_912_n N_VPWR_c_913_n N_VPWR_c_931_n
+ N_VPWR_c_914_n N_VPWR_c_915_n VPWR N_VPWR_c_916_n N_VPWR_c_917_n
+ N_VPWR_c_918_n N_VPWR_c_919_n N_VPWR_c_906_n N_VPWR_c_921_n N_VPWR_c_922_n
+ N_VPWR_c_923_n PM_SKY130_FD_SC_LP__FA_1%VPWR
x_PM_SKY130_FD_SC_LP__FA_1%A_417_457# N_A_417_457#_M1015_d N_A_417_457#_M1012_d
+ N_A_417_457#_c_1010_n N_A_417_457#_c_1011_n
+ PM_SKY130_FD_SC_LP__FA_1%A_417_457#
x_PM_SKY130_FD_SC_LP__FA_1%A_854_411# N_A_854_411#_M1002_d N_A_854_411#_M1010_d
+ N_A_854_411#_c_1034_n N_A_854_411#_c_1035_n N_A_854_411#_c_1036_n
+ N_A_854_411#_c_1037_n PM_SKY130_FD_SC_LP__FA_1%A_854_411#
x_PM_SKY130_FD_SC_LP__FA_1%SUM N_SUM_M1023_d N_SUM_M1013_d N_SUM_c_1071_n
+ N_SUM_c_1072_n N_SUM_c_1068_n SUM SUM N_SUM_c_1070_n
+ PM_SKY130_FD_SC_LP__FA_1%SUM
x_PM_SKY130_FD_SC_LP__FA_1%VGND N_VGND_M1016_d N_VGND_M1020_d N_VGND_M1022_s
+ N_VGND_M1024_d N_VGND_M1009_d N_VGND_c_1089_n N_VGND_c_1090_n N_VGND_c_1091_n
+ N_VGND_c_1092_n N_VGND_c_1093_n N_VGND_c_1094_n N_VGND_c_1095_n
+ N_VGND_c_1096_n N_VGND_c_1097_n N_VGND_c_1098_n VGND N_VGND_c_1099_n
+ N_VGND_c_1100_n N_VGND_c_1101_n N_VGND_c_1102_n N_VGND_c_1103_n
+ N_VGND_c_1104_n N_VGND_c_1105_n PM_SKY130_FD_SC_LP__FA_1%VGND
x_PM_SKY130_FD_SC_LP__FA_1%A_431_137# N_A_431_137#_M1001_d N_A_431_137#_M1021_d
+ N_A_431_137#_c_1185_n N_A_431_137#_c_1186_n N_A_431_137#_c_1187_n
+ N_A_431_137#_c_1188_n PM_SKY130_FD_SC_LP__FA_1%A_431_137#
x_PM_SKY130_FD_SC_LP__FA_1%A_818_83# N_A_818_83#_M1022_d N_A_818_83#_M1007_d
+ N_A_818_83#_c_1229_n N_A_818_83#_c_1213_n N_A_818_83#_c_1214_n
+ N_A_818_83#_c_1215_n PM_SKY130_FD_SC_LP__FA_1%A_818_83#
cc_1 VNB N_A_80_27#_M1017_g 0.00610546f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=2.465
cc_2 VNB N_A_80_27#_M1025_g 0.0319803f $X=-0.19 $Y=-0.245 $X2=5.555 $Y2=0.835
cc_3 VNB N_A_80_27#_c_163_n 7.17345e-19 $X=-0.19 $Y=-0.245 $X2=0.675 $Y2=2.3
cc_4 VNB N_A_80_27#_c_164_n 0.00376293f $X=-0.19 $Y=-0.245 $X2=1.865 $Y2=0.895
cc_5 VNB N_A_80_27#_c_165_n 0.0220384f $X=-0.19 $Y=-0.245 $X2=5.535 $Y2=1.61
cc_6 VNB N_A_80_27#_c_166_n 0.0169481f $X=-0.19 $Y=-0.245 $X2=5.535 $Y2=1.61
cc_7 VNB N_A_80_27#_c_167_n 0.00228617f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.38
cc_8 VNB N_A_80_27#_c_168_n 0.0418465f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.38
cc_9 VNB N_A_80_27#_c_169_n 0.0224739f $X=-0.19 $Y=-0.245 $X2=0.597 $Y2=1.215
cc_10 VNB N_A_M1004_g 0.00169147f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_M1006_g 0.0235144f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.215
cc_12 VNB N_A_M1020_g 0.0358994f $X=-0.19 $Y=-0.245 $X2=5.515 $Y2=2.265
cc_13 VNB N_A_M1007_g 0.0211279f $X=-0.19 $Y=-0.245 $X2=5.555 $Y2=0.835
cc_14 VNB N_A_c_307_n 0.14503f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_c_308_n 0.011606f $X=-0.19 $Y=-0.245 $X2=0.675 $Y2=1.545
cc_16 VNB N_A_M1010_g 0.0193978f $X=-0.19 $Y=-0.245 $X2=0.795 $Y2=2.385
cc_17 VNB N_A_M1009_g 0.0376059f $X=-0.19 $Y=-0.245 $X2=1.81 $Y2=1.695
cc_18 VNB N_A_c_311_n 0.020407f $X=-0.19 $Y=-0.245 $X2=0.665 $Y2=1.38
cc_19 VNB N_A_c_312_n 0.0201515f $X=-0.19 $Y=-0.245 $X2=0.665 $Y2=1.545
cc_20 VNB N_A_c_313_n 0.0153466f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_c_314_n 0.00435611f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_c_315_n 0.0317688f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_c_316_n 0.00520653f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_B_M1026_g 0.0539365f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.215
cc_25 VNB N_B_c_515_n 0.0793804f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.685
cc_26 VNB N_B_c_516_n 0.0123287f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.685
cc_27 VNB N_B_M1021_g 0.0281142f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_B_M1012_g 0.0164389f $X=-0.19 $Y=-0.245 $X2=5.515 $Y2=2.265
cc_29 VNB N_B_c_519_n 0.0417825f $X=-0.19 $Y=-0.245 $X2=5.555 $Y2=1.445
cc_30 VNB N_B_c_520_n 0.0197799f $X=-0.19 $Y=-0.245 $X2=5.555 $Y2=0.835
cc_31 VNB N_B_c_521_n 0.0398538f $X=-0.19 $Y=-0.245 $X2=0.675 $Y2=2.3
cc_32 VNB N_B_M1022_g 0.0219998f $X=-0.19 $Y=-0.245 $X2=1.842 $Y2=1.525
cc_33 VNB N_B_c_523_n 0.0154619f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_B_c_524_n 0.00732516f $X=-0.19 $Y=-0.245 $X2=1.775 $Y2=2.385
cc_35 VNB N_B_c_525_n 0.00857305f $X=-0.19 $Y=-0.245 $X2=1.775 $Y2=2.3
cc_36 VNB N_B_c_526_n 0.0165086f $X=-0.19 $Y=-0.245 $X2=0.597 $Y2=1.215
cc_37 VNB N_B_c_527_n 0.0194455f $X=-0.19 $Y=-0.245 $X2=0.597 $Y2=1.545
cc_38 VNB N_B_c_528_n 6.27546e-19 $X=-0.19 $Y=-0.245 $X2=5.535 $Y2=1.445
cc_39 VNB N_B_c_529_n 0.0152556f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB B 0.00750919f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB B 0.00533638f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_B_c_532_n 0.0146049f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_B_c_533_n 0.0552852f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_CIN_M1001_g 0.0369358f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.215
cc_45 VNB N_CIN_M1024_g 0.0417777f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_CIN_M1003_g 7.01305e-19 $X=-0.19 $Y=-0.245 $X2=0.675 $Y2=1.545
cc_47 VNB N_CIN_M1027_g 0.0373263f $X=-0.19 $Y=-0.245 $X2=1.842 $Y2=0.895
cc_48 VNB N_CIN_c_685_n 0.0206586f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.38
cc_49 VNB N_A_1118_411#_M1013_g 0.00739951f $X=-0.19 $Y=-0.245 $X2=0.485
+ $Y2=2.465
cc_50 VNB N_A_1118_411#_c_814_n 7.90942e-19 $X=-0.19 $Y=-0.245 $X2=0.795
+ $Y2=2.385
cc_51 VNB N_A_1118_411#_c_815_n 0.00393636f $X=-0.19 $Y=-0.245 $X2=5.535
+ $Y2=1.61
cc_52 VNB N_A_1118_411#_c_816_n 0.034501f $X=-0.19 $Y=-0.245 $X2=5.535 $Y2=1.61
cc_53 VNB N_A_1118_411#_c_817_n 0.00115022f $X=-0.19 $Y=-0.245 $X2=5.535
+ $Y2=1.61
cc_54 VNB N_A_1118_411#_c_818_n 0.0202345f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.38
cc_55 VNB N_COUT_c_890_n 0.0639583f $X=-0.19 $Y=-0.245 $X2=0.675 $Y2=1.545
cc_56 VNB N_VPWR_c_906_n 0.342803f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_SUM_c_1068_n 0.0318113f $X=-0.19 $Y=-0.245 $X2=5.515 $Y2=2.265
cc_58 VNB SUM 0.00992243f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_SUM_c_1070_n 0.0264241f $X=-0.19 $Y=-0.245 $X2=0.675 $Y2=1.545
cc_60 VNB N_VGND_c_1089_n 0.0137255f $X=-0.19 $Y=-0.245 $X2=5.555 $Y2=1.445
cc_61 VNB N_VGND_c_1090_n 0.0109783f $X=-0.19 $Y=-0.245 $X2=1.63 $Y2=2.385
cc_62 VNB N_VGND_c_1091_n 0.0148106f $X=-0.19 $Y=-0.245 $X2=1.865 $Y2=0.895
cc_63 VNB N_VGND_c_1092_n 0.0168587f $X=-0.19 $Y=-0.245 $X2=1.81 $Y2=1.695
cc_64 VNB N_VGND_c_1093_n 0.00225152f $X=-0.19 $Y=-0.245 $X2=5.535 $Y2=1.61
cc_65 VNB N_VGND_c_1094_n 0.00733085f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.38
cc_66 VNB N_VGND_c_1095_n 0.022189f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_1096_n 0.00577043f $X=-0.19 $Y=-0.245 $X2=0.665 $Y2=1.545
cc_68 VNB N_VGND_c_1097_n 0.0629727f $X=-0.19 $Y=-0.245 $X2=1.775 $Y2=2.3
cc_69 VNB N_VGND_c_1098_n 0.00513431f $X=-0.19 $Y=-0.245 $X2=1.775 $Y2=2.49
cc_70 VNB N_VGND_c_1099_n 0.0157034f $X=-0.19 $Y=-0.245 $X2=1.842 $Y2=1.61
cc_71 VNB N_VGND_c_1100_n 0.040649f $X=-0.19 $Y=-0.245 $X2=5.535 $Y2=1.445
cc_72 VNB N_VGND_c_1101_n 0.0189802f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_VGND_c_1102_n 0.414749f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_VGND_c_1103_n 0.0118535f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_VGND_c_1104_n 0.00512691f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_VGND_c_1105_n 0.00513431f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_A_431_137#_c_1185_n 0.00140877f $X=-0.19 $Y=-0.245 $X2=0.475
+ $Y2=0.685
cc_78 VNB N_A_431_137#_c_1186_n 0.00892937f $X=-0.19 $Y=-0.245 $X2=0.485
+ $Y2=2.465
cc_79 VNB N_A_431_137#_c_1187_n 0.00262604f $X=-0.19 $Y=-0.245 $X2=0.485
+ $Y2=2.465
cc_80 VNB N_A_431_137#_c_1188_n 0.0011457f $X=-0.19 $Y=-0.245 $X2=5.515
+ $Y2=2.265
cc_81 VNB N_A_818_83#_c_1213_n 0.00316739f $X=-0.19 $Y=-0.245 $X2=0.485
+ $Y2=2.465
cc_82 VNB N_A_818_83#_c_1214_n 0.00419356f $X=-0.19 $Y=-0.245 $X2=0.485
+ $Y2=2.465
cc_83 VNB N_A_818_83#_c_1215_n 0.00831244f $X=-0.19 $Y=-0.245 $X2=5.515
+ $Y2=1.775
cc_84 VPB N_A_80_27#_M1017_g 0.0251508f $X=-0.19 $Y=1.655 $X2=0.485 $Y2=2.465
cc_85 VPB N_A_80_27#_M1018_g 0.0243538f $X=-0.19 $Y=1.655 $X2=5.515 $Y2=2.265
cc_86 VPB N_A_80_27#_c_163_n 0.00140431f $X=-0.19 $Y=1.655 $X2=0.675 $Y2=2.3
cc_87 VPB N_A_80_27#_c_165_n 0.0224854f $X=-0.19 $Y=1.655 $X2=5.535 $Y2=1.61
cc_88 VPB N_A_80_27#_c_166_n 0.0125963f $X=-0.19 $Y=1.655 $X2=5.535 $Y2=1.61
cc_89 VPB N_A_80_27#_c_175_n 0.00584756f $X=-0.19 $Y=1.655 $X2=1.775 $Y2=2.3
cc_90 VPB N_A_80_27#_c_176_n 4.56748e-19 $X=-0.19 $Y=1.655 $X2=1.842 $Y2=1.61
cc_91 VPB N_A_M1004_g 0.0497084f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_92 VPB N_A_M1005_g 0.0192466f $X=-0.19 $Y=1.655 $X2=0.485 $Y2=2.465
cc_93 VPB N_A_M1020_g 0.00751904f $X=-0.19 $Y=1.655 $X2=5.515 $Y2=2.265
cc_94 VPB N_A_M1010_g 0.0273587f $X=-0.19 $Y=1.655 $X2=0.795 $Y2=2.385
cc_95 VPB N_A_M1019_g 0.0255252f $X=-0.19 $Y=1.655 $X2=5.535 $Y2=1.61
cc_96 VPB N_A_c_312_n 0.00238704f $X=-0.19 $Y=1.655 $X2=0.665 $Y2=1.545
cc_97 VPB N_A_c_323_n 0.0171562f $X=-0.19 $Y=1.655 $X2=1.775 $Y2=2.385
cc_98 VPB N_A_c_324_n 0.0135668f $X=-0.19 $Y=1.655 $X2=1.775 $Y2=2.3
cc_99 VPB N_A_c_325_n 0.00217111f $X=-0.19 $Y=1.655 $X2=1.775 $Y2=2.49
cc_100 VPB N_A_c_326_n 0.0275213f $X=-0.19 $Y=1.655 $X2=1.795 $Y2=2.49
cc_101 VPB N_A_c_327_n 0.00301794f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_102 VPB N_A_c_328_n 9.30636e-19 $X=-0.19 $Y=1.655 $X2=5.535 $Y2=1.61
cc_103 VPB N_A_c_314_n 0.00539133f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_104 VPB N_A_c_316_n 0.00420752f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_105 VPB N_A_c_331_n 0.0294334f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_106 VPB N_A_c_332_n 0.00614439f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_107 VPB N_B_M1026_g 0.0208789f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=1.215
cc_108 VPB N_B_M1012_g 0.0480523f $X=-0.19 $Y=1.655 $X2=5.515 $Y2=2.265
cc_109 VPB N_B_c_523_n 0.0142918f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_110 VPB N_B_c_537_n 0.0139712f $X=-0.19 $Y=1.655 $X2=1.81 $Y2=1.695
cc_111 VPB N_B_M1000_g 0.0251127f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=1.38
cc_112 VPB N_B_c_539_n 0.0284831f $X=-0.19 $Y=1.655 $X2=0.665 $Y2=1.545
cc_113 VPB N_B_c_540_n 0.0163004f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_114 VPB N_B_c_541_n 0.0154009f $X=-0.19 $Y=1.655 $X2=5.535 $Y2=1.61
cc_115 VPB B 0.00368673f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_116 VPB N_CIN_M1015_g 0.0300429f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_117 VPB N_CIN_M1001_g 0.0195836f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=1.215
cc_118 VPB N_CIN_c_688_n 0.104915f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.685
cc_119 VPB N_CIN_c_689_n 0.0134436f $X=-0.19 $Y=1.655 $X2=0.485 $Y2=1.545
cc_120 VPB N_CIN_c_690_n 0.0385772f $X=-0.19 $Y=1.655 $X2=0.485 $Y2=2.465
cc_121 VPB N_CIN_c_691_n 0.0570484f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_122 VPB N_CIN_M1003_g 0.0374701f $X=-0.19 $Y=1.655 $X2=0.675 $Y2=1.545
cc_123 VPB N_CIN_c_693_n 0.0880669f $X=-0.19 $Y=1.655 $X2=0.675 $Y2=2.3
cc_124 VPB N_CIN_M1027_g 0.0492213f $X=-0.19 $Y=1.655 $X2=1.842 $Y2=0.895
cc_125 VPB N_CIN_c_695_n 0.0122517f $X=-0.19 $Y=1.655 $X2=1.985 $Y2=1.61
cc_126 VPB N_CIN_c_696_n 0.0245214f $X=-0.19 $Y=1.655 $X2=5.535 $Y2=1.61
cc_127 VPB N_CIN_c_697_n 0.00661134f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_128 VPB N_CIN_c_698_n 0.0377669f $X=-0.19 $Y=1.655 $X2=1.775 $Y2=2.3
cc_129 VPB N_CIN_c_699_n 0.00476332f $X=-0.19 $Y=1.655 $X2=1.795 $Y2=2.49
cc_130 VPB CIN 0.0138078f $X=-0.19 $Y=1.655 $X2=0.597 $Y2=1.38
cc_131 VPB N_A_1118_411#_M1013_g 0.0250043f $X=-0.19 $Y=1.655 $X2=0.485
+ $Y2=2.465
cc_132 VPB N_A_1118_411#_c_814_n 0.00340679f $X=-0.19 $Y=1.655 $X2=0.795
+ $Y2=2.385
cc_133 VPB COUT 0.00628324f $X=-0.19 $Y=1.655 $X2=0.485 $Y2=2.465
cc_134 VPB N_COUT_c_890_n 0.00838036f $X=-0.19 $Y=1.655 $X2=0.675 $Y2=1.545
cc_135 VPB COUT 0.0437256f $X=-0.19 $Y=1.655 $X2=5.535 $Y2=1.61
cc_136 VPB N_VPWR_c_907_n 0.0142782f $X=-0.19 $Y=1.655 $X2=5.555 $Y2=1.445
cc_137 VPB N_VPWR_c_908_n 0.00982308f $X=-0.19 $Y=1.655 $X2=0.675 $Y2=1.545
cc_138 VPB N_VPWR_c_909_n 0.0198634f $X=-0.19 $Y=1.655 $X2=1.842 $Y2=1.525
cc_139 VPB N_VPWR_c_910_n 0.0236385f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_140 VPB N_VPWR_c_911_n 0.0206443f $X=-0.19 $Y=1.655 $X2=1.985 $Y2=1.61
cc_141 VPB N_VPWR_c_912_n 0.027879f $X=-0.19 $Y=1.655 $X2=5.535 $Y2=1.61
cc_142 VPB N_VPWR_c_913_n 0.00449427f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_143 VPB N_VPWR_c_914_n 0.0230073f $X=-0.19 $Y=1.655 $X2=1.775 $Y2=2.385
cc_144 VPB N_VPWR_c_915_n 0.00362871f $X=-0.19 $Y=1.655 $X2=1.775 $Y2=2.3
cc_145 VPB N_VPWR_c_916_n 0.0160483f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_146 VPB N_VPWR_c_917_n 0.0502858f $X=-0.19 $Y=1.655 $X2=5.535 $Y2=1.61
cc_147 VPB N_VPWR_c_918_n 0.0715359f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_148 VPB N_VPWR_c_919_n 0.0158241f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_149 VPB N_VPWR_c_906_n 0.108404f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_150 VPB N_VPWR_c_921_n 0.00522677f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_151 VPB N_VPWR_c_922_n 0.00473485f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_152 VPB N_VPWR_c_923_n 0.00522677f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_153 VPB N_A_854_411#_c_1034_n 3.97125e-19 $X=-0.19 $Y=1.655 $X2=0.475
+ $Y2=0.685
cc_154 VPB N_A_854_411#_c_1035_n 0.00946035f $X=-0.19 $Y=1.655 $X2=0.485
+ $Y2=2.465
cc_155 VPB N_A_854_411#_c_1036_n 0.00397907f $X=-0.19 $Y=1.655 $X2=0.485
+ $Y2=2.465
cc_156 VPB N_A_854_411#_c_1037_n 4.62516e-19 $X=-0.19 $Y=1.655 $X2=5.515
+ $Y2=2.265
cc_157 VPB N_SUM_c_1071_n 0.00743295f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=1.215
cc_158 VPB N_SUM_c_1072_n 0.043257f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.685
cc_159 VPB N_SUM_c_1068_n 0.00805538f $X=-0.19 $Y=1.655 $X2=5.515 $Y2=2.265
cc_160 N_A_80_27#_c_177_p N_A_M1004_g 0.0127939f $X=1.63 $Y=2.385 $X2=0 $Y2=0
cc_161 N_A_80_27#_c_178_p N_A_M1004_g 9.5866e-19 $X=1.775 $Y=2.385 $X2=0 $Y2=0
cc_162 N_A_80_27#_c_175_n N_A_M1004_g 7.56334e-19 $X=1.775 $Y=2.3 $X2=0 $Y2=0
cc_163 N_A_80_27#_c_164_n N_A_M1006_g 0.00213694f $X=1.865 $Y=0.895 $X2=0 $Y2=0
cc_164 N_A_80_27#_c_167_n N_A_M1006_g 4.61019e-19 $X=0.63 $Y=1.38 $X2=0 $Y2=0
cc_165 N_A_80_27#_c_168_n N_A_M1006_g 0.00274499f $X=0.63 $Y=1.38 $X2=0 $Y2=0
cc_166 N_A_80_27#_c_169_n N_A_M1006_g 0.00459178f $X=0.597 $Y=1.215 $X2=0 $Y2=0
cc_167 N_A_80_27#_c_165_n N_A_M1020_g 0.0108175f $X=5.535 $Y=1.61 $X2=0 $Y2=0
cc_168 N_A_80_27#_M1025_g N_A_M1007_g 0.00441558f $X=5.555 $Y=0.835 $X2=0 $Y2=0
cc_169 N_A_80_27#_M1025_g N_A_c_307_n 0.0089235f $X=5.555 $Y=0.835 $X2=0 $Y2=0
cc_170 N_A_80_27#_M1018_g N_A_M1010_g 0.0202074f $X=5.515 $Y=2.265 $X2=0 $Y2=0
cc_171 N_A_80_27#_c_165_n N_A_M1010_g 0.0098748f $X=5.535 $Y=1.61 $X2=0 $Y2=0
cc_172 N_A_80_27#_c_166_n N_A_M1010_g 0.022218f $X=5.535 $Y=1.61 $X2=0 $Y2=0
cc_173 N_A_80_27#_M1025_g N_A_c_311_n 0.0133836f $X=5.555 $Y=0.835 $X2=0 $Y2=0
cc_174 N_A_80_27#_c_165_n N_A_c_311_n 0.00106296f $X=5.535 $Y=1.61 $X2=0 $Y2=0
cc_175 N_A_80_27#_c_177_p N_A_c_324_n 0.0116765f $X=1.63 $Y=2.385 $X2=0 $Y2=0
cc_176 N_A_80_27#_c_165_n N_A_c_324_n 0.0117062f $X=5.535 $Y=1.61 $X2=0 $Y2=0
cc_177 N_A_80_27#_c_178_p N_A_c_324_n 0.00290703f $X=1.775 $Y=2.385 $X2=0 $Y2=0
cc_178 N_A_80_27#_c_175_n N_A_c_324_n 0.031114f $X=1.775 $Y=2.3 $X2=0 $Y2=0
cc_179 N_A_80_27#_c_176_n N_A_c_324_n 0.00310104f $X=1.842 $Y=1.61 $X2=0 $Y2=0
cc_180 N_A_80_27#_c_163_n N_A_c_325_n 0.00222863f $X=0.675 $Y=2.3 $X2=0 $Y2=0
cc_181 N_A_80_27#_c_177_p N_A_c_325_n 0.00773477f $X=1.63 $Y=2.385 $X2=0 $Y2=0
cc_182 N_A_80_27#_c_175_n N_A_c_325_n 0.00250724f $X=1.775 $Y=2.3 $X2=0 $Y2=0
cc_183 N_A_80_27#_M1018_g N_A_c_326_n 0.00848034f $X=5.515 $Y=2.265 $X2=0 $Y2=0
cc_184 N_A_80_27#_c_165_n N_A_c_326_n 0.0514942f $X=5.535 $Y=1.61 $X2=0 $Y2=0
cc_185 N_A_80_27#_c_166_n N_A_c_326_n 0.00289017f $X=5.535 $Y=1.61 $X2=0 $Y2=0
cc_186 N_A_80_27#_c_165_n N_A_c_327_n 0.00186707f $X=5.535 $Y=1.61 $X2=0 $Y2=0
cc_187 N_A_80_27#_c_175_n N_A_c_327_n 0.00102754f $X=1.775 $Y=2.3 $X2=0 $Y2=0
cc_188 N_A_80_27#_M1017_g N_A_c_315_n 0.0253357f $X=0.485 $Y=2.465 $X2=0 $Y2=0
cc_189 N_A_80_27#_c_163_n N_A_c_315_n 0.00815841f $X=0.675 $Y=2.3 $X2=0 $Y2=0
cc_190 N_A_80_27#_c_177_p N_A_c_315_n 4.12844e-19 $X=1.63 $Y=2.385 $X2=0 $Y2=0
cc_191 N_A_80_27#_c_164_n N_A_c_315_n 2.4134e-19 $X=1.865 $Y=0.895 $X2=0 $Y2=0
cc_192 N_A_80_27#_c_167_n N_A_c_315_n 8.71685e-19 $X=0.63 $Y=1.38 $X2=0 $Y2=0
cc_193 N_A_80_27#_c_168_n N_A_c_315_n 0.0154451f $X=0.63 $Y=1.38 $X2=0 $Y2=0
cc_194 N_A_80_27#_M1017_g N_A_c_316_n 5.42164e-19 $X=0.485 $Y=2.465 $X2=0 $Y2=0
cc_195 N_A_80_27#_c_177_p N_A_c_316_n 0.0206617f $X=1.63 $Y=2.385 $X2=0 $Y2=0
cc_196 N_A_80_27#_c_164_n N_A_c_316_n 0.0104227f $X=1.865 $Y=0.895 $X2=0 $Y2=0
cc_197 N_A_80_27#_c_167_n N_A_c_316_n 0.052215f $X=0.63 $Y=1.38 $X2=0 $Y2=0
cc_198 N_A_80_27#_c_168_n N_A_c_316_n 9.00408e-19 $X=0.63 $Y=1.38 $X2=0 $Y2=0
cc_199 N_A_80_27#_c_175_n N_A_c_316_n 0.0164188f $X=1.775 $Y=2.3 $X2=0 $Y2=0
cc_200 N_A_80_27#_c_176_n N_A_c_316_n 0.00822927f $X=1.842 $Y=1.61 $X2=0 $Y2=0
cc_201 N_A_80_27#_c_165_n N_A_c_331_n 0.00468135f $X=5.535 $Y=1.61 $X2=0 $Y2=0
cc_202 N_A_80_27#_c_165_n N_A_c_332_n 0.0283721f $X=5.535 $Y=1.61 $X2=0 $Y2=0
cc_203 N_A_80_27#_c_175_n N_A_c_332_n 0.007383f $X=1.775 $Y=2.3 $X2=0 $Y2=0
cc_204 N_A_80_27#_c_164_n N_B_M1026_g 0.0176876f $X=1.865 $Y=0.895 $X2=0 $Y2=0
cc_205 N_A_80_27#_c_175_n N_B_M1026_g 0.00795789f $X=1.775 $Y=2.3 $X2=0 $Y2=0
cc_206 N_A_80_27#_c_176_n N_B_M1026_g 0.00443765f $X=1.842 $Y=1.61 $X2=0 $Y2=0
cc_207 N_A_80_27#_c_164_n N_B_c_515_n 0.00304194f $X=1.865 $Y=0.895 $X2=0 $Y2=0
cc_208 N_A_80_27#_c_165_n N_B_M1012_g 0.0146583f $X=5.535 $Y=1.61 $X2=0 $Y2=0
cc_209 N_A_80_27#_c_165_n N_B_c_520_n 0.0155f $X=5.535 $Y=1.61 $X2=0 $Y2=0
cc_210 N_A_80_27#_c_165_n N_B_c_523_n 0.0134704f $X=5.535 $Y=1.61 $X2=0 $Y2=0
cc_211 N_A_80_27#_c_177_p N_B_c_539_n 0.00950387f $X=1.63 $Y=2.385 $X2=0 $Y2=0
cc_212 N_A_80_27#_c_178_p N_B_c_539_n 0.00525753f $X=1.775 $Y=2.385 $X2=0 $Y2=0
cc_213 N_A_80_27#_c_175_n N_B_c_539_n 0.00578524f $X=1.775 $Y=2.3 $X2=0 $Y2=0
cc_214 N_A_80_27#_c_165_n N_B_c_525_n 0.0025745f $X=5.535 $Y=1.61 $X2=0 $Y2=0
cc_215 N_A_80_27#_c_165_n N_B_c_540_n 0.00452662f $X=5.535 $Y=1.61 $X2=0 $Y2=0
cc_216 N_A_80_27#_c_165_n N_B_c_528_n 0.0255627f $X=5.535 $Y=1.61 $X2=0 $Y2=0
cc_217 N_A_80_27#_M1025_g N_B_c_529_n 0.0034772f $X=5.555 $Y=0.835 $X2=0 $Y2=0
cc_218 N_A_80_27#_c_165_n N_B_c_529_n 0.120746f $X=5.535 $Y=1.61 $X2=0 $Y2=0
cc_219 N_A_80_27#_c_166_n N_B_c_529_n 0.00289308f $X=5.535 $Y=1.61 $X2=0 $Y2=0
cc_220 N_A_80_27#_M1025_g B 0.0118362f $X=5.555 $Y=0.835 $X2=0 $Y2=0
cc_221 N_A_80_27#_c_165_n B 0.0137856f $X=5.535 $Y=1.61 $X2=0 $Y2=0
cc_222 N_A_80_27#_c_166_n B 0.0017253f $X=5.535 $Y=1.61 $X2=0 $Y2=0
cc_223 N_A_80_27#_M1018_g B 2.89637e-19 $X=5.515 $Y=2.265 $X2=0 $Y2=0
cc_224 N_A_80_27#_M1025_g B 5.50344e-19 $X=5.555 $Y=0.835 $X2=0 $Y2=0
cc_225 N_A_80_27#_c_165_n B 0.0118072f $X=5.535 $Y=1.61 $X2=0 $Y2=0
cc_226 N_A_80_27#_c_166_n B 0.00133981f $X=5.535 $Y=1.61 $X2=0 $Y2=0
cc_227 N_A_80_27#_c_164_n N_CIN_M1001_g 0.00669551f $X=1.865 $Y=0.895 $X2=0
+ $Y2=0
cc_228 N_A_80_27#_c_165_n N_CIN_M1001_g 0.0158733f $X=5.535 $Y=1.61 $X2=0 $Y2=0
cc_229 N_A_80_27#_c_175_n N_CIN_M1001_g 0.00594283f $X=1.775 $Y=2.3 $X2=0 $Y2=0
cc_230 N_A_80_27#_c_165_n N_CIN_M1003_g 0.0036468f $X=5.535 $Y=1.61 $X2=0 $Y2=0
cc_231 N_A_80_27#_M1018_g N_CIN_c_693_n 0.0108224f $X=5.515 $Y=2.265 $X2=0 $Y2=0
cc_232 N_A_80_27#_M1018_g N_CIN_M1027_g 0.0187002f $X=5.515 $Y=2.265 $X2=0 $Y2=0
cc_233 N_A_80_27#_M1025_g N_CIN_M1027_g 0.0260719f $X=5.555 $Y=0.835 $X2=0 $Y2=0
cc_234 N_A_80_27#_c_165_n N_CIN_M1027_g 5.06854e-19 $X=5.535 $Y=1.61 $X2=0 $Y2=0
cc_235 N_A_80_27#_c_166_n N_CIN_M1027_g 0.020278f $X=5.535 $Y=1.61 $X2=0 $Y2=0
cc_236 N_A_80_27#_c_165_n N_CIN_c_695_n 4.99272e-19 $X=5.535 $Y=1.61 $X2=0 $Y2=0
cc_237 N_A_80_27#_c_175_n N_CIN_c_695_n 0.00477622f $X=1.775 $Y=2.3 $X2=0 $Y2=0
cc_238 N_A_80_27#_c_176_n N_CIN_c_695_n 0.00156296f $X=1.842 $Y=1.61 $X2=0 $Y2=0
cc_239 N_A_80_27#_c_165_n N_CIN_c_685_n 0.0121227f $X=5.535 $Y=1.61 $X2=0 $Y2=0
cc_240 N_A_80_27#_c_165_n N_CIN_c_698_n 0.00293788f $X=5.535 $Y=1.61 $X2=0 $Y2=0
cc_241 N_A_80_27#_c_165_n N_CIN_c_699_n 0.023907f $X=5.535 $Y=1.61 $X2=0 $Y2=0
cc_242 N_A_80_27#_c_165_n N_A_1118_411#_c_821_n 0.00189815f $X=5.535 $Y=1.61
+ $X2=0 $Y2=0
cc_243 N_A_80_27#_c_166_n N_A_1118_411#_c_821_n 0.00189784f $X=5.535 $Y=1.61
+ $X2=0 $Y2=0
cc_244 N_A_80_27#_M1017_g COUT 0.00339457f $X=0.485 $Y=2.465 $X2=0 $Y2=0
cc_245 N_A_80_27#_c_163_n COUT 0.0172653f $X=0.675 $Y=2.3 $X2=0 $Y2=0
cc_246 N_A_80_27#_M1017_g N_COUT_c_890_n 0.00615752f $X=0.485 $Y=2.465 $X2=0
+ $Y2=0
cc_247 N_A_80_27#_c_163_n N_COUT_c_890_n 0.0188867f $X=0.675 $Y=2.3 $X2=0 $Y2=0
cc_248 N_A_80_27#_c_167_n N_COUT_c_890_n 0.0253306f $X=0.63 $Y=1.38 $X2=0 $Y2=0
cc_249 N_A_80_27#_c_169_n N_COUT_c_890_n 0.0168865f $X=0.597 $Y=1.215 $X2=0
+ $Y2=0
cc_250 N_A_80_27#_c_163_n N_VPWR_M1017_d 0.00593664f $X=0.675 $Y=2.3 $X2=-0.19
+ $Y2=-0.245
cc_251 N_A_80_27#_c_177_p N_VPWR_M1017_d 0.00830189f $X=1.63 $Y=2.385 $X2=-0.19
+ $Y2=-0.245
cc_252 N_A_80_27#_c_269_p N_VPWR_M1017_d 0.00245241f $X=0.795 $Y=2.385 $X2=-0.19
+ $Y2=-0.245
cc_253 N_A_80_27#_M1017_g N_VPWR_c_907_n 0.0128021f $X=0.485 $Y=2.465 $X2=0
+ $Y2=0
cc_254 N_A_80_27#_c_177_p N_VPWR_c_907_n 0.00705916f $X=1.63 $Y=2.385 $X2=0
+ $Y2=0
cc_255 N_A_80_27#_c_269_p N_VPWR_c_907_n 0.0159364f $X=0.795 $Y=2.385 $X2=0
+ $Y2=0
cc_256 N_A_80_27#_c_165_n N_VPWR_c_909_n 0.00528664f $X=5.535 $Y=1.61 $X2=0
+ $Y2=0
cc_257 N_A_80_27#_M1018_g N_VPWR_c_931_n 7.79229e-19 $X=5.515 $Y=2.265 $X2=0
+ $Y2=0
cc_258 N_A_80_27#_M1017_g N_VPWR_c_916_n 0.00564095f $X=0.485 $Y=2.465 $X2=0
+ $Y2=0
cc_259 N_A_80_27#_c_178_p N_VPWR_c_917_n 0.00417623f $X=1.775 $Y=2.385 $X2=0
+ $Y2=0
cc_260 N_A_80_27#_M1017_g N_VPWR_c_906_n 0.0104249f $X=0.485 $Y=2.465 $X2=0
+ $Y2=0
cc_261 N_A_80_27#_c_177_p N_VPWR_c_906_n 0.0246741f $X=1.63 $Y=2.385 $X2=0 $Y2=0
cc_262 N_A_80_27#_c_269_p N_VPWR_c_906_n 8.41524e-19 $X=0.795 $Y=2.385 $X2=0
+ $Y2=0
cc_263 N_A_80_27#_c_178_p N_VPWR_c_906_n 0.0083854f $X=1.775 $Y=2.385 $X2=0
+ $Y2=0
cc_264 N_A_80_27#_c_177_p A_231_457# 0.00737854f $X=1.63 $Y=2.385 $X2=-0.19
+ $Y2=-0.245
cc_265 N_A_80_27#_c_165_n N_A_417_457#_c_1010_n 0.00567252f $X=5.535 $Y=1.61
+ $X2=0 $Y2=0
cc_266 N_A_80_27#_c_165_n N_A_417_457#_c_1011_n 0.00268957f $X=5.535 $Y=1.61
+ $X2=0 $Y2=0
cc_267 N_A_80_27#_M1018_g N_A_854_411#_c_1035_n 0.00518877f $X=5.515 $Y=2.265
+ $X2=0 $Y2=0
cc_268 N_A_80_27#_c_165_n N_A_854_411#_c_1035_n 0.0621609f $X=5.535 $Y=1.61
+ $X2=0 $Y2=0
cc_269 N_A_80_27#_c_166_n N_A_854_411#_c_1035_n 0.00165659f $X=5.535 $Y=1.61
+ $X2=0 $Y2=0
cc_270 N_A_80_27#_c_165_n N_A_854_411#_c_1036_n 0.0190116f $X=5.535 $Y=1.61
+ $X2=0 $Y2=0
cc_271 N_A_80_27#_M1018_g N_A_854_411#_c_1037_n 9.29291e-19 $X=5.515 $Y=2.265
+ $X2=0 $Y2=0
cc_272 N_A_80_27#_c_164_n N_VGND_c_1089_n 0.0102502f $X=1.865 $Y=0.895 $X2=0
+ $Y2=0
cc_273 N_A_80_27#_c_167_n N_VGND_c_1089_n 0.0198162f $X=0.63 $Y=1.38 $X2=0 $Y2=0
cc_274 N_A_80_27#_c_168_n N_VGND_c_1089_n 0.00175752f $X=0.63 $Y=1.38 $X2=0
+ $Y2=0
cc_275 N_A_80_27#_c_169_n N_VGND_c_1089_n 0.015703f $X=0.597 $Y=1.215 $X2=0
+ $Y2=0
cc_276 N_A_80_27#_c_169_n N_VGND_c_1099_n 0.00498035f $X=0.597 $Y=1.215 $X2=0
+ $Y2=0
cc_277 N_A_80_27#_c_164_n N_VGND_c_1100_n 0.00368812f $X=1.865 $Y=0.895 $X2=0
+ $Y2=0
cc_278 N_A_80_27#_M1025_g N_VGND_c_1102_n 8.6132e-19 $X=5.555 $Y=0.835 $X2=0
+ $Y2=0
cc_279 N_A_80_27#_c_164_n N_VGND_c_1102_n 0.00684741f $X=1.865 $Y=0.895 $X2=0
+ $Y2=0
cc_280 N_A_80_27#_c_169_n N_VGND_c_1102_n 0.00961125f $X=0.597 $Y=1.215 $X2=0
+ $Y2=0
cc_281 N_A_80_27#_c_164_n N_A_431_137#_c_1185_n 0.0205239f $X=1.865 $Y=0.895
+ $X2=0 $Y2=0
cc_282 N_A_80_27#_c_165_n N_A_431_137#_c_1186_n 0.0637422f $X=5.535 $Y=1.61
+ $X2=0 $Y2=0
cc_283 N_A_80_27#_c_164_n N_A_431_137#_c_1187_n 0.0141076f $X=1.865 $Y=0.895
+ $X2=0 $Y2=0
cc_284 N_A_80_27#_c_165_n N_A_431_137#_c_1187_n 0.0192098f $X=5.535 $Y=1.61
+ $X2=0 $Y2=0
cc_285 N_A_80_27#_M1025_g N_A_818_83#_c_1215_n 0.00984869f $X=5.555 $Y=0.835
+ $X2=0 $Y2=0
cc_286 N_A_M1004_g N_B_M1026_g 0.0105378f $X=1.08 $Y=2.495 $X2=0 $Y2=0
cc_287 N_A_M1006_g N_B_M1026_g 0.0546252f $X=1.26 $Y=0.895 $X2=0 $Y2=0
cc_288 N_A_c_324_n N_B_M1026_g 0.00609722f $X=2.495 $Y=2.035 $X2=0 $Y2=0
cc_289 N_A_c_325_n N_B_M1026_g 6.94707e-19 $X=1.345 $Y=2.035 $X2=0 $Y2=0
cc_290 N_A_c_316_n N_B_M1026_g 0.00581311f $X=1.17 $Y=1.46 $X2=0 $Y2=0
cc_291 N_A_M1020_g N_B_c_515_n 0.00903575f $X=2.51 $Y=0.895 $X2=0 $Y2=0
cc_292 N_A_M1020_g N_B_M1021_g 0.0222413f $X=2.51 $Y=0.895 $X2=0 $Y2=0
cc_293 N_A_M1005_g N_B_M1012_g 0.017253f $X=2.44 $Y=2.495 $X2=0 $Y2=0
cc_294 N_A_M1020_g N_B_M1012_g 0.0131459f $X=2.51 $Y=0.895 $X2=0 $Y2=0
cc_295 N_A_c_326_n N_B_M1012_g 0.00547785f $X=6.815 $Y=2.035 $X2=0 $Y2=0
cc_296 N_A_c_327_n N_B_M1012_g 3.41389e-19 $X=2.785 $Y=2.035 $X2=0 $Y2=0
cc_297 N_A_c_331_n N_B_M1012_g 0.0167567f $X=2.53 $Y=1.96 $X2=0 $Y2=0
cc_298 N_A_c_332_n N_B_M1012_g 0.00243411f $X=2.53 $Y=1.96 $X2=0 $Y2=0
cc_299 N_A_c_326_n N_B_c_537_n 0.0069658f $X=6.815 $Y=2.035 $X2=0 $Y2=0
cc_300 N_A_c_323_n N_B_M1000_g 0.0229648f $X=7.035 $Y=1.855 $X2=0 $Y2=0
cc_301 N_A_c_326_n N_B_M1000_g 0.00547722f $X=6.815 $Y=2.035 $X2=0 $Y2=0
cc_302 N_A_c_328_n N_B_M1000_g 0.00126133f $X=6.96 $Y=2.035 $X2=0 $Y2=0
cc_303 N_A_c_314_n N_B_M1000_g 0.00414925f $X=7.035 $Y=1.35 $X2=0 $Y2=0
cc_304 N_A_M1004_g N_B_c_539_n 0.0278617f $X=1.08 $Y=2.495 $X2=0 $Y2=0
cc_305 N_A_c_324_n N_B_c_539_n 0.00293812f $X=2.495 $Y=2.035 $X2=0 $Y2=0
cc_306 N_A_c_325_n N_B_c_539_n 7.26499e-19 $X=1.345 $Y=2.035 $X2=0 $Y2=0
cc_307 N_A_c_316_n N_B_c_539_n 5.31406e-19 $X=1.17 $Y=1.46 $X2=0 $Y2=0
cc_308 N_A_c_326_n N_B_c_540_n 0.00381304f $X=6.815 $Y=2.035 $X2=0 $Y2=0
cc_309 N_A_c_307_n N_B_c_526_n 0.00839432f $X=6.87 $Y=0.18 $X2=0 $Y2=0
cc_310 N_A_M1009_g N_B_c_526_n 0.0191905f $X=6.945 $Y=0.835 $X2=0 $Y2=0
cc_311 N_A_c_313_n N_B_c_527_n 0.0122837f $X=7.035 $Y=1.35 $X2=0 $Y2=0
cc_312 N_A_c_312_n N_B_c_541_n 0.0122837f $X=7.035 $Y=1.69 $X2=0 $Y2=0
cc_313 N_A_c_326_n N_B_c_541_n 0.00503397f $X=6.815 $Y=2.035 $X2=0 $Y2=0
cc_314 N_A_M1010_g N_B_c_529_n 0.00578214f $X=5.085 $Y=2.265 $X2=0 $Y2=0
cc_315 N_A_c_311_n N_B_c_529_n 0.0122819f $X=5.085 $Y=1.195 $X2=0 $Y2=0
cc_316 N_A_c_326_n B 0.00665353f $X=6.815 $Y=2.035 $X2=0 $Y2=0
cc_317 N_A_c_326_n B 0.0218046f $X=6.815 $Y=2.035 $X2=0 $Y2=0
cc_318 N_A_c_313_n B 7.30898e-19 $X=7.035 $Y=1.35 $X2=0 $Y2=0
cc_319 N_A_c_314_n B 0.0489229f $X=7.035 $Y=1.35 $X2=0 $Y2=0
cc_320 N_A_M1009_g N_B_c_532_n 0.0122837f $X=6.945 $Y=0.835 $X2=0 $Y2=0
cc_321 N_A_c_314_n N_B_c_532_n 0.00218025f $X=7.035 $Y=1.35 $X2=0 $Y2=0
cc_322 N_A_M1005_g N_CIN_M1015_g 0.0108378f $X=2.44 $Y=2.495 $X2=0 $Y2=0
cc_323 N_A_M1020_g N_CIN_M1001_g 0.0377066f $X=2.51 $Y=0.895 $X2=0 $Y2=0
cc_324 N_A_c_324_n N_CIN_M1001_g 0.0031357f $X=2.495 $Y=2.035 $X2=0 $Y2=0
cc_325 N_A_c_331_n N_CIN_M1001_g 0.0132852f $X=2.53 $Y=1.96 $X2=0 $Y2=0
cc_326 N_A_c_332_n N_CIN_M1001_g 0.00108066f $X=2.53 $Y=1.96 $X2=0 $Y2=0
cc_327 N_A_M1005_g N_CIN_c_688_n 0.0100585f $X=2.44 $Y=2.495 $X2=0 $Y2=0
cc_328 N_A_M1007_g N_CIN_M1024_g 0.0295644f $X=4.895 $Y=0.625 $X2=0 $Y2=0
cc_329 N_A_M1010_g N_CIN_M1024_g 0.00554897f $X=5.085 $Y=2.265 $X2=0 $Y2=0
cc_330 N_A_c_326_n N_CIN_M1003_g 0.00601956f $X=6.815 $Y=2.035 $X2=0 $Y2=0
cc_331 N_A_M1010_g N_CIN_c_693_n 0.0106495f $X=5.085 $Y=2.265 $X2=0 $Y2=0
cc_332 N_A_c_307_n N_CIN_M1027_g 0.00839432f $X=6.87 $Y=0.18 $X2=0 $Y2=0
cc_333 N_A_c_326_n N_CIN_M1027_g 0.00485619f $X=6.815 $Y=2.035 $X2=0 $Y2=0
cc_334 N_A_M1005_g N_CIN_c_695_n 0.0132852f $X=2.44 $Y=2.495 $X2=0 $Y2=0
cc_335 N_A_c_324_n N_CIN_c_695_n 0.00828298f $X=2.495 $Y=2.035 $X2=0 $Y2=0
cc_336 N_A_M1010_g N_CIN_c_685_n 0.0355732f $X=5.085 $Y=2.265 $X2=0 $Y2=0
cc_337 N_A_c_326_n N_CIN_c_698_n 8.37852e-19 $X=6.815 $Y=2.035 $X2=0 $Y2=0
cc_338 N_A_c_326_n N_CIN_c_699_n 0.0241042f $X=6.815 $Y=2.035 $X2=0 $Y2=0
cc_339 N_A_c_327_n N_CIN_c_699_n 3.49882e-19 $X=2.785 $Y=2.035 $X2=0 $Y2=0
cc_340 N_A_c_332_n N_CIN_c_699_n 0.00488371f $X=2.53 $Y=1.96 $X2=0 $Y2=0
cc_341 N_A_c_326_n CIN 0.0045248f $X=6.815 $Y=2.035 $X2=0 $Y2=0
cc_342 N_A_c_326_n N_A_1118_411#_M1018_d 7.62208e-19 $X=6.815 $Y=2.035 $X2=0
+ $Y2=0
cc_343 N_A_M1019_g N_A_1118_411#_M1013_g 0.0116342f $X=6.945 $Y=2.265 $X2=0
+ $Y2=0
cc_344 N_A_c_312_n N_A_1118_411#_M1013_g 0.00819385f $X=7.035 $Y=1.69 $X2=0
+ $Y2=0
cc_345 N_A_c_314_n N_A_1118_411#_M1013_g 8.22149e-19 $X=7.035 $Y=1.35 $X2=0
+ $Y2=0
cc_346 N_A_c_307_n N_A_1118_411#_c_827_n 0.0142703f $X=6.87 $Y=0.18 $X2=0 $Y2=0
cc_347 N_A_M1019_g N_A_1118_411#_c_828_n 0.0133803f $X=6.945 $Y=2.265 $X2=0
+ $Y2=0
cc_348 N_A_c_323_n N_A_1118_411#_c_828_n 0.00279161f $X=7.035 $Y=1.855 $X2=0
+ $Y2=0
cc_349 N_A_c_326_n N_A_1118_411#_c_828_n 0.0288774f $X=6.815 $Y=2.035 $X2=0
+ $Y2=0
cc_350 N_A_c_328_n N_A_1118_411#_c_828_n 0.0076218f $X=6.96 $Y=2.035 $X2=0 $Y2=0
cc_351 N_A_c_314_n N_A_1118_411#_c_828_n 0.0139905f $X=7.035 $Y=1.35 $X2=0 $Y2=0
cc_352 N_A_M1009_g N_A_1118_411#_c_833_n 0.00530305f $X=6.945 $Y=0.835 $X2=0
+ $Y2=0
cc_353 N_A_c_313_n N_A_1118_411#_c_833_n 0.00389518f $X=7.035 $Y=1.35 $X2=0
+ $Y2=0
cc_354 N_A_M1019_g N_A_1118_411#_c_814_n 0.00487209f $X=6.945 $Y=2.265 $X2=0
+ $Y2=0
cc_355 N_A_c_323_n N_A_1118_411#_c_814_n 0.0018081f $X=7.035 $Y=1.855 $X2=0
+ $Y2=0
cc_356 N_A_c_328_n N_A_1118_411#_c_814_n 0.00260008f $X=6.96 $Y=2.035 $X2=0
+ $Y2=0
cc_357 N_A_c_326_n N_A_1118_411#_c_821_n 0.0184663f $X=6.815 $Y=2.035 $X2=0
+ $Y2=0
cc_358 N_A_M1009_g N_A_1118_411#_c_839_n 0.0153422f $X=6.945 $Y=0.835 $X2=0
+ $Y2=0
cc_359 N_A_c_314_n N_A_1118_411#_c_839_n 0.0197795f $X=7.035 $Y=1.35 $X2=0 $Y2=0
cc_360 N_A_c_312_n N_A_1118_411#_c_815_n 0.0018081f $X=7.035 $Y=1.69 $X2=0 $Y2=0
cc_361 N_A_c_313_n N_A_1118_411#_c_816_n 0.0204036f $X=7.035 $Y=1.35 $X2=0 $Y2=0
cc_362 N_A_c_314_n N_A_1118_411#_c_816_n 2.8795e-19 $X=7.035 $Y=1.35 $X2=0 $Y2=0
cc_363 N_A_M1009_g N_A_1118_411#_c_817_n 0.00334111f $X=6.945 $Y=0.835 $X2=0
+ $Y2=0
cc_364 N_A_c_313_n N_A_1118_411#_c_817_n 0.0018081f $X=7.035 $Y=1.35 $X2=0 $Y2=0
cc_365 N_A_c_314_n N_A_1118_411#_c_817_n 0.0736973f $X=7.035 $Y=1.35 $X2=0 $Y2=0
cc_366 N_A_c_307_n N_A_1118_411#_c_818_n 0.0210733f $X=6.87 $Y=0.18 $X2=0 $Y2=0
cc_367 N_A_c_313_n N_A_1118_411#_c_818_n 2.25951e-19 $X=7.035 $Y=1.35 $X2=0
+ $Y2=0
cc_368 N_A_c_326_n N_VPWR_M1002_s 0.00117908f $X=6.815 $Y=2.035 $X2=0 $Y2=0
cc_369 N_A_c_326_n N_VPWR_M1003_d 0.00207468f $X=6.815 $Y=2.035 $X2=0 $Y2=0
cc_370 N_A_c_328_n N_VPWR_M1019_d 8.61335e-19 $X=6.96 $Y=2.035 $X2=0 $Y2=0
cc_371 N_A_c_314_n N_VPWR_M1019_d 0.00100824f $X=7.035 $Y=1.35 $X2=0 $Y2=0
cc_372 N_A_M1004_g N_VPWR_c_907_n 0.00522923f $X=1.08 $Y=2.495 $X2=0 $Y2=0
cc_373 N_A_M1005_g N_VPWR_c_908_n 0.00415974f $X=2.44 $Y=2.495 $X2=0 $Y2=0
cc_374 N_A_c_326_n N_VPWR_c_909_n 0.015229f $X=6.815 $Y=2.035 $X2=0 $Y2=0
cc_375 N_A_M1010_g N_VPWR_c_910_n 0.00354658f $X=5.085 $Y=2.265 $X2=0 $Y2=0
cc_376 N_A_M1010_g N_VPWR_c_931_n 0.00331461f $X=5.085 $Y=2.265 $X2=0 $Y2=0
cc_377 N_A_c_326_n N_VPWR_c_931_n 0.00898092f $X=6.815 $Y=2.035 $X2=0 $Y2=0
cc_378 N_A_M1004_g N_VPWR_c_917_n 0.00415323f $X=1.08 $Y=2.495 $X2=0 $Y2=0
cc_379 N_A_M1019_g N_VPWR_c_918_n 0.00312414f $X=6.945 $Y=2.265 $X2=0 $Y2=0
cc_380 N_A_M1004_g N_VPWR_c_906_n 0.00469432f $X=1.08 $Y=2.495 $X2=0 $Y2=0
cc_381 N_A_M1005_g N_VPWR_c_906_n 9.03773e-19 $X=2.44 $Y=2.495 $X2=0 $Y2=0
cc_382 N_A_M1019_g N_VPWR_c_906_n 0.00410284f $X=6.945 $Y=2.265 $X2=0 $Y2=0
cc_383 N_A_M1005_g N_A_417_457#_c_1010_n 0.00898883f $X=2.44 $Y=2.495 $X2=0
+ $Y2=0
cc_384 N_A_c_324_n N_A_417_457#_c_1010_n 7.11786e-19 $X=2.495 $Y=2.035 $X2=0
+ $Y2=0
cc_385 N_A_c_326_n N_A_417_457#_c_1010_n 0.0160712f $X=6.815 $Y=2.035 $X2=0
+ $Y2=0
cc_386 N_A_c_327_n N_A_417_457#_c_1010_n 0.00806415f $X=2.785 $Y=2.035 $X2=0
+ $Y2=0
cc_387 N_A_c_331_n N_A_417_457#_c_1010_n 0.00112211f $X=2.53 $Y=1.96 $X2=0 $Y2=0
cc_388 N_A_c_332_n N_A_417_457#_c_1010_n 0.0237974f $X=2.53 $Y=1.96 $X2=0 $Y2=0
cc_389 N_A_M1005_g N_A_417_457#_c_1011_n 0.00528074f $X=2.44 $Y=2.495 $X2=0
+ $Y2=0
cc_390 N_A_c_324_n N_A_417_457#_c_1011_n 0.00856133f $X=2.495 $Y=2.035 $X2=0
+ $Y2=0
cc_391 N_A_c_332_n N_A_417_457#_c_1011_n 0.00159758f $X=2.53 $Y=1.96 $X2=0 $Y2=0
cc_392 N_A_c_326_n N_A_854_411#_M1002_d 0.00232013f $X=6.815 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_393 N_A_c_326_n N_A_854_411#_M1010_d 0.0016355f $X=6.815 $Y=2.035 $X2=0 $Y2=0
cc_394 N_A_c_326_n N_A_854_411#_c_1034_n 0.0167141f $X=6.815 $Y=2.035 $X2=0
+ $Y2=0
cc_395 N_A_M1010_g N_A_854_411#_c_1035_n 0.0111697f $X=5.085 $Y=2.265 $X2=0
+ $Y2=0
cc_396 N_A_c_326_n N_A_854_411#_c_1035_n 0.0273317f $X=6.815 $Y=2.035 $X2=0
+ $Y2=0
cc_397 N_A_c_326_n N_A_854_411#_c_1036_n 0.00663803f $X=6.815 $Y=2.035 $X2=0
+ $Y2=0
cc_398 N_A_M1010_g N_A_854_411#_c_1037_n 4.77646e-19 $X=5.085 $Y=2.265 $X2=0
+ $Y2=0
cc_399 N_A_c_326_n N_A_854_411#_c_1037_n 0.0165515f $X=6.815 $Y=2.035 $X2=0
+ $Y2=0
cc_400 N_A_c_326_n A_1212_411# 0.0019473f $X=6.815 $Y=2.035 $X2=-0.19 $Y2=-0.245
cc_401 N_A_c_326_n A_1290_411# 0.00310638f $X=6.815 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_402 N_A_c_328_n A_1290_411# 0.00124983f $X=6.96 $Y=2.035 $X2=-0.19 $Y2=-0.245
cc_403 N_A_M1006_g N_VGND_c_1089_n 0.0113927f $X=1.26 $Y=0.895 $X2=0 $Y2=0
cc_404 N_A_c_315_n N_VGND_c_1089_n 0.00112957f $X=1.17 $Y=1.46 $X2=0 $Y2=0
cc_405 N_A_c_316_n N_VGND_c_1089_n 0.0105138f $X=1.17 $Y=1.46 $X2=0 $Y2=0
cc_406 N_A_M1020_g N_VGND_c_1090_n 0.00836611f $X=2.51 $Y=0.895 $X2=0 $Y2=0
cc_407 N_A_M1007_g N_VGND_c_1093_n 0.0115381f $X=4.895 $Y=0.625 $X2=0 $Y2=0
cc_408 N_A_c_308_n N_VGND_c_1093_n 0.00763335f $X=4.97 $Y=0.18 $X2=0 $Y2=0
cc_409 N_A_c_307_n N_VGND_c_1094_n 0.0142976f $X=6.87 $Y=0.18 $X2=0 $Y2=0
cc_410 N_A_c_308_n N_VGND_c_1097_n 0.058408f $X=4.97 $Y=0.18 $X2=0 $Y2=0
cc_411 N_A_M1006_g N_VGND_c_1100_n 0.00345748f $X=1.26 $Y=0.895 $X2=0 $Y2=0
cc_412 N_A_M1006_g N_VGND_c_1102_n 0.00410867f $X=1.26 $Y=0.895 $X2=0 $Y2=0
cc_413 N_A_M1020_g N_VGND_c_1102_n 7.40973e-19 $X=2.51 $Y=0.895 $X2=0 $Y2=0
cc_414 N_A_c_307_n N_VGND_c_1102_n 0.0578582f $X=6.87 $Y=0.18 $X2=0 $Y2=0
cc_415 N_A_c_308_n N_VGND_c_1102_n 0.00373117f $X=4.97 $Y=0.18 $X2=0 $Y2=0
cc_416 N_A_M1020_g N_A_431_137#_c_1185_n 0.00116371f $X=2.51 $Y=0.895 $X2=0
+ $Y2=0
cc_417 N_A_M1020_g N_A_431_137#_c_1186_n 0.0140415f $X=2.51 $Y=0.895 $X2=0 $Y2=0
cc_418 N_A_M1007_g N_A_818_83#_c_1213_n 0.0112534f $X=4.895 $Y=0.625 $X2=0 $Y2=0
cc_419 N_A_c_311_n N_A_818_83#_c_1213_n 9.44079e-19 $X=5.085 $Y=1.195 $X2=0
+ $Y2=0
cc_420 N_A_M1007_g N_A_818_83#_c_1215_n 0.0018698f $X=4.895 $Y=0.625 $X2=0 $Y2=0
cc_421 N_A_c_307_n N_A_818_83#_c_1215_n 0.00977102f $X=6.87 $Y=0.18 $X2=0 $Y2=0
cc_422 N_A_c_311_n N_A_818_83#_c_1215_n 0.00411816f $X=5.085 $Y=1.195 $X2=0
+ $Y2=0
cc_423 N_B_c_539_n N_CIN_M1015_g 0.0105483f $X=1.615 $Y=2.21 $X2=0 $Y2=0
cc_424 N_B_M1026_g N_CIN_M1001_g 0.0476941f $X=1.65 $Y=0.895 $X2=0 $Y2=0
cc_425 N_B_c_515_n N_CIN_M1001_g 0.00918179f $X=2.865 $Y=0.24 $X2=0 $Y2=0
cc_426 N_B_M1012_g N_CIN_c_688_n 0.0100585f $X=3.03 $Y=2.495 $X2=0 $Y2=0
cc_427 N_B_M1012_g N_CIN_c_690_n 0.0118548f $X=3.03 $Y=2.495 $X2=0 $Y2=0
cc_428 N_B_c_537_n N_CIN_c_691_n 0.0108224f $X=4.195 $Y=1.98 $X2=0 $Y2=0
cc_429 N_B_M1022_g N_CIN_M1024_g 0.017977f $X=4.015 $Y=0.625 $X2=0 $Y2=0
cc_430 N_B_c_529_n N_CIN_M1024_g 0.011529f $X=5.495 $Y=1.27 $X2=0 $Y2=0
cc_431 N_B_c_533_n N_CIN_M1024_g 0.0180349f $X=4.015 $Y=1.23 $X2=0 $Y2=0
cc_432 N_B_c_523_n N_CIN_M1003_g 0.00389438f $X=4.09 $Y=1.83 $X2=0 $Y2=0
cc_433 N_B_c_540_n N_CIN_M1003_g 0.0152022f $X=4.195 $Y=1.905 $X2=0 $Y2=0
cc_434 N_B_c_526_n N_CIN_M1027_g 0.11826f $X=6.465 $Y=1.155 $X2=0 $Y2=0
cc_435 B N_CIN_M1027_g 0.00202331f $X=5.915 $Y=1.21 $X2=0 $Y2=0
cc_436 B N_CIN_M1027_g 0.0260253f $X=6.395 $Y=1.21 $X2=0 $Y2=0
cc_437 N_B_c_539_n N_CIN_c_695_n 0.00930541f $X=1.615 $Y=2.21 $X2=0 $Y2=0
cc_438 N_B_c_523_n N_CIN_c_685_n 0.0180349f $X=4.09 $Y=1.83 $X2=0 $Y2=0
cc_439 N_B_c_529_n N_CIN_c_685_n 0.00529209f $X=5.495 $Y=1.27 $X2=0 $Y2=0
cc_440 N_B_M1012_g N_CIN_c_698_n 0.0168745f $X=3.03 $Y=2.495 $X2=0 $Y2=0
cc_441 N_B_c_520_n N_CIN_c_698_n 0.00946893f $X=3.45 $Y=1.35 $X2=0 $Y2=0
cc_442 N_B_c_523_n N_CIN_c_698_n 0.00766264f $X=4.09 $Y=1.83 $X2=0 $Y2=0
cc_443 N_B_c_537_n N_CIN_c_698_n 0.010611f $X=4.195 $Y=1.98 $X2=0 $Y2=0
cc_444 N_B_M1012_g N_CIN_c_699_n 0.00111486f $X=3.03 $Y=2.495 $X2=0 $Y2=0
cc_445 N_B_c_537_n N_CIN_c_699_n 5.82851e-19 $X=4.195 $Y=1.98 $X2=0 $Y2=0
cc_446 N_B_c_540_n N_CIN_c_699_n 0.00100768f $X=4.195 $Y=1.905 $X2=0 $Y2=0
cc_447 N_B_M1012_g CIN 0.00436759f $X=3.03 $Y=2.495 $X2=0 $Y2=0
cc_448 N_B_c_526_n N_A_1118_411#_c_827_n 0.0185207f $X=6.465 $Y=1.155 $X2=0
+ $Y2=0
cc_449 B N_A_1118_411#_c_827_n 0.0682366f $X=5.915 $Y=1.21 $X2=0 $Y2=0
cc_450 N_B_c_532_n N_A_1118_411#_c_827_n 0.00475889f $X=6.465 $Y=1.32 $X2=0
+ $Y2=0
cc_451 N_B_M1000_g N_A_1118_411#_c_828_n 0.0132268f $X=6.375 $Y=2.265 $X2=0
+ $Y2=0
cc_452 N_B_c_541_n N_A_1118_411#_c_828_n 0.00349396f $X=6.465 $Y=1.825 $X2=0
+ $Y2=0
cc_453 B N_A_1118_411#_c_828_n 0.0101121f $X=6.395 $Y=1.21 $X2=0 $Y2=0
cc_454 N_B_M1012_g N_VPWR_c_908_n 0.00243468f $X=3.03 $Y=2.495 $X2=0 $Y2=0
cc_455 N_B_c_537_n N_VPWR_c_909_n 0.00387809f $X=4.195 $Y=1.98 $X2=0 $Y2=0
cc_456 N_B_c_540_n N_VPWR_c_909_n 0.00224377f $X=4.195 $Y=1.905 $X2=0 $Y2=0
cc_457 N_B_c_539_n N_VPWR_c_917_n 0.004006f $X=1.615 $Y=2.21 $X2=0 $Y2=0
cc_458 N_B_M1000_g N_VPWR_c_918_n 0.00312414f $X=6.375 $Y=2.265 $X2=0 $Y2=0
cc_459 N_B_M1012_g N_VPWR_c_906_n 9.03773e-19 $X=3.03 $Y=2.495 $X2=0 $Y2=0
cc_460 N_B_M1000_g N_VPWR_c_906_n 0.00410284f $X=6.375 $Y=2.265 $X2=0 $Y2=0
cc_461 N_B_c_539_n N_VPWR_c_906_n 0.00469432f $X=1.615 $Y=2.21 $X2=0 $Y2=0
cc_462 N_B_M1012_g N_A_417_457#_c_1010_n 0.0150607f $X=3.03 $Y=2.495 $X2=0 $Y2=0
cc_463 N_B_M1012_g N_A_417_457#_c_1011_n 8.54391e-19 $X=3.03 $Y=2.495 $X2=0
+ $Y2=0
cc_464 N_B_c_537_n N_A_854_411#_c_1034_n 4.73302e-19 $X=4.195 $Y=1.98 $X2=0
+ $Y2=0
cc_465 N_B_c_540_n N_A_854_411#_c_1036_n 0.00266927f $X=4.195 $Y=1.905 $X2=0
+ $Y2=0
cc_466 N_B_M1026_g N_VGND_c_1089_n 0.0017151f $X=1.65 $Y=0.895 $X2=0 $Y2=0
cc_467 N_B_c_516_n N_VGND_c_1089_n 0.0123346f $X=1.725 $Y=0.24 $X2=0 $Y2=0
cc_468 N_B_c_515_n N_VGND_c_1090_n 0.0201525f $X=2.865 $Y=0.24 $X2=0 $Y2=0
cc_469 N_B_M1021_g N_VGND_c_1090_n 0.0209635f $X=2.94 $Y=0.895 $X2=0 $Y2=0
cc_470 N_B_c_521_n N_VGND_c_1090_n 0.00152606f $X=3.525 $Y=1.035 $X2=0 $Y2=0
cc_471 N_B_c_524_n N_VGND_c_1090_n 0.00606056f $X=2.94 $Y=0.24 $X2=0 $Y2=0
cc_472 N_B_c_519_n N_VGND_c_1091_n 0.0186888f $X=3.45 $Y=0.24 $X2=0 $Y2=0
cc_473 N_B_M1022_g N_VGND_c_1091_n 0.00211334f $X=4.015 $Y=0.625 $X2=0 $Y2=0
cc_474 N_B_c_528_n N_VGND_c_1091_n 0.00892881f $X=3.805 $Y=1.225 $X2=0 $Y2=0
cc_475 N_B_c_529_n N_VGND_c_1091_n 0.00528921f $X=5.495 $Y=1.27 $X2=0 $Y2=0
cc_476 N_B_c_533_n N_VGND_c_1091_n 0.00383536f $X=4.015 $Y=1.23 $X2=0 $Y2=0
cc_477 N_B_M1022_g N_VGND_c_1092_n 0.00545098f $X=4.015 $Y=0.625 $X2=0 $Y2=0
cc_478 N_B_M1022_g N_VGND_c_1093_n 5.13269e-19 $X=4.015 $Y=0.625 $X2=0 $Y2=0
cc_479 N_B_c_524_n N_VGND_c_1095_n 0.0220223f $X=2.94 $Y=0.24 $X2=0 $Y2=0
cc_480 N_B_c_516_n N_VGND_c_1100_n 0.0273241f $X=1.725 $Y=0.24 $X2=0 $Y2=0
cc_481 N_B_c_515_n N_VGND_c_1102_n 0.0269567f $X=2.865 $Y=0.24 $X2=0 $Y2=0
cc_482 N_B_c_516_n N_VGND_c_1102_n 0.00991645f $X=1.725 $Y=0.24 $X2=0 $Y2=0
cc_483 N_B_c_519_n N_VGND_c_1102_n 0.029643f $X=3.45 $Y=0.24 $X2=0 $Y2=0
cc_484 N_B_M1022_g N_VGND_c_1102_n 0.005315f $X=4.015 $Y=0.625 $X2=0 $Y2=0
cc_485 N_B_c_524_n N_VGND_c_1102_n 0.00755648f $X=2.94 $Y=0.24 $X2=0 $Y2=0
cc_486 N_B_c_526_n N_VGND_c_1102_n 9.49986e-19 $X=6.465 $Y=1.155 $X2=0 $Y2=0
cc_487 N_B_c_515_n N_A_431_137#_c_1185_n 0.00405167f $X=2.865 $Y=0.24 $X2=0
+ $Y2=0
cc_488 N_B_M1021_g N_A_431_137#_c_1186_n 0.00819573f $X=2.94 $Y=0.895 $X2=0
+ $Y2=0
cc_489 N_B_c_520_n N_A_431_137#_c_1186_n 0.0082752f $X=3.45 $Y=1.35 $X2=0 $Y2=0
cc_490 N_B_c_525_n N_A_431_137#_c_1186_n 0.00540779f $X=2.985 $Y=1.35 $X2=0
+ $Y2=0
cc_491 N_B_c_528_n N_A_431_137#_c_1186_n 0.0147131f $X=3.805 $Y=1.225 $X2=0
+ $Y2=0
cc_492 N_B_M1021_g N_A_431_137#_c_1188_n 0.00133795f $X=2.94 $Y=0.895 $X2=0
+ $Y2=0
cc_493 N_B_c_519_n N_A_431_137#_c_1188_n 0.0033301f $X=3.45 $Y=0.24 $X2=0 $Y2=0
cc_494 N_B_c_521_n N_A_431_137#_c_1188_n 0.00773587f $X=3.525 $Y=1.035 $X2=0
+ $Y2=0
cc_495 N_B_c_528_n N_A_431_137#_c_1188_n 0.00704938f $X=3.805 $Y=1.225 $X2=0
+ $Y2=0
cc_496 N_B_c_533_n N_A_431_137#_c_1188_n 3.26879e-19 $X=4.015 $Y=1.23 $X2=0
+ $Y2=0
cc_497 N_B_c_529_n N_A_818_83#_c_1213_n 0.048652f $X=5.495 $Y=1.27 $X2=0 $Y2=0
cc_498 N_B_M1022_g N_A_818_83#_c_1214_n 0.00534941f $X=4.015 $Y=0.625 $X2=0
+ $Y2=0
cc_499 N_B_c_529_n N_A_818_83#_c_1214_n 0.0198853f $X=5.495 $Y=1.27 $X2=0 $Y2=0
cc_500 N_B_c_533_n N_A_818_83#_c_1214_n 0.00176202f $X=4.015 $Y=1.23 $X2=0 $Y2=0
cc_501 N_B_c_529_n N_A_818_83#_c_1215_n 0.036589f $X=5.495 $Y=1.27 $X2=0 $Y2=0
cc_502 N_CIN_M1027_g N_A_1118_411#_c_827_n 0.0129579f $X=5.985 $Y=0.835 $X2=0
+ $Y2=0
cc_503 N_CIN_M1027_g N_A_1118_411#_c_828_n 0.010782f $X=5.985 $Y=0.835 $X2=0
+ $Y2=0
cc_504 N_CIN_c_693_n N_A_1118_411#_c_821_n 0.00598936f $X=5.91 $Y=2.89 $X2=0
+ $Y2=0
cc_505 N_CIN_M1015_g N_VPWR_c_908_n 0.00586615f $X=2.01 $Y=2.495 $X2=0 $Y2=0
cc_506 N_CIN_c_688_n N_VPWR_c_908_n 0.0268152f $X=3.545 $Y=3.12 $X2=0 $Y2=0
cc_507 N_CIN_c_690_n N_VPWR_c_908_n 6.12907e-19 $X=3.62 $Y=2.815 $X2=0 $Y2=0
cc_508 N_CIN_c_696_n N_VPWR_c_908_n 0.00249565f $X=3.62 $Y=2.89 $X2=0 $Y2=0
cc_509 CIN N_VPWR_c_908_n 0.00848307f $X=3.515 $Y=2.32 $X2=0 $Y2=0
cc_510 N_CIN_c_691_n N_VPWR_c_909_n 0.0236583f $X=4.58 $Y=2.89 $X2=0 $Y2=0
cc_511 N_CIN_M1003_g N_VPWR_c_909_n 0.00345876f $X=4.655 $Y=2.265 $X2=0 $Y2=0
cc_512 N_CIN_c_696_n N_VPWR_c_909_n 0.00770416f $X=3.62 $Y=2.89 $X2=0 $Y2=0
cc_513 N_CIN_c_698_n N_VPWR_c_909_n 0.00324352f $X=3.53 $Y=1.96 $X2=0 $Y2=0
cc_514 N_CIN_c_699_n N_VPWR_c_909_n 0.00148292f $X=3.61 $Y=1.992 $X2=0 $Y2=0
cc_515 CIN N_VPWR_c_909_n 0.0628228f $X=3.515 $Y=2.32 $X2=0 $Y2=0
cc_516 N_CIN_M1003_g N_VPWR_c_910_n 0.011416f $X=4.655 $Y=2.265 $X2=0 $Y2=0
cc_517 N_CIN_c_693_n N_VPWR_c_910_n 0.0242822f $X=5.91 $Y=2.89 $X2=0 $Y2=0
cc_518 N_CIN_c_688_n N_VPWR_c_912_n 0.0224731f $X=3.545 $Y=3.12 $X2=0 $Y2=0
cc_519 N_CIN_c_691_n N_VPWR_c_912_n 0.00536658f $X=4.58 $Y=2.89 $X2=0 $Y2=0
cc_520 CIN N_VPWR_c_912_n 0.00750212f $X=3.515 $Y=2.32 $X2=0 $Y2=0
cc_521 N_CIN_M1003_g N_VPWR_c_931_n 0.00388695f $X=4.655 $Y=2.265 $X2=0 $Y2=0
cc_522 N_CIN_c_693_n N_VPWR_c_931_n 7.50704e-19 $X=5.91 $Y=2.89 $X2=0 $Y2=0
cc_523 N_CIN_c_691_n N_VPWR_c_914_n 0.0211062f $X=4.58 $Y=2.89 $X2=0 $Y2=0
cc_524 N_CIN_c_689_n N_VPWR_c_917_n 0.0190918f $X=2.085 $Y=3.12 $X2=0 $Y2=0
cc_525 N_CIN_c_693_n N_VPWR_c_918_n 0.0284356f $X=5.91 $Y=2.89 $X2=0 $Y2=0
cc_526 N_CIN_c_688_n N_VPWR_c_906_n 0.0367652f $X=3.545 $Y=3.12 $X2=0 $Y2=0
cc_527 N_CIN_c_689_n N_VPWR_c_906_n 0.0111398f $X=2.085 $Y=3.12 $X2=0 $Y2=0
cc_528 N_CIN_c_691_n N_VPWR_c_906_n 0.0567958f $X=4.58 $Y=2.89 $X2=0 $Y2=0
cc_529 N_CIN_c_696_n N_VPWR_c_906_n 0.00568549f $X=3.62 $Y=2.89 $X2=0 $Y2=0
cc_530 CIN N_VPWR_c_906_n 0.0065542f $X=3.515 $Y=2.32 $X2=0 $Y2=0
cc_531 N_CIN_c_688_n N_A_417_457#_c_1010_n 0.00587421f $X=3.545 $Y=3.12 $X2=0
+ $Y2=0
cc_532 N_CIN_c_690_n N_A_417_457#_c_1010_n 0.00124724f $X=3.62 $Y=2.815 $X2=0
+ $Y2=0
cc_533 CIN N_A_417_457#_c_1010_n 0.0278878f $X=3.515 $Y=2.32 $X2=0 $Y2=0
cc_534 N_CIN_c_688_n N_A_417_457#_c_1011_n 0.00331374f $X=3.545 $Y=3.12 $X2=0
+ $Y2=0
cc_535 N_CIN_c_695_n N_A_417_457#_c_1011_n 0.00180746f $X=2.045 $Y=2.21 $X2=0
+ $Y2=0
cc_536 N_CIN_c_691_n N_A_854_411#_c_1034_n 0.00565055f $X=4.58 $Y=2.89 $X2=0
+ $Y2=0
cc_537 N_CIN_M1003_g N_A_854_411#_c_1034_n 4.92491e-19 $X=4.655 $Y=2.265 $X2=0
+ $Y2=0
cc_538 N_CIN_c_699_n N_A_854_411#_c_1034_n 9.92335e-19 $X=3.61 $Y=1.992 $X2=0
+ $Y2=0
cc_539 N_CIN_M1003_g N_A_854_411#_c_1035_n 0.0114325f $X=4.655 $Y=2.265 $X2=0
+ $Y2=0
cc_540 N_CIN_c_685_n N_A_854_411#_c_1035_n 2.68316e-19 $X=4.655 $Y=1.555 $X2=0
+ $Y2=0
cc_541 N_CIN_c_685_n N_A_854_411#_c_1036_n 0.00103626f $X=4.655 $Y=1.555 $X2=0
+ $Y2=0
cc_542 N_CIN_c_699_n N_A_854_411#_c_1036_n 0.00506255f $X=3.61 $Y=1.992 $X2=0
+ $Y2=0
cc_543 N_CIN_c_693_n N_A_854_411#_c_1037_n 0.00609577f $X=5.91 $Y=2.89 $X2=0
+ $Y2=0
cc_544 N_CIN_M1001_g N_VGND_c_1090_n 8.69157e-19 $X=2.08 $Y=0.895 $X2=0 $Y2=0
cc_545 N_CIN_M1024_g N_VGND_c_1092_n 0.00507464f $X=4.45 $Y=0.625 $X2=0 $Y2=0
cc_546 N_CIN_M1024_g N_VGND_c_1093_n 0.006721f $X=4.45 $Y=0.625 $X2=0 $Y2=0
cc_547 N_CIN_M1001_g N_VGND_c_1102_n 8.82111e-19 $X=2.08 $Y=0.895 $X2=0 $Y2=0
cc_548 N_CIN_M1024_g N_VGND_c_1102_n 0.0049961f $X=4.45 $Y=0.625 $X2=0 $Y2=0
cc_549 N_CIN_M1027_g N_VGND_c_1102_n 9.49986e-19 $X=5.985 $Y=0.835 $X2=0 $Y2=0
cc_550 N_CIN_M1001_g N_A_431_137#_c_1185_n 7.117e-19 $X=2.08 $Y=0.895 $X2=0
+ $Y2=0
cc_551 N_CIN_M1001_g N_A_431_137#_c_1187_n 0.00154364f $X=2.08 $Y=0.895 $X2=0
+ $Y2=0
cc_552 N_CIN_M1024_g N_A_818_83#_c_1213_n 0.0114589f $X=4.45 $Y=0.625 $X2=0
+ $Y2=0
cc_553 N_CIN_M1027_g N_A_818_83#_c_1215_n 7.48399e-19 $X=5.985 $Y=0.835 $X2=0
+ $Y2=0
cc_554 N_A_1118_411#_c_828_n N_VPWR_M1019_d 0.0142304f $X=7.29 $Y=2.385 $X2=0
+ $Y2=0
cc_555 N_A_1118_411#_c_814_n N_VPWR_M1019_d 0.00553387f $X=7.457 $Y=2.3 $X2=0
+ $Y2=0
cc_556 N_A_1118_411#_M1013_g N_VPWR_c_911_n 0.0126992f $X=7.685 $Y=2.465 $X2=0
+ $Y2=0
cc_557 N_A_1118_411#_c_828_n N_VPWR_c_911_n 0.0234911f $X=7.29 $Y=2.385 $X2=0
+ $Y2=0
cc_558 N_A_1118_411#_M1013_g N_VPWR_c_919_n 0.00564095f $X=7.685 $Y=2.465 $X2=0
+ $Y2=0
cc_559 N_A_1118_411#_M1013_g N_VPWR_c_906_n 0.0100928f $X=7.685 $Y=2.465 $X2=0
+ $Y2=0
cc_560 N_A_1118_411#_c_828_n N_VPWR_c_906_n 0.0478893f $X=7.29 $Y=2.385 $X2=0
+ $Y2=0
cc_561 N_A_1118_411#_c_821_n N_VPWR_c_906_n 0.00978655f $X=5.77 $Y=2.265 $X2=0
+ $Y2=0
cc_562 N_A_1118_411#_c_828_n A_1212_411# 0.00448144f $X=7.29 $Y=2.385 $X2=-0.19
+ $Y2=-0.245
cc_563 N_A_1118_411#_c_828_n A_1290_411# 0.0108055f $X=7.29 $Y=2.385 $X2=-0.19
+ $Y2=-0.245
cc_564 N_A_1118_411#_M1013_g N_SUM_c_1071_n 0.00339074f $X=7.685 $Y=2.465 $X2=0
+ $Y2=0
cc_565 N_A_1118_411#_c_814_n N_SUM_c_1071_n 0.0189738f $X=7.457 $Y=2.3 $X2=0
+ $Y2=0
cc_566 N_A_1118_411#_c_814_n N_SUM_c_1068_n 0.0190171f $X=7.457 $Y=2.3 $X2=0
+ $Y2=0
cc_567 N_A_1118_411#_c_815_n N_SUM_c_1068_n 0.0245628f $X=7.575 $Y=1.355 $X2=0
+ $Y2=0
cc_568 N_A_1118_411#_c_816_n N_SUM_c_1068_n 0.0149618f $X=7.575 $Y=1.355 $X2=0
+ $Y2=0
cc_569 N_A_1118_411#_c_817_n N_SUM_c_1068_n 0.0069059f $X=7.475 $Y=1.19 $X2=0
+ $Y2=0
cc_570 N_A_1118_411#_c_818_n N_SUM_c_1068_n 0.00286205f $X=7.585 $Y=1.19 $X2=0
+ $Y2=0
cc_571 N_A_1118_411#_c_815_n SUM 9.98037e-19 $X=7.575 $Y=1.355 $X2=0 $Y2=0
cc_572 N_A_1118_411#_c_816_n SUM 0.00499436f $X=7.575 $Y=1.355 $X2=0 $Y2=0
cc_573 N_A_1118_411#_c_833_n N_VGND_M1009_d 0.00917294f $X=7.29 $Y=0.93 $X2=0
+ $Y2=0
cc_574 N_A_1118_411#_c_817_n N_VGND_M1009_d 7.44326e-19 $X=7.475 $Y=1.19 $X2=0
+ $Y2=0
cc_575 N_A_1118_411#_c_833_n N_VGND_c_1094_n 0.0223954f $X=7.29 $Y=0.93 $X2=0
+ $Y2=0
cc_576 N_A_1118_411#_c_839_n N_VGND_c_1094_n 7.41633e-19 $X=6.97 $Y=0.84 $X2=0
+ $Y2=0
cc_577 N_A_1118_411#_c_818_n N_VGND_c_1094_n 0.0120547f $X=7.585 $Y=1.19 $X2=0
+ $Y2=0
cc_578 N_A_1118_411#_c_827_n N_VGND_c_1097_n 0.019428f $X=6.795 $Y=0.84 $X2=0
+ $Y2=0
cc_579 N_A_1118_411#_c_818_n N_VGND_c_1101_n 0.00486043f $X=7.585 $Y=1.19 $X2=0
+ $Y2=0
cc_580 N_A_1118_411#_c_827_n N_VGND_c_1102_n 0.0319253f $X=6.795 $Y=0.84 $X2=0
+ $Y2=0
cc_581 N_A_1118_411#_c_833_n N_VGND_c_1102_n 0.00662452f $X=7.29 $Y=0.93 $X2=0
+ $Y2=0
cc_582 N_A_1118_411#_c_818_n N_VGND_c_1102_n 0.00930295f $X=7.585 $Y=1.19 $X2=0
+ $Y2=0
cc_583 N_A_1118_411#_c_827_n A_1212_125# 0.00323555f $X=6.795 $Y=0.84 $X2=-0.19
+ $Y2=-0.245
cc_584 N_A_1118_411#_c_827_n A_1290_125# 0.013294f $X=6.795 $Y=0.84 $X2=-0.19
+ $Y2=-0.245
cc_585 N_A_1118_411#_c_839_n A_1290_125# 0.00108193f $X=6.97 $Y=0.84 $X2=-0.19
+ $Y2=-0.245
cc_586 COUT N_VPWR_c_916_n 0.0195996f $X=0.24 $Y=2.035 $X2=0 $Y2=0
cc_587 N_COUT_M1017_s N_VPWR_c_906_n 0.00336915f $X=0.145 $Y=1.835 $X2=0 $Y2=0
cc_588 COUT N_VPWR_c_906_n 0.0111968f $X=0.24 $Y=2.035 $X2=0 $Y2=0
cc_589 N_COUT_c_890_n N_VGND_c_1089_n 0.0333587f $X=0.26 $Y=0.42 $X2=0 $Y2=0
cc_590 N_COUT_c_890_n N_VGND_c_1099_n 0.0199289f $X=0.26 $Y=0.42 $X2=0 $Y2=0
cc_591 N_COUT_c_890_n N_VGND_c_1102_n 0.010808f $X=0.26 $Y=0.42 $X2=0 $Y2=0
cc_592 N_VPWR_M1005_d N_A_417_457#_c_1010_n 0.00752482f $X=2.515 $Y=2.285 $X2=0
+ $Y2=0
cc_593 N_VPWR_c_908_n N_A_417_457#_c_1010_n 0.0249794f $X=2.735 $Y=2.755 $X2=0
+ $Y2=0
cc_594 N_VPWR_c_912_n N_A_417_457#_c_1010_n 0.00382193f $X=3.885 $Y=3.33 $X2=0
+ $Y2=0
cc_595 N_VPWR_c_906_n N_A_417_457#_c_1010_n 0.0173462f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_596 N_VPWR_c_917_n N_A_417_457#_c_1011_n 0.00417657f $X=2.57 $Y=3.33 $X2=0
+ $Y2=0
cc_597 N_VPWR_c_906_n N_A_417_457#_c_1011_n 0.00735281f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_598 N_VPWR_c_909_n N_A_854_411#_c_1034_n 0.013111f $X=3.98 $Y=2.265 $X2=0
+ $Y2=0
cc_599 N_VPWR_c_931_n N_A_854_411#_c_1035_n 0.0185457f $X=4.87 $Y=2.305 $X2=0
+ $Y2=0
cc_600 N_VPWR_c_906_n N_SUM_M1013_d 0.00336915f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_601 N_VPWR_c_919_n N_SUM_c_1072_n 0.0188828f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_602 N_VPWR_c_906_n N_SUM_c_1072_n 0.010808f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_603 N_SUM_c_1070_n N_VGND_c_1101_n 0.0303288f $X=7.755 $Y=0.42 $X2=0 $Y2=0
cc_604 N_SUM_M1023_d N_VGND_c_1102_n 0.00388458f $X=7.595 $Y=0.235 $X2=0 $Y2=0
cc_605 N_SUM_c_1070_n N_VGND_c_1102_n 0.016834f $X=7.755 $Y=0.42 $X2=0 $Y2=0
cc_606 N_VGND_c_1100_n N_A_431_137#_c_1185_n 0.00312836f $X=2.56 $Y=0 $X2=0
+ $Y2=0
cc_607 N_VGND_c_1102_n N_A_431_137#_c_1185_n 0.0056606f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_608 N_VGND_c_1090_n N_A_431_137#_c_1186_n 0.0216087f $X=2.725 $Y=0.895 $X2=0
+ $Y2=0
cc_609 N_VGND_c_1091_n N_A_431_137#_c_1188_n 0.00302314f $X=3.8 $Y=0.63 $X2=0
+ $Y2=0
cc_610 N_VGND_c_1095_n N_A_431_137#_c_1188_n 0.00334465f $X=3.635 $Y=0 $X2=0
+ $Y2=0
cc_611 N_VGND_c_1102_n N_A_431_137#_c_1188_n 0.00529619f $X=7.92 $Y=0 $X2=0
+ $Y2=0
cc_612 N_VGND_c_1092_n N_A_818_83#_c_1229_n 0.00598645f $X=4.515 $Y=0 $X2=0
+ $Y2=0
cc_613 N_VGND_c_1102_n N_A_818_83#_c_1229_n 0.00807755f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_614 N_VGND_M1024_d N_A_818_83#_c_1213_n 0.00189577f $X=4.525 $Y=0.415 $X2=0
+ $Y2=0
cc_615 N_VGND_c_1093_n N_A_818_83#_c_1213_n 0.0167557f $X=4.68 $Y=0.54 $X2=0
+ $Y2=0
cc_616 N_VGND_c_1102_n N_A_818_83#_c_1213_n 0.0114528f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_617 N_VGND_c_1093_n N_A_818_83#_c_1215_n 0.0114079f $X=4.68 $Y=0.54 $X2=0
+ $Y2=0
cc_618 N_VGND_c_1097_n N_A_818_83#_c_1215_n 0.0185312f $X=7.14 $Y=0 $X2=0 $Y2=0
cc_619 N_VGND_c_1102_n N_A_818_83#_c_1215_n 0.0152915f $X=7.92 $Y=0 $X2=0 $Y2=0
