* File: sky130_fd_sc_lp__sdfxbp_2.pex.spice
* Created: Wed Sep  2 10:36:16 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__SDFXBP_2%SCD 3 6 9 10 11 12 13 14 25
c31 14 0 1.20585e-19 $X=0.72 $Y=2.035
r32 13 14 6.29568 $w=7.17e-07 $l=3.7e-07 $layer=LI1_cond $X=0.445 $Y=1.665
+ $X2=0.445 $Y2=2.035
r33 12 13 6.29568 $w=7.17e-07 $l=3.7e-07 $layer=LI1_cond $X=0.445 $Y=1.295
+ $X2=0.445 $Y2=1.665
r34 12 25 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.385
+ $Y=1.295 $X2=0.385 $Y2=1.295
r35 10 25 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.385 $Y=1.635
+ $X2=0.385 $Y2=1.295
r36 10 11 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.385 $Y=1.635
+ $X2=0.385 $Y2=1.8
r37 9 25 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.385 $Y=1.13
+ $X2=0.385 $Y2=1.295
r38 6 11 494.819 $w=1.5e-07 $l=9.65e-07 $layer=POLY_cond $X=0.475 $Y=2.765
+ $X2=0.475 $Y2=1.8
r39 3 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.475 $Y=0.81
+ $X2=0.475 $Y2=1.13
.ends

.subckt PM_SKY130_FD_SC_LP__SDFXBP_2%D 3 7 11 12 13 15 22
c45 7 0 1.20585e-19 $X=1.305 $Y=2.765
r46 22 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.285
+ $Y=1.47 $X2=1.285 $Y2=1.47
r47 15 23 6.4279 $w=7.33e-07 $l=3.95e-07 $layer=LI1_cond $X=1.68 $Y=1.752
+ $X2=1.285 $Y2=1.752
r48 13 23 1.38322 $w=7.33e-07 $l=8.5e-08 $layer=LI1_cond $X=1.2 $Y=1.752
+ $X2=1.285 $Y2=1.752
r49 11 22 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.285 $Y=1.81
+ $X2=1.285 $Y2=1.47
r50 11 12 38.6168 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.285 $Y=1.81
+ $X2=1.285 $Y2=1.975
r51 10 22 38.6168 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.285 $Y=1.305
+ $X2=1.285 $Y2=1.47
r52 7 12 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.305 $Y=2.765
+ $X2=1.305 $Y2=1.975
r53 3 10 253.819 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=1.265 $Y=0.81
+ $X2=1.265 $Y2=1.305
.ends

.subckt PM_SKY130_FD_SC_LP__SDFXBP_2%A_332_94# 1 2 9 13 15 17 19 25 26
c59 26 0 1.59813e-19 $X=2.73 $Y=1.555
r60 25 28 53.334 $w=2.13e-07 $l=9.95e-07 $layer=LI1_cond $X=2.742 $Y=1.555
+ $X2=2.742 $Y2=2.55
r61 25 26 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.73
+ $Y=1.555 $X2=2.73 $Y2=1.555
r62 23 25 37.2534 $w=2.13e-07 $l=6.95e-07 $layer=LI1_cond $X=2.742 $Y=0.86
+ $X2=2.742 $Y2=1.555
r63 19 23 6.97049 $w=2.8e-07 $l=1.85957e-07 $layer=LI1_cond $X=2.635 $Y=0.72
+ $X2=2.742 $Y2=0.86
r64 19 21 7.20277 $w=2.78e-07 $l=1.75e-07 $layer=LI1_cond $X=2.635 $Y=0.72
+ $X2=2.46 $Y2=0.72
r65 18 26 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=2.73 $Y=1.54
+ $X2=2.73 $Y2=1.555
r66 16 17 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.81 $Y=1.465
+ $X2=1.735 $Y2=1.465
r67 15 18 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=2.565 $Y=1.465
+ $X2=2.73 $Y2=1.54
r68 15 16 387.138 $w=1.5e-07 $l=7.55e-07 $layer=POLY_cond $X=2.565 $Y=1.465
+ $X2=1.81 $Y2=1.465
r69 11 17 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.735 $Y=1.54
+ $X2=1.735 $Y2=1.465
r70 11 13 628.138 $w=1.5e-07 $l=1.225e-06 $layer=POLY_cond $X=1.735 $Y=1.54
+ $X2=1.735 $Y2=2.765
r71 7 17 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.735 $Y=1.39
+ $X2=1.735 $Y2=1.465
r72 7 9 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=1.735 $Y=1.39
+ $X2=1.735 $Y2=0.81
r73 2 28 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=2.64
+ $Y=2.405 $X2=2.765 $Y2=2.55
r74 1 21 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=2.32
+ $Y=0.6 $X2=2.46 $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_LP__SDFXBP_2%SCE 4 5 7 8 9 12 14 18 22 24 27 28 29 30 35
+ 36
r78 35 36 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.12
+ $Y=0.43 $X2=3.12 $Y2=0.43
r79 29 30 16.0907 $w=2.63e-07 $l=3.7e-07 $layer=LI1_cond $X=3.152 $Y=0.925
+ $X2=3.152 $Y2=1.295
r80 28 29 16.0907 $w=2.63e-07 $l=3.7e-07 $layer=LI1_cond $X=3.152 $Y=0.555
+ $X2=3.152 $Y2=0.925
r81 28 36 5.43605 $w=2.63e-07 $l=1.25e-07 $layer=LI1_cond $X=3.152 $Y=0.555
+ $X2=3.152 $Y2=0.43
r82 26 35 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=3.12 $Y=0.77
+ $X2=3.12 $Y2=0.43
r83 26 27 41.8716 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.12 $Y=0.77
+ $X2=3.12 $Y2=0.935
r84 25 35 29.7264 $w=3.3e-07 $l=1.7e-07 $layer=POLY_cond $X=3.12 $Y=0.26
+ $X2=3.12 $Y2=0.43
r85 20 22 56.4043 $w=1.5e-07 $l=1.1e-07 $layer=POLY_cond $X=0.835 $Y=2.26
+ $X2=0.945 $Y2=2.26
r86 18 27 917.851 $w=1.5e-07 $l=1.79e-06 $layer=POLY_cond $X=3.18 $Y=2.725
+ $X2=3.18 $Y2=0.935
r87 15 24 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.32 $Y=0.185
+ $X2=2.245 $Y2=0.185
r88 14 25 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=2.955 $Y=0.185
+ $X2=3.12 $Y2=0.26
r89 14 15 325.606 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.955 $Y=0.185
+ $X2=2.32 $Y2=0.185
r90 10 24 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.245 $Y=0.26
+ $X2=2.245 $Y2=0.185
r91 10 12 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=2.245 $Y=0.26
+ $X2=2.245 $Y2=0.81
r92 8 24 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.17 $Y=0.185
+ $X2=2.245 $Y2=0.185
r93 8 9 646.085 $w=1.5e-07 $l=1.26e-06 $layer=POLY_cond $X=2.17 $Y=0.185
+ $X2=0.91 $Y2=0.185
r94 5 22 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.945 $Y=2.335
+ $X2=0.945 $Y2=2.26
r95 5 7 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=0.945 $Y=2.335
+ $X2=0.945 $Y2=2.765
r96 2 20 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.835 $Y=2.185
+ $X2=0.835 $Y2=2.26
r97 2 4 705.053 $w=1.5e-07 $l=1.375e-06 $layer=POLY_cond $X=0.835 $Y=2.185
+ $X2=0.835 $Y2=0.81
r98 1 9 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.835 $Y=0.26
+ $X2=0.91 $Y2=0.185
r99 1 4 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=0.835 $Y=0.26
+ $X2=0.835 $Y2=0.81
.ends

.subckt PM_SKY130_FD_SC_LP__SDFXBP_2%A_778_399# 1 2 3 4 15 19 21 23 25 27 28 29
+ 32 33 34 37 45
c114 34 0 9.00427e-20 $X=6.795 $Y=2.45
c115 29 0 3.30294e-20 $X=6.625 $Y=1.76
c116 28 0 1.55846e-19 $X=4.98 $Y=2.035
c117 15 0 1.89499e-19 $X=4.89 $Y=2.335
r118 45 46 14.5084 $w=2.99e-07 $l=9e-08 $layer=POLY_cond $X=4.98 $Y=1.74
+ $X2=4.89 $Y2=1.74
r119 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.98
+ $Y=1.76 $X2=4.98 $Y2=1.76
r120 37 40 53.4113 $w=2.58e-07 $l=1.205e-06 $layer=LI1_cond $X=9.745 $Y=0.825
+ $X2=9.745 $Y2=2.03
r121 35 40 14.8488 $w=2.58e-07 $l=3.35e-07 $layer=LI1_cond $X=9.745 $Y=2.365
+ $X2=9.745 $Y2=2.03
r122 33 35 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=9.615 $Y=2.45
+ $X2=9.745 $Y2=2.365
r123 33 34 183.979 $w=1.68e-07 $l=2.82e-06 $layer=LI1_cond $X=9.615 $Y=2.45
+ $X2=6.795 $Y2=2.45
r124 32 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.71 $Y=2.365
+ $X2=6.795 $Y2=2.45
r125 31 32 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=6.71 $Y=1.845
+ $X2=6.71 $Y2=2.365
r126 30 44 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.145 $Y=1.76
+ $X2=4.98 $Y2=1.76
r127 29 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.625 $Y=1.76
+ $X2=6.71 $Y2=1.845
r128 29 30 96.5562 $w=1.68e-07 $l=1.48e-06 $layer=LI1_cond $X=6.625 $Y=1.76
+ $X2=5.145 $Y2=1.76
r129 27 44 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.98 $Y=1.845
+ $X2=4.98 $Y2=1.76
r130 27 28 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=4.98 $Y=1.845
+ $X2=4.98 $Y2=2.035
r131 26 42 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.2 $Y=2.12
+ $X2=4.035 $Y2=2.12
r132 25 28 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.815 $Y=2.12
+ $X2=4.98 $Y2=2.035
r133 25 26 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=4.815 $Y=2.12
+ $X2=4.2 $Y2=2.12
r134 21 42 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.035 $Y=2.035
+ $X2=4.035 $Y2=2.12
r135 21 23 44.8754 $w=3.28e-07 $l=1.285e-06 $layer=LI1_cond $X=4.035 $Y=2.035
+ $X2=4.035 $Y2=0.75
r136 17 45 39.495 $w=2.99e-07 $l=3.24577e-07 $layer=POLY_cond $X=5.225 $Y=1.555
+ $X2=4.98 $Y2=1.74
r137 17 19 384.574 $w=1.5e-07 $l=7.5e-07 $layer=POLY_cond $X=5.225 $Y=1.555
+ $X2=5.225 $Y2=0.805
r138 13 46 18.89 $w=1.5e-07 $l=1.85e-07 $layer=POLY_cond $X=4.89 $Y=1.925
+ $X2=4.89 $Y2=1.74
r139 13 15 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=4.89 $Y=1.925
+ $X2=4.89 $Y2=2.335
r140 4 40 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=9.635
+ $Y=1.895 $X2=9.78 $Y2=2.03
r141 3 42 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=3.89
+ $Y=1.995 $X2=4.035 $Y2=2.12
r142 2 37 182 $w=1.7e-07 $l=2.7037e-07 $layer=licon1_NDIFF $count=1 $X=9.625
+ $Y=0.61 $X2=9.75 $Y2=0.825
r143 1 23 91 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=2 $X=3.91
+ $Y=0.595 $X2=4.035 $Y2=0.75
.ends

.subckt PM_SKY130_FD_SC_LP__SDFXBP_2%A_733_21# 1 2 8 10 11 12 13 15 16 17 19 20
+ 22 23 26 27 28 30 33 37 39 40 43 48 49
c127 48 0 2.74945e-19 $X=6.66 $Y=0.35
c128 30 0 1.89499e-19 $X=6.115 $Y=2.11
c129 20 0 1.55846e-19 $X=4.365 $Y=3.075
r130 48 49 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.66
+ $Y=0.35 $X2=6.66 $Y2=0.35
r131 41 43 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=6.28 $Y=2.205
+ $X2=6.28 $Y2=2.65
r132 39 48 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.495 $Y=0.35
+ $X2=6.66 $Y2=0.35
r133 39 40 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=6.495 $Y=0.35
+ $X2=5.92 $Y2=0.35
r134 35 40 7.39867 $w=1.7e-07 $l=1.80566e-07 $layer=LI1_cond $X=5.777 $Y=0.435
+ $X2=5.92 $Y2=0.35
r135 35 37 14.7594 $w=2.83e-07 $l=3.65e-07 $layer=LI1_cond $X=5.777 $Y=0.435
+ $X2=5.777 $Y2=0.8
r136 33 54 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.565 $Y=2.11
+ $X2=5.565 $Y2=2.275
r137 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.565
+ $Y=2.11 $X2=5.565 $Y2=2.11
r138 30 41 7.47963 $w=1.9e-07 $l=2.07123e-07 $layer=LI1_cond $X=6.115 $Y=2.11
+ $X2=6.28 $Y2=2.205
r139 30 32 32.1053 $w=1.88e-07 $l=5.5e-07 $layer=LI1_cond $X=6.115 $Y=2.11
+ $X2=5.565 $Y2=2.11
r140 29 49 16.6118 $w=3.3e-07 $l=9.5e-08 $layer=POLY_cond $X=6.66 $Y=0.255
+ $X2=6.66 $Y2=0.35
r141 26 54 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=5.475 $Y=3.075
+ $X2=5.475 $Y2=2.275
r142 24 28 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.44 $Y=3.15
+ $X2=4.365 $Y2=3.15
r143 23 26 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.4 $Y=3.15
+ $X2=5.475 $Y2=3.075
r144 23 24 492.255 $w=1.5e-07 $l=9.6e-07 $layer=POLY_cond $X=5.4 $Y=3.15
+ $X2=4.44 $Y2=3.15
r145 20 28 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.365 $Y=3.075
+ $X2=4.365 $Y2=3.15
r146 20 22 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=4.365 $Y=3.075
+ $X2=4.365 $Y2=2.545
r147 17 19 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=4.25 $Y=1.345
+ $X2=4.25 $Y2=0.915
r148 15 28 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.29 $Y=3.15
+ $X2=4.365 $Y2=3.15
r149 15 16 243.564 $w=1.5e-07 $l=4.75e-07 $layer=POLY_cond $X=4.29 $Y=3.15
+ $X2=3.815 $Y2=3.15
r150 14 27 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.815 $Y=1.42
+ $X2=3.74 $Y2=1.42
r151 13 17 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.175 $Y=1.42
+ $X2=4.25 $Y2=1.345
r152 13 14 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=4.175 $Y=1.42
+ $X2=3.815 $Y2=1.42
r153 11 29 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=6.495 $Y=0.18
+ $X2=6.66 $Y2=0.255
r154 11 12 1374.21 $w=1.5e-07 $l=2.68e-06 $layer=POLY_cond $X=6.495 $Y=0.18
+ $X2=3.815 $Y2=0.18
r155 10 16 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.74 $Y=3.075
+ $X2=3.815 $Y2=3.15
r156 9 27 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.74 $Y=1.495
+ $X2=3.74 $Y2=1.42
r157 9 10 810.17 $w=1.5e-07 $l=1.58e-06 $layer=POLY_cond $X=3.74 $Y=1.495
+ $X2=3.74 $Y2=3.075
r158 8 27 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.74 $Y=1.345
+ $X2=3.74 $Y2=1.42
r159 7 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.74 $Y=0.255
+ $X2=3.815 $Y2=0.18
r160 7 8 558.915 $w=1.5e-07 $l=1.09e-06 $layer=POLY_cond $X=3.74 $Y=0.255
+ $X2=3.74 $Y2=1.345
r161 2 43 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=6.14
+ $Y=2.505 $X2=6.28 $Y2=2.65
r162 1 37 182 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_NDIFF $count=1 $X=5.66
+ $Y=0.595 $X2=5.8 $Y2=0.8
.ends

.subckt PM_SKY130_FD_SC_LP__SDFXBP_2%A_1102_93# 1 2 9 11 12 15 19 23 25 29 31 32
+ 34 35 36 40 41 42 44 48 51 57 59
c148 59 0 3.08584e-19 $X=7.23 $Y=0.18
c149 35 0 1.59193e-19 $X=6.065 $Y=1.59
c150 15 0 9.74678e-20 $X=6.065 $Y=2.715
r151 54 55 8.28399 $w=3.98e-07 $l=1.65e-07 $layer=LI1_cond $X=7.195 $Y=0.805
+ $X2=7.195 $Y2=0.97
r152 52 59 29.7264 $w=3.3e-07 $l=1.7e-07 $layer=POLY_cond $X=7.23 $Y=0.35
+ $X2=7.23 $Y2=0.18
r153 51 54 13.109 $w=3.98e-07 $l=4.55e-07 $layer=LI1_cond $X=7.195 $Y=0.35
+ $X2=7.195 $Y2=0.805
r154 51 52 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.23
+ $Y=0.35 $X2=7.23 $Y2=0.35
r155 46 54 1.86583 $w=3.3e-07 $l=2e-07 $layer=LI1_cond $X=7.395 $Y=0.805
+ $X2=7.195 $Y2=0.805
r156 46 48 8.20679 $w=3.28e-07 $l=2.35e-07 $layer=LI1_cond $X=7.395 $Y=0.805
+ $X2=7.63 $Y2=0.805
r157 42 44 7.90892 $w=2.53e-07 $l=1.75e-07 $layer=LI1_cond $X=7.175 $Y=2.067
+ $X2=7.35 $Y2=2.067
r158 41 57 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.09 $Y=1.65
+ $X2=6.925 $Y2=1.65
r159 40 55 41.899 $w=1.78e-07 $l=6.8e-07 $layer=LI1_cond $X=7.085 $Y=1.65
+ $X2=7.085 $Y2=0.97
r160 40 41 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.09
+ $Y=1.65 $X2=7.09 $Y2=1.65
r161 38 42 7.08339 $w=2.55e-07 $l=1.66009e-07 $layer=LI1_cond $X=7.085 $Y=1.94
+ $X2=7.175 $Y2=2.067
r162 38 40 17.8687 $w=1.78e-07 $l=2.9e-07 $layer=LI1_cond $X=7.085 $Y=1.94
+ $X2=7.085 $Y2=1.65
r163 33 34 1446 $w=1.5e-07 $l=2.82e-06 $layer=POLY_cond $X=11.96 $Y=0.255
+ $X2=11.96 $Y2=3.075
r164 31 34 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=11.885 $Y=3.15
+ $X2=11.96 $Y2=3.075
r165 31 32 669.16 $w=1.5e-07 $l=1.305e-06 $layer=POLY_cond $X=11.885 $Y=3.15
+ $X2=10.58 $Y2=3.15
r166 27 32 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=10.505 $Y=3.075
+ $X2=10.58 $Y2=3.15
r167 27 29 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=10.505 $Y=3.075
+ $X2=10.505 $Y2=2.525
r168 26 36 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=10.04 $Y=0.18
+ $X2=9.965 $Y2=0.18
r169 25 33 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=11.885 $Y=0.18
+ $X2=11.96 $Y2=0.255
r170 25 26 946.053 $w=1.5e-07 $l=1.845e-06 $layer=POLY_cond $X=11.885 $Y=0.18
+ $X2=10.04 $Y2=0.18
r171 21 36 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.965 $Y=0.255
+ $X2=9.965 $Y2=0.18
r172 21 23 289.713 $w=1.5e-07 $l=5.65e-07 $layer=POLY_cond $X=9.965 $Y=0.255
+ $X2=9.965 $Y2=0.82
r173 20 59 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.395 $Y=0.18
+ $X2=7.23 $Y2=0.18
r174 19 36 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.89 $Y=0.18
+ $X2=9.965 $Y2=0.18
r175 19 20 1279.35 $w=1.5e-07 $l=2.495e-06 $layer=POLY_cond $X=9.89 $Y=0.18
+ $X2=7.395 $Y2=0.18
r176 18 35 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.14 $Y=1.59
+ $X2=6.065 $Y2=1.59
r177 18 57 402.521 $w=1.5e-07 $l=7.85e-07 $layer=POLY_cond $X=6.14 $Y=1.59
+ $X2=6.925 $Y2=1.59
r178 13 35 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.065 $Y=1.665
+ $X2=6.065 $Y2=1.59
r179 13 15 538.404 $w=1.5e-07 $l=1.05e-06 $layer=POLY_cond $X=6.065 $Y=1.665
+ $X2=6.065 $Y2=2.715
r180 11 35 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.99 $Y=1.59
+ $X2=6.065 $Y2=1.59
r181 11 12 169.213 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=5.99 $Y=1.59
+ $X2=5.66 $Y2=1.59
r182 7 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.585 $Y=1.515
+ $X2=5.66 $Y2=1.59
r183 7 9 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=5.585 $Y=1.515
+ $X2=5.585 $Y2=0.805
r184 2 44 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=7.205
+ $Y=1.975 $X2=7.35 $Y2=2.11
r185 1 48 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=7.505
+ $Y=0.595 $X2=7.63 $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_LP__SDFXBP_2%A_1188_93# 1 2 7 9 10 11 12 14 15 16 21 23
+ 25 27 28 32 34 36 38 41 43 45 48 50 52 54 61 62 66
c151 32 0 1.73239e-19 $X=9.995 $Y=2.315
c152 10 0 3.30294e-20 $X=7.59 $Y=1.2
r153 70 71 67.0401 $w=3.5e-07 $l=2.9e-07 $layer=POLY_cond $X=8.88 $Y=1.445
+ $X2=8.88 $Y2=1.735
r154 62 70 35.4469 $w=3.5e-07 $l=2.15e-07 $layer=POLY_cond $X=8.88 $Y=1.23
+ $X2=8.88 $Y2=1.445
r155 61 62 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=8.89
+ $Y=1.23 $X2=8.89 $Y2=1.23
r156 59 61 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=8.885 $Y=1.565
+ $X2=8.885 $Y2=1.23
r157 58 61 9.07985 $w=3.28e-07 $l=2.6e-07 $layer=LI1_cond $X=8.885 $Y=0.97
+ $X2=8.885 $Y2=1.23
r158 54 58 6.81649 $w=3.3e-07 $l=2.33345e-07 $layer=LI1_cond $X=8.72 $Y=0.805
+ $X2=8.885 $Y2=0.97
r159 54 56 8.03218 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=8.72 $Y=0.805
+ $X2=8.49 $Y2=0.805
r160 50 59 26.3784 $w=1.85e-07 $l=4e-07 $layer=LI1_cond $X=8.485 $Y=1.667
+ $X2=8.885 $Y2=1.667
r161 50 52 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=8.485 $Y=1.77
+ $X2=8.485 $Y2=2.11
r162 48 67 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.755 $Y=1.65
+ $X2=7.755 $Y2=1.815
r163 48 66 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.755 $Y=1.65
+ $X2=7.755 $Y2=1.485
r164 47 48 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.755
+ $Y=1.65 $X2=7.755 $Y2=1.65
r165 45 50 9.96163 $w=2.05e-07 $l=1.65e-07 $layer=LI1_cond $X=8.32 $Y=1.667
+ $X2=8.485 $Y2=1.667
r166 45 47 30.5676 $w=2.03e-07 $l=5.65e-07 $layer=LI1_cond $X=8.32 $Y=1.667
+ $X2=7.755 $Y2=1.667
r167 40 41 92.2979 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=7.665 $Y=1.2
+ $X2=7.845 $Y2=1.2
r168 36 44 80.7822 $w=1.72e-07 $l=2.98672e-07 $layer=POLY_cond $X=10.41 $Y=1.16
+ $X2=10.382 $Y2=1.445
r169 36 38 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=10.41 $Y=1.16
+ $X2=10.41 $Y2=0.82
r170 35 43 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=10.07 $Y=1.445
+ $X2=9.995 $Y2=1.445
r171 34 44 6.07713 $w=1.5e-07 $l=1.02e-07 $layer=POLY_cond $X=10.28 $Y=1.445
+ $X2=10.382 $Y2=1.445
r172 34 35 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=10.28 $Y=1.445
+ $X2=10.07 $Y2=1.445
r173 30 43 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.995 $Y=1.52
+ $X2=9.995 $Y2=1.445
r174 30 32 407.649 $w=1.5e-07 $l=7.95e-07 $layer=POLY_cond $X=9.995 $Y=1.52
+ $X2=9.995 $Y2=2.315
r175 29 70 22.6286 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=9.055 $Y=1.445
+ $X2=8.88 $Y2=1.445
r176 28 43 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.92 $Y=1.445
+ $X2=9.995 $Y2=1.445
r177 28 29 443.543 $w=1.5e-07 $l=8.65e-07 $layer=POLY_cond $X=9.92 $Y=1.445
+ $X2=9.055 $Y2=1.445
r178 27 71 666.596 $w=1.5e-07 $l=1.3e-06 $layer=POLY_cond $X=8.78 $Y=3.035
+ $X2=8.78 $Y2=1.735
r179 23 41 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.845 $Y=1.125
+ $X2=7.845 $Y2=1.2
r180 23 25 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=7.845 $Y=1.125
+ $X2=7.845 $Y2=0.805
r181 21 67 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=7.68 $Y=2.295
+ $X2=7.68 $Y2=1.815
r182 17 40 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.665 $Y=1.275
+ $X2=7.665 $Y2=1.2
r183 17 66 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=7.665 $Y=1.275
+ $X2=7.665 $Y2=1.485
r184 15 27 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.705 $Y=3.11
+ $X2=8.78 $Y2=3.035
r185 15 16 1094.76 $w=1.5e-07 $l=2.135e-06 $layer=POLY_cond $X=8.705 $Y=3.11
+ $X2=6.57 $Y2=3.11
r186 12 16 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.495 $Y=3.035
+ $X2=6.57 $Y2=3.11
r187 12 14 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=6.495 $Y=3.035
+ $X2=6.495 $Y2=2.715
r188 10 40 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.59 $Y=1.2
+ $X2=7.665 $Y2=1.2
r189 10 11 769.149 $w=1.5e-07 $l=1.5e-06 $layer=POLY_cond $X=7.59 $Y=1.2
+ $X2=6.09 $Y2=1.2
r190 7 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.015 $Y=1.125
+ $X2=6.09 $Y2=1.2
r191 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=6.015 $Y=1.125
+ $X2=6.015 $Y2=0.805
r192 2 52 600 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_PDIFF $count=1 $X=8.345
+ $Y=1.975 $X2=8.485 $Y2=2.11
r193 1 56 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=8.35
+ $Y=0.595 $X2=8.49 $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_LP__SDFXBP_2%CLK 3 7 8 9 10 15 17
c44 10 0 3.3639e-20 $X=8.4 $Y=1.295
r45 15 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.325 $Y=1.295
+ $X2=8.325 $Y2=1.46
r46 15 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.325 $Y=1.295
+ $X2=8.325 $Y2=1.13
r47 10 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.325
+ $Y=1.295 $X2=8.325 $Y2=1.295
r48 9 10 18.3035 $w=2.53e-07 $l=4.05e-07 $layer=LI1_cond $X=7.92 $Y=1.267
+ $X2=8.325 $Y2=1.267
r49 8 9 21.693 $w=2.53e-07 $l=4.8e-07 $layer=LI1_cond $X=7.44 $Y=1.267 $X2=7.92
+ $Y2=1.267
r50 7 17 104.433 $w=1.5e-07 $l=3.25e-07 $layer=POLY_cond $X=8.275 $Y=0.805
+ $X2=8.275 $Y2=1.13
r51 3 18 428.16 $w=1.5e-07 $l=8.35e-07 $layer=POLY_cond $X=8.27 $Y=2.295
+ $X2=8.27 $Y2=1.46
.ends

.subckt PM_SKY130_FD_SC_LP__SDFXBP_2%A_2122_329# 1 2 9 13 17 21 25 29 31 32 35
+ 39 41 46 48 49 50 51 57 60 61 65 67 69 72 73
c154 67 0 1.73239e-19 $X=10.94 $Y=1.847
c155 60 0 1.68636e-19 $X=13.69 $Y=1.49
r156 83 84 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=13.475 $Y=1.49
+ $X2=13.495 $Y2=1.49
r157 80 81 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=12.95 $Y=1.49
+ $X2=12.97 $Y2=1.49
r158 79 80 71.6931 $w=3.3e-07 $l=4.1e-07 $layer=POLY_cond $X=12.54 $Y=1.49
+ $X2=12.95 $Y2=1.49
r159 77 79 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=12.52 $Y=1.49
+ $X2=12.54 $Y2=1.49
r160 69 71 14.3578 $w=4.18e-07 $l=4.55e-07 $layer=LI1_cond $X=11.73 $Y=0.755
+ $X2=11.73 $Y2=1.21
r161 65 76 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=10.775 $Y=1.81
+ $X2=10.775 $Y2=1.975
r162 65 75 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=10.775 $Y=1.81
+ $X2=10.775 $Y2=1.645
r163 64 67 8.46863 $w=2.53e-07 $l=1.65e-07 $layer=LI1_cond $X=10.775 $Y=1.847
+ $X2=10.94 $Y2=1.847
r164 64 65 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.775
+ $Y=1.81 $X2=10.775 $Y2=1.81
r165 61 84 34.0979 $w=3.3e-07 $l=1.95e-07 $layer=POLY_cond $X=13.69 $Y=1.49
+ $X2=13.495 $Y2=1.49
r166 60 61 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=13.69
+ $Y=1.49 $X2=13.69 $Y2=1.49
r167 58 73 4.23118 $w=2.15e-07 $l=1.00995e-07 $layer=LI1_cond $X=13.32 $Y=1.495
+ $X2=13.235 $Y2=1.53
r168 58 60 22.798 $w=1.78e-07 $l=3.7e-07 $layer=LI1_cond $X=13.32 $Y=1.495
+ $X2=13.69 $Y2=1.495
r169 56 73 2.20034 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=13.235 $Y=1.655
+ $X2=13.235 $Y2=1.53
r170 56 57 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=13.235 $Y=1.655
+ $X2=13.235 $Y2=2.375
r171 54 81 6.99445 $w=3.3e-07 $l=4e-08 $layer=POLY_cond $X=13.01 $Y=1.49
+ $X2=12.97 $Y2=1.49
r172 53 54 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=13.01
+ $Y=1.49 $X2=13.01 $Y2=1.49
r173 51 73 4.23118 $w=2.15e-07 $l=8.5e-08 $layer=LI1_cond $X=13.15 $Y=1.53
+ $X2=13.235 $Y2=1.53
r174 51 53 6.45368 $w=2.48e-07 $l=1.4e-07 $layer=LI1_cond $X=13.15 $Y=1.53
+ $X2=13.01 $Y2=1.53
r175 49 57 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=13.15 $Y=2.46
+ $X2=13.235 $Y2=2.375
r176 49 50 78.9412 $w=1.68e-07 $l=1.21e-06 $layer=LI1_cond $X=13.15 $Y=2.46
+ $X2=11.94 $Y2=2.46
r177 48 72 3.17288 $w=3.15e-07 $l=1.1811e-07 $layer=LI1_cond $X=11.815 $Y=1.795
+ $X2=11.75 $Y2=1.885
r178 48 71 26.9672 $w=2.48e-07 $l=5.85e-07 $layer=LI1_cond $X=11.815 $Y=1.795
+ $X2=11.815 $Y2=1.21
r179 44 50 8.19669 $w=1.7e-07 $l=2.28583e-07 $layer=LI1_cond $X=11.75 $Y=2.375
+ $X2=11.94 $Y2=2.46
r180 44 46 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=11.75 $Y=2.375
+ $X2=11.75 $Y2=2.04
r181 43 72 3.17288 $w=3.15e-07 $l=9e-08 $layer=LI1_cond $X=11.75 $Y=1.975
+ $X2=11.75 $Y2=1.885
r182 43 46 1.97128 $w=3.78e-07 $l=6.5e-08 $layer=LI1_cond $X=11.75 $Y=1.975
+ $X2=11.75 $Y2=2.04
r183 41 72 3.41642 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=11.56 $Y=1.885
+ $X2=11.75 $Y2=1.885
r184 41 67 38.202 $w=1.78e-07 $l=6.2e-07 $layer=LI1_cond $X=11.56 $Y=1.885
+ $X2=10.94 $Y2=1.885
r185 37 84 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=13.495 $Y=1.655
+ $X2=13.495 $Y2=1.49
r186 37 39 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=13.495 $Y=1.655
+ $X2=13.495 $Y2=2.155
r187 33 83 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=13.475 $Y=1.325
+ $X2=13.475 $Y2=1.49
r188 33 35 428.16 $w=1.5e-07 $l=8.35e-07 $layer=POLY_cond $X=13.475 $Y=1.325
+ $X2=13.475 $Y2=0.49
r189 32 54 6.12014 $w=3.3e-07 $l=3.5e-08 $layer=POLY_cond $X=13.045 $Y=1.49
+ $X2=13.01 $Y2=1.49
r190 31 83 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=13.4 $Y=1.49
+ $X2=13.475 $Y2=1.49
r191 31 32 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=13.4 $Y=1.49
+ $X2=13.045 $Y2=1.49
r192 27 81 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=12.97 $Y=1.655
+ $X2=12.97 $Y2=1.49
r193 27 29 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=12.97 $Y=1.655
+ $X2=12.97 $Y2=2.465
r194 23 80 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=12.95 $Y=1.325
+ $X2=12.95 $Y2=1.49
r195 23 25 320.479 $w=1.5e-07 $l=6.25e-07 $layer=POLY_cond $X=12.95 $Y=1.325
+ $X2=12.95 $Y2=0.7
r196 19 79 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=12.54 $Y=1.655
+ $X2=12.54 $Y2=1.49
r197 19 21 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=12.54 $Y=1.655
+ $X2=12.54 $Y2=2.465
r198 15 77 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=12.52 $Y=1.325
+ $X2=12.52 $Y2=1.49
r199 15 17 320.479 $w=1.5e-07 $l=6.25e-07 $layer=POLY_cond $X=12.52 $Y=1.325
+ $X2=12.52 $Y2=0.7
r200 13 76 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=10.865 $Y=2.525
+ $X2=10.865 $Y2=1.975
r201 9 75 423.032 $w=1.5e-07 $l=8.25e-07 $layer=POLY_cond $X=10.77 $Y=0.82
+ $X2=10.77 $Y2=1.645
r202 2 46 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=11.515
+ $Y=1.895 $X2=11.655 $Y2=2.04
r203 1 69 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=11.545
+ $Y=0.61 $X2=11.685 $Y2=0.755
.ends

.subckt PM_SKY130_FD_SC_LP__SDFXBP_2%A_2008_122# 1 2 9 13 16 20 26 28 29 30 33
r67 29 34 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=11.362 $Y=1.53
+ $X2=11.362 $Y2=1.695
r68 29 33 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=11.362 $Y=1.53
+ $X2=11.362 $Y2=1.365
r69 28 30 8.85254 $w=2.43e-07 $l=1.65e-07 $layer=LI1_cond $X=11.345 $Y=1.502
+ $X2=11.18 $Y2=1.502
r70 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.345
+ $Y=1.53 $X2=11.345 $Y2=1.53
r71 25 26 3.63293 $w=1.7e-07 $l=1.58e-07 $layer=LI1_cond $X=10.36 $Y=1.465
+ $X2=10.202 $Y2=1.465
r72 25 30 53.4973 $w=1.68e-07 $l=8.2e-07 $layer=LI1_cond $X=10.36 $Y=1.465
+ $X2=11.18 $Y2=1.465
r73 20 22 21.5854 $w=3.13e-07 $l=5.9e-07 $layer=LI1_cond $X=10.202 $Y=2.02
+ $X2=10.202 $Y2=2.61
r74 18 26 3.01263 $w=3.15e-07 $l=8.5e-08 $layer=LI1_cond $X=10.202 $Y=1.55
+ $X2=10.202 $Y2=1.465
r75 18 20 17.1952 $w=3.13e-07 $l=4.7e-07 $layer=LI1_cond $X=10.202 $Y=1.55
+ $X2=10.202 $Y2=2.02
r76 14 26 3.01263 $w=3.15e-07 $l=8.5e-08 $layer=LI1_cond $X=10.202 $Y=1.38
+ $X2=10.202 $Y2=1.465
r77 14 16 20.3049 $w=3.13e-07 $l=5.55e-07 $layer=LI1_cond $X=10.202 $Y=1.38
+ $X2=10.202 $Y2=0.825
r78 13 33 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=11.47 $Y=0.93
+ $X2=11.47 $Y2=1.365
r79 9 34 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=11.44 $Y=2.315
+ $X2=11.44 $Y2=1.695
r80 2 22 600 $w=1.7e-07 $l=7.81873e-07 $layer=licon1_PDIFF $count=1 $X=10.07
+ $Y=1.895 $X2=10.21 $Y2=2.61
r81 2 20 600 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=10.07
+ $Y=1.895 $X2=10.21 $Y2=2.02
r82 1 16 182 $w=1.7e-07 $l=2.82046e-07 $layer=licon1_NDIFF $count=1 $X=10.04
+ $Y=0.61 $X2=10.195 $Y2=0.825
.ends

.subckt PM_SKY130_FD_SC_LP__SDFXBP_2%A_2710_56# 1 2 7 9 12 14 16 19 23 27 29 30
+ 32 45
c65 45 0 1.13888e-19 $X=14.875 $Y=1.35
c66 12 0 5.47483e-20 $X=14.445 $Y=2.465
r67 44 45 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=14.445 $Y=1.35
+ $X2=14.875 $Y2=1.35
r68 33 44 27.1035 $w=3.3e-07 $l=1.55e-07 $layer=POLY_cond $X=14.29 $Y=1.35
+ $X2=14.445 $Y2=1.35
r69 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=14.29
+ $Y=1.35 $X2=14.29 $Y2=1.35
r70 30 32 13.3354 $w=3.48e-07 $l=4.05e-07 $layer=LI1_cond $X=14.2 $Y=1.755
+ $X2=14.2 $Y2=1.35
r71 29 32 4.11587 $w=3.48e-07 $l=1.25e-07 $layer=LI1_cond $X=14.2 $Y=1.225
+ $X2=14.2 $Y2=1.35
r72 25 29 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=13.705 $Y=1.14
+ $X2=14.2 $Y2=1.14
r73 25 27 21.7043 $w=2.98e-07 $l=5.65e-07 $layer=LI1_cond $X=13.705 $Y=1.055
+ $X2=13.705 $Y2=0.49
r74 21 30 31.9679 $w=1.68e-07 $l=4.9e-07 $layer=LI1_cond $X=13.71 $Y=1.84
+ $X2=14.2 $Y2=1.84
r75 21 23 1.92074 $w=3.28e-07 $l=5.5e-08 $layer=LI1_cond $X=13.71 $Y=1.925
+ $X2=13.71 $Y2=1.98
r76 17 45 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=14.875 $Y=1.515
+ $X2=14.875 $Y2=1.35
r77 17 19 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=14.875 $Y=1.515
+ $X2=14.875 $Y2=2.465
r78 14 45 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=14.875 $Y=1.185
+ $X2=14.875 $Y2=1.35
r79 14 16 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=14.875 $Y=1.185
+ $X2=14.875 $Y2=0.655
r80 10 44 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=14.445 $Y=1.515
+ $X2=14.445 $Y2=1.35
r81 10 12 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=14.445 $Y=1.515
+ $X2=14.445 $Y2=2.465
r82 7 44 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=14.445 $Y=1.185
+ $X2=14.445 $Y2=1.35
r83 7 9 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=14.445 $Y=1.185
+ $X2=14.445 $Y2=0.655
r84 2 23 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=13.57
+ $Y=1.835 $X2=13.71 $Y2=1.98
r85 1 27 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=13.55
+ $Y=0.28 $X2=13.69 $Y2=0.49
.ends

.subckt PM_SKY130_FD_SC_LP__SDFXBP_2%A_27_489# 1 2 9 11 12 13
r33 13 16 8.3814 $w=3.28e-07 $l=2.4e-07 $layer=LI1_cond $X=1.95 $Y=2.375
+ $X2=1.95 $Y2=2.615
r34 11 13 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.785 $Y=2.375
+ $X2=1.95 $Y2=2.375
r35 11 12 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=1.785 $Y=2.375
+ $X2=0.425 $Y2=2.375
r36 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.26 $Y=2.46
+ $X2=0.425 $Y2=2.375
r37 7 9 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=0.26 $Y=2.46 $X2=0.26
+ $Y2=2.59
r38 2 16 600 $w=1.7e-07 $l=2.29565e-07 $layer=licon1_PDIFF $count=1 $X=1.81
+ $Y=2.445 $X2=1.95 $Y2=2.615
r39 1 9 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.445 $X2=0.26 $Y2=2.59
.ends

.subckt PM_SKY130_FD_SC_LP__SDFXBP_2%VPWR 1 2 3 4 5 6 7 8 9 30 34 38 42 46 48 52
+ 56 58 62 66 68 73 74 75 77 89 93 101 109 114 120 123 126 129 132 135 138 142
r164 141 142 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=15.12 $Y=3.33
+ $X2=15.12 $Y2=3.33
r165 138 139 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=14.16 $Y=3.33
+ $X2=14.16 $Y2=3.33
r166 136 139 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=13.2 $Y=3.33
+ $X2=14.16 $Y2=3.33
r167 135 136 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.2 $Y=3.33
+ $X2=13.2 $Y2=3.33
r168 132 133 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=12.24 $Y=3.33
+ $X2=12.24 $Y2=3.33
r169 130 133 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=11.28 $Y=3.33
+ $X2=12.24 $Y2=3.33
r170 129 130 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.28 $Y=3.33
+ $X2=11.28 $Y2=3.33
r171 126 127 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r172 123 124 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r173 120 121 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r174 118 142 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=14.64 $Y=3.33
+ $X2=15.12 $Y2=3.33
r175 118 139 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=14.64 $Y=3.33
+ $X2=14.16 $Y2=3.33
r176 117 118 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.64 $Y=3.33
+ $X2=14.64 $Y2=3.33
r177 115 138 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=14.335 $Y=3.33
+ $X2=14.23 $Y2=3.33
r178 115 117 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=14.335 $Y=3.33
+ $X2=14.64 $Y2=3.33
r179 114 141 4.20444 $w=1.7e-07 $l=1.87e-07 $layer=LI1_cond $X=14.985 $Y=3.33
+ $X2=15.172 $Y2=3.33
r180 114 117 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=14.985 $Y=3.33
+ $X2=14.64 $Y2=3.33
r181 113 136 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.72 $Y=3.33
+ $X2=13.2 $Y2=3.33
r182 113 133 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.72 $Y=3.33
+ $X2=12.24 $Y2=3.33
r183 112 113 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.72 $Y=3.33
+ $X2=12.72 $Y2=3.33
r184 110 132 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.49 $Y=3.33
+ $X2=12.325 $Y2=3.33
r185 110 112 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=12.49 $Y=3.33
+ $X2=12.72 $Y2=3.33
r186 109 135 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.02 $Y=3.33
+ $X2=13.185 $Y2=3.33
r187 109 112 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=13.02 $Y=3.33
+ $X2=12.72 $Y2=3.33
r188 108 130 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.8 $Y=3.33
+ $X2=11.28 $Y2=3.33
r189 107 108 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=10.8 $Y=3.33
+ $X2=10.8 $Y2=3.33
r190 105 108 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=10.8 $Y2=3.33
r191 105 127 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=7.92 $Y2=3.33
r192 104 107 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=8.4 $Y=3.33
+ $X2=10.8 $Y2=3.33
r193 104 105 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r194 102 126 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.14 $Y=3.33
+ $X2=7.975 $Y2=3.33
r195 102 104 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=8.14 $Y=3.33
+ $X2=8.4 $Y2=3.33
r196 101 129 10.9443 $w=1.7e-07 $l=2.37e-07 $layer=LI1_cond $X=10.915 $Y=3.33
+ $X2=11.152 $Y2=3.33
r197 101 107 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=10.915 $Y=3.33
+ $X2=10.8 $Y2=3.33
r198 99 100 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r199 97 100 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=7.44 $Y2=3.33
r200 97 124 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=4.56 $Y2=3.33
r201 96 99 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=5.04 $Y=3.33
+ $X2=7.44 $Y2=3.33
r202 96 97 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r203 94 123 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.745 $Y=3.33
+ $X2=4.58 $Y2=3.33
r204 94 96 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=4.745 $Y=3.33
+ $X2=5.04 $Y2=3.33
r205 93 126 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.81 $Y=3.33
+ $X2=7.975 $Y2=3.33
r206 93 99 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=7.81 $Y=3.33
+ $X2=7.44 $Y2=3.33
r207 92 124 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r208 91 92 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r209 89 123 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.415 $Y=3.33
+ $X2=4.58 $Y2=3.33
r210 89 91 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=4.415 $Y=3.33
+ $X2=4.08 $Y2=3.33
r211 88 92 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=4.08 $Y2=3.33
r212 87 88 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r213 85 88 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=3.12 $Y2=3.33
r214 85 121 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r215 84 87 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=3.12 $Y2=3.33
r216 84 85 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r217 82 120 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=0.875 $Y=3.33
+ $X2=0.735 $Y2=3.33
r218 82 84 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.875 $Y=3.33
+ $X2=1.2 $Y2=3.33
r219 80 121 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r220 79 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r221 77 120 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=0.595 $Y=3.33
+ $X2=0.735 $Y2=3.33
r222 77 79 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=0.595 $Y=3.33
+ $X2=0.24 $Y2=3.33
r223 75 127 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=7.68 $Y=3.33
+ $X2=7.92 $Y2=3.33
r224 75 100 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=7.68 $Y=3.33
+ $X2=7.44 $Y2=3.33
r225 73 87 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=3.36 $Y=3.33
+ $X2=3.12 $Y2=3.33
r226 73 74 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.36 $Y=3.33
+ $X2=3.485 $Y2=3.33
r227 72 91 30.6631 $w=1.68e-07 $l=4.7e-07 $layer=LI1_cond $X=3.61 $Y=3.33
+ $X2=4.08 $Y2=3.33
r228 72 74 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.61 $Y=3.33
+ $X2=3.485 $Y2=3.33
r229 68 71 41.4026 $w=2.68e-07 $l=9.7e-07 $layer=LI1_cond $X=15.12 $Y=1.98
+ $X2=15.12 $Y2=2.95
r230 66 141 3.08026 $w=2.7e-07 $l=1.07912e-07 $layer=LI1_cond $X=15.12 $Y=3.245
+ $X2=15.172 $Y2=3.33
r231 66 71 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=15.12 $Y=3.245
+ $X2=15.12 $Y2=2.95
r232 62 65 35.9134 $w=2.08e-07 $l=6.8e-07 $layer=LI1_cond $X=14.23 $Y=2.27
+ $X2=14.23 $Y2=2.95
r233 60 138 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=14.23 $Y=3.245
+ $X2=14.23 $Y2=3.33
r234 60 65 15.5801 $w=2.08e-07 $l=2.95e-07 $layer=LI1_cond $X=14.23 $Y=3.245
+ $X2=14.23 $Y2=2.95
r235 59 135 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.35 $Y=3.33
+ $X2=13.185 $Y2=3.33
r236 58 138 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=14.125 $Y=3.33
+ $X2=14.23 $Y2=3.33
r237 58 59 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=14.125 $Y=3.33
+ $X2=13.35 $Y2=3.33
r238 54 135 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=13.185 $Y=3.245
+ $X2=13.185 $Y2=3.33
r239 54 56 14.8421 $w=3.28e-07 $l=4.25e-07 $layer=LI1_cond $X=13.185 $Y=3.245
+ $X2=13.185 $Y2=2.82
r240 50 132 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=12.325 $Y=3.245
+ $X2=12.325 $Y2=3.33
r241 50 52 14.8421 $w=3.28e-07 $l=4.25e-07 $layer=LI1_cond $X=12.325 $Y=3.245
+ $X2=12.325 $Y2=2.82
r242 49 129 10.9443 $w=1.7e-07 $l=2.38e-07 $layer=LI1_cond $X=11.39 $Y=3.33
+ $X2=11.152 $Y2=3.33
r243 48 132 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.16 $Y=3.33
+ $X2=12.325 $Y2=3.33
r244 48 49 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=12.16 $Y=3.33
+ $X2=11.39 $Y2=3.33
r245 44 129 1.94084 $w=4.75e-07 $l=8.5e-08 $layer=LI1_cond $X=11.152 $Y=3.245
+ $X2=11.152 $Y2=3.33
r246 44 46 25.5583 $w=4.73e-07 $l=1.015e-06 $layer=LI1_cond $X=11.152 $Y=3.245
+ $X2=11.152 $Y2=2.23
r247 40 126 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.975 $Y=3.245
+ $X2=7.975 $Y2=3.33
r248 40 42 15.8897 $w=3.28e-07 $l=4.55e-07 $layer=LI1_cond $X=7.975 $Y=3.245
+ $X2=7.975 $Y2=2.79
r249 36 123 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.58 $Y=3.245
+ $X2=4.58 $Y2=3.33
r250 36 38 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=4.58 $Y=3.245
+ $X2=4.58 $Y2=2.8
r251 32 74 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.485 $Y=3.245
+ $X2=3.485 $Y2=3.33
r252 32 34 16.8257 $w=2.48e-07 $l=3.65e-07 $layer=LI1_cond $X=3.485 $Y=3.245
+ $X2=3.485 $Y2=2.88
r253 28 120 0.375625 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=0.735 $Y=3.245
+ $X2=0.735 $Y2=3.33
r254 28 30 18.5214 $w=2.78e-07 $l=4.5e-07 $layer=LI1_cond $X=0.735 $Y=3.245
+ $X2=0.735 $Y2=2.795
r255 9 71 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=14.95
+ $Y=1.835 $X2=15.09 $Y2=2.95
r256 9 68 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=14.95
+ $Y=1.835 $X2=15.09 $Y2=1.98
r257 8 65 400 $w=1.7e-07 $l=1.17584e-06 $layer=licon1_PDIFF $count=1 $X=14.105
+ $Y=1.835 $X2=14.23 $Y2=2.95
r258 8 62 400 $w=1.7e-07 $l=4.93559e-07 $layer=licon1_PDIFF $count=1 $X=14.105
+ $Y=1.835 $X2=14.23 $Y2=2.27
r259 7 56 600 $w=1.7e-07 $l=1.05268e-06 $layer=licon1_PDIFF $count=1 $X=13.045
+ $Y=1.835 $X2=13.185 $Y2=2.82
r260 6 52 600 $w=1.7e-07 $l=1.04563e-06 $layer=licon1_PDIFF $count=1 $X=12.2
+ $Y=1.835 $X2=12.325 $Y2=2.82
r261 5 46 300 $w=1.7e-07 $l=3.24731e-07 $layer=licon1_PDIFF $count=2 $X=10.94
+ $Y=2.315 $X2=11.225 $Y2=2.23
r262 4 42 600 $w=1.7e-07 $l=9.18436e-07 $layer=licon1_PDIFF $count=1 $X=7.755
+ $Y=1.975 $X2=7.975 $Y2=2.79
r263 3 38 600 $w=1.7e-07 $l=7.41704e-07 $layer=licon1_PDIFF $count=1 $X=4.44
+ $Y=2.125 $X2=4.58 $Y2=2.8
r264 2 34 600 $w=1.7e-07 $l=5.62028e-07 $layer=licon1_PDIFF $count=1 $X=3.255
+ $Y=2.405 $X2=3.445 $Y2=2.88
r265 1 30 600 $w=1.7e-07 $l=4.22493e-07 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=2.445 $X2=0.71 $Y2=2.795
.ends

.subckt PM_SKY130_FD_SC_LP__SDFXBP_2%A_182_120# 1 2 3 4 13 17 19 20 22 23 26 28
+ 29 30 31 34 35 36 39 42 44 48 49
c164 48 0 1.59813e-19 $X=3.69 $Y=2.29
r165 49 52 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=5.77 $Y=2.46
+ $X2=5.77 $Y2=2.65
r166 47 48 7.70264 $w=5.08e-07 $l=8.5e-08 $layer=LI1_cond $X=3.605 $Y=2.29
+ $X2=3.69 $Y2=2.29
r167 45 47 11.7263 $w=5.08e-07 $l=5e-07 $layer=LI1_cond $X=3.105 $Y=2.29
+ $X2=3.605 $Y2=2.29
r168 42 43 12.688 $w=3e-07 $l=3.12e-07 $layer=LI1_cond $X=1.05 $Y=0.81 $X2=1.05
+ $Y2=1.122
r169 37 39 25.7461 $w=2.33e-07 $l=5.25e-07 $layer=LI1_cond $X=6.207 $Y=1.335
+ $X2=6.207 $Y2=0.81
r170 35 37 7.04737 $w=1.7e-07 $l=1.53734e-07 $layer=LI1_cond $X=6.09 $Y=1.42
+ $X2=6.207 $Y2=1.335
r171 35 36 101.123 $w=1.68e-07 $l=1.55e-06 $layer=LI1_cond $X=6.09 $Y=1.42
+ $X2=4.54 $Y2=1.42
r172 34 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.455 $Y=1.335
+ $X2=4.54 $Y2=1.42
r173 33 34 56.7594 $w=1.68e-07 $l=8.7e-07 $layer=LI1_cond $X=4.455 $Y=0.465
+ $X2=4.455 $Y2=1.335
r174 31 49 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.605 $Y=2.46
+ $X2=5.77 $Y2=2.46
r175 31 48 124.936 $w=1.68e-07 $l=1.915e-06 $layer=LI1_cond $X=5.605 $Y=2.46
+ $X2=3.69 $Y2=2.46
r176 29 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.37 $Y=0.38
+ $X2=4.455 $Y2=0.465
r177 29 30 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=4.37 $Y=0.38
+ $X2=3.69 $Y2=0.38
r178 28 47 7.28118 $w=1.7e-07 $l=2.55e-07 $layer=LI1_cond $X=3.605 $Y=2.035
+ $X2=3.605 $Y2=2.29
r179 27 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.605 $Y=0.465
+ $X2=3.69 $Y2=0.38
r180 27 28 102.428 $w=1.68e-07 $l=1.57e-06 $layer=LI1_cond $X=3.605 $Y=0.465
+ $X2=3.605 $Y2=2.035
r181 25 45 7.28118 $w=1.7e-07 $l=2.55e-07 $layer=LI1_cond $X=3.105 $Y=2.545
+ $X2=3.105 $Y2=2.29
r182 25 26 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=3.105 $Y=2.545
+ $X2=3.105 $Y2=2.905
r183 24 44 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.465 $Y=2.99
+ $X2=2.38 $Y2=2.99
r184 23 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.02 $Y=2.99
+ $X2=3.105 $Y2=2.905
r185 23 24 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=3.02 $Y=2.99
+ $X2=2.465 $Y2=2.99
r186 22 44 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.38 $Y=2.905
+ $X2=2.38 $Y2=2.99
r187 21 22 110.257 $w=1.68e-07 $l=1.69e-06 $layer=LI1_cond $X=2.38 $Y=1.215
+ $X2=2.38 $Y2=2.905
r188 19 44 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.295 $Y=2.99
+ $X2=2.38 $Y2=2.99
r189 19 20 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=2.295 $Y=2.99
+ $X2=1.615 $Y2=2.99
r190 15 20 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=1.485 $Y=2.905
+ $X2=1.615 $Y2=2.99
r191 15 17 4.87572 $w=2.58e-07 $l=1.1e-07 $layer=LI1_cond $X=1.485 $Y=2.905
+ $X2=1.485 $Y2=2.795
r192 14 43 3.58581 $w=1.85e-07 $l=1.65e-07 $layer=LI1_cond $X=1.215 $Y=1.122
+ $X2=1.05 $Y2=1.122
r193 13 21 6.83233 $w=1.85e-07 $l=1.28662e-07 $layer=LI1_cond $X=2.295 $Y=1.122
+ $X2=2.38 $Y2=1.215
r194 13 14 64.7469 $w=1.83e-07 $l=1.08e-06 $layer=LI1_cond $X=2.295 $Y=1.122
+ $X2=1.215 $Y2=1.122
r195 4 52 600 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=5.625
+ $Y=2.505 $X2=5.77 $Y2=2.65
r196 3 17 600 $w=1.7e-07 $l=4.14126e-07 $layer=licon1_PDIFF $count=1 $X=1.38
+ $Y=2.445 $X2=1.52 $Y2=2.795
r197 2 39 182 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_NDIFF $count=1 $X=6.09
+ $Y=0.595 $X2=6.23 $Y2=0.81
r198 1 42 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.91
+ $Y=0.6 $X2=1.05 $Y2=0.81
.ends

.subckt PM_SKY130_FD_SC_LP__SDFXBP_2%A_993_425# 1 2 7 10 15
c35 15 0 7.42513e-21 $X=6.79 $Y=2.79
r36 15 17 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=6.79 $Y=2.79 $X2=6.79
+ $Y2=2.99
r37 10 12 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=5.2 $Y=2.8 $X2=5.2
+ $Y2=2.99
r38 8 12 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.365 $Y=2.99 $X2=5.2
+ $Y2=2.99
r39 7 17 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.625 $Y=2.99
+ $X2=6.79 $Y2=2.99
r40 7 8 82.2032 $w=1.68e-07 $l=1.26e-06 $layer=LI1_cond $X=6.625 $Y=2.99
+ $X2=5.365 $Y2=2.99
r41 2 15 600 $w=1.7e-07 $l=3.79374e-07 $layer=licon1_PDIFF $count=1 $X=6.57
+ $Y=2.505 $X2=6.79 $Y2=2.79
r42 1 10 600 $w=1.7e-07 $l=7.83741e-07 $layer=licon1_PDIFF $count=1 $X=4.965
+ $Y=2.125 $X2=5.2 $Y2=2.8
.ends

.subckt PM_SKY130_FD_SC_LP__SDFXBP_2%Q 1 2 7 9 11 15 18 21 23
r44 21 23 3.84148 $w=2.23e-07 $l=7.5e-08 $layer=LI1_cond $X=12.222 $Y=1.22
+ $X2=12.222 $Y2=1.295
r45 18 21 3.00067 $w=2.25e-07 $l=8.5e-08 $layer=LI1_cond $X=12.222 $Y=1.135
+ $X2=12.222 $Y2=1.22
r46 18 23 0.256098 $w=2.23e-07 $l=5e-09 $layer=LI1_cond $X=12.222 $Y=1.3
+ $X2=12.222 $Y2=1.295
r47 17 18 29.4513 $w=2.23e-07 $l=5.75e-07 $layer=LI1_cond $X=12.222 $Y=1.875
+ $X2=12.222 $Y2=1.3
r48 13 15 31.3164 $w=2.28e-07 $l=6.25e-07 $layer=LI1_cond $X=12.755 $Y=1.05
+ $X2=12.755 $Y2=0.425
r49 9 17 7.1387 $w=3.3e-07 $l=2.14173e-07 $layer=LI1_cond $X=12.335 $Y=2.04
+ $X2=12.222 $Y2=1.875
r50 9 11 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=12.335 $Y=2.04
+ $X2=12.755 $Y2=2.04
r51 8 18 3.98913 $w=1.7e-07 $l=1.13e-07 $layer=LI1_cond $X=12.335 $Y=1.135
+ $X2=12.222 $Y2=1.135
r52 7 13 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=12.64 $Y=1.135
+ $X2=12.755 $Y2=1.05
r53 7 8 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=12.64 $Y=1.135
+ $X2=12.335 $Y2=1.135
r54 2 11 600 $w=1.7e-07 $l=3.07124e-07 $layer=licon1_PDIFF $count=1 $X=12.615
+ $Y=1.835 $X2=12.755 $Y2=2.08
r55 1 15 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=12.595
+ $Y=0.28 $X2=12.735 $Y2=0.425
.ends

.subckt PM_SKY130_FD_SC_LP__SDFXBP_2%Q_N 1 2 7 8 9 10 11 12 13 22
r18 13 40 5.98384 $w=2.58e-07 $l=1.35e-07 $layer=LI1_cond $X=14.685 $Y=2.775
+ $X2=14.685 $Y2=2.91
r19 12 13 16.4002 $w=2.58e-07 $l=3.7e-07 $layer=LI1_cond $X=14.685 $Y=2.405
+ $X2=14.685 $Y2=2.775
r20 11 12 17.2866 $w=2.58e-07 $l=3.9e-07 $layer=LI1_cond $X=14.685 $Y=2.015
+ $X2=14.685 $Y2=2.405
r21 10 11 15.5137 $w=2.58e-07 $l=3.5e-07 $layer=LI1_cond $X=14.685 $Y=1.665
+ $X2=14.685 $Y2=2.015
r22 9 10 16.4002 $w=2.58e-07 $l=3.7e-07 $layer=LI1_cond $X=14.685 $Y=1.295
+ $X2=14.685 $Y2=1.665
r23 8 9 16.4002 $w=2.58e-07 $l=3.7e-07 $layer=LI1_cond $X=14.685 $Y=0.925
+ $X2=14.685 $Y2=1.295
r24 7 8 16.4002 $w=2.58e-07 $l=3.7e-07 $layer=LI1_cond $X=14.685 $Y=0.555
+ $X2=14.685 $Y2=0.925
r25 7 22 5.98384 $w=2.58e-07 $l=1.35e-07 $layer=LI1_cond $X=14.685 $Y=0.555
+ $X2=14.685 $Y2=0.42
r26 2 40 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=14.52
+ $Y=1.835 $X2=14.66 $Y2=2.91
r27 2 11 400 $w=1.7e-07 $l=2.4e-07 $layer=licon1_PDIFF $count=1 $X=14.52
+ $Y=1.835 $X2=14.66 $Y2=2.015
r28 1 22 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=14.52
+ $Y=0.235 $X2=14.66 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__SDFXBP_2%VGND 1 2 3 4 5 6 7 8 9 28 30 34 38 42 46 50
+ 54 60 62 64 67 68 70 71 73 74 76 77 78 105 109 114 119 128 131 134 138
r163 137 138 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=15.12 $Y=0
+ $X2=15.12 $Y2=0
r164 134 135 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.16 $Y=0
+ $X2=14.16 $Y2=0
r165 131 132 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.2 $Y=0
+ $X2=13.2 $Y2=0
r166 128 129 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.24 $Y=0
+ $X2=12.24 $Y2=0
r167 125 126 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0
+ $X2=0.24 $Y2=0
r168 123 138 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=14.64 $Y=0
+ $X2=15.12 $Y2=0
r169 123 135 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=14.64 $Y=0
+ $X2=14.16 $Y2=0
r170 122 123 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.64 $Y=0
+ $X2=14.64 $Y2=0
r171 120 134 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=14.375 $Y=0
+ $X2=14.21 $Y2=0
r172 120 122 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=14.375 $Y=0
+ $X2=14.64 $Y2=0
r173 119 137 4.20444 $w=1.7e-07 $l=1.87e-07 $layer=LI1_cond $X=14.985 $Y=0
+ $X2=15.172 $Y2=0
r174 119 122 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=14.985 $Y=0
+ $X2=14.64 $Y2=0
r175 118 135 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.68 $Y=0
+ $X2=14.16 $Y2=0
r176 118 132 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.68 $Y=0
+ $X2=13.2 $Y2=0
r177 117 118 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.68 $Y=0
+ $X2=13.68 $Y2=0
r178 115 131 8.88104 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=13.385 $Y=0
+ $X2=13.212 $Y2=0
r179 115 117 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=13.385 $Y=0
+ $X2=13.68 $Y2=0
r180 114 134 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=14.045 $Y=0
+ $X2=14.21 $Y2=0
r181 114 117 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=14.045 $Y=0
+ $X2=13.68 $Y2=0
r182 113 132 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.72 $Y=0
+ $X2=13.2 $Y2=0
r183 113 129 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.72 $Y=0
+ $X2=12.24 $Y2=0
r184 112 113 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.72 $Y=0
+ $X2=12.72 $Y2=0
r185 110 128 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.47 $Y=0
+ $X2=12.305 $Y2=0
r186 110 112 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=12.47 $Y=0
+ $X2=12.72 $Y2=0
r187 109 131 8.88104 $w=1.7e-07 $l=1.72e-07 $layer=LI1_cond $X=13.04 $Y=0
+ $X2=13.212 $Y2=0
r188 109 112 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=13.04 $Y=0
+ $X2=12.72 $Y2=0
r189 108 129 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.76 $Y=0
+ $X2=12.24 $Y2=0
r190 107 108 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.76 $Y=0
+ $X2=11.76 $Y2=0
r191 105 128 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.14 $Y=0
+ $X2=12.305 $Y2=0
r192 105 107 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=12.14 $Y=0
+ $X2=11.76 $Y2=0
r193 104 108 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=10.8 $Y=0
+ $X2=11.76 $Y2=0
r194 103 104 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=10.8 $Y=0
+ $X2=10.8 $Y2=0
r195 101 104 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=8.4 $Y=0
+ $X2=10.8 $Y2=0
r196 100 103 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=8.4 $Y=0 $X2=10.8
+ $Y2=0
r197 100 101 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r198 98 101 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=8.4
+ $Y2=0
r199 97 98 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=7.92 $Y=0
+ $X2=7.92 $Y2=0
r200 94 97 187.893 $w=1.68e-07 $l=2.88e-06 $layer=LI1_cond $X=5.04 $Y=0 $X2=7.92
+ $Y2=0
r201 94 95 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=5.04 $Y=0
+ $X2=5.04 $Y2=0
r202 92 95 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.04
+ $Y2=0
r203 91 92 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r204 89 92 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=2.16 $Y=0 $X2=4.56
+ $Y2=0
r205 88 91 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=2.16 $Y=0 $X2=4.56
+ $Y2=0
r206 88 89 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r207 86 89 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r208 85 86 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r209 83 86 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r210 83 126 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0
+ $X2=0.24 $Y2=0
r211 82 85 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r212 82 83 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r213 80 125 4.78091 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=0
+ $X2=0.212 $Y2=0
r214 80 82 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.425 $Y=0 $X2=0.72
+ $Y2=0
r215 78 98 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=7.68 $Y=0
+ $X2=7.92 $Y2=0
r216 78 95 0.73586 $w=4.9e-07 $l=2.64e-06 $layer=MET1_cond $X=7.68 $Y=0 $X2=5.04
+ $Y2=0
r217 76 103 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=11.01 $Y=0
+ $X2=10.8 $Y2=0
r218 76 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.01 $Y=0
+ $X2=11.175 $Y2=0
r219 75 107 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=11.34 $Y=0
+ $X2=11.76 $Y2=0
r220 75 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.34 $Y=0
+ $X2=11.175 $Y2=0
r221 73 97 0.652406 $w=1.68e-07 $l=1e-08 $layer=LI1_cond $X=7.93 $Y=0 $X2=7.92
+ $Y2=0
r222 73 74 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.93 $Y=0 $X2=8.055
+ $Y2=0
r223 72 100 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=8.18 $Y=0 $X2=8.4
+ $Y2=0
r224 72 74 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.18 $Y=0 $X2=8.055
+ $Y2=0
r225 71 94 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.875 $Y=0 $X2=5.04
+ $Y2=0
r226 70 91 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=4.71 $Y=0 $X2=4.56
+ $Y2=0
r227 70 71 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.71 $Y=0 $X2=4.875
+ $Y2=0
r228 67 85 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=1.785 $Y=0
+ $X2=1.68 $Y2=0
r229 67 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.785 $Y=0 $X2=1.95
+ $Y2=0
r230 66 88 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=2.115 $Y=0 $X2=2.16
+ $Y2=0
r231 66 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.115 $Y=0 $X2=1.95
+ $Y2=0
r232 62 137 3.08026 $w=2.7e-07 $l=1.07912e-07 $layer=LI1_cond $X=15.12 $Y=0.085
+ $X2=15.172 $Y2=0
r233 62 64 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=15.12 $Y=0.085
+ $X2=15.12 $Y2=0.38
r234 58 134 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=14.21 $Y=0.085
+ $X2=14.21 $Y2=0
r235 58 60 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=14.21 $Y=0.085
+ $X2=14.21 $Y2=0.38
r236 54 56 18.3723 $w=3.43e-07 $l=5.5e-07 $layer=LI1_cond $X=13.212 $Y=0.425
+ $X2=13.212 $Y2=0.975
r237 52 131 1.03204 $w=3.45e-07 $l=8.5e-08 $layer=LI1_cond $X=13.212 $Y=0.085
+ $X2=13.212 $Y2=0
r238 52 54 11.3574 $w=3.43e-07 $l=3.4e-07 $layer=LI1_cond $X=13.212 $Y=0.085
+ $X2=13.212 $Y2=0.425
r239 48 128 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=12.305 $Y=0.085
+ $X2=12.305 $Y2=0
r240 48 50 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=12.305 $Y=0.085
+ $X2=12.305 $Y2=0.425
r241 44 77 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=11.175 $Y=0.085
+ $X2=11.175 $Y2=0
r242 44 46 23.3981 $w=3.28e-07 $l=6.7e-07 $layer=LI1_cond $X=11.175 $Y=0.085
+ $X2=11.175 $Y2=0.755
r243 40 74 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=8.055 $Y=0.085
+ $X2=8.055 $Y2=0
r244 40 42 33.1904 $w=2.48e-07 $l=7.2e-07 $layer=LI1_cond $X=8.055 $Y=0.085
+ $X2=8.055 $Y2=0.805
r245 36 71 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.875 $Y=0.085
+ $X2=4.875 $Y2=0
r246 36 38 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=4.875 $Y=0.085
+ $X2=4.875 $Y2=0.72
r247 32 68 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.95 $Y=0.085
+ $X2=1.95 $Y2=0
r248 32 34 23.2235 $w=3.28e-07 $l=6.65e-07 $layer=LI1_cond $X=1.95 $Y=0.085
+ $X2=1.95 $Y2=0.75
r249 28 125 2.98526 $w=3.3e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.212 $Y2=0
r250 28 30 25.3188 $w=3.28e-07 $l=7.25e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.26 $Y2=0.81
r251 9 64 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=14.95
+ $Y=0.235 $X2=15.09 $Y2=0.38
r252 8 60 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=14.085
+ $Y=0.235 $X2=14.21 $Y2=0.38
r253 7 56 182 $w=1.7e-07 $l=7.61791e-07 $layer=licon1_NDIFF $count=1 $X=13.025
+ $Y=0.28 $X2=13.165 $Y2=0.975
r254 7 54 182 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_NDIFF $count=1 $X=13.025
+ $Y=0.28 $X2=13.26 $Y2=0.425
r255 6 50 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=12.18
+ $Y=0.28 $X2=12.305 $Y2=0.425
r256 5 46 91 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=2 $X=10.845
+ $Y=0.61 $X2=11.12 $Y2=0.755
r257 4 42 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=7.92
+ $Y=0.595 $X2=8.06 $Y2=0.805
r258 3 38 91 $w=1.7e-07 $l=6.09303e-07 $layer=licon1_NDIFF $count=2 $X=4.325
+ $Y=0.595 $X2=4.875 $Y2=0.72
r259 2 34 182 $w=1.7e-07 $l=2.08567e-07 $layer=licon1_NDIFF $count=1 $X=1.81
+ $Y=0.6 $X2=1.95 $Y2=0.75
r260 1 30 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.6 $X2=0.26 $Y2=0.81
.ends

