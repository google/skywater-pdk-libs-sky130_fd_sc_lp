* NGSPICE file created from sky130_fd_sc_lp__nand2b_m.ext - technology: sky130A

.subckt sky130_fd_sc_lp__nand2b_m A_N B VGND VNB VPB VPWR Y
M1000 VPWR a_46_54# Y VPB phighvt w=420000u l=150000u
+  ad=2.289e+11p pd=2.77e+06u as=1.176e+11p ps=1.4e+06u
M1001 a_282_54# B VGND VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=2.583e+11p ps=2.07e+06u
M1002 Y a_46_54# a_282_54# VNB nshort w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1003 Y B VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VGND A_N a_46_54# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1005 VPWR A_N a_46_54# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
.ends

