# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__buflp_4
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__buflp_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.280000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.965000 1.180000 4.430000 1.515000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  1.352400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 0.975000 2.945000 1.145000 ;
        RECT 0.125000 1.145000 0.355000 1.780000 ;
        RECT 0.185000 1.780000 0.355000 1.815000 ;
        RECT 0.185000 1.815000 3.235000 1.985000 ;
        RECT 1.835000 0.595000 2.085000 0.975000 ;
        RECT 1.905000 1.985000 2.235000 2.735000 ;
        RECT 2.775000 0.595000 2.945000 0.975000 ;
        RECT 2.905000 1.985000 3.235000 2.735000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 5.280000 0.085000 ;
        RECT 0.115000  0.085000 0.365000 0.805000 ;
        RECT 0.975000  0.085000 1.305000 0.465000 ;
        RECT 3.625000  0.085000 3.955000 0.670000 ;
      LAYER mcon ;
        RECT 0.155000 -0.085000 0.325000 0.085000 ;
        RECT 0.635000 -0.085000 0.805000 0.085000 ;
        RECT 1.115000 -0.085000 1.285000 0.085000 ;
        RECT 1.595000 -0.085000 1.765000 0.085000 ;
        RECT 2.075000 -0.085000 2.245000 0.085000 ;
        RECT 2.555000 -0.085000 2.725000 0.085000 ;
        RECT 3.035000 -0.085000 3.205000 0.085000 ;
        RECT 3.515000 -0.085000 3.685000 0.085000 ;
        RECT 3.995000 -0.085000 4.165000 0.085000 ;
        RECT 4.475000 -0.085000 4.645000 0.085000 ;
        RECT 4.955000 -0.085000 5.125000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 5.280000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.245000 5.280000 3.415000 ;
        RECT 0.115000 2.155000 0.365000 3.245000 ;
        RECT 1.055000 2.495000 1.225000 3.245000 ;
        RECT 3.905000 1.815000 4.235000 3.245000 ;
      LAYER mcon ;
        RECT 0.155000 3.245000 0.325000 3.415000 ;
        RECT 0.635000 3.245000 0.805000 3.415000 ;
        RECT 1.115000 3.245000 1.285000 3.415000 ;
        RECT 1.595000 3.245000 1.765000 3.415000 ;
        RECT 2.075000 3.245000 2.245000 3.415000 ;
        RECT 2.555000 3.245000 2.725000 3.415000 ;
        RECT 3.035000 3.245000 3.205000 3.415000 ;
        RECT 3.515000 3.245000 3.685000 3.415000 ;
        RECT 3.995000 3.245000 4.165000 3.415000 ;
        RECT 4.475000 3.245000 4.645000 3.415000 ;
        RECT 4.955000 3.245000 5.125000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 5.280000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.545000 0.255000 0.795000 0.635000 ;
      RECT 0.545000 0.635000 1.655000 0.805000 ;
      RECT 0.545000 2.155000 1.735000 2.325000 ;
      RECT 0.545000 2.325000 0.875000 3.075000 ;
      RECT 0.745000 1.315000 3.795000 1.645000 ;
      RECT 1.405000 2.325000 1.735000 2.905000 ;
      RECT 1.405000 2.905000 3.735000 3.075000 ;
      RECT 1.485000 0.255000 3.455000 0.425000 ;
      RECT 1.485000 0.425000 1.655000 0.635000 ;
      RECT 2.265000 0.425000 2.595000 0.805000 ;
      RECT 2.405000 2.155000 2.735000 2.905000 ;
      RECT 3.125000 0.425000 3.455000 1.095000 ;
      RECT 3.405000 1.815000 3.735000 2.905000 ;
      RECT 3.625000 0.840000 5.125000 1.010000 ;
      RECT 3.625000 1.010000 3.795000 1.315000 ;
      RECT 4.795000 0.255000 5.125000 0.840000 ;
      RECT 4.795000 1.010000 5.125000 3.075000 ;
  END
END sky130_fd_sc_lp__buflp_4
