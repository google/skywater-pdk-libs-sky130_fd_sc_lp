* File: sky130_fd_sc_lp__and3b_lp.spice
* Created: Wed Sep  2 09:32:25 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__and3b_lp.pex.spice"
.subckt sky130_fd_sc_lp__and3b_lp  VNB VPB A_N B C VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* C	C
* B	B
* A_N	A_N
* VPB	VPB
* VNB	VNB
MM1005 A_114_57# N_A_N_M1005_g N_VGND_M1005_s VNB NSHORT L=0.15 W=0.42 AD=0.0504
+ AS=0.1197 PD=0.66 PS=1.41 NRD=18.564 NRS=0 M=1 R=2.8 SA=75000.2 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1011 N_A_137_408#_M1011_d N_A_N_M1011_g A_114_57# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0504 PD=1.41 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1001 A_391_57# N_A_137_408#_M1001_g N_A_248_409#_M1001_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0504 AS=0.1197 PD=0.66 PS=1.41 NRD=18.564 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.9 A=0.063 P=1.14 MULT=1
MM1006 A_469_57# N_B_M1006_g A_391_57# VNB NSHORT L=0.15 W=0.42 AD=0.0504
+ AS=0.0504 PD=0.66 PS=0.66 NRD=18.564 NRS=18.564 M=1 R=2.8 SA=75000.6
+ SB=75001.6 A=0.063 P=1.14 MULT=1
MM1007 N_VGND_M1007_d N_C_M1007_g A_469_57# VNB NSHORT L=0.15 W=0.42 AD=0.09345
+ AS=0.0504 PD=0.865 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75001 SB=75001.2
+ A=0.063 P=1.14 MULT=1
MM1000 A_666_57# N_A_248_409#_M1000_g N_VGND_M1007_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.09345 PD=0.63 PS=0.865 NRD=14.28 NRS=47.136 M=1 R=2.8
+ SA=75001.6 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1002 N_X_M1002_d N_A_248_409#_M1002_g A_666_57# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.9
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1009 N_A_137_408#_M1009_d N_A_N_M1009_g N_VPWR_M1009_s VPB PHIGHVT L=0.25 W=1
+ AD=0.285 AS=0.285 PD=2.57 PS=2.57 NRD=0 NRS=0 M=1 R=4 SA=125000 SB=125000
+ A=0.25 P=2.5 MULT=1
MM1008 N_VPWR_M1008_d N_A_137_408#_M1008_g N_A_248_409#_M1008_s VPB PHIGHVT
+ L=0.25 W=1 AD=0.14 AS=0.285 PD=1.28 PS=2.57 NRD=0 NRS=0 M=1 R=4 SA=125000
+ SB=125002 A=0.25 P=2.5 MULT=1
MM1003 N_A_248_409#_M1003_d N_B_M1003_g N_VPWR_M1008_d VPB PHIGHVT L=0.25 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125001 SB=125001 A=0.25
+ P=2.5 MULT=1
MM1010 N_VPWR_M1010_d N_C_M1010_g N_A_248_409#_M1003_d VPB PHIGHVT L=0.25 W=1
+ AD=0.1925 AS=0.14 PD=1.385 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125001 SB=125001
+ A=0.25 P=2.5 MULT=1
MM1004 N_X_M1004_d N_A_248_409#_M1004_g N_VPWR_M1010_d VPB PHIGHVT L=0.25 W=1
+ AD=0.285 AS=0.1925 PD=2.57 PS=1.385 NRD=0 NRS=20.685 M=1 R=4 SA=125002
+ SB=125000 A=0.25 P=2.5 MULT=1
DX12_noxref VNB VPB NWDIODE A=8.7655 P=13.13
*
.include "sky130_fd_sc_lp__and3b_lp.pxi.spice"
*
.ends
*
*
