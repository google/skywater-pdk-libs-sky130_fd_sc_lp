* File: sky130_fd_sc_lp__nand2b_1.pxi.spice
* Created: Wed Sep  2 10:03:26 2020
* 
x_PM_SKY130_FD_SC_LP__NAND2B_1%A_N N_A_N_M1004_g N_A_N_M1000_g N_A_N_c_49_n
+ N_A_N_c_50_n A_N N_A_N_c_51_n N_A_N_c_52_n PM_SKY130_FD_SC_LP__NAND2B_1%A_N
x_PM_SKY130_FD_SC_LP__NAND2B_1%B N_B_M1002_g N_B_c_79_n N_B_M1003_g B B
+ N_B_c_81_n PM_SKY130_FD_SC_LP__NAND2B_1%B
x_PM_SKY130_FD_SC_LP__NAND2B_1%A_40_367# N_A_40_367#_M1000_s N_A_40_367#_M1004_s
+ N_A_40_367#_M1005_g N_A_40_367#_M1001_g N_A_40_367#_c_122_n
+ N_A_40_367#_c_123_n N_A_40_367#_c_124_n N_A_40_367#_c_134_n
+ N_A_40_367#_c_125_n N_A_40_367#_c_126_n N_A_40_367#_c_127_n
+ N_A_40_367#_c_128_n N_A_40_367#_c_129_n N_A_40_367#_c_130_n
+ N_A_40_367#_c_131_n N_A_40_367#_c_132_n PM_SKY130_FD_SC_LP__NAND2B_1%A_40_367#
x_PM_SKY130_FD_SC_LP__NAND2B_1%VPWR N_VPWR_M1004_d N_VPWR_M1005_d N_VPWR_c_204_n
+ N_VPWR_c_205_n VPWR N_VPWR_c_206_n N_VPWR_c_207_n N_VPWR_c_203_n
+ N_VPWR_c_209_n N_VPWR_c_210_n PM_SKY130_FD_SC_LP__NAND2B_1%VPWR
x_PM_SKY130_FD_SC_LP__NAND2B_1%Y N_Y_M1001_d N_Y_M1002_d N_Y_c_231_n N_Y_c_228_n
+ N_Y_c_229_n N_Y_c_233_n N_Y_c_230_n Y Y PM_SKY130_FD_SC_LP__NAND2B_1%Y
x_PM_SKY130_FD_SC_LP__NAND2B_1%VGND N_VGND_M1000_d N_VGND_c_259_n N_VGND_c_260_n
+ N_VGND_c_261_n VGND N_VGND_c_262_n N_VGND_c_263_n
+ PM_SKY130_FD_SC_LP__NAND2B_1%VGND
cc_1 VNB N_A_N_M1004_g 0.00391126f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=2.045
cc_2 VNB N_A_N_M1000_g 0.0219095f $X=-0.19 $Y=-0.245 $X2=0.76 $Y2=0.445
cc_3 VNB N_A_N_c_49_n 0.047376f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=0.945
cc_4 VNB N_A_N_c_50_n 0.0364142f $X=-0.19 $Y=-0.245 $X2=0.37 $Y2=1.605
cc_5 VNB N_A_N_c_51_n 0.0451207f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.1
cc_6 VNB N_A_N_c_52_n 0.0223567f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.1
cc_7 VNB N_B_M1002_g 0.00768469f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=2.045
cc_8 VNB N_B_c_79_n 0.016616f $X=-0.19 $Y=-0.245 $X2=0.76 $Y2=0.795
cc_9 VNB B 0.00939957f $X=-0.19 $Y=-0.245 $X2=0.37 $Y2=0.945
cc_10 VNB N_B_c_81_n 0.0412395f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_40_367#_c_122_n 0.0122431f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_40_367#_c_123_n 0.0201197f $X=-0.19 $Y=-0.245 $X2=0.37 $Y2=1.1
cc_13 VNB N_A_40_367#_c_124_n 0.0185076f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.1
cc_14 VNB N_A_40_367#_c_125_n 0.0152117f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_40_367#_c_126_n 0.00235232f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_40_367#_c_127_n 0.0048873f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_40_367#_c_128_n 0.00557475f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_40_367#_c_129_n 0.00135177f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_40_367#_c_130_n 0.00116587f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_40_367#_c_131_n 0.00569552f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_40_367#_c_132_n 0.0176228f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_VPWR_c_203_n 0.103974f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_Y_c_228_n 0.0305318f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=0.945
cc_24 VNB N_Y_c_229_n 0.0289506f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_25 VNB N_Y_c_230_n 0.0206818f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.1
cc_26 VNB N_VGND_c_259_n 0.002833f $X=-0.19 $Y=-0.245 $X2=0.76 $Y2=0.445
cc_27 VNB N_VGND_c_260_n 0.0238547f $X=-0.19 $Y=-0.245 $X2=0.37 $Y2=0.945
cc_28 VNB N_VGND_c_261_n 0.00510363f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=0.795
cc_29 VNB N_VGND_c_262_n 0.0353786f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_263_n 0.15629f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.27
cc_31 VPB N_A_N_M1004_g 0.0310631f $X=-0.19 $Y=1.655 $X2=0.54 $Y2=2.045
cc_32 VPB N_B_M1002_g 0.0223182f $X=-0.19 $Y=1.655 $X2=0.54 $Y2=2.045
cc_33 VPB N_A_40_367#_c_122_n 0.0342319f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_34 VPB N_A_40_367#_c_134_n 0.0148521f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_35 VPB N_A_40_367#_c_128_n 0.00596438f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_36 VPB N_A_40_367#_c_129_n 0.0100772f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_37 VPB N_A_40_367#_c_131_n 0.0013059f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_38 VPB N_VPWR_c_204_n 0.0325139f $X=-0.19 $Y=1.655 $X2=0.48 $Y2=0.945
cc_39 VPB N_VPWR_c_205_n 0.0341734f $X=-0.19 $Y=1.655 $X2=0.29 $Y2=1.1
cc_40 VPB N_VPWR_c_206_n 0.0154314f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_41 VPB N_VPWR_c_207_n 0.0188498f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_42 VPB N_VPWR_c_203_n 0.0857654f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_43 VPB N_VPWR_c_209_n 0.0289132f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_44 VPB N_VPWR_c_210_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_45 VPB N_Y_c_231_n 0.0331841f $X=-0.19 $Y=1.655 $X2=0.76 $Y2=0.445
cc_46 VPB N_Y_c_229_n 0.0163055f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_47 N_A_N_c_50_n N_B_M1002_g 0.0202416f $X=0.37 $Y=1.605 $X2=0 $Y2=0
cc_48 N_A_N_M1000_g N_B_c_79_n 0.0221142f $X=0.76 $Y=0.445 $X2=0 $Y2=0
cc_49 N_A_N_c_51_n N_B_c_79_n 0.00435973f $X=0.29 $Y=1.1 $X2=0 $Y2=0
cc_50 N_A_N_c_49_n B 0.00586842f $X=0.48 $Y=0.945 $X2=0 $Y2=0
cc_51 N_A_N_c_51_n B 0.00503276f $X=0.29 $Y=1.1 $X2=0 $Y2=0
cc_52 N_A_N_c_52_n B 0.0355695f $X=0.29 $Y=1.1 $X2=0 $Y2=0
cc_53 N_A_N_c_51_n N_B_c_81_n 0.0162358f $X=0.29 $Y=1.1 $X2=0 $Y2=0
cc_54 N_A_N_c_52_n N_B_c_81_n 5.69533e-19 $X=0.29 $Y=1.1 $X2=0 $Y2=0
cc_55 N_A_N_M1004_g N_A_40_367#_c_134_n 0.00621462f $X=0.54 $Y=2.045 $X2=0 $Y2=0
cc_56 N_A_N_M1000_g N_A_40_367#_c_125_n 0.00107237f $X=0.76 $Y=0.445 $X2=0 $Y2=0
cc_57 N_A_N_M1000_g N_A_40_367#_c_126_n 0.00905216f $X=0.76 $Y=0.445 $X2=0 $Y2=0
cc_58 N_A_N_c_49_n N_A_40_367#_c_126_n 0.00386171f $X=0.48 $Y=0.945 $X2=0 $Y2=0
cc_59 N_A_N_c_49_n N_A_40_367#_c_127_n 0.0191306f $X=0.48 $Y=0.945 $X2=0 $Y2=0
cc_60 N_A_N_c_52_n N_A_40_367#_c_127_n 0.00609484f $X=0.29 $Y=1.1 $X2=0 $Y2=0
cc_61 N_A_N_M1004_g N_A_40_367#_c_129_n 0.0247185f $X=0.54 $Y=2.045 $X2=0 $Y2=0
cc_62 N_A_N_c_49_n N_A_40_367#_c_129_n 3.73644e-19 $X=0.48 $Y=0.945 $X2=0 $Y2=0
cc_63 N_A_N_c_50_n N_A_40_367#_c_129_n 0.00950705f $X=0.37 $Y=1.605 $X2=0 $Y2=0
cc_64 N_A_N_c_52_n N_A_40_367#_c_129_n 0.0250801f $X=0.29 $Y=1.1 $X2=0 $Y2=0
cc_65 N_A_N_M1004_g N_VPWR_c_204_n 0.00615905f $X=0.54 $Y=2.045 $X2=0 $Y2=0
cc_66 N_A_N_M1004_g N_Y_c_233_n 2.95428e-19 $X=0.54 $Y=2.045 $X2=0 $Y2=0
cc_67 N_A_N_M1000_g N_VGND_c_259_n 0.00927153f $X=0.76 $Y=0.445 $X2=0 $Y2=0
cc_68 N_A_N_M1000_g N_VGND_c_260_n 0.00358332f $X=0.76 $Y=0.445 $X2=0 $Y2=0
cc_69 N_A_N_M1000_g N_VGND_c_263_n 0.00547277f $X=0.76 $Y=0.445 $X2=0 $Y2=0
cc_70 N_A_N_c_49_n N_VGND_c_263_n 0.00673004f $X=0.48 $Y=0.945 $X2=0 $Y2=0
cc_71 N_B_M1002_g N_A_40_367#_c_122_n 0.0225616f $X=1.065 $Y=2.465 $X2=0 $Y2=0
cc_72 B N_A_40_367#_c_123_n 3.20537e-19 $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_73 N_B_c_81_n N_A_40_367#_c_123_n 0.0439857f $X=1.065 $Y=1.35 $X2=0 $Y2=0
cc_74 N_B_c_79_n N_A_40_367#_c_124_n 0.0379232f $X=1.27 $Y=1.185 $X2=0 $Y2=0
cc_75 B N_A_40_367#_c_124_n 2.97937e-19 $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_76 N_B_M1002_g N_A_40_367#_c_134_n 6.22473e-19 $X=1.065 $Y=2.465 $X2=0 $Y2=0
cc_77 N_B_c_79_n N_A_40_367#_c_126_n 0.013599f $X=1.27 $Y=1.185 $X2=0 $Y2=0
cc_78 B N_A_40_367#_c_126_n 0.0454673f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_79 N_B_c_81_n N_A_40_367#_c_126_n 0.00137707f $X=1.065 $Y=1.35 $X2=0 $Y2=0
cc_80 B N_A_40_367#_c_127_n 0.00126545f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_81 N_B_M1002_g N_A_40_367#_c_128_n 0.0147147f $X=1.065 $Y=2.465 $X2=0 $Y2=0
cc_82 B N_A_40_367#_c_128_n 0.0388114f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_83 N_B_c_81_n N_A_40_367#_c_128_n 0.00714203f $X=1.065 $Y=1.35 $X2=0 $Y2=0
cc_84 N_B_M1002_g N_A_40_367#_c_129_n 0.00237622f $X=1.065 $Y=2.465 $X2=0 $Y2=0
cc_85 B N_A_40_367#_c_129_n 0.0129789f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_86 N_B_c_79_n N_A_40_367#_c_130_n 0.00510375f $X=1.27 $Y=1.185 $X2=0 $Y2=0
cc_87 B N_A_40_367#_c_130_n 0.0204901f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_88 N_B_M1002_g N_A_40_367#_c_131_n 0.00150108f $X=1.065 $Y=2.465 $X2=0 $Y2=0
cc_89 B N_A_40_367#_c_131_n 0.0141307f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_90 N_B_c_81_n N_A_40_367#_c_131_n 0.00268658f $X=1.065 $Y=1.35 $X2=0 $Y2=0
cc_91 N_B_M1002_g N_A_40_367#_c_132_n 0.00142794f $X=1.065 $Y=2.465 $X2=0 $Y2=0
cc_92 N_B_M1002_g N_VPWR_c_204_n 0.00318541f $X=1.065 $Y=2.465 $X2=0 $Y2=0
cc_93 N_B_M1002_g N_VPWR_c_205_n 7.21976e-19 $X=1.065 $Y=2.465 $X2=0 $Y2=0
cc_94 N_B_M1002_g N_VPWR_c_206_n 0.0054895f $X=1.065 $Y=2.465 $X2=0 $Y2=0
cc_95 N_B_M1002_g N_VPWR_c_203_n 0.0110907f $X=1.065 $Y=2.465 $X2=0 $Y2=0
cc_96 N_B_M1002_g N_Y_c_233_n 0.00292711f $X=1.065 $Y=2.465 $X2=0 $Y2=0
cc_97 N_B_M1002_g Y 0.0112401f $X=1.065 $Y=2.465 $X2=0 $Y2=0
cc_98 B N_VGND_M1000_d 0.00211465f $X=1.115 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_99 N_B_c_79_n N_VGND_c_259_n 0.00443027f $X=1.27 $Y=1.185 $X2=0 $Y2=0
cc_100 N_B_c_79_n N_VGND_c_262_n 0.00430895f $X=1.27 $Y=1.185 $X2=0 $Y2=0
cc_101 N_B_c_79_n N_VGND_c_263_n 0.00605595f $X=1.27 $Y=1.185 $X2=0 $Y2=0
cc_102 N_A_40_367#_c_129_n N_VPWR_M1004_d 0.00199132f $X=0.78 $Y=1.69 $X2=-0.19
+ $Y2=-0.245
cc_103 N_A_40_367#_c_134_n N_VPWR_c_204_n 0.0120001f $X=0.325 $Y=2.045 $X2=0
+ $Y2=0
cc_104 N_A_40_367#_c_128_n N_VPWR_c_204_n 0.00959225f $X=1.455 $Y=1.69 $X2=0
+ $Y2=0
cc_105 N_A_40_367#_c_129_n N_VPWR_c_204_n 0.00791206f $X=0.78 $Y=1.69 $X2=0
+ $Y2=0
cc_106 N_A_40_367#_c_122_n N_VPWR_c_205_n 0.0164616f $X=1.66 $Y=1.725 $X2=0
+ $Y2=0
cc_107 N_A_40_367#_c_122_n N_VPWR_c_206_n 0.00486043f $X=1.66 $Y=1.725 $X2=0
+ $Y2=0
cc_108 N_A_40_367#_c_122_n N_VPWR_c_203_n 0.0082726f $X=1.66 $Y=1.725 $X2=0
+ $Y2=0
cc_109 N_A_40_367#_c_122_n N_Y_c_231_n 0.0213441f $X=1.66 $Y=1.725 $X2=0 $Y2=0
cc_110 N_A_40_367#_c_128_n N_Y_c_231_n 0.0039988f $X=1.455 $Y=1.69 $X2=0 $Y2=0
cc_111 N_A_40_367#_c_131_n N_Y_c_231_n 0.0236738f $X=1.735 $Y=1.44 $X2=0 $Y2=0
cc_112 N_A_40_367#_c_124_n N_Y_c_228_n 0.0107571f $X=1.727 $Y=1.185 $X2=0 $Y2=0
cc_113 N_A_40_367#_c_126_n N_Y_c_228_n 0.0144456f $X=1.455 $Y=0.76 $X2=0 $Y2=0
cc_114 N_A_40_367#_c_122_n N_Y_c_229_n 0.00785484f $X=1.66 $Y=1.725 $X2=0 $Y2=0
cc_115 N_A_40_367#_c_123_n N_Y_c_229_n 0.00471902f $X=1.727 $Y=1.357 $X2=0 $Y2=0
cc_116 N_A_40_367#_c_124_n N_Y_c_229_n 0.00157144f $X=1.727 $Y=1.185 $X2=0 $Y2=0
cc_117 N_A_40_367#_c_130_n N_Y_c_229_n 0.00641851f $X=1.54 $Y=1.275 $X2=0 $Y2=0
cc_118 N_A_40_367#_c_131_n N_Y_c_229_n 0.0332374f $X=1.735 $Y=1.44 $X2=0 $Y2=0
cc_119 N_A_40_367#_c_134_n N_Y_c_233_n 0.00242868f $X=0.325 $Y=2.045 $X2=0 $Y2=0
cc_120 N_A_40_367#_c_128_n N_Y_c_233_n 0.0181975f $X=1.455 $Y=1.69 $X2=0 $Y2=0
cc_121 N_A_40_367#_c_123_n N_Y_c_230_n 0.0029616f $X=1.727 $Y=1.357 $X2=0 $Y2=0
cc_122 N_A_40_367#_c_130_n N_Y_c_230_n 0.0192004f $X=1.54 $Y=1.275 $X2=0 $Y2=0
cc_123 N_A_40_367#_c_131_n N_Y_c_230_n 0.00843873f $X=1.735 $Y=1.44 $X2=0 $Y2=0
cc_124 N_A_40_367#_c_126_n N_VGND_M1000_d 0.00371103f $X=1.455 $Y=0.76 $X2=-0.19
+ $Y2=-0.245
cc_125 N_A_40_367#_c_126_n N_VGND_c_259_n 0.0227013f $X=1.455 $Y=0.76 $X2=0
+ $Y2=0
cc_126 N_A_40_367#_c_125_n N_VGND_c_260_n 0.0151488f $X=0.545 $Y=0.445 $X2=0
+ $Y2=0
cc_127 N_A_40_367#_c_126_n N_VGND_c_260_n 0.00260179f $X=1.455 $Y=0.76 $X2=0
+ $Y2=0
cc_128 N_A_40_367#_c_124_n N_VGND_c_262_n 0.00513223f $X=1.727 $Y=1.185 $X2=0
+ $Y2=0
cc_129 N_A_40_367#_c_126_n N_VGND_c_262_n 0.00646913f $X=1.455 $Y=0.76 $X2=0
+ $Y2=0
cc_130 N_A_40_367#_M1000_s N_VGND_c_263_n 0.00234689f $X=0.42 $Y=0.235 $X2=0
+ $Y2=0
cc_131 N_A_40_367#_c_124_n N_VGND_c_263_n 0.00955383f $X=1.727 $Y=1.185 $X2=0
+ $Y2=0
cc_132 N_A_40_367#_c_125_n N_VGND_c_263_n 0.00985676f $X=0.545 $Y=0.445 $X2=0
+ $Y2=0
cc_133 N_A_40_367#_c_126_n N_VGND_c_263_n 0.0180823f $X=1.455 $Y=0.76 $X2=0
+ $Y2=0
cc_134 N_A_40_367#_c_126_n A_269_47# 0.00375224f $X=1.455 $Y=0.76 $X2=-0.19
+ $Y2=-0.245
cc_135 N_A_40_367#_c_130_n A_269_47# 0.00238932f $X=1.54 $Y=1.275 $X2=-0.19
+ $Y2=-0.245
cc_136 N_VPWR_c_203_n N_Y_M1002_d 0.00380103f $X=2.16 $Y=3.33 $X2=0 $Y2=0
cc_137 N_VPWR_M1005_d N_Y_c_231_n 0.00533633f $X=1.57 $Y=1.835 $X2=0 $Y2=0
cc_138 N_VPWR_c_205_n N_Y_c_231_n 0.0220026f $X=1.71 $Y=2.415 $X2=0 $Y2=0
cc_139 N_VPWR_c_206_n Y 0.015688f $X=1.545 $Y=3.33 $X2=0 $Y2=0
cc_140 N_VPWR_c_203_n Y 0.00984745f $X=2.16 $Y=3.33 $X2=0 $Y2=0
cc_141 N_Y_c_228_n N_VGND_c_262_n 0.0367916f $X=1.88 $Y=0.42 $X2=0 $Y2=0
cc_142 N_Y_M1001_d N_VGND_c_263_n 0.0059108f $X=1.705 $Y=0.235 $X2=0 $Y2=0
cc_143 N_Y_c_228_n N_VGND_c_263_n 0.0201386f $X=1.88 $Y=0.42 $X2=0 $Y2=0
cc_144 N_VGND_c_263_n A_269_47# 0.00256287f $X=2.16 $Y=0 $X2=-0.19 $Y2=-0.245
