* File: sky130_fd_sc_lp__sleep_pargate_plv_21.pex.spice
* Created: Wed Sep  2 10:37:41 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__SLEEP_PARGATE_PLV_21%SLEEP 1 3 4 6 7 9 13 15 16 17
+ 18 19 26 29
r55 29 30 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=8.42
+ $Y=2.665 $X2=8.42 $Y2=2.665
r56 19 30 5.86755 $w=5.28e-07 $l=2.6e-07 $layer=LI1_cond $X=8.52 $Y=2.405
+ $X2=8.52 $Y2=2.665
r57 18 19 9.47836 $w=5.28e-07 $l=4.2e-07 $layer=LI1_cond $X=8.52 $Y=1.985
+ $X2=8.52 $Y2=2.405
r58 18 26 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=8.42
+ $Y=1.985 $X2=8.42 $Y2=1.985
r59 17 18 7.22161 $w=5.28e-07 $l=3.2e-07 $layer=LI1_cond $X=8.52 $Y=1.665
+ $X2=8.52 $Y2=1.985
r60 16 17 8.34998 $w=5.28e-07 $l=3.7e-07 $layer=LI1_cond $X=8.52 $Y=1.295
+ $X2=8.52 $Y2=1.665
r61 15 16 8.34998 $w=5.28e-07 $l=3.7e-07 $layer=LI1_cond $X=8.52 $Y=0.925
+ $X2=8.52 $Y2=1.295
r62 14 29 2.01019 $w=4.15e-07 $l=1.5e-08 $layer=POLY_cond $X=8.377 $Y=2.68
+ $X2=8.377 $Y2=2.665
r63 12 29 35.5134 $w=4.15e-07 $l=2.65e-07 $layer=POLY_cond $X=8.377 $Y=2.4
+ $X2=8.377 $Y2=2.665
r64 12 13 8.21244 $w=4.15e-07 $l=7.5e-08 $layer=POLY_cond $X=8.377 $Y=2.4
+ $X2=8.377 $Y2=2.325
r65 11 26 35.5134 $w=4.15e-07 $l=2.65e-07 $layer=POLY_cond $X=8.377 $Y=2.25
+ $X2=8.377 $Y2=1.985
r66 11 13 8.21244 $w=4.15e-07 $l=7.5e-08 $layer=POLY_cond $X=8.377 $Y=2.25
+ $X2=8.377 $Y2=2.325
r67 10 26 2.01019 $w=4.15e-07 $l=1.5e-08 $layer=POLY_cond $X=8.377 $Y=1.97
+ $X2=8.377 $Y2=1.985
r68 7 14 35.4752 $w=1.5e-07 $l=2.41607e-07 $layer=POLY_cond $X=8.17 $Y=2.755
+ $X2=8.377 $Y2=2.68
r69 7 9 1161.62 $w=1.5e-07 $l=3.615e-06 $layer=POLY_cond $X=8.17 $Y=2.755
+ $X2=4.555 $Y2=2.755
r70 4 13 20.4038 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=8.17 $Y=2.325
+ $X2=8.377 $Y2=2.325
r71 4 6 1161.62 $w=1.5e-07 $l=3.615e-06 $layer=POLY_cond $X=8.17 $Y=2.325
+ $X2=4.555 $Y2=2.325
r72 1 10 35.4752 $w=1.5e-07 $l=2.41607e-07 $layer=POLY_cond $X=8.17 $Y=1.895
+ $X2=8.377 $Y2=1.97
r73 1 3 1161.62 $w=1.5e-07 $l=3.615e-06 $layer=POLY_cond $X=8.17 $Y=1.895
+ $X2=4.555 $Y2=1.895
.ends

.subckt PM_SKY130_FD_SC_LP__SLEEP_PARGATE_PLV_21%VPWR 1 2 7 25 45 50 56 62 68 74
+ 75
c92 68 0 9.06808e-20 $X=6.2 $Y=1.68
c93 62 0 9.06808e-20 $X=4.645 $Y=1.68
c94 56 0 9.06808e-20 $X=3.09 $Y=1.68
c95 1 0 1.81343e-19 $X=1.055 $Y=1.555
r96 74 75 1.125 $w=1.5e-07 $l=6e-07 $layer=via $count=4 $X=7.775 $Y=1.68
+ $X2=7.775 $Y2=1.68
r97 69 75 0.0591216 $w=3.33e-06 $l=1.575e-06 $layer=MET2_cond $X=6.2 $Y=1.665
+ $X2=7.775 $Y2=1.665
r98 68 69 1.125 $w=1.5e-07 $l=6e-07 $layer=via $count=4 $X=6.2 $Y=1.68 $X2=6.2
+ $Y2=1.68
r99 63 69 0.0583709 $w=3.33e-06 $l=1.555e-06 $layer=MET2_cond $X=4.645 $Y=1.665
+ $X2=6.2 $Y2=1.665
r100 62 63 1.125 $w=1.5e-07 $l=6e-07 $layer=via $count=4 $X=4.645 $Y=1.68
+ $X2=4.645 $Y2=1.68
r101 56 57 1.125 $w=1.5e-07 $l=6e-07 $layer=via $count=4 $X=3.09 $Y=1.68
+ $X2=3.09 $Y2=1.68
r102 51 57 0.0579955 $w=3.33e-06 $l=1.545e-06 $layer=MET2_cond $X=1.545 $Y=1.665
+ $X2=3.09 $Y2=1.665
r103 50 51 1.125 $w=1.5e-07 $l=6e-07 $layer=via $count=4 $X=1.545 $Y=1.68
+ $X2=1.545 $Y2=1.68
r104 47 74 0.173696 $w=6.5e-07 $l=8.6e-07 $layer=MET1_cond $X=7.62 $Y=2.54
+ $X2=7.62 $Y2=1.68
r105 45 47 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.8 $Y=2.54
+ $X2=7.8 $Y2=2.54
r106 43 68 0.173696 $w=6.5e-07 $l=8.6e-07 $layer=MET1_cond $X=6.045 $Y=2.54
+ $X2=6.045 $Y2=1.68
r107 42 45 69.1466 $w=2.58e-07 $l=1.56e-06 $layer=LI1_cond $X=6.225 $Y=2.54
+ $X2=7.785 $Y2=2.54
r108 42 43 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.225 $Y=2.54
+ $X2=6.225 $Y2=2.54
r109 40 62 0.173696 $w=6.5e-07 $l=8.6e-07 $layer=MET1_cond $X=4.49 $Y=2.54
+ $X2=4.49 $Y2=1.68
r110 39 42 68.925 $w=2.58e-07 $l=1.555e-06 $layer=LI1_cond $X=4.67 $Y=2.54
+ $X2=6.225 $Y2=2.54
r111 39 40 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.67 $Y=2.54
+ $X2=4.67 $Y2=2.54
r112 37 56 0.173696 $w=6.5e-07 $l=8.6e-07 $layer=MET1_cond $X=2.935 $Y=2.54
+ $X2=2.935 $Y2=1.68
r113 36 39 68.925 $w=2.58e-07 $l=1.555e-06 $layer=LI1_cond $X=3.115 $Y=2.54
+ $X2=4.67 $Y2=2.54
r114 36 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.115 $Y=2.54
+ $X2=3.115 $Y2=2.54
r115 34 50 0.173696 $w=6.5e-07 $l=8.6e-07 $layer=MET1_cond $X=1.38 $Y=2.54
+ $X2=1.38 $Y2=1.68
r116 33 36 68.925 $w=2.58e-07 $l=1.555e-06 $layer=LI1_cond $X=1.56 $Y=2.54
+ $X2=3.115 $Y2=2.54
r117 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.56 $Y=2.54
+ $X2=1.56 $Y2=2.54
r118 30 33 10.4163 $w=2.58e-07 $l=2.35e-07 $layer=LI1_cond $X=1.325 $Y=2.54
+ $X2=1.56 $Y2=2.54
r119 25 74 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.8 $Y=1.68
+ $X2=7.8 $Y2=1.68
r120 22 25 69.1466 $w=2.58e-07 $l=1.56e-06 $layer=LI1_cond $X=6.225 $Y=1.68
+ $X2=7.785 $Y2=1.68
r121 22 68 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.225 $Y=1.68
+ $X2=6.225 $Y2=1.68
r122 19 22 68.925 $w=2.58e-07 $l=1.555e-06 $layer=LI1_cond $X=4.67 $Y=1.68
+ $X2=6.225 $Y2=1.68
r123 19 62 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.67 $Y=1.68
+ $X2=4.67 $Y2=1.68
r124 16 19 68.925 $w=2.58e-07 $l=1.555e-06 $layer=LI1_cond $X=3.115 $Y=1.68
+ $X2=4.67 $Y2=1.68
r125 16 56 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.115 $Y=1.68
+ $X2=3.115 $Y2=1.68
r126 13 16 68.925 $w=2.58e-07 $l=1.555e-06 $layer=LI1_cond $X=1.56 $Y=1.68
+ $X2=3.115 $Y2=1.68
r127 13 50 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.56 $Y=1.68
+ $X2=1.56 $Y2=1.68
r128 10 13 10.4163 $w=2.58e-07 $l=2.35e-07 $layer=LI1_cond $X=1.325 $Y=1.68
+ $X2=1.56 $Y2=1.68
r129 7 63 0.00319069 $w=3.33e-06 $l=8.5e-08 $layer=MET2_cond $X=4.56 $Y=1.665
+ $X2=4.645 $Y2=1.665
r130 7 57 0.0551802 $w=3.33e-06 $l=1.47e-06 $layer=MET2_cond $X=4.56 $Y=1.665
+ $X2=3.09 $Y2=1.665
r131 2 45 60 $w=1.7e-07 $l=6.79964e-06 $layer=licon1_PDIFF $count=10 $X=1.055
+ $Y=2.4 $X2=7.785 $Y2=2.54
r132 2 30 60 $w=1.7e-07 $l=3.32716e-07 $layer=licon1_PDIFF $count=10 $X=1.055
+ $Y=2.4 $X2=1.325 $Y2=2.54
r133 1 25 60 $w=1.7e-07 $l=6.79221e-06 $layer=licon1_PDIFF $count=10 $X=1.055
+ $Y=1.555 $X2=7.785 $Y2=1.68
r134 1 10 60 $w=1.7e-07 $l=3.26573e-07 $layer=licon1_PDIFF $count=10 $X=1.055
+ $Y=1.555 $X2=1.325 $Y2=1.68
.ends

.subckt PM_SKY130_FD_SC_LP__SLEEP_PARGATE_PLV_21%VIRTPWR 1 2 7 11 12 30 66 69 72
+ 75 77 81 82 89 90 95 99 104 105
c100 105 0 1.43534e-19 $X=6.51 $Y=3.33
c101 99 0 1.43534e-19 $X=4.955 $Y=3.33
c102 95 0 1.43534e-19 $X=3.4 $Y=3.33
c103 75 0 4.53393e-20 $X=7.005 $Y=2.11
c104 72 0 4.53347e-20 $X=5.45 $Y=2.11
c105 69 0 4.53347e-20 $X=3.895 $Y=2.11
c106 66 0 4.53347e-20 $X=2.34 $Y=2.11
c107 12 0 3.89769e-19 $X=0 $Y=3.085
c108 1 0 2.72043e-19 $X=1.055 $Y=1.97
r109 99 104 0.0432039 $w=4.9e-07 $l=1.55e-07 $layer=MET1_cond $X=4.955 $Y=3.33
+ $X2=4.8 $Y2=3.33
r110 88 109 0.213232 $w=4.9e-07 $l=7.65e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=7.155 $Y2=3.33
r111 87 89 9.36939 $w=5.73e-07 $l=1.35e-07 $layer=LI1_cond $X=7.92 $Y=3.127
+ $X2=8.055 $Y2=3.127
r112 87 88 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r113 85 87 2.80818 $w=5.73e-07 $l=1.35e-07 $layer=LI1_cond $X=7.785 $Y=3.127
+ $X2=7.92 $Y2=3.127
r114 81 89 53.8235 $w=1.68e-07 $l=8.25e-07 $layer=LI1_cond $X=8.88 $Y=3.33
+ $X2=8.055 $Y2=3.33
r115 81 82 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r116 74 77 34.5733 $w=2.58e-07 $l=7.8e-07 $layer=LI1_cond $X=7.005 $Y=2.11
+ $X2=7.785 $Y2=2.11
r117 74 75 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.005 $Y=2.11
+ $X2=7.005 $Y2=2.11
r118 71 74 68.925 $w=2.58e-07 $l=1.555e-06 $layer=LI1_cond $X=5.45 $Y=2.11
+ $X2=7.005 $Y2=2.11
r119 71 72 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.45 $Y=2.11
+ $X2=5.45 $Y2=2.11
r120 68 71 68.925 $w=2.58e-07 $l=1.555e-06 $layer=LI1_cond $X=3.895 $Y=2.11
+ $X2=5.45 $Y2=2.11
r121 68 69 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.895 $Y=2.11
+ $X2=3.895 $Y2=2.11
r122 65 68 68.925 $w=2.58e-07 $l=1.555e-06 $layer=LI1_cond $X=2.34 $Y=2.11
+ $X2=3.895 $Y2=2.11
r123 65 66 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.34 $Y=2.11
+ $X2=2.34 $Y2=2.11
r124 62 65 44.9896 $w=2.58e-07 $l=1.015e-06 $layer=LI1_cond $X=1.325 $Y=2.11
+ $X2=2.34 $Y2=2.11
r125 60 75 0.175043 $w=6.45e-07 $l=8.6e-07 $layer=MET1_cond $X=6.832 $Y=2.97
+ $X2=6.832 $Y2=2.11
r126 59 60 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=7.005 $Y=2.97
+ $X2=7.005 $Y2=2.97
r127 57 105 0.00836204 $w=4.9e-07 $l=3e-08 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=6.51 $Y2=3.33
r128 56 59 10.9207 $w=5.73e-07 $l=5.25e-07 $layer=LI1_cond $X=6.48 $Y=3.127
+ $X2=7.005 $Y2=3.127
r129 56 57 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r130 53 56 19.9693 $w=5.73e-07 $l=9.6e-07 $layer=LI1_cond $X=5.52 $Y=3.127
+ $X2=6.48 $Y2=3.127
r131 51 72 0.180644 $w=6.25e-07 $l=8.6e-07 $layer=MET1_cond $X=5.267 $Y=2.97
+ $X2=5.267 $Y2=2.11
r132 50 53 1.4561 $w=5.73e-07 $l=7e-08 $layer=LI1_cond $X=5.45 $Y=3.127 $X2=5.52
+ $Y2=3.127
r133 50 51 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=5.45 $Y=2.97
+ $X2=5.45 $Y2=2.97
r134 48 104 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=4.8 $Y2=3.33
r135 47 50 18.5132 $w=5.73e-07 $l=8.9e-07 $layer=LI1_cond $X=4.56 $Y=3.127
+ $X2=5.45 $Y2=3.127
r136 47 48 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r137 45 69 0.180644 $w=6.25e-07 $l=8.6e-07 $layer=MET1_cond $X=3.712 $Y=2.97
+ $X2=3.712 $Y2=2.11
r138 44 47 13.8329 $w=5.73e-07 $l=6.65e-07 $layer=LI1_cond $X=3.895 $Y=3.127
+ $X2=4.56 $Y2=3.127
r139 44 45 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.895 $Y=2.97
+ $X2=3.895 $Y2=2.97
r140 42 95 0.0780457 $w=4.9e-07 $l=2.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.4 $Y2=3.33
r141 41 44 16.1211 $w=5.73e-07 $l=7.75e-07 $layer=LI1_cond $X=3.12 $Y=3.127
+ $X2=3.895 $Y2=3.127
r142 41 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r143 38 41 16.2251 $w=5.73e-07 $l=7.8e-07 $layer=LI1_cond $X=2.34 $Y=3.127
+ $X2=3.12 $Y2=3.127
r144 36 66 0.180644 $w=6.25e-07 $l=8.6e-07 $layer=MET1_cond $X=2.157 $Y=2.97
+ $X2=2.157 $Y2=2.11
r145 36 38 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.34 $Y=2.97
+ $X2=2.34 $Y2=2.97
r146 35 38 7.48849 $w=5.73e-07 $l=3.6e-07 $layer=LI1_cond $X=1.98 $Y=3.127
+ $X2=2.34 $Y2=3.127
r147 35 36 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.98 $Y=2.97
+ $X2=1.98 $Y2=2.97
r148 33 90 0.0459912 $w=4.9e-07 $l=1.65e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.845 $Y2=3.33
r149 32 35 6.24041 $w=5.73e-07 $l=3e-07 $layer=LI1_cond $X=1.68 $Y=3.127
+ $X2=1.98 $Y2=3.127
r150 32 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r151 30 85 0.353623 $w=5.73e-07 $l=1.7e-08 $layer=LI1_cond $X=7.768 $Y=3.127
+ $X2=7.785 $Y2=3.127
r152 30 59 15.8714 $w=5.73e-07 $l=7.63e-07 $layer=LI1_cond $X=7.768 $Y=3.127
+ $X2=7.005 $Y2=3.127
r153 27 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r154 12 105 0.0661031 $w=4.9e-07 $l=3.22e-07 $layer=MET1_cond $X=6.832 $Y=3.33
+ $X2=6.51 $Y2=3.33
r155 12 109 0.0661031 $w=4.9e-07 $l=3.23e-07 $layer=MET1_cond $X=6.832 $Y=3.33
+ $X2=7.155 $Y2=3.33
r156 12 99 0.0644858 $w=4.9e-07 $l=3.12e-07 $layer=MET1_cond $X=5.267 $Y=3.33
+ $X2=4.955 $Y2=3.33
r157 12 106 0.0644858 $w=4.9e-07 $l=3.13e-07 $layer=MET1_cond $X=5.267 $Y=3.33
+ $X2=5.58 $Y2=3.33
r158 12 95 0.0644858 $w=4.9e-07 $l=3.12e-07 $layer=MET1_cond $X=3.712 $Y=3.33
+ $X2=3.4 $Y2=3.33
r159 12 100 0.0644858 $w=4.9e-07 $l=3.13e-07 $layer=MET1_cond $X=3.712 $Y=3.33
+ $X2=4.025 $Y2=3.33
r160 12 90 0.0644858 $w=4.9e-07 $l=3.12e-07 $layer=MET1_cond $X=2.157 $Y=3.33
+ $X2=1.845 $Y2=3.33
r161 12 96 0.0644858 $w=4.9e-07 $l=3.13e-07 $layer=MET1_cond $X=2.157 $Y=3.33
+ $X2=2.47 $Y2=3.33
r162 12 60 0.044502 $w=1.29e-06 $l=1.15e-07 $layer=MET1_cond $X=6.832 $Y=3.085
+ $X2=6.832 $Y2=2.97
r163 12 51 0.0448765 $w=1.25e-06 $l=1.15e-07 $layer=MET1_cond $X=5.267 $Y=3.085
+ $X2=5.267 $Y2=2.97
r164 12 45 0.0448765 $w=1.25e-06 $l=1.15e-07 $layer=MET1_cond $X=3.712 $Y=3.085
+ $X2=3.712 $Y2=2.97
r165 12 36 0.0448765 $w=1.25e-06 $l=1.15e-07 $layer=MET1_cond $X=2.157 $Y=3.085
+ $X2=2.157 $Y2=2.97
r166 12 82 0.2071 $w=4.9e-07 $l=7.43e-07 $layer=MET1_cond $X=8.137 $Y=3.33
+ $X2=8.88 $Y2=3.33
r167 12 88 0.0604854 $w=4.9e-07 $l=2.17e-07 $layer=MET1_cond $X=8.137 $Y=3.33
+ $X2=7.92 $Y2=3.33
r168 12 57 0.12125 $w=4.9e-07 $l=4.35e-07 $layer=MET1_cond $X=6.045 $Y=3.33
+ $X2=6.48 $Y2=3.33
r169 12 106 0.129612 $w=4.9e-07 $l=4.65e-07 $layer=MET1_cond $X=6.045 $Y=3.33
+ $X2=5.58 $Y2=3.33
r170 12 48 0.0195114 $w=4.9e-07 $l=7e-08 $layer=MET1_cond $X=4.49 $Y=3.33
+ $X2=4.56 $Y2=3.33
r171 12 100 0.129612 $w=4.9e-07 $l=4.65e-07 $layer=MET1_cond $X=4.49 $Y=3.33
+ $X2=4.025 $Y2=3.33
r172 12 42 0.0515659 $w=4.9e-07 $l=1.85e-07 $layer=MET1_cond $X=2.935 $Y=3.33
+ $X2=3.12 $Y2=3.33
r173 12 96 0.129612 $w=4.9e-07 $l=4.65e-07 $layer=MET1_cond $X=2.935 $Y=3.33
+ $X2=2.47 $Y2=3.33
r174 12 33 0.211281 $w=4.9e-07 $l=7.58e-07 $layer=MET1_cond $X=0.922 $Y=3.33
+ $X2=1.68 $Y2=3.33
r175 12 28 0.0563044 $w=4.9e-07 $l=2.02e-07 $layer=MET1_cond $X=0.922 $Y=3.33
+ $X2=0.72 $Y2=3.33
r176 12 53 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r177 11 27 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.055 $Y=3.33
+ $X2=0.72 $Y2=3.33
r178 10 11 12.1776 $w=5.73e-07 $l=2.7e-07 $layer=LI1_cond $X=1.325 $Y=3.127
+ $X2=1.055 $Y2=3.127
r179 7 32 7.03086 $w=5.73e-07 $l=3.38e-07 $layer=LI1_cond $X=1.342 $Y=3.127
+ $X2=1.68 $Y2=3.127
r180 7 10 0.353623 $w=5.73e-07 $l=1.7e-08 $layer=LI1_cond $X=1.342 $Y=3.127
+ $X2=1.325 $Y2=3.127
r181 2 85 60 $w=1.7e-07 $l=6.79964e-06 $layer=licon1_PDIFF $count=10 $X=1.055
+ $Y=2.83 $X2=7.785 $Y2=2.97
r182 2 10 60 $w=1.7e-07 $l=3.32716e-07 $layer=licon1_PDIFF $count=10 $X=1.055
+ $Y=2.83 $X2=1.325 $Y2=2.97
r183 1 77 60 $w=1.7e-07 $l=6.79964e-06 $layer=licon1_PDIFF $count=10 $X=1.055
+ $Y=1.97 $X2=7.785 $Y2=2.11
r184 1 62 60 $w=1.7e-07 $l=3.32716e-07 $layer=licon1_PDIFF $count=10 $X=1.055
+ $Y=1.97 $X2=1.325 $Y2=2.11
.ends

