* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__nor4bb_1 A B C_N D_N VGND VNB VPB VPWR Y
X0 a_513_367# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X1 VGND a_27_508# Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X2 VGND B Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X3 a_405_367# B a_513_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X4 a_333_367# a_375_269# a_405_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X5 Y A VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X6 a_27_508# D_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X7 VGND C_N a_375_269# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 VPWR C_N a_375_269# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X9 Y a_27_508# a_333_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X10 Y a_375_269# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X11 a_27_508# D_N VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
