* File: sky130_fd_sc_lp__o2bb2ai_2.pxi.spice
* Created: Wed Sep  2 10:22:17 2020
* 
x_PM_SKY130_FD_SC_LP__O2BB2AI_2%A1_N N_A1_N_M1015_g N_A1_N_M1001_g
+ N_A1_N_M1017_g N_A1_N_M1007_g N_A1_N_c_113_p N_A1_N_c_101_n N_A1_N_c_102_n
+ A1_N N_A1_N_c_103_n N_A1_N_c_104_n N_A1_N_c_105_n
+ PM_SKY130_FD_SC_LP__O2BB2AI_2%A1_N
x_PM_SKY130_FD_SC_LP__O2BB2AI_2%A2_N N_A2_N_c_183_n N_A2_N_M1008_g
+ N_A2_N_M1009_g N_A2_N_c_185_n N_A2_N_M1018_g N_A2_N_M1014_g A2_N A2_N
+ N_A2_N_c_188_n PM_SKY130_FD_SC_LP__O2BB2AI_2%A2_N
x_PM_SKY130_FD_SC_LP__O2BB2AI_2%A_125_367# N_A_125_367#_M1008_s
+ N_A_125_367#_M1001_s N_A_125_367#_M1014_d N_A_125_367#_c_233_n
+ N_A_125_367#_c_234_n N_A_125_367#_M1000_g N_A_125_367#_M1004_g
+ N_A_125_367#_c_236_n N_A_125_367#_c_237_n N_A_125_367#_M1006_g
+ N_A_125_367#_M1019_g N_A_125_367#_c_239_n N_A_125_367#_c_240_n
+ N_A_125_367#_c_253_n N_A_125_367#_c_241_n N_A_125_367#_c_303_p
+ N_A_125_367#_c_257_n N_A_125_367#_c_242_n N_A_125_367#_c_243_n
+ N_A_125_367#_c_266_n N_A_125_367#_c_268_n N_A_125_367#_c_244_n
+ N_A_125_367#_c_245_n PM_SKY130_FD_SC_LP__O2BB2AI_2%A_125_367#
x_PM_SKY130_FD_SC_LP__O2BB2AI_2%B1 N_B1_M1011_g N_B1_M1012_g N_B1_c_343_n
+ N_B1_M1016_g N_B1_M1013_g N_B1_c_345_n N_B1_c_346_n N_B1_c_347_n N_B1_c_354_n
+ N_B1_c_361_n B1 N_B1_c_348_n N_B1_c_349_n PM_SKY130_FD_SC_LP__O2BB2AI_2%B1
x_PM_SKY130_FD_SC_LP__O2BB2AI_2%B2 N_B2_M1002_g N_B2_c_427_n N_B2_M1003_g
+ N_B2_c_428_n N_B2_M1010_g N_B2_M1005_g B2 B2 B2 N_B2_c_431_n
+ PM_SKY130_FD_SC_LP__O2BB2AI_2%B2
x_PM_SKY130_FD_SC_LP__O2BB2AI_2%VPWR N_VPWR_M1001_d N_VPWR_M1009_s
+ N_VPWR_M1007_d N_VPWR_M1019_s N_VPWR_M1013_d N_VPWR_c_483_n N_VPWR_c_484_n
+ N_VPWR_c_485_n N_VPWR_c_486_n N_VPWR_c_487_n N_VPWR_c_488_n N_VPWR_c_489_n
+ N_VPWR_c_490_n N_VPWR_c_491_n VPWR N_VPWR_c_492_n N_VPWR_c_493_n
+ N_VPWR_c_482_n N_VPWR_c_495_n N_VPWR_c_496_n N_VPWR_c_497_n N_VPWR_c_498_n
+ PM_SKY130_FD_SC_LP__O2BB2AI_2%VPWR
x_PM_SKY130_FD_SC_LP__O2BB2AI_2%Y N_Y_M1000_d N_Y_M1004_d N_Y_M1002_s
+ N_Y_c_576_n Y Y Y Y Y Y N_Y_c_581_n PM_SKY130_FD_SC_LP__O2BB2AI_2%Y
x_PM_SKY130_FD_SC_LP__O2BB2AI_2%A_765_367# N_A_765_367#_M1011_s
+ N_A_765_367#_M1005_d N_A_765_367#_c_621_n N_A_765_367#_c_623_n
+ PM_SKY130_FD_SC_LP__O2BB2AI_2%A_765_367#
x_PM_SKY130_FD_SC_LP__O2BB2AI_2%VGND N_VGND_M1015_d N_VGND_M1017_d
+ N_VGND_M1012_d N_VGND_M1010_s N_VGND_c_635_n N_VGND_c_636_n N_VGND_c_637_n
+ N_VGND_c_638_n N_VGND_c_639_n N_VGND_c_640_n N_VGND_c_641_n VGND
+ N_VGND_c_642_n N_VGND_c_643_n N_VGND_c_644_n N_VGND_c_645_n N_VGND_c_646_n
+ N_VGND_c_647_n PM_SKY130_FD_SC_LP__O2BB2AI_2%VGND
x_PM_SKY130_FD_SC_LP__O2BB2AI_2%A_125_69# N_A_125_69#_M1015_s
+ N_A_125_69#_M1018_d N_A_125_69#_c_708_n N_A_125_69#_c_711_n
+ N_A_125_69#_c_709_n PM_SKY130_FD_SC_LP__O2BB2AI_2%A_125_69#
x_PM_SKY130_FD_SC_LP__O2BB2AI_2%A_502_69# N_A_502_69#_M1000_s
+ N_A_502_69#_M1006_s N_A_502_69#_M1003_d N_A_502_69#_M1016_s
+ N_A_502_69#_c_725_n N_A_502_69#_c_726_n N_A_502_69#_c_727_n
+ N_A_502_69#_c_741_n N_A_502_69#_c_743_n N_A_502_69#_c_728_n
+ N_A_502_69#_c_729_n N_A_502_69#_c_730_n N_A_502_69#_c_755_n
+ PM_SKY130_FD_SC_LP__O2BB2AI_2%A_502_69#
cc_1 VNB N_A1_N_M1015_g 0.0251081f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=0.765
cc_2 VNB N_A1_N_M1007_g 0.00167964f $X=-0.19 $Y=-0.245 $X2=1.84 $Y2=2.465
cc_3 VNB N_A1_N_c_101_n 0.00226717f $X=-0.19 $Y=-0.245 $X2=1.86 $Y2=1.46
cc_4 VNB N_A1_N_c_102_n 0.0327391f $X=-0.19 $Y=-0.245 $X2=1.86 $Y2=1.46
cc_5 VNB N_A1_N_c_103_n 0.0289656f $X=-0.19 $Y=-0.245 $X2=0.46 $Y2=1.51
cc_6 VNB N_A1_N_c_104_n 0.0208031f $X=-0.19 $Y=-0.245 $X2=0.46 $Y2=1.51
cc_7 VNB N_A1_N_c_105_n 0.0194157f $X=-0.19 $Y=-0.245 $X2=1.86 $Y2=1.295
cc_8 VNB N_A2_N_c_183_n 0.0165934f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=1.345
cc_9 VNB N_A2_N_M1009_g 0.00139356f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=2.465
cc_10 VNB N_A2_N_c_185_n 0.0165929f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A2_N_M1014_g 0.00139629f $X=-0.19 $Y=-0.245 $X2=1.84 $Y2=2.465
cc_12 VNB A2_N 0.00261899f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A2_N_c_188_n 0.0380555f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_125_367#_c_233_n 0.0152293f $X=-0.19 $Y=-0.245 $X2=1.84 $Y2=0.765
cc_15 VNB N_A_125_367#_c_234_n 0.0187492f $X=-0.19 $Y=-0.245 $X2=1.84 $Y2=1.625
cc_16 VNB N_A_125_367#_M1004_g 0.00945531f $X=-0.19 $Y=-0.245 $X2=0.805
+ $Y2=2.005
cc_17 VNB N_A_125_367#_c_236_n 0.0101534f $X=-0.19 $Y=-0.245 $X2=1.852 $Y2=1.46
cc_18 VNB N_A_125_367#_c_237_n 0.0166736f $X=-0.19 $Y=-0.245 $X2=1.86 $Y2=1.46
cc_19 VNB N_A_125_367#_M1019_g 0.00948431f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_125_367#_c_239_n 0.0023879f $X=-0.19 $Y=-0.245 $X2=0.46 $Y2=1.51
cc_21 VNB N_A_125_367#_c_240_n 0.00523885f $X=-0.19 $Y=-0.245 $X2=0.46 $Y2=1.51
cc_22 VNB N_A_125_367#_c_241_n 0.00569718f $X=-0.19 $Y=-0.245 $X2=1.86 $Y2=1.625
cc_23 VNB N_A_125_367#_c_242_n 0.00580866f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_125_367#_c_243_n 6.63536e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_125_367#_c_244_n 0.00320857f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_125_367#_c_245_n 0.0428654f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_B1_M1012_g 0.0203481f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=2.465
cc_28 VNB N_B1_c_343_n 0.0208765f $X=-0.19 $Y=-0.245 $X2=1.84 $Y2=1.295
cc_29 VNB N_B1_M1013_g 0.00167964f $X=-0.19 $Y=-0.245 $X2=1.84 $Y2=2.465
cc_30 VNB N_B1_c_345_n 0.00892116f $X=-0.19 $Y=-0.245 $X2=0.805 $Y2=2.005
cc_31 VNB N_B1_c_346_n 0.00175536f $X=-0.19 $Y=-0.245 $X2=1.86 $Y2=1.46
cc_32 VNB N_B1_c_347_n 0.0262028f $X=-0.19 $Y=-0.245 $X2=1.86 $Y2=1.46
cc_33 VNB N_B1_c_348_n 0.0544889f $X=-0.19 $Y=-0.245 $X2=0.46 $Y2=1.51
cc_34 VNB N_B1_c_349_n 0.0238734f $X=-0.19 $Y=-0.245 $X2=0.46 $Y2=1.345
cc_35 VNB N_B2_M1002_g 0.00118886f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=0.765
cc_36 VNB N_B2_c_427_n 0.0157642f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=1.675
cc_37 VNB N_B2_c_428_n 0.0157642f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_B2_M1005_g 0.00128054f $X=-0.19 $Y=-0.245 $X2=1.84 $Y2=2.465
cc_39 VNB B2 0.0136759f $X=-0.19 $Y=-0.245 $X2=1.852 $Y2=1.46
cc_40 VNB N_B2_c_431_n 0.041414f $X=-0.19 $Y=-0.245 $X2=1.86 $Y2=1.295
cc_41 VNB N_VPWR_c_482_n 0.243291f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_635_n 0.0134903f $X=-0.19 $Y=-0.245 $X2=1.84 $Y2=2.465
cc_43 VNB N_VGND_c_636_n 0.0469788f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_637_n 0.00951602f $X=-0.19 $Y=-0.245 $X2=1.852 $Y2=1.46
cc_45 VNB N_VGND_c_638_n 0.00270988f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_46 VNB N_VGND_c_639_n 0.00270988f $X=-0.19 $Y=-0.245 $X2=0.46 $Y2=1.51
cc_47 VNB N_VGND_c_640_n 0.0146145f $X=-0.19 $Y=-0.245 $X2=0.46 $Y2=1.345
cc_48 VNB N_VGND_c_641_n 0.00573719f $X=-0.19 $Y=-0.245 $X2=0.46 $Y2=1.675
cc_49 VNB N_VGND_c_642_n 0.0355699f $X=-0.19 $Y=-0.245 $X2=1.86 $Y2=1.625
cc_50 VNB N_VGND_c_643_n 0.0400809f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_644_n 0.0229341f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_645_n 0.33141f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_646_n 0.00596836f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_647_n 0.00573719f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_125_69#_c_708_n 0.00205439f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=2.465
cc_56 VNB N_A_125_69#_c_709_n 0.00461081f $X=-0.19 $Y=-0.245 $X2=1.84 $Y2=2.465
cc_57 VNB N_A_502_69#_c_725_n 0.00216574f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_502_69#_c_726_n 0.00552922f $X=-0.19 $Y=-0.245 $X2=0.805 $Y2=2.005
cc_59 VNB N_A_502_69#_c_727_n 0.00262397f $X=-0.19 $Y=-0.245 $X2=1.852 $Y2=1.92
cc_60 VNB N_A_502_69#_c_728_n 0.00189378f $X=-0.19 $Y=-0.245 $X2=0.46 $Y2=1.51
cc_61 VNB N_A_502_69#_c_729_n 0.00746084f $X=-0.19 $Y=-0.245 $X2=0.46 $Y2=1.51
cc_62 VNB N_A_502_69#_c_730_n 0.0228642f $X=-0.19 $Y=-0.245 $X2=1.86 $Y2=1.295
cc_63 VPB N_A1_N_M1001_g 0.0216476f $X=-0.19 $Y=1.655 $X2=0.55 $Y2=2.465
cc_64 VPB N_A1_N_M1007_g 0.0237302f $X=-0.19 $Y=1.655 $X2=1.84 $Y2=2.465
cc_65 VPB N_A1_N_c_101_n 0.00323442f $X=-0.19 $Y=1.655 $X2=1.86 $Y2=1.46
cc_66 VPB N_A1_N_c_103_n 0.00668482f $X=-0.19 $Y=1.655 $X2=0.46 $Y2=1.51
cc_67 VPB N_A1_N_c_104_n 0.0244981f $X=-0.19 $Y=1.655 $X2=0.46 $Y2=1.51
cc_68 VPB N_A2_N_M1009_g 0.01952f $X=-0.19 $Y=1.655 $X2=0.55 $Y2=2.465
cc_69 VPB N_A2_N_M1014_g 0.0195354f $X=-0.19 $Y=1.655 $X2=1.84 $Y2=2.465
cc_70 VPB A2_N 0.00261899f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_71 VPB N_A_125_367#_M1004_g 0.0232544f $X=-0.19 $Y=1.655 $X2=0.805 $Y2=2.005
cc_72 VPB N_A_125_367#_M1019_g 0.0197381f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_73 VPB N_A_125_367#_c_243_n 0.00317291f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_74 VPB N_B1_M1011_g 0.0188701f $X=-0.19 $Y=1.655 $X2=0.55 $Y2=0.765
cc_75 VPB N_B1_M1013_g 0.0228758f $X=-0.19 $Y=1.655 $X2=1.84 $Y2=2.465
cc_76 VPB N_B1_c_346_n 0.00124473f $X=-0.19 $Y=1.655 $X2=1.86 $Y2=1.46
cc_77 VPB N_B1_c_347_n 0.00633982f $X=-0.19 $Y=1.655 $X2=1.86 $Y2=1.46
cc_78 VPB N_B1_c_354_n 0.0176489f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_79 VPB N_B1_c_349_n 0.0125481f $X=-0.19 $Y=1.655 $X2=0.46 $Y2=1.345
cc_80 VPB N_B2_M1002_g 0.0196555f $X=-0.19 $Y=1.655 $X2=0.55 $Y2=0.765
cc_81 VPB N_B2_M1005_g 0.0197305f $X=-0.19 $Y=1.655 $X2=1.84 $Y2=2.465
cc_82 VPB B2 0.00812039f $X=-0.19 $Y=1.655 $X2=1.852 $Y2=1.46
cc_83 VPB N_VPWR_c_483_n 0.0127321f $X=-0.19 $Y=1.655 $X2=1.695 $Y2=2.005
cc_84 VPB N_VPWR_c_484_n 0.0348213f $X=-0.19 $Y=1.655 $X2=1.852 $Y2=1.92
cc_85 VPB N_VPWR_c_485_n 3.15043e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_86 VPB N_VPWR_c_486_n 0.0025093f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_87 VPB N_VPWR_c_487_n 0.00443685f $X=-0.19 $Y=1.655 $X2=0.46 $Y2=1.345
cc_88 VPB N_VPWR_c_488_n 0.0352283f $X=-0.19 $Y=1.655 $X2=1.86 $Y2=1.625
cc_89 VPB N_VPWR_c_489_n 0.0116899f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_90 VPB N_VPWR_c_490_n 0.0348216f $X=-0.19 $Y=1.655 $X2=0.445 $Y2=1.665
cc_91 VPB N_VPWR_c_491_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_92 VPB N_VPWR_c_492_n 0.0129398f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_93 VPB N_VPWR_c_493_n 0.0173273f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_94 VPB N_VPWR_c_482_n 0.0554576f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_95 VPB N_VPWR_c_495_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_96 VPB N_VPWR_c_496_n 0.0147711f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_97 VPB N_VPWR_c_497_n 0.0225077f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_98 VPB N_VPWR_c_498_n 0.00439057f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_99 N_A1_N_M1015_g N_A2_N_c_183_n 0.02258f $X=0.55 $Y=0.765 $X2=-0.19
+ $Y2=-0.245
cc_100 N_A1_N_M1001_g N_A2_N_M1009_g 0.02258f $X=0.55 $Y=2.465 $X2=0 $Y2=0
cc_101 N_A1_N_c_113_p N_A2_N_M1009_g 0.0119819f $X=1.695 $Y=2.005 $X2=0 $Y2=0
cc_102 N_A1_N_c_104_n N_A2_N_M1009_g 2.38631e-19 $X=0.46 $Y=1.51 $X2=0 $Y2=0
cc_103 N_A1_N_c_105_n N_A2_N_c_185_n 0.0341037f $X=1.86 $Y=1.295 $X2=0 $Y2=0
cc_104 N_A1_N_M1007_g N_A2_N_M1014_g 0.0351988f $X=1.84 $Y=2.465 $X2=0 $Y2=0
cc_105 N_A1_N_c_113_p N_A2_N_M1014_g 0.0113413f $X=1.695 $Y=2.005 $X2=0 $Y2=0
cc_106 N_A1_N_c_101_n N_A2_N_M1014_g 0.00454413f $X=1.86 $Y=1.46 $X2=0 $Y2=0
cc_107 N_A1_N_M1015_g A2_N 8.8105e-19 $X=0.55 $Y=0.765 $X2=0 $Y2=0
cc_108 N_A1_N_c_113_p A2_N 0.0327208f $X=1.695 $Y=2.005 $X2=0 $Y2=0
cc_109 N_A1_N_c_101_n A2_N 0.0270443f $X=1.86 $Y=1.46 $X2=0 $Y2=0
cc_110 N_A1_N_c_102_n A2_N 0.00109715f $X=1.86 $Y=1.46 $X2=0 $Y2=0
cc_111 N_A1_N_c_103_n A2_N 3.14592e-19 $X=0.46 $Y=1.51 $X2=0 $Y2=0
cc_112 N_A1_N_c_104_n A2_N 0.0310094f $X=0.46 $Y=1.51 $X2=0 $Y2=0
cc_113 N_A1_N_c_105_n A2_N 4.91346e-19 $X=1.86 $Y=1.295 $X2=0 $Y2=0
cc_114 N_A1_N_c_113_p N_A2_N_c_188_n 5.14635e-19 $X=1.695 $Y=2.005 $X2=0 $Y2=0
cc_115 N_A1_N_c_101_n N_A2_N_c_188_n 0.00130569f $X=1.86 $Y=1.46 $X2=0 $Y2=0
cc_116 N_A1_N_c_102_n N_A2_N_c_188_n 0.021113f $X=1.86 $Y=1.46 $X2=0 $Y2=0
cc_117 N_A1_N_c_103_n N_A2_N_c_188_n 0.02258f $X=0.46 $Y=1.51 $X2=0 $Y2=0
cc_118 N_A1_N_c_104_n N_A2_N_c_188_n 0.00828688f $X=0.46 $Y=1.51 $X2=0 $Y2=0
cc_119 N_A1_N_c_113_p N_A_125_367#_M1001_s 0.00250501f $X=1.695 $Y=2.005 $X2=0
+ $Y2=0
cc_120 N_A1_N_c_104_n N_A_125_367#_M1001_s 0.00289273f $X=0.46 $Y=1.51 $X2=0
+ $Y2=0
cc_121 N_A1_N_c_113_p N_A_125_367#_M1014_d 0.00754823f $X=1.695 $Y=2.005 $X2=0
+ $Y2=0
cc_122 N_A1_N_c_101_n N_A_125_367#_M1014_d 0.00107999f $X=1.86 $Y=1.46 $X2=0
+ $Y2=0
cc_123 N_A1_N_c_113_p N_A_125_367#_c_253_n 0.0323235f $X=1.695 $Y=2.005 $X2=0
+ $Y2=0
cc_124 N_A1_N_c_101_n N_A_125_367#_c_241_n 0.014698f $X=1.86 $Y=1.46 $X2=0 $Y2=0
cc_125 N_A1_N_c_102_n N_A_125_367#_c_241_n 0.00131694f $X=1.86 $Y=1.46 $X2=0
+ $Y2=0
cc_126 N_A1_N_c_105_n N_A_125_367#_c_241_n 0.0157763f $X=1.86 $Y=1.295 $X2=0
+ $Y2=0
cc_127 N_A1_N_M1007_g N_A_125_367#_c_257_n 0.0154716f $X=1.84 $Y=2.465 $X2=0
+ $Y2=0
cc_128 N_A1_N_c_113_p N_A_125_367#_c_257_n 0.0145499f $X=1.695 $Y=2.005 $X2=0
+ $Y2=0
cc_129 N_A1_N_c_102_n N_A_125_367#_c_257_n 5.73398e-19 $X=1.86 $Y=1.46 $X2=0
+ $Y2=0
cc_130 N_A1_N_c_101_n N_A_125_367#_c_242_n 0.0059911f $X=1.86 $Y=1.46 $X2=0
+ $Y2=0
cc_131 N_A1_N_c_102_n N_A_125_367#_c_242_n 4.34657e-19 $X=1.86 $Y=1.46 $X2=0
+ $Y2=0
cc_132 N_A1_N_c_105_n N_A_125_367#_c_242_n 0.0078543f $X=1.86 $Y=1.295 $X2=0
+ $Y2=0
cc_133 N_A1_N_M1007_g N_A_125_367#_c_243_n 0.00784643f $X=1.84 $Y=2.465 $X2=0
+ $Y2=0
cc_134 N_A1_N_c_113_p N_A_125_367#_c_243_n 0.0138309f $X=1.695 $Y=2.005 $X2=0
+ $Y2=0
cc_135 N_A1_N_c_101_n N_A_125_367#_c_243_n 0.0230194f $X=1.86 $Y=1.46 $X2=0
+ $Y2=0
cc_136 N_A1_N_c_113_p N_A_125_367#_c_266_n 0.00349842f $X=1.695 $Y=2.005 $X2=0
+ $Y2=0
cc_137 N_A1_N_c_104_n N_A_125_367#_c_266_n 0.0110408f $X=0.46 $Y=1.51 $X2=0
+ $Y2=0
cc_138 N_A1_N_c_113_p N_A_125_367#_c_268_n 0.0135384f $X=1.695 $Y=2.005 $X2=0
+ $Y2=0
cc_139 N_A1_N_c_101_n N_A_125_367#_c_244_n 0.0198998f $X=1.86 $Y=1.46 $X2=0
+ $Y2=0
cc_140 N_A1_N_c_102_n N_A_125_367#_c_244_n 0.00146344f $X=1.86 $Y=1.46 $X2=0
+ $Y2=0
cc_141 N_A1_N_c_101_n N_A_125_367#_c_245_n 3.55515e-19 $X=1.86 $Y=1.46 $X2=0
+ $Y2=0
cc_142 N_A1_N_c_102_n N_A_125_367#_c_245_n 0.0206497f $X=1.86 $Y=1.46 $X2=0
+ $Y2=0
cc_143 N_A1_N_c_104_n N_VPWR_M1001_d 0.00346745f $X=0.46 $Y=1.51 $X2=-0.19
+ $Y2=-0.245
cc_144 N_A1_N_c_113_p N_VPWR_M1009_s 0.0033464f $X=1.695 $Y=2.005 $X2=0 $Y2=0
cc_145 N_A1_N_c_113_p N_VPWR_M1007_d 0.00229635f $X=1.695 $Y=2.005 $X2=0 $Y2=0
cc_146 N_A1_N_c_101_n N_VPWR_M1007_d 9.12275e-19 $X=1.86 $Y=1.46 $X2=0 $Y2=0
cc_147 N_A1_N_M1001_g N_VPWR_c_484_n 0.0172637f $X=0.55 $Y=2.465 $X2=0 $Y2=0
cc_148 N_A1_N_c_103_n N_VPWR_c_484_n 5.32653e-19 $X=0.46 $Y=1.51 $X2=0 $Y2=0
cc_149 N_A1_N_c_104_n N_VPWR_c_484_n 0.0234591f $X=0.46 $Y=1.51 $X2=0 $Y2=0
cc_150 N_A1_N_M1001_g N_VPWR_c_485_n 5.84303e-19 $X=0.55 $Y=2.465 $X2=0 $Y2=0
cc_151 N_A1_N_M1007_g N_VPWR_c_485_n 5.9812e-19 $X=1.84 $Y=2.465 $X2=0 $Y2=0
cc_152 N_A1_N_M1007_g N_VPWR_c_486_n 0.00424227f $X=1.84 $Y=2.465 $X2=0 $Y2=0
cc_153 N_A1_N_M1001_g N_VPWR_c_492_n 0.00486043f $X=0.55 $Y=2.465 $X2=0 $Y2=0
cc_154 N_A1_N_M1001_g N_VPWR_c_482_n 0.0082726f $X=0.55 $Y=2.465 $X2=0 $Y2=0
cc_155 N_A1_N_M1007_g N_VPWR_c_482_n 0.0120521f $X=1.84 $Y=2.465 $X2=0 $Y2=0
cc_156 N_A1_N_M1007_g N_VPWR_c_496_n 0.00585385f $X=1.84 $Y=2.465 $X2=0 $Y2=0
cc_157 N_A1_N_M1007_g N_VPWR_c_497_n 0.00581385f $X=1.84 $Y=2.465 $X2=0 $Y2=0
cc_158 N_A1_N_M1015_g N_VGND_c_636_n 0.00882391f $X=0.55 $Y=0.765 $X2=0 $Y2=0
cc_159 N_A1_N_c_103_n N_VGND_c_636_n 0.0043204f $X=0.46 $Y=1.51 $X2=0 $Y2=0
cc_160 N_A1_N_c_104_n N_VGND_c_636_n 0.0276786f $X=0.46 $Y=1.51 $X2=0 $Y2=0
cc_161 N_A1_N_c_105_n N_VGND_c_637_n 0.00883307f $X=1.86 $Y=1.295 $X2=0 $Y2=0
cc_162 N_A1_N_M1015_g N_VGND_c_642_n 0.00480781f $X=0.55 $Y=0.765 $X2=0 $Y2=0
cc_163 N_A1_N_c_105_n N_VGND_c_642_n 0.00400407f $X=1.86 $Y=1.295 $X2=0 $Y2=0
cc_164 N_A1_N_M1015_g N_VGND_c_645_n 0.00964789f $X=0.55 $Y=0.765 $X2=0 $Y2=0
cc_165 N_A1_N_c_105_n N_VGND_c_645_n 0.00399422f $X=1.86 $Y=1.295 $X2=0 $Y2=0
cc_166 N_A1_N_M1015_g N_A_125_69#_c_708_n 3.43767e-19 $X=0.55 $Y=0.765 $X2=0
+ $Y2=0
cc_167 N_A1_N_c_104_n N_A_125_69#_c_711_n 0.00893916f $X=0.46 $Y=1.51 $X2=0
+ $Y2=0
cc_168 N_A1_N_c_105_n N_A_125_69#_c_709_n 3.19063e-19 $X=1.86 $Y=1.295 $X2=0
+ $Y2=0
cc_169 N_A1_N_c_105_n N_A_502_69#_c_725_n 0.00386652f $X=1.86 $Y=1.295 $X2=0
+ $Y2=0
cc_170 N_A1_N_c_105_n N_A_502_69#_c_727_n 5.76893e-19 $X=1.86 $Y=1.295 $X2=0
+ $Y2=0
cc_171 N_A2_N_M1009_g N_A_125_367#_c_253_n 0.0122595f $X=0.98 $Y=2.465 $X2=0
+ $Y2=0
cc_172 N_A2_N_M1014_g N_A_125_367#_c_253_n 0.0122129f $X=1.41 $Y=2.465 $X2=0
+ $Y2=0
cc_173 N_A2_N_c_183_n N_A_125_367#_c_241_n 0.00277239f $X=0.98 $Y=1.295 $X2=0
+ $Y2=0
cc_174 N_A2_N_c_185_n N_A_125_367#_c_241_n 0.0104276f $X=1.41 $Y=1.295 $X2=0
+ $Y2=0
cc_175 A2_N N_A_125_367#_c_241_n 0.0297194f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_176 N_A2_N_c_188_n N_A_125_367#_c_241_n 5.72878e-19 $X=1.41 $Y=1.46 $X2=0
+ $Y2=0
cc_177 N_A2_N_M1009_g N_VPWR_c_484_n 6.32678e-19 $X=0.98 $Y=2.465 $X2=0 $Y2=0
cc_178 N_A2_N_M1009_g N_VPWR_c_485_n 0.0112346f $X=0.98 $Y=2.465 $X2=0 $Y2=0
cc_179 N_A2_N_M1014_g N_VPWR_c_485_n 0.0113129f $X=1.41 $Y=2.465 $X2=0 $Y2=0
cc_180 N_A2_N_M1009_g N_VPWR_c_492_n 0.00486043f $X=0.98 $Y=2.465 $X2=0 $Y2=0
cc_181 N_A2_N_M1009_g N_VPWR_c_482_n 0.0082726f $X=0.98 $Y=2.465 $X2=0 $Y2=0
cc_182 N_A2_N_M1014_g N_VPWR_c_482_n 0.0082726f $X=1.41 $Y=2.465 $X2=0 $Y2=0
cc_183 N_A2_N_M1014_g N_VPWR_c_496_n 0.00486043f $X=1.41 $Y=2.465 $X2=0 $Y2=0
cc_184 N_A2_N_c_185_n N_VGND_c_637_n 6.51314e-19 $X=1.41 $Y=1.295 $X2=0 $Y2=0
cc_185 N_A2_N_c_183_n N_VGND_c_642_n 0.0029912f $X=0.98 $Y=1.295 $X2=0 $Y2=0
cc_186 N_A2_N_c_185_n N_VGND_c_642_n 0.0029912f $X=1.41 $Y=1.295 $X2=0 $Y2=0
cc_187 N_A2_N_c_183_n N_VGND_c_645_n 0.00401096f $X=0.98 $Y=1.295 $X2=0 $Y2=0
cc_188 N_A2_N_c_185_n N_VGND_c_645_n 0.00401096f $X=1.41 $Y=1.295 $X2=0 $Y2=0
cc_189 N_A2_N_c_183_n N_A_125_69#_c_709_n 0.0160837f $X=0.98 $Y=1.295 $X2=0
+ $Y2=0
cc_190 N_A2_N_c_185_n N_A_125_69#_c_709_n 0.0127734f $X=1.41 $Y=1.295 $X2=0
+ $Y2=0
cc_191 A2_N N_A_125_69#_c_709_n 0.00131813f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_192 N_A_125_367#_M1019_g N_B1_M1011_g 0.0446345f $X=3.28 $Y=2.465 $X2=0 $Y2=0
cc_193 N_A_125_367#_c_237_n N_B1_M1012_g 0.013726f $X=3.28 $Y=1.295 $X2=0 $Y2=0
cc_194 N_A_125_367#_M1019_g N_B1_c_346_n 0.00185009f $X=3.28 $Y=2.465 $X2=0
+ $Y2=0
cc_195 N_A_125_367#_c_240_n N_B1_c_346_n 0.00120569f $X=3.28 $Y=1.37 $X2=0 $Y2=0
cc_196 N_A_125_367#_c_240_n N_B1_c_347_n 0.0201462f $X=3.28 $Y=1.37 $X2=0 $Y2=0
cc_197 N_A_125_367#_M1019_g N_B1_c_361_n 0.00147829f $X=3.28 $Y=2.465 $X2=0
+ $Y2=0
cc_198 N_A_125_367#_c_253_n N_VPWR_M1009_s 0.0034506f $X=1.53 $Y=2.345 $X2=0
+ $Y2=0
cc_199 N_A_125_367#_c_257_n N_VPWR_M1007_d 0.0151467f $X=2.18 $Y=2.355 $X2=0
+ $Y2=0
cc_200 N_A_125_367#_c_243_n N_VPWR_M1007_d 0.0121568f $X=2.265 $Y=2.26 $X2=0
+ $Y2=0
cc_201 N_A_125_367#_c_253_n N_VPWR_c_485_n 0.0170777f $X=1.53 $Y=2.345 $X2=0
+ $Y2=0
cc_202 N_A_125_367#_c_233_n N_VPWR_c_486_n 0.00329096f $X=2.775 $Y=1.37 $X2=0
+ $Y2=0
cc_203 N_A_125_367#_M1004_g N_VPWR_c_486_n 0.00286486f $X=2.85 $Y=2.465 $X2=0
+ $Y2=0
cc_204 N_A_125_367#_c_257_n N_VPWR_c_486_n 0.0156812f $X=2.18 $Y=2.355 $X2=0
+ $Y2=0
cc_205 N_A_125_367#_c_243_n N_VPWR_c_486_n 0.0328601f $X=2.265 $Y=2.26 $X2=0
+ $Y2=0
cc_206 N_A_125_367#_c_244_n N_VPWR_c_486_n 0.00334988f $X=2.4 $Y=1.46 $X2=0
+ $Y2=0
cc_207 N_A_125_367#_c_245_n N_VPWR_c_486_n 0.00101476f $X=2.4 $Y=1.37 $X2=0
+ $Y2=0
cc_208 N_A_125_367#_M1019_g N_VPWR_c_487_n 0.00161646f $X=3.28 $Y=2.465 $X2=0
+ $Y2=0
cc_209 N_A_125_367#_c_266_n N_VPWR_c_492_n 0.0124525f $X=0.765 $Y=2.425 $X2=0
+ $Y2=0
cc_210 N_A_125_367#_M1004_g N_VPWR_c_493_n 0.0054895f $X=2.85 $Y=2.465 $X2=0
+ $Y2=0
cc_211 N_A_125_367#_M1019_g N_VPWR_c_493_n 0.00427694f $X=3.28 $Y=2.465 $X2=0
+ $Y2=0
cc_212 N_A_125_367#_M1001_s N_VPWR_c_482_n 0.00536646f $X=0.625 $Y=1.835 $X2=0
+ $Y2=0
cc_213 N_A_125_367#_M1014_d N_VPWR_c_482_n 0.0041489f $X=1.485 $Y=1.835 $X2=0
+ $Y2=0
cc_214 N_A_125_367#_M1004_g N_VPWR_c_482_n 0.0110627f $X=2.85 $Y=2.465 $X2=0
+ $Y2=0
cc_215 N_A_125_367#_M1019_g N_VPWR_c_482_n 0.00595547f $X=3.28 $Y=2.465 $X2=0
+ $Y2=0
cc_216 N_A_125_367#_c_303_p N_VPWR_c_482_n 0.00866972f $X=1.625 $Y=2.91 $X2=0
+ $Y2=0
cc_217 N_A_125_367#_c_266_n N_VPWR_c_482_n 0.00730901f $X=0.765 $Y=2.425 $X2=0
+ $Y2=0
cc_218 N_A_125_367#_c_303_p N_VPWR_c_496_n 0.0136943f $X=1.625 $Y=2.91 $X2=0
+ $Y2=0
cc_219 N_A_125_367#_M1004_g N_VPWR_c_497_n 0.00507123f $X=2.85 $Y=2.465 $X2=0
+ $Y2=0
cc_220 N_A_125_367#_c_257_n N_VPWR_c_497_n 0.0321086f $X=2.18 $Y=2.355 $X2=0
+ $Y2=0
cc_221 N_A_125_367#_M1019_g N_Y_c_576_n 0.0172047f $X=3.28 $Y=2.465 $X2=0 $Y2=0
cc_222 N_A_125_367#_M1004_g Y 0.00352951f $X=2.85 $Y=2.465 $X2=0 $Y2=0
cc_223 N_A_125_367#_M1019_g Y 7.45782e-19 $X=3.28 $Y=2.465 $X2=0 $Y2=0
cc_224 N_A_125_367#_M1004_g Y 0.00635596f $X=2.85 $Y=2.465 $X2=0 $Y2=0
cc_225 N_A_125_367#_M1019_g Y 0.00759475f $X=3.28 $Y=2.465 $X2=0 $Y2=0
cc_226 N_A_125_367#_c_234_n N_Y_c_581_n 0.00989882f $X=2.85 $Y=1.295 $X2=0 $Y2=0
cc_227 N_A_125_367#_M1004_g N_Y_c_581_n 0.0166193f $X=2.85 $Y=2.465 $X2=0 $Y2=0
cc_228 N_A_125_367#_c_236_n N_Y_c_581_n 0.00871516f $X=3.205 $Y=1.37 $X2=0 $Y2=0
cc_229 N_A_125_367#_c_237_n N_Y_c_581_n 0.011207f $X=3.28 $Y=1.295 $X2=0 $Y2=0
cc_230 N_A_125_367#_M1019_g N_Y_c_581_n 0.0177444f $X=3.28 $Y=2.465 $X2=0 $Y2=0
cc_231 N_A_125_367#_c_239_n N_Y_c_581_n 0.0038948f $X=2.85 $Y=1.37 $X2=0 $Y2=0
cc_232 N_A_125_367#_c_240_n N_Y_c_581_n 0.00234261f $X=3.28 $Y=1.37 $X2=0 $Y2=0
cc_233 N_A_125_367#_c_242_n N_Y_c_581_n 0.00495017f $X=2.265 $Y=1.375 $X2=0
+ $Y2=0
cc_234 N_A_125_367#_c_243_n N_Y_c_581_n 0.00588093f $X=2.265 $Y=2.26 $X2=0 $Y2=0
cc_235 N_A_125_367#_c_244_n N_Y_c_581_n 0.0109451f $X=2.4 $Y=1.46 $X2=0 $Y2=0
cc_236 N_A_125_367#_c_241_n N_VGND_M1017_d 0.00975961f $X=2.18 $Y=0.935 $X2=0
+ $Y2=0
cc_237 N_A_125_367#_c_234_n N_VGND_c_637_n 0.00123939f $X=2.85 $Y=1.295 $X2=0
+ $Y2=0
cc_238 N_A_125_367#_c_241_n N_VGND_c_637_n 0.022011f $X=2.18 $Y=0.935 $X2=0
+ $Y2=0
cc_239 N_A_125_367#_c_237_n N_VGND_c_638_n 3.3717e-19 $X=3.28 $Y=1.295 $X2=0
+ $Y2=0
cc_240 N_A_125_367#_c_234_n N_VGND_c_643_n 0.0029147f $X=2.85 $Y=1.295 $X2=0
+ $Y2=0
cc_241 N_A_125_367#_c_237_n N_VGND_c_643_n 0.0029147f $X=3.28 $Y=1.295 $X2=0
+ $Y2=0
cc_242 N_A_125_367#_c_234_n N_VGND_c_645_n 0.00428625f $X=2.85 $Y=1.295 $X2=0
+ $Y2=0
cc_243 N_A_125_367#_c_237_n N_VGND_c_645_n 0.0040339f $X=3.28 $Y=1.295 $X2=0
+ $Y2=0
cc_244 N_A_125_367#_c_241_n N_VGND_c_645_n 0.0126575f $X=2.18 $Y=0.935 $X2=0
+ $Y2=0
cc_245 N_A_125_367#_c_241_n N_A_125_69#_M1018_d 0.00790574f $X=2.18 $Y=0.935
+ $X2=0 $Y2=0
cc_246 N_A_125_367#_M1008_s N_A_125_69#_c_709_n 0.00172464f $X=1.055 $Y=0.345
+ $X2=0 $Y2=0
cc_247 N_A_125_367#_c_241_n N_A_125_69#_c_709_n 0.0376092f $X=2.18 $Y=0.935
+ $X2=0 $Y2=0
cc_248 N_A_125_367#_c_234_n N_A_502_69#_c_725_n 0.00354271f $X=2.85 $Y=1.295
+ $X2=0 $Y2=0
cc_249 N_A_125_367#_c_241_n N_A_502_69#_c_725_n 0.0177033f $X=2.18 $Y=0.935
+ $X2=0 $Y2=0
cc_250 N_A_125_367#_c_242_n N_A_502_69#_c_725_n 0.0123874f $X=2.265 $Y=1.375
+ $X2=0 $Y2=0
cc_251 N_A_125_367#_c_244_n N_A_502_69#_c_725_n 0.00364116f $X=2.4 $Y=1.46 $X2=0
+ $Y2=0
cc_252 N_A_125_367#_c_245_n N_A_502_69#_c_725_n 0.00589524f $X=2.4 $Y=1.37 $X2=0
+ $Y2=0
cc_253 N_A_125_367#_c_234_n N_A_502_69#_c_726_n 0.012797f $X=2.85 $Y=1.295 $X2=0
+ $Y2=0
cc_254 N_A_125_367#_c_237_n N_A_502_69#_c_726_n 0.0121331f $X=3.28 $Y=1.295
+ $X2=0 $Y2=0
cc_255 N_B1_M1011_g N_B2_M1002_g 0.0541449f $X=3.75 $Y=2.465 $X2=0 $Y2=0
cc_256 N_B1_c_346_n N_B2_M1002_g 0.00104941f $X=3.73 $Y=1.51 $X2=0 $Y2=0
cc_257 N_B1_c_354_n N_B2_M1002_g 0.0106797f $X=5.325 $Y=2.005 $X2=0 $Y2=0
cc_258 N_B1_M1012_g N_B2_c_427_n 0.0313168f $X=3.79 $Y=0.765 $X2=0 $Y2=0
cc_259 N_B1_c_343_n N_B2_c_428_n 0.0316897f $X=5.08 $Y=1.295 $X2=0 $Y2=0
cc_260 N_B1_M1013_g N_B2_M1005_g 0.0387451f $X=5.08 $Y=2.465 $X2=0 $Y2=0
cc_261 N_B1_c_354_n N_B2_M1005_g 0.0128139f $X=5.325 $Y=2.005 $X2=0 $Y2=0
cc_262 N_B1_M1011_g B2 4.82035e-19 $X=3.75 $Y=2.465 $X2=0 $Y2=0
cc_263 N_B1_M1012_g B2 0.00384422f $X=3.79 $Y=0.765 $X2=0 $Y2=0
cc_264 N_B1_c_343_n B2 0.00551249f $X=5.08 $Y=1.295 $X2=0 $Y2=0
cc_265 N_B1_M1013_g B2 0.00533139f $X=5.08 $Y=2.465 $X2=0 $Y2=0
cc_266 N_B1_c_345_n B2 0.0127478f $X=5.08 $Y=1.46 $X2=0 $Y2=0
cc_267 N_B1_c_346_n B2 0.0319914f $X=3.73 $Y=1.51 $X2=0 $Y2=0
cc_268 N_B1_c_347_n B2 0.00239443f $X=3.73 $Y=1.51 $X2=0 $Y2=0
cc_269 N_B1_c_354_n B2 0.0807349f $X=5.325 $Y=2.005 $X2=0 $Y2=0
cc_270 N_B1_c_349_n B2 0.0368644f $X=5.49 $Y=1.46 $X2=0 $Y2=0
cc_271 N_B1_M1012_g N_B2_c_431_n 0.00246605f $X=3.79 $Y=0.765 $X2=0 $Y2=0
cc_272 N_B1_c_345_n N_B2_c_431_n 0.0192676f $X=5.08 $Y=1.46 $X2=0 $Y2=0
cc_273 N_B1_c_346_n N_B2_c_431_n 3.70738e-19 $X=3.73 $Y=1.51 $X2=0 $Y2=0
cc_274 N_B1_c_347_n N_B2_c_431_n 0.0204654f $X=3.73 $Y=1.51 $X2=0 $Y2=0
cc_275 N_B1_c_354_n N_B2_c_431_n 7.19152e-19 $X=5.325 $Y=2.005 $X2=0 $Y2=0
cc_276 N_B1_c_346_n N_VPWR_M1019_s 9.55176e-19 $X=3.73 $Y=1.51 $X2=0 $Y2=0
cc_277 N_B1_c_361_n N_VPWR_M1019_s 0.00257041f $X=3.815 $Y=2.005 $X2=0 $Y2=0
cc_278 N_B1_c_354_n N_VPWR_M1013_d 0.0044646f $X=5.325 $Y=2.005 $X2=0 $Y2=0
cc_279 N_B1_c_349_n N_VPWR_M1013_d 0.00145825f $X=5.49 $Y=1.46 $X2=0 $Y2=0
cc_280 N_B1_M1011_g N_VPWR_c_487_n 0.0029183f $X=3.75 $Y=2.465 $X2=0 $Y2=0
cc_281 N_B1_M1013_g N_VPWR_c_488_n 0.0189346f $X=5.08 $Y=2.465 $X2=0 $Y2=0
cc_282 N_B1_c_354_n N_VPWR_c_488_n 0.0231176f $X=5.325 $Y=2.005 $X2=0 $Y2=0
cc_283 N_B1_c_348_n N_VPWR_c_488_n 5.80941e-19 $X=5.49 $Y=1.46 $X2=0 $Y2=0
cc_284 N_B1_M1011_g N_VPWR_c_490_n 0.00426211f $X=3.75 $Y=2.465 $X2=0 $Y2=0
cc_285 N_B1_M1013_g N_VPWR_c_490_n 0.00486043f $X=5.08 $Y=2.465 $X2=0 $Y2=0
cc_286 N_B1_M1011_g N_VPWR_c_482_n 0.00602171f $X=3.75 $Y=2.465 $X2=0 $Y2=0
cc_287 N_B1_M1013_g N_VPWR_c_482_n 0.0082726f $X=5.08 $Y=2.465 $X2=0 $Y2=0
cc_288 N_B1_c_354_n N_Y_M1002_s 0.00412744f $X=5.325 $Y=2.005 $X2=0 $Y2=0
cc_289 N_B1_M1011_g N_Y_c_576_n 0.0183823f $X=3.75 $Y=2.465 $X2=0 $Y2=0
cc_290 N_B1_c_347_n N_Y_c_576_n 2.77545e-19 $X=3.73 $Y=1.51 $X2=0 $Y2=0
cc_291 N_B1_c_354_n N_Y_c_576_n 0.0397835f $X=5.325 $Y=2.005 $X2=0 $Y2=0
cc_292 N_B1_c_361_n N_Y_c_576_n 0.0156021f $X=3.815 $Y=2.005 $X2=0 $Y2=0
cc_293 N_B1_M1011_g Y 8.23998e-19 $X=3.75 $Y=2.465 $X2=0 $Y2=0
cc_294 N_B1_M1011_g N_Y_c_581_n 0.00120174f $X=3.75 $Y=2.465 $X2=0 $Y2=0
cc_295 N_B1_M1012_g N_Y_c_581_n 0.00135911f $X=3.79 $Y=0.765 $X2=0 $Y2=0
cc_296 N_B1_c_346_n N_Y_c_581_n 0.0253457f $X=3.73 $Y=1.51 $X2=0 $Y2=0
cc_297 N_B1_c_347_n N_Y_c_581_n 9.52884e-19 $X=3.73 $Y=1.51 $X2=0 $Y2=0
cc_298 N_B1_c_361_n N_Y_c_581_n 0.00833522f $X=3.815 $Y=2.005 $X2=0 $Y2=0
cc_299 N_B1_c_354_n N_A_765_367#_M1011_s 0.00630874f $X=5.325 $Y=2.005 $X2=-0.19
+ $Y2=-0.245
cc_300 N_B1_c_354_n N_A_765_367#_M1005_d 0.00353353f $X=5.325 $Y=2.005 $X2=0
+ $Y2=0
cc_301 N_B1_M1011_g N_A_765_367#_c_621_n 0.003728f $X=3.75 $Y=2.465 $X2=0 $Y2=0
cc_302 N_B1_c_354_n N_A_765_367#_c_621_n 0.00326627f $X=5.325 $Y=2.005 $X2=0
+ $Y2=0
cc_303 N_B1_c_354_n N_A_765_367#_c_623_n 0.0137681f $X=5.325 $Y=2.005 $X2=0
+ $Y2=0
cc_304 N_B1_M1012_g N_VGND_c_638_n 0.00812868f $X=3.79 $Y=0.765 $X2=0 $Y2=0
cc_305 N_B1_c_343_n N_VGND_c_639_n 0.0108625f $X=5.08 $Y=1.295 $X2=0 $Y2=0
cc_306 N_B1_M1012_g N_VGND_c_643_n 0.00400407f $X=3.79 $Y=0.765 $X2=0 $Y2=0
cc_307 N_B1_c_343_n N_VGND_c_644_n 0.00400407f $X=5.08 $Y=1.295 $X2=0 $Y2=0
cc_308 N_B1_M1012_g N_VGND_c_645_n 0.00779262f $X=3.79 $Y=0.765 $X2=0 $Y2=0
cc_309 N_B1_c_343_n N_VGND_c_645_n 0.00799365f $X=5.08 $Y=1.295 $X2=0 $Y2=0
cc_310 N_B1_M1012_g N_A_502_69#_c_726_n 8.32438e-19 $X=3.79 $Y=0.765 $X2=0 $Y2=0
cc_311 N_B1_M1012_g N_A_502_69#_c_741_n 0.0140269f $X=3.79 $Y=0.765 $X2=0 $Y2=0
cc_312 N_B1_c_346_n N_A_502_69#_c_741_n 0.00587907f $X=3.73 $Y=1.51 $X2=0 $Y2=0
cc_313 N_B1_c_346_n N_A_502_69#_c_743_n 0.005434f $X=3.73 $Y=1.51 $X2=0 $Y2=0
cc_314 N_B1_c_347_n N_A_502_69#_c_743_n 7.17863e-19 $X=3.73 $Y=1.51 $X2=0 $Y2=0
cc_315 N_B1_c_343_n N_A_502_69#_c_729_n 0.0120345f $X=5.08 $Y=1.295 $X2=0 $Y2=0
cc_316 N_B1_c_348_n N_A_502_69#_c_729_n 0.00585131f $X=5.49 $Y=1.46 $X2=0 $Y2=0
cc_317 N_B1_c_349_n N_A_502_69#_c_729_n 0.00866423f $X=5.49 $Y=1.46 $X2=0 $Y2=0
cc_318 N_B1_c_343_n N_A_502_69#_c_730_n 4.46816e-19 $X=5.08 $Y=1.295 $X2=0 $Y2=0
cc_319 N_B2_M1005_g N_VPWR_c_488_n 0.0013781f $X=4.65 $Y=2.465 $X2=0 $Y2=0
cc_320 N_B2_M1002_g N_VPWR_c_490_n 0.00357877f $X=4.18 $Y=2.465 $X2=0 $Y2=0
cc_321 N_B2_M1005_g N_VPWR_c_490_n 0.0035787f $X=4.65 $Y=2.465 $X2=0 $Y2=0
cc_322 N_B2_M1002_g N_VPWR_c_482_n 0.00551666f $X=4.18 $Y=2.465 $X2=0 $Y2=0
cc_323 N_B2_M1005_g N_VPWR_c_482_n 0.00544851f $X=4.65 $Y=2.465 $X2=0 $Y2=0
cc_324 N_B2_M1002_g N_Y_c_576_n 0.0126151f $X=4.18 $Y=2.465 $X2=0 $Y2=0
cc_325 N_B2_M1002_g N_A_765_367#_c_621_n 0.0118408f $X=4.18 $Y=2.465 $X2=0 $Y2=0
cc_326 N_B2_M1005_g N_A_765_367#_c_621_n 0.0140573f $X=4.65 $Y=2.465 $X2=0 $Y2=0
cc_327 N_B2_M1002_g N_A_765_367#_c_623_n 7.2395e-19 $X=4.18 $Y=2.465 $X2=0 $Y2=0
cc_328 N_B2_M1005_g N_A_765_367#_c_623_n 0.00657933f $X=4.65 $Y=2.465 $X2=0
+ $Y2=0
cc_329 N_B2_c_427_n N_VGND_c_638_n 0.00833189f $X=4.22 $Y=1.295 $X2=0 $Y2=0
cc_330 N_B2_c_428_n N_VGND_c_638_n 4.39455e-19 $X=4.65 $Y=1.295 $X2=0 $Y2=0
cc_331 N_B2_c_427_n N_VGND_c_639_n 4.39455e-19 $X=4.22 $Y=1.295 $X2=0 $Y2=0
cc_332 N_B2_c_428_n N_VGND_c_639_n 0.00833189f $X=4.65 $Y=1.295 $X2=0 $Y2=0
cc_333 N_B2_c_427_n N_VGND_c_640_n 0.00400407f $X=4.22 $Y=1.295 $X2=0 $Y2=0
cc_334 N_B2_c_428_n N_VGND_c_640_n 0.00400407f $X=4.65 $Y=1.295 $X2=0 $Y2=0
cc_335 N_B2_c_427_n N_VGND_c_645_n 0.00774504f $X=4.22 $Y=1.295 $X2=0 $Y2=0
cc_336 N_B2_c_428_n N_VGND_c_645_n 0.00774504f $X=4.65 $Y=1.295 $X2=0 $Y2=0
cc_337 N_B2_c_427_n N_A_502_69#_c_741_n 0.0120345f $X=4.22 $Y=1.295 $X2=0 $Y2=0
cc_338 B2 N_A_502_69#_c_741_n 0.0232416f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_339 N_B2_c_427_n N_A_502_69#_c_728_n 4.63537e-19 $X=4.22 $Y=1.295 $X2=0 $Y2=0
cc_340 N_B2_c_428_n N_A_502_69#_c_728_n 4.63537e-19 $X=4.65 $Y=1.295 $X2=0 $Y2=0
cc_341 N_B2_c_428_n N_A_502_69#_c_729_n 0.0120345f $X=4.65 $Y=1.295 $X2=0 $Y2=0
cc_342 B2 N_A_502_69#_c_729_n 0.0428415f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_343 B2 N_A_502_69#_c_755_n 0.0160632f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_344 N_B2_c_431_n N_A_502_69#_c_755_n 6.37488e-19 $X=4.65 $Y=1.46 $X2=0 $Y2=0
cc_345 N_VPWR_c_482_n N_Y_M1004_d 0.00223559f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_346 N_VPWR_c_482_n N_Y_M1002_s 0.00257355f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_347 N_VPWR_M1019_s N_Y_c_576_n 0.00902219f $X=3.355 $Y=1.835 $X2=0 $Y2=0
cc_348 N_VPWR_c_487_n N_Y_c_576_n 0.0169036f $X=3.515 $Y=2.925 $X2=0 $Y2=0
cc_349 N_VPWR_c_490_n N_Y_c_576_n 0.00201952f $X=5.13 $Y=3.33 $X2=0 $Y2=0
cc_350 N_VPWR_c_493_n N_Y_c_576_n 0.00201346f $X=3.4 $Y=3.33 $X2=0 $Y2=0
cc_351 N_VPWR_c_482_n N_Y_c_576_n 0.0101116f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_352 N_VPWR_c_493_n Y 0.0189236f $X=3.4 $Y=3.33 $X2=0 $Y2=0
cc_353 N_VPWR_c_482_n Y 0.0123859f $X=5.52 $Y=3.33 $X2=0 $Y2=0
cc_354 N_VPWR_c_486_n N_Y_c_581_n 0.0173981f $X=2.635 $Y=1.98 $X2=0 $Y2=0
cc_355 N_VPWR_c_482_n N_A_765_367#_M1011_s 0.00223577f $X=5.52 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_356 N_VPWR_c_482_n N_A_765_367#_M1005_d 0.00411411f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_357 N_VPWR_c_490_n N_A_765_367#_c_621_n 0.0671356f $X=5.13 $Y=3.33 $X2=0
+ $Y2=0
cc_358 N_VPWR_c_482_n N_A_765_367#_c_621_n 0.0422944f $X=5.52 $Y=3.33 $X2=0
+ $Y2=0
cc_359 N_VPWR_c_486_n N_A_502_69#_c_725_n 0.00621462f $X=2.635 $Y=1.98 $X2=0
+ $Y2=0
cc_360 N_Y_c_576_n N_A_765_367#_M1011_s 0.00355644f $X=4.415 $Y=2.425 $X2=1.055
+ $Y2=0.345
cc_361 N_Y_M1002_s N_A_765_367#_c_621_n 0.00420878f $X=4.255 $Y=1.835 $X2=0
+ $Y2=0
cc_362 N_Y_c_576_n N_A_765_367#_c_621_n 0.0411635f $X=4.415 $Y=2.425 $X2=0 $Y2=0
cc_363 N_Y_c_581_n N_A_502_69#_c_725_n 0.0236268f $X=3.065 $Y=0.68 $X2=2.85
+ $Y2=1.445
cc_364 N_Y_M1000_d N_A_502_69#_c_726_n 0.00176461f $X=2.925 $Y=0.345 $X2=2.85
+ $Y2=2.465
cc_365 N_Y_c_581_n N_A_502_69#_c_726_n 0.0159805f $X=3.065 $Y=0.68 $X2=2.85
+ $Y2=2.465
cc_366 N_VGND_c_636_n N_A_125_69#_c_708_n 0.0164324f $X=0.335 $Y=0.49 $X2=0
+ $Y2=0
cc_367 N_VGND_c_642_n N_A_125_69#_c_708_n 0.0116964f $X=1.89 $Y=0 $X2=0 $Y2=0
cc_368 N_VGND_c_645_n N_A_125_69#_c_708_n 0.00814876f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_369 N_VGND_c_637_n N_A_125_69#_c_709_n 0.0144096f $X=2.055 $Y=0.535 $X2=0
+ $Y2=0
cc_370 N_VGND_c_642_n N_A_125_69#_c_709_n 0.0429744f $X=1.89 $Y=0 $X2=0 $Y2=0
cc_371 N_VGND_c_645_n N_A_125_69#_c_709_n 0.0301682f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_372 N_VGND_c_637_n N_A_502_69#_c_725_n 0.0123762f $X=2.055 $Y=0.535 $X2=0
+ $Y2=0
cc_373 N_VGND_c_638_n N_A_502_69#_c_726_n 0.0105582f $X=4.005 $Y=0.575 $X2=0
+ $Y2=0
cc_374 N_VGND_c_643_n N_A_502_69#_c_726_n 0.0615114f $X=3.84 $Y=0 $X2=0 $Y2=0
cc_375 N_VGND_c_645_n N_A_502_69#_c_726_n 0.0343015f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_376 N_VGND_c_637_n N_A_502_69#_c_727_n 0.00997144f $X=2.055 $Y=0.535 $X2=0
+ $Y2=0
cc_377 N_VGND_c_643_n N_A_502_69#_c_727_n 0.0150542f $X=3.84 $Y=0 $X2=0 $Y2=0
cc_378 N_VGND_c_645_n N_A_502_69#_c_727_n 0.00816431f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_379 N_VGND_M1012_d N_A_502_69#_c_741_n 0.00554099f $X=3.865 $Y=0.345 $X2=0
+ $Y2=0
cc_380 N_VGND_c_638_n N_A_502_69#_c_741_n 0.0170777f $X=4.005 $Y=0.575 $X2=0
+ $Y2=0
cc_381 N_VGND_c_638_n N_A_502_69#_c_728_n 0.0147979f $X=4.005 $Y=0.575 $X2=0
+ $Y2=0
cc_382 N_VGND_c_639_n N_A_502_69#_c_728_n 0.0147979f $X=4.865 $Y=0.575 $X2=0
+ $Y2=0
cc_383 N_VGND_c_640_n N_A_502_69#_c_728_n 0.00935612f $X=4.7 $Y=0 $X2=0 $Y2=0
cc_384 N_VGND_c_645_n N_A_502_69#_c_728_n 0.00705762f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_385 N_VGND_M1010_s N_A_502_69#_c_729_n 0.00353353f $X=4.725 $Y=0.345 $X2=0
+ $Y2=0
cc_386 N_VGND_c_639_n N_A_502_69#_c_729_n 0.0170777f $X=4.865 $Y=0.575 $X2=0
+ $Y2=0
cc_387 N_VGND_c_639_n N_A_502_69#_c_730_n 0.0148334f $X=4.865 $Y=0.575 $X2=0
+ $Y2=0
cc_388 N_VGND_c_644_n N_A_502_69#_c_730_n 0.0128398f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_389 N_VGND_c_645_n N_A_502_69#_c_730_n 0.00968545f $X=5.52 $Y=0 $X2=0 $Y2=0
