* File: sky130_fd_sc_lp__ha_1.pxi.spice
* Created: Wed Sep  2 09:54:23 2020
* 
x_PM_SKY130_FD_SC_LP__HA_1%A_80_30# N_A_80_30#_M1007_s N_A_80_30#_M1008_d
+ N_A_80_30#_M1009_g N_A_80_30#_M1003_g N_A_80_30#_c_101_n N_A_80_30#_c_102_n
+ N_A_80_30#_c_103_n N_A_80_30#_c_104_n N_A_80_30#_c_105_n N_A_80_30#_c_106_n
+ N_A_80_30#_c_107_n N_A_80_30#_c_118_p N_A_80_30#_c_108_n
+ PM_SKY130_FD_SC_LP__HA_1%A_80_30#
x_PM_SKY130_FD_SC_LP__HA_1%A_223_320# N_A_223_320#_M1010_s N_A_223_320#_M1006_d
+ N_A_223_320#_M1007_g N_A_223_320#_M1008_g N_A_223_320#_M1013_g
+ N_A_223_320#_M1001_g N_A_223_320#_c_164_n N_A_223_320#_c_176_n
+ N_A_223_320#_c_177_n N_A_223_320#_c_178_n N_A_223_320#_c_179_n
+ N_A_223_320#_c_180_n N_A_223_320#_c_165_n N_A_223_320#_c_181_n
+ N_A_223_320#_c_166_n N_A_223_320#_c_167_n N_A_223_320#_c_168_n
+ N_A_223_320#_c_169_n N_A_223_320#_c_183_n N_A_223_320#_c_170_n
+ N_A_223_320#_c_171_n N_A_223_320#_c_172_n PM_SKY130_FD_SC_LP__HA_1%A_223_320#
x_PM_SKY130_FD_SC_LP__HA_1%B N_B_M1012_g N_B_M1002_g N_B_c_299_n N_B_M1010_g
+ N_B_M1006_g N_B_c_301_n N_B_c_310_n N_B_c_302_n N_B_c_303_n N_B_c_304_n B
+ N_B_c_305_n N_B_c_306_n PM_SKY130_FD_SC_LP__HA_1%B
x_PM_SKY130_FD_SC_LP__HA_1%A N_A_c_386_n N_A_M1004_g N_A_M1011_g N_A_c_387_n
+ N_A_c_388_n N_A_c_389_n N_A_c_390_n N_A_c_391_n N_A_M1005_g N_A_M1000_g
+ N_A_c_399_n A N_A_c_394_n N_A_c_395_n PM_SKY130_FD_SC_LP__HA_1%A
x_PM_SKY130_FD_SC_LP__HA_1%SUM N_SUM_M1009_s N_SUM_M1003_s SUM SUM SUM SUM SUM
+ SUM SUM N_SUM_c_477_n SUM N_SUM_c_480_n PM_SKY130_FD_SC_LP__HA_1%SUM
x_PM_SKY130_FD_SC_LP__HA_1%VPWR N_VPWR_M1003_d N_VPWR_M1011_d N_VPWR_M1000_d
+ N_VPWR_c_494_n N_VPWR_c_495_n N_VPWR_c_496_n N_VPWR_c_497_n N_VPWR_c_498_n
+ VPWR N_VPWR_c_499_n N_VPWR_c_500_n N_VPWR_c_501_n N_VPWR_c_493_n
+ N_VPWR_c_503_n N_VPWR_c_504_n PM_SKY130_FD_SC_LP__HA_1%VPWR
x_PM_SKY130_FD_SC_LP__HA_1%COUT N_COUT_M1013_d N_COUT_M1001_d COUT COUT COUT
+ COUT COUT COUT COUT N_COUT_c_554_n COUT PM_SKY130_FD_SC_LP__HA_1%COUT
x_PM_SKY130_FD_SC_LP__HA_1%VGND N_VGND_M1009_d N_VGND_M1012_d N_VGND_M1005_d
+ N_VGND_c_569_n N_VGND_c_570_n N_VGND_c_571_n N_VGND_c_572_n N_VGND_c_573_n
+ VGND N_VGND_c_574_n N_VGND_c_575_n N_VGND_c_576_n N_VGND_c_577_n
+ N_VGND_c_578_n N_VGND_c_579_n PM_SKY130_FD_SC_LP__HA_1%VGND
x_PM_SKY130_FD_SC_LP__HA_1%A_307_62# N_A_307_62#_M1007_d N_A_307_62#_M1004_d
+ N_A_307_62#_c_624_n N_A_307_62#_c_625_n N_A_307_62#_c_626_n
+ N_A_307_62#_c_627_n PM_SKY130_FD_SC_LP__HA_1%A_307_62#
cc_1 VNB N_A_80_30#_M1003_g 0.00614907f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=2.465
cc_2 VNB N_A_80_30#_c_101_n 0.0138405f $X=-0.19 $Y=-0.245 $X2=1.08 $Y2=1.315
cc_3 VNB N_A_80_30#_c_102_n 0.0168321f $X=-0.19 $Y=-0.245 $X2=1.245 $Y2=0.52
cc_4 VNB N_A_80_30#_c_103_n 0.00364487f $X=-0.19 $Y=-0.245 $X2=1.545 $Y2=1.315
cc_5 VNB N_A_80_30#_c_104_n 0.0037274f $X=-0.19 $Y=-0.245 $X2=1.63 $Y2=2.175
cc_6 VNB N_A_80_30#_c_105_n 0.00433346f $X=-0.19 $Y=-0.245 $X2=0.665 $Y2=1.315
cc_7 VNB N_A_80_30#_c_106_n 0.0445031f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.395
cc_8 VNB N_A_80_30#_c_107_n 0.00432084f $X=-0.19 $Y=-0.245 $X2=1.225 $Y2=1.315
cc_9 VNB N_A_80_30#_c_108_n 0.0222826f $X=-0.19 $Y=-0.245 $X2=0.597 $Y2=1.23
cc_10 VNB N_A_223_320#_M1007_g 0.0628344f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.7
cc_11 VNB N_A_223_320#_M1001_g 0.00397561f $X=-0.19 $Y=-0.245 $X2=1.545
+ $Y2=1.315
cc_12 VNB N_A_223_320#_c_164_n 0.00166723f $X=-0.19 $Y=-0.245 $X2=0.665
+ $Y2=1.315
cc_13 VNB N_A_223_320#_c_165_n 0.00372035f $X=-0.19 $Y=-0.245 $X2=1.715 $Y2=2.34
cc_14 VNB N_A_223_320#_c_166_n 9.0175e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_223_320#_c_167_n 3.73364e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_223_320#_c_168_n 0.0061012f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_223_320#_c_169_n 0.0382984f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_223_320#_c_170_n 0.00195478f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_223_320#_c_171_n 0.0122026f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_223_320#_c_172_n 0.0208659f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_B_M1012_g 0.0341127f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_B_c_299_n 0.0166942f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.7
cc_23 VNB N_B_M1006_g 0.00343759f $X=-0.19 $Y=-0.245 $X2=1.08 $Y2=1.315
cc_24 VNB N_B_c_301_n 0.0219776f $X=-0.19 $Y=-0.245 $X2=1.245 $Y2=0.52
cc_25 VNB N_B_c_302_n 0.0196709f $X=-0.19 $Y=-0.245 $X2=1.63 $Y2=1.4
cc_26 VNB N_B_c_303_n 0.00221373f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_B_c_304_n 0.0160237f $X=-0.19 $Y=-0.245 $X2=0.665 $Y2=1.395
cc_28 VNB N_B_c_305_n 4.08926e-19 $X=-0.19 $Y=-0.245 $X2=1.715 $Y2=2.34
cc_29 VNB N_B_c_306_n 0.0425417f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_c_386_n 0.0175152f $X=-0.19 $Y=-0.245 $X2=1.12 $Y2=0.31
cc_31 VNB N_A_c_387_n 0.02028f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=1.56
cc_32 VNB N_A_c_388_n 0.0120216f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=2.465
cc_33 VNB N_A_c_389_n 0.0331906f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_c_390_n 0.0600564f $X=-0.19 $Y=-0.245 $X2=1.08 $Y2=1.315
cc_35 VNB N_A_c_391_n 0.0103145f $X=-0.19 $Y=-0.245 $X2=0.795 $Y2=1.315
cc_36 VNB N_A_M1005_g 0.0488476f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB A 0.00216615f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_c_394_n 0.0149168f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_c_395_n 0.0299847f $X=-0.19 $Y=-0.245 $X2=1.715 $Y2=2.34
cc_40 VNB N_SUM_c_477_n 0.0632793f $X=-0.19 $Y=-0.245 $X2=0.665 $Y2=1.315
cc_41 VNB N_VPWR_c_493_n 0.203486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB COUT 0.0307111f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.7
cc_43 VNB N_COUT_c_554_n 0.0298043f $X=-0.19 $Y=-0.245 $X2=0.665 $Y2=1.315
cc_44 VNB COUT 0.00856429f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_569_n 0.012484f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=2.465
cc_46 VNB N_VGND_c_570_n 0.00242f $X=-0.19 $Y=-0.245 $X2=1.225 $Y2=1.23
cc_47 VNB N_VGND_c_571_n 0.0107126f $X=-0.19 $Y=-0.245 $X2=1.545 $Y2=1.315
cc_48 VNB N_VGND_c_572_n 0.0433081f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_573_n 0.00640763f $X=-0.19 $Y=-0.245 $X2=0.665 $Y2=1.395
cc_50 VNB N_VGND_c_574_n 0.0159208f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_575_n 0.0299186f $X=-0.19 $Y=-0.245 $X2=1.715 $Y2=2.34
cc_52 VNB N_VGND_c_576_n 0.0187066f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_577_n 0.274799f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_578_n 0.0053257f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_579_n 0.00531f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_307_62#_c_624_n 0.00192983f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.7
cc_57 VNB N_A_307_62#_c_625_n 0.00966742f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=2.465
cc_58 VNB N_A_307_62#_c_626_n 0.00553528f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=2.465
cc_59 VNB N_A_307_62#_c_627_n 0.00604786f $X=-0.19 $Y=-0.245 $X2=0.795 $Y2=1.315
cc_60 VPB N_A_80_30#_M1003_g 0.0270606f $X=-0.19 $Y=1.655 $X2=0.615 $Y2=2.465
cc_61 VPB N_A_80_30#_c_104_n 0.00456337f $X=-0.19 $Y=1.655 $X2=1.63 $Y2=2.175
cc_62 VPB N_A_223_320#_M1008_g 0.0221654f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_63 VPB N_A_223_320#_M1001_g 0.0260557f $X=-0.19 $Y=1.655 $X2=1.545 $Y2=1.315
cc_64 VPB N_A_223_320#_c_164_n 0.00499468f $X=-0.19 $Y=1.655 $X2=0.665 $Y2=1.315
cc_65 VPB N_A_223_320#_c_176_n 0.0284617f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=1.395
cc_66 VPB N_A_223_320#_c_177_n 0.0037045f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=1.395
cc_67 VPB N_A_223_320#_c_178_n 0.00160392f $X=-0.19 $Y=1.655 $X2=1.225 $Y2=1.315
cc_68 VPB N_A_223_320#_c_179_n 0.0200034f $X=-0.19 $Y=1.655 $X2=1.63 $Y2=2.34
cc_69 VPB N_A_223_320#_c_180_n 0.00265684f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_70 VPB N_A_223_320#_c_181_n 3.62765e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_71 VPB N_A_223_320#_c_167_n 0.00221245f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_72 VPB N_A_223_320#_c_183_n 7.58183e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_73 VPB N_A_223_320#_c_171_n 0.0372415f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_74 VPB N_B_M1002_g 0.0252468f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=1.23
cc_75 VPB N_B_M1006_g 0.0404155f $X=-0.19 $Y=1.655 $X2=1.08 $Y2=1.315
cc_76 VPB N_B_c_301_n 0.00569565f $X=-0.19 $Y=1.655 $X2=1.245 $Y2=0.52
cc_77 VPB N_B_c_310_n 0.0206012f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_78 VPB N_B_c_305_n 0.00312283f $X=-0.19 $Y=1.655 $X2=1.715 $Y2=2.34
cc_79 VPB N_A_M1011_g 0.031429f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.7
cc_80 VPB N_A_M1005_g 0.00914566f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_81 VPB N_A_M1000_g 0.0210266f $X=-0.19 $Y=1.655 $X2=1.63 $Y2=1.4
cc_82 VPB N_A_c_399_n 0.0104874f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=1.395
cc_83 VPB A 0.00270009f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_84 VPB N_A_c_394_n 0.0168794f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_85 VPB SUM 0.0134994f $X=-0.19 $Y=1.655 $X2=0.615 $Y2=1.56
cc_86 VPB N_SUM_c_477_n 0.00471859f $X=-0.19 $Y=1.655 $X2=0.665 $Y2=1.315
cc_87 VPB N_SUM_c_480_n 0.0519868f $X=-0.19 $Y=1.655 $X2=0.597 $Y2=1.23
cc_88 VPB N_VPWR_c_494_n 0.0237779f $X=-0.19 $Y=1.655 $X2=0.615 $Y2=2.465
cc_89 VPB N_VPWR_c_495_n 0.0326204f $X=-0.19 $Y=1.655 $X2=1.545 $Y2=1.315
cc_90 VPB N_VPWR_c_496_n 0.0174131f $X=-0.19 $Y=1.655 $X2=0.665 $Y2=1.315
cc_91 VPB N_VPWR_c_497_n 0.0213759f $X=-0.19 $Y=1.655 $X2=1.63 $Y2=2.34
cc_92 VPB N_VPWR_c_498_n 0.00574453f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_93 VPB N_VPWR_c_499_n 0.0430759f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_94 VPB N_VPWR_c_500_n 0.0190296f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_95 VPB N_VPWR_c_501_n 0.0164025f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_96 VPB N_VPWR_c_493_n 0.0823937f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_97 VPB N_VPWR_c_503_n 0.0117073f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_98 VPB N_VPWR_c_504_n 0.00609234f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_99 VPB COUT 0.0606284f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.7
cc_100 N_A_80_30#_M1003_g N_A_223_320#_M1007_g 8.52072e-19 $X=0.615 $Y=2.465
+ $X2=0 $Y2=0
cc_101 N_A_80_30#_c_102_n N_A_223_320#_M1007_g 0.0156444f $X=1.245 $Y=0.52 $X2=0
+ $Y2=0
cc_102 N_A_80_30#_c_103_n N_A_223_320#_M1007_g 0.0201365f $X=1.545 $Y=1.315
+ $X2=0 $Y2=0
cc_103 N_A_80_30#_c_104_n N_A_223_320#_M1007_g 0.00666449f $X=1.63 $Y=2.175
+ $X2=0 $Y2=0
cc_104 N_A_80_30#_c_105_n N_A_223_320#_M1007_g 9.04632e-19 $X=0.665 $Y=1.315
+ $X2=0 $Y2=0
cc_105 N_A_80_30#_c_106_n N_A_223_320#_M1007_g 0.00603418f $X=0.63 $Y=1.395
+ $X2=0 $Y2=0
cc_106 N_A_80_30#_c_104_n N_A_223_320#_M1008_g 0.00438381f $X=1.63 $Y=2.175
+ $X2=0 $Y2=0
cc_107 N_A_80_30#_c_118_p N_A_223_320#_M1008_g 0.00418655f $X=1.715 $Y=2.34
+ $X2=0 $Y2=0
cc_108 N_A_80_30#_M1003_g N_A_223_320#_c_164_n 0.00108886f $X=0.615 $Y=2.465
+ $X2=0 $Y2=0
cc_109 N_A_80_30#_c_104_n N_A_223_320#_c_164_n 0.0387478f $X=1.63 $Y=2.175 $X2=0
+ $Y2=0
cc_110 N_A_80_30#_c_107_n N_A_223_320#_c_164_n 0.013243f $X=1.225 $Y=1.315 $X2=0
+ $Y2=0
cc_111 N_A_80_30#_c_118_p N_A_223_320#_c_164_n 0.023309f $X=1.715 $Y=2.34 $X2=0
+ $Y2=0
cc_112 N_A_80_30#_c_118_p N_A_223_320#_c_176_n 0.0209672f $X=1.715 $Y=2.34 $X2=0
+ $Y2=0
cc_113 N_A_80_30#_c_104_n N_A_223_320#_c_178_n 0.00225421f $X=1.63 $Y=2.175
+ $X2=0 $Y2=0
cc_114 N_A_80_30#_c_118_p N_A_223_320#_c_178_n 0.0120846f $X=1.715 $Y=2.34 $X2=0
+ $Y2=0
cc_115 N_A_80_30#_c_104_n N_A_223_320#_c_180_n 0.00601104f $X=1.63 $Y=2.175
+ $X2=0 $Y2=0
cc_116 N_A_80_30#_M1003_g N_A_223_320#_c_171_n 0.00802512f $X=0.615 $Y=2.465
+ $X2=0 $Y2=0
cc_117 N_A_80_30#_c_103_n N_A_223_320#_c_171_n 8.47085e-19 $X=1.545 $Y=1.315
+ $X2=0 $Y2=0
cc_118 N_A_80_30#_c_104_n N_A_223_320#_c_171_n 0.00414416f $X=1.63 $Y=2.175
+ $X2=0 $Y2=0
cc_119 N_A_80_30#_c_107_n N_A_223_320#_c_171_n 0.005046f $X=1.225 $Y=1.315 $X2=0
+ $Y2=0
cc_120 N_A_80_30#_c_104_n N_B_M1002_g 0.00306132f $X=1.63 $Y=2.175 $X2=0 $Y2=0
cc_121 N_A_80_30#_c_118_p N_B_M1002_g 0.00670105f $X=1.715 $Y=2.34 $X2=0 $Y2=0
cc_122 N_A_80_30#_c_104_n N_B_c_301_n 0.0042927f $X=1.63 $Y=2.175 $X2=0 $Y2=0
cc_123 N_A_80_30#_c_102_n N_B_c_303_n 0.0016525f $X=1.245 $Y=0.52 $X2=0 $Y2=0
cc_124 N_A_80_30#_c_103_n N_B_c_303_n 0.0151125f $X=1.545 $Y=1.315 $X2=0 $Y2=0
cc_125 N_A_80_30#_c_104_n N_B_c_303_n 0.0331017f $X=1.63 $Y=2.175 $X2=0 $Y2=0
cc_126 N_A_80_30#_c_103_n N_B_c_304_n 0.00137199f $X=1.545 $Y=1.315 $X2=0 $Y2=0
cc_127 N_A_80_30#_c_118_p N_A_M1011_g 3.16646e-19 $X=1.715 $Y=2.34 $X2=0 $Y2=0
cc_128 N_A_80_30#_M1003_g SUM 0.00672799f $X=0.615 $Y=2.465 $X2=0 $Y2=0
cc_129 N_A_80_30#_c_106_n SUM 0.00497804f $X=0.63 $Y=1.395 $X2=0 $Y2=0
cc_130 N_A_80_30#_M1003_g N_SUM_c_477_n 0.0064424f $X=0.615 $Y=2.465 $X2=0 $Y2=0
cc_131 N_A_80_30#_c_105_n N_SUM_c_477_n 0.025257f $X=0.665 $Y=1.315 $X2=0 $Y2=0
cc_132 N_A_80_30#_c_108_n N_SUM_c_477_n 0.0172808f $X=0.597 $Y=1.23 $X2=0 $Y2=0
cc_133 N_A_80_30#_M1003_g N_VPWR_c_494_n 0.00864197f $X=0.615 $Y=2.465 $X2=0
+ $Y2=0
cc_134 N_A_80_30#_c_101_n N_VPWR_c_494_n 0.0104152f $X=1.08 $Y=1.315 $X2=0 $Y2=0
cc_135 N_A_80_30#_c_105_n N_VPWR_c_494_n 0.00425239f $X=0.665 $Y=1.315 $X2=0
+ $Y2=0
cc_136 N_A_80_30#_c_106_n N_VPWR_c_494_n 5.12317e-19 $X=0.63 $Y=1.395 $X2=0
+ $Y2=0
cc_137 N_A_80_30#_M1003_g N_VPWR_c_497_n 0.00585385f $X=0.615 $Y=2.465 $X2=0
+ $Y2=0
cc_138 N_A_80_30#_M1003_g N_VPWR_c_493_n 0.0129312f $X=0.615 $Y=2.465 $X2=0
+ $Y2=0
cc_139 N_A_80_30#_c_101_n N_VGND_c_569_n 0.00494775f $X=1.08 $Y=1.315 $X2=0
+ $Y2=0
cc_140 N_A_80_30#_c_102_n N_VGND_c_569_n 0.0476791f $X=1.245 $Y=0.52 $X2=0 $Y2=0
cc_141 N_A_80_30#_c_105_n N_VGND_c_569_n 0.0187623f $X=0.665 $Y=1.315 $X2=0
+ $Y2=0
cc_142 N_A_80_30#_c_106_n N_VGND_c_569_n 0.00174523f $X=0.63 $Y=1.395 $X2=0
+ $Y2=0
cc_143 N_A_80_30#_c_108_n N_VGND_c_569_n 0.0152646f $X=0.597 $Y=1.23 $X2=0 $Y2=0
cc_144 N_A_80_30#_c_108_n N_VGND_c_574_n 0.00485045f $X=0.597 $Y=1.23 $X2=0
+ $Y2=0
cc_145 N_A_80_30#_c_102_n N_VGND_c_575_n 0.0114791f $X=1.245 $Y=0.52 $X2=0 $Y2=0
cc_146 N_A_80_30#_c_102_n N_VGND_c_577_n 0.0106048f $X=1.245 $Y=0.52 $X2=0 $Y2=0
cc_147 N_A_80_30#_c_108_n N_VGND_c_577_n 0.00942718f $X=0.597 $Y=1.23 $X2=0
+ $Y2=0
cc_148 N_A_80_30#_c_102_n N_A_307_62#_c_624_n 0.00870118f $X=1.245 $Y=0.52 $X2=0
+ $Y2=0
cc_149 N_A_80_30#_c_102_n N_A_307_62#_c_626_n 0.0148899f $X=1.245 $Y=0.52 $X2=0
+ $Y2=0
cc_150 N_A_80_30#_c_103_n N_A_307_62#_c_626_n 0.0135554f $X=1.545 $Y=1.315 $X2=0
+ $Y2=0
cc_151 N_A_223_320#_M1007_g N_B_M1012_g 0.024921f $X=1.46 $Y=0.52 $X2=0 $Y2=0
cc_152 N_A_223_320#_c_176_n N_B_M1002_g 0.00931885f $X=2.3 $Y=2.78 $X2=0 $Y2=0
cc_153 N_A_223_320#_c_178_n N_B_M1002_g 0.0062319f $X=2.385 $Y=2.675 $X2=0 $Y2=0
cc_154 N_A_223_320#_c_180_n N_B_M1002_g 0.00180152f $X=2.47 $Y=2.015 $X2=0 $Y2=0
cc_155 N_A_223_320#_c_171_n N_B_M1002_g 0.0170374f $X=1.46 $Y=1.765 $X2=0 $Y2=0
cc_156 N_A_223_320#_c_165_n N_B_c_299_n 0.0154956f $X=3.44 $Y=0.907 $X2=0 $Y2=0
cc_157 N_A_223_320#_c_166_n N_B_c_299_n 0.00412394f $X=3.53 $Y=1.26 $X2=0 $Y2=0
cc_158 N_A_223_320#_c_179_n N_B_M1006_g 0.0186695f $X=3.42 $Y=2.015 $X2=0 $Y2=0
cc_159 N_A_223_320#_c_181_n N_B_M1006_g 0.00102623f $X=3.515 $Y=2.34 $X2=0 $Y2=0
cc_160 N_A_223_320#_c_167_n N_B_M1006_g 0.00527343f $X=3.56 $Y=1.93 $X2=0 $Y2=0
cc_161 N_A_223_320#_c_171_n N_B_c_301_n 0.024921f $X=1.46 $Y=1.765 $X2=0 $Y2=0
cc_162 N_A_223_320#_c_171_n N_B_c_310_n 0.00627075f $X=1.46 $Y=1.765 $X2=0 $Y2=0
cc_163 N_A_223_320#_c_179_n N_B_c_302_n 0.00579113f $X=3.42 $Y=2.015 $X2=0 $Y2=0
cc_164 N_A_223_320#_c_180_n N_B_c_302_n 5.74729e-19 $X=2.47 $Y=2.015 $X2=0 $Y2=0
cc_165 N_A_223_320#_c_165_n N_B_c_302_n 0.0267699f $X=3.44 $Y=0.907 $X2=0 $Y2=0
cc_166 N_A_223_320#_c_166_n N_B_c_302_n 0.00232685f $X=3.53 $Y=1.26 $X2=0 $Y2=0
cc_167 N_A_223_320#_c_170_n N_B_c_302_n 0.01248f $X=3.56 $Y=1.425 $X2=0 $Y2=0
cc_168 N_A_223_320#_M1007_g N_B_c_303_n 3.09492e-19 $X=1.46 $Y=0.52 $X2=0 $Y2=0
cc_169 N_A_223_320#_c_179_n N_B_c_305_n 0.0251263f $X=3.42 $Y=2.015 $X2=0 $Y2=0
cc_170 N_A_223_320#_c_167_n N_B_c_305_n 0.0129813f $X=3.56 $Y=1.93 $X2=0 $Y2=0
cc_171 N_A_223_320#_c_170_n N_B_c_305_n 0.0159155f $X=3.56 $Y=1.425 $X2=0 $Y2=0
cc_172 N_A_223_320#_c_179_n N_B_c_306_n 0.00137262f $X=3.42 $Y=2.015 $X2=0 $Y2=0
cc_173 N_A_223_320#_c_165_n N_B_c_306_n 0.00170917f $X=3.44 $Y=0.907 $X2=0 $Y2=0
cc_174 N_A_223_320#_c_170_n N_B_c_306_n 0.00274728f $X=3.56 $Y=1.425 $X2=0 $Y2=0
cc_175 N_A_223_320#_c_176_n N_A_M1011_g 0.00199767f $X=2.3 $Y=2.78 $X2=0 $Y2=0
cc_176 N_A_223_320#_c_178_n N_A_M1011_g 0.0180359f $X=2.385 $Y=2.675 $X2=0 $Y2=0
cc_177 N_A_223_320#_c_179_n N_A_M1011_g 0.00805279f $X=3.42 $Y=2.015 $X2=0 $Y2=0
cc_178 N_A_223_320#_c_180_n N_A_M1011_g 0.00391502f $X=2.47 $Y=2.015 $X2=0 $Y2=0
cc_179 N_A_223_320#_c_165_n N_A_c_389_n 0.00269921f $X=3.44 $Y=0.907 $X2=0 $Y2=0
cc_180 N_A_223_320#_c_165_n N_A_c_390_n 0.00742702f $X=3.44 $Y=0.907 $X2=0 $Y2=0
cc_181 N_A_223_320#_c_172_n N_A_c_390_n 0.0133616f $X=4.172 $Y=1.26 $X2=0 $Y2=0
cc_182 N_A_223_320#_M1001_g N_A_M1005_g 0.00541683f $X=4.295 $Y=2.465 $X2=0
+ $Y2=0
cc_183 N_A_223_320#_c_165_n N_A_M1005_g 0.00594375f $X=3.44 $Y=0.907 $X2=0 $Y2=0
cc_184 N_A_223_320#_c_166_n N_A_M1005_g 0.00453448f $X=3.53 $Y=1.26 $X2=0 $Y2=0
cc_185 N_A_223_320#_c_167_n N_A_M1005_g 0.00706087f $X=3.56 $Y=1.93 $X2=0 $Y2=0
cc_186 N_A_223_320#_c_168_n N_A_M1005_g 0.0135551f $X=4.14 $Y=1.425 $X2=0 $Y2=0
cc_187 N_A_223_320#_c_169_n N_A_M1005_g 0.0213545f $X=4.14 $Y=1.425 $X2=0 $Y2=0
cc_188 N_A_223_320#_c_170_n N_A_M1005_g 0.00745611f $X=3.56 $Y=1.425 $X2=0 $Y2=0
cc_189 N_A_223_320#_c_181_n N_A_M1000_g 0.00513831f $X=3.515 $Y=2.34 $X2=0 $Y2=0
cc_190 N_A_223_320#_c_183_n N_A_M1000_g 0.00263145f $X=3.55 $Y=2.015 $X2=0 $Y2=0
cc_191 N_A_223_320#_M1001_g N_A_c_399_n 0.0120108f $X=4.295 $Y=2.465 $X2=0 $Y2=0
cc_192 N_A_223_320#_c_167_n N_A_c_399_n 0.00209681f $X=3.56 $Y=1.93 $X2=0 $Y2=0
cc_193 N_A_223_320#_c_168_n N_A_c_399_n 0.00164608f $X=4.14 $Y=1.425 $X2=0 $Y2=0
cc_194 N_A_223_320#_c_183_n N_A_c_399_n 0.00213079f $X=3.55 $Y=2.015 $X2=0 $Y2=0
cc_195 N_A_223_320#_c_179_n A 0.0230841f $X=3.42 $Y=2.015 $X2=0 $Y2=0
cc_196 N_A_223_320#_c_180_n A 0.0124822f $X=2.47 $Y=2.015 $X2=0 $Y2=0
cc_197 N_A_223_320#_c_179_n N_A_c_394_n 0.00438376f $X=3.42 $Y=2.015 $X2=0 $Y2=0
cc_198 N_A_223_320#_c_165_n N_A_c_395_n 0.00124723f $X=3.44 $Y=0.907 $X2=0 $Y2=0
cc_199 N_A_223_320#_c_164_n N_VPWR_M1003_d 0.0110977f $X=1.28 $Y=1.765 $X2=-0.19
+ $Y2=-0.245
cc_200 N_A_223_320#_M1008_g N_VPWR_c_494_n 0.00128334f $X=1.5 $Y=2.35 $X2=0
+ $Y2=0
cc_201 N_A_223_320#_c_164_n N_VPWR_c_494_n 0.0660085f $X=1.28 $Y=1.765 $X2=0
+ $Y2=0
cc_202 N_A_223_320#_c_177_n N_VPWR_c_494_n 0.018451f $X=1.365 $Y=2.78 $X2=0
+ $Y2=0
cc_203 N_A_223_320#_c_171_n N_VPWR_c_494_n 0.00117087f $X=1.46 $Y=1.765 $X2=0
+ $Y2=0
cc_204 N_A_223_320#_c_176_n N_VPWR_c_495_n 0.0193623f $X=2.3 $Y=2.78 $X2=0 $Y2=0
cc_205 N_A_223_320#_c_178_n N_VPWR_c_495_n 0.0316866f $X=2.385 $Y=2.675 $X2=0
+ $Y2=0
cc_206 N_A_223_320#_c_179_n N_VPWR_c_495_n 0.0475186f $X=3.42 $Y=2.015 $X2=0
+ $Y2=0
cc_207 N_A_223_320#_M1001_g N_VPWR_c_496_n 0.0265739f $X=4.295 $Y=2.465 $X2=0
+ $Y2=0
cc_208 N_A_223_320#_c_181_n N_VPWR_c_496_n 0.0162695f $X=3.515 $Y=2.34 $X2=0
+ $Y2=0
cc_209 N_A_223_320#_c_167_n N_VPWR_c_496_n 0.00891608f $X=3.56 $Y=1.93 $X2=0
+ $Y2=0
cc_210 N_A_223_320#_c_168_n N_VPWR_c_496_n 0.0260167f $X=4.14 $Y=1.425 $X2=0
+ $Y2=0
cc_211 N_A_223_320#_c_169_n N_VPWR_c_496_n 0.00584123f $X=4.14 $Y=1.425 $X2=0
+ $Y2=0
cc_212 N_A_223_320#_c_183_n N_VPWR_c_496_n 0.0143601f $X=3.55 $Y=2.015 $X2=0
+ $Y2=0
cc_213 N_A_223_320#_M1008_g N_VPWR_c_499_n 4.99308e-19 $X=1.5 $Y=2.35 $X2=0
+ $Y2=0
cc_214 N_A_223_320#_c_176_n N_VPWR_c_499_n 0.0331204f $X=2.3 $Y=2.78 $X2=0 $Y2=0
cc_215 N_A_223_320#_c_177_n N_VPWR_c_499_n 0.00547657f $X=1.365 $Y=2.78 $X2=0
+ $Y2=0
cc_216 N_A_223_320#_M1001_g N_VPWR_c_501_n 0.00564095f $X=4.295 $Y=2.465 $X2=0
+ $Y2=0
cc_217 N_A_223_320#_M1001_g N_VPWR_c_493_n 0.0104427f $X=4.295 $Y=2.465 $X2=0
+ $Y2=0
cc_218 N_A_223_320#_c_176_n N_VPWR_c_493_n 0.0369964f $X=2.3 $Y=2.78 $X2=0 $Y2=0
cc_219 N_A_223_320#_c_177_n N_VPWR_c_493_n 0.00590738f $X=1.365 $Y=2.78 $X2=0
+ $Y2=0
cc_220 N_A_223_320#_c_181_n N_VPWR_c_493_n 0.0101636f $X=3.515 $Y=2.34 $X2=0
+ $Y2=0
cc_221 N_A_223_320#_c_178_n A_401_428# 0.00545531f $X=2.385 $Y=2.675 $X2=-0.19
+ $Y2=-0.245
cc_222 N_A_223_320#_c_168_n COUT 0.0274565f $X=4.14 $Y=1.425 $X2=0 $Y2=0
cc_223 N_A_223_320#_c_169_n COUT 0.0224678f $X=4.14 $Y=1.425 $X2=0 $Y2=0
cc_224 N_A_223_320#_c_172_n COUT 0.00615806f $X=4.172 $Y=1.26 $X2=0 $Y2=0
cc_225 N_A_223_320#_c_172_n N_COUT_c_554_n 0.00202488f $X=4.172 $Y=1.26 $X2=0
+ $Y2=0
cc_226 N_A_223_320#_c_169_n COUT 0.00162091f $X=4.14 $Y=1.425 $X2=0 $Y2=0
cc_227 N_A_223_320#_M1007_g N_VGND_c_569_n 0.00461526f $X=1.46 $Y=0.52 $X2=0
+ $Y2=0
cc_228 N_A_223_320#_M1007_g N_VGND_c_570_n 0.00106196f $X=1.46 $Y=0.52 $X2=0
+ $Y2=0
cc_229 N_A_223_320#_c_168_n N_VGND_c_571_n 0.0267028f $X=4.14 $Y=1.425 $X2=0
+ $Y2=0
cc_230 N_A_223_320#_c_169_n N_VGND_c_571_n 0.0036701f $X=4.14 $Y=1.425 $X2=0
+ $Y2=0
cc_231 N_A_223_320#_c_172_n N_VGND_c_571_n 0.014715f $X=4.172 $Y=1.26 $X2=0
+ $Y2=0
cc_232 N_A_223_320#_c_165_n N_VGND_c_572_n 0.00868768f $X=3.44 $Y=0.907 $X2=0
+ $Y2=0
cc_233 N_A_223_320#_M1007_g N_VGND_c_575_n 0.00512921f $X=1.46 $Y=0.52 $X2=0
+ $Y2=0
cc_234 N_A_223_320#_c_172_n N_VGND_c_576_n 0.00460072f $X=4.172 $Y=1.26 $X2=0
+ $Y2=0
cc_235 N_A_223_320#_M1007_g N_VGND_c_577_n 0.0108108f $X=1.46 $Y=0.52 $X2=0
+ $Y2=0
cc_236 N_A_223_320#_c_165_n N_VGND_c_577_n 0.0159622f $X=3.44 $Y=0.907 $X2=0
+ $Y2=0
cc_237 N_A_223_320#_c_172_n N_VGND_c_577_n 0.00910138f $X=4.172 $Y=1.26 $X2=0
+ $Y2=0
cc_238 N_A_223_320#_M1007_g N_A_307_62#_c_624_n 9.4255e-19 $X=1.46 $Y=0.52 $X2=0
+ $Y2=0
cc_239 N_A_223_320#_c_165_n N_A_307_62#_c_625_n 0.0125932f $X=3.44 $Y=0.907
+ $X2=0 $Y2=0
cc_240 N_A_223_320#_M1007_g N_A_307_62#_c_626_n 0.00152707f $X=1.46 $Y=0.52
+ $X2=0 $Y2=0
cc_241 N_A_223_320#_c_165_n N_A_307_62#_c_627_n 0.0060671f $X=3.44 $Y=0.907
+ $X2=0 $Y2=0
cc_242 N_A_223_320#_c_165_n A_675_146# 0.00245672f $X=3.44 $Y=0.907 $X2=-0.19
+ $Y2=-0.245
cc_243 N_A_223_320#_c_166_n A_675_146# 9.87179e-19 $X=3.53 $Y=1.26 $X2=-0.19
+ $Y2=-0.245
cc_244 N_B_M1012_g N_A_c_386_n 0.0185387f $X=1.89 $Y=0.52 $X2=-0.19 $Y2=-0.245
cc_245 N_B_M1002_g N_A_M1011_g 0.0218311f $X=1.93 $Y=2.35 $X2=0 $Y2=0
cc_246 N_B_M1006_g N_A_M1011_g 0.00818402f $X=3.3 $Y=2.35 $X2=0 $Y2=0
cc_247 N_B_c_310_n N_A_M1011_g 0.0132278f $X=1.98 $Y=1.9 $X2=0 $Y2=0
cc_248 N_B_c_302_n N_A_c_387_n 0.00747118f $X=2.96 $Y=1.315 $X2=0 $Y2=0
cc_249 N_B_c_302_n N_A_c_388_n 8.80528e-19 $X=2.96 $Y=1.315 $X2=0 $Y2=0
cc_250 N_B_c_299_n N_A_c_389_n 0.00901525f $X=3.3 $Y=1.26 $X2=0 $Y2=0
cc_251 N_B_c_299_n N_A_c_390_n 0.00855642f $X=3.3 $Y=1.26 $X2=0 $Y2=0
cc_252 N_B_c_299_n N_A_M1005_g 0.0357538f $X=3.3 $Y=1.26 $X2=0 $Y2=0
cc_253 N_B_c_305_n N_A_M1005_g 2.89108e-19 $X=3.12 $Y=1.425 $X2=0 $Y2=0
cc_254 N_B_M1006_g N_A_M1000_g 0.0135468f $X=3.3 $Y=2.35 $X2=0 $Y2=0
cc_255 N_B_c_306_n N_A_c_399_n 0.0357538f $X=3.3 $Y=1.425 $X2=0 $Y2=0
cc_256 N_B_M1006_g A 4.05191e-19 $X=3.3 $Y=2.35 $X2=0 $Y2=0
cc_257 N_B_c_301_n A 0.00117289f $X=1.98 $Y=1.735 $X2=0 $Y2=0
cc_258 N_B_c_302_n A 0.034245f $X=2.96 $Y=1.315 $X2=0 $Y2=0
cc_259 N_B_c_303_n A 0.0151037f $X=1.98 $Y=1.345 $X2=0 $Y2=0
cc_260 N_B_c_305_n A 0.0160164f $X=3.12 $Y=1.425 $X2=0 $Y2=0
cc_261 N_B_M1006_g N_A_c_394_n 0.00535252f $X=3.3 $Y=2.35 $X2=0 $Y2=0
cc_262 N_B_c_301_n N_A_c_394_n 0.0132278f $X=1.98 $Y=1.735 $X2=0 $Y2=0
cc_263 N_B_c_302_n N_A_c_394_n 0.00182961f $X=2.96 $Y=1.315 $X2=0 $Y2=0
cc_264 N_B_c_303_n N_A_c_394_n 8.32463e-19 $X=1.98 $Y=1.345 $X2=0 $Y2=0
cc_265 N_B_c_305_n N_A_c_394_n 0.00108143f $X=3.12 $Y=1.425 $X2=0 $Y2=0
cc_266 N_B_c_306_n N_A_c_394_n 0.00528225f $X=3.3 $Y=1.425 $X2=0 $Y2=0
cc_267 N_B_M1012_g N_A_c_395_n 0.00647268f $X=1.89 $Y=0.52 $X2=0 $Y2=0
cc_268 N_B_c_299_n N_A_c_395_n 0.00379313f $X=3.3 $Y=1.26 $X2=0 $Y2=0
cc_269 N_B_c_302_n N_A_c_395_n 0.0112772f $X=2.96 $Y=1.315 $X2=0 $Y2=0
cc_270 N_B_c_303_n N_A_c_395_n 0.00146699f $X=1.98 $Y=1.345 $X2=0 $Y2=0
cc_271 N_B_c_304_n N_A_c_395_n 0.0132278f $X=1.98 $Y=1.345 $X2=0 $Y2=0
cc_272 N_B_c_305_n N_A_c_395_n 5.56007e-19 $X=3.12 $Y=1.425 $X2=0 $Y2=0
cc_273 N_B_c_306_n N_A_c_395_n 0.00683264f $X=3.3 $Y=1.425 $X2=0 $Y2=0
cc_274 N_B_M1006_g N_VPWR_c_495_n 0.00931588f $X=3.3 $Y=2.35 $X2=0 $Y2=0
cc_275 N_B_M1002_g N_VPWR_c_499_n 4.99308e-19 $X=1.93 $Y=2.35 $X2=0 $Y2=0
cc_276 N_B_M1006_g N_VPWR_c_500_n 0.0028805f $X=3.3 $Y=2.35 $X2=0 $Y2=0
cc_277 N_B_M1006_g N_VPWR_c_493_n 0.00362163f $X=3.3 $Y=2.35 $X2=0 $Y2=0
cc_278 N_B_M1012_g N_VGND_c_570_n 0.00909521f $X=1.89 $Y=0.52 $X2=0 $Y2=0
cc_279 N_B_M1012_g N_VGND_c_575_n 0.00425877f $X=1.89 $Y=0.52 $X2=0 $Y2=0
cc_280 N_B_M1012_g N_VGND_c_577_n 0.00424416f $X=1.89 $Y=0.52 $X2=0 $Y2=0
cc_281 N_B_c_299_n N_VGND_c_577_n 8.36174e-19 $X=3.3 $Y=1.26 $X2=0 $Y2=0
cc_282 N_B_M1012_g N_A_307_62#_c_624_n 0.00157803f $X=1.89 $Y=0.52 $X2=0 $Y2=0
cc_283 N_B_M1012_g N_A_307_62#_c_625_n 0.0135398f $X=1.89 $Y=0.52 $X2=0 $Y2=0
cc_284 N_B_c_302_n N_A_307_62#_c_625_n 0.0355114f $X=2.96 $Y=1.315 $X2=0 $Y2=0
cc_285 N_B_c_303_n N_A_307_62#_c_625_n 0.0204544f $X=1.98 $Y=1.345 $X2=0 $Y2=0
cc_286 N_B_c_304_n N_A_307_62#_c_625_n 0.00125196f $X=1.98 $Y=1.345 $X2=0 $Y2=0
cc_287 N_A_M1011_g N_VPWR_c_495_n 0.00244614f $X=2.46 $Y=2.35 $X2=0 $Y2=0
cc_288 N_A_M1000_g N_VPWR_c_495_n 4.92982e-19 $X=3.73 $Y=2.35 $X2=0 $Y2=0
cc_289 N_A_c_399_n N_VPWR_c_496_n 0.0055923f $X=3.71 $Y=1.98 $X2=0 $Y2=0
cc_290 N_A_M1011_g N_VPWR_c_499_n 0.00178413f $X=2.46 $Y=2.35 $X2=0 $Y2=0
cc_291 N_A_M1000_g N_VPWR_c_500_n 0.0034649f $X=3.73 $Y=2.35 $X2=0 $Y2=0
cc_292 N_A_M1011_g N_VPWR_c_493_n 0.0018683f $X=2.46 $Y=2.35 $X2=0 $Y2=0
cc_293 N_A_M1000_g N_VPWR_c_493_n 0.00431146f $X=3.73 $Y=2.35 $X2=0 $Y2=0
cc_294 N_A_c_386_n N_VGND_c_570_n 0.00922324f $X=2.32 $Y=0.84 $X2=0 $Y2=0
cc_295 N_A_c_391_n N_VGND_c_570_n 9.68607e-19 $X=2.885 $Y=0.285 $X2=0 $Y2=0
cc_296 N_A_c_390_n N_VGND_c_571_n 0.0156873f $X=3.615 $Y=0.285 $X2=0 $Y2=0
cc_297 N_A_c_386_n N_VGND_c_572_n 0.00425877f $X=2.32 $Y=0.84 $X2=0 $Y2=0
cc_298 N_A_c_391_n N_VGND_c_572_n 0.0257186f $X=2.885 $Y=0.285 $X2=0 $Y2=0
cc_299 N_A_c_386_n N_VGND_c_577_n 0.00457129f $X=2.32 $Y=0.84 $X2=0 $Y2=0
cc_300 N_A_c_390_n N_VGND_c_577_n 0.0311405f $X=3.615 $Y=0.285 $X2=0 $Y2=0
cc_301 N_A_c_391_n N_VGND_c_577_n 0.0094611f $X=2.885 $Y=0.285 $X2=0 $Y2=0
cc_302 N_A_c_387_n N_A_307_62#_c_625_n 0.00763828f $X=2.735 $Y=0.915 $X2=0 $Y2=0
cc_303 N_A_c_388_n N_A_307_62#_c_625_n 0.0132743f $X=2.535 $Y=0.915 $X2=0 $Y2=0
cc_304 N_A_c_395_n N_A_307_62#_c_625_n 0.00322408f $X=2.55 $Y=1.5 $X2=0 $Y2=0
cc_305 N_A_c_386_n N_A_307_62#_c_627_n 0.0017013f $X=2.32 $Y=0.84 $X2=0 $Y2=0
cc_306 N_A_c_391_n N_A_307_62#_c_627_n 0.0117389f $X=2.885 $Y=0.285 $X2=0 $Y2=0
cc_307 SUM N_VPWR_c_494_n 0.00133185f $X=0.155 $Y=1.58 $X2=0 $Y2=0
cc_308 N_SUM_c_480_n N_VPWR_c_497_n 0.028202f $X=0.4 $Y=1.98 $X2=0 $Y2=0
cc_309 N_SUM_M1003_s N_VPWR_c_493_n 0.00336915f $X=0.275 $Y=1.835 $X2=0 $Y2=0
cc_310 N_SUM_c_480_n N_VPWR_c_493_n 0.0158621f $X=0.4 $Y=1.98 $X2=0 $Y2=0
cc_311 N_SUM_c_477_n N_VGND_c_569_n 0.0306436f $X=0.26 $Y=0.425 $X2=0 $Y2=0
cc_312 N_SUM_c_477_n N_VGND_c_574_n 0.0186238f $X=0.26 $Y=0.425 $X2=0 $Y2=0
cc_313 N_SUM_c_477_n N_VGND_c_577_n 0.0103947f $X=0.26 $Y=0.425 $X2=0 $Y2=0
cc_314 N_VPWR_c_493_n N_COUT_M1001_d 0.00302127f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_315 N_VPWR_c_496_n COUT 0.0489991f $X=4.08 $Y=1.98 $X2=0 $Y2=0
cc_316 N_VPWR_c_501_n COUT 0.0213882f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_317 N_VPWR_c_493_n COUT 0.0123631f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_318 N_COUT_c_554_n N_VGND_c_571_n 0.0312953f $X=4.43 $Y=0.455 $X2=0 $Y2=0
cc_319 N_COUT_c_554_n N_VGND_c_576_n 0.0227613f $X=4.43 $Y=0.455 $X2=0 $Y2=0
cc_320 N_COUT_c_554_n N_VGND_c_577_n 0.0148244f $X=4.43 $Y=0.455 $X2=0 $Y2=0
cc_321 N_VGND_c_575_n N_A_307_62#_c_624_n 0.00843997f $X=1.94 $Y=0 $X2=0 $Y2=0
cc_322 N_VGND_c_577_n N_A_307_62#_c_624_n 0.00838461f $X=4.56 $Y=0 $X2=0 $Y2=0
cc_323 N_VGND_c_570_n N_A_307_62#_c_625_n 0.0210115f $X=2.105 $Y=0.52 $X2=0
+ $Y2=0
cc_324 N_VGND_c_577_n N_A_307_62#_c_625_n 0.0108697f $X=4.56 $Y=0 $X2=0 $Y2=0
cc_325 N_VGND_c_572_n N_A_307_62#_c_627_n 0.0107764f $X=3.79 $Y=0 $X2=0 $Y2=0
cc_326 N_VGND_c_577_n N_A_307_62#_c_627_n 0.00948785f $X=4.56 $Y=0 $X2=0 $Y2=0
