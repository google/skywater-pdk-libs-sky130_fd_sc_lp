* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
X0 X a_84_28# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X1 VGND A1 a_494_51# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X2 a_84_28# A2 a_584_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X3 a_84_28# a_281_138# a_494_51# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X4 VGND B1_N a_281_138# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 a_494_51# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X6 X a_84_28# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X7 VPWR B1_N a_281_138# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X8 a_584_367# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X9 VPWR a_281_138# a_84_28# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
.ends
