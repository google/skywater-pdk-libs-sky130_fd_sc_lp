# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__o21bai_2
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__o21bai_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.320000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.015000 1.425000 2.580000 1.920000 ;
        RECT 2.015000 1.920000 3.695000 2.120000 ;
        RECT 3.515000 1.425000 3.990000 1.645000 ;
        RECT 3.515000 1.645000 3.695000 1.920000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.800000 1.425000 3.345000 1.750000 ;
    END
  END A2
  PIN B1_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.840000 0.425000 1.510000 ;
    END
  END B1_N
  PIN Y
    ANTENNADIFFAREA  0.940800 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.555000 0.595000 1.885000 1.145000 ;
        RECT 1.595000 1.815000 1.845000 2.290000 ;
        RECT 1.595000 2.290000 3.185000 2.620000 ;
        RECT 1.595000 2.620000 1.825000 3.075000 ;
        RECT 1.625000 1.145000 1.845000 1.815000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.320000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.320000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.320000 0.085000 ;
      RECT 0.000000  3.245000 4.320000 3.415000 ;
      RECT 0.095000  0.085000 0.425000 0.670000 ;
      RECT 0.460000  1.755000 0.795000 2.210000 ;
      RECT 0.595000  0.355000 0.855000 1.355000 ;
      RECT 0.595000  1.355000 1.455000 1.605000 ;
      RECT 0.595000  1.605000 0.795000 1.755000 ;
      RECT 0.965000  1.815000 1.425000 3.245000 ;
      RECT 1.125000  0.255000 2.265000 0.425000 ;
      RECT 1.125000  0.425000 1.375000 1.185000 ;
      RECT 1.995000  2.790000 2.325000 3.245000 ;
      RECT 2.065000  0.425000 2.265000 1.085000 ;
      RECT 2.065000  1.085000 4.135000 1.255000 ;
      RECT 2.435000  0.085000 2.765000 0.915000 ;
      RECT 2.495000  2.800000 3.685000 3.075000 ;
      RECT 2.935000  0.305000 3.185000 1.085000 ;
      RECT 3.355000  0.085000 3.685000 0.915000 ;
      RECT 3.355000  2.290000 3.685000 2.800000 ;
      RECT 3.855000  0.305000 4.135000 1.085000 ;
      RECT 3.865000  1.815000 4.115000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
  END
END sky130_fd_sc_lp__o21bai_2
END LIBRARY
