# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__nand4b_4
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__nand4b_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.120000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A_N
    ANTENNAGATEAREA  0.315000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 1.365000 0.435000 1.760000 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.010000 1.425000 4.700000 1.605000 ;
        RECT 3.845000 1.605000 4.700000 1.780000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.230000 1.425000 6.920000 1.595000 ;
        RECT 5.230000 1.595000 6.085000 1.750000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.210000 1.425000 9.020000 1.595000 ;
        RECT 7.785000 1.595000 9.020000 1.750000 ;
    END
  END D
  PIN Y
    ANTENNADIFFAREA  3.292800 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.345000 1.775000 3.670000 1.945000 ;
        RECT 1.345000 1.945000 1.615000 3.075000 ;
        RECT 1.510000 0.595000 1.735000 1.075000 ;
        RECT 1.510000 1.075000 5.050000 1.255000 ;
        RECT 2.285000 1.945000 2.515000 3.075000 ;
        RECT 2.405000 0.595000 2.595000 1.075000 ;
        RECT 3.185000 1.945000 3.670000 1.950000 ;
        RECT 3.185000 1.950000 6.425000 2.120000 ;
        RECT 3.185000 2.120000 3.395000 3.075000 ;
        RECT 4.065000 2.120000 4.255000 3.075000 ;
        RECT 4.880000 1.255000 5.050000 1.920000 ;
        RECT 4.880000 1.920000 7.615000 1.930000 ;
        RECT 4.880000 1.930000 8.405000 1.935000 ;
        RECT 4.880000 1.935000 6.425000 1.950000 ;
        RECT 5.265000 2.120000 5.455000 3.075000 ;
        RECT 6.125000 2.120000 6.425000 3.075000 ;
        RECT 6.255000 1.765000 7.615000 1.920000 ;
        RECT 7.355000 1.935000 8.405000 2.100000 ;
        RECT 7.355000 2.100000 7.535000 3.075000 ;
        RECT 8.215000 2.100000 8.405000 3.075000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 9.120000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 9.120000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 9.120000 0.085000 ;
      RECT 0.000000  3.245000 9.120000 3.415000 ;
      RECT 0.095000  0.255000 0.345000 1.025000 ;
      RECT 0.095000  1.025000 0.855000 1.195000 ;
      RECT 0.445000  1.930000 0.775000 3.075000 ;
      RECT 0.525000  0.085000 0.855000 0.855000 ;
      RECT 0.605000  1.195000 0.855000 1.425000 ;
      RECT 0.605000  1.425000 2.800000 1.595000 ;
      RECT 0.605000  1.595000 0.775000 1.930000 ;
      RECT 0.945000  1.815000 1.175000 3.245000 ;
      RECT 1.045000  0.255000 4.895000 0.425000 ;
      RECT 1.045000  0.425000 1.340000 1.115000 ;
      RECT 1.785000  2.125000 2.115000 3.245000 ;
      RECT 1.905000  0.425000 2.235000 0.905000 ;
      RECT 2.685000  2.115000 3.015000 3.245000 ;
      RECT 2.765000  0.425000 4.895000 0.515000 ;
      RECT 2.765000  0.515000 3.095000 0.905000 ;
      RECT 3.275000  0.685000 4.465000 0.725000 ;
      RECT 3.275000  0.725000 5.795000 0.905000 ;
      RECT 3.565000  2.290000 3.895000 3.245000 ;
      RECT 4.425000  2.290000 5.095000 3.245000 ;
      RECT 5.105000  0.255000 7.165000 0.435000 ;
      RECT 5.105000  0.435000 6.295000 0.555000 ;
      RECT 5.530000  0.905000 5.795000 1.075000 ;
      RECT 5.530000  1.075000 6.805000 1.255000 ;
      RECT 5.625000  2.290000 5.955000 3.245000 ;
      RECT 5.965000  0.555000 6.295000 0.905000 ;
      RECT 6.475000  0.605000 6.805000 1.075000 ;
      RECT 6.595000  2.105000 7.185000 3.245000 ;
      RECT 6.975000  0.435000 7.165000 1.075000 ;
      RECT 6.975000  1.075000 8.955000 1.245000 ;
      RECT 7.335000  0.085000 7.665000 0.905000 ;
      RECT 7.715000  2.270000 8.045000 3.245000 ;
      RECT 7.835000  0.305000 8.025000 1.075000 ;
      RECT 8.195000  0.085000 8.525000 0.895000 ;
      RECT 8.575000  1.920000 8.905000 3.245000 ;
      RECT 8.695000  0.305000 8.955000 1.075000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
      RECT 8.315000 -0.085000 8.485000 0.085000 ;
      RECT 8.315000  3.245000 8.485000 3.415000 ;
      RECT 8.795000 -0.085000 8.965000 0.085000 ;
      RECT 8.795000  3.245000 8.965000 3.415000 ;
  END
END sky130_fd_sc_lp__nand4b_4
END LIBRARY
