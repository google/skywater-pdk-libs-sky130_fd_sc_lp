* NGSPICE file created from sky130_fd_sc_lp__nor2b_m.ext - technology: sky130A

.subckt sky130_fd_sc_lp__nor2b_m A B_N VGND VNB VPB VPWR Y
M1000 Y a_47_70# a_328_492# VPB phighvt w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=8.82e+10p ps=1.26e+06u
M1001 a_328_492# A VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.827e+11p ps=1.71e+06u
M1002 VGND a_47_70# Y VNB nshort w=420000u l=150000u
+  ad=3.549e+11p pd=3.37e+06u as=1.176e+11p ps=1.4e+06u
M1003 VGND B_N a_47_70# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1004 VPWR B_N a_47_70# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1005 Y A VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

