* File: sky130_fd_sc_lp__nor4b_4.pex.spice
* Created: Wed Sep  2 10:11:09 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__NOR4B_4%D_N 3 7 9 12 13
r31 12 15 46.3065 $w=3.4e-07 $l=1.65e-07 $layer=POLY_cond $X=0.39 $Y=1.46
+ $X2=0.39 $Y2=1.625
r32 12 14 46.3065 $w=3.4e-07 $l=1.65e-07 $layer=POLY_cond $X=0.39 $Y=1.46
+ $X2=0.39 $Y2=1.295
r33 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.385
+ $Y=1.46 $X2=0.385 $Y2=1.46
r34 9 13 5.27303 $w=4.63e-07 $l=2.05e-07 $layer=LI1_cond $X=0.317 $Y=1.665
+ $X2=0.317 $Y2=1.46
r35 7 14 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=0.485 $Y=0.655
+ $X2=0.485 $Y2=1.295
r36 3 15 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=0.475 $Y=2.465
+ $X2=0.475 $Y2=1.625
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4B_4%A_27_367# 1 2 9 13 17 21 25 29 33 37 39 41
+ 45 47 49 50 52 54 60 65 76
r127 73 74 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=2.285 $Y=1.4
+ $X2=2.305 $Y2=1.4
r128 72 73 71.6931 $w=3.3e-07 $l=4.1e-07 $layer=POLY_cond $X=1.875 $Y=1.4
+ $X2=2.285 $Y2=1.4
r129 71 72 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=1.855 $Y=1.4
+ $X2=1.875 $Y2=1.4
r130 70 71 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=1.425 $Y=1.4
+ $X2=1.855 $Y2=1.4
r131 69 70 5.24584 $w=3.3e-07 $l=3e-08 $layer=POLY_cond $X=1.395 $Y=1.4
+ $X2=1.425 $Y2=1.4
r132 68 69 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=0.965 $Y=1.4
+ $X2=1.395 $Y2=1.4
r133 61 76 13.9889 $w=3.3e-07 $l=8e-08 $layer=POLY_cond $X=2.635 $Y=1.4
+ $X2=2.715 $Y2=1.4
r134 61 74 57.7042 $w=3.3e-07 $l=3.3e-07 $layer=POLY_cond $X=2.635 $Y=1.4
+ $X2=2.305 $Y2=1.4
r135 60 61 48.4267 $w=1.7e-07 $l=5.1e-07 $layer=licon1_POLY $count=3 $X=2.635
+ $Y=1.4 $X2=2.635 $Y2=1.4
r136 58 68 5.24584 $w=3.3e-07 $l=3e-08 $layer=POLY_cond $X=0.935 $Y=1.4
+ $X2=0.965 $Y2=1.4
r137 57 60 110.909 $w=1.68e-07 $l=1.7e-06 $layer=LI1_cond $X=0.935 $Y=1.4
+ $X2=2.635 $Y2=1.4
r138 57 58 48.4267 $w=1.7e-07 $l=5.1e-07 $layer=licon1_POLY $count=3 $X=0.935
+ $Y=1.4 $X2=0.935 $Y2=1.4
r139 55 65 2.0246 $w=1.7e-07 $l=1.03e-07 $layer=LI1_cond $X=0.925 $Y=1.4
+ $X2=0.822 $Y2=1.4
r140 55 57 0.652406 $w=1.68e-07 $l=1e-08 $layer=LI1_cond $X=0.925 $Y=1.4
+ $X2=0.935 $Y2=1.4
r141 53 65 4.40882 $w=2.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.822 $Y=1.485
+ $X2=0.822 $Y2=1.4
r142 53 54 24.0754 $w=2.03e-07 $l=4.45e-07 $layer=LI1_cond $X=0.822 $Y=1.485
+ $X2=0.822 $Y2=1.93
r143 52 65 4.40882 $w=2.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.822 $Y=1.315
+ $X2=0.822 $Y2=1.4
r144 51 52 8.65632 $w=2.03e-07 $l=1.6e-07 $layer=LI1_cond $X=0.822 $Y=1.155
+ $X2=0.822 $Y2=1.315
r145 49 51 6.89401 $w=1.7e-07 $l=1.38109e-07 $layer=LI1_cond $X=0.72 $Y=1.07
+ $X2=0.822 $Y2=1.155
r146 49 50 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=0.72 $Y=1.07
+ $X2=0.365 $Y2=1.07
r147 48 64 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.355 $Y=2.015
+ $X2=0.225 $Y2=2.015
r148 47 54 6.89401 $w=1.7e-07 $l=1.38109e-07 $layer=LI1_cond $X=0.72 $Y=2.015
+ $X2=0.822 $Y2=1.93
r149 47 48 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.72 $Y=2.015
+ $X2=0.355 $Y2=2.015
r150 43 50 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=0.235 $Y=0.985
+ $X2=0.365 $Y2=1.07
r151 43 45 25.0435 $w=2.58e-07 $l=5.65e-07 $layer=LI1_cond $X=0.235 $Y=0.985
+ $X2=0.235 $Y2=0.42
r152 39 64 2.85134 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=0.225 $Y=2.1
+ $X2=0.225 $Y2=2.015
r153 39 41 35.903 $w=2.58e-07 $l=8.1e-07 $layer=LI1_cond $X=0.225 $Y=2.1
+ $X2=0.225 $Y2=2.91
r154 35 76 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.715 $Y=1.565
+ $X2=2.715 $Y2=1.4
r155 35 37 461.489 $w=1.5e-07 $l=9e-07 $layer=POLY_cond $X=2.715 $Y=1.565
+ $X2=2.715 $Y2=2.465
r156 31 74 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.305 $Y=1.235
+ $X2=2.305 $Y2=1.4
r157 31 33 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=2.305 $Y=1.235
+ $X2=2.305 $Y2=0.655
r158 27 73 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.285 $Y=1.565
+ $X2=2.285 $Y2=1.4
r159 27 29 461.489 $w=1.5e-07 $l=9e-07 $layer=POLY_cond $X=2.285 $Y=1.565
+ $X2=2.285 $Y2=2.465
r160 23 72 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.875 $Y=1.235
+ $X2=1.875 $Y2=1.4
r161 23 25 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=1.875 $Y=1.235
+ $X2=1.875 $Y2=0.655
r162 19 71 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.855 $Y=1.565
+ $X2=1.855 $Y2=1.4
r163 19 21 461.489 $w=1.5e-07 $l=9e-07 $layer=POLY_cond $X=1.855 $Y=1.565
+ $X2=1.855 $Y2=2.465
r164 15 70 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.425 $Y=1.565
+ $X2=1.425 $Y2=1.4
r165 15 17 461.489 $w=1.5e-07 $l=9e-07 $layer=POLY_cond $X=1.425 $Y=1.565
+ $X2=1.425 $Y2=2.465
r166 11 69 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.395 $Y=1.235
+ $X2=1.395 $Y2=1.4
r167 11 13 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=1.395 $Y=1.235
+ $X2=1.395 $Y2=0.655
r168 7 68 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.965 $Y=1.235
+ $X2=0.965 $Y2=1.4
r169 7 9 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=0.965 $Y=1.235
+ $X2=0.965 $Y2=0.655
r170 2 64 400 $w=1.7e-07 $l=3.16386e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.835 $X2=0.26 $Y2=2.095
r171 2 41 400 $w=1.7e-07 $l=1.13578e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.835 $X2=0.26 $Y2=2.91
r172 1 45 91 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=2 $X=0.145
+ $Y=0.235 $X2=0.27 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4B_4%C 3 7 11 15 19 23 27 31 41 42 61 64 66 74
r87 64 66 2.43061 $w=2.73e-07 $l=5.8e-08 $layer=LI1_cond $X=4.022 $Y=1.347
+ $X2=4.08 $Y2=1.347
r88 61 62 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.535
+ $Y=1.4 $X2=4.535 $Y2=1.4
r89 59 61 17.4861 $w=3.3e-07 $l=1e-07 $layer=POLY_cond $X=4.435 $Y=1.4 $X2=4.535
+ $Y2=1.4
r90 58 59 10.4917 $w=3.3e-07 $l=6e-08 $layer=POLY_cond $X=4.375 $Y=1.4 $X2=4.435
+ $Y2=1.4
r91 57 62 14.2484 $w=2.73e-07 $l=3.4e-07 $layer=LI1_cond $X=4.195 $Y=1.347
+ $X2=4.535 $Y2=1.347
r92 56 58 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=4.195 $Y=1.4
+ $X2=4.375 $Y2=1.4
r93 56 57 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.195
+ $Y=1.4 $X2=4.195 $Y2=1.4
r94 54 56 33.2236 $w=3.3e-07 $l=1.9e-07 $layer=POLY_cond $X=4.005 $Y=1.4
+ $X2=4.195 $Y2=1.4
r95 53 54 10.4917 $w=3.3e-07 $l=6e-08 $layer=POLY_cond $X=3.945 $Y=1.4 $X2=4.005
+ $Y2=1.4
r96 50 51 10.4917 $w=3.3e-07 $l=6e-08 $layer=POLY_cond $X=3.515 $Y=1.4 $X2=3.575
+ $Y2=1.4
r97 46 48 10.4917 $w=3.3e-07 $l=6e-08 $layer=POLY_cond $X=3.085 $Y=1.4 $X2=3.145
+ $Y2=1.4
r98 42 62 1.04768 $w=2.73e-07 $l=2.5e-08 $layer=LI1_cond $X=4.56 $Y=1.347
+ $X2=4.535 $Y2=1.347
r99 41 64 0.586698 $w=2.73e-07 $l=1.4e-08 $layer=LI1_cond $X=4.008 $Y=1.347
+ $X2=4.022 $Y2=1.347
r100 41 74 6.82415 $w=2.73e-07 $l=1.23e-07 $layer=LI1_cond $X=4.008 $Y=1.347
+ $X2=3.885 $Y2=1.347
r101 41 57 4.27452 $w=2.73e-07 $l=1.02e-07 $layer=LI1_cond $X=4.093 $Y=1.347
+ $X2=4.195 $Y2=1.347
r102 41 66 0.544791 $w=2.73e-07 $l=1.3e-08 $layer=LI1_cond $X=4.093 $Y=1.347
+ $X2=4.08 $Y2=1.347
r103 40 53 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=3.855 $Y=1.4
+ $X2=3.945 $Y2=1.4
r104 40 51 48.9612 $w=3.3e-07 $l=2.8e-07 $layer=POLY_cond $X=3.855 $Y=1.4
+ $X2=3.575 $Y2=1.4
r105 39 74 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=3.855 $Y=1.4
+ $X2=3.885 $Y2=1.4
r106 39 40 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=3.855
+ $Y=1.4 $X2=3.855 $Y2=1.4
r107 36 50 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=3.175 $Y=1.4
+ $X2=3.515 $Y2=1.4
r108 36 48 5.24584 $w=3.3e-07 $l=3e-08 $layer=POLY_cond $X=3.175 $Y=1.4
+ $X2=3.145 $Y2=1.4
r109 35 39 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=3.175 $Y=1.4
+ $X2=3.855 $Y2=1.4
r110 35 36 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=3.175
+ $Y=1.4 $X2=3.175 $Y2=1.4
r111 29 59 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.435 $Y=1.565
+ $X2=4.435 $Y2=1.4
r112 29 31 461.489 $w=1.5e-07 $l=9e-07 $layer=POLY_cond $X=4.435 $Y=1.565
+ $X2=4.435 $Y2=2.465
r113 25 58 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.375 $Y=1.235
+ $X2=4.375 $Y2=1.4
r114 25 27 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=4.375 $Y=1.235
+ $X2=4.375 $Y2=0.655
r115 21 54 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.005 $Y=1.565
+ $X2=4.005 $Y2=1.4
r116 21 23 461.489 $w=1.5e-07 $l=9e-07 $layer=POLY_cond $X=4.005 $Y=1.565
+ $X2=4.005 $Y2=2.465
r117 17 53 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.945 $Y=1.235
+ $X2=3.945 $Y2=1.4
r118 17 19 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=3.945 $Y=1.235
+ $X2=3.945 $Y2=0.655
r119 13 51 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.575 $Y=1.565
+ $X2=3.575 $Y2=1.4
r120 13 15 461.489 $w=1.5e-07 $l=9e-07 $layer=POLY_cond $X=3.575 $Y=1.565
+ $X2=3.575 $Y2=2.465
r121 9 50 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.515 $Y=1.235
+ $X2=3.515 $Y2=1.4
r122 9 11 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=3.515 $Y=1.235
+ $X2=3.515 $Y2=0.655
r123 5 48 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.145 $Y=1.565
+ $X2=3.145 $Y2=1.4
r124 5 7 461.489 $w=1.5e-07 $l=9e-07 $layer=POLY_cond $X=3.145 $Y=1.565
+ $X2=3.145 $Y2=2.465
r125 1 46 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.085 $Y=1.235
+ $X2=3.085 $Y2=1.4
r126 1 3 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=3.085 $Y=1.235
+ $X2=3.085 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4B_4%B 3 7 11 15 19 23 27 31 33 34 35 53
c88 53 0 5.10287e-20 $X=6.675 $Y=1.51
r89 52 53 13.9889 $w=3.3e-07 $l=8e-08 $layer=POLY_cond $X=6.595 $Y=1.51
+ $X2=6.675 $Y2=1.51
r90 50 52 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=6.415 $Y=1.51
+ $X2=6.595 $Y2=1.51
r91 50 51 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.415
+ $Y=1.51 $X2=6.415 $Y2=1.51
r92 48 50 29.7264 $w=3.3e-07 $l=1.7e-07 $layer=POLY_cond $X=6.245 $Y=1.51
+ $X2=6.415 $Y2=1.51
r93 47 48 13.9889 $w=3.3e-07 $l=8e-08 $layer=POLY_cond $X=6.165 $Y=1.51
+ $X2=6.245 $Y2=1.51
r94 46 47 61.2015 $w=3.3e-07 $l=3.5e-07 $layer=POLY_cond $X=5.815 $Y=1.51
+ $X2=6.165 $Y2=1.51
r95 45 46 13.9889 $w=3.3e-07 $l=8e-08 $layer=POLY_cond $X=5.735 $Y=1.51
+ $X2=5.815 $Y2=1.51
r96 43 45 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=5.395 $Y=1.51
+ $X2=5.735 $Y2=1.51
r97 43 44 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.395
+ $Y=1.51 $X2=5.395 $Y2=1.51
r98 41 43 1.74861 $w=3.3e-07 $l=1e-08 $layer=POLY_cond $X=5.385 $Y=1.51
+ $X2=5.395 $Y2=1.51
r99 39 41 13.9889 $w=3.3e-07 $l=8e-08 $layer=POLY_cond $X=5.305 $Y=1.51
+ $X2=5.385 $Y2=1.51
r100 35 51 1.61969 $w=4.78e-07 $l=6.5e-08 $layer=LI1_cond $X=6.48 $Y=1.595
+ $X2=6.415 $Y2=1.595
r101 34 51 10.3411 $w=4.78e-07 $l=4.15e-07 $layer=LI1_cond $X=6 $Y=1.595
+ $X2=6.415 $Y2=1.595
r102 33 34 11.9608 $w=4.78e-07 $l=4.8e-07 $layer=LI1_cond $X=5.52 $Y=1.595 $X2=6
+ $Y2=1.595
r103 33 44 3.11479 $w=4.78e-07 $l=1.25e-07 $layer=LI1_cond $X=5.52 $Y=1.595
+ $X2=5.395 $Y2=1.595
r104 29 53 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.675 $Y=1.675
+ $X2=6.675 $Y2=1.51
r105 29 31 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=6.675 $Y=1.675
+ $X2=6.675 $Y2=2.465
r106 25 52 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.595 $Y=1.345
+ $X2=6.595 $Y2=1.51
r107 25 27 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=6.595 $Y=1.345
+ $X2=6.595 $Y2=0.655
r108 21 48 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.245 $Y=1.675
+ $X2=6.245 $Y2=1.51
r109 21 23 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=6.245 $Y=1.675
+ $X2=6.245 $Y2=2.465
r110 17 47 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.165 $Y=1.345
+ $X2=6.165 $Y2=1.51
r111 17 19 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=6.165 $Y=1.345
+ $X2=6.165 $Y2=0.655
r112 13 46 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.815 $Y=1.675
+ $X2=5.815 $Y2=1.51
r113 13 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=5.815 $Y=1.675
+ $X2=5.815 $Y2=2.465
r114 9 45 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.735 $Y=1.345
+ $X2=5.735 $Y2=1.51
r115 9 11 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=5.735 $Y=1.345
+ $X2=5.735 $Y2=0.655
r116 5 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.385 $Y=1.675
+ $X2=5.385 $Y2=1.51
r117 5 7 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=5.385 $Y=1.675
+ $X2=5.385 $Y2=2.465
r118 1 39 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.305 $Y=1.345
+ $X2=5.305 $Y2=1.51
r119 1 3 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=5.305 $Y=1.345
+ $X2=5.305 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4B_4%A 3 7 11 15 19 23 27 31 38 39 40 45 47 66 68
+ 78
c83 11 0 8.13651e-20 $X=7.495 $Y=0.655
r84 66 68 1.02439 $w=3.13e-07 $l=2.8e-08 $layer=LI1_cond $X=7.892 $Y=1.367
+ $X2=7.92 $Y2=1.367
r85 64 65 6.99445 $w=3.3e-07 $l=4e-08 $layer=POLY_cond $X=8.355 $Y=1.44
+ $X2=8.395 $Y2=1.44
r86 62 64 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=8.145 $Y=1.44
+ $X2=8.355 $Y2=1.44
r87 62 63 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.145
+ $Y=1.44 $X2=8.145 $Y2=1.44
r88 60 62 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=7.965 $Y=1.44
+ $X2=8.145 $Y2=1.44
r89 59 60 6.99445 $w=3.3e-07 $l=4e-08 $layer=POLY_cond $X=7.925 $Y=1.44
+ $X2=7.965 $Y2=1.44
r90 58 78 4.98695 $w=3.13e-07 $l=7e-08 $layer=LI1_cond $X=7.805 $Y=1.367
+ $X2=7.735 $Y2=1.367
r91 57 59 20.9834 $w=3.3e-07 $l=1.2e-07 $layer=POLY_cond $X=7.805 $Y=1.44
+ $X2=7.925 $Y2=1.44
r92 57 58 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=7.805
+ $Y=1.44 $X2=7.805 $Y2=1.44
r93 55 57 47.2125 $w=3.3e-07 $l=2.7e-07 $layer=POLY_cond $X=7.535 $Y=1.44
+ $X2=7.805 $Y2=1.44
r94 54 55 6.99445 $w=3.3e-07 $l=4e-08 $layer=POLY_cond $X=7.495 $Y=1.44
+ $X2=7.535 $Y2=1.44
r95 50 52 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=7.035 $Y=1.44
+ $X2=7.105 $Y2=1.44
r96 47 48 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=8.825
+ $Y=1.44 $X2=8.825 $Y2=1.44
r97 45 65 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=8.47 $Y=1.44
+ $X2=8.395 $Y2=1.44
r98 45 47 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=8.47 $Y=1.44
+ $X2=8.825 $Y2=1.44
r99 40 48 2.0122 $w=3.13e-07 $l=5.5e-08 $layer=LI1_cond $X=8.88 $Y=1.367
+ $X2=8.825 $Y2=1.367
r100 39 48 15.5488 $w=3.13e-07 $l=4.25e-07 $layer=LI1_cond $X=8.4 $Y=1.367
+ $X2=8.825 $Y2=1.367
r101 39 63 9.3293 $w=3.13e-07 $l=2.55e-07 $layer=LI1_cond $X=8.4 $Y=1.367
+ $X2=8.145 $Y2=1.367
r102 38 66 1.06098 $w=3.13e-07 $l=2.9e-08 $layer=LI1_cond $X=7.863 $Y=1.367
+ $X2=7.892 $Y2=1.367
r103 38 58 2.12196 $w=3.13e-07 $l=5.8e-08 $layer=LI1_cond $X=7.863 $Y=1.367
+ $X2=7.805 $Y2=1.367
r104 38 63 7.20734 $w=3.13e-07 $l=1.97e-07 $layer=LI1_cond $X=7.948 $Y=1.367
+ $X2=8.145 $Y2=1.367
r105 38 68 1.02439 $w=3.13e-07 $l=2.8e-08 $layer=LI1_cond $X=7.948 $Y=1.367
+ $X2=7.92 $Y2=1.367
r106 36 54 64.6987 $w=3.3e-07 $l=3.7e-07 $layer=POLY_cond $X=7.125 $Y=1.44
+ $X2=7.495 $Y2=1.44
r107 36 52 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=7.125 $Y=1.44
+ $X2=7.105 $Y2=1.44
r108 35 78 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=7.125 $Y=1.44
+ $X2=7.735 $Y2=1.44
r109 35 36 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=7.125
+ $Y=1.44 $X2=7.125 $Y2=1.44
r110 29 65 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.395 $Y=1.605
+ $X2=8.395 $Y2=1.44
r111 29 31 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=8.395 $Y=1.605
+ $X2=8.395 $Y2=2.465
r112 25 64 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.355 $Y=1.275
+ $X2=8.355 $Y2=1.44
r113 25 27 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=8.355 $Y=1.275
+ $X2=8.355 $Y2=0.655
r114 21 60 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.965 $Y=1.605
+ $X2=7.965 $Y2=1.44
r115 21 23 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=7.965 $Y=1.605
+ $X2=7.965 $Y2=2.465
r116 17 59 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.925 $Y=1.275
+ $X2=7.925 $Y2=1.44
r117 17 19 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=7.925 $Y=1.275
+ $X2=7.925 $Y2=0.655
r118 13 55 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.535 $Y=1.605
+ $X2=7.535 $Y2=1.44
r119 13 15 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=7.535 $Y=1.605
+ $X2=7.535 $Y2=2.465
r120 9 54 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.495 $Y=1.275
+ $X2=7.495 $Y2=1.44
r121 9 11 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=7.495 $Y=1.275
+ $X2=7.495 $Y2=0.655
r122 5 52 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.105 $Y=1.605
+ $X2=7.105 $Y2=1.44
r123 5 7 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=7.105 $Y=1.605
+ $X2=7.105 $Y2=2.465
r124 1 50 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.035 $Y=1.275
+ $X2=7.035 $Y2=1.44
r125 1 3 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=7.035 $Y=1.275
+ $X2=7.035 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4B_4%VPWR 1 2 3 12 16 22 27 28 30 31 32 34 50 51
+ 54
r113 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r114 50 51 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r115 48 51 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=8.88 $Y2=3.33
r116 47 48 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r117 45 48 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=7.92 $Y2=3.33
r118 44 45 1.43077 $w=1.7e-07 $l=1.105e-06 $layer=mcon $count=6 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r119 42 55 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r120 41 44 375.786 $w=1.68e-07 $l=5.76e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=6.96 $Y2=3.33
r121 41 42 1.43077 $w=1.7e-07 $l=1.105e-06 $layer=mcon $count=6 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r122 39 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.855 $Y=3.33
+ $X2=0.69 $Y2=3.33
r123 39 41 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.855 $Y=3.33
+ $X2=1.2 $Y2=3.33
r124 37 55 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r125 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r126 34 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.525 $Y=3.33
+ $X2=0.69 $Y2=3.33
r127 34 36 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.525 $Y=3.33
+ $X2=0.24 $Y2=3.33
r128 32 45 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=6.96 $Y2=3.33
r129 32 42 0.936549 $w=4.9e-07 $l=3.36e-06 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=1.2 $Y2=3.33
r130 30 47 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=8.015 $Y=3.33
+ $X2=7.92 $Y2=3.33
r131 30 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.015 $Y=3.33
+ $X2=8.18 $Y2=3.33
r132 29 50 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=8.345 $Y=3.33
+ $X2=8.88 $Y2=3.33
r133 29 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.345 $Y=3.33
+ $X2=8.18 $Y2=3.33
r134 27 44 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=7.155 $Y=3.33
+ $X2=6.96 $Y2=3.33
r135 27 28 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.155 $Y=3.33
+ $X2=7.32 $Y2=3.33
r136 26 47 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=7.485 $Y=3.33
+ $X2=7.92 $Y2=3.33
r137 26 28 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.485 $Y=3.33
+ $X2=7.32 $Y2=3.33
r138 22 25 26.5411 $w=3.28e-07 $l=7.6e-07 $layer=LI1_cond $X=8.18 $Y=2.19
+ $X2=8.18 $Y2=2.95
r139 20 31 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.18 $Y=3.245
+ $X2=8.18 $Y2=3.33
r140 20 25 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=8.18 $Y=3.245
+ $X2=8.18 $Y2=2.95
r141 16 19 26.5411 $w=3.28e-07 $l=7.6e-07 $layer=LI1_cond $X=7.32 $Y=2.19
+ $X2=7.32 $Y2=2.95
r142 14 28 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.32 $Y=3.245
+ $X2=7.32 $Y2=3.33
r143 14 19 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=7.32 $Y=3.245
+ $X2=7.32 $Y2=2.95
r144 10 54 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=3.245
+ $X2=0.69 $Y2=3.33
r145 10 12 29.5095 $w=3.28e-07 $l=8.45e-07 $layer=LI1_cond $X=0.69 $Y=3.245
+ $X2=0.69 $Y2=2.4
r146 3 25 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=8.04
+ $Y=1.835 $X2=8.18 $Y2=2.95
r147 3 22 400 $w=1.7e-07 $l=4.19196e-07 $layer=licon1_PDIFF $count=1 $X=8.04
+ $Y=1.835 $X2=8.18 $Y2=2.19
r148 2 19 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=7.18
+ $Y=1.835 $X2=7.32 $Y2=2.95
r149 2 16 400 $w=1.7e-07 $l=4.19196e-07 $layer=licon1_PDIFF $count=1 $X=7.18
+ $Y=1.835 $X2=7.32 $Y2=2.19
r150 1 12 300 $w=1.7e-07 $l=6.3113e-07 $layer=licon1_PDIFF $count=2 $X=0.55
+ $Y=1.835 $X2=0.69 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4B_4%A_217_367# 1 2 3 4 5 16 18 20 24 26 30 32 36
+ 38 42 47 49 50
r60 40 42 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=4.65 $Y=2.905
+ $X2=4.65 $Y2=2.46
r61 39 50 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=3.895 $Y=2.99 $X2=3.795
+ $Y2=2.99
r62 38 40 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.485 $Y=2.99
+ $X2=4.65 $Y2=2.905
r63 38 39 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=4.485 $Y=2.99
+ $X2=3.895 $Y2=2.99
r64 34 50 0.764409 $w=2e-07 $l=8.5e-08 $layer=LI1_cond $X=3.795 $Y=2.905
+ $X2=3.795 $Y2=2.99
r65 34 36 21.35 $w=1.98e-07 $l=3.85e-07 $layer=LI1_cond $X=3.795 $Y=2.905
+ $X2=3.795 $Y2=2.52
r66 33 49 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=3.025 $Y=2.99
+ $X2=2.93 $Y2=2.99
r67 32 50 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=3.695 $Y=2.99 $X2=3.795
+ $Y2=2.99
r68 32 33 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.695 $Y=2.99
+ $X2=3.025 $Y2=2.99
r69 28 49 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=2.93 $Y=2.905
+ $X2=2.93 $Y2=2.99
r70 28 30 42.9043 $w=1.88e-07 $l=7.35e-07 $layer=LI1_cond $X=2.93 $Y=2.905
+ $X2=2.93 $Y2=2.17
r71 27 47 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.165 $Y=2.99
+ $X2=2.07 $Y2=2.99
r72 26 49 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.835 $Y=2.99
+ $X2=2.93 $Y2=2.99
r73 26 27 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.835 $Y=2.99
+ $X2=2.165 $Y2=2.99
r74 22 47 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=2.07 $Y=2.905
+ $X2=2.07 $Y2=2.99
r75 22 24 42.9043 $w=1.88e-07 $l=7.35e-07 $layer=LI1_cond $X=2.07 $Y=2.905
+ $X2=2.07 $Y2=2.17
r76 21 45 3.82155 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.305 $Y=2.99
+ $X2=1.2 $Y2=2.99
r77 20 47 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.975 $Y=2.99
+ $X2=2.07 $Y2=2.99
r78 20 21 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.975 $Y=2.99
+ $X2=1.305 $Y2=2.99
r79 16 45 3.09364 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=1.2 $Y=2.905 $X2=1.2
+ $Y2=2.99
r80 16 18 48.8528 $w=2.08e-07 $l=9.25e-07 $layer=LI1_cond $X=1.2 $Y=2.905
+ $X2=1.2 $Y2=1.98
r81 5 42 300 $w=1.7e-07 $l=6.91466e-07 $layer=licon1_PDIFF $count=2 $X=4.51
+ $Y=1.835 $X2=4.65 $Y2=2.46
r82 4 36 300 $w=1.7e-07 $l=7.51748e-07 $layer=licon1_PDIFF $count=2 $X=3.65
+ $Y=1.835 $X2=3.79 $Y2=2.52
r83 3 49 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=2.79
+ $Y=1.835 $X2=2.93 $Y2=2.91
r84 3 30 400 $w=1.7e-07 $l=3.98905e-07 $layer=licon1_PDIFF $count=1 $X=2.79
+ $Y=1.835 $X2=2.93 $Y2=2.17
r85 2 47 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=1.93
+ $Y=1.835 $X2=2.07 $Y2=2.91
r86 2 24 400 $w=1.7e-07 $l=3.98905e-07 $layer=licon1_PDIFF $count=1 $X=1.93
+ $Y=1.835 $X2=2.07 $Y2=2.17
r87 1 45 400 $w=1.7e-07 $l=1.13578e-06 $layer=licon1_PDIFF $count=1 $X=1.085
+ $Y=1.835 $X2=1.21 $Y2=2.91
r88 1 18 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=1.085
+ $Y=1.835 $X2=1.21 $Y2=1.98
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4B_4%Y 1 2 3 4 5 6 7 8 9 10 33 35 36 39 43 44 47
+ 49 53 57 61 64 65 69 71 75 77 81 83 84 87 88 89 93 94 95 96 105 107 111 116
+ 121
c172 71 0 8.13651e-20 $X=7.145 $Y=1.095
c173 57 0 2.17431e-19 $X=4.87 $Y=1.75
r174 96 111 3.91717 $w=2.62e-07 $l=9.5e-08 $layer=LI1_cond $X=5.52 $Y=1.012
+ $X2=5.425 $Y2=1.012
r175 96 121 16.0017 $w=3.58e-07 $l=4.2e-07 $layer=LI1_cond $X=5.52 $Y=0.84
+ $X2=5.52 $Y2=0.42
r176 95 107 3.79035 $w=2.72e-07 $l=1.25956e-07 $layer=LI1_cond $X=4.965 $Y=1.012
+ $X2=4.87 $Y2=0.94
r177 95 112 3.79035 $w=2.72e-07 $l=9.5e-08 $layer=LI1_cond $X=4.965 $Y=1.012
+ $X2=5.06 $Y2=1.012
r178 95 111 11.1236 $w=3.43e-07 $l=3.33e-07 $layer=LI1_cond $X=5.092 $Y=1.012
+ $X2=5.425 $Y2=1.012
r179 95 112 1.06893 $w=3.43e-07 $l=3.2e-08 $layer=LI1_cond $X=5.092 $Y=1.012
+ $X2=5.06 $Y2=1.012
r180 94 107 17.1909 $w=1.98e-07 $l=3.1e-07 $layer=LI1_cond $X=4.56 $Y=0.94
+ $X2=4.87 $Y2=0.94
r181 94 108 16.9136 $w=1.98e-07 $l=3.05e-07 $layer=LI1_cond $X=4.56 $Y=0.94
+ $X2=4.255 $Y2=0.94
r182 93 105 4.9491 $w=2e-07 $l=9.5e-08 $layer=LI1_cond $X=4.16 $Y=0.94 $X2=4.065
+ $Y2=0.94
r183 93 108 4.9491 $w=2e-07 $l=9.5e-08 $layer=LI1_cond $X=4.16 $Y=0.94 $X2=4.255
+ $Y2=0.94
r184 93 116 18.0604 $w=2.88e-07 $l=4.2e-07 $layer=LI1_cond $X=4.16 $Y=0.84
+ $X2=4.16 $Y2=0.42
r185 93 105 1.94091 $w=1.98e-07 $l=3.5e-08 $layer=LI1_cond $X=4.03 $Y=0.94
+ $X2=4.065 $Y2=0.94
r186 89 91 5.76222 $w=2.78e-07 $l=1.4e-07 $layer=LI1_cond $X=7.285 $Y=0.955
+ $X2=7.285 $Y2=1.095
r187 89 90 3.90007 $w=2.78e-07 $l=8.5e-08 $layer=LI1_cond $X=7.285 $Y=0.955
+ $X2=7.285 $Y2=0.87
r188 85 93 34.6591 $w=1.98e-07 $l=6.25e-07 $layer=LI1_cond $X=3.405 $Y=0.94
+ $X2=4.03 $Y2=0.94
r189 85 87 5.16603 $w=1.9e-07 $l=1.23288e-07 $layer=LI1_cond $X=3.405 $Y=0.94
+ $X2=3.305 $Y2=0.992
r190 79 81 26.2679 $w=1.88e-07 $l=4.5e-07 $layer=LI1_cond $X=8.14 $Y=0.87
+ $X2=8.14 $Y2=0.42
r191 78 89 3.65648 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=7.425 $Y=0.955
+ $X2=7.285 $Y2=0.955
r192 77 79 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=8.045 $Y=0.955
+ $X2=8.14 $Y2=0.87
r193 77 78 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=8.045 $Y=0.955
+ $X2=7.425 $Y2=0.955
r194 75 90 22.5478 $w=2.28e-07 $l=4.5e-07 $layer=LI1_cond $X=7.26 $Y=0.42
+ $X2=7.26 $Y2=0.87
r195 72 88 5.40251 $w=1.8e-07 $l=9.5e-08 $layer=LI1_cond $X=6.475 $Y=1.095
+ $X2=6.38 $Y2=1.095
r196 71 91 3.32261 $w=1.8e-07 $l=1.4e-07 $layer=LI1_cond $X=7.145 $Y=1.095
+ $X2=7.285 $Y2=1.095
r197 71 72 41.2828 $w=1.78e-07 $l=6.7e-07 $layer=LI1_cond $X=7.145 $Y=1.095
+ $X2=6.475 $Y2=1.095
r198 67 88 1.14861 $w=1.9e-07 $l=9e-08 $layer=LI1_cond $X=6.38 $Y=1.005 $X2=6.38
+ $Y2=1.095
r199 67 69 34.1483 $w=1.88e-07 $l=5.85e-07 $layer=LI1_cond $X=6.38 $Y=1.005
+ $X2=6.38 $Y2=0.42
r200 66 96 3.91717 $w=2.62e-07 $l=1.30038e-07 $layer=LI1_cond $X=5.615 $Y=1.095
+ $X2=5.52 $Y2=1.012
r201 65 88 5.40251 $w=1.8e-07 $l=9.5e-08 $layer=LI1_cond $X=6.285 $Y=1.095
+ $X2=6.38 $Y2=1.095
r202 65 66 41.2828 $w=1.78e-07 $l=6.7e-07 $layer=LI1_cond $X=6.285 $Y=1.095
+ $X2=5.615 $Y2=1.095
r203 63 95 2.66798 $w=1.9e-07 $l=1.73e-07 $layer=LI1_cond $X=4.965 $Y=1.185
+ $X2=4.965 $Y2=1.012
r204 63 64 28.0191 $w=1.88e-07 $l=4.8e-07 $layer=LI1_cond $X=4.965 $Y=1.185
+ $X2=4.965 $Y2=1.665
r205 59 87 1.34256 $w=1.9e-07 $l=1.5448e-07 $layer=LI1_cond $X=3.3 $Y=0.84
+ $X2=3.305 $Y2=0.992
r206 59 61 24.5167 $w=1.88e-07 $l=4.2e-07 $layer=LI1_cond $X=3.3 $Y=0.84 $X2=3.3
+ $Y2=0.42
r207 58 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.665 $Y=1.75
+ $X2=2.5 $Y2=1.75
r208 57 64 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=4.87 $Y=1.75
+ $X2=4.965 $Y2=1.665
r209 57 58 143.856 $w=1.68e-07 $l=2.205e-06 $layer=LI1_cond $X=4.87 $Y=1.75
+ $X2=2.665 $Y2=1.75
r210 53 55 24.0965 $w=3.28e-07 $l=6.9e-07 $layer=LI1_cond $X=2.5 $Y=1.96 $X2=2.5
+ $Y2=2.65
r211 51 84 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.5 $Y=1.835 $X2=2.5
+ $Y2=1.75
r212 51 53 4.36531 $w=3.28e-07 $l=1.25e-07 $layer=LI1_cond $X=2.5 $Y=1.835
+ $X2=2.5 $Y2=1.96
r213 50 83 6.08426 $w=1.8e-07 $l=1.1e-07 $layer=LI1_cond $X=2.185 $Y=1.055
+ $X2=2.075 $Y2=1.055
r214 49 87 5.16603 $w=1.9e-07 $l=1.27671e-07 $layer=LI1_cond $X=3.205 $Y=1.055
+ $X2=3.305 $Y2=0.992
r215 49 50 62.8485 $w=1.78e-07 $l=1.02e-06 $layer=LI1_cond $X=3.205 $Y=1.055
+ $X2=2.185 $Y2=1.055
r216 45 83 0.630948 $w=2.2e-07 $l=9e-08 $layer=LI1_cond $X=2.075 $Y=0.965
+ $X2=2.075 $Y2=1.055
r217 45 47 28.5492 $w=2.18e-07 $l=5.45e-07 $layer=LI1_cond $X=2.075 $Y=0.965
+ $X2=2.075 $Y2=0.42
r218 43 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.335 $Y=1.75
+ $X2=2.5 $Y2=1.75
r219 43 44 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=2.335 $Y=1.75
+ $X2=1.805 $Y2=1.75
r220 39 41 24.0965 $w=3.28e-07 $l=6.9e-07 $layer=LI1_cond $X=1.64 $Y=1.96
+ $X2=1.64 $Y2=2.65
r221 37 44 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.64 $Y=1.835
+ $X2=1.805 $Y2=1.75
r222 37 39 4.36531 $w=3.28e-07 $l=1.25e-07 $layer=LI1_cond $X=1.64 $Y=1.835
+ $X2=1.64 $Y2=1.96
r223 35 83 6.08426 $w=1.8e-07 $l=1.1e-07 $layer=LI1_cond $X=1.965 $Y=1.055
+ $X2=2.075 $Y2=1.055
r224 35 36 41.2828 $w=1.78e-07 $l=6.7e-07 $layer=LI1_cond $X=1.965 $Y=1.055
+ $X2=1.295 $Y2=1.055
r225 31 36 6.84108 $w=1.8e-07 $l=1.3784e-07 $layer=LI1_cond $X=1.195 $Y=0.965
+ $X2=1.295 $Y2=1.055
r226 31 33 30.2227 $w=1.98e-07 $l=5.45e-07 $layer=LI1_cond $X=1.195 $Y=0.965
+ $X2=1.195 $Y2=0.42
r227 10 55 400 $w=1.7e-07 $l=8.82227e-07 $layer=licon1_PDIFF $count=1 $X=2.36
+ $Y=1.835 $X2=2.5 $Y2=2.65
r228 10 53 400 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=2.36
+ $Y=1.835 $X2=2.5 $Y2=1.96
r229 9 41 400 $w=1.7e-07 $l=8.82227e-07 $layer=licon1_PDIFF $count=1 $X=1.5
+ $Y=1.835 $X2=1.64 $Y2=2.65
r230 9 39 400 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=1.5
+ $Y=1.835 $X2=1.64 $Y2=1.96
r231 8 81 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=8
+ $Y=0.235 $X2=8.14 $Y2=0.42
r232 7 75 91 $w=1.7e-07 $l=2.48948e-07 $layer=licon1_NDIFF $count=2 $X=7.11
+ $Y=0.235 $X2=7.26 $Y2=0.42
r233 6 69 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=6.24
+ $Y=0.235 $X2=6.38 $Y2=0.42
r234 5 121 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=5.38
+ $Y=0.235 $X2=5.52 $Y2=0.42
r235 4 116 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=4.02
+ $Y=0.235 $X2=4.16 $Y2=0.42
r236 3 87 182 $w=1.7e-07 $l=7.61791e-07 $layer=licon1_NDIFF $count=1 $X=3.16
+ $Y=0.235 $X2=3.3 $Y2=0.93
r237 3 61 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=3.16
+ $Y=0.235 $X2=3.3 $Y2=0.42
r238 2 47 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=1.95
+ $Y=0.235 $X2=2.09 $Y2=0.42
r239 1 33 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=1.04
+ $Y=0.235 $X2=1.18 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4B_4%A_644_367# 1 2 3 4 15 19 21 25 27 32 34 36
+ 38
r45 28 36 6.19399 $w=1.8e-07 $l=1.13e-07 $layer=LI1_cond $X=5.73 $Y=2.095
+ $X2=5.617 $Y2=2.095
r46 27 38 4.92601 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=6.295 $Y=2.095
+ $X2=6.46 $Y2=2.095
r47 27 28 34.8131 $w=1.78e-07 $l=5.65e-07 $layer=LI1_cond $X=6.295 $Y=2.095
+ $X2=5.73 $Y2=2.095
r48 23 36 0.552779 $w=2.25e-07 $l=9e-08 $layer=LI1_cond $X=5.617 $Y=2.185
+ $X2=5.617 $Y2=2.095
r49 23 25 19.7196 $w=2.23e-07 $l=3.85e-07 $layer=LI1_cond $X=5.617 $Y=2.185
+ $X2=5.617 $Y2=2.57
r50 22 34 5.63431 $w=1.8e-07 $l=1e-07 $layer=LI1_cond $X=4.315 $Y=2.095
+ $X2=4.215 $Y2=2.095
r51 21 36 6.19399 $w=1.8e-07 $l=1.12e-07 $layer=LI1_cond $X=5.505 $Y=2.095
+ $X2=5.617 $Y2=2.095
r52 21 22 73.3232 $w=1.78e-07 $l=1.19e-06 $layer=LI1_cond $X=5.505 $Y=2.095
+ $X2=4.315 $Y2=2.095
r53 17 34 0.966048 $w=2e-07 $l=9e-08 $layer=LI1_cond $X=4.215 $Y=2.185 $X2=4.215
+ $Y2=2.095
r54 17 19 21.35 $w=1.98e-07 $l=3.85e-07 $layer=LI1_cond $X=4.215 $Y=2.185
+ $X2=4.215 $Y2=2.57
r55 16 32 4.92601 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=3.525 $Y=2.095
+ $X2=3.36 $Y2=2.095
r56 15 34 5.63431 $w=1.8e-07 $l=1e-07 $layer=LI1_cond $X=4.115 $Y=2.095
+ $X2=4.215 $Y2=2.095
r57 15 16 36.3535 $w=1.78e-07 $l=5.9e-07 $layer=LI1_cond $X=4.115 $Y=2.095
+ $X2=3.525 $Y2=2.095
r58 4 38 300 $w=1.7e-07 $l=3.27605e-07 $layer=licon1_PDIFF $count=2 $X=6.32
+ $Y=1.835 $X2=6.46 $Y2=2.1
r59 3 36 600 $w=1.7e-07 $l=3.27605e-07 $layer=licon1_PDIFF $count=1 $X=5.46
+ $Y=1.835 $X2=5.6 $Y2=2.1
r60 3 25 600 $w=1.7e-07 $l=8.01951e-07 $layer=licon1_PDIFF $count=1 $X=5.46
+ $Y=1.835 $X2=5.6 $Y2=2.57
r61 2 34 600 $w=1.7e-07 $l=3.27605e-07 $layer=licon1_PDIFF $count=1 $X=4.08
+ $Y=1.835 $X2=4.22 $Y2=2.1
r62 2 19 600 $w=1.7e-07 $l=8.01951e-07 $layer=licon1_PDIFF $count=1 $X=4.08
+ $Y=1.835 $X2=4.22 $Y2=2.57
r63 1 32 300 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=2 $X=3.22
+ $Y=1.835 $X2=3.36 $Y2=2.11
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4B_4%A_1009_367# 1 2 3 4 5 18 20 21 24 26 29 32
+ 33 36 40 44 48 51
c65 1 0 1.66402e-19 $X=5.045 $Y=1.835
r66 44 46 41.222 $w=2.58e-07 $l=9.3e-07 $layer=LI1_cond $X=8.645 $Y=1.98
+ $X2=8.645 $Y2=2.91
r67 42 44 2.43786 $w=2.58e-07 $l=5.5e-08 $layer=LI1_cond $X=8.645 $Y=1.925
+ $X2=8.645 $Y2=1.98
r68 41 51 4.39427 $w=2.3e-07 $l=9.5e-08 $layer=LI1_cond $X=7.845 $Y=1.81
+ $X2=7.75 $Y2=1.81
r69 40 42 6.84978 $w=2.3e-07 $l=1.78466e-07 $layer=LI1_cond $X=8.515 $Y=1.81
+ $X2=8.645 $Y2=1.925
r70 40 41 33.5712 $w=2.28e-07 $l=6.7e-07 $layer=LI1_cond $X=8.515 $Y=1.81
+ $X2=7.845 $Y2=1.81
r71 36 38 54.2871 $w=1.88e-07 $l=9.3e-07 $layer=LI1_cond $X=7.75 $Y=1.98
+ $X2=7.75 $Y2=2.91
r72 34 51 2.03875 $w=1.9e-07 $l=1.15e-07 $layer=LI1_cond $X=7.75 $Y=1.925
+ $X2=7.75 $Y2=1.81
r73 34 36 3.21053 $w=1.88e-07 $l=5.5e-08 $layer=LI1_cond $X=7.75 $Y=1.925
+ $X2=7.75 $Y2=1.98
r74 32 51 4.39427 $w=2.3e-07 $l=9.5e-08 $layer=LI1_cond $X=7.655 $Y=1.81
+ $X2=7.75 $Y2=1.81
r75 32 33 33.5712 $w=2.28e-07 $l=6.7e-07 $layer=LI1_cond $X=7.655 $Y=1.81
+ $X2=6.985 $Y2=1.81
r76 29 50 3.23184 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=6.89 $Y=2.905
+ $X2=6.89 $Y2=2.99
r77 29 31 53.9952 $w=1.88e-07 $l=9.25e-07 $layer=LI1_cond $X=6.89 $Y=2.905
+ $X2=6.89 $Y2=1.98
r78 28 33 6.89722 $w=2.3e-07 $l=1.55403e-07 $layer=LI1_cond $X=6.89 $Y=1.925
+ $X2=6.985 $Y2=1.81
r79 28 31 3.21053 $w=1.88e-07 $l=5.5e-08 $layer=LI1_cond $X=6.89 $Y=1.925
+ $X2=6.89 $Y2=1.98
r80 27 48 6.47928 $w=1.7e-07 $l=1.13e-07 $layer=LI1_cond $X=6.125 $Y=2.99
+ $X2=6.012 $Y2=2.99
r81 26 50 3.61205 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=6.795 $Y=2.99
+ $X2=6.89 $Y2=2.99
r82 26 27 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=6.795 $Y=2.99
+ $X2=6.125 $Y2=2.99
r83 22 48 0.355529 $w=2.25e-07 $l=8.5e-08 $layer=LI1_cond $X=6.012 $Y=2.905
+ $X2=6.012 $Y2=2.99
r84 22 24 19.7196 $w=2.23e-07 $l=3.85e-07 $layer=LI1_cond $X=6.012 $Y=2.905
+ $X2=6.012 $Y2=2.52
r85 20 48 6.47928 $w=1.7e-07 $l=1.12e-07 $layer=LI1_cond $X=5.9 $Y=2.99
+ $X2=6.012 $Y2=2.99
r86 20 21 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=5.9 $Y=2.99
+ $X2=5.335 $Y2=2.99
r87 16 21 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.17 $Y=2.905
+ $X2=5.335 $Y2=2.99
r88 16 18 15.1913 $w=3.28e-07 $l=4.35e-07 $layer=LI1_cond $X=5.17 $Y=2.905
+ $X2=5.17 $Y2=2.47
r89 5 46 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=8.47
+ $Y=1.835 $X2=8.61 $Y2=2.91
r90 5 44 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=8.47
+ $Y=1.835 $X2=8.61 $Y2=1.98
r91 4 38 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=7.61
+ $Y=1.835 $X2=7.75 $Y2=2.91
r92 4 36 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=7.61
+ $Y=1.835 $X2=7.75 $Y2=1.98
r93 3 50 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=6.75
+ $Y=1.835 $X2=6.89 $Y2=2.91
r94 3 31 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=6.75
+ $Y=1.835 $X2=6.89 $Y2=1.98
r95 2 24 300 $w=1.7e-07 $l=7.51748e-07 $layer=licon1_PDIFF $count=2 $X=5.89
+ $Y=1.835 $X2=6.03 $Y2=2.52
r96 1 18 300 $w=1.7e-07 $l=6.94694e-07 $layer=licon1_PDIFF $count=2 $X=5.045
+ $Y=1.835 $X2=5.17 $Y2=2.47
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4B_4%VGND 1 2 3 4 5 6 7 8 9 30 34 38 40 44 48 52
+ 56 60 63 64 66 67 69 70 71 73 78 83 93 109 110 113 116 119 122 127 133 135
r148 135 136 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6
+ $Y2=0
r149 132 133 11.1544 $w=7.53e-07 $l=1.65e-07 $layer=LI1_cond $X=5.09 $Y=0.292
+ $X2=5.255 $Y2=0.292
r150 129 132 0.792105 $w=7.53e-07 $l=5e-08 $layer=LI1_cond $X=5.04 $Y=0.292
+ $X2=5.09 $Y2=0.292
r151 129 130 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0
+ $X2=5.04 $Y2=0
r152 125 129 7.60421 $w=7.53e-07 $l=4.8e-07 $layer=LI1_cond $X=4.56 $Y=0.292
+ $X2=5.04 $Y2=0.292
r153 125 127 10.6792 $w=7.53e-07 $l=1.35e-07 $layer=LI1_cond $X=4.56 $Y=0.292
+ $X2=4.425 $Y2=0.292
r154 122 123 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r155 120 123 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0
+ $X2=3.6 $Y2=0
r156 119 120 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0
+ $X2=2.64 $Y2=0
r157 116 117 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0
+ $X2=1.68 $Y2=0
r158 113 114 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0
+ $X2=0.72 $Y2=0
r159 109 110 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=0
+ $X2=8.88 $Y2=0
r160 107 110 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=0
+ $X2=8.88 $Y2=0
r161 106 107 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r162 104 107 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.44 $Y=0
+ $X2=8.4 $Y2=0
r163 103 104 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=0
+ $X2=7.44 $Y2=0
r164 101 104 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.48 $Y=0
+ $X2=7.44 $Y2=0
r165 101 136 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6
+ $Y2=0
r166 100 101 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=0
+ $X2=6.48 $Y2=0
r167 98 135 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.115 $Y=0
+ $X2=5.95 $Y2=0
r168 98 100 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=6.115 $Y=0
+ $X2=6.48 $Y2=0
r169 97 136 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=6
+ $Y2=0
r170 97 130 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0
+ $X2=5.04 $Y2=0
r171 96 133 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=5.52 $Y=0
+ $X2=5.255 $Y2=0
r172 96 97 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r173 93 135 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.785 $Y=0
+ $X2=5.95 $Y2=0
r174 93 96 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=5.785 $Y=0
+ $X2=5.52 $Y2=0
r175 92 123 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.6
+ $Y2=0
r176 91 127 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=4.08 $Y=0
+ $X2=4.425 $Y2=0
r177 91 92 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r178 89 122 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.895 $Y=0
+ $X2=3.73 $Y2=0
r179 89 91 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=3.895 $Y=0
+ $X2=4.08 $Y2=0
r180 87 120 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0
+ $X2=2.64 $Y2=0
r181 87 117 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0
+ $X2=1.68 $Y2=0
r182 86 87 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r183 84 116 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.795 $Y=0
+ $X2=1.63 $Y2=0
r184 84 86 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=1.795 $Y=0
+ $X2=2.16 $Y2=0
r185 83 119 13.4521 $w=1.7e-07 $l=3.4e-07 $layer=LI1_cond $X=2.355 $Y=0
+ $X2=2.695 $Y2=0
r186 83 86 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=2.355 $Y=0
+ $X2=2.16 $Y2=0
r187 82 117 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r188 82 114 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r189 81 82 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r190 79 113 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.865 $Y=0 $X2=0.7
+ $Y2=0
r191 79 81 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=0.865 $Y=0 $X2=1.2
+ $Y2=0
r192 78 116 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.465 $Y=0
+ $X2=1.63 $Y2=0
r193 78 81 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=1.465 $Y=0 $X2=1.2
+ $Y2=0
r194 76 114 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0
+ $X2=0.72 $Y2=0
r195 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r196 73 113 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.535 $Y=0 $X2=0.7
+ $Y2=0
r197 73 75 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.535 $Y=0 $X2=0.24
+ $Y2=0
r198 71 130 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0
+ $X2=5.04 $Y2=0
r199 71 92 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=4.08
+ $Y2=0
r200 71 125 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r201 69 106 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=8.405 $Y=0 $X2=8.4
+ $Y2=0
r202 69 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.405 $Y=0 $X2=8.57
+ $Y2=0
r203 68 109 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=8.735 $Y=0
+ $X2=8.88 $Y2=0
r204 68 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.735 $Y=0 $X2=8.57
+ $Y2=0
r205 66 103 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=7.545 $Y=0
+ $X2=7.44 $Y2=0
r206 66 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.545 $Y=0 $X2=7.71
+ $Y2=0
r207 65 106 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=7.875 $Y=0
+ $X2=8.4 $Y2=0
r208 65 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.875 $Y=0 $X2=7.71
+ $Y2=0
r209 63 100 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=6.645 $Y=0
+ $X2=6.48 $Y2=0
r210 63 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.645 $Y=0 $X2=6.81
+ $Y2=0
r211 62 103 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=6.975 $Y=0
+ $X2=7.44 $Y2=0
r212 62 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.975 $Y=0 $X2=6.81
+ $Y2=0
r213 58 70 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.57 $Y=0.085
+ $X2=8.57 $Y2=0
r214 58 60 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=8.57 $Y=0.085
+ $X2=8.57 $Y2=0.38
r215 54 67 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.71 $Y=0.085
+ $X2=7.71 $Y2=0
r216 54 56 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=7.71 $Y=0.085
+ $X2=7.71 $Y2=0.535
r217 50 64 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.81 $Y=0.085
+ $X2=6.81 $Y2=0
r218 50 52 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=6.81 $Y=0.085
+ $X2=6.81 $Y2=0.38
r219 46 135 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.95 $Y=0.085
+ $X2=5.95 $Y2=0
r220 46 48 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=5.95 $Y=0.085
+ $X2=5.95 $Y2=0.38
r221 42 122 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.73 $Y=0.085
+ $X2=3.73 $Y2=0
r222 42 44 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=3.73 $Y=0.085
+ $X2=3.73 $Y2=0.55
r223 41 119 13.4521 $w=1.7e-07 $l=3.4e-07 $layer=LI1_cond $X=3.035 $Y=0
+ $X2=2.695 $Y2=0
r224 40 122 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.565 $Y=0
+ $X2=3.73 $Y2=0
r225 40 41 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=3.565 $Y=0
+ $X2=3.035 $Y2=0
r226 36 119 2.80049 $w=6.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.695 $Y=0.085
+ $X2=2.695 $Y2=0
r227 36 38 4.83708 $w=6.78e-07 $l=2.75e-07 $layer=LI1_cond $X=2.695 $Y=0.085
+ $X2=2.695 $Y2=0.36
r228 32 116 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.63 $Y=0.085
+ $X2=1.63 $Y2=0
r229 32 34 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=1.63 $Y=0.085
+ $X2=1.63 $Y2=0.36
r230 28 113 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.7 $Y=0.085
+ $X2=0.7 $Y2=0
r231 28 30 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=0.7 $Y=0.085
+ $X2=0.7 $Y2=0.36
r232 9 60 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=8.43
+ $Y=0.235 $X2=8.57 $Y2=0.38
r233 8 56 182 $w=1.7e-07 $l=3.63318e-07 $layer=licon1_NDIFF $count=1 $X=7.57
+ $Y=0.235 $X2=7.71 $Y2=0.535
r234 7 52 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.67
+ $Y=0.235 $X2=6.81 $Y2=0.38
r235 6 48 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.81
+ $Y=0.235 $X2=5.95 $Y2=0.38
r236 5 132 91 $w=1.7e-07 $l=7.73563e-07 $layer=licon1_NDIFF $count=2 $X=4.45
+ $Y=0.235 $X2=5.09 $Y2=0.53
r237 4 44 182 $w=1.7e-07 $l=3.78583e-07 $layer=licon1_NDIFF $count=1 $X=3.59
+ $Y=0.235 $X2=3.73 $Y2=0.55
r238 3 38 45.5 $w=1.7e-07 $l=5.48954e-07 $layer=licon1_NDIFF $count=4 $X=2.38
+ $Y=0.235 $X2=2.87 $Y2=0.36
r239 2 34 91 $w=1.7e-07 $l=2.13542e-07 $layer=licon1_NDIFF $count=2 $X=1.47
+ $Y=0.235 $X2=1.63 $Y2=0.36
r240 1 30 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=0.56
+ $Y=0.235 $X2=0.7 $Y2=0.36
.ends

