* NGSPICE file created from sky130_fd_sc_lp__diode_1.ext - technology: sky130A

.subckt sky130_fd_sc_lp__diode_1 DIODE VGND VNB VPB VPWR
.ends

