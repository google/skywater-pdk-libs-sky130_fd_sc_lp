* File: sky130_fd_sc_lp__mux2_4.pex.spice
* Created: Wed Sep  2 10:00:19 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__MUX2_4%S 1 3 5 7 8 10 13 17 20 21 22 23 30 33 39
c94 21 0 1.31789e-19 $X=0.69 $Y=1.78
c95 13 0 3.37017e-20 $X=3.305 $Y=2.465
r96 33 39 0.987808 $w=3.48e-07 $l=3e-08 $layer=LI1_cond $X=3.08 $Y=1.695
+ $X2=3.08 $Y2=1.665
r97 28 30 41.0035 $w=2.88e-07 $l=2.45e-07 $layer=POLY_cond $X=2.825 $Y=1.35
+ $X2=3.07 $Y2=1.35
r98 23 33 2.59474 $w=3.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.08 $Y=1.78 $X2=3.08
+ $Y2=1.695
r99 23 39 0.921954 $w=3.48e-07 $l=2.8e-08 $layer=LI1_cond $X=3.08 $Y=1.637
+ $X2=3.08 $Y2=1.665
r100 22 23 11.261 $w=3.48e-07 $l=3.42e-07 $layer=LI1_cond $X=3.08 $Y=1.295
+ $X2=3.08 $Y2=1.637
r101 22 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.07
+ $Y=1.35 $X2=3.07 $Y2=1.35
r102 20 23 5.34211 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=2.905 $Y=1.78
+ $X2=3.08 $Y2=1.78
r103 20 21 144.508 $w=1.68e-07 $l=2.215e-06 $layer=LI1_cond $X=2.905 $Y=1.78
+ $X2=0.69 $Y2=1.78
r104 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.525
+ $Y=1.5 $X2=0.525 $Y2=1.5
r105 15 21 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=0.56 $Y=1.695
+ $X2=0.69 $Y2=1.78
r106 15 17 8.64332 $w=2.58e-07 $l=1.95e-07 $layer=LI1_cond $X=0.56 $Y=1.695
+ $X2=0.56 $Y2=1.5
r107 11 30 39.3299 $w=2.88e-07 $l=3.06594e-07 $layer=POLY_cond $X=3.305 $Y=1.515
+ $X2=3.07 $Y2=1.35
r108 11 13 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=3.305 $Y=1.515
+ $X2=3.305 $Y2=2.465
r109 8 28 18.0107 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.825 $Y=1.185
+ $X2=2.825 $Y2=1.35
r110 8 10 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.825 $Y=1.185
+ $X2=2.825 $Y2=0.655
r111 5 18 58.0228 $w=3.87e-07 $l=3.96068e-07 $layer=POLY_cond $X=0.8 $Y=1.185
+ $X2=0.617 $Y2=1.5
r112 5 7 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.8 $Y=1.185 $X2=0.8
+ $Y2=0.655
r113 1 18 39.3407 $w=3.87e-07 $l=1.9775e-07 $layer=POLY_cond $X=0.545 $Y=1.665
+ $X2=0.617 $Y2=1.5
r114 1 3 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=0.545 $Y=1.665
+ $X2=0.545 $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__MUX2_4%A_41_367# 1 2 7 9 12 16 22 24 28 29 31 33 34
c56 28 0 7.98639e-21 $X=1.25 $Y=1.43
c57 24 0 1.82641e-19 $X=1.085 $Y=1.07
r58 33 34 8.46614 $w=3.33e-07 $l=1.65e-07 $layer=LI1_cond $X=0.257 $Y=2.2
+ $X2=0.257 $Y2=2.035
r59 29 37 15.0625 $w=3.52e-07 $l=1.1e-07 $layer=POLY_cond $X=1.25 $Y=1.495
+ $X2=1.36 $Y2=1.495
r60 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.25
+ $Y=1.43 $X2=1.25 $Y2=1.43
r61 26 28 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=1.25 $Y=1.155
+ $X2=1.25 $Y2=1.43
r62 25 31 4.4465 $w=1.7e-07 $l=3.05e-07 $layer=LI1_cond $X=0.7 $Y=1.07 $X2=0.395
+ $Y2=1.07
r63 24 26 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.085 $Y=1.07
+ $X2=1.25 $Y2=1.155
r64 24 25 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=1.085 $Y=1.07
+ $X2=0.7 $Y2=1.07
r65 20 33 0.0688026 $w=3.33e-07 $l=2e-09 $layer=LI1_cond $X=0.257 $Y=2.202
+ $X2=0.257 $Y2=2.2
r66 20 22 24.3561 $w=3.33e-07 $l=7.08e-07 $layer=LI1_cond $X=0.257 $Y=2.202
+ $X2=0.257 $Y2=2.91
r67 18 31 2.47594 $w=3.9e-07 $l=2.59037e-07 $layer=LI1_cond $X=0.175 $Y=1.155
+ $X2=0.395 $Y2=1.07
r68 18 34 57.4118 $w=1.68e-07 $l=8.8e-07 $layer=LI1_cond $X=0.175 $Y=1.155
+ $X2=0.175 $Y2=2.035
r69 14 31 2.47594 $w=3.9e-07 $l=8.5e-08 $layer=LI1_cond $X=0.395 $Y=0.985
+ $X2=0.395 $Y2=1.07
r70 14 16 11.0784 $w=6.08e-07 $l=5.65e-07 $layer=LI1_cond $X=0.395 $Y=0.985
+ $X2=0.395 $Y2=0.42
r71 10 37 22.7654 $w=1.5e-07 $l=2.3e-07 $layer=POLY_cond $X=1.36 $Y=1.265
+ $X2=1.36 $Y2=1.495
r72 10 12 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.36 $Y=1.265
+ $X2=1.36 $Y2=0.655
r73 7 29 37.6562 $w=3.52e-07 $l=3.72659e-07 $layer=POLY_cond $X=0.975 $Y=1.725
+ $X2=1.25 $Y2=1.495
r74 7 9 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=0.975 $Y=1.725
+ $X2=0.975 $Y2=2.465
r75 2 33 400 $w=1.7e-07 $l=4.22907e-07 $layer=licon1_PDIFF $count=1 $X=0.205
+ $Y=1.835 $X2=0.33 $Y2=2.2
r76 2 22 400 $w=1.7e-07 $l=1.13578e-06 $layer=licon1_PDIFF $count=1 $X=0.205
+ $Y=1.835 $X2=0.33 $Y2=2.91
r77 1 16 91 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=2 $X=0.46
+ $Y=0.235 $X2=0.585 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__MUX2_4%A0 1 3 6 8 9 10 19
c41 8 0 6.38927e-21 $X=1.68 $Y=0.555
c42 6 0 7.98639e-21 $X=1.925 $Y=2.465
c43 1 0 1.82641e-19 $X=1.72 $Y=1.185
r44 17 19 20.109 $w=3.3e-07 $l=1.15e-07 $layer=POLY_cond $X=1.81 $Y=1.35
+ $X2=1.925 $Y2=1.35
r45 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.81
+ $Y=1.35 $X2=1.81 $Y2=1.35
r46 14 17 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=1.72 $Y=1.35 $X2=1.81
+ $Y2=1.35
r47 10 18 1.98076 $w=3.18e-07 $l=5.5e-08 $layer=LI1_cond $X=1.745 $Y=1.295
+ $X2=1.745 $Y2=1.35
r48 9 10 13.3251 $w=3.18e-07 $l=3.7e-07 $layer=LI1_cond $X=1.745 $Y=0.925
+ $X2=1.745 $Y2=1.295
r49 8 9 13.3251 $w=3.18e-07 $l=3.7e-07 $layer=LI1_cond $X=1.745 $Y=0.555
+ $X2=1.745 $Y2=0.925
r50 4 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.925 $Y=1.515
+ $X2=1.925 $Y2=1.35
r51 4 6 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=1.925 $Y=1.515
+ $X2=1.925 $Y2=2.465
r52 1 14 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.72 $Y=1.185
+ $X2=1.72 $Y2=1.35
r53 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.72 $Y=1.185 $X2=1.72
+ $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__MUX2_4%A1 3 7 8 9 13 15
c38 9 0 3.37017e-20 $X=2.64 $Y=1.295
c39 3 0 6.38927e-21 $X=2.355 $Y=2.465
r40 13 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.375 $Y=1.35
+ $X2=2.375 $Y2=1.515
r41 13 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.375 $Y=1.35
+ $X2=2.375 $Y2=1.185
r42 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.375
+ $Y=1.35 $X2=2.375 $Y2=1.35
r43 9 14 9.39684 $w=3.23e-07 $l=2.65e-07 $layer=LI1_cond $X=2.64 $Y=1.362
+ $X2=2.375 $Y2=1.362
r44 8 14 7.62385 $w=3.23e-07 $l=2.15e-07 $layer=LI1_cond $X=2.16 $Y=1.362
+ $X2=2.375 $Y2=1.362
r45 7 15 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.465 $Y=0.655
+ $X2=2.465 $Y2=1.185
r46 3 16 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=2.355 $Y=2.465
+ $X2=2.355 $Y2=1.515
.ends

.subckt PM_SKY130_FD_SC_LP__MUX2_4%A_359_47# 1 2 9 13 17 21 25 29 33 37 41 43 45
+ 46 48 50 56 57 62 63
r136 72 73 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=4.955 $Y=1.5
+ $X2=5.025 $Y2=1.5
r137 71 72 62.9501 $w=3.3e-07 $l=3.6e-07 $layer=POLY_cond $X=4.595 $Y=1.5
+ $X2=4.955 $Y2=1.5
r138 70 71 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=4.525 $Y=1.5
+ $X2=4.595 $Y2=1.5
r139 69 70 62.9501 $w=3.3e-07 $l=3.6e-07 $layer=POLY_cond $X=4.165 $Y=1.5
+ $X2=4.525 $Y2=1.5
r140 68 69 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=4.095 $Y=1.5
+ $X2=4.165 $Y2=1.5
r141 64 66 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=3.665 $Y=1.5
+ $X2=3.735 $Y2=1.5
r142 60 62 8.16804 $w=2.98e-07 $l=1.65e-07 $layer=LI1_cond $X=2.14 $Y=2.185
+ $X2=2.305 $Y2=2.185
r143 57 73 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=5.115 $Y=1.5
+ $X2=5.025 $Y2=1.5
r144 56 57 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=5.115
+ $Y=1.5 $X2=5.115 $Y2=1.5
r145 54 68 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=3.755 $Y=1.5
+ $X2=4.095 $Y2=1.5
r146 54 66 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=3.755 $Y=1.5
+ $X2=3.735 $Y2=1.5
r147 53 56 83.798 $w=1.78e-07 $l=1.36e-06 $layer=LI1_cond $X=3.755 $Y=1.495
+ $X2=5.115 $Y2=1.495
r148 53 54 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=3.755
+ $Y=1.5 $X2=3.755 $Y2=1.5
r149 51 63 1.6787 $w=1.8e-07 $l=1.13e-07 $layer=LI1_cond $X=3.65 $Y=1.495
+ $X2=3.537 $Y2=1.495
r150 51 53 6.4697 $w=1.78e-07 $l=1.05e-07 $layer=LI1_cond $X=3.65 $Y=1.495
+ $X2=3.755 $Y2=1.495
r151 49 63 4.77889 $w=1.97e-07 $l=9e-08 $layer=LI1_cond $X=3.537 $Y=1.585
+ $X2=3.537 $Y2=1.495
r152 49 50 23.0489 $w=2.23e-07 $l=4.5e-07 $layer=LI1_cond $X=3.537 $Y=1.585
+ $X2=3.537 $Y2=2.035
r153 48 63 4.77889 $w=1.97e-07 $l=1.02616e-07 $layer=LI1_cond $X=3.51 $Y=1.405
+ $X2=3.537 $Y2=1.495
r154 47 48 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=3.51 $Y=1.03
+ $X2=3.51 $Y2=1.405
r155 45 47 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.425 $Y=0.945
+ $X2=3.51 $Y2=1.03
r156 45 46 58.3904 $w=1.68e-07 $l=8.95e-07 $layer=LI1_cond $X=3.425 $Y=0.945
+ $X2=2.53 $Y2=0.945
r157 43 50 6.92652 $w=1.8e-07 $l=1.50413e-07 $layer=LI1_cond $X=3.425 $Y=2.125
+ $X2=3.537 $Y2=2.035
r158 43 62 69.0101 $w=1.78e-07 $l=1.12e-06 $layer=LI1_cond $X=3.425 $Y=2.125
+ $X2=2.305 $Y2=2.125
r159 39 46 8.76165 $w=1.7e-07 $l=2.62076e-07 $layer=LI1_cond $X=2.307 $Y=0.86
+ $X2=2.53 $Y2=0.945
r160 39 41 12.9488 $w=4.43e-07 $l=5e-07 $layer=LI1_cond $X=2.307 $Y=0.86
+ $X2=2.307 $Y2=0.36
r161 35 73 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.025 $Y=1.665
+ $X2=5.025 $Y2=1.5
r162 35 37 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=5.025 $Y=1.665
+ $X2=5.025 $Y2=2.465
r163 31 72 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.955 $Y=1.335
+ $X2=4.955 $Y2=1.5
r164 31 33 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=4.955 $Y=1.335
+ $X2=4.955 $Y2=0.655
r165 27 71 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.595 $Y=1.665
+ $X2=4.595 $Y2=1.5
r166 27 29 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=4.595 $Y=1.665
+ $X2=4.595 $Y2=2.465
r167 23 70 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.525 $Y=1.335
+ $X2=4.525 $Y2=1.5
r168 23 25 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=4.525 $Y=1.335
+ $X2=4.525 $Y2=0.655
r169 19 69 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.165 $Y=1.665
+ $X2=4.165 $Y2=1.5
r170 19 21 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=4.165 $Y=1.665
+ $X2=4.165 $Y2=2.465
r171 15 68 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.095 $Y=1.335
+ $X2=4.095 $Y2=1.5
r172 15 17 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=4.095 $Y=1.335
+ $X2=4.095 $Y2=0.655
r173 11 66 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.735 $Y=1.665
+ $X2=3.735 $Y2=1.5
r174 11 13 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=3.735 $Y=1.665
+ $X2=3.735 $Y2=2.465
r175 7 64 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.665 $Y=1.335
+ $X2=3.665 $Y2=1.5
r176 7 9 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=3.665 $Y=1.335
+ $X2=3.665 $Y2=0.655
r177 2 60 600 $w=1.7e-07 $l=3.98905e-07 $layer=licon1_PDIFF $count=1 $X=2
+ $Y=1.835 $X2=2.14 $Y2=2.17
r178 1 41 91 $w=1.7e-07 $l=5.13712e-07 $layer=licon1_NDIFF $count=2 $X=1.795
+ $Y=0.235 $X2=2.25 $Y2=0.36
.ends

.subckt PM_SKY130_FD_SC_LP__MUX2_4%VPWR 1 2 3 4 15 21 25 31 36 37 39 40 41 43 48
+ 64 65 68 71
c77 1 0 1.31789e-19 $X=0.62 $Y=1.835
r78 71 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r79 68 69 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r80 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r81 62 65 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=5.52 $Y2=3.33
r82 61 62 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r83 59 62 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=5.04 $Y2=3.33
r84 59 72 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.6 $Y2=3.33
r85 58 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r86 56 71 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.685 $Y=3.33
+ $X2=3.52 $Y2=3.33
r87 56 58 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=3.685 $Y=3.33
+ $X2=4.08 $Y2=3.33
r88 55 72 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r89 54 55 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r90 52 69 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r91 51 54 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=3.12 $Y2=3.33
r92 51 52 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r93 49 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.925 $Y=3.33
+ $X2=0.76 $Y2=3.33
r94 49 51 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.925 $Y=3.33
+ $X2=1.2 $Y2=3.33
r95 48 71 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.355 $Y=3.33
+ $X2=3.52 $Y2=3.33
r96 48 54 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=3.355 $Y=3.33
+ $X2=3.12 $Y2=3.33
r97 46 69 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r98 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r99 43 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.595 $Y=3.33
+ $X2=0.76 $Y2=3.33
r100 43 45 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=0.595 $Y=3.33
+ $X2=0.24 $Y2=3.33
r101 41 55 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.88 $Y=3.33
+ $X2=3.12 $Y2=3.33
r102 41 52 0.468274 $w=4.9e-07 $l=1.68e-06 $layer=MET1_cond $X=2.88 $Y=3.33
+ $X2=1.2 $Y2=3.33
r103 39 61 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=5.075 $Y=3.33
+ $X2=5.04 $Y2=3.33
r104 39 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.075 $Y=3.33
+ $X2=5.24 $Y2=3.33
r105 38 64 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=5.405 $Y=3.33
+ $X2=5.52 $Y2=3.33
r106 38 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.405 $Y=3.33
+ $X2=5.24 $Y2=3.33
r107 36 58 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=4.215 $Y=3.33
+ $X2=4.08 $Y2=3.33
r108 36 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.215 $Y=3.33
+ $X2=4.38 $Y2=3.33
r109 35 61 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=4.545 $Y=3.33
+ $X2=5.04 $Y2=3.33
r110 35 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.545 $Y=3.33
+ $X2=4.38 $Y2=3.33
r111 31 34 26.8903 $w=3.28e-07 $l=7.7e-07 $layer=LI1_cond $X=5.24 $Y=2.18
+ $X2=5.24 $Y2=2.95
r112 29 40 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.24 $Y=3.245
+ $X2=5.24 $Y2=3.33
r113 29 34 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=5.24 $Y=3.245
+ $X2=5.24 $Y2=2.95
r114 25 28 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=4.38 $Y=2.18
+ $X2=4.38 $Y2=2.97
r115 23 37 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.38 $Y=3.245
+ $X2=4.38 $Y2=3.33
r116 23 28 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=4.38 $Y=3.245
+ $X2=4.38 $Y2=2.97
r117 19 71 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.52 $Y=3.245
+ $X2=3.52 $Y2=3.33
r118 19 21 24.9696 $w=3.28e-07 $l=7.15e-07 $layer=LI1_cond $X=3.52 $Y=3.245
+ $X2=3.52 $Y2=2.53
r119 15 18 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=0.76 $Y=2.12
+ $X2=0.76 $Y2=2.95
r120 13 68 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.76 $Y=3.245
+ $X2=0.76 $Y2=3.33
r121 13 18 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.76 $Y=3.245
+ $X2=0.76 $Y2=2.95
r122 4 34 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=5.1
+ $Y=1.835 $X2=5.24 $Y2=2.95
r123 4 31 400 $w=1.7e-07 $l=4.09054e-07 $layer=licon1_PDIFF $count=1 $X=5.1
+ $Y=1.835 $X2=5.24 $Y2=2.18
r124 3 28 400 $w=1.7e-07 $l=1.20297e-06 $layer=licon1_PDIFF $count=1 $X=4.24
+ $Y=1.835 $X2=4.38 $Y2=2.97
r125 3 25 400 $w=1.7e-07 $l=4.09054e-07 $layer=licon1_PDIFF $count=1 $X=4.24
+ $Y=1.835 $X2=4.38 $Y2=2.18
r126 2 21 300 $w=1.7e-07 $l=7.61791e-07 $layer=licon1_PDIFF $count=2 $X=3.38
+ $Y=1.835 $X2=3.52 $Y2=2.53
r127 1 18 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=0.62
+ $Y=1.835 $X2=0.76 $Y2=2.95
r128 1 15 400 $w=1.7e-07 $l=3.4803e-07 $layer=licon1_PDIFF $count=1 $X=0.62
+ $Y=1.835 $X2=0.76 $Y2=2.12
.ends

.subckt PM_SKY130_FD_SC_LP__MUX2_4%A_210_367# 1 2 9 14 16 17
r29 16 17 9.07524 $w=2.28e-07 $l=1.65e-07 $layer=LI1_cond $X=2.57 $Y=2.96
+ $X2=2.405 $Y2=2.96
r30 14 17 68.5027 $w=1.68e-07 $l=1.05e-06 $layer=LI1_cond $X=1.355 $Y=2.99
+ $X2=2.405 $Y2=2.99
r31 9 12 30.1408 $w=2.58e-07 $l=6.8e-07 $layer=LI1_cond $X=1.225 $Y=2.22
+ $X2=1.225 $Y2=2.9
r32 7 14 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=1.225 $Y=2.905
+ $X2=1.355 $Y2=2.99
r33 7 12 0.221624 $w=2.58e-07 $l=5e-09 $layer=LI1_cond $X=1.225 $Y=2.905
+ $X2=1.225 $Y2=2.9
r34 2 16 600 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=2.43
+ $Y=1.835 $X2=2.57 $Y2=2.95
r35 1 12 400 $w=1.7e-07 $l=1.13284e-06 $layer=licon1_PDIFF $count=1 $X=1.05
+ $Y=1.835 $X2=1.19 $Y2=2.9
r36 1 9 400 $w=1.7e-07 $l=4.49583e-07 $layer=licon1_PDIFF $count=1 $X=1.05
+ $Y=1.835 $X2=1.19 $Y2=2.22
.ends

.subckt PM_SKY130_FD_SC_LP__MUX2_4%A_317_367# 1 2 9 11 12 16
r30 11 16 4.09051 $w=1.7e-07 $l=1.57162e-07 $layer=LI1_cond $X=2.925 $Y=2.59
+ $X2=3.055 $Y2=2.53
r31 11 12 73.0695 $w=1.68e-07 $l=1.12e-06 $layer=LI1_cond $X=2.925 $Y=2.59
+ $X2=1.805 $Y2=2.59
r32 7 12 8.23557 $w=1.88e-07 $l=1.67183e-07 $layer=LI1_cond $X=1.675 $Y=2.505
+ $X2=1.805 $Y2=2.59
r33 7 9 13.519 $w=2.58e-07 $l=3.05e-07 $layer=LI1_cond $X=1.675 $Y=2.505
+ $X2=1.675 $Y2=2.2
r34 2 16 300 $w=1.7e-07 $l=7.74984e-07 $layer=licon1_PDIFF $count=2 $X=2.965
+ $Y=1.835 $X2=3.09 $Y2=2.55
r35 1 9 300 $w=1.7e-07 $l=4.22907e-07 $layer=licon1_PDIFF $count=2 $X=1.585
+ $Y=1.835 $X2=1.71 $Y2=2.2
.ends

.subckt PM_SKY130_FD_SC_LP__MUX2_4%X 1 2 3 4 15 19 23 24 25 26 29 33 37 39 42 43
+ 44 46 47 48
r66 47 48 18.9513 $w=2.23e-07 $l=3.7e-07 $layer=LI1_cond $X=5.547 $Y=0.555
+ $X2=5.547 $Y2=0.925
r67 45 48 7.17076 $w=2.23e-07 $l=1.4e-07 $layer=LI1_cond $X=5.547 $Y=1.065
+ $X2=5.547 $Y2=0.925
r68 45 46 4.27425 $w=2.12e-07 $l=8.5e-08 $layer=LI1_cond $X=5.547 $Y=1.065
+ $X2=5.547 $Y2=1.15
r69 41 46 4.27425 $w=2.12e-07 $l=9.12688e-08 $layer=LI1_cond $X=5.56 $Y=1.235
+ $X2=5.547 $Y2=1.15
r70 41 42 28.8364 $w=1.98e-07 $l=5.2e-07 $layer=LI1_cond $X=5.56 $Y=1.235
+ $X2=5.56 $Y2=1.755
r71 40 44 5.41628 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=4.895 $Y=1.84 $X2=4.805
+ $Y2=1.84
r72 39 42 6.87494 $w=1.7e-07 $l=1.36015e-07 $layer=LI1_cond $X=5.46 $Y=1.84
+ $X2=5.56 $Y2=1.755
r73 39 40 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=5.46 $Y=1.84
+ $X2=4.895 $Y2=1.84
r74 38 43 6.47928 $w=1.7e-07 $l=1.13e-07 $layer=LI1_cond $X=4.87 $Y=1.15
+ $X2=4.757 $Y2=1.15
r75 37 46 2.15711 $w=1.7e-07 $l=1.12e-07 $layer=LI1_cond $X=5.435 $Y=1.15
+ $X2=5.547 $Y2=1.15
r76 37 38 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=5.435 $Y=1.15
+ $X2=4.87 $Y2=1.15
r77 33 35 57.303 $w=1.78e-07 $l=9.3e-07 $layer=LI1_cond $X=4.805 $Y=1.98
+ $X2=4.805 $Y2=2.91
r78 31 44 1.13756 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=4.805 $Y=1.925
+ $X2=4.805 $Y2=1.84
r79 31 33 3.38889 $w=1.78e-07 $l=5.5e-08 $layer=LI1_cond $X=4.805 $Y=1.925
+ $X2=4.805 $Y2=1.98
r80 27 43 0.355529 $w=2.25e-07 $l=8.5e-08 $layer=LI1_cond $X=4.757 $Y=1.065
+ $X2=4.757 $Y2=1.15
r81 27 29 33.0367 $w=2.23e-07 $l=6.45e-07 $layer=LI1_cond $X=4.757 $Y=1.065
+ $X2=4.757 $Y2=0.42
r82 25 44 5.41628 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=4.715 $Y=1.84 $X2=4.805
+ $Y2=1.84
r83 25 26 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.715 $Y=1.84
+ $X2=4.045 $Y2=1.84
r84 23 43 6.47928 $w=1.7e-07 $l=1.12e-07 $layer=LI1_cond $X=4.645 $Y=1.15
+ $X2=4.757 $Y2=1.15
r85 23 24 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.645 $Y=1.15
+ $X2=3.975 $Y2=1.15
r86 19 21 54.2871 $w=1.88e-07 $l=9.3e-07 $layer=LI1_cond $X=3.95 $Y=1.98
+ $X2=3.95 $Y2=2.91
r87 17 26 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=3.95 $Y=1.925
+ $X2=4.045 $Y2=1.84
r88 17 19 3.21053 $w=1.88e-07 $l=5.5e-08 $layer=LI1_cond $X=3.95 $Y=1.925
+ $X2=3.95 $Y2=1.98
r89 13 24 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=3.87 $Y=1.065
+ $X2=3.975 $Y2=1.15
r90 13 15 34.0649 $w=2.08e-07 $l=6.45e-07 $layer=LI1_cond $X=3.87 $Y=1.065
+ $X2=3.87 $Y2=0.42
r91 4 35 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=4.67
+ $Y=1.835 $X2=4.81 $Y2=2.91
r92 4 33 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=4.67
+ $Y=1.835 $X2=4.81 $Y2=1.98
r93 3 21 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=3.81
+ $Y=1.835 $X2=3.95 $Y2=2.91
r94 3 19 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=3.81
+ $Y=1.835 $X2=3.95 $Y2=1.98
r95 2 29 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=4.6
+ $Y=0.235 $X2=4.74 $Y2=0.42
r96 1 15 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=3.74
+ $Y=0.235 $X2=3.88 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__MUX2_4%VGND 1 2 3 4 15 19 21 25 27 28 29 31 50 51 54
+ 59 62 64
r75 64 65 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r76 61 62 10.9708 $w=7.73e-07 $l=1.45e-07 $layer=LI1_cond $X=3.45 $Y=0.302
+ $X2=3.595 $Y2=0.302
r77 57 61 5.09298 $w=7.73e-07 $l=3.3e-07 $layer=LI1_cond $X=3.12 $Y=0.302
+ $X2=3.45 $Y2=0.302
r78 57 59 12.5141 $w=7.73e-07 $l=2.45e-07 $layer=LI1_cond $X=3.12 $Y=0.302
+ $X2=2.875 $Y2=0.302
r79 57 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r80 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r81 51 65 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=5.04
+ $Y2=0
r82 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r83 48 64 6.47928 $w=1.7e-07 $l=1.13e-07 $layer=LI1_cond $X=5.265 $Y=0 $X2=5.152
+ $Y2=0
r84 48 50 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=5.265 $Y=0 $X2=5.52
+ $Y2=0
r85 47 65 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=5.04
+ $Y2=0
r86 47 58 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.12
+ $Y2=0
r87 46 62 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=4.08 $Y=0 $X2=3.595
+ $Y2=0
r88 46 47 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r89 42 59 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=2.64 $Y=0 $X2=2.875
+ $Y2=0
r90 42 43 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r91 40 43 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r92 40 55 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r93 39 42 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r94 39 40 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r95 37 54 10.7288 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=1.33 $Y=0 $X2=1.1
+ $Y2=0
r96 37 39 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=1.33 $Y=0 $X2=1.68
+ $Y2=0
r97 34 55 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r98 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r99 31 54 10.7288 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=0.87 $Y=0 $X2=1.1
+ $Y2=0
r100 31 33 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=0.87 $Y=0 $X2=0.72
+ $Y2=0
r101 29 58 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.88 $Y=0
+ $X2=3.12 $Y2=0
r102 29 43 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.88 $Y=0
+ $X2=2.64 $Y2=0
r103 27 46 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=4.145 $Y=0 $X2=4.08
+ $Y2=0
r104 27 28 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.145 $Y=0 $X2=4.31
+ $Y2=0
r105 23 64 0.355529 $w=2.25e-07 $l=8.5e-08 $layer=LI1_cond $X=5.152 $Y=0.085
+ $X2=5.152 $Y2=0
r106 23 25 15.1098 $w=2.23e-07 $l=2.95e-07 $layer=LI1_cond $X=5.152 $Y=0.085
+ $X2=5.152 $Y2=0.38
r107 22 28 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.475 $Y=0 $X2=4.31
+ $Y2=0
r108 21 64 6.47928 $w=1.7e-07 $l=1.12e-07 $layer=LI1_cond $X=5.04 $Y=0 $X2=5.152
+ $Y2=0
r109 21 22 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=5.04 $Y=0 $X2=4.475
+ $Y2=0
r110 17 28 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.31 $Y=0.085
+ $X2=4.31 $Y2=0
r111 17 19 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=4.31 $Y=0.085
+ $X2=4.31 $Y2=0.38
r112 13 54 1.85547 $w=4.6e-07 $l=8.5e-08 $layer=LI1_cond $X=1.1 $Y=0.085 $X2=1.1
+ $Y2=0
r113 13 15 7.15047 $w=4.58e-07 $l=2.75e-07 $layer=LI1_cond $X=1.1 $Y=0.085
+ $X2=1.1 $Y2=0.36
r114 4 25 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.03
+ $Y=0.235 $X2=5.17 $Y2=0.38
r115 3 19 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.17
+ $Y=0.235 $X2=4.31 $Y2=0.38
r116 2 61 91 $w=1.7e-07 $l=6.79706e-07 $layer=licon1_NDIFF $count=2 $X=2.9
+ $Y=0.235 $X2=3.45 $Y2=0.525
r117 1 15 91 $w=1.7e-07 $l=2.60096e-07 $layer=licon1_NDIFF $count=2 $X=0.875
+ $Y=0.235 $X2=1.08 $Y2=0.36
.ends

