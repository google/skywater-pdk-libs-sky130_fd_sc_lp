* File: sky130_fd_sc_lp__or4_lp.spice
* Created: Fri Aug 28 11:25:18 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__or4_lp.pex.spice"
.subckt sky130_fd_sc_lp__or4_lp  VNB VPB D C B A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* B	B
* C	C
* D	D
* VPB	VPB
* VNB	VNB
MM1004 A_114_47# N_D_M1004_g N_A_27_47#_M1004_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1197 PD=0.63 PS=1.41 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1014 N_VGND_M1014_d N_D_M1014_g A_114_47# VNB NSHORT L=0.15 W=0.42 AD=0.0588
+ AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6 SB=75001.1
+ A=0.063 P=1.14 MULT=1
MM1005 A_272_47# N_C_M1005_g N_VGND_M1014_d VNB NSHORT L=0.15 W=0.42 AD=0.0441
+ AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75001 SB=75000.6 A=0.063
+ P=1.14 MULT=1
MM1006 N_A_27_47#_M1006_d N_C_M1006_g A_272_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.1533 AS=0.0441 PD=1.57 PS=0.63 NRD=22.848 NRS=14.28 M=1 R=2.8 SA=75001.4
+ SB=75000.3 A=0.063 P=1.14 MULT=1
MM1011 A_465_185# N_B_M1011_g N_VGND_M1011_s VNB NSHORT L=0.15 W=0.42
+ AD=0.076125 AS=0.1197 PD=0.835 PS=1.41 NRD=36.06 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.8 A=0.063 P=1.14 MULT=1
MM1010 N_A_27_47#_M1010_d N_B_M1010_g A_465_185# VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.076125 PD=0.7 PS=0.835 NRD=0 NRS=36.06 M=1 R=2.8 SA=75000.6
+ SB=75001.8 A=0.063 P=1.14 MULT=1
MM1003 A_646_167# N_A_M1003_g N_A_27_47#_M1010_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75001
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1000 N_VGND_M1000_d N_A_M1000_g A_646_167# VNB NSHORT L=0.15 W=0.42 AD=0.0588
+ AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.4 SB=75001 A=0.063
+ P=1.14 MULT=1
MM1002 A_804_167# N_A_27_47#_M1002_g N_VGND_M1000_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75001.8
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1013 N_X_M1013_d N_A_27_47#_M1013_g A_804_167# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75002.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1001 A_154_419# N_D_M1001_g N_A_27_47#_M1001_s VPB PHIGHVT L=0.25 W=1 AD=0.12
+ AS=0.285 PD=1.24 PS=2.57 NRD=12.7853 NRS=0 M=1 R=4 SA=125000 SB=125003 A=0.25
+ P=2.5 MULT=1
MM1009 A_252_419# N_C_M1009_g A_154_419# VPB PHIGHVT L=0.25 W=1 AD=0.16 AS=0.12
+ PD=1.32 PS=1.24 NRD=20.6653 NRS=12.7853 M=1 R=4 SA=125001 SB=125003 A=0.25
+ P=2.5 MULT=1
MM1007 A_366_419# N_B_M1007_g A_252_419# VPB PHIGHVT L=0.25 W=1 AD=0.605 AS=0.16
+ PD=2.21 PS=1.32 NRD=108.33 NRS=20.6653 M=1 R=4 SA=125001 SB=125002 A=0.25
+ P=2.5 MULT=1
MM1012 N_VPWR_M1012_d N_A_M1012_g A_366_419# VPB PHIGHVT L=0.25 W=1 AD=0.2825
+ AS=0.605 PD=1.565 PS=2.21 NRD=56.145 NRS=108.33 M=1 R=4 SA=125003 SB=125001
+ A=0.25 P=2.5 MULT=1
MM1008 N_X_M1008_d N_A_27_47#_M1008_g N_VPWR_M1012_d VPB PHIGHVT L=0.25 W=1
+ AD=0.285 AS=0.2825 PD=2.57 PS=1.565 NRD=0 NRS=0 M=1 R=4 SA=125003 SB=125000
+ A=0.25 P=2.5 MULT=1
DX15_noxref VNB VPB NWDIODE A=9.0679 P=14.61
*
.include "sky130_fd_sc_lp__or4_lp.pxi.spice"
*
.ends
*
*
