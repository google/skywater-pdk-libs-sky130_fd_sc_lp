* File: sky130_fd_sc_lp__a22o_lp.pxi.spice
* Created: Wed Sep  2 09:22:46 2020
* 
x_PM_SKY130_FD_SC_LP__A22O_LP%A1 N_A1_M1009_g N_A1_M1008_g N_A1_c_73_n
+ N_A1_c_74_n N_A1_c_75_n N_A1_c_76_n A1 A1 N_A1_c_78_n
+ PM_SKY130_FD_SC_LP__A22O_LP%A1
x_PM_SKY130_FD_SC_LP__A22O_LP%B2 N_B2_M1006_g N_B2_M1005_g N_B2_c_134_n
+ N_B2_c_139_n B2 N_B2_c_136_n PM_SKY130_FD_SC_LP__A22O_LP%B2
x_PM_SKY130_FD_SC_LP__A22O_LP%B1 N_B1_M1004_g N_B1_c_178_n N_B1_M1000_g
+ N_B1_c_179_n N_B1_c_180_n B1 B1 N_B1_c_182_n PM_SKY130_FD_SC_LP__A22O_LP%B1
x_PM_SKY130_FD_SC_LP__A22O_LP%A2 N_A2_c_233_n N_A2_M1007_g N_A2_M1001_g
+ N_A2_c_230_n A2 A2 N_A2_c_232_n PM_SKY130_FD_SC_LP__A22O_LP%A2
x_PM_SKY130_FD_SC_LP__A22O_LP%A_243_409# N_A_243_409#_M1004_d
+ N_A_243_409#_M1006_d N_A_243_409#_c_276_n N_A_243_409#_M1002_g
+ N_A_243_409#_M1010_g N_A_243_409#_M1003_g N_A_243_409#_c_278_n
+ N_A_243_409#_c_279_n N_A_243_409#_c_301_n N_A_243_409#_c_280_n
+ N_A_243_409#_c_289_n N_A_243_409#_c_290_n N_A_243_409#_c_281_n
+ N_A_243_409#_c_349_p N_A_243_409#_c_282_n N_A_243_409#_c_283_n
+ N_A_243_409#_c_284_n N_A_243_409#_c_285_n N_A_243_409#_c_286_n
+ N_A_243_409#_c_287_n PM_SKY130_FD_SC_LP__A22O_LP%A_243_409#
x_PM_SKY130_FD_SC_LP__A22O_LP%VPWR N_VPWR_M1009_s N_VPWR_M1007_d N_VPWR_c_379_n
+ N_VPWR_c_380_n N_VPWR_c_381_n VPWR N_VPWR_c_382_n N_VPWR_c_383_n
+ N_VPWR_c_378_n N_VPWR_c_385_n PM_SKY130_FD_SC_LP__A22O_LP%VPWR
x_PM_SKY130_FD_SC_LP__A22O_LP%A_137_409# N_A_137_409#_M1009_d
+ N_A_137_409#_M1000_d N_A_137_409#_c_416_n N_A_137_409#_c_419_n
+ N_A_137_409#_c_417_n N_A_137_409#_c_426_n
+ PM_SKY130_FD_SC_LP__A22O_LP%A_137_409#
x_PM_SKY130_FD_SC_LP__A22O_LP%X N_X_M1003_d N_X_M1010_d N_X_c_444_n N_X_c_445_n
+ X X X N_X_c_448_n PM_SKY130_FD_SC_LP__A22O_LP%X
x_PM_SKY130_FD_SC_LP__A22O_LP%VGND N_VGND_M1005_s N_VGND_M1001_d N_VGND_c_468_n
+ N_VGND_c_469_n N_VGND_c_470_n N_VGND_c_471_n VGND N_VGND_c_472_n
+ N_VGND_c_473_n N_VGND_c_474_n PM_SKY130_FD_SC_LP__A22O_LP%VGND
cc_1 VNB N_A1_M1008_g 0.0225013f $X=-0.19 $Y=-0.245 $X2=1.87 $Y2=0.445
cc_2 VNB N_A1_c_73_n 0.0023438f $X=-0.19 $Y=-0.245 $X2=0.42 $Y2=1.625
cc_3 VNB N_A1_c_74_n 0.0296981f $X=-0.19 $Y=-0.245 $X2=1.795 $Y2=0.94
cc_4 VNB N_A1_c_75_n 0.00443866f $X=-0.19 $Y=-0.245 $X2=1.96 $Y2=0.94
cc_5 VNB N_A1_c_76_n 0.0332563f $X=-0.19 $Y=-0.245 $X2=1.96 $Y2=1.02
cc_6 VNB A1 0.0526351f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_7 VNB N_A1_c_78_n 0.0490126f $X=-0.19 $Y=-0.245 $X2=0.42 $Y2=1.285
cc_8 VNB N_B2_M1005_g 0.0488336f $X=-0.19 $Y=-0.245 $X2=1.87 $Y2=0.445
cc_9 VNB N_B2_c_134_n 0.017356f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=0.94
cc_10 VNB B2 0.00843345f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_B2_c_136_n 0.0145509f $X=-0.19 $Y=-0.245 $X2=1.96 $Y2=1.02
cc_12 VNB N_B1_c_178_n 0.035232f $X=-0.19 $Y=-0.245 $X2=1.87 $Y2=0.855
cc_13 VNB N_B1_c_179_n 0.014304f $X=-0.19 $Y=-0.245 $X2=1.795 $Y2=0.94
cc_14 VNB N_B1_c_180_n 0.0120969f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=0.94
cc_15 VNB B1 0.00966382f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_B1_c_182_n 0.0331683f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_17 VNB N_A2_M1001_g 0.0375775f $X=-0.19 $Y=-0.245 $X2=1.87 $Y2=0.445
cc_18 VNB N_A2_c_230_n 0.0312946f $X=-0.19 $Y=-0.245 $X2=0.42 $Y2=1.625
cc_19 VNB A2 0.00257517f $X=-0.19 $Y=-0.245 $X2=1.795 $Y2=0.94
cc_20 VNB N_A2_c_232_n 0.0298934f $X=-0.19 $Y=-0.245 $X2=1.96 $Y2=1.02
cc_21 VNB N_A_243_409#_c_276_n 0.0322144f $X=-0.19 $Y=-0.245 $X2=1.87 $Y2=0.445
cc_22 VNB N_A_243_409#_M1010_g 0.0135888f $X=-0.19 $Y=-0.245 $X2=1.96 $Y2=0.94
cc_23 VNB N_A_243_409#_c_278_n 0.0219435f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_24 VNB N_A_243_409#_c_279_n 0.0181343f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_243_409#_c_280_n 0.00739286f $X=-0.19 $Y=-0.245 $X2=1.96 $Y2=1.02
cc_26 VNB N_A_243_409#_c_281_n 0.0121136f $X=-0.19 $Y=-0.245 $X2=0.355 $Y2=1.285
cc_27 VNB N_A_243_409#_c_282_n 0.0031548f $X=-0.19 $Y=-0.245 $X2=0.355 $Y2=1.665
cc_28 VNB N_A_243_409#_c_283_n 0.00128319f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_243_409#_c_284_n 0.002408f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_243_409#_c_285_n 0.00489436f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_243_409#_c_286_n 0.0302797f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_243_409#_c_287_n 0.00182462f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VPWR_c_378_n 0.163682f $X=-0.19 $Y=-0.245 $X2=0.355 $Y2=1.285
cc_34 VNB N_X_c_444_n 0.0493798f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_X_c_445_n 0.0126713f $X=-0.19 $Y=-0.245 $X2=1.795 $Y2=0.94
cc_36 VNB N_VGND_c_468_n 0.022137f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=0.94
cc_37 VNB N_VGND_c_469_n 0.00240024f $X=-0.19 $Y=-0.245 $X2=1.96 $Y2=1.02
cc_38 VNB N_VGND_c_470_n 0.0449204f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_39 VNB N_VGND_c_471_n 0.00356964f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_40 VNB N_VGND_c_472_n 0.027824f $X=-0.19 $Y=-0.245 $X2=0.355 $Y2=1.285
cc_41 VNB N_VGND_c_473_n 0.22561f $X=-0.19 $Y=-0.245 $X2=0.355 $Y2=1.295
cc_42 VNB N_VGND_c_474_n 0.0285983f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VPB N_A1_M1009_g 0.0292395f $X=-0.19 $Y=1.655 $X2=0.56 $Y2=2.545
cc_44 VPB N_A1_c_73_n 0.0328914f $X=-0.19 $Y=1.655 $X2=0.42 $Y2=1.625
cc_45 VPB A1 0.009783f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_46 VPB N_B2_M1006_g 0.0295436f $X=-0.19 $Y=1.655 $X2=0.56 $Y2=2.545
cc_47 VPB N_B2_c_134_n 0.00361493f $X=-0.19 $Y=1.655 $X2=0.585 $Y2=0.94
cc_48 VPB N_B2_c_139_n 0.0134174f $X=-0.19 $Y=1.655 $X2=1.96 $Y2=0.94
cc_49 VPB B2 0.007911f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_50 VPB N_B1_M1000_g 0.0263559f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_51 VPB B1 0.00569959f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_52 VPB N_B1_c_182_n 0.0253978f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_53 VPB N_A2_c_233_n 0.0243801f $X=-0.19 $Y=1.655 $X2=0.56 $Y2=1.915
cc_54 VPB N_A2_c_230_n 0.0292302f $X=-0.19 $Y=1.655 $X2=0.42 $Y2=1.625
cc_55 VPB A2 0.00195292f $X=-0.19 $Y=1.655 $X2=1.795 $Y2=0.94
cc_56 VPB N_A_243_409#_M1010_g 0.0462863f $X=-0.19 $Y=1.655 $X2=1.96 $Y2=0.94
cc_57 VPB N_A_243_409#_c_289_n 0.0118733f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_58 VPB N_A_243_409#_c_290_n 0.00370004f $X=-0.19 $Y=1.655 $X2=0.585 $Y2=0.94
cc_59 VPB N_A_243_409#_c_283_n 0.00292443f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_60 VPB N_VPWR_c_379_n 0.0118353f $X=-0.19 $Y=1.655 $X2=1.87 $Y2=0.445
cc_61 VPB N_VPWR_c_380_n 0.0467213f $X=-0.19 $Y=1.655 $X2=0.42 $Y2=1.625
cc_62 VPB N_VPWR_c_381_n 0.00423313f $X=-0.19 $Y=1.655 $X2=1.96 $Y2=1.02
cc_63 VPB N_VPWR_c_382_n 0.0495494f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_64 VPB N_VPWR_c_383_n 0.0287692f $X=-0.19 $Y=1.655 $X2=0.585 $Y2=0.94
cc_65 VPB N_VPWR_c_378_n 0.0656179f $X=-0.19 $Y=1.655 $X2=0.355 $Y2=1.285
cc_66 VPB N_VPWR_c_385_n 0.00548753f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_67 VPB N_A_137_409#_c_416_n 0.00207453f $X=-0.19 $Y=1.655 $X2=1.87 $Y2=0.445
cc_68 VPB N_A_137_409#_c_417_n 0.00647109f $X=-0.19 $Y=1.655 $X2=0.585 $Y2=0.94
cc_69 VPB N_X_c_444_n 0.0129405f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_70 VPB X 0.0378954f $X=-0.19 $Y=1.655 $X2=1.96 $Y2=1.02
cc_71 VPB N_X_c_448_n 0.020717f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_72 N_A1_c_73_n N_B2_M1006_g 0.0156939f $X=0.42 $Y=1.625 $X2=0 $Y2=0
cc_73 N_A1_c_74_n N_B2_M1005_g 0.0138282f $X=1.795 $Y=0.94 $X2=0 $Y2=0
cc_74 A1 N_B2_M1005_g 0.00306983f $X=0.155 $Y=1.58 $X2=0 $Y2=0
cc_75 N_A1_c_78_n N_B2_M1005_g 0.0022955f $X=0.42 $Y=1.285 $X2=0 $Y2=0
cc_76 N_A1_c_73_n N_B2_c_134_n 0.0116189f $X=0.42 $Y=1.625 $X2=0 $Y2=0
cc_77 N_A1_c_73_n N_B2_c_139_n 0.00525144f $X=0.42 $Y=1.625 $X2=0 $Y2=0
cc_78 N_A1_c_73_n B2 5.83977e-19 $X=0.42 $Y=1.625 $X2=0 $Y2=0
cc_79 N_A1_c_74_n B2 0.0318021f $X=1.795 $Y=0.94 $X2=0 $Y2=0
cc_80 A1 B2 0.0284109f $X=0.155 $Y=1.58 $X2=0 $Y2=0
cc_81 N_A1_c_78_n B2 7.45647e-19 $X=0.42 $Y=1.285 $X2=0 $Y2=0
cc_82 N_A1_c_74_n N_B2_c_136_n 0.00468021f $X=1.795 $Y=0.94 $X2=0 $Y2=0
cc_83 A1 N_B2_c_136_n 7.44797e-19 $X=0.155 $Y=1.58 $X2=0 $Y2=0
cc_84 N_A1_c_78_n N_B2_c_136_n 0.0116189f $X=0.42 $Y=1.285 $X2=0 $Y2=0
cc_85 N_A1_c_74_n N_B1_c_178_n 0.0110666f $X=1.795 $Y=0.94 $X2=0 $Y2=0
cc_86 N_A1_c_75_n N_B1_c_178_n 0.00107336f $X=1.96 $Y=0.94 $X2=0 $Y2=0
cc_87 N_A1_c_76_n N_B1_c_178_n 0.0148465f $X=1.96 $Y=1.02 $X2=0 $Y2=0
cc_88 N_A1_M1008_g N_B1_c_179_n 0.0116433f $X=1.87 $Y=0.445 $X2=0 $Y2=0
cc_89 N_A1_M1008_g N_B1_c_180_n 0.0148465f $X=1.87 $Y=0.445 $X2=0 $Y2=0
cc_90 N_A1_c_74_n N_B1_c_180_n 0.00618001f $X=1.795 $Y=0.94 $X2=0 $Y2=0
cc_91 N_A1_c_74_n B1 0.00863458f $X=1.795 $Y=0.94 $X2=0 $Y2=0
cc_92 N_A1_c_75_n B1 0.0180619f $X=1.96 $Y=0.94 $X2=0 $Y2=0
cc_93 N_A1_c_76_n B1 0.00115092f $X=1.96 $Y=1.02 $X2=0 $Y2=0
cc_94 N_A1_c_74_n N_B1_c_182_n 0.0038114f $X=1.795 $Y=0.94 $X2=0 $Y2=0
cc_95 N_A1_c_75_n N_B1_c_182_n 6.81663e-19 $X=1.96 $Y=0.94 $X2=0 $Y2=0
cc_96 N_A1_c_76_n N_B1_c_182_n 0.00916657f $X=1.96 $Y=1.02 $X2=0 $Y2=0
cc_97 N_A1_M1008_g N_A2_M1001_g 0.0211718f $X=1.87 $Y=0.445 $X2=0 $Y2=0
cc_98 N_A1_c_75_n N_A2_M1001_g 0.00151074f $X=1.96 $Y=0.94 $X2=0 $Y2=0
cc_99 N_A1_c_76_n N_A2_M1001_g 0.0179896f $X=1.96 $Y=1.02 $X2=0 $Y2=0
cc_100 N_A1_c_75_n A2 0.00264671f $X=1.96 $Y=0.94 $X2=0 $Y2=0
cc_101 N_A1_M1008_g N_A_243_409#_c_280_n 0.00894269f $X=1.87 $Y=0.445 $X2=0
+ $Y2=0
cc_102 N_A1_c_75_n N_A_243_409#_c_280_n 0.0209137f $X=1.96 $Y=0.94 $X2=0 $Y2=0
cc_103 N_A1_c_76_n N_A_243_409#_c_280_n 0.00124625f $X=1.96 $Y=1.02 $X2=0 $Y2=0
cc_104 N_A1_M1008_g N_A_243_409#_c_284_n 0.00614365f $X=1.87 $Y=0.445 $X2=0
+ $Y2=0
cc_105 N_A1_c_74_n N_A_243_409#_c_284_n 0.022471f $X=1.795 $Y=0.94 $X2=0 $Y2=0
cc_106 N_A1_c_75_n N_A_243_409#_c_284_n 0.00163817f $X=1.96 $Y=0.94 $X2=0 $Y2=0
cc_107 N_A1_M1008_g N_A_243_409#_c_285_n 0.00328422f $X=1.87 $Y=0.445 $X2=0
+ $Y2=0
cc_108 N_A1_c_75_n N_A_243_409#_c_285_n 0.00647895f $X=1.96 $Y=0.94 $X2=0 $Y2=0
cc_109 N_A1_c_76_n N_A_243_409#_c_285_n 5.11076e-19 $X=1.96 $Y=1.02 $X2=0 $Y2=0
cc_110 N_A1_M1009_g N_VPWR_c_380_n 0.0238571f $X=0.56 $Y=2.545 $X2=0 $Y2=0
cc_111 N_A1_c_73_n N_VPWR_c_380_n 0.00135666f $X=0.42 $Y=1.625 $X2=0 $Y2=0
cc_112 A1 N_VPWR_c_380_n 0.02336f $X=0.155 $Y=1.58 $X2=0 $Y2=0
cc_113 N_A1_M1009_g N_VPWR_c_382_n 0.00767656f $X=0.56 $Y=2.545 $X2=0 $Y2=0
cc_114 N_A1_M1009_g N_VPWR_c_378_n 0.0134103f $X=0.56 $Y=2.545 $X2=0 $Y2=0
cc_115 N_A1_M1009_g N_A_137_409#_c_416_n 0.00348959f $X=0.56 $Y=2.545 $X2=0
+ $Y2=0
cc_116 N_A1_M1009_g N_A_137_409#_c_419_n 0.0157568f $X=0.56 $Y=2.545 $X2=0 $Y2=0
cc_117 N_A1_c_74_n N_VGND_c_468_n 0.0257555f $X=1.795 $Y=0.94 $X2=0 $Y2=0
cc_118 N_A1_M1008_g N_VGND_c_470_n 0.00399692f $X=1.87 $Y=0.445 $X2=0 $Y2=0
cc_119 N_A1_M1008_g N_VGND_c_473_n 0.00604037f $X=1.87 $Y=0.445 $X2=0 $Y2=0
cc_120 N_A1_c_74_n N_VGND_c_473_n 0.0193561f $X=1.795 $Y=0.94 $X2=0 $Y2=0
cc_121 N_A1_c_75_n N_VGND_c_473_n 4.57254e-19 $X=1.96 $Y=0.94 $X2=0 $Y2=0
cc_122 A1 N_VGND_c_473_n 0.00661595f $X=0.155 $Y=1.58 $X2=0 $Y2=0
cc_123 N_B2_M1005_g N_B1_c_178_n 0.013492f $X=1.05 $Y=0.445 $X2=0 $Y2=0
cc_124 B2 N_B1_c_178_n 0.0074215f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_125 N_B2_c_136_n N_B1_c_178_n 0.0119851f $X=1.06 $Y=1.37 $X2=0 $Y2=0
cc_126 N_B2_M1005_g N_B1_c_179_n 0.0415082f $X=1.05 $Y=0.445 $X2=0 $Y2=0
cc_127 N_B2_c_134_n B1 8.20615e-19 $X=1.06 $Y=1.71 $X2=0 $Y2=0
cc_128 B2 B1 0.0219668f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_129 N_B2_M1006_g N_B1_c_182_n 0.0177136f $X=1.09 $Y=2.545 $X2=0 $Y2=0
cc_130 N_B2_c_134_n N_B1_c_182_n 0.0170921f $X=1.06 $Y=1.71 $X2=0 $Y2=0
cc_131 N_B2_c_139_n N_B1_c_182_n 0.00149132f $X=1.06 $Y=1.875 $X2=0 $Y2=0
cc_132 B2 N_B1_c_182_n 0.00249351f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_133 N_B2_M1006_g N_A_243_409#_c_301_n 0.00635916f $X=1.09 $Y=2.545 $X2=0
+ $Y2=0
cc_134 N_B2_M1006_g N_A_243_409#_c_290_n 0.00328213f $X=1.09 $Y=2.545 $X2=0
+ $Y2=0
cc_135 N_B2_M1005_g N_A_243_409#_c_284_n 0.0010756f $X=1.05 $Y=0.445 $X2=0 $Y2=0
cc_136 N_B2_M1006_g N_VPWR_c_380_n 0.00103922f $X=1.09 $Y=2.545 $X2=0 $Y2=0
cc_137 N_B2_M1006_g N_VPWR_c_382_n 0.00546179f $X=1.09 $Y=2.545 $X2=0 $Y2=0
cc_138 N_B2_M1006_g N_VPWR_c_378_n 0.00782141f $X=1.09 $Y=2.545 $X2=0 $Y2=0
cc_139 N_B2_M1006_g N_A_137_409#_c_416_n 8.05528e-19 $X=1.09 $Y=2.545 $X2=0
+ $Y2=0
cc_140 N_B2_M1006_g N_A_137_409#_c_419_n 0.022245f $X=1.09 $Y=2.545 $X2=0 $Y2=0
cc_141 N_B2_c_139_n N_A_137_409#_c_419_n 0.00168897f $X=1.06 $Y=1.875 $X2=0
+ $Y2=0
cc_142 B2 N_A_137_409#_c_419_n 0.00525522f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_143 N_B2_M1006_g N_A_137_409#_c_417_n 0.0184508f $X=1.09 $Y=2.545 $X2=0 $Y2=0
cc_144 N_B2_M1005_g N_VGND_c_468_n 0.0146339f $X=1.05 $Y=0.445 $X2=0 $Y2=0
cc_145 N_B2_M1005_g N_VGND_c_470_n 0.00486043f $X=1.05 $Y=0.445 $X2=0 $Y2=0
cc_146 N_B2_M1005_g N_VGND_c_473_n 0.00456945f $X=1.05 $Y=0.445 $X2=0 $Y2=0
cc_147 N_B1_M1000_g N_A2_c_233_n 0.0162468f $X=1.925 $Y=2.545 $X2=-0.19
+ $Y2=-0.245
cc_148 B1 N_A2_c_230_n 0.00351359f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_149 N_B1_c_182_n N_A2_c_230_n 0.0250722f $X=1.785 $Y=1.615 $X2=0 $Y2=0
cc_150 B1 A2 0.0265518f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_151 N_B1_c_182_n A2 3.1711e-19 $X=1.785 $Y=1.615 $X2=0 $Y2=0
cc_152 N_B1_M1000_g N_A_243_409#_c_301_n 0.010498f $X=1.925 $Y=2.545 $X2=0 $Y2=0
cc_153 N_B1_M1000_g N_A_243_409#_c_289_n 0.0176036f $X=1.925 $Y=2.545 $X2=0
+ $Y2=0
cc_154 B1 N_A_243_409#_c_289_n 0.0309807f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_155 N_B1_M1000_g N_A_243_409#_c_290_n 0.00186615f $X=1.925 $Y=2.545 $X2=0
+ $Y2=0
cc_156 B1 N_A_243_409#_c_290_n 0.0198961f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_157 N_B1_c_182_n N_A_243_409#_c_290_n 0.00715407f $X=1.785 $Y=1.615 $X2=0
+ $Y2=0
cc_158 N_B1_c_179_n N_A_243_409#_c_284_n 0.00728765f $X=1.475 $Y=0.73 $X2=0
+ $Y2=0
cc_159 N_B1_c_180_n N_A_243_409#_c_284_n 0.00216596f $X=1.475 $Y=0.88 $X2=0
+ $Y2=0
cc_160 N_B1_M1000_g N_VPWR_c_381_n 8.6872e-19 $X=1.925 $Y=2.545 $X2=0 $Y2=0
cc_161 N_B1_M1000_g N_VPWR_c_382_n 0.00546179f $X=1.925 $Y=2.545 $X2=0 $Y2=0
cc_162 N_B1_M1000_g N_VPWR_c_378_n 0.00782141f $X=1.925 $Y=2.545 $X2=0 $Y2=0
cc_163 N_B1_M1000_g N_A_137_409#_c_417_n 0.0185321f $X=1.925 $Y=2.545 $X2=0
+ $Y2=0
cc_164 N_B1_M1000_g N_A_137_409#_c_426_n 0.015383f $X=1.925 $Y=2.545 $X2=0 $Y2=0
cc_165 N_B1_c_179_n N_VGND_c_468_n 0.0024608f $X=1.475 $Y=0.73 $X2=0 $Y2=0
cc_166 N_B1_c_179_n N_VGND_c_470_n 0.00550269f $X=1.475 $Y=0.73 $X2=0 $Y2=0
cc_167 N_B1_c_179_n N_VGND_c_473_n 0.00633508f $X=1.475 $Y=0.73 $X2=0 $Y2=0
cc_168 N_A2_M1001_g N_A_243_409#_c_276_n 0.0185847f $X=2.44 $Y=0.445 $X2=0 $Y2=0
cc_169 N_A2_c_230_n N_A_243_409#_M1010_g 0.0339811f $X=2.575 $Y=1.585 $X2=0
+ $Y2=0
cc_170 A2 N_A_243_409#_M1010_g 3.64151e-19 $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_171 N_A2_c_230_n N_A_243_409#_c_279_n 0.00772626f $X=2.575 $Y=1.585 $X2=0
+ $Y2=0
cc_172 N_A2_c_233_n N_A_243_409#_c_301_n 8.17244e-19 $X=2.455 $Y=1.92 $X2=0
+ $Y2=0
cc_173 N_A2_M1001_g N_A_243_409#_c_280_n 4.53244e-19 $X=2.44 $Y=0.445 $X2=0
+ $Y2=0
cc_174 N_A2_c_233_n N_A_243_409#_c_289_n 0.0256738f $X=2.455 $Y=1.92 $X2=0 $Y2=0
cc_175 N_A2_c_230_n N_A_243_409#_c_289_n 0.00140343f $X=2.575 $Y=1.585 $X2=0
+ $Y2=0
cc_176 A2 N_A_243_409#_c_289_n 0.0245995f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_177 N_A2_M1001_g N_A_243_409#_c_281_n 0.00521765f $X=2.44 $Y=0.445 $X2=0
+ $Y2=0
cc_178 A2 N_A_243_409#_c_281_n 0.0234643f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_179 N_A2_c_232_n N_A_243_409#_c_281_n 0.00185006f $X=2.62 $Y=1.29 $X2=0 $Y2=0
cc_180 N_A2_M1001_g N_A_243_409#_c_282_n 0.00345777f $X=2.44 $Y=0.445 $X2=0
+ $Y2=0
cc_181 A2 N_A_243_409#_c_282_n 0.0497339f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_182 N_A2_c_232_n N_A_243_409#_c_282_n 0.00223653f $X=2.62 $Y=1.29 $X2=0 $Y2=0
cc_183 N_A2_c_230_n N_A_243_409#_c_283_n 0.00323451f $X=2.575 $Y=1.585 $X2=0
+ $Y2=0
cc_184 N_A2_M1001_g N_A_243_409#_c_284_n 9.60447e-19 $X=2.44 $Y=0.445 $X2=0
+ $Y2=0
cc_185 N_A2_M1001_g N_A_243_409#_c_285_n 0.0179992f $X=2.44 $Y=0.445 $X2=0 $Y2=0
cc_186 A2 N_A_243_409#_c_285_n 0.00140639f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_187 N_A2_M1001_g N_A_243_409#_c_286_n 0.00410713f $X=2.44 $Y=0.445 $X2=0
+ $Y2=0
cc_188 A2 N_A_243_409#_c_286_n 3.53464e-19 $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_189 N_A2_c_232_n N_A_243_409#_c_286_n 0.00772626f $X=2.62 $Y=1.29 $X2=0 $Y2=0
cc_190 N_A2_c_230_n N_A_243_409#_c_287_n 0.00223653f $X=2.575 $Y=1.585 $X2=0
+ $Y2=0
cc_191 N_A2_c_233_n N_VPWR_c_381_n 0.0178662f $X=2.455 $Y=1.92 $X2=0 $Y2=0
cc_192 N_A2_c_233_n N_VPWR_c_382_n 0.00767656f $X=2.455 $Y=1.92 $X2=0 $Y2=0
cc_193 N_A2_c_233_n N_VPWR_c_378_n 0.0134103f $X=2.455 $Y=1.92 $X2=0 $Y2=0
cc_194 N_A2_c_233_n N_A_137_409#_c_417_n 0.00348959f $X=2.455 $Y=1.92 $X2=0
+ $Y2=0
cc_195 N_A2_c_233_n N_A_137_409#_c_426_n 0.0105402f $X=2.455 $Y=1.92 $X2=0 $Y2=0
cc_196 N_A2_M1001_g N_VGND_c_469_n 0.00951671f $X=2.44 $Y=0.445 $X2=0 $Y2=0
cc_197 N_A2_M1001_g N_VGND_c_470_n 0.00453961f $X=2.44 $Y=0.445 $X2=0 $Y2=0
cc_198 N_A2_M1001_g N_VGND_c_473_n 0.00647231f $X=2.44 $Y=0.445 $X2=0 $Y2=0
cc_199 N_A_243_409#_c_289_n N_VPWR_M1007_d 0.00963132f $X=2.965 $Y=2.06 $X2=0
+ $Y2=0
cc_200 N_A_243_409#_M1010_g N_VPWR_c_381_n 0.0105297f $X=3.215 $Y=2.545 $X2=0
+ $Y2=0
cc_201 N_A_243_409#_c_289_n N_VPWR_c_381_n 0.0209601f $X=2.965 $Y=2.06 $X2=0
+ $Y2=0
cc_202 N_A_243_409#_M1010_g N_VPWR_c_383_n 0.0086001f $X=3.215 $Y=2.545 $X2=0
+ $Y2=0
cc_203 N_A_243_409#_M1010_g N_VPWR_c_378_n 0.0167976f $X=3.215 $Y=2.545 $X2=0
+ $Y2=0
cc_204 N_A_243_409#_c_289_n N_A_137_409#_M1000_d 0.00180746f $X=2.965 $Y=2.06
+ $X2=0 $Y2=0
cc_205 N_A_243_409#_c_301_n N_A_137_409#_c_419_n 0.0189644f $X=1.66 $Y=2.19
+ $X2=0 $Y2=0
cc_206 N_A_243_409#_c_290_n N_A_137_409#_c_419_n 0.003186f $X=1.825 $Y=2.06
+ $X2=0 $Y2=0
cc_207 N_A_243_409#_M1006_d N_A_137_409#_c_417_n 0.0130537f $X=1.215 $Y=2.045
+ $X2=0 $Y2=0
cc_208 N_A_243_409#_c_301_n N_A_137_409#_c_417_n 0.0195297f $X=1.66 $Y=2.19
+ $X2=0 $Y2=0
cc_209 N_A_243_409#_c_301_n N_A_137_409#_c_426_n 0.0256974f $X=1.66 $Y=2.19
+ $X2=0 $Y2=0
cc_210 N_A_243_409#_c_289_n N_A_137_409#_c_426_n 0.0163515f $X=2.965 $Y=2.06
+ $X2=0 $Y2=0
cc_211 N_A_243_409#_c_276_n N_X_c_444_n 0.0223924f $X=2.955 $Y=0.735 $X2=0 $Y2=0
cc_212 N_A_243_409#_M1010_g N_X_c_444_n 0.010706f $X=3.215 $Y=2.545 $X2=0 $Y2=0
cc_213 N_A_243_409#_c_349_p N_X_c_444_n 0.0129665f $X=3.17 $Y=0.945 $X2=0 $Y2=0
cc_214 N_A_243_409#_c_282_n N_X_c_444_n 0.0364858f $X=3.17 $Y=1.24 $X2=0 $Y2=0
cc_215 N_A_243_409#_c_283_n N_X_c_444_n 0.0172578f $X=3.05 $Y=1.975 $X2=0 $Y2=0
cc_216 N_A_243_409#_c_276_n N_X_c_445_n 0.00771167f $X=2.955 $Y=0.735 $X2=0
+ $Y2=0
cc_217 N_A_243_409#_M1010_g X 0.0192609f $X=3.215 $Y=2.545 $X2=0 $Y2=0
cc_218 N_A_243_409#_M1010_g N_X_c_448_n 0.00957846f $X=3.215 $Y=2.545 $X2=0
+ $Y2=0
cc_219 N_A_243_409#_c_279_n N_X_c_448_n 0.00166869f $X=3.232 $Y=1.445 $X2=0
+ $Y2=0
cc_220 N_A_243_409#_c_289_n N_X_c_448_n 0.0117249f $X=2.965 $Y=2.06 $X2=0 $Y2=0
cc_221 N_A_243_409#_c_283_n N_X_c_448_n 0.00235233f $X=3.05 $Y=1.975 $X2=0 $Y2=0
cc_222 N_A_243_409#_c_287_n N_X_c_448_n 0.00195687f $X=3.17 $Y=1.445 $X2=0 $Y2=0
cc_223 N_A_243_409#_c_284_n N_VGND_c_468_n 0.0120387f $X=1.655 $Y=0.445 $X2=0
+ $Y2=0
cc_224 N_A_243_409#_c_276_n N_VGND_c_469_n 0.0131628f $X=2.955 $Y=0.735 $X2=0
+ $Y2=0
cc_225 N_A_243_409#_c_281_n N_VGND_c_469_n 0.0163712f $X=2.965 $Y=0.86 $X2=0
+ $Y2=0
cc_226 N_A_243_409#_c_285_n N_VGND_c_469_n 0.00623204f $X=2.39 $Y=0.59 $X2=0
+ $Y2=0
cc_227 N_A_243_409#_c_280_n N_VGND_c_470_n 0.0108713f $X=2.305 $Y=0.59 $X2=0
+ $Y2=0
cc_228 N_A_243_409#_c_284_n N_VGND_c_470_n 0.0146213f $X=1.655 $Y=0.445 $X2=0
+ $Y2=0
cc_229 N_A_243_409#_c_285_n N_VGND_c_470_n 0.00345258f $X=2.39 $Y=0.59 $X2=0
+ $Y2=0
cc_230 N_A_243_409#_c_276_n N_VGND_c_472_n 0.0103533f $X=2.955 $Y=0.735 $X2=0
+ $Y2=0
cc_231 N_A_243_409#_c_278_n N_VGND_c_472_n 0.0012347f $X=3.15 $Y=0.885 $X2=0
+ $Y2=0
cc_232 N_A_243_409#_M1004_d N_VGND_c_473_n 0.00227255f $X=1.515 $Y=0.235 $X2=0
+ $Y2=0
cc_233 N_A_243_409#_c_276_n N_VGND_c_473_n 0.0119912f $X=2.955 $Y=0.735 $X2=0
+ $Y2=0
cc_234 N_A_243_409#_c_278_n N_VGND_c_473_n 0.00163161f $X=3.15 $Y=0.885 $X2=0
+ $Y2=0
cc_235 N_A_243_409#_c_280_n N_VGND_c_473_n 0.014696f $X=2.305 $Y=0.59 $X2=0
+ $Y2=0
cc_236 N_A_243_409#_c_281_n N_VGND_c_473_n 0.00899998f $X=2.965 $Y=0.86 $X2=0
+ $Y2=0
cc_237 N_A_243_409#_c_349_p N_VGND_c_473_n 0.0148337f $X=3.17 $Y=0.945 $X2=0
+ $Y2=0
cc_238 N_A_243_409#_c_284_n N_VGND_c_473_n 0.0120479f $X=1.655 $Y=0.445 $X2=0
+ $Y2=0
cc_239 N_A_243_409#_c_285_n N_VGND_c_473_n 0.00493958f $X=2.39 $Y=0.59 $X2=0
+ $Y2=0
cc_240 N_A_243_409#_c_280_n A_389_47# 0.00529815f $X=2.305 $Y=0.59 $X2=-0.19
+ $Y2=-0.245
cc_241 N_A_243_409#_c_285_n A_389_47# 3.8464e-19 $X=2.39 $Y=0.59 $X2=-0.19
+ $Y2=-0.245
cc_242 N_VPWR_c_380_n N_A_137_409#_c_416_n 0.0119061f $X=0.295 $Y=2.19 $X2=0
+ $Y2=0
cc_243 N_VPWR_c_382_n N_A_137_409#_c_416_n 0.0220769f $X=2.555 $Y=3.33 $X2=0
+ $Y2=0
cc_244 N_VPWR_c_378_n N_A_137_409#_c_416_n 0.0125384f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_245 N_VPWR_c_380_n N_A_137_409#_c_419_n 0.0553152f $X=0.295 $Y=2.19 $X2=0
+ $Y2=0
cc_246 N_VPWR_c_381_n N_A_137_409#_c_417_n 0.0119061f $X=2.72 $Y=2.49 $X2=0
+ $Y2=0
cc_247 N_VPWR_c_382_n N_A_137_409#_c_417_n 0.0834959f $X=2.555 $Y=3.33 $X2=0
+ $Y2=0
cc_248 N_VPWR_c_378_n N_A_137_409#_c_417_n 0.0491523f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_249 N_VPWR_c_381_n N_A_137_409#_c_426_n 0.0375247f $X=2.72 $Y=2.49 $X2=0
+ $Y2=0
cc_250 N_VPWR_c_381_n X 0.0285424f $X=2.72 $Y=2.49 $X2=0 $Y2=0
cc_251 N_VPWR_c_383_n X 0.0274261f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_252 N_VPWR_c_378_n X 0.0156763f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_253 N_X_c_445_n N_VGND_c_469_n 0.0102369f $X=3.56 $Y=0.43 $X2=0 $Y2=0
cc_254 N_X_c_445_n N_VGND_c_472_n 0.0194268f $X=3.56 $Y=0.43 $X2=0 $Y2=0
cc_255 N_X_M1003_d N_VGND_c_473_n 0.0023218f $X=3.42 $Y=0.235 $X2=0 $Y2=0
cc_256 N_X_c_445_n N_VGND_c_473_n 0.0123961f $X=3.56 $Y=0.43 $X2=0 $Y2=0
cc_257 N_VGND_c_473_n A_225_47# 0.00357568f $X=3.6 $Y=0 $X2=-0.19 $Y2=-0.245
cc_258 N_VGND_c_473_n A_389_47# 0.00414659f $X=3.6 $Y=0 $X2=-0.19 $Y2=-0.245
cc_259 N_VGND_c_473_n A_606_47# 0.00328451f $X=3.6 $Y=0 $X2=-0.19 $Y2=-0.245
