* NGSPICE file created from sky130_fd_sc_lp__inv_lp.ext - technology: sky130A

.subckt sky130_fd_sc_lp__inv_lp A VGND VNB VPB VPWR Y
M1000 a_124_67# A VGND VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=1.197e+11p ps=1.41e+06u
M1001 Y A VPWR VPB phighvt w=1e+06u l=250000u
+  ad=2.85e+11p pd=2.57e+06u as=2.85e+11p ps=2.57e+06u
M1002 Y A a_124_67# VNB nshort w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=0p ps=0u
.ends

