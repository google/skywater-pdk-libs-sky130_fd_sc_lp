* File: sky130_fd_sc_lp__nand3_0.pex.spice
* Created: Fri Aug 28 10:48:47 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__NAND3_0%C 2 5 9 13 15 18 20 21 22 23 29
r36 22 23 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.22 $Y=1.665
+ $X2=0.22 $Y2=2.035
r37 21 22 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.22 $Y=1.295
+ $X2=0.22 $Y2=1.665
r38 20 21 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.22 $Y=0.925
+ $X2=0.22 $Y2=1.295
r39 20 29 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.27
+ $Y=1.005 $X2=0.27 $Y2=1.005
r40 16 18 71.7872 $w=1.5e-07 $l=1.4e-07 $layer=POLY_cond $X=0.36 $Y=1.845
+ $X2=0.5 $Y2=1.845
r41 14 29 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.27 $Y=1.345
+ $X2=0.27 $Y2=1.005
r42 14 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.27 $Y=1.345
+ $X2=0.27 $Y2=1.51
r43 13 29 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=0.27 $Y=0.99
+ $X2=0.27 $Y2=1.005
r44 12 13 43.5886 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=0.345 $Y=0.84
+ $X2=0.345 $Y2=0.99
r45 9 12 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.51 $Y=0.445
+ $X2=0.51 $Y2=0.84
r46 3 18 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.5 $Y=1.92 $X2=0.5
+ $Y2=1.845
r47 3 5 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=0.5 $Y=1.92 $X2=0.5
+ $Y2=2.63
r48 2 16 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.36 $Y=1.77 $X2=0.36
+ $Y2=1.845
r49 2 15 133.319 $w=1.5e-07 $l=2.6e-07 $layer=POLY_cond $X=0.36 $Y=1.77 $X2=0.36
+ $Y2=1.51
.ends

.subckt PM_SKY130_FD_SC_LP__NAND3_0%B 3 7 9 10 11 16
c39 16 0 6.20581e-20 $X=0.84 $Y=1.365
c40 9 0 1.99346e-19 $X=0.72 $Y=0.925
r41 16 19 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.84 $Y=1.365
+ $X2=0.84 $Y2=1.53
r42 16 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.84 $Y=1.365
+ $X2=0.84 $Y2=1.2
r43 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.84
+ $Y=1.365 $X2=0.84 $Y2=1.365
r44 11 17 9.73895 $w=3.53e-07 $l=3e-07 $layer=LI1_cond $X=0.747 $Y=1.665
+ $X2=0.747 $Y2=1.365
r45 10 17 2.27242 $w=3.53e-07 $l=7e-08 $layer=LI1_cond $X=0.747 $Y=1.295
+ $X2=0.747 $Y2=1.365
r46 9 10 12.0114 $w=3.53e-07 $l=3.7e-07 $layer=LI1_cond $X=0.747 $Y=0.925
+ $X2=0.747 $Y2=1.295
r47 7 19 564.043 $w=1.5e-07 $l=1.1e-06 $layer=POLY_cond $X=0.93 $Y=2.63 $X2=0.93
+ $Y2=1.53
r48 3 18 387.138 $w=1.5e-07 $l=7.55e-07 $layer=POLY_cond $X=0.9 $Y=0.445 $X2=0.9
+ $Y2=1.2
.ends

.subckt PM_SKY130_FD_SC_LP__NAND3_0%A 3 7 11 12 13 14 15 20
c35 7 0 1.99346e-19 $X=1.36 $Y=2.63
r36 20 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.38
+ $Y=1.005 $X2=1.38 $Y2=1.005
r37 14 15 11.2212 $w=3.78e-07 $l=3.7e-07 $layer=LI1_cond $X=1.285 $Y=1.295
+ $X2=1.285 $Y2=1.665
r38 14 21 8.79496 $w=3.78e-07 $l=2.9e-07 $layer=LI1_cond $X=1.285 $Y=1.295
+ $X2=1.285 $Y2=1.005
r39 13 21 2.4262 $w=3.78e-07 $l=8e-08 $layer=LI1_cond $X=1.285 $Y=0.925
+ $X2=1.285 $Y2=1.005
r40 11 20 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.38 $Y=1.345
+ $X2=1.38 $Y2=1.005
r41 11 12 38.6168 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.38 $Y=1.345
+ $X2=1.38 $Y2=1.51
r42 10 20 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.38 $Y=0.84
+ $X2=1.38 $Y2=1.005
r43 7 12 574.298 $w=1.5e-07 $l=1.12e-06 $layer=POLY_cond $X=1.36 $Y=2.63
+ $X2=1.36 $Y2=1.51
r44 3 10 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=1.29 $Y=0.445
+ $X2=1.29 $Y2=0.84
.ends

.subckt PM_SKY130_FD_SC_LP__NAND3_0%VPWR 1 2 7 9 13 16 17 18 25 26
r27 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r28 25 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r29 23 30 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r30 22 23 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r31 20 29 4.40602 $w=1.7e-07 $l=2.08e-07 $layer=LI1_cond $X=0.415 $Y=3.33
+ $X2=0.207 $Y2=3.33
r32 20 22 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.415 $Y=3.33
+ $X2=0.72 $Y2=3.33
r33 18 26 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=0.96 $Y=3.33
+ $X2=1.68 $Y2=3.33
r34 18 23 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=0.96 $Y=3.33
+ $X2=0.72 $Y2=3.33
r35 16 22 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=1.01 $Y=3.33
+ $X2=0.72 $Y2=3.33
r36 16 17 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.01 $Y=3.33 $X2=1.14
+ $Y2=3.33
r37 15 25 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=1.27 $Y=3.33
+ $X2=1.68 $Y2=3.33
r38 15 17 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.27 $Y=3.33 $X2=1.14
+ $Y2=3.33
r39 11 17 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=1.14 $Y=3.245
+ $X2=1.14 $Y2=3.33
r40 11 13 35.0165 $w=2.58e-07 $l=7.9e-07 $layer=LI1_cond $X=1.14 $Y=3.245
+ $X2=1.14 $Y2=2.455
r41 7 29 3.0715 $w=2.95e-07 $l=1.11018e-07 $layer=LI1_cond $X=0.267 $Y=3.245
+ $X2=0.207 $Y2=3.33
r42 7 9 30.862 $w=2.93e-07 $l=7.9e-07 $layer=LI1_cond $X=0.267 $Y=3.245
+ $X2=0.267 $Y2=2.455
r43 2 13 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=1.005
+ $Y=2.31 $X2=1.145 $Y2=2.455
r44 1 9 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.16
+ $Y=2.31 $X2=0.285 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_LP__NAND3_0%Y 1 2 3 11 15 17 18 19 25 31 36
c41 25 0 6.20581e-20 $X=1.44 $Y=2.02
r42 19 25 2.74102 $w=2e-07 $l=1.97e-07 $layer=LI1_cond $X=1.637 $Y=2.02 $X2=1.44
+ $Y2=2.02
r43 19 36 8.18787 $w=5.63e-07 $l=3.35e-07 $layer=LI1_cond $X=1.637 $Y=2.12
+ $X2=1.637 $Y2=2.455
r44 18 25 13.3091 $w=1.98e-07 $l=2.4e-07 $layer=LI1_cond $X=1.2 $Y=2.02 $X2=1.44
+ $Y2=2.02
r45 18 26 19.9636 $w=1.98e-07 $l=3.6e-07 $layer=LI1_cond $X=1.2 $Y=2.02 $X2=0.84
+ $Y2=2.02
r46 17 26 3.89998 $w=2e-07 $l=1.28e-07 $layer=LI1_cond $X=0.712 $Y=2.02 $X2=0.84
+ $Y2=2.02
r47 17 31 10.9136 $w=4.23e-07 $l=3.35e-07 $layer=LI1_cond $X=0.712 $Y=2.12
+ $X2=0.712 $Y2=2.455
r48 13 15 8.20679 $w=3.28e-07 $l=2.35e-07 $layer=LI1_cond $X=1.505 $Y=0.445
+ $X2=1.74 $Y2=0.445
r49 11 19 3.7255 $w=2.92e-07 $l=1.44599e-07 $layer=LI1_cond $X=1.74 $Y=1.92
+ $X2=1.637 $Y2=2.02
r50 10 15 3.96751 $w=1.9e-07 $l=1.65e-07 $layer=LI1_cond $X=1.74 $Y=0.61
+ $X2=1.74 $Y2=0.445
r51 10 11 76.4689 $w=1.88e-07 $l=1.31e-06 $layer=LI1_cond $X=1.74 $Y=0.61
+ $X2=1.74 $Y2=1.92
r52 3 36 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=1.435
+ $Y=2.31 $X2=1.575 $Y2=2.455
r53 2 31 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=0.575
+ $Y=2.31 $X2=0.715 $Y2=2.455
r54 1 13 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.365
+ $Y=0.235 $X2=1.505 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__NAND3_0%VGND 1 4 6 8 15 16
r22 19 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r23 15 16 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r24 13 20 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r25 12 15 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r26 12 13 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r27 10 19 4.70058 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=0.46 $Y=0 $X2=0.23
+ $Y2=0
r28 10 12 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=0.46 $Y=0 $X2=0.72
+ $Y2=0
r29 8 16 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=0.96 $Y=0 $X2=1.68
+ $Y2=0
r30 8 13 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=0.96 $Y=0 $X2=0.72
+ $Y2=0
r31 4 19 3.0656 $w=3.3e-07 $l=1.12916e-07 $layer=LI1_cond $X=0.295 $Y=0.085
+ $X2=0.23 $Y2=0
r32 4 6 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=0.295 $Y=0.085
+ $X2=0.295 $Y2=0.445
r33 1 6 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.17
+ $Y=0.235 $X2=0.295 $Y2=0.445
.ends

