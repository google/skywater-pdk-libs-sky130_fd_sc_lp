# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__dlxbn_1
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__dlxbn_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.160000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.455000 1.205000 0.900000 1.875000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.556500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.805000 0.255000 8.065000 3.075000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.556500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.590000 1.805000 7.125000 3.075000 ;
        RECT 6.785000 0.995000 7.125000 1.805000 ;
    END
  END Q_N
  PIN GATE_N
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 1.060000 0.255000 1.775000 0.675000 ;
    END
  END GATE_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 8.160000 0.085000 ;
        RECT 0.675000  0.085000 0.890000 1.035000 ;
        RECT 2.315000  0.085000 2.645000 0.505000 ;
        RECT 4.290000  0.085000 4.600000 1.095000 ;
        RECT 6.065000  0.085000 6.275000 0.905000 ;
        RECT 7.305000  0.085000 7.635000 0.485000 ;
      LAYER mcon ;
        RECT 0.155000 -0.085000 0.325000 0.085000 ;
        RECT 0.635000 -0.085000 0.805000 0.085000 ;
        RECT 1.115000 -0.085000 1.285000 0.085000 ;
        RECT 1.595000 -0.085000 1.765000 0.085000 ;
        RECT 2.075000 -0.085000 2.245000 0.085000 ;
        RECT 2.555000 -0.085000 2.725000 0.085000 ;
        RECT 3.035000 -0.085000 3.205000 0.085000 ;
        RECT 3.515000 -0.085000 3.685000 0.085000 ;
        RECT 3.995000 -0.085000 4.165000 0.085000 ;
        RECT 4.475000 -0.085000 4.645000 0.085000 ;
        RECT 4.955000 -0.085000 5.125000 0.085000 ;
        RECT 5.435000 -0.085000 5.605000 0.085000 ;
        RECT 5.915000 -0.085000 6.085000 0.085000 ;
        RECT 6.395000 -0.085000 6.565000 0.085000 ;
        RECT 6.875000 -0.085000 7.045000 0.085000 ;
        RECT 7.355000 -0.085000 7.525000 0.085000 ;
        RECT 7.835000 -0.085000 8.005000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 8.160000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.245000 8.160000 3.415000 ;
        RECT 0.640000 2.455000 0.970000 3.245000 ;
        RECT 2.350000 2.825000 2.680000 3.245000 ;
        RECT 4.155000 2.425000 4.755000 3.245000 ;
        RECT 6.090000 1.805000 6.350000 3.245000 ;
        RECT 7.305000 1.815000 7.635000 3.245000 ;
      LAYER mcon ;
        RECT 0.155000 3.245000 0.325000 3.415000 ;
        RECT 0.635000 3.245000 0.805000 3.415000 ;
        RECT 1.115000 3.245000 1.285000 3.415000 ;
        RECT 1.595000 3.245000 1.765000 3.415000 ;
        RECT 2.075000 3.245000 2.245000 3.415000 ;
        RECT 2.555000 3.245000 2.725000 3.415000 ;
        RECT 3.035000 3.245000 3.205000 3.415000 ;
        RECT 3.515000 3.245000 3.685000 3.415000 ;
        RECT 3.995000 3.245000 4.165000 3.415000 ;
        RECT 4.475000 3.245000 4.645000 3.415000 ;
        RECT 4.955000 3.245000 5.125000 3.415000 ;
        RECT 5.435000 3.245000 5.605000 3.415000 ;
        RECT 5.915000 3.245000 6.085000 3.415000 ;
        RECT 6.395000 3.245000 6.565000 3.415000 ;
        RECT 6.875000 3.245000 7.045000 3.415000 ;
        RECT 7.355000 3.245000 7.525000 3.415000 ;
        RECT 7.835000 3.245000 8.005000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 8.160000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.105000 0.695000 0.505000 1.035000 ;
      RECT 0.105000 1.035000 0.275000 2.045000 ;
      RECT 0.105000 2.045000 0.460000 2.115000 ;
      RECT 0.105000 2.115000 2.770000 2.285000 ;
      RECT 0.105000 2.285000 0.460000 2.695000 ;
      RECT 1.070000 0.845000 1.515000 1.195000 ;
      RECT 1.070000 1.195000 3.240000 1.365000 ;
      RECT 1.070000 1.365000 2.200000 1.945000 ;
      RECT 1.775000 2.455000 3.145000 2.635000 ;
      RECT 1.775000 2.635000 2.105000 3.075000 ;
      RECT 1.945000 0.285000 2.135000 0.675000 ;
      RECT 1.945000 0.675000 3.780000 0.845000 ;
      RECT 2.440000 1.585000 2.770000 2.115000 ;
      RECT 2.975000 1.925000 3.580000 2.225000 ;
      RECT 2.975000 2.225000 3.145000 2.455000 ;
      RECT 2.980000 1.015000 3.240000 1.195000 ;
      RECT 2.980000 1.365000 3.240000 1.685000 ;
      RECT 3.165000 0.275000 4.120000 0.485000 ;
      RECT 3.315000 2.395000 3.930000 2.565000 ;
      RECT 3.315000 2.565000 3.730000 3.065000 ;
      RECT 3.410000 0.845000 3.780000 1.095000 ;
      RECT 3.410000 1.095000 3.580000 1.925000 ;
      RECT 3.760000 1.575000 4.120000 1.745000 ;
      RECT 3.760000 1.745000 3.930000 2.395000 ;
      RECT 3.950000 0.485000 4.120000 1.275000 ;
      RECT 3.950000 1.275000 4.845000 1.445000 ;
      RECT 3.950000 1.445000 4.120000 1.575000 ;
      RECT 4.100000 1.925000 5.240000 2.255000 ;
      RECT 4.585000 1.445000 4.845000 1.605000 ;
      RECT 4.770000 0.255000 5.895000 0.675000 ;
      RECT 4.770000 0.675000 5.195000 1.095000 ;
      RECT 4.925000 2.255000 5.240000 3.075000 ;
      RECT 5.015000 1.095000 5.195000 1.925000 ;
      RECT 5.365000 0.855000 5.555000 1.415000 ;
      RECT 5.365000 1.415000 6.615000 1.585000 ;
      RECT 5.590000 1.585000 6.615000 1.635000 ;
      RECT 5.590000 1.635000 5.920000 2.485000 ;
      RECT 5.725000 0.675000 5.895000 1.075000 ;
      RECT 5.725000 1.075000 6.615000 1.245000 ;
      RECT 6.445000 0.655000 7.625000 0.825000 ;
      RECT 6.445000 0.825000 6.615000 1.075000 ;
      RECT 7.295000 0.825000 7.625000 1.515000 ;
  END
END sky130_fd_sc_lp__dlxbn_1
