* File: sky130_fd_sc_lp__nor3_m.pxi.spice
* Created: Fri Aug 28 10:56:01 2020
* 
x_PM_SKY130_FD_SC_LP__NOR3_M%A N_A_c_47_n N_A_M1002_g N_A_c_54_n N_A_M1000_g
+ N_A_c_48_n N_A_c_49_n N_A_c_50_n N_A_c_55_n A A A A N_A_c_52_n
+ PM_SKY130_FD_SC_LP__NOR3_M%A
x_PM_SKY130_FD_SC_LP__NOR3_M%B N_B_M1001_g N_B_M1003_g N_B_c_85_n N_B_c_90_n B B
+ B B B N_B_c_87_n PM_SKY130_FD_SC_LP__NOR3_M%B
x_PM_SKY130_FD_SC_LP__NOR3_M%C N_C_M1005_g N_C_M1004_g N_C_c_129_n N_C_c_134_n C
+ C C N_C_c_131_n PM_SKY130_FD_SC_LP__NOR3_M%C
x_PM_SKY130_FD_SC_LP__NOR3_M%VPWR N_VPWR_M1000_s N_VPWR_c_163_n N_VPWR_c_164_n
+ VPWR N_VPWR_c_165_n N_VPWR_c_162_n PM_SKY130_FD_SC_LP__NOR3_M%VPWR
x_PM_SKY130_FD_SC_LP__NOR3_M%Y N_Y_M1002_d N_Y_M1004_d N_Y_M1005_d N_Y_c_182_n
+ N_Y_c_183_n N_Y_c_184_n N_Y_c_189_n N_Y_c_185_n Y N_Y_c_187_n
+ PM_SKY130_FD_SC_LP__NOR3_M%Y
x_PM_SKY130_FD_SC_LP__NOR3_M%VGND N_VGND_M1002_s N_VGND_M1001_d N_VGND_c_220_n
+ N_VGND_c_221_n N_VGND_c_222_n N_VGND_c_223_n N_VGND_c_224_n VGND
+ N_VGND_c_225_n N_VGND_c_226_n PM_SKY130_FD_SC_LP__NOR3_M%VGND
cc_1 VNB N_A_c_47_n 0.00799575f $X=-0.19 $Y=-0.245 $X2=0.36 $Y2=2.155
cc_2 VNB N_A_c_48_n 0.0213365f $X=-0.19 $Y=-0.245 $X2=0.34 $Y2=0.855
cc_3 VNB N_A_c_49_n 0.0363598f $X=-0.19 $Y=-0.245 $X2=0.34 $Y2=1.005
cc_4 VNB N_A_c_50_n 0.0236201f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.525
cc_5 VNB A 0.00732696f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_6 VNB N_A_c_52_n 0.0381798f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.02
cc_7 VNB N_B_M1001_g 0.0373822f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=0.855
cc_8 VNB N_B_c_85_n 0.0154125f $X=-0.19 $Y=-0.245 $X2=0.34 $Y2=1.005
cc_9 VNB B 0.00540434f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.525
cc_10 VNB N_B_c_87_n 0.0155602f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_C_M1004_g 0.0414246f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=2.625
cc_12 VNB N_C_c_129_n 0.0191305f $X=-0.19 $Y=-0.245 $X2=0.34 $Y2=1.005
cc_13 VNB C 0.00470398f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.525
cc_14 VNB N_C_c_131_n 0.0161667f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_15 VNB N_VPWR_c_162_n 0.0840719f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=2.23
cc_16 VNB N_Y_c_182_n 0.0100202f $X=-0.19 $Y=-0.245 $X2=0.34 $Y2=0.855
cc_17 VNB N_Y_c_183_n 0.0190501f $X=-0.19 $Y=-0.245 $X2=0.36 $Y2=2.23
cc_18 VNB N_Y_c_184_n 0.0307399f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_Y_c_185_n 0.0130139f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB Y 0.00389508f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_Y_c_187_n 0.00187043f $X=-0.19 $Y=-0.245 $X2=0.255 $Y2=0.925
cc_22 VNB N_VGND_c_220_n 0.0119573f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=2.625
cc_23 VNB N_VGND_c_221_n 0.00881971f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.005
cc_24 VNB N_VGND_c_222_n 0.00673153f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.525
cc_25 VNB N_VGND_c_223_n 0.0192456f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=2.23
cc_26 VNB N_VGND_c_224_n 0.00401463f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_225_n 0.0211964f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_226_n 0.138211f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.02
cc_29 VPB N_A_c_47_n 0.0330096f $X=-0.19 $Y=1.655 $X2=0.36 $Y2=2.155
cc_30 VPB N_A_c_54_n 0.0198492f $X=-0.19 $Y=1.655 $X2=0.54 $Y2=2.305
cc_31 VPB N_A_c_55_n 0.0317071f $X=-0.19 $Y=1.655 $X2=0.54 $Y2=2.23
cc_32 VPB A 0.0186508f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_33 VPB N_B_M1003_g 0.0346988f $X=-0.19 $Y=1.655 $X2=0.54 $Y2=2.625
cc_34 VPB N_B_c_85_n 0.0059376f $X=-0.19 $Y=1.655 $X2=0.34 $Y2=1.005
cc_35 VPB N_B_c_90_n 0.0156026f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.36
cc_36 VPB B 0.00915083f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.525
cc_37 VPB N_C_M1005_g 0.0446125f $X=-0.19 $Y=1.655 $X2=0.5 $Y2=0.855
cc_38 VPB N_C_c_129_n 0.00404552f $X=-0.19 $Y=1.655 $X2=0.34 $Y2=1.005
cc_39 VPB N_C_c_134_n 0.0168323f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.36
cc_40 VPB C 0.0121972f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.525
cc_41 VPB N_VPWR_c_163_n 0.0121156f $X=-0.19 $Y=1.655 $X2=0.5 $Y2=0.535
cc_42 VPB N_VPWR_c_164_n 0.0239699f $X=-0.19 $Y=1.655 $X2=0.54 $Y2=2.305
cc_43 VPB N_VPWR_c_165_n 0.0465858f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_44 VPB N_VPWR_c_162_n 0.0758722f $X=-0.19 $Y=1.655 $X2=0.54 $Y2=2.23
cc_45 VPB N_Y_c_184_n 0.0361723f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_46 VPB N_Y_c_189_n 0.0300079f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.95
cc_47 N_A_c_48_n N_B_M1001_g 0.0195444f $X=0.34 $Y=0.855 $X2=0 $Y2=0
cc_48 A N_B_M1001_g 0.00112841f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_49 N_A_c_52_n N_B_M1001_g 0.00734446f $X=0.27 $Y=1.02 $X2=0 $Y2=0
cc_50 N_A_c_47_n N_B_M1003_g 0.00547445f $X=0.36 $Y=2.155 $X2=0 $Y2=0
cc_51 N_A_c_55_n N_B_M1003_g 0.0405766f $X=0.54 $Y=2.23 $X2=0 $Y2=0
cc_52 N_A_c_50_n N_B_c_85_n 0.0114238f $X=0.27 $Y=1.525 $X2=0 $Y2=0
cc_53 N_A_c_47_n N_B_c_90_n 0.0114238f $X=0.36 $Y=2.155 $X2=0 $Y2=0
cc_54 N_A_c_55_n B 0.00882625f $X=0.54 $Y=2.23 $X2=0 $Y2=0
cc_55 A B 0.0474145f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_56 N_A_c_52_n B 0.00725628f $X=0.27 $Y=1.02 $X2=0 $Y2=0
cc_57 A N_B_c_87_n 7.14411e-19 $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_58 N_A_c_52_n N_B_c_87_n 0.0114238f $X=0.27 $Y=1.02 $X2=0 $Y2=0
cc_59 N_A_c_54_n N_VPWR_c_164_n 0.0070913f $X=0.54 $Y=2.305 $X2=0 $Y2=0
cc_60 N_A_c_55_n N_VPWR_c_164_n 0.00427524f $X=0.54 $Y=2.23 $X2=0 $Y2=0
cc_61 A N_VPWR_c_164_n 0.0106281f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_62 N_A_c_54_n N_VPWR_c_165_n 0.00490845f $X=0.54 $Y=2.305 $X2=0 $Y2=0
cc_63 N_A_c_54_n N_VPWR_c_162_n 0.00506877f $X=0.54 $Y=2.305 $X2=0 $Y2=0
cc_64 N_A_c_48_n Y 0.00187595f $X=0.34 $Y=0.855 $X2=0 $Y2=0
cc_65 A Y 0.0102802f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_66 N_A_c_48_n N_Y_c_187_n 0.00237894f $X=0.34 $Y=0.855 $X2=0 $Y2=0
cc_67 N_A_c_48_n N_VGND_c_221_n 0.00355982f $X=0.34 $Y=0.855 $X2=0 $Y2=0
cc_68 N_A_c_49_n N_VGND_c_221_n 0.00239837f $X=0.34 $Y=1.005 $X2=0 $Y2=0
cc_69 A N_VGND_c_221_n 0.0133587f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_70 N_A_c_48_n N_VGND_c_223_n 0.00499542f $X=0.34 $Y=0.855 $X2=0 $Y2=0
cc_71 N_A_c_48_n N_VGND_c_226_n 0.0101395f $X=0.34 $Y=0.855 $X2=0 $Y2=0
cc_72 N_A_c_49_n N_VGND_c_226_n 0.00219168f $X=0.34 $Y=1.005 $X2=0 $Y2=0
cc_73 A N_VGND_c_226_n 0.00167711f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_74 N_B_c_90_n N_C_M1005_g 0.0545157f $X=0.84 $Y=1.915 $X2=0 $Y2=0
cc_75 B N_C_M1005_g 0.0032103f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_76 N_B_M1001_g N_C_M1004_g 0.0297377f $X=0.93 $Y=0.535 $X2=0 $Y2=0
cc_77 N_B_c_87_n N_C_c_129_n 0.0137631f $X=0.84 $Y=1.41 $X2=0 $Y2=0
cc_78 N_B_c_85_n N_C_c_134_n 0.0137631f $X=0.84 $Y=1.75 $X2=0 $Y2=0
cc_79 N_B_M1001_g C 0.00605045f $X=0.93 $Y=0.535 $X2=0 $Y2=0
cc_80 B C 0.065811f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_81 N_B_M1001_g N_C_c_131_n 0.0137631f $X=0.93 $Y=0.535 $X2=0 $Y2=0
cc_82 B N_C_c_131_n 6.12778e-19 $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_83 B N_VPWR_c_164_n 0.0143303f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_84 N_B_M1003_g N_VPWR_c_165_n 0.00431881f $X=0.93 $Y=2.625 $X2=0 $Y2=0
cc_85 B N_VPWR_c_165_n 0.00845743f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_86 N_B_M1003_g N_VPWR_c_162_n 0.00506877f $X=0.93 $Y=2.625 $X2=0 $Y2=0
cc_87 B N_VPWR_c_162_n 0.009768f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_88 N_B_M1001_g N_Y_c_182_n 0.0139794f $X=0.93 $Y=0.535 $X2=0 $Y2=0
cc_89 B N_Y_c_182_n 0.00721302f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_90 N_B_c_87_n N_Y_c_182_n 2.13288e-19 $X=0.84 $Y=1.41 $X2=0 $Y2=0
cc_91 B N_Y_c_189_n 0.00730376f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_92 B Y 0.0151683f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_93 N_B_c_87_n Y 9.98363e-19 $X=0.84 $Y=1.41 $X2=0 $Y2=0
cc_94 N_B_M1001_g N_Y_c_187_n 0.00129206f $X=0.93 $Y=0.535 $X2=0 $Y2=0
cc_95 N_B_M1001_g N_VGND_c_222_n 0.00168203f $X=0.93 $Y=0.535 $X2=0 $Y2=0
cc_96 N_B_M1001_g N_VGND_c_223_n 0.00499542f $X=0.93 $Y=0.535 $X2=0 $Y2=0
cc_97 N_B_M1001_g N_VGND_c_226_n 0.00533443f $X=0.93 $Y=0.535 $X2=0 $Y2=0
cc_98 N_C_M1005_g N_VPWR_c_165_n 0.00490845f $X=1.32 $Y=2.625 $X2=0 $Y2=0
cc_99 N_C_M1005_g N_VPWR_c_162_n 0.00506877f $X=1.32 $Y=2.625 $X2=0 $Y2=0
cc_100 N_C_M1004_g N_Y_c_182_n 0.0135724f $X=1.36 $Y=0.535 $X2=0 $Y2=0
cc_101 C N_Y_c_182_n 0.0244746f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_102 N_C_c_131_n N_Y_c_182_n 8.8805e-19 $X=1.38 $Y=1.375 $X2=0 $Y2=0
cc_103 N_C_M1004_g N_Y_c_183_n 0.00284132f $X=1.36 $Y=0.535 $X2=0 $Y2=0
cc_104 N_C_M1005_g N_Y_c_184_n 0.0100508f $X=1.32 $Y=2.625 $X2=0 $Y2=0
cc_105 N_C_M1004_g N_Y_c_184_n 0.00652586f $X=1.36 $Y=0.535 $X2=0 $Y2=0
cc_106 C N_Y_c_184_n 0.0667321f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_107 N_C_c_131_n N_Y_c_184_n 0.0163648f $X=1.38 $Y=1.375 $X2=0 $Y2=0
cc_108 N_C_M1005_g N_Y_c_189_n 0.00136961f $X=1.32 $Y=2.625 $X2=0 $Y2=0
cc_109 N_C_c_134_n N_Y_c_189_n 0.00271709f $X=1.38 $Y=1.88 $X2=0 $Y2=0
cc_110 C N_Y_c_189_n 0.00219841f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_111 N_C_c_131_n N_Y_c_185_n 0.00339815f $X=1.38 $Y=1.375 $X2=0 $Y2=0
cc_112 N_C_M1004_g N_VGND_c_222_n 0.00309744f $X=1.36 $Y=0.535 $X2=0 $Y2=0
cc_113 N_C_M1004_g N_VGND_c_225_n 0.00499542f $X=1.36 $Y=0.535 $X2=0 $Y2=0
cc_114 N_C_M1004_g N_VGND_c_226_n 0.0057107f $X=1.36 $Y=0.535 $X2=0 $Y2=0
cc_115 N_VPWR_c_165_n N_Y_c_189_n 0.0107098f $X=1.68 $Y=3.33 $X2=0 $Y2=0
cc_116 N_VPWR_c_162_n N_Y_c_189_n 0.0127831f $X=1.68 $Y=3.33 $X2=0 $Y2=0
cc_117 N_Y_c_182_n N_VGND_c_222_n 0.0128647f $X=1.47 $Y=0.925 $X2=0 $Y2=0
cc_118 N_Y_c_187_n N_VGND_c_223_n 0.00599271f $X=0.715 $Y=0.6 $X2=0 $Y2=0
cc_119 N_Y_c_183_n N_VGND_c_225_n 0.0107695f $X=1.575 $Y=0.6 $X2=0 $Y2=0
cc_120 N_Y_c_182_n N_VGND_c_226_n 0.0138164f $X=1.47 $Y=0.925 $X2=0 $Y2=0
cc_121 N_Y_c_183_n N_VGND_c_226_n 0.01196f $X=1.575 $Y=0.6 $X2=0 $Y2=0
cc_122 N_Y_c_187_n N_VGND_c_226_n 0.00722947f $X=0.715 $Y=0.6 $X2=0 $Y2=0
