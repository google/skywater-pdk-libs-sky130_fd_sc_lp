* NGSPICE file created from sky130_fd_sc_lp__or4_m.ext - technology: sky130A

.subckt sky130_fd_sc_lp__or4_m A B C D VGND VNB VPB VPWR X
M1000 VPWR A a_343_397# VPB phighvt w=420000u l=150000u
+  ad=2.499e+11p pd=2.03e+06u as=8.82e+10p ps=1.26e+06u
M1001 a_116_397# B VGND VNB nshort w=420000u l=150000u
+  ad=2.352e+11p pd=2.8e+06u as=5.817e+11p ps=5.29e+06u
M1002 a_271_397# C a_199_397# VPB phighvt w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=8.82e+10p ps=1.26e+06u
M1003 a_199_397# D a_116_397# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1004 X a_116_397# VGND VNB nshort w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1005 a_343_397# B a_271_397# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_116_397# D VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND A a_116_397# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 X a_116_397# VPWR VPB phighvt w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1009 VGND C a_116_397# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

