* NGSPICE file created from sky130_fd_sc_lp__dfstp_1.ext - technology: sky130A

.subckt sky130_fd_sc_lp__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
M1000 Q a_1832_131# VGND VNB nshort w=840000u l=150000u
+  ad=2.226e+11p pd=2.21e+06u as=1.2149e+12p ps=1.126e+07u
M1001 a_486_119# a_202_463# a_400_119# VPB phighvt w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=1.176e+11p ps=1.4e+06u
M1002 VPWR a_1329_65# a_1092_417# VPB phighvt w=420000u l=150000u
+  ad=1.4619e+12p pd=1.374e+07u as=2.226e+11p ps=2.74e+06u
M1003 a_614_93# a_486_119# VPWR VPB phighvt w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=0p ps=0u
M1004 a_985_379# a_33_463# a_1175_417# VPB phighvt w=840000u l=150000u
+  ad=5.625e+11p pd=4.91e+06u as=3.801e+11p ps=3.8e+06u
M1005 a_400_119# D VGND VNB nshort w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=0p ps=0u
M1006 Q a_1832_131# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=3.339e+11p pd=3.05e+06u as=0p ps=0u
M1007 a_985_379# a_486_119# VPWR VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND SET_B a_1359_91# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1009 a_400_119# D VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_1329_65# a_1175_417# VPWR VPB phighvt w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1011 VGND a_1175_417# a_1832_131# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1012 VPWR CLK a_33_463# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.696e+11p ps=1.81e+06u
M1013 a_1175_417# a_202_463# a_1092_417# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_1287_91# a_33_463# a_1175_417# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=2.158e+11p ps=2.03e+06u
M1015 a_1359_91# a_1329_65# a_1287_91# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VGND SET_B a_853_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1017 VGND CLK a_33_463# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1018 a_202_463# a_33_463# VGND VNB nshort w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1019 a_1329_65# a_1175_417# VGND VNB nshort w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=0p ps=0u
M1020 a_582_463# a_33_463# a_486_119# VPB phighvt w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1021 a_1175_417# SET_B VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VGND a_614_93# a_572_119# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1023 VPWR a_614_93# a_582_463# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_202_463# a_33_463# VPWR VPB phighvt w=640000u l=150000u
+  ad=1.696e+11p pd=1.81e+06u as=0p ps=0u
M1025 VPWR SET_B a_614_93# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 VPWR a_1175_417# a_1832_131# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.696e+11p ps=1.81e+06u
M1027 a_853_47# a_486_119# a_614_93# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1028 a_486_119# a_33_463# a_400_119# VNB nshort w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=0p ps=0u
M1029 a_1110_47# a_486_119# VGND VNB nshort w=640000u l=150000u
+  ad=1.344e+11p pd=1.7e+06u as=0p ps=0u
M1030 a_572_119# a_202_463# a_486_119# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_1175_417# a_202_463# a_1110_47# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

