* File: sky130_fd_sc_lp__o211a_1.pex.spice
* Created: Wed Sep  2 10:13:45 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O211A_1%A_80_237# 1 2 3 10 12 15 17 20 23 24 26 27
+ 30 32 36 38 40 42 44
c93 20 0 1.40531e-19 $X=0.925 $Y=1.35
r94 38 46 2.66522 $w=3.2e-07 $l=8.5e-08 $layer=LI1_cond $X=3.41 $Y=2.09 $X2=3.41
+ $Y2=2.005
r95 38 40 29.5314 $w=3.18e-07 $l=8.2e-07 $layer=LI1_cond $X=3.41 $Y=2.09
+ $X2=3.41 $Y2=2.91
r96 34 36 21.1281 $w=3.28e-07 $l=6.05e-07 $layer=LI1_cond $X=3.405 $Y=1.025
+ $X2=3.405 $Y2=0.42
r97 33 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.545 $Y=2.005
+ $X2=2.38 $Y2=2.005
r98 32 46 5.01689 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=3.25 $Y=2.005
+ $X2=3.41 $Y2=2.005
r99 32 33 45.9947 $w=1.68e-07 $l=7.05e-07 $layer=LI1_cond $X=3.25 $Y=2.005
+ $X2=2.545 $Y2=2.005
r100 28 44 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.38 $Y=2.09
+ $X2=2.38 $Y2=2.005
r101 28 30 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=2.38 $Y=2.09
+ $X2=2.38 $Y2=2.475
r102 26 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.215 $Y=2.005
+ $X2=2.38 $Y2=2.005
r103 26 27 58.0642 $w=1.68e-07 $l=8.9e-07 $layer=LI1_cond $X=2.215 $Y=2.005
+ $X2=1.325 $Y2=2.005
r104 25 42 4.9928 $w=2.5e-07 $l=2.1166e-07 $layer=LI1_cond $X=1.325 $Y=1.11
+ $X2=1.205 $Y2=1.27
r105 24 34 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.24 $Y=1.11
+ $X2=3.405 $Y2=1.025
r106 24 25 124.936 $w=1.68e-07 $l=1.915e-06 $layer=LI1_cond $X=3.24 $Y=1.11
+ $X2=1.325 $Y2=1.11
r107 23 27 7.07814 $w=1.7e-07 $l=1.56844e-07 $layer=LI1_cond $X=1.205 $Y=1.92
+ $X2=1.325 $Y2=2.005
r108 22 42 1.48997 $w=2.4e-07 $l=2.45e-07 $layer=LI1_cond $X=1.205 $Y=1.515
+ $X2=1.205 $Y2=1.27
r109 22 23 19.4475 $w=2.38e-07 $l=4.05e-07 $layer=LI1_cond $X=1.205 $Y=1.515
+ $X2=1.205 $Y2=1.92
r110 20 49 8.00906 $w=3.31e-07 $l=5.5e-08 $layer=POLY_cond $X=0.925 $Y=1.352
+ $X2=0.98 $Y2=1.352
r111 20 47 56.7915 $w=3.31e-07 $l=3.9e-07 $layer=POLY_cond $X=0.925 $Y=1.352
+ $X2=0.535 $Y2=1.352
r112 19 20 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.925
+ $Y=1.35 $X2=0.925 $Y2=1.35
r113 17 42 4.9928 $w=2.5e-07 $l=1.54919e-07 $layer=LI1_cond $X=1.085 $Y=1.35
+ $X2=1.205 $Y2=1.27
r114 17 19 5.5876 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=1.085 $Y=1.35
+ $X2=0.925 $Y2=1.35
r115 13 49 21.295 $w=1.5e-07 $l=1.68e-07 $layer=POLY_cond $X=0.98 $Y=1.52
+ $X2=0.98 $Y2=1.352
r116 13 15 484.564 $w=1.5e-07 $l=9.45e-07 $layer=POLY_cond $X=0.98 $Y=1.52
+ $X2=0.98 $Y2=2.465
r117 10 47 21.295 $w=1.5e-07 $l=1.67e-07 $layer=POLY_cond $X=0.535 $Y=1.185
+ $X2=0.535 $Y2=1.352
r118 10 12 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.535 $Y=1.185
+ $X2=0.535 $Y2=0.655
r119 3 46 400 $w=1.7e-07 $l=2.29565e-07 $layer=licon1_PDIFF $count=1 $X=3.265
+ $Y=1.835 $X2=3.405 $Y2=2.005
r120 3 40 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=3.265
+ $Y=1.835 $X2=3.405 $Y2=2.91
r121 2 44 600 $w=1.7e-07 $l=2.66786e-07 $layer=licon1_PDIFF $count=1 $X=2.185
+ $Y=1.835 $X2=2.38 $Y2=2.005
r122 2 30 300 $w=1.7e-07 $l=7.31027e-07 $layer=licon1_PDIFF $count=2 $X=2.185
+ $Y=1.835 $X2=2.38 $Y2=2.475
r123 1 36 91 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=2 $X=3.265
+ $Y=0.245 $X2=3.405 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__O211A_1%A1 3 7 9 12 13
c37 13 0 1.40531e-19 $X=1.66 $Y=1.51
r38 12 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.66 $Y=1.51
+ $X2=1.66 $Y2=1.675
r39 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.66 $Y=1.51
+ $X2=1.66 $Y2=1.345
r40 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.66
+ $Y=1.51 $X2=1.66 $Y2=1.51
r41 9 13 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=1.66 $Y=1.665
+ $X2=1.66 $Y2=1.51
r42 7 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.75 $Y=2.465
+ $X2=1.75 $Y2=1.675
r43 3 14 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=1.67 $Y=0.665
+ $X2=1.67 $Y2=1.345
.ends

.subckt PM_SKY130_FD_SC_LP__O211A_1%A2 3 7 9 12 13
r34 12 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.2 $Y=1.51 $X2=2.2
+ $Y2=1.675
r35 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.2 $Y=1.51 $X2=2.2
+ $Y2=1.345
r36 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.2
+ $Y=1.51 $X2=2.2 $Y2=1.51
r37 9 13 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=2.2 $Y=1.665 $X2=2.2
+ $Y2=1.51
r38 7 14 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=2.29 $Y=0.665
+ $X2=2.29 $Y2=1.345
r39 3 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.11 $Y=2.465
+ $X2=2.11 $Y2=1.675
.ends

.subckt PM_SKY130_FD_SC_LP__O211A_1%B1 3 7 9 10 14
c33 14 0 1.35912e-19 $X=2.74 $Y=1.51
r34 14 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.74 $Y=1.51
+ $X2=2.74 $Y2=1.675
r35 14 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.74 $Y=1.51
+ $X2=2.74 $Y2=1.345
r36 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.74
+ $Y=1.51 $X2=2.74 $Y2=1.51
r37 10 15 11.3748 $w=3.83e-07 $l=3.8e-07 $layer=LI1_cond $X=3.12 $Y=1.557
+ $X2=2.74 $Y2=1.557
r38 9 15 2.99336 $w=3.83e-07 $l=1e-07 $layer=LI1_cond $X=2.64 $Y=1.557 $X2=2.74
+ $Y2=1.557
r39 7 16 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=2.83 $Y=0.665
+ $X2=2.83 $Y2=1.345
r40 3 17 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.65 $Y=2.465
+ $X2=2.65 $Y2=1.675
.ends

.subckt PM_SKY130_FD_SC_LP__O211A_1%C1 3 7 10 11 14 15
c27 15 0 1.35912e-19 $X=3.55 $Y=1.46
r28 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.55
+ $Y=1.46 $X2=3.55 $Y2=1.46
r29 11 15 6.38516 $w=3.68e-07 $l=2.05e-07 $layer=LI1_cond $X=3.57 $Y=1.665
+ $X2=3.57 $Y2=1.46
r30 9 14 49.8355 $w=3.3e-07 $l=2.85e-07 $layer=POLY_cond $X=3.265 $Y=1.46
+ $X2=3.55 $Y2=1.46
r31 9 10 5.03009 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=3.265 $Y=1.46
+ $X2=3.19 $Y2=1.46
r32 5 10 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.19 $Y=1.625
+ $X2=3.19 $Y2=1.46
r33 5 7 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=3.19 $Y=1.625 $X2=3.19
+ $Y2=2.465
r34 1 10 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.19 $Y=1.295
+ $X2=3.19 $Y2=1.46
r35 1 3 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=3.19 $Y=1.295 $X2=3.19
+ $Y2=0.665
.ends

.subckt PM_SKY130_FD_SC_LP__O211A_1%X 1 2 7 8 9 10 11 12 13 24 45 48
r19 48 49 8.63019 $w=7.73e-07 $l=1.65e-07 $layer=LI1_cond $X=0.472 $Y=1.98
+ $X2=0.472 $Y2=1.815
r20 45 46 3.40798 $w=3.28e-07 $l=7.5e-08 $layer=LI1_cond $X=0.25 $Y=0.925
+ $X2=0.25 $Y2=1
r21 13 41 2.08349 $w=7.73e-07 $l=1.35e-07 $layer=LI1_cond $X=0.472 $Y=2.775
+ $X2=0.472 $Y2=2.91
r22 12 13 5.71031 $w=7.73e-07 $l=3.7e-07 $layer=LI1_cond $X=0.472 $Y=2.405
+ $X2=0.472 $Y2=2.775
r23 12 35 3.13295 $w=7.73e-07 $l=2.03e-07 $layer=LI1_cond $X=0.472 $Y=2.405
+ $X2=0.472 $Y2=2.202
r24 11 35 2.57736 $w=7.73e-07 $l=1.67e-07 $layer=LI1_cond $X=0.472 $Y=2.035
+ $X2=0.472 $Y2=2.202
r25 11 48 0.84883 $w=7.73e-07 $l=5.5e-08 $layer=LI1_cond $X=0.472 $Y=2.035
+ $X2=0.472 $Y2=1.98
r26 10 49 7.05577 $w=2.43e-07 $l=1.5e-07 $layer=LI1_cond $X=0.207 $Y=1.665
+ $X2=0.207 $Y2=1.815
r27 9 10 17.4042 $w=2.43e-07 $l=3.7e-07 $layer=LI1_cond $X=0.207 $Y=1.295
+ $X2=0.207 $Y2=1.665
r28 8 45 0.174613 $w=3.28e-07 $l=5e-09 $layer=LI1_cond $X=0.25 $Y=0.92 $X2=0.25
+ $Y2=0.925
r29 8 22 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=0.25 $Y=0.92 $X2=0.25
+ $Y2=0.835
r30 8 9 13.6412 $w=2.43e-07 $l=2.9e-07 $layer=LI1_cond $X=0.207 $Y=1.005
+ $X2=0.207 $Y2=1.295
r31 8 46 0.235192 $w=2.43e-07 $l=5e-09 $layer=LI1_cond $X=0.207 $Y=1.005
+ $X2=0.207 $Y2=1
r32 7 22 9.7783 $w=3.28e-07 $l=2.8e-07 $layer=LI1_cond $X=0.25 $Y=0.555 $X2=0.25
+ $Y2=0.835
r33 7 24 4.71454 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=0.25 $Y=0.555
+ $X2=0.25 $Y2=0.42
r34 2 48 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.64
+ $Y=1.835 $X2=0.765 $Y2=1.98
r35 2 41 400 $w=1.7e-07 $l=1.13578e-06 $layer=licon1_PDIFF $count=1 $X=0.64
+ $Y=1.835 $X2=0.765 $Y2=2.91
r36 1 24 91 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=2 $X=0.195
+ $Y=0.235 $X2=0.32 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__O211A_1%VPWR 1 2 9 13 16 17 18 20 30 31 34
r41 35 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r42 34 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r43 34 35 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r44 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r45 28 31 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r46 27 28 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r47 25 34 13.3456 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=1.7 $Y=3.33
+ $X2=1.365 $Y2=3.33
r48 25 27 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=1.7 $Y=3.33 $X2=2.64
+ $Y2=3.33
r49 23 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r50 22 23 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r51 20 34 13.3456 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=1.03 $Y=3.33
+ $X2=1.365 $Y2=3.33
r52 20 22 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=1.03 $Y=3.33
+ $X2=0.72 $Y2=3.33
r53 18 28 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=2.64 $Y2=3.33
r54 18 35 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=1.68 $Y2=3.33
r55 16 27 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=2.75 $Y=3.33
+ $X2=2.64 $Y2=3.33
r56 16 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.75 $Y=3.33
+ $X2=2.915 $Y2=3.33
r57 15 30 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=3.08 $Y=3.33 $X2=3.6
+ $Y2=3.33
r58 15 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.08 $Y=3.33
+ $X2=2.915 $Y2=3.33
r59 11 17 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.915 $Y=3.245
+ $X2=2.915 $Y2=3.33
r60 11 13 30.7318 $w=3.28e-07 $l=8.8e-07 $layer=LI1_cond $X=2.915 $Y=3.245
+ $X2=2.915 $Y2=2.365
r61 7 34 2.76849 $w=6.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.365 $Y=3.245
+ $X2=1.365 $Y2=3.33
r62 7 9 15.7097 $w=6.68e-07 $l=8.8e-07 $layer=LI1_cond $X=1.365 $Y=3.245
+ $X2=1.365 $Y2=2.365
r63 2 13 300 $w=1.7e-07 $l=6.17738e-07 $layer=licon1_PDIFF $count=2 $X=2.725
+ $Y=1.835 $X2=2.915 $Y2=2.365
r64 1 9 150 $w=1.7e-07 $l=7.31642e-07 $layer=licon1_PDIFF $count=4 $X=1.055
+ $Y=1.835 $X2=1.535 $Y2=2.365
.ends

.subckt PM_SKY130_FD_SC_LP__O211A_1%VGND 1 2 9 13 16 17 18 20 33 34 37
r47 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r48 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r49 31 34 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.6
+ $Y2=0
r50 30 33 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=2.16 $Y=0 $X2=3.6
+ $Y2=0
r51 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r52 28 38 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=0.72
+ $Y2=0
r53 27 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r54 25 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.915 $Y=0 $X2=0.75
+ $Y2=0
r55 25 27 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=0.915 $Y=0 $X2=1.68
+ $Y2=0
r56 23 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r57 22 23 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r58 20 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.585 $Y=0 $X2=0.75
+ $Y2=0
r59 20 22 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.585 $Y=0 $X2=0.24
+ $Y2=0
r60 18 31 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=2.16
+ $Y2=0
r61 18 28 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=1.68
+ $Y2=0
r62 16 27 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=1.815 $Y=0 $X2=1.68
+ $Y2=0
r63 16 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.815 $Y=0 $X2=1.98
+ $Y2=0
r64 15 30 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=2.145 $Y=0 $X2=2.16
+ $Y2=0
r65 15 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.145 $Y=0 $X2=1.98
+ $Y2=0
r66 11 17 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.98 $Y=0.085
+ $X2=1.98 $Y2=0
r67 11 13 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=1.98 $Y=0.085
+ $X2=1.98 $Y2=0.41
r68 7 37 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.75 $Y=0.085 $X2=0.75
+ $Y2=0
r69 7 9 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.75 $Y=0.085
+ $X2=0.75 $Y2=0.38
r70 2 13 182 $w=1.7e-07 $l=3.06594e-07 $layer=licon1_NDIFF $count=1 $X=1.745
+ $Y=0.245 $X2=1.98 $Y2=0.41
r71 1 9 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=0.61
+ $Y=0.235 $X2=0.75 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_LP__O211A_1%A_266_49# 1 2 9 11 12 13 15
r29 13 18 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.56 $Y=0.685 $X2=2.56
+ $Y2=0.77
r30 13 15 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=2.56 $Y=0.685
+ $X2=2.56 $Y2=0.4
r31 11 18 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.395 $Y=0.77
+ $X2=2.56 $Y2=0.77
r32 11 12 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=2.395 $Y=0.77
+ $X2=1.62 $Y2=0.77
r33 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.455 $Y=0.685
+ $X2=1.62 $Y2=0.77
r34 7 9 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=1.455 $Y=0.685
+ $X2=1.455 $Y2=0.4
r35 2 18 182 $w=1.7e-07 $l=6.14817e-07 $layer=licon1_NDIFF $count=1 $X=2.365
+ $Y=0.245 $X2=2.56 $Y2=0.77
r36 2 15 182 $w=1.7e-07 $l=2.61247e-07 $layer=licon1_NDIFF $count=1 $X=2.365
+ $Y=0.245 $X2=2.56 $Y2=0.4
r37 1 9 91 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=2 $X=1.33
+ $Y=0.245 $X2=1.455 $Y2=0.4
.ends

