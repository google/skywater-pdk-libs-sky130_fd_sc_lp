# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__a32o_lp
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__a32o_lp ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.320000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.313000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.495000 1.235000 1.825000 1.905000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.313000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.045000 0.810000 2.395000 1.905000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.313000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.925000 1.550000 3.255000 1.880000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.313000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.925000 1.235000 1.315000 1.905000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.313000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.235000 0.685000 1.905000 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  0.442500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.865000 0.440000 4.205000 3.065000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 4.320000 0.085000 ;
        RECT 0.230000  0.085000 0.560000 1.055000 ;
        RECT 2.925000  0.085000 3.175000 1.020000 ;
      LAYER mcon ;
        RECT 0.155000 -0.085000 0.325000 0.085000 ;
        RECT 0.635000 -0.085000 0.805000 0.085000 ;
        RECT 1.115000 -0.085000 1.285000 0.085000 ;
        RECT 1.595000 -0.085000 1.765000 0.085000 ;
        RECT 2.075000 -0.085000 2.245000 0.085000 ;
        RECT 2.555000 -0.085000 2.725000 0.085000 ;
        RECT 3.035000 -0.085000 3.205000 0.085000 ;
        RECT 3.515000 -0.085000 3.685000 0.085000 ;
        RECT 3.995000 -0.085000 4.165000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.320000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.245000 4.320000 3.415000 ;
        RECT 1.720000 2.785000 2.050000 3.245000 ;
        RECT 2.925000 2.075000 3.255000 3.245000 ;
      LAYER mcon ;
        RECT 0.155000 3.245000 0.325000 3.415000 ;
        RECT 0.635000 3.245000 0.805000 3.415000 ;
        RECT 1.115000 3.245000 1.285000 3.415000 ;
        RECT 1.595000 3.245000 1.765000 3.415000 ;
        RECT 2.075000 3.245000 2.245000 3.415000 ;
        RECT 2.555000 3.245000 2.725000 3.415000 ;
        RECT 3.035000 3.245000 3.205000 3.415000 ;
        RECT 3.515000 3.245000 3.685000 3.415000 ;
        RECT 3.995000 3.245000 4.165000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 4.320000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.130000 2.085000 0.460000 2.895000 ;
      RECT 0.130000 2.895000 1.520000 3.065000 ;
      RECT 0.660000 2.085000 2.745000 2.255000 ;
      RECT 0.660000 2.255000 0.990000 2.715000 ;
      RECT 1.190000 0.460000 2.745000 0.630000 ;
      RECT 1.190000 0.630000 1.520000 1.055000 ;
      RECT 1.190000 2.435000 2.660000 2.605000 ;
      RECT 1.190000 2.605000 1.520000 2.895000 ;
      RECT 2.330000 2.605000 2.660000 3.065000 ;
      RECT 2.575000 0.630000 2.745000 1.200000 ;
      RECT 2.575000 1.200000 3.685000 1.370000 ;
      RECT 2.575000 1.370000 2.745000 2.085000 ;
      RECT 3.355000 0.265000 3.685000 1.200000 ;
  END
END sky130_fd_sc_lp__a32o_lp
