* File: sky130_fd_sc_lp__bufinv_16.pxi.spice
* Created: Wed Sep  2 09:35:42 2020
* 
x_PM_SKY130_FD_SC_LP__BUFINV_16%A N_A_M1006_g N_A_M1008_g N_A_M1017_g
+ N_A_M1022_g N_A_M1040_g N_A_M1026_g A A A N_A_c_202_n N_A_c_203_n N_A_c_204_n
+ PM_SKY130_FD_SC_LP__BUFINV_16%A
x_PM_SKY130_FD_SC_LP__BUFINV_16%A_63_49# N_A_63_49#_M1006_d N_A_63_49#_M1017_d
+ N_A_63_49#_M1008_d N_A_63_49#_M1022_d N_A_63_49#_M1001_g N_A_63_49#_M1004_g
+ N_A_63_49#_M1005_g N_A_63_49#_M1010_g N_A_63_49#_M1020_g N_A_63_49#_M1018_g
+ N_A_63_49#_M1035_g N_A_63_49#_M1033_g N_A_63_49#_M1037_g N_A_63_49#_M1042_g
+ N_A_63_49#_M1041_g N_A_63_49#_M1049_g N_A_63_49#_c_265_n N_A_63_49#_c_280_n
+ N_A_63_49#_c_281_n N_A_63_49#_c_266_n N_A_63_49#_c_267_n N_A_63_49#_c_295_n
+ N_A_63_49#_c_391_p N_A_63_49#_c_361_p N_A_63_49#_c_268_n N_A_63_49#_c_301_n
+ N_A_63_49#_c_269_n N_A_63_49#_c_270_n N_A_63_49#_c_318_p N_A_63_49#_c_271_n
+ N_A_63_49#_c_308_n N_A_63_49#_c_272_n N_A_63_49#_c_273_n
+ PM_SKY130_FD_SC_LP__BUFINV_16%A_63_49#
x_PM_SKY130_FD_SC_LP__BUFINV_16%A_413_49# N_A_413_49#_M1001_s
+ N_A_413_49#_M1020_s N_A_413_49#_M1037_s N_A_413_49#_M1004_d
+ N_A_413_49#_M1018_d N_A_413_49#_M1042_d N_A_413_49#_M1002_g
+ N_A_413_49#_M1000_g N_A_413_49#_M1003_g N_A_413_49#_M1007_g
+ N_A_413_49#_M1011_g N_A_413_49#_M1009_g N_A_413_49#_M1013_g
+ N_A_413_49#_M1012_g N_A_413_49#_M1014_g N_A_413_49#_M1015_g
+ N_A_413_49#_M1016_g N_A_413_49#_M1019_g N_A_413_49#_M1021_g
+ N_A_413_49#_M1024_g N_A_413_49#_M1023_g N_A_413_49#_M1025_g
+ N_A_413_49#_M1030_g N_A_413_49#_M1027_g N_A_413_49#_M1031_g
+ N_A_413_49#_M1028_g N_A_413_49#_M1032_g N_A_413_49#_M1029_g
+ N_A_413_49#_M1036_g N_A_413_49#_M1034_g N_A_413_49#_M1038_g
+ N_A_413_49#_M1039_g N_A_413_49#_M1044_g N_A_413_49#_M1043_g
+ N_A_413_49#_M1045_g N_A_413_49#_M1046_g N_A_413_49#_M1048_g
+ N_A_413_49#_M1047_g N_A_413_49#_c_756_p N_A_413_49#_c_582_p
+ N_A_413_49#_c_433_n N_A_413_49#_c_434_n N_A_413_49#_c_465_n
+ N_A_413_49#_c_466_n N_A_413_49#_c_746_p N_A_413_49#_c_572_p
+ N_A_413_49#_c_435_n N_A_413_49#_c_467_n N_A_413_49#_c_747_p
+ N_A_413_49#_c_573_p N_A_413_49#_c_436_n N_A_413_49#_c_468_n
+ N_A_413_49#_c_437_n N_A_413_49#_c_469_n N_A_413_49#_c_438_n
+ N_A_413_49#_c_470_n N_A_413_49#_c_439_n N_A_413_49#_c_440_n
+ N_A_413_49#_c_441_n N_A_413_49#_c_442_n N_A_413_49#_c_443_n
+ N_A_413_49#_c_444_n N_A_413_49#_c_445_n N_A_413_49#_c_446_n
+ N_A_413_49#_c_447_n N_A_413_49#_c_448_n
+ PM_SKY130_FD_SC_LP__BUFINV_16%A_413_49#
x_PM_SKY130_FD_SC_LP__BUFINV_16%VPWR N_VPWR_M1008_s N_VPWR_M1026_s
+ N_VPWR_M1010_s N_VPWR_M1033_s N_VPWR_M1049_s N_VPWR_M1007_s N_VPWR_M1012_s
+ N_VPWR_M1019_s N_VPWR_M1025_s N_VPWR_M1028_s N_VPWR_M1034_s N_VPWR_M1043_s
+ N_VPWR_M1047_s N_VPWR_c_784_n N_VPWR_c_785_n N_VPWR_c_786_n N_VPWR_c_787_n
+ N_VPWR_c_788_n N_VPWR_c_789_n N_VPWR_c_790_n N_VPWR_c_791_n N_VPWR_c_792_n
+ N_VPWR_c_793_n N_VPWR_c_794_n N_VPWR_c_795_n N_VPWR_c_796_n N_VPWR_c_797_n
+ N_VPWR_c_798_n N_VPWR_c_799_n N_VPWR_c_800_n N_VPWR_c_801_n N_VPWR_c_802_n
+ N_VPWR_c_803_n N_VPWR_c_804_n N_VPWR_c_805_n N_VPWR_c_806_n N_VPWR_c_807_n
+ N_VPWR_c_808_n N_VPWR_c_809_n N_VPWR_c_810_n N_VPWR_c_811_n N_VPWR_c_812_n
+ N_VPWR_c_813_n N_VPWR_c_814_n VPWR N_VPWR_c_815_n N_VPWR_c_816_n
+ N_VPWR_c_817_n N_VPWR_c_818_n N_VPWR_c_819_n N_VPWR_c_820_n N_VPWR_c_821_n
+ N_VPWR_c_822_n N_VPWR_c_783_n PM_SKY130_FD_SC_LP__BUFINV_16%VPWR
x_PM_SKY130_FD_SC_LP__BUFINV_16%Y N_Y_M1002_s N_Y_M1011_s N_Y_M1014_s
+ N_Y_M1021_s N_Y_M1030_s N_Y_M1032_s N_Y_M1038_s N_Y_M1045_s N_Y_M1000_d
+ N_Y_M1009_d N_Y_M1015_d N_Y_M1024_d N_Y_M1027_d N_Y_M1029_d N_Y_M1039_d
+ N_Y_M1046_d Y N_Y_c_1002_n N_Y_c_1003_n N_Y_c_1004_n N_Y_c_1005_n N_Y_c_1006_n
+ N_Y_c_1007_n N_Y_c_1008_n N_Y_c_1009_n N_Y_c_1018_n
+ PM_SKY130_FD_SC_LP__BUFINV_16%Y
x_PM_SKY130_FD_SC_LP__BUFINV_16%VGND N_VGND_M1006_s N_VGND_M1040_s
+ N_VGND_M1005_d N_VGND_M1035_d N_VGND_M1041_d N_VGND_M1003_d N_VGND_M1013_d
+ N_VGND_M1016_d N_VGND_M1023_d N_VGND_M1031_d N_VGND_M1036_d N_VGND_M1044_d
+ N_VGND_M1048_d N_VGND_c_1187_n N_VGND_c_1188_n N_VGND_c_1189_n N_VGND_c_1190_n
+ N_VGND_c_1191_n N_VGND_c_1192_n N_VGND_c_1193_n N_VGND_c_1194_n
+ N_VGND_c_1195_n N_VGND_c_1196_n N_VGND_c_1197_n N_VGND_c_1198_n
+ N_VGND_c_1199_n N_VGND_c_1200_n N_VGND_c_1201_n N_VGND_c_1202_n
+ N_VGND_c_1203_n N_VGND_c_1204_n N_VGND_c_1205_n N_VGND_c_1206_n
+ N_VGND_c_1207_n N_VGND_c_1208_n N_VGND_c_1209_n N_VGND_c_1210_n
+ N_VGND_c_1211_n N_VGND_c_1212_n N_VGND_c_1213_n N_VGND_c_1214_n
+ N_VGND_c_1215_n N_VGND_c_1216_n N_VGND_c_1217_n VGND N_VGND_c_1218_n
+ N_VGND_c_1219_n N_VGND_c_1220_n N_VGND_c_1221_n N_VGND_c_1222_n
+ N_VGND_c_1223_n N_VGND_c_1224_n N_VGND_c_1225_n N_VGND_c_1226_n
+ PM_SKY130_FD_SC_LP__BUFINV_16%VGND
cc_1 VNB N_A_M1006_g 0.0304968f $X=-0.19 $Y=-0.245 $X2=0.655 $Y2=0.665
cc_2 VNB N_A_M1017_g 0.0224424f $X=-0.19 $Y=-0.245 $X2=1.085 $Y2=0.665
cc_3 VNB N_A_M1040_g 0.0232243f $X=-0.19 $Y=-0.245 $X2=1.515 $Y2=0.665
cc_4 VNB N_A_c_202_n 0.0324653f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=1.51
cc_5 VNB N_A_c_203_n 0.0144179f $X=-0.19 $Y=-0.245 $X2=1.405 $Y2=1.51
cc_6 VNB N_A_c_204_n 0.0431533f $X=-0.19 $Y=-0.245 $X2=1.515 $Y2=1.51
cc_7 VNB N_A_63_49#_M1001_g 0.0224522f $X=-0.19 $Y=-0.245 $X2=1.085 $Y2=2.465
cc_8 VNB N_A_63_49#_M1005_g 0.0216055f $X=-0.19 $Y=-0.245 $X2=1.515 $Y2=2.465
cc_9 VNB N_A_63_49#_M1020_g 0.021612f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=1.51
cc_10 VNB N_A_63_49#_M1035_g 0.021612f $X=-0.19 $Y=-0.245 $X2=1.065 $Y2=1.51
cc_11 VNB N_A_63_49#_M1037_g 0.0215919f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_63_49#_M1041_g 0.0217958f $X=-0.19 $Y=-0.245 $X2=1.405 $Y2=1.587
cc_13 VNB N_A_63_49#_c_265_n 0.0293109f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_63_49#_c_266_n 0.00237397f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_63_49#_c_267_n 0.00940068f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_63_49#_c_268_n 0.0055449f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_63_49#_c_269_n 0.00141111f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_63_49#_c_270_n 4.19138e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_63_49#_c_271_n 0.00210048f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_63_49#_c_272_n 0.00128659f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_63_49#_c_273_n 0.109392f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_413_49#_M1002_g 0.0227106f $X=-0.19 $Y=-0.245 $X2=1.515 $Y2=1.675
cc_23 VNB N_A_413_49#_M1003_g 0.0237342f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_413_49#_M1011_g 0.0237342f $X=-0.19 $Y=-0.245 $X2=1.065 $Y2=1.51
cc_25 VNB N_A_413_49#_M1013_g 0.0237342f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_413_49#_M1014_g 0.0237342f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=1.587
cc_27 VNB N_A_413_49#_M1016_g 0.0237342f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_413_49#_M1021_g 0.0237342f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_413_49#_M1023_g 0.0237342f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_413_49#_M1030_g 0.0237342f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_413_49#_M1031_g 0.0237342f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_413_49#_M1032_g 0.0237342f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_413_49#_M1036_g 0.0237342f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_413_49#_M1038_g 0.0237342f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_413_49#_M1044_g 0.0237342f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_413_49#_M1045_g 0.0237342f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_413_49#_M1048_g 0.034068f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_413_49#_c_433_n 0.00240399f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_413_49#_c_434_n 0.00309169f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_413_49#_c_435_n 0.00240399f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_413_49#_c_436_n 0.00158938f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_413_49#_c_437_n 0.00210048f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_413_49#_c_438_n 0.00210048f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_413_49#_c_439_n 0.00353166f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_413_49#_c_440_n 0.00180974f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_413_49#_c_441_n 0.00109967f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_413_49#_c_442_n 0.00109967f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_413_49#_c_443_n 0.00109967f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_413_49#_c_444_n 0.00109967f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_413_49#_c_445_n 0.00109967f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_413_49#_c_446_n 0.00109967f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_413_49#_c_447_n 0.00109967f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_413_49#_c_448_n 0.281281f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_VPWR_c_783_n 0.48212f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_Y_c_1002_n 0.00422413f $X=-0.19 $Y=-0.245 $X2=1.065 $Y2=1.587
cc_56 VNB N_Y_c_1003_n 0.00495171f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_Y_c_1004_n 0.00495171f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_Y_c_1005_n 0.00495171f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_Y_c_1006_n 0.00495171f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_Y_c_1007_n 0.00495171f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_Y_c_1008_n 0.00495171f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_Y_c_1009_n 0.00531707f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_VGND_c_1187_n 0.00492713f $X=-0.19 $Y=-0.245 $X2=1.405 $Y2=1.51
cc_64 VNB N_VGND_c_1188_n 0.0168711f $X=-0.19 $Y=-0.245 $X2=1.515 $Y2=1.51
cc_65 VNB N_VGND_c_1189_n 0.00438473f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_VGND_c_1190_n 0.00432463f $X=-0.19 $Y=-0.245 $X2=1.065 $Y2=1.587
cc_67 VNB N_VGND_c_1191_n 0.00428049f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_VGND_c_1192_n 0.00428049f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_VGND_c_1193_n 0.00428049f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_VGND_c_1194_n 0.0168711f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_VGND_c_1195_n 0.00428049f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_VGND_c_1196_n 0.00428049f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_VGND_c_1197_n 0.00428049f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_VGND_c_1198_n 0.00428049f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_VGND_c_1199_n 0.00428049f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_VGND_c_1200_n 0.0168711f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_VGND_c_1201_n 0.00428049f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_VGND_c_1202_n 0.0117031f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_VGND_c_1203_n 0.0386371f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_VGND_c_1204_n 0.0232402f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_VGND_c_1205_n 0.00500104f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_VGND_c_1206_n 0.0168711f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_VGND_c_1207_n 0.00500104f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_VGND_c_1208_n 0.0168711f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_VGND_c_1209_n 0.00500104f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_VGND_c_1210_n 0.0171639f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_VGND_c_1211_n 0.00500104f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_VGND_c_1212_n 0.0168711f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_VGND_c_1213_n 0.00500104f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_VGND_c_1214_n 0.0168711f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_VGND_c_1215_n 0.00500104f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_VGND_c_1216_n 0.0168711f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_93 VNB N_VGND_c_1217_n 0.00500104f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_94 VNB N_VGND_c_1218_n 0.0181103f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_95 VNB N_VGND_c_1219_n 0.0168711f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_96 VNB N_VGND_c_1220_n 0.0168711f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_97 VNB N_VGND_c_1221_n 0.00519339f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_98 VNB N_VGND_c_1222_n 0.00500104f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_99 VNB N_VGND_c_1223_n 0.00500104f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_100 VNB N_VGND_c_1224_n 0.00500104f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_101 VNB N_VGND_c_1225_n 0.00500104f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_102 VNB N_VGND_c_1226_n 0.535877f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_103 VPB N_A_M1008_g 0.024227f $X=-0.19 $Y=1.655 $X2=0.655 $Y2=2.465
cc_104 VPB N_A_M1022_g 0.0180527f $X=-0.19 $Y=1.655 $X2=1.085 $Y2=2.465
cc_105 VPB N_A_M1026_g 0.0191551f $X=-0.19 $Y=1.655 $X2=1.515 $Y2=2.465
cc_106 VPB N_A_c_202_n 0.0115962f $X=-0.19 $Y=1.655 $X2=0.58 $Y2=1.51
cc_107 VPB N_A_c_203_n 0.0190145f $X=-0.19 $Y=1.655 $X2=1.405 $Y2=1.51
cc_108 VPB N_A_c_204_n 0.00829008f $X=-0.19 $Y=1.655 $X2=1.515 $Y2=1.51
cc_109 VPB N_A_63_49#_M1004_g 0.0195772f $X=-0.19 $Y=1.655 $X2=1.515 $Y2=0.665
cc_110 VPB N_A_63_49#_M1010_g 0.0190558f $X=-0.19 $Y=1.655 $X2=1.115 $Y2=1.58
cc_111 VPB N_A_63_49#_M1018_g 0.0190623f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_112 VPB N_A_63_49#_M1033_g 0.0190623f $X=-0.19 $Y=1.655 $X2=1.405 $Y2=1.51
cc_113 VPB N_A_63_49#_M1042_g 0.0190422f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_114 VPB N_A_63_49#_M1049_g 0.0192418f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_115 VPB N_A_63_49#_c_280_n 0.0074315f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_116 VPB N_A_63_49#_c_281_n 0.035609f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_117 VPB N_A_63_49#_c_270_n 0.00135637f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_118 VPB N_A_63_49#_c_273_n 0.0149705f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_119 VPB N_A_413_49#_M1000_g 0.0176802f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_120 VPB N_A_413_49#_M1007_g 0.0178841f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.51
cc_121 VPB N_A_413_49#_M1009_g 0.0178841f $X=-0.19 $Y=1.655 $X2=1.405 $Y2=1.51
cc_122 VPB N_A_413_49#_M1012_g 0.0178841f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.587
cc_123 VPB N_A_413_49#_M1015_g 0.0178841f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_124 VPB N_A_413_49#_M1019_g 0.0178841f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_125 VPB N_A_413_49#_M1024_g 0.0178841f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_126 VPB N_A_413_49#_M1025_g 0.0178841f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_127 VPB N_A_413_49#_M1027_g 0.0178841f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_128 VPB N_A_413_49#_M1028_g 0.0178841f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_129 VPB N_A_413_49#_M1029_g 0.0178841f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_130 VPB N_A_413_49#_M1034_g 0.0178841f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_131 VPB N_A_413_49#_M1039_g 0.0178841f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_132 VPB N_A_413_49#_M1043_g 0.0178841f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_133 VPB N_A_413_49#_M1046_g 0.018271f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_134 VPB N_A_413_49#_M1047_g 0.0260532f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_135 VPB N_A_413_49#_c_465_n 0.00240399f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_136 VPB N_A_413_49#_c_466_n 0.00259519f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_137 VPB N_A_413_49#_c_467_n 0.00240399f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_138 VPB N_A_413_49#_c_468_n 0.00146241f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_139 VPB N_A_413_49#_c_469_n 0.00210048f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_140 VPB N_A_413_49#_c_470_n 0.00210048f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_141 VPB N_A_413_49#_c_439_n 0.00126819f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_142 VPB N_A_413_49#_c_440_n 0.00419141f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_143 VPB N_A_413_49#_c_441_n 0.00269492f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_144 VPB N_A_413_49#_c_442_n 0.00269492f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_145 VPB N_A_413_49#_c_443_n 0.00269492f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_146 VPB N_A_413_49#_c_444_n 0.00269492f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_147 VPB N_A_413_49#_c_445_n 0.00269492f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_148 VPB N_A_413_49#_c_446_n 0.00269492f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_149 VPB N_A_413_49#_c_447_n 0.00269492f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_150 VPB N_A_413_49#_c_448_n 0.0582637f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_151 VPB N_VPWR_c_784_n 0.00461568f $X=-0.19 $Y=1.655 $X2=1.405 $Y2=1.51
cc_152 VPB N_VPWR_c_785_n 0.0168284f $X=-0.19 $Y=1.655 $X2=1.515 $Y2=1.51
cc_153 VPB N_VPWR_c_786_n 0.00425796f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_154 VPB N_VPWR_c_787_n 0.00400996f $X=-0.19 $Y=1.655 $X2=1.065 $Y2=1.587
cc_155 VPB N_VPWR_c_788_n 0.00400996f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_156 VPB N_VPWR_c_789_n 0.00400996f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_157 VPB N_VPWR_c_790_n 0.00400996f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_158 VPB N_VPWR_c_791_n 0.0168284f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_159 VPB N_VPWR_c_792_n 0.00400996f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_160 VPB N_VPWR_c_793_n 0.00400996f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_161 VPB N_VPWR_c_794_n 0.00400996f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_162 VPB N_VPWR_c_795_n 0.00400996f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_163 VPB N_VPWR_c_796_n 0.00400996f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_164 VPB N_VPWR_c_797_n 0.0168284f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_165 VPB N_VPWR_c_798_n 0.00400996f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_166 VPB N_VPWR_c_799_n 0.0116772f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_167 VPB N_VPWR_c_800_n 0.0497254f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_168 VPB N_VPWR_c_801_n 0.0231918f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_169 VPB N_VPWR_c_802_n 0.00497514f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_170 VPB N_VPWR_c_803_n 0.0168284f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_171 VPB N_VPWR_c_804_n 0.00497514f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_172 VPB N_VPWR_c_805_n 0.0168284f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_173 VPB N_VPWR_c_806_n 0.00497514f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_174 VPB N_VPWR_c_807_n 0.017127f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_175 VPB N_VPWR_c_808_n 0.00497514f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_176 VPB N_VPWR_c_809_n 0.0168284f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_177 VPB N_VPWR_c_810_n 0.00497514f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_178 VPB N_VPWR_c_811_n 0.0168284f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_179 VPB N_VPWR_c_812_n 0.00497514f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_180 VPB N_VPWR_c_813_n 0.0168284f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_181 VPB N_VPWR_c_814_n 0.00497514f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_182 VPB N_VPWR_c_815_n 0.0169564f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_183 VPB N_VPWR_c_816_n 0.0168284f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_184 VPB N_VPWR_c_817_n 0.0168284f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_185 VPB N_VPWR_c_818_n 0.00584071f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_186 VPB N_VPWR_c_819_n 0.00497514f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_187 VPB N_VPWR_c_820_n 0.00497514f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_188 VPB N_VPWR_c_821_n 0.00497514f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_189 VPB N_VPWR_c_822_n 0.00497514f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_190 VPB N_VPWR_c_783_n 0.0537326f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_191 VPB N_Y_c_1002_n 0.00145261f $X=-0.19 $Y=1.655 $X2=1.065 $Y2=1.587
cc_192 VPB N_Y_c_1003_n 0.00156948f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_193 VPB N_Y_c_1004_n 0.00156948f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_194 VPB N_Y_c_1005_n 0.00156948f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_195 VPB N_Y_c_1006_n 0.00156948f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_196 VPB N_Y_c_1007_n 0.00156948f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_197 VPB N_Y_c_1008_n 0.00156948f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_198 VPB N_Y_c_1009_n 0.00242769f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_199 N_A_M1040_g N_A_63_49#_M1001_g 0.0193336f $X=1.515 $Y=0.665 $X2=0 $Y2=0
cc_200 N_A_c_204_n N_A_63_49#_M1004_g 0.0294881f $X=1.515 $Y=1.51 $X2=0 $Y2=0
cc_201 N_A_c_202_n N_A_63_49#_c_280_n 0.00176049f $X=0.58 $Y=1.51 $X2=0 $Y2=0
cc_202 N_A_c_203_n N_A_63_49#_c_280_n 0.0236178f $X=1.405 $Y=1.51 $X2=0 $Y2=0
cc_203 N_A_M1006_g N_A_63_49#_c_266_n 0.0164614f $X=0.655 $Y=0.665 $X2=0 $Y2=0
cc_204 N_A_M1017_g N_A_63_49#_c_266_n 0.0150738f $X=1.085 $Y=0.665 $X2=0 $Y2=0
cc_205 N_A_c_202_n N_A_63_49#_c_266_n 2.19188e-19 $X=0.58 $Y=1.51 $X2=0 $Y2=0
cc_206 N_A_c_203_n N_A_63_49#_c_266_n 0.0440138f $X=1.405 $Y=1.51 $X2=0 $Y2=0
cc_207 N_A_c_204_n N_A_63_49#_c_266_n 0.00243542f $X=1.515 $Y=1.51 $X2=0 $Y2=0
cc_208 N_A_c_202_n N_A_63_49#_c_267_n 0.00748177f $X=0.58 $Y=1.51 $X2=0 $Y2=0
cc_209 N_A_c_203_n N_A_63_49#_c_267_n 0.0249518f $X=1.405 $Y=1.51 $X2=0 $Y2=0
cc_210 N_A_M1008_g N_A_63_49#_c_295_n 0.0129934f $X=0.655 $Y=2.465 $X2=0 $Y2=0
cc_211 N_A_M1022_g N_A_63_49#_c_295_n 0.0129934f $X=1.085 $Y=2.465 $X2=0 $Y2=0
cc_212 N_A_c_203_n N_A_63_49#_c_295_n 0.0400361f $X=1.405 $Y=1.51 $X2=0 $Y2=0
cc_213 N_A_c_204_n N_A_63_49#_c_295_n 5.64665e-19 $X=1.515 $Y=1.51 $X2=0 $Y2=0
cc_214 N_A_M1040_g N_A_63_49#_c_268_n 0.0158897f $X=1.515 $Y=0.665 $X2=0 $Y2=0
cc_215 N_A_c_203_n N_A_63_49#_c_268_n 0.0100336f $X=1.405 $Y=1.51 $X2=0 $Y2=0
cc_216 N_A_M1026_g N_A_63_49#_c_301_n 0.0138093f $X=1.515 $Y=2.465 $X2=0 $Y2=0
cc_217 N_A_c_203_n N_A_63_49#_c_301_n 0.00970221f $X=1.405 $Y=1.51 $X2=0 $Y2=0
cc_218 N_A_M1040_g N_A_63_49#_c_269_n 0.00314254f $X=1.515 $Y=0.665 $X2=0 $Y2=0
cc_219 N_A_c_203_n N_A_63_49#_c_270_n 0.0132367f $X=1.405 $Y=1.51 $X2=0 $Y2=0
cc_220 N_A_c_204_n N_A_63_49#_c_270_n 0.00474671f $X=1.515 $Y=1.51 $X2=0 $Y2=0
cc_221 N_A_c_203_n N_A_63_49#_c_271_n 0.0219959f $X=1.405 $Y=1.51 $X2=0 $Y2=0
cc_222 N_A_c_204_n N_A_63_49#_c_271_n 0.00253619f $X=1.515 $Y=1.51 $X2=0 $Y2=0
cc_223 N_A_c_203_n N_A_63_49#_c_308_n 0.018394f $X=1.405 $Y=1.51 $X2=0 $Y2=0
cc_224 N_A_c_204_n N_A_63_49#_c_308_n 6.37898e-19 $X=1.515 $Y=1.51 $X2=0 $Y2=0
cc_225 N_A_c_203_n N_A_63_49#_c_272_n 0.0144259f $X=1.405 $Y=1.51 $X2=0 $Y2=0
cc_226 N_A_c_204_n N_A_63_49#_c_272_n 0.00177913f $X=1.515 $Y=1.51 $X2=0 $Y2=0
cc_227 N_A_M1040_g N_A_63_49#_c_273_n 0.0217639f $X=1.515 $Y=0.665 $X2=0 $Y2=0
cc_228 N_A_c_203_n N_A_63_49#_c_273_n 2.59735e-19 $X=1.405 $Y=1.51 $X2=0 $Y2=0
cc_229 N_A_M1008_g N_VPWR_c_784_n 0.00367019f $X=0.655 $Y=2.465 $X2=0 $Y2=0
cc_230 N_A_M1022_g N_VPWR_c_784_n 0.00220704f $X=1.085 $Y=2.465 $X2=0 $Y2=0
cc_231 N_A_M1022_g N_VPWR_c_785_n 0.00585385f $X=1.085 $Y=2.465 $X2=0 $Y2=0
cc_232 N_A_M1026_g N_VPWR_c_785_n 0.00585385f $X=1.515 $Y=2.465 $X2=0 $Y2=0
cc_233 N_A_M1026_g N_VPWR_c_786_n 0.00238131f $X=1.515 $Y=2.465 $X2=0 $Y2=0
cc_234 N_A_M1008_g N_VPWR_c_801_n 0.00585385f $X=0.655 $Y=2.465 $X2=0 $Y2=0
cc_235 N_A_M1008_g N_VPWR_c_783_n 0.0118835f $X=0.655 $Y=2.465 $X2=0 $Y2=0
cc_236 N_A_M1022_g N_VPWR_c_783_n 0.0107375f $X=1.085 $Y=2.465 $X2=0 $Y2=0
cc_237 N_A_M1026_g N_VPWR_c_783_n 0.0108778f $X=1.515 $Y=2.465 $X2=0 $Y2=0
cc_238 N_A_M1006_g N_VGND_c_1187_n 0.003002f $X=0.655 $Y=0.665 $X2=0 $Y2=0
cc_239 N_A_M1017_g N_VGND_c_1187_n 0.00159325f $X=1.085 $Y=0.665 $X2=0 $Y2=0
cc_240 N_A_M1017_g N_VGND_c_1188_n 0.00575161f $X=1.085 $Y=0.665 $X2=0 $Y2=0
cc_241 N_A_M1040_g N_VGND_c_1188_n 0.00575161f $X=1.515 $Y=0.665 $X2=0 $Y2=0
cc_242 N_A_M1040_g N_VGND_c_1189_n 0.0016716f $X=1.515 $Y=0.665 $X2=0 $Y2=0
cc_243 N_A_M1006_g N_VGND_c_1204_n 0.00575161f $X=0.655 $Y=0.665 $X2=0 $Y2=0
cc_244 N_A_M1006_g N_VGND_c_1226_n 0.0116456f $X=0.655 $Y=0.665 $X2=0 $Y2=0
cc_245 N_A_M1017_g N_VGND_c_1226_n 0.0105815f $X=1.085 $Y=0.665 $X2=0 $Y2=0
cc_246 N_A_M1040_g N_VGND_c_1226_n 0.0107118f $X=1.515 $Y=0.665 $X2=0 $Y2=0
cc_247 N_A_63_49#_M1041_g N_A_413_49#_M1002_g 0.0211204f $X=4.14 $Y=0.665 $X2=0
+ $Y2=0
cc_248 N_A_63_49#_M1049_g N_A_413_49#_M1000_g 0.0211204f $X=4.14 $Y=2.465 $X2=0
+ $Y2=0
cc_249 N_A_63_49#_M1005_g N_A_413_49#_c_433_n 0.0146866f $X=2.42 $Y=0.665 $X2=0
+ $Y2=0
cc_250 N_A_63_49#_M1020_g N_A_413_49#_c_433_n 0.0150272f $X=2.85 $Y=0.665 $X2=0
+ $Y2=0
cc_251 N_A_63_49#_c_318_p N_A_413_49#_c_433_n 0.0420697f $X=4.005 $Y=1.49 $X2=0
+ $Y2=0
cc_252 N_A_63_49#_c_273_n N_A_413_49#_c_433_n 0.00243542f $X=4.14 $Y=1.49 $X2=0
+ $Y2=0
cc_253 N_A_63_49#_M1001_g N_A_413_49#_c_434_n 0.00133232f $X=1.99 $Y=0.665 $X2=0
+ $Y2=0
cc_254 N_A_63_49#_c_268_n N_A_413_49#_c_434_n 0.0128561f $X=1.75 $Y=1.16 $X2=0
+ $Y2=0
cc_255 N_A_63_49#_c_318_p N_A_413_49#_c_434_n 0.0199136f $X=4.005 $Y=1.49 $X2=0
+ $Y2=0
cc_256 N_A_63_49#_c_273_n N_A_413_49#_c_434_n 0.00253619f $X=4.14 $Y=1.49 $X2=0
+ $Y2=0
cc_257 N_A_63_49#_M1010_g N_A_413_49#_c_465_n 0.0144087f $X=2.42 $Y=2.465 $X2=0
+ $Y2=0
cc_258 N_A_63_49#_M1018_g N_A_413_49#_c_465_n 0.0146941f $X=2.85 $Y=2.465 $X2=0
+ $Y2=0
cc_259 N_A_63_49#_c_318_p N_A_413_49#_c_465_n 0.0420697f $X=4.005 $Y=1.49 $X2=0
+ $Y2=0
cc_260 N_A_63_49#_c_273_n N_A_413_49#_c_465_n 0.00243542f $X=4.14 $Y=1.49 $X2=0
+ $Y2=0
cc_261 N_A_63_49#_M1004_g N_A_413_49#_c_466_n 9.76207e-19 $X=1.99 $Y=2.465 $X2=0
+ $Y2=0
cc_262 N_A_63_49#_c_270_n N_A_413_49#_c_466_n 0.00947157f $X=1.835 $Y=1.93 $X2=0
+ $Y2=0
cc_263 N_A_63_49#_c_318_p N_A_413_49#_c_466_n 0.0199136f $X=4.005 $Y=1.49 $X2=0
+ $Y2=0
cc_264 N_A_63_49#_c_273_n N_A_413_49#_c_466_n 0.00253619f $X=4.14 $Y=1.49 $X2=0
+ $Y2=0
cc_265 N_A_63_49#_M1035_g N_A_413_49#_c_435_n 0.0150738f $X=3.28 $Y=0.665 $X2=0
+ $Y2=0
cc_266 N_A_63_49#_M1037_g N_A_413_49#_c_435_n 0.0150738f $X=3.71 $Y=0.665 $X2=0
+ $Y2=0
cc_267 N_A_63_49#_c_318_p N_A_413_49#_c_435_n 0.0420697f $X=4.005 $Y=1.49 $X2=0
+ $Y2=0
cc_268 N_A_63_49#_c_273_n N_A_413_49#_c_435_n 0.00243542f $X=4.14 $Y=1.49 $X2=0
+ $Y2=0
cc_269 N_A_63_49#_M1033_g N_A_413_49#_c_467_n 0.0147406f $X=3.28 $Y=2.465 $X2=0
+ $Y2=0
cc_270 N_A_63_49#_M1042_g N_A_413_49#_c_467_n 0.0147406f $X=3.71 $Y=2.465 $X2=0
+ $Y2=0
cc_271 N_A_63_49#_c_318_p N_A_413_49#_c_467_n 0.0420697f $X=4.005 $Y=1.49 $X2=0
+ $Y2=0
cc_272 N_A_63_49#_c_273_n N_A_413_49#_c_467_n 0.00243542f $X=4.14 $Y=1.49 $X2=0
+ $Y2=0
cc_273 N_A_63_49#_M1041_g N_A_413_49#_c_436_n 0.015528f $X=4.14 $Y=0.665 $X2=0
+ $Y2=0
cc_274 N_A_63_49#_c_318_p N_A_413_49#_c_436_n 0.00786198f $X=4.005 $Y=1.49 $X2=0
+ $Y2=0
cc_275 N_A_63_49#_M1049_g N_A_413_49#_c_468_n 0.0151482f $X=4.14 $Y=2.465 $X2=0
+ $Y2=0
cc_276 N_A_63_49#_c_318_p N_A_413_49#_c_468_n 0.00786198f $X=4.005 $Y=1.49 $X2=0
+ $Y2=0
cc_277 N_A_63_49#_c_318_p N_A_413_49#_c_437_n 0.021133f $X=4.005 $Y=1.49 $X2=0
+ $Y2=0
cc_278 N_A_63_49#_c_273_n N_A_413_49#_c_437_n 0.00253619f $X=4.14 $Y=1.49 $X2=0
+ $Y2=0
cc_279 N_A_63_49#_c_318_p N_A_413_49#_c_469_n 0.021133f $X=4.005 $Y=1.49 $X2=0
+ $Y2=0
cc_280 N_A_63_49#_c_273_n N_A_413_49#_c_469_n 0.00253619f $X=4.14 $Y=1.49 $X2=0
+ $Y2=0
cc_281 N_A_63_49#_c_318_p N_A_413_49#_c_438_n 0.021133f $X=4.005 $Y=1.49 $X2=0
+ $Y2=0
cc_282 N_A_63_49#_c_273_n N_A_413_49#_c_438_n 0.00253619f $X=4.14 $Y=1.49 $X2=0
+ $Y2=0
cc_283 N_A_63_49#_c_318_p N_A_413_49#_c_470_n 0.021133f $X=4.005 $Y=1.49 $X2=0
+ $Y2=0
cc_284 N_A_63_49#_c_273_n N_A_413_49#_c_470_n 0.00253619f $X=4.14 $Y=1.49 $X2=0
+ $Y2=0
cc_285 N_A_63_49#_M1041_g N_A_413_49#_c_439_n 0.00854994f $X=4.14 $Y=0.665 $X2=0
+ $Y2=0
cc_286 N_A_63_49#_c_318_p N_A_413_49#_c_439_n 0.0147047f $X=4.005 $Y=1.49 $X2=0
+ $Y2=0
cc_287 N_A_63_49#_c_318_p N_A_413_49#_c_440_n 0.0012111f $X=4.005 $Y=1.49 $X2=0
+ $Y2=0
cc_288 N_A_63_49#_c_273_n N_A_413_49#_c_440_n 0.00444749f $X=4.14 $Y=1.49 $X2=0
+ $Y2=0
cc_289 N_A_63_49#_c_273_n N_A_413_49#_c_448_n 0.0211204f $X=4.14 $Y=1.49 $X2=0
+ $Y2=0
cc_290 N_A_63_49#_c_295_n N_VPWR_M1008_s 0.00333177f $X=1.17 $Y=2.015 $X2=-0.19
+ $Y2=-0.245
cc_291 N_A_63_49#_c_301_n N_VPWR_M1026_s 0.00616023f $X=1.75 $Y=2.015 $X2=0
+ $Y2=0
cc_292 N_A_63_49#_c_270_n N_VPWR_M1026_s 0.00108319f $X=1.835 $Y=1.93 $X2=0
+ $Y2=0
cc_293 N_A_63_49#_c_295_n N_VPWR_c_784_n 0.0135055f $X=1.17 $Y=2.015 $X2=0 $Y2=0
cc_294 N_A_63_49#_c_361_p N_VPWR_c_785_n 0.0113476f $X=1.3 $Y=2.86 $X2=0 $Y2=0
cc_295 N_A_63_49#_M1004_g N_VPWR_c_786_n 0.00238131f $X=1.99 $Y=2.465 $X2=0
+ $Y2=0
cc_296 N_A_63_49#_c_301_n N_VPWR_c_786_n 0.0180358f $X=1.75 $Y=2.015 $X2=0 $Y2=0
cc_297 N_A_63_49#_c_273_n N_VPWR_c_786_n 2.74829e-19 $X=4.14 $Y=1.49 $X2=0 $Y2=0
cc_298 N_A_63_49#_M1010_g N_VPWR_c_787_n 0.0016342f $X=2.42 $Y=2.465 $X2=0 $Y2=0
cc_299 N_A_63_49#_M1018_g N_VPWR_c_787_n 0.0016342f $X=2.85 $Y=2.465 $X2=0 $Y2=0
cc_300 N_A_63_49#_M1033_g N_VPWR_c_788_n 0.0016342f $X=3.28 $Y=2.465 $X2=0 $Y2=0
cc_301 N_A_63_49#_M1042_g N_VPWR_c_788_n 0.0016342f $X=3.71 $Y=2.465 $X2=0 $Y2=0
cc_302 N_A_63_49#_M1049_g N_VPWR_c_789_n 0.0016342f $X=4.14 $Y=2.465 $X2=0 $Y2=0
cc_303 N_A_63_49#_c_281_n N_VPWR_c_801_n 0.0144351f $X=0.44 $Y=2.86 $X2=0 $Y2=0
cc_304 N_A_63_49#_M1018_g N_VPWR_c_803_n 0.00585385f $X=2.85 $Y=2.465 $X2=0
+ $Y2=0
cc_305 N_A_63_49#_M1033_g N_VPWR_c_803_n 0.00585385f $X=3.28 $Y=2.465 $X2=0
+ $Y2=0
cc_306 N_A_63_49#_M1042_g N_VPWR_c_805_n 0.00585385f $X=3.71 $Y=2.465 $X2=0
+ $Y2=0
cc_307 N_A_63_49#_M1049_g N_VPWR_c_805_n 0.00585385f $X=4.14 $Y=2.465 $X2=0
+ $Y2=0
cc_308 N_A_63_49#_M1004_g N_VPWR_c_815_n 0.00585385f $X=1.99 $Y=2.465 $X2=0
+ $Y2=0
cc_309 N_A_63_49#_M1010_g N_VPWR_c_815_n 0.00585385f $X=2.42 $Y=2.465 $X2=0
+ $Y2=0
cc_310 N_A_63_49#_M1008_d N_VPWR_c_783_n 0.00256983f $X=0.315 $Y=1.835 $X2=0
+ $Y2=0
cc_311 N_A_63_49#_M1022_d N_VPWR_c_783_n 0.00304497f $X=1.16 $Y=1.835 $X2=0
+ $Y2=0
cc_312 N_A_63_49#_M1004_g N_VPWR_c_783_n 0.0108778f $X=1.99 $Y=2.465 $X2=0 $Y2=0
cc_313 N_A_63_49#_M1010_g N_VPWR_c_783_n 0.0106302f $X=2.42 $Y=2.465 $X2=0 $Y2=0
cc_314 N_A_63_49#_M1018_g N_VPWR_c_783_n 0.0106302f $X=2.85 $Y=2.465 $X2=0 $Y2=0
cc_315 N_A_63_49#_M1033_g N_VPWR_c_783_n 0.0106302f $X=3.28 $Y=2.465 $X2=0 $Y2=0
cc_316 N_A_63_49#_M1042_g N_VPWR_c_783_n 0.0106302f $X=3.71 $Y=2.465 $X2=0 $Y2=0
cc_317 N_A_63_49#_M1049_g N_VPWR_c_783_n 0.0106555f $X=4.14 $Y=2.465 $X2=0 $Y2=0
cc_318 N_A_63_49#_c_281_n N_VPWR_c_783_n 0.0111051f $X=0.44 $Y=2.86 $X2=0 $Y2=0
cc_319 N_A_63_49#_c_361_p N_VPWR_c_783_n 0.00977851f $X=1.3 $Y=2.86 $X2=0 $Y2=0
cc_320 N_A_63_49#_M1049_g N_Y_c_1018_n 7.85395e-19 $X=4.14 $Y=2.465 $X2=0 $Y2=0
cc_321 N_A_63_49#_c_266_n N_VGND_M1006_s 0.00176461f $X=1.17 $Y=1.16 $X2=-0.19
+ $Y2=-0.245
cc_322 N_A_63_49#_c_268_n N_VGND_M1040_s 0.00227943f $X=1.75 $Y=1.16 $X2=0 $Y2=0
cc_323 N_A_63_49#_c_266_n N_VGND_c_1187_n 0.0135055f $X=1.17 $Y=1.16 $X2=0 $Y2=0
cc_324 N_A_63_49#_c_391_p N_VGND_c_1188_n 0.0108254f $X=1.3 $Y=0.48 $X2=0 $Y2=0
cc_325 N_A_63_49#_M1001_g N_VGND_c_1189_n 0.00156508f $X=1.99 $Y=0.665 $X2=0
+ $Y2=0
cc_326 N_A_63_49#_c_268_n N_VGND_c_1189_n 0.0180809f $X=1.75 $Y=1.16 $X2=0 $Y2=0
cc_327 N_A_63_49#_c_273_n N_VGND_c_1189_n 2.92189e-19 $X=4.14 $Y=1.49 $X2=0
+ $Y2=0
cc_328 N_A_63_49#_M1005_g N_VGND_c_1190_n 0.00163847f $X=2.42 $Y=0.665 $X2=0
+ $Y2=0
cc_329 N_A_63_49#_M1020_g N_VGND_c_1190_n 0.00159325f $X=2.85 $Y=0.665 $X2=0
+ $Y2=0
cc_330 N_A_63_49#_M1035_g N_VGND_c_1191_n 0.00159325f $X=3.28 $Y=0.665 $X2=0
+ $Y2=0
cc_331 N_A_63_49#_M1037_g N_VGND_c_1191_n 0.00159325f $X=3.71 $Y=0.665 $X2=0
+ $Y2=0
cc_332 N_A_63_49#_M1041_g N_VGND_c_1192_n 0.00159325f $X=4.14 $Y=0.665 $X2=0
+ $Y2=0
cc_333 N_A_63_49#_c_265_n N_VGND_c_1204_n 0.0137633f $X=0.44 $Y=0.48 $X2=0 $Y2=0
cc_334 N_A_63_49#_M1020_g N_VGND_c_1206_n 0.00575161f $X=2.85 $Y=0.665 $X2=0
+ $Y2=0
cc_335 N_A_63_49#_M1035_g N_VGND_c_1206_n 0.00575161f $X=3.28 $Y=0.665 $X2=0
+ $Y2=0
cc_336 N_A_63_49#_M1037_g N_VGND_c_1208_n 0.00575161f $X=3.71 $Y=0.665 $X2=0
+ $Y2=0
cc_337 N_A_63_49#_M1041_g N_VGND_c_1208_n 0.00575161f $X=4.14 $Y=0.665 $X2=0
+ $Y2=0
cc_338 N_A_63_49#_M1001_g N_VGND_c_1218_n 0.00575161f $X=1.99 $Y=0.665 $X2=0
+ $Y2=0
cc_339 N_A_63_49#_M1005_g N_VGND_c_1218_n 0.00575161f $X=2.42 $Y=0.665 $X2=0
+ $Y2=0
cc_340 N_A_63_49#_M1006_d N_VGND_c_1226_n 0.00255136f $X=0.315 $Y=0.245 $X2=0
+ $Y2=0
cc_341 N_A_63_49#_M1017_d N_VGND_c_1226_n 0.00305524f $X=1.16 $Y=0.245 $X2=0
+ $Y2=0
cc_342 N_A_63_49#_M1001_g N_VGND_c_1226_n 0.0108075f $X=1.99 $Y=0.665 $X2=0
+ $Y2=0
cc_343 N_A_63_49#_M1005_g N_VGND_c_1226_n 0.0105815f $X=2.42 $Y=0.665 $X2=0
+ $Y2=0
cc_344 N_A_63_49#_M1020_g N_VGND_c_1226_n 0.0105815f $X=2.85 $Y=0.665 $X2=0
+ $Y2=0
cc_345 N_A_63_49#_M1035_g N_VGND_c_1226_n 0.0105815f $X=3.28 $Y=0.665 $X2=0
+ $Y2=0
cc_346 N_A_63_49#_M1037_g N_VGND_c_1226_n 0.0105815f $X=3.71 $Y=0.665 $X2=0
+ $Y2=0
cc_347 N_A_63_49#_M1041_g N_VGND_c_1226_n 0.0106069f $X=4.14 $Y=0.665 $X2=0
+ $Y2=0
cc_348 N_A_63_49#_c_265_n N_VGND_c_1226_n 0.0110438f $X=0.44 $Y=0.48 $X2=0 $Y2=0
cc_349 N_A_63_49#_c_391_p N_VGND_c_1226_n 0.00972454f $X=1.3 $Y=0.48 $X2=0 $Y2=0
cc_350 N_A_413_49#_c_465_n N_VPWR_M1010_s 0.00180746f $X=2.935 $Y=1.84 $X2=0
+ $Y2=0
cc_351 N_A_413_49#_c_467_n N_VPWR_M1033_s 0.00180746f $X=3.795 $Y=1.84 $X2=0
+ $Y2=0
cc_352 N_A_413_49#_c_468_n N_VPWR_M1049_s 0.00184059f $X=4.34 $Y=1.84 $X2=0
+ $Y2=0
cc_353 N_A_413_49#_c_465_n N_VPWR_c_787_n 0.0129403f $X=2.935 $Y=1.84 $X2=0
+ $Y2=0
cc_354 N_A_413_49#_c_467_n N_VPWR_c_788_n 0.0129403f $X=3.795 $Y=1.84 $X2=0
+ $Y2=0
cc_355 N_A_413_49#_M1000_g N_VPWR_c_789_n 0.0016342f $X=4.57 $Y=2.465 $X2=0
+ $Y2=0
cc_356 N_A_413_49#_c_468_n N_VPWR_c_789_n 0.0128326f $X=4.34 $Y=1.84 $X2=0 $Y2=0
cc_357 N_A_413_49#_c_440_n N_VPWR_c_789_n 0.0011754f $X=10.375 $Y=1.665 $X2=0
+ $Y2=0
cc_358 N_A_413_49#_M1007_g N_VPWR_c_790_n 0.00195587f $X=5 $Y=2.465 $X2=0 $Y2=0
cc_359 N_A_413_49#_M1009_g N_VPWR_c_790_n 0.00195587f $X=5.43 $Y=2.465 $X2=0
+ $Y2=0
cc_360 N_A_413_49#_c_440_n N_VPWR_c_790_n 2.64819e-19 $X=10.375 $Y=1.665 $X2=0
+ $Y2=0
cc_361 N_A_413_49#_c_441_n N_VPWR_c_790_n 0.0167299f $X=5.215 $Y=1.51 $X2=0
+ $Y2=0
cc_362 N_A_413_49#_c_448_n N_VPWR_c_790_n 5.09955e-19 $X=11.02 $Y=1.51 $X2=0
+ $Y2=0
cc_363 N_A_413_49#_M1009_g N_VPWR_c_791_n 0.00585385f $X=5.43 $Y=2.465 $X2=0
+ $Y2=0
cc_364 N_A_413_49#_M1012_g N_VPWR_c_791_n 0.00585385f $X=5.86 $Y=2.465 $X2=0
+ $Y2=0
cc_365 N_A_413_49#_M1012_g N_VPWR_c_792_n 0.00195587f $X=5.86 $Y=2.465 $X2=0
+ $Y2=0
cc_366 N_A_413_49#_M1015_g N_VPWR_c_792_n 0.00195587f $X=6.29 $Y=2.465 $X2=0
+ $Y2=0
cc_367 N_A_413_49#_c_440_n N_VPWR_c_792_n 2.64819e-19 $X=10.375 $Y=1.665 $X2=0
+ $Y2=0
cc_368 N_A_413_49#_c_442_n N_VPWR_c_792_n 0.0167299f $X=6.075 $Y=1.51 $X2=0
+ $Y2=0
cc_369 N_A_413_49#_c_448_n N_VPWR_c_792_n 5.09955e-19 $X=11.02 $Y=1.51 $X2=0
+ $Y2=0
cc_370 N_A_413_49#_M1019_g N_VPWR_c_793_n 0.00195587f $X=6.72 $Y=2.465 $X2=0
+ $Y2=0
cc_371 N_A_413_49#_M1024_g N_VPWR_c_793_n 0.00195587f $X=7.15 $Y=2.465 $X2=0
+ $Y2=0
cc_372 N_A_413_49#_c_440_n N_VPWR_c_793_n 2.64819e-19 $X=10.375 $Y=1.665 $X2=0
+ $Y2=0
cc_373 N_A_413_49#_c_443_n N_VPWR_c_793_n 0.0167299f $X=6.935 $Y=1.51 $X2=0
+ $Y2=0
cc_374 N_A_413_49#_c_448_n N_VPWR_c_793_n 5.09955e-19 $X=11.02 $Y=1.51 $X2=0
+ $Y2=0
cc_375 N_A_413_49#_M1025_g N_VPWR_c_794_n 0.00195587f $X=7.58 $Y=2.465 $X2=0
+ $Y2=0
cc_376 N_A_413_49#_M1027_g N_VPWR_c_794_n 0.00195587f $X=8.01 $Y=2.465 $X2=0
+ $Y2=0
cc_377 N_A_413_49#_c_440_n N_VPWR_c_794_n 2.64819e-19 $X=10.375 $Y=1.665 $X2=0
+ $Y2=0
cc_378 N_A_413_49#_c_444_n N_VPWR_c_794_n 0.0167299f $X=7.795 $Y=1.51 $X2=0
+ $Y2=0
cc_379 N_A_413_49#_c_448_n N_VPWR_c_794_n 5.09955e-19 $X=11.02 $Y=1.51 $X2=0
+ $Y2=0
cc_380 N_A_413_49#_M1028_g N_VPWR_c_795_n 0.00195587f $X=8.44 $Y=2.465 $X2=0
+ $Y2=0
cc_381 N_A_413_49#_M1029_g N_VPWR_c_795_n 0.00195587f $X=8.87 $Y=2.465 $X2=0
+ $Y2=0
cc_382 N_A_413_49#_c_440_n N_VPWR_c_795_n 2.64819e-19 $X=10.375 $Y=1.665 $X2=0
+ $Y2=0
cc_383 N_A_413_49#_c_445_n N_VPWR_c_795_n 0.0167299f $X=8.655 $Y=1.51 $X2=0
+ $Y2=0
cc_384 N_A_413_49#_c_448_n N_VPWR_c_795_n 5.09955e-19 $X=11.02 $Y=1.51 $X2=0
+ $Y2=0
cc_385 N_A_413_49#_M1034_g N_VPWR_c_796_n 0.00195587f $X=9.3 $Y=2.465 $X2=0
+ $Y2=0
cc_386 N_A_413_49#_M1039_g N_VPWR_c_796_n 0.00195587f $X=9.73 $Y=2.465 $X2=0
+ $Y2=0
cc_387 N_A_413_49#_c_440_n N_VPWR_c_796_n 2.64819e-19 $X=10.375 $Y=1.665 $X2=0
+ $Y2=0
cc_388 N_A_413_49#_c_446_n N_VPWR_c_796_n 0.0167299f $X=9.515 $Y=1.51 $X2=0
+ $Y2=0
cc_389 N_A_413_49#_c_448_n N_VPWR_c_796_n 5.09955e-19 $X=11.02 $Y=1.51 $X2=0
+ $Y2=0
cc_390 N_A_413_49#_M1039_g N_VPWR_c_797_n 0.00585385f $X=9.73 $Y=2.465 $X2=0
+ $Y2=0
cc_391 N_A_413_49#_M1043_g N_VPWR_c_797_n 0.00585385f $X=10.16 $Y=2.465 $X2=0
+ $Y2=0
cc_392 N_A_413_49#_M1043_g N_VPWR_c_798_n 0.00195587f $X=10.16 $Y=2.465 $X2=0
+ $Y2=0
cc_393 N_A_413_49#_M1046_g N_VPWR_c_798_n 0.00195587f $X=10.59 $Y=2.465 $X2=0
+ $Y2=0
cc_394 N_A_413_49#_c_440_n N_VPWR_c_798_n 2.64819e-19 $X=10.375 $Y=1.665 $X2=0
+ $Y2=0
cc_395 N_A_413_49#_c_447_n N_VPWR_c_798_n 0.0167299f $X=10.375 $Y=1.51 $X2=0
+ $Y2=0
cc_396 N_A_413_49#_c_448_n N_VPWR_c_798_n 5.09955e-19 $X=11.02 $Y=1.51 $X2=0
+ $Y2=0
cc_397 N_A_413_49#_M1047_g N_VPWR_c_800_n 0.00363905f $X=11.02 $Y=2.465 $X2=0
+ $Y2=0
cc_398 N_A_413_49#_c_572_p N_VPWR_c_803_n 0.0113476f $X=3.065 $Y=2.095 $X2=0
+ $Y2=0
cc_399 N_A_413_49#_c_573_p N_VPWR_c_805_n 0.0113476f $X=3.925 $Y=2.095 $X2=0
+ $Y2=0
cc_400 N_A_413_49#_M1000_g N_VPWR_c_807_n 0.00585385f $X=4.57 $Y=2.465 $X2=0
+ $Y2=0
cc_401 N_A_413_49#_M1007_g N_VPWR_c_807_n 0.00585385f $X=5 $Y=2.465 $X2=0 $Y2=0
cc_402 N_A_413_49#_M1024_g N_VPWR_c_809_n 0.00585385f $X=7.15 $Y=2.465 $X2=0
+ $Y2=0
cc_403 N_A_413_49#_M1025_g N_VPWR_c_809_n 0.00585385f $X=7.58 $Y=2.465 $X2=0
+ $Y2=0
cc_404 N_A_413_49#_M1027_g N_VPWR_c_811_n 0.00585385f $X=8.01 $Y=2.465 $X2=0
+ $Y2=0
cc_405 N_A_413_49#_M1028_g N_VPWR_c_811_n 0.00585385f $X=8.44 $Y=2.465 $X2=0
+ $Y2=0
cc_406 N_A_413_49#_M1029_g N_VPWR_c_813_n 0.00585385f $X=8.87 $Y=2.465 $X2=0
+ $Y2=0
cc_407 N_A_413_49#_M1034_g N_VPWR_c_813_n 0.00585385f $X=9.3 $Y=2.465 $X2=0
+ $Y2=0
cc_408 N_A_413_49#_c_582_p N_VPWR_c_815_n 0.0109351f $X=2.205 $Y=2.095 $X2=0
+ $Y2=0
cc_409 N_A_413_49#_M1015_g N_VPWR_c_816_n 0.00585385f $X=6.29 $Y=2.465 $X2=0
+ $Y2=0
cc_410 N_A_413_49#_M1019_g N_VPWR_c_816_n 0.00585385f $X=6.72 $Y=2.465 $X2=0
+ $Y2=0
cc_411 N_A_413_49#_M1046_g N_VPWR_c_817_n 0.00585385f $X=10.59 $Y=2.465 $X2=0
+ $Y2=0
cc_412 N_A_413_49#_M1047_g N_VPWR_c_817_n 0.00585385f $X=11.02 $Y=2.465 $X2=0
+ $Y2=0
cc_413 N_A_413_49#_M1004_d N_VPWR_c_783_n 0.00356516f $X=2.065 $Y=1.835 $X2=0
+ $Y2=0
cc_414 N_A_413_49#_M1018_d N_VPWR_c_783_n 0.00304497f $X=2.925 $Y=1.835 $X2=0
+ $Y2=0
cc_415 N_A_413_49#_M1042_d N_VPWR_c_783_n 0.00304497f $X=3.785 $Y=1.835 $X2=0
+ $Y2=0
cc_416 N_A_413_49#_M1000_g N_VPWR_c_783_n 0.0106555f $X=4.57 $Y=2.465 $X2=0
+ $Y2=0
cc_417 N_A_413_49#_M1007_g N_VPWR_c_783_n 0.0106302f $X=5 $Y=2.465 $X2=0 $Y2=0
cc_418 N_A_413_49#_M1009_g N_VPWR_c_783_n 0.0106302f $X=5.43 $Y=2.465 $X2=0
+ $Y2=0
cc_419 N_A_413_49#_M1012_g N_VPWR_c_783_n 0.0106302f $X=5.86 $Y=2.465 $X2=0
+ $Y2=0
cc_420 N_A_413_49#_M1015_g N_VPWR_c_783_n 0.0106302f $X=6.29 $Y=2.465 $X2=0
+ $Y2=0
cc_421 N_A_413_49#_M1019_g N_VPWR_c_783_n 0.0106302f $X=6.72 $Y=2.465 $X2=0
+ $Y2=0
cc_422 N_A_413_49#_M1024_g N_VPWR_c_783_n 0.0106302f $X=7.15 $Y=2.465 $X2=0
+ $Y2=0
cc_423 N_A_413_49#_M1025_g N_VPWR_c_783_n 0.0106302f $X=7.58 $Y=2.465 $X2=0
+ $Y2=0
cc_424 N_A_413_49#_M1027_g N_VPWR_c_783_n 0.0106302f $X=8.01 $Y=2.465 $X2=0
+ $Y2=0
cc_425 N_A_413_49#_M1028_g N_VPWR_c_783_n 0.0106302f $X=8.44 $Y=2.465 $X2=0
+ $Y2=0
cc_426 N_A_413_49#_M1029_g N_VPWR_c_783_n 0.0106302f $X=8.87 $Y=2.465 $X2=0
+ $Y2=0
cc_427 N_A_413_49#_M1034_g N_VPWR_c_783_n 0.0106302f $X=9.3 $Y=2.465 $X2=0 $Y2=0
cc_428 N_A_413_49#_M1039_g N_VPWR_c_783_n 0.0106302f $X=9.73 $Y=2.465 $X2=0
+ $Y2=0
cc_429 N_A_413_49#_M1043_g N_VPWR_c_783_n 0.0106302f $X=10.16 $Y=2.465 $X2=0
+ $Y2=0
cc_430 N_A_413_49#_M1046_g N_VPWR_c_783_n 0.0104456f $X=10.59 $Y=2.465 $X2=0
+ $Y2=0
cc_431 N_A_413_49#_M1047_g N_VPWR_c_783_n 0.0115856f $X=11.02 $Y=2.465 $X2=0
+ $Y2=0
cc_432 N_A_413_49#_c_582_p N_VPWR_c_783_n 0.00920999f $X=2.205 $Y=2.095 $X2=0
+ $Y2=0
cc_433 N_A_413_49#_c_572_p N_VPWR_c_783_n 0.00977851f $X=3.065 $Y=2.095 $X2=0
+ $Y2=0
cc_434 N_A_413_49#_c_573_p N_VPWR_c_783_n 0.00977851f $X=3.925 $Y=2.095 $X2=0
+ $Y2=0
cc_435 N_A_413_49#_M1002_g N_Y_c_1002_n 0.0020667f $X=4.57 $Y=0.665 $X2=0 $Y2=0
cc_436 N_A_413_49#_M1000_g N_Y_c_1002_n 0.00202698f $X=4.57 $Y=2.465 $X2=0 $Y2=0
cc_437 N_A_413_49#_M1003_g N_Y_c_1002_n 0.00383412f $X=5 $Y=0.665 $X2=0 $Y2=0
cc_438 N_A_413_49#_M1007_g N_Y_c_1002_n 0.00209454f $X=5 $Y=2.465 $X2=0 $Y2=0
cc_439 N_A_413_49#_c_436_n N_Y_c_1002_n 0.0126411f $X=4.34 $Y=1.14 $X2=0 $Y2=0
cc_440 N_A_413_49#_c_468_n N_Y_c_1002_n 0.0100042f $X=4.34 $Y=1.84 $X2=0 $Y2=0
cc_441 N_A_413_49#_c_439_n N_Y_c_1002_n 0.0365452f $X=4.435 $Y=1.665 $X2=0 $Y2=0
cc_442 N_A_413_49#_c_440_n N_Y_c_1002_n 0.0255158f $X=10.375 $Y=1.665 $X2=0
+ $Y2=0
cc_443 N_A_413_49#_c_441_n N_Y_c_1002_n 0.0306919f $X=5.215 $Y=1.51 $X2=0 $Y2=0
cc_444 N_A_413_49#_c_448_n N_Y_c_1002_n 0.0192745f $X=11.02 $Y=1.51 $X2=0 $Y2=0
cc_445 N_A_413_49#_M1011_g N_Y_c_1003_n 0.00391701f $X=5.43 $Y=0.665 $X2=0 $Y2=0
cc_446 N_A_413_49#_M1009_g N_Y_c_1003_n 0.00212348f $X=5.43 $Y=2.465 $X2=0 $Y2=0
cc_447 N_A_413_49#_M1013_g N_Y_c_1003_n 0.00391701f $X=5.86 $Y=0.665 $X2=0 $Y2=0
cc_448 N_A_413_49#_M1012_g N_Y_c_1003_n 0.00212348f $X=5.86 $Y=2.465 $X2=0 $Y2=0
cc_449 N_A_413_49#_c_440_n N_Y_c_1003_n 0.028855f $X=10.375 $Y=1.665 $X2=0 $Y2=0
cc_450 N_A_413_49#_c_441_n N_Y_c_1003_n 0.0308809f $X=5.215 $Y=1.51 $X2=0 $Y2=0
cc_451 N_A_413_49#_c_442_n N_Y_c_1003_n 0.0308809f $X=6.075 $Y=1.51 $X2=0 $Y2=0
cc_452 N_A_413_49#_c_448_n N_Y_c_1003_n 0.0205422f $X=11.02 $Y=1.51 $X2=0 $Y2=0
cc_453 N_A_413_49#_M1014_g N_Y_c_1004_n 0.00391701f $X=6.29 $Y=0.665 $X2=0 $Y2=0
cc_454 N_A_413_49#_M1015_g N_Y_c_1004_n 0.00212348f $X=6.29 $Y=2.465 $X2=0 $Y2=0
cc_455 N_A_413_49#_M1016_g N_Y_c_1004_n 0.00391701f $X=6.72 $Y=0.665 $X2=0 $Y2=0
cc_456 N_A_413_49#_M1019_g N_Y_c_1004_n 0.00212348f $X=6.72 $Y=2.465 $X2=0 $Y2=0
cc_457 N_A_413_49#_c_440_n N_Y_c_1004_n 0.028855f $X=10.375 $Y=1.665 $X2=0 $Y2=0
cc_458 N_A_413_49#_c_442_n N_Y_c_1004_n 0.0308809f $X=6.075 $Y=1.51 $X2=0 $Y2=0
cc_459 N_A_413_49#_c_443_n N_Y_c_1004_n 0.0308809f $X=6.935 $Y=1.51 $X2=0 $Y2=0
cc_460 N_A_413_49#_c_448_n N_Y_c_1004_n 0.0205422f $X=11.02 $Y=1.51 $X2=0 $Y2=0
cc_461 N_A_413_49#_M1021_g N_Y_c_1005_n 0.00391701f $X=7.15 $Y=0.665 $X2=0 $Y2=0
cc_462 N_A_413_49#_M1024_g N_Y_c_1005_n 0.00212348f $X=7.15 $Y=2.465 $X2=0 $Y2=0
cc_463 N_A_413_49#_M1023_g N_Y_c_1005_n 0.00391701f $X=7.58 $Y=0.665 $X2=0 $Y2=0
cc_464 N_A_413_49#_M1025_g N_Y_c_1005_n 0.00212348f $X=7.58 $Y=2.465 $X2=0 $Y2=0
cc_465 N_A_413_49#_c_440_n N_Y_c_1005_n 0.028855f $X=10.375 $Y=1.665 $X2=0 $Y2=0
cc_466 N_A_413_49#_c_443_n N_Y_c_1005_n 0.0308809f $X=6.935 $Y=1.51 $X2=0 $Y2=0
cc_467 N_A_413_49#_c_444_n N_Y_c_1005_n 0.0308809f $X=7.795 $Y=1.51 $X2=0 $Y2=0
cc_468 N_A_413_49#_c_448_n N_Y_c_1005_n 0.0205422f $X=11.02 $Y=1.51 $X2=0 $Y2=0
cc_469 N_A_413_49#_M1030_g N_Y_c_1006_n 0.00391701f $X=8.01 $Y=0.665 $X2=0 $Y2=0
cc_470 N_A_413_49#_M1027_g N_Y_c_1006_n 0.00212348f $X=8.01 $Y=2.465 $X2=0 $Y2=0
cc_471 N_A_413_49#_M1031_g N_Y_c_1006_n 0.00391701f $X=8.44 $Y=0.665 $X2=0 $Y2=0
cc_472 N_A_413_49#_M1028_g N_Y_c_1006_n 0.00212348f $X=8.44 $Y=2.465 $X2=0 $Y2=0
cc_473 N_A_413_49#_c_440_n N_Y_c_1006_n 0.028855f $X=10.375 $Y=1.665 $X2=0 $Y2=0
cc_474 N_A_413_49#_c_444_n N_Y_c_1006_n 0.0308809f $X=7.795 $Y=1.51 $X2=0 $Y2=0
cc_475 N_A_413_49#_c_445_n N_Y_c_1006_n 0.0308809f $X=8.655 $Y=1.51 $X2=0 $Y2=0
cc_476 N_A_413_49#_c_448_n N_Y_c_1006_n 0.0205422f $X=11.02 $Y=1.51 $X2=0 $Y2=0
cc_477 N_A_413_49#_M1032_g N_Y_c_1007_n 0.00391701f $X=8.87 $Y=0.665 $X2=0 $Y2=0
cc_478 N_A_413_49#_M1029_g N_Y_c_1007_n 0.00212348f $X=8.87 $Y=2.465 $X2=0 $Y2=0
cc_479 N_A_413_49#_M1036_g N_Y_c_1007_n 0.00391701f $X=9.3 $Y=0.665 $X2=0 $Y2=0
cc_480 N_A_413_49#_M1034_g N_Y_c_1007_n 0.00212348f $X=9.3 $Y=2.465 $X2=0 $Y2=0
cc_481 N_A_413_49#_c_440_n N_Y_c_1007_n 0.028855f $X=10.375 $Y=1.665 $X2=0 $Y2=0
cc_482 N_A_413_49#_c_445_n N_Y_c_1007_n 0.0308809f $X=8.655 $Y=1.51 $X2=0 $Y2=0
cc_483 N_A_413_49#_c_446_n N_Y_c_1007_n 0.0308809f $X=9.515 $Y=1.51 $X2=0 $Y2=0
cc_484 N_A_413_49#_c_448_n N_Y_c_1007_n 0.0205422f $X=11.02 $Y=1.51 $X2=0 $Y2=0
cc_485 N_A_413_49#_M1038_g N_Y_c_1008_n 0.00391701f $X=9.73 $Y=0.665 $X2=0 $Y2=0
cc_486 N_A_413_49#_M1039_g N_Y_c_1008_n 0.00212348f $X=9.73 $Y=2.465 $X2=0 $Y2=0
cc_487 N_A_413_49#_M1044_g N_Y_c_1008_n 0.00391701f $X=10.16 $Y=0.665 $X2=0
+ $Y2=0
cc_488 N_A_413_49#_M1043_g N_Y_c_1008_n 0.00212348f $X=10.16 $Y=2.465 $X2=0
+ $Y2=0
cc_489 N_A_413_49#_c_440_n N_Y_c_1008_n 0.028855f $X=10.375 $Y=1.665 $X2=0 $Y2=0
cc_490 N_A_413_49#_c_446_n N_Y_c_1008_n 0.0308809f $X=9.515 $Y=1.51 $X2=0 $Y2=0
cc_491 N_A_413_49#_c_447_n N_Y_c_1008_n 0.0308809f $X=10.375 $Y=1.51 $X2=0 $Y2=0
cc_492 N_A_413_49#_c_448_n N_Y_c_1008_n 0.0205422f $X=11.02 $Y=1.51 $X2=0 $Y2=0
cc_493 N_A_413_49#_M1045_g N_Y_c_1009_n 0.00391701f $X=10.59 $Y=0.665 $X2=0
+ $Y2=0
cc_494 N_A_413_49#_M1046_g N_Y_c_1009_n 0.00223604f $X=10.59 $Y=2.465 $X2=0
+ $Y2=0
cc_495 N_A_413_49#_M1048_g N_Y_c_1009_n 0.00728339f $X=11.02 $Y=0.665 $X2=0
+ $Y2=0
cc_496 N_A_413_49#_M1047_g N_Y_c_1009_n 0.00519805f $X=11.02 $Y=2.465 $X2=0
+ $Y2=0
cc_497 N_A_413_49#_c_440_n N_Y_c_1009_n 0.0068091f $X=10.375 $Y=1.665 $X2=0
+ $Y2=0
cc_498 N_A_413_49#_c_447_n N_Y_c_1009_n 0.0300917f $X=10.375 $Y=1.51 $X2=0 $Y2=0
cc_499 N_A_413_49#_c_448_n N_Y_c_1009_n 0.0308284f $X=11.02 $Y=1.51 $X2=0 $Y2=0
cc_500 N_A_413_49#_M1000_g N_Y_c_1018_n 0.00297851f $X=4.57 $Y=2.465 $X2=0 $Y2=0
cc_501 N_A_413_49#_M1007_g N_Y_c_1018_n 0.00770847f $X=5 $Y=2.465 $X2=0 $Y2=0
cc_502 N_A_413_49#_M1009_g N_Y_c_1018_n 0.00770847f $X=5.43 $Y=2.465 $X2=0 $Y2=0
cc_503 N_A_413_49#_M1012_g N_Y_c_1018_n 0.00770847f $X=5.86 $Y=2.465 $X2=0 $Y2=0
cc_504 N_A_413_49#_M1015_g N_Y_c_1018_n 0.00770847f $X=6.29 $Y=2.465 $X2=0 $Y2=0
cc_505 N_A_413_49#_M1019_g N_Y_c_1018_n 0.00770847f $X=6.72 $Y=2.465 $X2=0 $Y2=0
cc_506 N_A_413_49#_M1024_g N_Y_c_1018_n 0.00770847f $X=7.15 $Y=2.465 $X2=0 $Y2=0
cc_507 N_A_413_49#_M1025_g N_Y_c_1018_n 0.00770847f $X=7.58 $Y=2.465 $X2=0 $Y2=0
cc_508 N_A_413_49#_M1027_g N_Y_c_1018_n 0.00770847f $X=8.01 $Y=2.465 $X2=0 $Y2=0
cc_509 N_A_413_49#_M1028_g N_Y_c_1018_n 0.00770847f $X=8.44 $Y=2.465 $X2=0 $Y2=0
cc_510 N_A_413_49#_M1029_g N_Y_c_1018_n 0.00770847f $X=8.87 $Y=2.465 $X2=0 $Y2=0
cc_511 N_A_413_49#_M1034_g N_Y_c_1018_n 0.00770847f $X=9.3 $Y=2.465 $X2=0 $Y2=0
cc_512 N_A_413_49#_M1039_g N_Y_c_1018_n 0.00770847f $X=9.73 $Y=2.465 $X2=0 $Y2=0
cc_513 N_A_413_49#_M1043_g N_Y_c_1018_n 0.00770847f $X=10.16 $Y=2.465 $X2=0
+ $Y2=0
cc_514 N_A_413_49#_M1046_g N_Y_c_1018_n 0.0124653f $X=10.59 $Y=2.465 $X2=0 $Y2=0
cc_515 N_A_413_49#_M1047_g N_Y_c_1018_n 0.00307468f $X=11.02 $Y=2.465 $X2=0
+ $Y2=0
cc_516 N_A_413_49#_c_573_p N_Y_c_1018_n 0.00396634f $X=3.925 $Y=2.095 $X2=0
+ $Y2=0
cc_517 N_A_413_49#_c_440_n N_Y_c_1018_n 0.5714f $X=10.375 $Y=1.665 $X2=0 $Y2=0
cc_518 N_A_413_49#_c_441_n N_Y_c_1018_n 0.00167386f $X=5.215 $Y=1.51 $X2=0 $Y2=0
cc_519 N_A_413_49#_c_442_n N_Y_c_1018_n 0.00167386f $X=6.075 $Y=1.51 $X2=0 $Y2=0
cc_520 N_A_413_49#_c_443_n N_Y_c_1018_n 0.00167386f $X=6.935 $Y=1.51 $X2=0 $Y2=0
cc_521 N_A_413_49#_c_444_n N_Y_c_1018_n 0.00167386f $X=7.795 $Y=1.51 $X2=0 $Y2=0
cc_522 N_A_413_49#_c_445_n N_Y_c_1018_n 0.00167386f $X=8.655 $Y=1.51 $X2=0 $Y2=0
cc_523 N_A_413_49#_c_446_n N_Y_c_1018_n 0.00167386f $X=9.515 $Y=1.51 $X2=0 $Y2=0
cc_524 N_A_413_49#_c_447_n N_Y_c_1018_n 0.00167386f $X=10.375 $Y=1.51 $X2=0
+ $Y2=0
cc_525 N_A_413_49#_c_433_n N_VGND_M1005_d 0.00176461f $X=2.935 $Y=1.14 $X2=0
+ $Y2=0
cc_526 N_A_413_49#_c_435_n N_VGND_M1035_d 0.00176461f $X=3.795 $Y=1.14 $X2=0
+ $Y2=0
cc_527 N_A_413_49#_c_436_n N_VGND_M1041_d 0.00179671f $X=4.34 $Y=1.14 $X2=0
+ $Y2=0
cc_528 N_A_413_49#_c_433_n N_VGND_c_1190_n 0.0135055f $X=2.935 $Y=1.14 $X2=0
+ $Y2=0
cc_529 N_A_413_49#_c_435_n N_VGND_c_1191_n 0.0135055f $X=3.795 $Y=1.14 $X2=0
+ $Y2=0
cc_530 N_A_413_49#_M1002_g N_VGND_c_1192_n 0.00159325f $X=4.57 $Y=0.665 $X2=0
+ $Y2=0
cc_531 N_A_413_49#_c_436_n N_VGND_c_1192_n 0.0143318f $X=4.34 $Y=1.14 $X2=0
+ $Y2=0
cc_532 N_A_413_49#_M1003_g N_VGND_c_1193_n 0.00194012f $X=5 $Y=0.665 $X2=0 $Y2=0
cc_533 N_A_413_49#_M1011_g N_VGND_c_1193_n 0.00194012f $X=5.43 $Y=0.665 $X2=0
+ $Y2=0
cc_534 N_A_413_49#_c_440_n N_VGND_c_1193_n 0.00146999f $X=10.375 $Y=1.665 $X2=0
+ $Y2=0
cc_535 N_A_413_49#_c_441_n N_VGND_c_1193_n 0.0114862f $X=5.215 $Y=1.51 $X2=0
+ $Y2=0
cc_536 N_A_413_49#_c_448_n N_VGND_c_1193_n 7.49903e-19 $X=11.02 $Y=1.51 $X2=0
+ $Y2=0
cc_537 N_A_413_49#_M1011_g N_VGND_c_1194_n 0.00575161f $X=5.43 $Y=0.665 $X2=0
+ $Y2=0
cc_538 N_A_413_49#_M1013_g N_VGND_c_1194_n 0.00575161f $X=5.86 $Y=0.665 $X2=0
+ $Y2=0
cc_539 N_A_413_49#_M1013_g N_VGND_c_1195_n 0.00194012f $X=5.86 $Y=0.665 $X2=0
+ $Y2=0
cc_540 N_A_413_49#_M1014_g N_VGND_c_1195_n 0.00194012f $X=6.29 $Y=0.665 $X2=0
+ $Y2=0
cc_541 N_A_413_49#_c_440_n N_VGND_c_1195_n 0.00146999f $X=10.375 $Y=1.665 $X2=0
+ $Y2=0
cc_542 N_A_413_49#_c_442_n N_VGND_c_1195_n 0.0114862f $X=6.075 $Y=1.51 $X2=0
+ $Y2=0
cc_543 N_A_413_49#_c_448_n N_VGND_c_1195_n 7.49903e-19 $X=11.02 $Y=1.51 $X2=0
+ $Y2=0
cc_544 N_A_413_49#_M1016_g N_VGND_c_1196_n 0.00194012f $X=6.72 $Y=0.665 $X2=0
+ $Y2=0
cc_545 N_A_413_49#_M1021_g N_VGND_c_1196_n 0.00194012f $X=7.15 $Y=0.665 $X2=0
+ $Y2=0
cc_546 N_A_413_49#_c_440_n N_VGND_c_1196_n 0.00146999f $X=10.375 $Y=1.665 $X2=0
+ $Y2=0
cc_547 N_A_413_49#_c_443_n N_VGND_c_1196_n 0.0114862f $X=6.935 $Y=1.51 $X2=0
+ $Y2=0
cc_548 N_A_413_49#_c_448_n N_VGND_c_1196_n 7.49903e-19 $X=11.02 $Y=1.51 $X2=0
+ $Y2=0
cc_549 N_A_413_49#_M1023_g N_VGND_c_1197_n 0.00194012f $X=7.58 $Y=0.665 $X2=0
+ $Y2=0
cc_550 N_A_413_49#_M1030_g N_VGND_c_1197_n 0.00194012f $X=8.01 $Y=0.665 $X2=0
+ $Y2=0
cc_551 N_A_413_49#_c_440_n N_VGND_c_1197_n 0.00146999f $X=10.375 $Y=1.665 $X2=0
+ $Y2=0
cc_552 N_A_413_49#_c_444_n N_VGND_c_1197_n 0.0114862f $X=7.795 $Y=1.51 $X2=0
+ $Y2=0
cc_553 N_A_413_49#_c_448_n N_VGND_c_1197_n 7.49903e-19 $X=11.02 $Y=1.51 $X2=0
+ $Y2=0
cc_554 N_A_413_49#_M1031_g N_VGND_c_1198_n 0.00194012f $X=8.44 $Y=0.665 $X2=0
+ $Y2=0
cc_555 N_A_413_49#_M1032_g N_VGND_c_1198_n 0.00194012f $X=8.87 $Y=0.665 $X2=0
+ $Y2=0
cc_556 N_A_413_49#_c_440_n N_VGND_c_1198_n 0.00146999f $X=10.375 $Y=1.665 $X2=0
+ $Y2=0
cc_557 N_A_413_49#_c_445_n N_VGND_c_1198_n 0.0114862f $X=8.655 $Y=1.51 $X2=0
+ $Y2=0
cc_558 N_A_413_49#_c_448_n N_VGND_c_1198_n 7.49903e-19 $X=11.02 $Y=1.51 $X2=0
+ $Y2=0
cc_559 N_A_413_49#_M1036_g N_VGND_c_1199_n 0.00194012f $X=9.3 $Y=0.665 $X2=0
+ $Y2=0
cc_560 N_A_413_49#_M1038_g N_VGND_c_1199_n 0.00194012f $X=9.73 $Y=0.665 $X2=0
+ $Y2=0
cc_561 N_A_413_49#_c_440_n N_VGND_c_1199_n 0.00146999f $X=10.375 $Y=1.665 $X2=0
+ $Y2=0
cc_562 N_A_413_49#_c_446_n N_VGND_c_1199_n 0.0114862f $X=9.515 $Y=1.51 $X2=0
+ $Y2=0
cc_563 N_A_413_49#_c_448_n N_VGND_c_1199_n 7.49903e-19 $X=11.02 $Y=1.51 $X2=0
+ $Y2=0
cc_564 N_A_413_49#_M1038_g N_VGND_c_1200_n 0.00575161f $X=9.73 $Y=0.665 $X2=0
+ $Y2=0
cc_565 N_A_413_49#_M1044_g N_VGND_c_1200_n 0.00575161f $X=10.16 $Y=0.665 $X2=0
+ $Y2=0
cc_566 N_A_413_49#_M1044_g N_VGND_c_1201_n 0.00194012f $X=10.16 $Y=0.665 $X2=0
+ $Y2=0
cc_567 N_A_413_49#_M1045_g N_VGND_c_1201_n 0.00194012f $X=10.59 $Y=0.665 $X2=0
+ $Y2=0
cc_568 N_A_413_49#_c_440_n N_VGND_c_1201_n 0.00146999f $X=10.375 $Y=1.665 $X2=0
+ $Y2=0
cc_569 N_A_413_49#_c_447_n N_VGND_c_1201_n 0.0114862f $X=10.375 $Y=1.51 $X2=0
+ $Y2=0
cc_570 N_A_413_49#_c_448_n N_VGND_c_1201_n 7.49903e-19 $X=11.02 $Y=1.51 $X2=0
+ $Y2=0
cc_571 N_A_413_49#_M1048_g N_VGND_c_1203_n 0.00490597f $X=11.02 $Y=0.665 $X2=0
+ $Y2=0
cc_572 N_A_413_49#_c_746_p N_VGND_c_1206_n 0.0108254f $X=3.065 $Y=0.48 $X2=0
+ $Y2=0
cc_573 N_A_413_49#_c_747_p N_VGND_c_1208_n 0.0108254f $X=3.925 $Y=0.48 $X2=0
+ $Y2=0
cc_574 N_A_413_49#_M1002_g N_VGND_c_1210_n 0.00575161f $X=4.57 $Y=0.665 $X2=0
+ $Y2=0
cc_575 N_A_413_49#_M1003_g N_VGND_c_1210_n 0.00575161f $X=5 $Y=0.665 $X2=0 $Y2=0
cc_576 N_A_413_49#_M1021_g N_VGND_c_1212_n 0.00575161f $X=7.15 $Y=0.665 $X2=0
+ $Y2=0
cc_577 N_A_413_49#_M1023_g N_VGND_c_1212_n 0.00575161f $X=7.58 $Y=0.665 $X2=0
+ $Y2=0
cc_578 N_A_413_49#_M1030_g N_VGND_c_1214_n 0.00575161f $X=8.01 $Y=0.665 $X2=0
+ $Y2=0
cc_579 N_A_413_49#_M1031_g N_VGND_c_1214_n 0.00575161f $X=8.44 $Y=0.665 $X2=0
+ $Y2=0
cc_580 N_A_413_49#_M1032_g N_VGND_c_1216_n 0.00575161f $X=8.87 $Y=0.665 $X2=0
+ $Y2=0
cc_581 N_A_413_49#_M1036_g N_VGND_c_1216_n 0.00575161f $X=9.3 $Y=0.665 $X2=0
+ $Y2=0
cc_582 N_A_413_49#_c_756_p N_VGND_c_1218_n 0.0104304f $X=2.205 $Y=0.48 $X2=0
+ $Y2=0
cc_583 N_A_413_49#_M1014_g N_VGND_c_1219_n 0.00575161f $X=6.29 $Y=0.665 $X2=0
+ $Y2=0
cc_584 N_A_413_49#_M1016_g N_VGND_c_1219_n 0.00575161f $X=6.72 $Y=0.665 $X2=0
+ $Y2=0
cc_585 N_A_413_49#_M1045_g N_VGND_c_1220_n 0.00575161f $X=10.59 $Y=0.665 $X2=0
+ $Y2=0
cc_586 N_A_413_49#_M1048_g N_VGND_c_1220_n 0.00575161f $X=11.02 $Y=0.665 $X2=0
+ $Y2=0
cc_587 N_A_413_49#_M1001_s N_VGND_c_1226_n 0.00357483f $X=2.065 $Y=0.245 $X2=0
+ $Y2=0
cc_588 N_A_413_49#_M1020_s N_VGND_c_1226_n 0.00305524f $X=2.925 $Y=0.245 $X2=0
+ $Y2=0
cc_589 N_A_413_49#_M1037_s N_VGND_c_1226_n 0.00305524f $X=3.785 $Y=0.245 $X2=0
+ $Y2=0
cc_590 N_A_413_49#_M1002_g N_VGND_c_1226_n 0.0106069f $X=4.57 $Y=0.665 $X2=0
+ $Y2=0
cc_591 N_A_413_49#_M1003_g N_VGND_c_1226_n 0.0106277f $X=5 $Y=0.665 $X2=0 $Y2=0
cc_592 N_A_413_49#_M1011_g N_VGND_c_1226_n 0.0106277f $X=5.43 $Y=0.665 $X2=0
+ $Y2=0
cc_593 N_A_413_49#_M1013_g N_VGND_c_1226_n 0.0106277f $X=5.86 $Y=0.665 $X2=0
+ $Y2=0
cc_594 N_A_413_49#_M1014_g N_VGND_c_1226_n 0.0106277f $X=6.29 $Y=0.665 $X2=0
+ $Y2=0
cc_595 N_A_413_49#_M1016_g N_VGND_c_1226_n 0.0106277f $X=6.72 $Y=0.665 $X2=0
+ $Y2=0
cc_596 N_A_413_49#_M1021_g N_VGND_c_1226_n 0.0106277f $X=7.15 $Y=0.665 $X2=0
+ $Y2=0
cc_597 N_A_413_49#_M1023_g N_VGND_c_1226_n 0.0106277f $X=7.58 $Y=0.665 $X2=0
+ $Y2=0
cc_598 N_A_413_49#_M1030_g N_VGND_c_1226_n 0.0106277f $X=8.01 $Y=0.665 $X2=0
+ $Y2=0
cc_599 N_A_413_49#_M1031_g N_VGND_c_1226_n 0.0106277f $X=8.44 $Y=0.665 $X2=0
+ $Y2=0
cc_600 N_A_413_49#_M1032_g N_VGND_c_1226_n 0.0106277f $X=8.87 $Y=0.665 $X2=0
+ $Y2=0
cc_601 N_A_413_49#_M1036_g N_VGND_c_1226_n 0.0106277f $X=9.3 $Y=0.665 $X2=0
+ $Y2=0
cc_602 N_A_413_49#_M1038_g N_VGND_c_1226_n 0.0106277f $X=9.73 $Y=0.665 $X2=0
+ $Y2=0
cc_603 N_A_413_49#_M1044_g N_VGND_c_1226_n 0.0106277f $X=10.16 $Y=0.665 $X2=0
+ $Y2=0
cc_604 N_A_413_49#_M1045_g N_VGND_c_1226_n 0.0106277f $X=10.59 $Y=0.665 $X2=0
+ $Y2=0
cc_605 N_A_413_49#_M1048_g N_VGND_c_1226_n 0.0115831f $X=11.02 $Y=0.665 $X2=0
+ $Y2=0
cc_606 N_A_413_49#_c_756_p N_VGND_c_1226_n 0.00915916f $X=2.205 $Y=0.48 $X2=0
+ $Y2=0
cc_607 N_A_413_49#_c_746_p N_VGND_c_1226_n 0.00972454f $X=3.065 $Y=0.48 $X2=0
+ $Y2=0
cc_608 N_A_413_49#_c_747_p N_VGND_c_1226_n 0.00972454f $X=3.925 $Y=0.48 $X2=0
+ $Y2=0
cc_609 N_VPWR_c_783_n N_Y_M1000_d 0.00425874f $X=11.28 $Y=3.33 $X2=0 $Y2=0
cc_610 N_VPWR_c_783_n N_Y_M1009_d 0.00304497f $X=11.28 $Y=3.33 $X2=0 $Y2=0
cc_611 N_VPWR_c_783_n N_Y_M1015_d 0.00304497f $X=11.28 $Y=3.33 $X2=0 $Y2=0
cc_612 N_VPWR_c_783_n N_Y_M1024_d 0.00304497f $X=11.28 $Y=3.33 $X2=0 $Y2=0
cc_613 N_VPWR_c_783_n N_Y_M1027_d 0.00304497f $X=11.28 $Y=3.33 $X2=0 $Y2=0
cc_614 N_VPWR_c_783_n N_Y_M1029_d 0.00304497f $X=11.28 $Y=3.33 $X2=0 $Y2=0
cc_615 N_VPWR_c_783_n N_Y_M1039_d 0.00304497f $X=11.28 $Y=3.33 $X2=0 $Y2=0
cc_616 N_VPWR_c_783_n N_Y_M1046_d 0.00304497f $X=11.28 $Y=3.33 $X2=0 $Y2=0
cc_617 N_VPWR_c_790_n N_Y_c_1002_n 0.00695484f $X=5.215 $Y=2.12 $X2=0 $Y2=0
cc_618 N_VPWR_c_807_n N_Y_c_1002_n 0.0103851f $X=5.085 $Y=3.33 $X2=0 $Y2=0
cc_619 N_VPWR_c_783_n N_Y_c_1002_n 0.00845197f $X=11.28 $Y=3.33 $X2=0 $Y2=0
cc_620 N_VPWR_c_790_n N_Y_c_1003_n 0.00697067f $X=5.215 $Y=2.12 $X2=0 $Y2=0
cc_621 N_VPWR_c_791_n N_Y_c_1003_n 0.0113476f $X=5.945 $Y=3.33 $X2=0 $Y2=0
cc_622 N_VPWR_c_792_n N_Y_c_1003_n 0.00697067f $X=6.075 $Y=2.12 $X2=0 $Y2=0
cc_623 N_VPWR_c_783_n N_Y_c_1003_n 0.00977851f $X=11.28 $Y=3.33 $X2=0 $Y2=0
cc_624 N_VPWR_c_792_n N_Y_c_1004_n 0.00697067f $X=6.075 $Y=2.12 $X2=0 $Y2=0
cc_625 N_VPWR_c_793_n N_Y_c_1004_n 0.00697067f $X=6.935 $Y=2.12 $X2=0 $Y2=0
cc_626 N_VPWR_c_816_n N_Y_c_1004_n 0.0113476f $X=6.805 $Y=3.33 $X2=0 $Y2=0
cc_627 N_VPWR_c_783_n N_Y_c_1004_n 0.00977851f $X=11.28 $Y=3.33 $X2=0 $Y2=0
cc_628 N_VPWR_c_793_n N_Y_c_1005_n 0.00697067f $X=6.935 $Y=2.12 $X2=0 $Y2=0
cc_629 N_VPWR_c_794_n N_Y_c_1005_n 0.00697067f $X=7.795 $Y=2.12 $X2=0 $Y2=0
cc_630 N_VPWR_c_809_n N_Y_c_1005_n 0.0113476f $X=7.665 $Y=3.33 $X2=0 $Y2=0
cc_631 N_VPWR_c_783_n N_Y_c_1005_n 0.00977851f $X=11.28 $Y=3.33 $X2=0 $Y2=0
cc_632 N_VPWR_c_794_n N_Y_c_1006_n 0.00697067f $X=7.795 $Y=2.12 $X2=0 $Y2=0
cc_633 N_VPWR_c_795_n N_Y_c_1006_n 0.00697067f $X=8.655 $Y=2.12 $X2=0 $Y2=0
cc_634 N_VPWR_c_811_n N_Y_c_1006_n 0.0113476f $X=8.525 $Y=3.33 $X2=0 $Y2=0
cc_635 N_VPWR_c_783_n N_Y_c_1006_n 0.00977851f $X=11.28 $Y=3.33 $X2=0 $Y2=0
cc_636 N_VPWR_c_795_n N_Y_c_1007_n 0.00697067f $X=8.655 $Y=2.12 $X2=0 $Y2=0
cc_637 N_VPWR_c_796_n N_Y_c_1007_n 0.00697067f $X=9.515 $Y=2.12 $X2=0 $Y2=0
cc_638 N_VPWR_c_813_n N_Y_c_1007_n 0.0113476f $X=9.385 $Y=3.33 $X2=0 $Y2=0
cc_639 N_VPWR_c_783_n N_Y_c_1007_n 0.00977851f $X=11.28 $Y=3.33 $X2=0 $Y2=0
cc_640 N_VPWR_c_796_n N_Y_c_1008_n 0.00697067f $X=9.515 $Y=2.12 $X2=0 $Y2=0
cc_641 N_VPWR_c_797_n N_Y_c_1008_n 0.0113476f $X=10.245 $Y=3.33 $X2=0 $Y2=0
cc_642 N_VPWR_c_798_n N_Y_c_1008_n 0.00697067f $X=10.375 $Y=2.12 $X2=0 $Y2=0
cc_643 N_VPWR_c_783_n N_Y_c_1008_n 0.00977851f $X=11.28 $Y=3.33 $X2=0 $Y2=0
cc_644 N_VPWR_c_798_n N_Y_c_1009_n 0.00697067f $X=10.375 $Y=2.12 $X2=0 $Y2=0
cc_645 N_VPWR_c_817_n N_Y_c_1009_n 0.0113476f $X=11.105 $Y=3.33 $X2=0 $Y2=0
cc_646 N_VPWR_c_783_n N_Y_c_1009_n 0.00977851f $X=11.28 $Y=3.33 $X2=0 $Y2=0
cc_647 N_VPWR_M1007_s N_Y_c_1018_n 0.00191566f $X=5.075 $Y=1.835 $X2=0 $Y2=0
cc_648 N_VPWR_M1012_s N_Y_c_1018_n 0.00191566f $X=5.935 $Y=1.835 $X2=0 $Y2=0
cc_649 N_VPWR_M1019_s N_Y_c_1018_n 0.00191566f $X=6.795 $Y=1.835 $X2=0 $Y2=0
cc_650 N_VPWR_M1025_s N_Y_c_1018_n 0.00191566f $X=7.655 $Y=1.835 $X2=0 $Y2=0
cc_651 N_VPWR_M1028_s N_Y_c_1018_n 0.00191566f $X=8.515 $Y=1.835 $X2=0 $Y2=0
cc_652 N_VPWR_M1034_s N_Y_c_1018_n 0.00191566f $X=9.375 $Y=1.835 $X2=0 $Y2=0
cc_653 N_VPWR_M1043_s N_Y_c_1018_n 0.00191566f $X=10.235 $Y=1.835 $X2=0 $Y2=0
cc_654 N_VPWR_c_789_n N_Y_c_1018_n 0.00137712f $X=4.355 $Y=2.27 $X2=0 $Y2=0
cc_655 N_VPWR_c_790_n N_Y_c_1018_n 0.0245913f $X=5.215 $Y=2.12 $X2=0 $Y2=0
cc_656 N_VPWR_c_792_n N_Y_c_1018_n 0.0245913f $X=6.075 $Y=2.12 $X2=0 $Y2=0
cc_657 N_VPWR_c_793_n N_Y_c_1018_n 0.0245913f $X=6.935 $Y=2.12 $X2=0 $Y2=0
cc_658 N_VPWR_c_794_n N_Y_c_1018_n 0.0245913f $X=7.795 $Y=2.12 $X2=0 $Y2=0
cc_659 N_VPWR_c_795_n N_Y_c_1018_n 0.0245913f $X=8.655 $Y=2.12 $X2=0 $Y2=0
cc_660 N_VPWR_c_796_n N_Y_c_1018_n 0.0245913f $X=9.515 $Y=2.12 $X2=0 $Y2=0
cc_661 N_VPWR_c_798_n N_Y_c_1018_n 0.0245913f $X=10.375 $Y=2.12 $X2=0 $Y2=0
cc_662 N_VPWR_c_800_n N_Y_c_1018_n 0.00586406f $X=11.235 $Y=2.12 $X2=0 $Y2=0
cc_663 N_Y_c_1003_n N_VGND_c_1194_n 0.0108254f $X=5.645 $Y=0.48 $X2=0 $Y2=0
cc_664 N_Y_c_1008_n N_VGND_c_1200_n 0.0108254f $X=9.945 $Y=0.48 $X2=0 $Y2=0
cc_665 N_Y_c_1002_n N_VGND_c_1210_n 0.00990367f $X=4.785 $Y=0.48 $X2=0 $Y2=0
cc_666 N_Y_c_1005_n N_VGND_c_1212_n 0.0108254f $X=7.365 $Y=0.48 $X2=0 $Y2=0
cc_667 N_Y_c_1006_n N_VGND_c_1214_n 0.0108254f $X=8.225 $Y=0.48 $X2=0 $Y2=0
cc_668 N_Y_c_1007_n N_VGND_c_1216_n 0.0108254f $X=9.085 $Y=0.48 $X2=0 $Y2=0
cc_669 N_Y_c_1004_n N_VGND_c_1219_n 0.0108254f $X=6.505 $Y=0.48 $X2=0 $Y2=0
cc_670 N_Y_c_1009_n N_VGND_c_1220_n 0.0108254f $X=10.805 $Y=0.48 $X2=0 $Y2=0
cc_671 N_Y_M1002_s N_VGND_c_1226_n 0.00426761f $X=4.645 $Y=0.245 $X2=0 $Y2=0
cc_672 N_Y_M1011_s N_VGND_c_1226_n 0.00305524f $X=5.505 $Y=0.245 $X2=0 $Y2=0
cc_673 N_Y_M1014_s N_VGND_c_1226_n 0.00305524f $X=6.365 $Y=0.245 $X2=0 $Y2=0
cc_674 N_Y_M1021_s N_VGND_c_1226_n 0.00305524f $X=7.225 $Y=0.245 $X2=0 $Y2=0
cc_675 N_Y_M1030_s N_VGND_c_1226_n 0.00305524f $X=8.085 $Y=0.245 $X2=0 $Y2=0
cc_676 N_Y_M1032_s N_VGND_c_1226_n 0.00305524f $X=8.945 $Y=0.245 $X2=0 $Y2=0
cc_677 N_Y_M1038_s N_VGND_c_1226_n 0.00305524f $X=9.805 $Y=0.245 $X2=0 $Y2=0
cc_678 N_Y_M1045_s N_VGND_c_1226_n 0.00305524f $X=10.665 $Y=0.245 $X2=0 $Y2=0
cc_679 N_Y_c_1002_n N_VGND_c_1226_n 0.00840532f $X=4.785 $Y=0.48 $X2=0 $Y2=0
cc_680 N_Y_c_1003_n N_VGND_c_1226_n 0.00972454f $X=5.645 $Y=0.48 $X2=0 $Y2=0
cc_681 N_Y_c_1004_n N_VGND_c_1226_n 0.00972454f $X=6.505 $Y=0.48 $X2=0 $Y2=0
cc_682 N_Y_c_1005_n N_VGND_c_1226_n 0.00972454f $X=7.365 $Y=0.48 $X2=0 $Y2=0
cc_683 N_Y_c_1006_n N_VGND_c_1226_n 0.00972454f $X=8.225 $Y=0.48 $X2=0 $Y2=0
cc_684 N_Y_c_1007_n N_VGND_c_1226_n 0.00972454f $X=9.085 $Y=0.48 $X2=0 $Y2=0
cc_685 N_Y_c_1008_n N_VGND_c_1226_n 0.00972454f $X=9.945 $Y=0.48 $X2=0 $Y2=0
cc_686 N_Y_c_1009_n N_VGND_c_1226_n 0.00972454f $X=10.805 $Y=0.48 $X2=0 $Y2=0
