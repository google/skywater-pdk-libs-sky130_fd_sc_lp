* NGSPICE file created from sky130_fd_sc_lp__a221o_4.ext - technology: sky130A

.subckt sky130_fd_sc_lp__a221o_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
M1000 a_457_47# A2 VGND VNB nshort w=840000u l=150000u
+  ad=4.704e+11p pd=4.48e+06u as=1.386e+12p ps=1.338e+07u
M1001 VGND C1 a_83_21# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=9.156e+11p ps=8.9e+06u
M1002 a_457_367# A2 VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=1.4112e+12p pd=1.232e+07u as=1.7262e+12p ps=1.534e+07u
M1003 X a_83_21# VGND VNB nshort w=840000u l=150000u
+  ad=4.704e+11p pd=4.48e+06u as=0p ps=0u
M1004 a_457_367# B1 a_822_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=1.3734e+12p ps=1.226e+07u
M1005 a_83_21# B1 a_1077_47# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=6.804e+11p ps=6.66e+06u
M1006 VGND B2 a_1077_47# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR a_83_21# X VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=7.056e+11p ps=6.16e+06u
M1008 VPWR a_83_21# X VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND A2 a_457_47# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_457_367# B2 a_822_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_83_21# C1 VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VGND a_83_21# X VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_457_47# A1 a_83_21# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 X a_83_21# VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VPWR A1 a_457_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_822_367# C1 a_83_21# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=3.528e+11p ps=3.08e+06u
M1017 VPWR A2 a_457_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 X a_83_21# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_822_367# B1 a_457_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_83_21# A1 a_457_47# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VGND a_83_21# X VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_1077_47# B2 VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 X a_83_21# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_1077_47# B1 a_83_21# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_457_367# A1 VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_83_21# C1 a_822_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_822_367# B2 a_457_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

