* File: sky130_fd_sc_lp__or3_0.pex.spice
* Created: Wed Sep  2 10:30:20 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__OR3_0%C 3 9 11 12 13 14 15 20
r37 20 22 45.5639 $w=3.95e-07 $l=1.65e-07 $layer=POLY_cond $X=0.607 $Y=1.245
+ $X2=0.607 $Y2=1.08
r38 14 15 15.6137 $w=3.08e-07 $l=4.2e-07 $layer=LI1_cond $X=0.71 $Y=1.245
+ $X2=0.71 $Y2=1.665
r39 14 20 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.64
+ $Y=1.245 $X2=0.64 $Y2=1.245
r40 13 14 11.8962 $w=3.08e-07 $l=3.2e-07 $layer=LI1_cond $X=0.71 $Y=0.925
+ $X2=0.71 $Y2=1.245
r41 11 12 43.452 $w=3.95e-07 $l=1.5e-07 $layer=POLY_cond $X=0.682 $Y=1.715
+ $X2=0.682 $Y2=1.865
r42 9 12 384.574 $w=1.5e-07 $l=7.5e-07 $layer=POLY_cond $X=0.88 $Y=2.615
+ $X2=0.88 $Y2=1.865
r43 5 20 4.50555 $w=3.95e-07 $l=3.2e-08 $layer=POLY_cond $X=0.607 $Y=1.277
+ $X2=0.607 $Y2=1.245
r44 5 11 61.6697 $w=3.95e-07 $l=4.38e-07 $layer=POLY_cond $X=0.607 $Y=1.277
+ $X2=0.607 $Y2=1.715
r45 3 22 305.096 $w=1.5e-07 $l=5.95e-07 $layer=POLY_cond $X=0.485 $Y=0.485
+ $X2=0.485 $Y2=1.08
.ends

.subckt PM_SKY130_FD_SC_LP__OR3_0%B 3 7 9 10 11 12 13 20 25
c58 13 0 1.57783e-19 $X=1.2 $Y=1.665
r59 23 25 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.18 $Y=1.31
+ $X2=1.18 $Y2=1.475
r60 20 23 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.18 $Y=0.97
+ $X2=1.18 $Y2=1.31
r61 12 37 4.58814 $w=3.18e-07 $l=1.17e-07 $layer=LI1_cond $X=1.195 $Y=1.252
+ $X2=1.195 $Y2=1.135
r62 12 13 13.3251 $w=3.18e-07 $l=3.7e-07 $layer=LI1_cond $X=1.195 $Y=1.295
+ $X2=1.195 $Y2=1.665
r63 12 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.18
+ $Y=1.31 $X2=1.18 $Y2=1.31
r64 11 37 9.13257 $w=2.63e-07 $l=2.1e-07 $layer=LI1_cond $X=1.167 $Y=0.925
+ $X2=1.167 $Y2=1.135
r65 11 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.18
+ $Y=0.97 $X2=1.18 $Y2=0.97
r66 10 20 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=1.18 $Y=0.955
+ $X2=1.18 $Y2=0.97
r67 9 10 43.5886 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=1.237 $Y=0.805
+ $X2=1.237 $Y2=0.955
r68 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.385 $Y=0.485
+ $X2=1.385 $Y2=0.805
r69 3 25 584.553 $w=1.5e-07 $l=1.14e-06 $layer=POLY_cond $X=1.24 $Y=2.615
+ $X2=1.24 $Y2=1.475
.ends

.subckt PM_SKY130_FD_SC_LP__OR3_0%A 3 7 10 11 14 15 19
c51 11 0 1.77888e-19 $X=1.72 $Y=1.865
r52 14 15 13.755 $w=3.08e-07 $l=3.7e-07 $layer=LI1_cond $X=1.68 $Y=1.295
+ $X2=1.68 $Y2=1.665
r53 14 19 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.75
+ $Y=1.36 $X2=1.75 $Y2=1.36
r54 13 19 42.4377 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.75 $Y=1.195
+ $X2=1.75 $Y2=1.36
r55 10 19 56.8299 $w=3.3e-07 $l=3.25e-07 $layer=POLY_cond $X=1.75 $Y=1.685
+ $X2=1.75 $Y2=1.36
r56 10 11 48.8344 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=1.72 $Y=1.685
+ $X2=1.72 $Y2=1.865
r57 7 13 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=1.815 $Y=0.485
+ $X2=1.815 $Y2=1.195
r58 3 11 384.574 $w=1.5e-07 $l=7.5e-07 $layer=POLY_cond $X=1.6 $Y=2.615 $X2=1.6
+ $Y2=1.865
.ends

.subckt PM_SKY130_FD_SC_LP__OR3_0%A_29_55# 1 2 3 12 16 20 21 24 28 30 34 36 37
+ 41 45 47 48 49
c86 37 0 1.77888e-19 $X=1.73 $Y=0.912
c87 24 0 1.57783e-19 $X=0.27 $Y=0.485
r88 47 49 8.51103 $w=3.58e-07 $l=1.65e-07 $layer=LI1_cond $X=2.195 $Y=1.71
+ $X2=2.195 $Y2=1.545
r89 47 48 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.29
+ $Y=1.71 $X2=2.29 $Y2=1.71
r90 44 45 8.15436 $w=3.03e-07 $l=1.65e-07 $layer=LI1_cond $X=0.665 $Y=2.187
+ $X2=0.83 $Y2=2.187
r91 40 47 0.480185 $w=3.58e-07 $l=1.5e-08 $layer=LI1_cond $X=2.195 $Y=1.725
+ $X2=2.195 $Y2=1.71
r92 40 41 9.92381 $w=3.58e-07 $l=3.1e-07 $layer=LI1_cond $X=2.195 $Y=1.725
+ $X2=2.195 $Y2=2.035
r93 38 49 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=2.1 $Y=1.005 $X2=2.1
+ $Y2=1.545
r94 36 38 6.83233 $w=1.85e-07 $l=1.28662e-07 $layer=LI1_cond $X=2.015 $Y=0.912
+ $X2=2.1 $Y2=1.005
r95 36 37 17.086 $w=1.83e-07 $l=2.85e-07 $layer=LI1_cond $X=2.015 $Y=0.912
+ $X2=1.73 $Y2=0.912
r96 32 37 7.07139 $w=1.85e-07 $l=1.69882e-07 $layer=LI1_cond $X=1.6 $Y=0.82
+ $X2=1.73 $Y2=0.912
r97 32 34 14.8488 $w=2.58e-07 $l=3.35e-07 $layer=LI1_cond $X=1.6 $Y=0.82 $X2=1.6
+ $Y2=0.485
r98 30 41 7.85115 $w=1.8e-07 $l=2.20454e-07 $layer=LI1_cond $X=2.015 $Y=2.125
+ $X2=2.195 $Y2=2.035
r99 30 45 73.0152 $w=1.78e-07 $l=1.185e-06 $layer=LI1_cond $X=2.015 $Y=2.125
+ $X2=0.83 $Y2=2.125
r100 26 44 0.230243 $w=3.3e-07 $l=1.53e-07 $layer=LI1_cond $X=0.665 $Y=2.34
+ $X2=0.665 $Y2=2.187
r101 26 28 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=0.665 $Y=2.34
+ $X2=0.665 $Y2=2.615
r102 22 44 15.8697 $w=3.03e-07 $l=4.2e-07 $layer=LI1_cond $X=0.245 $Y=2.187
+ $X2=0.665 $Y2=2.187
r103 22 24 63.796 $w=2.78e-07 $l=1.55e-06 $layer=LI1_cond $X=0.245 $Y=2.035
+ $X2=0.245 $Y2=0.485
r104 20 48 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.29 $Y=2.05
+ $X2=2.29 $Y2=1.71
r105 20 21 44.4756 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.29 $Y=2.05
+ $X2=2.29 $Y2=2.215
r106 19 48 40.425 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.29 $Y=1.545
+ $X2=2.29 $Y2=1.71
r107 16 21 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=2.37 $Y=2.725
+ $X2=2.37 $Y2=2.215
r108 12 19 543.532 $w=1.5e-07 $l=1.06e-06 $layer=POLY_cond $X=2.245 $Y=0.485
+ $X2=2.245 $Y2=1.545
r109 3 28 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=0.54
+ $Y=2.405 $X2=0.665 $Y2=2.615
r110 2 34 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.46
+ $Y=0.275 $X2=1.6 $Y2=0.485
r111 1 24 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.145
+ $Y=0.275 $X2=0.27 $Y2=0.485
.ends

.subckt PM_SKY130_FD_SC_LP__OR3_0%VPWR 1 6 8 10 17 18 21
r24 22 24 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r25 21 24 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r26 21 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r27 18 22 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r28 17 18 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r29 15 21 12.3804 $w=1.7e-07 $l=2.93e-07 $layer=LI1_cond $X=2.25 $Y=3.33
+ $X2=1.957 $Y2=3.33
r30 15 17 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=2.25 $Y=3.33
+ $X2=2.64 $Y2=3.33
r31 12 13 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r32 10 21 12.3804 $w=1.7e-07 $l=2.92e-07 $layer=LI1_cond $X=1.665 $Y=3.33
+ $X2=1.957 $Y2=3.33
r33 10 12 92.9679 $w=1.68e-07 $l=1.425e-06 $layer=LI1_cond $X=1.665 $Y=3.33
+ $X2=0.24 $Y2=3.33
r34 8 24 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=1.68 $Y2=3.33
r35 8 13 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=0.24 $Y2=3.33
r36 4 21 2.46141 $w=5.85e-07 $l=8.5e-08 $layer=LI1_cond $X=1.957 $Y=3.245
+ $X2=1.957 $Y2=3.33
r37 4 6 14.2098 $w=5.83e-07 $l=6.95e-07 $layer=LI1_cond $X=1.957 $Y=3.245
+ $X2=1.957 $Y2=2.55
r38 1 6 200 $w=1.7e-07 $l=5.47723e-07 $layer=licon1_PDIFF $count=3 $X=1.675
+ $Y=2.405 $X2=2.155 $Y2=2.55
.ends

.subckt PM_SKY130_FD_SC_LP__OR3_0%X 1 2 7 8 9 10 11 12 13 42 45
r20 45 46 1.89813 $w=3.73e-07 $l=2e-08 $layer=LI1_cond $X=2.607 $Y=2.405
+ $X2=2.607 $Y2=2.385
r21 33 49 0.6761 $w=3.73e-07 $l=2.2e-08 $layer=LI1_cond $X=2.607 $Y=2.572
+ $X2=2.607 $Y2=2.55
r22 22 42 2.36532 $w=2.5e-07 $l=1.65e-07 $layer=LI1_cond $X=2.67 $Y=0.65
+ $X2=2.67 $Y2=0.485
r23 13 33 6.23856 $w=3.73e-07 $l=2.03e-07 $layer=LI1_cond $X=2.607 $Y=2.775
+ $X2=2.607 $Y2=2.572
r24 12 49 3.47269 $w=3.73e-07 $l=1.13e-07 $layer=LI1_cond $X=2.607 $Y=2.437
+ $X2=2.607 $Y2=2.55
r25 12 45 0.983418 $w=3.73e-07 $l=3.2e-08 $layer=LI1_cond $X=2.607 $Y=2.437
+ $X2=2.607 $Y2=2.405
r26 12 46 1.52122 $w=2.48e-07 $l=3.3e-08 $layer=LI1_cond $X=2.67 $Y=2.352
+ $X2=2.67 $Y2=2.385
r27 11 12 14.613 $w=2.48e-07 $l=3.17e-07 $layer=LI1_cond $X=2.67 $Y=2.035
+ $X2=2.67 $Y2=2.352
r28 10 11 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=2.67 $Y=1.665
+ $X2=2.67 $Y2=2.035
r29 9 10 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=2.67 $Y=1.295
+ $X2=2.67 $Y2=1.665
r30 8 9 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=2.67 $Y=0.925 $X2=2.67
+ $Y2=1.295
r31 8 22 12.6769 $w=2.48e-07 $l=2.75e-07 $layer=LI1_cond $X=2.67 $Y=0.925
+ $X2=2.67 $Y2=0.65
r32 7 42 1.04768 $w=3.28e-07 $l=3e-08 $layer=LI1_cond $X=2.64 $Y=0.485 $X2=2.67
+ $Y2=0.485
r33 7 38 4.88915 $w=3.28e-07 $l=1.4e-07 $layer=LI1_cond $X=2.64 $Y=0.485 $X2=2.5
+ $Y2=0.485
r34 2 49 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=2.445
+ $Y=2.405 $X2=2.585 $Y2=2.55
r35 1 38 182 $w=1.7e-07 $l=2.86182e-07 $layer=licon1_NDIFF $count=1 $X=2.32
+ $Y=0.275 $X2=2.5 $Y2=0.485
.ends

.subckt PM_SKY130_FD_SC_LP__OR3_0%VGND 1 2 9 12 13 14 26 27 32 38
r34 36 38 9.85322 $w=7.18e-07 $l=1e-07 $layer=LI1_cond $X=1.2 $Y=0.275 $X2=1.3
+ $Y2=0.275
r35 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r36 34 36 0.498366 $w=7.18e-07 $l=3e-08 $layer=LI1_cond $X=1.17 $Y=0.275 $X2=1.2
+ $Y2=0.275
r37 31 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r38 30 34 7.47549 $w=7.18e-07 $l=4.5e-07 $layer=LI1_cond $X=0.72 $Y=0.275
+ $X2=1.17 $Y2=0.275
r39 30 32 10.933 $w=7.18e-07 $l=1.65e-07 $layer=LI1_cond $X=0.72 $Y=0.275
+ $X2=0.555 $Y2=0.275
r40 30 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r41 26 27 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r42 24 27 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r43 23 38 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=1.68 $Y=0 $X2=1.3
+ $Y2=0
r44 23 24 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r45 19 31 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r46 18 32 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.24 $Y=0 $X2=0.555
+ $Y2=0
r47 18 19 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r48 14 24 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=1.68
+ $Y2=0
r49 14 37 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=1.2
+ $Y2=0
r50 12 23 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=1.9 $Y=0 $X2=1.68
+ $Y2=0
r51 12 13 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.9 $Y=0 $X2=2.03
+ $Y2=0
r52 11 26 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r53 11 13 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.16 $Y=0 $X2=2.03
+ $Y2=0
r54 7 13 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=2.03 $Y=0.085
+ $X2=2.03 $Y2=0
r55 7 9 17.7299 $w=2.58e-07 $l=4e-07 $layer=LI1_cond $X=2.03 $Y=0.085 $X2=2.03
+ $Y2=0.485
r56 2 9 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.89
+ $Y=0.275 $X2=2.03 $Y2=0.485
r57 1 34 91 $w=1.7e-07 $l=7.0075e-07 $layer=licon1_NDIFF $count=2 $X=0.56
+ $Y=0.275 $X2=1.17 $Y2=0.47
.ends

