* File: sky130_fd_sc_lp__sdlclkp_1.pex.spice
* Created: Wed Sep  2 10:37:03 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__SDLCLKP_1%SCE 3 7 9 10 12 13 14 15 16 17 24
c37 9 0 1.68929e-19 $X=0.437 $Y=0.875
r38 24 25 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.27
+ $Y=1.04 $X2=0.27 $Y2=1.04
r39 16 17 11.2212 $w=3.78e-07 $l=3.7e-07 $layer=LI1_cond $X=0.275 $Y=2.035
+ $X2=0.275 $Y2=2.405
r40 15 16 11.2212 $w=3.78e-07 $l=3.7e-07 $layer=LI1_cond $X=0.275 $Y=1.665
+ $X2=0.275 $Y2=2.035
r41 14 15 11.2212 $w=3.78e-07 $l=3.7e-07 $layer=LI1_cond $X=0.275 $Y=1.295
+ $X2=0.275 $Y2=1.665
r42 14 25 7.7335 $w=3.78e-07 $l=2.55e-07 $layer=LI1_cond $X=0.275 $Y=1.295
+ $X2=0.275 $Y2=1.04
r43 13 25 3.48766 $w=3.78e-07 $l=1.15e-07 $layer=LI1_cond $X=0.275 $Y=0.925
+ $X2=0.275 $Y2=1.04
r44 11 24 35.3689 $w=4.45e-07 $l=2.83e-07 $layer=POLY_cond $X=0.327 $Y=1.323
+ $X2=0.327 $Y2=1.04
r45 11 12 53.9265 $w=4.45e-07 $l=2.22e-07 $layer=POLY_cond $X=0.327 $Y=1.323
+ $X2=0.327 $Y2=1.545
r46 10 24 1.87468 $w=4.45e-07 $l=1.5e-08 $layer=POLY_cond $X=0.327 $Y=1.025
+ $X2=0.327 $Y2=1.04
r47 9 10 44.9281 $w=4.45e-07 $l=1.5e-07 $layer=POLY_cond $X=0.437 $Y=0.875
+ $X2=0.437 $Y2=1.025
r48 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.695 $Y=0.555
+ $X2=0.695 $Y2=0.875
r49 3 12 571.734 $w=1.5e-07 $l=1.115e-06 $layer=POLY_cond $X=0.475 $Y=2.66
+ $X2=0.475 $Y2=1.545
.ends

.subckt PM_SKY130_FD_SC_LP__SDLCLKP_1%GATE 3 7 11 14 15 16 17 22
c52 15 0 1.68929e-19 $X=1.2 $Y=0.925
r53 22 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.145
+ $Y=1.04 $X2=1.145 $Y2=1.04
r54 16 17 13.9805 $w=3.03e-07 $l=3.7e-07 $layer=LI1_cond $X=1.212 $Y=1.295
+ $X2=1.212 $Y2=1.665
r55 16 23 9.63518 $w=3.03e-07 $l=2.55e-07 $layer=LI1_cond $X=1.212 $Y=1.295
+ $X2=1.212 $Y2=1.04
r56 15 23 4.34528 $w=3.03e-07 $l=1.15e-07 $layer=LI1_cond $X=1.212 $Y=0.925
+ $X2=1.212 $Y2=1.04
r57 14 22 38.6168 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.145 $Y=0.875
+ $X2=1.145 $Y2=1.04
r58 11 22 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=1.145 $Y=1.395
+ $X2=1.145 $Y2=1.04
r59 8 11 158.957 $w=1.5e-07 $l=3.1e-07 $layer=POLY_cond $X=0.835 $Y=1.47
+ $X2=1.145 $Y2=1.47
r60 7 14 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.125 $Y=0.555
+ $X2=1.125 $Y2=0.875
r61 1 8 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.835 $Y=1.545
+ $X2=0.835 $Y2=1.47
r62 1 3 571.734 $w=1.5e-07 $l=1.115e-06 $layer=POLY_cond $X=0.835 $Y=1.545
+ $X2=0.835 $Y2=2.66
.ends

.subckt PM_SKY130_FD_SC_LP__SDLCLKP_1%A_334_69# 1 2 7 9 13 16 19 23 27 30 33 36
+ 38 39
c81 39 0 1.18174e-19 $X=2.535 $Y=1.72
c82 7 0 1.08032e-19 $X=3.325 $Y=1.66
r83 39 41 11.3858 $w=2.54e-07 $l=6e-08 $layer=POLY_cond $X=2.535 $Y=1.72
+ $X2=2.535 $Y2=1.66
r84 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.535
+ $Y=1.72 $X2=2.535 $Y2=1.72
r85 35 38 6.46067 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=2.35 $Y=1.72
+ $X2=2.535 $Y2=1.72
r86 35 36 6.00906 $w=3.28e-07 $l=1.25e-07 $layer=LI1_cond $X=2.35 $Y=1.72
+ $X2=2.225 $Y2=1.72
r87 31 35 2.36532 $w=2.5e-07 $l=1.65e-07 $layer=LI1_cond $X=2.35 $Y=1.885
+ $X2=2.35 $Y2=1.72
r88 31 33 14.0598 $w=2.48e-07 $l=3.05e-07 $layer=LI1_cond $X=2.35 $Y=1.885
+ $X2=2.35 $Y2=2.19
r89 30 36 13.5255 $w=2.03e-07 $l=2.5e-07 $layer=LI1_cond $X=1.975 $Y=1.657
+ $X2=2.225 $Y2=1.657
r90 25 30 7.31195 $w=2.05e-07 $l=2.09893e-07 $layer=LI1_cond $X=1.81 $Y=1.555
+ $X2=1.975 $Y2=1.657
r91 25 27 34.9225 $w=3.28e-07 $l=1e-06 $layer=LI1_cond $X=1.81 $Y=1.555 $X2=1.81
+ $Y2=0.555
r92 21 23 66.6596 $w=1.5e-07 $l=1.3e-07 $layer=POLY_cond $X=3.4 $Y=1.33 $X2=3.53
+ $Y2=1.33
r93 17 23 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.53 $Y=1.255
+ $X2=3.53 $Y2=1.33
r94 17 19 194.851 $w=1.5e-07 $l=3.8e-07 $layer=POLY_cond $X=3.53 $Y=1.255
+ $X2=3.53 $Y2=0.875
r95 15 21 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.4 $Y=1.405 $X2=3.4
+ $Y2=1.33
r96 15 16 92.2979 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=3.4 $Y=1.405 $X2=3.4
+ $Y2=1.585
r97 11 13 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=3.175 $Y=2.125
+ $X2=3.175 $Y2=2.525
r98 10 39 62.622 $w=2.54e-07 $l=4.04166e-07 $layer=POLY_cond $X=2.7 $Y=2.05
+ $X2=2.535 $Y2=1.72
r99 9 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.1 $Y=2.05
+ $X2=3.175 $Y2=2.125
r100 9 10 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=3.1 $Y=2.05 $X2=2.7
+ $Y2=2.05
r101 8 41 15.087 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.7 $Y=1.66
+ $X2=2.535 $Y2=1.66
r102 7 16 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.325 $Y=1.66
+ $X2=3.4 $Y2=1.585
r103 7 8 320.479 $w=1.5e-07 $l=6.25e-07 $layer=POLY_cond $X=3.325 $Y=1.66
+ $X2=2.7 $Y2=1.66
r104 2 33 300 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=2 $X=2.16
+ $Y=2.045 $X2=2.31 $Y2=2.19
r105 1 27 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.67
+ $Y=0.345 $X2=1.81 $Y2=0.555
.ends

.subckt PM_SKY130_FD_SC_LP__SDLCLKP_1%A_254_357# 1 2 8 9 10 11 12 15 17 18 20 21
+ 23 24 26 28 31 34 35 38 39 41 42 43 47 52 57 58
c151 38 0 1.18174e-19 $X=2.24 $Y=0.84
c152 20 0 5.31542e-20 $X=2.085 $Y=1.785
c153 17 0 6.36077e-20 $X=2.01 $Y=1.27
r154 57 58 6.90023 $w=3.28e-07 $l=1.75e-07 $layer=LI1_cond $X=5.275 $Y=1.97
+ $X2=5.275 $Y2=1.795
r155 55 58 51.7423 $w=2.43e-07 $l=1.1e-06 $layer=LI1_cond $X=5.232 $Y=0.695
+ $X2=5.232 $Y2=1.795
r156 54 55 3.75023 $w=2.68e-07 $l=8.5e-08 $layer=LI1_cond $X=5.22 $Y=0.61
+ $X2=5.22 $Y2=0.695
r157 52 54 5.97563 $w=2.68e-07 $l=1.4e-07 $layer=LI1_cond $X=5.22 $Y=0.47
+ $X2=5.22 $Y2=0.61
r158 47 49 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=3.765 $Y=0.455
+ $X2=3.765 $Y2=0.61
r159 44 49 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.85 $Y=0.61
+ $X2=3.765 $Y2=0.61
r160 43 54 3.44395 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=5.085 $Y=0.61
+ $X2=5.22 $Y2=0.61
r161 43 44 80.5722 $w=1.68e-07 $l=1.235e-06 $layer=LI1_cond $X=5.085 $Y=0.61
+ $X2=3.85 $Y2=0.61
r162 41 47 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.68 $Y=0.455
+ $X2=3.765 $Y2=0.455
r163 41 42 83.1818 $w=1.68e-07 $l=1.275e-06 $layer=LI1_cond $X=3.68 $Y=0.455
+ $X2=2.405 $Y2=0.455
r164 38 39 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.24
+ $Y=0.84 $X2=2.24 $Y2=0.84
r165 36 42 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=2.275 $Y=0.54
+ $X2=2.405 $Y2=0.455
r166 36 38 13.2974 $w=2.58e-07 $l=3e-07 $layer=LI1_cond $X=2.275 $Y=0.54
+ $X2=2.275 $Y2=0.84
r167 33 39 49.9834 $w=3.95e-07 $l=3.55e-07 $layer=POLY_cond $X=2.207 $Y=1.195
+ $X2=2.207 $Y2=0.84
r168 33 34 5.72943 $w=3.95e-07 $l=7.5e-08 $layer=POLY_cond $X=2.207 $Y=1.195
+ $X2=2.207 $Y2=1.27
r169 29 31 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=3.605 $Y=3.075
+ $X2=3.605 $Y2=2.525
r170 26 28 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=3.04 $Y=1.195
+ $X2=3.04 $Y2=0.875
r171 25 34 19.8978 $w=1.5e-07 $l=1.98e-07 $layer=POLY_cond $X=2.405 $Y=1.27
+ $X2=2.207 $Y2=1.27
r172 24 26 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.965 $Y=1.27
+ $X2=3.04 $Y2=1.195
r173 24 25 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=2.965 $Y=1.27
+ $X2=2.405 $Y2=1.27
r174 21 35 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.085 $Y=1.935
+ $X2=2.085 $Y2=1.86
r175 21 23 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=2.085 $Y=1.935
+ $X2=2.085 $Y2=2.365
r176 20 35 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.085 $Y=1.785
+ $X2=2.085 $Y2=1.86
r177 19 34 5.72943 $w=1.5e-07 $l=1.55029e-07 $layer=POLY_cond $X=2.085 $Y=1.345
+ $X2=2.207 $Y2=1.27
r178 19 20 225.617 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=2.085 $Y=1.345
+ $X2=2.085 $Y2=1.785
r179 17 34 19.8978 $w=1.5e-07 $l=1.97e-07 $layer=POLY_cond $X=2.01 $Y=1.27
+ $X2=2.207 $Y2=1.27
r180 17 18 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=2.01 $Y=1.27
+ $X2=1.67 $Y2=1.27
r181 13 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.595 $Y=1.195
+ $X2=1.67 $Y2=1.27
r182 13 15 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=1.595 $Y=1.195
+ $X2=1.595 $Y2=0.555
r183 11 29 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.53 $Y=3.15
+ $X2=3.605 $Y2=3.075
r184 11 12 1081.94 $w=1.5e-07 $l=2.11e-06 $layer=POLY_cond $X=3.53 $Y=3.15
+ $X2=1.42 $Y2=3.15
r185 9 35 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.01 $Y=1.86
+ $X2=2.085 $Y2=1.86
r186 9 10 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=2.01 $Y=1.86
+ $X2=1.42 $Y2=1.86
r187 8 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.345 $Y=3.075
+ $X2=1.42 $Y2=3.15
r188 7 10 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.345 $Y=1.935
+ $X2=1.42 $Y2=1.86
r189 7 8 584.553 $w=1.5e-07 $l=1.14e-06 $layer=POLY_cond $X=1.345 $Y=1.935
+ $X2=1.345 $Y2=3.075
r190 2 57 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=5.13
+ $Y=1.835 $X2=5.275 $Y2=1.97
r191 1 52 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=5.125
+ $Y=0.26 $X2=5.25 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_LP__SDLCLKP_1%A_737_329# 1 2 9 13 15 17 22 26 28 33 36
+ 39 40 43 44 45 46 50 55 57 58 60 61 69
c134 60 0 2.75113e-19 $X=6.53 $Y=1.51
c135 57 0 8.36873e-20 $X=4.782 $Y=1.73
c136 46 0 1.08032e-19 $X=3.825 $Y=1.73
c137 26 0 8.28063e-20 $X=6.44 $Y=0.865
c138 9 0 3.05678e-20 $X=3.89 $Y=0.875
r139 61 70 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.53 $Y=1.51
+ $X2=6.53 $Y2=1.675
r140 61 69 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.53 $Y=1.51
+ $X2=6.53 $Y2=1.345
r141 60 61 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.53
+ $Y=1.51 $X2=6.53 $Y2=1.51
r142 53 55 7.20277 $w=2.38e-07 $l=1.5e-07 $layer=LI1_cond $X=4.695 $Y=0.985
+ $X2=4.845 $Y2=0.985
r143 50 67 46.504 $w=3.55e-07 $l=1.65e-07 $layer=POLY_cond $X=3.862 $Y=1.81
+ $X2=3.862 $Y2=1.975
r144 50 66 46.504 $w=3.55e-07 $l=1.65e-07 $layer=POLY_cond $X=3.862 $Y=1.81
+ $X2=3.862 $Y2=1.645
r145 49 50 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.85
+ $Y=1.81 $X2=3.85 $Y2=1.81
r146 46 49 3.29269 $w=2.78e-07 $l=8e-08 $layer=LI1_cond $X=3.825 $Y=1.73
+ $X2=3.825 $Y2=1.81
r147 44 60 5.87094 $w=2.63e-07 $l=1.35e-07 $layer=LI1_cond $X=6.497 $Y=1.645
+ $X2=6.497 $Y2=1.51
r148 44 45 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=6.365 $Y=1.645
+ $X2=5.79 $Y2=1.645
r149 42 45 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.705 $Y=1.73
+ $X2=5.79 $Y2=1.645
r150 42 43 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=5.705 $Y=1.73
+ $X2=5.705 $Y2=2.225
r151 41 58 3.3845 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=4.93 $Y=2.31
+ $X2=4.782 $Y2=2.31
r152 40 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.62 $Y=2.31
+ $X2=5.705 $Y2=2.225
r153 40 41 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=5.62 $Y=2.31
+ $X2=4.93 $Y2=2.31
r154 39 57 3.95216 $w=2.32e-07 $l=1.12161e-07 $layer=LI1_cond $X=4.845 $Y=1.645
+ $X2=4.782 $Y2=1.73
r155 38 55 2.75731 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=4.845 $Y=1.105
+ $X2=4.845 $Y2=0.985
r156 38 39 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=4.845 $Y=1.105
+ $X2=4.845 $Y2=1.645
r157 34 58 3.19717 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=4.782 $Y=2.395
+ $X2=4.782 $Y2=2.31
r158 34 36 20.1189 $w=2.93e-07 $l=5.15e-07 $layer=LI1_cond $X=4.782 $Y=2.395
+ $X2=4.782 $Y2=2.91
r159 31 58 3.19717 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=4.782 $Y=2.225
+ $X2=4.782 $Y2=2.31
r160 31 33 10.7431 $w=2.93e-07 $l=2.75e-07 $layer=LI1_cond $X=4.782 $Y=2.225
+ $X2=4.782 $Y2=1.95
r161 30 57 3.95216 $w=2.32e-07 $l=8.5e-08 $layer=LI1_cond $X=4.782 $Y=1.815
+ $X2=4.782 $Y2=1.73
r162 30 33 5.27389 $w=2.93e-07 $l=1.35e-07 $layer=LI1_cond $X=4.782 $Y=1.815
+ $X2=4.782 $Y2=1.95
r163 29 46 3.65648 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=3.965 $Y=1.73
+ $X2=3.825 $Y2=1.73
r164 28 57 2.49072 $w=1.7e-07 $l=1.47e-07 $layer=LI1_cond $X=4.635 $Y=1.73
+ $X2=4.782 $Y2=1.73
r165 28 29 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.635 $Y=1.73
+ $X2=3.965 $Y2=1.73
r166 24 26 94.8617 $w=1.5e-07 $l=1.85e-07 $layer=POLY_cond $X=6.255 $Y=0.865
+ $X2=6.44 $Y2=0.865
r167 22 70 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=6.51 $Y=2.155
+ $X2=6.51 $Y2=1.675
r168 18 26 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.44 $Y=0.94
+ $X2=6.44 $Y2=0.865
r169 18 69 207.67 $w=1.5e-07 $l=4.05e-07 $layer=POLY_cond $X=6.44 $Y=0.94
+ $X2=6.44 $Y2=1.345
r170 15 24 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.255 $Y=0.79
+ $X2=6.255 $Y2=0.865
r171 15 17 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=6.255 $Y=0.79
+ $X2=6.255 $Y2=0.47
r172 13 67 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=3.965 $Y=2.525
+ $X2=3.965 $Y2=1.975
r173 9 66 394.83 $w=1.5e-07 $l=7.7e-07 $layer=POLY_cond $X=3.89 $Y=0.875
+ $X2=3.89 $Y2=1.645
r174 2 36 400 $w=1.7e-07 $l=1.17291e-06 $layer=licon1_PDIFF $count=1 $X=4.59
+ $Y=1.805 $X2=4.73 $Y2=2.91
r175 2 33 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=4.59
+ $Y=1.805 $X2=4.73 $Y2=1.95
r176 1 53 182 $w=1.7e-07 $l=7.71832e-07 $layer=licon1_NDIFF $count=1 $X=4.555
+ $Y=0.245 $X2=4.695 $Y2=0.95
.ends

.subckt PM_SKY130_FD_SC_LP__SDLCLKP_1%A_623_133# 1 2 9 12 16 20 24 25 27 29
r67 25 30 46.3065 $w=3.4e-07 $l=1.65e-07 $layer=POLY_cond $X=4.42 $Y=1.36
+ $X2=4.42 $Y2=1.525
r68 25 29 46.3065 $w=3.4e-07 $l=1.65e-07 $layer=POLY_cond $X=4.42 $Y=1.36
+ $X2=4.42 $Y2=1.195
r69 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.415
+ $Y=1.36 $X2=4.415 $Y2=1.36
r70 22 27 2.80448 $w=2e-07 $l=4.01902e-07 $layer=LI1_cond $X=3.495 $Y=1.375
+ $X2=3.14 $Y2=1.275
r71 22 24 51.0182 $w=1.98e-07 $l=9.2e-07 $layer=LI1_cond $X=3.495 $Y=1.375
+ $X2=4.415 $Y2=1.375
r72 18 27 3.66998 $w=2.97e-07 $l=3.19726e-07 $layer=LI1_cond $X=3.375 $Y=1.475
+ $X2=3.14 $Y2=1.275
r73 18 20 50.4194 $w=2.38e-07 $l=1.05e-06 $layer=LI1_cond $X=3.375 $Y=1.475
+ $X2=3.375 $Y2=2.525
r74 14 27 3.66998 $w=2.97e-07 $l=1.77e-07 $layer=LI1_cond $X=3.317 $Y=1.275
+ $X2=3.14 $Y2=1.275
r75 14 16 12.9853 $w=3.53e-07 $l=4e-07 $layer=LI1_cond $X=3.317 $Y=1.275
+ $X2=3.317 $Y2=0.875
r76 12 30 466.617 $w=1.5e-07 $l=9.1e-07 $layer=POLY_cond $X=4.515 $Y=2.435
+ $X2=4.515 $Y2=1.525
r77 9 29 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=4.48 $Y=0.665
+ $X2=4.48 $Y2=1.195
r78 2 20 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=3.25
+ $Y=2.315 $X2=3.39 $Y2=2.525
r79 1 16 182 $w=1.7e-07 $l=2.93428e-07 $layer=licon1_NDIFF $count=1 $X=3.115
+ $Y=0.665 $X2=3.315 $Y2=0.875
.ends

.subckt PM_SKY130_FD_SC_LP__SDLCLKP_1%CLK 1 3 6 8 10 13 15 16 24
c55 24 0 1.5317e-19 $X=5.895 $Y=1.125
c56 13 0 1.19488e-19 $X=6.08 $Y=2.155
c57 6 0 8.36873e-20 $X=5.49 $Y=2.155
r58 22 24 7.97426 $w=5.44e-07 $l=9e-08 $layer=POLY_cond $X=5.805 $Y=1.125
+ $X2=5.895 $Y2=1.125
r59 22 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.805
+ $Y=0.955 $X2=5.805 $Y2=0.955
r60 20 22 27.9099 $w=5.44e-07 $l=3.15e-07 $layer=POLY_cond $X=5.49 $Y=1.125
+ $X2=5.805 $Y2=1.125
r61 19 20 2.21507 $w=5.44e-07 $l=2.5e-08 $layer=POLY_cond $X=5.465 $Y=1.125
+ $X2=5.49 $Y2=1.125
r62 16 23 7.32733 $w=5.53e-07 $l=3.4e-07 $layer=LI1_cond $X=5.917 $Y=1.295
+ $X2=5.917 $Y2=0.955
r63 15 23 0.646529 $w=5.53e-07 $l=3e-08 $layer=LI1_cond $X=5.917 $Y=0.925
+ $X2=5.917 $Y2=0.955
r64 11 24 16.3915 $w=5.44e-07 $l=4.17373e-07 $layer=POLY_cond $X=6.08 $Y=1.46
+ $X2=5.895 $Y2=1.125
r65 11 13 356.372 $w=1.5e-07 $l=6.95e-07 $layer=POLY_cond $X=6.08 $Y=1.46
+ $X2=6.08 $Y2=2.155
r66 8 24 33.5519 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=5.895 $Y=0.79
+ $X2=5.895 $Y2=1.125
r67 8 10 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=5.895 $Y=0.79
+ $X2=5.895 $Y2=0.47
r68 4 20 33.5519 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=5.49 $Y=1.46
+ $X2=5.49 $Y2=1.125
r69 4 6 356.372 $w=1.5e-07 $l=6.95e-07 $layer=POLY_cond $X=5.49 $Y=1.46 $X2=5.49
+ $Y2=2.155
r70 1 19 33.5519 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=5.465 $Y=0.79
+ $X2=5.465 $Y2=1.125
r71 1 3 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=5.465 $Y=0.79
+ $X2=5.465 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_LP__SDLCLKP_1%A_1231_367# 1 2 9 11 13 18 20 23 25 27 34
c57 34 0 1.55625e-19 $X=7.205 $Y=1.35
c58 27 0 1.5317e-19 $X=6.885 $Y=1.335
r59 30 34 23.6063 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=7.07 $Y=1.35
+ $X2=7.205 $Y2=1.35
r60 30 31 8.74306 $w=3.3e-07 $l=5e-08 $layer=POLY_cond $X=7.07 $Y=1.35 $X2=7.02
+ $Y2=1.35
r61 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.07
+ $Y=1.35 $X2=7.07 $Y2=1.35
r62 27 29 7.94718 $w=2.84e-07 $l=1.85e-07 $layer=LI1_cond $X=6.885 $Y=1.335
+ $X2=7.07 $Y2=1.335
r63 22 27 3.73949 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=6.885 $Y=1.515
+ $X2=6.885 $Y2=1.335
r64 22 23 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=6.885 $Y=1.515
+ $X2=6.885 $Y2=1.91
r65 21 25 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.46 $Y=1.995
+ $X2=6.295 $Y2=1.995
r66 20 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.8 $Y=1.995
+ $X2=6.885 $Y2=1.91
r67 20 21 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=6.8 $Y=1.995
+ $X2=6.46 $Y2=1.995
r68 16 27 16.5387 $w=2.84e-07 $l=5.31954e-07 $layer=LI1_cond $X=6.5 $Y=0.985
+ $X2=6.885 $Y2=1.335
r69 16 18 21.9818 $w=2.68e-07 $l=5.15e-07 $layer=LI1_cond $X=6.5 $Y=0.985
+ $X2=6.5 $Y2=0.47
r70 11 34 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.205 $Y=1.185
+ $X2=7.205 $Y2=1.35
r71 11 13 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=7.205 $Y=1.185
+ $X2=7.205 $Y2=0.655
r72 7 31 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.02 $Y=1.515
+ $X2=7.02 $Y2=1.35
r73 7 9 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=7.02 $Y=1.515 $X2=7.02
+ $Y2=2.465
r74 2 25 300 $w=1.7e-07 $l=2.19089e-07 $layer=licon1_PDIFF $count=2 $X=6.155
+ $Y=1.835 $X2=6.295 $Y2=1.995
r75 1 18 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=6.33
+ $Y=0.26 $X2=6.47 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_LP__SDLCLKP_1%VPWR 1 2 3 4 5 16 18 22 26 34 38 43 44 46
+ 47 49 50 51 53 72 73 79
r85 79 80 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r86 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r87 72 73 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r88 70 73 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=7.44 $Y2=3.33
r89 69 70 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r90 67 70 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=6.48 $Y2=3.33
r91 66 67 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r92 64 67 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.52 $Y2=3.33
r93 63 66 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=4.56 $Y=3.33 $X2=5.52
+ $Y2=3.33
r94 63 64 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r95 61 64 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r96 60 61 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r97 58 79 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.715 $Y=3.33
+ $X2=1.585 $Y2=3.33
r98 58 60 154.294 $w=1.68e-07 $l=2.365e-06 $layer=LI1_cond $X=1.715 $Y=3.33
+ $X2=4.08 $Y2=3.33
r99 57 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r100 57 77 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.24 $Y2=3.33
r101 56 57 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r102 54 76 4.78091 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=3.33
+ $X2=0.212 $Y2=3.33
r103 54 56 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=0.425 $Y=3.33
+ $X2=1.2 $Y2=3.33
r104 53 79 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.455 $Y=3.33
+ $X2=1.585 $Y2=3.33
r105 53 56 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=1.455 $Y=3.33
+ $X2=1.2 $Y2=3.33
r106 51 61 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.84 $Y=3.33
+ $X2=4.08 $Y2=3.33
r107 51 80 0.602067 $w=4.9e-07 $l=2.16e-06 $layer=MET1_cond $X=3.84 $Y=3.33
+ $X2=1.68 $Y2=3.33
r108 49 69 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=6.64 $Y=3.33
+ $X2=6.48 $Y2=3.33
r109 49 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.64 $Y=3.33
+ $X2=6.805 $Y2=3.33
r110 48 72 30.6631 $w=1.68e-07 $l=4.7e-07 $layer=LI1_cond $X=6.97 $Y=3.33
+ $X2=7.44 $Y2=3.33
r111 48 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.97 $Y=3.33
+ $X2=6.805 $Y2=3.33
r112 46 66 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=5.62 $Y=3.33 $X2=5.52
+ $Y2=3.33
r113 46 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.62 $Y=3.33
+ $X2=5.785 $Y2=3.33
r114 45 69 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=5.95 $Y=3.33
+ $X2=6.48 $Y2=3.33
r115 45 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.95 $Y=3.33
+ $X2=5.785 $Y2=3.33
r116 43 60 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=4.135 $Y=3.33
+ $X2=4.08 $Y2=3.33
r117 43 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.135 $Y=3.33
+ $X2=4.3 $Y2=3.33
r118 42 63 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=4.465 $Y=3.33
+ $X2=4.56 $Y2=3.33
r119 42 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.465 $Y=3.33
+ $X2=4.3 $Y2=3.33
r120 38 41 20.0804 $w=3.28e-07 $l=5.75e-07 $layer=LI1_cond $X=6.805 $Y=2.335
+ $X2=6.805 $Y2=2.91
r121 36 50 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.805 $Y=3.245
+ $X2=6.805 $Y2=3.33
r122 36 41 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=6.805 $Y=3.245
+ $X2=6.805 $Y2=2.91
r123 32 47 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.785 $Y=3.245
+ $X2=5.785 $Y2=3.33
r124 32 34 20.7789 $w=3.28e-07 $l=5.95e-07 $layer=LI1_cond $X=5.785 $Y=3.245
+ $X2=5.785 $Y2=2.65
r125 29 31 14.8421 $w=3.28e-07 $l=4.25e-07 $layer=LI1_cond $X=4.3 $Y=2.495
+ $X2=4.3 $Y2=2.92
r126 26 29 14.8421 $w=3.28e-07 $l=4.25e-07 $layer=LI1_cond $X=4.3 $Y=2.07
+ $X2=4.3 $Y2=2.495
r127 24 44 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.3 $Y=3.245 $X2=4.3
+ $Y2=3.33
r128 24 31 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=4.3 $Y=3.245
+ $X2=4.3 $Y2=2.92
r129 20 79 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=1.585 $Y=3.245
+ $X2=1.585 $Y2=3.33
r130 20 22 35.903 $w=2.58e-07 $l=8.1e-07 $layer=LI1_cond $X=1.585 $Y=3.245
+ $X2=1.585 $Y2=2.435
r131 16 76 2.98526 $w=3.3e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.26 $Y=3.245
+ $X2=0.212 $Y2=3.33
r132 16 18 16.0644 $w=3.28e-07 $l=4.6e-07 $layer=LI1_cond $X=0.26 $Y=3.245
+ $X2=0.26 $Y2=2.785
r133 5 41 600 $w=1.7e-07 $l=1.17988e-06 $layer=licon1_PDIFF $count=1 $X=6.585
+ $Y=1.835 $X2=6.805 $Y2=2.91
r134 5 38 600 $w=1.7e-07 $l=6e-07 $layer=licon1_PDIFF $count=1 $X=6.585 $Y=1.835
+ $X2=6.805 $Y2=2.335
r135 4 34 600 $w=1.7e-07 $l=9.18436e-07 $layer=licon1_PDIFF $count=1 $X=5.565
+ $Y=1.835 $X2=5.785 $Y2=2.65
r136 3 31 600 $w=1.7e-07 $l=7.23412e-07 $layer=licon1_PDIFF $count=1 $X=4.04
+ $Y=2.315 $X2=4.3 $Y2=2.92
r137 3 29 600 $w=1.7e-07 $l=3.38231e-07 $layer=licon1_PDIFF $count=1 $X=4.04
+ $Y=2.315 $X2=4.3 $Y2=2.495
r138 3 26 600 $w=1.7e-07 $l=3.62353e-07 $layer=licon1_PDIFF $count=1 $X=4.04
+ $Y=2.315 $X2=4.3 $Y2=2.07
r139 2 22 600 $w=1.7e-07 $l=4.52493e-07 $layer=licon1_PDIFF $count=1 $X=1.495
+ $Y=2.045 $X2=1.63 $Y2=2.435
r140 1 18 600 $w=1.7e-07 $l=5.03637e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.34 $X2=0.26 $Y2=2.785
.ends

.subckt PM_SKY130_FD_SC_LP__SDLCLKP_1%A_154_69# 1 2 3 4 14 17 19 22 23 24 27 30
+ 34 36 38 41
c99 27 0 5.31542e-20 $X=2.942 $Y=1.642
c100 19 0 6.36077e-20 $X=1.885 $Y=2.015
r101 40 41 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=2.885 $Y=1.04
+ $X2=2.885 $Y2=1.5
r102 38 40 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=2.805 $Y=0.875
+ $X2=2.805 $Y2=1.04
r103 31 34 4.73325 $w=2.78e-07 $l=1.15e-07 $layer=LI1_cond $X=0.795 $Y=0.53
+ $X2=0.91 $Y2=0.53
r104 28 30 14.1528 $w=2.83e-07 $l=3.5e-07 $layer=LI1_cond $X=2.942 $Y=2.875
+ $X2=2.942 $Y2=2.525
r105 27 41 7.60349 $w=2.83e-07 $l=1.42e-07 $layer=LI1_cond $X=2.942 $Y=1.642
+ $X2=2.942 $Y2=1.5
r106 27 30 35.7055 $w=2.83e-07 $l=8.83e-07 $layer=LI1_cond $X=2.942 $Y=1.642
+ $X2=2.942 $Y2=2.525
r107 23 28 7.39867 $w=1.7e-07 $l=1.79538e-07 $layer=LI1_cond $X=2.8 $Y=2.96
+ $X2=2.942 $Y2=2.875
r108 23 24 48.6043 $w=1.68e-07 $l=7.45e-07 $layer=LI1_cond $X=2.8 $Y=2.96
+ $X2=2.055 $Y2=2.96
r109 22 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.97 $Y=2.875
+ $X2=2.055 $Y2=2.96
r110 21 22 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=1.97 $Y=2.1
+ $X2=1.97 $Y2=2.875
r111 20 36 3.89502 $w=1.7e-07 $l=2.53e-07 $layer=LI1_cond $X=1.215 $Y=2.015
+ $X2=0.962 $Y2=2.015
r112 19 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.885 $Y=2.015
+ $X2=1.97 $Y2=2.1
r113 19 20 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.885 $Y=2.015
+ $X2=1.215 $Y2=2.015
r114 15 36 2.82881 $w=3.37e-07 $l=8.5e-08 $layer=LI1_cond $X=0.962 $Y=2.1
+ $X2=0.962 $Y2=2.015
r115 15 17 9.11862 $w=5.03e-07 $l=3.85e-07 $layer=LI1_cond $X=0.962 $Y=2.1
+ $X2=0.962 $Y2=2.485
r116 14 36 2.82881 $w=3.37e-07 $l=2.05144e-07 $layer=LI1_cond $X=0.795 $Y=1.93
+ $X2=0.962 $Y2=2.015
r117 13 31 3.65648 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=0.795 $Y=0.67
+ $X2=0.795 $Y2=0.53
r118 13 14 82.2032 $w=1.68e-07 $l=1.26e-06 $layer=LI1_cond $X=0.795 $Y=0.67
+ $X2=0.795 $Y2=1.93
r119 4 30 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=2.835
+ $Y=2.315 $X2=2.96 $Y2=2.525
r120 3 17 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=0.91
+ $Y=2.34 $X2=1.05 $Y2=2.485
r121 2 38 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=2.66
+ $Y=0.665 $X2=2.805 $Y2=0.875
r122 1 34 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.77
+ $Y=0.345 $X2=0.91 $Y2=0.555
.ends

.subckt PM_SKY130_FD_SC_LP__SDLCLKP_1%GCLK 1 2 7 8 9 10 11 12 13 24 48
r14 46 48 0.517952 $w=4.43e-07 $l=2e-08 $layer=LI1_cond $X=7.372 $Y=2.015
+ $X2=7.372 $Y2=2.035
r15 34 48 0.958211 $w=4.43e-07 $l=3.7e-08 $layer=LI1_cond $X=7.372 $Y=2.072
+ $X2=7.372 $Y2=2.035
r16 13 41 3.49618 $w=4.43e-07 $l=1.35e-07 $layer=LI1_cond $X=7.372 $Y=2.775
+ $X2=7.372 $Y2=2.91
r17 12 13 9.58211 $w=4.43e-07 $l=3.7e-07 $layer=LI1_cond $X=7.372 $Y=2.405
+ $X2=7.372 $Y2=2.775
r18 11 46 0.10359 $w=4.43e-07 $l=4e-09 $layer=LI1_cond $X=7.372 $Y=2.011
+ $X2=7.372 $Y2=2.015
r19 11 44 5.93877 $w=4.43e-07 $l=1.61e-07 $layer=LI1_cond $X=7.372 $Y=2.011
+ $X2=7.372 $Y2=1.85
r20 11 12 8.00236 $w=4.43e-07 $l=3.09e-07 $layer=LI1_cond $X=7.372 $Y=2.096
+ $X2=7.372 $Y2=2.405
r21 11 34 0.621542 $w=4.43e-07 $l=2.4e-08 $layer=LI1_cond $X=7.372 $Y=2.096
+ $X2=7.372 $Y2=2.072
r22 10 44 7.89637 $w=2.68e-07 $l=1.85e-07 $layer=LI1_cond $X=7.46 $Y=1.665
+ $X2=7.46 $Y2=1.85
r23 9 10 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=7.46 $Y=1.295
+ $X2=7.46 $Y2=1.665
r24 8 9 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=7.46 $Y=0.925 $X2=7.46
+ $Y2=1.295
r25 7 8 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=7.46 $Y=0.555 $X2=7.46
+ $Y2=0.925
r26 7 24 5.76222 $w=2.68e-07 $l=1.35e-07 $layer=LI1_cond $X=7.46 $Y=0.555
+ $X2=7.46 $Y2=0.42
r27 2 46 400 $w=1.7e-07 $l=2.4e-07 $layer=licon1_PDIFF $count=1 $X=7.095
+ $Y=1.835 $X2=7.235 $Y2=2.015
r28 2 41 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=7.095
+ $Y=1.835 $X2=7.235 $Y2=2.91
r29 1 24 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=7.28
+ $Y=0.235 $X2=7.42 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__SDLCLKP_1%VGND 1 2 3 4 5 18 22 26 30 33 34 36 37 39
+ 40 41 49 60 66 67 71 77
c84 67 0 3.05678e-20 $X=7.44 $Y=0
c85 30 0 8.28063e-20 $X=6.99 $Y=0.38
r86 77 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r87 71 74 9.07985 $w=3.28e-07 $l=2.6e-07 $layer=LI1_cond $X=4.185 $Y=0 $X2=4.185
+ $Y2=0.26
r88 71 72 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r89 67 78 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0 $X2=6.96
+ $Y2=0
r90 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r91 64 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.155 $Y=0 $X2=6.99
+ $Y2=0
r92 64 66 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=7.155 $Y=0 $X2=7.44
+ $Y2=0
r93 63 78 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6.96
+ $Y2=0
r94 62 63 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r95 60 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.825 $Y=0 $X2=6.99
+ $Y2=0
r96 60 62 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=6.825 $Y=0 $X2=6.48
+ $Y2=0
r97 59 63 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=6.48
+ $Y2=0
r98 58 59 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r99 56 59 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.52
+ $Y2=0
r100 56 72 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=4.08
+ $Y2=0
r101 55 58 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=4.56 $Y=0 $X2=5.52
+ $Y2=0
r102 55 56 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r103 53 71 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.35 $Y=0 $X2=4.185
+ $Y2=0
r104 53 55 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=4.35 $Y=0 $X2=4.56
+ $Y2=0
r105 51 52 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r106 49 71 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.02 $Y=0 $X2=4.185
+ $Y2=0
r107 49 51 152.663 $w=1.68e-07 $l=2.34e-06 $layer=LI1_cond $X=4.02 $Y=0 $X2=1.68
+ $Y2=0
r108 48 52 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r109 47 48 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r110 45 48 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r111 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r112 41 72 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.84 $Y=0
+ $X2=4.08 $Y2=0
r113 41 52 0.602067 $w=4.9e-07 $l=2.16e-06 $layer=MET1_cond $X=3.84 $Y=0
+ $X2=1.68 $Y2=0
r114 39 58 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=5.575 $Y=0 $X2=5.52
+ $Y2=0
r115 39 40 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=5.575 $Y=0 $X2=5.68
+ $Y2=0
r116 38 62 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=5.785 $Y=0
+ $X2=6.48 $Y2=0
r117 38 40 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=5.785 $Y=0 $X2=5.68
+ $Y2=0
r118 36 47 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=1.245 $Y=0 $X2=1.2
+ $Y2=0
r119 36 37 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=1.245 $Y=0 $X2=1.36
+ $Y2=0
r120 35 51 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=1.475 $Y=0
+ $X2=1.68 $Y2=0
r121 35 37 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=1.475 $Y=0 $X2=1.36
+ $Y2=0
r122 33 44 3.58824 $w=1.7e-07 $l=5e-08 $layer=LI1_cond $X=0.29 $Y=0 $X2=0.24
+ $Y2=0
r123 33 34 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.29 $Y=0 $X2=0.415
+ $Y2=0
r124 32 47 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=0.54 $Y=0 $X2=1.2
+ $Y2=0
r125 32 34 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.54 $Y=0 $X2=0.415
+ $Y2=0
r126 28 77 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.99 $Y=0.085
+ $X2=6.99 $Y2=0
r127 28 30 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=6.99 $Y=0.085
+ $X2=6.99 $Y2=0.38
r128 24 40 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=5.68 $Y=0.085
+ $X2=5.68 $Y2=0
r129 24 26 20.3333 $w=2.08e-07 $l=3.85e-07 $layer=LI1_cond $X=5.68 $Y=0.085
+ $X2=5.68 $Y2=0.47
r130 20 37 0.280307 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.36 $Y=0.085
+ $X2=1.36 $Y2=0
r131 20 22 21.0446 $w=2.28e-07 $l=4.2e-07 $layer=LI1_cond $X=1.36 $Y=0.085
+ $X2=1.36 $Y2=0.505
r132 16 34 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.415 $Y=0.085
+ $X2=0.415 $Y2=0
r133 16 18 19.361 $w=2.48e-07 $l=4.2e-07 $layer=LI1_cond $X=0.415 $Y=0.085
+ $X2=0.415 $Y2=0.505
r134 5 30 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=6.865
+ $Y=0.235 $X2=6.99 $Y2=0.38
r135 4 26 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=5.54
+ $Y=0.26 $X2=5.68 $Y2=0.47
r136 3 74 182 $w=1.7e-07 $l=5.03115e-07 $layer=licon1_NDIFF $count=1 $X=3.965
+ $Y=0.665 $X2=4.185 $Y2=0.26
r137 2 22 182 $w=1.7e-07 $l=2.26274e-07 $layer=licon1_NDIFF $count=1 $X=1.2
+ $Y=0.345 $X2=1.36 $Y2=0.505
r138 1 18 182 $w=1.7e-07 $l=2.17256e-07 $layer=licon1_NDIFF $count=1 $X=0.32
+ $Y=0.345 $X2=0.455 $Y2=0.505
.ends

