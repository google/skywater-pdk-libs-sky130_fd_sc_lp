# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_lp__sdfrtp_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  15.36000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.050000 1.570000 2.325000 1.760000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  1.209600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 13.665000 0.255000 13.855000 1.045000 ;
        RECT 13.665000 1.045000 14.790000 1.055000 ;
        RECT 13.665000 1.055000 15.260000 1.225000 ;
        RECT 13.665000 1.735000 15.260000 1.985000 ;
        RECT 13.665000 1.985000 13.875000 3.075000 ;
        RECT 14.525000 0.255000 14.790000 1.045000 ;
        RECT 14.545000 1.985000 14.745000 3.075000 ;
        RECT 15.000000 1.225000 15.260000 1.735000 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  0.411000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.210000 1.895000 6.580000 2.130000 ;
        RECT 6.410000 2.130000 6.580000 2.285000 ;
        RECT 6.410000 2.285000 7.370000 2.455000 ;
        RECT 7.200000 2.455000 7.370000 2.725000 ;
        RECT 7.200000 2.725000 8.360000 2.895000 ;
        RECT 8.190000 2.485000 9.690000 2.655000 ;
        RECT 8.190000 2.655000 8.360000 2.725000 ;
        RECT 9.360000 2.245000 9.690000 2.485000 ;
    END
  END RESET_B
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.025000 1.290000 3.475000 2.125000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.550000 1.205000 2.805000 1.400000 ;
        RECT 0.550000 1.400000 0.880000 1.760000 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.315000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 12.155000 1.525000 12.570000 2.525000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 15.360000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.500000 0.500000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.800000 0.500000 3.300000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 15.360000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 15.360000 0.085000 ;
      RECT  0.000000  3.245000 15.360000 3.415000 ;
      RECT  0.155000  0.415000  0.355000 0.795000 ;
      RECT  0.155000  0.795000  1.500000 1.030000 ;
      RECT  0.155000  1.030000  0.380000 1.930000 ;
      RECT  0.155000  1.930000  2.855000 2.125000 ;
      RECT  0.155000  2.125000  1.450000 2.275000 ;
      RECT  0.525000  0.085000  0.855000 0.625000 ;
      RECT  1.045000  0.255000  3.185000 0.425000 ;
      RECT  1.045000  0.425000  1.375000 0.625000 ;
      RECT  1.150000  2.275000  1.450000 2.975000 ;
      RECT  1.620000  2.295000  1.910000 3.245000 ;
      RECT  1.950000  0.595000  2.280000 0.815000 ;
      RECT  1.950000  0.815000  3.075000 0.895000 ;
      RECT  1.950000  0.895000  4.875000 0.970000 ;
      RECT  1.950000  0.970000  4.235000 0.985000 ;
      RECT  2.370000  2.295000  4.235000 2.475000 ;
      RECT  2.370000  2.475000  2.700000 2.975000 ;
      RECT  2.605000  1.770000  2.855000 1.930000 ;
      RECT  2.855000  0.425000  3.185000 0.645000 ;
      RECT  2.905000  0.985000  4.235000 1.065000 ;
      RECT  3.355000  0.085000  3.615000 0.725000 ;
      RECT  3.355000  2.645000  3.685000 3.245000 ;
      RECT  3.780000  1.065000  4.235000 2.295000 ;
      RECT  3.785000  0.640000  4.875000 0.895000 ;
      RECT  3.855000  2.475000  4.235000 2.905000 ;
      RECT  4.405000  1.140000  4.645000 1.880000 ;
      RECT  4.405000  2.135000  6.040000 2.305000 ;
      RECT  4.405000  2.305000  4.825000 2.775000 ;
      RECT  4.815000  1.210000  5.215000 1.380000 ;
      RECT  4.815000  1.380000  4.995000 2.135000 ;
      RECT  5.045000  0.640000  5.955000 0.955000 ;
      RECT  5.045000  0.955000  5.215000 1.210000 ;
      RECT  5.265000  1.665000  7.315000 1.725000 ;
      RECT  5.265000  1.725000  6.040000 1.965000 ;
      RECT  5.360000  2.475000  5.700000 3.245000 ;
      RECT  5.385000  1.125000  5.615000 1.455000 ;
      RECT  5.785000  0.955000  5.955000 1.165000 ;
      RECT  5.785000  1.165000  6.935000 1.385000 ;
      RECT  5.870000  1.555000  7.315000 1.665000 ;
      RECT  5.870000  2.305000  6.040000 2.360000 ;
      RECT  5.870000  2.360000  6.240000 2.690000 ;
      RECT  6.435000  0.085000  6.765000 0.995000 ;
      RECT  6.690000  2.625000  7.020000 3.245000 ;
      RECT  7.105000  0.335000  7.315000 1.555000 ;
      RECT  7.115000  1.725000  7.315000 1.900000 ;
      RECT  7.115000  1.900000  7.565000 2.115000 ;
      RECT  7.485000  0.395000  8.710000 0.945000 ;
      RECT  7.485000  0.945000  7.655000 1.560000 ;
      RECT  7.485000  1.560000  8.020000 1.730000 ;
      RECT  7.735000  1.730000  8.020000 2.545000 ;
      RECT  7.835000  1.175000  8.360000 1.380000 ;
      RECT  8.190000  1.380000  8.360000 2.055000 ;
      RECT  8.190000  2.055000  8.540000 2.315000 ;
      RECT  8.530000  1.485000  8.790000 1.555000 ;
      RECT  8.530000  1.555000 10.390000 1.725000 ;
      RECT  8.530000  1.725000  8.790000 1.815000 ;
      RECT  8.540000  0.945000  8.710000 1.135000 ;
      RECT  8.540000  1.135000 10.485000 1.305000 ;
      RECT  8.820000  2.055000 10.040000 2.075000 ;
      RECT  8.820000  2.075000  9.150000 2.315000 ;
      RECT  8.955000  0.085000  9.285000 0.965000 ;
      RECT  8.980000  1.905000 10.040000 2.055000 ;
      RECT  9.005000  2.825000  9.335000 3.245000 ;
      RECT  9.595000  2.825000 10.040000 3.045000 ;
      RECT  9.720000  1.305000 10.485000 1.375000 ;
      RECT  9.845000  0.255000 10.575000 0.455000 ;
      RECT  9.845000  0.455000 10.145000 0.965000 ;
      RECT  9.870000  2.075000 10.040000 2.825000 ;
      RECT 10.210000  2.665000 10.410000 3.245000 ;
      RECT 10.220000  1.725000 10.390000 2.325000 ;
      RECT 10.220000  2.325000 11.260000 2.495000 ;
      RECT 10.315000  0.625000 12.470000 0.795000 ;
      RECT 10.315000  0.795000 10.485000 1.135000 ;
      RECT 10.665000  0.965000 10.995000 1.165000 ;
      RECT 10.665000  1.165000 10.920000 2.145000 ;
      RECT 11.090000  1.345000 11.985000 1.675000 ;
      RECT 11.090000  1.675000 11.260000 2.325000 ;
      RECT 11.095000  2.665000 11.610000 3.245000 ;
      RECT 11.175000  0.085000 11.505000 0.455000 ;
      RECT 11.430000  2.105000 11.610000 2.665000 ;
      RECT 11.790000  0.975000 12.120000 1.165000 ;
      RECT 11.790000  1.165000 11.985000 1.345000 ;
      RECT 11.805000  1.675000 11.985000 2.670000 ;
      RECT 11.805000  2.670000 12.060000 3.000000 ;
      RECT 12.300000  0.795000 12.470000 1.185000 ;
      RECT 12.300000  1.185000 13.135000 1.355000 ;
      RECT 12.735000  0.255000 12.995000 0.835000 ;
      RECT 12.735000  0.835000 13.475000 1.015000 ;
      RECT 12.740000  1.755000 13.475000 1.925000 ;
      RECT 12.740000  1.925000 12.995000 3.075000 ;
      RECT 12.860000  1.355000 13.135000 1.515000 ;
      RECT 13.165000  0.085000 13.495000 0.665000 ;
      RECT 13.165000  2.095000 13.495000 3.245000 ;
      RECT 13.305000  1.015000 13.475000 1.395000 ;
      RECT 13.305000  1.395000 14.820000 1.565000 ;
      RECT 13.305000  1.565000 13.475000 1.755000 ;
      RECT 14.025000  0.085000 14.355000 0.875000 ;
      RECT 14.045000  2.155000 14.375000 3.245000 ;
      RECT 14.925000  2.155000 15.255000 3.245000 ;
      RECT 14.960000  0.085000 15.255000 0.885000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  1.210000  4.645000 1.380000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  1.210000  5.605000 1.380000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  1.210000  8.005000 1.380000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  1.210000 10.885000 1.380000 ;
      RECT 10.715000  3.245000 10.885000 3.415000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  3.245000 11.365000 3.415000 ;
      RECT 11.675000 -0.085000 11.845000 0.085000 ;
      RECT 11.675000  3.245000 11.845000 3.415000 ;
      RECT 12.155000 -0.085000 12.325000 0.085000 ;
      RECT 12.155000  3.245000 12.325000 3.415000 ;
      RECT 12.635000 -0.085000 12.805000 0.085000 ;
      RECT 12.635000  3.245000 12.805000 3.415000 ;
      RECT 13.115000 -0.085000 13.285000 0.085000 ;
      RECT 13.115000  3.245000 13.285000 3.415000 ;
      RECT 13.595000 -0.085000 13.765000 0.085000 ;
      RECT 13.595000  3.245000 13.765000 3.415000 ;
      RECT 14.075000 -0.085000 14.245000 0.085000 ;
      RECT 14.075000  3.245000 14.245000 3.415000 ;
      RECT 14.555000 -0.085000 14.725000 0.085000 ;
      RECT 14.555000  3.245000 14.725000 3.415000 ;
      RECT 15.035000 -0.085000 15.205000 0.085000 ;
      RECT 15.035000  3.245000 15.205000 3.415000 ;
    LAYER met1 ;
      RECT  4.415000 1.180000  4.705000 1.225000 ;
      RECT  4.415000 1.225000 10.945000 1.365000 ;
      RECT  4.415000 1.365000  4.705000 1.410000 ;
      RECT  5.375000 1.180000  5.665000 1.225000 ;
      RECT  5.375000 1.365000  5.665000 1.410000 ;
      RECT  7.775000 1.180000  8.065000 1.225000 ;
      RECT  7.775000 1.365000  8.065000 1.410000 ;
      RECT 10.655000 1.180000 10.945000 1.225000 ;
      RECT 10.655000 1.365000 10.945000 1.410000 ;
  END
END sky130_fd_sc_lp__sdfrtp_4
