* File: sky130_fd_sc_lp__o22a_2.pxi.spice
* Created: Fri Aug 28 11:09:43 2020
* 
x_PM_SKY130_FD_SC_LP__O22A_2%A_80_23# N_A_80_23#_M1008_d N_A_80_23#_M1011_d
+ N_A_80_23#_M1005_g N_A_80_23#_M1000_g N_A_80_23#_M1007_g N_A_80_23#_M1003_g
+ N_A_80_23#_c_67_n N_A_80_23#_c_68_n N_A_80_23#_c_69_n N_A_80_23#_c_79_p
+ N_A_80_23#_c_106_p N_A_80_23#_c_148_p N_A_80_23#_c_92_p N_A_80_23#_c_80_p
+ N_A_80_23#_c_70_n PM_SKY130_FD_SC_LP__O22A_2%A_80_23#
x_PM_SKY130_FD_SC_LP__O22A_2%B1 N_B1_M1008_g N_B1_M1010_g B1 N_B1_c_153_n
+ N_B1_c_154_n PM_SKY130_FD_SC_LP__O22A_2%B1
x_PM_SKY130_FD_SC_LP__O22A_2%B2 N_B2_M1011_g N_B2_M1009_g B2 N_B2_c_191_n
+ N_B2_c_192_n PM_SKY130_FD_SC_LP__O22A_2%B2
x_PM_SKY130_FD_SC_LP__O22A_2%A2 N_A2_M1004_g N_A2_M1001_g A2 A2 A2 A2
+ N_A2_c_231_n N_A2_c_232_n PM_SKY130_FD_SC_LP__O22A_2%A2
x_PM_SKY130_FD_SC_LP__O22A_2%A1 N_A1_M1002_g N_A1_M1006_g A1 N_A1_c_270_n
+ N_A1_c_271_n PM_SKY130_FD_SC_LP__O22A_2%A1
x_PM_SKY130_FD_SC_LP__O22A_2%VPWR N_VPWR_M1000_s N_VPWR_M1003_s N_VPWR_M1006_d
+ N_VPWR_c_292_n N_VPWR_c_293_n N_VPWR_c_294_n N_VPWR_c_295_n N_VPWR_c_296_n
+ VPWR N_VPWR_c_297_n N_VPWR_c_298_n N_VPWR_c_299_n N_VPWR_c_291_n
+ PM_SKY130_FD_SC_LP__O22A_2%VPWR
x_PM_SKY130_FD_SC_LP__O22A_2%X N_X_M1005_d N_X_M1000_d N_X_c_342_n X X X X X X X
+ PM_SKY130_FD_SC_LP__O22A_2%X
x_PM_SKY130_FD_SC_LP__O22A_2%VGND N_VGND_M1005_s N_VGND_M1007_s N_VGND_M1001_d
+ N_VGND_c_364_n N_VGND_c_365_n N_VGND_c_366_n N_VGND_c_367_n VGND
+ N_VGND_c_368_n N_VGND_c_369_n N_VGND_c_370_n N_VGND_c_371_n N_VGND_c_372_n
+ N_VGND_c_373_n PM_SKY130_FD_SC_LP__O22A_2%VGND
x_PM_SKY130_FD_SC_LP__O22A_2%A_303_49# N_A_303_49#_M1008_s N_A_303_49#_M1009_d
+ N_A_303_49#_M1002_d N_A_303_49#_c_419_n N_A_303_49#_c_449_n
+ N_A_303_49#_c_426_n N_A_303_49#_c_414_n N_A_303_49#_c_415_n
+ N_A_303_49#_c_416_n N_A_303_49#_c_417_n PM_SKY130_FD_SC_LP__O22A_2%A_303_49#
cc_1 VNB N_A_80_23#_M1005_g 0.0249076f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.665
cc_2 VNB N_A_80_23#_M1000_g 0.0059873f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=2.465
cc_3 VNB N_A_80_23#_M1007_g 0.0204627f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=0.665
cc_4 VNB N_A_80_23#_M1003_g 0.00417304f $X=-0.19 $Y=-0.245 $X2=1.01 $Y2=2.465
cc_5 VNB N_A_80_23#_c_67_n 5.05386e-19 $X=-0.19 $Y=-0.245 $X2=1.145 $Y2=1.41
cc_6 VNB N_A_80_23#_c_68_n 0.0229762f $X=-0.19 $Y=-0.245 $X2=1.975 $Y2=1.16
cc_7 VNB N_A_80_23#_c_69_n 0.00237388f $X=-0.19 $Y=-0.245 $X2=1.31 $Y2=1.16
cc_8 VNB N_A_80_23#_c_70_n 0.0815074f $X=-0.19 $Y=-0.245 $X2=1.01 $Y2=1.41
cc_9 VNB N_B1_M1008_g 0.028841f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_B1_c_153_n 0.0270933f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=2.465
cc_11 VNB N_B1_c_154_n 0.00226038f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=2.465
cc_12 VNB N_B2_M1009_g 0.025235f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.245
cc_13 VNB N_B2_c_191_n 0.0249085f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=2.465
cc_14 VNB N_B2_c_192_n 0.00201521f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=2.465
cc_15 VNB N_A2_M1001_g 0.0258939f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.245
cc_16 VNB N_A2_c_231_n 0.024482f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A2_c_232_n 0.0054781f $X=-0.19 $Y=-0.245 $X2=1.01 $Y2=1.575
cc_18 VNB N_A1_M1002_g 0.0297643f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A1_M1006_g 0.00156062f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.245
cc_20 VNB N_A1_c_270_n 0.0521161f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A1_c_271_n 0.0122379f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=1.245
cc_22 VNB N_VPWR_c_291_n 0.163682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB X 4.5117e-19 $X=-0.19 $Y=-0.245 $X2=1.145 $Y2=1.41
cc_24 VNB N_VGND_c_364_n 0.0104214f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_365_n 0.0486435f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=2.465
cc_26 VNB N_VGND_c_366_n 0.00930818f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=0.665
cc_27 VNB N_VGND_c_367_n 0.00594753f $X=-0.19 $Y=-0.245 $X2=1.01 $Y2=2.465
cc_28 VNB N_VGND_c_368_n 0.0153705f $X=-0.19 $Y=-0.245 $X2=1.18 $Y2=1.93
cc_29 VNB N_VGND_c_369_n 0.0386612f $X=-0.19 $Y=-0.245 $X2=1.31 $Y2=1.16
cc_30 VNB N_VGND_c_370_n 0.0192865f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_371_n 0.218394f $X=-0.19 $Y=-0.245 $X2=2.417 $Y2=2.015
cc_32 VNB N_VGND_c_372_n 0.00521013f $X=-0.19 $Y=-0.245 $X2=1.145 $Y2=1.41
cc_33 VNB N_VGND_c_373_n 0.00634414f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_303_49#_c_414_n 0.0132728f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=0.665
cc_35 VNB N_A_303_49#_c_415_n 0.00946976f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=0.665
cc_36 VNB N_A_303_49#_c_416_n 0.0287349f $X=-0.19 $Y=-0.245 $X2=1.01 $Y2=2.465
cc_37 VNB N_A_303_49#_c_417_n 0.00638276f $X=-0.19 $Y=-0.245 $X2=1.18 $Y2=1.245
cc_38 VPB N_A_80_23#_M1000_g 0.0270121f $X=-0.19 $Y=1.655 $X2=0.58 $Y2=2.465
cc_39 VPB N_A_80_23#_M1003_g 0.021927f $X=-0.19 $Y=1.655 $X2=1.01 $Y2=2.465
cc_40 VPB N_A_80_23#_c_67_n 0.00190788f $X=-0.19 $Y=1.655 $X2=1.145 $Y2=1.41
cc_41 VPB N_B1_M1010_g 0.0209699f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=1.245
cc_42 VPB N_B1_c_153_n 0.00764776f $X=-0.19 $Y=1.655 $X2=0.58 $Y2=2.465
cc_43 VPB N_B1_c_154_n 0.00348126f $X=-0.19 $Y=1.655 $X2=0.58 $Y2=2.465
cc_44 VPB N_B2_M1011_g 0.0188007f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_45 VPB N_B2_c_191_n 0.00634975f $X=-0.19 $Y=1.655 $X2=0.58 $Y2=2.465
cc_46 VPB N_B2_c_192_n 0.00343467f $X=-0.19 $Y=1.655 $X2=0.58 $Y2=2.465
cc_47 VPB N_A2_M1004_g 0.0208208f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_48 VPB N_A2_c_231_n 0.00639522f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_49 VPB N_A2_c_232_n 0.00148588f $X=-0.19 $Y=1.655 $X2=1.01 $Y2=1.575
cc_50 VPB N_A1_M1006_g 0.0260227f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=1.245
cc_51 VPB N_A1_c_271_n 0.00942784f $X=-0.19 $Y=1.655 $X2=0.905 $Y2=1.245
cc_52 VPB N_VPWR_c_292_n 0.0133601f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_53 VPB N_VPWR_c_293_n 0.0450759f $X=-0.19 $Y=1.655 $X2=0.58 $Y2=2.465
cc_54 VPB N_VPWR_c_294_n 0.00226008f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_55 VPB N_VPWR_c_295_n 0.0118944f $X=-0.19 $Y=1.655 $X2=1.01 $Y2=2.465
cc_56 VPB N_VPWR_c_296_n 0.048095f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_57 VPB N_VPWR_c_297_n 0.0157463f $X=-0.19 $Y=1.655 $X2=1.975 $Y2=1.16
cc_58 VPB N_VPWR_c_298_n 0.0412428f $X=-0.19 $Y=1.655 $X2=2.09 $Y2=0.76
cc_59 VPB N_VPWR_c_299_n 0.0118777f $X=-0.19 $Y=1.655 $X2=1.01 $Y2=1.41
cc_60 VPB N_VPWR_c_291_n 0.0502638f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_61 VPB X 0.00108671f $X=-0.19 $Y=1.655 $X2=0.58 $Y2=1.41
cc_62 N_A_80_23#_c_67_n N_B1_M1008_g 5.428e-19 $X=1.145 $Y=1.41 $X2=0 $Y2=0
cc_63 N_A_80_23#_c_68_n N_B1_M1008_g 0.0152633f $X=1.975 $Y=1.16 $X2=0 $Y2=0
cc_64 N_A_80_23#_c_70_n N_B1_M1008_g 0.00301504f $X=1.01 $Y=1.41 $X2=0 $Y2=0
cc_65 N_A_80_23#_M1003_g N_B1_M1010_g 0.00911082f $X=1.01 $Y=2.465 $X2=0 $Y2=0
cc_66 N_A_80_23#_c_67_n N_B1_M1010_g 0.00342798f $X=1.145 $Y=1.41 $X2=0 $Y2=0
cc_67 N_A_80_23#_c_79_p N_B1_M1010_g 0.0164337f $X=2.245 $Y=2.015 $X2=0 $Y2=0
cc_68 N_A_80_23#_c_80_p N_B1_M1010_g 0.00314636f $X=2.48 $Y=2.91 $X2=0 $Y2=0
cc_69 N_A_80_23#_M1003_g N_B1_c_153_n 0.00206286f $X=1.01 $Y=2.465 $X2=0 $Y2=0
cc_70 N_A_80_23#_c_67_n N_B1_c_153_n 0.00103952f $X=1.145 $Y=1.41 $X2=0 $Y2=0
cc_71 N_A_80_23#_c_68_n N_B1_c_153_n 0.00526249f $X=1.975 $Y=1.16 $X2=0 $Y2=0
cc_72 N_A_80_23#_c_79_p N_B1_c_153_n 0.00112247f $X=2.245 $Y=2.015 $X2=0 $Y2=0
cc_73 N_A_80_23#_c_70_n N_B1_c_153_n 0.0125f $X=1.01 $Y=1.41 $X2=0 $Y2=0
cc_74 N_A_80_23#_M1003_g N_B1_c_154_n 4.59054e-19 $X=1.01 $Y=2.465 $X2=0 $Y2=0
cc_75 N_A_80_23#_c_67_n N_B1_c_154_n 0.0264585f $X=1.145 $Y=1.41 $X2=0 $Y2=0
cc_76 N_A_80_23#_c_68_n N_B1_c_154_n 0.0297527f $X=1.975 $Y=1.16 $X2=0 $Y2=0
cc_77 N_A_80_23#_c_79_p N_B1_c_154_n 0.0282508f $X=2.245 $Y=2.015 $X2=0 $Y2=0
cc_78 N_A_80_23#_c_70_n N_B1_c_154_n 0.00106277f $X=1.01 $Y=1.41 $X2=0 $Y2=0
cc_79 N_A_80_23#_c_79_p N_B2_M1011_g 0.00921181f $X=2.245 $Y=2.015 $X2=0 $Y2=0
cc_80 N_A_80_23#_c_92_p N_B2_M1011_g 0.00135946f $X=2.417 $Y=2.1 $X2=0 $Y2=0
cc_81 N_A_80_23#_c_80_p N_B2_M1011_g 0.0176284f $X=2.48 $Y=2.91 $X2=0 $Y2=0
cc_82 N_A_80_23#_c_68_n N_B2_M1009_g 0.00340201f $X=1.975 $Y=1.16 $X2=0 $Y2=0
cc_83 N_A_80_23#_c_68_n N_B2_c_191_n 0.00193086f $X=1.975 $Y=1.16 $X2=0 $Y2=0
cc_84 N_A_80_23#_c_92_p N_B2_c_191_n 0.00100362f $X=2.417 $Y=2.1 $X2=0 $Y2=0
cc_85 N_A_80_23#_c_68_n N_B2_c_192_n 0.0106845f $X=1.975 $Y=1.16 $X2=0 $Y2=0
cc_86 N_A_80_23#_c_79_p N_B2_c_192_n 0.0099672f $X=2.245 $Y=2.015 $X2=0 $Y2=0
cc_87 N_A_80_23#_c_92_p N_B2_c_192_n 0.0158761f $X=2.417 $Y=2.1 $X2=0 $Y2=0
cc_88 N_A_80_23#_c_92_p N_A2_M1004_g 0.00149839f $X=2.417 $Y=2.1 $X2=0 $Y2=0
cc_89 N_A_80_23#_c_80_p N_A2_M1004_g 0.0106413f $X=2.48 $Y=2.91 $X2=0 $Y2=0
cc_90 N_A_80_23#_c_92_p N_A2_c_232_n 0.0143384f $X=2.417 $Y=2.1 $X2=0 $Y2=0
cc_91 N_A_80_23#_c_80_p N_A2_c_232_n 0.0668636f $X=2.48 $Y=2.91 $X2=0 $Y2=0
cc_92 N_A_80_23#_c_67_n N_VPWR_M1003_s 0.00171332f $X=1.145 $Y=1.41 $X2=0 $Y2=0
cc_93 N_A_80_23#_c_79_p N_VPWR_M1003_s 0.01586f $X=2.245 $Y=2.015 $X2=0 $Y2=0
cc_94 N_A_80_23#_c_106_p N_VPWR_M1003_s 0.00227149f $X=1.31 $Y=2.015 $X2=0 $Y2=0
cc_95 N_A_80_23#_M1000_g N_VPWR_c_293_n 0.00360788f $X=0.58 $Y=2.465 $X2=0 $Y2=0
cc_96 N_A_80_23#_c_70_n N_VPWR_c_293_n 0.00150165f $X=1.01 $Y=1.41 $X2=0 $Y2=0
cc_97 N_A_80_23#_M1000_g N_VPWR_c_294_n 7.77257e-19 $X=0.58 $Y=2.465 $X2=0 $Y2=0
cc_98 N_A_80_23#_M1003_g N_VPWR_c_294_n 0.0177593f $X=1.01 $Y=2.465 $X2=0 $Y2=0
cc_99 N_A_80_23#_c_79_p N_VPWR_c_294_n 0.0353507f $X=2.245 $Y=2.015 $X2=0 $Y2=0
cc_100 N_A_80_23#_c_106_p N_VPWR_c_294_n 0.0170914f $X=1.31 $Y=2.015 $X2=0 $Y2=0
cc_101 N_A_80_23#_c_80_p N_VPWR_c_294_n 0.0297119f $X=2.48 $Y=2.91 $X2=0 $Y2=0
cc_102 N_A_80_23#_c_70_n N_VPWR_c_294_n 5.725e-19 $X=1.01 $Y=1.41 $X2=0 $Y2=0
cc_103 N_A_80_23#_M1000_g N_VPWR_c_297_n 0.00533769f $X=0.58 $Y=2.465 $X2=0
+ $Y2=0
cc_104 N_A_80_23#_M1003_g N_VPWR_c_297_n 0.00486043f $X=1.01 $Y=2.465 $X2=0
+ $Y2=0
cc_105 N_A_80_23#_c_80_p N_VPWR_c_298_n 0.022005f $X=2.48 $Y=2.91 $X2=0 $Y2=0
cc_106 N_A_80_23#_M1011_d N_VPWR_c_291_n 0.00630397f $X=2.29 $Y=1.835 $X2=0
+ $Y2=0
cc_107 N_A_80_23#_M1000_g N_VPWR_c_291_n 0.0104403f $X=0.58 $Y=2.465 $X2=0 $Y2=0
cc_108 N_A_80_23#_M1003_g N_VPWR_c_291_n 0.00824727f $X=1.01 $Y=2.465 $X2=0
+ $Y2=0
cc_109 N_A_80_23#_c_80_p N_VPWR_c_291_n 0.0130605f $X=2.48 $Y=2.91 $X2=0 $Y2=0
cc_110 N_A_80_23#_M1005_g N_X_c_342_n 0.00945765f $X=0.475 $Y=0.665 $X2=0 $Y2=0
cc_111 N_A_80_23#_M1005_g X 0.00814229f $X=0.475 $Y=0.665 $X2=0 $Y2=0
cc_112 N_A_80_23#_M1007_g X 0.0064766f $X=0.905 $Y=0.665 $X2=0 $Y2=0
cc_113 N_A_80_23#_c_69_n X 0.0143231f $X=1.31 $Y=1.16 $X2=0 $Y2=0
cc_114 N_A_80_23#_c_70_n X 0.00257836f $X=1.01 $Y=1.41 $X2=0 $Y2=0
cc_115 N_A_80_23#_M1000_g X 0.0212414f $X=0.58 $Y=2.465 $X2=0 $Y2=0
cc_116 N_A_80_23#_M1000_g X 0.00458512f $X=0.58 $Y=2.465 $X2=0 $Y2=0
cc_117 N_A_80_23#_M1003_g X 0.00255352f $X=1.01 $Y=2.465 $X2=0 $Y2=0
cc_118 N_A_80_23#_c_67_n X 0.0476929f $X=1.145 $Y=1.41 $X2=0 $Y2=0
cc_119 N_A_80_23#_c_70_n X 0.0309312f $X=1.01 $Y=1.41 $X2=0 $Y2=0
cc_120 N_A_80_23#_M1000_g X 0.0147196f $X=0.58 $Y=2.465 $X2=0 $Y2=0
cc_121 N_A_80_23#_c_79_p A_386_367# 0.007135f $X=2.245 $Y=2.015 $X2=-0.19
+ $Y2=-0.245
cc_122 N_A_80_23#_c_69_n N_VGND_M1007_s 0.00224282f $X=1.31 $Y=1.16 $X2=0 $Y2=0
cc_123 N_A_80_23#_M1005_g N_VGND_c_365_n 0.00679052f $X=0.475 $Y=0.665 $X2=0
+ $Y2=0
cc_124 N_A_80_23#_M1005_g N_VGND_c_366_n 7.07396e-19 $X=0.475 $Y=0.665 $X2=0
+ $Y2=0
cc_125 N_A_80_23#_M1007_g N_VGND_c_366_n 0.0137712f $X=0.905 $Y=0.665 $X2=0
+ $Y2=0
cc_126 N_A_80_23#_c_69_n N_VGND_c_366_n 0.0212355f $X=1.31 $Y=1.16 $X2=0 $Y2=0
cc_127 N_A_80_23#_c_70_n N_VGND_c_366_n 0.00290778f $X=1.01 $Y=1.41 $X2=0 $Y2=0
cc_128 N_A_80_23#_M1005_g N_VGND_c_368_n 0.00554241f $X=0.475 $Y=0.665 $X2=0
+ $Y2=0
cc_129 N_A_80_23#_M1007_g N_VGND_c_368_n 0.00477554f $X=0.905 $Y=0.665 $X2=0
+ $Y2=0
cc_130 N_A_80_23#_M1008_d N_VGND_c_371_n 0.0024127f $X=1.93 $Y=0.245 $X2=0 $Y2=0
cc_131 N_A_80_23#_M1005_g N_VGND_c_371_n 0.0110545f $X=0.475 $Y=0.665 $X2=0
+ $Y2=0
cc_132 N_A_80_23#_M1007_g N_VGND_c_371_n 0.00825815f $X=0.905 $Y=0.665 $X2=0
+ $Y2=0
cc_133 N_A_80_23#_c_68_n N_A_303_49#_M1008_s 0.00230711f $X=1.975 $Y=1.16
+ $X2=-0.19 $Y2=-0.245
cc_134 N_A_80_23#_M1008_d N_A_303_49#_c_419_n 0.00372385f $X=1.93 $Y=0.245 $X2=0
+ $Y2=0
cc_135 N_A_80_23#_c_68_n N_A_303_49#_c_419_n 0.00275981f $X=1.975 $Y=1.16 $X2=0
+ $Y2=0
cc_136 N_A_80_23#_c_148_p N_A_303_49#_c_419_n 0.0141078f $X=2.09 $Y=0.76 $X2=0
+ $Y2=0
cc_137 N_A_80_23#_c_68_n N_A_303_49#_c_415_n 0.00750769f $X=1.975 $Y=1.16 $X2=0
+ $Y2=0
cc_138 N_A_80_23#_M1007_g N_A_303_49#_c_417_n 8.23216e-19 $X=0.905 $Y=0.665
+ $X2=0 $Y2=0
cc_139 N_A_80_23#_c_68_n N_A_303_49#_c_417_n 0.0209786f $X=1.975 $Y=1.16 $X2=0
+ $Y2=0
cc_140 N_B1_M1010_g N_B2_M1011_g 0.0574653f $X=1.855 $Y=2.465 $X2=0 $Y2=0
cc_141 N_B1_M1008_g N_B2_M1009_g 0.033498f $X=1.855 $Y=0.665 $X2=0 $Y2=0
cc_142 N_B1_c_153_n N_B2_c_191_n 0.0574653f $X=1.73 $Y=1.51 $X2=0 $Y2=0
cc_143 N_B1_c_154_n N_B2_c_191_n 3.36937e-19 $X=1.73 $Y=1.51 $X2=0 $Y2=0
cc_144 N_B1_c_153_n N_B2_c_192_n 0.00198723f $X=1.73 $Y=1.51 $X2=0 $Y2=0
cc_145 N_B1_c_154_n N_B2_c_192_n 0.0253746f $X=1.73 $Y=1.51 $X2=0 $Y2=0
cc_146 N_B1_M1010_g N_VPWR_c_294_n 0.0229907f $X=1.855 $Y=2.465 $X2=0 $Y2=0
cc_147 N_B1_M1010_g N_VPWR_c_298_n 0.00486043f $X=1.855 $Y=2.465 $X2=0 $Y2=0
cc_148 N_B1_M1010_g N_VPWR_c_291_n 0.00818711f $X=1.855 $Y=2.465 $X2=0 $Y2=0
cc_149 N_B1_M1008_g N_VGND_c_366_n 0.00328094f $X=1.855 $Y=0.665 $X2=0 $Y2=0
cc_150 N_B1_M1008_g N_VGND_c_369_n 0.00351191f $X=1.855 $Y=0.665 $X2=0 $Y2=0
cc_151 N_B1_M1008_g N_VGND_c_371_n 0.00667569f $X=1.855 $Y=0.665 $X2=0 $Y2=0
cc_152 N_B1_M1008_g N_A_303_49#_c_419_n 0.00860303f $X=1.855 $Y=0.665 $X2=0
+ $Y2=0
cc_153 N_B1_M1008_g N_A_303_49#_c_426_n 5.28929e-19 $X=1.855 $Y=0.665 $X2=0
+ $Y2=0
cc_154 N_B1_M1008_g N_A_303_49#_c_417_n 0.00764405f $X=1.855 $Y=0.665 $X2=0
+ $Y2=0
cc_155 N_B2_M1011_g N_A2_M1004_g 0.0249548f $X=2.215 $Y=2.465 $X2=0 $Y2=0
cc_156 N_B2_c_192_n N_A2_M1004_g 6.05978e-19 $X=2.305 $Y=1.51 $X2=0 $Y2=0
cc_157 N_B2_M1009_g N_A2_M1001_g 0.0203038f $X=2.305 $Y=0.665 $X2=0 $Y2=0
cc_158 N_B2_c_191_n N_A2_c_231_n 0.0209411f $X=2.305 $Y=1.51 $X2=0 $Y2=0
cc_159 N_B2_c_192_n N_A2_c_231_n 9.23418e-19 $X=2.305 $Y=1.51 $X2=0 $Y2=0
cc_160 N_B2_M1011_g N_A2_c_232_n 0.00114415f $X=2.215 $Y=2.465 $X2=0 $Y2=0
cc_161 N_B2_c_191_n N_A2_c_232_n 0.0012428f $X=2.305 $Y=1.51 $X2=0 $Y2=0
cc_162 N_B2_c_192_n N_A2_c_232_n 0.016807f $X=2.305 $Y=1.51 $X2=0 $Y2=0
cc_163 N_B2_M1011_g N_VPWR_c_294_n 0.00345877f $X=2.215 $Y=2.465 $X2=0 $Y2=0
cc_164 N_B2_M1011_g N_VPWR_c_298_n 0.00518588f $X=2.215 $Y=2.465 $X2=0 $Y2=0
cc_165 N_B2_M1011_g N_VPWR_c_291_n 0.00937901f $X=2.215 $Y=2.465 $X2=0 $Y2=0
cc_166 N_B2_M1009_g N_VGND_c_369_n 0.00351219f $X=2.305 $Y=0.665 $X2=0 $Y2=0
cc_167 N_B2_M1009_g N_VGND_c_371_n 0.00546994f $X=2.305 $Y=0.665 $X2=0 $Y2=0
cc_168 N_B2_M1009_g N_A_303_49#_c_419_n 0.0119295f $X=2.305 $Y=0.665 $X2=0 $Y2=0
cc_169 N_B2_M1009_g N_A_303_49#_c_426_n 0.00788452f $X=2.305 $Y=0.665 $X2=0
+ $Y2=0
cc_170 N_B2_M1009_g N_A_303_49#_c_415_n 0.00262489f $X=2.305 $Y=0.665 $X2=0
+ $Y2=0
cc_171 N_B2_c_191_n N_A_303_49#_c_415_n 0.00221754f $X=2.305 $Y=1.51 $X2=0 $Y2=0
cc_172 N_B2_c_192_n N_A_303_49#_c_415_n 0.00576337f $X=2.305 $Y=1.51 $X2=0 $Y2=0
cc_173 N_B2_M1009_g N_A_303_49#_c_417_n 5.25011e-19 $X=2.305 $Y=0.665 $X2=0
+ $Y2=0
cc_174 N_A2_M1001_g N_A1_M1002_g 0.0185126f $X=2.78 $Y=0.665 $X2=0 $Y2=0
cc_175 N_A2_M1004_g N_A1_M1006_g 0.0384123f $X=2.755 $Y=2.465 $X2=0 $Y2=0
cc_176 N_A2_c_231_n N_A1_c_270_n 0.0188788f $X=2.845 $Y=1.51 $X2=0 $Y2=0
cc_177 N_A2_c_232_n N_A1_c_270_n 0.0135158f $X=2.845 $Y=1.51 $X2=0 $Y2=0
cc_178 N_A2_c_232_n N_A1_c_271_n 0.0298773f $X=2.845 $Y=1.51 $X2=0 $Y2=0
cc_179 N_A2_M1004_g N_VPWR_c_296_n 0.00219295f $X=2.755 $Y=2.465 $X2=0 $Y2=0
cc_180 N_A2_M1004_g N_VPWR_c_298_n 0.00492889f $X=2.755 $Y=2.465 $X2=0 $Y2=0
cc_181 N_A2_c_232_n N_VPWR_c_298_n 0.0149608f $X=2.845 $Y=1.51 $X2=0 $Y2=0
cc_182 N_A2_M1004_g N_VPWR_c_291_n 0.00907969f $X=2.755 $Y=2.465 $X2=0 $Y2=0
cc_183 N_A2_c_232_n N_VPWR_c_291_n 0.0156226f $X=2.845 $Y=1.51 $X2=0 $Y2=0
cc_184 N_A2_c_232_n A_566_367# 0.0138018f $X=2.845 $Y=1.51 $X2=-0.19 $Y2=-0.245
cc_185 N_A2_M1001_g N_VGND_c_367_n 0.00317194f $X=2.78 $Y=0.665 $X2=0 $Y2=0
cc_186 N_A2_M1001_g N_VGND_c_369_n 0.00575161f $X=2.78 $Y=0.665 $X2=0 $Y2=0
cc_187 N_A2_M1001_g N_VGND_c_371_n 0.0109404f $X=2.78 $Y=0.665 $X2=0 $Y2=0
cc_188 N_A2_M1001_g N_A_303_49#_c_414_n 0.0151828f $X=2.78 $Y=0.665 $X2=0 $Y2=0
cc_189 N_A2_c_231_n N_A_303_49#_c_414_n 0.00107915f $X=2.845 $Y=1.51 $X2=0 $Y2=0
cc_190 N_A2_c_232_n N_A_303_49#_c_414_n 0.0344321f $X=2.845 $Y=1.51 $X2=0 $Y2=0
cc_191 N_A2_M1001_g N_A_303_49#_c_415_n 0.00102684f $X=2.78 $Y=0.665 $X2=0 $Y2=0
cc_192 N_A2_c_231_n N_A_303_49#_c_415_n 0.00119665f $X=2.845 $Y=1.51 $X2=0 $Y2=0
cc_193 N_A2_M1001_g N_A_303_49#_c_416_n 3.82057e-19 $X=2.78 $Y=0.665 $X2=0 $Y2=0
cc_194 N_A1_M1006_g N_VPWR_c_296_n 0.0199532f $X=3.31 $Y=2.465 $X2=0 $Y2=0
cc_195 N_A1_c_270_n N_VPWR_c_296_n 0.00163033f $X=3.55 $Y=1.46 $X2=0 $Y2=0
cc_196 N_A1_c_271_n N_VPWR_c_296_n 0.0241836f $X=3.55 $Y=1.46 $X2=0 $Y2=0
cc_197 N_A1_M1006_g N_VPWR_c_298_n 0.00544582f $X=3.31 $Y=2.465 $X2=0 $Y2=0
cc_198 N_A1_M1006_g N_VPWR_c_291_n 0.00960156f $X=3.31 $Y=2.465 $X2=0 $Y2=0
cc_199 N_A1_M1002_g N_VGND_c_367_n 0.00311027f $X=3.31 $Y=0.665 $X2=0 $Y2=0
cc_200 N_A1_M1002_g N_VGND_c_370_n 0.00561712f $X=3.31 $Y=0.665 $X2=0 $Y2=0
cc_201 N_A1_M1002_g N_VGND_c_371_n 0.0115216f $X=3.31 $Y=0.665 $X2=0 $Y2=0
cc_202 N_A1_M1002_g N_A_303_49#_c_414_n 0.0192432f $X=3.31 $Y=0.665 $X2=0 $Y2=0
cc_203 N_A1_c_270_n N_A_303_49#_c_414_n 0.00768886f $X=3.55 $Y=1.46 $X2=0 $Y2=0
cc_204 N_A1_c_271_n N_A_303_49#_c_414_n 0.0221569f $X=3.55 $Y=1.46 $X2=0 $Y2=0
cc_205 N_A1_M1002_g N_A_303_49#_c_416_n 0.0111962f $X=3.31 $Y=0.665 $X2=0 $Y2=0
cc_206 N_VPWR_c_291_n N_X_M1000_d 0.0041489f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_207 N_VPWR_c_297_n X 0.016015f $X=1.06 $Y=3.33 $X2=0 $Y2=0
cc_208 N_VPWR_c_291_n X 0.00979641f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_209 N_VPWR_c_291_n A_386_367# 0.00899413f $X=3.6 $Y=3.33 $X2=-0.19 $Y2=-0.245
cc_210 N_VPWR_c_291_n A_566_367# 0.00458283f $X=3.6 $Y=3.33 $X2=-0.19 $Y2=-0.245
cc_211 N_X_c_342_n N_VGND_c_365_n 0.0311671f $X=0.69 $Y=0.42 $X2=0 $Y2=0
cc_212 N_X_c_342_n N_VGND_c_368_n 0.0146515f $X=0.69 $Y=0.42 $X2=0 $Y2=0
cc_213 N_X_M1005_d N_VGND_c_371_n 0.0041489f $X=0.55 $Y=0.245 $X2=0 $Y2=0
cc_214 N_X_c_342_n N_VGND_c_371_n 0.00911037f $X=0.69 $Y=0.42 $X2=0 $Y2=0
cc_215 N_VGND_c_371_n N_A_303_49#_M1008_s 0.00212301f $X=3.6 $Y=0 $X2=-0.19
+ $Y2=-0.245
cc_216 N_VGND_c_371_n N_A_303_49#_M1009_d 0.00259746f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_217 N_VGND_c_371_n N_A_303_49#_M1002_d 0.00212301f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_218 N_VGND_c_369_n N_A_303_49#_c_419_n 0.0323652f $X=2.875 $Y=0 $X2=0 $Y2=0
cc_219 N_VGND_c_371_n N_A_303_49#_c_419_n 0.0201952f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_220 N_VGND_c_369_n N_A_303_49#_c_449_n 0.019189f $X=2.875 $Y=0 $X2=0 $Y2=0
cc_221 N_VGND_c_371_n N_A_303_49#_c_449_n 0.0126947f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_222 N_VGND_M1001_d N_A_303_49#_c_414_n 0.00292615f $X=2.855 $Y=0.245 $X2=0
+ $Y2=0
cc_223 N_VGND_c_367_n N_A_303_49#_c_414_n 0.0216414f $X=3.04 $Y=0.37 $X2=0 $Y2=0
cc_224 N_VGND_c_370_n N_A_303_49#_c_416_n 0.0200241f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_225 N_VGND_c_371_n N_A_303_49#_c_416_n 0.0120544f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_226 N_VGND_c_366_n N_A_303_49#_c_417_n 0.0500526f $X=1.12 $Y=0.39 $X2=0 $Y2=0
cc_227 N_VGND_c_369_n N_A_303_49#_c_417_n 0.021102f $X=2.875 $Y=0 $X2=0 $Y2=0
cc_228 N_VGND_c_371_n N_A_303_49#_c_417_n 0.0126219f $X=3.6 $Y=0 $X2=0 $Y2=0
