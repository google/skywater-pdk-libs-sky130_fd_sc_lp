* File: sky130_fd_sc_lp__a21bo_1.pex.spice
* Created: Wed Sep  2 09:18:41 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A21BO_1%A_80_43# 1 2 9 12 17 18 19 20 21 26 30 33 34
+ 35 38 39 44
c88 17 0 1.80672e-19 $X=0.74 $Y=2.32
c89 12 0 1.82154e-19 $X=0.585 $Y=2.465
r90 39 41 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=2.41 $Y=0.72
+ $X2=2.41 $Y2=0.93
r91 34 45 45.5639 $w=3.95e-07 $l=1.65e-07 $layer=POLY_cond $X=0.597 $Y=1.46
+ $X2=0.597 $Y2=1.625
r92 34 44 45.5639 $w=3.95e-07 $l=1.65e-07 $layer=POLY_cond $X=0.597 $Y=1.46
+ $X2=0.597 $Y2=1.295
r93 33 36 8.51388 $w=2.88e-07 $l=1.65e-07 $layer=LI1_cond $X=0.68 $Y=1.46
+ $X2=0.68 $Y2=1.625
r94 33 35 8.51388 $w=2.88e-07 $l=1.65e-07 $layer=LI1_cond $X=0.68 $Y=1.46
+ $X2=0.68 $Y2=1.295
r95 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.63
+ $Y=1.46 $X2=0.63 $Y2=1.46
r96 28 39 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=2.41 $Y=0.635
+ $X2=2.41 $Y2=0.72
r97 28 30 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=2.41 $Y=0.635
+ $X2=2.41 $Y2=0.38
r98 24 38 3.58051 $w=2.6e-07 $l=1.03078e-07 $layer=LI1_cond $X=1.915 $Y=2.32
+ $X2=1.875 $Y2=2.405
r99 24 26 16.239 $w=2.18e-07 $l=3.1e-07 $layer=LI1_cond $X=1.915 $Y=2.32
+ $X2=1.915 $Y2=2.01
r100 20 38 2.90867 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=1.725 $Y=2.405
+ $X2=1.875 $Y2=2.405
r101 20 21 58.7166 $w=1.68e-07 $l=9e-07 $layer=LI1_cond $X=1.725 $Y=2.405
+ $X2=0.825 $Y2=2.405
r102 18 39 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.245 $Y=0.72
+ $X2=2.41 $Y2=0.72
r103 18 19 92.6417 $w=1.68e-07 $l=1.42e-06 $layer=LI1_cond $X=2.245 $Y=0.72
+ $X2=0.825 $Y2=0.72
r104 17 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.74 $Y=2.32
+ $X2=0.825 $Y2=2.405
r105 17 36 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=0.74 $Y=2.32
+ $X2=0.74 $Y2=1.625
r106 14 19 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.74 $Y=0.805
+ $X2=0.825 $Y2=0.72
r107 14 35 31.9679 $w=1.68e-07 $l=4.9e-07 $layer=LI1_cond $X=0.74 $Y=0.805
+ $X2=0.74 $Y2=1.295
r108 12 45 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=0.585 $Y=2.465
+ $X2=0.585 $Y2=1.625
r109 9 44 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.475 $Y=0.765
+ $X2=0.475 $Y2=1.295
r110 2 38 300 $w=1.7e-07 $l=6.79632e-07 $layer=licon1_PDIFF $count=2 $X=1.765
+ $Y=1.835 $X2=1.89 $Y2=2.455
r111 2 26 600 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=1.765
+ $Y=1.835 $X2=1.89 $Y2=2.01
r112 1 41 182 $w=1.7e-07 $l=8.01795e-07 $layer=licon1_NDIFF $count=1 $X=2.18
+ $Y=0.235 $X2=2.41 $Y2=0.93
r113 1 30 182 $w=1.7e-07 $l=2.93684e-07 $layer=licon1_NDIFF $count=1 $X=2.18
+ $Y=0.235 $X2=2.41 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_LP__A21BO_1%B1_N 3 7 9 12 13
r36 12 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.2 $Y=1.51 $X2=1.2
+ $Y2=1.675
r37 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.2 $Y=1.51 $X2=1.2
+ $Y2=1.345
r38 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.2
+ $Y=1.51 $X2=1.2 $Y2=1.51
r39 9 13 6.3796 $w=2.78e-07 $l=1.55e-07 $layer=LI1_cond $X=1.145 $Y=1.665
+ $X2=1.145 $Y2=1.51
r40 7 14 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=1.135 $Y=0.975
+ $X2=1.135 $Y2=1.345
r41 3 15 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=1.11 $Y=2.045
+ $X2=1.11 $Y2=1.675
.ends

.subckt PM_SKY130_FD_SC_LP__A21BO_1%A_237_367# 1 2 9 13 15 16 17 21 26 28 32
c65 17 0 1.82154e-19 $X=1.465 $Y=2.035
r66 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.81
+ $Y=1.51 $X2=1.81 $Y2=1.51
r67 29 32 9.07985 $w=3.28e-07 $l=2.6e-07 $layer=LI1_cond $X=1.55 $Y=1.51
+ $X2=1.81 $Y2=1.51
r68 27 29 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.55 $Y=1.675
+ $X2=1.55 $Y2=1.51
r69 27 28 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=1.55 $Y=1.675
+ $X2=1.55 $Y2=1.93
r70 26 29 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.55 $Y=1.345
+ $X2=1.55 $Y2=1.51
r71 25 26 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.55 $Y=1.175
+ $X2=1.55 $Y2=1.345
r72 21 25 6.87494 $w=2e-07 $l=1.36015e-07 $layer=LI1_cond $X=1.465 $Y=1.075
+ $X2=1.55 $Y2=1.175
r73 21 23 6.37727 $w=1.98e-07 $l=1.15e-07 $layer=LI1_cond $X=1.465 $Y=1.075
+ $X2=1.35 $Y2=1.075
r74 17 28 6.91519 $w=2.1e-07 $l=1.41244e-07 $layer=LI1_cond $X=1.465 $Y=2.035
+ $X2=1.55 $Y2=1.93
r75 17 19 7.39394 $w=2.08e-07 $l=1.4e-07 $layer=LI1_cond $X=1.465 $Y=2.035
+ $X2=1.325 $Y2=2.035
r76 15 33 38.4695 $w=3.3e-07 $l=2.2e-07 $layer=POLY_cond $X=2.03 $Y=1.51
+ $X2=1.81 $Y2=1.51
r77 15 16 5.03009 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=2.03 $Y=1.51
+ $X2=2.105 $Y2=1.51
r78 11 16 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.105 $Y=1.675
+ $X2=2.105 $Y2=1.51
r79 11 13 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.105 $Y=1.675
+ $X2=2.105 $Y2=2.465
r80 7 16 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.105 $Y=1.345
+ $X2=2.105 $Y2=1.51
r81 7 9 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.105 $Y=1.345
+ $X2=2.105 $Y2=0.655
r82 2 19 600 $w=1.7e-07 $l=2.60768e-07 $layer=licon1_PDIFF $count=1 $X=1.185
+ $Y=1.835 $X2=1.325 $Y2=2.035
r83 1 23 182 $w=1.7e-07 $l=3.58225e-07 $layer=licon1_NDIFF $count=1 $X=1.21
+ $Y=0.765 $X2=1.35 $Y2=1.06
.ends

.subckt PM_SKY130_FD_SC_LP__A21BO_1%A1 3 7 8 9 13 15
c35 13 0 1.24501e-19 $X=2.615 $Y=1.35
r36 13 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.615 $Y=1.35
+ $X2=2.615 $Y2=1.515
r37 13 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.615 $Y=1.35
+ $X2=2.615 $Y2=1.185
r38 9 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.615
+ $Y=1.35 $X2=2.615 $Y2=1.35
r39 8 9 20.9745 $w=2.48e-07 $l=4.55e-07 $layer=LI1_cond $X=2.16 $Y=1.335
+ $X2=2.615 $Y2=1.335
r40 7 15 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.705 $Y=0.655
+ $X2=2.705 $Y2=1.185
r41 3 16 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=2.535 $Y=2.465
+ $X2=2.535 $Y2=1.515
.ends

.subckt PM_SKY130_FD_SC_LP__A21BO_1%A2 3 6 8 9 13 15
r23 13 16 46.5827 $w=3.6e-07 $l=1.65e-07 $layer=POLY_cond $X=3.17 $Y=1.35
+ $X2=3.17 $Y2=1.515
r24 13 15 46.5827 $w=3.6e-07 $l=1.65e-07 $layer=POLY_cond $X=3.17 $Y=1.35
+ $X2=3.17 $Y2=1.185
r25 8 9 22.1269 $w=2.48e-07 $l=4.8e-07 $layer=LI1_cond $X=3.12 $Y=1.335 $X2=3.6
+ $Y2=1.335
r26 8 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.185
+ $Y=1.35 $X2=3.185 $Y2=1.35
r27 6 16 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=3.065 $Y=2.465
+ $X2=3.065 $Y2=1.515
r28 3 15 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=3.065 $Y=0.655
+ $X2=3.065 $Y2=1.185
.ends

.subckt PM_SKY130_FD_SC_LP__A21BO_1%X 1 2 7 8 9 10 11 12 33
r18 31 43 0.758186 $w=3.78e-07 $l=2.5e-08 $layer=LI1_cond $X=0.275 $Y=2.005
+ $X2=0.275 $Y2=1.98
r19 31 33 0.909823 $w=3.78e-07 $l=3e-08 $layer=LI1_cond $X=0.275 $Y=2.005
+ $X2=0.275 $Y2=2.035
r20 12 38 15.3154 $w=3.78e-07 $l=5.05e-07 $layer=LI1_cond $X=0.275 $Y=2.405
+ $X2=0.275 $Y2=2.91
r21 11 43 0.0909823 $w=3.78e-07 $l=3e-09 $layer=LI1_cond $X=0.275 $Y=1.977
+ $X2=0.275 $Y2=1.98
r22 11 41 5.73404 $w=3.78e-07 $l=1.62e-07 $layer=LI1_cond $X=0.275 $Y=1.977
+ $X2=0.275 $Y2=1.815
r23 11 12 10.4023 $w=3.78e-07 $l=3.43e-07 $layer=LI1_cond $X=0.275 $Y=2.062
+ $X2=0.275 $Y2=2.405
r24 11 33 0.818841 $w=3.78e-07 $l=2.7e-08 $layer=LI1_cond $X=0.275 $Y=2.062
+ $X2=0.275 $Y2=2.035
r25 10 41 6.1738 $w=2.78e-07 $l=1.5e-07 $layer=LI1_cond $X=0.225 $Y=1.665
+ $X2=0.225 $Y2=1.815
r26 9 10 15.2287 $w=2.78e-07 $l=3.7e-07 $layer=LI1_cond $X=0.225 $Y=1.295
+ $X2=0.225 $Y2=1.665
r27 8 9 15.2287 $w=2.78e-07 $l=3.7e-07 $layer=LI1_cond $X=0.225 $Y=0.925
+ $X2=0.225 $Y2=1.295
r28 7 8 17.904 $w=2.78e-07 $l=4.35e-07 $layer=LI1_cond $X=0.225 $Y=0.49
+ $X2=0.225 $Y2=0.925
r29 2 43 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.245
+ $Y=1.835 $X2=0.37 $Y2=1.98
r30 2 38 400 $w=1.7e-07 $l=1.13578e-06 $layer=licon1_PDIFF $count=1 $X=0.245
+ $Y=1.835 $X2=0.37 $Y2=2.91
r31 1 7 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.345 $X2=0.26 $Y2=0.49
.ends

.subckt PM_SKY130_FD_SC_LP__A21BO_1%VPWR 1 2 9 13 17 19 24 31 32 35 38
r40 38 39 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r41 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r42 32 39 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=2.64 $Y2=3.33
r43 31 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r44 29 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.965 $Y=3.33
+ $X2=2.8 $Y2=3.33
r45 29 31 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=2.965 $Y=3.33
+ $X2=3.6 $Y2=3.33
r46 28 36 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r47 27 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r48 25 35 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.965 $Y=3.33
+ $X2=0.8 $Y2=3.33
r49 25 27 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=0.965 $Y=3.33
+ $X2=1.2 $Y2=3.33
r50 24 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.635 $Y=3.33
+ $X2=2.8 $Y2=3.33
r51 24 27 93.6203 $w=1.68e-07 $l=1.435e-06 $layer=LI1_cond $X=2.635 $Y=3.33
+ $X2=1.2 $Y2=3.33
r52 22 36 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r53 21 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r54 19 35 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.635 $Y=3.33
+ $X2=0.8 $Y2=3.33
r55 19 21 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=0.635 $Y=3.33
+ $X2=0.24 $Y2=3.33
r56 17 39 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=2.64 $Y2=3.33
r57 17 28 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=1.2 $Y2=3.33
r58 13 16 31.2557 $w=3.28e-07 $l=8.95e-07 $layer=LI1_cond $X=2.8 $Y=2.055
+ $X2=2.8 $Y2=2.95
r59 11 38 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.8 $Y=3.245 $X2=2.8
+ $Y2=3.33
r60 11 16 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.8 $Y=3.245
+ $X2=2.8 $Y2=2.95
r61 7 35 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.8 $Y=3.245 $X2=0.8
+ $Y2=3.33
r62 7 9 16.0644 $w=3.28e-07 $l=4.6e-07 $layer=LI1_cond $X=0.8 $Y=3.245 $X2=0.8
+ $Y2=2.785
r63 2 16 400 $w=1.7e-07 $l=1.20626e-06 $layer=licon1_PDIFF $count=1 $X=2.61
+ $Y=1.835 $X2=2.8 $Y2=2.95
r64 2 13 400 $w=1.7e-07 $l=3.00333e-07 $layer=licon1_PDIFF $count=1 $X=2.61
+ $Y=1.835 $X2=2.8 $Y2=2.055
r65 1 9 600 $w=1.7e-07 $l=1.0176e-06 $layer=licon1_PDIFF $count=1 $X=0.66
+ $Y=1.835 $X2=0.8 $Y2=2.785
.ends

.subckt PM_SKY130_FD_SC_LP__A21BO_1%A_436_367# 1 2 9 13 14 17
c27 14 0 1.24501e-19 $X=2.455 $Y=1.715
r28 17 19 44.6572 $w=2.38e-07 $l=9.3e-07 $layer=LI1_cond $X=3.295 $Y=1.98
+ $X2=3.295 $Y2=2.91
r29 15 17 8.64332 $w=2.38e-07 $l=1.8e-07 $layer=LI1_cond $X=3.295 $Y=1.8
+ $X2=3.295 $Y2=1.98
r30 13 15 7.07814 $w=1.7e-07 $l=1.56844e-07 $layer=LI1_cond $X=3.175 $Y=1.715
+ $X2=3.295 $Y2=1.8
r31 13 14 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=3.175 $Y=1.715
+ $X2=2.455 $Y2=1.715
r32 9 11 41.222 $w=2.58e-07 $l=9.3e-07 $layer=LI1_cond $X=2.325 $Y=1.98
+ $X2=2.325 $Y2=2.91
r33 7 14 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=2.325 $Y=1.8
+ $X2=2.455 $Y2=1.715
r34 7 9 7.97845 $w=2.58e-07 $l=1.8e-07 $layer=LI1_cond $X=2.325 $Y=1.8 $X2=2.325
+ $Y2=1.98
r35 2 19 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=3.14
+ $Y=1.835 $X2=3.28 $Y2=2.91
r36 2 17 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=3.14
+ $Y=1.835 $X2=3.28 $Y2=1.98
r37 1 11 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=2.18
+ $Y=1.835 $X2=2.32 $Y2=2.91
r38 1 9 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.18
+ $Y=1.835 $X2=2.32 $Y2=1.98
.ends

.subckt PM_SKY130_FD_SC_LP__A21BO_1%VGND 1 2 3 14 18 22 25 26 27 33 39 40 43 46
r46 46 47 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r47 43 44 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r48 40 47 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=3.12
+ $Y2=0
r49 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r50 37 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.445 $Y=0 $X2=3.28
+ $Y2=0
r51 37 39 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=3.445 $Y=0 $X2=3.6
+ $Y2=0
r52 36 47 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r53 35 36 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r54 33 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.115 $Y=0 $X2=3.28
+ $Y2=0
r55 33 35 62.3048 $w=1.68e-07 $l=9.55e-07 $layer=LI1_cond $X=3.115 $Y=0 $X2=2.16
+ $Y2=0
r56 32 44 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=0.72
+ $Y2=0
r57 31 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r58 29 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.97 $Y=0 $X2=0.805
+ $Y2=0
r59 29 31 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=0.97 $Y=0 $X2=1.68
+ $Y2=0
r60 27 36 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=2.16
+ $Y2=0
r61 27 32 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=1.68
+ $Y2=0
r62 25 31 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=1.725 $Y=0 $X2=1.68
+ $Y2=0
r63 25 26 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.725 $Y=0 $X2=1.89
+ $Y2=0
r64 24 35 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=2.055 $Y=0 $X2=2.16
+ $Y2=0
r65 24 26 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.055 $Y=0 $X2=1.89
+ $Y2=0
r66 20 46 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.28 $Y=0.085
+ $X2=3.28 $Y2=0
r67 20 22 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=3.28 $Y=0.085
+ $X2=3.28 $Y2=0.38
r68 16 26 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.89 $Y=0.085
+ $X2=1.89 $Y2=0
r69 16 18 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.89 $Y=0.085
+ $X2=1.89 $Y2=0.38
r70 12 43 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.805 $Y=0.085
+ $X2=0.805 $Y2=0
r71 12 14 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.805 $Y=0.085
+ $X2=0.805 $Y2=0.38
r72 3 22 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.14
+ $Y=0.235 $X2=3.28 $Y2=0.38
r73 2 18 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=1.765
+ $Y=0.235 $X2=1.89 $Y2=0.38
r74 1 14 182 $w=1.7e-07 $l=2.71937e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.345 $X2=0.805 $Y2=0.38
.ends

