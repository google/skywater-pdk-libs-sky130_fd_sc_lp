* NGSPICE file created from sky130_fd_sc_lp__nand4b_1.ext - technology: sky130A

.subckt sky130_fd_sc_lp__nand4b_1 A_N B C D VGND VNB VPB VPWR Y
M1000 Y a_71_131# a_442_47# VNB nshort w=840000u l=150000u
+  ad=2.226e+11p pd=2.21e+06u as=3.276e+11p ps=2.46e+06u
M1001 Y D VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=7.056e+11p pd=6.16e+06u as=1.2621e+12p ps=9.73e+06u
M1002 Y B VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 VGND A_N a_71_131# VNB nshort w=420000u l=150000u
+  ad=2.814e+11p pd=2.46e+06u as=1.113e+11p ps=1.37e+06u
M1004 a_262_47# D VGND VNB nshort w=840000u l=150000u
+  ad=1.764e+11p pd=2.1e+06u as=0p ps=0u
M1005 a_334_47# C a_262_47# VNB nshort w=840000u l=150000u
+  ad=3.276e+11p pd=2.46e+06u as=0p ps=0u
M1006 VPWR A_N a_71_131# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1007 a_442_47# B a_334_47# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPWR C Y VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR a_71_131# Y VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

