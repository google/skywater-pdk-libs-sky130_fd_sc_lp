* File: sky130_fd_sc_lp__o21ba_0.pxi.spice
* Created: Fri Aug 28 11:05:28 2020
* 
x_PM_SKY130_FD_SC_LP__O21BA_0%A_80_225# N_A_80_225#_M1004_s N_A_80_225#_M1005_d
+ N_A_80_225#_c_77_n N_A_80_225#_M1001_g N_A_80_225#_M1002_g N_A_80_225#_c_79_n
+ N_A_80_225#_c_80_n N_A_80_225#_c_81_n N_A_80_225#_c_82_n N_A_80_225#_c_87_n
+ N_A_80_225#_c_88_n N_A_80_225#_c_89_n N_A_80_225#_c_83_n N_A_80_225#_c_91_n
+ N_A_80_225#_c_92_n PM_SKY130_FD_SC_LP__O21BA_0%A_80_225#
x_PM_SKY130_FD_SC_LP__O21BA_0%B1_N N_B1_N_c_165_n N_B1_N_M1007_g N_B1_N_M1006_g
+ N_B1_N_c_167_n B1_N B1_N N_B1_N_c_169_n N_B1_N_c_170_n
+ PM_SKY130_FD_SC_LP__O21BA_0%B1_N
x_PM_SKY130_FD_SC_LP__O21BA_0%A_258_397# N_A_258_397#_M1006_d
+ N_A_258_397#_M1007_d N_A_258_397#_c_206_n N_A_258_397#_M1005_g
+ N_A_258_397#_c_208_n N_A_258_397#_M1004_g N_A_258_397#_c_209_n
+ N_A_258_397#_c_210_n N_A_258_397#_c_214_n N_A_258_397#_c_211_n
+ PM_SKY130_FD_SC_LP__O21BA_0%A_258_397#
x_PM_SKY130_FD_SC_LP__O21BA_0%A2 N_A2_M1003_g N_A2_M1008_g N_A2_c_256_n
+ N_A2_c_260_n A2 A2 A2 N_A2_c_258_n PM_SKY130_FD_SC_LP__O21BA_0%A2
x_PM_SKY130_FD_SC_LP__O21BA_0%A1 N_A1_M1009_g N_A1_M1000_g N_A1_c_302_n
+ N_A1_c_303_n A1 A1 A1 N_A1_c_300_n PM_SKY130_FD_SC_LP__O21BA_0%A1
x_PM_SKY130_FD_SC_LP__O21BA_0%X N_X_M1002_s N_X_M1001_s X X X X X X X
+ N_X_c_332_n X PM_SKY130_FD_SC_LP__O21BA_0%X
x_PM_SKY130_FD_SC_LP__O21BA_0%VPWR N_VPWR_M1001_d N_VPWR_M1005_s N_VPWR_M1009_d
+ N_VPWR_c_352_n N_VPWR_c_353_n N_VPWR_c_354_n N_VPWR_c_355_n N_VPWR_c_356_n
+ VPWR N_VPWR_c_357_n N_VPWR_c_358_n N_VPWR_c_359_n N_VPWR_c_351_n
+ N_VPWR_c_361_n N_VPWR_c_362_n PM_SKY130_FD_SC_LP__O21BA_0%VPWR
x_PM_SKY130_FD_SC_LP__O21BA_0%VGND N_VGND_M1002_d N_VGND_M1008_d N_VGND_c_399_n
+ N_VGND_c_400_n N_VGND_c_401_n VGND N_VGND_c_402_n N_VGND_c_403_n
+ N_VGND_c_404_n N_VGND_c_405_n PM_SKY130_FD_SC_LP__O21BA_0%VGND
x_PM_SKY130_FD_SC_LP__O21BA_0%A_499_47# N_A_499_47#_M1004_d N_A_499_47#_M1000_d
+ N_A_499_47#_c_445_n N_A_499_47#_c_446_n N_A_499_47#_c_447_n
+ N_A_499_47#_c_448_n PM_SKY130_FD_SC_LP__O21BA_0%A_499_47#
cc_1 VNB N_A_80_225#_c_77_n 0.0259883f $X=-0.19 $Y=-0.245 $X2=0.577 $Y2=1.618
cc_2 VNB N_A_80_225#_M1002_g 0.0435781f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=0.445
cc_3 VNB N_A_80_225#_c_79_n 0.00293306f $X=-0.19 $Y=-0.245 $X2=0.577 $Y2=1.795
cc_4 VNB N_A_80_225#_c_80_n 0.0014441f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.29
cc_5 VNB N_A_80_225#_c_81_n 0.0213581f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.29
cc_6 VNB N_A_80_225#_c_82_n 0.00942331f $X=-0.19 $Y=-0.245 $X2=0.975 $Y2=1.71
cc_7 VNB N_A_80_225#_c_83_n 0.00426176f $X=-0.19 $Y=-0.245 $X2=2.205 $Y2=0.445
cc_8 VNB N_B1_N_c_165_n 0.0205784f $X=-0.19 $Y=-0.245 $X2=2.355 $Y2=2.435
cc_9 VNB N_B1_N_M1007_g 0.0132002f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_B1_N_c_167_n 0.0222896f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.305
cc_11 VNB B1_N 0.0106053f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.305
cc_12 VNB N_B1_N_c_169_n 0.022628f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_B1_N_c_170_n 0.0216231f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.625
cc_14 VNB N_A_258_397#_c_206_n 0.128694f $X=-0.19 $Y=-0.245 $X2=0.577 $Y2=1.302
cc_15 VNB N_A_258_397#_M1005_g 0.00737173f $X=-0.19 $Y=-0.245 $X2=0.475
+ $Y2=1.795
cc_16 VNB N_A_258_397#_c_208_n 0.0194536f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.305
cc_17 VNB N_A_258_397#_c_209_n 0.00855127f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_258_397#_c_210_n 0.00226931f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.29
cc_19 VNB N_A_258_397#_c_211_n 0.0159106f $X=-0.19 $Y=-0.245 $X2=1.06 $Y2=2.465
cc_20 VNB N_A2_M1008_g 0.0366696f $X=-0.19 $Y=-0.245 $X2=0.577 $Y2=1.302
cc_21 VNB N_A2_c_256_n 0.0218404f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.305
cc_22 VNB A2 0.00568593f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.125
cc_23 VNB N_A2_c_258_n 0.0160096f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.29
cc_24 VNB N_A1_M1000_g 0.0687408f $X=-0.19 $Y=-0.245 $X2=0.577 $Y2=1.302
cc_25 VNB A1 0.0273666f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=0.445
cc_26 VNB N_A1_c_300_n 0.0134109f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.29
cc_27 VNB X 0.0550659f $X=-0.19 $Y=-0.245 $X2=0.577 $Y2=1.302
cc_28 VNB N_X_c_332_n 0.0160437f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VPWR_c_351_n 0.163682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_399_n 0.00524934f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.795
cc_31 VNB N_VGND_c_400_n 0.0440432f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_401_n 0.00507191f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.125
cc_33 VNB N_VGND_c_402_n 0.0198779f $X=-0.19 $Y=-0.245 $X2=2.217 $Y2=2.395
cc_34 VNB N_VGND_c_403_n 0.218955f $X=-0.19 $Y=-0.245 $X2=2.217 $Y2=0.445
cc_35 VNB N_VGND_c_404_n 0.0178959f $X=-0.19 $Y=-0.245 $X2=2.217 $Y2=2.515
cc_36 VNB N_VGND_c_405_n 0.0123963f $X=-0.19 $Y=-0.245 $X2=0.577 $Y2=1.125
cc_37 VNB N_A_499_47#_c_445_n 0.00208349f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.795
cc_38 VNB N_A_499_47#_c_446_n 0.0223f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.305
cc_39 VNB N_A_499_47#_c_447_n 0.00349038f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_499_47#_c_448_n 0.020711f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=0.445
cc_41 VPB N_A_80_225#_M1001_g 0.0255802f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.305
cc_42 VPB N_A_80_225#_c_79_n 0.016779f $X=-0.19 $Y=1.655 $X2=0.577 $Y2=1.795
cc_43 VPB N_A_80_225#_c_82_n 0.00640873f $X=-0.19 $Y=1.655 $X2=0.975 $Y2=1.71
cc_44 VPB N_A_80_225#_c_87_n 0.00191139f $X=-0.19 $Y=1.655 $X2=0.755 $Y2=1.71
cc_45 VPB N_A_80_225#_c_88_n 0.00246218f $X=-0.19 $Y=1.655 $X2=1.06 $Y2=2.465
cc_46 VPB N_A_80_225#_c_89_n 0.00361791f $X=-0.19 $Y=1.655 $X2=1.145 $Y2=2.55
cc_47 VPB N_A_80_225#_c_83_n 0.0117537f $X=-0.19 $Y=1.655 $X2=2.205 $Y2=0.445
cc_48 VPB N_A_80_225#_c_91_n 0.0239419f $X=-0.19 $Y=1.655 $X2=2.1 $Y2=2.515
cc_49 VPB N_A_80_225#_c_92_n 0.00962067f $X=-0.19 $Y=1.655 $X2=2.495 $Y2=2.57
cc_50 VPB N_B1_N_M1007_g 0.033169f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_51 VPB N_A_258_397#_M1005_g 0.0615029f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=1.795
cc_52 VPB N_A_258_397#_c_210_n 0.00853491f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=1.29
cc_53 VPB N_A_258_397#_c_214_n 0.0115378f $X=-0.19 $Y=1.655 $X2=0.975 $Y2=1.71
cc_54 VPB N_A2_M1003_g 0.0392429f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_55 VPB N_A2_c_260_n 0.0179231f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_56 VPB A2 0.00941198f $X=-0.19 $Y=1.655 $X2=0.585 $Y2=1.125
cc_57 VPB N_A1_M1009_g 0.0295652f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_58 VPB N_A1_c_302_n 0.027826f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.305
cc_59 VPB N_A1_c_303_n 0.0266337f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.305
cc_60 VPB A1 0.0314411f $X=-0.19 $Y=1.655 $X2=0.585 $Y2=0.445
cc_61 VPB N_A1_c_300_n 0.00413656f $X=-0.19 $Y=1.655 $X2=0.59 $Y2=1.29
cc_62 VPB X 0.0167868f $X=-0.19 $Y=1.655 $X2=0.577 $Y2=1.302
cc_63 VPB X 0.0387744f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.305
cc_64 VPB X 0.00605788f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_352_n 0.0336592f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_353_n 0.014639f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_67 VPB N_VPWR_c_354_n 0.031297f $X=-0.19 $Y=1.655 $X2=0.59 $Y2=1.29
cc_68 VPB N_VPWR_c_355_n 0.024593f $X=-0.19 $Y=1.655 $X2=0.975 $Y2=1.71
cc_69 VPB N_VPWR_c_356_n 0.00526006f $X=-0.19 $Y=1.655 $X2=0.755 $Y2=1.71
cc_70 VPB N_VPWR_c_357_n 0.0169331f $X=-0.19 $Y=1.655 $X2=2.1 $Y2=2.55
cc_71 VPB N_VPWR_c_358_n 0.0305797f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_72 VPB N_VPWR_c_359_n 0.0135992f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_73 VPB N_VPWR_c_351_n 0.0905683f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_74 VPB N_VPWR_c_361_n 0.00535984f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_75 VPB N_VPWR_c_362_n 0.00535996f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_76 N_A_80_225#_c_80_n N_B1_N_c_165_n 3.72222e-19 $X=0.59 $Y=1.29 $X2=0 $Y2=0
cc_77 N_A_80_225#_c_81_n N_B1_N_c_165_n 0.00679362f $X=0.59 $Y=1.29 $X2=0 $Y2=0
cc_78 N_A_80_225#_c_77_n N_B1_N_M1007_g 0.0115334f $X=0.577 $Y=1.618 $X2=0 $Y2=0
cc_79 N_A_80_225#_M1001_g N_B1_N_M1007_g 0.00650042f $X=0.475 $Y=2.305 $X2=0
+ $Y2=0
cc_80 N_A_80_225#_c_80_n N_B1_N_M1007_g 0.00109777f $X=0.59 $Y=1.29 $X2=0 $Y2=0
cc_81 N_A_80_225#_c_82_n N_B1_N_M1007_g 0.00491215f $X=0.975 $Y=1.71 $X2=0 $Y2=0
cc_82 N_A_80_225#_c_88_n N_B1_N_M1007_g 0.0206896f $X=1.06 $Y=2.465 $X2=0 $Y2=0
cc_83 N_A_80_225#_c_89_n N_B1_N_M1007_g 0.00103411f $X=1.145 $Y=2.55 $X2=0 $Y2=0
cc_84 N_A_80_225#_c_91_n N_B1_N_M1007_g 0.0113025f $X=2.1 $Y=2.515 $X2=0 $Y2=0
cc_85 N_A_80_225#_c_77_n N_B1_N_c_167_n 0.00679362f $X=0.577 $Y=1.618 $X2=0
+ $Y2=0
cc_86 N_A_80_225#_c_82_n N_B1_N_c_167_n 8.10838e-19 $X=0.975 $Y=1.71 $X2=0 $Y2=0
cc_87 N_A_80_225#_M1002_g B1_N 0.00331382f $X=0.585 $Y=0.445 $X2=0 $Y2=0
cc_88 N_A_80_225#_c_80_n B1_N 0.0184808f $X=0.59 $Y=1.29 $X2=0 $Y2=0
cc_89 N_A_80_225#_c_81_n B1_N 0.00203219f $X=0.59 $Y=1.29 $X2=0 $Y2=0
cc_90 N_A_80_225#_c_82_n B1_N 0.012353f $X=0.975 $Y=1.71 $X2=0 $Y2=0
cc_91 N_A_80_225#_M1002_g N_B1_N_c_169_n 0.0101728f $X=0.585 $Y=0.445 $X2=0
+ $Y2=0
cc_92 N_A_80_225#_M1002_g N_B1_N_c_170_n 0.00487596f $X=0.585 $Y=0.445 $X2=0
+ $Y2=0
cc_93 N_A_80_225#_c_83_n N_A_258_397#_c_206_n 0.040704f $X=2.205 $Y=0.445 $X2=0
+ $Y2=0
cc_94 N_A_80_225#_c_83_n N_A_258_397#_M1005_g 0.0307306f $X=2.205 $Y=0.445 $X2=0
+ $Y2=0
cc_95 N_A_80_225#_c_92_n N_A_258_397#_M1005_g 0.0138738f $X=2.495 $Y=2.57 $X2=0
+ $Y2=0
cc_96 N_A_80_225#_c_83_n N_A_258_397#_c_208_n 0.00285568f $X=2.205 $Y=0.445
+ $X2=0 $Y2=0
cc_97 N_A_80_225#_c_83_n N_A_258_397#_c_209_n 0.0268773f $X=2.205 $Y=0.445 $X2=0
+ $Y2=0
cc_98 N_A_80_225#_c_82_n N_A_258_397#_c_210_n 0.00851171f $X=0.975 $Y=1.71 $X2=0
+ $Y2=0
cc_99 N_A_80_225#_c_88_n N_A_258_397#_c_210_n 0.00770794f $X=1.06 $Y=2.465 $X2=0
+ $Y2=0
cc_100 N_A_80_225#_c_83_n N_A_258_397#_c_210_n 0.0208631f $X=2.205 $Y=0.445
+ $X2=0 $Y2=0
cc_101 N_A_80_225#_c_88_n N_A_258_397#_c_214_n 0.0119534f $X=1.06 $Y=2.465 $X2=0
+ $Y2=0
cc_102 N_A_80_225#_c_83_n N_A_258_397#_c_214_n 0.0165502f $X=2.205 $Y=0.445
+ $X2=0 $Y2=0
cc_103 N_A_80_225#_c_91_n N_A_258_397#_c_214_n 0.032797f $X=2.1 $Y=2.515 $X2=0
+ $Y2=0
cc_104 N_A_80_225#_c_83_n N_A_258_397#_c_211_n 0.0502712f $X=2.205 $Y=0.445
+ $X2=0 $Y2=0
cc_105 N_A_80_225#_c_83_n N_A2_M1003_g 0.00152611f $X=2.205 $Y=0.445 $X2=0 $Y2=0
cc_106 N_A_80_225#_c_92_n N_A2_M1003_g 0.0125016f $X=2.495 $Y=2.57 $X2=0 $Y2=0
cc_107 N_A_80_225#_c_83_n N_A2_M1008_g 0.00109041f $X=2.205 $Y=0.445 $X2=0 $Y2=0
cc_108 N_A_80_225#_c_83_n A2 0.0831939f $X=2.205 $Y=0.445 $X2=0 $Y2=0
cc_109 N_A_80_225#_c_92_n A2 0.0120967f $X=2.495 $Y=2.57 $X2=0 $Y2=0
cc_110 N_A_80_225#_c_83_n N_A2_c_258_n 6.93002e-19 $X=2.205 $Y=0.445 $X2=0 $Y2=0
cc_111 N_A_80_225#_c_92_n N_A1_M1009_g 0.00195818f $X=2.495 $Y=2.57 $X2=0 $Y2=0
cc_112 N_A_80_225#_M1002_g X 0.0137994f $X=0.585 $Y=0.445 $X2=0 $Y2=0
cc_113 N_A_80_225#_c_80_n X 0.0378187f $X=0.59 $Y=1.29 $X2=0 $Y2=0
cc_114 N_A_80_225#_c_81_n X 0.0223685f $X=0.59 $Y=1.29 $X2=0 $Y2=0
cc_115 N_A_80_225#_c_87_n X 0.0139057f $X=0.755 $Y=1.71 $X2=0 $Y2=0
cc_116 N_A_80_225#_c_88_n X 0.00515787f $X=1.06 $Y=2.465 $X2=0 $Y2=0
cc_117 N_A_80_225#_c_81_n N_X_c_332_n 0.00184058f $X=0.59 $Y=1.29 $X2=0 $Y2=0
cc_118 N_A_80_225#_M1001_g X 0.00314712f $X=0.475 $Y=2.305 $X2=0 $Y2=0
cc_119 N_A_80_225#_c_88_n N_VPWR_M1001_d 0.00387773f $X=1.06 $Y=2.465 $X2=-0.19
+ $Y2=-0.245
cc_120 N_A_80_225#_c_91_n N_VPWR_M1005_s 0.00965384f $X=2.1 $Y=2.515 $X2=0 $Y2=0
cc_121 N_A_80_225#_c_92_n N_VPWR_M1005_s 0.00182295f $X=2.495 $Y=2.57 $X2=0
+ $Y2=0
cc_122 N_A_80_225#_M1001_g N_VPWR_c_352_n 0.0121315f $X=0.475 $Y=2.305 $X2=0
+ $Y2=0
cc_123 N_A_80_225#_c_79_n N_VPWR_c_352_n 0.00160397f $X=0.577 $Y=1.795 $X2=0
+ $Y2=0
cc_124 N_A_80_225#_c_82_n N_VPWR_c_352_n 0.00410075f $X=0.975 $Y=1.71 $X2=0
+ $Y2=0
cc_125 N_A_80_225#_c_87_n N_VPWR_c_352_n 0.0202866f $X=0.755 $Y=1.71 $X2=0 $Y2=0
cc_126 N_A_80_225#_c_88_n N_VPWR_c_352_n 0.0378233f $X=1.06 $Y=2.465 $X2=0 $Y2=0
cc_127 N_A_80_225#_c_89_n N_VPWR_c_352_n 0.0146274f $X=1.145 $Y=2.55 $X2=0 $Y2=0
cc_128 N_A_80_225#_c_91_n N_VPWR_c_353_n 0.0211422f $X=2.1 $Y=2.515 $X2=0 $Y2=0
cc_129 N_A_80_225#_c_92_n N_VPWR_c_354_n 0.0210986f $X=2.495 $Y=2.57 $X2=0 $Y2=0
cc_130 N_A_80_225#_c_92_n N_VPWR_c_355_n 0.0183199f $X=2.495 $Y=2.57 $X2=0 $Y2=0
cc_131 N_A_80_225#_M1001_g N_VPWR_c_357_n 0.0031218f $X=0.475 $Y=2.305 $X2=0
+ $Y2=0
cc_132 N_A_80_225#_c_89_n N_VPWR_c_358_n 0.00305473f $X=1.145 $Y=2.55 $X2=0
+ $Y2=0
cc_133 N_A_80_225#_c_91_n N_VPWR_c_358_n 0.0118334f $X=2.1 $Y=2.515 $X2=0 $Y2=0
cc_134 N_A_80_225#_M1001_g N_VPWR_c_351_n 0.00376215f $X=0.475 $Y=2.305 $X2=0
+ $Y2=0
cc_135 N_A_80_225#_c_89_n N_VPWR_c_351_n 0.00493499f $X=1.145 $Y=2.55 $X2=0
+ $Y2=0
cc_136 N_A_80_225#_c_91_n N_VPWR_c_351_n 0.0214112f $X=2.1 $Y=2.515 $X2=0 $Y2=0
cc_137 N_A_80_225#_c_92_n N_VPWR_c_351_n 0.0146173f $X=2.495 $Y=2.57 $X2=0 $Y2=0
cc_138 N_A_80_225#_c_83_n N_VGND_c_400_n 0.0127469f $X=2.205 $Y=0.445 $X2=0
+ $Y2=0
cc_139 N_A_80_225#_M1004_s N_VGND_c_403_n 0.00255938f $X=2.08 $Y=0.235 $X2=0
+ $Y2=0
cc_140 N_A_80_225#_M1002_g N_VGND_c_403_n 0.00940608f $X=0.585 $Y=0.445 $X2=0
+ $Y2=0
cc_141 N_A_80_225#_c_83_n N_VGND_c_403_n 0.00894849f $X=2.205 $Y=0.445 $X2=0
+ $Y2=0
cc_142 N_A_80_225#_M1002_g N_VGND_c_404_n 0.00486043f $X=0.585 $Y=0.445 $X2=0
+ $Y2=0
cc_143 N_A_80_225#_M1002_g N_VGND_c_405_n 0.0120127f $X=0.585 $Y=0.445 $X2=0
+ $Y2=0
cc_144 N_A_80_225#_c_80_n N_VGND_c_405_n 0.00307386f $X=0.59 $Y=1.29 $X2=0 $Y2=0
cc_145 N_A_80_225#_c_81_n N_VGND_c_405_n 3.60729e-19 $X=0.59 $Y=1.29 $X2=0 $Y2=0
cc_146 N_A_80_225#_c_83_n N_A_499_47#_c_445_n 0.00977775f $X=2.205 $Y=0.445
+ $X2=0 $Y2=0
cc_147 N_A_80_225#_c_83_n N_A_499_47#_c_447_n 0.0148338f $X=2.205 $Y=0.445 $X2=0
+ $Y2=0
cc_148 N_B1_N_M1007_g N_A_258_397#_c_206_n 0.00266839f $X=1.215 $Y=2.195 $X2=0
+ $Y2=0
cc_149 B1_N N_A_258_397#_c_206_n 4.21255e-19 $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_150 N_B1_N_c_169_n N_A_258_397#_c_206_n 0.0300465f $X=1.2 $Y=0.93 $X2=0 $Y2=0
cc_151 B1_N N_A_258_397#_c_209_n 0.0536937f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_152 N_B1_N_c_170_n N_A_258_397#_c_209_n 0.00609944f $X=1.232 $Y=0.765 $X2=0
+ $Y2=0
cc_153 N_B1_N_M1007_g N_A_258_397#_c_214_n 4.42647e-19 $X=1.215 $Y=2.195 $X2=0
+ $Y2=0
cc_154 N_B1_N_c_167_n N_A_258_397#_c_214_n 0.0035018f $X=1.232 $Y=1.435 $X2=0
+ $Y2=0
cc_155 N_B1_N_c_165_n N_A_258_397#_c_211_n 0.00609944f $X=1.232 $Y=1.238 $X2=0
+ $Y2=0
cc_156 N_B1_N_M1007_g N_A_258_397#_c_211_n 0.012873f $X=1.215 $Y=2.195 $X2=0
+ $Y2=0
cc_157 B1_N X 0.0112046f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_158 N_B1_N_M1007_g N_VPWR_c_352_n 0.00162615f $X=1.215 $Y=2.195 $X2=0 $Y2=0
cc_159 N_B1_N_c_170_n N_VGND_c_400_n 0.00486043f $X=1.232 $Y=0.765 $X2=0 $Y2=0
cc_160 B1_N N_VGND_c_403_n 0.00115705f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_161 N_B1_N_c_170_n N_VGND_c_403_n 0.00970589f $X=1.232 $Y=0.765 $X2=0 $Y2=0
cc_162 B1_N N_VGND_c_405_n 0.0234201f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_163 N_B1_N_c_169_n N_VGND_c_405_n 0.00173431f $X=1.2 $Y=0.93 $X2=0 $Y2=0
cc_164 N_B1_N_c_170_n N_VGND_c_405_n 0.0116648f $X=1.232 $Y=0.765 $X2=0 $Y2=0
cc_165 N_A_258_397#_M1005_g N_A2_M1003_g 0.0320718f $X=2.28 $Y=2.755 $X2=0 $Y2=0
cc_166 N_A_258_397#_c_206_n N_A2_M1008_g 0.00750834f $X=2.28 $Y=1.535 $X2=0
+ $Y2=0
cc_167 N_A_258_397#_c_208_n N_A2_M1008_g 0.0179309f $X=2.42 $Y=0.765 $X2=0 $Y2=0
cc_168 N_A_258_397#_M1005_g N_A2_c_256_n 0.0177019f $X=2.28 $Y=2.755 $X2=0 $Y2=0
cc_169 N_A_258_397#_c_206_n A2 0.00687243f $X=2.28 $Y=1.535 $X2=0 $Y2=0
cc_170 N_A_258_397#_c_206_n N_A2_c_258_n 0.0177019f $X=2.28 $Y=1.535 $X2=0 $Y2=0
cc_171 N_A_258_397#_M1005_g N_VPWR_c_353_n 0.00756704f $X=2.28 $Y=2.755 $X2=0
+ $Y2=0
cc_172 N_A_258_397#_M1005_g N_VPWR_c_355_n 0.00402217f $X=2.28 $Y=2.755 $X2=0
+ $Y2=0
cc_173 N_A_258_397#_M1005_g N_VPWR_c_351_n 0.0048345f $X=2.28 $Y=2.755 $X2=0
+ $Y2=0
cc_174 N_A_258_397#_c_206_n N_VGND_c_400_n 5.03696e-19 $X=2.28 $Y=1.535 $X2=0
+ $Y2=0
cc_175 N_A_258_397#_c_208_n N_VGND_c_400_n 0.00585385f $X=2.42 $Y=0.765 $X2=0
+ $Y2=0
cc_176 N_A_258_397#_c_209_n N_VGND_c_400_n 0.0153489f $X=1.57 $Y=0.445 $X2=0
+ $Y2=0
cc_177 N_A_258_397#_M1006_d N_VGND_c_403_n 0.00376753f $X=1.43 $Y=0.235 $X2=0
+ $Y2=0
cc_178 N_A_258_397#_c_206_n N_VGND_c_403_n 0.00459292f $X=2.28 $Y=1.535 $X2=0
+ $Y2=0
cc_179 N_A_258_397#_c_208_n N_VGND_c_403_n 0.0124078f $X=2.42 $Y=0.765 $X2=0
+ $Y2=0
cc_180 N_A_258_397#_c_209_n N_VGND_c_403_n 0.00990863f $X=1.57 $Y=0.445 $X2=0
+ $Y2=0
cc_181 N_A_258_397#_c_211_n N_VGND_c_403_n 0.00671959f $X=1.835 $Y=1.03 $X2=0
+ $Y2=0
cc_182 N_A_258_397#_c_208_n N_A_499_47#_c_445_n 0.00106926f $X=2.42 $Y=0.765
+ $X2=0 $Y2=0
cc_183 N_A_258_397#_c_206_n N_A_499_47#_c_447_n 0.00182092f $X=2.28 $Y=1.535
+ $X2=0 $Y2=0
cc_184 N_A2_M1008_g N_A1_M1000_g 0.0471841f $X=2.85 $Y=0.445 $X2=0 $Y2=0
cc_185 A2 N_A1_M1000_g 3.45134e-19 $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_186 N_A2_M1003_g N_A1_c_302_n 0.00716063f $X=2.71 $Y=2.755 $X2=0 $Y2=0
cc_187 N_A2_c_260_n N_A1_c_302_n 0.00726874f $X=2.76 $Y=1.825 $X2=0 $Y2=0
cc_188 A2 N_A1_c_302_n 6.40651e-19 $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_189 N_A2_M1003_g N_A1_c_303_n 0.0590135f $X=2.71 $Y=2.755 $X2=0 $Y2=0
cc_190 A2 N_A1_c_303_n 4.64512e-19 $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_191 N_A2_M1003_g A1 0.00153389f $X=2.71 $Y=2.755 $X2=0 $Y2=0
cc_192 N_A2_M1008_g A1 0.0053828f $X=2.85 $Y=0.445 $X2=0 $Y2=0
cc_193 A2 A1 0.0899594f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_194 N_A2_c_256_n N_A1_c_300_n 0.00726874f $X=2.76 $Y=1.66 $X2=0 $Y2=0
cc_195 A2 N_A1_c_300_n 2.37863e-19 $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_196 N_A2_M1003_g N_VPWR_c_353_n 9.35354e-19 $X=2.71 $Y=2.755 $X2=0 $Y2=0
cc_197 N_A2_M1003_g N_VPWR_c_354_n 0.00289441f $X=2.71 $Y=2.755 $X2=0 $Y2=0
cc_198 N_A2_M1003_g N_VPWR_c_355_n 0.00528829f $X=2.71 $Y=2.755 $X2=0 $Y2=0
cc_199 N_A2_M1003_g N_VPWR_c_351_n 0.0097789f $X=2.71 $Y=2.755 $X2=0 $Y2=0
cc_200 N_A2_M1008_g N_VGND_c_399_n 0.00316751f $X=2.85 $Y=0.445 $X2=0 $Y2=0
cc_201 N_A2_M1008_g N_VGND_c_400_n 0.00585385f $X=2.85 $Y=0.445 $X2=0 $Y2=0
cc_202 N_A2_M1008_g N_VGND_c_403_n 0.00619488f $X=2.85 $Y=0.445 $X2=0 $Y2=0
cc_203 N_A2_M1008_g N_A_499_47#_c_445_n 0.00185841f $X=2.85 $Y=0.445 $X2=0 $Y2=0
cc_204 N_A2_M1008_g N_A_499_47#_c_446_n 0.0143743f $X=2.85 $Y=0.445 $X2=0 $Y2=0
cc_205 A2 N_A_499_47#_c_446_n 0.0060865f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_206 A2 N_A_499_47#_c_447_n 0.0242648f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_207 N_A2_c_258_n N_A_499_47#_c_447_n 0.00123457f $X=2.76 $Y=1.32 $X2=0 $Y2=0
cc_208 N_A1_M1009_g N_VPWR_c_354_n 0.0175008f $X=3.1 $Y=2.755 $X2=0 $Y2=0
cc_209 N_A1_c_303_n N_VPWR_c_354_n 0.00233232f $X=3.26 $Y=2.215 $X2=0 $Y2=0
cc_210 A1 N_VPWR_c_354_n 0.0257447f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_211 N_A1_M1009_g N_VPWR_c_355_n 0.00469214f $X=3.1 $Y=2.755 $X2=0 $Y2=0
cc_212 N_A1_M1009_g N_VPWR_c_351_n 0.00818361f $X=3.1 $Y=2.755 $X2=0 $Y2=0
cc_213 N_A1_M1000_g N_VGND_c_399_n 0.00319852f $X=3.28 $Y=0.445 $X2=0 $Y2=0
cc_214 N_A1_M1000_g N_VGND_c_402_n 0.00585385f $X=3.28 $Y=0.445 $X2=0 $Y2=0
cc_215 N_A1_M1000_g N_VGND_c_403_n 0.00723478f $X=3.28 $Y=0.445 $X2=0 $Y2=0
cc_216 N_A1_M1000_g N_A_499_47#_c_446_n 0.0135841f $X=3.28 $Y=0.445 $X2=0 $Y2=0
cc_217 A1 N_A_499_47#_c_446_n 0.0445654f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_218 N_A1_c_300_n N_A_499_47#_c_446_n 5.81926e-19 $X=3.33 $Y=1.71 $X2=0 $Y2=0
cc_219 N_A1_M1000_g N_A_499_47#_c_448_n 0.00403231f $X=3.28 $Y=0.445 $X2=0 $Y2=0
cc_220 X N_VPWR_c_352_n 6.66668e-19 $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_221 X N_VPWR_c_352_n 0.0486901f $X=0.24 $Y=2.035 $X2=0 $Y2=0
cc_222 X N_VPWR_c_357_n 0.010123f $X=0.155 $Y=1.95 $X2=0 $Y2=0
cc_223 X N_VPWR_c_351_n 0.00962496f $X=0.155 $Y=1.95 $X2=0 $Y2=0
cc_224 N_X_M1002_s N_VGND_c_403_n 0.00373326f $X=0.245 $Y=0.235 $X2=0 $Y2=0
cc_225 N_X_c_332_n N_VGND_c_403_n 0.0143005f $X=0.37 $Y=0.445 $X2=0 $Y2=0
cc_226 N_X_c_332_n N_VGND_c_404_n 0.021604f $X=0.37 $Y=0.445 $X2=0 $Y2=0
cc_227 N_VGND_c_403_n N_A_499_47#_M1004_d 0.00269268f $X=3.6 $Y=0 $X2=-0.19
+ $Y2=-0.245
cc_228 N_VGND_c_403_n N_A_499_47#_M1000_d 0.00224632f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_229 N_VGND_c_400_n N_A_499_47#_c_445_n 0.0128989f $X=2.935 $Y=0 $X2=0 $Y2=0
cc_230 N_VGND_c_403_n N_A_499_47#_c_445_n 0.00990863f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_231 N_VGND_c_399_n N_A_499_47#_c_446_n 0.0168902f $X=3.065 $Y=0.445 $X2=0
+ $Y2=0
cc_232 N_VGND_c_403_n N_A_499_47#_c_446_n 0.0111518f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_233 N_VGND_c_402_n N_A_499_47#_c_448_n 0.0162773f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_234 N_VGND_c_403_n N_A_499_47#_c_448_n 0.0110608f $X=3.6 $Y=0 $X2=0 $Y2=0
