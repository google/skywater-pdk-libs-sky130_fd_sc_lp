* File: sky130_fd_sc_lp__fa_2.pex.spice
* Created: Wed Sep  2 09:53:16 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__FA_2%A_84_21# 1 2 9 13 15 19 23 25 26 31 34 35 37 38
+ 39 41 43 47 51 58 63
c151 63 0 4.16358e-19 $X=4.41 $Y=2.24
c152 37 0 1.39673e-19 $X=3.605 $Y=1.87
c153 23 0 1.55518e-19 $X=0.925 $Y=2.465
c154 15 0 1.80747e-19 $X=0.85 $Y=1.42
c155 9 0 7.53306e-20 $X=0.495 $Y=0.655
r156 58 60 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=3.69 $Y=1.87
+ $X2=3.69 $Y2=2.16
r157 51 53 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=2.955 $Y=1.17
+ $X2=2.955 $Y2=1.315
r158 47 49 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=1.575 $Y=1.315
+ $X2=1.575 $Y2=1.51
r159 44 60 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.775 $Y=2.16
+ $X2=3.69 $Y2=2.16
r160 43 63 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=4.245 $Y=2.16
+ $X2=4.375 $Y2=2.16
r161 43 44 30.6631 $w=1.68e-07 $l=4.7e-07 $layer=LI1_cond $X=4.245 $Y=2.16
+ $X2=3.775 $Y2=2.16
r162 39 56 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=3.63 $Y=0.805
+ $X2=3.63 $Y2=1.17
r163 39 41 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=3.715 $Y=0.805
+ $X2=4.41 $Y2=0.805
r164 37 58 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.605 $Y=1.87
+ $X2=3.69 $Y2=1.87
r165 37 38 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=3.605 $Y=1.87
+ $X2=3.04 $Y2=1.87
r166 36 51 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.04 $Y=1.17
+ $X2=2.955 $Y2=1.17
r167 35 56 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.545 $Y=1.17
+ $X2=3.63 $Y2=1.17
r168 35 36 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=3.545 $Y=1.17
+ $X2=3.04 $Y2=1.17
r169 34 38 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.955 $Y=1.785
+ $X2=3.04 $Y2=1.87
r170 33 53 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=2.955 $Y=1.4
+ $X2=2.955 $Y2=1.315
r171 33 34 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=2.955 $Y=1.4
+ $X2=2.955 $Y2=1.785
r172 32 47 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.66 $Y=1.315
+ $X2=1.575 $Y2=1.315
r173 31 53 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.87 $Y=1.315
+ $X2=2.955 $Y2=1.315
r174 31 32 78.9412 $w=1.68e-07 $l=1.21e-06 $layer=LI1_cond $X=2.87 $Y=1.315
+ $X2=1.66 $Y2=1.315
r175 29 67 46.255 $w=3.35e-07 $l=1.65e-07 $layer=POLY_cond $X=1.017 $Y=1.51
+ $X2=1.017 $Y2=1.675
r176 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.02
+ $Y=1.51 $X2=1.02 $Y2=1.51
r177 26 49 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.49 $Y=1.51
+ $X2=1.575 $Y2=1.51
r178 26 28 30.6631 $w=1.68e-07 $l=4.7e-07 $layer=LI1_cond $X=1.49 $Y=1.51
+ $X2=1.02 $Y2=1.51
r179 23 67 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=0.925 $Y=2.465
+ $X2=0.925 $Y2=1.675
r180 19 65 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=0.925 $Y=0.655
+ $X2=0.925 $Y2=1.345
r181 16 25 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.57 $Y=1.42
+ $X2=0.495 $Y2=1.42
r182 15 29 15.5026 $w=3.35e-07 $l=9e-08 $layer=POLY_cond $X=1.017 $Y=1.42
+ $X2=1.017 $Y2=1.51
r183 15 65 30.7523 $w=3.35e-07 $l=7.5e-08 $layer=POLY_cond $X=1.017 $Y=1.42
+ $X2=1.017 $Y2=1.345
r184 15 16 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=0.85 $Y=1.42
+ $X2=0.57 $Y2=1.42
r185 11 25 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.495 $Y=1.495
+ $X2=0.495 $Y2=1.42
r186 11 13 497.383 $w=1.5e-07 $l=9.7e-07 $layer=POLY_cond $X=0.495 $Y=1.495
+ $X2=0.495 $Y2=2.465
r187 7 25 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.495 $Y=1.345
+ $X2=0.495 $Y2=1.42
r188 7 9 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=0.495 $Y=1.345
+ $X2=0.495 $Y2=0.655
r189 2 63 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=4.27
+ $Y=2.095 $X2=4.41 $Y2=2.24
r190 1 41 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=4.27
+ $Y=0.595 $X2=4.41 $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_LP__FA_2%A 3 7 11 15 19 23 27 31 33 38 41 42 43 44 47 48
+ 49 50 56 57 59 60 67 73 74
c210 43 0 1.43592e-19 $X=5.475 $Y=1.93
c211 38 0 1.83475e-19 $X=5.305 $Y=1.42
c212 19 0 6.9935e-20 $X=6.19 $Y=2.54
c213 15 0 3.16332e-20 $X=3.475 $Y=2.415
r214 73 76 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.1 $Y=1.51
+ $X2=8.1 $Y2=1.675
r215 73 75 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.1 $Y=1.51
+ $X2=8.1 $Y2=1.345
r216 73 74 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.1
+ $Y=1.51 $X2=8.1 $Y2=1.51
r217 63 65 13.9889 $w=3.3e-07 $l=8e-08 $layer=POLY_cond $X=2.965 $Y=1.52
+ $X2=3.045 $Y2=1.52
r218 60 74 6.19223 $w=3.33e-07 $l=1.8e-07 $layer=LI1_cond $X=7.92 $Y=1.582
+ $X2=8.1 $Y2=1.582
r219 60 79 0.344013 $w=3.33e-07 $l=1e-08 $layer=LI1_cond $X=7.92 $Y=1.582
+ $X2=7.91 $Y2=1.582
r220 60 79 4.05585 $w=1.9e-07 $l=1.68e-07 $layer=LI1_cond $X=7.91 $Y=1.75
+ $X2=7.91 $Y2=1.582
r221 59 60 19.7652 $w=3.58e-07 $l=5.75e-07 $layer=LI1_cond $X=7.91 $Y=2.325
+ $X2=7.91 $Y2=1.75
r222 57 58 3.47987 $w=2.98e-07 $l=8.5e-08 $layer=LI1_cond $X=6.28 $Y=1.93
+ $X2=6.28 $Y2=2.015
r223 56 71 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.28 $Y=1.77
+ $X2=6.28 $Y2=1.935
r224 56 70 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.28 $Y=1.77
+ $X2=6.28 $Y2=1.605
r225 55 57 6.55034 $w=2.98e-07 $l=1.6e-07 $layer=LI1_cond $X=6.28 $Y=1.77
+ $X2=6.28 $Y2=1.93
r226 55 56 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.28
+ $Y=1.77 $X2=6.28 $Y2=1.77
r227 50 52 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=4.41 $Y=1.42
+ $X2=4.41 $Y2=1.525
r228 48 59 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=7.815 $Y=2.41
+ $X2=7.91 $Y2=2.325
r229 48 49 57.4118 $w=1.68e-07 $l=8.8e-07 $layer=LI1_cond $X=7.815 $Y=2.41
+ $X2=6.935 $Y2=2.41
r230 47 49 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.85 $Y=2.325
+ $X2=6.935 $Y2=2.41
r231 46 47 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=6.85 $Y=2.1
+ $X2=6.85 $Y2=2.325
r232 45 58 4.02169 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.445 $Y=2.015
+ $X2=6.28 $Y2=2.015
r233 44 46 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.765 $Y=2.015
+ $X2=6.85 $Y2=2.1
r234 44 45 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=6.765 $Y=2.015
+ $X2=6.445 $Y2=2.015
r235 42 57 4.02169 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.115 $Y=1.93
+ $X2=6.28 $Y2=1.93
r236 42 43 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=6.115 $Y=1.93
+ $X2=5.475 $Y2=1.93
r237 41 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.39 $Y=1.845
+ $X2=5.475 $Y2=1.93
r238 40 41 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=5.39 $Y=1.505
+ $X2=5.39 $Y2=1.845
r239 39 50 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.495 $Y=1.42
+ $X2=4.41 $Y2=1.42
r240 38 40 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.305 $Y=1.42
+ $X2=5.39 $Y2=1.505
r241 38 39 52.8449 $w=1.68e-07 $l=8.1e-07 $layer=LI1_cond $X=5.305 $Y=1.42
+ $X2=4.495 $Y2=1.42
r242 36 67 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=3.385 $Y=1.52
+ $X2=3.475 $Y2=1.52
r243 36 65 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=3.385 $Y=1.52
+ $X2=3.045 $Y2=1.52
r244 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.385
+ $Y=1.52 $X2=3.385 $Y2=1.52
r245 33 52 0.364908 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=4.325 $Y=1.525
+ $X2=4.41 $Y2=1.525
r246 33 35 57.9192 $w=1.78e-07 $l=9.4e-07 $layer=LI1_cond $X=4.325 $Y=1.525
+ $X2=3.385 $Y2=1.525
r247 31 76 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=8.19 $Y=2.155
+ $X2=8.19 $Y2=1.675
r248 27 75 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=8.19 $Y=0.895
+ $X2=8.19 $Y2=1.345
r249 23 70 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=6.29 $Y=0.805
+ $X2=6.29 $Y2=1.605
r250 19 71 310.223 $w=1.5e-07 $l=6.05e-07 $layer=POLY_cond $X=6.19 $Y=2.54
+ $X2=6.19 $Y2=1.935
r251 13 67 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.475 $Y=1.685
+ $X2=3.475 $Y2=1.52
r252 13 15 374.319 $w=1.5e-07 $l=7.3e-07 $layer=POLY_cond $X=3.475 $Y=1.685
+ $X2=3.475 $Y2=2.415
r253 9 67 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.475 $Y=1.355
+ $X2=3.475 $Y2=1.52
r254 9 11 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=3.475 $Y=1.355
+ $X2=3.475 $Y2=0.805
r255 5 65 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.045 $Y=1.355
+ $X2=3.045 $Y2=1.52
r256 5 7 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=3.045 $Y=1.355
+ $X2=3.045 $Y2=0.805
r257 1 63 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.965 $Y=1.685
+ $X2=2.965 $Y2=1.52
r258 1 3 374.319 $w=1.5e-07 $l=7.3e-07 $layer=POLY_cond $X=2.965 $Y=1.685
+ $X2=2.965 $Y2=2.415
.ends

.subckt PM_SKY130_FD_SC_LP__FA_2%A_395_398# 1 2 3 4 15 19 21 23 26 30 32 35 37
+ 39 40 41 42 48 49 51 52 53 54 58 60 62 68 71 72 73 74 83 90 91 94 104
c270 90 0 7.70653e-20 $X=4.84 $Y=1.77
c271 60 0 8.15636e-20 $X=2.115 $Y=2.135
c272 54 0 7.53306e-20 $X=1.14 $Y=0.965
c273 19 0 2.9941e-19 $X=4.63 $Y=2.415
r274 93 95 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=7.345 $Y=1.38
+ $X2=7.415 $Y2=1.38
r275 93 94 30.474 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=7.345 $Y=1.38
+ $X2=7.27 $Y2=1.38
r276 90 91 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.84
+ $Y=1.77 $X2=4.84 $Y2=1.77
r277 88 90 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=4.63 $Y=1.77
+ $X2=4.84 $Y2=1.77
r278 86 88 0.874306 $w=3.3e-07 $l=5e-09 $layer=POLY_cond $X=4.625 $Y=1.77
+ $X2=4.63 $Y2=1.77
r279 83 104 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=2.035
+ $X2=8.88 $Y2=2.035
r280 81 91 7.04357 $w=4.48e-07 $l=2.65e-07 $layer=LI1_cond $X=4.9 $Y=2.035
+ $X2=4.9 $Y2=1.77
r281 80 81 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=2.035
+ $X2=5.04 $Y2=2.035
r282 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=2.035
+ $X2=0.72 $Y2=2.035
r283 74 80 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.185 $Y=2.035
+ $X2=5.04 $Y2=2.035
r284 73 83 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.735 $Y=2.035
+ $X2=8.88 $Y2=2.035
r285 73 74 4.39356 $w=1.4e-07 $l=3.55e-06 $layer=MET1_cond $X=8.735 $Y=2.035
+ $X2=5.185 $Y2=2.035
r286 72 76 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.865 $Y=2.035
+ $X2=0.72 $Y2=2.035
r287 71 80 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.895 $Y=2.035
+ $X2=5.04 $Y2=2.035
r288 71 72 4.98761 $w=1.4e-07 $l=4.03e-06 $layer=MET1_cond $X=4.895 $Y=2.035
+ $X2=0.865 $Y2=2.035
r289 66 104 24.8861 $w=3.43e-07 $l=7.45e-07 $layer=LI1_cond $X=8.852 $Y=1.245
+ $X2=8.852 $Y2=1.99
r290 62 64 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=2.31 $Y=0.875
+ $X2=2.31 $Y2=0.965
r291 58 77 65.1381 $w=2.28e-07 $l=1.3e-06 $layer=LI1_cond $X=2.02 $Y=2.035
+ $X2=0.72 $Y2=2.035
r292 58 60 3.63458 $w=2.3e-07 $l=1.3e-07 $layer=LI1_cond $X=2.02 $Y=2.035
+ $X2=2.15 $Y2=2.035
r293 54 56 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=1.14 $Y=0.965
+ $X2=1.14 $Y2=1.16
r294 53 77 1.75372 $w=2.28e-07 $l=3.5e-08 $layer=LI1_cond $X=0.685 $Y=2.035
+ $X2=0.72 $Y2=2.035
r295 51 66 2.83935 $w=3.43e-07 $l=8.5e-08 $layer=LI1_cond $X=8.852 $Y=1.16
+ $X2=8.852 $Y2=1.245
r296 51 68 6.68083 $w=3.43e-07 $l=2e-07 $layer=LI1_cond $X=8.852 $Y=1.16
+ $X2=8.852 $Y2=0.96
r297 51 52 67.5241 $w=1.68e-07 $l=1.035e-06 $layer=LI1_cond $X=8.68 $Y=1.16
+ $X2=7.645 $Y2=1.16
r298 49 95 25.3549 $w=3.3e-07 $l=1.45e-07 $layer=POLY_cond $X=7.56 $Y=1.38
+ $X2=7.415 $Y2=1.38
r299 48 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.56
+ $Y=1.38 $X2=7.56 $Y2=1.38
r300 46 52 6.82373 $w=1.7e-07 $l=1.25499e-07 $layer=LI1_cond $X=7.555 $Y=1.245
+ $X2=7.645 $Y2=1.16
r301 46 48 8.31818 $w=1.78e-07 $l=1.35e-07 $layer=LI1_cond $X=7.555 $Y=1.245
+ $X2=7.555 $Y2=1.38
r302 43 54 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.225 $Y=0.965
+ $X2=1.14 $Y2=0.965
r303 42 64 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.145 $Y=0.965
+ $X2=2.31 $Y2=0.965
r304 42 43 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=2.145 $Y=0.965
+ $X2=1.225 $Y2=0.965
r305 40 56 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.055 $Y=1.16
+ $X2=1.14 $Y2=1.16
r306 40 41 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=1.055 $Y=1.16
+ $X2=0.685 $Y2=1.16
r307 39 53 6.94918 $w=2.3e-07 $l=1.53542e-07 $layer=LI1_cond $X=0.595 $Y=1.92
+ $X2=0.685 $Y2=2.035
r308 38 41 6.82373 $w=1.7e-07 $l=1.25499e-07 $layer=LI1_cond $X=0.595 $Y=1.245
+ $X2=0.685 $Y2=1.16
r309 38 39 41.5909 $w=1.78e-07 $l=6.75e-07 $layer=LI1_cond $X=0.595 $Y=1.245
+ $X2=0.595 $Y2=1.92
r310 33 95 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.415 $Y=1.545
+ $X2=7.415 $Y2=1.38
r311 33 35 471.745 $w=1.5e-07 $l=9.2e-07 $layer=POLY_cond $X=7.415 $Y=1.545
+ $X2=7.415 $Y2=2.465
r312 30 93 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.345 $Y=1.215
+ $X2=7.345 $Y2=1.38
r313 30 32 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=7.345 $Y=1.215
+ $X2=7.345 $Y2=0.685
r314 29 37 5.30422 $w=1.5e-07 $l=1.1e-07 $layer=POLY_cond $X=7.06 $Y=1.29
+ $X2=6.95 $Y2=1.29
r315 29 94 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=7.06 $Y=1.29
+ $X2=7.27 $Y2=1.29
r316 24 37 20.4101 $w=1.5e-07 $l=9.08295e-08 $layer=POLY_cond $X=6.985 $Y=1.365
+ $X2=6.95 $Y2=1.29
r317 24 26 564.043 $w=1.5e-07 $l=1.1e-06 $layer=POLY_cond $X=6.985 $Y=1.365
+ $X2=6.985 $Y2=2.465
r318 21 37 20.4101 $w=1.5e-07 $l=9.08295e-08 $layer=POLY_cond $X=6.915 $Y=1.215
+ $X2=6.95 $Y2=1.29
r319 21 23 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=6.915 $Y=1.215
+ $X2=6.915 $Y2=0.685
r320 17 88 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.63 $Y=1.935
+ $X2=4.63 $Y2=1.77
r321 17 19 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=4.63 $Y=1.935
+ $X2=4.63 $Y2=2.415
r322 13 86 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.625 $Y=1.605
+ $X2=4.625 $Y2=1.77
r323 13 15 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=4.625 $Y=1.605
+ $X2=4.625 $Y2=0.805
r324 4 104 300 $w=1.7e-07 $l=2.24499e-07 $layer=licon1_PDIFF $count=2 $X=8.625
+ $Y=1.835 $X2=8.785 $Y2=1.99
r325 3 60 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=1.975
+ $Y=1.99 $X2=2.115 $Y2=2.135
r326 2 68 182 $w=1.7e-07 $l=3.745e-07 $layer=licon1_NDIFF $count=1 $X=8.625
+ $Y=0.685 $X2=8.86 $Y2=0.96
r327 1 62 182 $w=1.7e-07 $l=2.81425e-07 $layer=licon1_NDIFF $count=1 $X=2.17
+ $Y=0.655 $X2=2.31 $Y2=0.875
.ends

.subckt PM_SKY130_FD_SC_LP__FA_2%CIN 3 7 10 11 12 15 18 19 23 28 29 32 34 42
c110 3 0 8.15636e-20 $X=1.9 $Y=2.31
r111 40 42 29.7264 $w=3.3e-07 $l=1.7e-07 $layer=POLY_cond $X=2.24 $Y=1.665
+ $X2=2.41 $Y2=1.665
r112 38 40 25.3549 $w=3.3e-07 $l=1.45e-07 $layer=POLY_cond $X=2.095 $Y=1.665
+ $X2=2.24 $Y2=1.665
r113 36 38 34.0979 $w=3.3e-07 $l=1.95e-07 $layer=POLY_cond $X=1.9 $Y=1.665
+ $X2=2.095 $Y2=1.665
r114 34 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.24
+ $Y=1.665 $X2=2.24 $Y2=1.665
r115 30 32 120.5 $w=1.5e-07 $l=2.35e-07 $layer=POLY_cond $X=5.055 $Y=1.29
+ $X2=5.29 $Y2=1.29
r116 26 28 274.33 $w=1.5e-07 $l=5.35e-07 $layer=POLY_cond $X=5.29 $Y=3.075
+ $X2=5.29 $Y2=2.54
r117 25 32 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.29 $Y=1.365
+ $X2=5.29 $Y2=1.29
r118 25 28 602.5 $w=1.5e-07 $l=1.175e-06 $layer=POLY_cond $X=5.29 $Y=1.365
+ $X2=5.29 $Y2=2.54
r119 21 30 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.055 $Y=1.215
+ $X2=5.055 $Y2=1.29
r120 21 23 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=5.055 $Y=1.215
+ $X2=5.055 $Y2=0.805
r121 20 29 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.27 $Y=3.15
+ $X2=4.195 $Y2=3.15
r122 19 26 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.215 $Y=3.15
+ $X2=5.29 $Y2=3.075
r123 19 20 484.564 $w=1.5e-07 $l=9.45e-07 $layer=POLY_cond $X=5.215 $Y=3.15
+ $X2=4.27 $Y2=3.15
r124 15 18 825.553 $w=1.5e-07 $l=1.61e-06 $layer=POLY_cond $X=4.195 $Y=0.805
+ $X2=4.195 $Y2=2.415
r125 13 29 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.195 $Y=3.075
+ $X2=4.195 $Y2=3.15
r126 13 18 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.195 $Y=3.075
+ $X2=4.195 $Y2=2.415
r127 11 29 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.12 $Y=3.15
+ $X2=4.195 $Y2=3.15
r128 11 12 838.372 $w=1.5e-07 $l=1.635e-06 $layer=POLY_cond $X=4.12 $Y=3.15
+ $X2=2.485 $Y2=3.15
r129 10 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.41 $Y=3.075
+ $X2=2.485 $Y2=3.15
r130 9 42 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.41 $Y=1.83
+ $X2=2.41 $Y2=1.665
r131 9 10 638.394 $w=1.5e-07 $l=1.245e-06 $layer=POLY_cond $X=2.41 $Y=1.83
+ $X2=2.41 $Y2=3.075
r132 5 38 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.095 $Y=1.5
+ $X2=2.095 $Y2=1.665
r133 5 7 325.606 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.095 $Y=1.5
+ $X2=2.095 $Y2=0.865
r134 1 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.9 $Y=1.83 $X2=1.9
+ $Y2=1.665
r135 1 3 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.9 $Y=1.83 $X2=1.9
+ $Y2=2.31
.ends

.subckt PM_SKY130_FD_SC_LP__FA_2%B 3 5 7 8 11 13 15 17 19 24 28 31 33 35 36 39
+ 41 42 48 54 58
c167 19 0 7.37335e-20 $X=5.76 $Y=2.54
c168 11 0 1.39673e-19 $X=3.835 $Y=0.805
c169 3 0 1.63187e-19 $X=1.47 $Y=0.865
r170 55 58 8.83531 $w=4.38e-07 $l=1.65e-07 $layer=LI1_cond $X=8.665 $Y=0.475
+ $X2=8.5 $Y2=0.475
r171 54 55 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.665
+ $Y=0.41 $X2=8.665 $Y2=0.41
r172 51 54 20.109 $w=3.3e-07 $l=1.15e-07 $layer=POLY_cond $X=8.55 $Y=0.41
+ $X2=8.665 $Y2=0.41
r173 48 55 5.63126 $w=4.38e-07 $l=2.15e-07 $layer=LI1_cond $X=8.88 $Y=0.475
+ $X2=8.665 $Y2=0.475
r174 45 46 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.74
+ $Y=1.5 $X2=5.74 $Y2=1.5
r175 42 45 3.54598 $w=2.58e-07 $l=8e-08 $layer=LI1_cond $X=5.775 $Y=1.42
+ $X2=5.775 $Y2=1.5
r176 41 58 117.759 $w=1.68e-07 $l=1.805e-06 $layer=LI1_cond $X=6.695 $Y=0.61
+ $X2=8.5 $Y2=0.61
r177 38 41 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.61 $Y=0.695
+ $X2=6.695 $Y2=0.61
r178 38 39 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=6.61 $Y=0.695
+ $X2=6.61 $Y2=1.335
r179 37 42 3.22376 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=5.905 $Y=1.42
+ $X2=5.775 $Y2=1.42
r180 36 39 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.525 $Y=1.42
+ $X2=6.61 $Y2=1.335
r181 36 37 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=6.525 $Y=1.42
+ $X2=5.905 $Y2=1.42
r182 34 35 58.3064 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=8.565 $Y=1.215
+ $X2=8.565 $Y2=1.365
r183 31 35 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=8.55 $Y=2.155
+ $X2=8.55 $Y2=1.365
r184 28 34 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=8.55 $Y=0.895
+ $X2=8.55 $Y2=1.215
r185 25 51 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.55 $Y=0.575
+ $X2=8.55 $Y2=0.41
r186 25 28 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=8.55 $Y=0.575
+ $X2=8.55 $Y2=0.895
r187 22 46 76.7137 $w=2.68e-07 $l=4.24264e-07 $layer=POLY_cond $X=5.86 $Y=1.125
+ $X2=5.755 $Y2=1.5
r188 22 24 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=5.86 $Y=1.125
+ $X2=5.86 $Y2=0.805
r189 21 24 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=5.86 $Y=0.255
+ $X2=5.86 $Y2=0.805
r190 17 46 38.945 $w=2.68e-07 $l=1.67481e-07 $layer=POLY_cond $X=5.76 $Y=1.665
+ $X2=5.755 $Y2=1.5
r191 17 19 448.67 $w=1.5e-07 $l=8.75e-07 $layer=POLY_cond $X=5.76 $Y=1.665
+ $X2=5.76 $Y2=2.54
r192 16 33 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.91 $Y=0.18
+ $X2=3.835 $Y2=0.18
r193 15 21 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.785 $Y=0.18
+ $X2=5.86 $Y2=0.255
r194 15 16 961.436 $w=1.5e-07 $l=1.875e-06 $layer=POLY_cond $X=5.785 $Y=0.18
+ $X2=3.91 $Y2=0.18
r195 11 13 825.553 $w=1.5e-07 $l=1.61e-06 $layer=POLY_cond $X=3.835 $Y=0.805
+ $X2=3.835 $Y2=2.415
r196 9 33 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.835 $Y=0.255
+ $X2=3.835 $Y2=0.18
r197 9 11 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=3.835 $Y=0.255
+ $X2=3.835 $Y2=0.805
r198 7 33 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.76 $Y=0.18
+ $X2=3.835 $Y2=0.18
r199 7 8 1135.78 $w=1.5e-07 $l=2.215e-06 $layer=POLY_cond $X=3.76 $Y=0.18
+ $X2=1.545 $Y2=0.18
r200 3 5 740.947 $w=1.5e-07 $l=1.445e-06 $layer=POLY_cond $X=1.47 $Y=0.865
+ $X2=1.47 $Y2=2.31
r201 1 8 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.47 $Y=0.255
+ $X2=1.545 $Y2=0.18
r202 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.47 $Y=0.255
+ $X2=1.47 $Y2=0.865
.ends

.subckt PM_SKY130_FD_SC_LP__FA_2%VPWR 1 2 3 4 5 6 19 21 25 31 35 39 43 46 47 48
+ 50 55 60 68 81 82 88 91 94 97
r129 97 98 6.15565 $w=6.93e-07 $l=1.65e-07 $layer=LI1_cond $X=6.587 $Y=2.83
+ $X2=6.587 $Y2=2.665
r130 94 95 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r131 91 92 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r132 88 89 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r133 85 86 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r134 81 82 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r135 79 82 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=8.88 $Y2=3.33
r136 78 81 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=7.92 $Y=3.33
+ $X2=8.88 $Y2=3.33
r137 78 79 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r138 76 79 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=7.92 $Y2=3.33
r139 76 101 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=6.48 $Y2=3.33
r140 75 76 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r141 73 75 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=6.935 $Y=3.33
+ $X2=7.44 $Y2=3.33
r142 72 101 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33
+ $X2=6.48 $Y2=3.33
r143 72 95 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=5.52
+ $Y2=3.33
r144 71 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r145 69 94 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.685 $Y=3.33
+ $X2=5.52 $Y2=3.33
r146 69 71 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=5.685 $Y=3.33
+ $X2=6 $Y2=3.33
r147 68 73 9.27432 $w=1.7e-07 $l=3.48e-07 $layer=LI1_cond $X=6.587 $Y=3.33
+ $X2=6.935 $Y2=3.33
r148 68 101 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r149 68 97 8.60488 $w=6.93e-07 $l=5e-07 $layer=LI1_cond $X=6.587 $Y=3.33
+ $X2=6.587 $Y2=2.83
r150 68 71 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=6.24 $Y=3.33 $X2=6
+ $Y2=3.33
r151 67 95 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=5.52 $Y2=3.33
r152 66 67 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r153 64 92 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=3.12 $Y2=3.33
r154 63 66 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=3.6 $Y=3.33
+ $X2=5.04 $Y2=3.33
r155 63 64 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r156 61 91 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.425 $Y=3.33
+ $X2=3.26 $Y2=3.33
r157 61 63 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=3.425 $Y=3.33
+ $X2=3.6 $Y2=3.33
r158 60 94 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.355 $Y=3.33
+ $X2=5.52 $Y2=3.33
r159 60 66 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=5.355 $Y=3.33
+ $X2=5.04 $Y2=3.33
r160 59 92 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=3.12 $Y2=3.33
r161 59 89 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r162 58 59 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r163 56 88 9.39981 $w=1.7e-07 $l=1.88e-07 $layer=LI1_cond $X=1.35 $Y=3.33
+ $X2=1.162 $Y2=3.33
r164 56 58 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=1.35 $Y=3.33
+ $X2=1.68 $Y2=3.33
r165 55 91 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.095 $Y=3.33
+ $X2=3.26 $Y2=3.33
r166 55 58 92.3155 $w=1.68e-07 $l=1.415e-06 $layer=LI1_cond $X=3.095 $Y=3.33
+ $X2=1.68 $Y2=3.33
r167 54 89 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r168 54 86 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r169 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r170 51 85 4.73185 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=3.33
+ $X2=0.222 $Y2=3.33
r171 51 53 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.445 $Y=3.33
+ $X2=0.72 $Y2=3.33
r172 50 88 9.39981 $w=1.7e-07 $l=1.87e-07 $layer=LI1_cond $X=0.975 $Y=3.33
+ $X2=1.162 $Y2=3.33
r173 50 53 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.975 $Y=3.33
+ $X2=0.72 $Y2=3.33
r174 48 67 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.04 $Y2=3.33
r175 48 64 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=3.6 $Y2=3.33
r176 46 75 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=7.465 $Y=3.33
+ $X2=7.44 $Y2=3.33
r177 46 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.465 $Y=3.33
+ $X2=7.63 $Y2=3.33
r178 45 78 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=7.795 $Y=3.33
+ $X2=7.92 $Y2=3.33
r179 45 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.795 $Y=3.33
+ $X2=7.63 $Y2=3.33
r180 41 47 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.63 $Y=3.245
+ $X2=7.63 $Y2=3.33
r181 41 43 15.8897 $w=3.28e-07 $l=4.55e-07 $layer=LI1_cond $X=7.63 $Y=3.245
+ $X2=7.63 $Y2=2.79
r182 39 98 10.826 $w=3.28e-07 $l=3.1e-07 $layer=LI1_cond $X=6.405 $Y=2.355
+ $X2=6.405 $Y2=2.665
r183 33 94 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.52 $Y=3.245
+ $X2=5.52 $Y2=3.33
r184 33 35 17.8105 $w=3.28e-07 $l=5.1e-07 $layer=LI1_cond $X=5.52 $Y=3.245
+ $X2=5.52 $Y2=2.735
r185 29 91 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.26 $Y=3.245
+ $X2=3.26 $Y2=3.33
r186 29 31 34.7479 $w=3.28e-07 $l=9.95e-07 $layer=LI1_cond $X=3.26 $Y=3.245
+ $X2=3.26 $Y2=2.25
r187 25 28 16.1342 $w=3.73e-07 $l=5.25e-07 $layer=LI1_cond $X=1.162 $Y=2.425
+ $X2=1.162 $Y2=2.95
r188 23 88 1.28102 $w=3.75e-07 $l=8.5e-08 $layer=LI1_cond $X=1.162 $Y=3.245
+ $X2=1.162 $Y2=3.33
r189 23 28 9.06588 $w=3.73e-07 $l=2.95e-07 $layer=LI1_cond $X=1.162 $Y=3.245
+ $X2=1.162 $Y2=2.95
r190 19 85 3.03433 $w=3.3e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.222 $Y2=3.33
r191 19 21 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.28 $Y2=2.825
r192 6 43 600 $w=1.7e-07 $l=1.02261e-06 $layer=licon1_PDIFF $count=1 $X=7.49
+ $Y=1.835 $X2=7.63 $Y2=2.79
r193 5 97 600 $w=1.7e-07 $l=8.24712e-07 $layer=licon1_PDIFF $count=1 $X=6.265
+ $Y=2.22 $X2=6.77 $Y2=2.83
r194 5 39 300 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_PDIFF $count=2 $X=6.265
+ $Y=2.22 $X2=6.405 $Y2=2.355
r195 4 35 600 $w=1.7e-07 $l=5.8741e-07 $layer=licon1_PDIFF $count=1 $X=5.365
+ $Y=2.22 $X2=5.52 $Y2=2.735
r196 3 31 300 $w=1.7e-07 $l=2.87228e-07 $layer=licon1_PDIFF $count=2 $X=3.04
+ $Y=2.095 $X2=3.26 $Y2=2.25
r197 2 28 600 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=1
+ $Y=1.835 $X2=1.14 $Y2=2.95
r198 2 25 600 $w=1.7e-07 $l=6.76203e-07 $layer=licon1_PDIFF $count=1 $X=1
+ $Y=1.835 $X2=1.185 $Y2=2.425
r199 1 21 600 $w=1.7e-07 $l=1.05064e-06 $layer=licon1_PDIFF $count=1 $X=0.155
+ $Y=1.835 $X2=0.28 $Y2=2.825
.ends

.subckt PM_SKY130_FD_SC_LP__FA_2%SUM 1 2 7 9 13 18 19 20 21 22 23 31 34
c50 13 0 1.63187e-19 $X=0.71 $Y=0.38
r51 31 34 0.921954 $w=2.48e-07 $l=2e-08 $layer=LI1_cond $X=0.21 $Y=0.905
+ $X2=0.21 $Y2=0.925
r52 22 23 9.69311 $w=4.18e-07 $l=2.85e-07 $layer=LI1_cond $X=0.21 $Y=2.035
+ $X2=0.21 $Y2=2.32
r53 21 22 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=0.21 $Y=1.665
+ $X2=0.21 $Y2=2.035
r54 20 21 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=0.21 $Y=1.295
+ $X2=0.21 $Y2=1.665
r55 19 31 2.95288 $w=2.5e-07 $l=9e-08 $layer=LI1_cond $X=0.21 $Y=0.815 $X2=0.21
+ $Y2=0.905
r56 19 20 15.581 $w=2.48e-07 $l=3.38e-07 $layer=LI1_cond $X=0.21 $Y=0.957
+ $X2=0.21 $Y2=1.295
r57 19 34 1.47513 $w=2.48e-07 $l=3.2e-08 $layer=LI1_cond $X=0.21 $Y=0.957
+ $X2=0.21 $Y2=0.925
r58 11 13 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=0.71 $Y=0.725
+ $X2=0.71 $Y2=0.38
r59 10 23 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.335 $Y=2.405
+ $X2=0.21 $Y2=2.405
r60 9 18 3.61205 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=0.615 $Y=2.405
+ $X2=0.71 $Y2=2.405
r61 9 10 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=0.615 $Y=2.405
+ $X2=0.335 $Y2=2.405
r62 8 19 4.10122 $w=1.8e-07 $l=1.25e-07 $layer=LI1_cond $X=0.335 $Y=0.815
+ $X2=0.21 $Y2=0.815
r63 7 11 7.61292 $w=1.8e-07 $l=2.05122e-07 $layer=LI1_cond $X=0.545 $Y=0.815
+ $X2=0.71 $Y2=0.725
r64 7 8 12.9394 $w=1.78e-07 $l=2.1e-07 $layer=LI1_cond $X=0.545 $Y=0.815
+ $X2=0.335 $Y2=0.815
r65 2 18 300 $w=1.7e-07 $l=7.16589e-07 $layer=licon1_PDIFF $count=2 $X=0.57
+ $Y=1.835 $X2=0.71 $Y2=2.485
r66 1 13 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=0.57
+ $Y=0.235 $X2=0.71 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_LP__FA_2%A_309_398# 1 2 9 11 12 15
c32 11 0 3.16332e-20 $X=2.585 $Y=2.905
c33 9 0 1.55518e-19 $X=1.685 $Y=2.425
r34 13 15 19.9058 $w=3.28e-07 $l=5.7e-07 $layer=LI1_cond $X=2.75 $Y=2.82
+ $X2=2.75 $Y2=2.25
r35 11 13 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.585 $Y=2.905
+ $X2=2.75 $Y2=2.82
r36 11 12 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=2.585 $Y=2.905
+ $X2=1.85 $Y2=2.905
r37 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.685 $Y=2.82
+ $X2=1.85 $Y2=2.905
r38 7 9 13.7944 $w=3.28e-07 $l=3.95e-07 $layer=LI1_cond $X=1.685 $Y=2.82
+ $X2=1.685 $Y2=2.425
r39 2 15 300 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_PDIFF $count=2 $X=2.625
+ $Y=2.095 $X2=2.75 $Y2=2.25
r40 1 9 600 $w=1.7e-07 $l=5.00125e-07 $layer=licon1_PDIFF $count=1 $X=1.545
+ $Y=1.99 $X2=1.685 $Y2=2.425
.ends

.subckt PM_SKY130_FD_SC_LP__FA_2%A_941_419# 1 2 9 11 13 16
c36 13 0 1.43669e-19 $X=5.975 $Y=2.705
r37 11 18 3.25649 $w=2.15e-07 $l=1.45585e-07 $layer=LI1_cond $X=5.962 $Y=2.47
+ $X2=5.94 $Y2=2.335
r38 11 13 12.5965 $w=2.13e-07 $l=2.35e-07 $layer=LI1_cond $X=5.962 $Y=2.47
+ $X2=5.962 $Y2=2.705
r39 10 16 4.92601 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=5.125 $Y=2.38
+ $X2=4.96 $Y2=2.38
r40 9 18 3.62984 $w=1.8e-07 $l=1.50831e-07 $layer=LI1_cond $X=5.81 $Y=2.38
+ $X2=5.94 $Y2=2.335
r41 9 10 42.2071 $w=1.78e-07 $l=6.85e-07 $layer=LI1_cond $X=5.81 $Y=2.38
+ $X2=5.125 $Y2=2.38
r42 2 18 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=5.835
+ $Y=2.22 $X2=5.975 $Y2=2.365
r43 2 13 600 $w=1.7e-07 $l=5.50568e-07 $layer=licon1_PDIFF $count=1 $X=5.835
+ $Y=2.22 $X2=5.975 $Y2=2.705
r44 1 16 300 $w=1.7e-07 $l=3.8704e-07 $layer=licon1_PDIFF $count=2 $X=4.705
+ $Y=2.095 $X2=4.96 $Y2=2.375
.ends

.subckt PM_SKY130_FD_SC_LP__FA_2%COUT 1 2 7 8 13 18
r32 18 20 14.0769 $w=2.73e-07 $l=3.15e-07 $layer=LI1_cond $X=7.115 $Y=1.665
+ $X2=7.115 $Y2=1.98
r33 11 18 5.30813 $w=4.3e-07 $l=1.46458e-07 $layer=LI1_cond $X=7.08 $Y=1.535
+ $X2=7.115 $Y2=1.665
r34 8 18 3.50848 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=6.96 $Y=1.665
+ $X2=7.115 $Y2=1.665
r35 7 11 6.43224 $w=4.28e-07 $l=2.4e-07 $layer=LI1_cond $X=7.08 $Y=1.295
+ $X2=7.08 $Y2=1.535
r36 7 13 8.71033 $w=4.28e-07 $l=3.25e-07 $layer=LI1_cond $X=7.08 $Y=1.295
+ $X2=7.08 $Y2=0.97
r37 2 20 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=7.06
+ $Y=1.835 $X2=7.2 $Y2=1.98
r38 1 13 182 $w=1.7e-07 $l=7.71832e-07 $layer=licon1_NDIFF $count=1 $X=6.99
+ $Y=0.265 $X2=7.13 $Y2=0.97
.ends

.subckt PM_SKY130_FD_SC_LP__FA_2%VGND 1 2 3 4 5 6 19 21 25 29 33 35 38 39 40 41
+ 47 49 61 76 77 83 86 90
c107 25 0 1.80747e-19 $X=1.16 $Y=0.545
r108 90 93 9.07985 $w=3.28e-07 $l=2.6e-07 $layer=LI1_cond $X=6.62 $Y=0 $X2=6.62
+ $Y2=0.26
r109 90 91 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r110 87 91 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=6.48
+ $Y2=0
r111 86 87 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r112 83 84 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r113 80 81 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r114 76 77 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.88 $Y=0 $X2=8.88
+ $Y2=0
r115 74 77 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=8.88
+ $Y2=0
r116 73 76 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=7.92 $Y=0 $X2=8.88
+ $Y2=0
r117 73 74 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r118 71 74 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0 $X2=7.92
+ $Y2=0
r119 71 91 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.44 $Y=0 $X2=6.48
+ $Y2=0
r120 70 71 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r121 68 90 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.785 $Y=0 $X2=6.62
+ $Y2=0
r122 68 70 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=6.785 $Y=0
+ $X2=7.44 $Y2=0
r123 67 87 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=5.52
+ $Y2=0
r124 66 67 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r125 63 66 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=3.6 $Y=0 $X2=5.04
+ $Y2=0
r126 63 64 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r127 61 86 13.7128 $w=1.7e-07 $l=3.52e-07 $layer=LI1_cond $X=5.105 $Y=0
+ $X2=5.457 $Y2=0
r128 61 66 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=5.105 $Y=0 $X2=5.04
+ $Y2=0
r129 60 64 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r130 59 60 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r131 57 60 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.68 $Y=0
+ $X2=3.12 $Y2=0
r132 57 84 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r133 56 59 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.68 $Y=0 $X2=3.12
+ $Y2=0
r134 56 57 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r135 54 83 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=1.325 $Y=0 $X2=1.185
+ $Y2=0
r136 54 56 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=1.325 $Y=0
+ $X2=1.68 $Y2=0
r137 53 84 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r138 53 81 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r139 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r140 50 80 4.09637 $w=1.7e-07 $l=1.88e-07 $layer=LI1_cond $X=0.375 $Y=0
+ $X2=0.187 $Y2=0
r141 50 52 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.375 $Y=0 $X2=0.72
+ $Y2=0
r142 49 83 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=1.045 $Y=0 $X2=1.185
+ $Y2=0
r143 49 52 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=1.045 $Y=0
+ $X2=0.72 $Y2=0
r144 47 67 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.04
+ $Y2=0
r145 47 64 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=3.6
+ $Y2=0
r146 43 73 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=7.805 $Y=0
+ $X2=7.92 $Y2=0
r147 41 70 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=7.475 $Y=0 $X2=7.44
+ $Y2=0
r148 40 45 9.07985 $w=3.28e-07 $l=2.6e-07 $layer=LI1_cond $X=7.64 $Y=0 $X2=7.64
+ $Y2=0.26
r149 40 43 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.64 $Y=0 $X2=7.805
+ $Y2=0
r150 40 41 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.64 $Y=0 $X2=7.475
+ $Y2=0
r151 38 59 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=3.165 $Y=0 $X2=3.12
+ $Y2=0
r152 38 39 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=3.165 $Y=0 $X2=3.27
+ $Y2=0
r153 37 63 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=3.375 $Y=0 $X2=3.6
+ $Y2=0
r154 37 39 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=3.375 $Y=0 $X2=3.27
+ $Y2=0
r155 36 86 13.7128 $w=1.7e-07 $l=3.53e-07 $layer=LI1_cond $X=5.81 $Y=0 $X2=5.457
+ $Y2=0
r156 35 90 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.455 $Y=0 $X2=6.62
+ $Y2=0
r157 35 36 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=6.455 $Y=0
+ $X2=5.81 $Y2=0
r158 31 86 2.87722 $w=7.05e-07 $l=8.5e-08 $layer=LI1_cond $X=5.457 $Y=0.085
+ $X2=5.457 $Y2=0
r159 31 33 11.1125 $w=7.03e-07 $l=6.55e-07 $layer=LI1_cond $X=5.457 $Y=0.085
+ $X2=5.457 $Y2=0.74
r160 27 39 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=3.27 $Y=0.085
+ $X2=3.27 $Y2=0
r161 27 29 35.1212 $w=2.08e-07 $l=6.65e-07 $layer=LI1_cond $X=3.27 $Y=0.085
+ $X2=3.27 $Y2=0.75
r162 23 83 0.375625 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=1.185 $Y=0.085
+ $X2=1.185 $Y2=0
r163 23 25 18.933 $w=2.78e-07 $l=4.6e-07 $layer=LI1_cond $X=1.185 $Y=0.085
+ $X2=1.185 $Y2=0.545
r164 19 80 3.11585 $w=2.6e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.245 $Y=0.085
+ $X2=0.187 $Y2=0
r165 19 21 13.519 $w=2.58e-07 $l=3.05e-07 $layer=LI1_cond $X=0.245 $Y=0.085
+ $X2=0.245 $Y2=0.39
r166 6 45 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=7.42
+ $Y=0.265 $X2=7.64 $Y2=0.26
r167 5 93 182 $w=1.7e-07 $l=4.44578e-07 $layer=licon1_NDIFF $count=1 $X=6.365
+ $Y=0.595 $X2=6.62 $Y2=0.26
r168 4 33 91 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_NDIFF $count=2 $X=5.13
+ $Y=0.595 $X2=5.645 $Y2=0.74
r169 3 29 182 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=1 $X=3.12
+ $Y=0.595 $X2=3.26 $Y2=0.75
r170 2 25 182 $w=1.7e-07 $l=3.81707e-07 $layer=licon1_NDIFF $count=1 $X=1
+ $Y=0.235 $X2=1.16 $Y2=0.545
r171 1 21 182 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=1 $X=0.155
+ $Y=0.235 $X2=0.28 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_LP__FA_2%A_309_131# 1 2 7 11 13
r26 13 16 5.5876 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=1.8 $Y=0.455 $X2=1.8
+ $Y2=0.615
r27 9 11 9.25447 $w=3.28e-07 $l=2.65e-07 $layer=LI1_cond $X=2.83 $Y=0.54
+ $X2=2.83 $Y2=0.805
r28 8 13 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.965 $Y=0.455
+ $X2=1.8 $Y2=0.455
r29 7 9 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.665 $Y=0.455
+ $X2=2.83 $Y2=0.54
r30 7 8 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=2.665 $Y=0.455 $X2=1.965
+ $Y2=0.455
r31 2 11 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=2.705
+ $Y=0.595 $X2=2.83 $Y2=0.805
r32 1 16 182 $w=1.7e-07 $l=2.74272e-07 $layer=licon1_NDIFF $count=1 $X=1.545
+ $Y=0.655 $X2=1.8 $Y2=0.615
.ends

.subckt PM_SKY130_FD_SC_LP__FA_2%A_940_119# 1 2 9 11 12 15
r20 13 15 6.93182 $w=1.98e-07 $l=1.25e-07 $layer=LI1_cond $X=6.08 $Y=0.995
+ $X2=6.08 $Y2=0.87
r21 11 13 6.87494 $w=1.7e-07 $l=1.36015e-07 $layer=LI1_cond $X=5.98 $Y=1.08
+ $X2=6.08 $Y2=0.995
r22 11 12 68.1765 $w=1.68e-07 $l=1.045e-06 $layer=LI1_cond $X=5.98 $Y=1.08
+ $X2=4.935 $Y2=1.08
r23 7 12 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=4.82 $Y=0.995
+ $X2=4.935 $Y2=1.08
r24 7 9 9.52018 $w=2.28e-07 $l=1.9e-07 $layer=LI1_cond $X=4.82 $Y=0.995 $X2=4.82
+ $Y2=0.805
r25 2 15 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=5.935
+ $Y=0.595 $X2=6.075 $Y2=0.87
r26 1 9 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=4.7
+ $Y=0.595 $X2=4.84 $Y2=0.805
.ends

