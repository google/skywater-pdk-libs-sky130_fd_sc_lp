* File: sky130_fd_sc_lp__dlymetal6s2s_1.spice
* Created: Wed Sep  2 09:50:18 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__dlymetal6s2s_1.pex.spice"
.subckt sky130_fd_sc_lp__dlymetal6s2s_1  VNB VPB A X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* A	A
* VPB	VPB
* VNB	VNB
MM1008 N_VGND_M1008_d N_A_M1008_g N_A_27_131#_M1008_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0847 AS=0.1113 PD=0.786667 PS=1.37 NRD=18.564 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1006 N_X_M1006_d N_A_27_131#_M1006_g N_VGND_M1008_d VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1694 PD=2.21 PS=1.57333 NRD=0 NRS=0 M=1 R=5.6 SA=75000.4
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1011 N_VGND_M1011_d N_X_M1011_g N_A_315_131#_M1011_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0847 AS=0.1113 PD=0.786667 PS=1.37 NRD=18.564 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1002 N_A_496_47#_M1002_d N_A_315_131#_M1002_g N_VGND_M1011_d VNB NSHORT L=0.15
+ W=0.84 AD=0.2226 AS=0.1694 PD=2.21 PS=1.57333 NRD=0 NRS=0 M=1 R=5.6 SA=75000.4
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1004 N_VGND_M1004_d N_A_496_47#_M1004_g N_A_603_131#_M1004_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0847 AS=0.1113 PD=0.786667 PS=1.37 NRD=18.564 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1009 N_A_784_47#_M1009_d N_A_603_131#_M1009_g N_VGND_M1004_d VNB NSHORT L=0.15
+ W=0.84 AD=0.2226 AS=0.1694 PD=2.21 PS=1.57333 NRD=0 NRS=0 M=1 R=5.6 SA=75000.4
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1010 N_VPWR_M1010_d N_A_M1010_g N_A_27_131#_M1010_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.09135 AS=0.1113 PD=0.8 PS=1.37 NRD=76.2193 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1001 N_X_M1001_d N_A_27_131#_M1001_g N_VPWR_M1010_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.27405 PD=3.05 PS=2.4 NRD=0 NRS=0 M=1 R=8.4 SA=75000.4
+ SB=75000.2 A=0.189 P=2.82 MULT=1
MM1005 N_VPWR_M1005_d N_X_M1005_g N_A_315_131#_M1005_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.09135 AS=0.1113 PD=0.8 PS=1.37 NRD=76.2193 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1000 N_A_496_47#_M1000_d N_A_315_131#_M1000_g N_VPWR_M1005_d VPB PHIGHVT
+ L=0.15 W=1.26 AD=0.3339 AS=0.27405 PD=3.05 PS=2.4 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.4 SB=75000.2 A=0.189 P=2.82 MULT=1
MM1003 N_VPWR_M1003_d N_A_496_47#_M1003_g N_A_603_131#_M1003_s VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.09135 AS=0.1113 PD=0.8 PS=1.37 NRD=76.2193 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1007 N_A_784_47#_M1007_d N_A_603_131#_M1007_g N_VPWR_M1003_d VPB PHIGHVT
+ L=0.15 W=1.26 AD=0.3339 AS=0.27405 PD=3.05 PS=2.4 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.4 SB=75000.2 A=0.189 P=2.82 MULT=1
DX12_noxref VNB VPB NWDIODE A=8.7655 P=13.13
*
.include "sky130_fd_sc_lp__dlymetal6s2s_1.pxi.spice"
*
.ends
*
*
