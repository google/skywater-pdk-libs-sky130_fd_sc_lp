* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__a311oi_m A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
X0 VPWR A1 a_191_535# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X1 a_199_51# A2 a_271_51# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 Y B1 VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 VGND C1 Y VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 a_191_535# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X5 VPWR A3 a_191_535# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X6 a_449_535# C1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X7 VGND A3 a_199_51# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 a_271_51# A1 Y VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 a_191_535# B1 a_449_535# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
.ends
