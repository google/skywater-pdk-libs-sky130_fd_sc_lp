* File: sky130_fd_sc_lp__o22a_0.pxi.spice
* Created: Fri Aug 28 11:09:15 2020
* 
x_PM_SKY130_FD_SC_LP__O22A_0%A_80_313# N_A_80_313#_M1003_d N_A_80_313#_M1001_d
+ N_A_80_313#_c_91_n N_A_80_313#_M1006_g N_A_80_313#_M1000_g N_A_80_313#_c_93_n
+ N_A_80_313#_c_84_n N_A_80_313#_c_85_n N_A_80_313#_c_95_n N_A_80_313#_c_96_n
+ N_A_80_313#_c_169_p N_A_80_313#_c_86_n N_A_80_313#_c_97_n N_A_80_313#_c_87_n
+ N_A_80_313#_c_88_n N_A_80_313#_c_89_n N_A_80_313#_c_100_n N_A_80_313#_c_101_n
+ N_A_80_313#_c_90_n N_A_80_313#_c_102_n PM_SKY130_FD_SC_LP__O22A_0%A_80_313#
x_PM_SKY130_FD_SC_LP__O22A_0%A1 N_A1_c_208_n N_A1_M1002_g N_A1_M1005_g
+ N_A1_c_209_n N_A1_c_210_n N_A1_c_216_n N_A1_c_217_n N_A1_c_218_n N_A1_c_219_n
+ A1 A1 A1 N_A1_c_211_n N_A1_c_212_n N_A1_c_213_n A1
+ PM_SKY130_FD_SC_LP__O22A_0%A1
x_PM_SKY130_FD_SC_LP__O22A_0%B1 N_B1_M1003_g N_B1_M1007_g N_B1_c_294_n
+ N_B1_c_295_n B1 B1 PM_SKY130_FD_SC_LP__O22A_0%B1
x_PM_SKY130_FD_SC_LP__O22A_0%B2 N_B2_M1001_g N_B2_M1004_g N_B2_c_342_n
+ N_B2_c_347_n B2 B2 N_B2_c_344_n PM_SKY130_FD_SC_LP__O22A_0%B2
x_PM_SKY130_FD_SC_LP__O22A_0%A2 N_A2_c_392_n N_A2_M1009_g N_A2_c_387_n
+ N_A2_M1008_g N_A2_c_388_n N_A2_c_394_n N_A2_c_389_n A2 N_A2_c_391_n
+ PM_SKY130_FD_SC_LP__O22A_0%A2
x_PM_SKY130_FD_SC_LP__O22A_0%X N_X_M1000_s N_X_M1006_s X X X X X X X N_X_c_434_n
+ PM_SKY130_FD_SC_LP__O22A_0%X
x_PM_SKY130_FD_SC_LP__O22A_0%VPWR N_VPWR_M1006_d N_VPWR_M1005_d N_VPWR_c_458_n
+ N_VPWR_c_459_n N_VPWR_c_460_n N_VPWR_c_461_n N_VPWR_c_462_n VPWR
+ N_VPWR_c_463_n N_VPWR_c_464_n N_VPWR_c_457_n N_VPWR_c_466_n
+ PM_SKY130_FD_SC_LP__O22A_0%VPWR
x_PM_SKY130_FD_SC_LP__O22A_0%VGND N_VGND_M1000_d N_VGND_M1008_d N_VGND_c_509_n
+ N_VGND_c_510_n N_VGND_c_519_n VGND N_VGND_c_511_n N_VGND_c_512_n
+ N_VGND_c_513_n N_VGND_c_514_n N_VGND_c_515_n PM_SKY130_FD_SC_LP__O22A_0%VGND
x_PM_SKY130_FD_SC_LP__O22A_0%A_286_125# N_A_286_125#_M1002_d
+ N_A_286_125#_M1004_d N_A_286_125#_c_559_n N_A_286_125#_c_552_n
+ N_A_286_125#_c_553_n N_A_286_125#_c_554_n
+ PM_SKY130_FD_SC_LP__O22A_0%A_286_125#
cc_1 VNB N_A_80_313#_M1000_g 0.0521843f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=0.835
cc_2 VNB N_A_80_313#_c_84_n 2.20794e-19 $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=1.73
cc_3 VNB N_A_80_313#_c_85_n 0.0141364f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=1.73
cc_4 VNB N_A_80_313#_c_86_n 0.006219f $X=-0.19 $Y=-0.245 $X2=2.905 $Y2=1.12
cc_5 VNB N_A_80_313#_c_87_n 0.00397678f $X=-0.19 $Y=-0.245 $X2=2.99 $Y2=1.585
cc_6 VNB N_A_80_313#_c_88_n 0.00900726f $X=-0.19 $Y=-0.245 $X2=3.54 $Y2=1.67
cc_7 VNB N_A_80_313#_c_89_n 4.16132e-19 $X=-0.19 $Y=-0.245 $X2=3.075 $Y2=1.67
cc_8 VNB N_A_80_313#_c_90_n 0.00538771f $X=-0.19 $Y=-0.245 $X2=2.02 $Y2=0.89
cc_9 VNB N_A1_c_208_n 0.017134f $X=-0.19 $Y=-0.245 $X2=1.86 $Y2=0.625
cc_10 VNB N_A1_c_209_n 0.00995212f $X=-0.19 $Y=-0.245 $X2=0.572 $Y2=2.063
cc_11 VNB N_A1_c_210_n 0.00693719f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.765
cc_12 VNB N_A1_c_211_n 0.0623709f $X=-0.19 $Y=-0.245 $X2=3.54 $Y2=2.52
cc_13 VNB N_A1_c_212_n 0.00216559f $X=-0.19 $Y=-0.245 $X2=3.075 $Y2=1.67
cc_14 VNB N_A1_c_213_n 0.00778126f $X=-0.19 $Y=-0.245 $X2=3.642 $Y2=1.755
cc_15 VNB A1 0.0015732f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=2.15
cc_16 VNB N_B1_M1003_g 0.03797f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_B1_c_294_n 0.0302668f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.235
cc_18 VNB N_B1_c_295_n 0.00306581f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.765
cc_19 VNB B1 0.00254083f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.765
cc_20 VNB N_B2_M1004_g 0.0235f $X=-0.19 $Y=-0.245 $X2=0.572 $Y2=1.737
cc_21 VNB N_B2_c_342_n 0.0107125f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.765
cc_22 VNB B2 0.00554832f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=0.835
cc_23 VNB N_B2_c_344_n 0.0151434f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=2.065
cc_24 VNB N_A2_c_387_n 0.0181104f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A2_c_388_n 0.00827939f $X=-0.19 $Y=-0.245 $X2=0.572 $Y2=2.063
cc_26 VNB N_A2_c_389_n 0.0110208f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=0.835
cc_27 VNB A2 0.0326281f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=0.835
cc_28 VNB N_A2_c_391_n 0.0802932f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=2.065
cc_29 VNB X 0.0378616f $X=-0.19 $Y=-0.245 $X2=0.572 $Y2=1.737
cc_30 VNB N_X_c_434_n 0.0197266f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VPWR_c_457_n 0.163682f $X=-0.19 $Y=-0.245 $X2=3.54 $Y2=1.67
cc_32 VNB N_VGND_c_509_n 0.0169501f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.765
cc_33 VNB N_VGND_c_510_n 0.0428316f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=1.565
cc_34 VNB N_VGND_c_511_n 0.0537213f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_512_n 0.0223503f $X=-0.19 $Y=-0.245 $X2=2.555 $Y2=2.52
cc_36 VNB N_VGND_c_513_n 0.25821f $X=-0.19 $Y=-0.245 $X2=2.99 $Y2=1.205
cc_37 VNB N_VGND_c_514_n 0.0243387f $X=-0.19 $Y=-0.245 $X2=3.075 $Y2=1.67
cc_38 VNB N_VGND_c_515_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=2.15
cc_39 VNB N_A_286_125#_c_552_n 0.0111239f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.765
cc_40 VNB N_A_286_125#_c_553_n 0.00363339f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_286_125#_c_554_n 0.00419926f $X=-0.19 $Y=-0.245 $X2=0.575
+ $Y2=1.565
cc_42 VPB N_A_80_313#_c_91_n 0.0248094f $X=-0.19 $Y=1.655 $X2=0.572 $Y2=2.063
cc_43 VPB N_A_80_313#_M1006_g 0.0283047f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.765
cc_44 VPB N_A_80_313#_c_93_n 0.0188066f $X=-0.19 $Y=1.655 $X2=0.572 $Y2=2.235
cc_45 VPB N_A_80_313#_c_85_n 0.00627891f $X=-0.19 $Y=1.655 $X2=0.58 $Y2=1.73
cc_46 VPB N_A_80_313#_c_95_n 0.00833763f $X=-0.19 $Y=1.655 $X2=0.68 $Y2=2.435
cc_47 VPB N_A_80_313#_c_96_n 0.0146475f $X=-0.19 $Y=1.655 $X2=2.225 $Y2=2.52
cc_48 VPB N_A_80_313#_c_97_n 0.0215754f $X=-0.19 $Y=1.655 $X2=3.54 $Y2=2.52
cc_49 VPB N_A_80_313#_c_88_n 0.013578f $X=-0.19 $Y=1.655 $X2=3.54 $Y2=1.67
cc_50 VPB N_A_80_313#_c_89_n 0.00313636f $X=-0.19 $Y=1.655 $X2=3.075 $Y2=1.67
cc_51 VPB N_A_80_313#_c_100_n 0.0388784f $X=-0.19 $Y=1.655 $X2=3.642 $Y2=2.435
cc_52 VPB N_A_80_313#_c_101_n 0.00196682f $X=-0.19 $Y=1.655 $X2=0.68 $Y2=2.15
cc_53 VPB N_A_80_313#_c_102_n 0.00222846f $X=-0.19 $Y=1.655 $X2=2.39 $Y2=2.59
cc_54 VPB N_A1_M1005_g 0.0238864f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_55 VPB N_A1_c_216_n 0.0177421f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_56 VPB N_A1_c_217_n 0.00281821f $X=-0.19 $Y=1.655 $X2=0.575 $Y2=1.565
cc_57 VPB N_A1_c_218_n 0.00367795f $X=-0.19 $Y=1.655 $X2=0.575 $Y2=0.835
cc_58 VPB N_A1_c_219_n 0.0357019f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_59 VPB N_B1_M1007_g 0.0281956f $X=-0.19 $Y=1.655 $X2=0.572 $Y2=1.737
cc_60 VPB N_B1_c_294_n 0.0771617f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.235
cc_61 VPB N_B1_c_295_n 0.0188876f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.765
cc_62 VPB B1 0.00286261f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.765
cc_63 VPB N_B2_M1001_g 0.0341223f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_64 VPB N_B2_c_342_n 0.00896588f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.765
cc_65 VPB N_B2_c_347_n 0.0148263f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_66 VPB B2 0.00506634f $X=-0.19 $Y=1.655 $X2=0.575 $Y2=0.835
cc_67 VPB N_A2_c_392_n 0.0173881f $X=-0.19 $Y=1.655 $X2=1.86 $Y2=0.625
cc_68 VPB N_A2_c_388_n 0.0314097f $X=-0.19 $Y=1.655 $X2=0.572 $Y2=2.063
cc_69 VPB N_A2_c_394_n 0.0167857f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.765
cc_70 VPB X 0.0381182f $X=-0.19 $Y=1.655 $X2=0.572 $Y2=1.737
cc_71 VPB X 0.00976767f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.765
cc_72 VPB X 0.0191418f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_73 VPB N_VPWR_c_458_n 0.0155155f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.235
cc_74 VPB N_VPWR_c_459_n 0.0100368f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.765
cc_75 VPB N_VPWR_c_460_n 0.0177734f $X=-0.19 $Y=1.655 $X2=0.575 $Y2=0.835
cc_76 VPB N_VPWR_c_461_n 0.0366193f $X=-0.19 $Y=1.655 $X2=0.572 $Y2=2.235
cc_77 VPB N_VPWR_c_462_n 0.0051822f $X=-0.19 $Y=1.655 $X2=0.58 $Y2=2.065
cc_78 VPB N_VPWR_c_463_n 0.0125043f $X=-0.19 $Y=1.655 $X2=2.225 $Y2=2.52
cc_79 VPB N_VPWR_c_464_n 0.0116336f $X=-0.19 $Y=1.655 $X2=2.99 $Y2=1.585
cc_80 VPB N_VPWR_c_457_n 0.0468121f $X=-0.19 $Y=1.655 $X2=3.54 $Y2=1.67
cc_81 VPB N_VPWR_c_466_n 0.00607282f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_82 N_A_80_313#_M1000_g N_A1_c_208_n 0.00600356f $X=0.575 $Y=0.835 $X2=-0.19
+ $Y2=-0.245
cc_83 N_A_80_313#_c_90_n N_A1_c_208_n 4.9641e-19 $X=2.02 $Y=0.89 $X2=-0.19
+ $Y2=-0.245
cc_84 N_A_80_313#_c_97_n N_A1_M1005_g 0.0142038f $X=3.54 $Y=2.52 $X2=0 $Y2=0
cc_85 N_A_80_313#_c_100_n N_A1_M1005_g 0.00498808f $X=3.642 $Y=2.435 $X2=0 $Y2=0
cc_86 N_A_80_313#_c_102_n N_A1_M1005_g 0.00172059f $X=2.39 $Y=2.59 $X2=0 $Y2=0
cc_87 N_A_80_313#_c_96_n N_A1_c_216_n 0.0385225f $X=2.225 $Y=2.52 $X2=0 $Y2=0
cc_88 N_A_80_313#_c_97_n N_A1_c_216_n 0.0365234f $X=3.54 $Y=2.52 $X2=0 $Y2=0
cc_89 N_A_80_313#_c_89_n N_A1_c_216_n 0.0081258f $X=3.075 $Y=1.67 $X2=0 $Y2=0
cc_90 N_A_80_313#_c_102_n N_A1_c_216_n 0.0273204f $X=2.39 $Y=2.59 $X2=0 $Y2=0
cc_91 N_A_80_313#_c_96_n N_A1_c_217_n 0.014356f $X=2.225 $Y=2.52 $X2=0 $Y2=0
cc_92 N_A_80_313#_c_97_n N_A1_c_218_n 0.022705f $X=3.54 $Y=2.52 $X2=0 $Y2=0
cc_93 N_A_80_313#_c_88_n N_A1_c_218_n 0.021227f $X=3.54 $Y=1.67 $X2=0 $Y2=0
cc_94 N_A_80_313#_c_89_n N_A1_c_218_n 0.00114157f $X=3.075 $Y=1.67 $X2=0 $Y2=0
cc_95 N_A_80_313#_c_100_n N_A1_c_218_n 0.0250415f $X=3.642 $Y=2.435 $X2=0 $Y2=0
cc_96 N_A_80_313#_c_97_n N_A1_c_219_n 0.00190976f $X=3.54 $Y=2.52 $X2=0 $Y2=0
cc_97 N_A_80_313#_c_88_n N_A1_c_219_n 0.00155081f $X=3.54 $Y=1.67 $X2=0 $Y2=0
cc_98 N_A_80_313#_c_100_n N_A1_c_219_n 0.00760768f $X=3.642 $Y=2.435 $X2=0 $Y2=0
cc_99 N_A_80_313#_M1000_g N_A1_c_211_n 6.64061e-19 $X=0.575 $Y=0.835 $X2=0 $Y2=0
cc_100 N_A_80_313#_M1000_g N_A1_c_213_n 0.00470519f $X=0.575 $Y=0.835 $X2=0
+ $Y2=0
cc_101 N_A_80_313#_c_90_n N_A1_c_213_n 0.00110287f $X=2.02 $Y=0.89 $X2=0 $Y2=0
cc_102 N_A_80_313#_M1000_g A1 0.00223814f $X=0.575 $Y=0.835 $X2=0 $Y2=0
cc_103 N_A_80_313#_c_90_n A1 0.00470173f $X=2.02 $Y=0.89 $X2=0 $Y2=0
cc_104 N_A_80_313#_c_90_n N_B1_M1003_g 0.00730323f $X=2.02 $Y=0.89 $X2=0 $Y2=0
cc_105 N_A_80_313#_c_96_n N_B1_M1007_g 0.0136814f $X=2.225 $Y=2.52 $X2=0 $Y2=0
cc_106 N_A_80_313#_c_102_n N_B1_M1007_g 0.0016906f $X=2.39 $Y=2.59 $X2=0 $Y2=0
cc_107 N_A_80_313#_c_84_n N_B1_c_294_n 0.00188305f $X=0.58 $Y=1.73 $X2=0 $Y2=0
cc_108 N_A_80_313#_c_85_n N_B1_c_294_n 0.04481f $X=0.58 $Y=1.73 $X2=0 $Y2=0
cc_109 N_A_80_313#_c_96_n N_B1_c_294_n 0.0140272f $X=2.225 $Y=2.52 $X2=0 $Y2=0
cc_110 N_A_80_313#_c_101_n N_B1_c_294_n 0.00123537f $X=0.68 $Y=2.15 $X2=0 $Y2=0
cc_111 N_A_80_313#_c_84_n B1 0.0180403f $X=0.58 $Y=1.73 $X2=0 $Y2=0
cc_112 N_A_80_313#_c_85_n B1 0.0015858f $X=0.58 $Y=1.73 $X2=0 $Y2=0
cc_113 N_A_80_313#_c_96_n B1 0.0203232f $X=2.225 $Y=2.52 $X2=0 $Y2=0
cc_114 N_A_80_313#_c_101_n B1 0.00873722f $X=0.68 $Y=2.15 $X2=0 $Y2=0
cc_115 N_A_80_313#_c_96_n N_B2_M1001_g 0.0085018f $X=2.225 $Y=2.52 $X2=0 $Y2=0
cc_116 N_A_80_313#_c_102_n N_B2_M1001_g 0.00898998f $X=2.39 $Y=2.59 $X2=0 $Y2=0
cc_117 N_A_80_313#_c_86_n N_B2_M1004_g 0.00943894f $X=2.905 $Y=1.12 $X2=0 $Y2=0
cc_118 N_A_80_313#_c_87_n N_B2_M1004_g 3.90743e-19 $X=2.99 $Y=1.585 $X2=0 $Y2=0
cc_119 N_A_80_313#_c_90_n N_B2_M1004_g 0.00769825f $X=2.02 $Y=0.89 $X2=0 $Y2=0
cc_120 N_A_80_313#_c_86_n B2 0.0414856f $X=2.905 $Y=1.12 $X2=0 $Y2=0
cc_121 N_A_80_313#_c_87_n B2 0.0154522f $X=2.99 $Y=1.585 $X2=0 $Y2=0
cc_122 N_A_80_313#_c_89_n B2 0.0151546f $X=3.075 $Y=1.67 $X2=0 $Y2=0
cc_123 N_A_80_313#_c_90_n B2 0.0189693f $X=2.02 $Y=0.89 $X2=0 $Y2=0
cc_124 N_A_80_313#_c_86_n N_B2_c_344_n 0.00339803f $X=2.905 $Y=1.12 $X2=0 $Y2=0
cc_125 N_A_80_313#_c_87_n N_B2_c_344_n 4.12354e-19 $X=2.99 $Y=1.585 $X2=0 $Y2=0
cc_126 N_A_80_313#_c_90_n N_B2_c_344_n 0.00176278f $X=2.02 $Y=0.89 $X2=0 $Y2=0
cc_127 N_A_80_313#_c_97_n N_A2_c_392_n 0.00927326f $X=3.54 $Y=2.52 $X2=-0.19
+ $Y2=-0.245
cc_128 N_A_80_313#_c_102_n N_A2_c_392_n 0.0102328f $X=2.39 $Y=2.59 $X2=-0.19
+ $Y2=-0.245
cc_129 N_A_80_313#_c_86_n N_A2_c_387_n 0.0112593f $X=2.905 $Y=1.12 $X2=0 $Y2=0
cc_130 N_A_80_313#_c_90_n N_A2_c_387_n 6.68528e-19 $X=2.02 $Y=0.89 $X2=0 $Y2=0
cc_131 N_A_80_313#_c_87_n N_A2_c_388_n 0.00209178f $X=2.99 $Y=1.585 $X2=0 $Y2=0
cc_132 N_A_80_313#_c_89_n N_A2_c_388_n 0.003767f $X=3.075 $Y=1.67 $X2=0 $Y2=0
cc_133 N_A_80_313#_c_97_n N_A2_c_394_n 0.00400478f $X=3.54 $Y=2.52 $X2=0 $Y2=0
cc_134 N_A_80_313#_c_86_n N_A2_c_389_n 0.006082f $X=2.905 $Y=1.12 $X2=0 $Y2=0
cc_135 N_A_80_313#_c_86_n A2 0.00771869f $X=2.905 $Y=1.12 $X2=0 $Y2=0
cc_136 N_A_80_313#_c_87_n A2 0.0155095f $X=2.99 $Y=1.585 $X2=0 $Y2=0
cc_137 N_A_80_313#_c_88_n A2 0.0397993f $X=3.54 $Y=1.67 $X2=0 $Y2=0
cc_138 N_A_80_313#_c_86_n N_A2_c_391_n 0.00943709f $X=2.905 $Y=1.12 $X2=0 $Y2=0
cc_139 N_A_80_313#_c_87_n N_A2_c_391_n 0.0178242f $X=2.99 $Y=1.585 $X2=0 $Y2=0
cc_140 N_A_80_313#_c_88_n N_A2_c_391_n 0.0104936f $X=3.54 $Y=1.67 $X2=0 $Y2=0
cc_141 N_A_80_313#_M1000_g X 0.0184063f $X=0.575 $Y=0.835 $X2=0 $Y2=0
cc_142 N_A_80_313#_c_84_n X 0.0366337f $X=0.58 $Y=1.73 $X2=0 $Y2=0
cc_143 N_A_80_313#_c_85_n X 0.0214706f $X=0.58 $Y=1.73 $X2=0 $Y2=0
cc_144 N_A_80_313#_c_95_n X 0.0106009f $X=0.68 $Y=2.435 $X2=0 $Y2=0
cc_145 N_A_80_313#_c_101_n X 0.0128377f $X=0.68 $Y=2.15 $X2=0 $Y2=0
cc_146 N_A_80_313#_M1006_g X 0.00343471f $X=0.475 $Y=2.765 $X2=0 $Y2=0
cc_147 N_A_80_313#_c_95_n X 7.15555e-19 $X=0.68 $Y=2.435 $X2=0 $Y2=0
cc_148 N_A_80_313#_c_169_p X 0.00682015f $X=0.765 $Y=2.52 $X2=0 $Y2=0
cc_149 N_A_80_313#_M1006_g X 0.0109006f $X=0.475 $Y=2.765 $X2=0 $Y2=0
cc_150 N_A_80_313#_M1000_g N_X_c_434_n 4.38513e-19 $X=0.575 $Y=0.835 $X2=0 $Y2=0
cc_151 N_A_80_313#_c_85_n N_X_c_434_n 0.00151548f $X=0.58 $Y=1.73 $X2=0 $Y2=0
cc_152 N_A_80_313#_c_96_n N_VPWR_M1006_d 0.0159395f $X=2.225 $Y=2.52 $X2=-0.19
+ $Y2=-0.245
cc_153 N_A_80_313#_c_169_p N_VPWR_M1006_d 0.00306607f $X=0.765 $Y=2.52 $X2=-0.19
+ $Y2=-0.245
cc_154 N_A_80_313#_c_97_n N_VPWR_M1005_d 0.00290405f $X=3.54 $Y=2.52 $X2=0 $Y2=0
cc_155 N_A_80_313#_c_97_n N_VPWR_c_458_n 0.0211535f $X=3.54 $Y=2.52 $X2=0 $Y2=0
cc_156 N_A_80_313#_c_102_n N_VPWR_c_458_n 0.00757892f $X=2.39 $Y=2.59 $X2=0
+ $Y2=0
cc_157 N_A_80_313#_M1006_g N_VPWR_c_459_n 0.00482245f $X=0.475 $Y=2.765 $X2=0
+ $Y2=0
cc_158 N_A_80_313#_c_93_n N_VPWR_c_459_n 5.18581e-19 $X=0.572 $Y=2.235 $X2=0
+ $Y2=0
cc_159 N_A_80_313#_c_96_n N_VPWR_c_459_n 0.0707605f $X=2.225 $Y=2.52 $X2=0 $Y2=0
cc_160 N_A_80_313#_c_169_p N_VPWR_c_459_n 0.0130203f $X=0.765 $Y=2.52 $X2=0
+ $Y2=0
cc_161 N_A_80_313#_M1006_g N_VPWR_c_460_n 0.00539298f $X=0.475 $Y=2.765 $X2=0
+ $Y2=0
cc_162 N_A_80_313#_c_96_n N_VPWR_c_461_n 0.00603158f $X=2.225 $Y=2.52 $X2=0
+ $Y2=0
cc_163 N_A_80_313#_c_97_n N_VPWR_c_461_n 0.00805425f $X=3.54 $Y=2.52 $X2=0 $Y2=0
cc_164 N_A_80_313#_c_102_n N_VPWR_c_461_n 0.0188581f $X=2.39 $Y=2.59 $X2=0 $Y2=0
cc_165 N_A_80_313#_c_97_n N_VPWR_c_464_n 0.00384571f $X=3.54 $Y=2.52 $X2=0 $Y2=0
cc_166 N_A_80_313#_M1001_d N_VPWR_c_457_n 0.00223559f $X=2.25 $Y=2.445 $X2=0
+ $Y2=0
cc_167 N_A_80_313#_M1006_g N_VPWR_c_457_n 0.0120083f $X=0.475 $Y=2.765 $X2=0
+ $Y2=0
cc_168 N_A_80_313#_c_96_n N_VPWR_c_457_n 0.0155146f $X=2.225 $Y=2.52 $X2=0 $Y2=0
cc_169 N_A_80_313#_c_169_p N_VPWR_c_457_n 7.0054e-19 $X=0.765 $Y=2.52 $X2=0
+ $Y2=0
cc_170 N_A_80_313#_c_97_n N_VPWR_c_457_n 0.0233321f $X=3.54 $Y=2.52 $X2=0 $Y2=0
cc_171 N_A_80_313#_c_102_n N_VPWR_c_457_n 0.0123659f $X=2.39 $Y=2.59 $X2=0 $Y2=0
cc_172 N_A_80_313#_c_102_n N_VPWR_c_466_n 0.0100461f $X=2.39 $Y=2.59 $X2=0 $Y2=0
cc_173 N_A_80_313#_c_96_n A_372_489# 0.00241572f $X=2.225 $Y=2.52 $X2=-0.19
+ $Y2=-0.245
cc_174 N_A_80_313#_c_97_n A_536_489# 0.00527588f $X=3.54 $Y=2.52 $X2=-0.19
+ $Y2=-0.245
cc_175 N_A_80_313#_c_86_n N_VGND_M1008_d 0.00262266f $X=2.905 $Y=1.12 $X2=0
+ $Y2=0
cc_176 N_A_80_313#_M1000_g N_VGND_c_509_n 0.00685449f $X=0.575 $Y=0.835 $X2=0
+ $Y2=0
cc_177 N_A_80_313#_c_86_n N_VGND_c_510_n 0.0176342f $X=2.905 $Y=1.12 $X2=0 $Y2=0
cc_178 N_A_80_313#_M1000_g N_VGND_c_519_n 0.00335494f $X=0.575 $Y=0.835 $X2=0
+ $Y2=0
cc_179 N_A_80_313#_c_84_n N_VGND_c_519_n 3.25389e-19 $X=0.58 $Y=1.73 $X2=0 $Y2=0
cc_180 N_A_80_313#_c_85_n N_VGND_c_519_n 0.00178465f $X=0.58 $Y=1.73 $X2=0 $Y2=0
cc_181 N_A_80_313#_M1000_g N_VGND_c_513_n 0.00456913f $X=0.575 $Y=0.835 $X2=0
+ $Y2=0
cc_182 N_A_80_313#_M1000_g N_VGND_c_514_n 0.00400585f $X=0.575 $Y=0.835 $X2=0
+ $Y2=0
cc_183 N_A_80_313#_c_86_n N_A_286_125#_M1004_d 0.00261503f $X=2.905 $Y=1.12
+ $X2=0 $Y2=0
cc_184 N_A_80_313#_c_86_n N_A_286_125#_c_552_n 0.0051905f $X=2.905 $Y=1.12 $X2=0
+ $Y2=0
cc_185 N_A_80_313#_c_90_n N_A_286_125#_c_552_n 0.0205552f $X=2.02 $Y=0.89 $X2=0
+ $Y2=0
cc_186 N_A_80_313#_c_86_n N_A_286_125#_c_554_n 0.0209703f $X=2.905 $Y=1.12 $X2=0
+ $Y2=0
cc_187 N_A1_c_209_n N_B1_M1003_g 0.00843215f $X=1.515 $Y=1.305 $X2=0 $Y2=0
cc_188 N_A1_c_210_n N_B1_M1003_g 0.00410117f $X=1.6 $Y=2.095 $X2=0 $Y2=0
cc_189 N_A1_c_211_n N_B1_M1003_g 0.0116175f $X=1.355 $Y=0.35 $X2=0 $Y2=0
cc_190 N_A1_c_213_n N_B1_M1003_g 8.28336e-19 $X=1.205 $Y=1.17 $X2=0 $Y2=0
cc_191 A1 N_B1_M1003_g 6.29036e-19 $X=1.2 $Y=0.555 $X2=0 $Y2=0
cc_192 N_A1_c_216_n N_B1_M1007_g 0.00324573f $X=3.06 $Y=2.18 $X2=0 $Y2=0
cc_193 N_A1_c_208_n N_B1_c_294_n 0.00417092f $X=1.355 $Y=0.515 $X2=0 $Y2=0
cc_194 N_A1_c_209_n N_B1_c_294_n 0.00571564f $X=1.515 $Y=1.305 $X2=0 $Y2=0
cc_195 N_A1_c_210_n N_B1_c_294_n 0.0257771f $X=1.6 $Y=2.095 $X2=0 $Y2=0
cc_196 N_A1_c_216_n N_B1_c_294_n 0.00160009f $X=3.06 $Y=2.18 $X2=0 $Y2=0
cc_197 N_A1_c_217_n N_B1_c_294_n 0.00673815f $X=1.685 $Y=2.18 $X2=0 $Y2=0
cc_198 N_A1_c_213_n N_B1_c_294_n 0.00457181f $X=1.205 $Y=1.17 $X2=0 $Y2=0
cc_199 N_A1_c_216_n N_B1_c_295_n 0.0100478f $X=3.06 $Y=2.18 $X2=0 $Y2=0
cc_200 N_A1_c_209_n B1 0.00388928f $X=1.515 $Y=1.305 $X2=0 $Y2=0
cc_201 N_A1_c_210_n B1 0.0374251f $X=1.6 $Y=2.095 $X2=0 $Y2=0
cc_202 N_A1_c_217_n B1 0.011072f $X=1.685 $Y=2.18 $X2=0 $Y2=0
cc_203 N_A1_c_213_n B1 0.0208619f $X=1.205 $Y=1.17 $X2=0 $Y2=0
cc_204 N_A1_c_216_n N_B2_M1001_g 0.0105167f $X=3.06 $Y=2.18 $X2=0 $Y2=0
cc_205 N_A1_c_210_n N_B2_c_342_n 2.88301e-19 $X=1.6 $Y=2.095 $X2=0 $Y2=0
cc_206 N_A1_c_210_n N_B2_c_347_n 7.92145e-19 $X=1.6 $Y=2.095 $X2=0 $Y2=0
cc_207 N_A1_c_216_n N_B2_c_347_n 0.00497948f $X=3.06 $Y=2.18 $X2=0 $Y2=0
cc_208 N_A1_c_209_n B2 6.09167e-19 $X=1.515 $Y=1.305 $X2=0 $Y2=0
cc_209 N_A1_c_210_n B2 0.0308767f $X=1.6 $Y=2.095 $X2=0 $Y2=0
cc_210 N_A1_c_216_n B2 0.0618018f $X=3.06 $Y=2.18 $X2=0 $Y2=0
cc_211 N_A1_M1005_g N_A2_c_392_n 0.0280146f $X=3.135 $Y=2.765 $X2=-0.19
+ $Y2=-0.245
cc_212 N_A1_c_216_n N_A2_c_388_n 0.00817868f $X=3.06 $Y=2.18 $X2=0 $Y2=0
cc_213 N_A1_c_218_n N_A2_c_388_n 0.00115257f $X=3.225 $Y=2.1 $X2=0 $Y2=0
cc_214 N_A1_c_219_n N_A2_c_388_n 0.011263f $X=3.225 $Y=2.1 $X2=0 $Y2=0
cc_215 N_A1_M1005_g N_A2_c_394_n 0.011263f $X=3.135 $Y=2.765 $X2=0 $Y2=0
cc_216 N_A1_c_216_n N_A2_c_394_n 0.00916887f $X=3.06 $Y=2.18 $X2=0 $Y2=0
cc_217 N_A1_c_216_n N_A2_c_391_n 0.00260674f $X=3.06 $Y=2.18 $X2=0 $Y2=0
cc_218 N_A1_c_219_n N_A2_c_391_n 0.00704939f $X=3.225 $Y=2.1 $X2=0 $Y2=0
cc_219 N_A1_c_213_n X 0.00731895f $X=1.205 $Y=1.17 $X2=0 $Y2=0
cc_220 N_A1_M1005_g N_VPWR_c_458_n 0.0122424f $X=3.135 $Y=2.765 $X2=0 $Y2=0
cc_221 N_A1_M1005_g N_VPWR_c_461_n 0.00356919f $X=3.135 $Y=2.765 $X2=0 $Y2=0
cc_222 N_A1_M1005_g N_VPWR_c_457_n 0.00457455f $X=3.135 $Y=2.765 $X2=0 $Y2=0
cc_223 A1 N_VGND_M1000_d 0.00428949f $X=1.2 $Y=0.555 $X2=-0.19 $Y2=-0.245
cc_224 N_A1_c_208_n N_VGND_c_509_n 5.35461e-19 $X=1.355 $Y=0.515 $X2=0 $Y2=0
cc_225 N_A1_c_211_n N_VGND_c_509_n 0.00434898f $X=1.355 $Y=0.35 $X2=0 $Y2=0
cc_226 N_A1_c_212_n N_VGND_c_509_n 0.0177911f $X=1.205 $Y=0.5 $X2=0 $Y2=0
cc_227 A1 N_VGND_c_509_n 0.0061579f $X=1.2 $Y=0.555 $X2=0 $Y2=0
cc_228 N_A1_c_208_n N_VGND_c_519_n 9.6204e-19 $X=1.355 $Y=0.515 $X2=0 $Y2=0
cc_229 A1 N_VGND_c_519_n 0.025106f $X=1.2 $Y=0.555 $X2=0 $Y2=0
cc_230 N_A1_c_211_n N_VGND_c_511_n 0.00989123f $X=1.355 $Y=0.35 $X2=0 $Y2=0
cc_231 N_A1_c_212_n N_VGND_c_511_n 0.0203878f $X=1.205 $Y=0.5 $X2=0 $Y2=0
cc_232 N_A1_c_211_n N_VGND_c_513_n 0.0165388f $X=1.355 $Y=0.35 $X2=0 $Y2=0
cc_233 N_A1_c_212_n N_VGND_c_513_n 0.0110914f $X=1.205 $Y=0.5 $X2=0 $Y2=0
cc_234 N_A1_c_209_n N_A_286_125#_c_559_n 0.014329f $X=1.515 $Y=1.305 $X2=0 $Y2=0
cc_235 N_A1_c_211_n N_A_286_125#_c_553_n 0.0024678f $X=1.355 $Y=0.35 $X2=0 $Y2=0
cc_236 N_A1_c_212_n N_A_286_125#_c_553_n 0.00409552f $X=1.205 $Y=0.5 $X2=0 $Y2=0
cc_237 A1 N_A_286_125#_c_553_n 0.0126446f $X=1.2 $Y=0.555 $X2=0 $Y2=0
cc_238 N_B1_M1003_g N_B2_M1004_g 0.0189399f $X=1.785 $Y=0.835 $X2=0 $Y2=0
cc_239 N_B1_c_295_n N_B2_c_342_n 0.0347805f $X=1.785 $Y=1.9 $X2=0 $Y2=0
cc_240 N_B1_M1007_g N_B2_c_347_n 0.0347805f $X=1.785 $Y=2.765 $X2=0 $Y2=0
cc_241 N_B1_M1003_g B2 0.00524471f $X=1.785 $Y=0.835 $X2=0 $Y2=0
cc_242 N_B1_M1003_g N_B2_c_344_n 0.0347805f $X=1.785 $Y=0.835 $X2=0 $Y2=0
cc_243 N_B1_M1007_g N_VPWR_c_461_n 0.00356919f $X=1.785 $Y=2.765 $X2=0 $Y2=0
cc_244 N_B1_M1007_g N_VPWR_c_457_n 0.00423442f $X=1.785 $Y=2.765 $X2=0 $Y2=0
cc_245 N_B1_M1007_g N_VPWR_c_466_n 0.0118918f $X=1.785 $Y=2.765 $X2=0 $Y2=0
cc_246 N_B1_M1003_g N_VGND_c_511_n 6.71716e-19 $X=1.785 $Y=0.835 $X2=0 $Y2=0
cc_247 N_B1_c_294_n N_A_286_125#_c_559_n 6.40452e-19 $X=1.71 $Y=1.9 $X2=0 $Y2=0
cc_248 N_B1_M1003_g N_A_286_125#_c_552_n 0.0129148f $X=1.785 $Y=0.835 $X2=0
+ $Y2=0
cc_249 N_B1_M1003_g N_A_286_125#_c_553_n 3.06931e-19 $X=1.785 $Y=0.835 $X2=0
+ $Y2=0
cc_250 N_B2_M1004_g N_A2_c_387_n 0.0213154f $X=2.235 $Y=0.835 $X2=0 $Y2=0
cc_251 N_B2_M1001_g N_A2_c_388_n 0.00651061f $X=2.175 $Y=2.765 $X2=0 $Y2=0
cc_252 N_B2_c_342_n N_A2_c_388_n 0.0188943f $X=2.265 $Y=1.81 $X2=0 $Y2=0
cc_253 B2 N_A2_c_388_n 0.0175286f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_254 N_B2_M1001_g N_A2_c_394_n 0.0194113f $X=2.175 $Y=2.765 $X2=0 $Y2=0
cc_255 B2 N_A2_c_394_n 8.49539e-19 $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_256 B2 N_A2_c_389_n 0.00403743f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_257 N_B2_c_344_n N_A2_c_389_n 0.0188943f $X=2.265 $Y=1.47 $X2=0 $Y2=0
cc_258 N_B2_M1001_g N_VPWR_c_461_n 0.0041769f $X=2.175 $Y=2.765 $X2=0 $Y2=0
cc_259 N_B2_M1001_g N_VPWR_c_457_n 0.00593058f $X=2.175 $Y=2.765 $X2=0 $Y2=0
cc_260 N_B2_M1001_g N_VPWR_c_466_n 0.00201585f $X=2.175 $Y=2.765 $X2=0 $Y2=0
cc_261 N_B2_M1004_g N_VGND_c_511_n 6.71716e-19 $X=2.235 $Y=0.835 $X2=0 $Y2=0
cc_262 N_B2_M1004_g N_A_286_125#_c_552_n 0.00930904f $X=2.235 $Y=0.835 $X2=0
+ $Y2=0
cc_263 N_B2_M1004_g N_A_286_125#_c_554_n 0.00183496f $X=2.235 $Y=0.835 $X2=0
+ $Y2=0
cc_264 N_A2_c_392_n N_VPWR_c_458_n 0.00185361f $X=2.605 $Y=2.335 $X2=0 $Y2=0
cc_265 N_A2_c_392_n N_VPWR_c_461_n 0.0041769f $X=2.605 $Y=2.335 $X2=0 $Y2=0
cc_266 N_A2_c_392_n N_VPWR_c_457_n 0.00625343f $X=2.605 $Y=2.335 $X2=0 $Y2=0
cc_267 N_A2_c_387_n N_VGND_c_510_n 0.00752728f $X=2.745 $Y=1.155 $X2=0 $Y2=0
cc_268 N_A2_c_391_n N_VGND_c_510_n 0.00622557f $X=3.42 $Y=1.32 $X2=0 $Y2=0
cc_269 N_A2_c_387_n N_VGND_c_511_n 0.00359608f $X=2.745 $Y=1.155 $X2=0 $Y2=0
cc_270 N_A2_c_387_n N_VGND_c_513_n 0.00394323f $X=2.745 $Y=1.155 $X2=0 $Y2=0
cc_271 N_A2_c_387_n N_A_286_125#_c_554_n 0.00631099f $X=2.745 $Y=1.155 $X2=0
+ $Y2=0
cc_272 X N_VPWR_c_460_n 0.0217542f $X=0.155 $Y=2.69 $X2=0 $Y2=0
cc_273 N_X_M1006_s N_VPWR_c_457_n 0.00212301f $X=0.135 $Y=2.445 $X2=0 $Y2=0
cc_274 X N_VPWR_c_457_n 0.0129532f $X=0.155 $Y=2.69 $X2=0 $Y2=0
cc_275 N_X_c_434_n N_VGND_c_509_n 0.00283769f $X=0.36 $Y=0.77 $X2=0 $Y2=0
cc_276 X N_VGND_c_519_n 0.0029717f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_277 N_X_c_434_n N_VGND_c_513_n 0.0114096f $X=0.36 $Y=0.77 $X2=0 $Y2=0
cc_278 N_X_c_434_n N_VGND_c_514_n 0.00775077f $X=0.36 $Y=0.77 $X2=0 $Y2=0
cc_279 N_VPWR_c_457_n A_372_489# 0.0031085f $X=3.6 $Y=3.33 $X2=-0.19 $Y2=-0.245
cc_280 N_VPWR_c_457_n A_536_489# 0.0049218f $X=3.6 $Y=3.33 $X2=-0.19 $Y2=-0.245
cc_281 N_VGND_c_511_n N_A_286_125#_c_552_n 0.0198324f $X=2.875 $Y=0 $X2=0 $Y2=0
cc_282 N_VGND_c_513_n N_A_286_125#_c_552_n 0.0224567f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_283 N_VGND_c_511_n N_A_286_125#_c_553_n 0.00664058f $X=2.875 $Y=0 $X2=0 $Y2=0
cc_284 N_VGND_c_513_n N_A_286_125#_c_553_n 0.00745183f $X=3.6 $Y=0 $X2=0 $Y2=0
cc_285 N_VGND_c_510_n N_A_286_125#_c_554_n 0.0224151f $X=3.04 $Y=0.77 $X2=0
+ $Y2=0
cc_286 N_VGND_c_511_n N_A_286_125#_c_554_n 0.0102106f $X=2.875 $Y=0 $X2=0 $Y2=0
cc_287 N_VGND_c_513_n N_A_286_125#_c_554_n 0.0111892f $X=3.6 $Y=0 $X2=0 $Y2=0
