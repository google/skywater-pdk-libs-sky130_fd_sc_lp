* File: sky130_fd_sc_lp__o2111a_2.pex.spice
* Created: Fri Aug 28 11:00:03 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O2111A_2%A_80_21# 1 2 3 10 12 13 15 16 18 19 21 23
+ 24 25 28 32 34 36 38 42 43 46
c80 43 0 1.11874e-19 $X=1.175 $Y=1.225
r81 49 51 42.6042 $w=5.4e-07 $l=4.3e-07 $layer=POLY_cond $X=0.475 $Y=1.455
+ $X2=0.905 $Y2=1.455
r82 42 51 15.3573 $w=5.4e-07 $l=1.55e-07 $layer=POLY_cond $X=1.06 $Y=1.455
+ $X2=0.905 $Y2=1.455
r83 41 43 4.99288 $w=2.81e-07 $l=1.15e-07 $layer=LI1_cond $X=1.06 $Y=1.225
+ $X2=1.175 $Y2=1.225
r84 41 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.06
+ $Y=1.35 $X2=1.06 $Y2=1.35
r85 36 48 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.03 $Y=2.125 $X2=3.03
+ $Y2=2.04
r86 36 38 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=3.03 $Y=2.125
+ $X2=3.03 $Y2=2.495
r87 35 46 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.155 $Y=2.04
+ $X2=2.03 $Y2=2.04
r88 34 48 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.865 $Y=2.04
+ $X2=3.03 $Y2=2.04
r89 34 35 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=2.865 $Y=2.04
+ $X2=2.155 $Y2=2.04
r90 30 46 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.03 $Y=2.125
+ $X2=2.03 $Y2=2.04
r91 30 32 15.6732 $w=2.48e-07 $l=3.4e-07 $layer=LI1_cond $X=2.03 $Y=2.125
+ $X2=2.03 $Y2=2.465
r92 26 43 19.7544 $w=2.81e-07 $l=5.47996e-07 $layer=LI1_cond $X=1.63 $Y=1.02
+ $X2=1.175 $Y2=1.225
r93 26 28 19.7562 $w=3.48e-07 $l=6e-07 $layer=LI1_cond $X=1.63 $Y=1.02 $X2=1.63
+ $Y2=0.42
r94 24 46 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.905 $Y=2.04
+ $X2=2.03 $Y2=2.04
r95 24 25 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=1.905 $Y=2.04
+ $X2=1.305 $Y2=2.04
r96 23 25 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=1.175 $Y=1.955
+ $X2=1.305 $Y2=2.04
r97 22 43 1.18573 $w=2.6e-07 $l=2.9e-07 $layer=LI1_cond $X=1.175 $Y=1.515
+ $X2=1.175 $Y2=1.225
r98 22 23 19.5029 $w=2.58e-07 $l=4.4e-07 $layer=LI1_cond $X=1.175 $Y=1.515
+ $X2=1.175 $Y2=1.955
r99 19 51 33.3633 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=0.905 $Y=1.725
+ $X2=0.905 $Y2=1.455
r100 19 21 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=0.905 $Y=1.725
+ $X2=0.905 $Y2=2.465
r101 16 51 33.3633 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=0.905 $Y=1.185
+ $X2=0.905 $Y2=1.455
r102 16 18 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.905 $Y=1.185
+ $X2=0.905 $Y2=0.655
r103 13 49 33.3633 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=0.475 $Y=1.725
+ $X2=0.475 $Y2=1.455
r104 13 15 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=0.475 $Y=1.725
+ $X2=0.475 $Y2=2.465
r105 10 49 33.3633 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=0.475 $Y=1.185
+ $X2=0.475 $Y2=1.455
r106 10 12 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.475 $Y=1.185
+ $X2=0.475 $Y2=0.655
r107 3 48 600 $w=1.7e-07 $l=2.88141e-07 $layer=licon1_PDIFF $count=1 $X=2.83
+ $Y=1.835 $X2=3.03 $Y2=2.04
r108 3 38 300 $w=1.7e-07 $l=7.53392e-07 $layer=licon1_PDIFF $count=2 $X=2.83
+ $Y=1.835 $X2=3.03 $Y2=2.495
r109 2 46 600 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=1 $X=1.86
+ $Y=1.835 $X2=2 $Y2=2.04
r110 2 32 300 $w=1.7e-07 $l=6.96491e-07 $layer=licon1_PDIFF $count=2 $X=1.86
+ $Y=1.835 $X2=2 $Y2=2.465
r111 1 28 91 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=2 $X=1.515
+ $Y=0.255 $X2=1.64 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__O2111A_2%D1 3 7 9 13 16
r34 15 16 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=1.785 $Y=1.51
+ $X2=1.855 $Y2=1.51
r35 12 15 25.3549 $w=3.3e-07 $l=1.45e-07 $layer=POLY_cond $X=1.64 $Y=1.51
+ $X2=1.785 $Y2=1.51
r36 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.64
+ $Y=1.51 $X2=1.64 $Y2=1.51
r37 9 13 4.89394 $w=3.63e-07 $l=1.55e-07 $layer=LI1_cond $X=1.657 $Y=1.665
+ $X2=1.657 $Y2=1.51
r38 5 16 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.855 $Y=1.345
+ $X2=1.855 $Y2=1.51
r39 5 7 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=1.855 $Y=1.345
+ $X2=1.855 $Y2=0.675
r40 1 15 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.785 $Y=1.675
+ $X2=1.785 $Y2=1.51
r41 1 3 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.785 $Y=1.675
+ $X2=1.785 $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__O2111A_2%C1 3 6 8 9 10 11 18 20 30
c43 20 0 1.11874e-19 $X=2.305 $Y=1.205
r44 22 30 1.51637 $w=3.78e-07 $l=5e-08 $layer=LI1_cond $X=2.2 $Y=1.345 $X2=2.2
+ $Y2=1.295
r45 18 21 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.305 $Y=1.37
+ $X2=2.305 $Y2=1.535
r46 18 20 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.305 $Y=1.37
+ $X2=2.305 $Y2=1.205
r47 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.305
+ $Y=1.37 $X2=2.305 $Y2=1.37
r48 11 19 10.5853 $w=3.4e-07 $l=2.95e-07 $layer=LI1_cond $X=2.2 $Y=1.665 $X2=2.2
+ $Y2=1.37
r49 10 19 0.287059 $w=3.4e-07 $l=8e-09 $layer=LI1_cond $X=2.2 $Y=1.362 $X2=2.2
+ $Y2=1.37
r50 10 22 0.7088 $w=3.8e-07 $l=1.7e-08 $layer=LI1_cond $X=2.2 $Y=1.362 $X2=2.2
+ $Y2=1.345
r51 10 30 0.545894 $w=3.78e-07 $l=1.8e-08 $layer=LI1_cond $X=2.2 $Y=1.277
+ $X2=2.2 $Y2=1.295
r52 9 10 10.6753 $w=3.78e-07 $l=3.52e-07 $layer=LI1_cond $X=2.2 $Y=0.925 $X2=2.2
+ $Y2=1.277
r53 8 9 11.2212 $w=3.78e-07 $l=3.7e-07 $layer=LI1_cond $X=2.2 $Y=0.555 $X2=2.2
+ $Y2=0.925
r54 6 21 476.872 $w=1.5e-07 $l=9.3e-07 $layer=POLY_cond $X=2.215 $Y=2.465
+ $X2=2.215 $Y2=1.535
r55 3 20 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.215 $Y=0.675
+ $X2=2.215 $Y2=1.205
.ends

.subckt PM_SKY130_FD_SC_LP__O2111A_2%B1 3 7 9 12
r34 12 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.845 $Y=1.51
+ $X2=2.845 $Y2=1.675
r35 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.845 $Y=1.51
+ $X2=2.845 $Y2=1.345
r36 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.845
+ $Y=1.51 $X2=2.845 $Y2=1.51
r37 9 13 7.88959 $w=3.17e-07 $l=2.05e-07 $layer=LI1_cond $X=2.64 $Y=1.605
+ $X2=2.845 $Y2=1.605
r38 7 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.755 $Y=2.465
+ $X2=2.755 $Y2=1.675
r39 3 14 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=2.755 $Y=0.675
+ $X2=2.755 $Y2=1.345
.ends

.subckt PM_SKY130_FD_SC_LP__O2111A_2%A2 3 7 9 10 11 12 19
r33 23 34 0.0129374 $w=2.8e-07 $l=1.25e-07 $layer=LI1_cond $X=3.575 $Y=1.675
+ $X2=3.575 $Y2=1.55
r34 20 34 8.75857 $w=2.48e-07 $l=1.9e-07 $layer=LI1_cond $X=3.385 $Y=1.55
+ $X2=3.575 $Y2=1.55
r35 19 22 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.385 $Y=1.51
+ $X2=3.385 $Y2=1.675
r36 19 21 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.385 $Y=1.51
+ $X2=3.385 $Y2=1.345
r37 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.385
+ $Y=1.51 $X2=3.385 $Y2=1.51
r38 11 12 15.2287 $w=2.78e-07 $l=3.7e-07 $layer=LI1_cond $X=3.575 $Y=2.405
+ $X2=3.575 $Y2=2.775
r39 10 11 15.2287 $w=2.78e-07 $l=3.7e-07 $layer=LI1_cond $X=3.575 $Y=2.035
+ $X2=3.575 $Y2=2.405
r40 9 34 1.15244 $w=2.48e-07 $l=2.5e-08 $layer=LI1_cond $X=3.6 $Y=1.55 $X2=3.575
+ $Y2=1.55
r41 9 10 13.2943 $w=2.78e-07 $l=3.23e-07 $layer=LI1_cond $X=3.575 $Y=1.712
+ $X2=3.575 $Y2=2.035
r42 9 23 1.52287 $w=2.78e-07 $l=3.7e-08 $layer=LI1_cond $X=3.575 $Y=1.712
+ $X2=3.575 $Y2=1.675
r43 7 22 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.295 $Y=2.465
+ $X2=3.295 $Y2=1.675
r44 3 21 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=3.295 $Y=0.675
+ $X2=3.295 $Y2=1.345
.ends

.subckt PM_SKY130_FD_SC_LP__O2111A_2%A1 3 7 9 14 15
r25 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.05
+ $Y=1.46 $X2=4.05 $Y2=1.46
r26 11 14 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=3.835 $Y=1.46
+ $X2=4.05 $Y2=1.46
r27 9 15 6.75002 $w=3.48e-07 $l=2.05e-07 $layer=LI1_cond $X=4.06 $Y=1.665
+ $X2=4.06 $Y2=1.46
r28 5 11 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.835 $Y=1.625
+ $X2=3.835 $Y2=1.46
r29 5 7 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=3.835 $Y=1.625
+ $X2=3.835 $Y2=2.465
r30 1 11 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.835 $Y=1.295
+ $X2=3.835 $Y2=1.46
r31 1 3 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=3.835 $Y=1.295
+ $X2=3.835 $Y2=0.675
.ends

.subckt PM_SKY130_FD_SC_LP__O2111A_2%VPWR 1 2 3 4 13 15 21 25 27 29 33 35 40 45
+ 54 57 61 68
r59 60 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r60 58 68 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.4 $Y2=3.33
r61 57 58 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r62 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r63 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r64 49 61 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r65 49 58 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=2.64 $Y2=3.33
r66 48 49 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r67 46 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.655 $Y=3.33
+ $X2=2.49 $Y2=3.33
r68 46 48 61.6524 $w=1.68e-07 $l=9.45e-07 $layer=LI1_cond $X=2.655 $Y=3.33
+ $X2=3.6 $Y2=3.33
r69 45 60 4.76062 $w=1.7e-07 $l=2.17e-07 $layer=LI1_cond $X=3.885 $Y=3.33
+ $X2=4.102 $Y2=3.33
r70 45 48 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=3.885 $Y=3.33
+ $X2=3.6 $Y2=3.33
r71 41 54 14.259 $w=1.7e-07 $l=3.8e-07 $layer=LI1_cond $X=1.735 $Y=3.33
+ $X2=1.355 $Y2=3.33
r72 41 43 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=1.735 $Y=3.33
+ $X2=2.16 $Y2=3.33
r73 40 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.325 $Y=3.33
+ $X2=2.49 $Y2=3.33
r74 40 43 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=2.325 $Y=3.33
+ $X2=2.16 $Y2=3.33
r75 39 55 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r76 39 52 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r77 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r78 36 51 4.45907 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=0.39 $Y=3.33
+ $X2=0.195 $Y2=3.33
r79 36 38 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=0.39 $Y=3.33
+ $X2=0.72 $Y2=3.33
r80 35 54 14.259 $w=1.7e-07 $l=3.8e-07 $layer=LI1_cond $X=0.975 $Y=3.33
+ $X2=1.355 $Y2=3.33
r81 35 38 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.975 $Y=3.33
+ $X2=0.72 $Y2=3.33
r82 33 68 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.4 $Y2=3.33
r83 33 55 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.2 $Y2=3.33
r84 33 43 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r85 29 32 33.0018 $w=3.28e-07 $l=9.45e-07 $layer=LI1_cond $X=4.05 $Y=2.005
+ $X2=4.05 $Y2=2.95
r86 27 60 3.00555 $w=3.3e-07 $l=1.07912e-07 $layer=LI1_cond $X=4.05 $Y=3.245
+ $X2=4.102 $Y2=3.33
r87 27 32 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=4.05 $Y=3.245
+ $X2=4.05 $Y2=2.95
r88 23 57 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.49 $Y=3.245
+ $X2=2.49 $Y2=3.33
r89 23 25 29.5095 $w=3.28e-07 $l=8.45e-07 $layer=LI1_cond $X=2.49 $Y=3.245
+ $X2=2.49 $Y2=2.4
r90 19 54 3.03114 $w=7.6e-07 $l=8.5e-08 $layer=LI1_cond $X=1.355 $Y=3.245
+ $X2=1.355 $Y2=3.33
r91 19 21 13.6133 $w=7.58e-07 $l=8.65e-07 $layer=LI1_cond $X=1.355 $Y=3.245
+ $X2=1.355 $Y2=2.38
r92 15 18 37.6986 $w=2.93e-07 $l=9.65e-07 $layer=LI1_cond $X=0.242 $Y=1.985
+ $X2=0.242 $Y2=2.95
r93 13 51 3.01845 $w=2.95e-07 $l=1.05924e-07 $layer=LI1_cond $X=0.242 $Y=3.245
+ $X2=0.195 $Y2=3.33
r94 13 18 11.5244 $w=2.93e-07 $l=2.95e-07 $layer=LI1_cond $X=0.242 $Y=3.245
+ $X2=0.242 $Y2=2.95
r95 4 32 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=3.91
+ $Y=1.835 $X2=4.05 $Y2=2.95
r96 4 29 400 $w=1.7e-07 $l=2.29565e-07 $layer=licon1_PDIFF $count=1 $X=3.91
+ $Y=1.835 $X2=4.05 $Y2=2.005
r97 3 25 300 $w=1.7e-07 $l=6.57438e-07 $layer=licon1_PDIFF $count=2 $X=2.29
+ $Y=1.835 $X2=2.49 $Y2=2.4
r98 2 21 150 $w=1.7e-07 $l=8.18321e-07 $layer=licon1_PDIFF $count=4 $X=0.98
+ $Y=1.835 $X2=1.57 $Y2=2.38
r99 1 18 400 $w=1.7e-07 $l=1.17584e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.835 $X2=0.26 $Y2=2.95
r100 1 15 400 $w=1.7e-07 $l=2.03101e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.835 $X2=0.26 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_LP__O2111A_2%X 1 2 7 8 9 10 11 12 13 22
r17 13 40 6.3502 $w=2.43e-07 $l=1.35e-07 $layer=LI1_cond $X=0.682 $Y=2.775
+ $X2=0.682 $Y2=2.91
r18 12 13 17.4042 $w=2.43e-07 $l=3.7e-07 $layer=LI1_cond $X=0.682 $Y=2.405
+ $X2=0.682 $Y2=2.775
r19 11 12 19.9914 $w=2.43e-07 $l=4.25e-07 $layer=LI1_cond $X=0.682 $Y=1.98
+ $X2=0.682 $Y2=2.405
r20 10 11 14.8171 $w=2.43e-07 $l=3.15e-07 $layer=LI1_cond $X=0.682 $Y=1.665
+ $X2=0.682 $Y2=1.98
r21 9 10 17.4042 $w=2.43e-07 $l=3.7e-07 $layer=LI1_cond $X=0.682 $Y=1.295
+ $X2=0.682 $Y2=1.665
r22 8 9 17.4042 $w=2.43e-07 $l=3.7e-07 $layer=LI1_cond $X=0.682 $Y=0.925
+ $X2=0.682 $Y2=1.295
r23 7 8 17.4042 $w=2.43e-07 $l=3.7e-07 $layer=LI1_cond $X=0.682 $Y=0.555
+ $X2=0.682 $Y2=0.925
r24 7 22 6.3502 $w=2.43e-07 $l=1.35e-07 $layer=LI1_cond $X=0.682 $Y=0.555
+ $X2=0.682 $Y2=0.42
r25 2 40 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=1.835 $X2=0.69 $Y2=2.91
r26 2 11 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=1.835 $X2=0.69 $Y2=1.98
r27 1 22 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=0.55
+ $Y=0.235 $X2=0.69 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__O2111A_2%VGND 1 2 3 10 12 16 20 22 24 29 39 40 46 49
+ 58
r48 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r49 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r50 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r51 40 50 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.6
+ $Y2=0
r52 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r53 37 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.715 $Y=0 $X2=3.55
+ $Y2=0
r54 37 39 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=3.715 $Y=0 $X2=4.08
+ $Y2=0
r55 36 50 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r56 36 58 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.4
+ $Y2=0
r57 35 36 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r58 33 47 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r59 32 35 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.68 $Y=0 $X2=3.12
+ $Y2=0
r60 32 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r61 30 46 8.23795 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=1.285 $Y=0 $X2=1.13
+ $Y2=0
r62 30 32 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=1.285 $Y=0 $X2=1.68
+ $Y2=0
r63 29 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.385 $Y=0 $X2=3.55
+ $Y2=0
r64 29 35 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=3.385 $Y=0 $X2=3.12
+ $Y2=0
r65 28 47 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r66 28 44 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r67 27 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r68 25 43 4.45907 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=0.39 $Y=0 $X2=0.195
+ $Y2=0
r69 25 27 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=0.39 $Y=0 $X2=0.72
+ $Y2=0
r70 24 46 8.23795 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=0.975 $Y=0 $X2=1.13
+ $Y2=0
r71 24 27 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.975 $Y=0 $X2=0.72
+ $Y2=0
r72 22 58 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.4
+ $Y2=0
r73 22 33 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.68
+ $Y2=0
r74 18 49 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.55 $Y=0.085
+ $X2=3.55 $Y2=0
r75 18 20 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=3.55 $Y=0.085
+ $X2=3.55 $Y2=0.4
r76 14 46 0.701276 $w=3.1e-07 $l=8.5e-08 $layer=LI1_cond $X=1.13 $Y=0.085
+ $X2=1.13 $Y2=0
r77 14 16 10.9668 $w=3.08e-07 $l=2.95e-07 $layer=LI1_cond $X=1.13 $Y=0.085
+ $X2=1.13 $Y2=0.38
r78 10 43 3.01845 $w=2.95e-07 $l=1.05924e-07 $layer=LI1_cond $X=0.242 $Y=0.085
+ $X2=0.195 $Y2=0
r79 10 12 11.5244 $w=2.93e-07 $l=2.95e-07 $layer=LI1_cond $X=0.242 $Y=0.085
+ $X2=0.242 $Y2=0.38
r80 3 20 91 $w=1.7e-07 $l=2.41868e-07 $layer=licon1_NDIFF $count=2 $X=3.37
+ $Y=0.255 $X2=3.55 $Y2=0.4
r81 2 16 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=0.98
+ $Y=0.235 $X2=1.12 $Y2=0.38
r82 1 12 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_LP__O2111A_2%A_566_51# 1 2 9 11 12 15
r22 13 15 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=4.05 $Y=1.035
+ $X2=4.05 $Y2=0.4
r23 11 13 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.885 $Y=1.12
+ $X2=4.05 $Y2=1.035
r24 11 12 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.885 $Y=1.12
+ $X2=3.195 $Y2=1.12
r25 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.03 $Y=1.035
+ $X2=3.195 $Y2=1.12
r26 7 9 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=3.03 $Y=1.035
+ $X2=3.03 $Y2=0.4
r27 2 15 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.91
+ $Y=0.255 $X2=4.05 $Y2=0.4
r28 1 9 91 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_NDIFF $count=2 $X=2.83
+ $Y=0.255 $X2=3.03 $Y2=0.4
.ends

