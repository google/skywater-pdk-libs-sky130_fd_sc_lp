* File: sky130_fd_sc_lp__dfstp_lp.pex.spice
* Created: Fri Aug 28 10:23:33 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__DFSTP_LP%D 1 3 8 10 12 16 18 19 23 24 25
c35 10 0 1.1902e-19 $X=0.835 $Y=0.78
r36 23 26 72.9334 $w=4.55e-07 $l=5.05e-07 $layer=POLY_cond $X=0.447 $Y=1.275
+ $X2=0.447 $Y2=1.78
r37 23 25 28.8071 $w=4.55e-07 $l=1.65e-07 $layer=POLY_cond $X=0.447 $Y=1.275
+ $X2=0.447 $Y2=1.11
r38 23 24 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.385
+ $Y=1.275 $X2=0.385 $Y2=1.275
r39 18 19 10.033 $w=4.23e-07 $l=3.7e-07 $layer=LI1_cond $X=0.337 $Y=1.295
+ $X2=0.337 $Y2=1.665
r40 18 24 0.542326 $w=4.23e-07 $l=2e-08 $layer=LI1_cond $X=0.337 $Y=1.295
+ $X2=0.337 $Y2=1.275
r41 10 16 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.835 $Y=0.78
+ $X2=0.835 $Y2=0.855
r42 10 12 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.835 $Y=0.78
+ $X2=0.835 $Y2=0.495
r43 8 26 190.067 $w=2.5e-07 $l=7.65e-07 $layer=POLY_cond $X=0.55 $Y=2.545
+ $X2=0.55 $Y2=1.78
r44 4 16 152.804 $w=1.5e-07 $l=2.98e-07 $layer=POLY_cond $X=0.537 $Y=0.855
+ $X2=0.835 $Y2=0.855
r45 4 13 31.7915 $w=1.5e-07 $l=6.2e-08 $layer=POLY_cond $X=0.537 $Y=0.855
+ $X2=0.475 $Y2=0.855
r46 4 25 39.2642 $w=2.75e-07 $l=1.8e-07 $layer=POLY_cond $X=0.537 $Y=0.93
+ $X2=0.537 $Y2=1.11
r47 1 13 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.475 $Y=0.78
+ $X2=0.475 $Y2=0.855
r48 1 3 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.475 $Y=0.78 $X2=0.475
+ $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__DFSTP_LP%CLK 3 5 7 10 12 14 15 16 19 21
c57 3 0 4.93603e-20 $X=1.74 $Y=2.545
r58 19 22 31.9397 $w=3.55e-07 $l=1.65e-07 $layer=POLY_cond $X=1.687 $Y=1.615
+ $X2=1.687 $Y2=1.78
r59 19 21 46.504 $w=3.55e-07 $l=1.65e-07 $layer=POLY_cond $X=1.687 $Y=1.615
+ $X2=1.687 $Y2=1.45
r60 16 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.675
+ $Y=1.615 $X2=1.675 $Y2=1.615
r61 12 14 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.15 $Y=1.04 $X2=2.15
+ $Y2=0.755
r62 11 15 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.865 $Y=1.115
+ $X2=1.79 $Y2=1.115
r63 10 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.075 $Y=1.115
+ $X2=2.15 $Y2=1.04
r64 10 11 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=2.075 $Y=1.115
+ $X2=1.865 $Y2=1.115
r65 8 15 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.79 $Y=1.19 $X2=1.79
+ $Y2=1.115
r66 8 21 133.319 $w=1.5e-07 $l=2.6e-07 $layer=POLY_cond $X=1.79 $Y=1.19 $X2=1.79
+ $Y2=1.45
r67 5 15 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.79 $Y=1.04 $X2=1.79
+ $Y2=1.115
r68 5 7 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=1.79 $Y=1.04 $X2=1.79
+ $Y2=0.755
r69 3 22 190.067 $w=2.5e-07 $l=7.65e-07 $layer=POLY_cond $X=1.74 $Y=2.545
+ $X2=1.74 $Y2=1.78
.ends

.subckt PM_SKY130_FD_SC_LP__DFSTP_LP%A_479_409# 1 2 9 11 13 17 21 23 25 27 32 35
+ 38 41 42 43 45 46 47 49 50 51 52 53 56 57 62 65 66 69 71 74
c233 74 0 2.60714e-19 $X=7.615 $Y=1.465
c234 52 0 8.79208e-20 $X=7.615 $Y=1.84
c235 51 0 1.93287e-19 $X=6.505 $Y=2.145
c236 42 0 4.4821e-20 $X=5.45 $Y=2.52
c237 23 0 4.93603e-20 $X=2.495 $Y=2.895
c238 11 0 1.26171e-20 $X=4.445 $Y=1.215
c239 9 0 5.35053e-20 $X=3.42 $Y=2.595
r240 74 80 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.615 $Y=1.465
+ $X2=7.615 $Y2=1.3
r241 73 74 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.615
+ $Y=1.465 $X2=7.615 $Y2=1.465
r242 69 77 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.38 $Y=1.675
+ $X2=3.38 $Y2=1.84
r243 68 70 9.6413 $w=5.18e-07 $l=1.65e-07 $layer=LI1_cond $X=3.41 $Y=1.675
+ $X2=3.41 $Y2=1.84
r244 68 69 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.38
+ $Y=1.675 $X2=3.38 $Y2=1.675
r245 65 68 6.0954 $w=5.18e-07 $l=2.65e-07 $layer=LI1_cond $X=3.41 $Y=1.41
+ $X2=3.41 $Y2=1.675
r246 65 66 9.6413 $w=5.18e-07 $l=1.65e-07 $layer=LI1_cond $X=3.41 $Y=1.41
+ $X2=3.41 $Y2=1.245
r247 64 66 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=3.235 $Y=0.985
+ $X2=3.235 $Y2=1.245
r248 62 64 9.16063 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=3.155 $Y=0.8
+ $X2=3.155 $Y2=0.985
r249 57 84 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.515 $Y=1.675
+ $X2=8.515 $Y2=1.84
r250 56 57 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.515
+ $Y=1.675 $X2=8.515 $Y2=1.675
r251 54 73 3.40825 $w=3.3e-07 $l=2.11069e-07 $layer=LI1_cond $X=7.78 $Y=1.675
+ $X2=7.615 $Y2=1.57
r252 54 56 25.668 $w=3.28e-07 $l=7.35e-07 $layer=LI1_cond $X=7.78 $Y=1.675
+ $X2=8.515 $Y2=1.675
r253 52 73 3.40825 $w=3.3e-07 $l=2.7e-07 $layer=LI1_cond $X=7.615 $Y=1.84
+ $X2=7.615 $Y2=1.57
r254 52 53 7.68295 $w=3.28e-07 $l=2.2e-07 $layer=LI1_cond $X=7.615 $Y=1.84
+ $X2=7.615 $Y2=2.06
r255 50 53 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=7.45 $Y=2.145
+ $X2=7.615 $Y2=2.06
r256 50 51 61.6524 $w=1.68e-07 $l=9.45e-07 $layer=LI1_cond $X=7.45 $Y=2.145
+ $X2=6.505 $Y2=2.145
r257 48 51 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.42 $Y=2.23
+ $X2=6.505 $Y2=2.145
r258 48 49 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=6.42 $Y=2.23
+ $X2=6.42 $Y2=2.895
r259 46 49 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.335 $Y=2.98
+ $X2=6.42 $Y2=2.895
r260 46 47 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=6.335 $Y=2.98
+ $X2=5.62 $Y2=2.98
r261 45 47 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.535 $Y=2.895
+ $X2=5.62 $Y2=2.98
r262 44 45 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=5.535 $Y=2.605
+ $X2=5.535 $Y2=2.895
r263 42 44 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.45 $Y=2.52
+ $X2=5.535 $Y2=2.605
r264 42 43 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=5.45 $Y=2.52
+ $X2=4.76 $Y2=2.52
r265 40 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.675 $Y=2.605
+ $X2=4.76 $Y2=2.52
r266 40 41 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=4.675 $Y=2.605
+ $X2=4.675 $Y2=2.895
r267 39 71 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.67 $Y=2.98
+ $X2=3.585 $Y2=2.98
r268 38 41 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.59 $Y=2.98
+ $X2=4.675 $Y2=2.895
r269 38 39 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=4.59 $Y=2.98
+ $X2=3.67 $Y2=2.98
r270 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.34
+ $Y=1.41 $X2=4.34 $Y2=1.41
r271 33 65 3.39791 $w=3.3e-07 $l=2.6e-07 $layer=LI1_cond $X=3.67 $Y=1.41
+ $X2=3.41 $Y2=1.41
r272 33 35 23.3981 $w=3.28e-07 $l=6.7e-07 $layer=LI1_cond $X=3.67 $Y=1.41
+ $X2=4.34 $Y2=1.41
r273 32 71 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.585 $Y=2.895
+ $X2=3.585 $Y2=2.98
r274 32 70 68.8289 $w=1.68e-07 $l=1.055e-06 $layer=LI1_cond $X=3.585 $Y=2.895
+ $X2=3.585 $Y2=1.84
r275 28 60 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.62 $Y=2.98
+ $X2=2.495 $Y2=2.98
r276 27 71 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.5 $Y=2.98
+ $X2=3.585 $Y2=2.98
r277 27 28 57.4118 $w=1.68e-07 $l=8.8e-07 $layer=LI1_cond $X=3.5 $Y=2.98
+ $X2=2.62 $Y2=2.98
r278 23 60 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.495 $Y=2.895
+ $X2=2.495 $Y2=2.98
r279 23 25 32.4989 $w=2.48e-07 $l=7.05e-07 $layer=LI1_cond $X=2.495 $Y=2.895
+ $X2=2.495 $Y2=2.19
r280 21 84 187.582 $w=2.5e-07 $l=7.55e-07 $layer=POLY_cond $X=8.505 $Y=2.595
+ $X2=8.505 $Y2=1.84
r281 17 80 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=7.555 $Y=0.835
+ $X2=7.555 $Y2=1.3
r282 11 36 42.9482 $w=3.36e-07 $l=2.39029e-07 $layer=POLY_cond $X=4.445 $Y=1.215
+ $X2=4.347 $Y2=1.41
r283 11 13 194.851 $w=1.5e-07 $l=3.8e-07 $layer=POLY_cond $X=4.445 $Y=1.215
+ $X2=4.445 $Y2=0.835
r284 9 77 187.582 $w=2.5e-07 $l=7.55e-07 $layer=POLY_cond $X=3.42 $Y=2.595
+ $X2=3.42 $Y2=1.84
r285 2 60 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=2.395
+ $Y=2.045 $X2=2.535 $Y2=2.9
r286 2 25 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.395
+ $Y=2.045 $X2=2.535 $Y2=2.19
r287 1 62 182 $w=1.7e-07 $l=3.17372e-07 $layer=licon1_NDIFF $count=1 $X=3.015
+ $Y=0.545 $X2=3.155 $Y2=0.8
.ends

.subckt PM_SKY130_FD_SC_LP__DFSTP_LP%A_943_321# 1 2 9 13 18 19 20 21 22 23 25 28
+ 33
c90 25 0 4.40676e-20 $X=5.78 $Y=1.225
c91 23 0 6.02731e-20 $X=5.365 $Y=2.17
c92 20 0 9.1185e-20 $X=5.695 $Y=1.31
c93 13 0 8.28843e-20 $X=4.805 $Y=0.835
r94 35 37 6.12014 $w=3.3e-07 $l=3.5e-08 $layer=POLY_cond $X=4.805 $Y=1.77
+ $X2=4.84 $Y2=1.77
r95 30 33 5.97563 $w=4.03e-07 $l=2.1e-07 $layer=LI1_cond $X=5.78 $Y=0.817
+ $X2=5.99 $Y2=0.817
r96 26 28 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=5.99 $Y=2.255
+ $X2=5.99 $Y2=2.4
r97 24 30 5.85399 $w=1.7e-07 $l=2.03e-07 $layer=LI1_cond $X=5.78 $Y=1.02
+ $X2=5.78 $Y2=0.817
r98 24 25 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=5.78 $Y=1.02
+ $X2=5.78 $Y2=1.225
r99 22 26 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.825 $Y=2.17
+ $X2=5.99 $Y2=2.255
r100 22 23 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=5.825 $Y=2.17
+ $X2=5.365 $Y2=2.17
r101 20 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.695 $Y=1.31
+ $X2=5.78 $Y2=1.225
r102 20 21 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=5.695 $Y=1.31
+ $X2=5.365 $Y2=1.31
r103 19 37 62.9501 $w=3.3e-07 $l=3.6e-07 $layer=POLY_cond $X=5.2 $Y=1.77
+ $X2=4.84 $Y2=1.77
r104 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.2
+ $Y=1.77 $X2=5.2 $Y2=1.77
r105 16 23 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.2 $Y=2.085
+ $X2=5.365 $Y2=2.17
r106 16 18 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=5.2 $Y=2.085
+ $X2=5.2 $Y2=1.77
r107 15 21 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.2 $Y=1.395
+ $X2=5.365 $Y2=1.31
r108 15 18 13.0959 $w=3.28e-07 $l=3.75e-07 $layer=LI1_cond $X=5.2 $Y=1.395
+ $X2=5.2 $Y2=1.77
r109 11 35 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.805 $Y=1.605
+ $X2=4.805 $Y2=1.77
r110 11 13 394.83 $w=1.5e-07 $l=7.7e-07 $layer=POLY_cond $X=4.805 $Y=1.605
+ $X2=4.805 $Y2=0.835
r111 7 37 9.34494 $w=2.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.84 $Y=1.935
+ $X2=4.84 $Y2=1.77
r112 7 9 163.979 $w=2.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.84 $Y=1.935
+ $X2=4.84 $Y2=2.595
r113 2 28 600 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_PDIFF $count=1 $X=5.85
+ $Y=2.095 $X2=5.99 $Y2=2.4
r114 1 33 182 $w=1.7e-07 $l=2.5229e-07 $layer=licon1_NDIFF $count=1 $X=5.845
+ $Y=0.625 $X2=5.99 $Y2=0.815
.ends

.subckt PM_SKY130_FD_SC_LP__DFSTP_LP%A_709_419# 1 2 9 13 14 15 17 20 24 28 29 32
+ 34 35 36 39 40 43 44 45 47 49 50 51 55 59 61 62 68 69 72
c198 69 0 8.79208e-20 $X=7.075 $Y=1.365
c199 68 0 8.70766e-20 $X=7.075 $Y=1.365
c200 55 0 8.28843e-20 $X=4.17 $Y=0.835
c201 35 0 1.26171e-20 $X=4.18 $Y=2.16
c202 20 0 5.61132e-20 $X=7.115 $Y=2.595
c203 9 0 1.93287e-19 $X=5.725 $Y=2.595
r204 68 69 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.075
+ $Y=1.365 $X2=7.075 $Y2=1.365
r205 64 66 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=6.13 $Y=1.285
+ $X2=6.42 $Y2=1.285
r206 62 73 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.74 $Y=1.74
+ $X2=5.74 $Y2=1.905
r207 62 72 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.74 $Y=1.74
+ $X2=5.74 $Y2=1.575
r208 61 63 18.881 $w=2.52e-07 $l=3.9e-07 $layer=LI1_cond $X=5.74 $Y=1.74
+ $X2=6.13 $Y2=1.74
r209 61 62 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.74
+ $Y=1.74 $X2=5.74 $Y2=1.74
r210 55 57 6.22319 $w=2.48e-07 $l=1.35e-07 $layer=LI1_cond $X=4.21 $Y=0.835
+ $X2=4.21 $Y2=0.97
r211 51 66 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=6.505 $Y=1.285
+ $X2=6.42 $Y2=1.285
r212 50 68 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.91 $Y=1.285
+ $X2=7.075 $Y2=1.285
r213 50 51 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=6.91 $Y=1.285
+ $X2=6.505 $Y2=1.285
r214 49 66 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.42 $Y=1.2
+ $X2=6.42 $Y2=1.285
r215 48 49 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=6.42 $Y=0.435
+ $X2=6.42 $Y2=1.2
r216 47 63 3.04159 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.13 $Y=1.575
+ $X2=6.13 $Y2=1.74
r217 46 64 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.13 $Y=1.37
+ $X2=6.13 $Y2=1.285
r218 46 47 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=6.13 $Y=1.37
+ $X2=6.13 $Y2=1.575
r219 44 48 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.335 $Y=0.35
+ $X2=6.42 $Y2=0.435
r220 44 45 53.4973 $w=1.68e-07 $l=8.2e-07 $layer=LI1_cond $X=6.335 $Y=0.35
+ $X2=5.515 $Y2=0.35
r221 42 45 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.43 $Y=0.435
+ $X2=5.515 $Y2=0.35
r222 42 43 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=5.43 $Y=0.435
+ $X2=5.43 $Y2=0.875
r223 41 59 4.92476 $w=1.8e-07 $l=8.9861e-08 $layer=LI1_cond $X=4.855 $Y=0.96
+ $X2=4.77 $Y2=0.97
r224 40 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.345 $Y=0.96
+ $X2=5.43 $Y2=0.875
r225 40 41 31.9679 $w=1.68e-07 $l=4.9e-07 $layer=LI1_cond $X=5.345 $Y=0.96
+ $X2=4.855 $Y2=0.96
r226 38 59 1.54918 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=4.77 $Y=1.065
+ $X2=4.77 $Y2=0.97
r227 38 39 65.8931 $w=1.68e-07 $l=1.01e-06 $layer=LI1_cond $X=4.77 $Y=1.065
+ $X2=4.77 $Y2=2.075
r228 37 57 2.34666 $w=1.9e-07 $l=1.25e-07 $layer=LI1_cond $X=4.335 $Y=0.97
+ $X2=4.21 $Y2=0.97
r229 36 59 4.92476 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=4.685 $Y=0.97
+ $X2=4.77 $Y2=0.97
r230 36 37 20.4306 $w=1.88e-07 $l=3.5e-07 $layer=LI1_cond $X=4.685 $Y=0.97
+ $X2=4.335 $Y2=0.97
r231 34 39 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.685 $Y=2.16
+ $X2=4.77 $Y2=2.075
r232 34 35 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=4.685 $Y=2.16
+ $X2=4.18 $Y2=2.16
r233 30 35 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.015 $Y=2.245
+ $X2=4.18 $Y2=2.16
r234 30 32 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=4.015 $Y=2.245
+ $X2=4.015 $Y2=2.395
r235 28 69 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=7.075 $Y=1.705
+ $X2=7.075 $Y2=1.365
r236 28 29 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.075 $Y=1.705
+ $X2=7.075 $Y2=1.87
r237 27 69 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.075 $Y=1.2
+ $X2=7.075 $Y2=1.365
r238 24 27 187.16 $w=1.5e-07 $l=3.65e-07 $layer=POLY_cond $X=7.165 $Y=0.835
+ $X2=7.165 $Y2=1.2
r239 20 29 180.129 $w=2.5e-07 $l=7.25e-07 $layer=POLY_cond $X=7.115 $Y=2.595
+ $X2=7.115 $Y2=1.87
r240 15 17 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=6.205 $Y=1.12
+ $X2=6.205 $Y2=0.835
r241 13 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.13 $Y=1.195
+ $X2=6.205 $Y2=1.12
r242 13 14 115.372 $w=1.5e-07 $l=2.25e-07 $layer=POLY_cond $X=6.13 $Y=1.195
+ $X2=5.905 $Y2=1.195
r243 11 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.83 $Y=1.27
+ $X2=5.905 $Y2=1.195
r244 11 72 156.394 $w=1.5e-07 $l=3.05e-07 $layer=POLY_cond $X=5.83 $Y=1.27
+ $X2=5.83 $Y2=1.575
r245 9 73 171.433 $w=2.5e-07 $l=6.9e-07 $layer=POLY_cond $X=5.725 $Y=2.595
+ $X2=5.725 $Y2=1.905
r246 2 32 600 $w=1.7e-07 $l=6.01581e-07 $layer=licon1_PDIFF $count=1 $X=3.545
+ $Y=2.095 $X2=4.015 $Y2=2.395
r247 1 55 182 $w=1.7e-07 $l=2.95212e-07 $layer=licon1_NDIFF $count=1 $X=3.965
+ $Y=0.625 $X2=4.17 $Y2=0.835
.ends

.subckt PM_SKY130_FD_SC_LP__DFSTP_LP%SET_B 3 7 9 11 12 13 16 20 21 24 26 33 36
+ 38 44
c131 24 0 5.61132e-20 $X=6.48 $Y=1.665
c132 20 0 3.62645e-19 $X=9.695 $Y=1.665
c133 7 0 1.35253e-19 $X=6.595 $Y=0.835
c134 3 0 4.4821e-20 $X=6.27 $Y=2.595
r135 36 39 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=9.865 $Y=1.675
+ $X2=9.865 $Y2=1.84
r136 36 38 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=9.865 $Y=1.675
+ $X2=9.865 $Y2=1.51
r137 36 44 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.865
+ $Y=1.675 $X2=9.865 $Y2=1.675
r138 31 33 10.4917 $w=3.3e-07 $l=6e-08 $layer=POLY_cond $X=6.535 $Y=1.715
+ $X2=6.595 $Y2=1.715
r139 28 31 46.3382 $w=3.3e-07 $l=2.65e-07 $layer=POLY_cond $X=6.27 $Y=1.715
+ $X2=6.535 $Y2=1.715
r140 26 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=1.665
+ $X2=9.84 $Y2=1.665
r141 24 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.535
+ $Y=1.715 $X2=6.535 $Y2=1.715
r142 23 24 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=1.665
+ $X2=6.48 $Y2=1.665
r143 21 23 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.625 $Y=1.665
+ $X2=6.48 $Y2=1.665
r144 20 26 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=9.695 $Y=1.665
+ $X2=9.84 $Y2=1.665
r145 20 21 3.7995 $w=1.4e-07 $l=3.07e-06 $layer=MET1_cond $X=9.695 $Y=1.665
+ $X2=6.625 $Y2=1.665
r146 18 38 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=9.955 $Y=1.27
+ $X2=9.955 $Y2=1.51
r147 16 39 187.582 $w=2.5e-07 $l=7.55e-07 $layer=POLY_cond $X=9.825 $Y=2.595
+ $X2=9.825 $Y2=1.84
r148 12 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.88 $Y=1.195
+ $X2=9.955 $Y2=1.27
r149 12 13 215.362 $w=1.5e-07 $l=4.2e-07 $layer=POLY_cond $X=9.88 $Y=1.195
+ $X2=9.46 $Y2=1.195
r150 9 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.385 $Y=1.12
+ $X2=9.46 $Y2=1.195
r151 9 11 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=9.385 $Y=1.12
+ $X2=9.385 $Y2=0.835
r152 5 33 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.595 $Y=1.55
+ $X2=6.595 $Y2=1.715
r153 5 7 366.628 $w=1.5e-07 $l=7.15e-07 $layer=POLY_cond $X=6.595 $Y=1.55
+ $X2=6.595 $Y2=0.835
r154 1 28 9.34494 $w=2.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.27 $Y=1.88
+ $X2=6.27 $Y2=1.715
r155 1 3 177.644 $w=2.5e-07 $l=7.15e-07 $layer=POLY_cond $X=6.27 $Y=1.88
+ $X2=6.27 $Y2=2.595
.ends

.subckt PM_SKY130_FD_SC_LP__DFSTP_LP%A_266_409# 1 2 9 13 16 17 21 23 26 30 31 32
+ 33 34 37 39 41 42 43 45 49 50 51 52 55 58 61 65 67 69 75 77 83
c207 83 0 5.35053e-20 $X=2.58 $Y=1.68
r208 78 83 47.2125 $w=3.3e-07 $l=2.7e-07 $layer=POLY_cond $X=2.31 $Y=1.68
+ $X2=2.58 $Y2=1.68
r209 78 80 6.99445 $w=3.3e-07 $l=4e-08 $layer=POLY_cond $X=2.31 $Y=1.68 $X2=2.27
+ $Y2=1.68
r210 77 78 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.31
+ $Y=1.68 $X2=2.31 $Y2=1.68
r211 70 75 3.75155 $w=1.7e-07 $l=2.4e-07 $layer=LI1_cond $X=1.64 $Y=2.045
+ $X2=1.4 $Y2=2.045
r212 69 77 13.8292 $w=3.22e-07 $l=4.64844e-07 $layer=LI1_cond $X=2.02 $Y=2.045
+ $X2=2.247 $Y2=1.68
r213 69 70 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=2.02 $Y=2.045
+ $X2=1.64 $Y2=2.045
r214 65 71 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=1.575 $Y=1.185
+ $X2=1.245 $Y2=1.185
r215 65 67 10.4768 $w=3.28e-07 $l=3e-07 $layer=LI1_cond $X=1.575 $Y=1.1
+ $X2=1.575 $Y2=0.8
r216 61 63 17.692 $w=4.78e-07 $l=7.1e-07 $layer=LI1_cond $X=1.4 $Y=2.19 $X2=1.4
+ $Y2=2.9
r217 59 75 2.92809 $w=3.25e-07 $l=8.5e-08 $layer=LI1_cond $X=1.4 $Y=2.13 $X2=1.4
+ $Y2=2.045
r218 59 61 1.4951 $w=4.78e-07 $l=6e-08 $layer=LI1_cond $X=1.4 $Y=2.13 $X2=1.4
+ $Y2=2.19
r219 58 75 2.92809 $w=3.25e-07 $l=1.92873e-07 $layer=LI1_cond $X=1.245 $Y=1.96
+ $X2=1.4 $Y2=2.045
r220 57 71 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.245 $Y=1.27
+ $X2=1.245 $Y2=1.185
r221 57 58 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.245 $Y=1.27
+ $X2=1.245 $Y2=1.96
r222 53 55 141.011 $w=1.5e-07 $l=2.75e-07 $layer=POLY_cond $X=8.065 $Y=1.195
+ $X2=8.34 $Y2=1.195
r223 47 55 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.34 $Y=1.12
+ $X2=8.34 $Y2=1.195
r224 47 49 146.138 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=8.34 $Y=1.12
+ $X2=8.34 $Y2=0.835
r225 46 49 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=8.34 $Y=0.255
+ $X2=8.34 $Y2=0.835
r226 44 53 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.065 $Y=1.27
+ $X2=8.065 $Y2=1.195
r227 44 45 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=8.065 $Y=1.27
+ $X2=8.065 $Y2=1.87
r228 42 45 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.99 $Y=1.945
+ $X2=8.065 $Y2=1.87
r229 42 43 133.319 $w=1.5e-07 $l=2.6e-07 $layer=POLY_cond $X=7.99 $Y=1.945
+ $X2=7.73 $Y2=1.945
r230 39 43 29.1797 $w=1.5e-07 $l=1.58114e-07 $layer=POLY_cond $X=7.605 $Y=2.02
+ $X2=7.73 $Y2=1.945
r231 39 41 110.86 $w=2.5e-07 $l=5.75e-07 $layer=POLY_cond $X=7.605 $Y=2.02
+ $X2=7.605 $Y2=2.595
r232 35 37 156.526 $w=2.5e-07 $l=6.3e-07 $layer=POLY_cond $X=4.28 $Y=1.965
+ $X2=4.28 $Y2=2.595
r233 33 46 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.265 $Y=0.18
+ $X2=8.34 $Y2=0.255
r234 33 34 2204.89 $w=1.5e-07 $l=4.3e-06 $layer=POLY_cond $X=8.265 $Y=0.18
+ $X2=3.965 $Y2=0.18
r235 31 35 29.1797 $w=1.5e-07 $l=1.58114e-07 $layer=POLY_cond $X=4.155 $Y=1.89
+ $X2=4.28 $Y2=1.965
r236 31 32 112.809 $w=1.5e-07 $l=2.2e-07 $layer=POLY_cond $X=4.155 $Y=1.89
+ $X2=3.935 $Y2=1.89
r237 28 52 20.4101 $w=1.5e-07 $l=8.21584e-08 $layer=POLY_cond $X=3.89 $Y=1.12
+ $X2=3.875 $Y2=1.195
r238 28 30 146.138 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.89 $Y=1.12
+ $X2=3.89 $Y2=0.835
r239 27 34 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.89 $Y=0.255
+ $X2=3.965 $Y2=0.18
r240 27 30 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=3.89 $Y=0.255
+ $X2=3.89 $Y2=0.835
r241 26 32 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.86 $Y=1.815
+ $X2=3.935 $Y2=1.89
r242 25 52 20.4101 $w=1.5e-07 $l=8.21584e-08 $layer=POLY_cond $X=3.86 $Y=1.27
+ $X2=3.875 $Y2=1.195
r243 25 26 279.457 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=3.86 $Y=1.27
+ $X2=3.86 $Y2=1.815
r244 24 51 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.015 $Y=1.195
+ $X2=2.94 $Y2=1.195
r245 23 52 5.30422 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.785 $Y=1.195
+ $X2=3.875 $Y2=1.195
r246 23 24 394.83 $w=1.5e-07 $l=7.7e-07 $layer=POLY_cond $X=3.785 $Y=1.195
+ $X2=3.015 $Y2=1.195
r247 19 51 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.94 $Y=1.12
+ $X2=2.94 $Y2=1.195
r248 19 21 187.16 $w=1.5e-07 $l=3.65e-07 $layer=POLY_cond $X=2.94 $Y=1.12
+ $X2=2.94 $Y2=0.755
r249 18 50 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.655 $Y=1.195
+ $X2=2.58 $Y2=1.195
r250 17 51 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.865 $Y=1.195
+ $X2=2.94 $Y2=1.195
r251 17 18 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=2.865 $Y=1.195
+ $X2=2.655 $Y2=1.195
r252 16 83 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.58 $Y=1.515
+ $X2=2.58 $Y2=1.68
r253 15 50 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.58 $Y=1.27
+ $X2=2.58 $Y2=1.195
r254 15 16 125.628 $w=1.5e-07 $l=2.45e-07 $layer=POLY_cond $X=2.58 $Y=1.27
+ $X2=2.58 $Y2=1.515
r255 11 50 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.58 $Y=1.12
+ $X2=2.58 $Y2=1.195
r256 11 13 187.16 $w=1.5e-07 $l=3.65e-07 $layer=POLY_cond $X=2.58 $Y=1.12
+ $X2=2.58 $Y2=0.755
r257 7 80 9.34494 $w=2.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.27 $Y=1.845
+ $X2=2.27 $Y2=1.68
r258 7 9 173.918 $w=2.5e-07 $l=7e-07 $layer=POLY_cond $X=2.27 $Y=1.845 $X2=2.27
+ $Y2=2.545
r259 2 63 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=1.33
+ $Y=2.045 $X2=1.475 $Y2=2.9
r260 2 61 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=1.33
+ $Y=2.045 $X2=1.475 $Y2=2.19
r261 1 67 182 $w=1.7e-07 $l=3.13329e-07 $layer=licon1_NDIFF $count=1 $X=1.445
+ $Y=0.545 $X2=1.575 $Y2=0.8
.ends

.subckt PM_SKY130_FD_SC_LP__DFSTP_LP%A_1731_99# 1 2 7 9 11 14 18 22 23 25 26 29
+ 33 35 40 42
c95 23 0 1.16491e-20 $X=9.325 $Y=1.675
r96 43 45 8.74306 $w=3.3e-07 $l=5e-08 $layer=POLY_cond $X=8.995 $Y=1.675
+ $X2=9.045 $Y2=1.675
r97 35 37 32.7294 $w=2.48e-07 $l=7.1e-07 $layer=LI1_cond $X=10.61 $Y=1.84
+ $X2=10.61 $Y2=2.55
r98 33 42 6.94937 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=10.61 $Y=1.8
+ $X2=10.61 $Y2=1.675
r99 33 35 1.84391 $w=2.48e-07 $l=4e-08 $layer=LI1_cond $X=10.61 $Y=1.8 $X2=10.61
+ $Y2=1.84
r100 31 40 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.57 $Y=1.33
+ $X2=10.57 $Y2=1.245
r101 31 42 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=10.57 $Y=1.33
+ $X2=10.57 $Y2=1.675
r102 27 40 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=10.23 $Y=1.245
+ $X2=10.57 $Y2=1.245
r103 27 29 24.0965 $w=3.28e-07 $l=6.9e-07 $layer=LI1_cond $X=10.23 $Y=1.16
+ $X2=10.23 $Y2=0.47
r104 25 27 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=10.065 $Y=1.245
+ $X2=10.23 $Y2=1.245
r105 25 26 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=10.065 $Y=1.245
+ $X2=9.49 $Y2=1.245
r106 23 45 48.9612 $w=3.3e-07 $l=2.8e-07 $layer=POLY_cond $X=9.325 $Y=1.675
+ $X2=9.045 $Y2=1.675
r107 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.325
+ $Y=1.675 $X2=9.325 $Y2=1.675
r108 20 26 7.55824 $w=1.7e-07 $l=1.90825e-07 $layer=LI1_cond $X=9.337 $Y=1.33
+ $X2=9.49 $Y2=1.245
r109 20 22 13.0358 $w=3.03e-07 $l=3.45e-07 $layer=LI1_cond $X=9.337 $Y=1.33
+ $X2=9.337 $Y2=1.675
r110 16 18 135.883 $w=1.5e-07 $l=2.65e-07 $layer=POLY_cond $X=8.73 $Y=1.195
+ $X2=8.995 $Y2=1.195
r111 12 45 9.34494 $w=2.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.045 $Y=1.84
+ $X2=9.045 $Y2=1.675
r112 12 14 187.582 $w=2.5e-07 $l=7.55e-07 $layer=POLY_cond $X=9.045 $Y=1.84
+ $X2=9.045 $Y2=2.595
r113 11 43 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.995 $Y=1.51
+ $X2=8.995 $Y2=1.675
r114 10 18 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.995 $Y=1.27
+ $X2=8.995 $Y2=1.195
r115 10 11 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=8.995 $Y=1.27
+ $X2=8.995 $Y2=1.51
r116 7 16 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.73 $Y=1.12
+ $X2=8.73 $Y2=1.195
r117 7 9 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=8.73 $Y=1.12 $X2=8.73
+ $Y2=0.835
r118 2 37 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=10.505
+ $Y=1.695 $X2=10.65 $Y2=2.55
r119 2 35 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=10.505
+ $Y=1.695 $X2=10.65 $Y2=1.84
r120 1 29 182 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_NDIFF $count=1 $X=10.085
+ $Y=0.235 $X2=10.23 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_LP__DFSTP_LP%A_1526_125# 1 2 3 10 12 13 14 15 17 20 22
+ 26 28 32 36 39 41 42 43 46 48 50 51 53 54 59 60 61 64 65 67 68 70 74
c180 67 0 1.56847e-19 $X=11 $Y=1.495
r181 70 72 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=8.125 $Y=0.835
+ $X2=8.125 $Y2=0.98
r182 67 68 91.3369 $w=1.68e-07 $l=1.4e-06 $layer=LI1_cond $X=11 $Y=1.495 $X2=11
+ $Y2=2.895
r183 64 65 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=11 $Y=0.99
+ $X2=11 $Y2=0.99
r184 62 67 7.1122 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=11 $Y=1.33 $X2=11
+ $Y2=1.495
r185 62 64 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=11 $Y=1.33 $X2=11
+ $Y2=0.99
r186 60 68 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.915 $Y=2.98
+ $X2=11 $Y2=2.895
r187 60 61 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=10.915 $Y=2.98
+ $X2=10.255 $Y2=2.98
r188 57 61 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=10.09 $Y=2.895
+ $X2=10.255 $Y2=2.98
r189 57 59 22.8742 $w=3.28e-07 $l=6.55e-07 $layer=LI1_cond $X=10.09 $Y=2.895
+ $X2=10.09 $Y2=2.24
r190 56 59 1.74613 $w=3.28e-07 $l=5e-08 $layer=LI1_cond $X=10.09 $Y=2.19
+ $X2=10.09 $Y2=2.24
r191 55 74 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.005 $Y=2.105
+ $X2=8.92 $Y2=2.105
r192 54 56 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=9.925 $Y=2.105
+ $X2=10.09 $Y2=2.19
r193 54 55 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=9.925 $Y=2.105
+ $X2=9.005 $Y2=2.105
r194 53 74 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.92 $Y=2.02
+ $X2=8.92 $Y2=2.105
r195 52 53 62.3048 $w=1.68e-07 $l=9.55e-07 $layer=LI1_cond $X=8.92 $Y=1.065
+ $X2=8.92 $Y2=2.02
r196 50 74 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.835 $Y=2.105
+ $X2=8.92 $Y2=2.105
r197 50 51 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=8.835 $Y=2.105
+ $X2=8.375 $Y2=2.105
r198 49 72 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.29 $Y=0.98
+ $X2=8.125 $Y2=0.98
r199 48 52 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.835 $Y=0.98
+ $X2=8.92 $Y2=1.065
r200 48 49 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=8.835 $Y=0.98
+ $X2=8.29 $Y2=0.98
r201 44 51 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=8.21 $Y=2.19
+ $X2=8.375 $Y2=2.105
r202 44 46 1.74613 $w=3.28e-07 $l=5e-08 $layer=LI1_cond $X=8.21 $Y=2.19 $X2=8.21
+ $Y2=2.24
r203 40 65 45.3873 $w=4.35e-07 $l=3.55e-07 $layer=POLY_cond $X=10.947 $Y=1.345
+ $X2=10.947 $Y2=0.99
r204 40 41 9.82482 $w=3.42e-07 $l=7.5e-08 $layer=POLY_cond $X=10.947 $Y=1.345
+ $X2=10.947 $Y2=1.42
r205 38 65 14.0637 $w=4.35e-07 $l=1.1e-07 $layer=POLY_cond $X=10.947 $Y=0.88
+ $X2=10.947 $Y2=0.99
r206 38 39 11.361 $w=2.92e-07 $l=2.82204e-07 $layer=POLY_cond $X=10.947 $Y=0.88
+ $X2=10.73 $Y2=0.73
r207 34 43 15.9654 $w=2e-07 $l=8.44097e-08 $layer=POLY_cond $X=12.155 $Y=1.345
+ $X2=12.175 $Y2=1.42
r208 34 36 392.266 $w=1.5e-07 $l=7.65e-07 $layer=POLY_cond $X=12.155 $Y=1.345
+ $X2=12.155 $Y2=0.58
r209 30 43 15.9654 $w=2e-07 $l=7.5e-08 $layer=POLY_cond $X=12.175 $Y=1.495
+ $X2=12.175 $Y2=1.42
r210 30 32 217.397 $w=2.5e-07 $l=8.75e-07 $layer=POLY_cond $X=12.175 $Y=1.495
+ $X2=12.175 $Y2=2.37
r211 29 42 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=11.87 $Y=1.42
+ $X2=11.795 $Y2=1.42
r212 28 43 9.46703 $w=1.5e-07 $l=1.25e-07 $layer=POLY_cond $X=12.05 $Y=1.42
+ $X2=12.175 $Y2=1.42
r213 28 29 92.2979 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=12.05 $Y=1.42
+ $X2=11.87 $Y2=1.42
r214 24 42 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=11.795 $Y=1.345
+ $X2=11.795 $Y2=1.42
r215 24 26 392.266 $w=1.5e-07 $l=7.65e-07 $layer=POLY_cond $X=11.795 $Y=1.345
+ $X2=11.795 $Y2=0.58
r216 23 41 17.4961 $w=1.5e-07 $l=2.18e-07 $layer=POLY_cond $X=11.165 $Y=1.42
+ $X2=10.947 $Y2=1.42
r217 22 42 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=11.72 $Y=1.42
+ $X2=11.795 $Y2=1.42
r218 22 23 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=11.72 $Y=1.42
+ $X2=11.165 $Y2=1.42
r219 18 41 9.82482 $w=3.42e-07 $l=8.95824e-08 $layer=POLY_cond $X=10.915
+ $Y=1.495 $X2=10.947 $Y2=1.42
r220 18 20 173.918 $w=2.5e-07 $l=7e-07 $layer=POLY_cond $X=10.915 $Y=1.495
+ $X2=10.915 $Y2=2.195
r221 15 39 11.361 $w=2.92e-07 $l=7.5e-08 $layer=POLY_cond $X=10.805 $Y=0.73
+ $X2=10.73 $Y2=0.73
r222 15 17 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=10.805 $Y=0.73
+ $X2=10.805 $Y2=0.445
r223 13 39 15.119 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=10.73 $Y=0.805
+ $X2=10.73 $Y2=0.73
r224 13 14 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=10.73 $Y=0.805
+ $X2=10.52 $Y2=0.805
r225 10 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=10.445 $Y=0.73
+ $X2=10.52 $Y2=0.805
r226 10 12 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=10.445 $Y=0.73
+ $X2=10.445 $Y2=0.445
r227 3 59 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=9.95
+ $Y=2.095 $X2=10.09 $Y2=2.24
r228 2 46 300 $w=1.7e-07 $l=5.47723e-07 $layer=licon1_PDIFF $count=2 $X=7.73
+ $Y=2.095 $X2=8.21 $Y2=2.24
r229 1 70 182 $w=1.7e-07 $l=5.90741e-07 $layer=licon1_NDIFF $count=1 $X=7.63
+ $Y=0.625 $X2=8.125 $Y2=0.835
.ends

.subckt PM_SKY130_FD_SC_LP__DFSTP_LP%A_2287_74# 1 2 9 13 17 23 26 28 31 35 39 40
+ 45 47
c72 47 0 2.21704e-19 $X=11.885 $Y=1.575
c73 26 0 7.71418e-20 $X=12.675 $Y=1.66
r74 43 45 5.20034 $w=4.58e-07 $l=2e-07 $layer=LI1_cond $X=11.58 $Y=0.58
+ $X2=11.78 $Y2=0.58
r75 39 40 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=12.675
+ $Y=1.155 $X2=12.675 $Y2=1.155
r76 37 39 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=12.675 $Y=1.49
+ $X2=12.675 $Y2=1.155
r77 36 47 3.11956 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=12.075 $Y=1.575
+ $X2=11.885 $Y2=1.575
r78 35 37 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=12.51 $Y=1.575
+ $X2=12.675 $Y2=1.49
r79 35 36 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=12.51 $Y=1.575
+ $X2=12.075 $Y2=1.575
r80 31 33 21.5325 $w=3.78e-07 $l=7.1e-07 $layer=LI1_cond $X=11.885 $Y=2.015
+ $X2=11.885 $Y2=2.725
r81 29 47 3.40559 $w=2.75e-07 $l=8.5e-08 $layer=LI1_cond $X=11.885 $Y=1.66
+ $X2=11.885 $Y2=1.575
r82 29 31 10.7662 $w=3.78e-07 $l=3.55e-07 $layer=LI1_cond $X=11.885 $Y=1.66
+ $X2=11.885 $Y2=2.015
r83 28 47 3.40559 $w=2.75e-07 $l=1.41244e-07 $layer=LI1_cond $X=11.78 $Y=1.49
+ $X2=11.885 $Y2=1.575
r84 27 45 6.6364 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=11.78 $Y=0.81
+ $X2=11.78 $Y2=0.58
r85 27 28 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=11.78 $Y=0.81
+ $X2=11.78 $Y2=1.49
r86 25 40 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=12.675 $Y=1.495
+ $X2=12.675 $Y2=1.155
r87 25 26 31.6748 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=12.675 $Y=1.495
+ $X2=12.675 $Y2=1.66
r88 22 40 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=12.675 $Y=1.14
+ $X2=12.675 $Y2=1.155
r89 22 23 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=12.675 $Y=1.065
+ $X2=12.945 $Y2=1.065
r90 19 22 46.1489 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=12.585 $Y=1.065
+ $X2=12.675 $Y2=1.065
r91 15 23 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=12.945 $Y=0.99
+ $X2=12.945 $Y2=1.065
r92 15 17 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=12.945 $Y=0.99
+ $X2=12.945 $Y2=0.58
r93 13 26 176.402 $w=2.5e-07 $l=7.1e-07 $layer=POLY_cond $X=12.705 $Y=2.37
+ $X2=12.705 $Y2=1.66
r94 7 19 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=12.585 $Y=0.99
+ $X2=12.585 $Y2=1.065
r95 7 9 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=12.585 $Y=0.99
+ $X2=12.585 $Y2=0.58
r96 2 33 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=11.765
+ $Y=1.87 $X2=11.91 $Y2=2.725
r97 2 31 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=11.765
+ $Y=1.87 $X2=11.91 $Y2=2.015
r98 1 43 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=11.435
+ $Y=0.37 $X2=11.58 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_LP__DFSTP_LP%VPWR 1 2 3 4 5 6 7 22 24 30 34 38 42 46 52
+ 57 58 59 61 69 74 82 87 97 98 104 107 110 113 116
r145 116 117 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.28 $Y=3.33
+ $X2=11.28 $Y2=3.33
r146 113 114 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r147 110 111 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r148 107 108 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r149 104 105 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r150 101 102 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r151 97 98 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=13.2 $Y=3.33
+ $X2=13.2 $Y2=3.33
r152 95 98 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=12.24 $Y=3.33
+ $X2=13.2 $Y2=3.33
r153 95 117 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=12.24 $Y=3.33
+ $X2=11.28 $Y2=3.33
r154 94 95 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=12.24 $Y=3.33
+ $X2=12.24 $Y2=3.33
r155 92 116 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=11.515 $Y=3.33
+ $X2=11.39 $Y2=3.33
r156 92 94 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=11.515 $Y=3.33
+ $X2=12.24 $Y2=3.33
r157 91 117 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=9.84 $Y=3.33
+ $X2=11.28 $Y2=3.33
r158 91 114 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.84 $Y=3.33
+ $X2=9.36 $Y2=3.33
r159 90 91 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r160 88 113 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.475 $Y=3.33
+ $X2=9.31 $Y2=3.33
r161 88 90 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=9.475 $Y=3.33
+ $X2=9.84 $Y2=3.33
r162 87 116 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=11.265 $Y=3.33
+ $X2=11.39 $Y2=3.33
r163 87 90 92.9679 $w=1.68e-07 $l=1.425e-06 $layer=LI1_cond $X=11.265 $Y=3.33
+ $X2=9.84 $Y2=3.33
r164 86 114 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=9.36 $Y2=3.33
r165 86 111 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=6.96 $Y2=3.33
r166 85 86 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r167 83 110 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.015 $Y=3.33
+ $X2=6.85 $Y2=3.33
r168 83 85 121.674 $w=1.68e-07 $l=1.865e-06 $layer=LI1_cond $X=7.015 $Y=3.33
+ $X2=8.88 $Y2=3.33
r169 82 113 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.145 $Y=3.33
+ $X2=9.31 $Y2=3.33
r170 82 85 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=9.145 $Y=3.33
+ $X2=8.88 $Y2=3.33
r171 80 81 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r172 78 81 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=6.48 $Y2=3.33
r173 78 108 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=5.04 $Y2=3.33
r174 77 80 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=5.52 $Y=3.33
+ $X2=6.48 $Y2=3.33
r175 77 78 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r176 75 107 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.27 $Y=3.33
+ $X2=5.105 $Y2=3.33
r177 75 77 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=5.27 $Y=3.33
+ $X2=5.52 $Y2=3.33
r178 74 110 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.685 $Y=3.33
+ $X2=6.85 $Y2=3.33
r179 74 80 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=6.685 $Y=3.33
+ $X2=6.48 $Y2=3.33
r180 73 108 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.04 $Y2=3.33
r181 73 105 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=2.16 $Y2=3.33
r182 72 73 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r183 70 104 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.17 $Y=3.33
+ $X2=2.005 $Y2=3.33
r184 70 72 155.925 $w=1.68e-07 $l=2.39e-06 $layer=LI1_cond $X=2.17 $Y=3.33
+ $X2=4.56 $Y2=3.33
r185 69 107 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.94 $Y=3.33
+ $X2=5.105 $Y2=3.33
r186 69 72 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=4.94 $Y=3.33
+ $X2=4.56 $Y2=3.33
r187 68 105 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r188 67 68 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r189 65 68 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r190 65 102 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r191 64 67 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r192 64 65 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r193 62 101 4.72267 $w=1.7e-07 $l=2.25e-07 $layer=LI1_cond $X=0.45 $Y=3.33
+ $X2=0.225 $Y2=3.33
r194 62 64 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=0.45 $Y=3.33
+ $X2=0.72 $Y2=3.33
r195 61 104 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.84 $Y=3.33
+ $X2=2.005 $Y2=3.33
r196 61 67 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=1.84 $Y=3.33
+ $X2=1.68 $Y2=3.33
r197 59 111 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=6.72 $Y=3.33
+ $X2=6.96 $Y2=3.33
r198 59 81 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=6.72 $Y=3.33
+ $X2=6.48 $Y2=3.33
r199 57 94 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=12.275 $Y=3.33
+ $X2=12.24 $Y2=3.33
r200 57 58 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.275 $Y=3.33
+ $X2=12.44 $Y2=3.33
r201 56 97 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=12.605 $Y=3.33
+ $X2=13.2 $Y2=3.33
r202 56 58 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.605 $Y=3.33
+ $X2=12.44 $Y2=3.33
r203 52 55 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=12.44 $Y=2.015
+ $X2=12.44 $Y2=2.725
r204 50 58 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=12.44 $Y=3.245
+ $X2=12.44 $Y2=3.33
r205 50 55 18.1597 $w=3.28e-07 $l=5.2e-07 $layer=LI1_cond $X=12.44 $Y=3.245
+ $X2=12.44 $Y2=2.725
r206 46 49 32.7294 $w=2.48e-07 $l=7.1e-07 $layer=LI1_cond $X=11.39 $Y=1.84
+ $X2=11.39 $Y2=2.55
r207 44 116 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=11.39 $Y=3.245
+ $X2=11.39 $Y2=3.33
r208 44 49 32.0379 $w=2.48e-07 $l=6.95e-07 $layer=LI1_cond $X=11.39 $Y=3.245
+ $X2=11.39 $Y2=2.55
r209 40 113 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.31 $Y=3.245
+ $X2=9.31 $Y2=3.33
r210 40 42 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=9.31 $Y=3.245
+ $X2=9.31 $Y2=2.535
r211 36 110 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.85 $Y=3.245
+ $X2=6.85 $Y2=3.33
r212 36 38 23.3981 $w=3.28e-07 $l=6.7e-07 $layer=LI1_cond $X=6.85 $Y=3.245
+ $X2=6.85 $Y2=2.575
r213 32 107 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.105 $Y=3.245
+ $X2=5.105 $Y2=3.33
r214 32 34 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=5.105 $Y=3.245
+ $X2=5.105 $Y2=2.95
r215 28 104 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.005 $Y=3.245
+ $X2=2.005 $Y2=3.33
r216 28 30 26.8903 $w=3.28e-07 $l=7.7e-07 $layer=LI1_cond $X=2.005 $Y=3.245
+ $X2=2.005 $Y2=2.475
r217 24 27 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=0.285 $Y=2.19
+ $X2=0.285 $Y2=2.9
r218 22 101 3.0435 $w=3.3e-07 $l=1.11018e-07 $layer=LI1_cond $X=0.285 $Y=3.245
+ $X2=0.225 $Y2=3.33
r219 22 27 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=0.285 $Y=3.245
+ $X2=0.285 $Y2=2.9
r220 7 55 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=12.3
+ $Y=1.87 $X2=12.44 $Y2=2.725
r221 7 52 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=12.3
+ $Y=1.87 $X2=12.44 $Y2=2.015
r222 6 49 400 $w=1.7e-07 $l=9.98036e-07 $layer=licon1_PDIFF $count=1 $X=11.04
+ $Y=1.695 $X2=11.35 $Y2=2.55
r223 6 46 400 $w=1.7e-07 $l=3.75566e-07 $layer=licon1_PDIFF $count=1 $X=11.04
+ $Y=1.695 $X2=11.35 $Y2=1.84
r224 5 42 300 $w=1.7e-07 $l=5.05173e-07 $layer=licon1_PDIFF $count=2 $X=9.17
+ $Y=2.095 $X2=9.31 $Y2=2.535
r225 4 38 300 $w=1.7e-07 $l=6.69925e-07 $layer=licon1_PDIFF $count=2 $X=6.395
+ $Y=2.095 $X2=6.85 $Y2=2.575
r226 3 34 600 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=4.965
+ $Y=2.095 $X2=5.105 $Y2=2.95
r227 2 30 300 $w=1.7e-07 $l=4.95076e-07 $layer=licon1_PDIFF $count=2 $X=1.865
+ $Y=2.045 $X2=2.005 $Y2=2.475
r228 1 27 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.14
+ $Y=2.045 $X2=0.285 $Y2=2.9
r229 1 24 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.14
+ $Y=2.045 $X2=0.285 $Y2=2.19
.ends

.subckt PM_SKY130_FD_SC_LP__DFSTP_LP%A_135_409# 1 2 3 4 15 17 21 24 26 27 28 30
+ 33 35 36 42 47
c106 21 0 1.1902e-19 $X=1.93 $Y=0.35
r107 44 47 5.04596 $w=6.38e-07 $l=2.7e-07 $layer=LI1_cond $X=2.885 $Y=2.395
+ $X2=3.155 $Y2=2.395
r108 42 43 9.73709 $w=2.13e-07 $l=1.7e-07 $layer=LI1_cond $X=2.715 $Y=1.217
+ $X2=2.885 $Y2=1.217
r109 41 42 40.0939 $w=2.13e-07 $l=7e-07 $layer=LI1_cond $X=2.015 $Y=1.217
+ $X2=2.715 $Y2=1.217
r110 39 40 10.5184 $w=4.03e-07 $l=2.3e-07 $layer=LI1_cond $X=1.012 $Y=0.495
+ $X2=1.012 $Y2=0.725
r111 36 39 4.12603 $w=4.03e-07 $l=1.45e-07 $layer=LI1_cond $X=1.012 $Y=0.35
+ $X2=1.012 $Y2=0.495
r112 35 40 84.8128 $w=1.68e-07 $l=1.3e-06 $layer=LI1_cond $X=0.895 $Y=2.025
+ $X2=0.895 $Y2=0.725
r113 31 33 13.969 $w=3.28e-07 $l=4e-07 $layer=LI1_cond $X=3.675 $Y=0.435
+ $X2=3.675 $Y2=0.835
r114 30 44 8.73481 $w=1.7e-07 $l=3.2e-07 $layer=LI1_cond $X=2.885 $Y=2.075
+ $X2=2.885 $Y2=2.395
r115 29 43 2.0603 $w=1.7e-07 $l=1.18e-07 $layer=LI1_cond $X=2.885 $Y=1.335
+ $X2=2.885 $Y2=1.217
r116 29 30 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=2.885 $Y=1.335
+ $X2=2.885 $Y2=2.075
r117 27 31 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.51 $Y=0.35
+ $X2=3.675 $Y2=0.435
r118 27 28 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=3.51 $Y=0.35
+ $X2=2.8 $Y2=0.35
r119 26 42 2.0603 $w=1.7e-07 $l=1.17e-07 $layer=LI1_cond $X=2.715 $Y=1.1
+ $X2=2.715 $Y2=1.217
r120 25 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.715 $Y=0.435
+ $X2=2.8 $Y2=0.35
r121 25 26 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=2.715 $Y=0.435
+ $X2=2.715 $Y2=1.1
r122 24 41 2.0603 $w=1.7e-07 $l=1.17e-07 $layer=LI1_cond $X=2.015 $Y=1.1
+ $X2=2.015 $Y2=1.217
r123 23 24 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=2.015 $Y=0.435
+ $X2=2.015 $Y2=1.1
r124 22 36 5.85399 $w=1.7e-07 $l=2.03e-07 $layer=LI1_cond $X=1.215 $Y=0.35
+ $X2=1.012 $Y2=0.35
r125 21 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.93 $Y=0.35
+ $X2=2.015 $Y2=0.435
r126 21 22 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=1.93 $Y=0.35
+ $X2=1.215 $Y2=0.35
r127 15 35 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.815 $Y=2.19
+ $X2=0.815 $Y2=2.025
r128 15 17 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=0.815 $Y=2.19
+ $X2=0.815 $Y2=2.9
r129 4 47 600 $w=1.7e-07 $l=3.65377e-07 $layer=licon1_PDIFF $count=1 $X=3.01
+ $Y=2.095 $X2=3.155 $Y2=2.395
r130 3 17 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=0.675
+ $Y=2.045 $X2=0.815 $Y2=2.9
r131 3 15 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.675
+ $Y=2.045 $X2=0.815 $Y2=2.19
r132 2 33 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=3.55
+ $Y=0.625 $X2=3.675 $Y2=0.835
r133 1 39 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.91
+ $Y=0.285 $X2=1.05 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__DFSTP_LP%Q 1 2 7 8 9 10 11 12 13 45 49
c22 45 0 7.71418e-20 $X=12.97 $Y=2.015
r23 45 46 7.29421 $w=5.18e-07 $l=1.65e-07 $layer=LI1_cond $X=13.065 $Y=2.015
+ $X2=13.065 $Y2=1.85
r24 30 49 1.72511 $w=5.18e-07 $l=7.5e-08 $layer=LI1_cond $X=13.065 $Y=2.11
+ $X2=13.065 $Y2=2.035
r25 13 35 1.15008 $w=5.18e-07 $l=5e-08 $layer=LI1_cond $X=13.065 $Y=2.775
+ $X2=13.065 $Y2=2.725
r26 12 35 7.36048 $w=5.18e-07 $l=3.2e-07 $layer=LI1_cond $X=13.065 $Y=2.405
+ $X2=13.065 $Y2=2.725
r27 11 49 0.115008 $w=5.18e-07 $l=5e-09 $layer=LI1_cond $X=13.065 $Y=2.03
+ $X2=13.065 $Y2=2.035
r28 11 45 0.345023 $w=5.18e-07 $l=1.5e-08 $layer=LI1_cond $X=13.065 $Y=2.03
+ $X2=13.065 $Y2=2.015
r29 11 12 6.67044 $w=5.18e-07 $l=2.9e-07 $layer=LI1_cond $X=13.065 $Y=2.115
+ $X2=13.065 $Y2=2.405
r30 11 30 0.115008 $w=5.18e-07 $l=5e-09 $layer=LI1_cond $X=13.065 $Y=2.115
+ $X2=13.065 $Y2=2.11
r31 10 46 8.88342 $w=2.38e-07 $l=1.85e-07 $layer=LI1_cond $X=13.205 $Y=1.665
+ $X2=13.205 $Y2=1.85
r32 9 10 17.7668 $w=2.38e-07 $l=3.7e-07 $layer=LI1_cond $X=13.205 $Y=1.295
+ $X2=13.205 $Y2=1.665
r33 8 9 17.7668 $w=2.38e-07 $l=3.7e-07 $layer=LI1_cond $X=13.205 $Y=0.925
+ $X2=13.205 $Y2=1.295
r34 8 43 5.52212 $w=2.38e-07 $l=1.15e-07 $layer=LI1_cond $X=13.205 $Y=0.925
+ $X2=13.205 $Y2=0.81
r35 7 43 9.78297 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=13.16 $Y=0.555
+ $X2=13.16 $Y2=0.81
r36 2 45 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=12.83
+ $Y=1.87 $X2=12.97 $Y2=2.015
r37 2 35 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=12.83
+ $Y=1.87 $X2=12.97 $Y2=2.725
r38 1 7 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=13.02
+ $Y=0.37 $X2=13.16 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_LP__DFSTP_LP%VGND 1 2 3 4 5 6 7 22 24 28 32 36 40 44 48
+ 51 52 54 55 57 58 59 68 75 93 99 100 106 109 112
c138 40 0 2.00657e-19 $X=9.6 $Y=0.79
r139 112 113 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=12.24 $Y=0
+ $X2=12.24 $Y2=0
r140 109 110 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=6.96 $Y=0
+ $X2=6.96 $Y2=0
r141 106 107 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0
+ $X2=5.04 $Y2=0
r142 103 104 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0
+ $X2=0.24 $Y2=0
r143 100 113 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=13.2 $Y=0
+ $X2=12.24 $Y2=0
r144 99 100 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=13.2 $Y=0
+ $X2=13.2 $Y2=0
r145 97 112 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.535 $Y=0
+ $X2=12.37 $Y2=0
r146 97 99 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=12.535 $Y=0
+ $X2=13.2 $Y2=0
r147 96 113 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=11.28 $Y=0
+ $X2=12.24 $Y2=0
r148 95 96 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=11.28 $Y=0
+ $X2=11.28 $Y2=0
r149 93 112 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.205 $Y=0
+ $X2=12.37 $Y2=0
r150 93 95 60.3476 $w=1.68e-07 $l=9.25e-07 $layer=LI1_cond $X=12.205 $Y=0
+ $X2=11.28 $Y2=0
r151 92 96 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.8 $Y=0
+ $X2=11.28 $Y2=0
r152 91 92 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=10.8 $Y=0 $X2=10.8
+ $Y2=0
r153 89 92 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=9.84 $Y=0 $X2=10.8
+ $Y2=0
r154 88 91 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=9.84 $Y=0 $X2=10.8
+ $Y2=0
r155 88 89 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=9.84 $Y=0 $X2=9.84
+ $Y2=0
r156 86 89 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=0 $X2=9.84
+ $Y2=0
r157 86 110 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=9.36 $Y=0
+ $X2=6.96 $Y2=0
r158 85 86 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=9.36 $Y=0 $X2=9.36
+ $Y2=0
r159 83 109 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.015 $Y=0
+ $X2=6.85 $Y2=0
r160 83 85 152.989 $w=1.68e-07 $l=2.345e-06 $layer=LI1_cond $X=7.015 $Y=0
+ $X2=9.36 $Y2=0
r161 81 82 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r162 79 82 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=6.48
+ $Y2=0
r163 79 107 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0
+ $X2=5.04 $Y2=0
r164 78 81 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=5.52 $Y=0 $X2=6.48
+ $Y2=0
r165 78 79 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r166 76 106 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.165 $Y=0
+ $X2=5.04 $Y2=0
r167 76 78 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=5.165 $Y=0
+ $X2=5.52 $Y2=0
r168 75 109 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.685 $Y=0
+ $X2=6.85 $Y2=0
r169 75 81 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=6.685 $Y=0
+ $X2=6.48 $Y2=0
r170 74 107 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0
+ $X2=5.04 $Y2=0
r171 73 74 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.56 $Y=0
+ $X2=4.56 $Y2=0
r172 71 74 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=2.64 $Y=0
+ $X2=4.56 $Y2=0
r173 70 73 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=2.64 $Y=0 $X2=4.56
+ $Y2=0
r174 70 71 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.64 $Y=0
+ $X2=2.64 $Y2=0
r175 68 106 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.915 $Y=0
+ $X2=5.04 $Y2=0
r176 68 73 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=4.915 $Y=0
+ $X2=4.56 $Y2=0
r177 67 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r178 66 67 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r179 64 67 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=0.72 $Y=0
+ $X2=2.16 $Y2=0
r180 64 104 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0
+ $X2=0.24 $Y2=0
r181 63 66 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=0.72 $Y=0 $X2=2.16
+ $Y2=0
r182 63 64 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r183 61 103 4.78091 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=0
+ $X2=0.212 $Y2=0
r184 61 63 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.425 $Y=0 $X2=0.72
+ $Y2=0
r185 59 110 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=6.72 $Y=0
+ $X2=6.96 $Y2=0
r186 59 82 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=6.72 $Y=0
+ $X2=6.48 $Y2=0
r187 57 91 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=10.855 $Y=0
+ $X2=10.8 $Y2=0
r188 57 58 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.855 $Y=0
+ $X2=11.02 $Y2=0
r189 56 95 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=11.185 $Y=0
+ $X2=11.28 $Y2=0
r190 56 58 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.185 $Y=0
+ $X2=11.02 $Y2=0
r191 54 85 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=9.435 $Y=0 $X2=9.36
+ $Y2=0
r192 54 55 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.435 $Y=0 $X2=9.6
+ $Y2=0
r193 53 88 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=9.765 $Y=0 $X2=9.84
+ $Y2=0
r194 53 55 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.765 $Y=0 $X2=9.6
+ $Y2=0
r195 51 66 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=2.28 $Y=0 $X2=2.16
+ $Y2=0
r196 51 52 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.28 $Y=0 $X2=2.365
+ $Y2=0
r197 50 70 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=2.45 $Y=0 $X2=2.64
+ $Y2=0
r198 50 52 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.45 $Y=0 $X2=2.365
+ $Y2=0
r199 46 112 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=12.37 $Y=0.085
+ $X2=12.37 $Y2=0
r200 46 48 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=12.37 $Y=0.085
+ $X2=12.37 $Y2=0.58
r201 42 58 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=11.02 $Y=0.085
+ $X2=11.02 $Y2=0
r202 42 44 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=11.02 $Y=0.085
+ $X2=11.02 $Y2=0.43
r203 38 55 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.6 $Y=0.085 $X2=9.6
+ $Y2=0
r204 38 40 24.6204 $w=3.28e-07 $l=7.05e-07 $layer=LI1_cond $X=9.6 $Y=0.085
+ $X2=9.6 $Y2=0.79
r205 34 109 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.85 $Y=0.085
+ $X2=6.85 $Y2=0
r206 34 36 25.3188 $w=3.28e-07 $l=7.25e-07 $layer=LI1_cond $X=6.85 $Y=0.085
+ $X2=6.85 $Y2=0.81
r207 30 106 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.04 $Y=0.085
+ $X2=5.04 $Y2=0
r208 30 32 20.5135 $w=2.48e-07 $l=4.45e-07 $layer=LI1_cond $X=5.04 $Y=0.085
+ $X2=5.04 $Y2=0.53
r209 26 52 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.365 $Y=0.085
+ $X2=2.365 $Y2=0
r210 26 28 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=2.365 $Y=0.085
+ $X2=2.365 $Y2=0.72
r211 22 103 2.98526 $w=3.3e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.212 $Y2=0
r212 22 24 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.26 $Y2=0.495
r213 7 48 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=12.23
+ $Y=0.37 $X2=12.37 $Y2=0.58
r214 6 44 182 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_NDIFF $count=1 $X=10.88
+ $Y=0.235 $X2=11.02 $Y2=0.43
r215 5 40 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=9.46
+ $Y=0.625 $X2=9.6 $Y2=0.79
r216 4 36 182 $w=1.7e-07 $l=2.59856e-07 $layer=licon1_NDIFF $count=1 $X=6.67
+ $Y=0.625 $X2=6.85 $Y2=0.81
r217 3 32 182 $w=1.7e-07 $l=2.42899e-07 $layer=licon1_NDIFF $count=1 $X=4.88
+ $Y=0.625 $X2=5.08 $Y2=0.53
r218 2 28 182 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=1 $X=2.225
+ $Y=0.545 $X2=2.365 $Y2=0.72
r219 1 24 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.285 $X2=0.26 $Y2=0.495
.ends

