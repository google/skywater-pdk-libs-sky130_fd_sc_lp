* File: sky130_fd_sc_lp__dlrtp_2.pxi.spice
* Created: Fri Aug 28 10:27:11 2020
* 
x_PM_SKY130_FD_SC_LP__DLRTP_2%D N_D_M1011_g N_D_c_153_n N_D_M1017_g N_D_c_155_n
+ D D D D D N_D_c_159_n N_D_c_160_n D PM_SKY130_FD_SC_LP__DLRTP_2%D
x_PM_SKY130_FD_SC_LP__DLRTP_2%GATE N_GATE_M1003_g N_GATE_M1019_g N_GATE_c_199_n
+ N_GATE_c_200_n GATE GATE GATE GATE N_GATE_c_202_n
+ PM_SKY130_FD_SC_LP__DLRTP_2%GATE
x_PM_SKY130_FD_SC_LP__DLRTP_2%A_251_475# N_A_251_475#_M1019_d
+ N_A_251_475#_M1003_d N_A_251_475#_c_264_n N_A_251_475#_M1020_g
+ N_A_251_475#_c_251_n N_A_251_475#_M1021_g N_A_251_475#_M1013_g
+ N_A_251_475#_c_252_n N_A_251_475#_c_253_n N_A_251_475#_M1015_g
+ N_A_251_475#_c_255_n N_A_251_475#_c_275_n N_A_251_475#_c_269_n
+ N_A_251_475#_c_270_n N_A_251_475#_c_292_p N_A_251_475#_c_256_n
+ N_A_251_475#_c_257_n N_A_251_475#_c_258_n N_A_251_475#_c_271_n
+ N_A_251_475#_c_315_p N_A_251_475#_c_259_n N_A_251_475#_c_260_n
+ N_A_251_475#_c_261_n N_A_251_475#_c_262_n N_A_251_475#_c_263_n
+ PM_SKY130_FD_SC_LP__DLRTP_2%A_251_475#
x_PM_SKY130_FD_SC_LP__DLRTP_2%A_40_54# N_A_40_54#_M1011_s N_A_40_54#_M1017_s
+ N_A_40_54#_M1004_g N_A_40_54#_M1010_g N_A_40_54#_c_406_n N_A_40_54#_c_410_n
+ N_A_40_54#_c_421_n N_A_40_54#_c_411_n N_A_40_54#_c_412_n N_A_40_54#_c_413_n
+ N_A_40_54#_c_414_n N_A_40_54#_c_415_n N_A_40_54#_c_416_n
+ PM_SKY130_FD_SC_LP__DLRTP_2%A_40_54#
x_PM_SKY130_FD_SC_LP__DLRTP_2%A_383_479# N_A_383_479#_M1021_s
+ N_A_383_479#_M1020_s N_A_383_479#_M1007_g N_A_383_479#_M1014_g
+ N_A_383_479#_c_496_n N_A_383_479#_c_505_n N_A_383_479#_c_497_n
+ N_A_383_479#_c_498_n N_A_383_479#_c_507_n N_A_383_479#_c_508_n
+ N_A_383_479#_c_584_n N_A_383_479#_c_509_n N_A_383_479#_c_499_n
+ N_A_383_479#_c_500_n N_A_383_479#_c_501_n N_A_383_479#_c_502_n
+ N_A_383_479#_c_503_n N_A_383_479#_c_512_n N_A_383_479#_c_513_n
+ PM_SKY130_FD_SC_LP__DLRTP_2%A_383_479#
x_PM_SKY130_FD_SC_LP__DLRTP_2%A_796_21# N_A_796_21#_M1008_s N_A_796_21#_M1012_d
+ N_A_796_21#_c_630_n N_A_796_21#_M1005_g N_A_796_21#_M1000_g
+ N_A_796_21#_M1006_g N_A_796_21#_M1001_g N_A_796_21#_c_632_n
+ N_A_796_21#_M1016_g N_A_796_21#_M1009_g N_A_796_21#_c_635_n
+ N_A_796_21#_c_636_n N_A_796_21#_c_644_n N_A_796_21#_c_645_n
+ N_A_796_21#_c_637_n N_A_796_21#_c_638_n N_A_796_21#_c_701_p
+ N_A_796_21#_c_647_n N_A_796_21#_c_668_p N_A_796_21#_c_672_p
+ N_A_796_21#_c_639_n N_A_796_21#_c_640_n PM_SKY130_FD_SC_LP__DLRTP_2%A_796_21#
x_PM_SKY130_FD_SC_LP__DLRTP_2%A_646_47# N_A_646_47#_M1007_d N_A_646_47#_M1013_d
+ N_A_646_47#_c_768_n N_A_646_47#_c_769_n N_A_646_47#_c_770_n
+ N_A_646_47#_c_771_n N_A_646_47#_c_772_n N_A_646_47#_M1008_g
+ N_A_646_47#_M1012_g N_A_646_47#_c_786_n N_A_646_47#_c_782_n
+ N_A_646_47#_c_773_n N_A_646_47#_c_793_n N_A_646_47#_c_774_n
+ N_A_646_47#_c_775_n N_A_646_47#_c_776_n N_A_646_47#_c_803_n
+ N_A_646_47#_c_777_n N_A_646_47#_c_778_n N_A_646_47#_c_779_n
+ PM_SKY130_FD_SC_LP__DLRTP_2%A_646_47#
x_PM_SKY130_FD_SC_LP__DLRTP_2%RESET_B N_RESET_B_M1002_g N_RESET_B_M1018_g
+ RESET_B RESET_B N_RESET_B_c_888_n N_RESET_B_c_889_n
+ PM_SKY130_FD_SC_LP__DLRTP_2%RESET_B
x_PM_SKY130_FD_SC_LP__DLRTP_2%VPWR N_VPWR_M1017_d N_VPWR_M1020_d N_VPWR_M1000_d
+ N_VPWR_M1018_d N_VPWR_M1009_d N_VPWR_c_926_n N_VPWR_c_927_n N_VPWR_c_928_n
+ N_VPWR_c_929_n N_VPWR_c_930_n N_VPWR_c_931_n N_VPWR_c_932_n N_VPWR_c_933_n
+ N_VPWR_c_934_n VPWR N_VPWR_c_935_n N_VPWR_c_936_n N_VPWR_c_937_n
+ N_VPWR_c_938_n N_VPWR_c_939_n N_VPWR_c_925_n PM_SKY130_FD_SC_LP__DLRTP_2%VPWR
x_PM_SKY130_FD_SC_LP__DLRTP_2%Q N_Q_M1006_d N_Q_M1001_s Q Q Q Q Q Q Q
+ N_Q_c_1024_n Q PM_SKY130_FD_SC_LP__DLRTP_2%Q
x_PM_SKY130_FD_SC_LP__DLRTP_2%VGND N_VGND_M1011_d N_VGND_M1021_d N_VGND_M1005_d
+ N_VGND_M1002_d N_VGND_M1016_s N_VGND_c_1046_n N_VGND_c_1047_n N_VGND_c_1048_n
+ N_VGND_c_1049_n N_VGND_c_1050_n N_VGND_c_1051_n N_VGND_c_1052_n
+ N_VGND_c_1053_n N_VGND_c_1054_n N_VGND_c_1055_n N_VGND_c_1056_n
+ N_VGND_c_1057_n VGND N_VGND_c_1058_n N_VGND_c_1059_n N_VGND_c_1060_n
+ N_VGND_c_1061_n PM_SKY130_FD_SC_LP__DLRTP_2%VGND
cc_1 VNB N_D_c_153_n 0.0215595f $X=-0.19 $Y=-0.245 $X2=0.652 $Y2=1.283
cc_2 VNB N_D_M1017_g 0.0104674f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=2.695
cc_3 VNB N_D_c_155_n 0.0201353f $X=-0.19 $Y=-0.245 $X2=0.652 $Y2=1.47
cc_4 VNB D 0.00127546f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.47
cc_5 VNB D 0.00170307f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.84
cc_6 VNB D 0.00421821f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_7 VNB N_D_c_159_n 0.0209671f $X=-0.19 $Y=-0.245 $X2=0.675 $Y2=0.965
cc_8 VNB N_D_c_160_n 0.021535f $X=-0.19 $Y=-0.245 $X2=0.652 $Y2=0.8
cc_9 VNB N_GATE_M1003_g 0.00766035f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=0.48
cc_10 VNB N_GATE_M1019_g 0.0240574f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=2.695
cc_11 VNB N_GATE_c_199_n 0.0237671f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.47
cc_12 VNB N_GATE_c_200_n 0.019187f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.84
cc_13 VNB GATE 0.00415422f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_14 VNB N_GATE_c_202_n 0.016847f $X=-0.19 $Y=-0.245 $X2=0.652 $Y2=0.965
cc_15 VNB N_A_251_475#_c_251_n 0.0197337f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.95
cc_16 VNB N_A_251_475#_c_252_n 0.015652f $X=-0.19 $Y=-0.245 $X2=0.652 $Y2=0.965
cc_17 VNB N_A_251_475#_c_253_n 0.00818056f $X=-0.19 $Y=-0.245 $X2=0.675
+ $Y2=0.965
cc_18 VNB N_A_251_475#_M1015_g 0.0347615f $X=-0.19 $Y=-0.245 $X2=0.692 $Y2=0.815
cc_19 VNB N_A_251_475#_c_255_n 0.0171948f $X=-0.19 $Y=-0.245 $X2=0.73 $Y2=0.965
cc_20 VNB N_A_251_475#_c_256_n 0.018674f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_251_475#_c_257_n 0.00223322f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_251_475#_c_258_n 0.0023489f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_251_475#_c_259_n 0.006828f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_251_475#_c_260_n 0.00482395f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_251_475#_c_261_n 0.0152321f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_251_475#_c_262_n 0.00968195f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_251_475#_c_263_n 0.120523f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_40_54#_M1004_g 0.0628642f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_40_54#_c_406_n 0.0633081f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_383_479#_M1007_g 0.0264823f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_383_479#_c_496_n 0.00746136f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_383_479#_c_497_n 0.00957103f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_383_479#_c_498_n 0.0050803f $X=-0.19 $Y=-0.245 $X2=0.675 $Y2=0.965
cc_34 VNB N_A_383_479#_c_499_n 0.00592012f $X=-0.19 $Y=-0.245 $X2=0.73 $Y2=1.665
cc_35 VNB N_A_383_479#_c_500_n 0.00252669f $X=-0.19 $Y=-0.245 $X2=0.73 $Y2=2.035
cc_36 VNB N_A_383_479#_c_501_n 0.00480244f $X=-0.19 $Y=-0.245 $X2=0.73 $Y2=0.815
cc_37 VNB N_A_383_479#_c_502_n 0.0333532f $X=-0.19 $Y=-0.245 $X2=0.73 $Y2=0.925
cc_38 VNB N_A_383_479#_c_503_n 0.00137822f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_796_21#_c_630_n 0.0164009f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=2.695
cc_40 VNB N_A_796_21#_M1006_g 0.0210063f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_796_21#_c_632_n 0.00705027f $X=-0.19 $Y=-0.245 $X2=0.675 $Y2=0.965
cc_42 VNB N_A_796_21#_M1016_g 0.0234029f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_796_21#_M1009_g 0.0127452f $X=-0.19 $Y=-0.245 $X2=0.73 $Y2=1.295
cc_44 VNB N_A_796_21#_c_635_n 0.0207553f $X=-0.19 $Y=-0.245 $X2=0.73 $Y2=2.035
cc_45 VNB N_A_796_21#_c_636_n 0.0180684f $X=-0.19 $Y=-0.245 $X2=0.73 $Y2=0.902
cc_46 VNB N_A_796_21#_c_637_n 0.00181497f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_796_21#_c_638_n 0.00372875f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_796_21#_c_639_n 0.0369087f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_796_21#_c_640_n 0.0239019f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_646_47#_c_768_n 0.0573702f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=2.695
cc_51 VNB N_A_646_47#_c_769_n 0.0324675f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_646_47#_c_770_n 0.0104628f $X=-0.19 $Y=-0.245 $X2=0.652 $Y2=1.47
cc_53 VNB N_A_646_47#_c_771_n 0.0136248f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.47
cc_54 VNB N_A_646_47#_c_772_n 0.0136423f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_55 VNB N_A_646_47#_c_773_n 0.00512737f $X=-0.19 $Y=-0.245 $X2=0.692 $Y2=0.815
cc_56 VNB N_A_646_47#_c_774_n 5.86216e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_646_47#_c_775_n 0.00753037f $X=-0.19 $Y=-0.245 $X2=0.73 $Y2=0.965
cc_58 VNB N_A_646_47#_c_776_n 0.00158194f $X=-0.19 $Y=-0.245 $X2=0.73 $Y2=0.965
cc_59 VNB N_A_646_47#_c_777_n 0.00425435f $X=-0.19 $Y=-0.245 $X2=0.73 $Y2=0.815
cc_60 VNB N_A_646_47#_c_778_n 0.026086f $X=-0.19 $Y=-0.245 $X2=0.73 $Y2=0.925
cc_61 VNB N_A_646_47#_c_779_n 0.00403922f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=0.925
cc_62 VNB N_RESET_B_M1018_g 3.97806e-19 $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=1.47
cc_63 VNB RESET_B 0.00910814f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=2.695
cc_64 VNB N_RESET_B_c_888_n 0.0326652f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_65 VNB N_RESET_B_c_889_n 0.0169003f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.95
cc_66 VNB N_VPWR_c_925_n 0.302998f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB Q 0.00385282f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_Q_c_1024_n 0.00321484f $X=-0.19 $Y=-0.245 $X2=0.675 $Y2=0.965
cc_69 VNB N_VGND_c_1046_n 0.0059352f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_VGND_c_1047_n 0.00250426f $X=-0.19 $Y=-0.245 $X2=0.652 $Y2=0.965
cc_71 VNB N_VGND_c_1048_n 0.00486219f $X=-0.19 $Y=-0.245 $X2=0.692 $Y2=0.815
cc_72 VNB N_VGND_c_1049_n 0.00971861f $X=-0.19 $Y=-0.245 $X2=0.73 $Y2=0.965
cc_73 VNB N_VGND_c_1050_n 0.0138678f $X=-0.19 $Y=-0.245 $X2=0.73 $Y2=1.295
cc_74 VNB N_VGND_c_1051_n 0.0479511f $X=-0.19 $Y=-0.245 $X2=0.73 $Y2=1.665
cc_75 VNB N_VGND_c_1052_n 0.0292292f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_VGND_c_1053_n 0.00384695f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_VGND_c_1054_n 0.0371766f $X=-0.19 $Y=-0.245 $X2=0.73 $Y2=0.815
cc_78 VNB N_VGND_c_1055_n 0.00381613f $X=-0.19 $Y=-0.245 $X2=0.73 $Y2=0.925
cc_79 VNB N_VGND_c_1056_n 0.0326753f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_VGND_c_1057_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_VGND_c_1058_n 0.0339529f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_VGND_c_1059_n 0.0222148f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_VGND_c_1060_n 0.00414071f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_VGND_c_1061_n 0.393918f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VPB N_D_M1017_g 0.0573947f $X=-0.19 $Y=1.655 $X2=0.54 $Y2=2.695
cc_86 VPB D 0.00712354f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_87 VPB N_GATE_M1003_g 0.0533468f $X=-0.19 $Y=1.655 $X2=0.54 $Y2=0.48
cc_88 VPB GATE 0.00860337f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_89 VPB N_A_251_475#_c_264_n 0.0348637f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_90 VPB N_A_251_475#_M1020_g 0.0252948f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_91 VPB N_A_251_475#_M1013_g 0.0526884f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_92 VPB N_A_251_475#_c_252_n 0.0103603f $X=-0.19 $Y=1.655 $X2=0.652 $Y2=0.965
cc_93 VPB N_A_251_475#_c_253_n 3.95601e-19 $X=-0.19 $Y=1.655 $X2=0.675 $Y2=0.965
cc_94 VPB N_A_251_475#_c_269_n 0.00310603f $X=-0.19 $Y=1.655 $X2=0.73 $Y2=2.035
cc_95 VPB N_A_251_475#_c_270_n 0.0347641f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_96 VPB N_A_251_475#_c_271_n 0.00993705f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_97 VPB N_A_251_475#_c_259_n 0.00143775f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_98 VPB N_A_251_475#_c_262_n 0.0125084f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_99 VPB N_A_40_54#_M1004_g 0.0159961f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_100 VPB N_A_40_54#_M1010_g 0.0211695f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_101 VPB N_A_40_54#_c_406_n 0.035558f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_102 VPB N_A_40_54#_c_410_n 0.0106282f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_103 VPB N_A_40_54#_c_411_n 0.0141936f $X=-0.19 $Y=1.655 $X2=0.652 $Y2=0.8
cc_104 VPB N_A_40_54#_c_412_n 9.19968e-19 $X=-0.19 $Y=1.655 $X2=0.692 $Y2=0.815
cc_105 VPB N_A_40_54#_c_413_n 0.00220368f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_106 VPB N_A_40_54#_c_414_n 0.0291297f $X=-0.19 $Y=1.655 $X2=0.73 $Y2=0.965
cc_107 VPB N_A_40_54#_c_415_n 0.00608141f $X=-0.19 $Y=1.655 $X2=0.73 $Y2=1.665
cc_108 VPB N_A_40_54#_c_416_n 0.0501766f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_109 VPB N_A_383_479#_M1014_g 0.0177929f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_110 VPB N_A_383_479#_c_505_n 0.0132903f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_111 VPB N_A_383_479#_c_497_n 0.00745922f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_112 VPB N_A_383_479#_c_507_n 0.00779991f $X=-0.19 $Y=1.655 $X2=0.692
+ $Y2=0.815
cc_113 VPB N_A_383_479#_c_508_n 0.00562272f $X=-0.19 $Y=1.655 $X2=0.692
+ $Y2=0.555
cc_114 VPB N_A_383_479#_c_509_n 0.00185535f $X=-0.19 $Y=1.655 $X2=0.73 $Y2=0.965
cc_115 VPB N_A_383_479#_c_500_n 0.00172823f $X=-0.19 $Y=1.655 $X2=0.73 $Y2=2.035
cc_116 VPB N_A_383_479#_c_503_n 5.34002e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_117 VPB N_A_383_479#_c_512_n 0.0312621f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_118 VPB N_A_383_479#_c_513_n 0.00334948f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_119 VPB N_A_796_21#_M1000_g 0.0225096f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_120 VPB N_A_796_21#_M1001_g 0.0203932f $X=-0.19 $Y=1.655 $X2=0.652 $Y2=0.965
cc_121 VPB N_A_796_21#_M1009_g 0.0264146f $X=-0.19 $Y=1.655 $X2=0.73 $Y2=1.295
cc_122 VPB N_A_796_21#_c_644_n 0.00657483f $X=-0.19 $Y=1.655 $X2=0.73 $Y2=0.925
cc_123 VPB N_A_796_21#_c_645_n 0.0332677f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_124 VPB N_A_796_21#_c_638_n 0.00181623f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_125 VPB N_A_796_21#_c_647_n 0.00153823f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_126 VPB N_A_796_21#_c_639_n 0.0183162f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_127 VPB N_A_796_21#_c_640_n 0.00795167f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_128 VPB N_A_646_47#_c_771_n 0.00765856f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=0.47
cc_129 VPB N_A_646_47#_M1012_g 0.02214f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_130 VPB N_A_646_47#_c_782_n 0.00585683f $X=-0.19 $Y=1.655 $X2=0.652 $Y2=0.8
cc_131 VPB N_A_646_47#_c_773_n 0.0111397f $X=-0.19 $Y=1.655 $X2=0.692 $Y2=0.815
cc_132 VPB N_A_646_47#_c_777_n 0.00312354f $X=-0.19 $Y=1.655 $X2=0.73 $Y2=0.815
cc_133 VPB N_A_646_47#_c_778_n 0.0105811f $X=-0.19 $Y=1.655 $X2=0.73 $Y2=0.925
cc_134 VPB N_RESET_B_M1018_g 0.0217307f $X=-0.19 $Y=1.655 $X2=0.54 $Y2=1.47
cc_135 VPB RESET_B 0.00308692f $X=-0.19 $Y=1.655 $X2=0.54 $Y2=2.695
cc_136 VPB N_VPWR_c_926_n 0.00434557f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_137 VPB N_VPWR_c_927_n 0.00755713f $X=-0.19 $Y=1.655 $X2=0.652 $Y2=0.965
cc_138 VPB N_VPWR_c_928_n 0.00509424f $X=-0.19 $Y=1.655 $X2=0.692 $Y2=0.815
cc_139 VPB N_VPWR_c_929_n 0.0114299f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_140 VPB N_VPWR_c_930_n 0.0594562f $X=-0.19 $Y=1.655 $X2=0.73 $Y2=0.965
cc_141 VPB N_VPWR_c_931_n 0.043913f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_142 VPB N_VPWR_c_932_n 0.00362871f $X=-0.19 $Y=1.655 $X2=0.73 $Y2=2.035
cc_143 VPB N_VPWR_c_933_n 0.0198787f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_144 VPB N_VPWR_c_934_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0.73 $Y2=0.902
cc_145 VPB N_VPWR_c_935_n 0.0184299f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=0.925
cc_146 VPB N_VPWR_c_936_n 0.0376809f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_147 VPB N_VPWR_c_937_n 0.0180584f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_148 VPB N_VPWR_c_938_n 0.00420726f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_149 VPB N_VPWR_c_939_n 0.029932f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_150 VPB N_VPWR_c_925_n 0.0844581f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_151 VPB Q 0.00356419f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_152 N_D_M1017_g N_GATE_M1003_g 0.0306399f $X=0.54 $Y=2.695 $X2=0 $Y2=0
cc_153 D N_GATE_M1003_g 0.00215018f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_154 D N_GATE_M1019_g 0.0018297f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_155 N_D_c_159_n N_GATE_M1019_g 0.00119515f $X=0.675 $Y=0.965 $X2=0 $Y2=0
cc_156 N_D_c_160_n N_GATE_M1019_g 0.00668735f $X=0.652 $Y=0.8 $X2=0 $Y2=0
cc_157 N_D_c_153_n N_GATE_c_199_n 0.0130946f $X=0.652 $Y=1.283 $X2=0 $Y2=0
cc_158 D N_GATE_c_199_n 0.00192047f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_159 N_D_M1017_g N_GATE_c_200_n 8.9634e-19 $X=0.54 $Y=2.695 $X2=0 $Y2=0
cc_160 N_D_c_155_n N_GATE_c_200_n 0.0130946f $X=0.652 $Y=1.47 $X2=0 $Y2=0
cc_161 N_D_M1017_g GATE 0.00134579f $X=0.54 $Y=2.695 $X2=0 $Y2=0
cc_162 D GATE 0.102865f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_163 N_D_c_159_n GATE 8.09896e-19 $X=0.675 $Y=0.965 $X2=0 $Y2=0
cc_164 D N_GATE_c_202_n 0.00192047f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_165 N_D_c_159_n N_GATE_c_202_n 0.0130946f $X=0.675 $Y=0.965 $X2=0 $Y2=0
cc_166 D N_A_251_475#_c_259_n 0.00432527f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_167 D N_A_40_54#_c_406_n 0.122737f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_168 N_D_c_160_n N_A_40_54#_c_406_n 0.044445f $X=0.652 $Y=0.8 $X2=0 $Y2=0
cc_169 N_D_M1017_g N_A_40_54#_c_410_n 0.0145484f $X=0.54 $Y=2.695 $X2=0 $Y2=0
cc_170 D N_A_40_54#_c_410_n 0.0197623f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_171 N_D_M1017_g N_A_40_54#_c_421_n 0.0012521f $X=0.54 $Y=2.695 $X2=0 $Y2=0
cc_172 N_D_M1017_g N_A_40_54#_c_412_n 3.62397e-19 $X=0.54 $Y=2.695 $X2=0 $Y2=0
cc_173 N_D_M1017_g N_A_40_54#_c_414_n 2.2485e-19 $X=0.54 $Y=2.695 $X2=0 $Y2=0
cc_174 N_D_M1017_g N_VPWR_c_926_n 0.00918319f $X=0.54 $Y=2.695 $X2=0 $Y2=0
cc_175 N_D_M1017_g N_VPWR_c_935_n 0.00456036f $X=0.54 $Y=2.695 $X2=0 $Y2=0
cc_176 N_D_M1017_g N_VPWR_c_925_n 0.00490792f $X=0.54 $Y=2.695 $X2=0 $Y2=0
cc_177 D N_VGND_M1011_d 0.00542875f $X=0.635 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_178 D N_VGND_c_1046_n 0.0247787f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_179 N_D_c_160_n N_VGND_c_1046_n 0.00358365f $X=0.652 $Y=0.8 $X2=0 $Y2=0
cc_180 D N_VGND_c_1052_n 0.00983876f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_181 N_D_c_160_n N_VGND_c_1052_n 0.00504079f $X=0.652 $Y=0.8 $X2=0 $Y2=0
cc_182 D N_VGND_c_1061_n 0.00824407f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_183 D N_VGND_c_1061_n 0.00284498f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_184 N_D_c_159_n N_VGND_c_1061_n 9.31712e-19 $X=0.675 $Y=0.965 $X2=0 $Y2=0
cc_185 N_D_c_160_n N_VGND_c_1061_n 0.0106406f $X=0.652 $Y=0.8 $X2=0 $Y2=0
cc_186 N_GATE_M1003_g N_A_251_475#_c_275_n 2.65919e-19 $X=1.18 $Y=2.695 $X2=0
+ $Y2=0
cc_187 N_GATE_M1003_g N_A_251_475#_c_269_n 0.00530813f $X=1.18 $Y=2.695 $X2=0
+ $Y2=0
cc_188 N_GATE_M1003_g N_A_251_475#_c_270_n 0.0217176f $X=1.18 $Y=2.695 $X2=0
+ $Y2=0
cc_189 GATE N_A_251_475#_c_270_n 0.00141857f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_190 N_GATE_M1003_g N_A_251_475#_c_271_n 0.00140139f $X=1.18 $Y=2.695 $X2=0
+ $Y2=0
cc_191 N_GATE_M1003_g N_A_251_475#_c_259_n 0.001172f $X=1.18 $Y=2.695 $X2=0
+ $Y2=0
cc_192 N_GATE_M1019_g N_A_251_475#_c_259_n 0.00292299f $X=1.295 $Y=0.48 $X2=0
+ $Y2=0
cc_193 GATE N_A_251_475#_c_259_n 0.0937519f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_194 N_GATE_c_202_n N_A_251_475#_c_259_n 0.00470804f $X=1.215 $Y=1.005 $X2=0
+ $Y2=0
cc_195 N_GATE_M1003_g N_A_251_475#_c_262_n 0.0107459f $X=1.18 $Y=2.695 $X2=0
+ $Y2=0
cc_196 N_GATE_c_199_n N_A_251_475#_c_262_n 0.0153786f $X=1.215 $Y=1.345 $X2=0
+ $Y2=0
cc_197 GATE N_A_251_475#_c_262_n 9.48102e-19 $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_198 N_GATE_M1019_g N_A_251_475#_c_263_n 0.00309855f $X=1.295 $Y=0.48 $X2=0
+ $Y2=0
cc_199 GATE N_A_251_475#_c_263_n 5.87087e-19 $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_200 N_GATE_c_202_n N_A_251_475#_c_263_n 0.0153786f $X=1.215 $Y=1.005 $X2=0
+ $Y2=0
cc_201 N_GATE_M1003_g N_A_40_54#_c_410_n 0.00691878f $X=1.18 $Y=2.695 $X2=0
+ $Y2=0
cc_202 GATE N_A_40_54#_c_410_n 0.00958738f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_203 N_GATE_M1003_g N_A_40_54#_c_421_n 0.0139095f $X=1.18 $Y=2.695 $X2=0 $Y2=0
cc_204 N_GATE_M1003_g N_A_40_54#_c_411_n 0.00837729f $X=1.18 $Y=2.695 $X2=0
+ $Y2=0
cc_205 N_GATE_M1003_g N_A_40_54#_c_412_n 0.0036468f $X=1.18 $Y=2.695 $X2=0 $Y2=0
cc_206 N_GATE_M1003_g N_A_383_479#_c_505_n 5.54363e-19 $X=1.18 $Y=2.695 $X2=0
+ $Y2=0
cc_207 N_GATE_M1019_g N_A_383_479#_c_499_n 0.00128819f $X=1.295 $Y=0.48 $X2=0
+ $Y2=0
cc_208 N_GATE_M1003_g N_VPWR_c_926_n 0.00275423f $X=1.18 $Y=2.695 $X2=0 $Y2=0
cc_209 N_GATE_M1003_g N_VPWR_c_931_n 0.00311439f $X=1.18 $Y=2.695 $X2=0 $Y2=0
cc_210 N_GATE_M1003_g N_VPWR_c_925_n 0.00533795f $X=1.18 $Y=2.695 $X2=0 $Y2=0
cc_211 N_GATE_M1019_g N_VGND_c_1046_n 0.00322794f $X=1.295 $Y=0.48 $X2=0 $Y2=0
cc_212 GATE N_VGND_c_1046_n 0.0105057f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_213 N_GATE_c_202_n N_VGND_c_1046_n 8.66294e-19 $X=1.215 $Y=1.005 $X2=0 $Y2=0
cc_214 N_GATE_M1019_g N_VGND_c_1058_n 0.00550375f $X=1.295 $Y=0.48 $X2=0 $Y2=0
cc_215 N_GATE_M1019_g N_VGND_c_1061_n 0.00962223f $X=1.295 $Y=0.48 $X2=0 $Y2=0
cc_216 GATE N_VGND_c_1061_n 0.00489131f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_217 N_GATE_c_202_n N_VGND_c_1061_n 2.5288e-19 $X=1.215 $Y=1.005 $X2=0 $Y2=0
cc_218 N_A_251_475#_c_251_n N_A_40_54#_M1004_g 0.0159908f $X=2.365 $Y=0.765
+ $X2=0 $Y2=0
cc_219 N_A_251_475#_c_253_n N_A_40_54#_M1004_g 0.00655854f $X=3.415 $Y=1.59
+ $X2=0 $Y2=0
cc_220 N_A_251_475#_c_292_p N_A_40_54#_M1004_g 0.00232573f $X=2.345 $Y=0.93
+ $X2=0 $Y2=0
cc_221 N_A_251_475#_c_256_n N_A_40_54#_M1004_g 0.0132675f $X=3.59 $Y=0.79 $X2=0
+ $Y2=0
cc_222 N_A_251_475#_c_263_n N_A_40_54#_M1004_g 0.0445622f $X=2.365 $Y=1.1 $X2=0
+ $Y2=0
cc_223 N_A_251_475#_M1020_g N_A_40_54#_M1010_g 0.00947684f $X=2.255 $Y=2.715
+ $X2=0 $Y2=0
cc_224 N_A_251_475#_c_271_n N_A_40_54#_c_410_n 0.0141001f $X=1.597 $Y=2.535
+ $X2=0 $Y2=0
cc_225 N_A_251_475#_c_271_n N_A_40_54#_c_421_n 0.0141042f $X=1.597 $Y=2.535
+ $X2=0 $Y2=0
cc_226 N_A_251_475#_M1003_d N_A_40_54#_c_411_n 0.00512462f $X=1.255 $Y=2.375
+ $X2=0 $Y2=0
cc_227 N_A_251_475#_c_264_n N_A_40_54#_c_411_n 6.49098e-19 $X=2.18 $Y=2.14 $X2=0
+ $Y2=0
cc_228 N_A_251_475#_M1020_g N_A_40_54#_c_411_n 0.0152235f $X=2.255 $Y=2.715
+ $X2=0 $Y2=0
cc_229 N_A_251_475#_c_270_n N_A_40_54#_c_411_n 0.00384991f $X=1.63 $Y=2.05 $X2=0
+ $Y2=0
cc_230 N_A_251_475#_c_271_n N_A_40_54#_c_411_n 0.0260862f $X=1.597 $Y=2.535
+ $X2=0 $Y2=0
cc_231 N_A_251_475#_M1020_g N_A_40_54#_c_413_n 0.0203403f $X=2.255 $Y=2.715
+ $X2=0 $Y2=0
cc_232 N_A_251_475#_c_264_n N_A_40_54#_c_415_n 0.00422387f $X=2.18 $Y=2.14 $X2=0
+ $Y2=0
cc_233 N_A_251_475#_M1020_g N_A_40_54#_c_415_n 2.14805e-19 $X=2.255 $Y=2.715
+ $X2=0 $Y2=0
cc_234 N_A_251_475#_c_264_n N_A_40_54#_c_416_n 0.0104165f $X=2.18 $Y=2.14 $X2=0
+ $Y2=0
cc_235 N_A_251_475#_M1013_g N_A_40_54#_c_416_n 0.0724072f $X=3.34 $Y=2.715 $X2=0
+ $Y2=0
cc_236 N_A_251_475#_M1015_g N_A_383_479#_M1007_g 0.0203292f $X=3.695 $Y=0.445
+ $X2=0 $Y2=0
cc_237 N_A_251_475#_c_256_n N_A_383_479#_M1007_g 0.0121786f $X=3.59 $Y=0.79
+ $X2=0 $Y2=0
cc_238 N_A_251_475#_c_258_n N_A_383_479#_M1007_g 0.00171438f $X=3.675 $Y=1.125
+ $X2=0 $Y2=0
cc_239 N_A_251_475#_M1013_g N_A_383_479#_M1014_g 0.0157481f $X=3.34 $Y=2.715
+ $X2=0 $Y2=0
cc_240 N_A_251_475#_c_251_n N_A_383_479#_c_496_n 0.00436289f $X=2.365 $Y=0.765
+ $X2=0 $Y2=0
cc_241 N_A_251_475#_c_292_p N_A_383_479#_c_496_n 0.0352413f $X=2.345 $Y=0.93
+ $X2=0 $Y2=0
cc_242 N_A_251_475#_c_257_n N_A_383_479#_c_496_n 0.0135498f $X=2.51 $Y=0.79
+ $X2=0 $Y2=0
cc_243 N_A_251_475#_c_315_p N_A_383_479#_c_496_n 0.0703689f $X=1.53 $Y=0.495
+ $X2=0 $Y2=0
cc_244 N_A_251_475#_c_262_n N_A_383_479#_c_496_n 2.25352e-19 $X=1.63 $Y=1.885
+ $X2=0 $Y2=0
cc_245 N_A_251_475#_c_263_n N_A_383_479#_c_496_n 0.0388362f $X=2.365 $Y=1.1
+ $X2=0 $Y2=0
cc_246 N_A_251_475#_c_264_n N_A_383_479#_c_505_n 0.0179137f $X=2.18 $Y=2.14
+ $X2=0 $Y2=0
cc_247 N_A_251_475#_M1020_g N_A_383_479#_c_505_n 0.00404045f $X=2.255 $Y=2.715
+ $X2=0 $Y2=0
cc_248 N_A_251_475#_c_275_n N_A_383_479#_c_505_n 0.0354218f $X=1.597 $Y=2.002
+ $X2=0 $Y2=0
cc_249 N_A_251_475#_c_271_n N_A_383_479#_c_505_n 0.0294977f $X=1.597 $Y=2.535
+ $X2=0 $Y2=0
cc_250 N_A_251_475#_c_259_n N_A_383_479#_c_505_n 0.010376f $X=1.597 $Y=1.885
+ $X2=0 $Y2=0
cc_251 N_A_251_475#_c_262_n N_A_383_479#_c_505_n 0.00621683f $X=1.63 $Y=1.885
+ $X2=0 $Y2=0
cc_252 N_A_251_475#_c_264_n N_A_383_479#_c_497_n 0.0035126f $X=2.18 $Y=2.14
+ $X2=0 $Y2=0
cc_253 N_A_251_475#_c_292_p N_A_383_479#_c_497_n 0.0261476f $X=2.345 $Y=0.93
+ $X2=0 $Y2=0
cc_254 N_A_251_475#_c_256_n N_A_383_479#_c_497_n 0.0133271f $X=3.59 $Y=0.79
+ $X2=0 $Y2=0
cc_255 N_A_251_475#_c_263_n N_A_383_479#_c_497_n 0.00842007f $X=2.365 $Y=1.1
+ $X2=0 $Y2=0
cc_256 N_A_251_475#_c_253_n N_A_383_479#_c_498_n 5.08546e-19 $X=3.415 $Y=1.59
+ $X2=0 $Y2=0
cc_257 N_A_251_475#_c_255_n N_A_383_479#_c_498_n 0.00409938f $X=3.785 $Y=1.515
+ $X2=0 $Y2=0
cc_258 N_A_251_475#_c_292_p N_A_383_479#_c_498_n 0.00201073f $X=2.345 $Y=0.93
+ $X2=0 $Y2=0
cc_259 N_A_251_475#_c_260_n N_A_383_479#_c_498_n 0.00341087f $X=3.785 $Y=1.29
+ $X2=0 $Y2=0
cc_260 N_A_251_475#_M1020_g N_A_383_479#_c_507_n 2.14464e-19 $X=2.255 $Y=2.715
+ $X2=0 $Y2=0
cc_261 N_A_251_475#_M1013_g N_A_383_479#_c_507_n 0.0100263f $X=3.34 $Y=2.715
+ $X2=0 $Y2=0
cc_262 N_A_251_475#_M1013_g N_A_383_479#_c_508_n 0.0131521f $X=3.34 $Y=2.715
+ $X2=0 $Y2=0
cc_263 N_A_251_475#_M1013_g N_A_383_479#_c_509_n 7.73147e-19 $X=3.34 $Y=2.715
+ $X2=0 $Y2=0
cc_264 N_A_251_475#_c_251_n N_A_383_479#_c_499_n 0.00243824f $X=2.365 $Y=0.765
+ $X2=0 $Y2=0
cc_265 N_A_251_475#_c_257_n N_A_383_479#_c_499_n 0.00711944f $X=2.51 $Y=0.79
+ $X2=0 $Y2=0
cc_266 N_A_251_475#_c_315_p N_A_383_479#_c_499_n 0.0167775f $X=1.53 $Y=0.495
+ $X2=0 $Y2=0
cc_267 N_A_251_475#_c_263_n N_A_383_479#_c_499_n 0.00823307f $X=2.365 $Y=1.1
+ $X2=0 $Y2=0
cc_268 N_A_251_475#_c_264_n N_A_383_479#_c_500_n 0.00159207f $X=2.18 $Y=2.14
+ $X2=0 $Y2=0
cc_269 N_A_251_475#_c_259_n N_A_383_479#_c_500_n 0.0137139f $X=1.597 $Y=1.885
+ $X2=0 $Y2=0
cc_270 N_A_251_475#_c_262_n N_A_383_479#_c_500_n 0.00406933f $X=1.63 $Y=1.885
+ $X2=0 $Y2=0
cc_271 N_A_251_475#_c_263_n N_A_383_479#_c_500_n 0.00458831f $X=2.365 $Y=1.1
+ $X2=0 $Y2=0
cc_272 N_A_251_475#_c_253_n N_A_383_479#_c_501_n 9.22588e-19 $X=3.415 $Y=1.59
+ $X2=0 $Y2=0
cc_273 N_A_251_475#_c_292_p N_A_383_479#_c_501_n 0.00931143f $X=2.345 $Y=0.93
+ $X2=0 $Y2=0
cc_274 N_A_251_475#_c_256_n N_A_383_479#_c_501_n 0.0296304f $X=3.59 $Y=0.79
+ $X2=0 $Y2=0
cc_275 N_A_251_475#_c_258_n N_A_383_479#_c_501_n 0.00580372f $X=3.675 $Y=1.125
+ $X2=0 $Y2=0
cc_276 N_A_251_475#_c_260_n N_A_383_479#_c_501_n 0.0139194f $X=3.785 $Y=1.29
+ $X2=0 $Y2=0
cc_277 N_A_251_475#_c_261_n N_A_383_479#_c_501_n 2.09038e-19 $X=3.785 $Y=1.29
+ $X2=0 $Y2=0
cc_278 N_A_251_475#_c_253_n N_A_383_479#_c_502_n 0.0100145f $X=3.415 $Y=1.59
+ $X2=0 $Y2=0
cc_279 N_A_251_475#_M1015_g N_A_383_479#_c_502_n 0.0211563f $X=3.695 $Y=0.445
+ $X2=0 $Y2=0
cc_280 N_A_251_475#_c_256_n N_A_383_479#_c_502_n 0.00438376f $X=3.59 $Y=0.79
+ $X2=0 $Y2=0
cc_281 N_A_251_475#_c_258_n N_A_383_479#_c_502_n 0.00166654f $X=3.675 $Y=1.125
+ $X2=0 $Y2=0
cc_282 N_A_251_475#_c_260_n N_A_383_479#_c_502_n 6.03139e-19 $X=3.785 $Y=1.29
+ $X2=0 $Y2=0
cc_283 N_A_251_475#_c_253_n N_A_383_479#_c_503_n 0.00226943f $X=3.415 $Y=1.59
+ $X2=0 $Y2=0
cc_284 N_A_251_475#_M1013_g N_A_383_479#_c_512_n 0.0203599f $X=3.34 $Y=2.715
+ $X2=0 $Y2=0
cc_285 N_A_251_475#_c_252_n N_A_383_479#_c_512_n 0.0176854f $X=3.62 $Y=1.59
+ $X2=0 $Y2=0
cc_286 N_A_251_475#_M1013_g N_A_383_479#_c_513_n 2.96597e-19 $X=3.34 $Y=2.715
+ $X2=0 $Y2=0
cc_287 N_A_251_475#_c_252_n N_A_383_479#_c_513_n 2.75229e-19 $X=3.62 $Y=1.59
+ $X2=0 $Y2=0
cc_288 N_A_251_475#_M1015_g N_A_796_21#_c_630_n 0.0508001f $X=3.695 $Y=0.445
+ $X2=0 $Y2=0
cc_289 N_A_251_475#_M1015_g N_A_796_21#_c_639_n 0.00651496f $X=3.695 $Y=0.445
+ $X2=0 $Y2=0
cc_290 N_A_251_475#_c_258_n N_A_796_21#_c_639_n 0.001192f $X=3.675 $Y=1.125
+ $X2=0 $Y2=0
cc_291 N_A_251_475#_c_260_n N_A_796_21#_c_639_n 9.7532e-19 $X=3.785 $Y=1.29
+ $X2=0 $Y2=0
cc_292 N_A_251_475#_c_261_n N_A_796_21#_c_639_n 0.0331542f $X=3.785 $Y=1.29
+ $X2=0 $Y2=0
cc_293 N_A_251_475#_M1015_g N_A_646_47#_c_786_n 0.00988926f $X=3.695 $Y=0.445
+ $X2=0 $Y2=0
cc_294 N_A_251_475#_c_256_n N_A_646_47#_c_786_n 0.0305295f $X=3.59 $Y=0.79 $X2=0
+ $Y2=0
cc_295 N_A_251_475#_c_260_n N_A_646_47#_c_786_n 0.00397417f $X=3.785 $Y=1.29
+ $X2=0 $Y2=0
cc_296 N_A_251_475#_c_261_n N_A_646_47#_c_786_n 0.00282605f $X=3.785 $Y=1.29
+ $X2=0 $Y2=0
cc_297 N_A_251_475#_M1013_g N_A_646_47#_c_782_n 0.0146263f $X=3.34 $Y=2.715
+ $X2=0 $Y2=0
cc_298 N_A_251_475#_c_252_n N_A_646_47#_c_773_n 0.0151802f $X=3.62 $Y=1.59 $X2=0
+ $Y2=0
cc_299 N_A_251_475#_c_260_n N_A_646_47#_c_773_n 0.0253089f $X=3.785 $Y=1.29
+ $X2=0 $Y2=0
cc_300 N_A_251_475#_M1013_g N_A_646_47#_c_793_n 0.00218095f $X=3.34 $Y=2.715
+ $X2=0 $Y2=0
cc_301 N_A_251_475#_c_252_n N_A_646_47#_c_793_n 0.00850434f $X=3.62 $Y=1.59
+ $X2=0 $Y2=0
cc_302 N_A_251_475#_c_253_n N_A_646_47#_c_793_n 0.00204239f $X=3.415 $Y=1.59
+ $X2=0 $Y2=0
cc_303 N_A_251_475#_M1015_g N_A_646_47#_c_774_n 0.00138212f $X=3.695 $Y=0.445
+ $X2=0 $Y2=0
cc_304 N_A_251_475#_c_256_n N_A_646_47#_c_774_n 0.00149399f $X=3.59 $Y=0.79
+ $X2=0 $Y2=0
cc_305 N_A_251_475#_M1015_g N_A_646_47#_c_776_n 9.78418e-19 $X=3.695 $Y=0.445
+ $X2=0 $Y2=0
cc_306 N_A_251_475#_c_256_n N_A_646_47#_c_776_n 0.0128337f $X=3.59 $Y=0.79 $X2=0
+ $Y2=0
cc_307 N_A_251_475#_c_258_n N_A_646_47#_c_776_n 0.00151728f $X=3.675 $Y=1.125
+ $X2=0 $Y2=0
cc_308 N_A_251_475#_c_260_n N_A_646_47#_c_776_n 6.58751e-19 $X=3.785 $Y=1.29
+ $X2=0 $Y2=0
cc_309 N_A_251_475#_c_261_n N_A_646_47#_c_776_n 2.47255e-19 $X=3.785 $Y=1.29
+ $X2=0 $Y2=0
cc_310 N_A_251_475#_M1013_g N_A_646_47#_c_803_n 0.00412621f $X=3.34 $Y=2.715
+ $X2=0 $Y2=0
cc_311 N_A_251_475#_c_260_n N_A_646_47#_c_779_n 0.00842803f $X=3.785 $Y=1.29
+ $X2=0 $Y2=0
cc_312 N_A_251_475#_M1020_g N_VPWR_c_927_n 0.00357685f $X=2.255 $Y=2.715 $X2=0
+ $Y2=0
cc_313 N_A_251_475#_M1020_g N_VPWR_c_931_n 0.00323385f $X=2.255 $Y=2.715 $X2=0
+ $Y2=0
cc_314 N_A_251_475#_M1013_g N_VPWR_c_936_n 0.00333662f $X=3.34 $Y=2.715 $X2=0
+ $Y2=0
cc_315 N_A_251_475#_M1020_g N_VPWR_c_925_n 0.00591839f $X=2.255 $Y=2.715 $X2=0
+ $Y2=0
cc_316 N_A_251_475#_M1013_g N_VPWR_c_925_n 0.00550332f $X=3.34 $Y=2.715 $X2=0
+ $Y2=0
cc_317 N_A_251_475#_c_251_n N_VGND_c_1047_n 0.00303181f $X=2.365 $Y=0.765 $X2=0
+ $Y2=0
cc_318 N_A_251_475#_c_256_n N_VGND_c_1047_n 0.0157463f $X=3.59 $Y=0.79 $X2=0
+ $Y2=0
cc_319 N_A_251_475#_c_257_n N_VGND_c_1047_n 0.00246711f $X=2.51 $Y=0.79 $X2=0
+ $Y2=0
cc_320 N_A_251_475#_c_263_n N_VGND_c_1047_n 2.09386e-19 $X=2.365 $Y=1.1 $X2=0
+ $Y2=0
cc_321 N_A_251_475#_M1015_g N_VGND_c_1054_n 0.00357877f $X=3.695 $Y=0.445 $X2=0
+ $Y2=0
cc_322 N_A_251_475#_c_256_n N_VGND_c_1054_n 0.00849173f $X=3.59 $Y=0.79 $X2=0
+ $Y2=0
cc_323 N_A_251_475#_c_251_n N_VGND_c_1058_n 0.004324f $X=2.365 $Y=0.765 $X2=0
+ $Y2=0
cc_324 N_A_251_475#_c_257_n N_VGND_c_1058_n 0.00265363f $X=2.51 $Y=0.79 $X2=0
+ $Y2=0
cc_325 N_A_251_475#_c_315_p N_VGND_c_1058_n 0.0103973f $X=1.53 $Y=0.495 $X2=0
+ $Y2=0
cc_326 N_A_251_475#_c_263_n N_VGND_c_1058_n 0.00348222f $X=2.365 $Y=1.1 $X2=0
+ $Y2=0
cc_327 N_A_251_475#_c_251_n N_VGND_c_1061_n 0.00710831f $X=2.365 $Y=0.765 $X2=0
+ $Y2=0
cc_328 N_A_251_475#_M1015_g N_VGND_c_1061_n 0.00545075f $X=3.695 $Y=0.445 $X2=0
+ $Y2=0
cc_329 N_A_251_475#_c_256_n N_VGND_c_1061_n 0.015478f $X=3.59 $Y=0.79 $X2=0
+ $Y2=0
cc_330 N_A_251_475#_c_257_n N_VGND_c_1061_n 0.00456282f $X=2.51 $Y=0.79 $X2=0
+ $Y2=0
cc_331 N_A_251_475#_c_315_p N_VGND_c_1061_n 0.00828371f $X=1.53 $Y=0.495 $X2=0
+ $Y2=0
cc_332 N_A_251_475#_c_263_n N_VGND_c_1061_n 0.00457574f $X=2.365 $Y=1.1 $X2=0
+ $Y2=0
cc_333 N_A_40_54#_c_411_n N_A_383_479#_M1020_s 0.00275621f $X=2.305 $Y=2.97
+ $X2=0 $Y2=0
cc_334 N_A_40_54#_M1004_g N_A_383_479#_M1007_g 0.0749616f $X=2.795 $Y=0.445
+ $X2=0 $Y2=0
cc_335 N_A_40_54#_M1004_g N_A_383_479#_c_505_n 0.00440096f $X=2.795 $Y=0.445
+ $X2=0 $Y2=0
cc_336 N_A_40_54#_c_411_n N_A_383_479#_c_505_n 0.0182001f $X=2.305 $Y=2.97 $X2=0
+ $Y2=0
cc_337 N_A_40_54#_c_413_n N_A_383_479#_c_505_n 0.023348f $X=2.39 $Y=2.885 $X2=0
+ $Y2=0
cc_338 N_A_40_54#_c_415_n N_A_383_479#_c_505_n 0.0265568f $X=2.705 $Y=2.06 $X2=0
+ $Y2=0
cc_339 N_A_40_54#_c_416_n N_A_383_479#_c_505_n 8.10792e-19 $X=2.795 $Y=2.06
+ $X2=0 $Y2=0
cc_340 N_A_40_54#_M1004_g N_A_383_479#_c_497_n 0.0160193f $X=2.795 $Y=0.445
+ $X2=0 $Y2=0
cc_341 N_A_40_54#_c_415_n N_A_383_479#_c_497_n 0.0371843f $X=2.705 $Y=2.06 $X2=0
+ $Y2=0
cc_342 N_A_40_54#_c_416_n N_A_383_479#_c_497_n 0.00829522f $X=2.795 $Y=2.06
+ $X2=0 $Y2=0
cc_343 N_A_40_54#_M1004_g N_A_383_479#_c_498_n 0.00718543f $X=2.795 $Y=0.445
+ $X2=0 $Y2=0
cc_344 N_A_40_54#_M1004_g N_A_383_479#_c_507_n 0.00579343f $X=2.795 $Y=0.445
+ $X2=0 $Y2=0
cc_345 N_A_40_54#_M1010_g N_A_383_479#_c_507_n 0.0116023f $X=2.98 $Y=2.715 $X2=0
+ $Y2=0
cc_346 N_A_40_54#_c_413_n N_A_383_479#_c_507_n 0.00516359f $X=2.39 $Y=2.885
+ $X2=0 $Y2=0
cc_347 N_A_40_54#_c_415_n N_A_383_479#_c_507_n 0.0251403f $X=2.705 $Y=2.06 $X2=0
+ $Y2=0
cc_348 N_A_40_54#_c_416_n N_A_383_479#_c_507_n 0.00463778f $X=2.795 $Y=2.06
+ $X2=0 $Y2=0
cc_349 N_A_40_54#_M1010_g N_A_383_479#_c_584_n 0.00414592f $X=2.98 $Y=2.715
+ $X2=0 $Y2=0
cc_350 N_A_40_54#_M1004_g N_A_383_479#_c_501_n 0.00260402f $X=2.795 $Y=0.445
+ $X2=0 $Y2=0
cc_351 N_A_40_54#_c_416_n N_A_646_47#_c_782_n 2.88863e-19 $X=2.795 $Y=2.06 $X2=0
+ $Y2=0
cc_352 N_A_40_54#_M1010_g N_A_646_47#_c_803_n 2.17258e-19 $X=2.98 $Y=2.715 $X2=0
+ $Y2=0
cc_353 N_A_40_54#_c_410_n N_VPWR_M1017_d 0.00623802f $X=1.02 $Y=2.44 $X2=-0.19
+ $Y2=-0.245
cc_354 N_A_40_54#_c_421_n N_VPWR_M1017_d 0.00422517f $X=1.105 $Y=2.885 $X2=-0.19
+ $Y2=-0.245
cc_355 N_A_40_54#_c_412_n N_VPWR_M1017_d 0.00124015f $X=1.19 $Y=2.97 $X2=-0.19
+ $Y2=-0.245
cc_356 N_A_40_54#_c_411_n N_VPWR_M1020_d 0.00144407f $X=2.305 $Y=2.97 $X2=0
+ $Y2=0
cc_357 N_A_40_54#_c_413_n N_VPWR_M1020_d 0.00452291f $X=2.39 $Y=2.885 $X2=0
+ $Y2=0
cc_358 N_A_40_54#_c_410_n N_VPWR_c_926_n 0.0151103f $X=1.02 $Y=2.44 $X2=0 $Y2=0
cc_359 N_A_40_54#_c_421_n N_VPWR_c_926_n 0.0141742f $X=1.105 $Y=2.885 $X2=0
+ $Y2=0
cc_360 N_A_40_54#_c_412_n N_VPWR_c_926_n 0.0143276f $X=1.19 $Y=2.97 $X2=0 $Y2=0
cc_361 N_A_40_54#_c_414_n N_VPWR_c_926_n 0.0122299f $X=0.325 $Y=2.52 $X2=0 $Y2=0
cc_362 N_A_40_54#_M1010_g N_VPWR_c_927_n 0.00563753f $X=2.98 $Y=2.715 $X2=0
+ $Y2=0
cc_363 N_A_40_54#_c_411_n N_VPWR_c_927_n 0.0139977f $X=2.305 $Y=2.97 $X2=0 $Y2=0
cc_364 N_A_40_54#_c_413_n N_VPWR_c_927_n 0.0358532f $X=2.39 $Y=2.885 $X2=0 $Y2=0
cc_365 N_A_40_54#_c_415_n N_VPWR_c_927_n 0.0155252f $X=2.705 $Y=2.06 $X2=0 $Y2=0
cc_366 N_A_40_54#_c_416_n N_VPWR_c_927_n 0.00482922f $X=2.795 $Y=2.06 $X2=0
+ $Y2=0
cc_367 N_A_40_54#_c_411_n N_VPWR_c_931_n 0.0740034f $X=2.305 $Y=2.97 $X2=0 $Y2=0
cc_368 N_A_40_54#_c_412_n N_VPWR_c_931_n 0.0105501f $X=1.19 $Y=2.97 $X2=0 $Y2=0
cc_369 N_A_40_54#_c_414_n N_VPWR_c_935_n 0.0145785f $X=0.325 $Y=2.52 $X2=0 $Y2=0
cc_370 N_A_40_54#_M1010_g N_VPWR_c_936_n 0.00462271f $X=2.98 $Y=2.715 $X2=0
+ $Y2=0
cc_371 N_A_40_54#_M1010_g N_VPWR_c_925_n 0.0086586f $X=2.98 $Y=2.715 $X2=0 $Y2=0
cc_372 N_A_40_54#_c_410_n N_VPWR_c_925_n 0.0119779f $X=1.02 $Y=2.44 $X2=0 $Y2=0
cc_373 N_A_40_54#_c_411_n N_VPWR_c_925_n 0.0469642f $X=2.305 $Y=2.97 $X2=0 $Y2=0
cc_374 N_A_40_54#_c_412_n N_VPWR_c_925_n 0.00615681f $X=1.19 $Y=2.97 $X2=0 $Y2=0
cc_375 N_A_40_54#_c_414_n N_VPWR_c_925_n 0.0101572f $X=0.325 $Y=2.52 $X2=0 $Y2=0
cc_376 N_A_40_54#_M1004_g N_VGND_c_1047_n 0.0101293f $X=2.795 $Y=0.445 $X2=0
+ $Y2=0
cc_377 N_A_40_54#_c_406_n N_VGND_c_1052_n 0.0125783f $X=0.325 $Y=0.48 $X2=0
+ $Y2=0
cc_378 N_A_40_54#_M1004_g N_VGND_c_1054_n 0.00361815f $X=2.795 $Y=0.445 $X2=0
+ $Y2=0
cc_379 N_A_40_54#_M1004_g N_VGND_c_1061_n 0.00416812f $X=2.795 $Y=0.445 $X2=0
+ $Y2=0
cc_380 N_A_40_54#_c_406_n N_VGND_c_1061_n 0.00934149f $X=0.325 $Y=0.48 $X2=0
+ $Y2=0
cc_381 N_A_383_479#_M1014_g N_A_796_21#_M1000_g 0.0348386f $X=3.85 $Y=2.605
+ $X2=0 $Y2=0
cc_382 N_A_383_479#_c_508_n N_A_796_21#_M1000_g 9.43202e-19 $X=3.9 $Y=2.91 $X2=0
+ $Y2=0
cc_383 N_A_383_479#_c_509_n N_A_796_21#_M1000_g 0.00708188f $X=3.985 $Y=2.825
+ $X2=0 $Y2=0
cc_384 N_A_383_479#_c_512_n N_A_796_21#_c_644_n 2.88089e-19 $X=3.79 $Y=2.07
+ $X2=0 $Y2=0
cc_385 N_A_383_479#_c_513_n N_A_796_21#_c_644_n 0.0278683f $X=3.985 $Y=2.07
+ $X2=0 $Y2=0
cc_386 N_A_383_479#_c_512_n N_A_796_21#_c_645_n 0.0204765f $X=3.79 $Y=2.07 $X2=0
+ $Y2=0
cc_387 N_A_383_479#_c_513_n N_A_796_21#_c_645_n 0.0021731f $X=3.985 $Y=2.07
+ $X2=0 $Y2=0
cc_388 N_A_383_479#_c_508_n N_A_646_47#_M1013_d 0.0041535f $X=3.9 $Y=2.91 $X2=0
+ $Y2=0
cc_389 N_A_383_479#_M1007_g N_A_646_47#_c_786_n 0.00432694f $X=3.155 $Y=0.445
+ $X2=0 $Y2=0
cc_390 N_A_383_479#_M1014_g N_A_646_47#_c_782_n 0.00125567f $X=3.85 $Y=2.605
+ $X2=0 $Y2=0
cc_391 N_A_383_479#_c_507_n N_A_646_47#_c_782_n 0.0465408f $X=3.09 $Y=2.825
+ $X2=0 $Y2=0
cc_392 N_A_383_479#_c_509_n N_A_646_47#_c_782_n 0.00671469f $X=3.985 $Y=2.825
+ $X2=0 $Y2=0
cc_393 N_A_383_479#_c_512_n N_A_646_47#_c_782_n 0.00207715f $X=3.79 $Y=2.07
+ $X2=0 $Y2=0
cc_394 N_A_383_479#_c_513_n N_A_646_47#_c_782_n 0.0239023f $X=3.985 $Y=2.07
+ $X2=0 $Y2=0
cc_395 N_A_383_479#_c_512_n N_A_646_47#_c_773_n 0.00324752f $X=3.79 $Y=2.07
+ $X2=0 $Y2=0
cc_396 N_A_383_479#_c_513_n N_A_646_47#_c_773_n 0.0267549f $X=3.985 $Y=2.07
+ $X2=0 $Y2=0
cc_397 N_A_383_479#_c_507_n N_A_646_47#_c_793_n 0.00149384f $X=3.09 $Y=2.825
+ $X2=0 $Y2=0
cc_398 N_A_383_479#_c_501_n N_A_646_47#_c_793_n 0.00316658f $X=3.245 $Y=1.14
+ $X2=0 $Y2=0
cc_399 N_A_383_479#_c_503_n N_A_646_47#_c_793_n 0.0127623f $X=3.09 $Y=1.62 $X2=0
+ $Y2=0
cc_400 N_A_383_479#_c_507_n N_A_646_47#_c_803_n 0.0177417f $X=3.09 $Y=2.825
+ $X2=0 $Y2=0
cc_401 N_A_383_479#_c_508_n N_A_646_47#_c_803_n 0.02165f $X=3.9 $Y=2.91 $X2=0
+ $Y2=0
cc_402 N_A_383_479#_c_512_n N_A_646_47#_c_803_n 0.00346876f $X=3.79 $Y=2.07
+ $X2=0 $Y2=0
cc_403 N_A_383_479#_c_513_n N_A_646_47#_c_803_n 0.00106301f $X=3.985 $Y=2.07
+ $X2=0 $Y2=0
cc_404 N_A_383_479#_c_507_n N_VPWR_c_927_n 0.0304165f $X=3.09 $Y=2.825 $X2=0
+ $Y2=0
cc_405 N_A_383_479#_c_584_n N_VPWR_c_927_n 0.013466f $X=3.175 $Y=2.91 $X2=0
+ $Y2=0
cc_406 N_A_383_479#_M1014_g N_VPWR_c_936_n 7.79124e-19 $X=3.85 $Y=2.605 $X2=0
+ $Y2=0
cc_407 N_A_383_479#_c_508_n N_VPWR_c_936_n 0.0364076f $X=3.9 $Y=2.91 $X2=0 $Y2=0
cc_408 N_A_383_479#_c_584_n N_VPWR_c_936_n 0.00647547f $X=3.175 $Y=2.91 $X2=0
+ $Y2=0
cc_409 N_A_383_479#_M1014_g N_VPWR_c_939_n 4.23432e-19 $X=3.85 $Y=2.605 $X2=0
+ $Y2=0
cc_410 N_A_383_479#_c_508_n N_VPWR_c_939_n 0.0127069f $X=3.9 $Y=2.91 $X2=0 $Y2=0
cc_411 N_A_383_479#_c_509_n N_VPWR_c_939_n 0.0244503f $X=3.985 $Y=2.825 $X2=0
+ $Y2=0
cc_412 N_A_383_479#_c_508_n N_VPWR_c_925_n 0.031515f $X=3.9 $Y=2.91 $X2=0 $Y2=0
cc_413 N_A_383_479#_c_584_n N_VPWR_c_925_n 0.00608328f $X=3.175 $Y=2.91 $X2=0
+ $Y2=0
cc_414 N_A_383_479#_c_507_n A_611_479# 0.00404206f $X=3.09 $Y=2.825 $X2=-0.19
+ $Y2=-0.245
cc_415 N_A_383_479#_c_508_n A_611_479# 0.00157486f $X=3.9 $Y=2.91 $X2=-0.19
+ $Y2=-0.245
cc_416 N_A_383_479#_c_584_n A_611_479# 7.1501e-19 $X=3.175 $Y=2.91 $X2=-0.19
+ $Y2=-0.245
cc_417 N_A_383_479#_c_509_n A_785_479# 0.00389099f $X=3.985 $Y=2.825 $X2=-0.19
+ $Y2=-0.245
cc_418 N_A_383_479#_c_499_n N_VGND_c_1046_n 0.00147674f $X=2.13 $Y=0.42 $X2=0
+ $Y2=0
cc_419 N_A_383_479#_M1007_g N_VGND_c_1047_n 0.00203054f $X=3.155 $Y=0.445 $X2=0
+ $Y2=0
cc_420 N_A_383_479#_M1007_g N_VGND_c_1054_n 0.00435108f $X=3.155 $Y=0.445 $X2=0
+ $Y2=0
cc_421 N_A_383_479#_c_499_n N_VGND_c_1058_n 0.0295908f $X=2.13 $Y=0.42 $X2=0
+ $Y2=0
cc_422 N_A_383_479#_M1021_s N_VGND_c_1061_n 0.00228716f $X=2.005 $Y=0.235 $X2=0
+ $Y2=0
cc_423 N_A_383_479#_M1007_g N_VGND_c_1061_n 0.00631645f $X=3.155 $Y=0.445 $X2=0
+ $Y2=0
cc_424 N_A_383_479#_c_499_n N_VGND_c_1061_n 0.0179621f $X=2.13 $Y=0.42 $X2=0
+ $Y2=0
cc_425 N_A_796_21#_c_635_n N_A_646_47#_c_768_n 0.0260981f $X=4.24 $Y=0.84 $X2=0
+ $Y2=0
cc_426 N_A_796_21#_c_637_n N_A_646_47#_c_768_n 0.0100288f $X=4.925 $Y=0.51 $X2=0
+ $Y2=0
cc_427 N_A_796_21#_c_638_n N_A_646_47#_c_768_n 0.00117407f $X=5.04 $Y=1.905
+ $X2=0 $Y2=0
cc_428 N_A_796_21#_c_637_n N_A_646_47#_c_769_n 0.00379632f $X=4.925 $Y=0.51
+ $X2=0 $Y2=0
cc_429 N_A_796_21#_c_630_n N_A_646_47#_c_770_n 0.0146041f $X=4.055 $Y=0.765
+ $X2=0 $Y2=0
cc_430 N_A_796_21#_c_638_n N_A_646_47#_c_771_n 0.0113957f $X=5.04 $Y=1.905 $X2=0
+ $Y2=0
cc_431 N_A_796_21#_c_668_p N_A_646_47#_c_771_n 0.00327631f $X=4.967 $Y=1.165
+ $X2=0 $Y2=0
cc_432 N_A_796_21#_c_637_n N_A_646_47#_c_772_n 0.0143781f $X=4.925 $Y=0.51 $X2=0
+ $Y2=0
cc_433 N_A_796_21#_c_638_n N_A_646_47#_c_772_n 0.00416646f $X=5.04 $Y=1.905
+ $X2=0 $Y2=0
cc_434 N_A_796_21#_c_668_p N_A_646_47#_c_772_n 0.00308101f $X=4.967 $Y=1.165
+ $X2=0 $Y2=0
cc_435 N_A_796_21#_c_672_p N_A_646_47#_c_772_n 3.28151e-19 $X=5.355 $Y=2.445
+ $X2=0 $Y2=0
cc_436 N_A_796_21#_c_645_n N_A_646_47#_M1012_g 0.00508394f $X=4.335 $Y=2.07
+ $X2=0 $Y2=0
cc_437 N_A_796_21#_c_638_n N_A_646_47#_M1012_g 0.00718227f $X=5.04 $Y=1.905
+ $X2=0 $Y2=0
cc_438 N_A_796_21#_c_672_p N_A_646_47#_M1012_g 0.0277419f $X=5.355 $Y=2.445
+ $X2=0 $Y2=0
cc_439 N_A_796_21#_c_630_n N_A_646_47#_c_786_n 0.00845782f $X=4.055 $Y=0.765
+ $X2=0 $Y2=0
cc_440 N_A_796_21#_c_639_n N_A_646_47#_c_782_n 0.00377268f $X=4.332 $Y=1.905
+ $X2=0 $Y2=0
cc_441 N_A_796_21#_c_635_n N_A_646_47#_c_773_n 0.00318545f $X=4.24 $Y=0.84 $X2=0
+ $Y2=0
cc_442 N_A_796_21#_c_644_n N_A_646_47#_c_773_n 0.0162742f $X=4.955 $Y=2.07 $X2=0
+ $Y2=0
cc_443 N_A_796_21#_c_645_n N_A_646_47#_c_773_n 0.00345287f $X=4.335 $Y=2.07
+ $X2=0 $Y2=0
cc_444 N_A_796_21#_c_639_n N_A_646_47#_c_773_n 0.0148286f $X=4.332 $Y=1.905
+ $X2=0 $Y2=0
cc_445 N_A_796_21#_c_630_n N_A_646_47#_c_774_n 0.00540311f $X=4.055 $Y=0.765
+ $X2=0 $Y2=0
cc_446 N_A_796_21#_c_630_n N_A_646_47#_c_775_n 0.00117218f $X=4.055 $Y=0.765
+ $X2=0 $Y2=0
cc_447 N_A_796_21#_c_635_n N_A_646_47#_c_775_n 0.0117781f $X=4.24 $Y=0.84 $X2=0
+ $Y2=0
cc_448 N_A_796_21#_c_637_n N_A_646_47#_c_775_n 0.0139928f $X=4.925 $Y=0.51 $X2=0
+ $Y2=0
cc_449 N_A_796_21#_c_630_n N_A_646_47#_c_776_n 5.74535e-19 $X=4.055 $Y=0.765
+ $X2=0 $Y2=0
cc_450 N_A_796_21#_c_635_n N_A_646_47#_c_776_n 0.00414293f $X=4.24 $Y=0.84 $X2=0
+ $Y2=0
cc_451 N_A_796_21#_c_644_n N_A_646_47#_c_777_n 0.0251337f $X=4.955 $Y=2.07 $X2=0
+ $Y2=0
cc_452 N_A_796_21#_c_645_n N_A_646_47#_c_777_n 6.72244e-19 $X=4.335 $Y=2.07
+ $X2=0 $Y2=0
cc_453 N_A_796_21#_c_638_n N_A_646_47#_c_777_n 0.0274632f $X=5.04 $Y=1.905 $X2=0
+ $Y2=0
cc_454 N_A_796_21#_c_639_n N_A_646_47#_c_777_n 0.00584257f $X=4.332 $Y=1.905
+ $X2=0 $Y2=0
cc_455 N_A_796_21#_c_644_n N_A_646_47#_c_778_n 0.00827028f $X=4.955 $Y=2.07
+ $X2=0 $Y2=0
cc_456 N_A_796_21#_c_638_n N_A_646_47#_c_778_n 0.00231029f $X=5.04 $Y=1.905
+ $X2=0 $Y2=0
cc_457 N_A_796_21#_c_668_p N_A_646_47#_c_778_n 0.00197328f $X=4.967 $Y=1.165
+ $X2=0 $Y2=0
cc_458 N_A_796_21#_c_639_n N_A_646_47#_c_778_n 0.0209826f $X=4.332 $Y=1.905
+ $X2=0 $Y2=0
cc_459 N_A_796_21#_c_635_n N_A_646_47#_c_779_n 0.00555793f $X=4.24 $Y=0.84 $X2=0
+ $Y2=0
cc_460 N_A_796_21#_c_637_n N_A_646_47#_c_779_n 0.0198294f $X=4.925 $Y=0.51 $X2=0
+ $Y2=0
cc_461 N_A_796_21#_c_638_n N_A_646_47#_c_779_n 0.00758407f $X=5.04 $Y=1.905
+ $X2=0 $Y2=0
cc_462 N_A_796_21#_M1001_g N_RESET_B_M1018_g 0.0249131f $X=6.265 $Y=2.465 $X2=0
+ $Y2=0
cc_463 N_A_796_21#_c_638_n N_RESET_B_M1018_g 7.25433e-19 $X=5.04 $Y=1.905 $X2=0
+ $Y2=0
cc_464 N_A_796_21#_c_701_p N_RESET_B_M1018_g 0.0140739f $X=5.965 $Y=2.01 $X2=0
+ $Y2=0
cc_465 N_A_796_21#_c_647_n N_RESET_B_M1018_g 0.00384636f $X=6.13 $Y=1.51 $X2=0
+ $Y2=0
cc_466 N_A_796_21#_c_640_n N_RESET_B_M1018_g 0.00109602f $X=6.34 $Y=1.51 $X2=0
+ $Y2=0
cc_467 N_A_796_21#_M1006_g RESET_B 0.0034f $X=6.04 $Y=0.785 $X2=0 $Y2=0
cc_468 N_A_796_21#_M1001_g RESET_B 2.25506e-19 $X=6.265 $Y=2.465 $X2=0 $Y2=0
cc_469 N_A_796_21#_c_638_n RESET_B 0.0335638f $X=5.04 $Y=1.905 $X2=0 $Y2=0
cc_470 N_A_796_21#_c_701_p RESET_B 0.0136198f $X=5.965 $Y=2.01 $X2=0 $Y2=0
cc_471 N_A_796_21#_c_647_n RESET_B 0.0204023f $X=6.13 $Y=1.51 $X2=0 $Y2=0
cc_472 N_A_796_21#_c_672_p RESET_B 0.0088626f $X=5.355 $Y=2.445 $X2=0 $Y2=0
cc_473 N_A_796_21#_c_640_n RESET_B 2.09162e-19 $X=6.34 $Y=1.51 $X2=0 $Y2=0
cc_474 N_A_796_21#_M1006_g N_RESET_B_c_888_n 0.021082f $X=6.04 $Y=0.785 $X2=0
+ $Y2=0
cc_475 N_A_796_21#_c_638_n N_RESET_B_c_888_n 8.05347e-19 $X=5.04 $Y=1.905 $X2=0
+ $Y2=0
cc_476 N_A_796_21#_c_701_p N_RESET_B_c_888_n 0.00227332f $X=5.965 $Y=2.01 $X2=0
+ $Y2=0
cc_477 N_A_796_21#_c_647_n N_RESET_B_c_888_n 0.00111105f $X=6.13 $Y=1.51 $X2=0
+ $Y2=0
cc_478 N_A_796_21#_M1006_g N_RESET_B_c_889_n 0.00894998f $X=6.04 $Y=0.785 $X2=0
+ $Y2=0
cc_479 N_A_796_21#_c_637_n N_RESET_B_c_889_n 0.00298394f $X=4.925 $Y=0.51 $X2=0
+ $Y2=0
cc_480 N_A_796_21#_c_644_n N_VPWR_M1000_d 0.00603993f $X=4.955 $Y=2.07 $X2=0
+ $Y2=0
cc_481 N_A_796_21#_c_638_n N_VPWR_M1000_d 0.00119436f $X=5.04 $Y=1.905 $X2=0
+ $Y2=0
cc_482 N_A_796_21#_c_672_p N_VPWR_M1000_d 0.0048328f $X=5.355 $Y=2.445 $X2=0
+ $Y2=0
cc_483 N_A_796_21#_c_701_p N_VPWR_M1018_d 0.0181805f $X=5.965 $Y=2.01 $X2=0
+ $Y2=0
cc_484 N_A_796_21#_c_647_n N_VPWR_M1018_d 0.00138878f $X=6.13 $Y=1.51 $X2=0
+ $Y2=0
cc_485 N_A_796_21#_M1001_g N_VPWR_c_928_n 0.0111903f $X=6.265 $Y=2.465 $X2=0
+ $Y2=0
cc_486 N_A_796_21#_c_701_p N_VPWR_c_928_n 0.0276076f $X=5.965 $Y=2.01 $X2=0
+ $Y2=0
cc_487 N_A_796_21#_c_640_n N_VPWR_c_928_n 3.77354e-19 $X=6.34 $Y=1.51 $X2=0
+ $Y2=0
cc_488 N_A_796_21#_M1001_g N_VPWR_c_930_n 8.786e-19 $X=6.265 $Y=2.465 $X2=0
+ $Y2=0
cc_489 N_A_796_21#_M1009_g N_VPWR_c_930_n 0.0242625f $X=6.695 $Y=2.465 $X2=0
+ $Y2=0
cc_490 N_A_796_21#_c_672_p N_VPWR_c_933_n 0.0145813f $X=5.355 $Y=2.445 $X2=0
+ $Y2=0
cc_491 N_A_796_21#_M1000_g N_VPWR_c_936_n 0.00397465f $X=4.24 $Y=2.605 $X2=0
+ $Y2=0
cc_492 N_A_796_21#_M1001_g N_VPWR_c_937_n 0.00585385f $X=6.265 $Y=2.465 $X2=0
+ $Y2=0
cc_493 N_A_796_21#_M1009_g N_VPWR_c_937_n 0.00447018f $X=6.695 $Y=2.465 $X2=0
+ $Y2=0
cc_494 N_A_796_21#_M1000_g N_VPWR_c_939_n 0.010106f $X=4.24 $Y=2.605 $X2=0 $Y2=0
cc_495 N_A_796_21#_c_644_n N_VPWR_c_939_n 0.0420141f $X=4.955 $Y=2.07 $X2=0
+ $Y2=0
cc_496 N_A_796_21#_c_645_n N_VPWR_c_939_n 0.00404012f $X=4.335 $Y=2.07 $X2=0
+ $Y2=0
cc_497 N_A_796_21#_c_672_p N_VPWR_c_939_n 0.00645883f $X=5.355 $Y=2.445 $X2=0
+ $Y2=0
cc_498 N_A_796_21#_M1012_d N_VPWR_c_925_n 0.00327921f $X=5.215 $Y=1.835 $X2=0
+ $Y2=0
cc_499 N_A_796_21#_M1000_g N_VPWR_c_925_n 0.00417428f $X=4.24 $Y=2.605 $X2=0
+ $Y2=0
cc_500 N_A_796_21#_M1001_g N_VPWR_c_925_n 0.0114504f $X=6.265 $Y=2.465 $X2=0
+ $Y2=0
cc_501 N_A_796_21#_M1009_g N_VPWR_c_925_n 0.00762944f $X=6.695 $Y=2.465 $X2=0
+ $Y2=0
cc_502 N_A_796_21#_c_672_p N_VPWR_c_925_n 0.00964167f $X=5.355 $Y=2.445 $X2=0
+ $Y2=0
cc_503 N_A_796_21#_M1016_g Q 0.00256193f $X=6.585 $Y=0.785 $X2=0 $Y2=0
cc_504 N_A_796_21#_c_647_n Q 0.00413663f $X=6.13 $Y=1.51 $X2=0 $Y2=0
cc_505 N_A_796_21#_c_640_n Q 0.0083201f $X=6.34 $Y=1.51 $X2=0 $Y2=0
cc_506 N_A_796_21#_M1006_g Q 0.00330001f $X=6.04 $Y=0.785 $X2=0 $Y2=0
cc_507 N_A_796_21#_c_632_n Q 0.00657641f $X=6.51 $Y=1.42 $X2=0 $Y2=0
cc_508 N_A_796_21#_M1016_g Q 0.00701066f $X=6.585 $Y=0.785 $X2=0 $Y2=0
cc_509 N_A_796_21#_M1009_g Q 0.00848518f $X=6.695 $Y=2.465 $X2=0 $Y2=0
cc_510 N_A_796_21#_c_636_n Q 0.0071612f $X=6.695 $Y=1.42 $X2=0 $Y2=0
cc_511 N_A_796_21#_c_647_n Q 0.0387788f $X=6.13 $Y=1.51 $X2=0 $Y2=0
cc_512 N_A_796_21#_c_640_n Q 0.00325596f $X=6.34 $Y=1.51 $X2=0 $Y2=0
cc_513 N_A_796_21#_M1006_g N_Q_c_1024_n 0.00487586f $X=6.04 $Y=0.785 $X2=0 $Y2=0
cc_514 N_A_796_21#_M1016_g N_Q_c_1024_n 0.010237f $X=6.585 $Y=0.785 $X2=0 $Y2=0
cc_515 N_A_796_21#_c_630_n N_VGND_c_1048_n 0.0051034f $X=4.055 $Y=0.765 $X2=0
+ $Y2=0
cc_516 N_A_796_21#_c_635_n N_VGND_c_1048_n 2.3658e-19 $X=4.24 $Y=0.84 $X2=0
+ $Y2=0
cc_517 N_A_796_21#_c_637_n N_VGND_c_1048_n 0.00995915f $X=4.925 $Y=0.51 $X2=0
+ $Y2=0
cc_518 N_A_796_21#_M1006_g N_VGND_c_1049_n 0.00370895f $X=6.04 $Y=0.785 $X2=0
+ $Y2=0
cc_519 N_A_796_21#_c_637_n N_VGND_c_1049_n 0.0114921f $X=4.925 $Y=0.51 $X2=0
+ $Y2=0
cc_520 N_A_796_21#_M1016_g N_VGND_c_1051_n 0.0106135f $X=6.585 $Y=0.785 $X2=0
+ $Y2=0
cc_521 N_A_796_21#_c_636_n N_VGND_c_1051_n 0.00120394f $X=6.695 $Y=1.42 $X2=0
+ $Y2=0
cc_522 N_A_796_21#_c_630_n N_VGND_c_1054_n 0.00368359f $X=4.055 $Y=0.765 $X2=0
+ $Y2=0
cc_523 N_A_796_21#_c_635_n N_VGND_c_1054_n 4.89446e-19 $X=4.24 $Y=0.84 $X2=0
+ $Y2=0
cc_524 N_A_796_21#_c_637_n N_VGND_c_1056_n 0.0140681f $X=4.925 $Y=0.51 $X2=0
+ $Y2=0
cc_525 N_A_796_21#_M1006_g N_VGND_c_1059_n 0.00465548f $X=6.04 $Y=0.785 $X2=0
+ $Y2=0
cc_526 N_A_796_21#_M1016_g N_VGND_c_1059_n 0.00403641f $X=6.585 $Y=0.785 $X2=0
+ $Y2=0
cc_527 N_A_796_21#_c_630_n N_VGND_c_1061_n 0.00576395f $X=4.055 $Y=0.765 $X2=0
+ $Y2=0
cc_528 N_A_796_21#_M1006_g N_VGND_c_1061_n 0.00919412f $X=6.04 $Y=0.785 $X2=0
+ $Y2=0
cc_529 N_A_796_21#_M1016_g N_VGND_c_1061_n 0.00729083f $X=6.585 $Y=0.785 $X2=0
+ $Y2=0
cc_530 N_A_796_21#_c_637_n N_VGND_c_1061_n 0.0102659f $X=4.925 $Y=0.51 $X2=0
+ $Y2=0
cc_531 N_A_646_47#_c_771_n N_RESET_B_M1018_g 0.0191745f $X=5.065 $Y=1.62 $X2=0
+ $Y2=0
cc_532 N_A_646_47#_c_771_n RESET_B 0.00158234f $X=5.065 $Y=1.62 $X2=0 $Y2=0
cc_533 N_A_646_47#_c_772_n RESET_B 7.8519e-19 $X=5.14 $Y=0.255 $X2=0 $Y2=0
cc_534 N_A_646_47#_c_771_n N_RESET_B_c_888_n 0.0065766f $X=5.065 $Y=1.62 $X2=0
+ $Y2=0
cc_535 N_A_646_47#_c_772_n N_RESET_B_c_888_n 0.0320383f $X=5.14 $Y=0.255 $X2=0
+ $Y2=0
cc_536 N_A_646_47#_c_778_n N_RESET_B_c_888_n 0.00297489f $X=4.69 $Y=1.5 $X2=0
+ $Y2=0
cc_537 N_A_646_47#_c_769_n N_RESET_B_c_889_n 0.0320383f $X=5.065 $Y=0.18 $X2=0
+ $Y2=0
cc_538 N_A_646_47#_M1012_g N_VPWR_c_933_n 0.00585385f $X=5.14 $Y=2.465 $X2=0
+ $Y2=0
cc_539 N_A_646_47#_M1012_g N_VPWR_c_939_n 0.0103899f $X=5.14 $Y=2.465 $X2=0
+ $Y2=0
cc_540 N_A_646_47#_M1012_g N_VPWR_c_925_n 0.0120657f $X=5.14 $Y=2.465 $X2=0
+ $Y2=0
cc_541 N_A_646_47#_c_786_n N_VGND_c_1047_n 0.00877218f $X=3.94 $Y=0.395 $X2=0
+ $Y2=0
cc_542 N_A_646_47#_c_770_n N_VGND_c_1048_n 0.0077975f $X=4.725 $Y=0.18 $X2=0
+ $Y2=0
cc_543 N_A_646_47#_c_786_n N_VGND_c_1048_n 0.0222597f $X=3.94 $Y=0.395 $X2=0
+ $Y2=0
cc_544 N_A_646_47#_c_774_n N_VGND_c_1048_n 0.00138813f $X=4.025 $Y=0.725 $X2=0
+ $Y2=0
cc_545 N_A_646_47#_c_775_n N_VGND_c_1048_n 0.0157746f $X=4.47 $Y=0.81 $X2=0
+ $Y2=0
cc_546 N_A_646_47#_c_769_n N_VGND_c_1049_n 0.00409708f $X=5.065 $Y=0.18 $X2=0
+ $Y2=0
cc_547 N_A_646_47#_c_786_n N_VGND_c_1054_n 0.0469293f $X=3.94 $Y=0.395 $X2=0
+ $Y2=0
cc_548 N_A_646_47#_c_775_n N_VGND_c_1054_n 0.00253464f $X=4.47 $Y=0.81 $X2=0
+ $Y2=0
cc_549 N_A_646_47#_c_770_n N_VGND_c_1056_n 0.0193242f $X=4.725 $Y=0.18 $X2=0
+ $Y2=0
cc_550 N_A_646_47#_c_775_n N_VGND_c_1056_n 0.0025622f $X=4.47 $Y=0.81 $X2=0
+ $Y2=0
cc_551 N_A_646_47#_M1007_d N_VGND_c_1061_n 0.00353059f $X=3.23 $Y=0.235 $X2=0
+ $Y2=0
cc_552 N_A_646_47#_c_769_n N_VGND_c_1061_n 0.0206334f $X=5.065 $Y=0.18 $X2=0
+ $Y2=0
cc_553 N_A_646_47#_c_770_n N_VGND_c_1061_n 0.00848199f $X=4.725 $Y=0.18 $X2=0
+ $Y2=0
cc_554 N_A_646_47#_c_786_n N_VGND_c_1061_n 0.0290017f $X=3.94 $Y=0.395 $X2=0
+ $Y2=0
cc_555 N_A_646_47#_c_775_n N_VGND_c_1061_n 0.00947637f $X=4.47 $Y=0.81 $X2=0
+ $Y2=0
cc_556 N_A_646_47#_c_786_n A_754_47# 0.00257434f $X=3.94 $Y=0.395 $X2=-0.19
+ $Y2=-0.245
cc_557 N_RESET_B_M1018_g N_VPWR_c_928_n 0.0124789f $X=5.57 $Y=2.465 $X2=0 $Y2=0
cc_558 N_RESET_B_M1018_g N_VPWR_c_933_n 0.00585385f $X=5.57 $Y=2.465 $X2=0 $Y2=0
cc_559 N_RESET_B_M1018_g N_VPWR_c_925_n 0.0114757f $X=5.57 $Y=2.465 $X2=0 $Y2=0
cc_560 RESET_B N_VGND_c_1049_n 0.00497483f $X=5.435 $Y=1.21 $X2=0 $Y2=0
cc_561 N_RESET_B_c_888_n N_VGND_c_1049_n 0.00356347f $X=5.59 $Y=1.48 $X2=0 $Y2=0
cc_562 N_RESET_B_c_889_n N_VGND_c_1049_n 0.00378434f $X=5.59 $Y=1.315 $X2=0
+ $Y2=0
cc_563 N_RESET_B_c_889_n N_VGND_c_1056_n 0.00465548f $X=5.59 $Y=1.315 $X2=0
+ $Y2=0
cc_564 N_RESET_B_c_889_n N_VGND_c_1061_n 0.00916139f $X=5.59 $Y=1.315 $X2=0
+ $Y2=0
cc_565 N_VPWR_c_925_n N_Q_M1001_s 0.00571434f $X=6.96 $Y=3.33 $X2=0 $Y2=0
cc_566 N_VPWR_c_930_n Q 0.0482158f $X=6.91 $Y=1.98 $X2=0 $Y2=0
cc_567 N_VPWR_c_937_n Q 0.0120977f $X=6.735 $Y=3.33 $X2=0 $Y2=0
cc_568 N_VPWR_c_925_n Q 0.00691495f $X=6.96 $Y=3.33 $X2=0 $Y2=0
cc_569 N_VPWR_c_930_n N_VGND_c_1051_n 0.00956613f $X=6.91 $Y=1.98 $X2=0 $Y2=0
cc_570 N_Q_c_1024_n N_VGND_c_1049_n 0.00131925f $X=6.325 $Y=0.51 $X2=0 $Y2=0
cc_571 N_Q_c_1024_n N_VGND_c_1051_n 0.0676849f $X=6.325 $Y=0.51 $X2=0 $Y2=0
cc_572 N_Q_c_1024_n N_VGND_c_1059_n 0.0181874f $X=6.325 $Y=0.51 $X2=0 $Y2=0
cc_573 N_Q_c_1024_n N_VGND_c_1061_n 0.0146688f $X=6.325 $Y=0.51 $X2=0 $Y2=0
cc_574 N_VGND_c_1061_n A_574_47# 0.00265743f $X=6.96 $Y=0 $X2=-0.19 $Y2=-0.245
cc_575 N_VGND_c_1061_n A_754_47# 0.00168887f $X=6.96 $Y=0 $X2=-0.19 $Y2=-0.245
