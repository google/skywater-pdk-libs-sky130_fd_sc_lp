# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_lp__o211ai_2
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.800000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.560000 1.420000 4.715000 1.590000 ;
        RECT 4.115000 1.210000 4.715000 1.420000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.075000 1.195000 2.735000 1.420000 ;
        RECT 2.075000 1.420000 3.280000 1.590000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.045000 1.210000 1.905000 1.525000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.210000 0.385000 1.285000 ;
        RECT 0.085000 1.285000 0.445000 1.750000 ;
    END
  END C1
  PIN Y
    ANTENNADIFFAREA  1.293600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.545000 0.595000 0.875000 1.145000 ;
        RECT 0.615000 1.145000 0.875000 1.760000 ;
        RECT 0.615000 1.760000 3.155000 1.930000 ;
        RECT 0.615000 1.930000 0.805000 3.075000 ;
        RECT 1.475000 1.930000 1.665000 3.075000 ;
        RECT 2.825000 1.930000 3.155000 2.735000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.800000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.500000 0.500000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.800000 0.500000 3.300000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.800000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.800000 0.085000 ;
      RECT 0.000000  3.245000 4.800000 3.415000 ;
      RECT 0.095000  0.255000 2.165000 0.425000 ;
      RECT 0.095000  0.425000 0.375000 1.040000 ;
      RECT 0.115000  1.920000 0.445000 3.245000 ;
      RECT 0.975000  2.100000 1.305000 3.245000 ;
      RECT 1.045000  0.425000 2.165000 0.645000 ;
      RECT 1.045000  0.645000 1.235000 1.040000 ;
      RECT 1.405000  0.815000 3.085000 1.025000 ;
      RECT 1.835000  2.100000 2.165000 3.245000 ;
      RECT 2.395000  0.085000 2.725000 0.645000 ;
      RECT 2.395000  2.100000 2.655000 2.905000 ;
      RECT 2.395000  2.905000 3.515000 3.075000 ;
      RECT 2.895000  0.255000 3.085000 0.815000 ;
      RECT 2.905000  1.025000 3.085000 1.080000 ;
      RECT 2.905000  1.080000 3.945000 1.250000 ;
      RECT 3.255000  0.085000 3.585000 0.910000 ;
      RECT 3.325000  1.760000 4.445000 1.930000 ;
      RECT 3.325000  1.930000 3.515000 2.905000 ;
      RECT 3.685000  2.100000 4.015000 3.245000 ;
      RECT 3.755000  0.255000 3.945000 1.080000 ;
      RECT 4.115000  0.085000 4.445000 1.040000 ;
      RECT 4.185000  1.930000 4.445000 3.075000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
  END
END sky130_fd_sc_lp__o211ai_2
END LIBRARY
