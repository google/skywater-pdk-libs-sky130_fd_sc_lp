* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__dlxbn_2 D GATE_N VGND VNB VPB VPWR Q Q_N
X0 VGND a_805_21# Q VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X1 a_769_491# a_805_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X2 VGND a_1138_153# Q_N VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X3 Q_N a_1138_153# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X4 a_589_491# a_354_47# a_619_47# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X5 VPWR a_619_47# a_805_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X6 VGND a_45_136# a_547_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 a_45_136# D VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 VPWR a_805_21# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X9 a_547_47# a_214_136# a_619_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 Q a_805_21# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X11 a_354_47# a_214_136# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X12 a_45_136# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X13 a_1138_153# a_805_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X14 Q a_805_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X15 VGND GATE_N a_214_136# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X16 VPWR a_1138_153# Q_N VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X17 a_354_47# a_214_136# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X18 a_619_47# a_354_47# a_737_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X19 a_619_47# a_214_136# a_769_491# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X20 a_1138_153# a_805_21# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X21 VPWR GATE_N a_214_136# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X22 VPWR a_45_136# a_589_491# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X23 Q_N a_1138_153# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X24 VGND a_619_47# a_805_21# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X25 a_737_47# a_805_21# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
