# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__o311a_4
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__o311a_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.160000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.285000 1.425000 8.075000 1.760000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.850000 1.425000 7.115000 1.760000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.955000 1.210000 5.680000 1.515000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.435000 1.195000 3.785000 1.525000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.965000 1.195000 3.265000 1.525000 ;
    END
  END C1
  PIN X
    ANTENNADIFFAREA  1.176000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.055000 0.790000 1.065000 ;
        RECT 0.085000 1.065000 1.690000 1.235000 ;
        RECT 0.085000 1.235000 0.360000 1.755000 ;
        RECT 0.085000 1.755000 2.025000 1.925000 ;
        RECT 0.600000 0.255000 0.790000 1.055000 ;
        RECT 0.975000 1.925000 1.165000 3.075000 ;
        RECT 1.460000 0.255000 1.690000 1.065000 ;
        RECT 1.835000 1.925000 2.025000 3.075000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 8.160000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 8.160000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.160000 0.085000 ;
      RECT 0.000000  3.245000 8.160000 3.415000 ;
      RECT 0.100000  0.085000 0.430000 0.885000 ;
      RECT 0.475000  2.095000 0.805000 3.245000 ;
      RECT 0.530000  1.405000 2.795000 1.585000 ;
      RECT 0.960000  0.085000 1.290000 0.895000 ;
      RECT 1.335000  2.105000 1.665000 3.245000 ;
      RECT 1.860000  0.085000 2.150000 1.105000 ;
      RECT 2.195000  1.585000 2.795000 1.705000 ;
      RECT 2.195000  1.705000 5.235000 1.875000 ;
      RECT 2.195000  2.045000 2.525000 3.245000 ;
      RECT 2.320000  0.765000 3.100000 1.015000 ;
      RECT 2.320000  1.015000 2.795000 1.405000 ;
      RECT 2.340000  0.255000 4.390000 0.435000 ;
      RECT 2.340000  0.435000 3.460000 0.595000 ;
      RECT 2.695000  1.875000 2.925000 3.075000 ;
      RECT 3.095000  2.045000 3.425000 3.245000 ;
      RECT 3.270000  0.595000 3.460000 1.025000 ;
      RECT 3.595000  1.875000 3.820000 3.075000 ;
      RECT 3.630000  0.615000 3.960000 0.855000 ;
      RECT 3.630000  0.855000 4.840000 0.870000 ;
      RECT 3.630000  0.870000 6.200000 1.025000 ;
      RECT 3.955000  1.025000 6.200000 1.040000 ;
      RECT 3.990000  2.045000 4.320000 3.245000 ;
      RECT 4.130000  0.435000 4.390000 0.685000 ;
      RECT 4.510000  2.045000 4.840000 2.905000 ;
      RECT 4.510000  2.905000 6.700000 3.075000 ;
      RECT 4.580000  0.255000 4.840000 0.855000 ;
      RECT 5.010000  0.085000 5.840000 0.700000 ;
      RECT 5.010000  1.875000 5.235000 2.735000 ;
      RECT 5.405000  1.705000 5.680000 2.905000 ;
      RECT 5.940000  1.930000 7.990000 2.100000 ;
      RECT 5.940000  2.100000 6.200000 2.735000 ;
      RECT 6.000000  1.040000 6.200000 1.085000 ;
      RECT 6.000000  1.085000 7.990000 1.255000 ;
      RECT 6.010000  0.255000 6.200000 0.870000 ;
      RECT 6.370000  0.085000 6.700000 0.915000 ;
      RECT 6.370000  2.270000 6.700000 2.905000 ;
      RECT 6.870000  0.255000 7.060000 1.085000 ;
      RECT 6.870000  2.100000 7.060000 3.075000 ;
      RECT 7.230000  0.085000 7.560000 0.915000 ;
      RECT 7.230000  2.270000 7.560000 3.245000 ;
      RECT 7.730000  0.255000 7.990000 1.085000 ;
      RECT 7.730000  2.100000 7.990000 3.075000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
  END
END sky130_fd_sc_lp__o311a_4
