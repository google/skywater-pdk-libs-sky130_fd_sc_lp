* File: sky130_fd_sc_lp__and4_4.spice
* Created: Wed Sep  2 09:32:59 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__and4_4.pex.spice"
.subckt sky130_fd_sc_lp__and4_4  VNB VPB A B C D VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* D	D
* C	C
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1009 A_141_47# N_A_M1009_g N_A_58_47#_M1009_s VNB NSHORT L=0.15 W=0.84
+ AD=0.0882 AS=0.2226 PD=1.05 PS=2.21 NRD=7.14 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75003.5 A=0.126 P=1.98 MULT=1
MM1003 A_213_47# N_B_M1003_g A_141_47# VNB NSHORT L=0.15 W=0.84 AD=0.1638
+ AS=0.0882 PD=1.23 PS=1.05 NRD=19.992 NRS=7.14 M=1 R=5.6 SA=75000.6 SB=75003.1
+ A=0.126 P=1.98 MULT=1
MM1008 A_321_47# N_C_M1008_g A_213_47# VNB NSHORT L=0.15 W=0.84 AD=0.1638
+ AS=0.1638 PD=1.23 PS=1.23 NRD=19.992 NRS=19.992 M=1 R=5.6 SA=75001.1
+ SB=75002.6 A=0.126 P=1.98 MULT=1
MM1015 N_VGND_M1015_d N_D_M1015_g A_321_47# VNB NSHORT L=0.15 W=0.84 AD=0.1785
+ AS=0.1638 PD=1.265 PS=1.23 NRD=8.568 NRS=19.992 M=1 R=5.6 SA=75001.6
+ SB=75002.1 A=0.126 P=1.98 MULT=1
MM1002 N_VGND_M1015_d N_A_58_47#_M1002_g N_X_M1002_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1785 AS=0.1176 PD=1.265 PS=1.12 NRD=12.132 NRS=0 M=1 R=5.6 SA=75002.2
+ SB=75001.5 A=0.126 P=1.98 MULT=1
MM1004 N_VGND_M1004_d N_A_58_47#_M1004_g N_X_M1002_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002.6
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1011 N_VGND_M1004_d N_A_58_47#_M1011_g N_X_M1011_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75003.1
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1014 N_VGND_M1014_d N_A_58_47#_M1014_g N_X_M1011_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75003.5
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1000 N_A_58_47#_M1000_d N_A_M1000_g N_VPWR_M1000_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75003.5 A=0.189 P=2.82 MULT=1
MM1007 N_VPWR_M1007_d N_B_M1007_g N_A_58_47#_M1000_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.2709 AS=0.1764 PD=1.69 PS=1.54 NRD=11.7215 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75003.1 A=0.189 P=2.82 MULT=1
MM1006 N_A_58_47#_M1006_d N_C_M1006_g N_VPWR_M1007_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.2709 PD=1.54 PS=1.69 NRD=0 NRS=11.7215 M=1 R=8.4 SA=75001.2
+ SB=75002.5 A=0.189 P=2.82 MULT=1
MM1012 N_VPWR_M1012_d N_D_M1012_g N_A_58_47#_M1006_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.26775 AS=0.1764 PD=1.685 PS=1.54 NRD=9.3772 NRS=0 M=1 R=8.4 SA=75001.6
+ SB=75002.1 A=0.189 P=2.82 MULT=1
MM1001 N_VPWR_M1012_d N_A_58_47#_M1001_g N_X_M1001_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.26775 AS=0.1764 PD=1.685 PS=1.54 NRD=13.2778 NRS=0 M=1 R=8.4 SA=75002.2
+ SB=75001.5 A=0.189 P=2.82 MULT=1
MM1005 N_VPWR_M1005_d N_A_58_47#_M1005_g N_X_M1001_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.6
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1010 N_VPWR_M1005_d N_A_58_47#_M1010_g N_X_M1010_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75003.1
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1013 N_VPWR_M1013_d N_A_58_47#_M1013_g N_X_M1010_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75003.5
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX16_noxref VNB VPB NWDIODE A=9.6607 P=14.09
*
.include "sky130_fd_sc_lp__and4_4.pxi.spice"
*
.ends
*
*
