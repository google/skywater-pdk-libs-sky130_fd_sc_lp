* File: sky130_fd_sc_lp__o31ai_0.spice
* Created: Wed Sep  2 10:25:06 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__o31ai_0.pex.spice"
.subckt sky130_fd_sc_lp__o31ai_0  VNB VPB A1 A2 A3 B1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B1	B1
* A3	A3
* A2	A2
* A1	A1
* VPB	VPB
* VNB	VNB
MM1006 N_A_138_65#_M1006_d N_A1_M1006_g N_VGND_M1006_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75001.9
+ A=0.063 P=1.14 MULT=1
MM1007 N_VGND_M1007_d N_A2_M1007_g N_A_138_65#_M1006_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0798 AS=0.0588 PD=0.8 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75001.5 A=0.063 P=1.14 MULT=1
MM1002 N_A_138_65#_M1002_d N_A3_M1002_g N_VGND_M1007_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0798 PD=0.7 PS=0.8 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.1
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1004 N_Y_M1004_d N_B1_M1004_g N_A_138_65#_M1002_d VNB NSHORT L=0.15 W=0.42
+ AD=0.2541 AS=0.0588 PD=2.05 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.6 SB=75000.5
+ A=0.063 P=1.14 MULT=1
MM1000 A_146_483# N_A1_M1000_g N_VPWR_M1000_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0768 AS=0.1696 PD=0.88 PS=1.81 NRD=19.9955 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75001.4 A=0.096 P=1.58 MULT=1
MM1001 A_224_483# N_A2_M1001_g A_146_483# VPB PHIGHVT L=0.15 W=0.64 AD=0.0768
+ AS=0.0768 PD=0.88 PS=0.88 NRD=19.9955 NRS=19.9955 M=1 R=4.26667 SA=75000.6
+ SB=75001 A=0.096 P=1.58 MULT=1
MM1005 N_Y_M1005_d N_A3_M1005_g A_224_483# VPB PHIGHVT L=0.15 W=0.64 AD=0.0896
+ AS=0.0768 PD=0.92 PS=0.88 NRD=0 NRS=19.9955 M=1 R=4.26667 SA=75001 SB=75000.6
+ A=0.096 P=1.58 MULT=1
MM1003 N_VPWR_M1003_d N_B1_M1003_g N_Y_M1005_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1696 AS=0.0896 PD=1.81 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667 SA=75001.4
+ SB=75000.2 A=0.096 P=1.58 MULT=1
DX8_noxref VNB VPB NWDIODE A=6.0799 P=10.25
c_35 VNB 0 1.95508e-19 $X=0 $Y=0
*
.include "sky130_fd_sc_lp__o31ai_0.pxi.spice"
*
.ends
*
*
