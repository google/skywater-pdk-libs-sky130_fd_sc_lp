* File: sky130_fd_sc_lp__sdfxtp_4.pex.spice
* Created: Fri Aug 28 11:30:57 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__SDFXTP_4%A_91_123# 1 2 9 13 16 17 21 22 27 31 32
c86 21 0 6.94633e-20 $X=2.215 $Y=2.13
r87 32 34 4.88247 $w=9.87e-07 $l=3.95e-07 $layer=LI1_cond $X=0.7 $Y=2.385
+ $X2=0.7 $Y2=2.78
r88 31 36 18.3619 $w=3.15e-07 $l=1.2e-07 $layer=POLY_cond $X=1.105 $Y=1.74
+ $X2=1.225 $Y2=1.74
r89 30 32 7.97264 $w=9.87e-07 $l=6.45e-07 $layer=LI1_cond $X=0.7 $Y=1.74 $X2=0.7
+ $Y2=2.385
r90 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.105
+ $Y=1.74 $X2=1.105 $Y2=1.74
r91 24 27 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=0.22 $Y=0.8 $X2=0.58
+ $Y2=0.8
r92 22 39 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.215 $Y=2.13
+ $X2=2.215 $Y2=2.295
r93 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.215
+ $Y=2.13 $X2=2.215 $Y2=2.13
r94 19 21 7.5352 $w=2.58e-07 $l=1.7e-07 $layer=LI1_cond $X=2.18 $Y=2.3 $X2=2.18
+ $Y2=2.13
r95 18 32 11.6346 $w=1.7e-07 $l=5.7e-07 $layer=LI1_cond $X=1.27 $Y=2.385 $X2=0.7
+ $Y2=2.385
r96 17 19 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=2.05 $Y=2.385
+ $X2=2.18 $Y2=2.3
r97 17 18 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=2.05 $Y=2.385
+ $X2=1.27 $Y2=2.385
r98 16 30 11.3536 $w=9.87e-07 $l=5.20769e-07 $layer=LI1_cond $X=0.22 $Y=1.655
+ $X2=0.7 $Y2=1.74
r99 15 24 4.28565 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=0.22 $Y=0.965
+ $X2=0.22 $Y2=0.8
r100 15 16 42.5152 $w=1.78e-07 $l=6.9e-07 $layer=LI1_cond $X=0.22 $Y=0.965
+ $X2=0.22 $Y2=1.655
r101 13 39 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.195 $Y=2.775
+ $X2=2.195 $Y2=2.295
r102 7 36 20.1192 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.225 $Y=1.575
+ $X2=1.225 $Y2=1.74
r103 7 9 384.574 $w=1.5e-07 $l=7.5e-07 $layer=POLY_cond $X=1.225 $Y=1.575
+ $X2=1.225 $Y2=0.825
r104 2 34 600 $w=1.7e-07 $l=3.82426e-07 $layer=licon1_PDIFF $count=1 $X=0.635
+ $Y=2.455 $X2=0.76 $Y2=2.78
r105 1 27 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=0.455
+ $Y=0.615 $X2=0.58 $Y2=0.8
.ends

.subckt PM_SKY130_FD_SC_LP__SDFXTP_4%D 3 6 9 10 11 12 13 14 15 16 23
c52 12 0 2.3436e-19 $X=1.68 $Y=0.555
c53 9 0 1.28145e-19 $X=1.675 $Y=1.145
r54 15 16 16.0907 $w=2.63e-07 $l=3.7e-07 $layer=LI1_cond $X=1.642 $Y=1.665
+ $X2=1.642 $Y2=2.035
r55 14 15 16.0907 $w=2.63e-07 $l=3.7e-07 $layer=LI1_cond $X=1.642 $Y=1.295
+ $X2=1.642 $Y2=1.665
r56 14 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.675
+ $Y=1.31 $X2=1.675 $Y2=1.31
r57 13 14 16.0907 $w=2.63e-07 $l=3.7e-07 $layer=LI1_cond $X=1.642 $Y=0.925
+ $X2=1.642 $Y2=1.295
r58 12 13 16.0907 $w=2.63e-07 $l=3.7e-07 $layer=LI1_cond $X=1.642 $Y=0.555
+ $X2=1.642 $Y2=0.925
r59 10 23 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.675 $Y=1.65
+ $X2=1.675 $Y2=1.31
r60 10 11 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.675 $Y=1.65
+ $X2=1.675 $Y2=1.815
r61 9 23 40.425 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.675 $Y=1.145
+ $X2=1.675 $Y2=1.31
r62 6 11 492.255 $w=1.5e-07 $l=9.6e-07 $layer=POLY_cond $X=1.765 $Y=2.775
+ $X2=1.765 $Y2=1.815
r63 3 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.72 $Y=0.825 $X2=1.72
+ $Y2=1.145
.ends

.subckt PM_SKY130_FD_SC_LP__SDFXTP_4%SCE 2 3 4 8 9 10 13 15 19 23 25 26 27 32
c69 15 0 1.3975e-19 $X=1.33 $Y=2.19
c70 8 0 9.46099e-20 $X=0.795 $Y=0.825
r71 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.565
+ $Y=1.31 $X2=0.565 $Y2=1.31
r72 30 32 15.7174 $w=2.76e-07 $l=9e-08 $layer=POLY_cond $X=0.475 $Y=1.31
+ $X2=0.565 $Y2=1.31
r73 26 27 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=0.72 $Y=1.31 $X2=1.2
+ $Y2=1.31
r74 26 33 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=0.72 $Y=1.31
+ $X2=0.565 $Y2=1.31
r75 21 23 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=2.34 $Y=0.275
+ $X2=2.34 $Y2=0.825
r76 17 19 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=1.405 $Y=2.265
+ $X2=1.405 $Y2=2.775
r77 16 25 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.05 $Y=2.19
+ $X2=0.975 $Y2=2.19
r78 15 17 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.33 $Y=2.19
+ $X2=1.405 $Y2=2.265
r79 15 16 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=1.33 $Y=2.19
+ $X2=1.05 $Y2=2.19
r80 11 25 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.975 $Y=2.265
+ $X2=0.975 $Y2=2.19
r81 11 13 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=0.975 $Y=2.265
+ $X2=0.975 $Y2=2.775
r82 9 21 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.265 $Y=0.2
+ $X2=2.34 $Y2=0.275
r83 9 10 715.309 $w=1.5e-07 $l=1.395e-06 $layer=POLY_cond $X=2.265 $Y=0.2
+ $X2=0.87 $Y2=0.2
r84 6 32 40.1667 $w=2.76e-07 $l=3.01413e-07 $layer=POLY_cond $X=0.795 $Y=1.145
+ $X2=0.565 $Y2=1.31
r85 6 8 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.795 $Y=1.145
+ $X2=0.795 $Y2=0.825
r86 5 10 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.795 $Y=0.275
+ $X2=0.87 $Y2=0.2
r87 5 8 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=0.795 $Y=0.275
+ $X2=0.795 $Y2=0.825
r88 3 25 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.9 $Y=2.19 $X2=0.975
+ $Y2=2.19
r89 3 4 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=0.9 $Y=2.19 $X2=0.55
+ $Y2=2.19
r90 2 4 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.475 $Y=2.115
+ $X2=0.55 $Y2=2.19
r91 1 30 17.0164 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=1.475
+ $X2=0.475 $Y2=1.31
r92 1 2 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=0.475 $Y=1.475
+ $X2=0.475 $Y2=2.115
.ends

.subckt PM_SKY130_FD_SC_LP__SDFXTP_4%SCD 3 7 9 10 14
c44 7 0 1.26524e-19 $X=2.7 $Y=0.825
r45 14 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.61 $Y=1.56
+ $X2=2.61 $Y2=1.725
r46 14 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.61 $Y=1.56
+ $X2=2.61 $Y2=1.395
r47 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.61
+ $Y=1.56 $X2=2.61 $Y2=1.56
r48 10 15 0.864332 $w=3.98e-07 $l=3e-08 $layer=LI1_cond $X=2.64 $Y=1.595
+ $X2=2.61 $Y2=1.595
r49 9 15 12.965 $w=3.98e-07 $l=4.5e-07 $layer=LI1_cond $X=2.16 $Y=1.595 $X2=2.61
+ $Y2=1.595
r50 7 16 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=2.7 $Y=0.825 $X2=2.7
+ $Y2=1.395
r51 3 17 538.404 $w=1.5e-07 $l=1.05e-06 $layer=POLY_cond $X=2.665 $Y=2.775
+ $X2=2.665 $Y2=1.725
.ends

.subckt PM_SKY130_FD_SC_LP__SDFXTP_4%CLK 3 7 9 10 11 16
c45 16 0 1.34012e-19 $X=3.34 $Y=1.375
c46 9 0 1.26524e-19 $X=3.6 $Y=1.295
r47 16 19 88.9594 $w=4.5e-07 $l=5.05e-07 $layer=POLY_cond $X=3.28 $Y=1.375
+ $X2=3.28 $Y2=1.88
r48 16 18 46.9389 $w=4.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.28 $Y=1.375
+ $X2=3.28 $Y2=1.21
r49 16 17 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.34
+ $Y=1.375 $X2=3.34 $Y2=1.375
r50 10 11 9.691 $w=4.38e-07 $l=3.7e-07 $layer=LI1_cond $X=3.475 $Y=1.665
+ $X2=3.475 $Y2=2.035
r51 10 17 7.59565 $w=4.38e-07 $l=2.9e-07 $layer=LI1_cond $X=3.475 $Y=1.665
+ $X2=3.475 $Y2=1.375
r52 9 17 2.09535 $w=4.38e-07 $l=8e-08 $layer=LI1_cond $X=3.475 $Y=1.295
+ $X2=3.475 $Y2=1.375
r53 7 19 458.926 $w=1.5e-07 $l=8.95e-07 $layer=POLY_cond $X=3.13 $Y=2.775
+ $X2=3.13 $Y2=1.88
r54 3 18 197.415 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=3.13 $Y=0.825
+ $X2=3.13 $Y2=1.21
.ends

.subckt PM_SKY130_FD_SC_LP__SDFXTP_4%A_641_123# 1 2 9 11 12 14 17 21 25 29 32 33
+ 34 37 39 40 43 47 49 50 52 53 54 56 57 60 61 64 67 68 72 75 76 81 83 88 91 93
c240 91 0 3.05834e-19 $X=7.6 $Y=1.93
c241 88 0 4.17627e-20 $X=7.435 $Y=1.92
c242 83 0 1.27388e-19 $X=5.96 $Y=2.72
c243 81 0 5.18384e-21 $X=5.96 $Y=1.68
c244 64 0 2.72499e-20 $X=7.89 $Y=1.825
c245 60 0 4.05543e-20 $X=7.515 $Y=2.635
c246 50 0 4.40926e-20 $X=4.082 $Y=2.3
c247 21 0 3.05678e-20 $X=5.92 $Y=2.455
c248 17 0 2.38548e-19 $X=5.19 $Y=0.835
r249 92 93 8.67109 $w=3.58e-07 $l=1.7e-07 $layer=LI1_cond $X=8.07 $Y=1.345
+ $X2=8.07 $Y2=1.515
r250 90 91 4.74668 $w=2.08e-07 $l=8.5e-08 $layer=LI1_cond $X=7.515 $Y=1.93
+ $X2=7.6 $Y2=1.93
r251 88 96 23.6063 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=7.435 $Y=1.92
+ $X2=7.3 $Y2=1.92
r252 87 90 4.22511 $w=2.08e-07 $l=8e-08 $layer=LI1_cond $X=7.435 $Y=1.93
+ $X2=7.515 $Y2=1.93
r253 87 88 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.435
+ $Y=1.92 $X2=7.435 $Y2=1.92
r254 83 84 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=5.96 $Y=2.72
+ $X2=5.96 $Y2=2.98
r255 78 81 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=5.83 $Y=1.68
+ $X2=5.96 $Y2=1.68
r256 78 79 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.83
+ $Y=1.68 $X2=5.83 $Y2=1.68
r257 74 75 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.085
+ $Y=0.95 $X2=4.085 $Y2=0.95
r258 70 72 11.39 $w=2.41e-07 $l=2.25e-07 $layer=LI1_cond $X=3.345 $Y=2.385
+ $X2=3.345 $Y2=2.61
r259 68 101 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.25 $Y=1.02
+ $X2=8.25 $Y2=0.855
r260 67 92 10.404 $w=3.58e-07 $l=3.25e-07 $layer=LI1_cond $X=8.155 $Y=1.02
+ $X2=8.155 $Y2=1.345
r261 67 68 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.25
+ $Y=1.02 $X2=8.25 $Y2=1.02
r262 64 93 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=7.89 $Y=1.825
+ $X2=7.89 $Y2=1.515
r263 61 64 6.82373 $w=1.8e-07 $l=1.25499e-07 $layer=LI1_cond $X=7.805 $Y=1.915
+ $X2=7.89 $Y2=1.825
r264 61 91 12.6313 $w=1.78e-07 $l=2.05e-07 $layer=LI1_cond $X=7.805 $Y=1.915
+ $X2=7.6 $Y2=1.915
r265 59 90 1.9771 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=7.515 $Y=2.035
+ $X2=7.515 $Y2=1.93
r266 59 60 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=7.515 $Y=2.035
+ $X2=7.515 $Y2=2.635
r267 58 83 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.045 $Y=2.72
+ $X2=5.96 $Y2=2.72
r268 57 60 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.43 $Y=2.72
+ $X2=7.515 $Y2=2.635
r269 57 58 90.3583 $w=1.68e-07 $l=1.385e-06 $layer=LI1_cond $X=7.43 $Y=2.72
+ $X2=6.045 $Y2=2.72
r270 56 83 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=5.96 $Y=2.635
+ $X2=5.96 $Y2=2.72
r271 55 81 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.96 $Y=1.845
+ $X2=5.96 $Y2=1.68
r272 55 56 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=5.96 $Y=1.845
+ $X2=5.96 $Y2=2.635
r273 53 84 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.875 $Y=2.98
+ $X2=5.96 $Y2=2.98
r274 53 54 102.754 $w=1.68e-07 $l=1.575e-06 $layer=LI1_cond $X=5.875 $Y=2.98
+ $X2=4.3 $Y2=2.98
r275 52 54 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.215 $Y=2.895
+ $X2=4.3 $Y2=2.98
r276 51 76 3.12539 $w=3.02e-07 $l=1.70276e-07 $layer=LI1_cond $X=4.215 $Y=2.47
+ $X2=4.082 $Y2=2.385
r277 51 52 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=4.215 $Y=2.47
+ $X2=4.215 $Y2=2.895
r278 50 76 3.12539 $w=3.02e-07 $l=8.5e-08 $layer=LI1_cond $X=4.082 $Y=2.3
+ $X2=4.082 $Y2=2.385
r279 49 74 2.69035 $w=4.35e-07 $l=1.18e-07 $layer=LI1_cond $X=4.082 $Y=1.02
+ $X2=4.082 $Y2=0.902
r280 49 50 33.911 $w=4.33e-07 $l=1.28e-06 $layer=LI1_cond $X=4.082 $Y=1.02
+ $X2=4.082 $Y2=2.3
r281 48 70 2.78154 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.51 $Y=2.385
+ $X2=3.345 $Y2=2.385
r282 47 76 3.47949 $w=1.7e-07 $l=2.17e-07 $layer=LI1_cond $X=3.865 $Y=2.385
+ $X2=4.082 $Y2=2.385
r283 47 48 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=3.865 $Y=2.385
+ $X2=3.51 $Y2=2.385
r284 43 74 4.9475 $w=2.35e-07 $l=2.17e-07 $layer=LI1_cond $X=3.865 $Y=0.902
+ $X2=4.082 $Y2=0.902
r285 43 45 20.8421 $w=2.33e-07 $l=4.25e-07 $layer=LI1_cond $X=3.865 $Y=0.902
+ $X2=3.44 $Y2=0.902
r286 40 79 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=5.845 $Y=1.68
+ $X2=5.83 $Y2=1.68
r287 39 79 98.7966 $w=3.3e-07 $l=5.65e-07 $layer=POLY_cond $X=5.265 $Y=1.68
+ $X2=5.83 $Y2=1.68
r288 35 37 89.734 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=4.175 $Y=2.22
+ $X2=4.35 $Y2=2.22
r289 33 75 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=4.085 $Y=1.29
+ $X2=4.085 $Y2=0.95
r290 33 34 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.085 $Y=1.29
+ $X2=4.085 $Y2=1.455
r291 32 75 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.085 $Y=0.785
+ $X2=4.085 $Y2=0.95
r292 29 101 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=8.275 $Y=0.515
+ $X2=8.275 $Y2=0.855
r293 23 96 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.3 $Y=2.085
+ $X2=7.3 $Y2=1.92
r294 23 25 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=7.3 $Y=2.085
+ $X2=7.3 $Y2=2.665
r295 19 40 32.1775 $w=3.3e-07 $l=1.98997e-07 $layer=POLY_cond $X=5.92 $Y=1.845
+ $X2=5.845 $Y2=1.68
r296 19 21 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=5.92 $Y=1.845
+ $X2=5.92 $Y2=2.455
r297 15 39 32.1775 $w=3.3e-07 $l=1.98997e-07 $layer=POLY_cond $X=5.19 $Y=1.515
+ $X2=5.265 $Y2=1.68
r298 15 17 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=5.19 $Y=1.515
+ $X2=5.19 $Y2=0.835
r299 12 37 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.35 $Y=2.295
+ $X2=4.35 $Y2=2.22
r300 12 14 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=4.35 $Y=2.295
+ $X2=4.35 $Y2=2.725
r301 11 35 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.175 $Y=2.145
+ $X2=4.175 $Y2=2.22
r302 11 34 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=4.175 $Y=2.145
+ $X2=4.175 $Y2=1.455
r303 9 32 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=4.175 $Y=0.465
+ $X2=4.175 $Y2=0.785
r304 2 72 300 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_PDIFF $count=2 $X=3.205
+ $Y=2.455 $X2=3.345 $Y2=2.61
r305 1 45 182 $w=1.7e-07 $l=3.745e-07 $layer=licon1_NDIFF $count=1 $X=3.205
+ $Y=0.615 $X2=3.44 $Y2=0.89
.ends

.subckt PM_SKY130_FD_SC_LP__SDFXTP_4%A_850_51# 1 2 8 9 10 11 13 14 16 19 21 22
+ 23 26 29 32 34 35 39 43 44 46 50 51 57 58 63 72
c175 39 0 8.05806e-20 $X=5.72 $Y=0.375
c176 26 0 1.10981e-19 $X=8.08 $Y=2.745
c177 21 0 1.52416e-19 $X=7.77 $Y=1.395
c178 14 0 2.07351e-19 $X=5.64 $Y=0.515
c179 11 0 1.28676e-19 $X=5.3 $Y=2.205
c180 10 0 4.40926e-20 $X=4.82 $Y=2.13
r181 63 65 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=6.85 $Y=0.34 $X2=6.85
+ $Y2=0.64
r182 56 57 4.3334 $w=3.38e-07 $l=9.8e-08 $layer=LI1_cond $X=4.567 $Y=0.425
+ $X2=4.665 $Y2=0.425
r183 54 56 5.99948 $w=3.38e-07 $l=1.77e-07 $layer=LI1_cond $X=4.39 $Y=0.425
+ $X2=4.567 $Y2=0.425
r184 51 73 46.3065 $w=3.4e-07 $l=1.65e-07 $layer=POLY_cond $X=7.705 $Y=1
+ $X2=7.705 $Y2=1.165
r185 51 72 46.3065 $w=3.4e-07 $l=1.65e-07 $layer=POLY_cond $X=7.705 $Y=1
+ $X2=7.705 $Y2=0.835
r186 50 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.71 $Y=1
+ $X2=7.71 $Y2=1
r187 48 50 35.4293 $w=1.78e-07 $l=5.75e-07 $layer=LI1_cond $X=7.705 $Y=0.425
+ $X2=7.705 $Y2=1
r188 47 63 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.935 $Y=0.34
+ $X2=6.85 $Y2=0.34
r189 46 48 6.82373 $w=1.7e-07 $l=1.25499e-07 $layer=LI1_cond $X=7.615 $Y=0.34
+ $X2=7.705 $Y2=0.425
r190 46 47 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=7.615 $Y=0.34
+ $X2=6.935 $Y2=0.34
r191 45 61 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.89 $Y=0.64
+ $X2=5.805 $Y2=0.64
r192 44 65 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.765 $Y=0.64
+ $X2=6.85 $Y2=0.64
r193 44 45 57.0856 $w=1.68e-07 $l=8.75e-07 $layer=LI1_cond $X=6.765 $Y=0.64
+ $X2=5.89 $Y2=0.64
r194 42 57 46.818 $w=2.38e-07 $l=9.75e-07 $layer=LI1_cond $X=5.64 $Y=0.375
+ $X2=4.665 $Y2=0.375
r195 42 43 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.64
+ $Y=0.35 $X2=5.64 $Y2=0.35
r196 39 61 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=5.805 $Y=0.375
+ $X2=5.805 $Y2=0.64
r197 39 42 3.84148 $w=2.38e-07 $l=8e-08 $layer=LI1_cond $X=5.72 $Y=0.375
+ $X2=5.64 $Y2=0.375
r198 34 37 47.7441 $w=2.78e-07 $l=1.16e-06 $layer=LI1_cond $X=4.61 $Y=1.4
+ $X2=4.61 $Y2=2.56
r199 34 35 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.655
+ $Y=1.4 $X2=4.655 $Y2=1.4
r200 32 58 6.83623 $w=2.78e-07 $l=1.4e-07 $layer=LI1_cond $X=4.61 $Y=1.375
+ $X2=4.61 $Y2=1.235
r201 32 34 1.02897 $w=2.78e-07 $l=2.5e-08 $layer=LI1_cond $X=4.61 $Y=1.375
+ $X2=4.61 $Y2=1.4
r202 30 56 4.00821 $w=1.95e-07 $l=1.7e-07 $layer=LI1_cond $X=4.567 $Y=0.595
+ $X2=4.567 $Y2=0.425
r203 30 58 36.4009 $w=1.93e-07 $l=6.4e-07 $layer=LI1_cond $X=4.567 $Y=0.595
+ $X2=4.567 $Y2=1.235
r204 28 35 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=4.655 $Y=1.74
+ $X2=4.655 $Y2=1.4
r205 28 29 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.655 $Y=1.74
+ $X2=4.655 $Y2=1.905
r206 24 26 615.319 $w=1.5e-07 $l=1.2e-06 $layer=POLY_cond $X=8.08 $Y=1.545
+ $X2=8.08 $Y2=2.745
r207 22 24 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.005 $Y=1.47
+ $X2=8.08 $Y2=1.545
r208 22 23 82.0426 $w=1.5e-07 $l=1.6e-07 $layer=POLY_cond $X=8.005 $Y=1.47
+ $X2=7.845 $Y2=1.47
r209 21 23 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.77 $Y=1.395
+ $X2=7.845 $Y2=1.47
r210 21 73 117.936 $w=1.5e-07 $l=2.3e-07 $layer=POLY_cond $X=7.77 $Y=1.395
+ $X2=7.77 $Y2=1.165
r211 19 72 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=7.61 $Y=0.515
+ $X2=7.61 $Y2=0.835
r212 14 43 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.64 $Y=0.515
+ $X2=5.64 $Y2=0.35
r213 14 16 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=5.64 $Y=0.515
+ $X2=5.64 $Y2=0.835
r214 11 13 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=5.3 $Y=2.205
+ $X2=5.3 $Y2=2.525
r215 9 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.225 $Y=2.13
+ $X2=5.3 $Y2=2.205
r216 9 10 207.67 $w=1.5e-07 $l=4.05e-07 $layer=POLY_cond $X=5.225 $Y=2.13
+ $X2=4.82 $Y2=2.13
r217 8 10 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.745 $Y=2.055
+ $X2=4.82 $Y2=2.13
r218 8 29 76.9149 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=4.745 $Y=2.055
+ $X2=4.745 $Y2=1.905
r219 2 37 600 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_PDIFF $count=1 $X=4.425
+ $Y=2.405 $X2=4.565 $Y2=2.56
r220 1 54 182 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=1 $X=4.25
+ $Y=0.255 $X2=4.39 $Y2=0.43
.ends

.subckt PM_SKY130_FD_SC_LP__SDFXTP_4%A_1203_99# 1 2 7 9 10 11 14 16 17 22 25 31
c66 14 0 1.27388e-19 $X=6.28 $Y=2.455
r67 31 33 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=7.28 $Y=0.72
+ $X2=7.28 $Y2=0.885
r68 25 33 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=7.36 $Y=1.475
+ $X2=7.36 $Y2=0.885
r69 22 25 6.82373 $w=1.8e-07 $l=1.25499e-07 $layer=LI1_cond $X=7.275 $Y=1.565
+ $X2=7.36 $Y2=1.475
r70 22 23 11.399 $w=1.78e-07 $l=1.85e-07 $layer=LI1_cond $X=7.275 $Y=1.565
+ $X2=7.09 $Y2=1.565
r71 17 29 34.2406 $w=2.12e-07 $l=5.95e-07 $layer=LI1_cond $X=7.085 $Y=1.775
+ $X2=7.085 $Y2=2.37
r72 17 23 12.0849 $w=2.12e-07 $l=2.1e-07 $layer=LI1_cond $X=7.085 $Y=1.775
+ $X2=7.085 $Y2=1.565
r73 17 19 10.5654 $w=5.98e-07 $l=5.3e-07 $layer=LI1_cond $X=6.92 $Y=1.775
+ $X2=6.39 $Y2=1.775
r74 14 16 194.851 $w=1.5e-07 $l=3.8e-07 $layer=POLY_cond $X=6.28 $Y=2.455
+ $X2=6.28 $Y2=2.075
r75 11 16 48.0802 $w=3.5e-07 $l=1.75e-07 $layer=POLY_cond $X=6.38 $Y=1.9
+ $X2=6.38 $Y2=2.075
r76 10 19 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.39
+ $Y=1.57 $X2=6.39 $Y2=1.57
r77 10 11 52.7581 $w=3.5e-07 $l=3.2e-07 $layer=POLY_cond $X=6.38 $Y=1.58
+ $X2=6.38 $Y2=1.9
r78 7 10 59.4809 $w=2.35e-07 $l=5.51249e-07 $layer=POLY_cond $X=6.09 $Y=1.155
+ $X2=6.38 $Y2=1.58
r79 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=6.09 $Y=1.155 $X2=6.09
+ $Y2=0.835
r80 2 29 600 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=6.945
+ $Y=2.245 $X2=7.085 $Y2=2.37
r81 1 31 182 $w=1.7e-07 $l=4.79922e-07 $layer=licon1_NDIFF $count=1 $X=7.14
+ $Y=0.305 $X2=7.28 $Y2=0.72
.ends

.subckt PM_SKY130_FD_SC_LP__SDFXTP_4%A_1053_125# 1 2 9 11 13 16 22 25 27 28 33
c71 16 0 2.98067e-19 $X=5.425 $Y=0.83
c72 9 0 2.35407e-19 $X=6.87 $Y=2.665
r73 27 28 11.1425 $w=3.43e-07 $l=2.55e-07 $layer=LI1_cond $X=5.532 $Y=2.48
+ $X2=5.532 $Y2=2.225
r74 23 33 23.6063 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=6.93 $Y=1.22
+ $X2=7.065 $Y2=1.22
r75 23 30 10.4917 $w=3.3e-07 $l=6e-08 $layer=POLY_cond $X=6.93 $Y=1.22 $X2=6.87
+ $Y2=1.22
r76 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.93
+ $Y=1.22 $X2=6.93 $Y2=1.22
r77 20 25 0.638687 $w=2.5e-07 $l=2.85745e-07 $layer=LI1_cond $X=5.55 $Y=1.18
+ $X2=5.32 $Y2=1.055
r78 20 22 63.6149 $w=2.48e-07 $l=1.38e-06 $layer=LI1_cond $X=5.55 $Y=1.18
+ $X2=6.93 $Y2=1.18
r79 18 25 6.0735 $w=2.05e-07 $l=3.08221e-07 $layer=LI1_cond $X=5.45 $Y=1.305
+ $X2=5.32 $Y2=1.055
r80 18 28 56.6869 $w=1.78e-07 $l=9.2e-07 $layer=LI1_cond $X=5.45 $Y=1.305
+ $X2=5.45 $Y2=2.225
r81 14 25 6.0735 $w=2.05e-07 $l=1.15e-07 $layer=LI1_cond $X=5.435 $Y=1.055
+ $X2=5.32 $Y2=1.055
r82 14 16 11.2739 $w=2.28e-07 $l=2.25e-07 $layer=LI1_cond $X=5.435 $Y=1.055
+ $X2=5.435 $Y2=0.83
r83 11 33 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.065 $Y=1.055
+ $X2=7.065 $Y2=1.22
r84 11 13 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=7.065 $Y=1.055
+ $X2=7.065 $Y2=0.625
r85 7 30 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.87 $Y=1.385
+ $X2=6.87 $Y2=1.22
r86 7 9 656.34 $w=1.5e-07 $l=1.28e-06 $layer=POLY_cond $X=6.87 $Y=1.385 $X2=6.87
+ $Y2=2.665
r87 2 27 600 $w=1.7e-07 $l=3.06594e-07 $layer=licon1_PDIFF $count=1 $X=5.375
+ $Y=2.315 $X2=5.61 $Y2=2.48
r88 1 16 182 $w=1.7e-07 $l=2.73542e-07 $layer=licon1_NDIFF $count=1 $X=5.265
+ $Y=0.625 $X2=5.425 $Y2=0.83
.ends

.subckt PM_SKY130_FD_SC_LP__SDFXTP_4%A_1673_409# 1 2 9 13 15 17 20 22 24 27 29
+ 31 34 36 38 41 43 47 51 54 58 64 67 73 74 75 76 82 88
c141 76 0 1.76576e-19 $X=10.15 $Y=1.37
c142 34 0 1.55372e-19 $X=11.085 $Y=2.465
c143 15 0 1.75356e-19 $X=10.225 $Y=1.205
c144 13 0 2.72499e-20 $X=8.7 $Y=0.515
r145 87 88 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=11.085 $Y=1.37
+ $X2=11.515 $Y2=1.37
r146 84 85 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=10.225 $Y=1.37
+ $X2=10.655 $Y2=1.37
r147 76 84 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=10.15 $Y=1.37
+ $X2=10.225 $Y2=1.37
r148 71 82 19.2347 $w=3.3e-07 $l=1.1e-07 $layer=POLY_cond $X=8.59 $Y=2.21
+ $X2=8.7 $Y2=2.21
r149 71 79 26.2292 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=8.59 $Y=2.21
+ $X2=8.44 $Y2=2.21
r150 70 71 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.59
+ $Y=2.21 $X2=8.59 $Y2=2.21
r151 67 70 4.0085 $w=2.28e-07 $l=8e-08 $layer=LI1_cond $X=8.61 $Y=2.13 $X2=8.61
+ $Y2=2.21
r152 65 87 41.0924 $w=3.3e-07 $l=2.35e-07 $layer=POLY_cond $X=10.85 $Y=1.37
+ $X2=11.085 $Y2=1.37
r153 65 85 34.0979 $w=3.3e-07 $l=1.95e-07 $layer=POLY_cond $X=10.85 $Y=1.37
+ $X2=10.655 $Y2=1.37
r154 64 65 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=10.85
+ $Y=1.37 $X2=10.85 $Y2=1.37
r155 62 76 55.9556 $w=3.3e-07 $l=3.2e-07 $layer=POLY_cond $X=9.83 $Y=1.37
+ $X2=10.15 $Y2=1.37
r156 61 64 56.5636 $w=1.98e-07 $l=1.02e-06 $layer=LI1_cond $X=9.83 $Y=1.385
+ $X2=10.85 $Y2=1.385
r157 61 62 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=9.83
+ $Y=1.37 $X2=9.83 $Y2=1.37
r158 59 75 1.25155 $w=2e-07 $l=1e-07 $layer=LI1_cond $X=9.605 $Y=1.385 $X2=9.505
+ $Y2=1.385
r159 59 61 12.4773 $w=1.98e-07 $l=2.25e-07 $layer=LI1_cond $X=9.605 $Y=1.385
+ $X2=9.83 $Y2=1.385
r160 56 74 4.60183 $w=1.95e-07 $l=8.74643e-08 $layer=LI1_cond $X=9.5 $Y=2.045
+ $X2=9.495 $Y2=2.13
r161 56 58 10.799 $w=1.88e-07 $l=1.85e-07 $layer=LI1_cond $X=9.5 $Y=2.045
+ $X2=9.5 $Y2=1.86
r162 55 75 5.27577 $w=1.95e-07 $l=1.0247e-07 $layer=LI1_cond $X=9.5 $Y=1.485
+ $X2=9.505 $Y2=1.385
r163 55 58 21.89 $w=1.88e-07 $l=3.75e-07 $layer=LI1_cond $X=9.5 $Y=1.485 $X2=9.5
+ $Y2=1.86
r164 54 75 5.27577 $w=1.95e-07 $l=1e-07 $layer=LI1_cond $X=9.505 $Y=1.285
+ $X2=9.505 $Y2=1.385
r165 54 73 15.5273 $w=1.98e-07 $l=2.8e-07 $layer=LI1_cond $X=9.505 $Y=1.285
+ $X2=9.505 $Y2=1.005
r166 49 74 4.60183 $w=1.95e-07 $l=8.5e-08 $layer=LI1_cond $X=9.495 $Y=2.215
+ $X2=9.495 $Y2=2.13
r167 49 51 6.65455 $w=1.98e-07 $l=1.2e-07 $layer=LI1_cond $X=9.495 $Y=2.215
+ $X2=9.495 $Y2=2.335
r168 45 73 6.4054 $w=2.58e-07 $l=1.3e-07 $layer=LI1_cond $X=9.475 $Y=0.875
+ $X2=9.475 $Y2=1.005
r169 45 47 20.1678 $w=2.58e-07 $l=4.55e-07 $layer=LI1_cond $X=9.475 $Y=0.875
+ $X2=9.475 $Y2=0.42
r170 44 67 2.50919 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=8.725 $Y=2.13
+ $X2=8.61 $Y2=2.13
r171 43 74 1.84097 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=9.395 $Y=2.13
+ $X2=9.495 $Y2=2.13
r172 43 44 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=9.395 $Y=2.13
+ $X2=8.725 $Y2=2.13
r173 39 88 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=11.515 $Y=1.535
+ $X2=11.515 $Y2=1.37
r174 39 41 476.872 $w=1.5e-07 $l=9.3e-07 $layer=POLY_cond $X=11.515 $Y=1.535
+ $X2=11.515 $Y2=2.465
r175 36 88 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=11.515 $Y=1.205
+ $X2=11.515 $Y2=1.37
r176 36 38 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=11.515 $Y=1.205
+ $X2=11.515 $Y2=0.675
r177 32 87 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=11.085 $Y=1.535
+ $X2=11.085 $Y2=1.37
r178 32 34 476.872 $w=1.5e-07 $l=9.3e-07 $layer=POLY_cond $X=11.085 $Y=1.535
+ $X2=11.085 $Y2=2.465
r179 29 87 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=11.085 $Y=1.205
+ $X2=11.085 $Y2=1.37
r180 29 31 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=11.085 $Y=1.205
+ $X2=11.085 $Y2=0.675
r181 25 85 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.655 $Y=1.535
+ $X2=10.655 $Y2=1.37
r182 25 27 476.872 $w=1.5e-07 $l=9.3e-07 $layer=POLY_cond $X=10.655 $Y=1.535
+ $X2=10.655 $Y2=2.465
r183 22 85 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.655 $Y=1.205
+ $X2=10.655 $Y2=1.37
r184 22 24 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=10.655 $Y=1.205
+ $X2=10.655 $Y2=0.675
r185 18 84 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.225 $Y=1.535
+ $X2=10.225 $Y2=1.37
r186 18 20 476.872 $w=1.5e-07 $l=9.3e-07 $layer=POLY_cond $X=10.225 $Y=1.535
+ $X2=10.225 $Y2=2.465
r187 15 84 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.225 $Y=1.205
+ $X2=10.225 $Y2=1.37
r188 15 17 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=10.225 $Y=1.205
+ $X2=10.225 $Y2=0.675
r189 11 82 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.7 $Y=2.045
+ $X2=8.7 $Y2=2.21
r190 11 13 784.532 $w=1.5e-07 $l=1.53e-06 $layer=POLY_cond $X=8.7 $Y=2.045
+ $X2=8.7 $Y2=0.515
r191 7 79 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.44 $Y=2.375
+ $X2=8.44 $Y2=2.21
r192 7 9 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=8.44 $Y=2.375
+ $X2=8.44 $Y2=2.745
r193 2 58 600 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_PDIFF $count=1 $X=9.35
+ $Y=1.695 $X2=9.49 $Y2=1.86
r194 2 51 300 $w=1.7e-07 $l=7.06541e-07 $layer=licon1_PDIFF $count=2 $X=9.35
+ $Y=1.695 $X2=9.49 $Y2=2.335
r195 1 47 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=9.3
+ $Y=0.235 $X2=9.44 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__SDFXTP_4%A_1475_449# 1 2 9 12 14 18 23 24 25 27 29
+ 32 33 35 37
c96 35 0 1.52416e-19 $X=8.6 $Y=1.35
c97 32 0 1.76576e-19 $X=9.15 $Y=1.35
c98 25 0 4.17627e-20 $X=8.325 $Y=1.78
r99 33 38 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=9.167 $Y=1.35
+ $X2=9.167 $Y2=1.515
r100 33 37 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=9.167 $Y=1.35
+ $X2=9.167 $Y2=1.185
r101 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.15
+ $Y=1.35 $X2=9.15 $Y2=1.35
r102 30 35 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.685 $Y=1.35
+ $X2=8.6 $Y2=1.35
r103 30 32 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=8.685 $Y=1.35
+ $X2=9.15 $Y2=1.35
r104 28 35 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.6 $Y=1.515
+ $X2=8.6 $Y2=1.35
r105 28 29 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=8.6 $Y=1.515
+ $X2=8.6 $Y2=1.695
r106 27 35 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.6 $Y=1.185
+ $X2=8.6 $Y2=1.35
r107 26 27 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=8.6 $Y=0.675
+ $X2=8.6 $Y2=1.185
r108 24 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.515 $Y=1.78
+ $X2=8.6 $Y2=1.695
r109 24 25 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=8.515 $Y=1.78
+ $X2=8.325 $Y2=1.78
r110 22 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.24 $Y=1.865
+ $X2=8.325 $Y2=1.78
r111 22 23 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=8.24 $Y=1.865
+ $X2=8.24 $Y2=2.58
r112 18 26 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=8.515 $Y=0.51
+ $X2=8.6 $Y2=0.675
r113 18 20 15.8897 $w=3.28e-07 $l=4.55e-07 $layer=LI1_cond $X=8.515 $Y=0.51
+ $X2=8.06 $Y2=0.51
r114 14 23 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=8.155 $Y=2.745
+ $X2=8.24 $Y2=2.58
r115 14 16 10.1275 $w=3.28e-07 $l=2.9e-07 $layer=LI1_cond $X=8.155 $Y=2.745
+ $X2=7.865 $Y2=2.745
r116 12 38 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=9.275 $Y=2.325
+ $X2=9.275 $Y2=1.515
r117 9 37 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=9.225 $Y=0.655
+ $X2=9.225 $Y2=1.185
r118 2 16 600 $w=1.7e-07 $l=7.03562e-07 $layer=licon1_PDIFF $count=1 $X=7.375
+ $Y=2.245 $X2=7.865 $Y2=2.745
r119 1 20 182 $w=1.7e-07 $l=4.66369e-07 $layer=licon1_NDIFF $count=1 $X=7.685
+ $Y=0.305 $X2=8.06 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_LP__SDFXTP_4%VPWR 1 2 3 4 5 6 7 8 27 31 35 39 45 49 51
+ 56 57 59 60 62 63 64 66 81 85 97 101 107 110 121 124 128
c154 128 0 3.05678e-20 $X=11.76 $Y=3.33
r155 127 128 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.76 $Y=3.33
+ $X2=11.76 $Y2=3.33
r156 124 125 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=3.33
+ $X2=10.8 $Y2=3.33
r157 121 122 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r158 119 121 10.8136 $w=6.6e-07 $l=5.85e-07 $layer=LI1_cond $X=8.86 $Y=2.745
+ $X2=8.86 $Y2=3.33
r159 117 119 4.71364 $w=6.6e-07 $l=3.40624e-07 $layer=LI1_cond $X=9.06 $Y=2.49
+ $X2=8.86 $Y2=2.745
r160 113 114 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r161 110 113 9.07985 $w=3.28e-07 $l=2.6e-07 $layer=LI1_cond $X=6.575 $Y=3.07
+ $X2=6.575 $Y2=3.33
r162 107 108 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r163 105 128 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=3.33
+ $X2=11.76 $Y2=3.33
r164 105 125 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=3.33
+ $X2=10.8 $Y2=3.33
r165 104 105 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.28 $Y=3.33
+ $X2=11.28 $Y2=3.33
r166 102 124 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.035 $Y=3.33
+ $X2=10.87 $Y2=3.33
r167 102 104 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=11.035 $Y=3.33
+ $X2=11.28 $Y2=3.33
r168 101 127 4.76062 $w=1.7e-07 $l=2.17e-07 $layer=LI1_cond $X=11.565 $Y=3.33
+ $X2=11.782 $Y2=3.33
r169 101 104 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=11.565 $Y=3.33
+ $X2=11.28 $Y2=3.33
r170 100 125 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=3.33
+ $X2=10.8 $Y2=3.33
r171 99 100 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.32 $Y=3.33
+ $X2=10.32 $Y2=3.33
r172 97 124 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.705 $Y=3.33
+ $X2=10.87 $Y2=3.33
r173 97 99 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=10.705 $Y=3.33
+ $X2=10.32 $Y2=3.33
r174 96 100 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.84 $Y=3.33
+ $X2=10.32 $Y2=3.33
r175 96 122 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=9.84 $Y=3.33
+ $X2=8.88 $Y2=3.33
r176 95 96 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r177 93 121 8.93547 $w=1.7e-07 $l=3.65e-07 $layer=LI1_cond $X=9.225 $Y=3.33
+ $X2=8.86 $Y2=3.33
r178 93 95 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=9.225 $Y=3.33
+ $X2=9.84 $Y2=3.33
r179 92 122 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=8.88 $Y2=3.33
r180 91 92 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r181 89 92 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=8.4 $Y2=3.33
r182 89 114 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=6.48 $Y2=3.33
r183 88 91 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=6.96 $Y=3.33
+ $X2=8.4 $Y2=3.33
r184 88 89 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r185 86 113 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.74 $Y=3.33
+ $X2=6.575 $Y2=3.33
r186 86 88 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=6.74 $Y=3.33
+ $X2=6.96 $Y2=3.33
r187 85 121 8.93547 $w=1.7e-07 $l=3.65e-07 $layer=LI1_cond $X=8.495 $Y=3.33
+ $X2=8.86 $Y2=3.33
r188 85 91 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=8.495 $Y=3.33
+ $X2=8.4 $Y2=3.33
r189 83 84 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r190 81 113 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.41 $Y=3.33
+ $X2=6.575 $Y2=3.33
r191 81 83 152.011 $w=1.68e-07 $l=2.33e-06 $layer=LI1_cond $X=6.41 $Y=3.33
+ $X2=4.08 $Y2=3.33
r192 80 84 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r193 79 80 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r194 77 80 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r195 76 77 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r196 74 77 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r197 74 108 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r198 73 76 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r199 73 74 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r200 71 107 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.355 $Y=3.33
+ $X2=1.19 $Y2=3.33
r201 71 73 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=1.355 $Y=3.33
+ $X2=1.68 $Y2=3.33
r202 69 108 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r203 68 69 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r204 66 107 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.025 $Y=3.33
+ $X2=1.19 $Y2=3.33
r205 66 68 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.025 $Y=3.33
+ $X2=0.72 $Y2=3.33
r206 64 114 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33
+ $X2=6.48 $Y2=3.33
r207 64 84 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r208 62 95 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=9.845 $Y=3.33
+ $X2=9.84 $Y2=3.33
r209 62 63 7.94884 $w=1.7e-07 $l=1.47e-07 $layer=LI1_cond $X=9.845 $Y=3.33
+ $X2=9.992 $Y2=3.33
r210 61 99 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=10.14 $Y=3.33
+ $X2=10.32 $Y2=3.33
r211 61 63 7.94884 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=10.14 $Y=3.33
+ $X2=9.992 $Y2=3.33
r212 59 79 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=3.7 $Y=3.33 $X2=3.6
+ $Y2=3.33
r213 59 60 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.7 $Y=3.33 $X2=3.83
+ $Y2=3.33
r214 58 83 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=3.96 $Y=3.33
+ $X2=4.08 $Y2=3.33
r215 58 60 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.96 $Y=3.33
+ $X2=3.83 $Y2=3.33
r216 56 76 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=2.82 $Y=3.33
+ $X2=2.64 $Y2=3.33
r217 56 57 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.82 $Y=3.33
+ $X2=2.915 $Y2=3.33
r218 55 79 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=3.01 $Y=3.33 $X2=3.6
+ $Y2=3.33
r219 55 57 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=3.01 $Y=3.33
+ $X2=2.915 $Y2=3.33
r220 51 54 26.8903 $w=3.28e-07 $l=7.7e-07 $layer=LI1_cond $X=11.73 $Y=2.18
+ $X2=11.73 $Y2=2.95
r221 49 127 3.00555 $w=3.3e-07 $l=1.07912e-07 $layer=LI1_cond $X=11.73 $Y=3.245
+ $X2=11.782 $Y2=3.33
r222 49 54 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=11.73 $Y=3.245
+ $X2=11.73 $Y2=2.95
r223 45 48 30.3826 $w=3.28e-07 $l=8.7e-07 $layer=LI1_cond $X=10.87 $Y=2.08
+ $X2=10.87 $Y2=2.95
r224 43 124 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.87 $Y=3.245
+ $X2=10.87 $Y2=3.33
r225 43 48 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=10.87 $Y=3.245
+ $X2=10.87 $Y2=2.95
r226 39 42 37.8939 $w=2.93e-07 $l=9.7e-07 $layer=LI1_cond $X=9.992 $Y=1.98
+ $X2=9.992 $Y2=2.95
r227 37 63 0.543863 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=9.992 $Y=3.245
+ $X2=9.992 $Y2=3.33
r228 37 42 11.5244 $w=2.93e-07 $l=2.95e-07 $layer=LI1_cond $X=9.992 $Y=3.245
+ $X2=9.992 $Y2=2.95
r229 33 60 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=3.83 $Y=3.245
+ $X2=3.83 $Y2=3.33
r230 33 35 19.5029 $w=2.58e-07 $l=4.4e-07 $layer=LI1_cond $X=3.83 $Y=3.245
+ $X2=3.83 $Y2=2.805
r231 29 57 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=2.915 $Y=3.245
+ $X2=2.915 $Y2=3.33
r232 29 31 24.5167 $w=1.88e-07 $l=4.2e-07 $layer=LI1_cond $X=2.915 $Y=3.245
+ $X2=2.915 $Y2=2.825
r233 25 107 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.19 $Y=3.245
+ $X2=1.19 $Y2=3.33
r234 25 27 15.3659 $w=3.28e-07 $l=4.4e-07 $layer=LI1_cond $X=1.19 $Y=3.245
+ $X2=1.19 $Y2=2.805
r235 8 54 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=11.59
+ $Y=1.835 $X2=11.73 $Y2=2.95
r236 8 51 400 $w=1.7e-07 $l=4.09054e-07 $layer=licon1_PDIFF $count=1 $X=11.59
+ $Y=1.835 $X2=11.73 $Y2=2.18
r237 7 48 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=10.73
+ $Y=1.835 $X2=10.87 $Y2=2.95
r238 7 45 400 $w=1.7e-07 $l=3.07124e-07 $layer=licon1_PDIFF $count=1 $X=10.73
+ $Y=1.835 $X2=10.87 $Y2=2.08
r239 6 42 400 $w=1.7e-07 $l=1.17584e-06 $layer=licon1_PDIFF $count=1 $X=9.885
+ $Y=1.835 $X2=10.01 $Y2=2.95
r240 6 39 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=9.885
+ $Y=1.835 $X2=10.01 $Y2=1.98
r241 5 119 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=8.515
+ $Y=2.535 $X2=8.655 $Y2=2.745
r242 5 117 300 $w=1.7e-07 $l=5.67054e-07 $layer=licon1_PDIFF $count=2 $X=8.515
+ $Y=2.535 $X2=9.06 $Y2=2.49
r243 4 110 600 $w=1.7e-07 $l=9.28507e-07 $layer=licon1_PDIFF $count=1 $X=6.355
+ $Y=2.245 $X2=6.575 $Y2=3.07
r244 3 35 600 $w=1.7e-07 $l=4.58258e-07 $layer=licon1_PDIFF $count=1 $X=3.74
+ $Y=2.405 $X2=3.865 $Y2=2.805
r245 2 31 600 $w=1.7e-07 $l=4.49055e-07 $layer=licon1_PDIFF $count=1 $X=2.74
+ $Y=2.455 $X2=2.915 $Y2=2.825
r246 1 27 600 $w=1.7e-07 $l=4.14126e-07 $layer=licon1_PDIFF $count=1 $X=1.05
+ $Y=2.455 $X2=1.19 $Y2=2.805
.ends

.subckt PM_SKY130_FD_SC_LP__SDFXTP_4%A_359_123# 1 2 3 4 13 19 21 22 24 26 30 33
+ 34 37 40 41 46
c113 46 0 9.22437e-20 $X=5.055 $Y=2.295
c114 40 0 1.28676e-19 $X=5.04 $Y=2.405
c115 34 0 6.94633e-20 $X=2.785 $Y=2.405
c116 30 0 1.09923e-19 $X=4.975 $Y=0.83
c117 21 0 1.34012e-19 $X=2.905 $Y=1.13
c118 19 0 1.8276e-19 $X=2.03 $Y=0.89
r119 41 46 4.98096 $w=2.68e-07 $l=1.1e-07 $layer=LI1_cond $X=5.055 $Y=2.405
+ $X2=5.055 $Y2=2.295
r120 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=2.405
+ $X2=5.04 $Y2=2.405
r121 37 44 16.305 $w=3.18e-07 $l=4.25e-07 $layer=LI1_cond $X=2.565 $Y=2.322
+ $X2=2.99 $Y2=2.322
r122 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=2.405
+ $X2=2.64 $Y2=2.405
r123 34 36 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.785 $Y=2.405
+ $X2=2.64 $Y2=2.405
r124 33 40 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.895 $Y=2.405
+ $X2=5.04 $Y2=2.405
r125 33 34 2.61138 $w=1.4e-07 $l=2.11e-06 $layer=MET1_cond $X=4.895 $Y=2.405
+ $X2=2.785 $Y2=2.405
r126 32 46 65.1381 $w=2.28e-07 $l=1.3e-06 $layer=LI1_cond $X=5.035 $Y=0.995
+ $X2=5.035 $Y2=2.295
r127 30 32 6.89702 $w=3.13e-07 $l=1.65e-07 $layer=LI1_cond $X=4.992 $Y=0.83
+ $X2=4.992 $Y2=0.995
r128 26 44 4.40442 $w=1.7e-07 $l=1.67e-07 $layer=LI1_cond $X=2.99 $Y=2.155
+ $X2=2.99 $Y2=2.322
r129 25 26 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=2.99 $Y=1.215
+ $X2=2.99 $Y2=2.155
r130 23 37 4.40442 $w=1.7e-07 $l=1.68e-07 $layer=LI1_cond $X=2.565 $Y=2.49
+ $X2=2.565 $Y2=2.322
r131 23 24 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=2.565 $Y=2.49
+ $X2=2.565 $Y2=2.64
r132 21 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.905 $Y=1.13
+ $X2=2.99 $Y2=1.215
r133 21 22 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=2.905 $Y=1.13
+ $X2=2.135 $Y2=1.13
r134 17 22 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=2.04 $Y=1.045
+ $X2=2.135 $Y2=1.13
r135 17 19 9.04785 $w=1.88e-07 $l=1.55e-07 $layer=LI1_cond $X=2.04 $Y=1.045
+ $X2=2.04 $Y2=0.89
r136 13 24 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.48 $Y=2.805
+ $X2=2.565 $Y2=2.64
r137 13 15 17.4613 $w=3.28e-07 $l=5e-07 $layer=LI1_cond $X=2.48 $Y=2.805
+ $X2=1.98 $Y2=2.805
r138 4 41 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=4.96
+ $Y=2.315 $X2=5.085 $Y2=2.46
r139 3 15 600 $w=1.7e-07 $l=4.14126e-07 $layer=licon1_PDIFF $count=1 $X=1.84
+ $Y=2.455 $X2=1.98 $Y2=2.805
r140 2 30 182 $w=1.7e-07 $l=2.60096e-07 $layer=licon1_NDIFF $count=1 $X=4.85
+ $Y=0.625 $X2=4.975 $Y2=0.83
r141 1 19 182 $w=1.7e-07 $l=3.745e-07 $layer=licon1_NDIFF $count=1 $X=1.795
+ $Y=0.615 $X2=2.03 $Y2=0.89
.ends

.subckt PM_SKY130_FD_SC_LP__SDFXTP_4%Q 1 2 3 4 15 19 23 24 25 26 29 33 38 40 41
c53 40 0 1.55372e-19 $X=11.195 $Y=1.655
c54 24 0 1.75356e-19 $X=10.535 $Y=1.03
c55 19 0 1.42881e-19 $X=10.44 $Y=1.98
r56 39 41 6.02221 $w=7.13e-07 $l=3.6e-07 $layer=LI1_cond $X=11.552 $Y=1.655
+ $X2=11.552 $Y2=1.295
r57 39 40 2.15548 $w=4.52e-07 $l=3.57e-07 $layer=LI1_cond $X=11.552 $Y=1.655
+ $X2=11.195 $Y2=1.655
r58 37 41 3.01111 $w=7.13e-07 $l=1.8e-07 $layer=LI1_cond $X=11.552 $Y=1.115
+ $X2=11.552 $Y2=1.295
r59 37 38 2.15548 $w=4.52e-07 $l=8.5e-08 $layer=LI1_cond $X=11.552 $Y=1.115
+ $X2=11.552 $Y2=1.03
r60 33 35 54.2871 $w=1.88e-07 $l=9.3e-07 $layer=LI1_cond $X=11.3 $Y=1.98
+ $X2=11.3 $Y2=2.91
r61 31 40 2.15548 $w=4.52e-07 $l=3.18198e-07 $layer=LI1_cond $X=11.3 $Y=1.925
+ $X2=11.195 $Y2=1.655
r62 31 33 3.21053 $w=1.88e-07 $l=5.5e-08 $layer=LI1_cond $X=11.3 $Y=1.925
+ $X2=11.3 $Y2=1.98
r63 27 38 2.15548 $w=4.52e-07 $l=2.91417e-07 $layer=LI1_cond $X=11.3 $Y=0.945
+ $X2=11.552 $Y2=1.03
r64 27 29 30.6459 $w=1.88e-07 $l=5.25e-07 $layer=LI1_cond $X=11.3 $Y=0.945
+ $X2=11.3 $Y2=0.42
r65 25 40 5.01601 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.195 $Y=1.74
+ $X2=11.195 $Y2=1.655
r66 25 26 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=11.195 $Y=1.74
+ $X2=10.535 $Y2=1.74
r67 23 38 5.01601 $w=1.7e-07 $l=3.57e-07 $layer=LI1_cond $X=11.195 $Y=1.03
+ $X2=11.552 $Y2=1.03
r68 23 24 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=11.195 $Y=1.03
+ $X2=10.535 $Y2=1.03
r69 19 21 47.6343 $w=2.23e-07 $l=9.3e-07 $layer=LI1_cond $X=10.422 $Y=1.98
+ $X2=10.422 $Y2=2.91
r70 17 26 6.9898 $w=1.7e-07 $l=1.49579e-07 $layer=LI1_cond $X=10.422 $Y=1.825
+ $X2=10.535 $Y2=1.74
r71 17 19 7.93905 $w=2.23e-07 $l=1.55e-07 $layer=LI1_cond $X=10.422 $Y=1.825
+ $X2=10.422 $Y2=1.98
r72 13 24 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=10.42 $Y=0.945
+ $X2=10.535 $Y2=1.03
r73 13 15 26.3058 $w=2.28e-07 $l=5.25e-07 $layer=LI1_cond $X=10.42 $Y=0.945
+ $X2=10.42 $Y2=0.42
r74 4 35 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=11.16
+ $Y=1.835 $X2=11.3 $Y2=2.91
r75 4 33 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=11.16
+ $Y=1.835 $X2=11.3 $Y2=1.98
r76 3 21 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=10.3
+ $Y=1.835 $X2=10.44 $Y2=2.91
r77 3 19 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=10.3
+ $Y=1.835 $X2=10.44 $Y2=1.98
r78 2 29 91 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=2 $X=11.16
+ $Y=0.255 $X2=11.3 $Y2=0.42
r79 1 15 91 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=2 $X=10.3
+ $Y=0.255 $X2=10.44 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__SDFXTP_4%VGND 1 2 3 4 5 6 7 8 27 31 35 39 45 49 51
+ 53 56 57 59 60 62 63 64 76 80 85 94 98 104 108 114 117 121
c137 121 0 1.28145e-19 $X=11.76 $Y=0
r138 120 121 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.76 $Y=0
+ $X2=11.76 $Y2=0
r139 117 118 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=0
+ $X2=10.8 $Y2=0
r140 114 115 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=8.88 $Y=0
+ $X2=8.88 $Y2=0
r141 108 111 10.1275 $w=3.28e-07 $l=2.9e-07 $layer=LI1_cond $X=6.42 $Y=0
+ $X2=6.42 $Y2=0.29
r142 108 109 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=0
+ $X2=6.48 $Y2=0
r143 104 105 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.08 $Y=0
+ $X2=4.08 $Y2=0
r144 102 121 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=0
+ $X2=11.76 $Y2=0
r145 102 118 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=0
+ $X2=10.8 $Y2=0
r146 101 102 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.28 $Y=0
+ $X2=11.28 $Y2=0
r147 99 117 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.035 $Y=0
+ $X2=10.87 $Y2=0
r148 99 101 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=11.035 $Y=0
+ $X2=11.28 $Y2=0
r149 98 120 4.76062 $w=1.7e-07 $l=2.17e-07 $layer=LI1_cond $X=11.565 $Y=0
+ $X2=11.782 $Y2=0
r150 98 101 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=11.565 $Y=0
+ $X2=11.28 $Y2=0
r151 97 118 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=0
+ $X2=10.8 $Y2=0
r152 96 97 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.32 $Y=0
+ $X2=10.32 $Y2=0
r153 94 117 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.705 $Y=0
+ $X2=10.87 $Y2=0
r154 94 96 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=10.705 $Y=0
+ $X2=10.32 $Y2=0
r155 93 97 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.84 $Y=0
+ $X2=10.32 $Y2=0
r156 93 115 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=9.84 $Y=0
+ $X2=8.88 $Y2=0
r157 92 93 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.84 $Y=0 $X2=9.84
+ $Y2=0
r158 90 114 8.42608 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=9.175 $Y=0
+ $X2=9.015 $Y2=0
r159 90 92 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=9.175 $Y=0 $X2=9.84
+ $Y2=0
r160 89 115 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=6.96 $Y=0
+ $X2=8.88 $Y2=0
r161 89 109 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0
+ $X2=6.48 $Y2=0
r162 88 89 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.96 $Y=0
+ $X2=6.96 $Y2=0
r163 86 108 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.585 $Y=0
+ $X2=6.42 $Y2=0
r164 86 88 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=6.585 $Y=0
+ $X2=6.96 $Y2=0
r165 85 114 8.42608 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=8.855 $Y=0
+ $X2=9.015 $Y2=0
r166 85 88 123.631 $w=1.68e-07 $l=1.895e-06 $layer=LI1_cond $X=8.855 $Y=0
+ $X2=6.96 $Y2=0
r167 81 104 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.125 $Y=0
+ $X2=3.96 $Y2=0
r168 81 83 122.326 $w=1.68e-07 $l=1.875e-06 $layer=LI1_cond $X=4.125 $Y=0 $X2=6
+ $Y2=0
r169 80 108 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.255 $Y=0
+ $X2=6.42 $Y2=0
r170 80 83 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=6.255 $Y=0 $X2=6
+ $Y2=0
r171 79 105 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r172 78 79 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r173 76 104 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.795 $Y=0
+ $X2=3.96 $Y2=0
r174 76 78 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=3.795 $Y=0 $X2=3.6
+ $Y2=0
r175 75 79 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r176 74 75 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r177 72 75 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.64
+ $Y2=0
r178 71 74 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.64
+ $Y2=0
r179 71 72 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r180 68 72 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r181 67 68 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r182 64 109 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.48
+ $Y2=0
r183 64 105 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=6 $Y=0 $X2=4.08
+ $Y2=0
r184 64 83 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6 $Y=0 $X2=6
+ $Y2=0
r185 62 92 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=9.845 $Y=0 $X2=9.84
+ $Y2=0
r186 62 63 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=9.845 $Y=0 $X2=9.99
+ $Y2=0
r187 61 96 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=10.135 $Y=0
+ $X2=10.32 $Y2=0
r188 61 63 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=10.135 $Y=0
+ $X2=9.99 $Y2=0
r189 59 74 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=2.75 $Y=0 $X2=2.64
+ $Y2=0
r190 59 60 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.75 $Y=0 $X2=2.915
+ $Y2=0
r191 58 78 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=3.08 $Y=0 $X2=3.6
+ $Y2=0
r192 58 60 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.08 $Y=0 $X2=2.915
+ $Y2=0
r193 56 67 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=0.845 $Y=0
+ $X2=0.72 $Y2=0
r194 56 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.845 $Y=0 $X2=1.01
+ $Y2=0
r195 55 71 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=1.175 $Y=0 $X2=1.2
+ $Y2=0
r196 55 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.175 $Y=0 $X2=1.01
+ $Y2=0
r197 51 120 3.00555 $w=3.3e-07 $l=1.07912e-07 $layer=LI1_cond $X=11.73 $Y=0.085
+ $X2=11.782 $Y2=0
r198 51 53 19.0328 $w=3.28e-07 $l=5.45e-07 $layer=LI1_cond $X=11.73 $Y=0.085
+ $X2=11.73 $Y2=0.63
r199 47 117 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.87 $Y=0.085
+ $X2=10.87 $Y2=0
r200 47 49 19.0328 $w=3.28e-07 $l=5.45e-07 $layer=LI1_cond $X=10.87 $Y=0.085
+ $X2=10.87 $Y2=0.63
r201 43 63 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=9.99 $Y=0.085
+ $X2=9.99 $Y2=0
r202 43 45 12.5179 $w=2.88e-07 $l=3.15e-07 $layer=LI1_cond $X=9.99 $Y=0.085
+ $X2=9.99 $Y2=0.4
r203 39 41 16.9265 $w=3.18e-07 $l=4.7e-07 $layer=LI1_cond $X=9.015 $Y=0.38
+ $X2=9.015 $Y2=0.85
r204 37 114 0.800721 $w=3.2e-07 $l=8.5e-08 $layer=LI1_cond $X=9.015 $Y=0.085
+ $X2=9.015 $Y2=0
r205 37 39 10.6241 $w=3.18e-07 $l=2.95e-07 $layer=LI1_cond $X=9.015 $Y=0.085
+ $X2=9.015 $Y2=0.38
r206 33 104 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.96 $Y=0.085
+ $X2=3.96 $Y2=0
r207 33 35 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=3.96 $Y=0.085
+ $X2=3.96 $Y2=0.45
r208 29 60 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.915 $Y=0.085
+ $X2=2.915 $Y2=0
r209 29 31 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=2.915 $Y=0.085
+ $X2=2.915 $Y2=0.76
r210 25 57 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.01 $Y=0.085
+ $X2=1.01 $Y2=0
r211 25 27 25.8427 $w=3.28e-07 $l=7.4e-07 $layer=LI1_cond $X=1.01 $Y=0.085
+ $X2=1.01 $Y2=0.825
r212 8 53 182 $w=1.7e-07 $l=4.3946e-07 $layer=licon1_NDIFF $count=1 $X=11.59
+ $Y=0.255 $X2=11.73 $Y2=0.63
r213 7 49 182 $w=1.7e-07 $l=4.3946e-07 $layer=licon1_NDIFF $count=1 $X=10.73
+ $Y=0.255 $X2=10.87 $Y2=0.63
r214 6 45 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=9.885
+ $Y=0.255 $X2=10.01 $Y2=0.4
r215 5 41 182 $w=1.7e-07 $l=6.51997e-07 $layer=licon1_NDIFF $count=1 $X=8.775
+ $Y=0.305 $X2=9.01 $Y2=0.85
r216 5 39 182 $w=1.7e-07 $l=2.69907e-07 $layer=licon1_NDIFF $count=1 $X=8.775
+ $Y=0.305 $X2=9.01 $Y2=0.38
r217 4 111 182 $w=1.7e-07 $l=4.44578e-07 $layer=licon1_NDIFF $count=1 $X=6.165
+ $Y=0.625 $X2=6.42 $Y2=0.29
r218 3 35 182 $w=1.7e-07 $l=2.498e-07 $layer=licon1_NDIFF $count=1 $X=3.835
+ $Y=0.255 $X2=3.96 $Y2=0.45
r219 2 31 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=2.775
+ $Y=0.615 $X2=2.915 $Y2=0.76
r220 1 27 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.87
+ $Y=0.615 $X2=1.01 $Y2=0.825
.ends

