* NGSPICE file created from sky130_fd_sc_lp__o21a_2.ext - technology: sky130A

.subckt sky130_fd_sc_lp__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
M1000 a_392_51# B1 a_86_21# VNB nshort w=840000u l=150000u
+  ad=4.578e+11p pd=4.45e+06u as=2.226e+11p ps=2.21e+06u
M1001 a_86_21# B1 VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=3.528e+11p pd=3.08e+06u as=1.6758e+12p ps=1.022e+07u
M1002 a_392_51# A1 VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=7.14e+11p ps=6.74e+06u
M1003 X a_86_21# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=3.528e+11p pd=3.08e+06u as=0p ps=0u
M1004 X a_86_21# VGND VNB nshort w=840000u l=150000u
+  ad=2.352e+11p pd=2.24e+06u as=0p ps=0u
M1005 VGND a_86_21# X VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND A2 a_392_51# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR A1 a_478_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=4.032e+11p ps=3.16e+06u
M1008 VPWR a_86_21# X VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_478_367# A2 a_86_21# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

