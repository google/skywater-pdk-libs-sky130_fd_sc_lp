* File: sky130_fd_sc_lp__o21ba_4.pex.spice
* Created: Wed Sep  2 10:16:57 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O21BA_4%B1_N 3 6 8 9 13 15
c36 13 0 2.56343e-20 $X=0.525 $Y=1.375
r37 13 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.525 $Y=1.375
+ $X2=0.525 $Y2=1.54
r38 13 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.525 $Y=1.375
+ $X2=0.525 $Y2=1.21
r39 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.525
+ $Y=1.375 $X2=0.525 $Y2=1.375
r40 9 14 7.68295 $w=4.33e-07 $l=2.9e-07 $layer=LI1_cond $X=0.647 $Y=1.665
+ $X2=0.647 $Y2=1.375
r41 8 14 2.11944 $w=4.33e-07 $l=8e-08 $layer=LI1_cond $X=0.647 $Y=1.295
+ $X2=0.647 $Y2=1.375
r42 6 16 474.309 $w=1.5e-07 $l=9.25e-07 $layer=POLY_cond $X=0.585 $Y=2.465
+ $X2=0.585 $Y2=1.54
r43 3 15 175.127 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=0.545 $Y=0.665
+ $X2=0.545 $Y2=1.21
.ends

.subckt PM_SKY130_FD_SC_LP__O21BA_4%A_180_23# 1 2 3 12 16 20 24 28 32 36 40 42
+ 51 52 53 56 62 64 67 68 70 72 81
c162 70 0 1.95334e-19 $X=4.96 $Y=2.035
c163 64 0 8.21834e-20 $X=4.525 $Y=1.16
r164 81 82 6.67385 $w=3.25e-07 $l=4.5e-08 $layer=POLY_cond $X=2.265 $Y=1.51
+ $X2=2.31 $Y2=1.51
r165 78 79 6.67385 $w=3.25e-07 $l=4.5e-08 $layer=POLY_cond $X=1.835 $Y=1.51
+ $X2=1.88 $Y2=1.51
r166 75 76 5.93231 $w=3.25e-07 $l=4e-08 $layer=POLY_cond $X=1.405 $Y=1.51
+ $X2=1.445 $Y2=1.51
r167 74 75 57.84 $w=3.25e-07 $l=3.9e-07 $layer=POLY_cond $X=1.015 $Y=1.51
+ $X2=1.405 $Y2=1.51
r168 73 74 5.93231 $w=3.25e-07 $l=4e-08 $layer=POLY_cond $X=0.975 $Y=1.51
+ $X2=1.015 $Y2=1.51
r169 68 70 13.9957 $w=2.08e-07 $l=2.65e-07 $layer=LI1_cond $X=4.695 $Y=2.035
+ $X2=4.96 $Y2=2.035
r170 67 68 6.91519 $w=2.1e-07 $l=1.41244e-07 $layer=LI1_cond $X=4.61 $Y=1.93
+ $X2=4.695 $Y2=2.035
r171 66 67 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=4.61 $Y=1.245
+ $X2=4.61 $Y2=1.93
r172 65 72 4.62853 $w=1.7e-07 $l=2.35e-07 $layer=LI1_cond $X=3.675 $Y=1.16
+ $X2=3.44 $Y2=1.16
r173 64 66 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.525 $Y=1.16
+ $X2=4.61 $Y2=1.245
r174 64 65 55.4545 $w=1.68e-07 $l=8.5e-07 $layer=LI1_cond $X=4.525 $Y=1.16
+ $X2=3.675 $Y2=1.16
r175 60 72 1.72426 $w=3.3e-07 $l=1.14782e-07 $layer=LI1_cond $X=3.51 $Y=1.075
+ $X2=3.44 $Y2=1.16
r176 60 62 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=3.51 $Y=1.075
+ $X2=3.51 $Y2=0.69
r177 56 58 48.7169 $w=2.18e-07 $l=9.3e-07 $layer=LI1_cond $X=3.315 $Y=1.98
+ $X2=3.315 $Y2=2.91
r178 54 72 1.72426 $w=2.2e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.315 $Y=1.245
+ $X2=3.44 $Y2=1.16
r179 54 56 38.5021 $w=2.18e-07 $l=7.35e-07 $layer=LI1_cond $X=3.315 $Y=1.245
+ $X2=3.315 $Y2=1.98
r180 52 72 4.62853 $w=1.7e-07 $l=2.35e-07 $layer=LI1_cond $X=3.205 $Y=1.16
+ $X2=3.44 $Y2=1.16
r181 52 53 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=3.205 $Y=1.16
+ $X2=2.485 $Y2=1.16
r182 50 53 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.4 $Y=1.245
+ $X2=2.485 $Y2=1.16
r183 50 51 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=2.4 $Y=1.245
+ $X2=2.4 $Y2=1.415
r184 49 81 6.67385 $w=3.25e-07 $l=4.5e-08 $layer=POLY_cond $X=2.22 $Y=1.51
+ $X2=2.265 $Y2=1.51
r185 49 79 50.4246 $w=3.25e-07 $l=3.4e-07 $layer=POLY_cond $X=2.22 $Y=1.51
+ $X2=1.88 $Y2=1.51
r186 48 49 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.22
+ $Y=1.51 $X2=2.22 $Y2=1.51
r187 45 78 43.7508 $w=3.25e-07 $l=2.95e-07 $layer=POLY_cond $X=1.54 $Y=1.51
+ $X2=1.835 $Y2=1.51
r188 45 76 14.0892 $w=3.25e-07 $l=9.5e-08 $layer=POLY_cond $X=1.54 $Y=1.51
+ $X2=1.445 $Y2=1.51
r189 44 48 39.6938 $w=1.88e-07 $l=6.8e-07 $layer=LI1_cond $X=1.54 $Y=1.51
+ $X2=2.22 $Y2=1.51
r190 44 45 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.54
+ $Y=1.51 $X2=1.54 $Y2=1.51
r191 42 51 6.84389 $w=1.9e-07 $l=1.30767e-07 $layer=LI1_cond $X=2.315 $Y=1.51
+ $X2=2.4 $Y2=1.415
r192 42 48 5.54545 $w=1.88e-07 $l=9.5e-08 $layer=LI1_cond $X=2.315 $Y=1.51
+ $X2=2.22 $Y2=1.51
r193 38 82 20.86 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.31 $Y=1.675
+ $X2=2.31 $Y2=1.51
r194 38 40 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.31 $Y=1.675
+ $X2=2.31 $Y2=2.465
r195 34 81 20.86 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.265 $Y=1.345
+ $X2=2.265 $Y2=1.51
r196 34 36 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=2.265 $Y=1.345
+ $X2=2.265 $Y2=0.665
r197 30 79 20.86 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.88 $Y=1.675
+ $X2=1.88 $Y2=1.51
r198 30 32 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.88 $Y=1.675
+ $X2=1.88 $Y2=2.465
r199 26 78 20.86 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.835 $Y=1.345
+ $X2=1.835 $Y2=1.51
r200 26 28 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=1.835 $Y=1.345
+ $X2=1.835 $Y2=0.665
r201 22 76 20.86 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.445 $Y=1.675
+ $X2=1.445 $Y2=1.51
r202 22 24 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.445 $Y=1.675
+ $X2=1.445 $Y2=2.465
r203 18 75 20.86 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.405 $Y=1.345
+ $X2=1.405 $Y2=1.51
r204 18 20 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=1.405 $Y=1.345
+ $X2=1.405 $Y2=0.665
r205 14 74 20.86 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.015 $Y=1.675
+ $X2=1.015 $Y2=1.51
r206 14 16 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.015 $Y=1.675
+ $X2=1.015 $Y2=2.465
r207 10 73 20.86 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.975 $Y=1.345
+ $X2=0.975 $Y2=1.51
r208 10 12 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=0.975 $Y=1.345
+ $X2=0.975 $Y2=0.665
r209 3 70 600 $w=1.7e-07 $l=2.60768e-07 $layer=licon1_PDIFF $count=1 $X=4.82
+ $Y=1.835 $X2=4.96 $Y2=2.035
r210 2 58 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=3.19
+ $Y=1.835 $X2=3.33 $Y2=2.91
r211 2 56 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=3.19
+ $Y=1.835 $X2=3.33 $Y2=1.98
r212 1 62 91 $w=1.7e-07 $l=4.29331e-07 $layer=licon1_NDIFF $count=2 $X=3.37
+ $Y=0.325 $X2=3.51 $Y2=0.69
.ends

.subckt PM_SKY130_FD_SC_LP__O21BA_4%A_37_49# 1 2 9 13 17 21 25 30 33 35 38 39 41
+ 44 46 47 48 56
r100 46 47 8.35844 $w=3.68e-07 $l=1.65e-07 $layer=LI1_cond $X=0.27 $Y=2.085
+ $X2=0.27 $Y2=1.92
r101 44 47 56.4052 $w=1.73e-07 $l=8.9e-07 $layer=LI1_cond $X=0.172 $Y=1.03
+ $X2=0.172 $Y2=1.92
r102 42 54 64.1084 $w=2.03e-07 $l=2.7e-07 $layer=POLY_cond $X=2.845 $Y=1.525
+ $X2=3.115 $Y2=1.525
r103 41 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.845
+ $Y=1.51 $X2=2.845 $Y2=1.51
r104 39 49 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=2.845 $Y=1.86
+ $X2=2.51 $Y2=1.86
r105 39 41 9.25447 $w=3.28e-07 $l=2.65e-07 $layer=LI1_cond $X=2.845 $Y=1.775
+ $X2=2.845 $Y2=1.51
r106 37 49 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.51 $Y=1.945
+ $X2=2.51 $Y2=1.86
r107 37 38 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=2.51 $Y=1.945
+ $X2=2.51 $Y2=2.43
r108 36 48 4.07856 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=0.465 $Y=2.52
+ $X2=0.275 $Y2=2.52
r109 35 38 6.82373 $w=1.8e-07 $l=1.25499e-07 $layer=LI1_cond $X=2.425 $Y=2.52
+ $X2=2.51 $Y2=2.43
r110 35 36 120.768 $w=1.78e-07 $l=1.96e-06 $layer=LI1_cond $X=2.425 $Y=2.52
+ $X2=0.465 $Y2=2.52
r111 31 48 2.70642 $w=3.75e-07 $l=9e-08 $layer=LI1_cond $X=0.275 $Y=2.61
+ $X2=0.275 $Y2=2.52
r112 31 33 9.09823 $w=3.78e-07 $l=3e-07 $layer=LI1_cond $X=0.275 $Y=2.61
+ $X2=0.275 $Y2=2.91
r113 30 48 2.70642 $w=3.75e-07 $l=9.24662e-08 $layer=LI1_cond $X=0.27 $Y=2.43
+ $X2=0.275 $Y2=2.52
r114 29 46 0.622942 $w=3.68e-07 $l=2e-08 $layer=LI1_cond $X=0.27 $Y=2.105
+ $X2=0.27 $Y2=2.085
r115 29 30 10.1228 $w=3.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.27 $Y=2.105
+ $X2=0.27 $Y2=2.43
r116 23 44 8.46734 $w=3.38e-07 $l=1.7e-07 $layer=LI1_cond $X=0.255 $Y=0.86
+ $X2=0.255 $Y2=1.03
r117 23 25 14.914 $w=3.38e-07 $l=4.4e-07 $layer=LI1_cond $X=0.255 $Y=0.86
+ $X2=0.255 $Y2=0.42
r118 19 56 42.7389 $w=2.03e-07 $l=1.8e-07 $layer=POLY_cond $X=3.725 $Y=1.525
+ $X2=3.545 $Y2=1.525
r119 19 21 399.957 $w=1.5e-07 $l=7.8e-07 $layer=POLY_cond $X=3.725 $Y=1.525
+ $X2=3.725 $Y2=0.745
r120 15 56 9.92004 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=3.545 $Y=1.675
+ $X2=3.545 $Y2=1.525
r121 15 17 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.545 $Y=1.675
+ $X2=3.545 $Y2=2.465
r122 11 56 59.3596 $w=2.03e-07 $l=2.5e-07 $layer=POLY_cond $X=3.295 $Y=1.525
+ $X2=3.545 $Y2=1.525
r123 11 54 42.7389 $w=2.03e-07 $l=1.8e-07 $layer=POLY_cond $X=3.295 $Y=1.525
+ $X2=3.115 $Y2=1.525
r124 11 13 399.957 $w=1.5e-07 $l=7.8e-07 $layer=POLY_cond $X=3.295 $Y=1.525
+ $X2=3.295 $Y2=0.745
r125 7 54 9.92004 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=3.115 $Y=1.675
+ $X2=3.115 $Y2=1.525
r126 7 9 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.115 $Y=1.675
+ $X2=3.115 $Y2=2.465
r127 2 46 300 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_PDIFF $count=2 $X=0.245
+ $Y=1.835 $X2=0.37 $Y2=2.085
r128 2 33 600 $w=1.7e-07 $l=1.13578e-06 $layer=licon1_PDIFF $count=1 $X=0.245
+ $Y=1.835 $X2=0.37 $Y2=2.91
r129 1 25 91 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_NDIFF $count=2 $X=0.185
+ $Y=0.245 $X2=0.31 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__O21BA_4%A1 3 7 11 15 18 20 22 23 26 30 31 33 34 35
c87 15 0 1.95334e-19 $X=5.605 $Y=2.465
r88 34 35 15.2014 $w=3.58e-07 $l=3.95e-07 $layer=LI1_cond $X=5.04 $Y=2.405
+ $X2=5.435 $Y2=2.405
r89 33 34 28.0191 $w=1.88e-07 $l=4.8e-07 $layer=LI1_cond $X=4.56 $Y=2.405
+ $X2=5.04 $Y2=2.405
r90 31 45 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.695 $Y=1.51
+ $X2=5.695 $Y2=1.675
r91 31 44 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.695 $Y=1.51
+ $X2=5.695 $Y2=1.345
r92 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.695
+ $Y=1.51 $X2=5.695 $Y2=1.51
r93 27 30 8.76859 $w=2.28e-07 $l=1.75e-07 $layer=LI1_cond $X=5.52 $Y=1.53
+ $X2=5.695 $Y2=1.53
r94 26 33 12.5502 $w=1.88e-07 $l=2.15e-07 $layer=LI1_cond $X=4.345 $Y=2.405
+ $X2=4.56 $Y2=2.405
r95 23 42 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=4.202 $Y=1.51
+ $X2=4.202 $Y2=1.675
r96 23 41 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=4.202 $Y=1.51
+ $X2=4.202 $Y2=1.345
r97 22 25 6.17723 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=4.18 $Y=1.51
+ $X2=4.18 $Y2=1.675
r98 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.18
+ $Y=1.51 $X2=4.18 $Y2=1.51
r99 20 35 3.61205 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=5.52 $Y=2.31 $X2=5.52
+ $Y2=2.405
r100 19 27 2.50919 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=5.52 $Y=1.645
+ $X2=5.52 $Y2=1.53
r101 19 20 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=5.52 $Y=1.645
+ $X2=5.52 $Y2=2.31
r102 18 26 7.08811 $w=1.9e-07 $l=1.7621e-07 $layer=LI1_cond $X=4.21 $Y=2.31
+ $X2=4.345 $Y2=2.405
r103 18 25 27.1038 $w=2.68e-07 $l=6.35e-07 $layer=LI1_cond $X=4.21 $Y=2.31
+ $X2=4.21 $Y2=1.675
r104 15 45 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=5.605 $Y=2.465
+ $X2=5.605 $Y2=1.675
r105 11 44 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=5.605 $Y=0.745
+ $X2=5.605 $Y2=1.345
r106 7 42 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=4.315 $Y=2.465
+ $X2=4.315 $Y2=1.675
r107 3 41 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=4.235 $Y=0.745
+ $X2=4.235 $Y2=1.345
.ends

.subckt PM_SKY130_FD_SC_LP__O21BA_4%A2 3 7 11 15 17 23 24
c59 11 0 8.21834e-20 $X=5.175 $Y=0.745
c60 3 0 6.61592e-20 $X=4.745 $Y=0.745
r61 22 24 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=5.085 $Y=1.51
+ $X2=5.175 $Y2=1.51
r62 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.085
+ $Y=1.51 $X2=5.085 $Y2=1.51
r63 19 22 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=4.745 $Y=1.51
+ $X2=5.085 $Y2=1.51
r64 17 23 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=5.085 $Y=1.665
+ $X2=5.085 $Y2=1.51
r65 13 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.175 $Y=1.675
+ $X2=5.175 $Y2=1.51
r66 13 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=5.175 $Y=1.675
+ $X2=5.175 $Y2=2.465
r67 9 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.175 $Y=1.345
+ $X2=5.175 $Y2=1.51
r68 9 11 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=5.175 $Y=1.345 $X2=5.175
+ $Y2=0.745
r69 5 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.745 $Y=1.675
+ $X2=4.745 $Y2=1.51
r70 5 7 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=4.745 $Y=1.675
+ $X2=4.745 $Y2=2.465
r71 1 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.745 $Y=1.345
+ $X2=4.745 $Y2=1.51
r72 1 3 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=4.745 $Y=1.345 $X2=4.745
+ $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_LP__O21BA_4%VPWR 1 2 3 4 5 18 22 26 32 34 36 40 42 47 57
+ 66 69 73 79 83 92 95
r102 94 95 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r103 91 92 10.3517 $w=6.28e-07 $l=1.65e-07 $layer=LI1_cond $X=4.1 $Y=3.1
+ $X2=4.265 $Y2=3.1
r104 88 91 0.379707 $w=6.28e-07 $l=2e-08 $layer=LI1_cond $X=4.08 $Y=3.1 $X2=4.1
+ $Y2=3.1
r105 88 89 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r106 86 88 6.07532 $w=6.28e-07 $l=3.2e-07 $layer=LI1_cond $X=3.76 $Y=3.1
+ $X2=4.08 $Y2=3.1
r107 84 86 0.189854 $w=6.28e-07 $l=1e-08 $layer=LI1_cond $X=3.75 $Y=3.1 $X2=3.76
+ $Y2=3.1
r108 82 89 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r109 81 84 2.84781 $w=6.28e-07 $l=1.5e-07 $layer=LI1_cond $X=3.6 $Y=3.1 $X2=3.75
+ $Y2=3.1
r110 81 83 7.31405 $w=6.28e-07 $l=5e-09 $layer=LI1_cond $X=3.6 $Y=3.1 $X2=3.595
+ $Y2=3.1
r111 81 82 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r112 79 83 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=3.035 $Y=3.33
+ $X2=3.595 $Y2=3.33
r113 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r114 72 75 2.16613 $w=6.33e-07 $l=1.15e-07 $layer=LI1_cond $X=2.525 $Y=3.097
+ $X2=2.64 $Y2=3.097
r115 72 73 10.3843 $w=6.33e-07 $l=1.65e-07 $layer=LI1_cond $X=2.525 $Y=3.097
+ $X2=2.36 $Y2=3.097
r116 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r117 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r118 64 95 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33 $X2=6
+ $Y2=3.33
r119 63 64 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r120 61 64 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.52 $Y2=3.33
r121 61 89 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=4.08 $Y2=3.33
r122 60 63 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=4.56 $Y=3.33
+ $X2=5.52 $Y2=3.33
r123 60 92 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=4.56 $Y=3.33
+ $X2=4.265 $Y2=3.33
r124 60 61 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r125 57 94 3.90852 $w=1.7e-07 $l=2.32e-07 $layer=LI1_cond $X=5.775 $Y=3.33
+ $X2=6.007 $Y2=3.33
r126 57 63 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=5.775 $Y=3.33
+ $X2=5.52 $Y2=3.33
r127 56 76 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r128 56 70 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r129 55 73 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=2.16 $Y=3.33 $X2=2.36
+ $Y2=3.33
r130 55 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r131 53 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.825 $Y=3.33
+ $X2=1.66 $Y2=3.33
r132 53 55 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.825 $Y=3.33
+ $X2=2.16 $Y2=3.33
r133 51 70 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r134 51 67 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r135 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r136 48 66 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.965 $Y=3.33
+ $X2=0.8 $Y2=3.33
r137 48 50 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=0.965 $Y=3.33
+ $X2=1.2 $Y2=3.33
r138 47 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.495 $Y=3.33
+ $X2=1.66 $Y2=3.33
r139 47 50 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.495 $Y=3.33
+ $X2=1.2 $Y2=3.33
r140 45 67 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r141 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r142 42 66 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.635 $Y=3.33
+ $X2=0.8 $Y2=3.33
r143 42 44 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=0.635 $Y=3.33
+ $X2=0.24 $Y2=3.33
r144 40 82 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r145 40 76 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.64 $Y2=3.33
r146 36 39 44.7148 $w=2.48e-07 $l=9.7e-07 $layer=LI1_cond $X=5.9 $Y=1.98 $X2=5.9
+ $Y2=2.95
r147 34 94 3.23464 $w=2.5e-07 $l=1.43332e-07 $layer=LI1_cond $X=5.9 $Y=3.245
+ $X2=6.007 $Y2=3.33
r148 34 39 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=5.9 $Y=3.245
+ $X2=5.9 $Y2=2.95
r149 30 84 4.89649 $w=3.1e-07 $l=3.15e-07 $layer=LI1_cond $X=3.75 $Y=2.785
+ $X2=3.75 $Y2=3.1
r150 30 32 29.9263 $w=3.08e-07 $l=8.05e-07 $layer=LI1_cond $X=3.75 $Y=2.785
+ $X2=3.75 $Y2=1.98
r151 24 79 9.81922 $w=6.33e-07 $l=1.35e-07 $layer=LI1_cond $X=2.9 $Y=3.097
+ $X2=3.035 $Y2=3.097
r152 24 75 4.89733 $w=6.33e-07 $l=2.6e-07 $layer=LI1_cond $X=2.9 $Y=3.097
+ $X2=2.64 $Y2=3.097
r153 24 26 21.3415 $w=2.68e-07 $l=5e-07 $layer=LI1_cond $X=2.9 $Y=2.78 $X2=2.9
+ $Y2=2.28
r154 20 69 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.66 $Y=3.245
+ $X2=1.66 $Y2=3.33
r155 20 22 12.2229 $w=3.28e-07 $l=3.5e-07 $layer=LI1_cond $X=1.66 $Y=3.245
+ $X2=1.66 $Y2=2.895
r156 16 66 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.8 $Y=3.245 $X2=0.8
+ $Y2=3.33
r157 16 18 12.2229 $w=3.28e-07 $l=3.5e-07 $layer=LI1_cond $X=0.8 $Y=3.245
+ $X2=0.8 $Y2=2.895
r158 5 39 400 $w=1.7e-07 $l=1.20163e-06 $layer=licon1_PDIFF $count=1 $X=5.68
+ $Y=1.835 $X2=5.86 $Y2=2.95
r159 5 36 400 $w=1.7e-07 $l=2.41868e-07 $layer=licon1_PDIFF $count=1 $X=5.68
+ $Y=1.835 $X2=5.86 $Y2=1.98
r160 4 91 600 $w=1.7e-07 $l=1.33358e-06 $layer=licon1_PDIFF $count=1 $X=3.62
+ $Y=1.835 $X2=4.1 $Y2=2.95
r161 4 86 600 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=3.62
+ $Y=1.835 $X2=3.76 $Y2=2.95
r162 4 32 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=3.62
+ $Y=1.835 $X2=3.76 $Y2=1.98
r163 3 24 600 $w=1.7e-07 $l=1.36848e-06 $layer=licon1_PDIFF $count=1 $X=2.385
+ $Y=1.835 $X2=2.9 $Y2=2.97
r164 3 72 600 $w=1.7e-07 $l=1.17792e-06 $layer=licon1_PDIFF $count=1 $X=2.385
+ $Y=1.835 $X2=2.525 $Y2=2.945
r165 3 26 300 $w=1.7e-07 $l=7.03136e-07 $layer=licon1_PDIFF $count=2 $X=2.385
+ $Y=1.835 $X2=2.9 $Y2=2.28
r166 2 22 600 $w=1.7e-07 $l=1.12783e-06 $layer=licon1_PDIFF $count=1 $X=1.52
+ $Y=1.835 $X2=1.66 $Y2=2.895
r167 1 18 600 $w=1.7e-07 $l=1.12783e-06 $layer=licon1_PDIFF $count=1 $X=0.66
+ $Y=1.835 $X2=0.8 $Y2=2.895
.ends

.subckt PM_SKY130_FD_SC_LP__O21BA_4%X 1 2 3 4 15 18 19 23 25 26 27 28 29 35
c51 25 0 2.56343e-20 $X=1.16 $Y=1.16
r52 28 29 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=1.68 $Y=2.095
+ $X2=2.095 $Y2=2.095
r53 27 35 2.84813 $w=3.35e-07 $l=8.5e-08 $layer=LI1_cond $X=1.12 $Y=2.09
+ $X2=1.035 $Y2=2.09
r54 27 39 2.84813 $w=3.35e-07 $l=8.74643e-08 $layer=LI1_cond $X=1.12 $Y=2.09
+ $X2=1.205 $Y2=2.095
r55 27 28 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=1.23 $Y=2.095
+ $X2=1.68 $Y2=2.095
r56 27 39 0.873063 $w=3.28e-07 $l=2.5e-08 $layer=LI1_cond $X=1.23 $Y=2.095
+ $X2=1.205 $Y2=2.095
r57 26 35 10.677 $w=3.38e-07 $l=3.15e-07 $layer=LI1_cond $X=0.72 $Y=2.09
+ $X2=1.035 $Y2=2.09
r58 21 23 38.2345 $w=1.88e-07 $l=6.55e-07 $layer=LI1_cond $X=2.05 $Y=1.075
+ $X2=2.05 $Y2=0.42
r59 20 25 2.11342 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.285 $Y=1.16
+ $X2=1.16 $Y2=1.16
r60 19 21 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=1.955 $Y=1.16
+ $X2=2.05 $Y2=1.075
r61 19 20 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.955 $Y=1.16
+ $X2=1.285 $Y2=1.16
r62 18 27 3.86674 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=1.12 $Y=1.92 $X2=1.12
+ $Y2=2.09
r63 17 25 4.3182 $w=2.1e-07 $l=1.03078e-07 $layer=LI1_cond $X=1.12 $Y=1.245
+ $X2=1.16 $Y2=1.16
r64 17 18 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=1.12 $Y=1.245
+ $X2=1.12 $Y2=1.92
r65 13 25 4.3182 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=1.16 $Y=1.075 $X2=1.16
+ $Y2=1.16
r66 13 15 30.194 $w=2.48e-07 $l=6.55e-07 $layer=LI1_cond $X=1.16 $Y=1.075
+ $X2=1.16 $Y2=0.42
r67 4 29 600 $w=1.7e-07 $l=3.2249e-07 $layer=licon1_PDIFF $count=1 $X=1.955
+ $Y=1.835 $X2=2.095 $Y2=2.095
r68 3 27 600 $w=1.7e-07 $l=3.2249e-07 $layer=licon1_PDIFF $count=1 $X=1.09
+ $Y=1.835 $X2=1.23 $Y2=2.095
r69 2 23 91 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=2 $X=1.91
+ $Y=0.245 $X2=2.05 $Y2=0.42
r70 1 15 91 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=2 $X=1.05
+ $Y=0.245 $X2=1.19 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__O21BA_4%A_878_367# 1 2 11
r14 8 11 30.0334 $w=3.28e-07 $l=8.6e-07 $layer=LI1_cond $X=4.53 $Y=2.835
+ $X2=5.39 $Y2=2.835
r15 2 11 600 $w=1.7e-07 $l=1.06771e-06 $layer=licon1_PDIFF $count=1 $X=5.25
+ $Y=1.835 $X2=5.39 $Y2=2.835
r16 1 8 600 $w=1.7e-07 $l=1.06771e-06 $layer=licon1_PDIFF $count=1 $X=4.39
+ $Y=1.835 $X2=4.53 $Y2=2.835
.ends

.subckt PM_SKY130_FD_SC_LP__O21BA_4%VGND 1 2 3 4 5 18 22 26 30 34 37 38 39 41 46
+ 51 56 66 67 70 73 76 79
r93 79 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r94 76 77 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r95 73 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r96 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r97 66 67 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=0 $X2=6 $Y2=0
r98 64 67 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=6
+ $Y2=0
r99 64 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=4.56
+ $Y2=0
r100 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r101 61 79 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=4.695 $Y=0 $X2=4.525
+ $Y2=0
r102 61 63 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=4.695 $Y=0 $X2=5.04
+ $Y2=0
r103 60 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=4.56
+ $Y2=0
r104 59 60 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r105 57 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.645 $Y=0 $X2=2.48
+ $Y2=0
r106 57 59 93.6203 $w=1.68e-07 $l=1.435e-06 $layer=LI1_cond $X=2.645 $Y=0
+ $X2=4.08 $Y2=0
r107 56 79 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=4.355 $Y=0 $X2=4.525
+ $Y2=0
r108 56 59 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=4.355 $Y=0
+ $X2=4.08 $Y2=0
r109 55 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r110 55 74 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.68
+ $Y2=0
r111 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r112 52 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.785 $Y=0 $X2=1.62
+ $Y2=0
r113 52 54 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.785 $Y=0
+ $X2=2.16 $Y2=0
r114 51 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.315 $Y=0 $X2=2.48
+ $Y2=0
r115 51 54 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=2.315 $Y=0
+ $X2=2.16 $Y2=0
r116 50 74 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r117 50 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r118 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r119 47 70 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=0.865 $Y=0 $X2=0.73
+ $Y2=0
r120 47 49 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=0.865 $Y=0 $X2=1.2
+ $Y2=0
r121 46 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.455 $Y=0 $X2=1.62
+ $Y2=0
r122 46 49 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=1.455 $Y=0 $X2=1.2
+ $Y2=0
r123 44 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r124 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r125 41 70 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=0.595 $Y=0 $X2=0.73
+ $Y2=0
r126 41 43 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=0.595 $Y=0
+ $X2=0.24 $Y2=0
r127 39 60 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=4.08
+ $Y2=0
r128 39 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.64
+ $Y2=0
r129 37 63 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=5.225 $Y=0
+ $X2=5.04 $Y2=0
r130 37 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.225 $Y=0 $X2=5.39
+ $Y2=0
r131 36 66 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=5.555 $Y=0 $X2=6
+ $Y2=0
r132 36 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.555 $Y=0 $X2=5.39
+ $Y2=0
r133 32 38 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.39 $Y=0.085
+ $X2=5.39 $Y2=0
r134 32 34 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=5.39 $Y=0.085
+ $X2=5.39 $Y2=0.45
r135 28 79 0.987631 $w=3.4e-07 $l=8.5e-08 $layer=LI1_cond $X=4.525 $Y=0.085
+ $X2=4.525 $Y2=0
r136 28 30 12.3718 $w=3.38e-07 $l=3.65e-07 $layer=LI1_cond $X=4.525 $Y=0.085
+ $X2=4.525 $Y2=0.45
r137 24 76 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.48 $Y=0.085
+ $X2=2.48 $Y2=0
r138 24 26 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=2.48 $Y=0.085
+ $X2=2.48 $Y2=0.39
r139 20 73 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.62 $Y=0.085
+ $X2=1.62 $Y2=0
r140 20 22 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=1.62 $Y=0.085
+ $X2=1.62 $Y2=0.39
r141 16 70 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=0.085
+ $X2=0.73 $Y2=0
r142 16 18 13.0183 $w=2.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.73 $Y=0.085
+ $X2=0.73 $Y2=0.39
r143 5 34 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=5.25
+ $Y=0.325 $X2=5.39 $Y2=0.45
r144 4 30 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=4.31
+ $Y=0.325 $X2=4.52 $Y2=0.45
r145 3 26 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.34
+ $Y=0.245 $X2=2.48 $Y2=0.39
r146 2 22 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.48
+ $Y=0.245 $X2=1.62 $Y2=0.39
r147 1 18 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=0.62
+ $Y=0.245 $X2=0.76 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_LP__O21BA_4%A_575_65# 1 2 3 4 15 17 18 22 23 24 27 33 34
+ 37
c59 17 0 6.61592e-20 $X=3.855 $Y=0.35
r60 35 37 25.8233 $w=2.68e-07 $l=6.05e-07 $layer=LI1_cond $X=5.87 $Y=1.075
+ $X2=5.87 $Y2=0.47
r61 33 35 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=5.735 $Y=1.16
+ $X2=5.87 $Y2=1.075
r62 33 34 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=5.735 $Y=1.16
+ $X2=5.055 $Y2=1.16
r63 30 34 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=4.96 $Y=1.075
+ $X2=5.055 $Y2=1.16
r64 30 32 3.21053 $w=1.88e-07 $l=5.5e-08 $layer=LI1_cond $X=4.96 $Y=1.075
+ $X2=4.96 $Y2=1.02
r65 29 39 4.70473 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=4.96 $Y=0.895
+ $X2=4.96 $Y2=0.81
r66 29 32 7.29665 $w=1.88e-07 $l=1.25e-07 $layer=LI1_cond $X=4.96 $Y=0.895
+ $X2=4.96 $Y2=1.02
r67 25 39 4.70473 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=4.96 $Y=0.725
+ $X2=4.96 $Y2=0.81
r68 25 27 15.4689 $w=1.88e-07 $l=2.65e-07 $layer=LI1_cond $X=4.96 $Y=0.725
+ $X2=4.96 $Y2=0.46
r69 23 39 1.74598 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=4.865 $Y=0.81
+ $X2=4.96 $Y2=0.81
r70 23 24 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=4.865 $Y=0.81
+ $X2=4.185 $Y2=0.81
r71 20 24 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.02 $Y=0.725
+ $X2=4.185 $Y2=0.81
r72 20 22 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=4.02 $Y=0.725
+ $X2=4.02 $Y2=0.45
r73 19 22 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=4.02 $Y=0.435
+ $X2=4.02 $Y2=0.45
r74 17 19 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.855 $Y=0.35
+ $X2=4.02 $Y2=0.435
r75 17 18 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=3.855 $Y=0.35
+ $X2=3.175 $Y2=0.35
r76 13 18 7.85115 $w=1.7e-07 $l=2.08207e-07 $layer=LI1_cond $X=3.005 $Y=0.435
+ $X2=3.175 $Y2=0.35
r77 13 15 1.18634 $w=3.38e-07 $l=3.5e-08 $layer=LI1_cond $X=3.005 $Y=0.435
+ $X2=3.005 $Y2=0.47
r78 4 37 91 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_NDIFF $count=2 $X=5.68
+ $Y=0.325 $X2=5.84 $Y2=0.47
r79 3 32 182 $w=1.7e-07 $l=7.61791e-07 $layer=licon1_NDIFF $count=1 $X=4.82
+ $Y=0.325 $X2=4.96 $Y2=1.02
r80 3 27 182 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_NDIFF $count=1 $X=4.82
+ $Y=0.325 $X2=4.96 $Y2=0.46
r81 2 22 91 $w=1.7e-07 $l=2.755e-07 $layer=licon1_NDIFF $count=2 $X=3.8 $Y=0.325
+ $X2=4.02 $Y2=0.45
r82 1 15 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=2.875
+ $Y=0.325 $X2=3.01 $Y2=0.47
.ends

