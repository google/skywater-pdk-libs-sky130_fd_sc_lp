* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__dlclkp_lp CLK GATE VGND VNB VPB VPWR GCLK
X0 a_1147_419# a_584_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X1 a_352_419# a_80_21# a_526_419# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X2 a_80_21# CLK a_923_185# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 VPWR GATE a_254_419# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X4 a_110_47# a_80_21# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 a_352_419# a_27_47# a_448_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 a_27_47# a_80_21# a_110_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 a_1284_47# a_1147_419# GCLK VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 VGND GATE a_284_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 a_254_419# a_27_47# a_352_419# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X10 a_80_21# CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X11 VGND a_1147_419# a_1284_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 VGND CLK a_1104_185# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X13 a_27_47# a_80_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X14 a_526_419# a_584_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X15 VPWR a_1147_419# GCLK VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X16 a_700_47# a_352_419# a_584_21# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X17 a_448_47# a_584_21# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X18 a_923_185# CLK VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X19 VGND a_352_419# a_700_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X20 VPWR CLK a_1147_419# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X21 a_1104_185# a_584_21# a_1147_419# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X22 a_284_47# a_80_21# a_352_419# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X23 VPWR a_352_419# a_584_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
.ends
