* File: sky130_fd_sc_lp__sdfxbp_2.spice
* Created: Fri Aug 28 11:30:24 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__sdfxbp_2.pex.spice"
.subckt sky130_fd_sc_lp__sdfxbp_2  VNB VPB SCD D SCE CLK VPWR Q Q_N VGND
* 
* VGND	VGND
* Q_N	Q_N
* Q	Q
* VPWR	VPWR
* CLK	CLK
* SCE	SCE
* D	D
* SCD	SCD
* VPB	VPB
* VNB	VNB
MM1035 A_110_120# N_SCD_M1035_g N_VGND_M1035_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1113 PD=0.63 PS=1.37 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002 A=0.063 P=1.14 MULT=1
MM1020 N_A_182_120#_M1020_d N_SCE_M1020_g A_110_120# VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6
+ SB=75001.6 A=0.063 P=1.14 MULT=1
MM1006 A_268_120# N_D_M1006_g N_A_182_120#_M1020_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0672 AS=0.0588 PD=0.74 PS=0.7 NRD=30 NRS=0 M=1 R=2.8 SA=75001 SB=75001.2
+ A=0.063 P=1.14 MULT=1
MM1026 N_VGND_M1026_d N_A_332_94#_M1026_g A_268_120# VNB NSHORT L=0.15 W=0.42
+ AD=0.0756 AS=0.0672 PD=0.78 PS=0.74 NRD=0 NRS=30 M=1 R=2.8 SA=75001.4
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1003 N_A_332_94#_M1003_d N_SCE_M1003_g N_VGND_M1026_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.0756 PD=1.37 PS=0.78 NRD=0 NRS=22.848 M=1 R=2.8 SA=75002
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1013 N_VGND_M1013_d N_A_733_21#_M1013_g N_A_778_399#_M1013_s VNB NSHORT L=0.15
+ W=0.64 AD=0.304181 AS=0.1696 PD=1.76906 PS=1.81 NRD=76.872 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75001.5 A=0.096 P=1.58 MULT=1
MM1031 A_1060_119# N_A_778_399#_M1031_g N_VGND_M1013_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.199619 PD=0.63 PS=1.16094 NRD=14.28 NRS=39.276 M=1 R=2.8
+ SA=75001.2 SB=75001 A=0.063 P=1.14 MULT=1
MM1017 N_A_733_21#_M1017_d N_A_1102_93#_M1017_g A_1060_119# VNB NSHORT L=0.15
+ W=0.42 AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.5
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1010 N_A_182_120#_M1010_d N_A_1188_93#_M1010_g N_A_733_21#_M1017_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8
+ SA=75002 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1016 N_VGND_M1016_d N_A_1188_93#_M1016_g N_A_1102_93#_M1016_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1018 N_A_1188_93#_M1018_d N_CLK_M1018_g N_VGND_M1016_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1021 N_A_2008_122#_M1021_d N_A_1102_93#_M1021_g N_A_778_399#_M1021_s VNB
+ NSHORT L=0.15 W=0.42 AD=0.06195 AS=0.1113 PD=0.715 PS=1.37 NRD=4.284 NRS=0 M=1
+ R=2.8 SA=75000.2 SB=75001.7 A=0.063 P=1.14 MULT=1
MM1015 A_2097_122# N_A_1188_93#_M1015_g N_A_2008_122#_M1021_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.06195 PD=0.63 PS=0.715 NRD=14.28 NRS=0 M=1 R=2.8
+ SA=75000.6 SB=75001.2 A=0.063 P=1.14 MULT=1
MM1000 N_VGND_M1000_d N_A_2122_329#_M1000_g A_2097_122# VNB NSHORT L=0.15 W=0.42
+ AD=0.121602 AS=0.0441 PD=0.943019 PS=0.63 NRD=47.136 NRS=14.28 M=1 R=2.8
+ SA=75001 SB=75000.9 A=0.063 P=1.14 MULT=1
MM1032 N_A_2122_329#_M1032_d N_A_2008_122#_M1032_g N_VGND_M1000_d VNB NSHORT
+ L=0.15 W=0.64 AD=0.1696 AS=0.185298 PD=1.81 PS=1.43698 NRD=0 NRS=20.148 M=1
+ R=4.26667 SA=75001.2 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1002 N_Q_M1002_d N_A_2122_329#_M1002_g N_VGND_M1002_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75000.9 A=0.126 P=1.98 MULT=1
MM1019 N_Q_M1002_d N_A_2122_329#_M1019_g N_VGND_M1019_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1792 PD=1.12 PS=1.62 NRD=0 NRS=6.78 M=1 R=5.6 SA=75000.6
+ SB=75000.5 A=0.126 P=1.98 MULT=1
MM1029 N_A_2710_56#_M1029_d N_A_2122_329#_M1029_g N_VGND_M1019_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.1113 AS=0.0896 PD=1.37 PS=0.81 NRD=0 NRS=0 M=1 R=2.8
+ SA=75001.1 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1012 N_Q_N_M1012_d N_A_2710_56#_M1012_g N_VGND_M1012_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.2394 PD=1.12 PS=2.25 NRD=0 NRS=2.856 M=1 R=5.6
+ SA=75000.2 SB=75000.6 A=0.126 P=1.98 MULT=1
MM1030 N_Q_N_M1012_d N_A_2710_56#_M1030_g N_VGND_M1030_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1023 N_VPWR_M1023_d N_SCD_M1023_g N_A_27_489#_M1023_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1024 AS=0.1696 PD=0.96 PS=1.81 NRD=6.1464 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75001.4 A=0.096 P=1.58 MULT=1
MM1009 A_204_489# N_SCE_M1009_g N_VPWR_M1023_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0672 AS=0.1024 PD=0.85 PS=0.96 NRD=15.3857 NRS=6.1464 M=1 R=4.26667
+ SA=75000.7 SB=75001 A=0.096 P=1.58 MULT=1
MM1014 N_A_182_120#_M1014_d N_D_M1014_g A_204_489# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0896 AS=0.0672 PD=0.92 PS=0.85 NRD=0 NRS=15.3857 M=1 R=4.26667 SA=75001
+ SB=75000.6 A=0.096 P=1.58 MULT=1
MM1038 N_A_27_489#_M1038_d N_A_332_94#_M1038_g N_A_182_120#_M1014_d VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.1696 AS=0.0896 PD=1.81 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75001.4 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1005 N_VPWR_M1005_d N_SCE_M1005_g N_A_332_94#_M1005_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.2144 AS=0.2976 PD=1.95 PS=2.21 NRD=15.3857 NRS=61.5625 M=1
+ R=4.26667 SA=75000.4 SB=75000.3 A=0.096 P=1.58 MULT=1
MM1004 N_VPWR_M1004_d N_A_733_21#_M1004_g N_A_778_399#_M1004_s VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.1792 AS=0.3737 PD=1.62 PS=2.74 NRD=0 NRS=28.1316 M=1 R=5.6
+ SA=75000.3 SB=75000.5 A=0.126 P=1.98 MULT=1
MM1033 N_A_993_425#_M1033_d N_A_778_399#_M1033_g N_VPWR_M1004_d VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.2252 AS=0.0896 PD=2.4 PS=0.81 NRD=225.683 NRS=74.2493 M=1
+ R=2.8 SA=75000.8 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1039 N_A_733_21#_M1039_d N_A_1102_93#_M1039_g N_A_182_120#_M1039_s VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.0588 AS=0.1533 PD=0.7 PS=1.57 NRD=0 NRS=37.5088 M=1 R=2.8
+ SA=75000.3 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1024 N_A_993_425#_M1024_d N_A_1188_93#_M1024_g N_A_733_21#_M1039_d VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.1533 AS=0.0588 PD=1.57 PS=0.7 NRD=37.5088 NRS=0 M=1 R=2.8
+ SA=75000.7 SB=75000.3 A=0.063 P=1.14 MULT=1
MM1027 N_VPWR_M1027_d N_A_1188_93#_M1027_g N_A_1102_93#_M1027_s VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.18575 AS=0.256 PD=1.39 PS=2.08 NRD=72.3975 NRS=35.3812 M=1
+ R=4.26667 SA=75000.3 SB=75000.8 A=0.096 P=1.58 MULT=1
MM1001 N_A_1188_93#_M1001_d N_CLK_M1001_g N_VPWR_M1027_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1824 AS=0.18575 PD=1.85 PS=1.39 NRD=0 NRS=72.3975 M=1 R=4.26667
+ SA=75000.9 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1011 N_A_2008_122#_M1011_d N_A_1188_93#_M1011_g N_A_778_399#_M1011_s VPB
+ PHIGHVT L=0.15 W=0.84 AD=0.1806 AS=0.2394 PD=1.6 PS=2.25 NRD=0 NRS=0 M=1 R=5.6
+ SA=75000.2 SB=75000.9 A=0.126 P=1.98 MULT=1
MM1034 A_2116_463# N_A_1102_93#_M1034_g N_A_2008_122#_M1011_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0441 AS=0.0903 PD=0.63 PS=0.8 NRD=23.443 NRS=37.5088 M=1 R=2.8
+ SA=75000.7 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1036 N_VPWR_M1036_d N_A_2122_329#_M1036_g A_2116_463# VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0966 AS=0.0441 PD=0.843333 PS=0.63 NRD=0 NRS=23.443 M=1 R=2.8
+ SA=75001.1 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1025 N_A_2122_329#_M1025_d N_A_2008_122#_M1025_g N_VPWR_M1036_d VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.2226 AS=0.1932 PD=2.21 PS=1.68667 NRD=0 NRS=17.0011 M=1
+ R=5.6 SA=75000.9 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1022 N_VPWR_M1022_d N_A_2122_329#_M1022_g N_Q_M1022_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75000.9 A=0.189 P=2.82 MULT=1
MM1037 N_VPWR_M1037_d N_A_2122_329#_M1037_g N_Q_M1022_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.268115 AS=0.1764 PD=2.16853 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.6 SB=75000.5 A=0.189 P=2.82 MULT=1
MM1007 N_A_2710_56#_M1007_d N_A_2122_329#_M1007_g N_VPWR_M1037_d VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.1696 AS=0.136185 PD=1.81 PS=1.10147 NRD=0 NRS=48.5605 M=1
+ R=4.26667 SA=75001.1 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1008 N_VPWR_M1008_d N_A_2710_56#_M1008_g N_Q_N_M1008_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1028 N_VPWR_M1028_d N_A_2710_56#_M1028_g N_Q_N_M1008_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX40_noxref VNB VPB NWDIODE A=29.3551 P=35.21
c_277 VPB 0 1.59193e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_lp__sdfxbp_2.pxi.spice"
*
.ends
*
*
