* NGSPICE file created from sky130_fd_sc_lp__sdfrtp_4.ext - technology: sky130A

.subckt sky130_fd_sc_lp__sdfrtp_4 CLK D RESET_B SCD SCE VGND VNB VPB VPWR Q
M1000 VGND SCE a_27_74# VNB nshort w=420000u l=150000u
+  ad=1.8964e+12p pd=1.655e+07u as=1.113e+11p ps=1.37e+06u
M1001 VGND RESET_B a_217_50# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=2.289e+11p ps=2.77e+06u
M1002 VPWR SCE a_27_74# VPB phighvt w=640000u l=150000u
+  ad=3.1901e+12p pd=2.491e+07u as=1.696e+11p ps=1.81e+06u
M1003 VPWR a_1047_369# a_1005_463# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1004 VPWR a_975_255# a_851_242# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=3.402e+11p ps=3.06e+06u
M1005 Q a_2555_47# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=7.056e+11p pd=6.16e+06u as=0p ps=0u
M1006 a_1705_113# a_975_255# a_1524_69# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=3.754e+11p ps=2.79e+06u
M1007 a_1005_463# a_975_255# a_881_463# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=3.087e+11p ps=3.15e+06u
M1008 VPWR a_2555_47# Q VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_881_463# RESET_B VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_1524_69# a_975_255# a_1047_369# VPB phighvt w=840000u l=150000u
+  ad=4.361e+11p pd=3.32e+06u as=2.352e+11p ps=2.24e+06u
M1011 a_975_255# CLK VGND VNB nshort w=840000u l=150000u
+  ad=2.394e+11p pd=2.25e+06u as=0p ps=0u
M1012 VPWR SCD a_565_463# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=2.048e+11p ps=1.92e+06u
M1013 a_1662_533# a_851_242# a_1524_69# VPB phighvt w=420000u l=150000u
+  ad=1.848e+11p pd=1.72e+06u as=0p ps=0u
M1014 VGND a_2555_47# Q VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=5.04e+11p ps=4.56e+06u
M1015 a_1047_369# a_881_463# VGND VNB nshort w=640000u l=150000u
+  ad=3.104e+11p pd=2.25e+06u as=0p ps=0u
M1016 a_1747_21# a_1524_69# a_1902_119# VNB nshort w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=8.82e+10p ps=1.26e+06u
M1017 a_881_463# a_851_242# a_372_50# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=3.95e+11p ps=3.87e+06u
M1018 a_1747_21# RESET_B VPWR VPB phighvt w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=0p ps=0u
M1019 a_1524_69# a_851_242# a_1047_369# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_565_463# a_27_74# a_372_50# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_300_50# a_27_74# a_217_50# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1022 a_1047_369# a_881_463# VPWR VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_372_50# D a_300_50# VNB nshort w=420000u l=150000u
+  ad=3.8515e+11p pd=3.61e+06u as=0p ps=0u
M1024 a_1107_119# a_851_242# a_881_463# VNB nshort w=420000u l=150000u
+  ad=1.344e+11p pd=1.48e+06u as=1.176e+11p ps=1.4e+06u
M1025 Q a_2555_47# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_1902_119# RESET_B VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 VGND a_2555_47# Q VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 VPWR a_1747_21# a_1662_533# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 a_504_81# SCE a_372_50# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1030 a_881_463# a_975_255# a_372_50# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 VGND a_975_255# a_851_242# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=2.394e+11p ps=2.25e+06u
M1032 a_217_50# SCD a_504_81# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 a_372_50# RESET_B VPWR VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1034 VPWR a_2555_47# Q VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1035 a_407_463# SCE VPWR VPB phighvt w=640000u l=150000u
+  ad=1.344e+11p pd=1.7e+06u as=0p ps=0u
M1036 VGND RESET_B a_1201_119# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1037 a_975_255# CLK VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=3.339e+11p pd=3.05e+06u as=0p ps=0u
M1038 a_372_50# D a_407_463# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1039 VGND a_1747_21# a_1705_113# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1040 Q a_2555_47# VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1041 VGND a_1524_69# a_2555_47# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=2.226e+11p ps=2.21e+06u
M1042 VPWR a_1524_69# a_1747_21# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1043 Q a_2555_47# VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1044 VPWR a_1524_69# a_2555_47# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=3.339e+11p ps=3.05e+06u
M1045 a_1201_119# a_1047_369# a_1107_119# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

