* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__srdlxtp_1 D GATE SLEEP_B KAPWR VGND VNB VPB VPWR Q
X0 a_84_153# GATE a_1289_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 a_1361_47# SLEEP_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 a_226_491# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X3 VGND a_226_491# a_476_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 a_861_47# a_831_21# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 KAPWR GATE a_84_153# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X6 a_476_47# a_114_179# a_590_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 VPWR a_1530_367# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X8 a_662_47# a_114_179# a_849_419# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X9 a_1289_47# SLEEP_B a_1361_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 a_226_491# D VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X11 a_476_47# a_84_153# a_621_491# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X12 a_783_47# a_831_21# a_861_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X13 a_849_419# a_831_21# KAPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X14 VGND a_1530_367# Q VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X15 a_1530_367# a_662_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X16 VGND a_84_153# a_114_179# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X17 a_621_491# a_84_153# a_662_47# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X18 a_84_153# SLEEP_B KAPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X19 a_831_21# a_662_47# KAPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X20 VPWR a_226_491# a_476_47# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X21 VPWR a_84_153# a_114_179# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X22 a_1530_367# a_662_47# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X23 a_590_47# a_114_179# a_662_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X24 a_662_47# a_84_153# a_783_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X25 VGND a_662_47# a_1019_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X26 a_1019_47# a_662_47# a_831_21# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
