* File: sky130_fd_sc_lp__xor2_0.spice
* Created: Wed Sep  2 10:40:59 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__xor2_0.pex.spice"
.subckt sky130_fd_sc_lp__xor2_0  VNB VPB B A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* B	B
* VPB	VPB
* VNB	VNB
MM1009 N_A_27_481#_M1009_d N_B_M1009_g N_VGND_M1009_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75002.4
+ A=0.063 P=1.14 MULT=1
MM1002 N_VGND_M1002_d N_A_M1002_g N_A_27_481#_M1009_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6 SB=75002
+ A=0.063 P=1.14 MULT=1
MM1004 A_317_85# N_A_M1004_g N_VGND_M1002_d VNB NSHORT L=0.15 W=0.42 AD=0.0504
+ AS=0.0588 PD=0.66 PS=0.7 NRD=18.564 NRS=0 M=1 R=2.8 SA=75001.1 SB=75001.6
+ A=0.063 P=1.14 MULT=1
MM1005 N_X_M1005_d N_B_M1005_g A_317_85# VNB NSHORT L=0.15 W=0.42 AD=0.17325
+ AS=0.0504 PD=1.245 PS=0.66 NRD=5.712 NRS=18.564 M=1 R=2.8 SA=75001.4
+ SB=75001.2 A=0.063 P=1.14 MULT=1
MM1008 N_VGND_M1008_d N_A_27_481#_M1008_g N_X_M1005_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.17325 PD=1.37 PS=1.245 NRD=0 NRS=2.856 M=1 R=2.8 SA=75002.4
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1001 A_110_481# N_B_M1001_g N_A_27_481#_M1001_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0768 AS=0.1696 PD=0.88 PS=1.81 NRD=19.9955 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75001.4 A=0.096 P=1.58 MULT=1
MM1003 N_VPWR_M1003_d N_A_M1003_g A_110_481# VPB PHIGHVT L=0.15 W=0.64 AD=0.0896
+ AS=0.0768 PD=0.92 PS=0.88 NRD=0 NRS=19.9955 M=1 R=4.26667 SA=75000.6
+ SB=75001.1 A=0.096 P=1.58 MULT=1
MM1000 N_A_274_481#_M1000_d N_A_M1000_g N_VPWR_M1003_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667 SA=75001
+ SB=75000.6 A=0.096 P=1.58 MULT=1
MM1006 N_VPWR_M1006_d N_B_M1006_g N_A_274_481#_M1000_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1696 AS=0.0896 PD=1.81 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667 SA=75001.4
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1007 N_A_274_481#_M1007_d N_A_27_481#_M1007_g N_X_M1007_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1696 AS=0.1696 PD=1.81 PS=1.81 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75000.2 A=0.096 P=1.58 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9751 P=11.21
*
.include "sky130_fd_sc_lp__xor2_0.pxi.spice"
*
.ends
*
*
