* NGSPICE file created from sky130_fd_sc_lp__a211oi_lp.ext - technology: sky130A

.subckt sky130_fd_sc_lp__a211oi_lp A1 A2 B1 C1 VGND VNB VPB VPWR Y
M1000 a_295_57# B1 VGND VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=2.373e+11p ps=2.81e+06u
M1001 Y B1 a_295_57# VNB nshort w=420000u l=150000u
+  ad=2.373e+11p pd=2.81e+06u as=0p ps=0u
M1002 a_279_409# B1 a_181_409# VPB phighvt w=1e+06u l=250000u
+  ad=6.05e+11p pd=5.21e+06u as=2.4e+11p ps=2.48e+06u
M1003 a_453_57# A1 Y VNB nshort w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=0p ps=0u
M1004 a_181_409# C1 Y VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=4.9e+11p ps=2.98e+06u
M1005 VGND C1 a_137_57# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1006 a_279_409# A2 VPWR VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=5.8e+11p ps=3.16e+06u
M1007 VPWR A1 a_279_409# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_137_57# C1 Y VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND A2 a_453_57# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

