* File: sky130_fd_sc_lp__clkbuflp_16.pex.spice
* Created: Wed Sep  2 09:38:53 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__CLKBUFLP_16%A 1 3 6 8 10 13 15 17 20 22 24 25 27 30
+ 32 34 37 39 41 44 46 48 49 50 51 72
r124 71 72 2.39565 $w=6.7e-07 $l=3e-08 $layer=POLY_cond $X=3.175 $Y=1.23
+ $X2=3.205 $Y2=1.23
r125 70 71 26.3522 $w=6.7e-07 $l=3.3e-07 $layer=POLY_cond $X=2.845 $Y=1.23
+ $X2=3.175 $Y2=1.23
r126 69 70 15.971 $w=6.7e-07 $l=2e-07 $layer=POLY_cond $X=2.645 $Y=1.23
+ $X2=2.845 $Y2=1.23
r127 68 69 18.3667 $w=6.7e-07 $l=2.3e-07 $layer=POLY_cond $X=2.415 $Y=1.23
+ $X2=2.645 $Y2=1.23
r128 67 68 23.9565 $w=6.7e-07 $l=3e-07 $layer=POLY_cond $X=2.115 $Y=1.23
+ $X2=2.415 $Y2=1.23
r129 66 67 4.79131 $w=6.7e-07 $l=6e-08 $layer=POLY_cond $X=2.055 $Y=1.23
+ $X2=2.115 $Y2=1.23
r130 65 66 34.3377 $w=6.7e-07 $l=4.3e-07 $layer=POLY_cond $X=1.625 $Y=1.23
+ $X2=2.055 $Y2=1.23
r131 64 65 3.19421 $w=6.7e-07 $l=4e-08 $layer=POLY_cond $X=1.585 $Y=1.23
+ $X2=1.625 $Y2=1.23
r132 63 64 25.5536 $w=6.7e-07 $l=3.2e-07 $layer=POLY_cond $X=1.265 $Y=1.23
+ $X2=1.585 $Y2=1.23
r133 62 63 16.7696 $w=6.7e-07 $l=2.1e-07 $layer=POLY_cond $X=1.055 $Y=1.23
+ $X2=1.265 $Y2=1.23
r134 61 62 17.5681 $w=6.7e-07 $l=2.2e-07 $layer=POLY_cond $X=0.835 $Y=1.23
+ $X2=1.055 $Y2=1.23
r135 59 61 21.5609 $w=6.7e-07 $l=2.7e-07 $layer=POLY_cond $X=0.565 $Y=1.23
+ $X2=0.835 $Y2=1.23
r136 59 60 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.565
+ $Y=1.06 $X2=0.565 $Y2=1.06
r137 57 59 3.19421 $w=6.7e-07 $l=4e-08 $layer=POLY_cond $X=0.525 $Y=1.23
+ $X2=0.565 $Y2=1.23
r138 55 57 3.99276 $w=6.7e-07 $l=5e-08 $layer=POLY_cond $X=0.475 $Y=1.23
+ $X2=0.525 $Y2=1.23
r139 50 51 9.13765 $w=4.94e-07 $l=4.4699e-07 $layer=LI1_cond $X=0.41 $Y=1.295
+ $X2=0.24 $Y2=1.665
r140 50 60 5.80364 $w=4.94e-07 $l=2.35e-07 $layer=LI1_cond $X=0.41 $Y=1.295
+ $X2=0.41 $Y2=1.06
r141 49 60 3.33401 $w=4.94e-07 $l=1.35e-07 $layer=LI1_cond $X=0.41 $Y=0.925
+ $X2=0.41 $Y2=1.06
r142 46 72 38.9565 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=3.205 $Y=0.895
+ $X2=3.205 $Y2=1.23
r143 46 48 123.713 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=3.205 $Y=0.895
+ $X2=3.205 $Y2=0.51
r144 42 71 25.9839 $w=2.5e-07 $l=3.35e-07 $layer=POLY_cond $X=3.175 $Y=1.565
+ $X2=3.175 $Y2=1.23
r145 42 44 253.423 $w=2.5e-07 $l=1.02e-06 $layer=POLY_cond $X=3.175 $Y=1.565
+ $X2=3.175 $Y2=2.585
r146 39 70 38.9565 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=2.845 $Y=0.895
+ $X2=2.845 $Y2=1.23
r147 39 41 123.713 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=2.845 $Y=0.895
+ $X2=2.845 $Y2=0.51
r148 35 69 25.9839 $w=2.5e-07 $l=3.35e-07 $layer=POLY_cond $X=2.645 $Y=1.565
+ $X2=2.645 $Y2=1.23
r149 35 37 253.423 $w=2.5e-07 $l=1.02e-06 $layer=POLY_cond $X=2.645 $Y=1.565
+ $X2=2.645 $Y2=2.585
r150 32 68 38.9565 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=2.415 $Y=0.895
+ $X2=2.415 $Y2=1.23
r151 32 34 123.713 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=2.415 $Y=0.895
+ $X2=2.415 $Y2=0.51
r152 28 67 25.9839 $w=2.5e-07 $l=3.35e-07 $layer=POLY_cond $X=2.115 $Y=1.565
+ $X2=2.115 $Y2=1.23
r153 28 30 253.423 $w=2.5e-07 $l=1.02e-06 $layer=POLY_cond $X=2.115 $Y=1.565
+ $X2=2.115 $Y2=2.585
r154 25 66 38.9565 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=2.055 $Y=0.895
+ $X2=2.055 $Y2=1.23
r155 25 27 123.713 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=2.055 $Y=0.895
+ $X2=2.055 $Y2=0.51
r156 22 65 38.9565 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=1.625 $Y=0.895
+ $X2=1.625 $Y2=1.23
r157 22 24 123.713 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=1.625 $Y=0.895
+ $X2=1.625 $Y2=0.51
r158 18 64 25.9839 $w=2.5e-07 $l=3.35e-07 $layer=POLY_cond $X=1.585 $Y=1.565
+ $X2=1.585 $Y2=1.23
r159 18 20 253.423 $w=2.5e-07 $l=1.02e-06 $layer=POLY_cond $X=1.585 $Y=1.565
+ $X2=1.585 $Y2=2.585
r160 15 63 38.9565 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=1.265 $Y=0.895
+ $X2=1.265 $Y2=1.23
r161 15 17 123.713 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=1.265 $Y=0.895
+ $X2=1.265 $Y2=0.51
r162 11 62 25.9839 $w=2.5e-07 $l=3.35e-07 $layer=POLY_cond $X=1.055 $Y=1.565
+ $X2=1.055 $Y2=1.23
r163 11 13 253.423 $w=2.5e-07 $l=1.02e-06 $layer=POLY_cond $X=1.055 $Y=1.565
+ $X2=1.055 $Y2=2.585
r164 8 61 38.9565 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=0.835 $Y=0.895
+ $X2=0.835 $Y2=1.23
r165 8 10 123.713 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=0.835 $Y=0.895
+ $X2=0.835 $Y2=0.51
r166 4 57 25.9839 $w=2.5e-07 $l=3.35e-07 $layer=POLY_cond $X=0.525 $Y=1.565
+ $X2=0.525 $Y2=1.23
r167 4 6 253.423 $w=2.5e-07 $l=1.02e-06 $layer=POLY_cond $X=0.525 $Y=1.565
+ $X2=0.525 $Y2=2.585
r168 1 55 38.9565 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=0.475 $Y=0.895
+ $X2=0.475 $Y2=1.23
r169 1 3 123.713 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=0.475 $Y=0.895
+ $X2=0.475 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_LP__CLKBUFLP_16%A_130_417# 1 2 3 4 5 18 22 26 30 34 38
+ 42 46 50 54 58 62 66 70 74 78 82 86 90 94 98 102 106 110 114 118 122 126 130
+ 134 138 142 146 150 154 158 162 166 170 174 182 186 191 192 193 194 195 197
+ 201 205 208 211 214 216 274 275
c431 154 0 3.2513e-20 $X=11.125 $Y=0.51
c432 102 0 8.52417e-20 $X=8.395 $Y=0.51
c433 98 0 3.40562e-20 $X=7.965 $Y=0.51
c434 46 0 4.0915e-20 $X=5.235 $Y=0.51
c435 42 0 3.223e-20 $X=4.805 $Y=0.51
r436 274 275 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=11.755
+ $Y=1.37 $X2=11.755 $Y2=1.37
r437 272 274 16.9718 $w=3.4e-07 $l=1e-07 $layer=POLY_cond $X=11.655 $Y=1.375
+ $X2=11.755 $Y2=1.375
r438 271 272 89.9507 $w=3.4e-07 $l=5.3e-07 $layer=POLY_cond $X=11.125 $Y=1.375
+ $X2=11.655 $Y2=1.375
r439 270 275 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=11.075 $Y=1.345
+ $X2=11.755 $Y2=1.345
r440 269 271 8.48592 $w=3.4e-07 $l=5e-08 $layer=POLY_cond $X=11.075 $Y=1.375
+ $X2=11.125 $Y2=1.375
r441 269 270 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.075
+ $Y=1.37 $X2=11.075 $Y2=1.37
r442 267 269 52.6127 $w=3.4e-07 $l=3.1e-07 $layer=POLY_cond $X=10.765 $Y=1.375
+ $X2=11.075 $Y2=1.375
r443 266 267 28.8521 $w=3.4e-07 $l=1.7e-07 $layer=POLY_cond $X=10.595 $Y=1.375
+ $X2=10.765 $Y2=1.375
r444 265 266 44.1268 $w=3.4e-07 $l=2.6e-07 $layer=POLY_cond $X=10.335 $Y=1.375
+ $X2=10.595 $Y2=1.375
r445 264 265 45.8239 $w=3.4e-07 $l=2.7e-07 $layer=POLY_cond $X=10.065 $Y=1.375
+ $X2=10.335 $Y2=1.375
r446 263 264 15.2746 $w=3.4e-07 $l=9e-08 $layer=POLY_cond $X=9.975 $Y=1.375
+ $X2=10.065 $Y2=1.375
r447 261 263 27.1549 $w=3.4e-07 $l=1.6e-07 $layer=POLY_cond $X=9.815 $Y=1.375
+ $X2=9.975 $Y2=1.375
r448 259 261 45.8239 $w=3.4e-07 $l=2.7e-07 $layer=POLY_cond $X=9.545 $Y=1.375
+ $X2=9.815 $Y2=1.375
r449 258 259 1.69718 $w=3.4e-07 $l=1e-08 $layer=POLY_cond $X=9.535 $Y=1.375
+ $X2=9.545 $Y2=1.375
r450 257 258 59.4014 $w=3.4e-07 $l=3.5e-07 $layer=POLY_cond $X=9.185 $Y=1.375
+ $X2=9.535 $Y2=1.375
r451 256 257 30.5493 $w=3.4e-07 $l=1.8e-07 $layer=POLY_cond $X=9.005 $Y=1.375
+ $X2=9.185 $Y2=1.375
r452 255 256 42.4296 $w=3.4e-07 $l=2.5e-07 $layer=POLY_cond $X=8.755 $Y=1.375
+ $X2=9.005 $Y2=1.375
r453 254 255 47.5211 $w=3.4e-07 $l=2.8e-07 $layer=POLY_cond $X=8.475 $Y=1.375
+ $X2=8.755 $Y2=1.375
r454 253 254 13.5775 $w=3.4e-07 $l=8e-08 $layer=POLY_cond $X=8.395 $Y=1.375
+ $X2=8.475 $Y2=1.375
r455 251 253 0.848592 $w=3.4e-07 $l=5e-09 $layer=POLY_cond $X=8.39 $Y=1.375
+ $X2=8.395 $Y2=1.375
r456 249 251 72.1303 $w=3.4e-07 $l=4.25e-07 $layer=POLY_cond $X=7.965 $Y=1.375
+ $X2=8.39 $Y2=1.375
r457 248 249 3.39437 $w=3.4e-07 $l=2e-08 $layer=POLY_cond $X=7.945 $Y=1.375
+ $X2=7.965 $Y2=1.375
r458 247 248 57.7042 $w=3.4e-07 $l=3.4e-07 $layer=POLY_cond $X=7.605 $Y=1.375
+ $X2=7.945 $Y2=1.375
r459 246 247 32.2465 $w=3.4e-07 $l=1.9e-07 $layer=POLY_cond $X=7.415 $Y=1.375
+ $X2=7.605 $Y2=1.375
r460 245 246 40.7324 $w=3.4e-07 $l=2.4e-07 $layer=POLY_cond $X=7.175 $Y=1.375
+ $X2=7.415 $Y2=1.375
r461 244 245 49.2183 $w=3.4e-07 $l=2.9e-07 $layer=POLY_cond $X=6.885 $Y=1.375
+ $X2=7.175 $Y2=1.375
r462 243 244 11.8803 $w=3.4e-07 $l=7e-08 $layer=POLY_cond $X=6.815 $Y=1.375
+ $X2=6.885 $Y2=1.375
r463 241 243 30.5493 $w=3.4e-07 $l=1.8e-07 $layer=POLY_cond $X=6.635 $Y=1.375
+ $X2=6.815 $Y2=1.375
r464 239 241 42.4296 $w=3.4e-07 $l=2.5e-07 $layer=POLY_cond $X=6.385 $Y=1.375
+ $X2=6.635 $Y2=1.375
r465 238 239 5.09155 $w=3.4e-07 $l=3e-08 $layer=POLY_cond $X=6.355 $Y=1.375
+ $X2=6.385 $Y2=1.375
r466 237 238 56.007 $w=3.4e-07 $l=3.3e-07 $layer=POLY_cond $X=6.025 $Y=1.375
+ $X2=6.355 $Y2=1.375
r467 236 237 33.9437 $w=3.4e-07 $l=2e-07 $layer=POLY_cond $X=5.825 $Y=1.375
+ $X2=6.025 $Y2=1.375
r468 235 236 39.0352 $w=3.4e-07 $l=2.3e-07 $layer=POLY_cond $X=5.595 $Y=1.375
+ $X2=5.825 $Y2=1.375
r469 234 235 50.9155 $w=3.4e-07 $l=3e-07 $layer=POLY_cond $X=5.295 $Y=1.375
+ $X2=5.595 $Y2=1.375
r470 233 234 10.1831 $w=3.4e-07 $l=6e-08 $layer=POLY_cond $X=5.235 $Y=1.375
+ $X2=5.295 $Y2=1.375
r471 231 233 1.69718 $w=3.4e-07 $l=1e-08 $layer=POLY_cond $X=5.225 $Y=1.375
+ $X2=5.235 $Y2=1.375
r472 231 232 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.225
+ $Y=1.37 $X2=5.225 $Y2=1.37
r473 229 231 71.2817 $w=3.4e-07 $l=4.2e-07 $layer=POLY_cond $X=4.805 $Y=1.375
+ $X2=5.225 $Y2=1.375
r474 228 229 6.78873 $w=3.4e-07 $l=4e-08 $layer=POLY_cond $X=4.765 $Y=1.375
+ $X2=4.805 $Y2=1.375
r475 227 228 54.3099 $w=3.4e-07 $l=3.2e-07 $layer=POLY_cond $X=4.445 $Y=1.375
+ $X2=4.765 $Y2=1.375
r476 226 227 35.6408 $w=3.4e-07 $l=2.1e-07 $layer=POLY_cond $X=4.235 $Y=1.375
+ $X2=4.445 $Y2=1.375
r477 225 226 37.338 $w=3.4e-07 $l=2.2e-07 $layer=POLY_cond $X=4.015 $Y=1.375
+ $X2=4.235 $Y2=1.375
r478 223 225 45.8239 $w=3.4e-07 $l=2.7e-07 $layer=POLY_cond $X=3.745 $Y=1.375
+ $X2=4.015 $Y2=1.375
r479 221 223 6.78873 $w=3.4e-07 $l=4e-08 $layer=POLY_cond $X=3.705 $Y=1.375
+ $X2=3.745 $Y2=1.375
r480 219 221 8.48592 $w=3.4e-07 $l=5e-08 $layer=POLY_cond $X=3.655 $Y=1.375
+ $X2=3.705 $Y2=1.375
r481 216 275 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.76 $Y=1.295
+ $X2=11.76 $Y2=1.295
r482 214 261 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.815
+ $Y=1.37 $X2=9.815 $Y2=1.37
r483 213 216 1.23188 $w=2.3e-07 $l=1.92e-06 $layer=MET1_cond $X=9.84 $Y=1.295
+ $X2=11.76 $Y2=1.295
r484 213 214 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=1.295
+ $X2=9.84 $Y2=1.295
r485 211 251 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=8.39
+ $Y=1.37 $X2=8.39 $Y2=1.37
r486 210 213 0.92391 $w=2.3e-07 $l=1.44e-06 $layer=MET1_cond $X=8.4 $Y=1.295
+ $X2=9.84 $Y2=1.295
r487 210 211 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.4 $Y=1.295
+ $X2=8.4 $Y2=1.295
r488 208 241 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.635
+ $Y=1.37 $X2=6.635 $Y2=1.37
r489 207 210 1.13243 $w=2.3e-07 $l=1.765e-06 $layer=MET1_cond $X=6.635 $Y=1.295
+ $X2=8.4 $Y2=1.295
r490 207 208 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.635 $Y=1.295
+ $X2=6.635 $Y2=1.295
r491 205 232 1.11436 $w=8.03e-07 $l=7.5e-08 $layer=LI1_cond $X=4.987 $Y=1.295
+ $X2=4.987 $Y2=1.37
r492 204 207 1.02336 $w=2.3e-07 $l=1.595e-06 $layer=MET1_cond $X=5.04 $Y=1.295
+ $X2=6.635 $Y2=1.295
r493 204 205 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=1.295
+ $X2=5.04 $Y2=1.295
r494 201 223 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.745
+ $Y=1.37 $X2=3.745 $Y2=1.37
r495 200 204 0.92391 $w=2.3e-07 $l=1.44e-06 $layer=MET1_cond $X=3.6 $Y=1.295
+ $X2=5.04 $Y2=1.295
r496 200 201 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=1.295
+ $X2=3.6 $Y2=1.295
r497 195 201 17.0432 $w=3.53e-07 $l=5.25e-07 $layer=LI1_cond $X=3.075 $Y=1.357
+ $X2=3.6 $Y2=1.357
r498 195 198 5.35643 $w=3.53e-07 $l=1.65e-07 $layer=LI1_cond $X=3.075 $Y=1.357
+ $X2=2.91 $Y2=1.357
r499 191 192 10.5802 $w=4.58e-07 $l=2.15e-07 $layer=LI1_cond $X=0.825 $Y=2.23
+ $X2=0.825 $Y2=2.015
r500 186 188 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=2.91 $Y=2.23
+ $X2=2.91 $Y2=2.91
r501 184 198 1.15789 $w=3.3e-07 $l=1.78e-07 $layer=LI1_cond $X=2.91 $Y=1.535
+ $X2=2.91 $Y2=1.357
r502 184 186 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=2.91 $Y=1.535
+ $X2=2.91 $Y2=2.23
r503 180 198 9.3494 $w=3.53e-07 $l=2.88e-07 $layer=LI1_cond $X=2.622 $Y=1.357
+ $X2=2.91 $Y2=1.357
r504 180 197 5.65824 $w=3.53e-07 $l=1.72e-07 $layer=LI1_cond $X=2.622 $Y=1.357
+ $X2=2.45 $Y2=1.357
r505 180 182 24.7191 $w=3.43e-07 $l=7.4e-07 $layer=LI1_cond $X=2.622 $Y=1.18
+ $X2=2.622 $Y2=0.44
r506 179 194 5.16603 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=2.015 $Y=1.37
+ $X2=1.85 $Y2=1.37
r507 179 197 15.1913 $w=3.28e-07 $l=4.35e-07 $layer=LI1_cond $X=2.015 $Y=1.37
+ $X2=2.45 $Y2=1.37
r508 174 176 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=1.85 $Y=2.23
+ $X2=1.85 $Y2=2.91
r509 172 194 1.34256 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=1.85 $Y=1.535
+ $X2=1.85 $Y2=1.37
r510 172 174 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=1.85 $Y=1.535
+ $X2=1.85 $Y2=2.23
r511 171 193 0.466467 $w=3.3e-07 $l=1.73e-07 $layer=LI1_cond $X=1.23 $Y=1.37
+ $X2=1.057 $Y2=1.37
r512 170 194 5.16603 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=1.685 $Y=1.37
+ $X2=1.85 $Y2=1.37
r513 170 171 15.8897 $w=3.28e-07 $l=4.55e-07 $layer=LI1_cond $X=1.685 $Y=1.37
+ $X2=1.23 $Y2=1.37
r514 168 193 6.31733 $w=2.57e-07 $l=2.03912e-07 $layer=LI1_cond $X=0.97 $Y=1.535
+ $X2=1.057 $Y2=1.37
r515 168 192 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=0.97 $Y=1.535
+ $X2=0.97 $Y2=2.015
r516 164 193 6.31733 $w=2.57e-07 $l=1.65e-07 $layer=LI1_cond $X=1.057 $Y=1.205
+ $X2=1.057 $Y2=1.37
r517 164 166 25.5542 $w=3.43e-07 $l=7.65e-07 $layer=LI1_cond $X=1.057 $Y=1.205
+ $X2=1.057 $Y2=0.44
r518 160 191 0.390026 $w=4.58e-07 $l=1.5e-08 $layer=LI1_cond $X=0.825 $Y=2.245
+ $X2=0.825 $Y2=2.23
r519 160 162 17.2911 $w=4.58e-07 $l=6.65e-07 $layer=LI1_cond $X=0.825 $Y=2.245
+ $X2=0.825 $Y2=2.91
r520 156 272 10.0333 $w=2.5e-07 $l=1.7e-07 $layer=POLY_cond $X=11.655 $Y=1.545
+ $X2=11.655 $Y2=1.375
r521 156 158 258.392 $w=2.5e-07 $l=1.04e-06 $layer=POLY_cond $X=11.655 $Y=1.545
+ $X2=11.655 $Y2=2.585
r522 152 271 21.9347 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=11.125 $Y=1.205
+ $X2=11.125 $Y2=1.375
r523 152 154 356.372 $w=1.5e-07 $l=6.95e-07 $layer=POLY_cond $X=11.125 $Y=1.205
+ $X2=11.125 $Y2=0.51
r524 148 271 10.0333 $w=2.5e-07 $l=1.7e-07 $layer=POLY_cond $X=11.125 $Y=1.545
+ $X2=11.125 $Y2=1.375
r525 148 150 258.392 $w=2.5e-07 $l=1.04e-06 $layer=POLY_cond $X=11.125 $Y=1.545
+ $X2=11.125 $Y2=2.585
r526 144 267 21.9347 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=10.765 $Y=1.205
+ $X2=10.765 $Y2=1.375
r527 144 146 356.372 $w=1.5e-07 $l=6.95e-07 $layer=POLY_cond $X=10.765 $Y=1.205
+ $X2=10.765 $Y2=0.51
r528 140 266 10.0333 $w=2.5e-07 $l=1.7e-07 $layer=POLY_cond $X=10.595 $Y=1.545
+ $X2=10.595 $Y2=1.375
r529 140 142 258.392 $w=2.5e-07 $l=1.04e-06 $layer=POLY_cond $X=10.595 $Y=1.545
+ $X2=10.595 $Y2=2.585
r530 136 265 21.9347 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=10.335 $Y=1.205
+ $X2=10.335 $Y2=1.375
r531 136 138 356.372 $w=1.5e-07 $l=6.95e-07 $layer=POLY_cond $X=10.335 $Y=1.205
+ $X2=10.335 $Y2=0.51
r532 132 264 10.0333 $w=2.5e-07 $l=1.7e-07 $layer=POLY_cond $X=10.065 $Y=1.545
+ $X2=10.065 $Y2=1.375
r533 132 134 258.392 $w=2.5e-07 $l=1.04e-06 $layer=POLY_cond $X=10.065 $Y=1.545
+ $X2=10.065 $Y2=2.585
r534 128 263 21.9347 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=9.975 $Y=1.205
+ $X2=9.975 $Y2=1.375
r535 128 130 356.372 $w=1.5e-07 $l=6.95e-07 $layer=POLY_cond $X=9.975 $Y=1.205
+ $X2=9.975 $Y2=0.51
r536 124 259 21.9347 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=9.545 $Y=1.205
+ $X2=9.545 $Y2=1.375
r537 124 126 356.372 $w=1.5e-07 $l=6.95e-07 $layer=POLY_cond $X=9.545 $Y=1.205
+ $X2=9.545 $Y2=0.51
r538 120 258 10.0333 $w=2.5e-07 $l=1.7e-07 $layer=POLY_cond $X=9.535 $Y=1.545
+ $X2=9.535 $Y2=1.375
r539 120 122 258.392 $w=2.5e-07 $l=1.04e-06 $layer=POLY_cond $X=9.535 $Y=1.545
+ $X2=9.535 $Y2=2.585
r540 116 257 21.9347 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=9.185 $Y=1.205
+ $X2=9.185 $Y2=1.375
r541 116 118 356.372 $w=1.5e-07 $l=6.95e-07 $layer=POLY_cond $X=9.185 $Y=1.205
+ $X2=9.185 $Y2=0.51
r542 112 256 10.0333 $w=2.5e-07 $l=1.7e-07 $layer=POLY_cond $X=9.005 $Y=1.545
+ $X2=9.005 $Y2=1.375
r543 112 114 258.392 $w=2.5e-07 $l=1.04e-06 $layer=POLY_cond $X=9.005 $Y=1.545
+ $X2=9.005 $Y2=2.585
r544 108 255 21.9347 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=8.755 $Y=1.205
+ $X2=8.755 $Y2=1.375
r545 108 110 356.372 $w=1.5e-07 $l=6.95e-07 $layer=POLY_cond $X=8.755 $Y=1.205
+ $X2=8.755 $Y2=0.51
r546 104 254 10.0333 $w=2.5e-07 $l=1.7e-07 $layer=POLY_cond $X=8.475 $Y=1.545
+ $X2=8.475 $Y2=1.375
r547 104 106 258.392 $w=2.5e-07 $l=1.04e-06 $layer=POLY_cond $X=8.475 $Y=1.545
+ $X2=8.475 $Y2=2.585
r548 100 253 21.9347 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=8.395 $Y=1.205
+ $X2=8.395 $Y2=1.375
r549 100 102 356.372 $w=1.5e-07 $l=6.95e-07 $layer=POLY_cond $X=8.395 $Y=1.205
+ $X2=8.395 $Y2=0.51
r550 96 249 21.9347 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=7.965 $Y=1.205
+ $X2=7.965 $Y2=1.375
r551 96 98 356.372 $w=1.5e-07 $l=6.95e-07 $layer=POLY_cond $X=7.965 $Y=1.205
+ $X2=7.965 $Y2=0.51
r552 92 248 10.0333 $w=2.5e-07 $l=1.7e-07 $layer=POLY_cond $X=7.945 $Y=1.545
+ $X2=7.945 $Y2=1.375
r553 92 94 258.392 $w=2.5e-07 $l=1.04e-06 $layer=POLY_cond $X=7.945 $Y=1.545
+ $X2=7.945 $Y2=2.585
r554 88 247 21.9347 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=7.605 $Y=1.205
+ $X2=7.605 $Y2=1.375
r555 88 90 356.372 $w=1.5e-07 $l=6.95e-07 $layer=POLY_cond $X=7.605 $Y=1.205
+ $X2=7.605 $Y2=0.51
r556 84 246 10.0333 $w=2.5e-07 $l=1.7e-07 $layer=POLY_cond $X=7.415 $Y=1.545
+ $X2=7.415 $Y2=1.375
r557 84 86 258.392 $w=2.5e-07 $l=1.04e-06 $layer=POLY_cond $X=7.415 $Y=1.545
+ $X2=7.415 $Y2=2.585
r558 80 245 21.9347 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=7.175 $Y=1.205
+ $X2=7.175 $Y2=1.375
r559 80 82 356.372 $w=1.5e-07 $l=6.95e-07 $layer=POLY_cond $X=7.175 $Y=1.205
+ $X2=7.175 $Y2=0.51
r560 76 244 10.0333 $w=2.5e-07 $l=1.7e-07 $layer=POLY_cond $X=6.885 $Y=1.545
+ $X2=6.885 $Y2=1.375
r561 76 78 258.392 $w=2.5e-07 $l=1.04e-06 $layer=POLY_cond $X=6.885 $Y=1.545
+ $X2=6.885 $Y2=2.585
r562 72 243 21.9347 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=6.815 $Y=1.205
+ $X2=6.815 $Y2=1.375
r563 72 74 356.372 $w=1.5e-07 $l=6.95e-07 $layer=POLY_cond $X=6.815 $Y=1.205
+ $X2=6.815 $Y2=0.51
r564 68 239 21.9347 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=6.385 $Y=1.205
+ $X2=6.385 $Y2=1.375
r565 68 70 356.372 $w=1.5e-07 $l=6.95e-07 $layer=POLY_cond $X=6.385 $Y=1.205
+ $X2=6.385 $Y2=0.51
r566 64 238 10.0333 $w=2.5e-07 $l=1.7e-07 $layer=POLY_cond $X=6.355 $Y=1.545
+ $X2=6.355 $Y2=1.375
r567 64 66 258.392 $w=2.5e-07 $l=1.04e-06 $layer=POLY_cond $X=6.355 $Y=1.545
+ $X2=6.355 $Y2=2.585
r568 60 237 21.9347 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=6.025 $Y=1.205
+ $X2=6.025 $Y2=1.375
r569 60 62 356.372 $w=1.5e-07 $l=6.95e-07 $layer=POLY_cond $X=6.025 $Y=1.205
+ $X2=6.025 $Y2=0.51
r570 56 236 10.0333 $w=2.5e-07 $l=1.7e-07 $layer=POLY_cond $X=5.825 $Y=1.545
+ $X2=5.825 $Y2=1.375
r571 56 58 258.392 $w=2.5e-07 $l=1.04e-06 $layer=POLY_cond $X=5.825 $Y=1.545
+ $X2=5.825 $Y2=2.585
r572 52 235 21.9347 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=5.595 $Y=1.205
+ $X2=5.595 $Y2=1.375
r573 52 54 356.372 $w=1.5e-07 $l=6.95e-07 $layer=POLY_cond $X=5.595 $Y=1.205
+ $X2=5.595 $Y2=0.51
r574 48 234 10.0333 $w=2.5e-07 $l=1.7e-07 $layer=POLY_cond $X=5.295 $Y=1.545
+ $X2=5.295 $Y2=1.375
r575 48 50 258.392 $w=2.5e-07 $l=1.04e-06 $layer=POLY_cond $X=5.295 $Y=1.545
+ $X2=5.295 $Y2=2.585
r576 44 233 21.9347 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=5.235 $Y=1.205
+ $X2=5.235 $Y2=1.375
r577 44 46 356.372 $w=1.5e-07 $l=6.95e-07 $layer=POLY_cond $X=5.235 $Y=1.205
+ $X2=5.235 $Y2=0.51
r578 40 229 21.9347 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=4.805 $Y=1.205
+ $X2=4.805 $Y2=1.375
r579 40 42 356.372 $w=1.5e-07 $l=6.95e-07 $layer=POLY_cond $X=4.805 $Y=1.205
+ $X2=4.805 $Y2=0.51
r580 36 228 10.0333 $w=2.5e-07 $l=1.7e-07 $layer=POLY_cond $X=4.765 $Y=1.545
+ $X2=4.765 $Y2=1.375
r581 36 38 258.392 $w=2.5e-07 $l=1.04e-06 $layer=POLY_cond $X=4.765 $Y=1.545
+ $X2=4.765 $Y2=2.585
r582 32 227 21.9347 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=4.445 $Y=1.205
+ $X2=4.445 $Y2=1.375
r583 32 34 356.372 $w=1.5e-07 $l=6.95e-07 $layer=POLY_cond $X=4.445 $Y=1.205
+ $X2=4.445 $Y2=0.51
r584 28 226 10.0333 $w=2.5e-07 $l=1.7e-07 $layer=POLY_cond $X=4.235 $Y=1.545
+ $X2=4.235 $Y2=1.375
r585 28 30 258.392 $w=2.5e-07 $l=1.04e-06 $layer=POLY_cond $X=4.235 $Y=1.545
+ $X2=4.235 $Y2=2.585
r586 24 225 21.9347 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=4.015 $Y=1.205
+ $X2=4.015 $Y2=1.375
r587 24 26 356.372 $w=1.5e-07 $l=6.95e-07 $layer=POLY_cond $X=4.015 $Y=1.205
+ $X2=4.015 $Y2=0.51
r588 20 221 10.0333 $w=2.5e-07 $l=1.7e-07 $layer=POLY_cond $X=3.705 $Y=1.545
+ $X2=3.705 $Y2=1.375
r589 20 22 258.392 $w=2.5e-07 $l=1.04e-06 $layer=POLY_cond $X=3.705 $Y=1.545
+ $X2=3.705 $Y2=2.585
r590 16 219 21.9347 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=3.655 $Y=1.205
+ $X2=3.655 $Y2=1.375
r591 16 18 356.372 $w=1.5e-07 $l=6.95e-07 $layer=POLY_cond $X=3.655 $Y=1.205
+ $X2=3.655 $Y2=0.51
r592 5 188 400 $w=1.7e-07 $l=8.92258e-07 $layer=licon1_PDIFF $count=1 $X=2.77
+ $Y=2.085 $X2=2.91 $Y2=2.91
r593 5 186 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.77
+ $Y=2.085 $X2=2.91 $Y2=2.23
r594 4 176 400 $w=1.7e-07 $l=8.92258e-07 $layer=licon1_PDIFF $count=1 $X=1.71
+ $Y=2.085 $X2=1.85 $Y2=2.91
r595 4 174 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.71
+ $Y=2.085 $X2=1.85 $Y2=2.23
r596 3 191 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.65
+ $Y=2.085 $X2=0.79 $Y2=2.23
r597 3 162 400 $w=1.7e-07 $l=8.92258e-07 $layer=licon1_PDIFF $count=1 $X=0.65
+ $Y=2.085 $X2=0.79 $Y2=2.91
r598 2 182 182 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_NDIFF $count=1 $X=2.49
+ $Y=0.235 $X2=2.63 $Y2=0.44
r599 1 166 182 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_NDIFF $count=1 $X=0.91
+ $Y=0.235 $X2=1.05 $Y2=0.44
.ends

.subckt PM_SKY130_FD_SC_LP__CLKBUFLP_16%VPWR 1 2 3 4 5 6 7 8 9 10 11 12 37 39 45
+ 51 57 63 69 73 77 83 89 95 101 105 109 114 115 117 118 120 121 123 124 126 127
+ 128 140 144 156 160 167 168 174 177 180 183 186 189
r214 189 190 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.76 $Y=3.33
+ $X2=11.76 $Y2=3.33
r215 187 190 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=10.8 $Y=3.33
+ $X2=11.76 $Y2=3.33
r216 186 187 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=3.33
+ $X2=10.8 $Y2=3.33
r217 183 184 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r218 180 181 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r219 177 178 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r220 174 175 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r221 171 172 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r222 168 190 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.24 $Y=3.33
+ $X2=11.76 $Y2=3.33
r223 167 168 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.24 $Y=3.33
+ $X2=12.24 $Y2=3.33
r224 165 189 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.085 $Y=3.33
+ $X2=11.92 $Y2=3.33
r225 165 167 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=12.085 $Y=3.33
+ $X2=12.24 $Y2=3.33
r226 164 187 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=3.33
+ $X2=10.8 $Y2=3.33
r227 164 184 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=3.33
+ $X2=9.84 $Y2=3.33
r228 163 164 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.32 $Y=3.33
+ $X2=10.32 $Y2=3.33
r229 161 183 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.965 $Y=3.33
+ $X2=9.8 $Y2=3.33
r230 161 163 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=9.965 $Y=3.33
+ $X2=10.32 $Y2=3.33
r231 160 186 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.695 $Y=3.33
+ $X2=10.86 $Y2=3.33
r232 160 163 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=10.695 $Y=3.33
+ $X2=10.32 $Y2=3.33
r233 159 184 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=9.84 $Y2=3.33
r234 158 159 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r235 156 183 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.635 $Y=3.33
+ $X2=9.8 $Y2=3.33
r236 156 158 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=9.635 $Y=3.33
+ $X2=9.36 $Y2=3.33
r237 155 159 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=9.36 $Y2=3.33
r238 154 155 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r239 152 155 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=8.4 $Y2=3.33
r240 152 181 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=6.48 $Y2=3.33
r241 151 152 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r242 149 180 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.785 $Y=3.33
+ $X2=6.62 $Y2=3.33
r243 149 151 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=6.785 $Y=3.33
+ $X2=7.44 $Y2=3.33
r244 148 178 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=5.52 $Y2=3.33
r245 148 175 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=4.56 $Y2=3.33
r246 147 148 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r247 145 174 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.665 $Y=3.33
+ $X2=4.5 $Y2=3.33
r248 145 147 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=4.665 $Y=3.33
+ $X2=5.04 $Y2=3.33
r249 144 177 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.395 $Y=3.33
+ $X2=5.56 $Y2=3.33
r250 144 147 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=5.395 $Y=3.33
+ $X2=5.04 $Y2=3.33
r251 143 175 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r252 142 143 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r253 140 174 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.335 $Y=3.33
+ $X2=4.5 $Y2=3.33
r254 140 142 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=4.335 $Y=3.33
+ $X2=4.08 $Y2=3.33
r255 139 143 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=4.08 $Y2=3.33
r256 138 139 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r257 136 139 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r258 135 136 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r259 133 136 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r260 133 172 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.24 $Y2=3.33
r261 132 133 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r262 130 171 4.78091 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=3.33
+ $X2=0.212 $Y2=3.33
r263 130 132 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=0.425 $Y=3.33
+ $X2=1.2 $Y2=3.33
r264 128 181 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=6.24 $Y=3.33
+ $X2=6.48 $Y2=3.33
r265 128 178 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=6.24 $Y=3.33
+ $X2=5.52 $Y2=3.33
r266 126 154 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=8.575 $Y=3.33
+ $X2=8.4 $Y2=3.33
r267 126 127 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.575 $Y=3.33
+ $X2=8.74 $Y2=3.33
r268 125 158 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=8.905 $Y=3.33
+ $X2=9.36 $Y2=3.33
r269 125 127 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.905 $Y=3.33
+ $X2=8.74 $Y2=3.33
r270 123 151 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=7.515 $Y=3.33
+ $X2=7.44 $Y2=3.33
r271 123 124 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.515 $Y=3.33
+ $X2=7.68 $Y2=3.33
r272 122 154 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=7.845 $Y=3.33
+ $X2=8.4 $Y2=3.33
r273 122 124 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.845 $Y=3.33
+ $X2=7.68 $Y2=3.33
r274 120 138 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=3.275 $Y=3.33
+ $X2=3.12 $Y2=3.33
r275 120 121 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.275 $Y=3.33
+ $X2=3.44 $Y2=3.33
r276 119 142 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=3.605 $Y=3.33
+ $X2=4.08 $Y2=3.33
r277 119 121 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.605 $Y=3.33
+ $X2=3.44 $Y2=3.33
r278 117 135 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=2.215 $Y=3.33
+ $X2=2.16 $Y2=3.33
r279 117 118 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.215 $Y=3.33
+ $X2=2.38 $Y2=3.33
r280 116 138 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=2.545 $Y=3.33
+ $X2=3.12 $Y2=3.33
r281 116 118 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.545 $Y=3.33
+ $X2=2.38 $Y2=3.33
r282 114 132 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=1.225 $Y=3.33
+ $X2=1.2 $Y2=3.33
r283 114 115 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.225 $Y=3.33
+ $X2=1.355 $Y2=3.33
r284 113 135 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=1.485 $Y=3.33
+ $X2=2.16 $Y2=3.33
r285 113 115 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.485 $Y=3.33
+ $X2=1.355 $Y2=3.33
r286 109 112 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=11.92 $Y=2.23
+ $X2=11.92 $Y2=2.91
r287 107 189 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=11.92 $Y=3.245
+ $X2=11.92 $Y2=3.33
r288 107 112 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=11.92 $Y=3.245
+ $X2=11.92 $Y2=2.91
r289 106 186 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.025 $Y=3.33
+ $X2=10.86 $Y2=3.33
r290 105 189 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.755 $Y=3.33
+ $X2=11.92 $Y2=3.33
r291 105 106 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=11.755 $Y=3.33
+ $X2=11.025 $Y2=3.33
r292 101 104 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=10.86 $Y=2.23
+ $X2=10.86 $Y2=2.91
r293 99 186 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.86 $Y=3.245
+ $X2=10.86 $Y2=3.33
r294 99 104 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=10.86 $Y=3.245
+ $X2=10.86 $Y2=2.91
r295 95 98 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=9.8 $Y=2.23 $X2=9.8
+ $Y2=2.91
r296 93 183 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.8 $Y=3.245
+ $X2=9.8 $Y2=3.33
r297 93 98 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=9.8 $Y=3.245
+ $X2=9.8 $Y2=2.91
r298 89 92 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=8.74 $Y=2.23
+ $X2=8.74 $Y2=2.91
r299 87 127 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.74 $Y=3.245
+ $X2=8.74 $Y2=3.33
r300 87 92 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=8.74 $Y=3.245
+ $X2=8.74 $Y2=2.91
r301 83 86 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=7.68 $Y=2.23
+ $X2=7.68 $Y2=2.91
r302 81 124 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.68 $Y=3.245
+ $X2=7.68 $Y2=3.33
r303 81 86 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=7.68 $Y=3.245
+ $X2=7.68 $Y2=2.91
r304 77 80 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=6.62 $Y=2.23
+ $X2=6.62 $Y2=2.91
r305 75 180 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.62 $Y=3.245
+ $X2=6.62 $Y2=3.33
r306 75 80 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=6.62 $Y=3.245
+ $X2=6.62 $Y2=2.91
r307 74 177 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.725 $Y=3.33
+ $X2=5.56 $Y2=3.33
r308 73 180 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.455 $Y=3.33
+ $X2=6.62 $Y2=3.33
r309 73 74 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=6.455 $Y=3.33
+ $X2=5.725 $Y2=3.33
r310 69 72 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=5.56 $Y=2.23
+ $X2=5.56 $Y2=2.91
r311 67 177 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.56 $Y=3.245
+ $X2=5.56 $Y2=3.33
r312 67 72 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=5.56 $Y=3.245
+ $X2=5.56 $Y2=2.91
r313 63 66 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=4.5 $Y=2.23 $X2=4.5
+ $Y2=2.91
r314 61 174 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.5 $Y=3.245
+ $X2=4.5 $Y2=3.33
r315 61 66 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=4.5 $Y=3.245
+ $X2=4.5 $Y2=2.91
r316 57 60 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=3.44 $Y=2.23
+ $X2=3.44 $Y2=2.91
r317 55 121 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.44 $Y=3.245
+ $X2=3.44 $Y2=3.33
r318 55 60 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=3.44 $Y=3.245
+ $X2=3.44 $Y2=2.91
r319 51 54 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=2.38 $Y=2.23
+ $X2=2.38 $Y2=2.91
r320 49 118 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.38 $Y=3.245
+ $X2=2.38 $Y2=3.33
r321 49 54 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=2.38 $Y=3.245
+ $X2=2.38 $Y2=2.91
r322 45 48 30.1408 $w=2.58e-07 $l=6.8e-07 $layer=LI1_cond $X=1.355 $Y=2.23
+ $X2=1.355 $Y2=2.91
r323 43 115 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=1.355 $Y=3.245
+ $X2=1.355 $Y2=3.33
r324 43 48 14.8488 $w=2.58e-07 $l=3.35e-07 $layer=LI1_cond $X=1.355 $Y=3.245
+ $X2=1.355 $Y2=2.91
r325 39 42 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=0.26 $Y=2.23
+ $X2=0.26 $Y2=2.91
r326 37 171 2.98526 $w=3.3e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.26 $Y=3.245
+ $X2=0.212 $Y2=3.33
r327 37 42 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=0.26 $Y=3.245
+ $X2=0.26 $Y2=2.91
r328 12 112 400 $w=1.7e-07 $l=8.92258e-07 $layer=licon1_PDIFF $count=1 $X=11.78
+ $Y=2.085 $X2=11.92 $Y2=2.91
r329 12 109 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=11.78
+ $Y=2.085 $X2=11.92 $Y2=2.23
r330 11 104 400 $w=1.7e-07 $l=8.92258e-07 $layer=licon1_PDIFF $count=1 $X=10.72
+ $Y=2.085 $X2=10.86 $Y2=2.91
r331 11 101 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=10.72
+ $Y=2.085 $X2=10.86 $Y2=2.23
r332 10 98 400 $w=1.7e-07 $l=8.92258e-07 $layer=licon1_PDIFF $count=1 $X=9.66
+ $Y=2.085 $X2=9.8 $Y2=2.91
r333 10 95 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=9.66
+ $Y=2.085 $X2=9.8 $Y2=2.23
r334 9 92 400 $w=1.7e-07 $l=8.92258e-07 $layer=licon1_PDIFF $count=1 $X=8.6
+ $Y=2.085 $X2=8.74 $Y2=2.91
r335 9 89 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=8.6
+ $Y=2.085 $X2=8.74 $Y2=2.23
r336 8 86 400 $w=1.7e-07 $l=8.92258e-07 $layer=licon1_PDIFF $count=1 $X=7.54
+ $Y=2.085 $X2=7.68 $Y2=2.91
r337 8 83 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=7.54
+ $Y=2.085 $X2=7.68 $Y2=2.23
r338 7 80 400 $w=1.7e-07 $l=8.92258e-07 $layer=licon1_PDIFF $count=1 $X=6.48
+ $Y=2.085 $X2=6.62 $Y2=2.91
r339 7 77 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=6.48
+ $Y=2.085 $X2=6.62 $Y2=2.23
r340 6 72 400 $w=1.7e-07 $l=8.92258e-07 $layer=licon1_PDIFF $count=1 $X=5.42
+ $Y=2.085 $X2=5.56 $Y2=2.91
r341 6 69 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=5.42
+ $Y=2.085 $X2=5.56 $Y2=2.23
r342 5 66 400 $w=1.7e-07 $l=8.92258e-07 $layer=licon1_PDIFF $count=1 $X=4.36
+ $Y=2.085 $X2=4.5 $Y2=2.91
r343 5 63 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=4.36
+ $Y=2.085 $X2=4.5 $Y2=2.23
r344 4 60 400 $w=1.7e-07 $l=8.92258e-07 $layer=licon1_PDIFF $count=1 $X=3.3
+ $Y=2.085 $X2=3.44 $Y2=2.91
r345 4 57 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=3.3
+ $Y=2.085 $X2=3.44 $Y2=2.23
r346 3 54 400 $w=1.7e-07 $l=8.92258e-07 $layer=licon1_PDIFF $count=1 $X=2.24
+ $Y=2.085 $X2=2.38 $Y2=2.91
r347 3 51 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.24
+ $Y=2.085 $X2=2.38 $Y2=2.23
r348 2 48 400 $w=1.7e-07 $l=8.92258e-07 $layer=licon1_PDIFF $count=1 $X=1.18
+ $Y=2.085 $X2=1.32 $Y2=2.91
r349 2 45 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.18
+ $Y=2.085 $X2=1.32 $Y2=2.23
r350 1 42 400 $w=1.7e-07 $l=8.85297e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.085 $X2=0.26 $Y2=2.91
r351 1 39 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.085 $X2=0.26 $Y2=2.23
.ends

.subckt PM_SKY130_FD_SC_LP__CLKBUFLP_16%X 1 2 3 4 5 6 7 8 9 10 11 12 13 42 45 48
+ 52 56 60 67 70 73 76 81 82 85 93 102 110 118 127 135 143 144
c238 81 0 3.2513e-20 $X=10.44 $Y=1.79
c239 76 0 8.52417e-20 $X=9.27 $Y=1.48
c240 73 0 3.40562e-20 $X=7.27 $Y=1.79
c241 70 0 4.0915e-20 $X=5.95 $Y=1.79
c242 45 0 3.223e-20 $X=4.237 $Y=1.705
r243 147 149 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=11.39 $Y=2.23
+ $X2=11.39 $Y2=2.91
r244 143 147 6.80989 $w=3.28e-07 $l=1.95e-07 $layer=LI1_cond $X=11.39 $Y=2.035
+ $X2=11.39 $Y2=2.23
r245 143 144 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.39 $Y=2.035
+ $X2=11.39 $Y2=2.035
r246 138 140 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=10.33 $Y=2.23
+ $X2=10.33 $Y2=2.91
r247 136 144 0.686517 $w=2.3e-07 $l=1.07e-06 $layer=MET1_cond $X=10.32 $Y=2.035
+ $X2=11.39 $Y2=2.035
r248 135 138 6.80989 $w=3.28e-07 $l=1.95e-07 $layer=LI1_cond $X=10.33 $Y=2.035
+ $X2=10.33 $Y2=2.23
r249 135 136 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.32 $Y=2.035
+ $X2=10.32 $Y2=2.035
r250 130 132 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=9.27 $Y=2.23
+ $X2=9.27 $Y2=2.91
r251 128 136 0.670477 $w=2.3e-07 $l=1.045e-06 $layer=MET1_cond $X=9.275 $Y=2.035
+ $X2=10.32 $Y2=2.035
r252 127 130 6.80989 $w=3.28e-07 $l=1.95e-07 $layer=LI1_cond $X=9.27 $Y=2.035
+ $X2=9.27 $Y2=2.23
r253 127 128 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.275 $Y=2.035
+ $X2=9.275 $Y2=2.035
r254 122 124 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=8.21 $Y=2.23
+ $X2=8.21 $Y2=2.91
r255 119 128 0.680101 $w=2.3e-07 $l=1.06e-06 $layer=MET1_cond $X=8.215 $Y=2.035
+ $X2=9.275 $Y2=2.035
r256 118 122 6.80989 $w=3.28e-07 $l=1.95e-07 $layer=LI1_cond $X=8.21 $Y=2.035
+ $X2=8.21 $Y2=2.23
r257 118 119 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.215 $Y=2.035
+ $X2=8.215 $Y2=2.035
r258 113 115 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=7.15 $Y=2.23
+ $X2=7.15 $Y2=2.91
r259 110 113 6.80989 $w=3.28e-07 $l=1.95e-07 $layer=LI1_cond $X=7.15 $Y=2.035
+ $X2=7.15 $Y2=2.23
r260 110 111 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.155 $Y=2.035
+ $X2=7.155 $Y2=2.035
r261 105 107 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=6.09 $Y=2.23
+ $X2=6.09 $Y2=2.91
r262 103 111 0.683309 $w=2.3e-07 $l=1.065e-06 $layer=MET1_cond $X=6.09 $Y=2.035
+ $X2=7.155 $Y2=2.035
r263 102 105 6.80989 $w=3.28e-07 $l=1.95e-07 $layer=LI1_cond $X=6.09 $Y=2.035
+ $X2=6.09 $Y2=2.23
r264 102 103 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.09 $Y=2.035
+ $X2=6.09 $Y2=2.035
r265 97 99 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=5.03 $Y=2.23
+ $X2=5.03 $Y2=2.91
r266 94 103 0.673685 $w=2.3e-07 $l=1.05e-06 $layer=MET1_cond $X=5.04 $Y=2.035
+ $X2=6.09 $Y2=2.035
r267 93 97 6.80989 $w=3.28e-07 $l=1.95e-07 $layer=LI1_cond $X=5.03 $Y=2.035
+ $X2=5.03 $Y2=2.23
r268 93 94 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=2.035
+ $X2=5.04 $Y2=2.035
r269 88 90 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=3.97 $Y=2.23
+ $X2=3.97 $Y2=2.91
r270 86 94 0.686517 $w=2.3e-07 $l=1.07e-06 $layer=MET1_cond $X=3.97 $Y=2.035
+ $X2=5.04 $Y2=2.035
r271 85 88 6.80989 $w=3.28e-07 $l=1.95e-07 $layer=LI1_cond $X=3.97 $Y=2.035
+ $X2=3.97 $Y2=2.23
r272 85 86 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.97 $Y=2.035
+ $X2=3.97 $Y2=2.035
r273 82 119 0.343258 $w=2.3e-07 $l=5.35e-07 $layer=MET1_cond $X=7.68 $Y=2.035
+ $X2=8.215 $Y2=2.035
r274 82 111 0.336842 $w=2.3e-07 $l=5.25e-07 $layer=MET1_cond $X=7.68 $Y=2.035
+ $X2=7.155 $Y2=2.035
r275 81 135 8.55602 $w=3.28e-07 $l=2.45e-07 $layer=LI1_cond $X=10.33 $Y=1.79
+ $X2=10.33 $Y2=2.035
r276 80 81 13.4831 $w=5.48e-07 $l=6.2e-07 $layer=LI1_cond $X=10.44 $Y=1.17
+ $X2=10.44 $Y2=1.79
r277 77 127 8.55602 $w=3.28e-07 $l=2.45e-07 $layer=LI1_cond $X=9.27 $Y=1.79
+ $X2=9.27 $Y2=2.035
r278 76 77 4.43028 $w=3.3e-07 $l=3.1e-07 $layer=LI1_cond $X=9.27 $Y=1.48
+ $X2=9.27 $Y2=1.79
r279 74 76 5.78748 $w=6.18e-07 $l=3e-07 $layer=LI1_cond $X=8.97 $Y=1.48 $X2=9.27
+ $Y2=1.48
r280 73 110 8.55602 $w=3.28e-07 $l=2.45e-07 $layer=LI1_cond $X=7.15 $Y=1.79
+ $X2=7.15 $Y2=2.035
r281 72 73 13.01 $w=5.68e-07 $l=6.2e-07 $layer=LI1_cond $X=7.27 $Y=1.17 $X2=7.27
+ $Y2=1.79
r282 70 102 8.55602 $w=3.28e-07 $l=2.45e-07 $layer=LI1_cond $X=6.09 $Y=1.79
+ $X2=6.09 $Y2=2.035
r283 69 70 12.1569 $w=6.08e-07 $l=6.2e-07 $layer=LI1_cond $X=5.95 $Y=1.17
+ $X2=5.95 $Y2=1.79
r284 63 85 5.5876 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=3.97 $Y=1.875
+ $X2=3.97 $Y2=2.035
r285 60 80 25.4934 $w=3.28e-07 $l=7.3e-07 $layer=LI1_cond $X=10.55 $Y=0.44
+ $X2=10.55 $Y2=1.17
r286 54 74 4.43028 $w=3.3e-07 $l=3.1e-07 $layer=LI1_cond $X=8.97 $Y=1.17
+ $X2=8.97 $Y2=1.48
r287 54 56 25.4934 $w=3.28e-07 $l=7.3e-07 $layer=LI1_cond $X=8.97 $Y=1.17
+ $X2=8.97 $Y2=0.44
r288 52 72 25.4934 $w=3.28e-07 $l=7.3e-07 $layer=LI1_cond $X=7.39 $Y=0.44
+ $X2=7.39 $Y2=1.17
r289 48 69 25.4934 $w=3.28e-07 $l=7.3e-07 $layer=LI1_cond $X=5.81 $Y=0.44
+ $X2=5.81 $Y2=1.17
r290 45 63 17.4193 $w=1.68e-07 $l=2.67e-07 $layer=LI1_cond $X=4.237 $Y=1.79
+ $X2=3.97 $Y2=1.79
r291 45 67 24.5123 $w=3.13e-07 $l=6.7e-07 $layer=LI1_cond $X=4.237 $Y=1.705
+ $X2=4.237 $Y2=1.035
r292 40 67 5.76222 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=4.23 $Y=0.87
+ $X2=4.23 $Y2=1.035
r293 40 42 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=4.23 $Y=0.87
+ $X2=4.23 $Y2=0.44
r294 13 149 400 $w=1.7e-07 $l=8.92258e-07 $layer=licon1_PDIFF $count=1 $X=11.25
+ $Y=2.085 $X2=11.39 $Y2=2.91
r295 13 147 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=11.25
+ $Y=2.085 $X2=11.39 $Y2=2.23
r296 12 140 400 $w=1.7e-07 $l=8.92258e-07 $layer=licon1_PDIFF $count=1 $X=10.19
+ $Y=2.085 $X2=10.33 $Y2=2.91
r297 12 138 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=10.19
+ $Y=2.085 $X2=10.33 $Y2=2.23
r298 11 132 400 $w=1.7e-07 $l=8.92258e-07 $layer=licon1_PDIFF $count=1 $X=9.13
+ $Y=2.085 $X2=9.27 $Y2=2.91
r299 11 130 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=9.13
+ $Y=2.085 $X2=9.27 $Y2=2.23
r300 10 124 400 $w=1.7e-07 $l=8.92258e-07 $layer=licon1_PDIFF $count=1 $X=8.07
+ $Y=2.085 $X2=8.21 $Y2=2.91
r301 10 122 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=8.07
+ $Y=2.085 $X2=8.21 $Y2=2.23
r302 9 115 400 $w=1.7e-07 $l=8.92258e-07 $layer=licon1_PDIFF $count=1 $X=7.01
+ $Y=2.085 $X2=7.15 $Y2=2.91
r303 9 113 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=7.01
+ $Y=2.085 $X2=7.15 $Y2=2.23
r304 8 107 400 $w=1.7e-07 $l=8.92258e-07 $layer=licon1_PDIFF $count=1 $X=5.95
+ $Y=2.085 $X2=6.09 $Y2=2.91
r305 8 105 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=5.95
+ $Y=2.085 $X2=6.09 $Y2=2.23
r306 7 99 400 $w=1.7e-07 $l=8.92258e-07 $layer=licon1_PDIFF $count=1 $X=4.89
+ $Y=2.085 $X2=5.03 $Y2=2.91
r307 7 97 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=4.89
+ $Y=2.085 $X2=5.03 $Y2=2.23
r308 6 90 400 $w=1.7e-07 $l=8.92258e-07 $layer=licon1_PDIFF $count=1 $X=3.83
+ $Y=2.085 $X2=3.97 $Y2=2.91
r309 6 88 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=3.83
+ $Y=2.085 $X2=3.97 $Y2=2.23
r310 5 60 182 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_NDIFF $count=1 $X=10.41
+ $Y=0.235 $X2=10.55 $Y2=0.44
r311 4 56 182 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_NDIFF $count=1 $X=8.83
+ $Y=0.235 $X2=8.97 $Y2=0.44
r312 3 52 182 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_NDIFF $count=1 $X=7.25
+ $Y=0.235 $X2=7.39 $Y2=0.44
r313 2 48 182 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_NDIFF $count=1 $X=5.67
+ $Y=0.235 $X2=5.81 $Y2=0.44
r314 1 42 182 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_NDIFF $count=1 $X=4.09
+ $Y=0.235 $X2=4.23 $Y2=0.44
.ends

.subckt PM_SKY130_FD_SC_LP__CLKBUFLP_16%VGND 1 2 3 4 5 6 7 8 25 27 31 35 39 43
+ 47 51 55 58 59 61 62 63 65 77 84 96 103 110 111 117 120 123 126 129
r181 129 130 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.28 $Y=0
+ $X2=11.28 $Y2=0
r182 126 127 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=0
+ $X2=9.84 $Y2=0
r183 123 124 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.48 $Y=0
+ $X2=6.48 $Y2=0
r184 120 121 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0
+ $X2=5.04 $Y2=0
r185 117 118 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0
+ $X2=1.68 $Y2=0
r186 114 115 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0
+ $X2=0.24 $Y2=0
r187 111 130 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=12.24 $Y=0
+ $X2=11.28 $Y2=0
r188 110 111 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=12.24 $Y=0
+ $X2=12.24 $Y2=0
r189 108 129 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.505 $Y=0
+ $X2=11.34 $Y2=0
r190 108 110 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=11.505 $Y=0
+ $X2=12.24 $Y2=0
r191 107 130 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.8 $Y=0
+ $X2=11.28 $Y2=0
r192 107 127 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=10.8 $Y=0
+ $X2=9.84 $Y2=0
r193 106 107 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.8 $Y=0
+ $X2=10.8 $Y2=0
r194 104 126 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.925 $Y=0
+ $X2=9.76 $Y2=0
r195 104 106 57.0856 $w=1.68e-07 $l=8.75e-07 $layer=LI1_cond $X=9.925 $Y=0
+ $X2=10.8 $Y2=0
r196 103 129 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.175 $Y=0
+ $X2=11.34 $Y2=0
r197 103 106 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=11.175 $Y=0
+ $X2=10.8 $Y2=0
r198 102 127 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=0
+ $X2=9.84 $Y2=0
r199 101 102 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=9.36 $Y=0
+ $X2=9.36 $Y2=0
r200 99 102 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=8.4 $Y=0 $X2=9.36
+ $Y2=0
r201 98 101 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=8.4 $Y=0 $X2=9.36
+ $Y2=0
r202 98 99 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r203 96 126 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.595 $Y=0
+ $X2=9.76 $Y2=0
r204 96 101 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=9.595 $Y=0
+ $X2=9.36 $Y2=0
r205 95 99 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=8.4
+ $Y2=0
r206 94 95 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r207 92 95 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=7.92
+ $Y2=0
r208 92 124 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0
+ $X2=6.48 $Y2=0
r209 91 94 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=6.96 $Y=0 $X2=7.92
+ $Y2=0
r210 91 92 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r211 89 123 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.765 $Y=0 $X2=6.6
+ $Y2=0
r212 89 91 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=6.765 $Y=0
+ $X2=6.96 $Y2=0
r213 88 121 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0
+ $X2=5.04 $Y2=0
r214 87 88 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r215 85 120 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.185 $Y=0
+ $X2=5.02 $Y2=0
r216 85 87 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=5.185 $Y=0
+ $X2=5.52 $Y2=0
r217 84 123 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.435 $Y=0 $X2=6.6
+ $Y2=0
r218 84 87 59.6952 $w=1.68e-07 $l=9.15e-07 $layer=LI1_cond $X=6.435 $Y=0
+ $X2=5.52 $Y2=0
r219 83 121 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0
+ $X2=5.04 $Y2=0
r220 82 83 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r221 80 83 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.56
+ $Y2=0
r222 79 82 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=3.6 $Y=0 $X2=4.56
+ $Y2=0
r223 79 80 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r224 77 120 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.855 $Y=0
+ $X2=5.02 $Y2=0
r225 77 82 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=4.855 $Y=0 $X2=4.56
+ $Y2=0
r226 76 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r227 75 76 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r228 73 76 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r229 73 118 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0
+ $X2=1.68 $Y2=0
r230 72 75 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r231 72 73 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r232 70 117 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.005 $Y=0
+ $X2=1.84 $Y2=0
r233 70 72 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=2.005 $Y=0
+ $X2=2.16 $Y2=0
r234 69 118 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0
+ $X2=1.68 $Y2=0
r235 69 115 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0
+ $X2=0.24 $Y2=0
r236 68 69 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r237 66 114 4.43563 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=0
+ $X2=0.212 $Y2=0
r238 66 68 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.425 $Y=0 $X2=0.72
+ $Y2=0
r239 65 117 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.675 $Y=0
+ $X2=1.84 $Y2=0
r240 65 68 62.3048 $w=1.68e-07 $l=9.55e-07 $layer=LI1_cond $X=1.675 $Y=0
+ $X2=0.72 $Y2=0
r241 63 124 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=6.24 $Y=0
+ $X2=6.48 $Y2=0
r242 63 88 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=6.24 $Y=0 $X2=5.52
+ $Y2=0
r243 61 94 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=8.015 $Y=0 $X2=7.92
+ $Y2=0
r244 61 62 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.015 $Y=0 $X2=8.18
+ $Y2=0
r245 60 98 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=8.345 $Y=0 $X2=8.4
+ $Y2=0
r246 60 62 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.345 $Y=0 $X2=8.18
+ $Y2=0
r247 58 75 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=3.255 $Y=0
+ $X2=3.12 $Y2=0
r248 58 59 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.255 $Y=0 $X2=3.42
+ $Y2=0
r249 57 79 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=3.585 $Y=0 $X2=3.6
+ $Y2=0
r250 57 59 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.585 $Y=0 $X2=3.42
+ $Y2=0
r251 53 129 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=11.34 $Y=0.085
+ $X2=11.34 $Y2=0
r252 53 55 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=11.34 $Y=0.085
+ $X2=11.34 $Y2=0.44
r253 49 126 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.76 $Y=0.085
+ $X2=9.76 $Y2=0
r254 49 51 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=9.76 $Y=0.085
+ $X2=9.76 $Y2=0.44
r255 45 62 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.18 $Y=0.085
+ $X2=8.18 $Y2=0
r256 45 47 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=8.18 $Y=0.085
+ $X2=8.18 $Y2=0.44
r257 41 123 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.6 $Y=0.085
+ $X2=6.6 $Y2=0
r258 41 43 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=6.6 $Y=0.085
+ $X2=6.6 $Y2=0.44
r259 37 120 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.02 $Y=0.085
+ $X2=5.02 $Y2=0
r260 37 39 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=5.02 $Y=0.085
+ $X2=5.02 $Y2=0.44
r261 33 59 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.42 $Y=0.085
+ $X2=3.42 $Y2=0
r262 33 35 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=3.42 $Y=0.085
+ $X2=3.42 $Y2=0.44
r263 29 117 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.84 $Y=0.085
+ $X2=1.84 $Y2=0
r264 29 31 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=1.84 $Y=0.085
+ $X2=1.84 $Y2=0.44
r265 25 114 3.08204 $w=3e-07 $l=1.12161e-07 $layer=LI1_cond $X=0.275 $Y=0.085
+ $X2=0.212 $Y2=0
r266 25 27 13.6372 $w=2.98e-07 $l=3.55e-07 $layer=LI1_cond $X=0.275 $Y=0.085
+ $X2=0.275 $Y2=0.44
r267 8 55 182 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_NDIFF $count=1 $X=11.2
+ $Y=0.235 $X2=11.34 $Y2=0.44
r268 7 51 182 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_NDIFF $count=1 $X=9.62
+ $Y=0.235 $X2=9.76 $Y2=0.44
r269 6 47 182 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_NDIFF $count=1 $X=8.04
+ $Y=0.235 $X2=8.18 $Y2=0.44
r270 5 43 182 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_NDIFF $count=1 $X=6.46
+ $Y=0.235 $X2=6.6 $Y2=0.44
r271 4 39 182 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_NDIFF $count=1 $X=4.88
+ $Y=0.235 $X2=5.02 $Y2=0.44
r272 3 35 182 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_NDIFF $count=1 $X=3.28
+ $Y=0.235 $X2=3.42 $Y2=0.44
r273 2 31 182 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_NDIFF $count=1 $X=1.7
+ $Y=0.235 $X2=1.84 $Y2=0.44
r274 1 27 182 $w=1.7e-07 $l=2.60096e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.44
.ends

