* File: sky130_fd_sc_lp__o311ai_1.pxi.spice
* Created: Fri Aug 28 11:14:26 2020
* 
x_PM_SKY130_FD_SC_LP__O311AI_1%A1 N_A1_M1000_g N_A1_M1009_g A1 A1 N_A1_c_57_n
+ PM_SKY130_FD_SC_LP__O311AI_1%A1
x_PM_SKY130_FD_SC_LP__O311AI_1%A2 N_A2_M1007_g N_A2_M1001_g A2 A2 A2 A2
+ N_A2_c_81_n N_A2_c_82_n PM_SKY130_FD_SC_LP__O311AI_1%A2
x_PM_SKY130_FD_SC_LP__O311AI_1%A3 N_A3_M1005_g N_A3_M1008_g A3 N_A3_c_116_n
+ N_A3_c_117_n PM_SKY130_FD_SC_LP__O311AI_1%A3
x_PM_SKY130_FD_SC_LP__O311AI_1%B1 N_B1_M1006_g N_B1_M1002_g B1 N_B1_c_148_n
+ N_B1_c_149_n PM_SKY130_FD_SC_LP__O311AI_1%B1
x_PM_SKY130_FD_SC_LP__O311AI_1%C1 N_C1_M1004_g N_C1_M1003_g C1 C1 N_C1_c_184_n
+ PM_SKY130_FD_SC_LP__O311AI_1%C1
x_PM_SKY130_FD_SC_LP__O311AI_1%VPWR N_VPWR_M1009_s N_VPWR_M1006_d N_VPWR_c_205_n
+ N_VPWR_c_206_n N_VPWR_c_207_n N_VPWR_c_208_n VPWR N_VPWR_c_209_n
+ N_VPWR_c_210_n N_VPWR_c_204_n N_VPWR_c_212_n PM_SKY130_FD_SC_LP__O311AI_1%VPWR
x_PM_SKY130_FD_SC_LP__O311AI_1%Y N_Y_M1004_d N_Y_M1005_d N_Y_M1003_d N_Y_c_253_n
+ N_Y_c_275_n N_Y_c_248_n N_Y_c_249_n Y Y Y N_Y_c_261_n
+ PM_SKY130_FD_SC_LP__O311AI_1%Y
x_PM_SKY130_FD_SC_LP__O311AI_1%VGND N_VGND_M1000_s N_VGND_M1007_d N_VGND_c_289_n
+ N_VGND_c_290_n N_VGND_c_291_n N_VGND_c_292_n N_VGND_c_293_n N_VGND_c_294_n
+ VGND N_VGND_c_295_n N_VGND_c_296_n PM_SKY130_FD_SC_LP__O311AI_1%VGND
x_PM_SKY130_FD_SC_LP__O311AI_1%A_173_47# N_A_173_47#_M1000_d N_A_173_47#_M1008_d
+ N_A_173_47#_c_327_n N_A_173_47#_c_325_n N_A_173_47#_c_326_n
+ N_A_173_47#_c_349_n PM_SKY130_FD_SC_LP__O311AI_1%A_173_47#
cc_1 VNB N_A1_M1000_g 0.0343536f $X=-0.19 $Y=-0.245 $X2=0.79 $Y2=0.655
cc_2 VNB A1 0.0294598f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_3 VNB N_A1_c_57_n 0.0305838f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.51
cc_4 VNB N_A2_M1007_g 0.0253396f $X=-0.19 $Y=-0.245 $X2=0.79 $Y2=0.655
cc_5 VNB N_A2_c_81_n 0.0240348f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.547
cc_6 VNB N_A2_c_82_n 0.0034924f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_A3_M1008_g 0.0293187f $X=-0.19 $Y=-0.245 $X2=0.79 $Y2=2.465
cc_8 VNB N_A3_c_116_n 0.0239053f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A3_c_117_n 0.00359211f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.51
cc_10 VNB N_B1_M1002_g 0.0280858f $X=-0.19 $Y=-0.245 $X2=0.79 $Y2=2.465
cc_11 VNB N_B1_c_148_n 0.0029417f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.51
cc_12 VNB N_B1_c_149_n 0.0294742f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.345
cc_13 VNB N_C1_M1004_g 0.023581f $X=-0.19 $Y=-0.245 $X2=0.79 $Y2=0.655
cc_14 VNB N_C1_M1003_g 0.00606684f $X=-0.19 $Y=-0.245 $X2=0.79 $Y2=2.465
cc_15 VNB C1 0.0215381f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_16 VNB N_C1_c_184_n 0.0496322f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.345
cc_17 VNB N_VPWR_c_204_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_Y_c_248_n 0.0105881f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.675
cc_19 VNB N_Y_c_249_n 0.0335135f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.547
cc_20 VNB N_VGND_c_289_n 0.0393518f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_21 VNB N_VGND_c_290_n 0.00505246f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.51
cc_22 VNB N_VGND_c_291_n 0.0151903f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.345
cc_23 VNB N_VGND_c_292_n 0.00500104f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.675
cc_24 VNB N_VGND_c_293_n 0.0175532f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_294_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_295_n 0.0449868f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_296_n 0.202338f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_173_47#_c_325_n 0.0156288f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_173_47#_c_326_n 0.00757151f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VPB N_A1_M1009_g 0.0242814f $X=-0.19 $Y=1.655 $X2=0.79 $Y2=2.465
cc_31 VPB A1 0.0200543f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_32 VPB N_A1_c_57_n 0.00674969f $X=-0.19 $Y=1.655 $X2=0.7 $Y2=1.51
cc_33 VPB N_A2_M1001_g 0.0179593f $X=-0.19 $Y=1.655 $X2=0.79 $Y2=2.465
cc_34 VPB N_A2_c_81_n 0.00752527f $X=-0.19 $Y=1.655 $X2=0.24 $Y2=1.547
cc_35 VPB N_A2_c_82_n 0.00275316f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_36 VPB N_A3_M1005_g 0.019705f $X=-0.19 $Y=1.655 $X2=0.79 $Y2=0.655
cc_37 VPB N_A3_c_116_n 0.00615968f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_38 VPB N_A3_c_117_n 0.00661962f $X=-0.19 $Y=1.655 $X2=0.7 $Y2=1.51
cc_39 VPB N_B1_M1006_g 0.0211287f $X=-0.19 $Y=1.655 $X2=0.79 $Y2=0.655
cc_40 VPB N_B1_c_148_n 0.0035173f $X=-0.19 $Y=1.655 $X2=0.7 $Y2=1.51
cc_41 VPB N_B1_c_149_n 0.00901244f $X=-0.19 $Y=1.655 $X2=0.7 $Y2=1.345
cc_42 VPB N_C1_M1003_g 0.0268802f $X=-0.19 $Y=1.655 $X2=0.79 $Y2=2.465
cc_43 VPB C1 0.00870122f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_44 VPB N_VPWR_c_205_n 0.0484537f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_45 VPB N_VPWR_c_206_n 0.00564356f $X=-0.19 $Y=1.655 $X2=0.7 $Y2=1.51
cc_46 VPB N_VPWR_c_207_n 0.0454687f $X=-0.19 $Y=1.655 $X2=0.24 $Y2=1.547
cc_47 VPB N_VPWR_c_208_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_48 VPB N_VPWR_c_209_n 0.0151903f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=1.547
cc_49 VPB N_VPWR_c_210_n 0.0192817f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_50 VPB N_VPWR_c_204_n 0.0570979f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_51 VPB N_VPWR_c_212_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_52 VPB N_Y_c_248_n 0.00334943f $X=-0.19 $Y=1.655 $X2=0.7 $Y2=1.675
cc_53 VPB Y 0.008504f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_54 VPB Y 0.0393706f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_55 N_A1_M1000_g N_A2_M1007_g 0.0240219f $X=0.79 $Y=0.655 $X2=0 $Y2=0
cc_56 N_A1_M1009_g N_A2_M1001_g 0.0618479f $X=0.79 $Y=2.465 $X2=0 $Y2=0
cc_57 A1 N_A2_c_81_n 3.69592e-19 $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_58 N_A1_c_57_n N_A2_c_81_n 0.0206141f $X=0.7 $Y=1.51 $X2=0 $Y2=0
cc_59 A1 N_A2_c_82_n 0.0337366f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_60 N_A1_c_57_n N_A2_c_82_n 0.0144965f $X=0.7 $Y=1.51 $X2=0 $Y2=0
cc_61 N_A1_M1009_g N_VPWR_c_205_n 0.0252947f $X=0.79 $Y=2.465 $X2=0 $Y2=0
cc_62 A1 N_VPWR_c_205_n 0.0261668f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_63 N_A1_c_57_n N_VPWR_c_205_n 0.00102542f $X=0.7 $Y=1.51 $X2=0 $Y2=0
cc_64 N_A1_M1009_g N_VPWR_c_207_n 0.00486043f $X=0.79 $Y=2.465 $X2=0 $Y2=0
cc_65 N_A1_M1009_g N_VPWR_c_204_n 0.00840826f $X=0.79 $Y=2.465 $X2=0 $Y2=0
cc_66 N_A1_M1000_g N_VGND_c_289_n 0.00678015f $X=0.79 $Y=0.655 $X2=0 $Y2=0
cc_67 A1 N_VGND_c_289_n 0.0170907f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_68 N_A1_c_57_n N_VGND_c_289_n 0.00298821f $X=0.7 $Y=1.51 $X2=0 $Y2=0
cc_69 N_A1_M1000_g N_VGND_c_293_n 0.00549284f $X=0.79 $Y=0.655 $X2=0 $Y2=0
cc_70 N_A1_M1000_g N_VGND_c_296_n 0.010916f $X=0.79 $Y=0.655 $X2=0 $Y2=0
cc_71 N_A1_M1000_g N_A_173_47#_c_327_n 0.00918705f $X=0.79 $Y=0.655 $X2=0 $Y2=0
cc_72 N_A1_M1000_g N_A_173_47#_c_326_n 0.00644255f $X=0.79 $Y=0.655 $X2=0 $Y2=0
cc_73 A1 N_A_173_47#_c_326_n 0.0016205f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_74 N_A2_M1001_g N_A3_M1005_g 0.0580927f $X=1.23 $Y=2.465 $X2=0 $Y2=0
cc_75 N_A2_c_82_n N_A3_M1005_g 0.00507952f $X=1.24 $Y=1.51 $X2=0 $Y2=0
cc_76 N_A2_M1007_g N_A3_M1008_g 0.019102f $X=1.22 $Y=0.655 $X2=0 $Y2=0
cc_77 N_A2_c_81_n N_A3_c_116_n 0.0204911f $X=1.24 $Y=1.51 $X2=0 $Y2=0
cc_78 N_A2_c_82_n N_A3_c_116_n 3.182e-19 $X=1.24 $Y=1.51 $X2=0 $Y2=0
cc_79 N_A2_M1001_g N_A3_c_117_n 3.2043e-19 $X=1.23 $Y=2.465 $X2=0 $Y2=0
cc_80 N_A2_c_81_n N_A3_c_117_n 0.00206266f $X=1.24 $Y=1.51 $X2=0 $Y2=0
cc_81 N_A2_c_82_n N_A3_c_117_n 0.0344815f $X=1.24 $Y=1.51 $X2=0 $Y2=0
cc_82 N_A2_M1001_g N_VPWR_c_205_n 0.0025368f $X=1.23 $Y=2.465 $X2=0 $Y2=0
cc_83 N_A2_c_82_n N_VPWR_c_205_n 0.0545787f $X=1.24 $Y=1.51 $X2=0 $Y2=0
cc_84 N_A2_M1001_g N_VPWR_c_207_n 0.00376756f $X=1.23 $Y=2.465 $X2=0 $Y2=0
cc_85 N_A2_c_82_n N_VPWR_c_207_n 0.0115833f $X=1.24 $Y=1.51 $X2=0 $Y2=0
cc_86 N_A2_M1001_g N_VPWR_c_204_n 0.00563467f $X=1.23 $Y=2.465 $X2=0 $Y2=0
cc_87 N_A2_c_82_n N_VPWR_c_204_n 0.011206f $X=1.24 $Y=1.51 $X2=0 $Y2=0
cc_88 N_A2_c_82_n A_173_367# 0.0130813f $X=1.24 $Y=1.51 $X2=-0.19 $Y2=-0.245
cc_89 N_A2_M1007_g N_VGND_c_290_n 0.00182632f $X=1.22 $Y=0.655 $X2=0 $Y2=0
cc_90 N_A2_M1007_g N_VGND_c_293_n 0.00585385f $X=1.22 $Y=0.655 $X2=0 $Y2=0
cc_91 N_A2_M1007_g N_VGND_c_296_n 0.0107676f $X=1.22 $Y=0.655 $X2=0 $Y2=0
cc_92 N_A2_M1007_g N_A_173_47#_c_325_n 0.0145349f $X=1.22 $Y=0.655 $X2=0 $Y2=0
cc_93 N_A2_c_81_n N_A_173_47#_c_325_n 0.00236392f $X=1.24 $Y=1.51 $X2=0 $Y2=0
cc_94 N_A2_c_82_n N_A_173_47#_c_325_n 0.0165031f $X=1.24 $Y=1.51 $X2=0 $Y2=0
cc_95 N_A2_c_81_n N_A_173_47#_c_326_n 5.14458e-19 $X=1.24 $Y=1.51 $X2=0 $Y2=0
cc_96 N_A2_c_82_n N_A_173_47#_c_326_n 0.00991774f $X=1.24 $Y=1.51 $X2=0 $Y2=0
cc_97 N_A3_M1005_g N_B1_M1006_g 0.012629f $X=1.69 $Y=2.465 $X2=0 $Y2=0
cc_98 N_A3_c_117_n N_B1_M1006_g 2.87075e-19 $X=1.78 $Y=1.51 $X2=0 $Y2=0
cc_99 N_A3_M1008_g N_B1_M1002_g 0.00873284f $X=1.73 $Y=0.655 $X2=0 $Y2=0
cc_100 N_A3_M1005_g N_B1_c_148_n 3.05546e-19 $X=1.69 $Y=2.465 $X2=0 $Y2=0
cc_101 N_A3_c_116_n N_B1_c_148_n 0.00220692f $X=1.78 $Y=1.51 $X2=0 $Y2=0
cc_102 N_A3_c_117_n N_B1_c_148_n 0.0349137f $X=1.78 $Y=1.51 $X2=0 $Y2=0
cc_103 N_A3_c_116_n N_B1_c_149_n 0.0204626f $X=1.78 $Y=1.51 $X2=0 $Y2=0
cc_104 N_A3_c_117_n N_B1_c_149_n 2.85635e-19 $X=1.78 $Y=1.51 $X2=0 $Y2=0
cc_105 N_A3_M1005_g N_VPWR_c_207_n 0.00585385f $X=1.69 $Y=2.465 $X2=0 $Y2=0
cc_106 N_A3_M1005_g N_VPWR_c_204_n 0.0112442f $X=1.69 $Y=2.465 $X2=0 $Y2=0
cc_107 N_A3_c_116_n N_Y_c_253_n 0.00357197f $X=1.78 $Y=1.51 $X2=0 $Y2=0
cc_108 N_A3_c_117_n N_Y_c_253_n 0.00480792f $X=1.78 $Y=1.51 $X2=0 $Y2=0
cc_109 N_A3_M1008_g N_VGND_c_290_n 0.00327036f $X=1.73 $Y=0.655 $X2=0 $Y2=0
cc_110 N_A3_M1008_g N_VGND_c_295_n 0.00585385f $X=1.73 $Y=0.655 $X2=0 $Y2=0
cc_111 N_A3_M1008_g N_VGND_c_296_n 0.0113834f $X=1.73 $Y=0.655 $X2=0 $Y2=0
cc_112 N_A3_M1008_g N_A_173_47#_c_325_n 0.0152811f $X=1.73 $Y=0.655 $X2=0 $Y2=0
cc_113 N_A3_c_116_n N_A_173_47#_c_325_n 0.00433842f $X=1.78 $Y=1.51 $X2=0 $Y2=0
cc_114 N_A3_c_117_n N_A_173_47#_c_325_n 0.0263322f $X=1.78 $Y=1.51 $X2=0 $Y2=0
cc_115 N_B1_M1002_g N_C1_M1004_g 0.0459181f $X=2.5 $Y=0.655 $X2=0 $Y2=0
cc_116 N_B1_M1006_g N_C1_M1003_g 0.0278533f $X=2.23 $Y=2.465 $X2=0 $Y2=0
cc_117 N_B1_c_149_n N_C1_c_184_n 0.0459181f $X=2.5 $Y=1.51 $X2=0 $Y2=0
cc_118 N_B1_M1006_g N_VPWR_c_206_n 0.0120173f $X=2.23 $Y=2.465 $X2=0 $Y2=0
cc_119 N_B1_M1006_g N_VPWR_c_207_n 0.00585385f $X=2.23 $Y=2.465 $X2=0 $Y2=0
cc_120 N_B1_M1006_g N_VPWR_c_204_n 0.0115408f $X=2.23 $Y=2.465 $X2=0 $Y2=0
cc_121 N_B1_c_148_n N_Y_c_253_n 0.00675081f $X=2.32 $Y=1.51 $X2=0 $Y2=0
cc_122 N_B1_M1006_g N_Y_c_248_n 0.00358764f $X=2.23 $Y=2.465 $X2=0 $Y2=0
cc_123 N_B1_M1002_g N_Y_c_248_n 0.0105406f $X=2.5 $Y=0.655 $X2=0 $Y2=0
cc_124 N_B1_c_148_n N_Y_c_248_n 0.0337002f $X=2.32 $Y=1.51 $X2=0 $Y2=0
cc_125 N_B1_M1006_g Y 2.34189e-19 $X=2.23 $Y=2.465 $X2=0 $Y2=0
cc_126 N_B1_M1006_g Y 9.08036e-19 $X=2.23 $Y=2.465 $X2=0 $Y2=0
cc_127 N_B1_M1006_g N_Y_c_261_n 0.0138701f $X=2.23 $Y=2.465 $X2=0 $Y2=0
cc_128 N_B1_c_148_n N_Y_c_261_n 0.0181259f $X=2.32 $Y=1.51 $X2=0 $Y2=0
cc_129 N_B1_c_149_n N_Y_c_261_n 0.00665691f $X=2.5 $Y=1.51 $X2=0 $Y2=0
cc_130 N_B1_M1002_g N_VGND_c_295_n 0.00585385f $X=2.5 $Y=0.655 $X2=0 $Y2=0
cc_131 N_B1_M1002_g N_VGND_c_296_n 0.0113463f $X=2.5 $Y=0.655 $X2=0 $Y2=0
cc_132 N_B1_M1002_g N_A_173_47#_c_325_n 0.00128014f $X=2.5 $Y=0.655 $X2=0 $Y2=0
cc_133 N_B1_c_148_n N_A_173_47#_c_325_n 0.0323195f $X=2.32 $Y=1.51 $X2=0 $Y2=0
cc_134 N_B1_c_149_n N_A_173_47#_c_325_n 0.00641554f $X=2.5 $Y=1.51 $X2=0 $Y2=0
cc_135 N_C1_M1003_g N_VPWR_c_206_n 0.0113301f $X=2.86 $Y=2.465 $X2=0 $Y2=0
cc_136 N_C1_M1003_g N_VPWR_c_210_n 0.0054895f $X=2.86 $Y=2.465 $X2=0 $Y2=0
cc_137 N_C1_M1003_g N_VPWR_c_204_n 0.0113763f $X=2.86 $Y=2.465 $X2=0 $Y2=0
cc_138 N_C1_M1004_g N_Y_c_248_n 0.0103187f $X=2.86 $Y=0.655 $X2=0 $Y2=0
cc_139 C1 N_Y_c_248_n 0.0434794f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_140 N_C1_M1004_g N_Y_c_249_n 0.0287429f $X=2.86 $Y=0.655 $X2=0 $Y2=0
cc_141 C1 N_Y_c_249_n 0.023654f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_142 N_C1_c_184_n N_Y_c_249_n 0.00222846f $X=3.09 $Y=1.375 $X2=0 $Y2=0
cc_143 N_C1_M1003_g Y 0.0178276f $X=2.86 $Y=2.465 $X2=0 $Y2=0
cc_144 C1 Y 0.0257895f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_145 N_C1_c_184_n Y 0.00125139f $X=3.09 $Y=1.375 $X2=0 $Y2=0
cc_146 N_C1_M1003_g Y 0.0146212f $X=2.86 $Y=2.465 $X2=0 $Y2=0
cc_147 N_C1_M1004_g N_VGND_c_295_n 0.00357668f $X=2.86 $Y=0.655 $X2=0 $Y2=0
cc_148 N_C1_M1004_g N_VGND_c_296_n 0.00613857f $X=2.86 $Y=0.655 $X2=0 $Y2=0
cc_149 N_VPWR_c_204_n A_173_367# 0.00814802f $X=3.12 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_150 N_VPWR_c_204_n A_261_367# 0.0115887f $X=3.12 $Y=3.33 $X2=-0.19 $Y2=-0.245
cc_151 N_VPWR_c_204_n N_Y_M1005_d 0.00521751f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_152 N_VPWR_c_204_n N_Y_M1003_d 0.00215158f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_153 N_VPWR_c_207_n N_Y_c_275_n 0.0212513f $X=2.38 $Y=3.33 $X2=0 $Y2=0
cc_154 N_VPWR_c_204_n N_Y_c_275_n 0.0127519f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_155 N_VPWR_M1006_d N_Y_c_248_n 0.00194138f $X=2.305 $Y=1.835 $X2=0 $Y2=0
cc_156 N_VPWR_M1006_d Y 0.00302499f $X=2.305 $Y=1.835 $X2=0 $Y2=0
cc_157 N_VPWR_c_206_n Y 0.0541709f $X=2.545 $Y=2.395 $X2=0 $Y2=0
cc_158 N_VPWR_c_210_n Y 0.0235557f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_159 N_VPWR_c_204_n Y 0.0139296f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_160 N_VPWR_M1006_d N_Y_c_261_n 0.00610506f $X=2.305 $Y=1.835 $X2=0 $Y2=0
cc_161 N_VPWR_c_206_n N_Y_c_261_n 0.0266544f $X=2.545 $Y=2.395 $X2=0 $Y2=0
cc_162 N_Y_c_249_n N_VGND_c_295_n 0.0403958f $X=3.075 $Y=0.38 $X2=0 $Y2=0
cc_163 N_Y_M1004_d N_VGND_c_296_n 0.00215158f $X=2.935 $Y=0.235 $X2=0 $Y2=0
cc_164 N_Y_c_249_n N_VGND_c_296_n 0.0250164f $X=3.075 $Y=0.38 $X2=0 $Y2=0
cc_165 N_Y_c_248_n N_A_173_47#_c_325_n 0.00841925f $X=2.67 $Y=1.94 $X2=0 $Y2=0
cc_166 N_Y_c_249_n A_515_47# 9.38685e-19 $X=3.075 $Y=0.38 $X2=-0.19 $Y2=-0.245
cc_167 N_VGND_c_296_n N_A_173_47#_M1000_d 0.00241208f $X=3.12 $Y=0 $X2=-0.19
+ $Y2=-0.245
cc_168 N_VGND_c_296_n N_A_173_47#_M1008_d 0.00593242f $X=3.12 $Y=0 $X2=0 $Y2=0
cc_169 N_VGND_c_293_n N_A_173_47#_c_327_n 0.0160895f $X=1.31 $Y=0 $X2=0 $Y2=0
cc_170 N_VGND_c_296_n N_A_173_47#_c_327_n 0.0113472f $X=3.12 $Y=0 $X2=0 $Y2=0
cc_171 N_VGND_M1007_d N_A_173_47#_c_325_n 0.00261503f $X=1.295 $Y=0.235 $X2=0
+ $Y2=0
cc_172 N_VGND_c_290_n N_A_173_47#_c_325_n 0.0200142f $X=1.475 $Y=0.36 $X2=0
+ $Y2=0
cc_173 N_VGND_c_289_n N_A_173_47#_c_326_n 0.00455684f $X=0.575 $Y=0.38 $X2=0
+ $Y2=0
cc_174 N_VGND_c_295_n N_A_173_47#_c_349_n 0.0363434f $X=3.12 $Y=0 $X2=0 $Y2=0
cc_175 N_VGND_c_296_n N_A_173_47#_c_349_n 0.022945f $X=3.12 $Y=0 $X2=0 $Y2=0
cc_176 N_VGND_c_296_n A_515_47# 0.00168071f $X=3.12 $Y=0 $X2=-0.19 $Y2=-0.245
