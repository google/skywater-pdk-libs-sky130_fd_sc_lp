# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__nand4_2
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__nand4_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.800000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.505000 1.425000 4.715000 1.750000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.005000 1.425000 3.335000 1.750000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.585000 1.165000 2.330000 1.435000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.555000 1.345000 0.845000 1.640000 ;
        RECT 0.555000 1.640000 0.805000 1.670000 ;
        RECT 0.625000 1.670000 0.805000 2.120000 ;
    END
  END D
  PIN Y
    ANTENNADIFFAREA  1.646400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.975000 1.755000 2.835000 1.920000 ;
        RECT 0.975000 1.920000 4.075000 1.925000 ;
        RECT 0.975000 1.925000 1.165000 3.075000 ;
        RECT 1.835000 1.925000 4.075000 2.090000 ;
        RECT 1.835000 2.090000 2.015000 3.075000 ;
        RECT 2.015000 1.605000 2.835000 1.755000 ;
        RECT 2.500000 1.075000 4.215000 1.245000 ;
        RECT 2.500000 1.245000 2.835000 1.605000 ;
        RECT 2.740000 2.090000 3.035000 3.075000 ;
        RECT 3.815000 2.090000 4.075000 3.075000 ;
        RECT 3.885000 0.595000 4.215000 1.075000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.800000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.800000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.800000 0.085000 ;
      RECT 0.000000  3.245000 4.800000 3.415000 ;
      RECT 0.135000  1.815000 0.455000 2.295000 ;
      RECT 0.135000  2.295000 0.805000 3.245000 ;
      RECT 0.305000  0.255000 0.565000 0.985000 ;
      RECT 0.305000  0.985000 1.415000 1.155000 ;
      RECT 0.735000  0.085000 1.065000 0.805000 ;
      RECT 1.235000  0.255000 2.385000 0.545000 ;
      RECT 1.235000  0.545000 1.415000 0.985000 ;
      RECT 1.335000  2.095000 1.665000 3.245000 ;
      RECT 1.625000  0.715000 3.355000 0.905000 ;
      RECT 1.625000  0.905000 1.955000 0.995000 ;
      RECT 2.240000  2.260000 2.570000 3.245000 ;
      RECT 2.595000  0.255000 4.645000 0.425000 ;
      RECT 2.595000  0.425000 3.715000 0.545000 ;
      RECT 3.260000  2.260000 3.590000 3.245000 ;
      RECT 3.525000  0.545000 3.715000 0.905000 ;
      RECT 4.245000  1.920000 4.575000 3.245000 ;
      RECT 4.385000  0.425000 4.645000 1.195000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
  END
END sky130_fd_sc_lp__nand4_2
