* File: sky130_fd_sc_lp__buflp_4.pex.spice
* Created: Fri Aug 28 10:12:39 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__BUFLP_4%A_84_21# 1 2 9 13 17 21 25 29 33 37 41 45 49
+ 53 57 61 65 69 71 77 78 79 82 86 93 108
c194 69 0 4.8492e-20 $X=3.785 $Y=2.465
c195 45 0 1.08995e-19 $X=2.285 $Y=2.465
r196 105 106 38.4695 $w=3.3e-07 $l=2.2e-07 $layer=POLY_cond $X=3.285 $Y=1.48
+ $X2=3.505 $Y2=1.48
r197 104 105 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=3.075 $Y=1.48
+ $X2=3.285 $Y2=1.48
r198 103 104 50.7098 $w=3.3e-07 $l=2.9e-07 $layer=POLY_cond $X=2.785 $Y=1.48
+ $X2=3.075 $Y2=1.48
r199 102 103 24.4806 $w=3.3e-07 $l=1.4e-07 $layer=POLY_cond $X=2.645 $Y=1.48
+ $X2=2.785 $Y2=1.48
r200 101 102 62.9501 $w=3.3e-07 $l=3.6e-07 $layer=POLY_cond $X=2.285 $Y=1.48
+ $X2=2.645 $Y2=1.48
r201 100 101 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=2.215 $Y=1.48
+ $X2=2.285 $Y2=1.48
r202 99 100 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=1.785 $Y=1.48
+ $X2=2.215 $Y2=1.48
r203 98 99 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=1.355 $Y=1.48
+ $X2=1.785 $Y2=1.48
r204 97 98 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=0.925 $Y=1.48
+ $X2=1.355 $Y2=1.48
r205 92 108 27.1035 $w=3.3e-07 $l=1.55e-07 $layer=POLY_cond $X=3.63 $Y=1.48
+ $X2=3.785 $Y2=1.48
r206 92 106 21.8577 $w=3.3e-07 $l=1.25e-07 $layer=POLY_cond $X=3.63 $Y=1.48
+ $X2=3.505 $Y2=1.48
r207 91 92 32.2844 $w=1.7e-07 $l=7.65e-07 $layer=licon1_POLY $count=4 $X=3.63
+ $Y=1.48 $X2=3.63 $Y2=1.48
r208 86 88 32.4779 $w=3.28e-07 $l=9.3e-07 $layer=LI1_cond $X=4.96 $Y=1.98
+ $X2=4.96 $Y2=2.91
r209 84 93 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.96 $Y=1.01
+ $X2=4.96 $Y2=0.925
r210 84 86 33.8748 $w=3.28e-07 $l=9.7e-07 $layer=LI1_cond $X=4.96 $Y=1.01
+ $X2=4.96 $Y2=1.98
r211 80 93 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.96 $Y=0.84
+ $X2=4.96 $Y2=0.925
r212 80 82 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=4.96 $Y=0.84
+ $X2=4.96 $Y2=0.42
r213 78 93 3.80956 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.795 $Y=0.925
+ $X2=4.96 $Y2=0.925
r214 78 79 65.2406 $w=1.68e-07 $l=1e-06 $layer=LI1_cond $X=4.795 $Y=0.925
+ $X2=3.795 $Y2=0.925
r215 77 91 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.71 $Y=1.315
+ $X2=3.71 $Y2=1.48
r216 76 79 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.71 $Y=1.01
+ $X2=3.795 $Y2=0.925
r217 76 77 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3.71 $Y=1.01
+ $X2=3.71 $Y2=1.315
r218 74 97 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=0.91 $Y=1.48
+ $X2=0.925 $Y2=1.48
r219 74 94 72.5674 $w=3.3e-07 $l=4.15e-07 $layer=POLY_cond $X=0.91 $Y=1.48
+ $X2=0.495 $Y2=1.48
r220 73 74 32.2844 $w=1.7e-07 $l=7.65e-07 $layer=licon1_POLY $count=4 $X=0.91
+ $Y=1.48 $X2=0.91 $Y2=1.48
r221 71 91 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.625 $Y=1.48
+ $X2=3.71 $Y2=1.48
r222 71 73 94.8146 $w=3.28e-07 $l=2.715e-06 $layer=LI1_cond $X=3.625 $Y=1.48
+ $X2=0.91 $Y2=1.48
r223 67 108 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.785 $Y=1.645
+ $X2=3.785 $Y2=1.48
r224 67 69 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=3.785 $Y=1.645
+ $X2=3.785 $Y2=2.465
r225 63 106 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.505 $Y=1.315
+ $X2=3.505 $Y2=1.48
r226 63 65 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.505 $Y=1.315
+ $X2=3.505 $Y2=0.655
r227 59 105 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.285 $Y=1.645
+ $X2=3.285 $Y2=1.48
r228 59 61 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=3.285 $Y=1.645
+ $X2=3.285 $Y2=2.465
r229 55 104 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.075 $Y=1.315
+ $X2=3.075 $Y2=1.48
r230 55 57 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.075 $Y=1.315
+ $X2=3.075 $Y2=0.655
r231 51 103 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.785 $Y=1.645
+ $X2=2.785 $Y2=1.48
r232 51 53 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=2.785 $Y=1.645
+ $X2=2.785 $Y2=2.465
r233 47 102 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.645 $Y=1.315
+ $X2=2.645 $Y2=1.48
r234 47 49 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.645 $Y=1.315
+ $X2=2.645 $Y2=0.655
r235 43 101 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.285 $Y=1.645
+ $X2=2.285 $Y2=1.48
r236 43 45 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=2.285 $Y=1.645
+ $X2=2.285 $Y2=2.465
r237 39 100 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.215 $Y=1.315
+ $X2=2.215 $Y2=1.48
r238 39 41 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.215 $Y=1.315
+ $X2=2.215 $Y2=0.655
r239 35 99 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.785 $Y=1.645
+ $X2=1.785 $Y2=1.48
r240 35 37 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=1.785 $Y=1.645
+ $X2=1.785 $Y2=2.465
r241 31 99 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.785 $Y=1.315
+ $X2=1.785 $Y2=1.48
r242 31 33 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.785 $Y=1.315
+ $X2=1.785 $Y2=0.655
r243 27 98 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.355 $Y=1.645
+ $X2=1.355 $Y2=1.48
r244 27 29 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=1.355 $Y=1.645
+ $X2=1.355 $Y2=2.465
r245 23 98 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.355 $Y=1.315
+ $X2=1.355 $Y2=1.48
r246 23 25 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.355 $Y=1.315
+ $X2=1.355 $Y2=0.655
r247 19 97 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.925 $Y=1.645
+ $X2=0.925 $Y2=1.48
r248 19 21 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=0.925 $Y=1.645
+ $X2=0.925 $Y2=2.465
r249 15 97 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.925 $Y=1.315
+ $X2=0.925 $Y2=1.48
r250 15 17 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.925 $Y=1.315
+ $X2=0.925 $Y2=0.655
r251 11 94 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=1.645
+ $X2=0.495 $Y2=1.48
r252 11 13 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=0.495 $Y=1.645
+ $X2=0.495 $Y2=2.465
r253 7 94 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=1.315
+ $X2=0.495 $Y2=1.48
r254 7 9 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.495 $Y=1.315
+ $X2=0.495 $Y2=0.655
r255 2 88 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=4.82
+ $Y=1.835 $X2=4.96 $Y2=2.91
r256 2 86 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=4.82
+ $Y=1.835 $X2=4.96 $Y2=1.98
r257 1 82 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=4.82
+ $Y=0.235 $X2=4.96 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__BUFLP_4%A 3 6 8 10 12 15 17 18 20 21 24
r45 23 25 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.265 $Y=1.35
+ $X2=4.265 $Y2=1.515
r46 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.265
+ $Y=1.35 $X2=4.265 $Y2=1.35
r47 20 23 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=4.265 $Y=1.26
+ $X2=4.265 $Y2=1.35
r48 20 21 30.474 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=4.265 $Y=1.26
+ $X2=4.265 $Y2=1.185
r49 18 24 6.36424 $w=3.33e-07 $l=1.85e-07 $layer=LI1_cond $X=4.08 $Y=1.347
+ $X2=4.265 $Y2=1.347
r50 13 17 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.745 $Y=1.335
+ $X2=4.745 $Y2=1.26
r51 13 15 579.426 $w=1.5e-07 $l=1.13e-06 $layer=POLY_cond $X=4.745 $Y=1.335
+ $X2=4.745 $Y2=2.465
r52 10 17 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.745 $Y=1.185
+ $X2=4.745 $Y2=1.26
r53 10 12 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=4.745 $Y=1.185
+ $X2=4.745 $Y2=0.655
r54 9 20 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.43 $Y=1.26
+ $X2=4.265 $Y2=1.26
r55 8 17 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.67 $Y=1.26
+ $X2=4.745 $Y2=1.26
r56 8 9 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=4.67 $Y=1.26 $X2=4.43
+ $Y2=1.26
r57 6 25 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=4.355 $Y=2.465
+ $X2=4.355 $Y2=1.515
r58 3 21 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=4.355 $Y=0.655
+ $X2=4.355 $Y2=1.185
.ends

.subckt PM_SKY130_FD_SC_LP__BUFLP_4%VPWR 1 2 3 10 12 16 20 24 26 31 38 39 45 48
c68 1 0 7.44113e-20 $X=0.135 $Y=1.835
r69 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r70 45 46 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r71 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r72 39 49 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=4.08 $Y2=3.33
r73 38 39 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r74 36 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.235 $Y=3.33
+ $X2=4.07 $Y2=3.33
r75 36 38 52.5187 $w=1.68e-07 $l=8.05e-07 $layer=LI1_cond $X=4.235 $Y=3.33
+ $X2=5.04 $Y2=3.33
r76 35 49 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r77 34 35 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r78 32 45 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.225 $Y=3.33
+ $X2=1.14 $Y2=3.33
r79 32 34 154.947 $w=1.68e-07 $l=2.375e-06 $layer=LI1_cond $X=1.225 $Y=3.33
+ $X2=3.6 $Y2=3.33
r80 31 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.905 $Y=3.33
+ $X2=4.07 $Y2=3.33
r81 31 34 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3.905 $Y=3.33
+ $X2=3.6 $Y2=3.33
r82 30 46 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r83 30 43 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r84 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r85 27 42 4.00981 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=0.365 $Y=3.33
+ $X2=0.182 $Y2=3.33
r86 27 29 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=0.365 $Y=3.33
+ $X2=0.72 $Y2=3.33
r87 26 45 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.055 $Y=3.33
+ $X2=1.14 $Y2=3.33
r88 26 29 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.055 $Y=3.33
+ $X2=0.72 $Y2=3.33
r89 24 35 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r90 24 46 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=1.2 $Y2=3.33
r91 20 23 33.8748 $w=3.28e-07 $l=9.7e-07 $layer=LI1_cond $X=4.07 $Y=1.98
+ $X2=4.07 $Y2=2.95
r92 18 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.07 $Y=3.245
+ $X2=4.07 $Y2=3.33
r93 18 23 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=4.07 $Y=3.245
+ $X2=4.07 $Y2=2.95
r94 14 45 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.14 $Y=3.245
+ $X2=1.14 $Y2=3.33
r95 14 16 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=1.14 $Y=3.245
+ $X2=1.14 $Y2=2.805
r96 10 42 3.13335 $w=2.5e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.24 $Y=3.245
+ $X2=0.182 $Y2=3.33
r97 10 12 42.6404 $w=2.48e-07 $l=9.25e-07 $layer=LI1_cond $X=0.24 $Y=3.245
+ $X2=0.24 $Y2=2.32
r98 3 23 400 $w=1.7e-07 $l=1.21547e-06 $layer=licon1_PDIFF $count=1 $X=3.86
+ $Y=1.835 $X2=4.07 $Y2=2.95
r99 3 20 400 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=1 $X=3.86
+ $Y=1.835 $X2=4.07 $Y2=1.98
r100 2 16 600 $w=1.7e-07 $l=1.03764e-06 $layer=licon1_PDIFF $count=1 $X=1
+ $Y=1.835 $X2=1.14 $Y2=2.805
r101 1 12 300 $w=1.7e-07 $l=5.52766e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.835 $X2=0.28 $Y2=2.32
.ends

.subckt PM_SKY130_FD_SC_LP__BUFLP_4%A_114_367# 1 2 3 4 15 17 18 19 20 23 25 27
+ 29 32 35
c58 17 0 1.08995e-19 $X=1.57 $Y=2.325
r59 27 37 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.57 $Y=2.905 $X2=3.57
+ $Y2=2.99
r60 27 29 32.3033 $w=3.28e-07 $l=9.25e-07 $layer=LI1_cond $X=3.57 $Y=2.905
+ $X2=3.57 $Y2=1.98
r61 26 35 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.735 $Y=2.99
+ $X2=2.57 $Y2=2.99
r62 25 37 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.405 $Y=2.99
+ $X2=3.57 $Y2=2.99
r63 25 26 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.405 $Y=2.99
+ $X2=2.735 $Y2=2.99
r64 21 35 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.57 $Y=2.905
+ $X2=2.57 $Y2=2.99
r65 21 23 20.4297 $w=3.28e-07 $l=5.85e-07 $layer=LI1_cond $X=2.57 $Y=2.905
+ $X2=2.57 $Y2=2.32
r66 19 35 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.405 $Y=2.99
+ $X2=2.57 $Y2=2.99
r67 19 20 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.405 $Y=2.99
+ $X2=1.735 $Y2=2.99
r68 18 20 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.57 $Y=2.905
+ $X2=1.735 $Y2=2.99
r69 17 34 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.57 $Y=2.325 $X2=1.57
+ $Y2=2.24
r70 17 18 20.2551 $w=3.28e-07 $l=5.8e-07 $layer=LI1_cond $X=1.57 $Y=2.325
+ $X2=1.57 $Y2=2.905
r71 16 32 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.875 $Y=2.24
+ $X2=0.71 $Y2=2.24
r72 15 34 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.405 $Y=2.24
+ $X2=1.57 $Y2=2.24
r73 15 16 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=1.405 $Y=2.24
+ $X2=0.875 $Y2=2.24
r74 4 37 400 $w=1.7e-07 $l=1.17532e-06 $layer=licon1_PDIFF $count=1 $X=3.36
+ $Y=1.835 $X2=3.57 $Y2=2.91
r75 4 29 400 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=1 $X=3.36
+ $Y=1.835 $X2=3.57 $Y2=1.98
r76 3 23 300 $w=1.7e-07 $l=5.80582e-07 $layer=licon1_PDIFF $count=2 $X=2.36
+ $Y=1.835 $X2=2.57 $Y2=2.32
r77 2 34 300 $w=1.7e-07 $l=5.50568e-07 $layer=licon1_PDIFF $count=2 $X=1.43
+ $Y=1.835 $X2=1.57 $Y2=2.32
r78 1 32 300 $w=1.7e-07 $l=5.50568e-07 $layer=licon1_PDIFF $count=2 $X=0.57
+ $Y=1.835 $X2=0.71 $Y2=2.32
.ends

.subckt PM_SKY130_FD_SC_LP__BUFLP_4%X 1 2 3 4 13 14 15 19 23 25 29 34 36 38 39
+ 40 49
c86 38 0 4.8492e-20 $X=3.07 $Y=1.98
c87 15 0 7.44113e-20 $X=1.905 $Y=1.9
c88 13 0 7.44113e-20 $X=1.835 $Y=1.06
r89 40 53 12.3277 $w=1.91e-07 $l=1.93e-07 $layer=LI1_cond $X=0.24 $Y=1.707
+ $X2=0.24 $Y2=1.9
r90 40 49 2.68272 $w=1.91e-07 $l=4.2e-08 $layer=LI1_cond $X=0.24 $Y=1.707
+ $X2=0.24 $Y2=1.665
r91 40 49 2.15457 $w=2.28e-07 $l=4.3e-08 $layer=LI1_cond $X=0.24 $Y=1.622
+ $X2=0.24 $Y2=1.665
r92 39 40 16.3847 $w=2.28e-07 $l=3.27e-07 $layer=LI1_cond $X=0.24 $Y=1.295
+ $X2=0.24 $Y2=1.622
r93 33 39 7.51593 $w=2.28e-07 $l=1.5e-07 $layer=LI1_cond $X=0.24 $Y=1.145
+ $X2=0.24 $Y2=1.295
r94 27 29 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=2.86 $Y=0.975
+ $X2=2.86 $Y2=0.845
r95 26 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.235 $Y=1.9
+ $X2=2.07 $Y2=1.9
r96 25 38 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.905 $Y=1.9
+ $X2=3.07 $Y2=1.9
r97 25 26 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.905 $Y=1.9
+ $X2=2.235 $Y2=1.9
r98 24 34 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.085 $Y=1.06
+ $X2=1.96 $Y2=1.06
r99 23 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.775 $Y=1.06
+ $X2=2.86 $Y2=0.975
r100 23 24 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.775 $Y=1.06
+ $X2=2.085 $Y2=1.06
r101 17 34 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.96 $Y=0.975
+ $X2=1.96 $Y2=1.06
r102 17 19 5.9927 $w=2.48e-07 $l=1.3e-07 $layer=LI1_cond $X=1.96 $Y=0.975
+ $X2=1.96 $Y2=0.845
r103 16 53 1.41722 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=0.355 $Y=1.9
+ $X2=0.24 $Y2=1.9
r104 15 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.905 $Y=1.9
+ $X2=2.07 $Y2=1.9
r105 15 16 101.123 $w=1.68e-07 $l=1.55e-06 $layer=LI1_cond $X=1.905 $Y=1.9
+ $X2=0.355 $Y2=1.9
r106 14 33 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=0.355 $Y=1.06
+ $X2=0.24 $Y2=1.145
r107 13 34 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.835 $Y=1.06
+ $X2=1.96 $Y2=1.06
r108 13 14 96.5562 $w=1.68e-07 $l=1.48e-06 $layer=LI1_cond $X=1.835 $Y=1.06
+ $X2=0.355 $Y2=1.06
r109 4 38 300 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=2 $X=2.86
+ $Y=1.835 $X2=3.07 $Y2=1.98
r110 3 36 300 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=2 $X=1.86
+ $Y=1.835 $X2=2.07 $Y2=1.98
r111 2 29 182 $w=1.7e-07 $l=6.76387e-07 $layer=licon1_NDIFF $count=1 $X=2.72
+ $Y=0.235 $X2=2.86 $Y2=0.845
r112 1 19 182 $w=1.7e-07 $l=6.76387e-07 $layer=licon1_NDIFF $count=1 $X=1.86
+ $Y=0.235 $X2=2 $Y2=0.845
.ends

.subckt PM_SKY130_FD_SC_LP__BUFLP_4%VGND 1 2 3 10 12 16 20 23 24 25 27 43 44 50
c76 1 0 7.44113e-20 $X=0.135 $Y=0.235
r77 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r78 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r79 43 44 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r80 41 44 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=5.04
+ $Y2=0
r81 40 43 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=4.08 $Y=0 $X2=5.04
+ $Y2=0
r82 40 41 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r83 38 41 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r84 37 38 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r85 35 51 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r86 34 37 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=1.68 $Y=0 $X2=3.6
+ $Y2=0
r87 34 35 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r88 32 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.305 $Y=0 $X2=1.14
+ $Y2=0
r89 32 34 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.305 $Y=0 $X2=1.68
+ $Y2=0
r90 31 51 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r91 31 48 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r92 30 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r93 28 47 4.00981 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=0.365 $Y=0 $X2=0.182
+ $Y2=0
r94 28 30 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=0.365 $Y=0 $X2=0.72
+ $Y2=0
r95 27 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.975 $Y=0 $X2=1.14
+ $Y2=0
r96 27 30 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.975 $Y=0 $X2=0.72
+ $Y2=0
r97 25 38 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r98 25 35 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=1.68
+ $Y2=0
r99 23 37 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=3.625 $Y=0 $X2=3.6
+ $Y2=0
r100 23 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.625 $Y=0 $X2=3.79
+ $Y2=0
r101 22 40 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=3.955 $Y=0
+ $X2=4.08 $Y2=0
r102 22 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.955 $Y=0 $X2=3.79
+ $Y2=0
r103 18 24 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.79 $Y=0.085
+ $X2=3.79 $Y2=0
r104 18 20 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=3.79 $Y=0.085
+ $X2=3.79 $Y2=0.44
r105 14 50 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.14 $Y=0.085
+ $X2=1.14 $Y2=0
r106 14 16 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.14 $Y=0.085
+ $X2=1.14 $Y2=0.38
r107 10 47 3.13335 $w=2.5e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.24 $Y=0.085
+ $X2=0.182 $Y2=0
r108 10 12 19.5915 $w=2.48e-07 $l=4.25e-07 $layer=LI1_cond $X=0.24 $Y=0.085
+ $X2=0.24 $Y2=0.51
r109 3 20 182 $w=1.7e-07 $l=2.95212e-07 $layer=licon1_NDIFF $count=1 $X=3.58
+ $Y=0.235 $X2=3.79 $Y2=0.44
r110 2 16 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=1
+ $Y=0.235 $X2=1.14 $Y2=0.38
r111 1 12 182 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.28 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_LP__BUFLP_4%A_114_47# 1 2 3 4 15 17 18 23 24 27 29 33 35
r56 30 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.595 $Y=0.34
+ $X2=2.43 $Y2=0.34
r57 29 35 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.125 $Y=0.34
+ $X2=3.29 $Y2=0.34
r58 29 30 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=3.125 $Y=0.34
+ $X2=2.595 $Y2=0.34
r59 25 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.43 $Y=0.425
+ $X2=2.43 $Y2=0.34
r60 25 27 3.66686 $w=3.28e-07 $l=1.05e-07 $layer=LI1_cond $X=2.43 $Y=0.425
+ $X2=2.43 $Y2=0.53
r61 23 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.265 $Y=0.34
+ $X2=2.43 $Y2=0.34
r62 23 24 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=2.265 $Y=0.34
+ $X2=1.655 $Y2=0.34
r63 20 22 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=1.57 $Y=0.635
+ $X2=1.57 $Y2=0.53
r64 19 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.57 $Y=0.425
+ $X2=1.655 $Y2=0.34
r65 19 22 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=1.57 $Y=0.425
+ $X2=1.57 $Y2=0.53
r66 17 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.485 $Y=0.72
+ $X2=1.57 $Y2=0.635
r67 17 18 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.485 $Y=0.72
+ $X2=0.795 $Y2=0.72
r68 13 18 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.67 $Y=0.635
+ $X2=0.795 $Y2=0.72
r69 13 15 4.84026 $w=2.48e-07 $l=1.05e-07 $layer=LI1_cond $X=0.67 $Y=0.635
+ $X2=0.67 $Y2=0.53
r70 4 35 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=3.15
+ $Y=0.235 $X2=3.29 $Y2=0.42
r71 3 27 182 $w=1.7e-07 $l=3.58225e-07 $layer=licon1_NDIFF $count=1 $X=2.29
+ $Y=0.235 $X2=2.43 $Y2=0.53
r72 2 22 182 $w=1.7e-07 $l=3.58225e-07 $layer=licon1_NDIFF $count=1 $X=1.43
+ $Y=0.235 $X2=1.57 $Y2=0.53
r73 1 15 182 $w=1.7e-07 $l=3.58225e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.235 $X2=0.71 $Y2=0.53
.ends

