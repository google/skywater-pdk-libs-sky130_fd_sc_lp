* NGSPICE file created from sky130_fd_sc_lp__einvn_1.ext - technology: sky130A

.subckt sky130_fd_sc_lp__einvn_1 A TE_B VGND VNB VPB VPWR Z
M1000 a_166_73# A Z VNB nshort w=840000u l=150000u
+  ad=2.016e+11p pd=2.16e+06u as=2.226e+11p ps=2.21e+06u
M1001 VGND a_214_21# a_166_73# VNB nshort w=840000u l=150000u
+  ad=3.906e+11p pd=2.95e+06u as=0p ps=0u
M1002 a_214_21# TE_B VGND VNB nshort w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1003 a_214_21# TE_B VPWR VPB phighvt w=640000u l=150000u
+  ad=1.696e+11p pd=1.81e+06u as=4.9845e+11p ps=3.43e+06u
M1004 a_166_367# A Z VPB phighvt w=1.26e+06u l=150000u
+  ad=3.024e+11p pd=3e+06u as=3.339e+11p ps=3.05e+06u
M1005 VPWR TE_B a_166_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

