* File: sky130_fd_sc_lp__a311oi_4.pex.spice
* Created: Fri Aug 28 09:58:36 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A311OI_4%A3 1 3 6 8 10 13 15 17 20 22 24 27 29 30 31
+ 32 49
r80 49 50 10.4783 $w=3.22e-07 $l=7e-08 $layer=POLY_cond $X=1.765 $Y=1.35
+ $X2=1.835 $Y2=1.35
r81 47 49 13.472 $w=3.22e-07 $l=9e-08 $layer=POLY_cond $X=1.675 $Y=1.35
+ $X2=1.765 $Y2=1.35
r82 45 47 40.4161 $w=3.22e-07 $l=2.7e-07 $layer=POLY_cond $X=1.405 $Y=1.35
+ $X2=1.675 $Y2=1.35
r83 44 45 10.4783 $w=3.22e-07 $l=7e-08 $layer=POLY_cond $X=1.335 $Y=1.35
+ $X2=1.405 $Y2=1.35
r84 43 44 53.8882 $w=3.22e-07 $l=3.6e-07 $layer=POLY_cond $X=0.975 $Y=1.35
+ $X2=1.335 $Y2=1.35
r85 42 43 10.4783 $w=3.22e-07 $l=7e-08 $layer=POLY_cond $X=0.905 $Y=1.35
+ $X2=0.975 $Y2=1.35
r86 41 42 53.8882 $w=3.22e-07 $l=3.6e-07 $layer=POLY_cond $X=0.545 $Y=1.35
+ $X2=0.905 $Y2=1.35
r87 40 41 10.4783 $w=3.22e-07 $l=7e-08 $layer=POLY_cond $X=0.475 $Y=1.35
+ $X2=0.545 $Y2=1.35
r88 38 40 23.9503 $w=3.22e-07 $l=1.6e-07 $layer=POLY_cond $X=0.315 $Y=1.35
+ $X2=0.475 $Y2=1.35
r89 32 47 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=1.675
+ $Y=1.35 $X2=1.675 $Y2=1.35
r90 31 32 24.3294 $w=2.23e-07 $l=4.75e-07 $layer=LI1_cond $X=1.2 $Y=1.322
+ $X2=1.675 $Y2=1.322
r91 30 31 24.5855 $w=2.23e-07 $l=4.8e-07 $layer=LI1_cond $X=0.72 $Y=1.322
+ $X2=1.2 $Y2=1.322
r92 29 30 24.5855 $w=2.23e-07 $l=4.8e-07 $layer=LI1_cond $X=0.24 $Y=1.322
+ $X2=0.72 $Y2=1.322
r93 29 38 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=0.315
+ $Y=1.35 $X2=0.315 $Y2=1.35
r94 25 50 20.6399 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.835 $Y=1.515
+ $X2=1.835 $Y2=1.35
r95 25 27 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=1.835 $Y=1.515
+ $X2=1.835 $Y2=2.465
r96 22 49 20.6399 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.765 $Y=1.185
+ $X2=1.765 $Y2=1.35
r97 22 24 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.765 $Y=1.185
+ $X2=1.765 $Y2=0.655
r98 18 45 20.6399 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.405 $Y=1.515
+ $X2=1.405 $Y2=1.35
r99 18 20 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=1.405 $Y=1.515
+ $X2=1.405 $Y2=2.465
r100 15 44 20.6399 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.335 $Y=1.185
+ $X2=1.335 $Y2=1.35
r101 15 17 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.335 $Y=1.185
+ $X2=1.335 $Y2=0.655
r102 11 43 20.6399 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.975 $Y=1.515
+ $X2=0.975 $Y2=1.35
r103 11 13 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=0.975 $Y=1.515
+ $X2=0.975 $Y2=2.465
r104 8 42 20.6399 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.905 $Y=1.185
+ $X2=0.905 $Y2=1.35
r105 8 10 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.905 $Y=1.185
+ $X2=0.905 $Y2=0.655
r106 4 41 20.6399 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.545 $Y=1.515
+ $X2=0.545 $Y2=1.35
r107 4 6 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=0.545 $Y=1.515
+ $X2=0.545 $Y2=2.465
r108 1 40 20.6399 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=1.185
+ $X2=0.475 $Y2=1.35
r109 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.475 $Y=1.185
+ $X2=0.475 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__A311OI_4%A2 1 3 6 8 10 13 15 17 20 22 24 27 29 30 31
+ 32 50
r87 48 50 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=3.555 $Y=1.35
+ $X2=3.645 $Y2=1.35
r88 47 48 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=3.485 $Y=1.35
+ $X2=3.555 $Y2=1.35
r89 46 47 62.9501 $w=3.3e-07 $l=3.6e-07 $layer=POLY_cond $X=3.125 $Y=1.35
+ $X2=3.485 $Y2=1.35
r90 45 46 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=3.055 $Y=1.35
+ $X2=3.125 $Y2=1.35
r91 44 45 62.9501 $w=3.3e-07 $l=3.6e-07 $layer=POLY_cond $X=2.695 $Y=1.35
+ $X2=3.055 $Y2=1.35
r92 43 44 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=2.625 $Y=1.35
+ $X2=2.695 $Y2=1.35
r93 41 43 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.285 $Y=1.35
+ $X2=2.625 $Y2=1.35
r94 41 42 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=2.285
+ $Y=1.35 $X2=2.285 $Y2=1.35
r95 39 41 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=2.265 $Y=1.35
+ $X2=2.285 $Y2=1.35
r96 37 39 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=2.195 $Y=1.35
+ $X2=2.265 $Y2=1.35
r97 32 50 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=3.645
+ $Y=1.35 $X2=3.645 $Y2=1.35
r98 31 32 24.5855 $w=2.23e-07 $l=4.8e-07 $layer=LI1_cond $X=3.12 $Y=1.322
+ $X2=3.6 $Y2=1.322
r99 30 31 24.5855 $w=2.23e-07 $l=4.8e-07 $layer=LI1_cond $X=2.64 $Y=1.322
+ $X2=3.12 $Y2=1.322
r100 30 42 18.183 $w=2.23e-07 $l=3.55e-07 $layer=LI1_cond $X=2.64 $Y=1.322
+ $X2=2.285 $Y2=1.322
r101 29 42 6.40246 $w=2.23e-07 $l=1.25e-07 $layer=LI1_cond $X=2.16 $Y=1.322
+ $X2=2.285 $Y2=1.322
r102 25 48 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.555 $Y=1.515
+ $X2=3.555 $Y2=1.35
r103 25 27 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=3.555 $Y=1.515
+ $X2=3.555 $Y2=2.465
r104 22 47 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.485 $Y=1.185
+ $X2=3.485 $Y2=1.35
r105 22 24 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=3.485 $Y=1.185
+ $X2=3.485 $Y2=0.655
r106 18 46 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.125 $Y=1.515
+ $X2=3.125 $Y2=1.35
r107 18 20 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=3.125 $Y=1.515
+ $X2=3.125 $Y2=2.465
r108 15 45 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.055 $Y=1.185
+ $X2=3.055 $Y2=1.35
r109 15 17 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=3.055 $Y=1.185
+ $X2=3.055 $Y2=0.655
r110 11 44 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.695 $Y=1.515
+ $X2=2.695 $Y2=1.35
r111 11 13 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=2.695 $Y=1.515
+ $X2=2.695 $Y2=2.465
r112 8 43 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.625 $Y=1.185
+ $X2=2.625 $Y2=1.35
r113 8 10 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.625 $Y=1.185
+ $X2=2.625 $Y2=0.655
r114 4 39 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.265 $Y=1.515
+ $X2=2.265 $Y2=1.35
r115 4 6 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=2.265 $Y=1.515
+ $X2=2.265 $Y2=2.465
r116 1 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.195 $Y=1.185
+ $X2=2.195 $Y2=1.35
r117 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.195 $Y=1.185
+ $X2=2.195 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__A311OI_4%A1 3 5 6 7 9 12 14 16 19 21 23 26 28 30 31
+ 32 33 47
c86 33 0 1.95594e-19 $X=5.52 $Y=1.295
c87 6 0 1.70462e-19 $X=4.17 $Y=1.59
r88 45 47 16.2158 $w=4.31e-07 $l=1.45e-07 $layer=POLY_cond $X=5.385 $Y=1.425
+ $X2=5.53 $Y2=1.425
r89 44 45 10.065 $w=4.31e-07 $l=9e-08 $layer=POLY_cond $X=5.295 $Y=1.425
+ $X2=5.385 $Y2=1.425
r90 43 44 38.0232 $w=4.31e-07 $l=3.4e-07 $layer=POLY_cond $X=4.955 $Y=1.425
+ $X2=5.295 $Y2=1.425
r91 42 43 10.065 $w=4.31e-07 $l=9e-08 $layer=POLY_cond $X=4.865 $Y=1.425
+ $X2=4.955 $Y2=1.425
r92 41 42 38.0232 $w=4.31e-07 $l=3.4e-07 $layer=POLY_cond $X=4.525 $Y=1.425
+ $X2=4.865 $Y2=1.425
r93 39 41 1.67749 $w=4.31e-07 $l=1.5e-08 $layer=POLY_cond $X=4.51 $Y=1.425
+ $X2=4.525 $Y2=1.425
r94 37 39 8.38747 $w=4.31e-07 $l=7.5e-08 $layer=POLY_cond $X=4.435 $Y=1.425
+ $X2=4.51 $Y2=1.425
r95 33 47 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.53
+ $Y=1.35 $X2=5.53 $Y2=1.35
r96 32 33 24.5855 $w=2.23e-07 $l=4.8e-07 $layer=LI1_cond $X=5.04 $Y=1.322
+ $X2=5.52 $Y2=1.322
r97 31 32 27.1464 $w=2.23e-07 $l=5.3e-07 $layer=LI1_cond $X=4.51 $Y=1.322
+ $X2=5.04 $Y2=1.322
r98 31 39 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.51
+ $Y=1.35 $X2=4.51 $Y2=1.35
r99 28 47 21.8074 $w=4.31e-07 $l=3.2311e-07 $layer=POLY_cond $X=5.725 $Y=1.185
+ $X2=5.53 $Y2=1.425
r100 28 30 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=5.725 $Y=1.185
+ $X2=5.725 $Y2=0.655
r101 24 45 27.6969 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=5.385 $Y=1.665
+ $X2=5.385 $Y2=1.425
r102 24 26 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=5.385 $Y=1.665
+ $X2=5.385 $Y2=2.465
r103 21 44 27.6969 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=5.295 $Y=1.185
+ $X2=5.295 $Y2=1.425
r104 21 23 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=5.295 $Y=1.185
+ $X2=5.295 $Y2=0.655
r105 17 43 27.6969 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=4.955 $Y=1.665
+ $X2=4.955 $Y2=1.425
r106 17 19 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=4.955 $Y=1.665
+ $X2=4.955 $Y2=2.465
r107 14 42 27.6969 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=4.865 $Y=1.185
+ $X2=4.865 $Y2=1.425
r108 14 16 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=4.865 $Y=1.185
+ $X2=4.865 $Y2=0.655
r109 10 41 27.6969 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=4.525 $Y=1.665
+ $X2=4.525 $Y2=1.425
r110 10 12 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=4.525 $Y=1.665
+ $X2=4.525 $Y2=2.465
r111 7 37 27.6969 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=4.435 $Y=1.185
+ $X2=4.435 $Y2=1.425
r112 7 9 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=4.435 $Y=1.185
+ $X2=4.435 $Y2=0.655
r113 5 37 31.8532 $w=4.31e-07 $l=2.05122e-07 $layer=POLY_cond $X=4.345 $Y=1.59
+ $X2=4.435 $Y2=1.425
r114 5 6 89.734 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=4.345 $Y=1.59
+ $X2=4.17 $Y2=1.59
r115 1 6 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.095 $Y=1.665
+ $X2=4.17 $Y2=1.59
r116 1 3 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=4.095 $Y=1.665
+ $X2=4.095 $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__A311OI_4%B1 1 3 6 8 10 13 15 17 20 22 24 27 29 30 31
+ 32 49 51
c89 51 0 1.95594e-19 $X=7.625 $Y=1.35
r90 50 51 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=7.555 $Y=1.35
+ $X2=7.625 $Y2=1.35
r91 48 50 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=7.535 $Y=1.35
+ $X2=7.555 $Y2=1.35
r92 48 49 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=7.535
+ $Y=1.35 $X2=7.535 $Y2=1.35
r93 46 48 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=7.195 $Y=1.35
+ $X2=7.535 $Y2=1.35
r94 45 46 29.7264 $w=3.3e-07 $l=1.7e-07 $layer=POLY_cond $X=7.025 $Y=1.35
+ $X2=7.195 $Y2=1.35
r95 44 45 45.4639 $w=3.3e-07 $l=2.6e-07 $layer=POLY_cond $X=6.765 $Y=1.35
+ $X2=7.025 $Y2=1.35
r96 43 44 29.7264 $w=3.3e-07 $l=1.7e-07 $layer=POLY_cond $X=6.595 $Y=1.35
+ $X2=6.765 $Y2=1.35
r97 42 43 45.4639 $w=3.3e-07 $l=2.6e-07 $layer=POLY_cond $X=6.335 $Y=1.35
+ $X2=6.595 $Y2=1.35
r98 40 42 27.9778 $w=3.3e-07 $l=1.6e-07 $layer=POLY_cond $X=6.175 $Y=1.35
+ $X2=6.335 $Y2=1.35
r99 40 41 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=6.175
+ $Y=1.35 $X2=6.175 $Y2=1.35
r100 37 40 1.74861 $w=3.3e-07 $l=1e-08 $layer=POLY_cond $X=6.165 $Y=1.35
+ $X2=6.175 $Y2=1.35
r101 32 49 4.86587 $w=2.23e-07 $l=9.5e-08 $layer=LI1_cond $X=7.44 $Y=1.322
+ $X2=7.535 $Y2=1.322
r102 31 32 24.5855 $w=2.23e-07 $l=4.8e-07 $layer=LI1_cond $X=6.96 $Y=1.322
+ $X2=7.44 $Y2=1.322
r103 30 31 24.5855 $w=2.23e-07 $l=4.8e-07 $layer=LI1_cond $X=6.48 $Y=1.322
+ $X2=6.96 $Y2=1.322
r104 30 41 15.622 $w=2.23e-07 $l=3.05e-07 $layer=LI1_cond $X=6.48 $Y=1.322
+ $X2=6.175 $Y2=1.322
r105 29 41 8.96345 $w=2.23e-07 $l=1.75e-07 $layer=LI1_cond $X=6 $Y=1.322
+ $X2=6.175 $Y2=1.322
r106 25 51 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.625 $Y=1.515
+ $X2=7.625 $Y2=1.35
r107 25 27 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=7.625 $Y=1.515
+ $X2=7.625 $Y2=2.465
r108 22 50 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.555 $Y=1.185
+ $X2=7.555 $Y2=1.35
r109 22 24 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=7.555 $Y=1.185
+ $X2=7.555 $Y2=0.655
r110 18 46 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.195 $Y=1.515
+ $X2=7.195 $Y2=1.35
r111 18 20 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=7.195 $Y=1.515
+ $X2=7.195 $Y2=2.465
r112 15 45 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.025 $Y=1.185
+ $X2=7.025 $Y2=1.35
r113 15 17 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=7.025 $Y=1.185
+ $X2=7.025 $Y2=0.655
r114 11 44 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.765 $Y=1.515
+ $X2=6.765 $Y2=1.35
r115 11 13 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=6.765 $Y=1.515
+ $X2=6.765 $Y2=2.465
r116 8 43 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.595 $Y=1.185
+ $X2=6.595 $Y2=1.35
r117 8 10 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=6.595 $Y=1.185
+ $X2=6.595 $Y2=0.655
r118 4 42 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.335 $Y=1.515
+ $X2=6.335 $Y2=1.35
r119 4 6 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=6.335 $Y=1.515
+ $X2=6.335 $Y2=2.465
r120 1 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.165 $Y=1.185
+ $X2=6.165 $Y2=1.35
r121 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=6.165 $Y=1.185
+ $X2=6.165 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__A311OI_4%C1 1 3 6 8 10 13 15 17 20 22 24 27 29 30 31
+ 32 37 39
r83 52 53 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=9.275 $Y=1.35
+ $X2=9.345 $Y2=1.35
r84 51 52 62.9501 $w=3.3e-07 $l=3.6e-07 $layer=POLY_cond $X=8.915 $Y=1.35
+ $X2=9.275 $Y2=1.35
r85 50 51 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=8.845 $Y=1.35
+ $X2=8.915 $Y2=1.35
r86 49 50 62.9501 $w=3.3e-07 $l=3.6e-07 $layer=POLY_cond $X=8.485 $Y=1.35
+ $X2=8.845 $Y2=1.35
r87 48 49 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=8.415 $Y=1.35
+ $X2=8.485 $Y2=1.35
r88 46 48 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=8.075 $Y=1.35
+ $X2=8.415 $Y2=1.35
r89 46 47 48.4267 $w=1.7e-07 $l=5.1e-07 $layer=licon1_POLY $count=3 $X=8.075
+ $Y=1.35 $X2=8.075 $Y2=1.35
r90 44 46 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=8.055 $Y=1.35
+ $X2=8.075 $Y2=1.35
r91 42 44 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=7.985 $Y=1.35
+ $X2=8.055 $Y2=1.35
r92 37 53 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=9.42 $Y=1.35
+ $X2=9.345 $Y2=1.35
r93 37 39 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=9.42 $Y=1.35
+ $X2=9.775 $Y2=1.35
r94 32 39 48.4267 $w=1.7e-07 $l=5.1e-07 $layer=licon1_POLY $count=3 $X=9.775
+ $Y=1.35 $X2=9.775 $Y2=1.35
r95 31 32 21.2562 $w=2.23e-07 $l=4.15e-07 $layer=LI1_cond $X=9.36 $Y=1.322
+ $X2=9.775 $Y2=1.322
r96 30 31 24.5855 $w=2.23e-07 $l=4.8e-07 $layer=LI1_cond $X=8.88 $Y=1.322
+ $X2=9.36 $Y2=1.322
r97 29 30 24.5855 $w=2.23e-07 $l=4.8e-07 $layer=LI1_cond $X=8.4 $Y=1.322
+ $X2=8.88 $Y2=1.322
r98 29 47 16.6464 $w=2.23e-07 $l=3.25e-07 $layer=LI1_cond $X=8.4 $Y=1.322
+ $X2=8.075 $Y2=1.322
r99 25 53 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.345 $Y=1.515
+ $X2=9.345 $Y2=1.35
r100 25 27 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=9.345 $Y=1.515
+ $X2=9.345 $Y2=2.465
r101 22 52 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.275 $Y=1.185
+ $X2=9.275 $Y2=1.35
r102 22 24 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=9.275 $Y=1.185
+ $X2=9.275 $Y2=0.655
r103 18 51 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.915 $Y=1.515
+ $X2=8.915 $Y2=1.35
r104 18 20 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=8.915 $Y=1.515
+ $X2=8.915 $Y2=2.465
r105 15 50 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.845 $Y=1.185
+ $X2=8.845 $Y2=1.35
r106 15 17 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=8.845 $Y=1.185
+ $X2=8.845 $Y2=0.655
r107 11 49 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.485 $Y=1.515
+ $X2=8.485 $Y2=1.35
r108 11 13 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=8.485 $Y=1.515
+ $X2=8.485 $Y2=2.465
r109 8 48 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.415 $Y=1.185
+ $X2=8.415 $Y2=1.35
r110 8 10 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=8.415 $Y=1.185
+ $X2=8.415 $Y2=0.655
r111 4 44 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.055 $Y=1.515
+ $X2=8.055 $Y2=1.35
r112 4 6 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=8.055 $Y=1.515
+ $X2=8.055 $Y2=2.465
r113 1 42 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.985 $Y=1.185
+ $X2=7.985 $Y2=1.35
r114 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=7.985 $Y=1.185
+ $X2=7.985 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__A311OI_4%VPWR 1 2 3 4 5 6 7 22 24 30 36 42 48 52 56
+ 59 60 62 63 65 66 68 69 70 72 90 99 100 106 109
r145 109 110 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r146 106 107 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r147 103 104 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r148 99 100 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r149 97 100 1.07034 $w=4.9e-07 $l=3.84e-06 $layer=MET1_cond $X=6 $Y=3.33
+ $X2=9.84 $Y2=3.33
r150 97 110 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33
+ $X2=5.52 $Y2=3.33
r151 96 99 250.524 $w=1.68e-07 $l=3.84e-06 $layer=LI1_cond $X=6 $Y=3.33 $X2=9.84
+ $Y2=3.33
r152 96 97 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=6 $Y=3.33
+ $X2=6 $Y2=3.33
r153 94 109 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.765 $Y=3.33
+ $X2=5.6 $Y2=3.33
r154 94 96 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=5.765 $Y=3.33
+ $X2=6 $Y2=3.33
r155 90 109 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.435 $Y=3.33
+ $X2=5.6 $Y2=3.33
r156 90 92 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=5.435 $Y=3.33
+ $X2=5.04 $Y2=3.33
r157 88 89 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r158 86 89 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.56 $Y2=3.33
r159 85 86 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r160 83 86 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r161 82 83 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r162 80 83 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r163 80 107 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r164 79 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r165 77 106 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.355 $Y=3.33
+ $X2=1.19 $Y2=3.33
r166 77 79 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=1.355 $Y=3.33
+ $X2=1.68 $Y2=3.33
r167 76 107 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r168 76 104 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r169 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r170 73 103 4.62984 $w=1.7e-07 $l=2.48e-07 $layer=LI1_cond $X=0.495 $Y=3.33
+ $X2=0.247 $Y2=3.33
r171 73 75 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=0.495 $Y=3.33
+ $X2=0.72 $Y2=3.33
r172 72 106 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.025 $Y=3.33
+ $X2=1.19 $Y2=3.33
r173 72 75 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.025 $Y=3.33
+ $X2=0.72 $Y2=3.33
r174 70 110 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=5.52 $Y2=3.33
r175 70 89 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=4.56 $Y2=3.33
r176 70 92 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r177 68 88 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=4.575 $Y=3.33
+ $X2=4.56 $Y2=3.33
r178 68 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.575 $Y=3.33
+ $X2=4.74 $Y2=3.33
r179 67 92 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=4.905 $Y=3.33
+ $X2=5.04 $Y2=3.33
r180 67 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.905 $Y=3.33
+ $X2=4.74 $Y2=3.33
r181 65 85 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=3.66 $Y=3.33 $X2=3.6
+ $Y2=3.33
r182 65 66 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.66 $Y=3.33
+ $X2=3.825 $Y2=3.33
r183 64 88 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=3.99 $Y=3.33
+ $X2=4.56 $Y2=3.33
r184 64 66 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.99 $Y=3.33
+ $X2=3.825 $Y2=3.33
r185 62 82 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=2.745 $Y=3.33
+ $X2=2.64 $Y2=3.33
r186 62 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.745 $Y=3.33
+ $X2=2.91 $Y2=3.33
r187 61 85 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=3.075 $Y=3.33
+ $X2=3.6 $Y2=3.33
r188 61 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.075 $Y=3.33
+ $X2=2.91 $Y2=3.33
r189 59 79 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=1.885 $Y=3.33
+ $X2=1.68 $Y2=3.33
r190 59 60 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.885 $Y=3.33
+ $X2=2.05 $Y2=3.33
r191 58 82 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=2.215 $Y=3.33
+ $X2=2.64 $Y2=3.33
r192 58 60 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.215 $Y=3.33
+ $X2=2.05 $Y2=3.33
r193 54 109 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.6 $Y=3.245
+ $X2=5.6 $Y2=3.33
r194 54 56 29.8588 $w=3.28e-07 $l=8.55e-07 $layer=LI1_cond $X=5.6 $Y=3.245
+ $X2=5.6 $Y2=2.39
r195 50 69 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.74 $Y=3.245
+ $X2=4.74 $Y2=3.33
r196 50 52 29.8588 $w=3.28e-07 $l=8.55e-07 $layer=LI1_cond $X=4.74 $Y=3.245
+ $X2=4.74 $Y2=2.39
r197 46 66 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.825 $Y=3.245
+ $X2=3.825 $Y2=3.33
r198 46 48 29.8588 $w=3.28e-07 $l=8.55e-07 $layer=LI1_cond $X=3.825 $Y=3.245
+ $X2=3.825 $Y2=2.39
r199 42 45 32.1287 $w=3.28e-07 $l=9.2e-07 $layer=LI1_cond $X=2.91 $Y=2.03
+ $X2=2.91 $Y2=2.95
r200 40 63 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.91 $Y=3.245
+ $X2=2.91 $Y2=3.33
r201 40 45 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.91 $Y=3.245
+ $X2=2.91 $Y2=2.95
r202 36 39 32.1287 $w=3.28e-07 $l=9.2e-07 $layer=LI1_cond $X=2.05 $Y=2.03
+ $X2=2.05 $Y2=2.95
r203 34 60 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.05 $Y=3.245
+ $X2=2.05 $Y2=3.33
r204 34 39 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.05 $Y=3.245
+ $X2=2.05 $Y2=2.95
r205 30 33 32.1287 $w=3.28e-07 $l=9.2e-07 $layer=LI1_cond $X=1.19 $Y=2.03
+ $X2=1.19 $Y2=2.95
r206 28 106 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.19 $Y=3.245
+ $X2=1.19 $Y2=3.33
r207 28 33 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.19 $Y=3.245
+ $X2=1.19 $Y2=2.95
r208 24 27 33.8748 $w=3.28e-07 $l=9.7e-07 $layer=LI1_cond $X=0.33 $Y=1.98
+ $X2=0.33 $Y2=2.95
r209 22 103 3.13634 $w=3.3e-07 $l=1.19499e-07 $layer=LI1_cond $X=0.33 $Y=3.245
+ $X2=0.247 $Y2=3.33
r210 22 27 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.33 $Y=3.245
+ $X2=0.33 $Y2=2.95
r211 7 56 300 $w=1.7e-07 $l=6.21068e-07 $layer=licon1_PDIFF $count=2 $X=5.46
+ $Y=1.835 $X2=5.6 $Y2=2.39
r212 6 52 300 $w=1.7e-07 $l=6.21068e-07 $layer=licon1_PDIFF $count=2 $X=4.6
+ $Y=1.835 $X2=4.74 $Y2=2.39
r213 5 48 300 $w=1.7e-07 $l=6.45174e-07 $layer=licon1_PDIFF $count=2 $X=3.63
+ $Y=1.835 $X2=3.825 $Y2=2.39
r214 4 45 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=2.77
+ $Y=1.835 $X2=2.91 $Y2=2.95
r215 4 42 400 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_PDIFF $count=1 $X=2.77
+ $Y=1.835 $X2=2.91 $Y2=2.03
r216 3 39 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=1.91
+ $Y=1.835 $X2=2.05 $Y2=2.95
r217 3 36 400 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_PDIFF $count=1 $X=1.91
+ $Y=1.835 $X2=2.05 $Y2=2.03
r218 2 33 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=1.05
+ $Y=1.835 $X2=1.19 $Y2=2.95
r219 2 30 400 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_PDIFF $count=1 $X=1.05
+ $Y=1.835 $X2=1.19 $Y2=2.03
r220 1 27 400 $w=1.7e-07 $l=1.17584e-06 $layer=licon1_PDIFF $count=1 $X=0.205
+ $Y=1.835 $X2=0.33 $Y2=2.95
r221 1 24 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.205
+ $Y=1.835 $X2=0.33 $Y2=1.98
.ends

.subckt PM_SKY130_FD_SC_LP__A311OI_4%A_124_367# 1 2 3 4 5 6 7 8 27 31 32 35 39
+ 43 47 50 53 55 59 61 65 67 71 73 77 78 80 82 84 86 88
c113 47 0 1.70462e-19 $X=3.245 $Y=1.69
r114 74 86 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=6.645 $Y=2.03
+ $X2=6.55 $Y2=2.03
r115 73 88 3.61205 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=7.315 $Y=2.03
+ $X2=7.41 $Y2=2.03
r116 73 74 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=7.315 $Y=2.03
+ $X2=6.645 $Y2=2.03
r117 69 86 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=6.55 $Y=2.115
+ $X2=6.55 $Y2=2.03
r118 69 71 26.5598 $w=1.88e-07 $l=4.55e-07 $layer=LI1_cond $X=6.55 $Y=2.115
+ $X2=6.55 $Y2=2.57
r119 68 84 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=5.265 $Y=2.03
+ $X2=5.17 $Y2=2.03
r120 67 86 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=6.455 $Y=2.03
+ $X2=6.55 $Y2=2.03
r121 67 68 77.6364 $w=1.68e-07 $l=1.19e-06 $layer=LI1_cond $X=6.455 $Y=2.03
+ $X2=5.265 $Y2=2.03
r122 63 84 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=5.17 $Y=2.115
+ $X2=5.17 $Y2=2.03
r123 63 65 23.3493 $w=1.88e-07 $l=4e-07 $layer=LI1_cond $X=5.17 $Y=2.115
+ $X2=5.17 $Y2=2.515
r124 62 82 6.92067 $w=1.7e-07 $l=1.23e-07 $layer=LI1_cond $X=4.405 $Y=2.03
+ $X2=4.282 $Y2=2.03
r125 61 84 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=5.075 $Y=2.03
+ $X2=5.17 $Y2=2.03
r126 61 62 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.075 $Y=2.03
+ $X2=4.405 $Y2=2.03
r127 57 82 0.066131 $w=2.45e-07 $l=8.5e-08 $layer=LI1_cond $X=4.282 $Y=2.115
+ $X2=4.282 $Y2=2.03
r128 57 59 18.8154 $w=2.43e-07 $l=4e-07 $layer=LI1_cond $X=4.282 $Y=2.115
+ $X2=4.282 $Y2=2.515
r129 56 80 2.79892 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.505 $Y=2.03
+ $X2=3.375 $Y2=2.03
r130 55 82 6.92067 $w=1.7e-07 $l=1.22e-07 $layer=LI1_cond $X=4.16 $Y=2.03
+ $X2=4.282 $Y2=2.03
r131 55 56 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=4.16 $Y=2.03
+ $X2=3.505 $Y2=2.03
r132 51 80 3.67481 $w=2.52e-07 $l=8.89101e-08 $layer=LI1_cond $X=3.367 $Y=2.115
+ $X2=3.375 $Y2=2.03
r133 51 53 37.3956 $w=2.43e-07 $l=7.95e-07 $layer=LI1_cond $X=3.367 $Y=2.115
+ $X2=3.367 $Y2=2.91
r134 50 80 3.67481 $w=2.52e-07 $l=8.5e-08 $layer=LI1_cond $X=3.375 $Y=1.945
+ $X2=3.375 $Y2=2.03
r135 49 50 7.5352 $w=2.58e-07 $l=1.7e-07 $layer=LI1_cond $X=3.375 $Y=1.775
+ $X2=3.375 $Y2=1.945
r136 48 78 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.575 $Y=1.69
+ $X2=2.48 $Y2=1.69
r137 47 49 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=3.245 $Y=1.69
+ $X2=3.375 $Y2=1.775
r138 47 48 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.245 $Y=1.69
+ $X2=2.575 $Y2=1.69
r139 43 45 54.2871 $w=1.88e-07 $l=9.3e-07 $layer=LI1_cond $X=2.48 $Y=1.98
+ $X2=2.48 $Y2=2.91
r140 41 78 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=2.48 $Y=1.775
+ $X2=2.48 $Y2=1.69
r141 41 43 11.9665 $w=1.88e-07 $l=2.05e-07 $layer=LI1_cond $X=2.48 $Y=1.775
+ $X2=2.48 $Y2=1.98
r142 40 77 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.715 $Y=1.69
+ $X2=1.62 $Y2=1.69
r143 39 78 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.385 $Y=1.69
+ $X2=2.48 $Y2=1.69
r144 39 40 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.385 $Y=1.69
+ $X2=1.715 $Y2=1.69
r145 35 37 54.2871 $w=1.88e-07 $l=9.3e-07 $layer=LI1_cond $X=1.62 $Y=1.98
+ $X2=1.62 $Y2=2.91
r146 33 77 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.62 $Y=1.775
+ $X2=1.62 $Y2=1.69
r147 33 35 11.9665 $w=1.88e-07 $l=2.05e-07 $layer=LI1_cond $X=1.62 $Y=1.775
+ $X2=1.62 $Y2=1.98
r148 31 77 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.525 $Y=1.69
+ $X2=1.62 $Y2=1.69
r149 31 32 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.525 $Y=1.69
+ $X2=0.855 $Y2=1.69
r150 27 29 54.2871 $w=1.88e-07 $l=9.3e-07 $layer=LI1_cond $X=0.76 $Y=1.98
+ $X2=0.76 $Y2=2.91
r151 25 32 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=0.76 $Y=1.775
+ $X2=0.855 $Y2=1.69
r152 25 27 11.9665 $w=1.88e-07 $l=2.05e-07 $layer=LI1_cond $X=0.76 $Y=1.775
+ $X2=0.76 $Y2=1.98
r153 8 88 300 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=2 $X=7.27
+ $Y=1.835 $X2=7.41 $Y2=2.11
r154 7 86 600 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_PDIFF $count=1 $X=6.41
+ $Y=1.835 $X2=6.55 $Y2=2.03
r155 7 71 600 $w=1.7e-07 $l=8.01951e-07 $layer=licon1_PDIFF $count=1 $X=6.41
+ $Y=1.835 $X2=6.55 $Y2=2.57
r156 6 84 600 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_PDIFF $count=1 $X=5.03
+ $Y=1.835 $X2=5.17 $Y2=2.03
r157 6 65 300 $w=1.7e-07 $l=7.46726e-07 $layer=licon1_PDIFF $count=2 $X=5.03
+ $Y=1.835 $X2=5.17 $Y2=2.515
r158 5 82 600 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_PDIFF $count=1 $X=4.17
+ $Y=1.835 $X2=4.31 $Y2=2.03
r159 5 59 300 $w=1.7e-07 $l=7.46726e-07 $layer=licon1_PDIFF $count=2 $X=4.17
+ $Y=1.835 $X2=4.31 $Y2=2.515
r160 4 80 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=3.2
+ $Y=1.835 $X2=3.34 $Y2=1.98
r161 4 53 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=3.2
+ $Y=1.835 $X2=3.34 $Y2=2.91
r162 3 45 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=2.34
+ $Y=1.835 $X2=2.48 $Y2=2.91
r163 3 43 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.34
+ $Y=1.835 $X2=2.48 $Y2=1.98
r164 2 37 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=1.48
+ $Y=1.835 $X2=1.62 $Y2=2.91
r165 2 35 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.48
+ $Y=1.835 $X2=1.62 $Y2=1.98
r166 1 29 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=0.62
+ $Y=1.835 $X2=0.76 $Y2=2.91
r167 1 27 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.62
+ $Y=1.835 $X2=0.76 $Y2=1.98
.ends

.subckt PM_SKY130_FD_SC_LP__A311OI_4%A_1199_367# 1 2 3 4 5 18 20 21 24 26 30 32
+ 36 38 40 42 44 46 48
r77 40 50 2.74877 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=9.58 $Y=2.905
+ $X2=9.58 $Y2=2.99
r78 40 42 36.759 $w=2.88e-07 $l=9.25e-07 $layer=LI1_cond $X=9.58 $Y=2.905
+ $X2=9.58 $Y2=1.98
r79 39 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.865 $Y=2.99
+ $X2=8.7 $Y2=2.99
r80 38 50 4.68908 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=9.435 $Y=2.99
+ $X2=9.58 $Y2=2.99
r81 38 39 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=9.435 $Y=2.99
+ $X2=8.865 $Y2=2.99
r82 34 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.7 $Y=2.905 $X2=8.7
+ $Y2=2.99
r83 34 36 30.5572 $w=3.28e-07 $l=8.75e-07 $layer=LI1_cond $X=8.7 $Y=2.905
+ $X2=8.7 $Y2=2.03
r84 33 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.005 $Y=2.99
+ $X2=7.84 $Y2=2.99
r85 32 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.535 $Y=2.99
+ $X2=8.7 $Y2=2.99
r86 32 33 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=8.535 $Y=2.99
+ $X2=8.005 $Y2=2.99
r87 28 46 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.84 $Y=2.905
+ $X2=7.84 $Y2=2.99
r88 28 30 30.5572 $w=3.28e-07 $l=8.75e-07 $layer=LI1_cond $X=7.84 $Y=2.905
+ $X2=7.84 $Y2=2.03
r89 27 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.145 $Y=2.99
+ $X2=6.98 $Y2=2.99
r90 26 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.675 $Y=2.99
+ $X2=7.84 $Y2=2.99
r91 26 27 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=7.675 $Y=2.99
+ $X2=7.145 $Y2=2.99
r92 22 44 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.98 $Y=2.905
+ $X2=6.98 $Y2=2.99
r93 22 24 17.9851 $w=3.28e-07 $l=5.15e-07 $layer=LI1_cond $X=6.98 $Y=2.905
+ $X2=6.98 $Y2=2.39
r94 20 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.815 $Y=2.99
+ $X2=6.98 $Y2=2.99
r95 20 21 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=6.815 $Y=2.99
+ $X2=6.285 $Y2=2.99
r96 16 21 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.12 $Y=2.905
+ $X2=6.285 $Y2=2.99
r97 16 18 17.9851 $w=3.28e-07 $l=5.15e-07 $layer=LI1_cond $X=6.12 $Y=2.905
+ $X2=6.12 $Y2=2.39
r98 5 50 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=9.42
+ $Y=1.835 $X2=9.56 $Y2=2.91
r99 5 42 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=9.42
+ $Y=1.835 $X2=9.56 $Y2=1.98
r100 4 48 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=8.56
+ $Y=1.835 $X2=8.7 $Y2=2.95
r101 4 36 400 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_PDIFF $count=1 $X=8.56
+ $Y=1.835 $X2=8.7 $Y2=2.03
r102 3 46 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=7.7
+ $Y=1.835 $X2=7.84 $Y2=2.95
r103 3 30 400 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_PDIFF $count=1 $X=7.7
+ $Y=1.835 $X2=7.84 $Y2=2.03
r104 2 24 300 $w=1.7e-07 $l=6.21068e-07 $layer=licon1_PDIFF $count=2 $X=6.84
+ $Y=1.835 $X2=6.98 $Y2=2.39
r105 1 18 300 $w=1.7e-07 $l=6.14329e-07 $layer=licon1_PDIFF $count=2 $X=5.995
+ $Y=1.835 $X2=6.12 $Y2=2.39
.ends

.subckt PM_SKY130_FD_SC_LP__A311OI_4%Y 1 2 3 4 5 6 7 8 9 28 29 30 32 36 38 42 44
+ 48 50 54 56 60 62 66 70 77 80 84 85 86 87 88 89
r144 80 82 5.98384 $w=2.58e-07 $l=1.35e-07 $layer=LI1_cond $X=5.08 $Y=0.82
+ $X2=5.08 $Y2=0.955
r145 78 89 19.101 $w=1.78e-07 $l=3.1e-07 $layer=LI1_cond $X=4.085 $Y=1.605
+ $X2=4.085 $Y2=1.295
r146 76 77 7.69093 $w=3.83e-07 $l=1.35e-07 $layer=LI1_cond $X=4.22 $Y=0.847
+ $X2=4.355 $Y2=0.847
r147 73 89 15.7121 $w=1.78e-07 $l=2.55e-07 $layer=LI1_cond $X=4.085 $Y=1.04
+ $X2=4.085 $Y2=1.295
r148 72 76 4.04103 $w=3.83e-07 $l=1.35e-07 $layer=LI1_cond $X=4.085 $Y=0.847
+ $X2=4.22 $Y2=0.847
r149 72 73 5.20241 $w=1.8e-07 $l=1.93e-07 $layer=LI1_cond $X=4.085 $Y=0.847
+ $X2=4.085 $Y2=1.04
r150 68 70 19.9461 $w=2.58e-07 $l=4.5e-07 $layer=LI1_cond $X=9.525 $Y=0.87
+ $X2=9.525 $Y2=0.42
r151 64 66 10.2718 $w=2.28e-07 $l=2.05e-07 $layer=LI1_cond $X=9.15 $Y=1.775
+ $X2=9.15 $Y2=1.98
r152 63 88 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=8.725 $Y=0.955
+ $X2=8.63 $Y2=0.955
r153 62 68 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=9.395 $Y=0.955
+ $X2=9.525 $Y2=0.87
r154 62 63 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=9.395 $Y=0.955
+ $X2=8.725 $Y2=0.955
r155 58 88 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=8.63 $Y=0.87
+ $X2=8.63 $Y2=0.955
r156 58 60 26.2679 $w=1.88e-07 $l=4.5e-07 $layer=LI1_cond $X=8.63 $Y=0.87
+ $X2=8.63 $Y2=0.42
r157 57 87 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=8.365 $Y=1.69
+ $X2=8.27 $Y2=1.69
r158 56 64 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=9.035 $Y=1.69
+ $X2=9.15 $Y2=1.775
r159 56 57 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=9.035 $Y=1.69
+ $X2=8.365 $Y2=1.69
r160 52 87 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=8.27 $Y=1.775
+ $X2=8.27 $Y2=1.69
r161 52 54 11.9665 $w=1.88e-07 $l=2.05e-07 $layer=LI1_cond $X=8.27 $Y=1.775
+ $X2=8.27 $Y2=1.98
r162 51 86 6.92067 $w=1.7e-07 $l=1.23e-07 $layer=LI1_cond $X=7.865 $Y=0.955
+ $X2=7.742 $Y2=0.955
r163 50 88 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=8.535 $Y=0.955
+ $X2=8.63 $Y2=0.955
r164 50 51 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=8.535 $Y=0.955
+ $X2=7.865 $Y2=0.955
r165 46 86 0.066131 $w=2.45e-07 $l=8.5e-08 $layer=LI1_cond $X=7.742 $Y=0.87
+ $X2=7.742 $Y2=0.955
r166 46 48 21.1673 $w=2.43e-07 $l=4.5e-07 $layer=LI1_cond $X=7.742 $Y=0.87
+ $X2=7.742 $Y2=0.42
r167 45 85 6.70225 $w=1.7e-07 $l=1.18e-07 $layer=LI1_cond $X=6.95 $Y=0.955
+ $X2=6.832 $Y2=0.955
r168 44 86 6.92067 $w=1.7e-07 $l=1.22e-07 $layer=LI1_cond $X=7.62 $Y=0.955
+ $X2=7.742 $Y2=0.955
r169 44 45 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=7.62 $Y=0.955
+ $X2=6.95 $Y2=0.955
r170 40 85 0.207053 $w=2.35e-07 $l=8.5e-08 $layer=LI1_cond $X=6.832 $Y=0.87
+ $X2=6.832 $Y2=0.955
r171 40 42 22.0681 $w=2.33e-07 $l=4.5e-07 $layer=LI1_cond $X=6.832 $Y=0.87
+ $X2=6.832 $Y2=0.42
r172 39 84 6.81202 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=6.045 $Y=0.955
+ $X2=5.925 $Y2=0.955
r173 38 85 6.70225 $w=1.7e-07 $l=1.17e-07 $layer=LI1_cond $X=6.715 $Y=0.955
+ $X2=6.832 $Y2=0.955
r174 38 39 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=6.715 $Y=0.955
+ $X2=6.045 $Y2=0.955
r175 34 84 0.135687 $w=2.4e-07 $l=8.5e-08 $layer=LI1_cond $X=5.925 $Y=0.87
+ $X2=5.925 $Y2=0.955
r176 34 36 21.6083 $w=2.38e-07 $l=4.5e-07 $layer=LI1_cond $X=5.925 $Y=0.87
+ $X2=5.925 $Y2=0.42
r177 33 82 3.22376 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=5.21 $Y=0.955
+ $X2=5.08 $Y2=0.955
r178 32 84 6.81202 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=5.805 $Y=0.955
+ $X2=5.925 $Y2=0.955
r179 32 33 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=5.805 $Y=0.955
+ $X2=5.21 $Y2=0.955
r180 30 82 3.22376 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=4.95 $Y=0.955
+ $X2=5.08 $Y2=0.955
r181 30 77 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=4.95 $Y=0.955
+ $X2=4.355 $Y2=0.955
r182 29 78 6.82373 $w=1.7e-07 $l=1.25499e-07 $layer=LI1_cond $X=4.175 $Y=1.69
+ $X2=4.085 $Y2=1.605
r183 28 87 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=8.175 $Y=1.69
+ $X2=8.27 $Y2=1.69
r184 28 29 260.963 $w=1.68e-07 $l=4e-06 $layer=LI1_cond $X=8.175 $Y=1.69
+ $X2=4.175 $Y2=1.69
r185 9 66 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=8.99
+ $Y=1.835 $X2=9.13 $Y2=1.98
r186 8 54 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=8.13
+ $Y=1.835 $X2=8.27 $Y2=1.98
r187 7 70 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=9.35
+ $Y=0.235 $X2=9.49 $Y2=0.42
r188 6 60 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=8.49
+ $Y=0.235 $X2=8.63 $Y2=0.42
r189 5 48 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=7.63
+ $Y=0.235 $X2=7.77 $Y2=0.42
r190 4 42 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=6.67
+ $Y=0.235 $X2=6.81 $Y2=0.42
r191 3 36 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=5.8
+ $Y=0.235 $X2=5.94 $Y2=0.42
r192 2 80 182 $w=1.7e-07 $l=6.51249e-07 $layer=licon1_NDIFF $count=1 $X=4.94
+ $Y=0.235 $X2=5.08 $Y2=0.82
r193 1 76 182 $w=1.7e-07 $l=6.44477e-07 $layer=licon1_NDIFF $count=1 $X=4.095
+ $Y=0.235 $X2=4.22 $Y2=0.82
.ends

.subckt PM_SKY130_FD_SC_LP__A311OI_4%A_27_47# 1 2 3 4 5 18 20 21 24 26 30 32 34
+ 36 37 39 44
r56 34 44 5.64923 $w=2.53e-07 $l=1.25e-07 $layer=LI1_cond $X=3.697 $Y=0.955
+ $X2=3.697 $Y2=0.83
r57 34 35 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=3.57 $Y=0.955
+ $X2=2.965 $Y2=0.955
r58 33 37 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=2.115 $Y=0.955 $X2=2
+ $Y2=0.955
r59 32 35 3.11056 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=2.837 $Y=0.955
+ $X2=2.965 $Y2=0.955
r60 32 39 5.64923 $w=2.53e-07 $l=1.25e-07 $layer=LI1_cond $X=2.837 $Y=0.955
+ $X2=2.837 $Y2=0.83
r61 32 33 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=2.71 $Y=0.955
+ $X2=2.115 $Y2=0.955
r62 28 37 0.280307 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2 $Y=0.87 $X2=2
+ $Y2=0.955
r63 28 30 22.5478 $w=2.28e-07 $l=4.5e-07 $layer=LI1_cond $X=2 $Y=0.87 $X2=2
+ $Y2=0.42
r64 27 36 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.215 $Y=0.955
+ $X2=1.12 $Y2=0.955
r65 26 37 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=1.885 $Y=0.955 $X2=2
+ $Y2=0.955
r66 26 27 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.885 $Y=0.955
+ $X2=1.215 $Y2=0.955
r67 22 36 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.12 $Y=0.87
+ $X2=1.12 $Y2=0.955
r68 22 24 26.2679 $w=1.88e-07 $l=4.5e-07 $layer=LI1_cond $X=1.12 $Y=0.87
+ $X2=1.12 $Y2=0.42
r69 20 36 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.025 $Y=0.955
+ $X2=1.12 $Y2=0.955
r70 20 21 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.025 $Y=0.955
+ $X2=0.355 $Y2=0.955
r71 16 21 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=0.225 $Y=0.87
+ $X2=0.355 $Y2=0.955
r72 16 18 19.9461 $w=2.58e-07 $l=4.5e-07 $layer=LI1_cond $X=0.225 $Y=0.87
+ $X2=0.225 $Y2=0.42
r73 5 44 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=3.56
+ $Y=0.235 $X2=3.7 $Y2=0.83
r74 4 39 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=2.7
+ $Y=0.235 $X2=2.84 $Y2=0.83
r75 3 30 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=1.84
+ $Y=0.235 $X2=1.98 $Y2=0.42
r76 2 24 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=0.98
+ $Y=0.235 $X2=1.12 $Y2=0.42
r77 1 18 91 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__A311OI_4%VGND 1 2 3 4 5 6 21 25 29 33 37 41 44 45 47
+ 48 50 51 53 54 55 57 62 81 82 85 88
r132 88 89 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r133 85 86 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r134 81 82 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.84 $Y=0 $X2=9.84
+ $Y2=0
r135 79 82 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=8.88 $Y=0 $X2=9.84
+ $Y2=0
r136 78 79 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.88 $Y=0 $X2=8.88
+ $Y2=0
r137 76 79 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=8.88
+ $Y2=0
r138 75 76 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r139 73 76 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=7.92
+ $Y2=0
r140 72 73 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r141 70 73 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.96
+ $Y2=0
r142 69 70 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=6 $Y=0 $X2=6 $Y2=0
r143 67 88 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.715 $Y=0 $X2=1.55
+ $Y2=0
r144 67 69 279.556 $w=1.68e-07 $l=4.285e-06 $layer=LI1_cond $X=1.715 $Y=0 $X2=6
+ $Y2=0
r145 66 89 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r146 66 86 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r147 65 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r148 63 85 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.855 $Y=0 $X2=0.69
+ $Y2=0
r149 63 65 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.855 $Y=0 $X2=1.2
+ $Y2=0
r150 62 88 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.385 $Y=0 $X2=1.55
+ $Y2=0
r151 62 65 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=1.385 $Y=0 $X2=1.2
+ $Y2=0
r152 60 86 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r153 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r154 57 85 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.525 $Y=0 $X2=0.69
+ $Y2=0
r155 57 59 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.525 $Y=0
+ $X2=0.24 $Y2=0
r156 55 70 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=6
+ $Y2=0
r157 55 89 0.936549 $w=4.9e-07 $l=3.36e-06 $layer=MET1_cond $X=5.04 $Y=0
+ $X2=1.68 $Y2=0
r158 53 78 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=8.895 $Y=0 $X2=8.88
+ $Y2=0
r159 53 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.895 $Y=0 $X2=9.06
+ $Y2=0
r160 52 81 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=9.225 $Y=0 $X2=9.84
+ $Y2=0
r161 52 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.225 $Y=0 $X2=9.06
+ $Y2=0
r162 50 75 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=8.035 $Y=0
+ $X2=7.92 $Y2=0
r163 50 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.035 $Y=0 $X2=8.2
+ $Y2=0
r164 49 78 33.5989 $w=1.68e-07 $l=5.15e-07 $layer=LI1_cond $X=8.365 $Y=0
+ $X2=8.88 $Y2=0
r165 49 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.365 $Y=0 $X2=8.2
+ $Y2=0
r166 47 72 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=7.12 $Y=0 $X2=6.96
+ $Y2=0
r167 47 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.12 $Y=0 $X2=7.285
+ $Y2=0
r168 46 75 30.6631 $w=1.68e-07 $l=4.7e-07 $layer=LI1_cond $X=7.45 $Y=0 $X2=7.92
+ $Y2=0
r169 46 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.45 $Y=0 $X2=7.285
+ $Y2=0
r170 44 69 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=6.215 $Y=0 $X2=6
+ $Y2=0
r171 44 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.215 $Y=0 $X2=6.38
+ $Y2=0
r172 43 72 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=6.545 $Y=0
+ $X2=6.96 $Y2=0
r173 43 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.545 $Y=0 $X2=6.38
+ $Y2=0
r174 39 54 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.06 $Y=0.085
+ $X2=9.06 $Y2=0
r175 39 41 17.112 $w=3.28e-07 $l=4.9e-07 $layer=LI1_cond $X=9.06 $Y=0.085
+ $X2=9.06 $Y2=0.575
r176 35 51 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.2 $Y=0.085 $X2=8.2
+ $Y2=0
r177 35 37 17.112 $w=3.28e-07 $l=4.9e-07 $layer=LI1_cond $X=8.2 $Y=0.085 $X2=8.2
+ $Y2=0.575
r178 31 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.285 $Y=0.085
+ $X2=7.285 $Y2=0
r179 31 33 17.112 $w=3.28e-07 $l=4.9e-07 $layer=LI1_cond $X=7.285 $Y=0.085
+ $X2=7.285 $Y2=0.575
r180 27 45 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.38 $Y=0.085
+ $X2=6.38 $Y2=0
r181 27 29 17.112 $w=3.28e-07 $l=4.9e-07 $layer=LI1_cond $X=6.38 $Y=0.085
+ $X2=6.38 $Y2=0.575
r182 23 88 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.55 $Y=0.085
+ $X2=1.55 $Y2=0
r183 23 25 17.112 $w=3.28e-07 $l=4.9e-07 $layer=LI1_cond $X=1.55 $Y=0.085
+ $X2=1.55 $Y2=0.575
r184 19 85 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=0.085
+ $X2=0.69 $Y2=0
r185 19 21 17.112 $w=3.28e-07 $l=4.9e-07 $layer=LI1_cond $X=0.69 $Y=0.085
+ $X2=0.69 $Y2=0.575
r186 6 41 182 $w=1.7e-07 $l=4.0398e-07 $layer=licon1_NDIFF $count=1 $X=8.92
+ $Y=0.235 $X2=9.06 $Y2=0.575
r187 5 37 182 $w=1.7e-07 $l=4.0398e-07 $layer=licon1_NDIFF $count=1 $X=8.06
+ $Y=0.235 $X2=8.2 $Y2=0.575
r188 4 33 182 $w=1.7e-07 $l=4.22493e-07 $layer=licon1_NDIFF $count=1 $X=7.1
+ $Y=0.235 $X2=7.285 $Y2=0.575
r189 3 29 182 $w=1.7e-07 $l=4.0398e-07 $layer=licon1_NDIFF $count=1 $X=6.24
+ $Y=0.235 $X2=6.38 $Y2=0.575
r190 2 25 182 $w=1.7e-07 $l=4.0398e-07 $layer=licon1_NDIFF $count=1 $X=1.41
+ $Y=0.235 $X2=1.55 $Y2=0.575
r191 1 21 182 $w=1.7e-07 $l=4.0398e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.235 $X2=0.69 $Y2=0.575
.ends

.subckt PM_SKY130_FD_SC_LP__A311OI_4%A_454_47# 1 2 3 4 13 15 17 19
r38 26 28 7.17559 $w=2.63e-07 $l=1.65e-07 $layer=LI1_cond $X=3.267 $Y=0.37
+ $X2=3.267 $Y2=0.535
r39 19 22 8.36086 $w=2.53e-07 $l=1.85e-07 $layer=LI1_cond $X=2.412 $Y=0.35
+ $X2=2.412 $Y2=0.535
r40 17 38 7.45698 $w=2.53e-07 $l=1.65e-07 $layer=LI1_cond $X=5.507 $Y=0.37
+ $X2=5.507 $Y2=0.535
r41 17 18 30.0637 $w=2.28e-07 $l=6e-07 $layer=LI1_cond $X=5.38 $Y=0.37 $X2=4.78
+ $Y2=0.37
r42 16 26 1.56657 $w=2.3e-07 $l=1.33e-07 $layer=LI1_cond $X=3.4 $Y=0.37
+ $X2=3.267 $Y2=0.37
r43 15 33 7.45698 $w=2.53e-07 $l=1.65e-07 $layer=LI1_cond $X=4.652 $Y=0.37
+ $X2=4.652 $Y2=0.535
r44 15 18 1.33812 $w=2.3e-07 $l=1.28e-07 $layer=LI1_cond $X=4.652 $Y=0.37
+ $X2=4.78 $Y2=0.37
r45 15 16 56.3695 $w=2.28e-07 $l=1.125e-06 $layer=LI1_cond $X=4.525 $Y=0.37
+ $X2=3.4 $Y2=0.37
r46 14 19 2.46227 $w=1.9e-07 $l=1.28e-07 $layer=LI1_cond $X=2.54 $Y=0.35
+ $X2=2.412 $Y2=0.35
r47 13 26 0.869768 $w=2.63e-07 $l=2e-08 $layer=LI1_cond $X=3.267 $Y=0.35
+ $X2=3.267 $Y2=0.37
r48 13 14 34.7321 $w=1.88e-07 $l=5.95e-07 $layer=LI1_cond $X=3.135 $Y=0.35
+ $X2=2.54 $Y2=0.35
r49 4 38 182 $w=1.7e-07 $l=3.63318e-07 $layer=licon1_NDIFF $count=1 $X=5.37
+ $Y=0.235 $X2=5.51 $Y2=0.535
r50 3 33 182 $w=1.7e-07 $l=3.63318e-07 $layer=licon1_NDIFF $count=1 $X=4.51
+ $Y=0.235 $X2=4.65 $Y2=0.535
r51 2 28 182 $w=1.7e-07 $l=3.63318e-07 $layer=licon1_NDIFF $count=1 $X=3.13
+ $Y=0.235 $X2=3.27 $Y2=0.535
r52 1 22 182 $w=1.7e-07 $l=3.63318e-07 $layer=licon1_NDIFF $count=1 $X=2.27
+ $Y=0.235 $X2=2.41 $Y2=0.535
.ends

