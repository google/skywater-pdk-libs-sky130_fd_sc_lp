* File: sky130_fd_sc_lp__nand2b_lp.spice
* Created: Fri Aug 28 10:48:31 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__nand2b_lp.pex.spice"
.subckt sky130_fd_sc_lp__nand2b_lp  VNB VPB A_N B VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B	B
* A_N	A_N
* VPB	VPB
* VNB	VNB
MM1000 A_119_51# N_A_N_M1000_g N_A_32_51#_M1000_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1197 PD=0.63 PS=1.41 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1005 N_VGND_M1005_d N_A_N_M1005_g A_119_51# VNB NSHORT L=0.15 W=0.42 AD=0.0588
+ AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6 SB=75001 A=0.063
+ P=1.14 MULT=1
MM1001 A_277_51# N_B_M1001_g N_VGND_M1005_d VNB NSHORT L=0.15 W=0.42 AD=0.0504
+ AS=0.0588 PD=0.66 PS=0.7 NRD=18.564 NRS=0 M=1 R=2.8 SA=75001 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1002 N_Y_M1002_d N_A_32_51#_M1002_g A_277_51# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0504 PD=1.41 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75001.4
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1003 N_VPWR_M1003_d N_A_N_M1003_g N_A_32_51#_M1003_s VPB PHIGHVT L=0.25 W=1
+ AD=0.14 AS=0.285 PD=1.28 PS=2.57 NRD=0 NRS=0 M=1 R=4 SA=125000 SB=125001
+ A=0.25 P=2.5 MULT=1
MM1006 N_Y_M1006_d N_B_M1006_g N_VPWR_M1003_d VPB PHIGHVT L=0.25 W=1 AD=0.14
+ AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125001 SB=125001 A=0.25 P=2.5
+ MULT=1
MM1004 N_VPWR_M1004_d N_A_32_51#_M1004_g N_Y_M1006_d VPB PHIGHVT L=0.25 W=1
+ AD=0.35 AS=0.14 PD=2.7 PS=1.28 NRD=12.7853 NRS=0 M=1 R=4 SA=125001 SB=125000
+ A=0.25 P=2.5 MULT=1
DX7_noxref VNB VPB NWDIODE A=5.1847 P=9.29
*
.include "sky130_fd_sc_lp__nand2b_lp.pxi.spice"
*
.ends
*
*
