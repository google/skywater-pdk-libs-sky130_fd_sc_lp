* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__a211o_lp A1 A2 B1 C1 VGND VNB VPB VPWR X
M1000 VPWR A1 a_29_409# VPB phighvt w=1e+06u l=250000u
+  ad=6.15e+11p pd=5.23e+06u as=5.65e+11p ps=5.13e+06u
M1001 a_130_57# A1 a_43_57# VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=2.373e+11p ps=2.81e+06u
M1002 a_294_57# B1 VGND VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=2.352e+11p ps=2.8e+06u
M1003 a_43_57# B1 a_294_57# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VGND C1 a_452_57# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1005 a_358_409# B1 a_29_409# VPB phighvt w=1e+06u l=250000u
+  ad=2.8e+11p pd=2.56e+06u as=0p ps=0u
M1006 X a_43_57# VPWR VPB phighvt w=1e+06u l=250000u
+  ad=2.85e+11p pd=2.57e+06u as=0p ps=0u
M1007 a_452_57# C1 a_43_57# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_610_57# a_43_57# VGND VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1009 a_29_409# A2 VPWR VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1010 X a_43_57# a_610_57# VNB nshort w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=0p ps=0u
M1011 a_43_57# C1 a_358_409# VPB phighvt w=1e+06u l=250000u
+  ad=2.85e+11p pd=2.57e+06u as=0p ps=0u
M1012 VGND A2 a_130_57# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
