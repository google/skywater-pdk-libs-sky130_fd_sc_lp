* File: sky130_fd_sc_lp__and3b_4.spice
* Created: Fri Aug 28 10:06:52 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__and3b_4.pex.spice"
.subckt sky130_fd_sc_lp__and3b_4  VNB VPB A_N C B VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* B	B
* C	C
* A_N	A_N
* VPB	VPB
* VNB	VNB
MM1015 N_VGND_M1015_d N_A_N_M1015_g N_A_49_133#_M1015_s VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.1197 PD=0.913333 PS=1.41 NRD=72.852 NRS=5.712 M=1 R=2.8
+ SA=75000.2 SB=75003.6 A=0.063 P=1.14 MULT=1
MM1002 N_X_M1002_d N_A_242_23#_M1002_g N_VGND_M1015_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2226 PD=1.12 PS=1.82667 NRD=0 NRS=0 M=1 R=5.6 SA=75000.5
+ SB=75003 A=0.126 P=1.98 MULT=1
MM1003 N_X_M1002_d N_A_242_23#_M1003_g N_VGND_M1003_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001 SB=75002.5
+ A=0.126 P=1.98 MULT=1
MM1008 N_X_M1008_d N_A_242_23#_M1008_g N_VGND_M1003_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.4
+ SB=75002.1 A=0.126 P=1.98 MULT=1
MM1012 N_X_M1008_d N_A_242_23#_M1012_g N_VGND_M1012_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1785 PD=1.12 PS=1.265 NRD=0 NRS=9.996 M=1 R=5.6 SA=75001.8
+ SB=75001.7 A=0.126 P=1.98 MULT=1
MM1011 A_645_49# N_C_M1011_g N_VGND_M1012_s VNB NSHORT L=0.15 W=0.84 AD=0.0882
+ AS=0.1785 PD=1.05 PS=1.265 NRD=7.14 NRS=10.704 M=1 R=5.6 SA=75002.4 SB=75001.1
+ A=0.126 P=1.98 MULT=1
MM1004 A_717_49# N_B_M1004_g A_645_49# VNB NSHORT L=0.15 W=0.84 AD=0.1638
+ AS=0.0882 PD=1.23 PS=1.05 NRD=19.992 NRS=7.14 M=1 R=5.6 SA=75002.8 SB=75000.7
+ A=0.126 P=1.98 MULT=1
MM1010 N_A_242_23#_M1010_d N_A_49_133#_M1010_g A_717_49# VNB NSHORT L=0.15
+ W=0.84 AD=0.2226 AS=0.1638 PD=2.21 PS=1.23 NRD=0 NRS=19.992 M=1 R=5.6
+ SA=75003.3 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1009 N_VPWR_M1009_d N_A_N_M1009_g N_A_49_133#_M1009_s VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1113 AS=0.1197 PD=0.895 PS=1.41 NRD=98.5 NRS=9.3772 M=1 R=2.8
+ SA=75000.2 SB=75003.7 A=0.063 P=1.14 MULT=1
MM1000 N_X_M1000_d N_A_242_23#_M1000_g N_VPWR_M1009_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.3339 PD=1.54 PS=2.685 NRD=0 NRS=0 M=1 R=8.4 SA=75000.4 SB=75003
+ A=0.189 P=2.82 MULT=1
MM1006 N_X_M1000_d N_A_242_23#_M1006_g N_VPWR_M1006_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.9
+ SB=75002.6 A=0.189 P=2.82 MULT=1
MM1013 N_X_M1013_d N_A_242_23#_M1013_g N_VPWR_M1006_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.3
+ SB=75002.1 A=0.189 P=2.82 MULT=1
MM1014 N_X_M1013_d N_A_242_23#_M1014_g N_VPWR_M1014_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.22365 PD=1.54 PS=1.615 NRD=0 NRS=0 M=1 R=8.4 SA=75001.7
+ SB=75001.7 A=0.189 P=2.82 MULT=1
MM1001 N_A_242_23#_M1001_d N_C_M1001_g N_VPWR_M1014_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.22365 PD=1.54 PS=1.615 NRD=0 NRS=11.7215 M=1 R=8.4 SA=75002.2
+ SB=75001.2 A=0.189 P=2.82 MULT=1
MM1005 N_VPWR_M1005_d N_B_M1005_g N_A_242_23#_M1001_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.26775 AS=0.1764 PD=1.685 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.6
+ SB=75000.8 A=0.189 P=2.82 MULT=1
MM1007 N_A_242_23#_M1007_d N_A_49_133#_M1007_g N_VPWR_M1005_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.26775 PD=3.05 PS=1.685 NRD=0 NRS=22.655 M=1 R=8.4
+ SA=75003.2 SB=75000.2 A=0.189 P=2.82 MULT=1
DX16_noxref VNB VPB NWDIODE A=9.6607 P=14.09
*
.include "sky130_fd_sc_lp__and3b_4.pxi.spice"
*
.ends
*
*
