* File: sky130_fd_sc_lp__a21bo_0.pxi.spice
* Created: Fri Aug 28 09:49:02 2020
* 
x_PM_SKY130_FD_SC_LP__A21BO_0%A_72_212# N_A_72_212#_M1004_d N_A_72_212#_M1001_s
+ N_A_72_212#_M1002_g N_A_72_212#_M1007_g N_A_72_212#_c_82_n N_A_72_212#_c_83_n
+ N_A_72_212#_c_84_n N_A_72_212#_c_85_n N_A_72_212#_c_86_n N_A_72_212#_c_92_n
+ N_A_72_212#_c_93_n N_A_72_212#_c_87_n N_A_72_212#_c_88_n N_A_72_212#_c_110_p
+ PM_SKY130_FD_SC_LP__A21BO_0%A_72_212#
x_PM_SKY130_FD_SC_LP__A21BO_0%B1_N N_B1_N_M1005_g N_B1_N_M1008_g N_B1_N_c_168_n
+ N_B1_N_c_169_n N_B1_N_c_170_n B1_N B1_N N_B1_N_c_172_n
+ PM_SKY130_FD_SC_LP__A21BO_0%B1_N
x_PM_SKY130_FD_SC_LP__A21BO_0%A_216_526# N_A_216_526#_M1008_d
+ N_A_216_526#_M1005_d N_A_216_526#_c_212_n N_A_216_526#_c_213_n
+ N_A_216_526#_c_214_n N_A_216_526#_M1004_g N_A_216_526#_c_215_n
+ N_A_216_526#_M1001_g N_A_216_526#_c_216_n N_A_216_526#_c_217_n
+ N_A_216_526#_c_224_n N_A_216_526#_c_225_n N_A_216_526#_c_218_n
+ N_A_216_526#_c_226_n N_A_216_526#_c_227_n N_A_216_526#_c_247_n
+ N_A_216_526#_c_219_n N_A_216_526#_c_220_n N_A_216_526#_c_221_n
+ PM_SKY130_FD_SC_LP__A21BO_0%A_216_526#
x_PM_SKY130_FD_SC_LP__A21BO_0%A1 N_A1_M1009_g N_A1_M1006_g N_A1_c_295_n
+ N_A1_c_296_n A1 A1 A1 N_A1_c_298_n PM_SKY130_FD_SC_LP__A21BO_0%A1
x_PM_SKY130_FD_SC_LP__A21BO_0%A2 N_A2_M1000_g N_A2_M1003_g N_A2_c_342_n
+ N_A2_c_343_n A2 A2 A2 N_A2_c_345_n PM_SKY130_FD_SC_LP__A21BO_0%A2
x_PM_SKY130_FD_SC_LP__A21BO_0%X N_X_M1007_s N_X_M1002_s N_X_c_372_n X X X X
+ PM_SKY130_FD_SC_LP__A21BO_0%X
x_PM_SKY130_FD_SC_LP__A21BO_0%VPWR N_VPWR_M1002_d N_VPWR_M1006_d N_VPWR_c_393_n
+ N_VPWR_c_394_n N_VPWR_c_395_n N_VPWR_c_396_n VPWR N_VPWR_c_397_n
+ N_VPWR_c_398_n N_VPWR_c_392_n N_VPWR_c_400_n PM_SKY130_FD_SC_LP__A21BO_0%VPWR
x_PM_SKY130_FD_SC_LP__A21BO_0%A_467_458# N_A_467_458#_M1001_d
+ N_A_467_458#_M1003_d N_A_467_458#_c_433_n N_A_467_458#_c_434_n
+ N_A_467_458#_c_435_n N_A_467_458#_c_436_n
+ PM_SKY130_FD_SC_LP__A21BO_0%A_467_458#
x_PM_SKY130_FD_SC_LP__A21BO_0%VGND N_VGND_M1007_d N_VGND_M1004_s N_VGND_M1000_d
+ N_VGND_c_459_n N_VGND_c_460_n N_VGND_c_461_n N_VGND_c_462_n N_VGND_c_463_n
+ N_VGND_c_464_n N_VGND_c_465_n VGND N_VGND_c_466_n N_VGND_c_467_n
+ N_VGND_c_468_n PM_SKY130_FD_SC_LP__A21BO_0%VGND
cc_1 VNB N_A_72_212#_M1007_g 0.0355703f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=0.47
cc_2 VNB N_A_72_212#_c_82_n 0.0235993f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.565
cc_3 VNB N_A_72_212#_c_83_n 0.00629928f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.73
cc_4 VNB N_A_72_212#_c_84_n 0.0057224f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.225
cc_5 VNB N_A_72_212#_c_85_n 0.0168779f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.225
cc_6 VNB N_A_72_212#_c_86_n 0.0187029f $X=-0.19 $Y=-0.245 $X2=1.88 $Y2=1.645
cc_7 VNB N_A_72_212#_c_87_n 0.00592257f $X=-0.19 $Y=-0.245 $X2=2.29 $Y2=1.56
cc_8 VNB N_A_72_212#_c_88_n 0.0066146f $X=-0.19 $Y=-0.245 $X2=2.29 $Y2=1.645
cc_9 VNB N_B1_N_M1005_g 0.0100234f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_B1_N_c_168_n 0.0202798f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=2.73
cc_11 VNB N_B1_N_c_169_n 0.0218043f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_B1_N_c_170_n 0.0156144f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=1.06
cc_13 VNB B1_N 0.00472648f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=0.47
cc_14 VNB N_B1_N_c_172_n 0.0158912f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.565
cc_15 VNB N_A_216_526#_c_212_n 0.0135561f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=2.73
cc_16 VNB N_A_216_526#_c_213_n 0.0194911f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_216_526#_c_214_n 0.0193229f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=1.06
cc_18 VNB N_A_216_526#_c_215_n 0.0329823f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.225
cc_19 VNB N_A_216_526#_c_216_n 0.0159487f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.225
cc_20 VNB N_A_216_526#_c_217_n 0.00421024f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_216_526#_c_218_n 0.0119833f $X=-0.19 $Y=-0.245 $X2=2.025 $Y2=1.645
cc_22 VNB N_A_216_526#_c_219_n 0.0244154f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_216_526#_c_220_n 0.00338374f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_216_526#_c_221_n 0.0112443f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A1_M1009_g 0.0203513f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A1_M1006_g 0.00664365f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=1.73
cc_27 VNB N_A1_c_295_n 0.0238502f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=1.06
cc_28 VNB N_A1_c_296_n 0.016991f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=0.47
cc_29 VNB A1 0.00462168f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=0.47
cc_30 VNB N_A1_c_298_n 0.0168496f $X=-0.19 $Y=-0.245 $X2=0.562 $Y2=1.225
cc_31 VNB N_A2_M1000_g 0.0258556f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A2_M1003_g 0.00832693f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=1.73
cc_33 VNB N_A2_c_342_n 0.0330084f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=1.06
cc_34 VNB N_A2_c_343_n 0.0212229f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=0.47
cc_35 VNB A2 0.0152232f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=0.47
cc_36 VNB N_A2_c_345_n 0.0212229f $X=-0.19 $Y=-0.245 $X2=0.562 $Y2=1.225
cc_37 VNB N_X_c_372_n 0.0174598f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=1.06
cc_38 VNB X 0.049522f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=0.47
cc_39 VNB N_VPWR_c_392_n 0.163682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_459_n 0.00594222f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_460_n 0.00592691f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.73
cc_42 VNB N_VGND_c_461_n 0.0200862f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.225
cc_43 VNB N_VGND_c_462_n 0.0234554f $X=-0.19 $Y=-0.245 $X2=0.695 $Y2=1.645
cc_44 VNB N_VGND_c_463_n 0.00372602f $X=-0.19 $Y=-0.245 $X2=2.025 $Y2=1.73
cc_45 VNB N_VGND_c_464_n 0.0323153f $X=-0.19 $Y=-0.245 $X2=2.045 $Y2=2.435
cc_46 VNB N_VGND_c_465_n 0.0052999f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_466_n 0.0129628f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_467_n 0.241707f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_468_n 0.0255686f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VPB N_A_72_212#_M1002_g 0.0582293f $X=-0.19 $Y=1.655 $X2=0.48 $Y2=2.73
cc_51 VPB N_A_72_212#_c_83_n 0.0103073f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=1.73
cc_52 VPB N_A_72_212#_c_86_n 0.0161409f $X=-0.19 $Y=1.655 $X2=1.88 $Y2=1.645
cc_53 VPB N_A_72_212#_c_92_n 0.00317908f $X=-0.19 $Y=1.655 $X2=0.695 $Y2=1.645
cc_54 VPB N_A_72_212#_c_93_n 0.0242003f $X=-0.19 $Y=1.655 $X2=2.045 $Y2=2.435
cc_55 VPB N_A_72_212#_c_88_n 0.00253518f $X=-0.19 $Y=1.655 $X2=2.29 $Y2=1.645
cc_56 VPB N_B1_N_M1005_g 0.0724155f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_57 VPB N_A_216_526#_c_215_n 0.00493101f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=1.225
cc_58 VPB N_A_216_526#_M1001_g 0.0371345f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=1.73
cc_59 VPB N_A_216_526#_c_224_n 0.0154509f $X=-0.19 $Y=1.655 $X2=2.025 $Y2=1.73
cc_60 VPB N_A_216_526#_c_225_n 0.0166466f $X=-0.19 $Y=1.655 $X2=2.29 $Y2=0.635
cc_61 VPB N_A_216_526#_c_226_n 0.00462017f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_62 VPB N_A_216_526#_c_227_n 0.0430854f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_63 VPB N_A_216_526#_c_221_n 0.010149f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_64 VPB N_A1_M1006_g 0.0424963f $X=-0.19 $Y=1.655 $X2=0.48 $Y2=1.73
cc_65 VPB A1 0.00225151f $X=-0.19 $Y=1.655 $X2=0.615 $Y2=0.47
cc_66 VPB N_A2_M1003_g 0.0548872f $X=-0.19 $Y=1.655 $X2=0.48 $Y2=1.73
cc_67 VPB A2 0.00711146f $X=-0.19 $Y=1.655 $X2=0.615 $Y2=0.47
cc_68 VPB X 0.0659299f $X=-0.19 $Y=1.655 $X2=0.615 $Y2=0.47
cc_69 VPB N_VPWR_c_393_n 0.0133765f $X=-0.19 $Y=1.655 $X2=0.48 $Y2=2.73
cc_70 VPB N_VPWR_c_394_n 0.0140579f $X=-0.19 $Y=1.655 $X2=0.615 $Y2=0.47
cc_71 VPB N_VPWR_c_395_n 0.0532353f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=1.06
cc_72 VPB N_VPWR_c_396_n 0.00507132f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=1.565
cc_73 VPB N_VPWR_c_397_n 0.0179217f $X=-0.19 $Y=1.655 $X2=0.562 $Y2=1.225
cc_74 VPB N_VPWR_c_398_n 0.0256438f $X=-0.19 $Y=1.655 $X2=2.29 $Y2=1.645
cc_75 VPB N_VPWR_c_392_n 0.100381f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_76 VPB N_VPWR_c_400_n 0.00564836f $X=-0.19 $Y=1.655 $X2=2.375 $Y2=0.47
cc_77 VPB N_A_467_458#_c_433_n 0.00588286f $X=-0.19 $Y=1.655 $X2=0.48 $Y2=2.73
cc_78 VPB N_A_467_458#_c_434_n 0.024605f $X=-0.19 $Y=1.655 $X2=0.615 $Y2=1.06
cc_79 VPB N_A_467_458#_c_435_n 0.00734383f $X=-0.19 $Y=1.655 $X2=0.615 $Y2=0.47
cc_80 VPB N_A_467_458#_c_436_n 0.0370539f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=1.225
cc_81 N_A_72_212#_M1002_g N_B1_N_M1005_g 0.0282084f $X=0.48 $Y=2.73 $X2=0 $Y2=0
cc_82 N_A_72_212#_c_83_n N_B1_N_M1005_g 0.0125353f $X=0.525 $Y=1.73 $X2=0 $Y2=0
cc_83 N_A_72_212#_c_86_n N_B1_N_M1005_g 0.0146286f $X=1.88 $Y=1.645 $X2=0 $Y2=0
cc_84 N_A_72_212#_M1007_g N_B1_N_c_168_n 0.0131561f $X=0.615 $Y=0.47 $X2=0 $Y2=0
cc_85 N_A_72_212#_c_84_n N_B1_N_c_169_n 0.00545465f $X=0.525 $Y=1.225 $X2=0
+ $Y2=0
cc_86 N_A_72_212#_c_85_n N_B1_N_c_169_n 0.0125353f $X=0.525 $Y=1.225 $X2=0 $Y2=0
cc_87 N_A_72_212#_c_82_n N_B1_N_c_170_n 0.0125353f $X=0.525 $Y=1.565 $X2=0 $Y2=0
cc_88 N_A_72_212#_c_86_n N_B1_N_c_170_n 0.00508709f $X=1.88 $Y=1.645 $X2=0 $Y2=0
cc_89 N_A_72_212#_M1007_g B1_N 9.31759e-19 $X=0.615 $Y=0.47 $X2=0 $Y2=0
cc_90 N_A_72_212#_c_84_n B1_N 0.0204107f $X=0.525 $Y=1.225 $X2=0 $Y2=0
cc_91 N_A_72_212#_c_85_n B1_N 4.16558e-19 $X=0.525 $Y=1.225 $X2=0 $Y2=0
cc_92 N_A_72_212#_c_86_n B1_N 0.0310654f $X=1.88 $Y=1.645 $X2=0 $Y2=0
cc_93 N_A_72_212#_M1007_g N_B1_N_c_172_n 0.0125353f $X=0.615 $Y=0.47 $X2=0 $Y2=0
cc_94 N_A_72_212#_c_88_n N_A_216_526#_c_212_n 0.00161104f $X=2.29 $Y=1.645 $X2=0
+ $Y2=0
cc_95 N_A_72_212#_c_87_n N_A_216_526#_c_214_n 0.00414077f $X=2.29 $Y=1.56 $X2=0
+ $Y2=0
cc_96 N_A_72_212#_c_110_p N_A_216_526#_c_214_n 0.00400798f $X=2.375 $Y=0.47
+ $X2=0 $Y2=0
cc_97 N_A_72_212#_c_93_n N_A_216_526#_c_215_n 8.49296e-19 $X=2.045 $Y=2.435
+ $X2=0 $Y2=0
cc_98 N_A_72_212#_c_87_n N_A_216_526#_c_215_n 0.0139769f $X=2.29 $Y=1.56 $X2=0
+ $Y2=0
cc_99 N_A_72_212#_c_88_n N_A_216_526#_c_215_n 0.0152582f $X=2.29 $Y=1.645 $X2=0
+ $Y2=0
cc_100 N_A_72_212#_c_93_n N_A_216_526#_M1001_g 0.00678366f $X=2.045 $Y=2.435
+ $X2=0 $Y2=0
cc_101 N_A_72_212#_c_86_n N_A_216_526#_c_216_n 0.00511067f $X=1.88 $Y=1.645
+ $X2=0 $Y2=0
cc_102 N_A_72_212#_c_87_n N_A_216_526#_c_217_n 0.00491673f $X=2.29 $Y=1.56 $X2=0
+ $Y2=0
cc_103 N_A_72_212#_c_93_n N_A_216_526#_c_224_n 0.00754027f $X=2.045 $Y=2.435
+ $X2=0 $Y2=0
cc_104 N_A_72_212#_c_88_n N_A_216_526#_c_224_n 0.00489055f $X=2.29 $Y=1.645
+ $X2=0 $Y2=0
cc_105 N_A_72_212#_M1002_g N_A_216_526#_c_225_n 8.80087e-19 $X=0.48 $Y=2.73
+ $X2=0 $Y2=0
cc_106 N_A_72_212#_c_93_n N_A_216_526#_c_225_n 0.0307105f $X=2.045 $Y=2.435
+ $X2=0 $Y2=0
cc_107 N_A_72_212#_M1002_g N_A_216_526#_c_226_n 8.75936e-19 $X=0.48 $Y=2.73
+ $X2=0 $Y2=0
cc_108 N_A_72_212#_c_86_n N_A_216_526#_c_226_n 0.0442204f $X=1.88 $Y=1.645 $X2=0
+ $Y2=0
cc_109 N_A_72_212#_c_93_n N_A_216_526#_c_226_n 0.0169026f $X=2.045 $Y=2.435
+ $X2=0 $Y2=0
cc_110 N_A_72_212#_c_86_n N_A_216_526#_c_227_n 0.00438376f $X=1.88 $Y=1.645
+ $X2=0 $Y2=0
cc_111 N_A_72_212#_c_93_n N_A_216_526#_c_227_n 0.00109062f $X=2.045 $Y=2.435
+ $X2=0 $Y2=0
cc_112 N_A_72_212#_c_86_n N_A_216_526#_c_247_n 0.0242594f $X=1.88 $Y=1.645 $X2=0
+ $Y2=0
cc_113 N_A_72_212#_c_87_n N_A_216_526#_c_247_n 0.0192035f $X=2.29 $Y=1.56 $X2=0
+ $Y2=0
cc_114 N_A_72_212#_c_87_n N_A_216_526#_c_219_n 0.00181323f $X=2.29 $Y=1.56 $X2=0
+ $Y2=0
cc_115 N_A_72_212#_c_87_n N_A_216_526#_c_220_n 0.00676077f $X=2.29 $Y=1.56 $X2=0
+ $Y2=0
cc_116 N_A_72_212#_c_86_n N_A_216_526#_c_221_n 0.0119634f $X=1.88 $Y=1.645 $X2=0
+ $Y2=0
cc_117 N_A_72_212#_c_93_n N_A_216_526#_c_221_n 0.00394943f $X=2.045 $Y=2.435
+ $X2=0 $Y2=0
cc_118 N_A_72_212#_c_87_n N_A_216_526#_c_221_n 4.57466e-19 $X=2.29 $Y=1.56 $X2=0
+ $Y2=0
cc_119 N_A_72_212#_c_87_n N_A1_M1009_g 0.00374311f $X=2.29 $Y=1.56 $X2=0 $Y2=0
cc_120 N_A_72_212#_c_110_p N_A1_M1009_g 0.00782453f $X=2.375 $Y=0.47 $X2=0 $Y2=0
cc_121 N_A_72_212#_c_93_n N_A1_M1006_g 6.83691e-19 $X=2.045 $Y=2.435 $X2=0 $Y2=0
cc_122 N_A_72_212#_c_88_n N_A1_M1006_g 6.11626e-19 $X=2.29 $Y=1.645 $X2=0 $Y2=0
cc_123 N_A_72_212#_c_93_n A1 0.00104416f $X=2.045 $Y=2.435 $X2=0 $Y2=0
cc_124 N_A_72_212#_c_87_n A1 0.0556488f $X=2.29 $Y=1.56 $X2=0 $Y2=0
cc_125 N_A_72_212#_c_88_n A1 0.0145695f $X=2.29 $Y=1.645 $X2=0 $Y2=0
cc_126 N_A_72_212#_c_87_n N_A1_c_298_n 0.00436826f $X=2.29 $Y=1.56 $X2=0 $Y2=0
cc_127 N_A_72_212#_c_110_p N_A2_M1000_g 0.00101943f $X=2.375 $Y=0.47 $X2=0 $Y2=0
cc_128 N_A_72_212#_c_84_n N_X_c_372_n 0.00314251f $X=0.525 $Y=1.225 $X2=0 $Y2=0
cc_129 N_A_72_212#_c_85_n N_X_c_372_n 0.00284789f $X=0.525 $Y=1.225 $X2=0 $Y2=0
cc_130 N_A_72_212#_M1002_g X 0.0328782f $X=0.48 $Y=2.73 $X2=0 $Y2=0
cc_131 N_A_72_212#_M1007_g X 0.010269f $X=0.615 $Y=0.47 $X2=0 $Y2=0
cc_132 N_A_72_212#_c_83_n X 0.00204649f $X=0.525 $Y=1.73 $X2=0 $Y2=0
cc_133 N_A_72_212#_c_84_n X 0.0368823f $X=0.525 $Y=1.225 $X2=0 $Y2=0
cc_134 N_A_72_212#_c_85_n X 0.0162713f $X=0.525 $Y=1.225 $X2=0 $Y2=0
cc_135 N_A_72_212#_c_92_n X 0.0135424f $X=0.695 $Y=1.645 $X2=0 $Y2=0
cc_136 N_A_72_212#_M1002_g N_VPWR_c_393_n 0.00311119f $X=0.48 $Y=2.73 $X2=0
+ $Y2=0
cc_137 N_A_72_212#_c_83_n N_VPWR_c_393_n 5.94709e-19 $X=0.525 $Y=1.73 $X2=0
+ $Y2=0
cc_138 N_A_72_212#_c_86_n N_VPWR_c_393_n 0.00609107f $X=1.88 $Y=1.645 $X2=0
+ $Y2=0
cc_139 N_A_72_212#_c_92_n N_VPWR_c_393_n 0.00326515f $X=0.695 $Y=1.645 $X2=0
+ $Y2=0
cc_140 N_A_72_212#_c_93_n N_VPWR_c_395_n 0.011068f $X=2.045 $Y=2.435 $X2=0 $Y2=0
cc_141 N_A_72_212#_M1002_g N_VPWR_c_397_n 0.00521236f $X=0.48 $Y=2.73 $X2=0
+ $Y2=0
cc_142 N_A_72_212#_M1002_g N_VPWR_c_392_n 0.0106484f $X=0.48 $Y=2.73 $X2=0 $Y2=0
cc_143 N_A_72_212#_c_93_n N_VPWR_c_392_n 0.0103764f $X=2.045 $Y=2.435 $X2=0
+ $Y2=0
cc_144 N_A_72_212#_c_93_n N_A_467_458#_c_433_n 0.0159835f $X=2.045 $Y=2.435
+ $X2=0 $Y2=0
cc_145 N_A_72_212#_c_93_n N_A_467_458#_c_435_n 0.0148899f $X=2.045 $Y=2.435
+ $X2=0 $Y2=0
cc_146 N_A_72_212#_c_88_n N_A_467_458#_c_435_n 0.00263564f $X=2.29 $Y=1.645
+ $X2=0 $Y2=0
cc_147 N_A_72_212#_M1007_g N_VGND_c_459_n 0.00307942f $X=0.615 $Y=0.47 $X2=0
+ $Y2=0
cc_148 N_A_72_212#_c_110_p N_VGND_c_461_n 0.00831198f $X=2.375 $Y=0.47 $X2=0
+ $Y2=0
cc_149 N_A_72_212#_c_110_p N_VGND_c_464_n 0.0140843f $X=2.375 $Y=0.47 $X2=0
+ $Y2=0
cc_150 N_A_72_212#_M1007_g N_VGND_c_467_n 0.0114189f $X=0.615 $Y=0.47 $X2=0
+ $Y2=0
cc_151 N_A_72_212#_c_110_p N_VGND_c_467_n 0.0121447f $X=2.375 $Y=0.47 $X2=0
+ $Y2=0
cc_152 N_A_72_212#_M1007_g N_VGND_c_468_n 0.00560159f $X=0.615 $Y=0.47 $X2=0
+ $Y2=0
cc_153 B1_N N_A_216_526#_c_213_n 0.00369604f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_154 N_B1_N_c_172_n N_A_216_526#_c_213_n 0.0122899f $X=1.095 $Y=0.955 $X2=0
+ $Y2=0
cc_155 N_B1_N_c_170_n N_A_216_526#_c_216_n 0.0122899f $X=1.095 $Y=1.46 $X2=0
+ $Y2=0
cc_156 N_B1_N_M1005_g N_A_216_526#_c_225_n 0.0210684f $X=1.005 $Y=2.84 $X2=0
+ $Y2=0
cc_157 B1_N N_A_216_526#_c_218_n 0.0127284f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_158 N_B1_N_c_172_n N_A_216_526#_c_218_n 0.00350863f $X=1.095 $Y=0.955 $X2=0
+ $Y2=0
cc_159 N_B1_N_M1005_g N_A_216_526#_c_226_n 0.00821217f $X=1.005 $Y=2.84 $X2=0
+ $Y2=0
cc_160 N_B1_N_M1005_g N_A_216_526#_c_227_n 0.0186055f $X=1.005 $Y=2.84 $X2=0
+ $Y2=0
cc_161 N_B1_N_c_169_n N_A_216_526#_c_247_n 2.0199e-19 $X=1.095 $Y=1.295 $X2=0
+ $Y2=0
cc_162 N_B1_N_c_170_n N_A_216_526#_c_247_n 2.0199e-19 $X=1.095 $Y=1.46 $X2=0
+ $Y2=0
cc_163 N_B1_N_c_169_n N_A_216_526#_c_219_n 0.0122899f $X=1.095 $Y=1.295 $X2=0
+ $Y2=0
cc_164 N_B1_N_c_168_n N_A_216_526#_c_220_n 0.00381397f $X=1.095 $Y=0.79 $X2=0
+ $Y2=0
cc_165 B1_N N_A_216_526#_c_220_n 0.0439104f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_166 N_B1_N_c_172_n N_A_216_526#_c_220_n 4.83844e-19 $X=1.095 $Y=0.955 $X2=0
+ $Y2=0
cc_167 N_B1_N_M1005_g N_A_216_526#_c_221_n 0.0113655f $X=1.005 $Y=2.84 $X2=0
+ $Y2=0
cc_168 N_B1_N_M1005_g X 0.00151684f $X=1.005 $Y=2.84 $X2=0 $Y2=0
cc_169 B1_N X 0.00608688f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_170 N_B1_N_M1005_g N_VPWR_c_393_n 0.00559626f $X=1.005 $Y=2.84 $X2=0 $Y2=0
cc_171 N_B1_N_M1005_g N_VPWR_c_395_n 0.00508863f $X=1.005 $Y=2.84 $X2=0 $Y2=0
cc_172 N_B1_N_M1005_g N_VPWR_c_392_n 0.0105749f $X=1.005 $Y=2.84 $X2=0 $Y2=0
cc_173 N_B1_N_c_168_n N_VGND_c_459_n 0.00307942f $X=1.095 $Y=0.79 $X2=0 $Y2=0
cc_174 N_B1_N_c_168_n N_VGND_c_462_n 0.00560159f $X=1.095 $Y=0.79 $X2=0 $Y2=0
cc_175 N_B1_N_c_168_n N_VGND_c_467_n 0.00717327f $X=1.095 $Y=0.79 $X2=0 $Y2=0
cc_176 B1_N N_VGND_c_467_n 0.00588921f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_177 N_B1_N_c_172_n N_VGND_c_467_n 5.51567e-19 $X=1.095 $Y=0.955 $X2=0 $Y2=0
cc_178 N_A_216_526#_c_214_n N_A1_M1009_g 0.0142203f $X=2.16 $Y=0.79 $X2=0 $Y2=0
cc_179 N_A_216_526#_c_215_n N_A1_M1006_g 0.00708813f $X=2.16 $Y=1.75 $X2=0 $Y2=0
cc_180 N_A_216_526#_c_224_n N_A1_M1006_g 0.0277628f $X=2.26 $Y=1.825 $X2=0 $Y2=0
cc_181 N_A_216_526#_c_215_n N_A1_c_295_n 0.0173838f $X=2.16 $Y=1.75 $X2=0 $Y2=0
cc_182 N_A_216_526#_c_215_n A1 7.26413e-19 $X=2.16 $Y=1.75 $X2=0 $Y2=0
cc_183 N_A_216_526#_c_217_n A1 6.27163e-19 $X=2.16 $Y=0.865 $X2=0 $Y2=0
cc_184 N_A_216_526#_c_217_n N_A1_c_298_n 0.0173838f $X=2.16 $Y=0.865 $X2=0 $Y2=0
cc_185 N_A_216_526#_c_225_n X 0.00601829f $X=1.22 $Y=2.84 $X2=0 $Y2=0
cc_186 N_A_216_526#_c_226_n X 0.00548507f $X=1.485 $Y=1.995 $X2=0 $Y2=0
cc_187 N_A_216_526#_c_225_n N_VPWR_c_393_n 0.0320683f $X=1.22 $Y=2.84 $X2=0
+ $Y2=0
cc_188 N_A_216_526#_M1001_g N_VPWR_c_395_n 0.0055601f $X=2.26 $Y=2.61 $X2=0
+ $Y2=0
cc_189 N_A_216_526#_c_225_n N_VPWR_c_395_n 0.0145217f $X=1.22 $Y=2.84 $X2=0
+ $Y2=0
cc_190 N_A_216_526#_M1001_g N_VPWR_c_392_n 0.00536257f $X=2.26 $Y=2.61 $X2=0
+ $Y2=0
cc_191 N_A_216_526#_c_225_n N_VPWR_c_392_n 0.012167f $X=1.22 $Y=2.84 $X2=0 $Y2=0
cc_192 N_A_216_526#_M1001_g N_A_467_458#_c_433_n 0.00160705f $X=2.26 $Y=2.61
+ $X2=0 $Y2=0
cc_193 N_A_216_526#_M1001_g N_A_467_458#_c_435_n 0.00152707f $X=2.26 $Y=2.61
+ $X2=0 $Y2=0
cc_194 N_A_216_526#_c_212_n N_VGND_c_460_n 0.00878893f $X=2.085 $Y=0.865 $X2=0
+ $Y2=0
cc_195 N_A_216_526#_c_214_n N_VGND_c_460_n 0.00474713f $X=2.16 $Y=0.79 $X2=0
+ $Y2=0
cc_196 N_A_216_526#_c_218_n N_VGND_c_460_n 0.0271814f $X=1.5 $Y=0.47 $X2=0 $Y2=0
cc_197 N_A_216_526#_c_218_n N_VGND_c_462_n 0.0270056f $X=1.5 $Y=0.47 $X2=0 $Y2=0
cc_198 N_A_216_526#_c_214_n N_VGND_c_464_n 0.00518341f $X=2.16 $Y=0.79 $X2=0
+ $Y2=0
cc_199 N_A_216_526#_c_213_n N_VGND_c_467_n 0.00579769f $X=1.83 $Y=0.865 $X2=0
+ $Y2=0
cc_200 N_A_216_526#_c_214_n N_VGND_c_467_n 0.0106264f $X=2.16 $Y=0.79 $X2=0
+ $Y2=0
cc_201 N_A_216_526#_c_218_n N_VGND_c_467_n 0.0203441f $X=1.5 $Y=0.47 $X2=0 $Y2=0
cc_202 N_A1_M1009_g N_A2_M1000_g 0.0222955f $X=2.59 $Y=0.47 $X2=0 $Y2=0
cc_203 N_A1_M1006_g N_A2_M1003_g 0.0397663f $X=2.69 $Y=2.61 $X2=0 $Y2=0
cc_204 A1 N_A2_M1003_g 6.7886e-19 $X=2.555 $Y=0.84 $X2=0 $Y2=0
cc_205 N_A1_c_295_n N_A2_c_342_n 0.0117125f $X=2.64 $Y=1.345 $X2=0 $Y2=0
cc_206 N_A1_c_296_n N_A2_c_343_n 0.0117125f $X=2.64 $Y=1.51 $X2=0 $Y2=0
cc_207 N_A1_M1006_g A2 9.50465e-19 $X=2.69 $Y=2.61 $X2=0 $Y2=0
cc_208 A1 A2 0.0760517f $X=2.555 $Y=0.84 $X2=0 $Y2=0
cc_209 N_A1_c_298_n A2 0.00420641f $X=2.64 $Y=1.005 $X2=0 $Y2=0
cc_210 A1 N_A2_c_345_n 7.16165e-19 $X=2.555 $Y=0.84 $X2=0 $Y2=0
cc_211 N_A1_c_298_n N_A2_c_345_n 0.0117125f $X=2.64 $Y=1.005 $X2=0 $Y2=0
cc_212 N_A1_M1006_g N_VPWR_c_394_n 0.00347719f $X=2.69 $Y=2.61 $X2=0 $Y2=0
cc_213 N_A1_M1006_g N_VPWR_c_395_n 0.0055601f $X=2.69 $Y=2.61 $X2=0 $Y2=0
cc_214 N_A1_M1006_g N_VPWR_c_392_n 0.00536257f $X=2.69 $Y=2.61 $X2=0 $Y2=0
cc_215 N_A1_M1006_g N_A_467_458#_c_433_n 0.00272031f $X=2.69 $Y=2.61 $X2=0 $Y2=0
cc_216 N_A1_M1006_g N_A_467_458#_c_434_n 0.0147234f $X=2.69 $Y=2.61 $X2=0 $Y2=0
cc_217 N_A1_c_296_n N_A_467_458#_c_434_n 5.21468e-19 $X=2.64 $Y=1.51 $X2=0 $Y2=0
cc_218 A1 N_A_467_458#_c_434_n 0.0147655f $X=2.555 $Y=0.84 $X2=0 $Y2=0
cc_219 N_A1_c_296_n N_A_467_458#_c_435_n 0.00287065f $X=2.64 $Y=1.51 $X2=0 $Y2=0
cc_220 A1 N_A_467_458#_c_435_n 0.00495584f $X=2.555 $Y=0.84 $X2=0 $Y2=0
cc_221 N_A1_M1009_g N_VGND_c_461_n 0.00208133f $X=2.59 $Y=0.47 $X2=0 $Y2=0
cc_222 N_A1_M1009_g N_VGND_c_464_n 0.00525311f $X=2.59 $Y=0.47 $X2=0 $Y2=0
cc_223 N_A1_M1009_g N_VGND_c_467_n 0.00642393f $X=2.59 $Y=0.47 $X2=0 $Y2=0
cc_224 A1 N_VGND_c_467_n 0.00916158f $X=2.555 $Y=0.84 $X2=0 $Y2=0
cc_225 N_A1_c_298_n N_VGND_c_467_n 2.78168e-19 $X=2.64 $Y=1.005 $X2=0 $Y2=0
cc_226 N_A2_M1003_g N_VPWR_c_394_n 0.00345435f $X=3.12 $Y=2.61 $X2=0 $Y2=0
cc_227 N_A2_M1003_g N_VPWR_c_398_n 0.0055601f $X=3.12 $Y=2.61 $X2=0 $Y2=0
cc_228 N_A2_M1003_g N_VPWR_c_392_n 0.00536257f $X=3.12 $Y=2.61 $X2=0 $Y2=0
cc_229 N_A2_M1003_g N_A_467_458#_c_434_n 0.0164086f $X=3.12 $Y=2.61 $X2=0 $Y2=0
cc_230 N_A2_c_343_n N_A_467_458#_c_434_n 7.97015e-19 $X=3.21 $Y=1.51 $X2=0 $Y2=0
cc_231 A2 N_A_467_458#_c_434_n 0.03474f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_232 N_A2_M1003_g N_A_467_458#_c_436_n 0.00590286f $X=3.12 $Y=2.61 $X2=0 $Y2=0
cc_233 N_A2_M1000_g N_VGND_c_461_n 0.0138046f $X=3.12 $Y=0.47 $X2=0 $Y2=0
cc_234 A2 N_VGND_c_461_n 0.0154125f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_235 N_A2_c_345_n N_VGND_c_461_n 0.00111259f $X=3.21 $Y=1.005 $X2=0 $Y2=0
cc_236 N_A2_M1000_g N_VGND_c_464_n 0.00465098f $X=3.12 $Y=0.47 $X2=0 $Y2=0
cc_237 N_A2_M1000_g N_VGND_c_467_n 0.00463525f $X=3.12 $Y=0.47 $X2=0 $Y2=0
cc_238 A2 N_VGND_c_467_n 0.00812866f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_239 X N_VPWR_c_393_n 0.0255011f $X=0.155 $Y=1.95 $X2=0 $Y2=0
cc_240 X N_VPWR_c_397_n 0.0214273f $X=0.155 $Y=1.95 $X2=0 $Y2=0
cc_241 X N_VPWR_c_392_n 0.0125957f $X=0.155 $Y=1.95 $X2=0 $Y2=0
cc_242 N_X_c_372_n N_VGND_c_467_n 0.016502f $X=0.4 $Y=0.47 $X2=0 $Y2=0
cc_243 N_X_c_372_n N_VGND_c_468_n 0.0213766f $X=0.4 $Y=0.47 $X2=0 $Y2=0
cc_244 N_VPWR_c_394_n N_A_467_458#_c_433_n 0.00144674f $X=2.905 $Y=2.445 $X2=0
+ $Y2=0
cc_245 N_VPWR_c_395_n N_A_467_458#_c_433_n 0.00991508f $X=2.77 $Y=3.33 $X2=0
+ $Y2=0
cc_246 N_VPWR_c_392_n N_A_467_458#_c_433_n 0.00929549f $X=3.6 $Y=3.33 $X2=0
+ $Y2=0
cc_247 N_VPWR_c_394_n N_A_467_458#_c_434_n 0.0213307f $X=2.905 $Y=2.445 $X2=0
+ $Y2=0
cc_248 N_VPWR_c_394_n N_A_467_458#_c_436_n 0.00146069f $X=2.905 $Y=2.445 $X2=0
+ $Y2=0
cc_249 N_VPWR_c_398_n N_A_467_458#_c_436_n 0.0112601f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_250 N_VPWR_c_392_n N_A_467_458#_c_436_n 0.0105565f $X=3.6 $Y=3.33 $X2=0 $Y2=0
