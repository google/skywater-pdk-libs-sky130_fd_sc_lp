* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__o2bb2a_m A1_N A2_N B1 B2 VGND VNB VPB VPWR X
M1000 a_85_187# a_209_535# VPWR VPB phighvt w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=5.565e+11p ps=5.17e+06u
M1001 VPWR a_85_187# X VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1002 VPWR A2_N a_209_535# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.176e+11p ps=1.4e+06u
M1003 a_487_167# a_209_535# a_85_187# VNB nshort w=420000u l=150000u
+  ad=2.289e+11p pd=2.77e+06u as=1.113e+11p ps=1.37e+06u
M1004 VGND B2 a_487_167# VNB nshort w=420000u l=150000u
+  ad=2.52e+11p pd=2.88e+06u as=0p ps=0u
M1005 a_487_167# B1 VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND a_85_187# X VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1007 a_223_47# A1_N VGND VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1008 a_209_535# A2_N a_223_47# VNB nshort w=420000u l=150000u
+  ad=2.172e+11p pd=2.02e+06u as=0p ps=0u
M1009 a_559_535# B2 a_85_187# VPB phighvt w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1010 VPWR B1 a_559_535# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_209_535# A1_N VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
