* File: sky130_fd_sc_lp__dfrtp_4.pex.spice
* Created: Fri Aug 28 10:22:30 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__DFRTP_4%CLK 3 7 12 13 14 15 16 21
r38 21 22 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.385
+ $Y=1.535 $X2=0.385 $Y2=1.535
r39 15 16 11.0754 $w=3.83e-07 $l=3.7e-07 $layer=LI1_cond $X=0.277 $Y=1.665
+ $X2=0.277 $Y2=2.035
r40 15 22 3.89137 $w=3.83e-07 $l=1.3e-07 $layer=LI1_cond $X=0.277 $Y=1.665
+ $X2=0.277 $Y2=1.535
r41 14 22 7.18406 $w=3.83e-07 $l=2.4e-07 $layer=LI1_cond $X=0.277 $Y=1.295
+ $X2=0.277 $Y2=1.535
r42 12 21 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=0.385 $Y=1.89
+ $X2=0.385 $Y2=1.535
r43 12 13 43.5886 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=0.435 $Y=1.89
+ $X2=0.435 $Y2=2.04
r44 10 21 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.385 $Y=1.37
+ $X2=0.385 $Y2=1.535
r45 7 13 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=0.575 $Y=2.63
+ $X2=0.575 $Y2=2.04
r46 3 10 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=0.475 $Y=0.66
+ $X2=0.475 $Y2=1.37
.ends

.subckt PM_SKY130_FD_SC_LP__DFRTP_4%A_27_90# 1 2 9 13 16 20 24 28 31 35 36 37 42
+ 43 45 47 48 49 51 52 53 55 56 57 60 62 66 67 70 71 74 75 76 78 79 80 82 83 89
+ 91 93 94 99 109
c293 66 0 1.34651e-19 $X=6.22 $Y=1.79
c294 62 0 1.44909e-19 $X=6.315 $Y=0.61
c295 49 0 1.11939e-19 $X=1.205 $Y=0.375
c296 43 0 1.55256e-19 $X=0.955 $Y=1.145
c297 16 0 2.0335e-20 $X=3.37 $Y=0.805
c298 9 0 6.36774e-20 $X=1.005 $Y=2.63
r299 94 109 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.26 $Y=0.39
+ $X2=7.26 $Y2=0.555
r300 93 96 7.68295 $w=3.28e-07 $l=2.2e-07 $layer=LI1_cond $X=7.26 $Y=0.39
+ $X2=7.26 $Y2=0.61
r301 93 94 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.26
+ $Y=0.39 $X2=7.26 $Y2=0.39
r302 87 89 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=6.22 $Y=1.33
+ $X2=6.4 $Y2=1.33
r303 83 85 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=4.225 $Y=0.45
+ $X2=4.225 $Y2=0.61
r304 79 103 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.46 $Y=1.4
+ $X2=3.46 $Y2=1.565
r305 79 102 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.46 $Y=1.4
+ $X2=3.46 $Y2=1.235
r306 78 80 9.16686 $w=2.23e-07 $l=1.65e-07 $layer=LI1_cond $X=3.477 $Y=1.4
+ $X2=3.477 $Y2=1.235
r307 78 79 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.46
+ $Y=1.4 $X2=3.46 $Y2=1.4
r308 72 91 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.485 $Y=0.61
+ $X2=6.4 $Y2=0.61
r309 71 96 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.095 $Y=0.61
+ $X2=7.26 $Y2=0.61
r310 71 72 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=7.095 $Y=0.61
+ $X2=6.485 $Y2=0.61
r311 70 89 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.4 $Y=1.245
+ $X2=6.4 $Y2=1.33
r312 69 91 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.4 $Y=0.695 $X2=6.4
+ $Y2=0.61
r313 69 70 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=6.4 $Y=0.695
+ $X2=6.4 $Y2=1.245
r314 67 106 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.22 $Y=1.79
+ $X2=6.22 $Y2=1.955
r315 66 67 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.22
+ $Y=1.79 $X2=6.22 $Y2=1.79
r316 64 87 0.0262452 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=6.22 $Y=1.415
+ $X2=6.22 $Y2=1.33
r317 64 66 21.89 $w=1.88e-07 $l=3.75e-07 $layer=LI1_cond $X=6.22 $Y=1.415
+ $X2=6.22 $Y2=1.79
r318 63 85 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.31 $Y=0.61
+ $X2=4.225 $Y2=0.61
r319 62 91 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.315 $Y=0.61
+ $X2=6.4 $Y2=0.61
r320 62 63 130.807 $w=1.68e-07 $l=2.005e-06 $layer=LI1_cond $X=6.315 $Y=0.61
+ $X2=4.31 $Y2=0.61
r321 61 82 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.59 $Y=0.45
+ $X2=3.505 $Y2=0.45
r322 60 83 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.14 $Y=0.45
+ $X2=4.225 $Y2=0.45
r323 60 61 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=4.14 $Y=0.45
+ $X2=3.59 $Y2=0.45
r324 58 82 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.505 $Y=0.535
+ $X2=3.505 $Y2=0.45
r325 58 80 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=3.505 $Y=0.535
+ $X2=3.505 $Y2=1.235
r326 56 82 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.42 $Y=0.45
+ $X2=3.505 $Y2=0.45
r327 56 57 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=3.42 $Y=0.45 $X2=2.82
+ $Y2=0.45
r328 54 57 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.735 $Y=0.535
+ $X2=2.82 $Y2=0.45
r329 54 55 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=2.735 $Y=0.535
+ $X2=2.735 $Y2=1.085
r330 52 55 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.65 $Y=1.17
+ $X2=2.735 $Y2=1.085
r331 52 53 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=2.65 $Y=1.17
+ $X2=2.065 $Y2=1.17
r332 51 53 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.98 $Y=1.085
+ $X2=2.065 $Y2=1.17
r333 50 51 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=1.98 $Y=0.46
+ $X2=1.98 $Y2=1.085
r334 48 50 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.895 $Y=0.375
+ $X2=1.98 $Y2=0.46
r335 48 49 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.895 $Y=0.375
+ $X2=1.205 $Y2=0.375
r336 47 75 3.10218 $w=3.05e-07 $l=1.72337e-07 $layer=LI1_cond $X=1.12 $Y=0.86
+ $X2=0.985 $Y2=0.945
r337 46 49 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.12 $Y=0.46
+ $X2=1.205 $Y2=0.375
r338 46 47 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=1.12 $Y=0.46 $X2=1.12
+ $Y2=0.86
r339 45 76 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=0.85 $Y=2.3
+ $X2=0.85 $Y2=1.65
r340 43 100 79.8068 $w=6e-07 $l=5.05e-07 $layer=POLY_cond $X=1.09 $Y=1.145
+ $X2=1.09 $Y2=1.65
r341 43 99 49.4885 $w=6e-07 $l=1.65e-07 $layer=POLY_cond $X=1.09 $Y=1.145
+ $X2=1.09 $Y2=0.98
r342 42 43 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.955
+ $Y=1.145 $X2=0.955 $Y2=1.145
r343 40 76 10.2759 $w=4.38e-07 $l=2.2e-07 $layer=LI1_cond $X=0.985 $Y=1.43
+ $X2=0.985 $Y2=1.65
r344 40 42 7.46469 $w=4.38e-07 $l=2.85e-07 $layer=LI1_cond $X=0.985 $Y=1.43
+ $X2=0.985 $Y2=1.145
r345 39 75 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.985 $Y=1.03
+ $X2=0.985 $Y2=0.945
r346 39 42 3.01207 $w=4.38e-07 $l=1.15e-07 $layer=LI1_cond $X=0.985 $Y=1.03
+ $X2=0.985 $Y2=1.145
r347 38 74 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.455 $Y=2.385
+ $X2=0.325 $Y2=2.385
r348 37 45 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.765 $Y=2.385
+ $X2=0.85 $Y2=2.3
r349 37 38 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=0.765 $Y=2.385
+ $X2=0.455 $Y2=2.385
r350 35 75 3.51065 $w=1.7e-07 $l=2.2e-07 $layer=LI1_cond $X=0.765 $Y=0.945
+ $X2=0.985 $Y2=0.945
r351 35 36 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=0.765 $Y=0.945
+ $X2=0.355 $Y2=0.945
r352 29 36 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=0.225 $Y=0.86
+ $X2=0.355 $Y2=0.945
r353 29 31 8.86495 $w=2.58e-07 $l=2e-07 $layer=LI1_cond $X=0.225 $Y=0.86
+ $X2=0.225 $Y2=0.66
r354 28 109 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=7.17 $Y=0.875
+ $X2=7.17 $Y2=0.555
r355 24 106 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=6.2 $Y=2.665
+ $X2=6.2 $Y2=1.955
r356 20 103 676.851 $w=1.5e-07 $l=1.32e-06 $layer=POLY_cond $X=3.37 $Y=2.885
+ $X2=3.37 $Y2=1.565
r357 16 102 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=3.37 $Y=0.805
+ $X2=3.37 $Y2=1.235
r358 13 99 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.315 $Y=0.66
+ $X2=1.315 $Y2=0.98
r359 9 100 502.511 $w=1.5e-07 $l=9.8e-07 $layer=POLY_cond $X=1.005 $Y=2.63
+ $X2=1.005 $Y2=1.65
r360 2 74 300 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_PDIFF $count=2 $X=0.235
+ $Y=2.31 $X2=0.36 $Y2=2.465
r361 1 31 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.45 $X2=0.26 $Y2=0.66
.ends

.subckt PM_SKY130_FD_SC_LP__DFRTP_4%D 5 9 11 12 13 14 15 16
c53 16 0 3.16933e-19 $X=2.64 $Y=1.665
c54 13 0 1.5785e-19 $X=2.455 $Y=2.175
r55 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.53
+ $Y=1.62 $X2=2.53 $Y2=1.62
r56 16 21 3.20933 $w=3.93e-07 $l=1.1e-07 $layer=LI1_cond $X=2.64 $Y=1.652
+ $X2=2.53 $Y2=1.652
r57 15 21 10.795 $w=3.93e-07 $l=3.7e-07 $layer=LI1_cond $X=2.16 $Y=1.652
+ $X2=2.53 $Y2=1.652
r58 14 20 58.5785 $w=3.3e-07 $l=3.35e-07 $layer=POLY_cond $X=2.865 $Y=1.62
+ $X2=2.53 $Y2=1.62
r59 12 13 58.3064 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=2.455 $Y=2.025
+ $X2=2.455 $Y2=2.175
r60 11 20 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=2.515 $Y=1.62
+ $X2=2.53 $Y2=1.62
r61 7 14 32.1775 $w=3.3e-07 $l=1.98997e-07 $layer=POLY_cond $X=2.94 $Y=1.455
+ $X2=2.865 $Y2=1.62
r62 7 9 333.298 $w=1.5e-07 $l=6.5e-07 $layer=POLY_cond $X=2.94 $Y=1.455 $X2=2.94
+ $Y2=0.805
r63 5 13 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=2.47 $Y=2.885
+ $X2=2.47 $Y2=2.175
r64 1 11 32.1775 $w=3.3e-07 $l=1.98997e-07 $layer=POLY_cond $X=2.44 $Y=1.785
+ $X2=2.515 $Y2=1.62
r65 1 12 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=2.44 $Y=1.785
+ $X2=2.44 $Y2=2.025
.ends

.subckt PM_SKY130_FD_SC_LP__DFRTP_4%A_216_462# 1 2 9 13 17 19 20 22 25 31 35 39
+ 40 42 43 44 45 54 55 58 59 68 82
c221 59 0 1.3691e-19 $X=4 $Y=1.31
c222 55 0 7.51852e-20 $X=6.96 $Y=2.035
c223 45 0 1.25615e-19 $X=4.225 $Y=2.035
c224 20 0 2.97539e-19 $X=6.385 $Y=1.235
c225 17 0 6.79976e-20 $X=6.31 $Y=0.625
c226 13 0 2.77228e-19 $X=4.07 $Y=0.805
r227 66 68 30.6007 $w=3.3e-07 $l=1.75e-07 $layer=POLY_cond $X=6.825 $Y=2.03
+ $X2=7 $Y2=2.03
r228 64 66 7.86876 $w=3.3e-07 $l=4.5e-08 $layer=POLY_cond $X=6.78 $Y=2.03
+ $X2=6.825 $Y2=2.03
r229 58 59 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4 $Y=1.31
+ $X2=4 $Y2=1.31
r230 55 68 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7 $Y=2.03
+ $X2=7 $Y2=2.03
r231 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=2.035
+ $X2=6.96 $Y2=2.035
r232 52 59 22.5817 $w=3.68e-07 $l=7.25e-07 $layer=LI1_cond $X=4.02 $Y=2.035
+ $X2=4.02 $Y2=1.31
r233 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=2.035
+ $X2=4.08 $Y2=2.035
r234 48 80 1.24964 $w=4.13e-07 $l=4.5e-08 $layer=LI1_cond $X=1.2 $Y=2.077
+ $X2=1.245 $Y2=2.077
r235 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=2.035
+ $X2=1.2 $Y2=2.035
r236 45 51 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.225 $Y=2.035
+ $X2=4.08 $Y2=2.035
r237 44 54 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.815 $Y=2.035
+ $X2=6.96 $Y2=2.035
r238 44 45 3.20544 $w=1.4e-07 $l=2.59e-06 $layer=MET1_cond $X=6.815 $Y=2.035
+ $X2=4.225 $Y2=2.035
r239 43 47 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.345 $Y=2.035
+ $X2=1.2 $Y2=2.035
r240 42 51 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.935 $Y=2.035
+ $X2=4.08 $Y2=2.035
r241 42 43 3.20544 $w=1.4e-07 $l=2.59e-06 $layer=MET1_cond $X=3.935 $Y=2.035
+ $X2=1.345 $Y2=2.035
r242 40 63 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.92 $Y=2.19
+ $X2=2.92 $Y2=2.355
r243 39 82 66.8227 $w=1.98e-07 $l=1.205e-06 $layer=LI1_cond $X=2.92 $Y=2.185
+ $X2=1.715 $Y2=2.185
r244 39 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.92
+ $Y=2.19 $X2=2.92 $Y2=2.19
r245 33 82 7.68553 $w=4.13e-07 $l=1.65e-07 $layer=LI1_cond $X=1.55 $Y=2.077
+ $X2=1.715 $Y2=2.077
r246 33 80 8.46976 $w=4.13e-07 $l=3.05e-07 $layer=LI1_cond $X=1.55 $Y=2.077
+ $X2=1.245 $Y2=2.077
r247 33 35 39.9863 $w=3.28e-07 $l=1.145e-06 $layer=LI1_cond $X=1.55 $Y=1.87
+ $X2=1.55 $Y2=0.725
r248 29 80 3.04077 $w=2.8e-07 $l=2.08e-07 $layer=LI1_cond $X=1.245 $Y=2.285
+ $X2=1.245 $Y2=2.077
r249 29 31 6.99698 $w=2.78e-07 $l=1.7e-07 $layer=LI1_cond $X=1.245 $Y=2.285
+ $X2=1.245 $Y2=2.455
r250 28 58 43.0552 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4 $Y=1.145 $X2=4
+ $Y2=1.31
r251 23 66 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.825 $Y=2.195
+ $X2=6.825 $Y2=2.03
r252 23 25 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=6.825 $Y=2.195
+ $X2=6.825 $Y2=2.65
r253 22 64 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.78 $Y=1.865
+ $X2=6.78 $Y2=2.03
r254 21 22 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=6.78 $Y=1.31
+ $X2=6.78 $Y2=1.865
r255 19 21 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.705 $Y=1.235
+ $X2=6.78 $Y2=1.31
r256 19 20 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=6.705 $Y=1.235
+ $X2=6.385 $Y2=1.235
r257 15 20 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.31 $Y=1.16
+ $X2=6.385 $Y2=1.235
r258 15 17 274.33 $w=1.5e-07 $l=5.35e-07 $layer=POLY_cond $X=6.31 $Y=1.16
+ $X2=6.31 $Y2=0.625
r259 13 28 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=4.07 $Y=0.805
+ $X2=4.07 $Y2=1.145
r260 9 63 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.9 $Y=2.885 $X2=2.9
+ $Y2=2.355
r261 2 31 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=1.08
+ $Y=2.31 $X2=1.22 $Y2=2.455
r262 1 35 182 $w=1.7e-07 $l=3.45868e-07 $layer=licon1_NDIFF $count=1 $X=1.39
+ $Y=0.45 $X2=1.55 $Y2=0.725
.ends

.subckt PM_SKY130_FD_SC_LP__DFRTP_4%A_731_405# 1 2 9 11 12 15 18 21 22 23 26 28
+ 30 31 38 40 44
c110 30 0 9.31515e-20 $X=4.54 $Y=1.31
c111 26 0 1.80912e-19 $X=5.87 $Y=1.485
c112 9 0 2.98772e-19 $X=3.73 $Y=2.885
r113 41 44 5.09734 $w=2.58e-07 $l=1.15e-07 $layer=LI1_cond $X=5.87 $Y=2.335
+ $X2=5.985 $Y2=2.335
r114 35 38 6.1 $w=1.98e-07 $l=1.1e-07 $layer=LI1_cond $X=5.87 $Y=0.965 $X2=5.98
+ $Y2=0.965
r115 30 33 9.07985 $w=3.28e-07 $l=2.6e-07 $layer=LI1_cond $X=4.54 $Y=1.31
+ $X2=4.54 $Y2=1.57
r116 30 31 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.54
+ $Y=1.31 $X2=4.54 $Y2=1.31
r117 28 41 3.22376 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=5.87 $Y=2.205
+ $X2=5.87 $Y2=2.335
r118 27 40 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.87 $Y=1.655
+ $X2=5.87 $Y2=1.57
r119 27 28 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=5.87 $Y=1.655
+ $X2=5.87 $Y2=2.205
r120 26 40 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.87 $Y=1.485
+ $X2=5.87 $Y2=1.57
r121 25 35 1.68994 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=5.87 $Y=1.065 $X2=5.87
+ $Y2=0.965
r122 25 26 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=5.87 $Y=1.065
+ $X2=5.87 $Y2=1.485
r123 24 33 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.705 $Y=1.57
+ $X2=4.54 $Y2=1.57
r124 23 40 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.785 $Y=1.57
+ $X2=5.87 $Y2=1.57
r125 23 24 70.4599 $w=1.68e-07 $l=1.08e-06 $layer=LI1_cond $X=5.785 $Y=1.57
+ $X2=4.705 $Y2=1.57
r126 21 31 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=4.54 $Y=1.65
+ $X2=4.54 $Y2=1.31
r127 21 22 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.54 $Y=1.65
+ $X2=4.54 $Y2=1.815
r128 20 31 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.54 $Y=1.145
+ $X2=4.54 $Y2=1.31
r129 18 22 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=4.45 $Y=2.025
+ $X2=4.45 $Y2=1.815
r130 15 20 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=4.45 $Y=0.805
+ $X2=4.45 $Y2=1.145
r131 11 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.375 $Y=2.1
+ $X2=4.45 $Y2=2.025
r132 11 12 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=4.375 $Y=2.1
+ $X2=3.805 $Y2=2.1
r133 7 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.73 $Y=2.175
+ $X2=3.805 $Y2=2.1
r134 7 9 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=3.73 $Y=2.175
+ $X2=3.73 $Y2=2.885
r135 2 44 600 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=5.845
+ $Y=2.245 $X2=5.985 $Y2=2.37
r136 1 38 182 $w=1.7e-07 $l=7.72043e-07 $layer=licon1_NDIFF $count=1 $X=5.725
+ $Y=0.305 $X2=5.98 $Y2=0.96
.ends

.subckt PM_SKY130_FD_SC_LP__DFRTP_4%RESET_B 3 5 6 9 11 15 17 18 22 25 29 31 34
+ 35 36 38 41 42 43 45 46 48 52 53 58 64 66
c209 29 0 4.01027e-20 $X=8.41 $Y=0.875
c210 18 0 1.25615e-19 $X=4.31 $Y=2.46
c211 17 0 9.31515e-20 $X=4.735 $Y=2.46
c212 11 0 1.76895e-19 $X=4.915 $Y=0.18
c213 9 0 1.61677e-19 $X=2.58 $Y=0.805
r214 64 66 1.26488 $w=4.08e-07 $l=4.5e-08 $layer=LI1_cond $X=8.36 $Y=1.62
+ $X2=8.36 $Y2=1.665
r215 52 64 2.47908 $w=4.1e-07 $l=8.5e-08 $layer=LI1_cond $X=8.36 $Y=1.535
+ $X2=8.36 $Y2=1.62
r216 52 53 9.83793 $w=4.08e-07 $l=3.5e-07 $layer=LI1_cond $X=8.36 $Y=1.685
+ $X2=8.36 $Y2=2.035
r217 52 66 0.562167 $w=4.08e-07 $l=2e-08 $layer=LI1_cond $X=8.36 $Y=1.685
+ $X2=8.36 $Y2=1.665
r218 52 58 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=8.32
+ $Y=1.615 $X2=8.32 $Y2=1.615
r219 48 50 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=5.87 $Y=2.72
+ $X2=5.87 $Y2=2.87
r220 46 62 19.2347 $w=3.3e-07 $l=1.1e-07 $layer=POLY_cond $X=4.9 $Y=2.35 $X2=4.9
+ $Y2=2.46
r221 46 61 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.9 $Y=2.35
+ $X2=4.9 $Y2=2.185
r222 45 47 18.2753 $w=2.47e-07 $l=3.7e-07 $layer=LI1_cond $X=4.9 $Y=2.35 $X2=4.9
+ $Y2=2.72
r223 45 46 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.9
+ $Y=2.35 $X2=4.9 $Y2=2.35
r224 42 52 5.97895 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=8.155 $Y=1.535
+ $X2=8.36 $Y2=1.535
r225 42 43 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=8.155 $Y=1.535
+ $X2=7.515 $Y2=1.535
r226 40 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.43 $Y=1.62
+ $X2=7.515 $Y2=1.535
r227 40 41 76.0053 $w=1.68e-07 $l=1.165e-06 $layer=LI1_cond $X=7.43 $Y=1.62
+ $X2=7.43 $Y2=2.785
r228 39 50 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.955 $Y=2.87
+ $X2=5.87 $Y2=2.87
r229 38 41 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.345 $Y=2.87
+ $X2=7.43 $Y2=2.785
r230 38 39 90.6845 $w=1.68e-07 $l=1.39e-06 $layer=LI1_cond $X=7.345 $Y=2.87
+ $X2=5.955 $Y2=2.87
r231 37 47 2.92482 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.065 $Y=2.72
+ $X2=4.9 $Y2=2.72
r232 36 48 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.785 $Y=2.72
+ $X2=5.87 $Y2=2.72
r233 36 37 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=5.785 $Y=2.72
+ $X2=5.065 $Y2=2.72
r234 34 58 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=8.32 $Y=1.955
+ $X2=8.32 $Y2=1.615
r235 34 35 37.7798 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.32 $Y=1.955
+ $X2=8.32 $Y2=2.12
r236 33 58 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.32 $Y=1.45
+ $X2=8.32 $Y2=1.615
r237 29 33 294.84 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=8.41 $Y=0.875
+ $X2=8.41 $Y2=1.45
r238 25 35 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=8.315 $Y=2.65
+ $X2=8.315 $Y2=2.12
r239 22 61 743.511 $w=1.5e-07 $l=1.45e-06 $layer=POLY_cond $X=4.99 $Y=0.735
+ $X2=4.99 $Y2=2.185
r240 19 22 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=4.99 $Y=0.255
+ $X2=4.99 $Y2=0.735
r241 17 62 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.735 $Y=2.46
+ $X2=4.9 $Y2=2.46
r242 17 18 217.926 $w=1.5e-07 $l=4.25e-07 $layer=POLY_cond $X=4.735 $Y=2.46
+ $X2=4.31 $Y2=2.46
r243 13 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.235 $Y=2.535
+ $X2=4.31 $Y2=2.46
r244 13 15 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=4.235 $Y=2.535
+ $X2=4.235 $Y2=2.885
r245 12 31 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.655 $Y=0.18
+ $X2=2.58 $Y2=0.18
r246 11 19 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.915 $Y=0.18
+ $X2=4.99 $Y2=0.255
r247 11 12 1158.85 $w=1.5e-07 $l=2.26e-06 $layer=POLY_cond $X=4.915 $Y=0.18
+ $X2=2.655 $Y2=0.18
r248 7 31 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.58 $Y=0.255
+ $X2=2.58 $Y2=0.18
r249 7 9 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=2.58 $Y=0.255
+ $X2=2.58 $Y2=0.805
r250 5 31 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.505 $Y=0.18
+ $X2=2.58 $Y2=0.18
r251 5 6 199.979 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=2.505 $Y=0.18
+ $X2=2.115 $Y2=0.18
r252 1 6 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.04 $Y=0.255
+ $X2=2.115 $Y2=0.18
r253 1 3 1348.57 $w=1.5e-07 $l=2.63e-06 $layer=POLY_cond $X=2.04 $Y=0.255
+ $X2=2.04 $Y2=2.885
.ends

.subckt PM_SKY130_FD_SC_LP__DFRTP_4%A_595_535# 1 2 3 11 12 14 17 19 24 25 26 27
+ 29 31 34 35 36 38 43 50 51 58
c147 51 0 1.80239e-20 $X=5.44 $Y=1.92
c148 43 0 6.79976e-20 $X=5.44 $Y=0.96
c149 38 0 1.26057e-19 $X=3.855 $Y=0.88
c150 27 0 1.76895e-19 $X=5.275 $Y=0.96
r151 51 60 17.0787 $w=2.54e-07 $l=9e-08 $layer=POLY_cond $X=5.44 $Y=1.92
+ $X2=5.35 $Y2=1.92
r152 50 53 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=5.44 $Y=1.92 $X2=5.44
+ $Y2=2
r153 50 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.44
+ $Y=1.92 $X2=5.44 $Y2=1.92
r154 47 58 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=5.44 $Y=1.22
+ $X2=5.65 $Y2=1.22
r155 47 55 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=5.44 $Y=1.22 $X2=5.35
+ $Y2=1.22
r156 46 47 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.44
+ $Y=1.22 $X2=5.44 $Y2=1.22
r157 43 46 9.07985 $w=3.28e-07 $l=2.6e-07 $layer=LI1_cond $X=5.44 $Y=0.96
+ $X2=5.44 $Y2=1.22
r158 38 40 4.43636 $w=1.98e-07 $l=8e-08 $layer=LI1_cond $X=3.86 $Y=0.88 $X2=3.86
+ $Y2=0.96
r159 35 53 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.275 $Y=2 $X2=5.44
+ $Y2=2
r160 35 36 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=5.275 $Y=2
+ $X2=4.545 $Y2=2
r161 34 42 5.3796 $w=2.42e-07 $l=8.89101e-08 $layer=LI1_cond $X=4.46 $Y=2.455
+ $X2=4.452 $Y2=2.54
r162 33 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.46 $Y=2.085
+ $X2=4.545 $Y2=2
r163 33 34 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=4.46 $Y=2.085
+ $X2=4.46 $Y2=2.455
r164 29 42 10.1053 $w=2.65e-07 $l=2.17e-07 $layer=LI1_cond $X=4.452 $Y=2.757
+ $X2=4.452 $Y2=2.54
r165 29 31 5.56652 $w=2.63e-07 $l=1.28e-07 $layer=LI1_cond $X=4.452 $Y=2.757
+ $X2=4.452 $Y2=2.885
r166 28 40 1.68994 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=3.96 $Y=0.96 $X2=3.86
+ $Y2=0.96
r167 27 43 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.275 $Y=0.96
+ $X2=5.44 $Y2=0.96
r168 27 28 85.7914 $w=1.68e-07 $l=1.315e-06 $layer=LI1_cond $X=5.275 $Y=0.96
+ $X2=3.96 $Y2=0.96
r169 25 42 2.80567 $w=1.7e-07 $l=1.32e-07 $layer=LI1_cond $X=4.32 $Y=2.54
+ $X2=4.452 $Y2=2.54
r170 25 26 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=4.32 $Y=2.54
+ $X2=3.765 $Y2=2.54
r171 23 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.68 $Y=2.625
+ $X2=3.765 $Y2=2.54
r172 23 24 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=3.68 $Y=2.625
+ $X2=3.68 $Y2=2.795
r173 19 24 7.36005 $w=2.8e-07 $l=1.77482e-07 $layer=LI1_cond $X=3.595 $Y=2.935
+ $X2=3.68 $Y2=2.795
r174 19 21 18.1098 $w=2.78e-07 $l=4.4e-07 $layer=LI1_cond $X=3.595 $Y=2.935
+ $X2=3.155 $Y2=2.935
r175 15 51 62.622 $w=2.54e-07 $l=4.04166e-07 $layer=POLY_cond $X=5.77 $Y=2.085
+ $X2=5.44 $Y2=1.92
r176 15 17 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=5.77 $Y=2.085
+ $X2=5.77 $Y2=2.665
r177 12 58 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.65 $Y=1.055
+ $X2=5.65 $Y2=1.22
r178 12 14 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=5.65 $Y=1.055
+ $X2=5.65 $Y2=0.625
r179 11 60 15.087 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.35 $Y=1.755
+ $X2=5.35 $Y2=1.92
r180 10 55 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.35 $Y=1.385
+ $X2=5.35 $Y2=1.22
r181 10 11 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=5.35 $Y=1.385
+ $X2=5.35 $Y2=1.755
r182 3 31 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=4.31
+ $Y=2.675 $X2=4.45 $Y2=2.885
r183 2 21 600 $w=1.7e-07 $l=3.1229e-07 $layer=licon1_PDIFF $count=1 $X=2.975
+ $Y=2.675 $X2=3.155 $Y2=2.91
r184 1 38 182 $w=1.7e-07 $l=5.33807e-07 $layer=licon1_NDIFF $count=1 $X=3.445
+ $Y=0.595 $X2=3.855 $Y2=0.88
.ends

.subckt PM_SKY130_FD_SC_LP__DFRTP_4%A_1475_426# 1 2 9 13 17 20 21 24 26 28 33 34
+ 36
c88 36 0 7.51852e-20 $X=7.71 $Y=2.115
c89 33 0 4.01027e-20 $X=9.21 $Y=2.3
c90 13 0 1.3753e-19 $X=7.71 $Y=0.875
r91 32 33 89.3797 $w=1.68e-07 $l=1.37e-06 $layer=LI1_cond $X=9.21 $Y=0.93
+ $X2=9.21 $Y2=2.3
r92 28 32 7.36005 $w=2.8e-07 $l=1.77482e-07 $layer=LI1_cond $X=9.125 $Y=0.79
+ $X2=9.21 $Y2=0.93
r93 28 30 4.93904 $w=2.78e-07 $l=1.2e-07 $layer=LI1_cond $X=9.125 $Y=0.79
+ $X2=9.005 $Y2=0.79
r94 27 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.695 $Y=2.385
+ $X2=8.53 $Y2=2.385
r95 26 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.125 $Y=2.385
+ $X2=9.21 $Y2=2.3
r96 26 27 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=9.125 $Y=2.385
+ $X2=8.695 $Y2=2.385
r97 22 34 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.53 $Y=2.47 $X2=8.53
+ $Y2=2.385
r98 22 24 6.28605 $w=3.28e-07 $l=1.8e-07 $layer=LI1_cond $X=8.53 $Y=2.47
+ $X2=8.53 $Y2=2.65
r99 20 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.365 $Y=2.385
+ $X2=8.53 $Y2=2.385
r100 20 21 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=8.365 $Y=2.385
+ $X2=7.945 $Y2=2.385
r101 18 36 11.9645 $w=2.82e-07 $l=7e-08 $layer=POLY_cond $X=7.78 $Y=2.115
+ $X2=7.71 $Y2=2.115
r102 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.78
+ $Y=2.115 $X2=7.78 $Y2=2.115
r103 15 21 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=7.815 $Y=2.3
+ $X2=7.945 $Y2=2.385
r104 15 17 8.20008 $w=2.58e-07 $l=1.85e-07 $layer=LI1_cond $X=7.815 $Y=2.3
+ $X2=7.815 $Y2=2.115
r105 11 36 17.5183 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.71 $Y=1.95
+ $X2=7.71 $Y2=2.115
r106 11 13 551.223 $w=1.5e-07 $l=1.075e-06 $layer=POLY_cond $X=7.71 $Y=1.95
+ $X2=7.71 $Y2=0.875
r107 7 36 44.4397 $w=2.82e-07 $l=3.32415e-07 $layer=POLY_cond $X=7.45 $Y=2.28
+ $X2=7.71 $Y2=2.115
r108 7 9 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=7.45 $Y=2.28 $X2=7.45
+ $Y2=2.65
r109 2 24 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=8.39
+ $Y=2.44 $X2=8.53 $Y2=2.65
r110 1 30 182 $w=1.7e-07 $l=2.22711e-07 $layer=licon1_NDIFF $count=1 $X=8.845
+ $Y=0.665 $X2=9.005 $Y2=0.815
.ends

.subckt PM_SKY130_FD_SC_LP__DFRTP_4%A_1255_449# 1 2 7 9 12 14 16 18 21 24 26 27
+ 31 32 36 37 40 41 45 48
c119 48 0 1.3753e-19 $X=6.82 $Y=0.96
r120 50 51 5.02519 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=6.82 $Y=1.185
+ $X2=6.82 $Y2=1.27
r121 48 50 7.85757 $w=3.28e-07 $l=2.25e-07 $layer=LI1_cond $X=6.82 $Y=0.96
+ $X2=6.82 $Y2=1.185
r122 43 45 11.6128 $w=1.68e-07 $l=1.78e-07 $layer=LI1_cond $X=6.572 $Y=1.68
+ $X2=6.75 $Y2=1.68
r123 40 41 8.29065 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=6.495 $Y=2.51
+ $X2=6.495 $Y2=2.345
r124 36 37 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=8.86
+ $Y=1.36 $X2=8.86 $Y2=1.36
r125 34 36 4.71454 $w=2.18e-07 $l=9e-08 $layer=LI1_cond $X=8.845 $Y=1.27
+ $X2=8.845 $Y2=1.36
r126 33 50 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.985 $Y=1.185
+ $X2=6.82 $Y2=1.185
r127 32 34 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=8.735 $Y=1.185
+ $X2=8.845 $Y2=1.27
r128 32 33 114.171 $w=1.68e-07 $l=1.75e-06 $layer=LI1_cond $X=8.735 $Y=1.185
+ $X2=6.985 $Y2=1.185
r129 31 45 0.0262452 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=6.75 $Y=1.595
+ $X2=6.75 $Y2=1.68
r130 31 51 18.9713 $w=1.88e-07 $l=3.25e-07 $layer=LI1_cond $X=6.75 $Y=1.595
+ $X2=6.75 $Y2=1.27
r131 28 43 0.574824 $w=1.75e-07 $l=8.5e-08 $layer=LI1_cond $X=6.572 $Y=1.765
+ $X2=6.572 $Y2=1.68
r132 28 41 36.7584 $w=1.73e-07 $l=5.8e-07 $layer=LI1_cond $X=6.572 $Y=1.765
+ $X2=6.572 $Y2=2.345
r133 25 37 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=8.86 $Y=1.7
+ $X2=8.86 $Y2=1.36
r134 25 26 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.86 $Y=1.7
+ $X2=8.86 $Y2=1.865
r135 23 37 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=8.86 $Y=1.345
+ $X2=8.86 $Y2=1.36
r136 23 24 13.5877 $w=2.4e-07 $l=7.5e-08 $layer=POLY_cond $X=8.86 $Y=1.345
+ $X2=8.86 $Y2=1.27
r137 19 27 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.795 $Y=1.345
+ $X2=9.795 $Y2=1.27
r138 19 21 574.298 $w=1.5e-07 $l=1.12e-06 $layer=POLY_cond $X=9.795 $Y=1.345
+ $X2=9.795 $Y2=2.465
r139 16 27 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.795 $Y=1.195
+ $X2=9.795 $Y2=1.27
r140 16 18 173.52 $w=1.5e-07 $l=5.4e-07 $layer=POLY_cond $X=9.795 $Y=1.195
+ $X2=9.795 $Y2=0.655
r141 15 24 12.1617 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.025 $Y=1.27
+ $X2=8.86 $Y2=1.27
r142 14 27 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.72 $Y=1.27
+ $X2=9.795 $Y2=1.27
r143 14 15 356.372 $w=1.5e-07 $l=6.95e-07 $layer=POLY_cond $X=9.72 $Y=1.27
+ $X2=9.025 $Y2=1.27
r144 12 26 402.521 $w=1.5e-07 $l=7.85e-07 $layer=POLY_cond $X=8.77 $Y=2.65
+ $X2=8.77 $Y2=1.865
r145 7 24 13.5877 $w=2.4e-07 $l=1.21861e-07 $layer=POLY_cond $X=8.77 $Y=1.195
+ $X2=8.86 $Y2=1.27
r146 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=8.77 $Y=1.195
+ $X2=8.77 $Y2=0.875
r147 2 40 600 $w=1.7e-07 $l=3.58504e-07 $layer=licon1_PDIFF $count=1 $X=6.275
+ $Y=2.245 $X2=6.495 $Y2=2.51
r148 1 48 182 $w=1.7e-07 $l=8.44956e-07 $layer=licon1_NDIFF $count=1 $X=6.385
+ $Y=0.305 $X2=6.82 $Y2=0.96
.ends

.subckt PM_SKY130_FD_SC_LP__DFRTP_4%A_1891_47# 1 2 9 13 17 21 25 29 33 37 41 45
+ 54 57 64
r99 61 62 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=10.655 $Y=1.49
+ $X2=11.085 $Y2=1.49
r100 55 64 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=11.335 $Y=1.49
+ $X2=11.515 $Y2=1.49
r101 55 62 43.7153 $w=3.3e-07 $l=2.5e-07 $layer=POLY_cond $X=11.335 $Y=1.49
+ $X2=11.085 $Y2=1.49
r102 54 55 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=11.335
+ $Y=1.49 $X2=11.335 $Y2=1.49
r103 52 61 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=10.315 $Y=1.49
+ $X2=10.655 $Y2=1.49
r104 52 58 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=10.315 $Y=1.49
+ $X2=10.225 $Y2=1.49
r105 51 54 62.8485 $w=1.78e-07 $l=1.02e-06 $layer=LI1_cond $X=10.315 $Y=1.495
+ $X2=11.335 $Y2=1.495
r106 51 52 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=10.315
+ $Y=1.49 $X2=10.315 $Y2=1.49
r107 49 57 2.47289 $w=1.8e-07 $l=1.23e-07 $layer=LI1_cond $X=9.71 $Y=1.495
+ $X2=9.587 $Y2=1.495
r108 49 51 37.2778 $w=1.78e-07 $l=6.05e-07 $layer=LI1_cond $X=9.71 $Y=1.495
+ $X2=10.315 $Y2=1.495
r109 45 47 43.7458 $w=2.43e-07 $l=9.3e-07 $layer=LI1_cond $X=9.587 $Y=1.98
+ $X2=9.587 $Y2=2.91
r110 43 57 3.96879 $w=2.45e-07 $l=9e-08 $layer=LI1_cond $X=9.587 $Y=1.585
+ $X2=9.587 $Y2=1.495
r111 43 45 18.5802 $w=2.43e-07 $l=3.95e-07 $layer=LI1_cond $X=9.587 $Y=1.585
+ $X2=9.587 $Y2=1.98
r112 39 57 3.96879 $w=2.45e-07 $l=9e-08 $layer=LI1_cond $X=9.587 $Y=1.405
+ $X2=9.587 $Y2=1.495
r113 39 41 46.3329 $w=2.43e-07 $l=9.85e-07 $layer=LI1_cond $X=9.587 $Y=1.405
+ $X2=9.587 $Y2=0.42
r114 35 64 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=11.515 $Y=1.655
+ $X2=11.515 $Y2=1.49
r115 35 37 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=11.515 $Y=1.655
+ $X2=11.515 $Y2=2.465
r116 31 64 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=11.515 $Y=1.325
+ $X2=11.515 $Y2=1.49
r117 31 33 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=11.515 $Y=1.325
+ $X2=11.515 $Y2=0.655
r118 27 62 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=11.085 $Y=1.655
+ $X2=11.085 $Y2=1.49
r119 27 29 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=11.085 $Y=1.655
+ $X2=11.085 $Y2=2.465
r120 23 62 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=11.085 $Y=1.325
+ $X2=11.085 $Y2=1.49
r121 23 25 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=11.085 $Y=1.325
+ $X2=11.085 $Y2=0.655
r122 19 61 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.655 $Y=1.655
+ $X2=10.655 $Y2=1.49
r123 19 21 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=10.655 $Y=1.655
+ $X2=10.655 $Y2=2.465
r124 15 61 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.655 $Y=1.325
+ $X2=10.655 $Y2=1.49
r125 15 17 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=10.655 $Y=1.325
+ $X2=10.655 $Y2=0.655
r126 11 58 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.225 $Y=1.655
+ $X2=10.225 $Y2=1.49
r127 11 13 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=10.225 $Y=1.655
+ $X2=10.225 $Y2=2.465
r128 7 58 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.225 $Y=1.325
+ $X2=10.225 $Y2=1.49
r129 7 9 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=10.225 $Y=1.325
+ $X2=10.225 $Y2=0.655
r130 2 47 400 $w=1.7e-07 $l=1.13578e-06 $layer=licon1_PDIFF $count=1 $X=9.455
+ $Y=1.835 $X2=9.58 $Y2=2.91
r131 2 45 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=9.455
+ $Y=1.835 $X2=9.58 $Y2=1.98
r132 1 41 91 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=2 $X=9.455
+ $Y=0.235 $X2=9.58 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__DFRTP_4%VPWR 1 2 3 4 5 6 7 8 9 30 34 38 42 44 48 52
+ 58 62 64 69 70 71 73 78 83 91 96 108 112 118 121 124 127 134 137 140 144
r165 143 144 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.76 $Y=3.33
+ $X2=11.76 $Y2=3.33
r166 140 141 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=3.33
+ $X2=10.8 $Y2=3.33
r167 137 138 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r168 135 138 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=8.88 $Y2=3.33
r169 134 135 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r170 130 131 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r171 127 130 9.07985 $w=3.28e-07 $l=2.6e-07 $layer=LI1_cond $X=5.44 $Y=3.07
+ $X2=5.44 $Y2=3.33
r172 124 125 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r173 121 122 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r174 118 119 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r175 116 144 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=3.33
+ $X2=11.76 $Y2=3.33
r176 116 141 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=3.33
+ $X2=10.8 $Y2=3.33
r177 115 116 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.28 $Y=3.33
+ $X2=11.28 $Y2=3.33
r178 113 140 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.035 $Y=3.33
+ $X2=10.87 $Y2=3.33
r179 113 115 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=11.035 $Y=3.33
+ $X2=11.28 $Y2=3.33
r180 112 143 4.76062 $w=1.7e-07 $l=2.17e-07 $layer=LI1_cond $X=11.565 $Y=3.33
+ $X2=11.782 $Y2=3.33
r181 112 115 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=11.565 $Y=3.33
+ $X2=11.28 $Y2=3.33
r182 111 141 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=3.33
+ $X2=10.8 $Y2=3.33
r183 110 111 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.32 $Y=3.33
+ $X2=10.32 $Y2=3.33
r184 108 140 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.705 $Y=3.33
+ $X2=10.87 $Y2=3.33
r185 108 110 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=10.705 $Y=3.33
+ $X2=10.32 $Y2=3.33
r186 107 111 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.84 $Y=3.33
+ $X2=10.32 $Y2=3.33
r187 107 138 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=9.84 $Y=3.33
+ $X2=8.88 $Y2=3.33
r188 106 107 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r189 104 137 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.205 $Y=3.33
+ $X2=9.04 $Y2=3.33
r190 104 106 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=9.205 $Y=3.33
+ $X2=9.84 $Y2=3.33
r191 103 135 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=7.92 $Y2=3.33
r192 102 103 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r193 99 102 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=6 $Y=3.33
+ $X2=7.44 $Y2=3.33
r194 97 130 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.605 $Y=3.33
+ $X2=5.44 $Y2=3.33
r195 97 99 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=5.605 $Y=3.33
+ $X2=6 $Y2=3.33
r196 96 134 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.715 $Y=3.33
+ $X2=7.88 $Y2=3.33
r197 96 102 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=7.715 $Y=3.33
+ $X2=7.44 $Y2=3.33
r198 95 131 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=5.52 $Y2=3.33
r199 95 125 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=4.08 $Y2=3.33
r200 94 95 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r201 92 124 6.25164 $w=1.7e-07 $l=1.08e-07 $layer=LI1_cond $X=4.15 $Y=3.33
+ $X2=4.042 $Y2=3.33
r202 92 94 58.0642 $w=1.68e-07 $l=8.9e-07 $layer=LI1_cond $X=4.15 $Y=3.33
+ $X2=5.04 $Y2=3.33
r203 91 130 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.275 $Y=3.33
+ $X2=5.44 $Y2=3.33
r204 91 94 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=5.275 $Y=3.33
+ $X2=5.04 $Y2=3.33
r205 90 125 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r206 89 90 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r207 87 90 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r208 87 122 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r209 86 89 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.64 $Y=3.33 $X2=3.6
+ $Y2=3.33
r210 86 87 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r211 84 121 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.42 $Y=3.33
+ $X2=2.255 $Y2=3.33
r212 84 86 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=2.42 $Y=3.33
+ $X2=2.64 $Y2=3.33
r213 83 124 6.25164 $w=1.7e-07 $l=1.07e-07 $layer=LI1_cond $X=3.935 $Y=3.33
+ $X2=4.042 $Y2=3.33
r214 83 89 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=3.935 $Y=3.33
+ $X2=3.6 $Y2=3.33
r215 82 122 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r216 82 119 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r217 81 82 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r218 79 118 8.23795 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=0.935 $Y=3.33
+ $X2=0.78 $Y2=3.33
r219 79 81 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.935 $Y=3.33
+ $X2=1.2 $Y2=3.33
r220 78 121 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.09 $Y=3.33
+ $X2=2.255 $Y2=3.33
r221 78 81 58.0642 $w=1.68e-07 $l=8.9e-07 $layer=LI1_cond $X=2.09 $Y=3.33
+ $X2=1.2 $Y2=3.33
r222 76 119 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r223 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r224 73 118 8.23795 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=0.625 $Y=3.33
+ $X2=0.78 $Y2=3.33
r225 73 75 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=0.625 $Y=3.33
+ $X2=0.24 $Y2=3.33
r226 71 103 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=6 $Y=3.33
+ $X2=7.44 $Y2=3.33
r227 71 131 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33
+ $X2=5.52 $Y2=3.33
r228 71 99 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r229 69 106 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=9.88 $Y=3.33
+ $X2=9.84 $Y2=3.33
r230 69 70 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=9.88 $Y=3.33
+ $X2=10.01 $Y2=3.33
r231 68 110 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=10.14 $Y=3.33
+ $X2=10.32 $Y2=3.33
r232 68 70 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=10.14 $Y=3.33
+ $X2=10.01 $Y2=3.33
r233 64 67 26.8903 $w=3.28e-07 $l=7.7e-07 $layer=LI1_cond $X=11.73 $Y=2.18
+ $X2=11.73 $Y2=2.95
r234 62 143 3.00555 $w=3.3e-07 $l=1.07912e-07 $layer=LI1_cond $X=11.73 $Y=3.245
+ $X2=11.782 $Y2=3.33
r235 62 67 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=11.73 $Y=3.245
+ $X2=11.73 $Y2=2.95
r236 58 61 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=10.87 $Y=2.18
+ $X2=10.87 $Y2=2.97
r237 56 140 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.87 $Y=3.245
+ $X2=10.87 $Y2=3.33
r238 56 61 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=10.87 $Y=3.245
+ $X2=10.87 $Y2=2.97
r239 52 55 43.8815 $w=2.58e-07 $l=9.9e-07 $layer=LI1_cond $X=10.01 $Y=1.98
+ $X2=10.01 $Y2=2.97
r240 50 70 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=10.01 $Y=3.245
+ $X2=10.01 $Y2=3.33
r241 50 55 12.1893 $w=2.58e-07 $l=2.75e-07 $layer=LI1_cond $X=10.01 $Y=3.245
+ $X2=10.01 $Y2=2.97
r242 46 137 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.04 $Y=3.245
+ $X2=9.04 $Y2=3.33
r243 46 48 17.8105 $w=3.28e-07 $l=5.1e-07 $layer=LI1_cond $X=9.04 $Y=3.245
+ $X2=9.04 $Y2=2.735
r244 45 134 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.045 $Y=3.33
+ $X2=7.88 $Y2=3.33
r245 44 137 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.875 $Y=3.33
+ $X2=9.04 $Y2=3.33
r246 44 45 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=8.875 $Y=3.33
+ $X2=8.045 $Y2=3.33
r247 40 134 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.88 $Y=3.245
+ $X2=7.88 $Y2=3.33
r248 40 42 17.8105 $w=3.28e-07 $l=5.1e-07 $layer=LI1_cond $X=7.88 $Y=3.245
+ $X2=7.88 $Y2=2.735
r249 36 124 0.512231 $w=2.15e-07 $l=8.5e-08 $layer=LI1_cond $X=4.042 $Y=3.245
+ $X2=4.042 $Y2=3.33
r250 36 38 15.2766 $w=2.13e-07 $l=2.85e-07 $layer=LI1_cond $X=4.042 $Y=3.245
+ $X2=4.042 $Y2=2.96
r251 32 121 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.255 $Y=3.245
+ $X2=2.255 $Y2=3.33
r252 32 34 11.5244 $w=3.28e-07 $l=3.3e-07 $layer=LI1_cond $X=2.255 $Y=3.245
+ $X2=2.255 $Y2=2.915
r253 28 118 0.701276 $w=3.1e-07 $l=8.5e-08 $layer=LI1_cond $X=0.78 $Y=3.245
+ $X2=0.78 $Y2=3.33
r254 28 30 16.3573 $w=3.08e-07 $l=4.4e-07 $layer=LI1_cond $X=0.78 $Y=3.245
+ $X2=0.78 $Y2=2.805
r255 9 67 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=11.59
+ $Y=1.835 $X2=11.73 $Y2=2.95
r256 9 64 400 $w=1.7e-07 $l=4.09054e-07 $layer=licon1_PDIFF $count=1 $X=11.59
+ $Y=1.835 $X2=11.73 $Y2=2.18
r257 8 61 400 $w=1.7e-07 $l=1.20297e-06 $layer=licon1_PDIFF $count=1 $X=10.73
+ $Y=1.835 $X2=10.87 $Y2=2.97
r258 8 58 400 $w=1.7e-07 $l=4.09054e-07 $layer=licon1_PDIFF $count=1 $X=10.73
+ $Y=1.835 $X2=10.87 $Y2=2.18
r259 7 55 400 $w=1.7e-07 $l=1.20297e-06 $layer=licon1_PDIFF $count=1 $X=9.87
+ $Y=1.835 $X2=10.01 $Y2=2.97
r260 7 52 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=9.87
+ $Y=1.835 $X2=10.01 $Y2=1.98
r261 6 48 600 $w=1.7e-07 $l=3.80197e-07 $layer=licon1_PDIFF $count=1 $X=8.845
+ $Y=2.44 $X2=9.04 $Y2=2.735
r262 5 42 600 $w=1.7e-07 $l=4.80364e-07 $layer=licon1_PDIFF $count=1 $X=7.525
+ $Y=2.44 $X2=7.88 $Y2=2.735
r263 4 127 600 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=5.295
+ $Y=2.245 $X2=5.44 $Y2=3.07
r264 3 38 600 $w=1.7e-07 $l=3.77492e-07 $layer=licon1_PDIFF $count=1 $X=3.805
+ $Y=2.675 $X2=4.02 $Y2=2.96
r265 2 34 600 $w=1.7e-07 $l=3.01993e-07 $layer=licon1_PDIFF $count=1 $X=2.115
+ $Y=2.675 $X2=2.255 $Y2=2.915
r266 1 30 600 $w=1.7e-07 $l=5.60647e-07 $layer=licon1_PDIFF $count=1 $X=0.65
+ $Y=2.31 $X2=0.79 $Y2=2.805
.ends

.subckt PM_SKY130_FD_SC_LP__DFRTP_4%A_340_535# 1 2 3 12 14 15 18 20 23 25 26 28
+ 33
c77 20 0 1.82197e-19 $X=3.255 $Y=2.54
c78 14 0 1.5785e-19 $X=2.59 $Y=2.54
r79 28 30 7.86138 $w=2.58e-07 $l=1.65e-07 $layer=LI1_cond $X=3.12 $Y=0.89
+ $X2=3.12 $Y2=1.055
r80 24 33 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.34 $Y=1.915
+ $X2=3.34 $Y2=1.83
r81 24 25 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=3.34 $Y=1.915
+ $X2=3.34 $Y2=2.455
r82 23 33 16.1797 $w=1.68e-07 $l=2.48e-07 $layer=LI1_cond $X=3.092 $Y=1.83
+ $X2=3.34 $Y2=1.83
r83 23 30 37.3304 $w=2.03e-07 $l=6.9e-07 $layer=LI1_cond $X=3.092 $Y=1.745
+ $X2=3.092 $Y2=1.055
r84 21 26 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=2.82 $Y=2.54
+ $X2=2.705 $Y2=2.54
r85 20 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.255 $Y=2.54
+ $X2=3.34 $Y2=2.455
r86 20 21 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=3.255 $Y=2.54
+ $X2=2.82 $Y2=2.54
r87 16 26 0.280307 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.705 $Y=2.625
+ $X2=2.705 $Y2=2.54
r88 16 18 13.0276 $w=2.28e-07 $l=2.6e-07 $layer=LI1_cond $X=2.705 $Y=2.625
+ $X2=2.705 $Y2=2.885
r89 14 26 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=2.59 $Y=2.54
+ $X2=2.705 $Y2=2.54
r90 14 15 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.59 $Y=2.54
+ $X2=1.92 $Y2=2.54
r91 10 15 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=1.79 $Y=2.625
+ $X2=1.92 $Y2=2.54
r92 10 12 11.5244 $w=2.58e-07 $l=2.6e-07 $layer=LI1_cond $X=1.79 $Y=2.625
+ $X2=1.79 $Y2=2.885
r93 3 18 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=2.545
+ $Y=2.675 $X2=2.685 $Y2=2.885
r94 2 12 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=1.7
+ $Y=2.675 $X2=1.825 $Y2=2.885
r95 1 28 182 $w=1.7e-07 $l=3.58225e-07 $layer=licon1_NDIFF $count=1 $X=3.015
+ $Y=0.595 $X2=3.155 $Y2=0.89
.ends

.subckt PM_SKY130_FD_SC_LP__DFRTP_4%Q 1 2 3 4 15 19 23 24 25 26 29 33 35 38 40
+ 41 42 45
r61 42 45 23.7544 $w=2.43e-07 $l=5.05e-07 $layer=LI1_cond $X=11.272 $Y=0.925
+ $X2=11.272 $Y2=0.42
r62 39 42 6.58539 $w=2.43e-07 $l=1.4e-07 $layer=LI1_cond $X=11.272 $Y=1.065
+ $X2=11.272 $Y2=0.925
r63 39 40 0.066131 $w=2.45e-07 $l=8.5e-08 $layer=LI1_cond $X=11.272 $Y=1.065
+ $X2=11.272 $Y2=1.15
r64 37 38 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=11.765 $Y=1.235
+ $X2=11.765 $Y2=1.755
r65 36 41 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=11.395 $Y=1.84
+ $X2=11.3 $Y2=1.84
r66 35 38 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=11.68 $Y=1.84
+ $X2=11.765 $Y2=1.755
r67 35 36 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=11.68 $Y=1.84
+ $X2=11.395 $Y2=1.84
r68 34 40 6.92067 $w=1.7e-07 $l=1.23e-07 $layer=LI1_cond $X=11.395 $Y=1.15
+ $X2=11.272 $Y2=1.15
r69 33 37 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=11.68 $Y=1.15
+ $X2=11.765 $Y2=1.235
r70 33 34 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=11.68 $Y=1.15
+ $X2=11.395 $Y2=1.15
r71 29 31 55.4545 $w=1.88e-07 $l=9.5e-07 $layer=LI1_cond $X=11.3 $Y=1.96
+ $X2=11.3 $Y2=2.91
r72 27 41 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=11.3 $Y=1.925
+ $X2=11.3 $Y2=1.84
r73 27 29 2.04306 $w=1.88e-07 $l=3.5e-08 $layer=LI1_cond $X=11.3 $Y=1.925
+ $X2=11.3 $Y2=1.96
r74 25 41 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=11.205 $Y=1.84
+ $X2=11.3 $Y2=1.84
r75 25 26 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=11.205 $Y=1.84
+ $X2=10.535 $Y2=1.84
r76 23 40 6.92067 $w=1.7e-07 $l=1.22e-07 $layer=LI1_cond $X=11.15 $Y=1.15
+ $X2=11.272 $Y2=1.15
r77 23 24 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=11.15 $Y=1.15
+ $X2=10.535 $Y2=1.15
r78 19 21 48.6587 $w=2.23e-07 $l=9.5e-07 $layer=LI1_cond $X=10.422 $Y=1.96
+ $X2=10.422 $Y2=2.91
r79 17 26 6.9898 $w=1.7e-07 $l=1.49579e-07 $layer=LI1_cond $X=10.422 $Y=1.925
+ $X2=10.535 $Y2=1.84
r80 17 19 1.79269 $w=2.23e-07 $l=3.5e-08 $layer=LI1_cond $X=10.422 $Y=1.925
+ $X2=10.422 $Y2=1.96
r81 13 24 6.9898 $w=1.7e-07 $l=1.49579e-07 $layer=LI1_cond $X=10.422 $Y=1.065
+ $X2=10.535 $Y2=1.15
r82 13 15 33.0367 $w=2.23e-07 $l=6.45e-07 $layer=LI1_cond $X=10.422 $Y=1.065
+ $X2=10.422 $Y2=0.42
r83 4 31 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=11.16
+ $Y=1.835 $X2=11.3 $Y2=2.91
r84 4 29 400 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=11.16
+ $Y=1.835 $X2=11.3 $Y2=1.96
r85 3 21 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=10.3
+ $Y=1.835 $X2=10.44 $Y2=2.91
r86 3 19 400 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=10.3
+ $Y=1.835 $X2=10.44 $Y2=1.96
r87 2 45 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=11.16
+ $Y=0.235 $X2=11.3 $Y2=0.42
r88 1 15 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=10.3
+ $Y=0.235 $X2=10.44 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__DFRTP_4%VGND 1 2 3 4 5 6 7 24 28 32 36 40 42 44 47
+ 48 49 50 57 58 59 61 79 90 94 100 103 106 110
c135 110 0 6.26159e-21 $X=11.76 $Y=0
c136 1 0 1.11939e-19 $X=0.55 $Y=0.45
r137 109 110 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.76 $Y=0
+ $X2=11.76 $Y2=0
r138 106 107 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=0
+ $X2=10.8 $Y2=0
r139 103 104 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=7.92 $Y=0
+ $X2=7.92 $Y2=0
r140 100 101 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0
+ $X2=0.72 $Y2=0
r141 98 110 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=0
+ $X2=11.76 $Y2=0
r142 98 107 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=0
+ $X2=10.8 $Y2=0
r143 97 98 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.28 $Y=0
+ $X2=11.28 $Y2=0
r144 95 106 7.54988 $w=1.7e-07 $l=1.38e-07 $layer=LI1_cond $X=10.98 $Y=0
+ $X2=10.842 $Y2=0
r145 95 97 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=10.98 $Y=0 $X2=11.28
+ $Y2=0
r146 94 109 4.76062 $w=1.7e-07 $l=2.17e-07 $layer=LI1_cond $X=11.565 $Y=0
+ $X2=11.782 $Y2=0
r147 94 97 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=11.565 $Y=0
+ $X2=11.28 $Y2=0
r148 93 107 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=0
+ $X2=10.8 $Y2=0
r149 92 93 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.32 $Y=0
+ $X2=10.32 $Y2=0
r150 90 106 7.54988 $w=1.7e-07 $l=1.37e-07 $layer=LI1_cond $X=10.705 $Y=0
+ $X2=10.842 $Y2=0
r151 90 92 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=10.705 $Y=0
+ $X2=10.32 $Y2=0
r152 89 93 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.84 $Y=0
+ $X2=10.32 $Y2=0
r153 88 89 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.84 $Y=0 $X2=9.84
+ $Y2=0
r154 86 89 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=8.4 $Y=0 $X2=9.84
+ $Y2=0
r155 86 104 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=0 $X2=7.92
+ $Y2=0
r156 85 88 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=8.4 $Y=0 $X2=9.84
+ $Y2=0
r157 85 86 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r158 83 103 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.225 $Y=0
+ $X2=8.06 $Y2=0
r159 83 85 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=8.225 $Y=0 $X2=8.4
+ $Y2=0
r160 81 82 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r161 79 103 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.895 $Y=0
+ $X2=8.06 $Y2=0
r162 79 81 154.947 $w=1.68e-07 $l=2.375e-06 $layer=LI1_cond $X=7.895 $Y=0
+ $X2=5.52 $Y2=0
r163 78 82 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=5.52
+ $Y2=0
r164 77 78 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r165 75 78 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=2.64 $Y=0 $X2=5.04
+ $Y2=0
r166 74 77 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=2.64 $Y=0 $X2=5.04
+ $Y2=0
r167 74 75 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r168 72 75 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r169 71 72 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r170 69 72 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r171 69 101 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r172 68 71 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r173 68 69 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r174 66 100 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=0.865 $Y=0
+ $X2=0.695 $Y2=0
r175 66 68 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=0.865 $Y=0 $X2=1.2
+ $Y2=0
r176 64 101 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0
+ $X2=0.72 $Y2=0
r177 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r178 61 100 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=0.525 $Y=0
+ $X2=0.695 $Y2=0
r179 61 63 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.525 $Y=0
+ $X2=0.24 $Y2=0
r180 59 104 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=6 $Y=0 $X2=7.92
+ $Y2=0
r181 59 82 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=5.52
+ $Y2=0
r182 57 88 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=9.88 $Y=0 $X2=9.84
+ $Y2=0
r183 57 58 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=9.88 $Y=0 $X2=10.01
+ $Y2=0
r184 56 92 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=10.14 $Y=0
+ $X2=10.32 $Y2=0
r185 56 58 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=10.14 $Y=0 $X2=10.01
+ $Y2=0
r186 52 81 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=5.485 $Y=0 $X2=5.52
+ $Y2=0
r187 50 77 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=5.155 $Y=0
+ $X2=5.04 $Y2=0
r188 49 54 9.07985 $w=3.28e-07 $l=2.6e-07 $layer=LI1_cond $X=5.32 $Y=0 $X2=5.32
+ $Y2=0.26
r189 49 52 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.32 $Y=0 $X2=5.485
+ $Y2=0
r190 49 50 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.32 $Y=0 $X2=5.155
+ $Y2=0
r191 47 71 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=2.235 $Y=0 $X2=2.16
+ $Y2=0
r192 47 48 6.92067 $w=1.7e-07 $l=1.22e-07 $layer=LI1_cond $X=2.235 $Y=0
+ $X2=2.357 $Y2=0
r193 46 74 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=2.48 $Y=0 $X2=2.64
+ $Y2=0
r194 46 48 6.92067 $w=1.7e-07 $l=1.23e-07 $layer=LI1_cond $X=2.48 $Y=0 $X2=2.357
+ $Y2=0
r195 42 109 3.00555 $w=3.3e-07 $l=1.07912e-07 $layer=LI1_cond $X=11.73 $Y=0.085
+ $X2=11.782 $Y2=0
r196 42 44 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=11.73 $Y=0.085
+ $X2=11.73 $Y2=0.38
r197 38 106 0.316938 $w=2.75e-07 $l=8.5e-08 $layer=LI1_cond $X=10.842 $Y=0.085
+ $X2=10.842 $Y2=0
r198 38 40 11.5244 $w=2.73e-07 $l=2.75e-07 $layer=LI1_cond $X=10.842 $Y=0.085
+ $X2=10.842 $Y2=0.36
r199 34 58 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=10.01 $Y=0.085
+ $X2=10.01 $Y2=0
r200 34 36 12.1893 $w=2.58e-07 $l=2.75e-07 $layer=LI1_cond $X=10.01 $Y=0.085
+ $X2=10.01 $Y2=0.36
r201 30 103 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.06 $Y=0.085
+ $X2=8.06 $Y2=0
r202 30 32 25.4934 $w=3.28e-07 $l=7.3e-07 $layer=LI1_cond $X=8.06 $Y=0.085
+ $X2=8.06 $Y2=0.815
r203 26 48 0.066131 $w=2.45e-07 $l=8.5e-08 $layer=LI1_cond $X=2.357 $Y=0.085
+ $X2=2.357 $Y2=0
r204 26 28 31.2806 $w=2.43e-07 $l=6.65e-07 $layer=LI1_cond $X=2.357 $Y=0.085
+ $X2=2.357 $Y2=0.75
r205 22 100 0.987631 $w=3.4e-07 $l=8.5e-08 $layer=LI1_cond $X=0.695 $Y=0.085
+ $X2=0.695 $Y2=0
r206 22 24 16.6087 $w=3.38e-07 $l=4.9e-07 $layer=LI1_cond $X=0.695 $Y=0.085
+ $X2=0.695 $Y2=0.575
r207 7 44 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=11.59
+ $Y=0.235 $X2=11.73 $Y2=0.38
r208 6 40 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=10.73
+ $Y=0.235 $X2=10.87 $Y2=0.36
r209 5 36 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=9.87
+ $Y=0.235 $X2=10.01 $Y2=0.36
r210 4 32 182 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_NDIFF $count=1 $X=7.785
+ $Y=0.665 $X2=8.06 $Y2=0.815
r211 3 54 182 $w=1.7e-07 $l=3.71214e-07 $layer=licon1_NDIFF $count=1 $X=5.065
+ $Y=0.525 $X2=5.32 $Y2=0.26
r212 2 28 182 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=1 $X=2.24
+ $Y=0.595 $X2=2.365 $Y2=0.75
r213 1 24 182 $w=1.7e-07 $l=2.03101e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.45 $X2=0.7 $Y2=0.575
.ends

