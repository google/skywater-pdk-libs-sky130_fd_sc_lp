* File: sky130_fd_sc_lp__dlrbp_1.spice
* Created: Fri Aug 28 10:25:55 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__dlrbp_1.pex.spice"
.subckt sky130_fd_sc_lp__dlrbp_1  VNB VPB GATE D RESET_B VPWR Q_N Q VGND
* 
* VGND	VGND
* Q	Q
* Q_N	Q_N
* VPWR	VPWR
* RESET_B	RESET_B
* D	D
* GATE	GATE
* VPB	VPB
* VNB	VNB
MM1004 N_VGND_M1004_d N_GATE_M1004_g N_A_49_93#_M1004_s VNB NSHORT L=0.15 W=0.42
+ AD=0.09135 AS=0.1113 PD=0.855 PS=1.37 NRD=22.848 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.8 A=0.063 P=1.14 MULT=1
MM1023 N_A_218_483#_M1023_d N_A_49_93#_M1023_g N_VGND_M1004_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1113 AS=0.09135 PD=1.37 PS=0.855 NRD=0 NRS=21.42 M=1 R=2.8
+ SA=75000.8 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1017 N_VGND_M1017_d N_D_M1017_g N_A_373_481#_M1017_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75001.9
+ A=0.063 P=1.14 MULT=1
MM1018 A_554_119# N_A_373_481#_M1018_g N_VGND_M1017_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75001.5 A=0.063 P=1.14 MULT=1
MM1015 N_A_626_119#_M1015_d N_A_218_483#_M1015_g A_554_119# VNB NSHORT L=0.15
+ W=0.42 AD=0.0819 AS=0.0441 PD=0.81 PS=0.63 NRD=15.708 NRS=14.28 M=1 R=2.8
+ SA=75001 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1021 A_734_119# N_A_49_93#_M1021_g N_A_626_119#_M1015_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.0819 PD=0.63 PS=0.81 NRD=14.28 NRS=15.708 M=1 R=2.8
+ SA=75001.5 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1019 N_VGND_M1019_d N_A_776_93#_M1019_g A_734_119# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.9
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1013 A_1000_47# N_A_626_119#_M1013_g N_A_776_93#_M1013_s VNB NSHORT L=0.15
+ W=0.84 AD=0.0882 AS=0.2226 PD=1.05 PS=2.21 NRD=7.14 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75000.8 A=0.126 P=1.98 MULT=1
MM1005 N_VGND_M1005_d N_RESET_B_M1005_g A_1000_47# VNB NSHORT L=0.15 W=0.84
+ AD=0.1988 AS=0.0882 PD=1.68667 PS=1.05 NRD=0 NRS=7.14 M=1 R=5.6 SA=75000.6
+ SB=75000.5 A=0.126 P=1.98 MULT=1
MM1007 N_A_1187_131#_M1007_d N_A_776_93#_M1007_g N_VGND_M1005_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.1113 AS=0.0994 PD=1.37 PS=0.843333 NRD=0 NRS=51.9 M=1 R=2.8
+ SA=75001.1 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1002 N_VGND_M1002_d N_A_1187_131#_M1002_g N_Q_N_M1002_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1239 AS=0.2226 PD=1.135 PS=2.21 NRD=2.136 NRS=0 M=1 R=5.6
+ SA=75000.2 SB=75000.6 A=0.126 P=1.98 MULT=1
MM1008 N_Q_M1008_d N_A_776_93#_M1008_g N_VGND_M1002_d VNB NSHORT L=0.15 W=0.84
+ AD=0.231 AS=0.1239 PD=2.23 PS=1.135 NRD=1.428 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1011 N_VPWR_M1011_d N_GATE_M1011_g N_A_49_93#_M1011_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.0896 AS=0.1696 PD=0.92 PS=1.81 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1020 N_A_218_483#_M1020_d N_A_49_93#_M1020_g N_VPWR_M1011_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1696 AS=0.0896 PD=1.81 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.6 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1003 N_VPWR_M1003_d N_D_M1003_g N_A_373_481#_M1003_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.176 AS=0.1696 PD=1.19 PS=1.81 NRD=83.0946 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75002.6 A=0.096 P=1.58 MULT=1
MM1009 A_596_481# N_A_373_481#_M1009_g N_VPWR_M1003_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0672 AS=0.176 PD=0.85 PS=1.19 NRD=15.3857 NRS=0 M=1 R=4.26667 SA=75000.9
+ SB=75001.9 A=0.096 P=1.58 MULT=1
MM1014 N_A_626_119#_M1014_d N_A_49_93#_M1014_g A_596_481# VPB PHIGHVT L=0.15
+ W=0.64 AD=0.130294 AS=0.0672 PD=1.22566 PS=0.85 NRD=0 NRS=15.3857 M=1
+ R=4.26667 SA=75001.2 SB=75001.5 A=0.096 P=1.58 MULT=1
MM1001 A_773_525# N_A_218_483#_M1001_g N_A_626_119#_M1014_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0924 AS=0.0855057 PD=0.86 PS=0.80434 NRD=77.3816 NRS=46.886 M=1
+ R=2.8 SA=75001.8 SB=75001.7 A=0.063 P=1.14 MULT=1
MM1010 N_VPWR_M1010_d N_A_776_93#_M1010_g A_773_525# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.095025 AS=0.0924 PD=0.8175 PS=0.86 NRD=44.5417 NRS=77.3816 M=1 R=2.8
+ SA=75002.4 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1006 N_A_776_93#_M1006_d N_A_626_119#_M1006_g N_VPWR_M1010_d VPB PHIGHVT
+ L=0.15 W=1.26 AD=0.1764 AS=0.285075 PD=1.54 PS=2.4525 NRD=0 NRS=0 M=1 R=8.4
+ SA=75001.1 SB=75000.9 A=0.189 P=2.82 MULT=1
MM1022 N_VPWR_M1022_d N_RESET_B_M1022_g N_A_776_93#_M1006_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.268115 AS=0.1764 PD=2.16853 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75001.5 SB=75000.5 A=0.189 P=2.82 MULT=1
MM1016 N_A_1187_131#_M1016_d N_A_776_93#_M1016_g N_VPWR_M1022_d VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.1696 AS=0.136185 PD=1.81 PS=1.10147 NRD=0 NRS=48.5605 M=1
+ R=4.26667 SA=75001.1 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1012 N_VPWR_M1012_d N_A_1187_131#_M1012_g N_Q_N_M1012_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1000 N_Q_M1000_d N_A_776_93#_M1000_g N_VPWR_M1012_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX24_noxref VNB VPB NWDIODE A=16.0268 P=20.91
*
.include "sky130_fd_sc_lp__dlrbp_1.pxi.spice"
*
.ends
*
*
