* File: sky130_fd_sc_lp__srdlrtp_1.pex.spice
* Created: Fri Aug 28 11:33:01 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__SRDLRTP_1%D 3 7 9 15
r22 12 15 39.3438 $w=3.3e-07 $l=2.25e-07 $layer=POLY_cond $X=0.27 $Y=1.245
+ $X2=0.495 $Y2=1.245
r23 9 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=1.245 $X2=0.27 $Y2=1.245
r24 5 15 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.245
r25 5 7 689.67 $w=1.5e-07 $l=1.345e-06 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=2.755
r26 1 15 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=1.08
+ $X2=0.495 $Y2=1.245
r27 1 3 197.415 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=0.495 $Y=1.08
+ $X2=0.495 $Y2=0.695
.ends

.subckt PM_SKY130_FD_SC_LP__SRDLRTP_1%RESET_B 3 7 11 13 16 18 19 20 21 26 29 32
+ 37 38
c157 20 0 8.42426e-21 $X=9.215 $Y=2.035
r158 38 46 4.32554 $w=7.28e-07 $l=2.65e-07 $layer=LI1_cond $X=9.59 $Y=1.77
+ $X2=9.59 $Y2=2.035
r159 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.39
+ $Y=1.77 $X2=9.39 $Y2=1.77
r160 35 37 40.2181 $w=3.3e-07 $l=2.3e-07 $layer=POLY_cond $X=9.16 $Y=1.77
+ $X2=9.39 $Y2=1.77
r161 33 35 8.74306 $w=3.3e-07 $l=5e-08 $layer=POLY_cond $X=9.11 $Y=1.77 $X2=9.16
+ $Y2=1.77
r162 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.11
+ $Y=2.09 $X2=1.11 $Y2=2.09
r163 29 31 19.8674 $w=2.79e-07 $l=1.15e-07 $layer=POLY_cond $X=0.995 $Y=2.09
+ $X2=1.11 $Y2=2.09
r164 26 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=2.035
+ $X2=9.36 $Y2=2.035
r165 23 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=2.035
+ $X2=1.2 $Y2=2.035
r166 21 23 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.345 $Y=2.035
+ $X2=1.2 $Y2=2.035
r167 20 26 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=9.215 $Y=2.035
+ $X2=9.36 $Y2=2.035
r168 20 21 9.74008 $w=1.4e-07 $l=7.87e-06 $layer=MET1_cond $X=9.215 $Y=2.035
+ $X2=1.345 $Y2=2.035
r169 18 19 53.9552 $w=1.9e-07 $l=1.5e-07 $layer=POLY_cond $X=9.09 $Y=0.765
+ $X2=9.09 $Y2=0.915
r170 14 35 9.34494 $w=2.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.16 $Y=1.935
+ $X2=9.16 $Y2=1.77
r171 14 16 163.979 $w=2.5e-07 $l=6.6e-07 $layer=POLY_cond $X=9.16 $Y=1.935
+ $X2=9.16 $Y2=2.595
r172 13 33 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.11 $Y=1.605
+ $X2=9.11 $Y2=1.77
r173 13 19 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=9.11 $Y=1.605
+ $X2=9.11 $Y2=0.915
r174 11 18 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=9.07 $Y=0.445
+ $X2=9.07 $Y2=0.765
r175 5 29 17.2686 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.995 $Y=2.255
+ $X2=0.995 $Y2=2.09
r176 5 7 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=0.995 $Y=2.255
+ $X2=0.995 $Y2=2.755
r177 1 29 24.1864 $w=2.79e-07 $l=2.24332e-07 $layer=POLY_cond $X=0.855 $Y=1.925
+ $X2=0.995 $Y2=2.09
r178 1 3 630.702 $w=1.5e-07 $l=1.23e-06 $layer=POLY_cond $X=0.855 $Y=1.925
+ $X2=0.855 $Y2=0.695
.ends

.subckt PM_SKY130_FD_SC_LP__SRDLRTP_1%A_27_97# 1 2 9 12 15 17 19 22 27 29 33 34
+ 37 39 40 41
r91 40 41 8.63679 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=0.775 $Y=2.425
+ $X2=0.775 $Y2=2.595
r92 33 34 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.305
+ $Y=1.18 $X2=1.305 $Y2=1.18
r93 31 33 13.969 $w=3.28e-07 $l=4e-07 $layer=LI1_cond $X=1.305 $Y=1.58 $X2=1.305
+ $Y2=1.18
r94 30 39 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.775 $Y=1.665
+ $X2=0.69 $Y2=1.665
r95 29 31 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.14 $Y=1.665
+ $X2=1.305 $Y2=1.58
r96 29 30 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=1.14 $Y=1.665
+ $X2=0.775 $Y2=1.665
r97 27 41 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=0.78 $Y=2.75
+ $X2=0.78 $Y2=2.595
r98 23 39 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=1.75 $X2=0.69
+ $Y2=1.665
r99 23 40 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=0.69 $Y=1.75
+ $X2=0.69 $Y2=2.425
r100 22 39 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=1.58
+ $X2=0.69 $Y2=1.665
r101 21 37 16.2932 $w=3.07e-07 $l=5.09441e-07 $layer=LI1_cond $X=0.69 $Y=0.91
+ $X2=0.28 $Y2=0.687
r102 21 22 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=0.69 $Y=0.91
+ $X2=0.69 $Y2=1.58
r103 17 34 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=1.305 $Y=1.535
+ $X2=1.305 $Y2=1.18
r104 17 19 156.394 $w=1.5e-07 $l=3.05e-07 $layer=POLY_cond $X=1.305 $Y=1.61
+ $X2=1.61 $Y2=1.61
r105 15 34 38.6168 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.305 $Y=1.015
+ $X2=1.305 $Y2=1.18
r106 10 19 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.61 $Y=1.685
+ $X2=1.61 $Y2=1.61
r107 10 12 548.66 $w=1.5e-07 $l=1.07e-06 $layer=POLY_cond $X=1.61 $Y=1.685
+ $X2=1.61 $Y2=2.755
r108 9 15 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.325 $Y=0.695
+ $X2=1.325 $Y2=1.015
r109 2 27 600 $w=1.7e-07 $l=4.06663e-07 $layer=licon1_PDIFF $count=1 $X=0.57
+ $Y=2.435 $X2=0.78 $Y2=2.75
r110 1 37 182 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.485 $X2=0.28 $Y2=0.685
.ends

.subckt PM_SKY130_FD_SC_LP__SRDLRTP_1%A_336_71# 1 2 9 11 12 15 19 23 24 25 27 28
+ 29 32 33 34 36 37 38 40 42 44 51 57 61 63
c198 63 0 8.42426e-21 $X=2.165 $Y=1.17
c199 57 0 1.21577e-19 $X=7.755 $Y=0.34
r200 63 64 30.474 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=2.165 $Y=1.17
+ $X2=2.165 $Y2=1.095
r201 61 69 32.0725 $w=3.45e-07 $l=1.65e-07 $layer=POLY_cond $X=7.747 $Y=0.42
+ $X2=7.747 $Y2=0.585
r202 60 61 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.755
+ $Y=0.42 $X2=7.755 $Y2=0.42
r203 57 60 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=7.755 $Y=0.34
+ $X2=7.755 $Y2=0.42
r204 54 56 2.02539 $w=5.12e-07 $l=8.5e-08 $layer=LI1_cond $X=4.217 $Y=0.61
+ $X2=4.217 $Y2=0.695
r205 53 54 6.43359 $w=5.12e-07 $l=2.7e-07 $layer=LI1_cond $X=4.217 $Y=0.34
+ $X2=4.217 $Y2=0.61
r206 49 51 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=3.805 $Y=2.04
+ $X2=3.985 $Y2=2.04
r207 44 46 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=2.925 $Y=0.34
+ $X2=2.925 $Y2=0.61
r208 41 63 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=2.165 $Y=1.26
+ $X2=2.165 $Y2=1.17
r209 40 42 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=2.165 $Y=1.26
+ $X2=2.165 $Y2=1.095
r210 40 41 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.165
+ $Y=1.26 $X2=2.165 $Y2=1.26
r211 37 57 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.59 $Y=0.34
+ $X2=7.755 $Y2=0.34
r212 37 38 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=7.59 $Y=0.34 $X2=7
+ $Y2=0.34
r213 35 38 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.915 $Y=0.425
+ $X2=7 $Y2=0.34
r214 35 36 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=6.915 $Y=0.425
+ $X2=6.915 $Y2=0.8
r215 33 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.83 $Y=0.885
+ $X2=6.915 $Y2=0.8
r216 33 34 55.7807 $w=1.68e-07 $l=8.55e-07 $layer=LI1_cond $X=6.83 $Y=0.885
+ $X2=5.975 $Y2=0.885
r217 32 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.89 $Y=0.8
+ $X2=5.975 $Y2=0.885
r218 31 32 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=5.89 $Y=0.425
+ $X2=5.89 $Y2=0.8
r219 30 53 7.30583 $w=1.7e-07 $l=3.18e-07 $layer=LI1_cond $X=4.535 $Y=0.34
+ $X2=4.217 $Y2=0.34
r220 29 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.805 $Y=0.34
+ $X2=5.89 $Y2=0.425
r221 29 30 82.8556 $w=1.68e-07 $l=1.27e-06 $layer=LI1_cond $X=5.805 $Y=0.34
+ $X2=4.535 $Y2=0.34
r222 28 51 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.985 $Y=1.955
+ $X2=3.985 $Y2=2.04
r223 27 56 11.3319 $w=5.12e-07 $l=3.2739e-07 $layer=LI1_cond $X=3.985 $Y=0.925
+ $X2=4.217 $Y2=0.695
r224 27 28 67.1979 $w=1.68e-07 $l=1.03e-06 $layer=LI1_cond $X=3.985 $Y=0.925
+ $X2=3.985 $Y2=1.955
r225 26 46 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.01 $Y=0.61
+ $X2=2.925 $Y2=0.61
r226 25 54 7.30583 $w=1.7e-07 $l=3.17e-07 $layer=LI1_cond $X=3.9 $Y=0.61
+ $X2=4.217 $Y2=0.61
r227 25 26 58.0642 $w=1.68e-07 $l=8.9e-07 $layer=LI1_cond $X=3.9 $Y=0.61
+ $X2=3.01 $Y2=0.61
r228 23 44 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.84 $Y=0.34
+ $X2=2.925 $Y2=0.34
r229 23 24 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.84 $Y=0.34
+ $X2=2.17 $Y2=0.34
r230 21 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.085 $Y=0.425
+ $X2=2.17 $Y2=0.34
r231 21 42 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.085 $Y=0.425
+ $X2=2.085 $Y2=1.095
r232 19 69 499.392 $w=2.5e-07 $l=2.01e-06 $layer=POLY_cond $X=7.7 $Y=2.595
+ $X2=7.7 $Y2=0.585
r233 15 64 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=2.115 $Y=0.695
+ $X2=2.115 $Y2=1.095
r234 11 63 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2 $Y=1.17
+ $X2=2.165 $Y2=1.17
r235 11 12 87.1702 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=2 $Y=1.17 $X2=1.83
+ $Y2=1.17
r236 7 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.755 $Y=1.095
+ $X2=1.83 $Y2=1.17
r237 7 9 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=1.755 $Y=1.095
+ $X2=1.755 $Y2=0.695
r238 2 49 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=3.66
+ $Y=1.9 $X2=3.805 $Y2=2.04
r239 1 56 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=4.23
+ $Y=0.485 $X2=4.37 $Y2=0.695
.ends

.subckt PM_SKY130_FD_SC_LP__SRDLRTP_1%A_612_71# 1 2 9 13 17 20 21 22 24 25 26 28
+ 29 30 32 34 35 39 42 46 52 53 55 57 59 65
c201 29 0 5.91988e-20 $X=7.93 $Y=2.99
c202 17 0 4.70163e-20 $X=8.16 $Y=2.595
r203 59 61 9.9374 $w=3.73e-07 $l=2.1e-07 $layer=LI1_cond $X=10.107 $Y=0.465
+ $X2=10.107 $Y2=0.675
r204 53 69 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.2 $Y=1.77
+ $X2=8.2 $Y2=1.935
r205 52 53 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.2
+ $Y=1.77 $X2=8.2 $Y2=1.77
r206 49 52 7.35179 $w=2.88e-07 $l=1.85e-07 $layer=LI1_cond $X=8.015 $Y=1.79
+ $X2=8.2 $Y2=1.79
r207 47 65 47.2125 $w=3.3e-07 $l=2.7e-07 $layer=POLY_cond $X=3.225 $Y=1.3
+ $X2=3.495 $Y2=1.3
r208 47 62 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=3.225 $Y=1.3
+ $X2=3.135 $Y2=1.3
r209 46 47 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.225
+ $Y=1.3 $X2=3.225 $Y2=1.3
r210 43 46 8.64332 $w=2.38e-07 $l=1.8e-07 $layer=LI1_cond $X=3.045 $Y=1.325
+ $X2=3.225 $Y2=1.325
r211 42 61 107.321 $w=1.68e-07 $l=1.645e-06 $layer=LI1_cond $X=10.21 $Y=2.32
+ $X2=10.21 $Y2=0.675
r212 40 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.705 $Y=2.405
+ $X2=9.54 $Y2=2.405
r213 39 42 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.125 $Y=2.405
+ $X2=10.21 $Y2=2.32
r214 39 40 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=10.125 $Y=2.405
+ $X2=9.705 $Y2=2.405
r215 36 55 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.1 $Y=2.405
+ $X2=8.015 $Y2=2.405
r216 35 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.375 $Y=2.405
+ $X2=9.54 $Y2=2.405
r217 35 36 83.1818 $w=1.68e-07 $l=1.275e-06 $layer=LI1_cond $X=9.375 $Y=2.405
+ $X2=8.1 $Y2=2.405
r218 33 55 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.015 $Y=2.49
+ $X2=8.015 $Y2=2.405
r219 33 34 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=8.015 $Y=2.49
+ $X2=8.015 $Y2=2.905
r220 32 55 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.015 $Y=2.32
+ $X2=8.015 $Y2=2.405
r221 31 49 3.86198 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=8.015 $Y=1.935
+ $X2=8.015 $Y2=1.79
r222 31 32 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=8.015 $Y=1.935
+ $X2=8.015 $Y2=2.32
r223 29 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.93 $Y=2.99
+ $X2=8.015 $Y2=2.905
r224 29 30 77.9626 $w=1.68e-07 $l=1.195e-06 $layer=LI1_cond $X=7.93 $Y=2.99
+ $X2=6.735 $Y2=2.99
r225 28 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.65 $Y=2.905
+ $X2=6.735 $Y2=2.99
r226 27 28 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=6.65 $Y=2.49
+ $X2=6.65 $Y2=2.905
r227 25 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.565 $Y=2.405
+ $X2=6.65 $Y2=2.49
r228 25 26 117.107 $w=1.68e-07 $l=1.795e-06 $layer=LI1_cond $X=6.565 $Y=2.405
+ $X2=4.77 $Y2=2.405
r229 23 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.685 $Y=2.49
+ $X2=4.77 $Y2=2.405
r230 23 24 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=4.685 $Y=2.49
+ $X2=4.685 $Y2=2.635
r231 21 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.6 $Y=2.72
+ $X2=4.685 $Y2=2.635
r232 21 22 95.9037 $w=1.68e-07 $l=1.47e-06 $layer=LI1_cond $X=4.6 $Y=2.72
+ $X2=3.13 $Y2=2.72
r233 20 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.045 $Y=2.635
+ $X2=3.13 $Y2=2.72
r234 19 43 2.75731 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=3.045 $Y=1.445
+ $X2=3.045 $Y2=1.325
r235 19 20 77.6364 $w=1.68e-07 $l=1.19e-06 $layer=LI1_cond $X=3.045 $Y=1.445
+ $X2=3.045 $Y2=2.635
r236 17 69 163.979 $w=2.5e-07 $l=6.6e-07 $layer=POLY_cond $X=8.16 $Y=2.595
+ $X2=8.16 $Y2=1.935
r237 11 65 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.495 $Y=1.135
+ $X2=3.495 $Y2=1.3
r238 11 13 225.617 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=3.495 $Y=1.135
+ $X2=3.495 $Y2=0.695
r239 7 62 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.135 $Y=1.135
+ $X2=3.135 $Y2=1.3
r240 7 9 225.617 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=3.135 $Y=1.135
+ $X2=3.135 $Y2=0.695
r241 2 57 300 $w=1.7e-07 $l=5.01548e-07 $layer=licon1_PDIFF $count=2 $X=9.285
+ $Y=2.095 $X2=9.54 $Y2=2.485
r242 1 59 182 $w=1.7e-07 $l=2.91719e-07 $layer=licon1_NDIFF $count=1 $X=9.945
+ $Y=0.235 $X2=10.085 $Y2=0.465
.ends

.subckt PM_SKY130_FD_SC_LP__SRDLRTP_1%A_393_335# 1 2 9 11 12 15 17 21 23 25 27
+ 30 32 33 35 38 40 43 45 49
c123 30 0 1.8278e-19 $X=4.155 $Y=0.695
c124 21 0 3.39925e-20 $X=2.775 $Y=0.695
r125 46 49 9.39684 $w=3.23e-07 $l=2.65e-07 $layer=LI1_cond $X=4.79 $Y=0.757
+ $X2=5.055 $Y2=0.757
r126 44 52 36.7822 $w=6.29e-07 $l=4.8e-07 $layer=POLY_cond $X=4.382 $Y=1.27
+ $X2=4.382 $Y2=1.75
r127 43 45 9.51712 $w=4.98e-07 $l=1.65e-07 $layer=LI1_cond $X=4.625 $Y=1.27
+ $X2=4.625 $Y2=1.105
r128 43 44 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.54
+ $Y=1.27 $X2=4.54 $Y2=1.27
r129 38 40 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=4.875 $Y=1.725
+ $X2=5.57 $Y2=1.725
r130 36 46 4.53325 $w=1.7e-07 $l=1.63e-07 $layer=LI1_cond $X=4.79 $Y=0.92
+ $X2=4.79 $Y2=0.757
r131 36 45 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=4.79 $Y=0.92
+ $X2=4.79 $Y2=1.105
r132 35 38 9.23067 $w=1.7e-07 $l=2.89396e-07 $layer=LI1_cond $X=4.625 $Y=1.64
+ $X2=4.875 $Y2=1.725
r133 34 43 2.03333 $w=4.98e-07 $l=8.5e-08 $layer=LI1_cond $X=4.625 $Y=1.355
+ $X2=4.625 $Y2=1.27
r134 34 35 6.81765 $w=4.98e-07 $l=2.85e-07 $layer=LI1_cond $X=4.625 $Y=1.355
+ $X2=4.625 $Y2=1.64
r135 28 44 45.3624 $w=6.29e-07 $l=2.98302e-07 $layer=POLY_cond $X=4.155 $Y=1.105
+ $X2=4.382 $Y2=1.27
r136 28 30 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=4.155 $Y=1.105
+ $X2=4.155 $Y2=0.695
r137 25 52 38.4657 $w=6.29e-07 $l=2.82018e-07 $layer=POLY_cond $X=4.135 $Y=1.825
+ $X2=4.382 $Y2=1.75
r138 25 27 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=4.135 $Y=1.825
+ $X2=4.135 $Y2=2.255
r139 24 33 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.85 $Y=1.75
+ $X2=2.775 $Y2=1.75
r140 23 52 37.3022 $w=1.5e-07 $l=3.22e-07 $layer=POLY_cond $X=4.06 $Y=1.75
+ $X2=4.382 $Y2=1.75
r141 23 24 620.447 $w=1.5e-07 $l=1.21e-06 $layer=POLY_cond $X=4.06 $Y=1.75
+ $X2=2.85 $Y2=1.75
r142 19 33 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.775 $Y=1.675
+ $X2=2.775 $Y2=1.75
r143 19 21 502.511 $w=1.5e-07 $l=9.8e-07 $layer=POLY_cond $X=2.775 $Y=1.675
+ $X2=2.775 $Y2=0.695
r144 18 32 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.475 $Y=1.75
+ $X2=2.4 $Y2=1.75
r145 17 33 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.7 $Y=1.75
+ $X2=2.775 $Y2=1.75
r146 17 18 115.372 $w=1.5e-07 $l=2.25e-07 $layer=POLY_cond $X=2.7 $Y=1.75
+ $X2=2.475 $Y2=1.75
r147 13 32 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.4 $Y=1.825
+ $X2=2.4 $Y2=1.75
r148 13 15 476.872 $w=1.5e-07 $l=9.3e-07 $layer=POLY_cond $X=2.4 $Y=1.825
+ $X2=2.4 $Y2=2.755
r149 11 32 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.325 $Y=1.75
+ $X2=2.4 $Y2=1.75
r150 11 12 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=2.325 $Y=1.75
+ $X2=2.115 $Y2=1.75
r151 7 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.04 $Y=1.825
+ $X2=2.115 $Y2=1.75
r152 7 9 476.872 $w=1.5e-07 $l=9.3e-07 $layer=POLY_cond $X=2.04 $Y=1.825
+ $X2=2.04 $Y2=2.755
r153 2 40 600 $w=1.7e-07 $l=7.21318e-07 $layer=licon1_PDIFF $count=1 $X=5.315
+ $Y=2.33 $X2=5.57 $Y2=1.725
r154 1 49 182 $w=1.7e-07 $l=2.93684e-07 $layer=licon1_NDIFF $count=1 $X=4.91
+ $Y=0.485 $X2=5.055 $Y2=0.715
.ends

.subckt PM_SKY130_FD_SC_LP__SRDLRTP_1%GATE 3 7 9 12
c42 12 0 1.90567e-19 $X=5.21 $Y=1.255
r43 12 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.21 $Y=1.255
+ $X2=5.21 $Y2=1.42
r44 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.21 $Y=1.255
+ $X2=5.21 $Y2=1.09
r45 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.21
+ $Y=1.255 $X2=5.21 $Y2=1.255
r46 9 13 10.826 $w=3.28e-07 $l=3.1e-07 $layer=LI1_cond $X=5.52 $Y=1.255 $X2=5.21
+ $Y2=1.255
r47 7 14 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=5.27 $Y=0.695
+ $X2=5.27 $Y2=1.09
r48 3 15 630.702 $w=1.5e-07 $l=1.23e-06 $layer=POLY_cond $X=5.24 $Y=2.65
+ $X2=5.24 $Y2=1.42
.ends

.subckt PM_SKY130_FD_SC_LP__SRDLRTP_1%SLEEP_B 3 7 11 15 19 21 22 25 27 28
c88 28 0 1.90567e-19 $X=6.48 $Y=1.295
r89 37 38 24.8454 $w=2.91e-07 $l=1.5e-07 $layer=POLY_cond $X=6.495 $Y=1.305
+ $X2=6.645 $Y2=1.305
r90 35 37 14.9072 $w=2.91e-07 $l=9e-08 $layer=POLY_cond $X=6.405 $Y=1.305
+ $X2=6.495 $Y2=1.305
r91 33 35 63.7698 $w=2.91e-07 $l=3.85e-07 $layer=POLY_cond $X=6.02 $Y=1.305
+ $X2=6.405 $Y2=1.305
r92 32 33 19.8763 $w=2.91e-07 $l=1.2e-07 $layer=POLY_cond $X=5.9 $Y=1.305
+ $X2=6.02 $Y2=1.305
r93 28 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.405
+ $Y=1.305 $X2=6.405 $Y2=1.305
r94 27 28 14.1436 $w=3.28e-07 $l=4.05e-07 $layer=LI1_cond $X=6 $Y=1.305
+ $X2=6.405 $Y2=1.305
r95 23 25 228.181 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=7.005 $Y=1.14
+ $X2=7.005 $Y2=0.695
r96 22 38 23.6999 $w=2.91e-07 $l=1.21861e-07 $layer=POLY_cond $X=6.72 $Y=1.215
+ $X2=6.645 $Y2=1.305
r97 21 23 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.93 $Y=1.215
+ $X2=7.005 $Y2=1.14
r98 21 22 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=6.93 $Y=1.215
+ $X2=6.72 $Y2=1.215
r99 17 38 18.2534 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.645 $Y=1.14
+ $X2=6.645 $Y2=1.305
r100 17 19 228.181 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=6.645 $Y=1.14
+ $X2=6.645 $Y2=0.695
r101 13 37 6.42794 $w=2.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.495 $Y=1.47
+ $X2=6.495 $Y2=1.305
r102 13 15 248.454 $w=2.5e-07 $l=1e-06 $layer=POLY_cond $X=6.495 $Y=1.47
+ $X2=6.495 $Y2=2.47
r103 9 33 18.2534 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.02 $Y=1.14
+ $X2=6.02 $Y2=1.305
r104 9 11 228.181 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=6.02 $Y=1.14
+ $X2=6.02 $Y2=0.695
r105 5 32 18.2534 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.9 $Y=1.47 $X2=5.9
+ $Y2=1.305
r106 5 7 605.064 $w=1.5e-07 $l=1.18e-06 $layer=POLY_cond $X=5.9 $Y=1.47 $X2=5.9
+ $Y2=2.65
r107 1 32 39.7526 $w=2.91e-07 $l=3.11769e-07 $layer=POLY_cond $X=5.66 $Y=1.14
+ $X2=5.9 $Y2=1.305
r108 1 3 228.181 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=5.66 $Y=1.14
+ $X2=5.66 $Y2=0.695
.ends

.subckt PM_SKY130_FD_SC_LP__SRDLRTP_1%A_1324_394# 1 2 9 11 13 16 19 21 23 27
c86 13 0 5.91988e-20 $X=8.7 $Y=2.595
c87 9 0 1.21577e-19 $X=8.48 $Y=0.445
r88 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.55
+ $Y=1.005 $X2=8.55 $Y2=1.005
r89 21 23 50.0869 $w=2.58e-07 $l=1.13e-06 $layer=LI1_cond $X=7.42 $Y=1.005
+ $X2=8.55 $Y2=1.005
r90 17 21 5.41659 $w=2.9e-07 $l=1.25996e-07 $layer=LI1_cond $X=7.295 $Y=1.007
+ $X2=7.42 $Y2=1.005
r91 17 19 5.30124 $w=2.48e-07 $l=1.15e-07 $layer=LI1_cond $X=7.295 $Y=0.875
+ $X2=7.295 $Y2=0.76
r92 16 27 0.716491 $w=1.7e-07 $l=1.18427e-07 $layer=LI1_cond $X=6.955 $Y=1.64
+ $X2=6.875 $Y2=1.725
r93 15 17 14.3034 $w=2.9e-07 $l=4.67568e-07 $layer=LI1_cond $X=6.955 $Y=1.31
+ $X2=7.295 $Y2=1.007
r94 15 16 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=6.955 $Y=1.31
+ $X2=6.955 $Y2=1.64
r95 11 24 44.0745 $w=3.72e-07 $l=3.44238e-07 $layer=POLY_cond $X=8.7 $Y=1.305
+ $X2=8.605 $Y2=1.005
r96 11 13 320.505 $w=2.5e-07 $l=1.29e-06 $layer=POLY_cond $X=8.7 $Y=1.305
+ $X2=8.7 $Y2=2.595
r97 7 24 39.087 $w=3.72e-07 $l=2.18746e-07 $layer=POLY_cond $X=8.48 $Y=0.84
+ $X2=8.605 $Y2=1.005
r98 7 9 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=8.48 $Y=0.84 $X2=8.48
+ $Y2=0.445
r99 2 27 600 $w=1.7e-07 $l=3.57071e-07 $layer=licon1_PDIFF $count=1 $X=6.62
+ $Y=1.97 $X2=6.875 $Y2=1.725
r100 1 19 182 $w=1.7e-07 $l=3.81772e-07 $layer=licon1_NDIFF $count=1 $X=7.08
+ $Y=0.485 $X2=7.335 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_LP__SRDLRTP_1%A_438_97# 1 2 3 12 16 20 22 23 26 30 32 33
+ 35 37 39 42 43 44 46 48 49 50 53 56 58 61 67 70 72 73 74
c226 56 0 4.70163e-20 $X=7.675 $Y=1.98
c227 39 0 1.8278e-19 $X=3.56 $Y=0.95
c228 32 0 4.70822e-20 $X=10.96 $Y=1.26
c229 12 0 3.05941e-20 $X=9.51 $Y=0.445
r230 77 78 7.90164 $w=3.05e-07 $l=5e-08 $layer=POLY_cond $X=9.87 $Y=1.2 $X2=9.92
+ $Y2=1.2
r231 73 74 8.63679 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=8.885 $Y=1.255
+ $X2=9.055 $Y2=1.255
r232 68 70 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=3.385 $Y=1.7
+ $X2=3.645 $Y2=1.7
r233 65 66 7.3123 $w=3.17e-07 $l=1.9e-07 $layer=LI1_cond $X=2.57 $Y=0.76
+ $X2=2.57 $Y2=0.95
r234 62 77 42.6689 $w=3.05e-07 $l=2.7e-07 $layer=POLY_cond $X=9.6 $Y=1.2
+ $X2=9.87 $Y2=1.2
r235 62 75 14.223 $w=3.05e-07 $l=9e-08 $layer=POLY_cond $X=9.6 $Y=1.2 $X2=9.51
+ $Y2=1.2
r236 61 74 19.0328 $w=3.28e-07 $l=5.45e-07 $layer=LI1_cond $X=9.6 $Y=1.2
+ $X2=9.055 $Y2=1.2
r237 61 62 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.6
+ $Y=1.2 $X2=9.6 $Y2=1.2
r238 58 73 73.3957 $w=1.68e-07 $l=1.125e-06 $layer=LI1_cond $X=7.76 $Y=1.39
+ $X2=8.885 $Y2=1.39
r239 56 72 2.88756 $w=3.3e-07 $l=1.9799e-07 $layer=LI1_cond $X=7.675 $Y=1.98
+ $X2=7.515 $Y2=2.065
r240 55 58 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.675 $Y=1.475
+ $X2=7.76 $Y2=1.39
r241 55 56 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=7.675 $Y=1.475
+ $X2=7.675 $Y2=1.98
r242 51 72 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.515 $Y=2.15
+ $X2=7.515 $Y2=2.065
r243 51 53 6.22449 $w=4.88e-07 $l=2.55e-07 $layer=LI1_cond $X=7.515 $Y=2.15
+ $X2=7.515 $Y2=2.405
r244 49 72 3.80956 $w=1.7e-07 $l=2.45e-07 $layer=LI1_cond $X=7.27 $Y=2.065
+ $X2=7.515 $Y2=2.065
r245 49 50 185.283 $w=1.68e-07 $l=2.84e-06 $layer=LI1_cond $X=7.27 $Y=2.065
+ $X2=4.43 $Y2=2.065
r246 47 50 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.345 $Y=2.15
+ $X2=4.43 $Y2=2.065
r247 47 48 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=4.345 $Y=2.15
+ $X2=4.345 $Y2=2.295
r248 46 70 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.645 $Y=1.615
+ $X2=3.645 $Y2=1.7
r249 45 46 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=3.645 $Y=1.035
+ $X2=3.645 $Y2=1.615
r250 43 48 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.26 $Y=2.38
+ $X2=4.345 $Y2=2.295
r251 43 44 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=4.26 $Y=2.38
+ $X2=3.47 $Y2=2.38
r252 42 44 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.385 $Y=2.295
+ $X2=3.47 $Y2=2.38
r253 41 68 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.385 $Y=1.785
+ $X2=3.385 $Y2=1.7
r254 41 42 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=3.385 $Y=1.785
+ $X2=3.385 $Y2=2.295
r255 40 66 4.38581 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=2.78 $Y=0.95
+ $X2=2.57 $Y2=0.95
r256 39 45 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.56 $Y=0.95
+ $X2=3.645 $Y2=1.035
r257 39 40 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=3.56 $Y=0.95
+ $X2=2.78 $Y2=0.95
r258 37 66 3.46775 $w=3.17e-07 $l=1.14782e-07 $layer=LI1_cond $X=2.64 $Y=1.035
+ $X2=2.57 $Y2=0.95
r259 37 67 56.799 $w=2.78e-07 $l=1.38e-06 $layer=LI1_cond $X=2.64 $Y=1.035
+ $X2=2.64 $Y2=2.415
r260 33 67 6.05995 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=2.615 $Y=2.58
+ $X2=2.615 $Y2=2.415
r261 33 35 5.76222 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=2.615 $Y=2.58
+ $X2=2.615 $Y2=2.745
r262 28 32 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=10.96 $Y=1.335
+ $X2=10.96 $Y2=1.26
r263 28 30 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=10.96 $Y=1.335
+ $X2=10.96 $Y2=2.155
r264 24 32 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=10.96 $Y=1.185
+ $X2=10.96 $Y2=1.26
r265 24 26 358.936 $w=1.5e-07 $l=7e-07 $layer=POLY_cond $X=10.96 $Y=1.185
+ $X2=10.96 $Y2=0.485
r266 23 78 32.2155 $w=3.05e-07 $l=1.52069e-07 $layer=POLY_cond $X=10.045 $Y=1.26
+ $X2=9.92 $Y2=1.2
r267 22 32 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=10.885 $Y=1.26
+ $X2=10.96 $Y2=1.26
r268 22 23 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=10.885 $Y=1.26
+ $X2=10.045 $Y2=1.26
r269 18 78 7.52206 $w=2.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.92 $Y=1.365
+ $X2=9.92 $Y2=1.2
r270 18 20 305.598 $w=2.5e-07 $l=1.23e-06 $layer=POLY_cond $X=9.92 $Y=1.365
+ $X2=9.92 $Y2=2.595
r271 14 77 19.3576 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.87 $Y=1.035
+ $X2=9.87 $Y2=1.2
r272 14 16 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=9.87 $Y=1.035
+ $X2=9.87 $Y2=0.445
r273 10 75 19.3576 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.51 $Y=1.035
+ $X2=9.51 $Y2=1.2
r274 10 12 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=9.51 $Y=1.035
+ $X2=9.51 $Y2=0.445
r275 3 53 600 $w=1.7e-07 $l=3.75566e-07 $layer=licon1_PDIFF $count=1 $X=7.29
+ $Y=2.095 $X2=7.435 $Y2=2.405
r276 2 35 600 $w=1.7e-07 $l=3.73497e-07 $layer=licon1_PDIFF $count=1 $X=2.475
+ $Y=2.435 $X2=2.615 $Y2=2.745
r277 1 65 182 $w=1.7e-07 $l=3.81772e-07 $layer=licon1_NDIFF $count=1 $X=2.19
+ $Y=0.485 $X2=2.445 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_LP__SRDLRTP_1%A_2120_55# 1 2 9 13 17 21 25 26 28
c50 28 0 4.70822e-20 $X=10.745 $Y=1.48
c51 21 0 1.20584e-19 $X=10.745 $Y=1.98
r52 26 31 46.255 $w=3.35e-07 $l=1.65e-07 $layer=POLY_cond $X=11.412 $Y=1.48
+ $X2=11.412 $Y2=1.645
r53 26 30 46.255 $w=3.35e-07 $l=1.65e-07 $layer=POLY_cond $X=11.412 $Y=1.48
+ $X2=11.412 $Y2=1.315
r54 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.41
+ $Y=1.48 $X2=11.41 $Y2=1.48
r55 23 28 1.34256 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=10.91 $Y=1.48
+ $X2=10.745 $Y2=1.48
r56 23 25 17.4613 $w=3.28e-07 $l=5e-07 $layer=LI1_cond $X=10.91 $Y=1.48
+ $X2=11.41 $Y2=1.48
r57 19 28 5.16603 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=10.745 $Y=1.645
+ $X2=10.745 $Y2=1.48
r58 19 21 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=10.745 $Y=1.645
+ $X2=10.745 $Y2=1.98
r59 15 28 5.16603 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=10.745 $Y=1.315
+ $X2=10.745 $Y2=1.48
r60 15 17 28.9857 $w=3.28e-07 $l=8.3e-07 $layer=LI1_cond $X=10.745 $Y=1.315
+ $X2=10.745 $Y2=0.485
r61 13 31 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=11.505 $Y=2.465
+ $X2=11.505 $Y2=1.645
r62 9 30 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=11.505 $Y=0.695
+ $X2=11.505 $Y2=1.315
r63 2 21 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=10.6
+ $Y=1.835 $X2=10.745 $Y2=1.98
r64 1 17 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=10.6
+ $Y=0.275 $X2=10.745 $Y2=0.485
.ends

.subckt PM_SKY130_FD_SC_LP__SRDLRTP_1%VPWR 1 2 3 4 13 15 17 21 25 29 31 39 46 47
+ 53 56 63
r120 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.28 $Y=3.33
+ $X2=11.28 $Y2=3.33
r121 59 60 1.32857 $w=1.7e-07 $l=1.19e-06 $layer=mcon $count=7 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r122 56 59 9.42908 $w=3.28e-07 $l=2.7e-07 $layer=LI1_cond $X=4.465 $Y=3.06
+ $X2=4.465 $Y2=3.33
r123 53 54 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r124 51 54 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.2 $Y2=3.33
r125 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r126 47 64 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.76 $Y=3.33
+ $X2=11.28 $Y2=3.33
r127 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.76 $Y=3.33
+ $X2=11.76 $Y2=3.33
r128 44 63 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=11.375 $Y=3.33
+ $X2=11.25 $Y2=3.33
r129 44 46 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=11.375 $Y=3.33
+ $X2=11.76 $Y2=3.33
r130 43 64 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.8 $Y=3.33
+ $X2=11.28 $Y2=3.33
r131 42 43 1.32857 $w=1.7e-07 $l=1.19e-06 $layer=mcon $count=7 $X=10.8 $Y=3.33
+ $X2=10.8 $Y2=3.33
r132 40 59 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.63 $Y=3.33
+ $X2=4.465 $Y2=3.33
r133 40 42 402.535 $w=1.68e-07 $l=6.17e-06 $layer=LI1_cond $X=4.63 $Y=3.33
+ $X2=10.8 $Y2=3.33
r134 39 63 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=11.125 $Y=3.33
+ $X2=11.25 $Y2=3.33
r135 39 42 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=11.125 $Y=3.33
+ $X2=10.8 $Y2=3.33
r136 38 60 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r137 37 38 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r138 35 38 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=4.08 $Y2=3.33
r139 35 54 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r140 34 37 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=1.68 $Y=3.33
+ $X2=4.08 $Y2=3.33
r141 34 35 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r142 32 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.49 $Y=3.33
+ $X2=1.325 $Y2=3.33
r143 32 34 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=1.49 $Y=3.33
+ $X2=1.68 $Y2=3.33
r144 31 59 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.3 $Y=3.33
+ $X2=4.465 $Y2=3.33
r145 31 37 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=4.3 $Y=3.33
+ $X2=4.08 $Y2=3.33
r146 29 43 1.33793 $w=4.9e-07 $l=4.8e-06 $layer=MET1_cond $X=6 $Y=3.33 $X2=10.8
+ $Y2=3.33
r147 29 60 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=6 $Y=3.33
+ $X2=4.56 $Y2=3.33
r148 25 28 22.3574 $w=2.48e-07 $l=4.85e-07 $layer=LI1_cond $X=11.25 $Y=1.98
+ $X2=11.25 $Y2=2.465
r149 23 63 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=11.25 $Y=3.245
+ $X2=11.25 $Y2=3.33
r150 23 28 35.9562 $w=2.48e-07 $l=7.8e-07 $layer=LI1_cond $X=11.25 $Y=3.245
+ $X2=11.25 $Y2=2.465
r151 19 53 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.325 $Y=3.245
+ $X2=1.325 $Y2=3.33
r152 19 21 22.8742 $w=3.28e-07 $l=6.55e-07 $layer=LI1_cond $X=1.325 $Y=3.245
+ $X2=1.325 $Y2=2.59
r153 18 50 4.73185 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=3.33
+ $X2=0.222 $Y2=3.33
r154 17 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.16 $Y=3.33
+ $X2=1.325 $Y2=3.33
r155 17 18 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=1.16 $Y=3.33
+ $X2=0.445 $Y2=3.33
r156 13 50 3.03433 $w=3.3e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.222 $Y2=3.33
r157 13 15 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.28 $Y2=2.93
r158 4 28 300 $w=1.7e-07 $l=7.46693e-07 $layer=licon1_PDIFF $count=2 $X=11.035
+ $Y=1.835 $X2=11.29 $Y2=2.465
r159 4 25 600 $w=1.7e-07 $l=3.19374e-07 $layer=licon1_PDIFF $count=1 $X=11.035
+ $Y=1.835 $X2=11.29 $Y2=1.98
r160 3 56 600 $w=1.7e-07 $l=1.24599e-06 $layer=licon1_PDIFF $count=1 $X=4.21
+ $Y=1.935 $X2=4.465 $Y2=3.06
r161 2 21 300 $w=1.7e-07 $l=3.23342e-07 $layer=licon1_PDIFF $count=2 $X=1.07
+ $Y=2.435 $X2=1.325 $Y2=2.59
r162 1 15 600 $w=1.7e-07 $l=5.6285e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.435 $X2=0.28 $Y2=2.93
.ends

.subckt PM_SKY130_FD_SC_LP__SRDLRTP_1%A_280_97# 1 2 9 11 16 18
r45 14 16 6.21713 $w=3.78e-07 $l=2.05e-07 $layer=LI1_cond $X=1.54 $Y=0.655
+ $X2=1.745 $Y2=0.655
r46 9 18 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=1.825 $Y=2.58
+ $X2=1.825 $Y2=2.415
r47 9 11 5.76222 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=1.825 $Y=2.58
+ $X2=1.825 $Y2=2.745
r48 7 16 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.745 $Y=0.845
+ $X2=1.745 $Y2=0.655
r49 7 18 102.428 $w=1.68e-07 $l=1.57e-06 $layer=LI1_cond $X=1.745 $Y=0.845
+ $X2=1.745 $Y2=2.415
r50 2 11 600 $w=1.7e-07 $l=3.73497e-07 $layer=licon1_PDIFF $count=1 $X=1.685
+ $Y=2.435 $X2=1.825 $Y2=2.745
r51 1 14 182 $w=1.7e-07 $l=2.29565e-07 $layer=licon1_NDIFF $count=1 $X=1.4
+ $Y=0.485 $X2=1.54 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__SRDLRTP_1%KAPWR 1 2 3 4 13 19 27 30 36 39
r103 36 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.32 $Y=2.82
+ $X2=10.32 $Y2=2.82
r104 31 39 1.04938 $w=2.7e-07 $l=1.92e-06 $layer=MET1_cond $X=8.4 $Y=2.81
+ $X2=10.32 $Y2=2.81
r105 30 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=2.82 $X2=8.4
+ $Y2=2.82
r106 23 27 8.03218 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=6 $Y=2.825 $X2=6.23
+ $Y2=2.825
r107 19 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=2.82
+ $X2=5.52 $Y2=2.82
r108 16 19 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=5.025 $Y=2.825
+ $X2=5.52 $Y2=2.825
r109 13 31 1.31172 $w=2.7e-07 $l=2.4e-06 $layer=MET1_cond $X=6 $Y=2.81 $X2=8.4
+ $Y2=2.81
r110 13 20 0.262345 $w=2.7e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=2.81 $X2=5.52
+ $Y2=2.81
r111 13 23 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=2.82 $X2=6
+ $Y2=2.82
r112 4 36 600 $w=1.7e-07 $l=8.37078e-07 $layer=licon1_PDIFF $count=1 $X=10.045
+ $Y=2.095 $X2=10.185 $Y2=2.865
r113 3 30 600 $w=1.7e-07 $l=8.41665e-07 $layer=licon1_PDIFF $count=1 $X=8.285
+ $Y=2.095 $X2=8.435 $Y2=2.865
r114 2 27 600 $w=1.7e-07 $l=6.09303e-07 $layer=licon1_PDIFF $count=1 $X=5.975
+ $Y=2.33 $X2=6.23 $Y2=2.825
r115 1 16 600 $w=1.7e-07 $l=5.6285e-07 $layer=licon1_PDIFF $count=1 $X=4.88
+ $Y=2.33 $X2=5.025 $Y2=2.825
.ends

.subckt PM_SKY130_FD_SC_LP__SRDLRTP_1%Q 1 2 9 14 15 16 17 23 29
r24 21 29 0.960369 $w=3.58e-07 $l=3e-08 $layer=LI1_cond $X=11.735 $Y=0.955
+ $X2=11.735 $Y2=0.925
r25 17 31 8.12688 $w=3.58e-07 $l=1.53e-07 $layer=LI1_cond $X=11.735 $Y=0.982
+ $X2=11.735 $Y2=1.135
r26 17 21 0.864332 $w=3.58e-07 $l=2.7e-08 $layer=LI1_cond $X=11.735 $Y=0.982
+ $X2=11.735 $Y2=0.955
r27 17 29 0.896345 $w=3.58e-07 $l=2.8e-08 $layer=LI1_cond $X=11.735 $Y=0.897
+ $X2=11.735 $Y2=0.925
r28 16 17 10.9482 $w=3.58e-07 $l=3.42e-07 $layer=LI1_cond $X=11.735 $Y=0.555
+ $X2=11.735 $Y2=0.897
r29 16 23 4.32166 $w=3.58e-07 $l=1.35e-07 $layer=LI1_cond $X=11.735 $Y=0.555
+ $X2=11.735 $Y2=0.42
r30 15 31 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=11.83 $Y=1.815
+ $X2=11.83 $Y2=1.135
r31 14 15 8.51103 $w=3.58e-07 $l=1.65e-07 $layer=LI1_cond $X=11.735 $Y=1.98
+ $X2=11.735 $Y2=1.815
r32 7 14 0.480185 $w=3.58e-07 $l=1.5e-08 $layer=LI1_cond $X=11.735 $Y=1.995
+ $X2=11.735 $Y2=1.98
r33 7 9 29.2913 $w=3.58e-07 $l=9.15e-07 $layer=LI1_cond $X=11.735 $Y=1.995
+ $X2=11.735 $Y2=2.91
r34 2 14 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=11.58
+ $Y=1.835 $X2=11.72 $Y2=1.98
r35 2 9 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=11.58
+ $Y=1.835 $X2=11.72 $Y2=2.91
r36 1 23 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=11.58
+ $Y=0.275 $X2=11.72 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__SRDLRTP_1%VGND 1 2 3 4 5 18 22 26 31 32 33 34 41 42
+ 43 61 68 75 76 80 86
c122 76 0 3.39925e-20 $X=11.76 $Y=0
r123 86 87 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.28 $Y=0
+ $X2=11.28 $Y2=0
r124 80 83 9.7783 $w=3.28e-07 $l=2.8e-07 $layer=LI1_cond $X=8.775 $Y=0 $X2=8.775
+ $Y2=0.28
r125 80 81 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=8.88 $Y=0
+ $X2=8.88 $Y2=0
r126 76 87 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.76 $Y=0
+ $X2=11.28 $Y2=0
r127 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.76 $Y=0
+ $X2=11.76 $Y2=0
r128 73 86 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=11.375 $Y=0
+ $X2=11.25 $Y2=0
r129 73 75 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=11.375 $Y=0
+ $X2=11.76 $Y2=0
r130 72 87 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.8 $Y=0
+ $X2=11.28 $Y2=0
r131 72 81 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=10.8 $Y=0
+ $X2=8.88 $Y2=0
r132 71 72 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=10.8 $Y=0
+ $X2=10.8 $Y2=0
r133 69 80 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.94 $Y=0 $X2=8.775
+ $Y2=0
r134 69 71 121.348 $w=1.68e-07 $l=1.86e-06 $layer=LI1_cond $X=8.94 $Y=0 $X2=10.8
+ $Y2=0
r135 68 86 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=11.125 $Y=0
+ $X2=11.25 $Y2=0
r136 68 71 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=11.125 $Y=0
+ $X2=10.8 $Y2=0
r137 67 81 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=0 $X2=8.88
+ $Y2=0
r138 66 67 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r139 64 67 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=6.48 $Y=0 $X2=8.4
+ $Y2=0
r140 63 66 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=6.48 $Y=0 $X2=8.4
+ $Y2=0
r141 63 64 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.48 $Y=0
+ $X2=6.48 $Y2=0
r142 61 80 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.61 $Y=0 $X2=8.775
+ $Y2=0
r143 61 66 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=8.61 $Y=0 $X2=8.4
+ $Y2=0
r144 56 59 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=4.08 $Y=0 $X2=6
+ $Y2=0
r145 56 57 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.08 $Y=0
+ $X2=4.08 $Y2=0
r146 54 57 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r147 53 54 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r148 51 54 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=1.2 $Y=0 $X2=3.6
+ $Y2=0
r149 50 53 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=3.6
+ $Y2=0
r150 50 51 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r151 47 51 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r152 46 47 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r153 43 64 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.48
+ $Y2=0
r154 43 57 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=6 $Y=0 $X2=4.08
+ $Y2=0
r155 43 59 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6 $Y=0 $X2=6
+ $Y2=0
r156 42 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.315 $Y=0 $X2=6.48
+ $Y2=0
r157 41 59 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=6.15 $Y=0 $X2=6
+ $Y2=0
r158 41 42 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.15 $Y=0 $X2=6.315
+ $Y2=0
r159 36 56 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=3.99 $Y=0 $X2=4.08
+ $Y2=0
r160 34 53 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=3.66 $Y=0 $X2=3.6
+ $Y2=0
r161 33 38 9.42908 $w=3.28e-07 $l=2.7e-07 $layer=LI1_cond $X=3.825 $Y=0
+ $X2=3.825 $Y2=0.27
r162 33 36 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.825 $Y=0 $X2=3.99
+ $Y2=0
r163 33 34 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.825 $Y=0 $X2=3.66
+ $Y2=0
r164 31 46 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=0.945 $Y=0
+ $X2=0.72 $Y2=0
r165 31 32 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.945 $Y=0 $X2=1.07
+ $Y2=0
r166 30 50 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=1.195 $Y=0 $X2=1.2
+ $Y2=0
r167 30 32 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.195 $Y=0 $X2=1.07
+ $Y2=0
r168 26 28 17.5171 $w=2.48e-07 $l=3.8e-07 $layer=LI1_cond $X=11.25 $Y=0.42
+ $X2=11.25 $Y2=0.8
r169 24 86 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=11.25 $Y=0.085
+ $X2=11.25 $Y2=0
r170 24 26 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=11.25 $Y=0.085
+ $X2=11.25 $Y2=0.42
r171 20 42 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.315 $Y=0.085
+ $X2=6.315 $Y2=0
r172 20 22 13.2706 $w=3.28e-07 $l=3.8e-07 $layer=LI1_cond $X=6.315 $Y=0.085
+ $X2=6.315 $Y2=0.465
r173 16 32 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.07 $Y=0.085
+ $X2=1.07 $Y2=0
r174 16 18 26.2757 $w=2.48e-07 $l=5.7e-07 $layer=LI1_cond $X=1.07 $Y=0.085
+ $X2=1.07 $Y2=0.655
r175 5 28 182 $w=1.7e-07 $l=6.39922e-07 $layer=licon1_NDIFF $count=1 $X=11.035
+ $Y=0.275 $X2=11.29 $Y2=0.8
r176 5 26 182 $w=1.7e-07 $l=3.19374e-07 $layer=licon1_NDIFF $count=1 $X=11.035
+ $Y=0.275 $X2=11.29 $Y2=0.42
r177 4 83 182 $w=1.7e-07 $l=2.41454e-07 $layer=licon1_NDIFF $count=1 $X=8.555
+ $Y=0.235 $X2=8.775 $Y2=0.28
r178 3 22 182 $w=1.7e-07 $l=2.29783e-07 $layer=licon1_NDIFF $count=1 $X=6.095
+ $Y=0.485 $X2=6.315 $Y2=0.465
r179 2 38 182 $w=1.7e-07 $l=3.46194e-07 $layer=licon1_NDIFF $count=1 $X=3.57
+ $Y=0.485 $X2=3.825 $Y2=0.27
r180 1 18 182 $w=1.7e-07 $l=2.50998e-07 $layer=licon1_NDIFF $count=1 $X=0.93
+ $Y=0.485 $X2=1.11 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__SRDLRTP_1%A_1624_47# 1 2 9 11 12 14
c38 11 0 3.05941e-20 $X=9.125 $Y=0.62
r39 14 16 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=9.29 $Y=0.465
+ $X2=9.29 $Y2=0.62
r40 11 16 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.125 $Y=0.62
+ $X2=9.29 $Y2=0.62
r41 11 12 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=9.125 $Y=0.62
+ $X2=8.43 $Y2=0.62
r42 7 12 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=8.305 $Y=0.535
+ $X2=8.43 $Y2=0.62
r43 7 9 3.22684 $w=2.48e-07 $l=7e-08 $layer=LI1_cond $X=8.305 $Y=0.535 $X2=8.305
+ $Y2=0.465
r44 2 14 182 $w=1.7e-07 $l=2.93684e-07 $layer=licon1_NDIFF $count=1 $X=9.145
+ $Y=0.235 $X2=9.29 $Y2=0.465
r45 1 9 182 $w=1.7e-07 $l=2.93684e-07 $layer=licon1_NDIFF $count=1 $X=8.12
+ $Y=0.235 $X2=8.265 $Y2=0.465
.ends

