* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__sdfstp_4 CLK D SCD SCE SET_B VGND VNB VPB VPWR Q
M1000 VGND a_346_93# a_304_119# VNB nshort w=420000u l=150000u
+  ad=1.7677e+12p pd=1.701e+07u as=8.82e+10p ps=1.26e+06u
M1001 a_346_93# SCE VGND VNB nshort w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1002 a_1751_379# a_773_409# a_1960_125# VPB phighvt w=840000u l=150000u
+  ad=4.452e+11p pd=4.42e+06u as=3.801e+11p ps=3.8e+06u
M1003 a_1960_125# SET_B VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=2.5593e+12p ps=2.281e+07u
M1004 VGND a_2638_53# Q VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=4.704e+11p ps=4.48e+06u
M1005 a_961_491# a_773_409# VGND VNB nshort w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1006 VPWR a_2638_53# Q VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=7.056e+11p ps=6.16e+06u
M1007 VGND a_1960_125# a_2638_53# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=2.226e+11p ps=2.21e+06u
M1008 a_1315_81# a_961_491# a_1211_463# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=1.176e+11p ps=1.4e+06u
M1009 a_218_119# SCE a_146_119# VNB nshort w=420000u l=150000u
+  ad=3.843e+11p pd=3.51e+06u as=8.82e+10p ps=1.26e+06u
M1010 a_1751_379# a_1211_463# VPWR VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND a_1339_331# a_1315_81# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_196_479# SCE VPWR VPB phighvt w=640000u l=150000u
+  ad=1.344e+11p pd=1.7e+06u as=0p ps=0u
M1013 a_304_119# D a_218_119# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_146_119# SCD VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_2205_231# a_1960_125# VPWR VPB phighvt w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1016 a_2248_125# a_2205_231# a_2163_125# VNB nshort w=420000u l=150000u
+  ad=1.365e+11p pd=1.49e+06u as=1.155e+11p ps=1.39e+06u
M1017 a_218_119# D a_196_479# VPB phighvt w=640000u l=150000u
+  ad=4.743e+11p pd=3.97e+06u as=0p ps=0u
M1018 VPWR SET_B a_1339_331# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.344e+11p ps=1.48e+06u
M1019 VPWR a_2205_231# a_1858_463# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=3e+11p ps=3.23e+06u
M1020 a_2163_125# a_773_409# a_1960_125# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=5.294e+11p ps=3.01e+06u
M1021 Q a_2638_53# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_1297_463# a_773_409# a_1211_463# VPB phighvt w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=1.176e+11p ps=1.4e+06u
M1023 a_961_491# a_773_409# VPWR VPB phighvt w=640000u l=150000u
+  ad=1.696e+11p pd=1.81e+06u as=0p ps=0u
M1024 VGND SET_B a_2248_125# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 VPWR a_1339_331# a_1297_463# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_1960_125# a_961_491# a_1858_463# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_1598_125# a_1211_463# a_1339_331# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=1.113e+11p ps=1.37e+06u
M1028 a_1888_125# a_1211_463# VGND VNB nshort w=640000u l=150000u
+  ad=1.344e+11p pd=1.7e+06u as=0p ps=0u
M1029 a_1339_331# a_1211_463# VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 Q a_2638_53# VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_27_479# a_346_93# a_218_119# VPB phighvt w=640000u l=150000u
+  ad=3.392e+11p pd=3.62e+06u as=0p ps=0u
M1032 VGND SET_B a_1598_125# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 a_1211_463# a_961_491# a_218_119# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1034 Q a_2638_53# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1035 a_1960_125# a_961_491# a_1888_125# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1036 Q a_2638_53# VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1037 VGND CLK a_773_409# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1038 VPWR SCD a_27_479# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1039 a_346_93# SCE VPWR VPB phighvt w=640000u l=150000u
+  ad=1.696e+11p pd=1.81e+06u as=0p ps=0u
M1040 VPWR a_1960_125# a_2638_53# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=3.339e+11p ps=3.05e+06u
M1041 a_1211_463# a_773_409# a_218_119# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1042 VPWR CLK a_773_409# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=3.329e+11p ps=2.82e+06u
M1043 a_2205_231# a_1960_125# VGND VNB nshort w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1044 VPWR a_2638_53# Q VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1045 VGND a_2638_53# Q VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
