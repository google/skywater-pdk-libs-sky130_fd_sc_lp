* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__a211o_0 A1 A2 B1 C1 VGND VNB VPB VPWR X
X0 X a_80_172# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 a_265_60# A1 a_80_172# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 VGND A2 a_265_60# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 X a_80_172# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X4 a_80_172# B1 VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 VPWR A1 a_224_482# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X6 a_224_482# B1 a_487_482# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X7 a_487_482# C1 a_80_172# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X8 VGND C1 a_80_172# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 a_224_482# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
.ends
