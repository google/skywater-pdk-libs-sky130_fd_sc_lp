* File: sky130_fd_sc_lp__dfsbp_lp.spice
* Created: Wed Sep  2 09:44:14 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__dfsbp_lp.pex.spice"
.subckt sky130_fd_sc_lp__dfsbp_lp  VNB VPB D CLK SET_B VPWR Q_N Q VGND
* 
* VGND	VGND
* Q	Q
* Q_N	Q_N
* VPWR	VPWR
* SET_B	SET_B
* CLK	CLK
* D	D
* VPB	VPB
* VNB	VNB
MM1019 A_110_57# N_D_M1019_g N_VGND_M1019_s VNB NSHORT L=0.15 W=0.42 AD=0.0441
+ AS=0.1113 PD=0.63 PS=1.37 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1010 N_A_145_409#_M1010_d N_D_M1010_g A_110_57# VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.0441 PD=1.37 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1036 A_373_113# N_CLK_M1036_g N_A_263_409#_M1036_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1134 PD=0.63 PS=1.38 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.3 A=0.063 P=1.14 MULT=1
MM1024 N_VGND_M1024_d N_CLK_M1024_g A_373_113# VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1028 A_531_113# N_A_263_409#_M1028_g N_VGND_M1024_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75001
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1021 N_A_476_409#_M1021_d N_A_263_409#_M1021_g A_531_113# VNB NSHORT L=0.15
+ W=0.42 AD=0.1113 AS=0.0441 PD=1.37 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8
+ SA=75001.3 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1020 N_A_712_419#_M1020_d N_A_263_409#_M1020_g N_A_145_409#_M1020_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.108 AS=0.1113 PD=1.005 PS=1.37 NRD=18.564 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1017 A_904_125# N_A_476_409#_M1017_g N_A_712_419#_M1020_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.108 PD=0.63 PS=1.005 NRD=14.28 NRS=17.136 M=1 R=2.8
+ SA=75000.5 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1008 N_VGND_M1008_d N_A_946_99#_M1008_g A_904_125# VNB NSHORT L=0.15 W=0.42
+ AD=0.2124 AS=0.0441 PD=2.03 PS=0.63 NRD=128.772 NRS=14.28 M=1 R=2.8 SA=75000.9
+ SB=75000.3 A=0.063 P=1.14 MULT=1
MM1034 A_1249_125# N_A_712_419#_M1034_g N_A_946_99#_M1034_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0504 AS=0.1197 PD=0.66 PS=1.41 NRD=18.564 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75002.3 A=0.063 P=1.14 MULT=1
MM1022 N_VGND_M1022_d N_SET_B_M1022_g A_1249_125# VNB NSHORT L=0.15 W=0.42
+ AD=0.0882 AS=0.0504 PD=0.84 PS=0.66 NRD=39.996 NRS=18.564 M=1 R=2.8 SA=75000.6
+ SB=75001.9 A=0.063 P=1.14 MULT=1
MM1029 A_1441_125# N_A_712_419#_M1029_g N_VGND_M1022_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.0882 PD=0.66 PS=0.84 NRD=18.564 NRS=0 M=1 R=2.8 SA=75001.2
+ SB=75001.3 A=0.063 P=1.14 MULT=1
MM1009 N_A_1519_125#_M1009_d N_A_476_409#_M1009_g A_1441_125# VNB NSHORT L=0.15
+ W=0.42 AD=0.0756 AS=0.0504 PD=0.78 PS=0.66 NRD=22.848 NRS=18.564 M=1 R=2.8
+ SA=75001.6 SB=75001 A=0.063 P=1.14 MULT=1
MM1000 A_1621_125# N_A_263_409#_M1000_g N_A_1519_125#_M1009_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0940625 AS=0.0756 PD=1.04 PS=0.78 NRD=48.264 NRS=0 M=1 R=2.8
+ SA=75002.1 SB=75000.4 A=0.063 P=1.14 MULT=1
MM1039 A_1716_66# N_A_1686_40#_M1039_g A_1621_125# VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.0940625 PD=0.66 PS=1.04 NRD=18.564 NRS=48.264 M=1 R=2.8
+ SA=75000.9 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1037 N_VGND_M1037_d N_SET_B_M1037_g A_1716_66# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0504 PD=1.41 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75001.3
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1006 A_2042_57# N_A_1519_125#_M1006_g N_A_1686_40#_M1006_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.1197 PD=0.63 PS=1.41 NRD=14.28 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.4 A=0.063 P=1.14 MULT=1
MM1035 N_VGND_M1035_d N_A_1519_125#_M1035_g A_2042_57# VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1011 A_2200_57# N_A_1519_125#_M1011_g N_VGND_M1035_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75001
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1012 N_Q_N_M1012_d N_A_1519_125#_M1012_g A_2200_57# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.4
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1023 A_2470_57# N_A_1519_125#_M1023_g N_A_2383_57#_M1023_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.1197 PD=0.63 PS=1.41 NRD=14.28 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.4 A=0.063 P=1.14 MULT=1
MM1025 N_VGND_M1025_d N_A_1519_125#_M1025_g A_2470_57# VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1040 A_2628_57# N_A_2383_57#_M1040_g N_VGND_M1025_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75001
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1031 N_Q_M1031_d N_A_2383_57#_M1031_g A_2628_57# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.4
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1002 N_A_145_409#_M1002_d N_D_M1002_g N_VPWR_M1002_s VPB PHIGHVT L=0.25 W=1
+ AD=0.285 AS=0.285 PD=2.57 PS=2.57 NRD=0 NRS=0 M=1 R=4 SA=125000 SB=125000
+ A=0.25 P=2.5 MULT=1
MM1001 N_VPWR_M1001_d N_CLK_M1001_g N_A_263_409#_M1001_s VPB PHIGHVT L=0.25 W=1
+ AD=0.14 AS=0.285 PD=1.28 PS=2.57 NRD=0 NRS=0 M=1 R=4 SA=125000 SB=125001
+ A=0.25 P=2.5 MULT=1
MM1026 N_A_476_409#_M1026_d N_A_263_409#_M1026_g N_VPWR_M1001_d VPB PHIGHVT
+ L=0.25 W=1 AD=0.285 AS=0.14 PD=2.57 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125001
+ SB=125000 A=0.25 P=2.5 MULT=1
MM1005 N_A_712_419#_M1005_d N_A_476_409#_M1005_g N_A_145_409#_M1005_s VPB
+ PHIGHVT L=0.25 W=1 AD=0.305 AS=0.285 PD=1.61 PS=2.57 NRD=65.01 NRS=0 M=1 R=4
+ SA=125000 SB=125006 A=0.25 P=2.5 MULT=1
MM1016 A_884_419# N_A_263_409#_M1016_g N_A_712_419#_M1005_d VPB PHIGHVT L=0.25
+ W=1 AD=0.17 AS=0.305 PD=1.34 PS=1.61 NRD=22.6353 NRS=0 M=1 R=4 SA=125001
+ SB=125006 A=0.25 P=2.5 MULT=1
MM1032 N_VPWR_M1032_d N_A_946_99#_M1032_g A_884_419# VPB PHIGHVT L=0.25 W=1
+ AD=0.325 AS=0.17 PD=1.65 PS=1.34 NRD=0 NRS=22.6353 M=1 R=4 SA=125002 SB=125005
+ A=0.25 P=2.5 MULT=1
MM1003 N_A_946_99#_M1003_d N_A_712_419#_M1003_g N_VPWR_M1032_d VPB PHIGHVT
+ L=0.25 W=1 AD=0.14 AS=0.325 PD=1.28 PS=1.65 NRD=0 NRS=72.8703 M=1 R=4
+ SA=125003 SB=125004 A=0.25 P=2.5 MULT=1
MM1027 N_VPWR_M1027_d N_SET_B_M1027_g N_A_946_99#_M1003_d VPB PHIGHVT L=0.25 W=1
+ AD=0.26765 AS=0.14 PD=1.585 PS=1.28 NRD=16.7253 NRS=0 M=1 R=4 SA=125003
+ SB=125004 A=0.25 P=2.5 MULT=1
MM1018 A_1441_419# N_A_712_419#_M1018_g N_VPWR_M1027_d VPB PHIGHVT L=0.25 W=1
+ AD=0.12 AS=0.26765 PD=1.24 PS=1.585 NRD=12.7853 NRS=31.5003 M=1 R=4 SA=125004
+ SB=125003 A=0.25 P=2.5 MULT=1
MM1038 N_A_1519_125#_M1038_d N_A_263_409#_M1038_g A_1441_419# VPB PHIGHVT L=0.25
+ W=1 AD=0.325 AS=0.12 PD=1.65 PS=1.24 NRD=26.5753 NRS=12.7853 M=1 R=4 SA=125004
+ SB=125002 A=0.25 P=2.5 MULT=1
MM1015 A_1719_419# N_A_476_409#_M1015_g N_A_1519_125#_M1038_d VPB PHIGHVT L=0.25
+ W=1 AD=0.145 AS=0.325 PD=1.29 PS=1.65 NRD=17.7103 NRS=46.2753 M=1 R=4
+ SA=125005 SB=125001 A=0.25 P=2.5 MULT=1
MM1033 N_VPWR_M1033_d N_A_1686_40#_M1033_g A_1719_419# VPB PHIGHVT L=0.25 W=1
+ AD=0.225 AS=0.145 PD=1.45 PS=1.29 NRD=0 NRS=17.7103 M=1 R=4 SA=125006
+ SB=125001 A=0.25 P=2.5 MULT=1
MM1013 N_A_1519_125#_M1013_d N_SET_B_M1013_g N_VPWR_M1033_d VPB PHIGHVT L=0.25
+ W=1 AD=0.28 AS=0.225 PD=2.56 PS=1.45 NRD=0 NRS=33.4703 M=1 R=4 SA=125006
+ SB=125000 A=0.25 P=2.5 MULT=1
MM1007 N_VPWR_M1007_d N_A_1519_125#_M1007_g N_A_1686_40#_M1007_s VPB PHIGHVT
+ L=0.25 W=1 AD=0.225 AS=0.285 PD=1.45 PS=2.57 NRD=33.4703 NRS=0 M=1 R=4
+ SA=125000 SB=125001 A=0.25 P=2.5 MULT=1
MM1014 N_Q_N_M1014_d N_A_1519_125#_M1014_g N_VPWR_M1007_d VPB PHIGHVT L=0.25 W=1
+ AD=0.285 AS=0.225 PD=2.57 PS=1.45 NRD=0 NRS=0 M=1 R=4 SA=125001 SB=125000
+ A=0.25 P=2.5 MULT=1
MM1004 N_VPWR_M1004_d N_A_1519_125#_M1004_g N_A_2383_57#_M1004_s VPB PHIGHVT
+ L=0.25 W=1 AD=0.14 AS=0.285 PD=1.28 PS=2.57 NRD=0 NRS=0 M=1 R=4 SA=125000
+ SB=125001 A=0.25 P=2.5 MULT=1
MM1030 N_Q_M1030_d N_A_2383_57#_M1030_g N_VPWR_M1004_d VPB PHIGHVT L=0.25 W=1
+ AD=0.285 AS=0.14 PD=2.57 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125001 SB=125000
+ A=0.25 P=2.5 MULT=1
DX41_noxref VNB VPB NWDIODE A=26.6695 P=32.33
c_279 VPB 0 6.93588e-20 $X=0 $Y=3.085
*
.include "sky130_fd_sc_lp__dfsbp_lp.pxi.spice"
*
.ends
*
*
