# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_lp__buflp_8
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  10.56000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  1.890000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.535000 1.180000 2.255000 1.185000 ;
        RECT 0.535000 1.185000 2.565000 1.515000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  2.822400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.235000 1.765000 10.435000 1.935000 ;
        RECT 6.235000 1.935000  6.565000 2.735000 ;
        RECT 6.405000 0.595000  6.575000 0.925000 ;
        RECT 6.405000 0.925000 10.435000 1.095000 ;
        RECT 7.235000 1.935000  7.565000 2.735000 ;
        RECT 7.265000 0.595000  7.515000 0.925000 ;
        RECT 8.185000 0.595000  8.515000 0.925000 ;
        RECT 8.235000 1.935000  8.565000 2.735000 ;
        RECT 9.185000 0.595000  9.515000 0.925000 ;
        RECT 9.235000 1.935000  9.565000 2.735000 ;
        RECT 9.995000 1.095000 10.435000 1.765000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 10.560000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.500000 0.500000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.800000 0.500000 3.300000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 10.560000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 10.560000 0.085000 ;
      RECT  0.000000  3.245000 10.560000 3.415000 ;
      RECT  0.115000  0.255000  0.365000 0.840000 ;
      RECT  0.115000  0.840000  1.375000 1.010000 ;
      RECT  0.115000  1.010000  0.365000 1.095000 ;
      RECT  0.115000  1.685000  2.985000 1.855000 ;
      RECT  0.115000  1.855000  0.365000 3.075000 ;
      RECT  0.195000  1.095000  0.365000 1.685000 ;
      RECT  0.545000  0.255000  1.725000 0.425000 ;
      RECT  0.545000  0.425000  0.875000 0.670000 ;
      RECT  0.545000  2.025000  0.875000 2.905000 ;
      RECT  0.545000  2.905000  1.735000 3.075000 ;
      RECT  1.045000  0.595000  1.375000 0.840000 ;
      RECT  1.055000  1.855000  1.225000 2.735000 ;
      RECT  1.405000  2.025000  2.595000 2.195000 ;
      RECT  1.405000  2.195000  1.735000 2.905000 ;
      RECT  1.555000  0.425000  1.725000 0.775000 ;
      RECT  1.555000  0.775000  2.665000 1.010000 ;
      RECT  1.905000  0.085000  2.155000 0.605000 ;
      RECT  1.915000  2.365000  2.085000 3.245000 ;
      RECT  2.265000  2.195000  2.595000 3.075000 ;
      RECT  2.335000  0.255000  2.665000 0.775000 ;
      RECT  2.335000  1.010000  2.665000 1.015000 ;
      RECT  2.775000  2.025000  2.945000 3.245000 ;
      RECT  2.815000  1.265000  9.820000 1.595000 ;
      RECT  2.815000  1.595000  2.985000 1.685000 ;
      RECT  2.845000  0.085000  3.015000 1.095000 ;
      RECT  3.155000  1.765000  6.065000 1.935000 ;
      RECT  3.155000  1.935000  3.485000 3.075000 ;
      RECT  3.195000  0.255000  3.445000 0.925000 ;
      RECT  3.195000  0.925000  6.225000 1.095000 ;
      RECT  3.625000  0.085000  3.875000 0.755000 ;
      RECT  3.665000  2.105000  3.835000 3.245000 ;
      RECT  4.015000  1.935000  4.345000 3.075000 ;
      RECT  4.055000  0.255000  4.305000 0.925000 ;
      RECT  4.485000  0.085000  4.815000 0.755000 ;
      RECT  4.525000  2.105000  4.695000 3.245000 ;
      RECT  4.875000  1.935000  5.205000 3.075000 ;
      RECT  5.035000  0.255000  5.285000 0.925000 ;
      RECT  5.385000  2.105000  5.555000 3.245000 ;
      RECT  5.465000  0.085000  5.715000 0.755000 ;
      RECT  5.735000  1.935000  6.065000 2.905000 ;
      RECT  5.735000  2.905000  9.915000 3.075000 ;
      RECT  5.895000  0.255000  9.945000 0.425000 ;
      RECT  5.895000  0.425000  6.225000 0.925000 ;
      RECT  6.735000  2.105000  7.065000 2.905000 ;
      RECT  6.755000  0.425000  7.085000 0.755000 ;
      RECT  7.685000  0.425000  8.015000 0.755000 ;
      RECT  7.735000  2.105000  8.065000 2.905000 ;
      RECT  8.685000  0.425000  9.015000 0.755000 ;
      RECT  8.735000  2.105000  9.065000 2.905000 ;
      RECT  9.695000  0.425000  9.945000 0.755000 ;
      RECT  9.745000  2.105000  9.915000 2.905000 ;
      RECT 10.095000  2.105000 10.425000 3.245000 ;
      RECT 10.115000  0.085000 10.445000 0.755000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
  END
END sky130_fd_sc_lp__buflp_8
END LIBRARY
