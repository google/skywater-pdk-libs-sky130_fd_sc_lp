* NGSPICE file created from sky130_fd_sc_lp__o311ai_m.ext - technology: sky130A

.subckt sky130_fd_sc_lp__o311ai_m A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
M1000 VPWR B1 Y VPB phighvt w=420000u l=150000u
+  ad=3.5825e+11p pd=3.42e+06u as=2.289e+11p ps=2.77e+06u
M1001 a_220_403# A2 a_148_403# VPB phighvt w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=8.82e+10p ps=1.26e+06u
M1002 Y A3 a_220_403# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 Y C1 VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_136_82# A3 VGND VNB nshort w=420000u l=150000u
+  ad=2.352e+11p pd=2.8e+06u as=2.289e+11p ps=2.77e+06u
M1005 a_148_403# A1 VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_394_82# B1 a_136_82# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1007 Y C1 a_394_82# VNB nshort w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1008 a_136_82# A1 VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND A2 a_136_82# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

