* File: sky130_fd_sc_lp__decap_6.pxi.spice
* Created: Fri Aug 28 10:20:04 2020
* 
x_PM_SKY130_FD_SC_LP__DECAP_6%VGND N_VGND_M1001_s N_VGND_c_24_n N_VGND_c_25_n
+ N_VGND_c_26_n N_VGND_c_27_n N_VGND_c_28_n N_VGND_c_29_n N_VGND_c_30_n VGND
+ N_VGND_M1000_g N_VGND_c_31_n N_VGND_c_32_n PM_SKY130_FD_SC_LP__DECAP_6%VGND
x_PM_SKY130_FD_SC_LP__DECAP_6%VPWR N_VPWR_M1000_s N_VPWR_c_53_n N_VPWR_c_54_n
+ N_VPWR_c_50_n N_VPWR_c_51_n N_VPWR_c_57_n N_VPWR_c_58_n VPWR N_VPWR_M1001_g
+ N_VPWR_c_59_n N_VPWR_c_52_n PM_SKY130_FD_SC_LP__DECAP_6%VPWR
cc_1 VNB N_VGND_c_24_n 0.012758f $X=-0.19 $Y=-0.245 $X2=0.335 $Y2=0.085
cc_2 VNB N_VGND_c_25_n 0.0651019f $X=-0.19 $Y=-0.245 $X2=0.335 $Y2=0.38
cc_3 VNB N_VGND_c_26_n 0.00211035f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=1.77
cc_4 VNB N_VGND_c_27_n 4.97259e-19 $X=-0.19 $Y=-0.245 $X2=0.915 $Y2=1.77
cc_5 VNB N_VGND_c_28_n 0.0193278f $X=-0.19 $Y=-0.245 $X2=0.915 $Y2=1.77
cc_6 VNB N_VGND_c_29_n 0.0105251f $X=-0.19 $Y=-0.245 $X2=2.615 $Y2=0.085
cc_7 VNB N_VGND_c_30_n 0.0403852f $X=-0.19 $Y=-0.245 $X2=2.615 $Y2=0.405
cc_8 VNB N_VGND_c_31_n 0.0598957f $X=-0.19 $Y=-0.245 $X2=2.45 $Y2=0
cc_9 VNB N_VGND_c_32_n 0.170588f $X=-0.19 $Y=-0.245 $X2=2.64 $Y2=0
cc_10 VNB N_VPWR_c_50_n 0.0155672f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=1.77
cc_11 VNB N_VPWR_c_51_n 0.216628f $X=-0.19 $Y=-0.245 $X2=0.915 $Y2=1.77
cc_12 VNB N_VPWR_c_52_n 0.123877f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=0
cc_13 VPB N_VGND_c_26_n 0.0140672f $X=-0.19 $Y=1.655 $X2=0.5 $Y2=1.77
cc_14 VPB N_VGND_c_27_n 0.00874558f $X=-0.19 $Y=1.655 $X2=0.915 $Y2=1.77
cc_15 VPB N_VGND_c_28_n 0.220836f $X=-0.19 $Y=1.655 $X2=0.915 $Y2=1.77
cc_16 VPB N_VPWR_c_53_n 0.0103989f $X=-0.19 $Y=1.655 $X2=0.335 $Y2=0.085
cc_17 VPB N_VPWR_c_54_n 0.0425694f $X=-0.19 $Y=1.655 $X2=0.335 $Y2=0.38
cc_18 VPB N_VPWR_c_50_n 8.51536e-19 $X=-0.19 $Y=1.655 $X2=0.5 $Y2=1.77
cc_19 VPB N_VPWR_c_51_n 0.0211573f $X=-0.19 $Y=1.655 $X2=0.915 $Y2=1.77
cc_20 VPB N_VPWR_c_57_n 0.0125726f $X=-0.19 $Y=1.655 $X2=2.615 $Y2=1.085
cc_21 VPB N_VPWR_c_58_n 0.0654031f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_22 VPB N_VPWR_c_59_n 0.0602139f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=0
cc_23 VPB N_VPWR_c_52_n 0.0463038f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=0
cc_24 N_VGND_c_26_n N_VPWR_c_54_n 0.0205458f $X=0.5 $Y=1.77 $X2=0 $Y2=0
cc_25 N_VGND_c_28_n N_VPWR_c_54_n 0.0546006f $X=0.915 $Y=1.77 $X2=0 $Y2=0
cc_26 N_VGND_c_27_n N_VPWR_c_50_n 0.0024823f $X=0.915 $Y=1.77 $X2=0 $Y2=0
cc_27 N_VGND_c_28_n N_VPWR_c_50_n 0.0064509f $X=0.915 $Y=1.77 $X2=0 $Y2=0
cc_28 N_VGND_c_30_n N_VPWR_c_50_n 0.0214376f $X=2.615 $Y=0.405 $X2=0 $Y2=0
cc_29 N_VGND_c_25_n N_VPWR_c_51_n 0.0654854f $X=0.335 $Y=0.38 $X2=0 $Y2=0
cc_30 N_VGND_c_27_n N_VPWR_c_51_n 0.00473507f $X=0.915 $Y=1.77 $X2=0 $Y2=0
cc_31 N_VGND_c_28_n N_VPWR_c_51_n 0.127834f $X=0.915 $Y=1.77 $X2=0 $Y2=0
cc_32 N_VGND_c_30_n N_VPWR_c_51_n 0.0532165f $X=2.615 $Y=0.405 $X2=0 $Y2=0
cc_33 N_VGND_c_31_n N_VPWR_c_51_n 0.0760645f $X=2.45 $Y=0 $X2=0 $Y2=0
cc_34 N_VGND_c_32_n N_VPWR_c_51_n 0.120027f $X=2.64 $Y=0 $X2=0 $Y2=0
cc_35 N_VGND_c_28_n N_VPWR_c_58_n 0.0710714f $X=0.915 $Y=1.77 $X2=0 $Y2=0
cc_36 N_VGND_c_28_n N_VPWR_c_59_n 0.0764547f $X=0.915 $Y=1.77 $X2=0 $Y2=0
cc_37 N_VGND_c_28_n N_VPWR_c_52_n 0.120644f $X=0.915 $Y=1.77 $X2=0 $Y2=0
