* NGSPICE file created from sky130_fd_sc_lp__dfstp_4.ext - technology: sky130A

.subckt sky130_fd_sc_lp__dfstp_4 CLK D SET_B VGND VNB VPB VPWR Q
M1000 a_690_463# a_30_99# a_562_119# VPB phighvt w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=1.176e+11p ps=1.4e+06u
M1001 a_230_465# a_30_99# VGND VNB nshort w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=1.8475e+12p ps=1.655e+07u
M1002 a_562_119# a_30_99# a_476_119# VNB nshort w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=1.176e+11p ps=1.4e+06u
M1003 VPWR SET_B a_690_93# VPB phighvt w=420000u l=150000u
+  ad=2.05945e+12p pd=1.957e+07u as=1.176e+11p ps=1.4e+06u
M1004 Q a_1989_49# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=7.056e+11p pd=6.16e+06u as=0p ps=0u
M1005 VPWR CLK a_30_99# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.824e+11p ps=1.85e+06u
M1006 VPWR a_690_93# a_690_463# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_914_47# a_562_119# a_690_93# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=1.113e+11p ps=1.37e+06u
M1008 a_1428_91# a_1398_65# a_1356_91# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=8.82e+10p ps=1.26e+06u
M1009 VGND SET_B a_914_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND a_1989_49# Q VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=4.704e+11p ps=4.48e+06u
M1011 VPWR a_1247_47# a_1989_49# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=3.339e+11p ps=3.05e+06u
M1012 VGND a_1247_47# a_1989_49# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=2.226e+11p ps=2.21e+06u
M1013 VGND CLK a_30_99# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1014 VPWR a_1398_65# a_1201_407# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=2.226e+11p ps=2.74e+06u
M1015 a_1175_47# a_562_119# VGND VNB nshort w=640000u l=150000u
+  ad=1.344e+11p pd=1.7e+06u as=0p ps=0u
M1016 a_690_93# a_562_119# VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VPWR a_1989_49# Q VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_1247_47# a_230_465# a_1175_47# VNB nshort w=640000u l=150000u
+  ad=2.242e+11p pd=2.07e+06u as=0p ps=0u
M1019 a_562_119# a_230_465# a_476_119# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.176e+11p ps=1.4e+06u
M1020 a_1094_379# a_562_119# VPWR VPB phighvt w=840000u l=150000u
+  ad=5.825e+11p pd=5.07e+06u as=0p ps=0u
M1021 a_1356_91# a_30_99# a_1247_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VPWR a_1989_49# Q VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 Q a_1989_49# VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_1398_65# a_1247_47# VPWR VPB phighvt w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1025 a_230_465# a_30_99# VPWR VPB phighvt w=640000u l=150000u
+  ad=1.696e+11p pd=1.81e+06u as=0p ps=0u
M1026 a_1094_379# a_30_99# a_1247_47# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=3.801e+11p ps=3.8e+06u
M1027 a_648_119# a_230_465# a_562_119# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1028 a_1398_65# a_1247_47# VGND VNB nshort w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1029 VGND a_1989_49# Q VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 Q a_1989_49# VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_476_119# D VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 a_1247_47# SET_B VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 Q a_1989_49# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1034 VGND SET_B a_1428_91# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1035 VGND a_690_93# a_648_119# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1036 a_1247_47# a_230_465# a_1201_407# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1037 a_476_119# D VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

