* File: sky130_fd_sc_lp__nand2b_m.pex.spice
* Created: Fri Aug 28 10:48:39 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__NAND2B_M%A_N 3 6 9 11 12 13 14 15 16 23
r38 23 25 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=0.682 $Y=1.205
+ $X2=0.682 $Y2=1.04
r39 23 24 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.705
+ $Y=1.205 $X2=0.705 $Y2=1.205
r40 15 16 22.1818 $w=1.83e-07 $l=3.7e-07 $layer=LI1_cond $X=0.712 $Y=1.665
+ $X2=0.712 $Y2=2.035
r41 14 15 22.1818 $w=1.83e-07 $l=3.7e-07 $layer=LI1_cond $X=0.712 $Y=1.295
+ $X2=0.712 $Y2=1.665
r42 14 24 5.39558 $w=1.83e-07 $l=9e-08 $layer=LI1_cond $X=0.712 $Y=1.295
+ $X2=0.712 $Y2=1.205
r43 13 24 16.7862 $w=1.83e-07 $l=2.8e-07 $layer=LI1_cond $X=0.712 $Y=0.925
+ $X2=0.712 $Y2=1.205
r44 12 13 22.1818 $w=1.83e-07 $l=3.7e-07 $layer=LI1_cond $X=0.712 $Y=0.555
+ $X2=0.712 $Y2=0.925
r45 9 11 594.809 $w=1.5e-07 $l=1.16e-06 $layer=POLY_cond $X=0.795 $Y=2.87
+ $X2=0.795 $Y2=1.71
r46 6 11 48.4185 $w=3.75e-07 $l=1.87e-07 $layer=POLY_cond $X=0.682 $Y=1.523
+ $X2=0.682 $Y2=1.71
r47 5 23 3.26277 $w=3.75e-07 $l=2.2e-08 $layer=POLY_cond $X=0.682 $Y=1.227
+ $X2=0.682 $Y2=1.205
r48 5 6 43.8991 $w=3.75e-07 $l=2.96e-07 $layer=POLY_cond $X=0.682 $Y=1.227
+ $X2=0.682 $Y2=1.523
r49 3 25 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=0.57 $Y=0.48 $X2=0.57
+ $Y2=1.04
.ends

.subckt PM_SKY130_FD_SC_LP__NAND2B_M%B 3 7 9 10 11 12 13 17
c46 3 0 2.89892e-19 $X=1.225 $Y=2.87
r47 12 13 19.8327 $w=2.13e-07 $l=3.7e-07 $layer=LI1_cond $X=1.222 $Y=0.925
+ $X2=1.222 $Y2=1.295
r48 12 17 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.245
+ $Y=0.965 $X2=1.245 $Y2=0.965
r49 10 17 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.245 $Y=1.305
+ $X2=1.245 $Y2=0.965
r50 10 11 38.6168 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.245 $Y=1.305
+ $X2=1.245 $Y2=1.47
r51 9 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.245 $Y=0.8
+ $X2=1.245 $Y2=0.965
r52 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.335 $Y=0.48
+ $X2=1.335 $Y2=0.8
r53 3 11 717.872 $w=1.5e-07 $l=1.4e-06 $layer=POLY_cond $X=1.225 $Y=2.87
+ $X2=1.225 $Y2=1.47
.ends

.subckt PM_SKY130_FD_SC_LP__NAND2B_M%A_46_54# 1 2 9 13 17 18 19 20 21 24 28 30
+ 31 32 36 37 42
c68 30 0 1.72444e-19 $X=0.985 $Y=2.385
r69 42 44 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.07 $Y=2.215
+ $X2=1.07 $Y2=2.385
r70 36 37 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.705
+ $Y=1.875 $X2=1.705 $Y2=1.875
r71 34 36 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=1.705 $Y=2.13
+ $X2=1.705 $Y2=1.875
r72 33 42 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.155 $Y=2.215
+ $X2=1.07 $Y2=2.215
r73 32 34 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.54 $Y=2.215
+ $X2=1.705 $Y2=2.13
r74 32 33 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=1.54 $Y=2.215
+ $X2=1.155 $Y2=2.215
r75 30 44 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.985 $Y=2.385
+ $X2=1.07 $Y2=2.385
r76 30 31 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=0.985 $Y=2.385
+ $X2=0.685 $Y2=2.385
r77 26 31 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=0.58 $Y=2.385
+ $X2=0.685 $Y2=2.385
r78 26 39 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=0.58 $Y=2.385
+ $X2=0.345 $Y2=2.385
r79 26 28 17.6926 $w=2.08e-07 $l=3.35e-07 $layer=LI1_cond $X=0.58 $Y=2.47
+ $X2=0.58 $Y2=2.805
r80 22 39 0.0262452 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=0.345 $Y=2.3
+ $X2=0.345 $Y2=2.385
r81 22 24 102.445 $w=1.88e-07 $l=1.755e-06 $layer=LI1_cond $X=0.345 $Y=2.3
+ $X2=0.345 $Y2=0.545
r82 20 21 58.3064 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=1.71 $Y=0.8 $X2=1.71
+ $Y2=0.95
r83 18 37 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.705 $Y=2.215
+ $X2=1.705 $Y2=1.875
r84 18 19 40.8701 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.705 $Y=2.215
+ $X2=1.705 $Y2=2.38
r85 17 37 38.6168 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.705 $Y=1.71
+ $X2=1.705 $Y2=1.875
r86 17 21 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=1.725 $Y=1.71
+ $X2=1.725 $Y2=0.95
r87 13 20 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.695 $Y=0.48
+ $X2=1.695 $Y2=0.8
r88 9 19 251.255 $w=1.5e-07 $l=4.9e-07 $layer=POLY_cond $X=1.655 $Y=2.87
+ $X2=1.655 $Y2=2.38
r89 2 28 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.455
+ $Y=2.66 $X2=0.58 $Y2=2.805
r90 1 24 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=0.23
+ $Y=0.27 $X2=0.355 $Y2=0.545
.ends

.subckt PM_SKY130_FD_SC_LP__NAND2B_M%VPWR 1 2 9 13 16 17 19 20 21 31 32
r34 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r35 29 32 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r36 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r37 24 25 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r38 21 29 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r39 21 25 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r40 19 28 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=1.705 $Y=3.33
+ $X2=1.68 $Y2=3.33
r41 19 20 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.705 $Y=3.33
+ $X2=1.87 $Y2=3.33
r42 18 31 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=2.035 $Y=3.33
+ $X2=2.16 $Y2=3.33
r43 18 20 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.035 $Y=3.33
+ $X2=1.87 $Y2=3.33
r44 16 24 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=0.905 $Y=3.33
+ $X2=0.72 $Y2=3.33
r45 16 17 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=0.905 $Y=3.33
+ $X2=1.01 $Y2=3.33
r46 15 28 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=1.115 $Y=3.33
+ $X2=1.68 $Y2=3.33
r47 15 17 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.115 $Y=3.33
+ $X2=1.01 $Y2=3.33
r48 11 20 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.87 $Y=3.245
+ $X2=1.87 $Y2=3.33
r49 11 13 10.826 $w=3.28e-07 $l=3.1e-07 $layer=LI1_cond $X=1.87 $Y=3.245
+ $X2=1.87 $Y2=2.935
r50 7 17 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=1.01 $Y=3.245
+ $X2=1.01 $Y2=3.33
r51 7 9 16.3723 $w=2.08e-07 $l=3.1e-07 $layer=LI1_cond $X=1.01 $Y=3.245 $X2=1.01
+ $Y2=2.935
r52 2 13 600 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=1 $X=1.73
+ $Y=2.66 $X2=1.87 $Y2=2.935
r53 1 9 600 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=1 $X=0.87
+ $Y=2.66 $X2=1.01 $Y2=2.935
.ends

.subckt PM_SKY130_FD_SC_LP__NAND2B_M%Y 1 2 9 11 12 13 14 15 16 17 27 28 39
c38 9 0 2.86763e-19 $X=1.44 $Y=2.805
r39 28 39 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=2.16 $Y=2.48
+ $X2=2.16 $Y2=2.405
r40 17 28 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.16 $Y=2.565
+ $X2=2.16 $Y2=2.48
r41 17 39 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=2.16 $Y=2.4 $X2=2.16
+ $Y2=2.405
r42 16 17 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=2.16 $Y=2.035
+ $X2=2.16 $Y2=2.4
r43 15 16 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=2.16 $Y=1.665
+ $X2=2.16 $Y2=2.035
r44 14 15 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=2.16 $Y=1.295
+ $X2=2.16 $Y2=1.665
r45 13 14 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=2.16 $Y=0.925
+ $X2=2.16 $Y2=1.295
r46 13 27 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=2.16 $Y=0.925
+ $X2=2.16 $Y2=0.65
r47 12 27 3.82155 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=2.16 $Y=0.545
+ $X2=2.16 $Y2=0.65
r48 12 42 7.29301 $w=3.78e-07 $l=1.65e-07 $layer=LI1_cond $X=2.075 $Y=0.545
+ $X2=1.91 $Y2=0.545
r49 11 17 33.9357 $w=1.78e-07 $l=5.5e-07 $layer=LI1_cond $X=1.525 $Y=2.565
+ $X2=2.075 $Y2=2.565
r50 7 11 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=1.43 $Y=2.65
+ $X2=1.525 $Y2=2.565
r51 7 9 9.04785 $w=1.88e-07 $l=1.55e-07 $layer=LI1_cond $X=1.43 $Y=2.65 $X2=1.43
+ $Y2=2.805
r52 2 9 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.3
+ $Y=2.66 $X2=1.44 $Y2=2.805
r53 1 42 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=1.77
+ $Y=0.27 $X2=1.91 $Y2=0.545
.ends

.subckt PM_SKY130_FD_SC_LP__NAND2B_M%VGND 1 6 9 10 11 21 22
r27 21 22 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r28 18 21 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r29 14 15 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r30 11 22 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r31 11 15 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r32 11 18 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r33 9 14 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.985 $Y=0 $X2=0.72
+ $Y2=0
r34 9 10 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=0.985 $Y=0 $X2=1.09
+ $Y2=0
r35 8 18 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=1.195 $Y=0 $X2=1.2
+ $Y2=0
r36 8 10 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.195 $Y=0 $X2=1.09
+ $Y2=0
r37 4 10 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=1.09 $Y=0.085
+ $X2=1.09 $Y2=0
r38 4 6 17.4286 $w=2.08e-07 $l=3.3e-07 $layer=LI1_cond $X=1.09 $Y=0.085 $X2=1.09
+ $Y2=0.415
r39 1 6 182 $w=1.7e-07 $l=5.12396e-07 $layer=licon1_NDIFF $count=1 $X=0.645
+ $Y=0.27 $X2=1.09 $Y2=0.415
.ends

