* NGSPICE file created from sky130_fd_sc_lp__a21oi_1.ext - technology: sky130A

.subckt sky130_fd_sc_lp__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
M1000 Y A1 a_110_69# VNB nshort w=840000u l=150000u
+  ad=3.276e+11p pd=2.46e+06u as=2.016e+11p ps=2.16e+06u
M1001 Y B1 a_27_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=3.339e+11p pd=3.05e+06u as=6.867e+11p ps=6.13e+06u
M1002 a_110_69# A2 VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=4.662e+11p ps=4.47e+06u
M1003 VGND B1 Y VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_27_367# A1 VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=4.41e+11p ps=3.22e+06u
M1005 VPWR A2 a_27_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

