* File: sky130_fd_sc_lp__o221ai_m.pex.spice
* Created: Wed Sep  2 10:19:33 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O221AI_M%C1 5 7 9 12 14 17 19
c44 12 0 1.05734e-19 $X=0.665 $Y=0.84
r45 17 20 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.67 $Y=2.035
+ $X2=0.67 $Y2=2.2
r46 17 19 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.67 $Y=2.035
+ $X2=0.67 $Y2=1.87
r47 14 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.67
+ $Y=2.035 $X2=0.67 $Y2=2.035
r48 10 12 43.5851 $w=1.5e-07 $l=8.5e-08 $layer=POLY_cond $X=0.58 $Y=0.84
+ $X2=0.665 $Y2=0.84
r49 7 12 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.665 $Y=0.765
+ $X2=0.665 $Y2=0.84
r50 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.665 $Y=0.765
+ $X2=0.665 $Y2=0.445
r51 5 20 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=0.6 $Y=2.61 $X2=0.6
+ $Y2=2.2
r52 1 10 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.58 $Y=0.915
+ $X2=0.58 $Y2=0.84
r53 1 19 489.691 $w=1.5e-07 $l=9.55e-07 $layer=POLY_cond $X=0.58 $Y=0.915
+ $X2=0.58 $Y2=1.87
.ends

.subckt PM_SKY130_FD_SC_LP__O221AI_M%B1 3 7 9 12
c47 12 0 1.22854e-19 $X=1.06 $Y=1.32
r48 12 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.06 $Y=1.32
+ $X2=1.06 $Y2=1.485
r49 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.06 $Y=1.32
+ $X2=1.06 $Y2=1.155
r50 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.06
+ $Y=1.32 $X2=1.06 $Y2=1.32
r51 9 13 7.9627 $w=1.93e-07 $l=1.4e-07 $layer=LI1_cond $X=1.2 $Y=1.307 $X2=1.06
+ $Y2=1.307
r52 7 15 576.862 $w=1.5e-07 $l=1.125e-06 $layer=POLY_cond $X=1.15 $Y=2.61
+ $X2=1.15 $Y2=1.485
r53 3 14 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=1.095 $Y=0.445
+ $X2=1.095 $Y2=1.155
.ends

.subckt PM_SKY130_FD_SC_LP__O221AI_M%A2 3 6 7 9 12 13 16 19
r45 19 20 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.63
+ $Y=1.08 $X2=1.63 $Y2=1.08
r46 16 20 1.17263 $w=5.08e-07 $l=5e-08 $layer=LI1_cond $X=1.68 $Y=1.25 $X2=1.63
+ $Y2=1.25
r47 12 19 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.63 $Y=1.42
+ $X2=1.63 $Y2=1.08
r48 12 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.63 $Y=1.42
+ $X2=1.63 $Y2=1.585
r49 11 19 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.63 $Y=0.915
+ $X2=1.63 $Y2=1.08
r50 7 9 106.04 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=2.13 $Y=2.195 $X2=2.13
+ $Y2=2.525
r51 6 7 101.866 $w=1.94e-07 $l=5.45206e-07 $layer=POLY_cond $X=1.72 $Y=1.88
+ $X2=2.13 $Y2=2.195
r52 6 13 151.266 $w=1.5e-07 $l=2.95e-07 $layer=POLY_cond $X=1.72 $Y=1.88
+ $X2=1.72 $Y2=1.585
r53 3 11 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=1.54 $Y=0.445 $X2=1.54
+ $Y2=0.915
.ends

.subckt PM_SKY130_FD_SC_LP__O221AI_M%A1 3 7 9 10 14
r34 14 16 28.2737 $w=3.58e-07 $l=2.1e-07 $layer=POLY_cond $X=2.49 $Y=1.812
+ $X2=2.7 $Y2=1.812
r35 9 10 23.5393 $w=2.33e-07 $l=4.8e-07 $layer=LI1_cond $X=2.64 $Y=2.002
+ $X2=3.12 $Y2=2.002
r36 9 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.7 $Y=1.97
+ $X2=2.7 $Y2=1.97
r37 5 14 23.1716 $w=1.5e-07 $l=3.23e-07 $layer=POLY_cond $X=2.49 $Y=2.135
+ $X2=2.49 $Y2=1.812
r38 5 7 199.979 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=2.49 $Y=2.135 $X2=2.49
+ $Y2=2.525
r39 1 14 51.162 $w=3.58e-07 $l=5.16488e-07 $layer=POLY_cond $X=2.11 $Y=1.49
+ $X2=2.49 $Y2=1.812
r40 1 3 535.84 $w=1.5e-07 $l=1.045e-06 $layer=POLY_cond $X=2.11 $Y=1.49 $X2=2.11
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__O221AI_M%B2 3 5 6 9 10 11 13 15 16 18 21
c55 15 0 9.3038e-20 $X=2.685 $Y=0.765
r56 21 22 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.74
+ $Y=0.93 $X2=2.74 $Y2=0.93
r57 18 22 0.164635 $w=3.48e-07 $l=5e-09 $layer=LI1_cond $X=2.73 $Y=0.925
+ $X2=2.73 $Y2=0.93
r58 17 21 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=2.74 $Y=1.285
+ $X2=2.74 $Y2=0.93
r59 16 21 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=2.74 $Y=0.915
+ $X2=2.74 $Y2=0.93
r60 15 16 43.5886 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=2.685 $Y=0.765
+ $X2=2.685 $Y2=0.915
r61 12 13 840.936 $w=1.5e-07 $l=1.64e-06 $layer=POLY_cond $X=3.18 $Y=1.435
+ $X2=3.18 $Y2=3.075
r62 11 17 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=2.905 $Y=1.36
+ $X2=2.74 $Y2=1.285
r63 10 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.105 $Y=1.36
+ $X2=3.18 $Y2=1.435
r64 10 11 102.553 $w=1.5e-07 $l=2e-07 $layer=POLY_cond $X=3.105 $Y=1.36
+ $X2=2.905 $Y2=1.36
r65 9 15 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.54 $Y=0.445
+ $X2=2.54 $Y2=0.765
r66 5 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.105 $Y=3.15
+ $X2=3.18 $Y2=3.075
r67 5 6 779.404 $w=1.5e-07 $l=1.52e-06 $layer=POLY_cond $X=3.105 $Y=3.15
+ $X2=1.585 $Y2=3.15
r68 1 6 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.51 $Y=3.075
+ $X2=1.585 $Y2=3.15
r69 1 3 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.51 $Y=3.075
+ $X2=1.51 $Y2=2.61
.ends

.subckt PM_SKY130_FD_SC_LP__O221AI_M%Y 1 2 3 10 12 17 18 19 20 21 22 23 53
r48 23 45 7.9123 $w=3.33e-07 $l=2.3e-07 $layer=LI1_cond $X=0.322 $Y=2.775
+ $X2=0.322 $Y2=2.545
r49 22 33 3.67481 $w=2.52e-07 $l=1.19143e-07 $layer=LI1_cond $X=0.322 $Y=2.385
+ $X2=0.24 $Y2=2.3
r50 22 42 3.67481 $w=2.52e-07 $l=8.5e-08 $layer=LI1_cond $X=0.322 $Y=2.385
+ $X2=0.322 $Y2=2.47
r51 22 45 2.23608 $w=3.33e-07 $l=6.5e-08 $layer=LI1_cond $X=0.322 $Y=2.48
+ $X2=0.322 $Y2=2.545
r52 22 42 0.344013 $w=3.33e-07 $l=1e-08 $layer=LI1_cond $X=0.322 $Y=2.48
+ $X2=0.322 $Y2=2.47
r53 21 33 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.24 $Y=2.035
+ $X2=0.24 $Y2=2.3
r54 20 21 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.24 $Y=1.665
+ $X2=0.24 $Y2=2.035
r55 19 20 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.24 $Y=1.295
+ $X2=0.24 $Y2=1.665
r56 18 19 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.24 $Y=0.925
+ $X2=0.24 $Y2=1.295
r57 18 32 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=0.24 $Y=0.925
+ $X2=0.24 $Y2=0.675
r58 17 53 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=0.24 $Y=0.51
+ $X2=0.45 $Y2=0.51
r59 17 32 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.24 $Y=0.51
+ $X2=0.24 $Y2=0.675
r60 12 15 4.22511 $w=2.08e-07 $l=8e-08 $layer=LI1_cond $X=1.82 $Y=2.385 $X2=1.82
+ $Y2=2.465
r61 11 22 2.79892 $w=1.7e-07 $l=1.68e-07 $layer=LI1_cond $X=0.49 $Y=2.385
+ $X2=0.322 $Y2=2.385
r62 10 12 1.9771 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.715 $Y=2.385
+ $X2=1.82 $Y2=2.385
r63 10 11 79.9198 $w=1.68e-07 $l=1.225e-06 $layer=LI1_cond $X=1.715 $Y=2.385
+ $X2=0.49 $Y2=2.385
r64 3 15 600 $w=1.7e-07 $l=2.65518e-07 $layer=licon1_PDIFF $count=1 $X=1.585
+ $Y=2.4 $X2=1.82 $Y2=2.465
r65 2 45 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.26
+ $Y=2.4 $X2=0.385 $Y2=2.545
r66 1 53 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=0.325
+ $Y=0.235 $X2=0.45 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_LP__O221AI_M%VPWR 1 2 11 15 17 19 29 30 33 36
r36 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r37 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r38 30 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.64 $Y2=3.33
r39 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r40 27 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.87 $Y=3.33
+ $X2=2.705 $Y2=3.33
r41 27 29 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=2.87 $Y=3.33
+ $X2=3.12 $Y2=3.33
r42 26 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r43 25 26 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r44 23 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r45 22 25 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=3.33 $X2=2.16
+ $Y2=3.33
r46 22 23 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r47 20 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.04 $Y=3.33
+ $X2=0.875 $Y2=3.33
r48 20 22 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=1.04 $Y=3.33 $X2=1.2
+ $Y2=3.33
r49 19 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.54 $Y=3.33
+ $X2=2.705 $Y2=3.33
r50 19 25 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=2.54 $Y=3.33
+ $X2=2.16 $Y2=3.33
r51 17 26 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r52 17 23 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r53 13 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.705 $Y=3.245
+ $X2=2.705 $Y2=3.33
r54 13 15 22.8742 $w=3.28e-07 $l=6.55e-07 $layer=LI1_cond $X=2.705 $Y=3.245
+ $X2=2.705 $Y2=2.59
r55 9 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.875 $Y=3.245
+ $X2=0.875 $Y2=3.33
r56 9 11 17.8105 $w=3.28e-07 $l=5.1e-07 $layer=LI1_cond $X=0.875 $Y=3.245
+ $X2=0.875 $Y2=2.735
r57 2 15 600 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=1 $X=2.565
+ $Y=2.315 $X2=2.705 $Y2=2.59
r58 1 11 600 $w=1.7e-07 $l=4.2335e-07 $layer=licon1_PDIFF $count=1 $X=0.675
+ $Y=2.4 $X2=0.875 $Y2=2.735
.ends

.subckt PM_SKY130_FD_SC_LP__O221AI_M%A_148_47# 1 2 8 9 10 11 13 15 17 19 24 29
+ 33
c85 19 0 9.3038e-20 $X=3.085 $Y=0.495
c86 9 0 1.05734e-19 $X=1.015 $Y=1.67
r87 33 35 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=2.06 $Y=1.62 $X2=2.06
+ $Y2=1.77
r88 29 31 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=1.1 $Y=1.67 $X2=1.1
+ $Y2=1.77
r89 23 24 57.0856 $w=1.68e-07 $l=8.75e-07 $layer=LI1_cond $X=3.17 $Y=0.66
+ $X2=3.17 $Y2=1.535
r90 19 23 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.085 $Y=0.495
+ $X2=3.17 $Y2=0.66
r91 19 21 11.5244 $w=3.28e-07 $l=3.3e-07 $layer=LI1_cond $X=3.085 $Y=0.495
+ $X2=2.755 $Y2=0.495
r92 18 33 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.145 $Y=1.62
+ $X2=2.06 $Y2=1.62
r93 17 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.085 $Y=1.62
+ $X2=3.17 $Y2=1.535
r94 17 18 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=3.085 $Y=1.62
+ $X2=2.145 $Y2=1.62
r95 16 31 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.185 $Y=1.77
+ $X2=1.1 $Y2=1.77
r96 15 35 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.975 $Y=1.77
+ $X2=2.06 $Y2=1.77
r97 15 16 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=1.975 $Y=1.77
+ $X2=1.185 $Y2=1.77
r98 11 25 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=0.88 $Y=0.945
+ $X2=0.63 $Y2=0.945
r99 11 13 18.4848 $w=2.08e-07 $l=3.5e-07 $layer=LI1_cond $X=0.88 $Y=0.86
+ $X2=0.88 $Y2=0.51
r100 9 29 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.015 $Y=1.67
+ $X2=1.1 $Y2=1.67
r101 9 10 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=1.015 $Y=1.67
+ $X2=0.715 $Y2=1.67
r102 8 10 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.63 $Y=1.585
+ $X2=0.715 $Y2=1.67
r103 7 25 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.63 $Y=1.03
+ $X2=0.63 $Y2=0.945
r104 7 8 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=0.63 $Y=1.03
+ $X2=0.63 $Y2=1.585
r105 2 21 182 $w=1.7e-07 $l=3.2249e-07 $layer=licon1_NDIFF $count=1 $X=2.615
+ $Y=0.235 $X2=2.755 $Y2=0.495
r106 1 13 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=0.74
+ $Y=0.235 $X2=0.88 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_LP__O221AI_M%A_234_47# 1 2 9 11 12 15
c23 12 0 1.22854e-19 $X=1.43 $Y=0.73
r24 13 15 7.68295 $w=2.23e-07 $l=1.5e-07 $layer=LI1_cond $X=2.317 $Y=0.645
+ $X2=2.317 $Y2=0.495
r25 11 13 11.9044 $w=1.15e-07 $l=1.4854e-07 $layer=LI1_cond $X=2.205 $Y=0.73
+ $X2=2.317 $Y2=0.645
r26 11 12 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=2.205 $Y=0.73
+ $X2=1.43 $Y2=0.73
r27 7 12 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=1.325 $Y=0.645
+ $X2=1.43 $Y2=0.73
r28 7 9 7.12987 $w=2.08e-07 $l=1.35e-07 $layer=LI1_cond $X=1.325 $Y=0.645
+ $X2=1.325 $Y2=0.51
r29 2 15 182 $w=1.7e-07 $l=3.2249e-07 $layer=licon1_NDIFF $count=1 $X=2.185
+ $Y=0.235 $X2=2.325 $Y2=0.495
r30 1 9 182 $w=1.7e-07 $l=3.43875e-07 $layer=licon1_NDIFF $count=1 $X=1.17
+ $Y=0.235 $X2=1.325 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_LP__O221AI_M%VGND 1 6 8 10 20 21 24
r44 20 21 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r45 18 21 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r46 17 20 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r47 17 18 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r48 15 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.94 $Y=0 $X2=1.775
+ $Y2=0
r49 15 17 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=1.94 $Y=0 $X2=2.16
+ $Y2=0
r50 12 13 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r51 10 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.61 $Y=0 $X2=1.775
+ $Y2=0
r52 10 12 89.3797 $w=1.68e-07 $l=1.37e-06 $layer=LI1_cond $X=1.61 $Y=0 $X2=0.24
+ $Y2=0
r53 8 18 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r54 8 13 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.68 $Y=0 $X2=0.24
+ $Y2=0
r55 8 24 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r56 4 24 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.775 $Y=0.085
+ $X2=1.775 $Y2=0
r57 4 6 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=1.775 $Y=0.085
+ $X2=1.775 $Y2=0.36
r58 1 6 182 $w=1.7e-07 $l=2.13542e-07 $layer=licon1_NDIFF $count=1 $X=1.615
+ $Y=0.235 $X2=1.775 $Y2=0.36
.ends

