* File: sky130_fd_sc_lp__a21bo_1.spice
* Created: Wed Sep  2 09:18:41 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__a21bo_1.pex.spice"
.subckt sky130_fd_sc_lp__a21bo_1  VNB VPB B1_N A1 A2 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* A2	A2
* A1	A1
* B1_N	B1_N
* VPB	VPB
* VNB	VNB
MM1005 N_VGND_M1005_d N_A_80_43#_M1005_g N_X_M1005_s VNB NSHORT L=0.15 W=0.84
+ AD=0.279933 AS=0.2226 PD=1.97333 PS=2.21 NRD=17.136 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1002 N_A_237_367#_M1002_d N_B1_N_M1002_g N_VGND_M1005_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1197 AS=0.139967 PD=1.41 PS=0.986667 NRD=0 NRS=79.5 M=1 R=2.8
+ SA=75000.8 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1007 N_A_80_43#_M1007_d N_A_237_367#_M1007_g N_VGND_M1007_s VNB NSHORT L=0.15
+ W=0.84 AD=0.189 AS=0.2226 PD=1.29 PS=2.21 NRD=12.852 NRS=0 M=1 R=5.6
+ SA=75000.2 SB=75001.1 A=0.126 P=1.98 MULT=1
MM1003 A_556_47# N_A1_M1003_g N_A_80_43#_M1007_d VNB NSHORT L=0.15 W=0.84
+ AD=0.0882 AS=0.189 PD=1.05 PS=1.29 NRD=7.14 NRS=11.424 M=1 R=5.6 SA=75000.8
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1008 N_VGND_M1008_d N_A2_M1008_g A_556_47# VNB NSHORT L=0.15 W=0.84 AD=0.2226
+ AS=0.0882 PD=2.21 PS=1.05 NRD=0 NRS=7.14 M=1 R=5.6 SA=75001.1 SB=75000.2
+ A=0.126 P=1.98 MULT=1
MM1009 N_VPWR_M1009_d N_A_80_43#_M1009_g N_X_M1009_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.285075 AS=0.3339 PD=2.4525 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75000.4 A=0.189 P=2.82 MULT=1
MM1006 N_A_237_367#_M1006_d N_B1_N_M1006_g N_VPWR_M1009_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1113 AS=0.095025 PD=1.37 PS=0.8175 NRD=0 NRS=80.3169 M=1 R=2.8
+ SA=75000.7 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1001 N_A_436_367#_M1001_d N_A_237_367#_M1001_g N_A_80_43#_M1001_s VPB PHIGHVT
+ L=0.15 W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.2 SB=75001.1 A=0.189 P=2.82 MULT=1
MM1004 N_VPWR_M1004_d N_A1_M1004_g N_A_436_367#_M1001_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.2394 AS=0.1764 PD=1.64 PS=1.54 NRD=7.8012 NRS=0 M=1 R=8.4
+ SA=75000.6 SB=75000.7 A=0.189 P=2.82 MULT=1
MM1000 N_A_436_367#_M1000_d N_A2_M1000_g N_VPWR_M1004_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.2394 PD=3.05 PS=1.64 NRD=0 NRS=7.8012 M=1 R=8.4
+ SA=75001.1 SB=75000.2 A=0.189 P=2.82 MULT=1
DX10_noxref VNB VPB NWDIODE A=7.8703 P=12.17
c_38 VNB 0 1.80672e-19 $X=0 $Y=0
*
.include "sky130_fd_sc_lp__a21bo_1.pxi.spice"
*
.ends
*
*
