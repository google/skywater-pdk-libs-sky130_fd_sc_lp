* File: sky130_fd_sc_lp__o32a_lp.pxi.spice
* Created: Wed Sep  2 10:26:19 2020
* 
x_PM_SKY130_FD_SC_LP__O32A_LP%B1 N_B1_c_78_n N_B1_c_83_n N_B1_M1005_g
+ N_B1_c_79_n N_B1_M1000_g N_B1_c_80_n N_B1_c_81_n B1 B1
+ PM_SKY130_FD_SC_LP__O32A_LP%B1
x_PM_SKY130_FD_SC_LP__O32A_LP%B2 N_B2_c_114_n N_B2_M1007_g N_B2_M1009_g
+ N_B2_c_115_n B2 B2 B2 B2 N_B2_c_112_n N_B2_c_113_n
+ PM_SKY130_FD_SC_LP__O32A_LP%B2
x_PM_SKY130_FD_SC_LP__O32A_LP%A3 N_A3_M1010_g N_A3_M1004_g N_A3_c_162_n
+ N_A3_c_163_n A3 N_A3_c_160_n N_A3_c_161_n PM_SKY130_FD_SC_LP__O32A_LP%A3
x_PM_SKY130_FD_SC_LP__O32A_LP%A2 N_A2_M1001_g N_A2_c_210_n N_A2_M1012_g
+ N_A2_c_211_n A2 N_A2_c_208_n N_A2_c_209_n PM_SKY130_FD_SC_LP__O32A_LP%A2
x_PM_SKY130_FD_SC_LP__O32A_LP%A1 N_A1_M1003_g N_A1_c_260_n N_A1_M1002_g
+ N_A1_c_255_n N_A1_c_256_n N_A1_c_261_n A1 N_A1_c_257_n N_A1_c_258_n
+ N_A1_c_259_n PM_SKY130_FD_SC_LP__O32A_LP%A1
x_PM_SKY130_FD_SC_LP__O32A_LP%A_134_101# N_A_134_101#_M1000_d
+ N_A_134_101#_M1007_d N_A_134_101#_c_303_n N_A_134_101#_M1008_g
+ N_A_134_101#_M1006_g N_A_134_101#_M1011_g N_A_134_101#_c_304_n
+ N_A_134_101#_c_305_n N_A_134_101#_c_306_n N_A_134_101#_c_307_n
+ N_A_134_101#_c_308_n N_A_134_101#_c_327_n N_A_134_101#_c_314_n
+ N_A_134_101#_c_315_n N_A_134_101#_c_309_n N_A_134_101#_c_310_n
+ N_A_134_101#_c_316_n N_A_134_101#_c_311_n
+ PM_SKY130_FD_SC_LP__O32A_LP%A_134_101#
x_PM_SKY130_FD_SC_LP__O32A_LP%VPWR N_VPWR_M1005_s N_VPWR_M1002_d N_VPWR_c_400_n
+ N_VPWR_c_401_n N_VPWR_c_402_n N_VPWR_c_403_n N_VPWR_c_404_n VPWR
+ N_VPWR_c_405_n N_VPWR_c_399_n PM_SKY130_FD_SC_LP__O32A_LP%VPWR
x_PM_SKY130_FD_SC_LP__O32A_LP%X N_X_M1011_d N_X_M1006_d N_X_c_447_n X X X
+ N_X_c_448_n X PM_SKY130_FD_SC_LP__O32A_LP%X
x_PM_SKY130_FD_SC_LP__O32A_LP%A_31_101# N_A_31_101#_M1000_s N_A_31_101#_M1009_d
+ N_A_31_101#_M1001_d N_A_31_101#_c_470_n N_A_31_101#_c_471_n
+ N_A_31_101#_c_472_n N_A_31_101#_c_479_n N_A_31_101#_c_485_n
+ N_A_31_101#_c_482_n N_A_31_101#_c_473_n PM_SKY130_FD_SC_LP__O32A_LP%A_31_101#
x_PM_SKY130_FD_SC_LP__O32A_LP%VGND N_VGND_M1010_d N_VGND_M1003_d N_VGND_c_512_n
+ N_VGND_c_513_n N_VGND_c_514_n VGND N_VGND_c_515_n N_VGND_c_516_n
+ N_VGND_c_517_n N_VGND_c_518_n N_VGND_c_519_n PM_SKY130_FD_SC_LP__O32A_LP%VGND
cc_1 VNB N_B1_c_78_n 0.0277102f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=1.51
cc_2 VNB N_B1_c_79_n 0.0173502f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=1
cc_3 VNB N_B1_c_80_n 0.0568418f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.345
cc_4 VNB N_B1_c_81_n 0.00704122f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.965
cc_5 VNB B1 0.0106118f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_6 VNB N_B2_M1009_g 0.0409294f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=0.715
cc_7 VNB N_B2_c_112_n 0.0196567f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.295
cc_8 VNB N_B2_c_113_n 0.00466456f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A3_M1010_g 0.0404396f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=2.09
cc_10 VNB N_A3_c_160_n 0.0212378f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A3_c_161_n 0.00383048f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.345
cc_12 VNB N_A2_M1001_g 0.037931f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=2.09
cc_13 VNB N_A2_c_208_n 0.0277451f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A2_c_209_n 0.00169237f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A1_c_255_n 0.0143672f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.965
cc_16 VNB N_A1_c_256_n 0.0105822f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_17 VNB N_A1_c_257_n 0.0224048f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.345
cc_18 VNB N_A1_c_258_n 0.00179875f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.345
cc_19 VNB N_A1_c_259_n 0.017037f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_134_101#_c_303_n 0.0322311f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=0.715
cc_21 VNB N_A_134_101#_c_304_n 0.0194634f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_134_101#_c_305_n 0.00706051f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_134_101#_c_306_n 0.00111332f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_134_101#_c_307_n 0.0457067f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_134_101#_c_308_n 0.00328862f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_134_101#_c_309_n 0.00395228f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_134_101#_c_310_n 0.0358605f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_134_101#_c_311_n 5.9093e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VPWR_c_399_n 0.163682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_X_c_447_n 0.0265294f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.345
cc_31 VNB N_X_c_448_n 0.0359441f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_31_101#_c_470_n 0.0232649f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_33 VNB N_A_31_101#_c_471_n 0.0131157f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_31_101#_c_472_n 0.0106428f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_31_101#_c_473_n 0.00229875f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.665
cc_36 VNB N_VGND_c_512_n 0.00853868f $X=-0.19 $Y=-0.245 $X2=0.587 $Y2=1.345
cc_37 VNB N_VGND_c_513_n 0.0168596f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.965
cc_38 VNB N_VGND_c_514_n 0.00765741f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_515_n 0.0418815f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_516_n 0.0286633f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_517_n 0.247807f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_518_n 0.0063135f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_519_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VPB N_B1_c_83_n 0.0314439f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=2.09
cc_45 VPB N_B1_c_81_n 0.0206838f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=1.965
cc_46 VPB B1 0.0125773f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_47 VPB N_B2_c_114_n 0.0253887f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=2.09
cc_48 VPB N_B2_c_115_n 0.0105439f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=1.345
cc_49 VPB N_B2_c_112_n 0.0101722f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.295
cc_50 VPB N_B2_c_113_n 0.00265984f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_51 VPB N_A3_c_162_n 0.00833772f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=1.345
cc_52 VPB N_A3_c_163_n 0.0356281f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=1.965
cc_53 VPB N_A3_c_160_n 0.00982257f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_54 VPB N_A3_c_161_n 0.00307809f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.345
cc_55 VPB N_A2_c_210_n 0.0237548f $X=-0.19 $Y=1.655 $X2=0.595 $Y2=0.715
cc_56 VPB N_A2_c_211_n 0.0158071f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=1.345
cc_57 VPB N_A2_c_208_n 0.00494057f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_58 VPB N_A2_c_209_n 0.00315145f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_59 VPB N_A1_c_260_n 0.0247534f $X=-0.19 $Y=1.655 $X2=0.595 $Y2=0.715
cc_60 VPB N_A1_c_261_n 0.0127338f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_61 VPB N_A1_c_257_n 0.00845822f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.345
cc_62 VPB N_A1_c_258_n 0.00214181f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.345
cc_63 VPB N_A_134_101#_M1006_g 0.0434556f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_64 VPB N_A_134_101#_c_305_n 0.00949863f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_65 VPB N_A_134_101#_c_314_n 0.0179697f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_66 VPB N_A_134_101#_c_315_n 0.0034064f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_67 VPB N_A_134_101#_c_316_n 0.00209378f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_68 VPB N_A_134_101#_c_311_n 5.32916e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_69 VPB N_VPWR_c_400_n 0.012885f $X=-0.19 $Y=1.655 $X2=0.595 $Y2=0.715
cc_70 VPB N_VPWR_c_401_n 0.0449796f $X=-0.19 $Y=1.655 $X2=0.587 $Y2=1.345
cc_71 VPB N_VPWR_c_402_n 4.89148e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_72 VPB N_VPWR_c_403_n 0.0689942f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.345
cc_73 VPB N_VPWR_c_404_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_74 VPB N_VPWR_c_405_n 0.0192736f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_75 VPB N_VPWR_c_399_n 0.048444f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_76 VPB X 0.0523424f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_77 VPB N_X_c_448_n 0.012463f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_78 N_B1_c_83_n N_B2_c_114_n 0.0703131f $X=0.63 $Y=2.09 $X2=0 $Y2=0
cc_79 N_B1_c_78_n N_B2_M1009_g 0.0106545f $X=0.58 $Y=1.51 $X2=0 $Y2=0
cc_80 N_B1_c_79_n N_B2_M1009_g 0.0177818f $X=0.595 $Y=1 $X2=0 $Y2=0
cc_81 B1 N_B2_M1009_g 9.74994e-19 $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_82 N_B1_c_81_n N_B2_c_115_n 0.00727746f $X=0.63 $Y=1.965 $X2=0 $Y2=0
cc_83 N_B1_c_78_n N_B2_c_112_n 0.0180819f $X=0.58 $Y=1.51 $X2=0 $Y2=0
cc_84 N_B1_c_78_n N_B2_c_113_n 0.00426616f $X=0.58 $Y=1.51 $X2=0 $Y2=0
cc_85 N_B1_c_83_n N_B2_c_113_n 0.037737f $X=0.63 $Y=2.09 $X2=0 $Y2=0
cc_86 N_B1_c_81_n N_B2_c_113_n 0.017346f $X=0.63 $Y=1.965 $X2=0 $Y2=0
cc_87 B1 N_B2_c_113_n 0.027773f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_88 N_B1_c_79_n N_A_134_101#_c_306_n 0.00606129f $X=0.595 $Y=1 $X2=0 $Y2=0
cc_89 N_B1_c_78_n N_A_134_101#_c_308_n 0.00944202f $X=0.58 $Y=1.51 $X2=0 $Y2=0
cc_90 N_B1_c_79_n N_A_134_101#_c_308_n 0.00116628f $X=0.595 $Y=1 $X2=0 $Y2=0
cc_91 N_B1_c_83_n N_VPWR_c_401_n 0.0116609f $X=0.63 $Y=2.09 $X2=0 $Y2=0
cc_92 N_B1_c_80_n N_VPWR_c_401_n 0.00112012f $X=0.505 $Y=1.345 $X2=0 $Y2=0
cc_93 B1 N_VPWR_c_401_n 0.0156483f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_94 N_B1_c_83_n N_VPWR_c_403_n 0.007977f $X=0.63 $Y=2.09 $X2=0 $Y2=0
cc_95 N_B1_c_83_n N_VPWR_c_399_n 0.0129312f $X=0.63 $Y=2.09 $X2=0 $Y2=0
cc_96 N_B1_c_79_n N_A_31_101#_c_470_n 0.0113909f $X=0.595 $Y=1 $X2=0 $Y2=0
cc_97 N_B1_c_80_n N_A_31_101#_c_470_n 0.00348761f $X=0.505 $Y=1.345 $X2=0 $Y2=0
cc_98 B1 N_A_31_101#_c_470_n 0.0206308f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_99 N_B1_c_78_n N_A_31_101#_c_471_n 4.12567e-19 $X=0.58 $Y=1.51 $X2=0 $Y2=0
cc_100 N_B1_c_79_n N_A_31_101#_c_471_n 0.0113073f $X=0.595 $Y=1 $X2=0 $Y2=0
cc_101 N_B1_c_79_n N_A_31_101#_c_479_n 7.73341e-19 $X=0.595 $Y=1 $X2=0 $Y2=0
cc_102 N_B1_c_79_n N_VGND_c_515_n 7.10185e-19 $X=0.595 $Y=1 $X2=0 $Y2=0
cc_103 N_B2_M1009_g N_A3_M1010_g 0.0340522f $X=1.105 $Y=0.655 $X2=0 $Y2=0
cc_104 N_B2_c_115_n N_A3_c_162_n 0.00434254f $X=1.12 $Y=1.965 $X2=0 $Y2=0
cc_105 N_B2_c_112_n N_A3_c_162_n 8.00009e-19 $X=1.06 $Y=1.59 $X2=0 $Y2=0
cc_106 N_B2_c_113_n N_A3_c_162_n 0.00409407f $X=1.06 $Y=1.59 $X2=0 $Y2=0
cc_107 N_B2_c_114_n N_A3_c_163_n 0.0245676f $X=1.12 $Y=2.09 $X2=0 $Y2=0
cc_108 N_B2_c_113_n N_A3_c_163_n 4.60479e-19 $X=1.06 $Y=1.59 $X2=0 $Y2=0
cc_109 N_B2_M1009_g N_A3_c_160_n 0.00155278f $X=1.105 $Y=0.655 $X2=0 $Y2=0
cc_110 N_B2_c_112_n N_A3_c_160_n 0.0182822f $X=1.06 $Y=1.59 $X2=0 $Y2=0
cc_111 N_B2_c_113_n N_A3_c_160_n 0.00104195f $X=1.06 $Y=1.59 $X2=0 $Y2=0
cc_112 N_B2_c_112_n N_A3_c_161_n 0.0012808f $X=1.06 $Y=1.59 $X2=0 $Y2=0
cc_113 N_B2_c_113_n N_A3_c_161_n 0.0241046f $X=1.06 $Y=1.59 $X2=0 $Y2=0
cc_114 N_B2_M1009_g N_A_134_101#_c_306_n 0.00449692f $X=1.105 $Y=0.655 $X2=0
+ $Y2=0
cc_115 N_B2_M1009_g N_A_134_101#_c_307_n 0.0129694f $X=1.105 $Y=0.655 $X2=0
+ $Y2=0
cc_116 N_B2_c_112_n N_A_134_101#_c_307_n 6.25529e-19 $X=1.06 $Y=1.59 $X2=0 $Y2=0
cc_117 N_B2_c_113_n N_A_134_101#_c_307_n 0.0132469f $X=1.06 $Y=1.59 $X2=0 $Y2=0
cc_118 N_B2_c_112_n N_A_134_101#_c_308_n 5.77235e-19 $X=1.06 $Y=1.59 $X2=0 $Y2=0
cc_119 N_B2_c_113_n N_A_134_101#_c_308_n 0.0211338f $X=1.06 $Y=1.59 $X2=0 $Y2=0
cc_120 N_B2_c_114_n N_A_134_101#_c_327_n 0.0100368f $X=1.12 $Y=2.09 $X2=0 $Y2=0
cc_121 N_B2_c_113_n N_A_134_101#_c_327_n 0.0579085f $X=1.06 $Y=1.59 $X2=0 $Y2=0
cc_122 N_B2_c_114_n N_A_134_101#_c_315_n 0.00136229f $X=1.12 $Y=2.09 $X2=0 $Y2=0
cc_123 N_B2_c_113_n N_A_134_101#_c_315_n 0.0142558f $X=1.06 $Y=1.59 $X2=0 $Y2=0
cc_124 N_B2_c_113_n N_VPWR_c_401_n 0.0621272f $X=1.06 $Y=1.59 $X2=0 $Y2=0
cc_125 N_B2_c_114_n N_VPWR_c_403_n 0.00682486f $X=1.12 $Y=2.09 $X2=0 $Y2=0
cc_126 N_B2_c_113_n N_VPWR_c_403_n 0.0169742f $X=1.06 $Y=1.59 $X2=0 $Y2=0
cc_127 N_B2_c_114_n N_VPWR_c_399_n 0.00915809f $X=1.12 $Y=2.09 $X2=0 $Y2=0
cc_128 N_B2_c_113_n N_VPWR_c_399_n 0.0193652f $X=1.06 $Y=1.59 $X2=0 $Y2=0
cc_129 N_B2_c_113_n A_151_419# 0.00175001f $X=1.06 $Y=1.59 $X2=-0.19 $Y2=-0.245
cc_130 N_B2_M1009_g N_A_31_101#_c_471_n 0.0108088f $X=1.105 $Y=0.655 $X2=0 $Y2=0
cc_131 N_B2_M1009_g N_A_31_101#_c_479_n 0.00372244f $X=1.105 $Y=0.655 $X2=0
+ $Y2=0
cc_132 N_B2_M1009_g N_A_31_101#_c_482_n 0.00214195f $X=1.105 $Y=0.655 $X2=0
+ $Y2=0
cc_133 N_B2_M1009_g N_VGND_c_515_n 8.47083e-19 $X=1.105 $Y=0.655 $X2=0 $Y2=0
cc_134 N_A3_M1010_g N_A2_M1001_g 0.0269111f $X=1.535 $Y=0.655 $X2=0 $Y2=0
cc_135 N_A3_c_163_n N_A2_c_210_n 0.0397239f $X=1.747 $Y=2.02 $X2=0 $Y2=0
cc_136 N_A3_c_163_n N_A2_c_211_n 0.0397239f $X=1.747 $Y=2.02 $X2=0 $Y2=0
cc_137 N_A3_c_160_n N_A2_c_211_n 0.00759044f $X=1.6 $Y=1.56 $X2=0 $Y2=0
cc_138 N_A3_c_161_n N_A2_c_211_n 3.28797e-19 $X=1.6 $Y=1.56 $X2=0 $Y2=0
cc_139 N_A3_M1010_g N_A2_c_208_n 0.00234323f $X=1.535 $Y=0.655 $X2=0 $Y2=0
cc_140 N_A3_c_160_n N_A2_c_208_n 0.0165914f $X=1.6 $Y=1.56 $X2=0 $Y2=0
cc_141 N_A3_c_161_n N_A2_c_208_n 0.00151402f $X=1.6 $Y=1.56 $X2=0 $Y2=0
cc_142 N_A3_M1010_g N_A2_c_209_n 3.79646e-19 $X=1.535 $Y=0.655 $X2=0 $Y2=0
cc_143 N_A3_c_160_n N_A2_c_209_n 7.333e-19 $X=1.6 $Y=1.56 $X2=0 $Y2=0
cc_144 N_A3_c_161_n N_A2_c_209_n 0.0298899f $X=1.6 $Y=1.56 $X2=0 $Y2=0
cc_145 N_A3_M1010_g N_A_134_101#_c_307_n 0.0116706f $X=1.535 $Y=0.655 $X2=0
+ $Y2=0
cc_146 N_A3_c_160_n N_A_134_101#_c_307_n 0.00115733f $X=1.6 $Y=1.56 $X2=0 $Y2=0
cc_147 N_A3_c_161_n N_A_134_101#_c_307_n 0.0203312f $X=1.6 $Y=1.56 $X2=0 $Y2=0
cc_148 N_A3_c_163_n N_A_134_101#_c_327_n 0.0211155f $X=1.747 $Y=2.02 $X2=0 $Y2=0
cc_149 N_A3_c_163_n N_A_134_101#_c_314_n 0.0201408f $X=1.747 $Y=2.02 $X2=0 $Y2=0
cc_150 N_A3_c_161_n N_A_134_101#_c_314_n 0.00973705f $X=1.6 $Y=1.56 $X2=0 $Y2=0
cc_151 N_A3_c_163_n N_A_134_101#_c_315_n 0.00292465f $X=1.747 $Y=2.02 $X2=0
+ $Y2=0
cc_152 N_A3_c_160_n N_A_134_101#_c_315_n 0.0012091f $X=1.6 $Y=1.56 $X2=0 $Y2=0
cc_153 N_A3_c_161_n N_A_134_101#_c_315_n 0.0185376f $X=1.6 $Y=1.56 $X2=0 $Y2=0
cc_154 N_A3_c_163_n N_VPWR_c_403_n 0.00939541f $X=1.747 $Y=2.02 $X2=0 $Y2=0
cc_155 N_A3_c_163_n N_VPWR_c_399_n 0.0163858f $X=1.747 $Y=2.02 $X2=0 $Y2=0
cc_156 N_A3_M1010_g N_A_31_101#_c_471_n 0.0030617f $X=1.535 $Y=0.655 $X2=0 $Y2=0
cc_157 N_A3_M1010_g N_A_31_101#_c_479_n 0.00394039f $X=1.535 $Y=0.655 $X2=0
+ $Y2=0
cc_158 N_A3_M1010_g N_A_31_101#_c_485_n 0.00897052f $X=1.535 $Y=0.655 $X2=0
+ $Y2=0
cc_159 N_A3_M1010_g N_A_31_101#_c_482_n 7.38868e-19 $X=1.535 $Y=0.655 $X2=0
+ $Y2=0
cc_160 N_A3_M1010_g N_A_31_101#_c_473_n 9.02326e-19 $X=1.535 $Y=0.655 $X2=0
+ $Y2=0
cc_161 N_A3_M1010_g N_VGND_c_512_n 0.00127271f $X=1.535 $Y=0.655 $X2=0 $Y2=0
cc_162 N_A3_M1010_g N_VGND_c_515_n 0.00348245f $X=1.535 $Y=0.655 $X2=0 $Y2=0
cc_163 N_A3_M1010_g N_VGND_c_517_n 0.004351f $X=1.535 $Y=0.655 $X2=0 $Y2=0
cc_164 N_A2_c_210_n N_A1_c_260_n 0.074393f $X=2.245 $Y=2.09 $X2=0 $Y2=0
cc_165 N_A2_M1001_g N_A1_c_255_n 0.0192187f $X=2.125 $Y=0.655 $X2=0 $Y2=0
cc_166 N_A2_c_211_n N_A1_c_261_n 0.00973769f $X=2.245 $Y=1.965 $X2=0 $Y2=0
cc_167 N_A2_c_211_n N_A1_c_257_n 0.00331863f $X=2.245 $Y=1.965 $X2=0 $Y2=0
cc_168 N_A2_c_208_n N_A1_c_257_n 0.0161493f $X=2.14 $Y=1.495 $X2=0 $Y2=0
cc_169 N_A2_c_209_n N_A1_c_257_n 0.00132255f $X=2.14 $Y=1.495 $X2=0 $Y2=0
cc_170 N_A2_c_211_n N_A1_c_258_n 2.73669e-19 $X=2.245 $Y=1.965 $X2=0 $Y2=0
cc_171 N_A2_c_208_n N_A1_c_258_n 9.2297e-19 $X=2.14 $Y=1.495 $X2=0 $Y2=0
cc_172 N_A2_c_209_n N_A1_c_258_n 0.0251343f $X=2.14 $Y=1.495 $X2=0 $Y2=0
cc_173 N_A2_M1001_g N_A1_c_259_n 0.00959448f $X=2.125 $Y=0.655 $X2=0 $Y2=0
cc_174 N_A2_c_208_n N_A1_c_259_n 0.00360906f $X=2.14 $Y=1.495 $X2=0 $Y2=0
cc_175 N_A2_c_209_n N_A1_c_259_n 4.18638e-19 $X=2.14 $Y=1.495 $X2=0 $Y2=0
cc_176 N_A2_M1001_g N_A_134_101#_c_307_n 0.0114004f $X=2.125 $Y=0.655 $X2=0
+ $Y2=0
cc_177 N_A2_c_208_n N_A_134_101#_c_307_n 0.00123291f $X=2.14 $Y=1.495 $X2=0
+ $Y2=0
cc_178 N_A2_c_209_n N_A_134_101#_c_307_n 0.0237277f $X=2.14 $Y=1.495 $X2=0 $Y2=0
cc_179 N_A2_c_210_n N_A_134_101#_c_327_n 0.00405544f $X=2.245 $Y=2.09 $X2=0
+ $Y2=0
cc_180 N_A2_c_210_n N_A_134_101#_c_314_n 0.0191967f $X=2.245 $Y=2.09 $X2=0 $Y2=0
cc_181 N_A2_c_211_n N_A_134_101#_c_314_n 0.00215083f $X=2.245 $Y=1.965 $X2=0
+ $Y2=0
cc_182 N_A2_c_208_n N_A_134_101#_c_314_n 8.24837e-19 $X=2.14 $Y=1.495 $X2=0
+ $Y2=0
cc_183 N_A2_c_209_n N_A_134_101#_c_314_n 0.024499f $X=2.14 $Y=1.495 $X2=0 $Y2=0
cc_184 N_A2_c_210_n N_VPWR_c_402_n 0.00429931f $X=2.245 $Y=2.09 $X2=0 $Y2=0
cc_185 N_A2_c_210_n N_VPWR_c_403_n 0.00975641f $X=2.245 $Y=2.09 $X2=0 $Y2=0
cc_186 N_A2_c_210_n N_VPWR_c_399_n 0.0170051f $X=2.245 $Y=2.09 $X2=0 $Y2=0
cc_187 N_A2_M1001_g N_A_31_101#_c_479_n 8.13476e-19 $X=2.125 $Y=0.655 $X2=0
+ $Y2=0
cc_188 N_A2_M1001_g N_A_31_101#_c_485_n 0.00951876f $X=2.125 $Y=0.655 $X2=0
+ $Y2=0
cc_189 N_A2_M1001_g N_A_31_101#_c_473_n 0.00556924f $X=2.125 $Y=0.655 $X2=0
+ $Y2=0
cc_190 N_A2_M1001_g N_VGND_c_512_n 0.00195394f $X=2.125 $Y=0.655 $X2=0 $Y2=0
cc_191 N_A2_M1001_g N_VGND_c_513_n 0.00398919f $X=2.125 $Y=0.655 $X2=0 $Y2=0
cc_192 N_A2_M1001_g N_VGND_c_514_n 4.55413e-19 $X=2.125 $Y=0.655 $X2=0 $Y2=0
cc_193 N_A2_M1001_g N_VGND_c_517_n 0.0052212f $X=2.125 $Y=0.655 $X2=0 $Y2=0
cc_194 N_A1_c_255_n N_A_134_101#_c_303_n 0.0126598f $X=2.587 $Y=0.94 $X2=0 $Y2=0
cc_195 N_A1_c_260_n N_A_134_101#_M1006_g 0.024325f $X=2.735 $Y=2.075 $X2=0 $Y2=0
cc_196 N_A1_c_261_n N_A_134_101#_M1006_g 0.0055728f $X=2.735 $Y=1.95 $X2=0 $Y2=0
cc_197 N_A1_c_256_n N_A_134_101#_c_304_n 0.0098589f $X=2.587 $Y=1.09 $X2=0 $Y2=0
cc_198 N_A1_c_261_n N_A_134_101#_c_305_n 6.1362e-19 $X=2.735 $Y=1.95 $X2=0 $Y2=0
cc_199 N_A1_c_256_n N_A_134_101#_c_307_n 0.0113299f $X=2.587 $Y=1.09 $X2=0 $Y2=0
cc_200 N_A1_c_257_n N_A_134_101#_c_307_n 0.00106681f $X=2.68 $Y=1.56 $X2=0 $Y2=0
cc_201 N_A1_c_258_n N_A_134_101#_c_307_n 0.0184631f $X=2.68 $Y=1.56 $X2=0 $Y2=0
cc_202 N_A1_c_259_n N_A_134_101#_c_307_n 0.00493169f $X=2.68 $Y=1.395 $X2=0
+ $Y2=0
cc_203 N_A1_c_260_n N_A_134_101#_c_314_n 0.021055f $X=2.735 $Y=2.075 $X2=0 $Y2=0
cc_204 N_A1_c_257_n N_A_134_101#_c_314_n 6.55073e-19 $X=2.68 $Y=1.56 $X2=0 $Y2=0
cc_205 N_A1_c_258_n N_A_134_101#_c_314_n 0.023873f $X=2.68 $Y=1.56 $X2=0 $Y2=0
cc_206 N_A1_c_257_n N_A_134_101#_c_309_n 0.00188269f $X=2.68 $Y=1.56 $X2=0 $Y2=0
cc_207 N_A1_c_258_n N_A_134_101#_c_309_n 0.0293695f $X=2.68 $Y=1.56 $X2=0 $Y2=0
cc_208 N_A1_c_259_n N_A_134_101#_c_309_n 0.00499481f $X=2.68 $Y=1.395 $X2=0
+ $Y2=0
cc_209 N_A1_c_257_n N_A_134_101#_c_310_n 0.0206365f $X=2.68 $Y=1.56 $X2=0 $Y2=0
cc_210 N_A1_c_258_n N_A_134_101#_c_310_n 3.93466e-19 $X=2.68 $Y=1.56 $X2=0 $Y2=0
cc_211 N_A1_c_259_n N_A_134_101#_c_310_n 0.0092569f $X=2.68 $Y=1.395 $X2=0 $Y2=0
cc_212 N_A1_c_261_n N_A_134_101#_c_316_n 0.00329356f $X=2.735 $Y=1.95 $X2=0
+ $Y2=0
cc_213 N_A1_c_260_n N_VPWR_c_402_n 0.021829f $X=2.735 $Y=2.075 $X2=0 $Y2=0
cc_214 N_A1_c_260_n N_VPWR_c_403_n 0.008763f $X=2.735 $Y=2.075 $X2=0 $Y2=0
cc_215 N_A1_c_260_n N_VPWR_c_399_n 0.0144563f $X=2.735 $Y=2.075 $X2=0 $Y2=0
cc_216 N_A1_c_260_n X 9.38255e-19 $X=2.735 $Y=2.075 $X2=0 $Y2=0
cc_217 N_A1_c_255_n N_VGND_c_513_n 0.00435433f $X=2.587 $Y=0.94 $X2=0 $Y2=0
cc_218 N_A1_c_255_n N_VGND_c_514_n 0.00830046f $X=2.587 $Y=0.94 $X2=0 $Y2=0
cc_219 N_A1_c_256_n N_VGND_c_514_n 0.00165177f $X=2.587 $Y=1.09 $X2=0 $Y2=0
cc_220 N_A1_c_255_n N_VGND_c_517_n 0.0043858f $X=2.587 $Y=0.94 $X2=0 $Y2=0
cc_221 N_A_134_101#_c_314_n N_VPWR_M1002_d 0.001936f $X=3.025 $Y=2.045 $X2=0
+ $Y2=0
cc_222 N_A_134_101#_M1006_g N_VPWR_c_402_n 0.0198402f $X=3.275 $Y=2.595 $X2=0
+ $Y2=0
cc_223 N_A_134_101#_c_305_n N_VPWR_c_402_n 2.47575e-19 $X=3.237 $Y=1.74 $X2=0
+ $Y2=0
cc_224 N_A_134_101#_c_314_n N_VPWR_c_402_n 0.0170535f $X=3.025 $Y=2.045 $X2=0
+ $Y2=0
cc_225 N_A_134_101#_c_327_n N_VPWR_c_403_n 0.014447f $X=1.49 $Y=2.24 $X2=0 $Y2=0
cc_226 N_A_134_101#_M1006_g N_VPWR_c_405_n 0.00879225f $X=3.275 $Y=2.595 $X2=0
+ $Y2=0
cc_227 N_A_134_101#_M1007_d N_VPWR_c_399_n 0.00869929f $X=1.245 $Y=2.095 $X2=0
+ $Y2=0
cc_228 N_A_134_101#_M1006_g N_VPWR_c_399_n 0.0151595f $X=3.275 $Y=2.595 $X2=0
+ $Y2=0
cc_229 N_A_134_101#_c_327_n N_VPWR_c_399_n 0.00941258f $X=1.49 $Y=2.24 $X2=0
+ $Y2=0
cc_230 N_A_134_101#_c_314_n A_376_419# 0.0048076f $X=3.025 $Y=2.045 $X2=-0.19
+ $Y2=-0.245
cc_231 N_A_134_101#_c_314_n A_474_419# 0.0048076f $X=3.025 $Y=2.045 $X2=-0.19
+ $Y2=-0.245
cc_232 N_A_134_101#_c_303_n N_X_c_447_n 0.011792f $X=2.985 $Y=0.94 $X2=0 $Y2=0
cc_233 N_A_134_101#_M1006_g X 0.0303836f $X=3.275 $Y=2.595 $X2=0 $Y2=0
cc_234 N_A_134_101#_c_305_n X 9.57316e-19 $X=3.237 $Y=1.74 $X2=0 $Y2=0
cc_235 N_A_134_101#_c_314_n X 0.0130043f $X=3.025 $Y=2.045 $X2=0 $Y2=0
cc_236 N_A_134_101#_c_316_n X 0.00271538f $X=3.11 $Y=1.96 $X2=0 $Y2=0
cc_237 N_A_134_101#_c_311_n X 6.45782e-19 $X=3.205 $Y=1.74 $X2=0 $Y2=0
cc_238 N_A_134_101#_c_303_n N_X_c_448_n 0.020136f $X=2.985 $Y=0.94 $X2=0 $Y2=0
cc_239 N_A_134_101#_M1006_g N_X_c_448_n 0.00303969f $X=3.275 $Y=2.595 $X2=0
+ $Y2=0
cc_240 N_A_134_101#_c_307_n N_X_c_448_n 0.0100814f $X=3.025 $Y=1.065 $X2=0 $Y2=0
cc_241 N_A_134_101#_c_309_n N_X_c_448_n 0.0426092f $X=3.22 $Y=1.235 $X2=0 $Y2=0
cc_242 N_A_134_101#_c_316_n N_X_c_448_n 0.00519041f $X=3.11 $Y=1.96 $X2=0 $Y2=0
cc_243 N_A_134_101#_c_306_n N_A_31_101#_c_470_n 0.0125869f $X=0.81 $Y=0.78 $X2=0
+ $Y2=0
cc_244 N_A_134_101#_c_306_n N_A_31_101#_c_471_n 0.0215434f $X=0.81 $Y=0.78 $X2=0
+ $Y2=0
cc_245 N_A_134_101#_c_307_n N_A_31_101#_c_471_n 0.00507493f $X=3.025 $Y=1.065
+ $X2=0 $Y2=0
cc_246 N_A_134_101#_c_307_n N_A_31_101#_c_485_n 0.0434123f $X=3.025 $Y=1.065
+ $X2=0 $Y2=0
cc_247 N_A_134_101#_c_307_n N_A_31_101#_c_482_n 0.0205422f $X=3.025 $Y=1.065
+ $X2=0 $Y2=0
cc_248 N_A_134_101#_c_307_n N_A_31_101#_c_473_n 0.0162934f $X=3.025 $Y=1.065
+ $X2=0 $Y2=0
cc_249 N_A_134_101#_c_303_n N_VGND_c_514_n 0.0118205f $X=2.985 $Y=0.94 $X2=0
+ $Y2=0
cc_250 N_A_134_101#_c_307_n N_VGND_c_514_n 0.0204691f $X=3.025 $Y=1.065 $X2=0
+ $Y2=0
cc_251 N_A_134_101#_c_303_n N_VGND_c_516_n 0.00936557f $X=2.985 $Y=0.94 $X2=0
+ $Y2=0
cc_252 N_A_134_101#_c_303_n N_VGND_c_517_n 0.009607f $X=2.985 $Y=0.94 $X2=0
+ $Y2=0
cc_253 N_VPWR_c_399_n A_151_419# 0.00219029f $X=3.6 $Y=3.33 $X2=-0.19 $Y2=-0.245
cc_254 N_VPWR_c_399_n A_376_419# 0.010279f $X=3.6 $Y=3.33 $X2=-0.19 $Y2=-0.245
cc_255 N_VPWR_c_399_n A_474_419# 0.010279f $X=3.6 $Y=3.33 $X2=-0.19 $Y2=-0.245
cc_256 N_VPWR_c_399_n N_X_M1006_d 0.0023218f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_257 N_VPWR_c_402_n X 0.0481682f $X=3 $Y=2.475 $X2=0 $Y2=0
cc_258 N_VPWR_c_405_n X 0.0217808f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_259 N_VPWR_c_399_n X 0.0136688f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_260 N_X_c_447_n N_VGND_c_514_n 0.0125752f $X=3.56 $Y=0.655 $X2=0 $Y2=0
cc_261 N_X_c_447_n N_VGND_c_516_n 0.0113525f $X=3.56 $Y=0.655 $X2=0 $Y2=0
cc_262 N_X_c_447_n N_VGND_c_517_n 0.0117944f $X=3.56 $Y=0.655 $X2=0 $Y2=0
cc_263 N_A_31_101#_c_485_n N_VGND_M1010_d 0.00758216f $X=2.175 $Y=0.715
+ $X2=-0.19 $Y2=-0.245
cc_264 N_A_31_101#_c_471_n N_VGND_c_512_n 0.0138885f $X=1.155 $Y=0.35 $X2=0
+ $Y2=0
cc_265 N_A_31_101#_c_479_n N_VGND_c_512_n 8.61411e-19 $X=1.32 $Y=0.61 $X2=0
+ $Y2=0
cc_266 N_A_31_101#_c_485_n N_VGND_c_512_n 0.0235796f $X=2.175 $Y=0.715 $X2=0
+ $Y2=0
cc_267 N_A_31_101#_c_473_n N_VGND_c_512_n 0.00161794f $X=2.34 $Y=0.61 $X2=0
+ $Y2=0
cc_268 N_A_31_101#_c_485_n N_VGND_c_513_n 0.00260066f $X=2.175 $Y=0.715 $X2=0
+ $Y2=0
cc_269 N_A_31_101#_c_473_n N_VGND_c_513_n 0.00808182f $X=2.34 $Y=0.61 $X2=0
+ $Y2=0
cc_270 N_A_31_101#_c_473_n N_VGND_c_514_n 0.0141685f $X=2.34 $Y=0.61 $X2=0 $Y2=0
cc_271 N_A_31_101#_c_471_n N_VGND_c_515_n 0.0636368f $X=1.155 $Y=0.35 $X2=0
+ $Y2=0
cc_272 N_A_31_101#_c_472_n N_VGND_c_515_n 0.0222501f $X=0.465 $Y=0.35 $X2=0
+ $Y2=0
cc_273 N_A_31_101#_c_485_n N_VGND_c_515_n 0.00259405f $X=2.175 $Y=0.715 $X2=0
+ $Y2=0
cc_274 N_A_31_101#_c_471_n N_VGND_c_517_n 0.0384659f $X=1.155 $Y=0.35 $X2=0
+ $Y2=0
cc_275 N_A_31_101#_c_472_n N_VGND_c_517_n 0.0127687f $X=0.465 $Y=0.35 $X2=0
+ $Y2=0
cc_276 N_A_31_101#_c_485_n N_VGND_c_517_n 0.011656f $X=2.175 $Y=0.715 $X2=0
+ $Y2=0
cc_277 N_A_31_101#_c_473_n N_VGND_c_517_n 0.00852167f $X=2.34 $Y=0.61 $X2=0
+ $Y2=0
