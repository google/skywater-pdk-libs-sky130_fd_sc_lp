* File: sky130_fd_sc_lp__a311o_4.pex.spice
* Created: Fri Aug 28 09:57:45 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A311O_4%C1 3 7 11 15 17 18 26
r47 25 26 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=0.48 $Y=1.375
+ $X2=0.91 $Y2=1.375
r48 22 25 27.1035 $w=3.3e-07 $l=1.55e-07 $layer=POLY_cond $X=0.325 $Y=1.375
+ $X2=0.48 $Y2=1.375
r49 17 18 12.3595 $w=3.43e-07 $l=3.7e-07 $layer=LI1_cond $X=0.257 $Y=1.295
+ $X2=0.257 $Y2=1.665
r50 17 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.325
+ $Y=1.375 $X2=0.325 $Y2=1.375
r51 13 26 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.91 $Y=1.54
+ $X2=0.91 $Y2=1.375
r52 13 15 474.309 $w=1.5e-07 $l=9.25e-07 $layer=POLY_cond $X=0.91 $Y=1.54
+ $X2=0.91 $Y2=2.465
r53 9 26 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.91 $Y=1.21
+ $X2=0.91 $Y2=1.375
r54 9 11 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=0.91 $Y=1.21
+ $X2=0.91 $Y2=0.655
r55 5 25 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.48 $Y=1.54
+ $X2=0.48 $Y2=1.375
r56 5 7 474.309 $w=1.5e-07 $l=9.25e-07 $layer=POLY_cond $X=0.48 $Y=1.54 $X2=0.48
+ $Y2=2.465
r57 1 25 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.48 $Y=1.21
+ $X2=0.48 $Y2=1.375
r58 1 3 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=0.48 $Y=1.21 $X2=0.48
+ $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__A311O_4%B1 3 7 9 11 15 17 18 26
c54 7 0 1.87962e-19 $X=1.38 $Y=0.655
r55 25 26 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.7 $Y=1.5
+ $X2=1.7 $Y2=1.5
r56 18 26 0.688026 $w=3.33e-07 $l=2e-08 $layer=LI1_cond $X=1.68 $Y=1.582 $X2=1.7
+ $Y2=1.582
r57 17 18 16.5126 $w=3.33e-07 $l=4.8e-07 $layer=LI1_cond $X=1.2 $Y=1.582
+ $X2=1.68 $Y2=1.582
r58 13 15 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=1.81 $Y=1.665 $X2=1.81
+ $Y2=2.465
r59 9 13 24.2915 $w=1.5e-07 $l=1.88e-07 $layer=POLY_cond $X=1.81 $Y=1.477
+ $X2=1.81 $Y2=1.665
r60 9 25 16.3138 $w=3.75e-07 $l=1.1e-07 $layer=POLY_cond $X=1.81 $Y=1.477
+ $X2=1.7 $Y2=1.477
r61 9 11 325.606 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.81 $Y=1.29
+ $X2=1.81 $Y2=0.655
r62 5 25 47.4585 $w=3.75e-07 $l=3.2e-07 $layer=POLY_cond $X=1.38 $Y=1.477
+ $X2=1.7 $Y2=1.477
r63 5 21 5.93231 $w=3.75e-07 $l=4e-08 $layer=POLY_cond $X=1.38 $Y=1.477 $X2=1.34
+ $Y2=1.477
r64 5 7 325.606 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.38 $Y=1.29 $X2=1.38
+ $Y2=0.655
r65 1 21 24.2915 $w=1.5e-07 $l=1.88e-07 $layer=POLY_cond $X=1.34 $Y=1.665
+ $X2=1.34 $Y2=1.477
r66 1 3 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=1.34 $Y=1.665 $X2=1.34
+ $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__A311O_4%A_111_47# 1 2 3 4 15 19 23 27 31 35 37 39 40
+ 41 44 48 52 54 58 60 62 65 71 74 75 76 79 82 84 85 86 91 93 99
c200 52 0 1.87962e-19 $X=0.695 $Y=2.095
c201 40 0 1.45841e-19 $X=4.465 $Y=1.625
r202 97 99 13.4452 $w=2.98e-07 $l=3.5e-07 $layer=LI1_cond $X=6.63 $Y=1.495
+ $X2=6.98 $Y2=1.495
r203 93 95 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=4.65 $Y=2.005
+ $X2=4.65 $Y2=2.27
r204 92 101 63.9691 $w=3.24e-07 $l=4.3e-07 $layer=POLY_cond $X=2.68 $Y=1.492
+ $X2=2.25 $Y2=1.492
r205 91 92 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.68
+ $Y=1.45 $X2=2.68 $Y2=1.45
r206 80 99 0.126616 $w=3.3e-07 $l=1.5e-07 $layer=LI1_cond $X=6.98 $Y=1.345
+ $X2=6.98 $Y2=1.495
r207 80 82 23.2235 $w=3.28e-07 $l=6.65e-07 $layer=LI1_cond $X=6.98 $Y=1.345
+ $X2=6.98 $Y2=0.68
r208 78 97 4.061 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=6.63 $Y=1.645 $X2=6.63
+ $Y2=1.495
r209 78 79 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=6.63 $Y=1.645
+ $X2=6.63 $Y2=1.92
r210 77 93 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.735 $Y=2.005
+ $X2=4.65 $Y2=2.005
r211 76 79 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.545 $Y=2.005
+ $X2=6.63 $Y2=1.92
r212 76 77 118.086 $w=1.68e-07 $l=1.81e-06 $layer=LI1_cond $X=6.545 $Y=2.005
+ $X2=4.735 $Y2=2.005
r213 74 95 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.565 $Y=2.27
+ $X2=4.65 $Y2=2.27
r214 74 75 114.497 $w=1.68e-07 $l=1.755e-06 $layer=LI1_cond $X=4.565 $Y=2.27
+ $X2=2.81 $Y2=2.27
r215 72 109 32.7284 $w=3.24e-07 $l=2.2e-07 $layer=POLY_cond $X=3.7 $Y=1.492
+ $X2=3.92 $Y2=1.492
r216 72 107 23.8025 $w=3.24e-07 $l=1.6e-07 $layer=POLY_cond $X=3.7 $Y=1.492
+ $X2=3.54 $Y2=1.492
r217 71 72 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=3.7
+ $Y=1.45 $X2=3.7 $Y2=1.45
r218 69 105 13.3889 $w=3.24e-07 $l=9e-08 $layer=POLY_cond $X=3.02 $Y=1.492
+ $X2=3.11 $Y2=1.492
r219 68 71 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=3.02 $Y=1.45
+ $X2=3.7 $Y2=1.45
r220 68 69 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=3.02
+ $Y=1.45 $X2=3.02 $Y2=1.45
r221 66 91 4.60183 $w=1.95e-07 $l=9.66954e-08 $layer=LI1_cond $X=2.81 $Y=1.45
+ $X2=2.725 $Y2=1.475
r222 66 68 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=2.81 $Y=1.45
+ $X2=3.02 $Y2=1.45
r223 65 75 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.725 $Y=2.185
+ $X2=2.81 $Y2=2.27
r224 64 91 1.84097 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=2.725 $Y=1.585
+ $X2=2.725 $Y2=1.475
r225 64 65 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=2.725 $Y=1.585
+ $X2=2.725 $Y2=2.185
r226 63 86 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=2.12 $Y=1.475
+ $X2=2.12 $Y2=1.16
r227 62 91 4.60183 $w=1.95e-07 $l=8.5e-08 $layer=LI1_cond $X=2.64 $Y=1.475
+ $X2=2.725 $Y2=1.475
r228 62 63 22.7869 $w=2.18e-07 $l=4.35e-07 $layer=LI1_cond $X=2.64 $Y=1.475
+ $X2=2.205 $Y2=1.475
r229 61 85 6.25164 $w=1.7e-07 $l=1.08e-07 $layer=LI1_cond $X=1.69 $Y=1.16
+ $X2=1.582 $Y2=1.16
r230 60 86 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.035 $Y=1.16
+ $X2=2.12 $Y2=1.16
r231 60 61 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=2.035 $Y=1.16
+ $X2=1.69 $Y2=1.16
r232 56 85 0.512231 $w=2.15e-07 $l=8.5e-08 $layer=LI1_cond $X=1.582 $Y=1.075
+ $X2=1.582 $Y2=1.16
r233 56 58 35.1093 $w=2.13e-07 $l=6.55e-07 $layer=LI1_cond $X=1.582 $Y=1.075
+ $X2=1.582 $Y2=0.42
r234 55 84 1.88765 $w=1.7e-07 $l=1.03e-07 $layer=LI1_cond $X=0.805 $Y=1.16
+ $X2=0.702 $Y2=1.16
r235 54 85 6.25164 $w=1.7e-07 $l=1.07e-07 $layer=LI1_cond $X=1.475 $Y=1.16
+ $X2=1.582 $Y2=1.16
r236 54 55 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.475 $Y=1.16
+ $X2=0.805 $Y2=1.16
r237 50 84 4.55203 $w=1.97e-07 $l=8.84308e-08 $layer=LI1_cond $X=0.695 $Y=1.245
+ $X2=0.702 $Y2=1.16
r238 50 52 49.6172 $w=1.88e-07 $l=8.5e-07 $layer=LI1_cond $X=0.695 $Y=1.245
+ $X2=0.695 $Y2=2.095
r239 46 84 4.55203 $w=1.97e-07 $l=8.5e-08 $layer=LI1_cond $X=0.702 $Y=1.075
+ $X2=0.702 $Y2=1.16
r240 46 48 35.4368 $w=2.03e-07 $l=6.55e-07 $layer=LI1_cond $X=0.702 $Y=1.075
+ $X2=0.702 $Y2=0.42
r241 42 44 392.266 $w=1.5e-07 $l=7.65e-07 $layer=POLY_cond $X=4.54 $Y=1.7
+ $X2=4.54 $Y2=2.465
r242 41 109 25.1772 $w=3.24e-07 $l=1.66325e-07 $layer=POLY_cond $X=3.995
+ $Y=1.625 $X2=3.92 $Y2=1.492
r243 40 42 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.465 $Y=1.625
+ $X2=4.54 $Y2=1.7
r244 40 41 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=4.465 $Y=1.625
+ $X2=3.995 $Y2=1.625
r245 37 109 20.7868 $w=1.5e-07 $l=2.08e-07 $layer=POLY_cond $X=3.92 $Y=1.7
+ $X2=3.92 $Y2=1.492
r246 37 39 226.54 $w=1.5e-07 $l=7.05e-07 $layer=POLY_cond $X=3.92 $Y=1.7
+ $X2=3.92 $Y2=2.405
r247 33 107 20.7868 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.54 $Y=1.285
+ $X2=3.54 $Y2=1.492
r248 33 35 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=3.54 $Y=1.285
+ $X2=3.54 $Y2=0.655
r249 29 107 25.2901 $w=3.24e-07 $l=1.7e-07 $layer=POLY_cond $X=3.37 $Y=1.492
+ $X2=3.54 $Y2=1.492
r250 29 105 38.679 $w=3.24e-07 $l=2.6e-07 $layer=POLY_cond $X=3.37 $Y=1.492
+ $X2=3.11 $Y2=1.492
r251 29 31 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.37 $Y=1.615
+ $X2=3.37 $Y2=2.405
r252 25 105 20.7868 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.11 $Y=1.285
+ $X2=3.11 $Y2=1.492
r253 25 27 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=3.11 $Y=1.285
+ $X2=3.11 $Y2=0.655
r254 21 69 11.9012 $w=3.24e-07 $l=8e-08 $layer=POLY_cond $X=2.94 $Y=1.492
+ $X2=3.02 $Y2=1.492
r255 21 92 38.679 $w=3.24e-07 $l=2.6e-07 $layer=POLY_cond $X=2.94 $Y=1.492
+ $X2=2.68 $Y2=1.492
r256 21 23 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.94 $Y=1.615
+ $X2=2.94 $Y2=2.405
r257 17 92 20.7868 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.68 $Y=1.285
+ $X2=2.68 $Y2=1.492
r258 17 19 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=2.68 $Y=1.285
+ $X2=2.68 $Y2=0.655
r259 13 101 20.7868 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.25 $Y=1.285
+ $X2=2.25 $Y2=1.492
r260 13 15 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=2.25 $Y=1.285
+ $X2=2.25 $Y2=0.655
r261 4 52 300 $w=1.7e-07 $l=3.2249e-07 $layer=licon1_PDIFF $count=2 $X=0.555
+ $Y=1.835 $X2=0.695 $Y2=2.095
r262 3 82 91 $w=1.7e-07 $l=3.98905e-07 $layer=licon1_NDIFF $count=2 $X=6.84
+ $Y=0.345 $X2=6.98 $Y2=0.68
r263 2 58 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=1.455
+ $Y=0.235 $X2=1.595 $Y2=0.42
r264 1 48 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=0.555
+ $Y=0.235 $X2=0.695 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__A311O_4%A3 1 3 4 5 6 8 11 15 17 18 24
r63 24 26 29.4403 $w=3.52e-07 $l=2.15e-07 $layer=POLY_cond $X=5.185 $Y=1.412
+ $X2=5.4 $Y2=1.412
r64 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.185
+ $Y=1.5 $X2=5.185 $Y2=1.5
r65 22 24 29.4403 $w=3.52e-07 $l=2.15e-07 $layer=POLY_cond $X=4.97 $Y=1.412
+ $X2=5.185 $Y2=1.412
r66 18 25 11.5244 $w=3.33e-07 $l=3.35e-07 $layer=LI1_cond $X=5.52 $Y=1.582
+ $X2=5.185 $Y2=1.582
r67 17 25 4.98819 $w=3.33e-07 $l=1.45e-07 $layer=LI1_cond $X=5.04 $Y=1.582
+ $X2=5.185 $Y2=1.582
r68 13 26 22.7654 $w=1.5e-07 $l=2.53e-07 $layer=POLY_cond $X=5.4 $Y=1.665
+ $X2=5.4 $Y2=1.412
r69 13 15 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=5.4 $Y=1.665 $X2=5.4
+ $Y2=2.465
r70 9 22 22.7654 $w=1.5e-07 $l=2.53e-07 $layer=POLY_cond $X=4.97 $Y=1.665
+ $X2=4.97 $Y2=1.412
r71 9 11 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=4.97 $Y=1.665 $X2=4.97
+ $Y2=2.465
r72 6 22 31.4943 $w=3.52e-07 $l=3.48517e-07 $layer=POLY_cond $X=4.74 $Y=1.16
+ $X2=4.97 $Y2=1.412
r73 6 8 162.273 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=4.74 $Y=1.16 $X2=4.74
+ $Y2=0.655
r74 4 6 21.7466 $w=3.52e-07 $l=1.21861e-07 $layer=POLY_cond $X=4.665 $Y=1.25
+ $X2=4.74 $Y2=1.16
r75 4 5 108.839 $w=1.8e-07 $l=2.8e-07 $layer=POLY_cond $X=4.665 $Y=1.25
+ $X2=4.385 $Y2=1.25
r76 1 5 23.1999 $w=1.93e-07 $l=1.21861e-07 $layer=POLY_cond $X=4.31 $Y=1.16
+ $X2=4.385 $Y2=1.25
r77 1 3 162.273 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=4.31 $Y=1.16 $X2=4.31
+ $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__A311O_4%A2 3 7 11 15 17 24 25
r48 23 25 9.61737 $w=3.3e-07 $l=5.5e-08 $layer=POLY_cond $X=6.28 $Y=1.51
+ $X2=6.335 $Y2=1.51
r49 23 24 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.28
+ $Y=1.51 $X2=6.28 $Y2=1.51
r50 21 23 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=6.26 $Y=1.51 $X2=6.28
+ $Y2=1.51
r51 19 21 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=5.83 $Y=1.51
+ $X2=6.26 $Y2=1.51
r52 17 24 3.08987 $w=5.98e-07 $l=1.55e-07 $layer=LI1_cond $X=6.075 $Y=1.665
+ $X2=6.075 $Y2=1.51
r53 13 25 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.335 $Y=1.345
+ $X2=6.335 $Y2=1.51
r54 13 15 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=6.335 $Y=1.345
+ $X2=6.335 $Y2=0.765
r55 9 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.26 $Y=1.675
+ $X2=6.26 $Y2=1.51
r56 9 11 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=6.26 $Y=1.675
+ $X2=6.26 $Y2=2.465
r57 5 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.83 $Y=1.675
+ $X2=5.83 $Y2=1.51
r58 5 7 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=5.83 $Y=1.675 $X2=5.83
+ $Y2=2.465
r59 1 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.83 $Y=1.345
+ $X2=5.83 $Y2=1.51
r60 1 3 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=5.83 $Y=1.345 $X2=5.83
+ $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_LP__A311O_4%A1 1 3 6 8 10 13 15 16 23
r47 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.41
+ $Y=1.46 $X2=7.41 $Y2=1.46
r48 21 23 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=7.195 $Y=1.46
+ $X2=7.41 $Y2=1.46
r49 19 21 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=6.765 $Y=1.46
+ $X2=7.195 $Y2=1.46
r50 16 24 8.43753 $w=2.78e-07 $l=2.05e-07 $layer=LI1_cond $X=7.455 $Y=1.665
+ $X2=7.455 $Y2=1.46
r51 15 24 6.79118 $w=2.78e-07 $l=1.65e-07 $layer=LI1_cond $X=7.455 $Y=1.295
+ $X2=7.455 $Y2=1.46
r52 11 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.195 $Y=1.625
+ $X2=7.195 $Y2=1.46
r53 11 13 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=7.195 $Y=1.625
+ $X2=7.195 $Y2=2.465
r54 8 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.195 $Y=1.295
+ $X2=7.195 $Y2=1.46
r55 8 10 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=7.195 $Y=1.295
+ $X2=7.195 $Y2=0.765
r56 4 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.765 $Y=1.625
+ $X2=6.765 $Y2=1.46
r57 4 6 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=6.765 $Y=1.625
+ $X2=6.765 $Y2=2.465
r58 1 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.765 $Y=1.295
+ $X2=6.765 $Y2=1.46
r59 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=6.765 $Y=1.295
+ $X2=6.765 $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_LP__A311O_4%A_28_367# 1 2 3 10 12 14 18 20 24 29
r43 22 24 21.2759 $w=2.58e-07 $l=4.8e-07 $layer=LI1_cond $X=1.99 $Y=2.905
+ $X2=1.99 $Y2=2.425
r44 21 29 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.29 $Y=2.99
+ $X2=1.125 $Y2=2.99
r45 20 22 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=1.86 $Y=2.99
+ $X2=1.99 $Y2=2.905
r46 20 21 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=1.86 $Y=2.99
+ $X2=1.29 $Y2=2.99
r47 16 29 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.125 $Y=2.905
+ $X2=1.125 $Y2=2.99
r48 16 18 31.4303 $w=3.28e-07 $l=9e-07 $layer=LI1_cond $X=1.125 $Y=2.905
+ $X2=1.125 $Y2=2.005
r49 15 27 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.43 $Y=2.99
+ $X2=0.265 $Y2=2.99
r50 14 29 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.96 $Y=2.99
+ $X2=1.125 $Y2=2.99
r51 14 15 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=0.96 $Y=2.99
+ $X2=0.43 $Y2=2.99
r52 10 27 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.265 $Y=2.905
+ $X2=0.265 $Y2=2.99
r53 10 12 31.4303 $w=3.28e-07 $l=9e-07 $layer=LI1_cond $X=0.265 $Y=2.905
+ $X2=0.265 $Y2=2.005
r54 3 24 300 $w=1.7e-07 $l=6.56277e-07 $layer=licon1_PDIFF $count=2 $X=1.885
+ $Y=1.835 $X2=2.025 $Y2=2.425
r55 2 29 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=0.985
+ $Y=1.835 $X2=1.125 $Y2=2.91
r56 2 18 400 $w=1.7e-07 $l=2.29565e-07 $layer=licon1_PDIFF $count=1 $X=0.985
+ $Y=1.835 $X2=1.125 $Y2=2.005
r57 1 27 400 $w=1.7e-07 $l=1.13578e-06 $layer=licon1_PDIFF $count=1 $X=0.14
+ $Y=1.835 $X2=0.265 $Y2=2.91
r58 1 12 400 $w=1.7e-07 $l=2.23942e-07 $layer=licon1_PDIFF $count=1 $X=0.14
+ $Y=1.835 $X2=0.265 $Y2=2.005
.ends

.subckt PM_SKY130_FD_SC_LP__A311O_4%A_283_367# 1 2 3 4 15 18 19 20 23 25 29 31
+ 35 39 42 44 49
c83 19 0 7.29344e-20 $X=5.02 $Y=2.61
r84 46 47 4.62437 $w=2.58e-07 $l=8.5e-08 $layer=LI1_cond $X=5.15 $Y=2.61
+ $X2=5.15 $Y2=2.695
r85 44 46 11.7461 $w=2.58e-07 $l=2.65e-07 $layer=LI1_cond $X=5.15 $Y=2.345
+ $X2=5.15 $Y2=2.61
r86 37 50 4.3182 $w=2.1e-07 $l=9.44722e-08 $layer=LI1_cond $X=6.98 $Y=2.26
+ $X2=6.96 $Y2=2.345
r87 37 39 16.3445 $w=1.88e-07 $l=2.8e-07 $layer=LI1_cond $X=6.98 $Y=2.26
+ $X2=6.98 $Y2=1.98
r88 33 50 4.3182 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=6.96 $Y=2.43 $X2=6.96
+ $Y2=2.345
r89 33 35 1.00212 $w=2.28e-07 $l=2e-08 $layer=LI1_cond $X=6.96 $Y=2.43 $X2=6.96
+ $Y2=2.45
r90 32 49 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=6.16 $Y=2.345
+ $X2=6.055 $Y2=2.345
r91 31 50 2.11342 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=6.845 $Y=2.345
+ $X2=6.96 $Y2=2.345
r92 31 32 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=6.845 $Y=2.345
+ $X2=6.16 $Y2=2.345
r93 27 49 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=6.055 $Y=2.43
+ $X2=6.055 $Y2=2.345
r94 27 29 25.3506 $w=2.08e-07 $l=4.8e-07 $layer=LI1_cond $X=6.055 $Y=2.43
+ $X2=6.055 $Y2=2.91
r95 26 44 3.22376 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=5.28 $Y=2.345
+ $X2=5.15 $Y2=2.345
r96 25 49 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=5.95 $Y=2.345
+ $X2=6.055 $Y2=2.345
r97 25 26 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.95 $Y=2.345
+ $X2=5.28 $Y2=2.345
r98 23 47 12.5502 $w=1.88e-07 $l=2.15e-07 $layer=LI1_cond $X=5.185 $Y=2.91
+ $X2=5.185 $Y2=2.695
r99 19 46 3.22376 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=5.02 $Y=2.61 $X2=5.15
+ $Y2=2.61
r100 19 20 167.016 $w=1.68e-07 $l=2.56e-06 $layer=LI1_cond $X=5.02 $Y=2.61
+ $X2=2.46 $Y2=2.61
r101 18 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.375 $Y=2.525
+ $X2=2.46 $Y2=2.61
r102 17 18 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=2.375 $Y=2.09
+ $X2=2.375 $Y2=2.525
r103 16 42 4.03528 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=1.69 $Y=2.005
+ $X2=1.575 $Y2=2.005
r104 15 17 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.29 $Y=2.005
+ $X2=2.375 $Y2=2.09
r105 15 16 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=2.29 $Y=2.005
+ $X2=1.69 $Y2=2.005
r106 4 39 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=6.84
+ $Y=1.835 $X2=6.98 $Y2=1.98
r107 4 35 300 $w=1.7e-07 $l=6.81414e-07 $layer=licon1_PDIFF $count=2 $X=6.84
+ $Y=1.835 $X2=6.98 $Y2=2.45
r108 3 49 600 $w=1.7e-07 $l=5.7576e-07 $layer=licon1_PDIFF $count=1 $X=5.905
+ $Y=1.835 $X2=6.045 $Y2=2.345
r109 3 29 600 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=5.905
+ $Y=1.835 $X2=6.045 $Y2=2.91
r110 2 44 600 $w=1.7e-07 $l=5.7576e-07 $layer=licon1_PDIFF $count=1 $X=5.045
+ $Y=1.835 $X2=5.185 $Y2=2.345
r111 2 23 600 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=5.045
+ $Y=1.835 $X2=5.185 $Y2=2.91
r112 1 42 300 $w=1.7e-07 $l=3.20156e-07 $layer=licon1_PDIFF $count=2 $X=1.415
+ $Y=1.835 $X2=1.575 $Y2=2.085
.ends

.subckt PM_SKY130_FD_SC_LP__A311O_4%VPWR 1 2 3 4 5 6 21 25 29 31 35 39 41 43 47
+ 48 49 51 59 68 73 79 82 85 88 92
c119 51 0 7.29344e-20 $X=2.465 $Y=3.33
r120 91 92 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r121 88 89 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r122 85 86 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r123 82 83 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r124 79 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r125 77 92 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=7.44 $Y2=3.33
r126 77 89 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=6.48 $Y2=3.33
r127 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r128 74 88 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.675 $Y=3.33
+ $X2=6.51 $Y2=3.33
r129 74 76 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=6.675 $Y=3.33
+ $X2=6.96 $Y2=3.33
r130 73 91 4.76062 $w=1.7e-07 $l=2.17e-07 $layer=LI1_cond $X=7.245 $Y=3.33
+ $X2=7.462 $Y2=3.33
r131 73 76 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=7.245 $Y=3.33
+ $X2=6.96 $Y2=3.33
r132 72 89 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=6.48
+ $Y2=3.33
r133 72 86 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=5.52
+ $Y2=3.33
r134 71 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r135 69 85 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.78 $Y=3.33
+ $X2=5.615 $Y2=3.33
r136 69 71 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=5.78 $Y=3.33 $X2=6
+ $Y2=3.33
r137 68 88 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.345 $Y=3.33
+ $X2=6.51 $Y2=3.33
r138 68 71 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=6.345 $Y=3.33 $X2=6
+ $Y2=3.33
r139 67 86 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.52 $Y2=3.33
r140 66 67 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r141 64 82 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.81 $Y=3.33
+ $X2=3.645 $Y2=3.33
r142 64 66 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=3.81 $Y=3.33
+ $X2=4.56 $Y2=3.33
r143 63 83 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r144 63 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.64 $Y2=3.33
r145 62 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r146 60 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.795 $Y=3.33
+ $X2=2.63 $Y2=3.33
r147 60 62 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=2.795 $Y=3.33
+ $X2=3.12 $Y2=3.33
r148 59 82 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.48 $Y=3.33
+ $X2=3.645 $Y2=3.33
r149 59 62 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=3.48 $Y=3.33
+ $X2=3.12 $Y2=3.33
r150 58 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r151 57 58 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r152 54 58 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=2.16 $Y2=3.33
r153 53 57 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=0.24 $Y=3.33
+ $X2=2.16 $Y2=3.33
r154 53 54 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r155 51 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.465 $Y=3.33
+ $X2=2.63 $Y2=3.33
r156 51 57 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.465 $Y=3.33
+ $X2=2.16 $Y2=3.33
r157 49 67 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=3.84 $Y=3.33
+ $X2=4.56 $Y2=3.33
r158 49 83 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.84 $Y=3.33
+ $X2=3.6 $Y2=3.33
r159 47 66 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=4.59 $Y=3.33 $X2=4.56
+ $Y2=3.33
r160 47 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.59 $Y=3.33
+ $X2=4.755 $Y2=3.33
r161 43 46 33.0018 $w=3.28e-07 $l=9.45e-07 $layer=LI1_cond $X=7.41 $Y=2.005
+ $X2=7.41 $Y2=2.95
r162 41 91 3.00555 $w=3.3e-07 $l=1.07912e-07 $layer=LI1_cond $X=7.41 $Y=3.245
+ $X2=7.462 $Y2=3.33
r163 41 46 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=7.41 $Y=3.245
+ $X2=7.41 $Y2=2.95
r164 37 88 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.51 $Y=3.245
+ $X2=6.51 $Y2=3.33
r165 37 39 18.1597 $w=3.28e-07 $l=5.2e-07 $layer=LI1_cond $X=6.51 $Y=3.245
+ $X2=6.51 $Y2=2.725
r166 33 85 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.615 $Y=3.245
+ $X2=5.615 $Y2=3.33
r167 33 35 18.1597 $w=3.28e-07 $l=5.2e-07 $layer=LI1_cond $X=5.615 $Y=3.245
+ $X2=5.615 $Y2=2.725
r168 32 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.92 $Y=3.33
+ $X2=4.755 $Y2=3.33
r169 31 85 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.45 $Y=3.33
+ $X2=5.615 $Y2=3.33
r170 31 32 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=5.45 $Y=3.33
+ $X2=4.92 $Y2=3.33
r171 27 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.755 $Y=3.245
+ $X2=4.755 $Y2=3.33
r172 27 29 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=4.755 $Y=3.245
+ $X2=4.755 $Y2=2.97
r173 23 82 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.645 $Y=3.245
+ $X2=3.645 $Y2=3.33
r174 23 25 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=3.645 $Y=3.245
+ $X2=3.645 $Y2=2.97
r175 19 79 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.63 $Y=3.245
+ $X2=2.63 $Y2=3.33
r176 19 21 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.63 $Y=3.245
+ $X2=2.63 $Y2=2.95
r177 6 46 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=7.27
+ $Y=1.835 $X2=7.41 $Y2=2.95
r178 6 43 400 $w=1.7e-07 $l=2.29565e-07 $layer=licon1_PDIFF $count=1 $X=7.27
+ $Y=1.835 $X2=7.41 $Y2=2.005
r179 5 39 600 $w=1.7e-07 $l=9.73576e-07 $layer=licon1_PDIFF $count=1 $X=6.335
+ $Y=1.835 $X2=6.51 $Y2=2.725
r180 4 35 600 $w=1.7e-07 $l=9.57445e-07 $layer=licon1_PDIFF $count=1 $X=5.475
+ $Y=1.835 $X2=5.615 $Y2=2.725
r181 3 29 600 $w=1.7e-07 $l=1.20297e-06 $layer=licon1_PDIFF $count=1 $X=4.615
+ $Y=1.835 $X2=4.755 $Y2=2.97
r182 2 25 600 $w=1.7e-07 $l=1.29113e-06 $layer=licon1_PDIFF $count=1 $X=3.445
+ $Y=1.775 $X2=3.645 $Y2=2.97
r183 1 21 600 $w=1.7e-07 $l=1.23592e-06 $layer=licon1_PDIFF $count=1 $X=2.505
+ $Y=1.775 $X2=2.63 $Y2=2.95
.ends

.subckt PM_SKY130_FD_SC_LP__A311O_4%X 1 2 3 4 15 17 18 19 25 27 30 31 32 36
r69 36 38 0.889827 $w=5.21e-07 $l=3.8e-08 $layer=LI1_cond $X=4.392 $Y=1.882
+ $X2=4.392 $Y2=1.92
r70 32 36 5.08138 $w=5.21e-07 $l=2.17e-07 $layer=LI1_cond $X=4.392 $Y=1.665
+ $X2=4.392 $Y2=1.882
r71 30 32 12.0651 $w=5.21e-07 $l=3.6307e-07 $layer=LI1_cond $X=4.145 $Y=1.405
+ $X2=4.392 $Y2=1.665
r72 29 30 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=4.145 $Y=1.195
+ $X2=4.145 $Y2=1.405
r73 28 31 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=3.42 $Y=1.11
+ $X2=3.325 $Y2=1.11
r74 27 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.06 $Y=1.11
+ $X2=4.145 $Y2=1.195
r75 27 28 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=4.06 $Y=1.11 $X2=3.42
+ $Y2=1.11
r76 23 31 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=3.325 $Y=1.025
+ $X2=3.325 $Y2=1.11
r77 23 25 35.3158 $w=1.88e-07 $l=6.05e-07 $layer=LI1_cond $X=3.325 $Y=1.025
+ $X2=3.325 $Y2=0.42
r78 19 36 4.71101 $w=2.65e-07 $l=3.32e-07 $layer=LI1_cond $X=4.06 $Y=1.882
+ $X2=4.392 $Y2=1.882
r79 19 21 39.357 $w=2.63e-07 $l=9.05e-07 $layer=LI1_cond $X=4.06 $Y=1.882
+ $X2=3.155 $Y2=1.882
r80 17 31 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=3.23 $Y=1.11
+ $X2=3.325 $Y2=1.11
r81 17 18 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.23 $Y=1.11
+ $X2=2.56 $Y2=1.11
r82 13 18 6.83233 $w=1.7e-07 $l=1.28662e-07 $layer=LI1_cond $X=2.467 $Y=1.025
+ $X2=2.56 $Y2=1.11
r83 13 15 36.2703 $w=1.83e-07 $l=6.05e-07 $layer=LI1_cond $X=2.467 $Y=1.025
+ $X2=2.467 $Y2=0.42
r84 4 38 600 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_PDIFF $count=1 $X=3.995
+ $Y=1.775 $X2=4.23 $Y2=1.92
r85 3 21 600 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=3.015
+ $Y=1.775 $X2=3.155 $Y2=1.9
r86 2 25 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=3.185
+ $Y=0.235 $X2=3.325 $Y2=0.42
r87 1 15 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=2.325
+ $Y=0.235 $X2=2.465 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__A311O_4%VGND 1 2 3 4 5 6 19 21 25 29 33 35 39 43 46
+ 47 48 49 50 52 64 71 72 78 81 86
r107 86 87 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r108 81 84 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r109 81 82 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r110 78 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r111 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r112 72 87 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=7.44 $Y=0 $X2=5.04
+ $Y2=0
r113 71 72 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r114 69 86 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.12 $Y=0 $X2=4.955
+ $Y2=0
r115 69 71 151.358 $w=1.68e-07 $l=2.32e-06 $layer=LI1_cond $X=5.12 $Y=0 $X2=7.44
+ $Y2=0
r116 68 87 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.04
+ $Y2=0
r117 68 82 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=4.08
+ $Y2=0
r118 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r119 65 81 13.3456 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=4.26 $Y=0 $X2=3.925
+ $Y2=0
r120 65 67 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=4.26 $Y=0 $X2=4.56
+ $Y2=0
r121 64 86 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.79 $Y=0 $X2=4.955
+ $Y2=0
r122 64 67 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=4.79 $Y=0 $X2=4.56
+ $Y2=0
r123 63 84 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r124 62 63 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r125 60 63 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r126 60 79 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r127 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r128 57 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.305 $Y=0 $X2=1.14
+ $Y2=0
r129 57 59 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.305 $Y=0
+ $X2=1.68 $Y2=0
r130 56 79 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r131 56 76 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r132 55 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r133 53 75 4.77065 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=0.43 $Y=0 $X2=0.215
+ $Y2=0
r134 53 55 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=0.43 $Y=0 $X2=0.72
+ $Y2=0
r135 52 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.975 $Y=0 $X2=1.14
+ $Y2=0
r136 52 55 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.975 $Y=0
+ $X2=0.72 $Y2=0
r137 50 82 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.84 $Y=0
+ $X2=4.08 $Y2=0
r138 50 84 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.84 $Y=0 $X2=3.6
+ $Y2=0
r139 48 62 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=2.73 $Y=0 $X2=2.64
+ $Y2=0
r140 48 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.73 $Y=0 $X2=2.895
+ $Y2=0
r141 46 59 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=1.86 $Y=0 $X2=1.68
+ $Y2=0
r142 46 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.86 $Y=0 $X2=2.025
+ $Y2=0
r143 45 62 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=2.19 $Y=0 $X2=2.64
+ $Y2=0
r144 45 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.19 $Y=0 $X2=2.025
+ $Y2=0
r145 41 86 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.955 $Y=0.085
+ $X2=4.955 $Y2=0
r146 41 43 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=4.955 $Y=0.085
+ $X2=4.955 $Y2=0.38
r147 37 81 2.76849 $w=6.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.925 $Y=0.085
+ $X2=3.925 $Y2=0
r148 37 39 5.26632 $w=6.68e-07 $l=2.95e-07 $layer=LI1_cond $X=3.925 $Y=0.085
+ $X2=3.925 $Y2=0.38
r149 36 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.06 $Y=0 $X2=2.895
+ $Y2=0
r150 35 81 13.3456 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=3.59 $Y=0 $X2=3.925
+ $Y2=0
r151 35 36 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=3.59 $Y=0 $X2=3.06
+ $Y2=0
r152 31 49 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.895 $Y=0.085
+ $X2=2.895 $Y2=0
r153 31 33 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.895 $Y=0.085
+ $X2=2.895 $Y2=0.38
r154 27 47 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.025 $Y=0.085
+ $X2=2.025 $Y2=0
r155 27 29 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.025 $Y=0.085
+ $X2=2.025 $Y2=0.38
r156 23 78 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.14 $Y=0.085
+ $X2=1.14 $Y2=0
r157 23 25 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=1.14 $Y=0.085
+ $X2=1.14 $Y2=0.36
r158 19 75 2.99552 $w=3.3e-07 $l=1.07121e-07 $layer=LI1_cond $X=0.265 $Y=0.085
+ $X2=0.215 $Y2=0
r159 19 21 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.265 $Y=0.085
+ $X2=0.265 $Y2=0.38
r160 6 43 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.815
+ $Y=0.235 $X2=4.955 $Y2=0.38
r161 5 39 45.5 $w=1.7e-07 $l=5.47723e-07 $layer=licon1_NDIFF $count=4 $X=3.615
+ $Y=0.235 $X2=4.095 $Y2=0.38
r162 4 33 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.755
+ $Y=0.235 $X2=2.895 $Y2=0.38
r163 3 29 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.885
+ $Y=0.235 $X2=2.025 $Y2=0.38
r164 2 25 91 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=2 $X=0.985
+ $Y=0.235 $X2=1.14 $Y2=0.36
r165 1 21 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.14
+ $Y=0.235 $X2=0.265 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_LP__A311O_4%A_877_47# 1 2 9 12 13 17 19 20
c32 12 0 1.45841e-19 $X=4.62 $Y=1.15
r33 19 20 8.51806 $w=2.28e-07 $l=1.7e-07 $layer=LI1_cond $X=5.21 $Y=1.12
+ $X2=5.38 $Y2=1.12
r34 15 17 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=6.08 $Y=1.005
+ $X2=6.08 $Y2=0.68
r35 13 15 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.915 $Y=1.09
+ $X2=6.08 $Y2=1.005
r36 13 20 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=5.915 $Y=1.09
+ $X2=5.38 $Y2=1.09
r37 12 19 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=4.62 $Y=1.15 $X2=5.21
+ $Y2=1.15
r38 7 12 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=4.525 $Y=1.065
+ $X2=4.62 $Y2=1.15
r39 7 9 37.6507 $w=1.88e-07 $l=6.45e-07 $layer=LI1_cond $X=4.525 $Y=1.065
+ $X2=4.525 $Y2=0.42
r40 2 17 91 $w=1.7e-07 $l=4.1334e-07 $layer=licon1_NDIFF $count=2 $X=5.905
+ $Y=0.345 $X2=6.08 $Y2=0.68
r41 1 9 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=4.385
+ $Y=0.235 $X2=4.525 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__A311O_4%A_1098_69# 1 2 3 12 14 15 18 20 24 26
r30 22 24 2.88111 $w=2.58e-07 $l=6.5e-08 $layer=LI1_cond $X=7.445 $Y=0.425
+ $X2=7.445 $Y2=0.49
r31 21 26 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=6.645 $Y=0.34
+ $X2=6.53 $Y2=0.34
r32 20 22 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=7.315 $Y=0.34
+ $X2=7.445 $Y2=0.425
r33 20 21 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=7.315 $Y=0.34
+ $X2=6.645 $Y2=0.34
r34 16 26 0.280307 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.53 $Y=0.425
+ $X2=6.53 $Y2=0.34
r35 16 18 3.2569 $w=2.28e-07 $l=6.5e-08 $layer=LI1_cond $X=6.53 $Y=0.425
+ $X2=6.53 $Y2=0.49
r36 14 26 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=6.415 $Y=0.34
+ $X2=6.53 $Y2=0.34
r37 14 15 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=6.415 $Y=0.34
+ $X2=5.745 $Y2=0.34
r38 10 15 7.47753 $w=1.7e-07 $l=1.85699e-07 $layer=LI1_cond $X=5.597 $Y=0.425
+ $X2=5.745 $Y2=0.34
r39 10 12 9.57114 $w=2.93e-07 $l=2.45e-07 $layer=LI1_cond $X=5.597 $Y=0.425
+ $X2=5.597 $Y2=0.67
r40 3 24 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=7.27
+ $Y=0.345 $X2=7.41 $Y2=0.49
r41 2 18 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.41
+ $Y=0.345 $X2=6.55 $Y2=0.49
r42 1 12 182 $w=1.7e-07 $l=3.82426e-07 $layer=licon1_NDIFF $count=1 $X=5.49
+ $Y=0.345 $X2=5.615 $Y2=0.67
.ends

