* File: sky130_fd_sc_lp__sdfrtn_1.pxi.spice
* Created: Wed Sep  2 10:34:28 2020
* 
x_PM_SKY130_FD_SC_LP__SDFRTN_1%A_113_63# N_A_113_63#_M1039_d N_A_113_63#_M1021_d
+ N_A_113_63#_c_267_n N_A_113_63#_M1032_g N_A_113_63#_M1015_g
+ N_A_113_63#_c_262_n N_A_113_63#_c_269_n N_A_113_63#_c_270_n
+ N_A_113_63#_c_263_n N_A_113_63#_c_264_n N_A_113_63#_c_272_n
+ N_A_113_63#_c_273_n N_A_113_63#_c_265_n N_A_113_63#_c_266_n
+ PM_SKY130_FD_SC_LP__SDFRTN_1%A_113_63#
x_PM_SKY130_FD_SC_LP__SDFRTN_1%SCD N_SCD_c_341_n N_SCD_c_342_n N_SCD_M1026_g
+ N_SCD_M1037_g N_SCD_c_343_n N_SCD_c_344_n N_SCD_c_345_n SCD SCD N_SCD_c_346_n
+ N_SCD_c_347_n PM_SKY130_FD_SC_LP__SDFRTN_1%SCD
x_PM_SKY130_FD_SC_LP__SDFRTN_1%SCE N_SCE_M1039_g N_SCE_M1021_g N_SCE_c_395_n
+ N_SCE_M1028_g N_SCE_M1014_g N_SCE_c_397_n N_SCE_c_398_n N_SCE_c_399_n SCE SCE
+ N_SCE_c_404_n PM_SKY130_FD_SC_LP__SDFRTN_1%SCE
x_PM_SKY130_FD_SC_LP__SDFRTN_1%D N_D_M1010_g N_D_c_466_n N_D_M1018_g D
+ PM_SKY130_FD_SC_LP__SDFRTN_1%D
x_PM_SKY130_FD_SC_LP__SDFRTN_1%RESET_B N_RESET_B_M1000_g N_RESET_B_M1034_g
+ N_RESET_B_c_525_n N_RESET_B_M1003_g N_RESET_B_M1009_g N_RESET_B_c_526_n
+ N_RESET_B_c_514_n N_RESET_B_M1033_g N_RESET_B_M1002_g N_RESET_B_c_516_n
+ N_RESET_B_c_530_n N_RESET_B_c_531_n N_RESET_B_c_532_n N_RESET_B_c_517_n
+ N_RESET_B_c_534_n N_RESET_B_c_602_p N_RESET_B_c_535_n N_RESET_B_c_571_p
+ N_RESET_B_c_518_n N_RESET_B_c_537_n N_RESET_B_c_519_n N_RESET_B_c_520_n
+ N_RESET_B_c_572_p RESET_B RESET_B N_RESET_B_c_540_n N_RESET_B_c_541_n
+ N_RESET_B_c_542_n N_RESET_B_c_543_n N_RESET_B_c_544_n N_RESET_B_c_521_n
+ N_RESET_B_c_522_n N_RESET_B_c_523_n RESET_B
+ PM_SKY130_FD_SC_LP__SDFRTN_1%RESET_B
x_PM_SKY130_FD_SC_LP__SDFRTN_1%CLK_N N_CLK_N_M1035_g N_CLK_N_M1023_g CLK_N
+ N_CLK_N_c_752_n N_CLK_N_c_753_n PM_SKY130_FD_SC_LP__SDFRTN_1%CLK_N
x_PM_SKY130_FD_SC_LP__SDFRTN_1%A_1080_47# N_A_1080_47#_M1019_d
+ N_A_1080_47#_M1022_d N_A_1080_47#_M1020_g N_A_1080_47#_M1027_g
+ N_A_1080_47#_M1006_g N_A_1080_47#_M1017_g N_A_1080_47#_c_792_n
+ N_A_1080_47#_c_793_n N_A_1080_47#_c_810_n N_A_1080_47#_c_794_n
+ N_A_1080_47#_c_795_n N_A_1080_47#_c_796_n N_A_1080_47#_c_797_n
+ N_A_1080_47#_c_820_n N_A_1080_47#_c_831_p N_A_1080_47#_c_798_n
+ N_A_1080_47#_c_799_n N_A_1080_47#_c_800_n N_A_1080_47#_c_801_n
+ N_A_1080_47#_c_802_n N_A_1080_47#_c_803_n N_A_1080_47#_c_812_n
+ N_A_1080_47#_c_804_n N_A_1080_47#_c_889_p N_A_1080_47#_c_813_n
+ N_A_1080_47#_c_814_n N_A_1080_47#_c_815_n N_A_1080_47#_c_805_n
+ N_A_1080_47#_c_806_n PM_SKY130_FD_SC_LP__SDFRTN_1%A_1080_47#
x_PM_SKY130_FD_SC_LP__SDFRTN_1%A_1406_399# N_A_1406_399#_M1001_d
+ N_A_1406_399#_M1038_d N_A_1406_399#_M1036_g N_A_1406_399#_M1007_g
+ N_A_1406_399#_c_968_n N_A_1406_399#_c_975_n N_A_1406_399#_c_969_n
+ N_A_1406_399#_c_970_n N_A_1406_399#_c_1014_n N_A_1406_399#_c_971_n
+ N_A_1406_399#_c_1000_n N_A_1406_399#_c_1003_n
+ PM_SKY130_FD_SC_LP__SDFRTN_1%A_1406_399#
x_PM_SKY130_FD_SC_LP__SDFRTN_1%A_1278_529# N_A_1278_529#_M1020_d
+ N_A_1278_529#_M1005_d N_A_1278_529#_M1003_d N_A_1278_529#_M1001_g
+ N_A_1278_529#_c_1058_n N_A_1278_529#_c_1059_n N_A_1278_529#_c_1060_n
+ N_A_1278_529#_M1038_g N_A_1278_529#_c_1061_n N_A_1278_529#_c_1056_n
+ N_A_1278_529#_c_1063_n N_A_1278_529#_c_1064_n N_A_1278_529#_c_1065_n
+ N_A_1278_529#_c_1066_n N_A_1278_529#_c_1067_n
+ PM_SKY130_FD_SC_LP__SDFRTN_1%A_1278_529#
x_PM_SKY130_FD_SC_LP__SDFRTN_1%A_857_367# N_A_857_367#_M1023_d
+ N_A_857_367#_M1035_d N_A_857_367#_M1019_g N_A_857_367#_M1022_g
+ N_A_857_367#_c_1171_n N_A_857_367#_c_1172_n N_A_857_367#_c_1173_n
+ N_A_857_367#_c_1187_n N_A_857_367#_M1005_g N_A_857_367#_M1008_g
+ N_A_857_367#_c_1175_n N_A_857_367#_c_1176_n N_A_857_367#_M1016_g
+ N_A_857_367#_c_1178_n N_A_857_367#_c_1179_n N_A_857_367#_M1024_g
+ N_A_857_367#_c_1181_n N_A_857_367#_c_1189_n N_A_857_367#_c_1190_n
+ N_A_857_367#_c_1182_n N_A_857_367#_c_1183_n N_A_857_367#_c_1184_n
+ PM_SKY130_FD_SC_LP__SDFRTN_1%A_857_367#
x_PM_SKY130_FD_SC_LP__SDFRTN_1%A_2064_101# N_A_2064_101#_M1030_d
+ N_A_2064_101#_M1033_d N_A_2064_101#_M1029_g N_A_2064_101#_M1012_g
+ N_A_2064_101#_c_1326_n N_A_2064_101#_c_1327_n N_A_2064_101#_c_1328_n
+ N_A_2064_101#_c_1329_n N_A_2064_101#_c_1330_n N_A_2064_101#_c_1331_n
+ N_A_2064_101#_c_1322_n N_A_2064_101#_c_1323_n N_A_2064_101#_c_1333_n
+ PM_SKY130_FD_SC_LP__SDFRTN_1%A_2064_101#
x_PM_SKY130_FD_SC_LP__SDFRTN_1%A_1870_127# N_A_1870_127#_M1016_d
+ N_A_1870_127#_M1006_d N_A_1870_127#_M1030_g N_A_1870_127#_M1013_g
+ N_A_1870_127#_c_1413_n N_A_1870_127#_c_1414_n N_A_1870_127#_M1004_g
+ N_A_1870_127#_c_1416_n N_A_1870_127#_M1011_g N_A_1870_127#_c_1417_n
+ N_A_1870_127#_c_1418_n N_A_1870_127#_c_1419_n N_A_1870_127#_c_1420_n
+ N_A_1870_127#_c_1421_n N_A_1870_127#_c_1422_n N_A_1870_127#_c_1423_n
+ N_A_1870_127#_c_1429_n N_A_1870_127#_c_1424_n N_A_1870_127#_c_1425_n
+ PM_SKY130_FD_SC_LP__SDFRTN_1%A_1870_127#
x_PM_SKY130_FD_SC_LP__SDFRTN_1%A_2370_351# N_A_2370_351#_M1011_s
+ N_A_2370_351#_M1004_s N_A_2370_351#_M1025_g N_A_2370_351#_M1031_g
+ N_A_2370_351#_c_1544_n N_A_2370_351#_c_1538_n N_A_2370_351#_c_1545_n
+ N_A_2370_351#_c_1539_n N_A_2370_351#_c_1540_n N_A_2370_351#_c_1541_n
+ N_A_2370_351#_c_1542_n PM_SKY130_FD_SC_LP__SDFRTN_1%A_2370_351#
x_PM_SKY130_FD_SC_LP__SDFRTN_1%VPWR N_VPWR_M1021_s N_VPWR_M1037_d N_VPWR_M1000_d
+ N_VPWR_M1022_s N_VPWR_M1036_d N_VPWR_M1038_s N_VPWR_M1012_d N_VPWR_M1013_d
+ N_VPWR_M1004_d N_VPWR_c_1598_n N_VPWR_c_1599_n N_VPWR_c_1600_n N_VPWR_c_1601_n
+ N_VPWR_c_1602_n N_VPWR_c_1603_n N_VPWR_c_1604_n N_VPWR_c_1605_n
+ N_VPWR_c_1606_n N_VPWR_c_1607_n N_VPWR_c_1608_n N_VPWR_c_1609_n
+ N_VPWR_c_1610_n N_VPWR_c_1611_n N_VPWR_c_1612_n N_VPWR_c_1613_n
+ N_VPWR_c_1614_n N_VPWR_c_1615_n VPWR N_VPWR_c_1616_n N_VPWR_c_1617_n
+ N_VPWR_c_1618_n N_VPWR_c_1619_n N_VPWR_c_1597_n N_VPWR_c_1621_n
+ N_VPWR_c_1622_n N_VPWR_c_1623_n N_VPWR_c_1624_n N_VPWR_c_1625_n
+ PM_SKY130_FD_SC_LP__SDFRTN_1%VPWR
x_PM_SKY130_FD_SC_LP__SDFRTN_1%A_229_491# N_A_229_491#_M1028_d
+ N_A_229_491#_M1020_s N_A_229_491#_M1032_s N_A_229_491#_M1018_d
+ N_A_229_491#_M1005_s N_A_229_491#_c_1781_n N_A_229_491#_c_1770_n
+ N_A_229_491#_c_1775_n N_A_229_491#_c_1771_n N_A_229_491#_c_1772_n
+ N_A_229_491#_c_1777_n N_A_229_491#_c_1778_n N_A_229_491#_c_1779_n
+ N_A_229_491#_c_1773_n N_A_229_491#_c_1780_n N_A_229_491#_c_1826_n
+ N_A_229_491#_c_1834_n N_A_229_491#_c_1774_n
+ PM_SKY130_FD_SC_LP__SDFRTN_1%A_229_491#
x_PM_SKY130_FD_SC_LP__SDFRTN_1%Q N_Q_M1031_d N_Q_M1025_d Q Q Q Q Q Q Q
+ N_Q_c_1923_n N_Q_c_1926_n Q PM_SKY130_FD_SC_LP__SDFRTN_1%Q
x_PM_SKY130_FD_SC_LP__SDFRTN_1%VGND N_VGND_M1039_s N_VGND_M1034_d N_VGND_M1019_s
+ N_VGND_M1009_d N_VGND_M1029_d N_VGND_M1011_d N_VGND_c_1942_n N_VGND_c_1943_n
+ N_VGND_c_1944_n N_VGND_c_1945_n N_VGND_c_1946_n N_VGND_c_1947_n
+ N_VGND_c_1948_n VGND N_VGND_c_1949_n N_VGND_c_1950_n N_VGND_c_1951_n
+ N_VGND_c_1952_n N_VGND_c_1953_n N_VGND_c_1954_n N_VGND_c_1955_n
+ N_VGND_c_1956_n N_VGND_c_1957_n N_VGND_c_1958_n N_VGND_c_1959_n
+ N_VGND_c_1960_n PM_SKY130_FD_SC_LP__SDFRTN_1%VGND
x_PM_SKY130_FD_SC_LP__SDFRTN_1%noxref_24 N_noxref_24_M1026_s N_noxref_24_M1015_d
+ N_noxref_24_c_2073_n N_noxref_24_c_2074_n N_noxref_24_c_2075_n
+ PM_SKY130_FD_SC_LP__SDFRTN_1%noxref_24
cc_1 VNB N_A_113_63#_M1015_g 0.0234979f $X=-0.19 $Y=-0.245 $X2=3.17 $Y2=0.505
cc_2 VNB N_A_113_63#_c_262_n 0.0269043f $X=-0.19 $Y=-0.245 $X2=0.672 $Y2=1.815
cc_3 VNB N_A_113_63#_c_263_n 0.00531001f $X=-0.19 $Y=-0.245 $X2=3.18 $Y2=2.02
cc_4 VNB N_A_113_63#_c_264_n 0.00784981f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=0.46
cc_5 VNB N_A_113_63#_c_265_n 0.0027201f $X=-0.19 $Y=-0.245 $X2=3.26 $Y2=1.12
cc_6 VNB N_A_113_63#_c_266_n 0.0351422f $X=-0.19 $Y=-0.245 $X2=3.26 $Y2=1.12
cc_7 VNB N_SCD_c_341_n 0.026977f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=0.315
cc_8 VNB N_SCD_c_342_n 0.0181208f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_SCD_c_343_n 0.00434237f $X=-0.19 $Y=-0.245 $X2=3.17 $Y2=0.955
cc_10 VNB N_SCD_c_344_n 0.0166036f $X=-0.19 $Y=-0.245 $X2=3.17 $Y2=0.505
cc_11 VNB N_SCD_c_345_n 0.00765776f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_SCD_c_346_n 0.0357695f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=0.43
cc_13 VNB N_SCD_c_347_n 0.0131659f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=2.33
cc_14 VNB N_SCE_M1039_g 0.0577911f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_SCE_M1021_g 0.0226377f $X=-0.19 $Y=-0.245 $X2=1.485 $Y2=2.345
cc_16 VNB N_SCE_c_395_n 0.0937901f $X=-0.19 $Y=-0.245 $X2=1.485 $Y2=2.775
cc_17 VNB N_SCE_M1028_g 0.0317425f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_SCE_c_397_n 0.0106787f $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=2.36
cc_19 VNB N_SCE_c_398_n 0.00638f $X=-0.19 $Y=-0.245 $X2=0.672 $Y2=0.43
cc_20 VNB N_SCE_c_399_n 0.0357747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB SCE 0.0102327f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_D_M1010_g 0.0317541f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_D_c_466_n 0.060329f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB D 0.00676984f $X=-0.19 $Y=-0.245 $X2=1.485 $Y2=2.775
cc_25 VNB N_RESET_B_M1034_g 0.0610647f $X=-0.19 $Y=-0.245 $X2=1.485 $Y2=2.345
cc_26 VNB N_RESET_B_M1009_g 0.030542f $X=-0.19 $Y=-0.245 $X2=0.672 $Y2=0.565
cc_27 VNB N_RESET_B_c_514_n 0.0111589f $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=2.36
cc_28 VNB N_RESET_B_M1002_g 0.0244015f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_RESET_B_c_516_n 0.0189328f $X=-0.19 $Y=-0.245 $X2=1.26 $Y2=2.205
cc_30 VNB N_RESET_B_c_517_n 0.00590095f $X=-0.19 $Y=-0.245 $X2=3.26 $Y2=1.12
cc_31 VNB N_RESET_B_c_518_n 0.00334871f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_RESET_B_c_519_n 0.0015053f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_RESET_B_c_520_n 0.0233424f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_RESET_B_c_521_n 0.00301754f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_RESET_B_c_522_n 0.0226175f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_RESET_B_c_523_n 0.00225256f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_CLK_N_M1023_g 0.0254414f $X=-0.19 $Y=-0.245 $X2=1.485 $Y2=2.345
cc_38 VNB N_CLK_N_c_752_n 0.0447173f $X=-0.19 $Y=-0.245 $X2=0.672 $Y2=1.815
cc_39 VNB N_CLK_N_c_753_n 0.00159439f $X=-0.19 $Y=-0.245 $X2=1.185 $Y2=2.205
cc_40 VNB N_A_1080_47#_c_792_n 0.00581801f $X=-0.19 $Y=-0.245 $X2=0.672 $Y2=0.43
cc_41 VNB N_A_1080_47#_c_793_n 0.0215439f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_1080_47#_c_794_n 0.0103855f $X=-0.19 $Y=-0.245 $X2=1.26 $Y2=2.205
cc_43 VNB N_A_1080_47#_c_795_n 0.00453692f $X=-0.19 $Y=-0.245 $X2=1.26 $Y2=2.13
cc_44 VNB N_A_1080_47#_c_796_n 0.0155175f $X=-0.19 $Y=-0.245 $X2=1.26 $Y2=2.13
cc_45 VNB N_A_1080_47#_c_797_n 0.00111447f $X=-0.19 $Y=-0.245 $X2=3.18 $Y2=1.12
cc_46 VNB N_A_1080_47#_c_798_n 0.00574474f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_1080_47#_c_799_n 0.00323794f $X=-0.19 $Y=-0.245 $X2=1.485
+ $Y2=2.345
cc_48 VNB N_A_1080_47#_c_800_n 0.00887346f $X=-0.19 $Y=-0.245 $X2=3.26 $Y2=1.12
cc_49 VNB N_A_1080_47#_c_801_n 0.0130844f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_1080_47#_c_802_n 0.0430832f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_1080_47#_c_803_n 0.0037057f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_1080_47#_c_804_n 0.0429625f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_1080_47#_c_805_n 0.0176468f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_1080_47#_c_806_n 0.0143693f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_1406_399#_M1007_g 0.0348348f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_1406_399#_c_968_n 0.00277969f $X=-0.19 $Y=-0.245 $X2=0.81
+ $Y2=2.205
cc_57 VNB N_A_1406_399#_c_969_n 0.0132051f $X=-0.19 $Y=-0.245 $X2=3.18 $Y2=1.205
cc_58 VNB N_A_1406_399#_c_970_n 0.00295782f $X=-0.19 $Y=-0.245 $X2=3.18 $Y2=2.02
cc_59 VNB N_A_1406_399#_c_971_n 0.00787368f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_1278_529#_M1001_g 0.0360849f $X=-0.19 $Y=-0.245 $X2=3.17 $Y2=0.505
cc_61 VNB N_A_1278_529#_c_1056_n 0.013303f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=1.98
cc_62 VNB N_A_857_367#_M1019_g 0.0294622f $X=-0.19 $Y=-0.245 $X2=1.485 $Y2=2.775
cc_63 VNB N_A_857_367#_M1022_g 0.00185418f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_A_857_367#_c_1171_n 0.0341218f $X=-0.19 $Y=-0.245 $X2=0.672
+ $Y2=1.815
cc_65 VNB N_A_857_367#_c_1172_n 0.00337036f $X=-0.19 $Y=-0.245 $X2=2.79 $Y2=2.36
cc_66 VNB N_A_857_367#_c_1173_n 0.0607317f $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=2.36
cc_67 VNB N_A_857_367#_M1008_g 0.0391829f $X=-0.19 $Y=-0.245 $X2=0.692 $Y2=2.155
cc_68 VNB N_A_857_367#_c_1175_n 0.15677f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=2.33
cc_69 VNB N_A_857_367#_c_1176_n 0.0113562f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=1.98
cc_70 VNB N_A_857_367#_M1016_g 0.0314682f $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=2.205
cc_71 VNB N_A_857_367#_c_1178_n 0.0510418f $X=-0.19 $Y=-0.245 $X2=3.18 $Y2=2.195
cc_72 VNB N_A_857_367#_c_1179_n 0.0128727f $X=-0.19 $Y=-0.245 $X2=3.18 $Y2=1.12
cc_73 VNB N_A_857_367#_M1024_g 0.00661793f $X=-0.19 $Y=-0.245 $X2=3.26 $Y2=1.12
cc_74 VNB N_A_857_367#_c_1181_n 0.00620718f $X=-0.19 $Y=-0.245 $X2=1.26
+ $Y2=2.155
cc_75 VNB N_A_857_367#_c_1182_n 0.014649f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_A_857_367#_c_1183_n 0.00305036f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_A_857_367#_c_1184_n 0.0426154f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_A_2064_101#_M1029_g 0.0412839f $X=-0.19 $Y=-0.245 $X2=1.485
+ $Y2=2.775
cc_79 VNB N_A_2064_101#_c_1322_n 0.00907321f $X=-0.19 $Y=-0.245 $X2=0.705
+ $Y2=2.33
cc_80 VNB N_A_2064_101#_c_1323_n 0.00720614f $X=-0.19 $Y=-0.245 $X2=1.425
+ $Y2=2.205
cc_81 VNB N_A_1870_127#_M1013_g 0.00965759f $X=-0.19 $Y=-0.245 $X2=3.17
+ $Y2=0.505
cc_82 VNB N_A_1870_127#_c_1413_n 0.0346559f $X=-0.19 $Y=-0.245 $X2=0.672
+ $Y2=0.565
cc_83 VNB N_A_1870_127#_c_1414_n 0.0102926f $X=-0.19 $Y=-0.245 $X2=0.81
+ $Y2=2.205
cc_84 VNB N_A_1870_127#_M1004_g 0.0138065f $X=-0.19 $Y=-0.245 $X2=3.18 $Y2=1.205
cc_85 VNB N_A_1870_127#_c_1416_n 0.0215031f $X=-0.19 $Y=-0.245 $X2=0.672
+ $Y2=0.43
cc_86 VNB N_A_1870_127#_c_1417_n 0.027366f $X=-0.19 $Y=-0.245 $X2=0.692
+ $Y2=2.155
cc_87 VNB N_A_1870_127#_c_1418_n 0.00550205f $X=-0.19 $Y=-0.245 $X2=0.705
+ $Y2=1.98
cc_88 VNB N_A_1870_127#_c_1419_n 0.00235891f $X=-0.19 $Y=-0.245 $X2=1.26
+ $Y2=2.13
cc_89 VNB N_A_1870_127#_c_1420_n 0.00323554f $X=-0.19 $Y=-0.245 $X2=3.18
+ $Y2=1.12
cc_90 VNB N_A_1870_127#_c_1421_n 0.0145941f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_A_1870_127#_c_1422_n 0.00125491f $X=-0.19 $Y=-0.245 $X2=1.26
+ $Y2=2.155
cc_92 VNB N_A_1870_127#_c_1423_n 0.00308386f $X=-0.19 $Y=-0.245 $X2=3.26
+ $Y2=0.955
cc_93 VNB N_A_1870_127#_c_1424_n 0.0283434f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_94 VNB N_A_1870_127#_c_1425_n 0.0180207f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_95 VNB N_A_2370_351#_M1025_g 0.00184036f $X=-0.19 $Y=-0.245 $X2=1.485
+ $Y2=2.775
cc_96 VNB N_A_2370_351#_c_1538_n 0.00696788f $X=-0.19 $Y=-0.245 $X2=3.18
+ $Y2=1.205
cc_97 VNB N_A_2370_351#_c_1539_n 0.00394723f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_98 VNB N_A_2370_351#_c_1540_n 0.0358601f $X=-0.19 $Y=-0.245 $X2=0.692
+ $Y2=2.155
cc_99 VNB N_A_2370_351#_c_1541_n 0.00188487f $X=-0.19 $Y=-0.245 $X2=0.705
+ $Y2=1.98
cc_100 VNB N_A_2370_351#_c_1542_n 0.0212406f $X=-0.19 $Y=-0.245 $X2=1.26
+ $Y2=2.13
cc_101 VNB N_VPWR_c_1597_n 0.561729f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_102 VNB N_A_229_491#_c_1770_n 0.0102152f $X=-0.19 $Y=-0.245 $X2=2.79 $Y2=2.36
cc_103 VNB N_A_229_491#_c_1771_n 0.014472f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_104 VNB N_A_229_491#_c_1772_n 0.0146245f $X=-0.19 $Y=-0.245 $X2=0.705
+ $Y2=0.43
cc_105 VNB N_A_229_491#_c_1773_n 0.00871578f $X=-0.19 $Y=-0.245 $X2=1.26
+ $Y2=2.155
cc_106 VNB N_A_229_491#_c_1774_n 0.00674342f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_107 VNB N_Q_c_1923_n 0.0609276f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=0.43
cc_108 VNB N_VGND_c_1942_n 0.0113841f $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=2.36
cc_109 VNB N_VGND_c_1943_n 0.025654f $X=-0.19 $Y=-0.245 $X2=3.18 $Y2=2.02
cc_110 VNB N_VGND_c_1944_n 0.00741811f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=0.46
cc_111 VNB N_VGND_c_1945_n 0.00632233f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=1.98
cc_112 VNB N_VGND_c_1946_n 0.0205679f $X=-0.19 $Y=-0.245 $X2=1.425 $Y2=2.205
cc_113 VNB N_VGND_c_1947_n 0.0258229f $X=-0.19 $Y=-0.245 $X2=3.26 $Y2=1.12
cc_114 VNB N_VGND_c_1948_n 0.00983248f $X=-0.19 $Y=-0.245 $X2=1.485 $Y2=2.345
cc_115 VNB N_VGND_c_1949_n 0.0847976f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_116 VNB N_VGND_c_1950_n 0.0201399f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_117 VNB N_VGND_c_1951_n 0.0721874f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_118 VNB N_VGND_c_1952_n 0.0542927f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_119 VNB N_VGND_c_1953_n 0.0477805f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_120 VNB N_VGND_c_1954_n 0.0160851f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_121 VNB N_VGND_c_1955_n 0.707492f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_122 VNB N_VGND_c_1956_n 0.00631381f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_123 VNB N_VGND_c_1957_n 0.00510065f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_124 VNB N_VGND_c_1958_n 0.00436638f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_125 VNB N_VGND_c_1959_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_126 VNB N_VGND_c_1960_n 0.00689498f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_127 VNB N_noxref_24_c_2073_n 0.00771805f $X=-0.19 $Y=-0.245 $X2=1.485
+ $Y2=2.775
cc_128 VNB N_noxref_24_c_2074_n 0.00257438f $X=-0.19 $Y=-0.245 $X2=0.672
+ $Y2=1.815
cc_129 VNB N_noxref_24_c_2075_n 0.00733364f $X=-0.19 $Y=-0.245 $X2=1.185
+ $Y2=2.205
cc_130 VPB N_A_113_63#_c_267_n 0.0189966f $X=-0.19 $Y=1.655 $X2=1.485 $Y2=2.345
cc_131 VPB N_A_113_63#_c_262_n 0.0150256f $X=-0.19 $Y=1.655 $X2=0.672 $Y2=1.815
cc_132 VPB N_A_113_63#_c_269_n 0.0171416f $X=-0.19 $Y=1.655 $X2=1.185 $Y2=2.205
cc_133 VPB N_A_113_63#_c_270_n 0.0314176f $X=-0.19 $Y=1.655 $X2=2.79 $Y2=2.36
cc_134 VPB N_A_113_63#_c_263_n 0.00211869f $X=-0.19 $Y=1.655 $X2=3.18 $Y2=2.02
cc_135 VPB N_A_113_63#_c_272_n 0.0552249f $X=-0.19 $Y=1.655 $X2=1.26 $Y2=2.13
cc_136 VPB N_A_113_63#_c_273_n 0.00482191f $X=-0.19 $Y=1.655 $X2=1.425 $Y2=2.205
cc_137 VPB N_SCD_M1037_g 0.0434328f $X=-0.19 $Y=1.655 $X2=1.485 $Y2=2.775
cc_138 VPB N_SCD_c_344_n 0.00155411f $X=-0.19 $Y=1.655 $X2=3.17 $Y2=0.505
cc_139 VPB N_SCD_c_345_n 0.037302f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_140 VPB N_SCE_M1021_g 0.0304981f $X=-0.19 $Y=1.655 $X2=1.485 $Y2=2.345
cc_141 VPB N_SCE_M1014_g 0.0296277f $X=-0.19 $Y=1.655 $X2=0.81 $Y2=2.205
cc_142 VPB SCE 0.00805642f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_143 VPB N_SCE_c_404_n 0.0541859f $X=-0.19 $Y=1.655 $X2=3.18 $Y2=2.195
cc_144 VPB N_D_c_466_n 0.00431327f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_145 VPB N_D_M1018_g 0.0483596f $X=-0.19 $Y=1.655 $X2=1.485 $Y2=2.345
cc_146 VPB N_RESET_B_M1000_g 0.0270753f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_147 VPB N_RESET_B_c_525_n 0.020329f $X=-0.19 $Y=1.655 $X2=1.485 $Y2=2.775
cc_148 VPB N_RESET_B_c_526_n 0.0330271f $X=-0.19 $Y=1.655 $X2=0.81 $Y2=2.205
cc_149 VPB N_RESET_B_c_514_n 0.00741429f $X=-0.19 $Y=1.655 $X2=1.425 $Y2=2.36
cc_150 VPB N_RESET_B_M1033_g 0.0461573f $X=-0.19 $Y=1.655 $X2=0.672 $Y2=0.43
cc_151 VPB N_RESET_B_c_516_n 0.00543348f $X=-0.19 $Y=1.655 $X2=1.26 $Y2=2.205
cc_152 VPB N_RESET_B_c_530_n 0.0167579f $X=-0.19 $Y=1.655 $X2=1.26 $Y2=2.13
cc_153 VPB N_RESET_B_c_531_n 0.0262021f $X=-0.19 $Y=1.655 $X2=3.18 $Y2=1.12
cc_154 VPB N_RESET_B_c_532_n 0.0225231f $X=-0.19 $Y=1.655 $X2=3.26 $Y2=1.12
cc_155 VPB N_RESET_B_c_517_n 0.00434666f $X=-0.19 $Y=1.655 $X2=3.26 $Y2=1.12
cc_156 VPB N_RESET_B_c_534_n 0.00627694f $X=-0.19 $Y=1.655 $X2=1.485 $Y2=2.345
cc_157 VPB N_RESET_B_c_535_n 0.00242886f $X=-0.19 $Y=1.655 $X2=3.26 $Y2=0.955
cc_158 VPB N_RESET_B_c_518_n 0.00185497f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_159 VPB N_RESET_B_c_537_n 0.0125732f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_160 VPB N_RESET_B_c_519_n 6.02119e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_161 VPB N_RESET_B_c_520_n 0.0135792f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_162 VPB N_RESET_B_c_540_n 0.0140414f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_163 VPB N_RESET_B_c_541_n 0.00141717f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_164 VPB N_RESET_B_c_542_n 0.00253242f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_165 VPB N_RESET_B_c_543_n 0.00405115f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_166 VPB N_RESET_B_c_544_n 0.0261462f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_167 VPB N_RESET_B_c_521_n 9.18866e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_168 VPB N_RESET_B_c_523_n 0.00172542f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_169 VPB N_CLK_N_M1035_g 0.025954f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_170 VPB N_CLK_N_c_752_n 0.0146659f $X=-0.19 $Y=1.655 $X2=0.672 $Y2=1.815
cc_171 VPB N_CLK_N_c_753_n 0.00272763f $X=-0.19 $Y=1.655 $X2=1.185 $Y2=2.205
cc_172 VPB N_A_1080_47#_M1027_g 0.0348331f $X=-0.19 $Y=1.655 $X2=3.17 $Y2=0.505
cc_173 VPB N_A_1080_47#_M1006_g 0.0203006f $X=-0.19 $Y=1.655 $X2=1.185 $Y2=2.205
cc_174 VPB N_A_1080_47#_c_792_n 0.00322844f $X=-0.19 $Y=1.655 $X2=0.672 $Y2=0.43
cc_175 VPB N_A_1080_47#_c_810_n 0.0066733f $X=-0.19 $Y=1.655 $X2=0.692 $Y2=2.155
cc_176 VPB N_A_1080_47#_c_799_n 0.00191231f $X=-0.19 $Y=1.655 $X2=1.485
+ $Y2=2.345
cc_177 VPB N_A_1080_47#_c_812_n 0.00982522f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_178 VPB N_A_1080_47#_c_813_n 0.00327917f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_179 VPB N_A_1080_47#_c_814_n 0.0348615f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_180 VPB N_A_1080_47#_c_815_n 0.0386757f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_181 VPB N_A_1406_399#_M1036_g 0.0358699f $X=-0.19 $Y=1.655 $X2=1.485
+ $Y2=2.775
cc_182 VPB N_A_1406_399#_M1007_g 0.00966633f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_183 VPB N_A_1406_399#_c_968_n 0.00463061f $X=-0.19 $Y=1.655 $X2=0.81
+ $Y2=2.205
cc_184 VPB N_A_1406_399#_c_975_n 0.0453338f $X=-0.19 $Y=1.655 $X2=2.79 $Y2=2.36
cc_185 VPB N_A_1406_399#_c_971_n 0.00637999f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_186 VPB N_A_1278_529#_M1001_g 0.0220024f $X=-0.19 $Y=1.655 $X2=3.17 $Y2=0.505
cc_187 VPB N_A_1278_529#_c_1058_n 0.0352218f $X=-0.19 $Y=1.655 $X2=0.672
+ $Y2=0.565
cc_188 VPB N_A_1278_529#_c_1059_n 0.0277071f $X=-0.19 $Y=1.655 $X2=0.672
+ $Y2=1.815
cc_189 VPB N_A_1278_529#_c_1060_n 0.0194972f $X=-0.19 $Y=1.655 $X2=1.185
+ $Y2=2.205
cc_190 VPB N_A_1278_529#_c_1061_n 0.00159197f $X=-0.19 $Y=1.655 $X2=0.705
+ $Y2=0.46
cc_191 VPB N_A_1278_529#_c_1056_n 0.00767492f $X=-0.19 $Y=1.655 $X2=0.705
+ $Y2=1.98
cc_192 VPB N_A_1278_529#_c_1063_n 0.00187663f $X=-0.19 $Y=1.655 $X2=3.18
+ $Y2=1.12
cc_193 VPB N_A_1278_529#_c_1064_n 0.0493662f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_194 VPB N_A_1278_529#_c_1065_n 0.00992066f $X=-0.19 $Y=1.655 $X2=1.485
+ $Y2=2.345
cc_195 VPB N_A_1278_529#_c_1066_n 0.00615419f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_196 VPB N_A_1278_529#_c_1067_n 0.0169385f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_197 VPB N_A_857_367#_M1022_g 0.0257951f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_198 VPB N_A_857_367#_c_1172_n 0.0410413f $X=-0.19 $Y=1.655 $X2=2.79 $Y2=2.36
cc_199 VPB N_A_857_367#_c_1187_n 0.019826f $X=-0.19 $Y=1.655 $X2=3.18 $Y2=2.02
cc_200 VPB N_A_857_367#_M1024_g 0.0599841f $X=-0.19 $Y=1.655 $X2=3.26 $Y2=1.12
cc_201 VPB N_A_857_367#_c_1189_n 0.0262737f $X=-0.19 $Y=1.655 $X2=3.26 $Y2=0.955
cc_202 VPB N_A_857_367#_c_1190_n 0.0200026f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_203 VPB N_A_857_367#_c_1183_n 0.00530238f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_204 VPB N_A_2064_101#_M1029_g 0.0238001f $X=-0.19 $Y=1.655 $X2=1.485
+ $Y2=2.775
cc_205 VPB N_A_2064_101#_M1012_g 0.020481f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_206 VPB N_A_2064_101#_c_1326_n 0.00413712f $X=-0.19 $Y=1.655 $X2=0.672
+ $Y2=1.815
cc_207 VPB N_A_2064_101#_c_1327_n 0.0380225f $X=-0.19 $Y=1.655 $X2=2.79 $Y2=2.36
cc_208 VPB N_A_2064_101#_c_1328_n 0.00152771f $X=-0.19 $Y=1.655 $X2=0.672
+ $Y2=0.43
cc_209 VPB N_A_2064_101#_c_1329_n 0.00193255f $X=-0.19 $Y=1.655 $X2=0.705
+ $Y2=0.46
cc_210 VPB N_A_2064_101#_c_1330_n 0.0133437f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_211 VPB N_A_2064_101#_c_1331_n 0.00332407f $X=-0.19 $Y=1.655 $X2=0.692
+ $Y2=2.155
cc_212 VPB N_A_2064_101#_c_1323_n 0.00446731f $X=-0.19 $Y=1.655 $X2=1.425
+ $Y2=2.205
cc_213 VPB N_A_2064_101#_c_1333_n 0.00405935f $X=-0.19 $Y=1.655 $X2=3.18
+ $Y2=2.195
cc_214 VPB N_A_1870_127#_M1013_g 0.0735001f $X=-0.19 $Y=1.655 $X2=3.17 $Y2=0.505
cc_215 VPB N_A_1870_127#_M1004_g 0.0250947f $X=-0.19 $Y=1.655 $X2=3.18 $Y2=1.205
cc_216 VPB N_A_1870_127#_c_1420_n 0.00502547f $X=-0.19 $Y=1.655 $X2=3.18
+ $Y2=1.12
cc_217 VPB N_A_1870_127#_c_1429_n 3.14067e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_218 VPB N_A_2370_351#_M1025_g 0.0294488f $X=-0.19 $Y=1.655 $X2=1.485
+ $Y2=2.775
cc_219 VPB N_A_2370_351#_c_1544_n 0.0144533f $X=-0.19 $Y=1.655 $X2=0.672
+ $Y2=0.565
cc_220 VPB N_A_2370_351#_c_1545_n 0.00311778f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_221 VPB N_A_2370_351#_c_1539_n 0.00555329f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_222 VPB N_A_2370_351#_c_1540_n 0.00302031f $X=-0.19 $Y=1.655 $X2=0.692
+ $Y2=2.155
cc_223 VPB N_A_2370_351#_c_1541_n 0.00320621f $X=-0.19 $Y=1.655 $X2=0.705
+ $Y2=1.98
cc_224 VPB N_VPWR_c_1598_n 0.0113582f $X=-0.19 $Y=1.655 $X2=0.705 $Y2=2.33
cc_225 VPB N_VPWR_c_1599_n 0.0911056f $X=-0.19 $Y=1.655 $X2=1.26 $Y2=2.205
cc_226 VPB N_VPWR_c_1600_n 0.00561719f $X=-0.19 $Y=1.655 $X2=3.18 $Y2=2.195
cc_227 VPB N_VPWR_c_1601_n 0.00883244f $X=-0.19 $Y=1.655 $X2=3.26 $Y2=1.12
cc_228 VPB N_VPWR_c_1602_n 0.00347957f $X=-0.19 $Y=1.655 $X2=3.26 $Y2=1.12
cc_229 VPB N_VPWR_c_1603_n 0.00602232f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_230 VPB N_VPWR_c_1604_n 0.0112102f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_231 VPB N_VPWR_c_1605_n 0.00708349f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_232 VPB N_VPWR_c_1606_n 0.00980965f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_233 VPB N_VPWR_c_1607_n 0.00130851f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_234 VPB N_VPWR_c_1608_n 0.0289797f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_235 VPB N_VPWR_c_1609_n 0.0063198f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_236 VPB N_VPWR_c_1610_n 0.0387988f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_237 VPB N_VPWR_c_1611_n 0.00632279f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_238 VPB N_VPWR_c_1612_n 0.018644f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_239 VPB N_VPWR_c_1613_n 0.00555326f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_240 VPB N_VPWR_c_1614_n 0.016802f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_241 VPB N_VPWR_c_1615_n 0.0065106f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_242 VPB N_VPWR_c_1616_n 0.0241492f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_243 VPB N_VPWR_c_1617_n 0.050384f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_244 VPB N_VPWR_c_1618_n 0.0293304f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_245 VPB N_VPWR_c_1619_n 0.0208865f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_246 VPB N_VPWR_c_1597_n 0.113951f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_247 VPB N_VPWR_c_1621_n 0.0440032f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_248 VPB N_VPWR_c_1622_n 0.0182264f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_249 VPB N_VPWR_c_1623_n 0.00510664f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_250 VPB N_VPWR_c_1624_n 0.00475884f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_251 VPB N_VPWR_c_1625_n 0.0142496f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_252 VPB N_A_229_491#_c_1775_n 0.00155109f $X=-0.19 $Y=1.655 $X2=3.18
+ $Y2=1.205
cc_253 VPB N_A_229_491#_c_1771_n 0.00698395f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_254 VPB N_A_229_491#_c_1777_n 0.0196501f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_255 VPB N_A_229_491#_c_1778_n 0.00641153f $X=-0.19 $Y=1.655 $X2=1.26
+ $Y2=2.205
cc_256 VPB N_A_229_491#_c_1779_n 0.014137f $X=-0.19 $Y=1.655 $X2=1.26 $Y2=2.13
cc_257 VPB N_A_229_491#_c_1780_n 0.00774262f $X=-0.19 $Y=1.655 $X2=1.485
+ $Y2=2.345
cc_258 VPB Q 0.0477912f $X=-0.19 $Y=1.655 $X2=3.17 $Y2=0.505
cc_259 VPB N_Q_c_1923_n 0.00876551f $X=-0.19 $Y=1.655 $X2=0.705 $Y2=0.43
cc_260 VPB N_Q_c_1926_n 0.0140998f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_261 N_A_113_63#_c_270_n N_SCD_M1037_g 0.0137148f $X=2.79 $Y=2.36 $X2=0 $Y2=0
cc_262 N_A_113_63#_c_272_n N_SCD_M1037_g 0.073973f $X=1.26 $Y=2.13 $X2=0 $Y2=0
cc_263 N_A_113_63#_c_273_n N_SCD_M1037_g 0.00147087f $X=1.425 $Y=2.205 $X2=0
+ $Y2=0
cc_264 N_A_113_63#_c_270_n N_SCD_c_344_n 0.0116288f $X=2.79 $Y=2.36 $X2=0 $Y2=0
cc_265 N_A_113_63#_c_270_n N_SCD_c_345_n 0.00242751f $X=2.79 $Y=2.36 $X2=0 $Y2=0
cc_266 N_A_113_63#_c_262_n N_SCD_c_346_n 0.00273378f $X=0.672 $Y=1.815 $X2=0
+ $Y2=0
cc_267 N_A_113_63#_c_262_n N_SCD_c_347_n 0.0273476f $X=0.672 $Y=1.815 $X2=0
+ $Y2=0
cc_268 N_A_113_63#_c_262_n N_SCE_M1039_g 0.0176558f $X=0.672 $Y=1.815 $X2=0
+ $Y2=0
cc_269 N_A_113_63#_c_264_n N_SCE_M1039_g 4.45351e-19 $X=0.705 $Y=0.46 $X2=0
+ $Y2=0
cc_270 N_A_113_63#_c_262_n N_SCE_M1021_g 0.0187148f $X=0.672 $Y=1.815 $X2=0
+ $Y2=0
cc_271 N_A_113_63#_c_262_n N_SCE_c_395_n 0.024008f $X=0.672 $Y=1.815 $X2=0 $Y2=0
cc_272 N_A_113_63#_c_269_n N_SCE_c_395_n 0.00888532f $X=1.185 $Y=2.205 $X2=0
+ $Y2=0
cc_273 N_A_113_63#_c_264_n N_SCE_c_395_n 0.00238483f $X=0.705 $Y=0.46 $X2=0
+ $Y2=0
cc_274 N_A_113_63#_c_272_n N_SCE_c_395_n 0.00758253f $X=1.26 $Y=2.13 $X2=0 $Y2=0
cc_275 N_A_113_63#_c_270_n N_SCE_M1014_g 0.0149942f $X=2.79 $Y=2.36 $X2=0 $Y2=0
cc_276 N_A_113_63#_c_270_n SCE 0.0570264f $X=2.79 $Y=2.36 $X2=0 $Y2=0
cc_277 N_A_113_63#_c_263_n SCE 0.0193845f $X=3.18 $Y=2.02 $X2=0 $Y2=0
cc_278 N_A_113_63#_c_273_n SCE 0.00445333f $X=1.425 $Y=2.205 $X2=0 $Y2=0
cc_279 N_A_113_63#_c_270_n N_SCE_c_404_n 0.0180328f $X=2.79 $Y=2.36 $X2=0 $Y2=0
cc_280 N_A_113_63#_c_263_n N_SCE_c_404_n 6.56813e-19 $X=3.18 $Y=2.02 $X2=0 $Y2=0
cc_281 N_A_113_63#_M1015_g N_D_M1010_g 0.0448884f $X=3.17 $Y=0.505 $X2=0 $Y2=0
cc_282 N_A_113_63#_c_265_n N_D_M1010_g 2.12577e-19 $X=3.26 $Y=1.12 $X2=0 $Y2=0
cc_283 N_A_113_63#_c_270_n N_D_c_466_n 0.00619798f $X=2.79 $Y=2.36 $X2=0 $Y2=0
cc_284 N_A_113_63#_c_263_n N_D_c_466_n 0.0109762f $X=3.18 $Y=2.02 $X2=0 $Y2=0
cc_285 N_A_113_63#_c_265_n N_D_c_466_n 2.04125e-19 $X=3.26 $Y=1.12 $X2=0 $Y2=0
cc_286 N_A_113_63#_c_266_n N_D_c_466_n 0.0179717f $X=3.26 $Y=1.12 $X2=0 $Y2=0
cc_287 N_A_113_63#_c_270_n N_D_M1018_g 0.0166529f $X=2.79 $Y=2.36 $X2=0 $Y2=0
cc_288 N_A_113_63#_c_263_n N_D_M1018_g 0.00794456f $X=3.18 $Y=2.02 $X2=0 $Y2=0
cc_289 N_A_113_63#_c_270_n D 0.00290708f $X=2.79 $Y=2.36 $X2=0 $Y2=0
cc_290 N_A_113_63#_c_263_n D 0.0126329f $X=3.18 $Y=2.02 $X2=0 $Y2=0
cc_291 N_A_113_63#_c_265_n D 0.00858464f $X=3.26 $Y=1.12 $X2=0 $Y2=0
cc_292 N_A_113_63#_c_266_n D 4.53999e-19 $X=3.26 $Y=1.12 $X2=0 $Y2=0
cc_293 N_A_113_63#_M1015_g N_RESET_B_M1034_g 0.0190248f $X=3.17 $Y=0.505 $X2=0
+ $Y2=0
cc_294 N_A_113_63#_c_263_n N_RESET_B_M1034_g 0.00431531f $X=3.18 $Y=2.02 $X2=0
+ $Y2=0
cc_295 N_A_113_63#_c_265_n N_RESET_B_M1034_g 6.05555e-19 $X=3.26 $Y=1.12 $X2=0
+ $Y2=0
cc_296 N_A_113_63#_c_266_n N_RESET_B_M1034_g 0.0203459f $X=3.26 $Y=1.12 $X2=0
+ $Y2=0
cc_297 N_A_113_63#_c_263_n N_RESET_B_c_516_n 0.0031056f $X=3.18 $Y=2.02 $X2=0
+ $Y2=0
cc_298 N_A_113_63#_c_265_n N_RESET_B_c_516_n 2.86732e-19 $X=3.26 $Y=1.12 $X2=0
+ $Y2=0
cc_299 N_A_113_63#_c_266_n N_RESET_B_c_516_n 0.00282203f $X=3.26 $Y=1.12 $X2=0
+ $Y2=0
cc_300 N_A_113_63#_c_270_n N_RESET_B_c_541_n 0.00362369f $X=2.79 $Y=2.36 $X2=0
+ $Y2=0
cc_301 N_A_113_63#_c_263_n N_RESET_B_c_541_n 0.00268572f $X=3.18 $Y=2.02 $X2=0
+ $Y2=0
cc_302 N_A_113_63#_c_270_n N_RESET_B_c_544_n 0.0012146f $X=2.79 $Y=2.36 $X2=0
+ $Y2=0
cc_303 N_A_113_63#_c_270_n N_RESET_B_c_521_n 0.0109444f $X=2.79 $Y=2.36 $X2=0
+ $Y2=0
cc_304 N_A_113_63#_c_263_n N_RESET_B_c_521_n 0.0314817f $X=3.18 $Y=2.02 $X2=0
+ $Y2=0
cc_305 N_A_113_63#_c_262_n N_VPWR_c_1599_n 0.00307081f $X=0.672 $Y=1.815 $X2=0
+ $Y2=0
cc_306 N_A_113_63#_c_267_n N_VPWR_c_1597_n 0.00698426f $X=1.485 $Y=2.345 $X2=0
+ $Y2=0
cc_307 N_A_113_63#_c_262_n N_VPWR_c_1597_n 0.00928629f $X=0.672 $Y=1.815 $X2=0
+ $Y2=0
cc_308 N_A_113_63#_c_267_n N_VPWR_c_1621_n 0.00407336f $X=1.485 $Y=2.345 $X2=0
+ $Y2=0
cc_309 N_A_113_63#_c_267_n N_A_229_491#_c_1781_n 0.00822819f $X=1.485 $Y=2.345
+ $X2=0 $Y2=0
cc_310 N_A_113_63#_c_270_n N_A_229_491#_c_1781_n 0.108587f $X=2.79 $Y=2.36 $X2=0
+ $Y2=0
cc_311 N_A_113_63#_M1015_g N_A_229_491#_c_1770_n 0.0112884f $X=3.17 $Y=0.505
+ $X2=0 $Y2=0
cc_312 N_A_113_63#_c_265_n N_A_229_491#_c_1770_n 0.0220435f $X=3.26 $Y=1.12
+ $X2=0 $Y2=0
cc_313 N_A_113_63#_c_266_n N_A_229_491#_c_1770_n 0.00440824f $X=3.26 $Y=1.12
+ $X2=0 $Y2=0
cc_314 N_A_113_63#_c_263_n N_A_229_491#_c_1771_n 0.00963159f $X=3.18 $Y=2.02
+ $X2=0 $Y2=0
cc_315 N_A_113_63#_c_265_n N_A_229_491#_c_1771_n 0.00618731f $X=3.26 $Y=1.12
+ $X2=0 $Y2=0
cc_316 N_A_113_63#_c_267_n N_A_229_491#_c_1779_n 0.00462341f $X=1.485 $Y=2.345
+ $X2=0 $Y2=0
cc_317 N_A_113_63#_c_269_n N_A_229_491#_c_1779_n 0.0253235f $X=1.185 $Y=2.205
+ $X2=0 $Y2=0
cc_318 N_A_113_63#_c_272_n N_A_229_491#_c_1779_n 0.00164817f $X=1.26 $Y=2.13
+ $X2=0 $Y2=0
cc_319 N_A_113_63#_c_270_n N_A_229_491#_c_1780_n 0.0120624f $X=2.79 $Y=2.36
+ $X2=0 $Y2=0
cc_320 N_A_113_63#_c_264_n N_VGND_c_1943_n 0.00147947f $X=0.705 $Y=0.46 $X2=0
+ $Y2=0
cc_321 N_A_113_63#_M1015_g N_VGND_c_1949_n 0.00321654f $X=3.17 $Y=0.505 $X2=0
+ $Y2=0
cc_322 N_A_113_63#_c_264_n N_VGND_c_1949_n 0.0156922f $X=0.705 $Y=0.46 $X2=0
+ $Y2=0
cc_323 N_A_113_63#_M1015_g N_VGND_c_1955_n 0.00492419f $X=3.17 $Y=0.505 $X2=0
+ $Y2=0
cc_324 N_A_113_63#_c_264_n N_VGND_c_1955_n 0.0109469f $X=0.705 $Y=0.46 $X2=0
+ $Y2=0
cc_325 N_A_113_63#_c_264_n N_noxref_24_c_2073_n 0.0100505f $X=0.705 $Y=0.46
+ $X2=0 $Y2=0
cc_326 N_A_113_63#_M1015_g N_noxref_24_c_2074_n 0.00270664f $X=3.17 $Y=0.505
+ $X2=0 $Y2=0
cc_327 N_A_113_63#_M1015_g N_noxref_24_c_2075_n 0.00689373f $X=3.17 $Y=0.505
+ $X2=0 $Y2=0
cc_328 N_SCD_c_346_n N_SCE_M1039_g 0.0083031f $X=1.28 $Y=0.83 $X2=0 $Y2=0
cc_329 N_SCD_c_341_n N_SCE_c_395_n 0.0241956f $X=1.655 $Y=0.9 $X2=0 $Y2=0
cc_330 N_SCD_c_344_n N_SCE_c_395_n 0.0184279f $X=1.8 $Y=1.79 $X2=0 $Y2=0
cc_331 N_SCD_c_345_n N_SCE_c_395_n 0.0191823f $X=1.8 $Y=1.79 $X2=0 $Y2=0
cc_332 N_SCD_c_346_n N_SCE_c_395_n 0.0163795f $X=1.28 $Y=0.83 $X2=0 $Y2=0
cc_333 N_SCD_c_347_n N_SCE_c_395_n 0.0167835f $X=1.64 $Y=0.92 $X2=0 $Y2=0
cc_334 N_SCD_c_342_n N_SCE_M1028_g 0.0507507f $X=1.73 $Y=0.825 $X2=0 $Y2=0
cc_335 N_SCD_c_343_n N_SCE_M1028_g 0.00881416f $X=1.762 $Y=1.095 $X2=0 $Y2=0
cc_336 N_SCD_c_343_n N_SCE_c_398_n 0.00333965f $X=1.762 $Y=1.095 $X2=0 $Y2=0
cc_337 N_SCD_c_344_n N_SCE_c_398_n 0.0368043f $X=1.8 $Y=1.79 $X2=0 $Y2=0
cc_338 N_SCD_c_344_n N_SCE_c_399_n 0.00331679f $X=1.8 $Y=1.79 $X2=0 $Y2=0
cc_339 N_SCD_M1037_g SCE 0.00213158f $X=1.845 $Y=2.775 $X2=0 $Y2=0
cc_340 N_SCD_c_344_n SCE 0.0314682f $X=1.8 $Y=1.79 $X2=0 $Y2=0
cc_341 N_SCD_c_345_n SCE 0.00665323f $X=1.8 $Y=1.79 $X2=0 $Y2=0
cc_342 N_SCD_M1037_g N_SCE_c_404_n 0.0104039f $X=1.845 $Y=2.775 $X2=0 $Y2=0
cc_343 N_SCD_c_345_n N_SCE_c_404_n 0.00521913f $X=1.8 $Y=1.79 $X2=0 $Y2=0
cc_344 N_SCD_M1037_g N_VPWR_c_1597_n 0.00686971f $X=1.845 $Y=2.775 $X2=0 $Y2=0
cc_345 N_SCD_M1037_g N_VPWR_c_1621_n 0.00411233f $X=1.845 $Y=2.775 $X2=0 $Y2=0
cc_346 N_SCD_M1037_g N_VPWR_c_1622_n 0.00768714f $X=1.845 $Y=2.775 $X2=0 $Y2=0
cc_347 N_SCD_M1037_g N_A_229_491#_c_1781_n 0.0129844f $X=1.845 $Y=2.775 $X2=0
+ $Y2=0
cc_348 N_SCD_M1037_g N_A_229_491#_c_1779_n 9.5959e-19 $X=1.845 $Y=2.775 $X2=0
+ $Y2=0
cc_349 N_SCD_c_343_n N_A_229_491#_c_1773_n 0.00591481f $X=1.762 $Y=1.095 $X2=0
+ $Y2=0
cc_350 N_SCD_c_342_n N_VGND_c_1949_n 0.00322088f $X=1.73 $Y=0.825 $X2=0 $Y2=0
cc_351 N_SCD_c_346_n N_VGND_c_1949_n 0.00503617f $X=1.28 $Y=0.83 $X2=0 $Y2=0
cc_352 N_SCD_c_347_n N_VGND_c_1949_n 0.00553491f $X=1.64 $Y=0.92 $X2=0 $Y2=0
cc_353 N_SCD_c_342_n N_VGND_c_1955_n 0.00545377f $X=1.73 $Y=0.825 $X2=0 $Y2=0
cc_354 N_SCD_c_343_n N_VGND_c_1955_n 7.91752e-19 $X=1.762 $Y=1.095 $X2=0 $Y2=0
cc_355 N_SCD_c_346_n N_VGND_c_1955_n 0.00828758f $X=1.28 $Y=0.83 $X2=0 $Y2=0
cc_356 N_SCD_c_347_n N_VGND_c_1955_n 0.0110843f $X=1.64 $Y=0.92 $X2=0 $Y2=0
cc_357 N_SCD_c_341_n N_noxref_24_c_2073_n 0.00168381f $X=1.655 $Y=0.9 $X2=0
+ $Y2=0
cc_358 N_SCD_c_342_n N_noxref_24_c_2073_n 0.00389622f $X=1.73 $Y=0.825 $X2=0
+ $Y2=0
cc_359 N_SCD_c_343_n N_noxref_24_c_2073_n 0.00210636f $X=1.762 $Y=1.095 $X2=0
+ $Y2=0
cc_360 N_SCD_c_347_n N_noxref_24_c_2073_n 0.0183778f $X=1.64 $Y=0.92 $X2=0 $Y2=0
cc_361 N_SCD_c_342_n N_noxref_24_c_2075_n 0.00733238f $X=1.73 $Y=0.825 $X2=0
+ $Y2=0
cc_362 N_SCD_c_343_n N_noxref_24_c_2075_n 0.00754899f $X=1.762 $Y=1.095 $X2=0
+ $Y2=0
cc_363 N_SCE_M1028_g N_D_M1010_g 0.0205076f $X=2.09 $Y=0.505 $X2=0 $Y2=0
cc_364 N_SCE_c_399_n N_D_M1010_g 5.88217e-19 $X=2.18 $Y=1.22 $X2=0 $Y2=0
cc_365 N_SCE_c_398_n N_D_c_466_n 0.00560173f $X=2.18 $Y=1.22 $X2=0 $Y2=0
cc_366 N_SCE_c_399_n N_D_c_466_n 0.0202498f $X=2.18 $Y=1.22 $X2=0 $Y2=0
cc_367 SCE N_D_c_466_n 0.00612149f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_368 N_SCE_c_404_n N_D_c_466_n 0.00551041f $X=2.37 $Y=2.02 $X2=0 $Y2=0
cc_369 SCE N_D_M1018_g 0.00427346f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_370 N_SCE_c_404_n N_D_M1018_g 0.0797826f $X=2.37 $Y=2.02 $X2=0 $Y2=0
cc_371 N_SCE_c_398_n D 0.0265515f $X=2.18 $Y=1.22 $X2=0 $Y2=0
cc_372 N_SCE_c_399_n D 0.00190231f $X=2.18 $Y=1.22 $X2=0 $Y2=0
cc_373 SCE D 0.022775f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_374 N_SCE_c_404_n D 3.67187e-19 $X=2.37 $Y=2.02 $X2=0 $Y2=0
cc_375 N_SCE_M1021_g N_VPWR_c_1599_n 0.00573078f $X=0.49 $Y=2.155 $X2=0 $Y2=0
cc_376 N_SCE_M1014_g N_VPWR_c_1608_n 0.00411233f $X=2.735 $Y=2.775 $X2=0 $Y2=0
cc_377 N_SCE_M1021_g N_VPWR_c_1597_n 0.00410284f $X=0.49 $Y=2.155 $X2=0 $Y2=0
cc_378 N_SCE_M1014_g N_VPWR_c_1597_n 0.00686971f $X=2.735 $Y=2.775 $X2=0 $Y2=0
cc_379 N_SCE_M1021_g N_VPWR_c_1621_n 0.00312414f $X=0.49 $Y=2.155 $X2=0 $Y2=0
cc_380 N_SCE_M1014_g N_VPWR_c_1622_n 0.00768714f $X=2.735 $Y=2.775 $X2=0 $Y2=0
cc_381 N_SCE_M1014_g N_A_229_491#_c_1781_n 0.0129836f $X=2.735 $Y=2.775 $X2=0
+ $Y2=0
cc_382 N_SCE_M1028_g N_A_229_491#_c_1773_n 0.00572407f $X=2.09 $Y=0.505 $X2=0
+ $Y2=0
cc_383 N_SCE_c_398_n N_A_229_491#_c_1773_n 0.00610527f $X=2.18 $Y=1.22 $X2=0
+ $Y2=0
cc_384 N_SCE_c_399_n N_A_229_491#_c_1773_n 8.18125e-19 $X=2.18 $Y=1.22 $X2=0
+ $Y2=0
cc_385 N_SCE_M1039_g N_VGND_c_1943_n 0.0052018f $X=0.49 $Y=0.525 $X2=0 $Y2=0
cc_386 N_SCE_M1039_g N_VGND_c_1949_n 0.00508422f $X=0.49 $Y=0.525 $X2=0 $Y2=0
cc_387 N_SCE_M1028_g N_VGND_c_1949_n 0.00321654f $X=2.09 $Y=0.505 $X2=0 $Y2=0
cc_388 N_SCE_M1039_g N_VGND_c_1955_n 0.0108828f $X=0.49 $Y=0.525 $X2=0 $Y2=0
cc_389 N_SCE_M1028_g N_VGND_c_1955_n 0.00495964f $X=2.09 $Y=0.505 $X2=0 $Y2=0
cc_390 N_SCE_M1028_g N_noxref_24_c_2073_n 6.28332e-19 $X=2.09 $Y=0.505 $X2=0
+ $Y2=0
cc_391 N_SCE_M1028_g N_noxref_24_c_2075_n 0.0128444f $X=2.09 $Y=0.505 $X2=0
+ $Y2=0
cc_392 N_SCE_c_398_n N_noxref_24_c_2075_n 0.00457627f $X=2.18 $Y=1.22 $X2=0
+ $Y2=0
cc_393 N_SCE_c_399_n N_noxref_24_c_2075_n 3.53301e-19 $X=2.18 $Y=1.22 $X2=0
+ $Y2=0
cc_394 N_D_M1018_g N_RESET_B_M1000_g 0.0192608f $X=3.095 $Y=2.775 $X2=0 $Y2=0
cc_395 N_D_c_466_n N_RESET_B_M1034_g 3.78951e-19 $X=3.095 $Y=1.675 $X2=0 $Y2=0
cc_396 N_D_c_466_n N_RESET_B_c_516_n 0.0207722f $X=3.095 $Y=1.675 $X2=0 $Y2=0
cc_397 N_D_M1018_g N_RESET_B_c_544_n 0.0207722f $X=3.095 $Y=2.775 $X2=0 $Y2=0
cc_398 N_D_c_466_n N_RESET_B_c_521_n 7.47921e-19 $X=3.095 $Y=1.675 $X2=0 $Y2=0
cc_399 N_D_M1018_g N_VPWR_c_1608_n 0.00411233f $X=3.095 $Y=2.775 $X2=0 $Y2=0
cc_400 N_D_M1018_g N_VPWR_c_1597_n 0.00584183f $X=3.095 $Y=2.775 $X2=0 $Y2=0
cc_401 N_D_M1018_g N_A_229_491#_c_1781_n 0.0101952f $X=3.095 $Y=2.775 $X2=0
+ $Y2=0
cc_402 N_D_M1010_g N_A_229_491#_c_1770_n 0.0118256f $X=2.75 $Y=0.505 $X2=0 $Y2=0
cc_403 N_D_c_466_n N_A_229_491#_c_1770_n 0.00623987f $X=3.095 $Y=1.675 $X2=0
+ $Y2=0
cc_404 N_D_M1010_g N_A_229_491#_c_1773_n 0.00225985f $X=2.75 $Y=0.505 $X2=0
+ $Y2=0
cc_405 N_D_c_466_n N_A_229_491#_c_1773_n 0.00261586f $X=3.095 $Y=1.675 $X2=0
+ $Y2=0
cc_406 D N_A_229_491#_c_1773_n 0.0233885f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_407 N_D_M1018_g N_A_229_491#_c_1780_n 0.00111668f $X=3.095 $Y=2.775 $X2=0
+ $Y2=0
cc_408 N_D_M1010_g N_VGND_c_1949_n 0.00321654f $X=2.75 $Y=0.505 $X2=0 $Y2=0
cc_409 N_D_M1010_g N_VGND_c_1955_n 0.00505612f $X=2.75 $Y=0.505 $X2=0 $Y2=0
cc_410 N_D_M1010_g N_noxref_24_c_2074_n 3.87543e-19 $X=2.75 $Y=0.505 $X2=0 $Y2=0
cc_411 N_D_M1010_g N_noxref_24_c_2075_n 0.0109254f $X=2.75 $Y=0.505 $X2=0 $Y2=0
cc_412 N_RESET_B_c_540_n N_CLK_N_M1035_g 0.0094764f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_413 N_RESET_B_c_544_n N_CLK_N_M1035_g 0.0368476f $X=3.545 $Y=1.69 $X2=0 $Y2=0
cc_414 N_RESET_B_M1034_g N_CLK_N_M1023_g 0.0219772f $X=3.71 $Y=0.505 $X2=0 $Y2=0
cc_415 N_RESET_B_M1034_g N_CLK_N_c_752_n 0.00508257f $X=3.71 $Y=0.505 $X2=0
+ $Y2=0
cc_416 N_RESET_B_c_516_n N_CLK_N_c_752_n 0.00521643f $X=3.597 $Y=1.675 $X2=0
+ $Y2=0
cc_417 N_RESET_B_c_540_n N_CLK_N_c_752_n 8.88908e-19 $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_418 N_RESET_B_c_540_n N_CLK_N_c_753_n 0.00127188f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_419 N_RESET_B_c_571_p N_A_1080_47#_M1006_g 0.0135215f $X=10.145 $Y=2.99 $X2=0
+ $Y2=0
cc_420 N_RESET_B_c_572_p N_A_1080_47#_M1006_g 0.004484f $X=9.18 $Y=2.72 $X2=0
+ $Y2=0
cc_421 N_RESET_B_c_540_n N_A_1080_47#_c_792_n 0.0022777f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_422 N_RESET_B_c_540_n N_A_1080_47#_c_810_n 0.0268885f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_423 N_RESET_B_M1009_g N_A_1080_47#_c_820_n 0.0119976f $X=7.83 $Y=0.845 $X2=0
+ $Y2=0
cc_424 N_RESET_B_c_540_n N_A_1080_47#_c_812_n 0.0413987f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_425 N_RESET_B_c_540_n N_A_1080_47#_c_815_n 0.00437533f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_426 N_RESET_B_c_571_p N_A_1406_399#_M1038_d 0.00336733f $X=10.145 $Y=2.99
+ $X2=0 $Y2=0
cc_427 N_RESET_B_c_572_p N_A_1406_399#_M1038_d 0.00460686f $X=9.18 $Y=2.72 $X2=0
+ $Y2=0
cc_428 N_RESET_B_c_526_n N_A_1406_399#_M1036_g 0.0057168f $X=7.83 $Y=2.385 $X2=0
+ $Y2=0
cc_429 N_RESET_B_c_531_n N_A_1406_399#_M1036_g 0.0192425f $X=7.83 $Y=2.46 $X2=0
+ $Y2=0
cc_430 N_RESET_B_M1009_g N_A_1406_399#_M1007_g 0.0510636f $X=7.83 $Y=0.845 $X2=0
+ $Y2=0
cc_431 N_RESET_B_c_519_n N_A_1406_399#_M1007_g 9.46926e-19 $X=7.89 $Y=1.745
+ $X2=0 $Y2=0
cc_432 N_RESET_B_c_543_n N_A_1406_399#_M1007_g 0.00140383f $X=7.92 $Y=2.035
+ $X2=0 $Y2=0
cc_433 N_RESET_B_M1009_g N_A_1406_399#_c_968_n 0.00113589f $X=7.83 $Y=0.845
+ $X2=0 $Y2=0
cc_434 N_RESET_B_c_526_n N_A_1406_399#_c_968_n 0.00122646f $X=7.83 $Y=2.385
+ $X2=0 $Y2=0
cc_435 N_RESET_B_c_519_n N_A_1406_399#_c_968_n 0.0212145f $X=7.89 $Y=1.745 $X2=0
+ $Y2=0
cc_436 N_RESET_B_c_520_n N_A_1406_399#_c_968_n 3.96797e-19 $X=8 $Y=1.58 $X2=0
+ $Y2=0
cc_437 N_RESET_B_c_540_n N_A_1406_399#_c_968_n 0.0296998f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_438 N_RESET_B_c_542_n N_A_1406_399#_c_968_n 5.83524e-19 $X=7.92 $Y=2.035
+ $X2=0 $Y2=0
cc_439 N_RESET_B_c_543_n N_A_1406_399#_c_968_n 0.0227583f $X=7.92 $Y=2.035 $X2=0
+ $Y2=0
cc_440 N_RESET_B_c_531_n N_A_1406_399#_c_975_n 0.00472229f $X=7.83 $Y=2.46 $X2=0
+ $Y2=0
cc_441 N_RESET_B_c_520_n N_A_1406_399#_c_975_n 0.0510636f $X=8 $Y=1.58 $X2=0
+ $Y2=0
cc_442 N_RESET_B_c_540_n N_A_1406_399#_c_975_n 0.00637976f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_443 N_RESET_B_M1009_g N_A_1406_399#_c_969_n 0.0126253f $X=7.83 $Y=0.845 $X2=0
+ $Y2=0
cc_444 N_RESET_B_c_517_n N_A_1406_399#_c_969_n 0.0505416f $X=8.545 $Y=1.587
+ $X2=0 $Y2=0
cc_445 N_RESET_B_c_519_n N_A_1406_399#_c_969_n 0.0212588f $X=7.89 $Y=1.745 $X2=0
+ $Y2=0
cc_446 N_RESET_B_c_520_n N_A_1406_399#_c_969_n 0.00595368f $X=8 $Y=1.58 $X2=0
+ $Y2=0
cc_447 N_RESET_B_c_517_n N_A_1406_399#_c_971_n 0.0218424f $X=8.545 $Y=1.587
+ $X2=0 $Y2=0
cc_448 N_RESET_B_c_534_n N_A_1406_399#_c_971_n 0.0309074f $X=8.63 $Y=2.635 $X2=0
+ $Y2=0
cc_449 N_RESET_B_c_534_n N_A_1406_399#_c_1000_n 0.0129318f $X=8.63 $Y=2.635
+ $X2=0 $Y2=0
cc_450 N_RESET_B_c_602_p N_A_1406_399#_c_1000_n 0.0072788f $X=9.095 $Y=2.72
+ $X2=0 $Y2=0
cc_451 N_RESET_B_c_572_p N_A_1406_399#_c_1000_n 0.00108073f $X=9.18 $Y=2.72
+ $X2=0 $Y2=0
cc_452 N_RESET_B_c_571_p N_A_1406_399#_c_1003_n 0.00489924f $X=10.145 $Y=2.99
+ $X2=0 $Y2=0
cc_453 N_RESET_B_c_572_p N_A_1406_399#_c_1003_n 0.00740686f $X=9.18 $Y=2.72
+ $X2=0 $Y2=0
cc_454 N_RESET_B_M1009_g N_A_1278_529#_M1001_g 0.0167491f $X=7.83 $Y=0.845 $X2=0
+ $Y2=0
cc_455 N_RESET_B_c_526_n N_A_1278_529#_M1001_g 0.00300142f $X=7.83 $Y=2.385
+ $X2=0 $Y2=0
cc_456 N_RESET_B_c_517_n N_A_1278_529#_M1001_g 0.0149041f $X=8.545 $Y=1.587
+ $X2=0 $Y2=0
cc_457 N_RESET_B_c_534_n N_A_1278_529#_M1001_g 0.0087214f $X=8.63 $Y=2.635 $X2=0
+ $Y2=0
cc_458 N_RESET_B_c_520_n N_A_1278_529#_M1001_g 0.0102878f $X=8 $Y=1.58 $X2=0
+ $Y2=0
cc_459 N_RESET_B_c_542_n N_A_1278_529#_M1001_g 9.67442e-19 $X=7.92 $Y=2.035
+ $X2=0 $Y2=0
cc_460 N_RESET_B_c_543_n N_A_1278_529#_M1001_g 0.00163058f $X=7.92 $Y=2.035
+ $X2=0 $Y2=0
cc_461 N_RESET_B_c_534_n N_A_1278_529#_c_1058_n 0.0037292f $X=8.63 $Y=2.635
+ $X2=0 $Y2=0
cc_462 N_RESET_B_c_602_p N_A_1278_529#_c_1058_n 0.00483221f $X=9.095 $Y=2.72
+ $X2=0 $Y2=0
cc_463 N_RESET_B_c_526_n N_A_1278_529#_c_1059_n 0.0177866f $X=7.83 $Y=2.385
+ $X2=0 $Y2=0
cc_464 N_RESET_B_c_517_n N_A_1278_529#_c_1059_n 0.00909251f $X=8.545 $Y=1.587
+ $X2=0 $Y2=0
cc_465 N_RESET_B_c_534_n N_A_1278_529#_c_1059_n 0.00742355f $X=8.63 $Y=2.635
+ $X2=0 $Y2=0
cc_466 N_RESET_B_c_520_n N_A_1278_529#_c_1059_n 0.00292537f $X=8 $Y=1.58 $X2=0
+ $Y2=0
cc_467 N_RESET_B_c_542_n N_A_1278_529#_c_1059_n 0.00338595f $X=7.92 $Y=2.035
+ $X2=0 $Y2=0
cc_468 N_RESET_B_c_543_n N_A_1278_529#_c_1059_n 0.0012688f $X=7.92 $Y=2.035
+ $X2=0 $Y2=0
cc_469 N_RESET_B_c_534_n N_A_1278_529#_c_1060_n 0.00452544f $X=8.63 $Y=2.635
+ $X2=0 $Y2=0
cc_470 N_RESET_B_c_602_p N_A_1278_529#_c_1060_n 0.00851662f $X=9.095 $Y=2.72
+ $X2=0 $Y2=0
cc_471 N_RESET_B_c_571_p N_A_1278_529#_c_1060_n 2.26329e-19 $X=10.145 $Y=2.99
+ $X2=0 $Y2=0
cc_472 N_RESET_B_c_572_p N_A_1278_529#_c_1060_n 0.0145981f $X=9.18 $Y=2.72 $X2=0
+ $Y2=0
cc_473 N_RESET_B_c_540_n N_A_1278_529#_c_1056_n 0.0139273f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_474 N_RESET_B_c_526_n N_A_1278_529#_c_1063_n 0.00111991f $X=7.83 $Y=2.385
+ $X2=0 $Y2=0
cc_475 N_RESET_B_c_517_n N_A_1278_529#_c_1063_n 0.0109695f $X=8.545 $Y=1.587
+ $X2=0 $Y2=0
cc_476 N_RESET_B_c_534_n N_A_1278_529#_c_1063_n 0.0251889f $X=8.63 $Y=2.635
+ $X2=0 $Y2=0
cc_477 N_RESET_B_c_542_n N_A_1278_529#_c_1063_n 0.00543717f $X=7.92 $Y=2.035
+ $X2=0 $Y2=0
cc_478 N_RESET_B_c_543_n N_A_1278_529#_c_1063_n 0.0126097f $X=7.92 $Y=2.035
+ $X2=0 $Y2=0
cc_479 N_RESET_B_c_525_n N_A_1278_529#_c_1064_n 0.00197737f $X=7.535 $Y=2.535
+ $X2=0 $Y2=0
cc_480 N_RESET_B_c_531_n N_A_1278_529#_c_1064_n 0.0177866f $X=7.83 $Y=2.46 $X2=0
+ $Y2=0
cc_481 N_RESET_B_c_534_n N_A_1278_529#_c_1064_n 0.00537706f $X=8.63 $Y=2.635
+ $X2=0 $Y2=0
cc_482 N_RESET_B_c_535_n N_A_1278_529#_c_1064_n 2.30674e-19 $X=8.715 $Y=2.72
+ $X2=0 $Y2=0
cc_483 N_RESET_B_c_540_n N_A_1278_529#_c_1065_n 0.00883728f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_484 N_RESET_B_c_531_n N_A_1278_529#_c_1066_n 0.00875772f $X=7.83 $Y=2.46
+ $X2=0 $Y2=0
cc_485 N_RESET_B_c_540_n N_A_1278_529#_c_1066_n 0.0198349f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_486 N_RESET_B_c_525_n N_A_1278_529#_c_1067_n 0.00411693f $X=7.535 $Y=2.535
+ $X2=0 $Y2=0
cc_487 N_RESET_B_c_526_n N_A_1278_529#_c_1067_n 0.00347304f $X=7.83 $Y=2.385
+ $X2=0 $Y2=0
cc_488 N_RESET_B_c_531_n N_A_1278_529#_c_1067_n 0.0137629f $X=7.83 $Y=2.46 $X2=0
+ $Y2=0
cc_489 N_RESET_B_c_517_n N_A_1278_529#_c_1067_n 0.00447308f $X=8.545 $Y=1.587
+ $X2=0 $Y2=0
cc_490 N_RESET_B_c_534_n N_A_1278_529#_c_1067_n 0.0226564f $X=8.63 $Y=2.635
+ $X2=0 $Y2=0
cc_491 N_RESET_B_c_535_n N_A_1278_529#_c_1067_n 0.0155904f $X=8.715 $Y=2.72
+ $X2=0 $Y2=0
cc_492 N_RESET_B_c_520_n N_A_1278_529#_c_1067_n 0.00204313f $X=8 $Y=1.58 $X2=0
+ $Y2=0
cc_493 N_RESET_B_c_542_n N_A_1278_529#_c_1067_n 0.00333404f $X=7.92 $Y=2.035
+ $X2=0 $Y2=0
cc_494 N_RESET_B_c_543_n N_A_1278_529#_c_1067_n 0.0215634f $X=7.92 $Y=2.035
+ $X2=0 $Y2=0
cc_495 N_RESET_B_c_540_n N_A_857_367#_M1035_d 8.52718e-19 $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_496 N_RESET_B_c_540_n N_A_857_367#_M1022_g 0.00977478f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_497 N_RESET_B_c_540_n N_A_857_367#_c_1173_n 0.00259255f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_498 N_RESET_B_M1009_g N_A_857_367#_c_1175_n 0.00807149f $X=7.83 $Y=0.845
+ $X2=0 $Y2=0
cc_499 N_RESET_B_c_518_n N_A_857_367#_c_1178_n 0.00457361f $X=10.23 $Y=1.965
+ $X2=0 $Y2=0
cc_500 N_RESET_B_c_571_p N_A_857_367#_M1024_g 0.0136259f $X=10.145 $Y=2.99 $X2=0
+ $Y2=0
cc_501 N_RESET_B_c_537_n N_A_857_367#_M1024_g 0.00533439f $X=10.23 $Y=2.905
+ $X2=0 $Y2=0
cc_502 N_RESET_B_c_540_n N_A_857_367#_c_1190_n 0.0532227f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_503 N_RESET_B_c_540_n N_A_857_367#_c_1184_n 7.79575e-19 $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_504 N_RESET_B_M1033_g N_A_2064_101#_M1029_g 0.00546707f $X=11.03 $Y=2.875
+ $X2=0 $Y2=0
cc_505 N_RESET_B_M1002_g N_A_2064_101#_M1029_g 0.0158993f $X=11.055 $Y=0.845
+ $X2=0 $Y2=0
cc_506 N_RESET_B_c_537_n N_A_2064_101#_M1029_g 0.0124636f $X=10.23 $Y=2.905
+ $X2=0 $Y2=0
cc_507 N_RESET_B_c_522_n N_A_2064_101#_M1029_g 0.0373897f $X=10.875 $Y=1.46
+ $X2=0 $Y2=0
cc_508 N_RESET_B_c_523_n N_A_2064_101#_M1029_g 0.0280023f $X=10.875 $Y=1.46
+ $X2=0 $Y2=0
cc_509 N_RESET_B_M1033_g N_A_2064_101#_M1012_g 0.0134546f $X=11.03 $Y=2.875
+ $X2=0 $Y2=0
cc_510 N_RESET_B_M1033_g N_A_2064_101#_c_1326_n 0.0131492f $X=11.03 $Y=2.875
+ $X2=0 $Y2=0
cc_511 N_RESET_B_c_532_n N_A_2064_101#_c_1326_n 0.00552356f $X=10.92 $Y=1.965
+ $X2=0 $Y2=0
cc_512 N_RESET_B_c_537_n N_A_2064_101#_c_1326_n 0.0250925f $X=10.23 $Y=2.905
+ $X2=0 $Y2=0
cc_513 N_RESET_B_c_523_n N_A_2064_101#_c_1326_n 0.038002f $X=10.875 $Y=1.46
+ $X2=0 $Y2=0
cc_514 N_RESET_B_M1033_g N_A_2064_101#_c_1327_n 0.0213635f $X=11.03 $Y=2.875
+ $X2=0 $Y2=0
cc_515 N_RESET_B_c_532_n N_A_2064_101#_c_1327_n 0.00225346f $X=10.92 $Y=1.965
+ $X2=0 $Y2=0
cc_516 N_RESET_B_c_523_n N_A_2064_101#_c_1327_n 0.00602838f $X=10.875 $Y=1.46
+ $X2=0 $Y2=0
cc_517 N_RESET_B_M1033_g N_A_2064_101#_c_1328_n 0.0104589f $X=11.03 $Y=2.875
+ $X2=0 $Y2=0
cc_518 N_RESET_B_M1033_g N_A_2064_101#_c_1329_n 0.00460684f $X=11.03 $Y=2.875
+ $X2=0 $Y2=0
cc_519 N_RESET_B_c_532_n N_A_2064_101#_c_1331_n 0.00143848f $X=10.92 $Y=1.965
+ $X2=0 $Y2=0
cc_520 N_RESET_B_c_523_n N_A_2064_101#_c_1331_n 0.0144899f $X=10.875 $Y=1.46
+ $X2=0 $Y2=0
cc_521 N_RESET_B_M1002_g N_A_2064_101#_c_1322_n 7.45426e-19 $X=11.055 $Y=0.845
+ $X2=0 $Y2=0
cc_522 N_RESET_B_M1033_g N_A_2064_101#_c_1333_n 0.0059248f $X=11.03 $Y=2.875
+ $X2=0 $Y2=0
cc_523 N_RESET_B_c_532_n N_A_2064_101#_c_1333_n 0.00115863f $X=10.92 $Y=1.965
+ $X2=0 $Y2=0
cc_524 N_RESET_B_c_571_p N_A_1870_127#_M1006_d 0.00537165f $X=10.145 $Y=2.99
+ $X2=0 $Y2=0
cc_525 N_RESET_B_M1033_g N_A_1870_127#_M1013_g 0.0374387f $X=11.03 $Y=2.875
+ $X2=0 $Y2=0
cc_526 N_RESET_B_c_522_n N_A_1870_127#_M1013_g 0.0235682f $X=10.875 $Y=1.46
+ $X2=0 $Y2=0
cc_527 N_RESET_B_c_523_n N_A_1870_127#_M1013_g 0.00170172f $X=10.875 $Y=1.46
+ $X2=0 $Y2=0
cc_528 N_RESET_B_c_518_n N_A_1870_127#_c_1420_n 0.0456388f $X=10.23 $Y=1.965
+ $X2=0 $Y2=0
cc_529 N_RESET_B_c_537_n N_A_1870_127#_c_1420_n 0.0301065f $X=10.23 $Y=2.905
+ $X2=0 $Y2=0
cc_530 N_RESET_B_M1002_g N_A_1870_127#_c_1421_n 0.0184292f $X=11.055 $Y=0.845
+ $X2=0 $Y2=0
cc_531 N_RESET_B_c_518_n N_A_1870_127#_c_1421_n 0.0144144f $X=10.23 $Y=1.965
+ $X2=0 $Y2=0
cc_532 N_RESET_B_c_522_n N_A_1870_127#_c_1421_n 0.0077193f $X=10.875 $Y=1.46
+ $X2=0 $Y2=0
cc_533 N_RESET_B_c_523_n N_A_1870_127#_c_1421_n 0.0575072f $X=10.875 $Y=1.46
+ $X2=0 $Y2=0
cc_534 N_RESET_B_M1002_g N_A_1870_127#_c_1422_n 0.00165133f $X=11.055 $Y=0.845
+ $X2=0 $Y2=0
cc_535 N_RESET_B_c_523_n N_A_1870_127#_c_1422_n 0.00591683f $X=10.875 $Y=1.46
+ $X2=0 $Y2=0
cc_536 N_RESET_B_c_571_p N_A_1870_127#_c_1429_n 0.0190131f $X=10.145 $Y=2.99
+ $X2=0 $Y2=0
cc_537 N_RESET_B_c_537_n N_A_1870_127#_c_1429_n 0.0212058f $X=10.23 $Y=2.905
+ $X2=0 $Y2=0
cc_538 N_RESET_B_c_522_n N_A_1870_127#_c_1424_n 0.0312031f $X=10.875 $Y=1.46
+ $X2=0 $Y2=0
cc_539 N_RESET_B_c_523_n N_A_1870_127#_c_1424_n 3.6133e-19 $X=10.875 $Y=1.46
+ $X2=0 $Y2=0
cc_540 N_RESET_B_M1002_g N_A_1870_127#_c_1425_n 0.0312031f $X=11.055 $Y=0.845
+ $X2=0 $Y2=0
cc_541 N_RESET_B_c_540_n N_VPWR_M1000_d 0.00479327f $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_542 N_RESET_B_c_540_n N_VPWR_M1022_s 8.86199e-19 $X=7.775 $Y=2.035 $X2=0
+ $Y2=0
cc_543 N_RESET_B_c_534_n N_VPWR_M1038_s 0.00622929f $X=8.63 $Y=2.635 $X2=0 $Y2=0
cc_544 N_RESET_B_c_602_p N_VPWR_M1038_s 0.0076234f $X=9.095 $Y=2.72 $X2=0 $Y2=0
cc_545 N_RESET_B_c_535_n N_VPWR_M1038_s 0.00219111f $X=8.715 $Y=2.72 $X2=0 $Y2=0
cc_546 N_RESET_B_M1000_g N_VPWR_c_1600_n 0.00515877f $X=3.635 $Y=2.775 $X2=0
+ $Y2=0
cc_547 N_RESET_B_c_525_n N_VPWR_c_1602_n 0.00322432f $X=7.535 $Y=2.535 $X2=0
+ $Y2=0
cc_548 N_RESET_B_M1033_g N_VPWR_c_1603_n 0.00685991f $X=11.03 $Y=2.875 $X2=0
+ $Y2=0
cc_549 N_RESET_B_M1000_g N_VPWR_c_1608_n 0.00438531f $X=3.635 $Y=2.775 $X2=0
+ $Y2=0
cc_550 N_RESET_B_c_602_p N_VPWR_c_1610_n 0.0034313f $X=9.095 $Y=2.72 $X2=0 $Y2=0
cc_551 N_RESET_B_c_571_p N_VPWR_c_1610_n 0.0588f $X=10.145 $Y=2.99 $X2=0 $Y2=0
cc_552 N_RESET_B_c_572_p N_VPWR_c_1610_n 0.00946397f $X=9.18 $Y=2.72 $X2=0 $Y2=0
cc_553 N_RESET_B_M1033_g N_VPWR_c_1612_n 0.00539298f $X=11.03 $Y=2.875 $X2=0
+ $Y2=0
cc_554 N_RESET_B_c_525_n N_VPWR_c_1618_n 0.00555245f $X=7.535 $Y=2.535 $X2=0
+ $Y2=0
cc_555 N_RESET_B_c_535_n N_VPWR_c_1618_n 0.00103822f $X=8.715 $Y=2.72 $X2=0
+ $Y2=0
cc_556 N_RESET_B_M1000_g N_VPWR_c_1597_n 0.0067597f $X=3.635 $Y=2.775 $X2=0
+ $Y2=0
cc_557 N_RESET_B_c_525_n N_VPWR_c_1597_n 0.00699218f $X=7.535 $Y=2.535 $X2=0
+ $Y2=0
cc_558 N_RESET_B_M1033_g N_VPWR_c_1597_n 0.00662615f $X=11.03 $Y=2.875 $X2=0
+ $Y2=0
cc_559 N_RESET_B_c_531_n N_VPWR_c_1597_n 3.13815e-19 $X=7.83 $Y=2.46 $X2=0 $Y2=0
cc_560 N_RESET_B_c_602_p N_VPWR_c_1597_n 0.00633129f $X=9.095 $Y=2.72 $X2=0
+ $Y2=0
cc_561 N_RESET_B_c_535_n N_VPWR_c_1597_n 0.00220142f $X=8.715 $Y=2.72 $X2=0
+ $Y2=0
cc_562 N_RESET_B_c_571_p N_VPWR_c_1597_n 0.0383155f $X=10.145 $Y=2.99 $X2=0
+ $Y2=0
cc_563 N_RESET_B_c_572_p N_VPWR_c_1597_n 0.00618975f $X=9.18 $Y=2.72 $X2=0 $Y2=0
cc_564 N_RESET_B_c_602_p N_VPWR_c_1625_n 0.013809f $X=9.095 $Y=2.72 $X2=0 $Y2=0
cc_565 N_RESET_B_c_535_n N_VPWR_c_1625_n 0.00991451f $X=8.715 $Y=2.72 $X2=0
+ $Y2=0
cc_566 N_RESET_B_c_572_p N_VPWR_c_1625_n 0.00637247f $X=9.18 $Y=2.72 $X2=0 $Y2=0
cc_567 N_RESET_B_M1034_g N_A_229_491#_c_1770_n 0.0168434f $X=3.71 $Y=0.505 $X2=0
+ $Y2=0
cc_568 N_RESET_B_c_516_n N_A_229_491#_c_1770_n 0.00233077f $X=3.597 $Y=1.675
+ $X2=0 $Y2=0
cc_569 N_RESET_B_c_521_n N_A_229_491#_c_1770_n 0.0062518f $X=3.545 $Y=1.69 $X2=0
+ $Y2=0
cc_570 N_RESET_B_M1000_g N_A_229_491#_c_1775_n 0.0142313f $X=3.635 $Y=2.775
+ $X2=0 $Y2=0
cc_571 N_RESET_B_c_516_n N_A_229_491#_c_1775_n 0.00250809f $X=3.597 $Y=1.675
+ $X2=0 $Y2=0
cc_572 N_RESET_B_c_530_n N_A_229_491#_c_1775_n 2.49654e-19 $X=3.545 $Y=2.195
+ $X2=0 $Y2=0
cc_573 N_RESET_B_c_540_n N_A_229_491#_c_1775_n 0.00510689f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_574 N_RESET_B_c_541_n N_A_229_491#_c_1775_n 0.00338285f $X=3.745 $Y=2.035
+ $X2=0 $Y2=0
cc_575 N_RESET_B_c_521_n N_A_229_491#_c_1775_n 0.0122367f $X=3.545 $Y=1.69 $X2=0
+ $Y2=0
cc_576 N_RESET_B_M1034_g N_A_229_491#_c_1771_n 0.0108942f $X=3.71 $Y=0.505 $X2=0
+ $Y2=0
cc_577 N_RESET_B_c_516_n N_A_229_491#_c_1771_n 0.00133496f $X=3.597 $Y=1.675
+ $X2=0 $Y2=0
cc_578 N_RESET_B_c_540_n N_A_229_491#_c_1771_n 0.0233297f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_579 N_RESET_B_c_541_n N_A_229_491#_c_1771_n 0.00272324f $X=3.745 $Y=2.035
+ $X2=0 $Y2=0
cc_580 N_RESET_B_c_544_n N_A_229_491#_c_1771_n 0.0076359f $X=3.545 $Y=1.69 $X2=0
+ $Y2=0
cc_581 N_RESET_B_c_521_n N_A_229_491#_c_1771_n 0.0473063f $X=3.545 $Y=1.69 $X2=0
+ $Y2=0
cc_582 N_RESET_B_c_540_n N_A_229_491#_c_1777_n 0.0253812f $X=7.775 $Y=2.035
+ $X2=0 $Y2=0
cc_583 N_RESET_B_M1000_g N_A_229_491#_c_1780_n 7.66845e-19 $X=3.635 $Y=2.775
+ $X2=0 $Y2=0
cc_584 N_RESET_B_c_530_n N_A_229_491#_c_1780_n 0.00436676f $X=3.545 $Y=2.195
+ $X2=0 $Y2=0
cc_585 N_RESET_B_c_541_n N_A_229_491#_c_1780_n 7.71471e-19 $X=3.745 $Y=2.035
+ $X2=0 $Y2=0
cc_586 N_RESET_B_c_521_n N_A_229_491#_c_1780_n 0.00512399f $X=3.545 $Y=1.69
+ $X2=0 $Y2=0
cc_587 N_RESET_B_M1034_g N_A_229_491#_c_1826_n 0.00197753f $X=3.71 $Y=0.505
+ $X2=0 $Y2=0
cc_588 N_RESET_B_c_571_p A_2022_533# 9.38685e-19 $X=10.145 $Y=2.99 $X2=-0.19
+ $Y2=-0.245
cc_589 N_RESET_B_c_537_n A_2022_533# 3.24131e-19 $X=10.23 $Y=2.905 $X2=-0.19
+ $Y2=-0.245
cc_590 N_RESET_B_M1034_g N_VGND_c_1944_n 0.00505774f $X=3.71 $Y=0.505 $X2=0
+ $Y2=0
cc_591 N_RESET_B_M1009_g N_VGND_c_1946_n 0.00114139f $X=7.83 $Y=0.845 $X2=0
+ $Y2=0
cc_592 N_RESET_B_M1002_g N_VGND_c_1947_n 0.00651061f $X=11.055 $Y=0.845 $X2=0
+ $Y2=0
cc_593 N_RESET_B_M1034_g N_VGND_c_1949_n 0.00383942f $X=3.71 $Y=0.505 $X2=0
+ $Y2=0
cc_594 N_RESET_B_M1002_g N_VGND_c_1953_n 0.00410092f $X=11.055 $Y=0.845 $X2=0
+ $Y2=0
cc_595 N_RESET_B_M1034_g N_VGND_c_1955_n 0.00621997f $X=3.71 $Y=0.505 $X2=0
+ $Y2=0
cc_596 N_RESET_B_M1009_g N_VGND_c_1955_n 9.53055e-19 $X=7.83 $Y=0.845 $X2=0
+ $Y2=0
cc_597 N_RESET_B_M1002_g N_VGND_c_1955_n 0.00466677f $X=11.055 $Y=0.845 $X2=0
+ $Y2=0
cc_598 N_RESET_B_M1034_g N_noxref_24_c_2074_n 0.00382334f $X=3.71 $Y=0.505 $X2=0
+ $Y2=0
cc_599 N_CLK_N_c_752_n N_A_857_367#_M1022_g 7.95293e-19 $X=4.56 $Y=1.51 $X2=0
+ $Y2=0
cc_600 N_CLK_N_c_752_n N_A_857_367#_c_1190_n 0.00968186f $X=4.56 $Y=1.51 $X2=0
+ $Y2=0
cc_601 N_CLK_N_c_753_n N_A_857_367#_c_1190_n 0.0122831f $X=4.56 $Y=1.51 $X2=0
+ $Y2=0
cc_602 N_CLK_N_M1023_g N_A_857_367#_c_1182_n 0.00426097f $X=4.335 $Y=0.765 $X2=0
+ $Y2=0
cc_603 N_CLK_N_c_752_n N_A_857_367#_c_1182_n 0.0057283f $X=4.56 $Y=1.51 $X2=0
+ $Y2=0
cc_604 N_CLK_N_c_753_n N_A_857_367#_c_1182_n 0.0122617f $X=4.56 $Y=1.51 $X2=0
+ $Y2=0
cc_605 N_CLK_N_M1023_g N_A_857_367#_c_1183_n 0.00275731f $X=4.335 $Y=0.765 $X2=0
+ $Y2=0
cc_606 N_CLK_N_c_752_n N_A_857_367#_c_1183_n 0.00153445f $X=4.56 $Y=1.51 $X2=0
+ $Y2=0
cc_607 N_CLK_N_c_753_n N_A_857_367#_c_1183_n 0.0145412f $X=4.56 $Y=1.51 $X2=0
+ $Y2=0
cc_608 N_CLK_N_M1023_g N_A_857_367#_c_1184_n 0.00122777f $X=4.335 $Y=0.765 $X2=0
+ $Y2=0
cc_609 N_CLK_N_c_752_n N_A_857_367#_c_1184_n 0.0163378f $X=4.56 $Y=1.51 $X2=0
+ $Y2=0
cc_610 N_CLK_N_c_753_n N_A_857_367#_c_1184_n 0.00105358f $X=4.56 $Y=1.51 $X2=0
+ $Y2=0
cc_611 N_CLK_N_M1035_g N_VPWR_c_1600_n 0.00510775f $X=4.21 $Y=2.465 $X2=0 $Y2=0
cc_612 N_CLK_N_M1035_g N_VPWR_c_1601_n 0.008718f $X=4.21 $Y=2.465 $X2=0 $Y2=0
cc_613 N_CLK_N_M1035_g N_VPWR_c_1616_n 0.00438531f $X=4.21 $Y=2.465 $X2=0 $Y2=0
cc_614 N_CLK_N_M1035_g N_VPWR_c_1597_n 0.00788496f $X=4.21 $Y=2.465 $X2=0 $Y2=0
cc_615 N_CLK_N_M1023_g N_A_229_491#_c_1771_n 0.0078265f $X=4.335 $Y=0.765 $X2=0
+ $Y2=0
cc_616 N_CLK_N_c_752_n N_A_229_491#_c_1771_n 0.0146218f $X=4.56 $Y=1.51 $X2=0
+ $Y2=0
cc_617 N_CLK_N_c_753_n N_A_229_491#_c_1771_n 0.0144884f $X=4.56 $Y=1.51 $X2=0
+ $Y2=0
cc_618 N_CLK_N_M1023_g N_A_229_491#_c_1772_n 0.0182872f $X=4.335 $Y=0.765 $X2=0
+ $Y2=0
cc_619 N_CLK_N_c_752_n N_A_229_491#_c_1772_n 0.00282525f $X=4.56 $Y=1.51 $X2=0
+ $Y2=0
cc_620 N_CLK_N_M1035_g N_A_229_491#_c_1777_n 0.0156777f $X=4.21 $Y=2.465 $X2=0
+ $Y2=0
cc_621 N_CLK_N_M1023_g N_A_229_491#_c_1826_n 0.00165394f $X=4.335 $Y=0.765 $X2=0
+ $Y2=0
cc_622 N_CLK_N_M1035_g N_A_229_491#_c_1834_n 0.00192845f $X=4.21 $Y=2.465 $X2=0
+ $Y2=0
cc_623 N_CLK_N_M1023_g N_VGND_c_1944_n 0.00436282f $X=4.335 $Y=0.765 $X2=0 $Y2=0
cc_624 N_CLK_N_M1023_g N_VGND_c_1945_n 0.00576575f $X=4.335 $Y=0.765 $X2=0 $Y2=0
cc_625 N_CLK_N_M1023_g N_VGND_c_1950_n 0.00341315f $X=4.335 $Y=0.765 $X2=0 $Y2=0
cc_626 N_CLK_N_M1023_g N_VGND_c_1955_n 0.00490366f $X=4.335 $Y=0.765 $X2=0 $Y2=0
cc_627 N_A_1080_47#_c_820_n N_A_1406_399#_M1001_d 0.0127541f $X=9.195 $Y=0.805
+ $X2=-0.19 $Y2=-0.245
cc_628 N_A_1080_47#_M1027_g N_A_1406_399#_M1036_g 0.0367956f $X=6.745 $Y=2.855
+ $X2=0 $Y2=0
cc_629 N_A_1080_47#_c_797_n N_A_1406_399#_M1007_g 0.00314207f $X=7.265 $Y=0.72
+ $X2=0 $Y2=0
cc_630 N_A_1080_47#_c_820_n N_A_1406_399#_M1007_g 0.0101654f $X=9.195 $Y=0.805
+ $X2=0 $Y2=0
cc_631 N_A_1080_47#_c_815_n N_A_1406_399#_c_968_n 3.1098e-19 $X=6.745 $Y=1.98
+ $X2=0 $Y2=0
cc_632 N_A_1080_47#_c_815_n N_A_1406_399#_c_975_n 0.046073f $X=6.745 $Y=1.98
+ $X2=0 $Y2=0
cc_633 N_A_1080_47#_c_820_n N_A_1406_399#_c_969_n 0.0870516f $X=9.195 $Y=0.805
+ $X2=0 $Y2=0
cc_634 N_A_1080_47#_c_820_n N_A_1406_399#_c_970_n 0.0135257f $X=9.195 $Y=0.805
+ $X2=0 $Y2=0
cc_635 N_A_1080_47#_c_831_p N_A_1406_399#_c_970_n 0.0106086f $X=7.35 $Y=0.805
+ $X2=0 $Y2=0
cc_636 N_A_1080_47#_c_820_n N_A_1406_399#_c_1014_n 0.013831f $X=9.195 $Y=0.805
+ $X2=0 $Y2=0
cc_637 N_A_1080_47#_c_799_n N_A_1406_399#_c_1014_n 0.015786f $X=9.365 $Y=1.755
+ $X2=0 $Y2=0
cc_638 N_A_1080_47#_M1006_g N_A_1406_399#_c_971_n 9.76774e-19 $X=9.51 $Y=2.665
+ $X2=0 $Y2=0
cc_639 N_A_1080_47#_c_799_n N_A_1406_399#_c_971_n 0.0361056f $X=9.365 $Y=1.755
+ $X2=0 $Y2=0
cc_640 N_A_1080_47#_c_813_n N_A_1406_399#_c_971_n 0.0258427f $X=9.53 $Y=1.92
+ $X2=0 $Y2=0
cc_641 N_A_1080_47#_c_814_n N_A_1406_399#_c_971_n 8.56979e-19 $X=9.53 $Y=1.92
+ $X2=0 $Y2=0
cc_642 N_A_1080_47#_M1006_g N_A_1406_399#_c_1003_n 0.00345894f $X=9.51 $Y=2.665
+ $X2=0 $Y2=0
cc_643 N_A_1080_47#_c_813_n N_A_1406_399#_c_1003_n 0.0110559f $X=9.53 $Y=1.92
+ $X2=0 $Y2=0
cc_644 N_A_1080_47#_c_814_n N_A_1406_399#_c_1003_n 0.00143126f $X=9.53 $Y=1.92
+ $X2=0 $Y2=0
cc_645 N_A_1080_47#_c_820_n N_A_1278_529#_M1001_g 0.0134774f $X=9.195 $Y=0.805
+ $X2=0 $Y2=0
cc_646 N_A_1080_47#_c_798_n N_A_1278_529#_M1001_g 0.0023956f $X=9.322 $Y=0.72
+ $X2=0 $Y2=0
cc_647 N_A_1080_47#_c_799_n N_A_1278_529#_M1001_g 9.66683e-19 $X=9.365 $Y=1.755
+ $X2=0 $Y2=0
cc_648 N_A_1080_47#_c_814_n N_A_1278_529#_M1001_g 0.00242397f $X=9.53 $Y=1.92
+ $X2=0 $Y2=0
cc_649 N_A_1080_47#_M1006_g N_A_1278_529#_c_1058_n 0.0357702f $X=9.51 $Y=2.665
+ $X2=0 $Y2=0
cc_650 N_A_1080_47#_c_813_n N_A_1278_529#_c_1058_n 6.78682e-19 $X=9.53 $Y=1.92
+ $X2=0 $Y2=0
cc_651 N_A_1080_47#_c_814_n N_A_1278_529#_c_1058_n 0.00659447f $X=9.53 $Y=1.92
+ $X2=0 $Y2=0
cc_652 N_A_1080_47#_M1027_g N_A_1278_529#_c_1061_n 0.00985362f $X=6.745 $Y=2.855
+ $X2=0 $Y2=0
cc_653 N_A_1080_47#_M1027_g N_A_1278_529#_c_1056_n 0.00512219f $X=6.745 $Y=2.855
+ $X2=0 $Y2=0
cc_654 N_A_1080_47#_c_793_n N_A_1278_529#_c_1056_n 0.0142454f $X=6.46 $Y=1.21
+ $X2=0 $Y2=0
cc_655 N_A_1080_47#_c_810_n N_A_1278_529#_c_1056_n 0.0240557f $X=6.545 $Y=1.98
+ $X2=0 $Y2=0
cc_656 N_A_1080_47#_c_795_n N_A_1278_529#_c_1056_n 0.0177082f $X=6.545 $Y=1.125
+ $X2=0 $Y2=0
cc_657 N_A_1080_47#_c_796_n N_A_1278_529#_c_1056_n 0.014755f $X=7.18 $Y=0.382
+ $X2=0 $Y2=0
cc_658 N_A_1080_47#_c_812_n N_A_1278_529#_c_1056_n 0.00326632f $X=6.16 $Y=2.037
+ $X2=0 $Y2=0
cc_659 N_A_1080_47#_c_815_n N_A_1278_529#_c_1056_n 0.00664756f $X=6.745 $Y=1.98
+ $X2=0 $Y2=0
cc_660 N_A_1080_47#_c_805_n N_A_1278_529#_c_1056_n 0.00100223f $X=6.625 $Y=0.525
+ $X2=0 $Y2=0
cc_661 N_A_1080_47#_M1027_g N_A_1278_529#_c_1065_n 0.0122403f $X=6.745 $Y=2.855
+ $X2=0 $Y2=0
cc_662 N_A_1080_47#_c_810_n N_A_1278_529#_c_1065_n 0.0165782f $X=6.545 $Y=1.98
+ $X2=0 $Y2=0
cc_663 N_A_1080_47#_c_815_n N_A_1278_529#_c_1065_n 0.00310507f $X=6.745 $Y=1.98
+ $X2=0 $Y2=0
cc_664 N_A_1080_47#_c_793_n N_A_857_367#_M1019_g 4.54798e-19 $X=6.46 $Y=1.21
+ $X2=0 $Y2=0
cc_665 N_A_1080_47#_c_803_n N_A_857_367#_M1019_g 0.0103032f $X=5.655 $Y=1.06
+ $X2=0 $Y2=0
cc_666 N_A_1080_47#_c_792_n N_A_857_367#_M1022_g 0.00507988f $X=5.607 $Y=1.815
+ $X2=0 $Y2=0
cc_667 N_A_1080_47#_c_812_n N_A_857_367#_M1022_g 0.00537011f $X=6.16 $Y=2.037
+ $X2=0 $Y2=0
cc_668 N_A_1080_47#_c_792_n N_A_857_367#_c_1171_n 0.0268583f $X=5.607 $Y=1.815
+ $X2=0 $Y2=0
cc_669 N_A_1080_47#_c_793_n N_A_857_367#_c_1171_n 0.0170957f $X=6.46 $Y=1.21
+ $X2=0 $Y2=0
cc_670 N_A_1080_47#_c_812_n N_A_857_367#_c_1171_n 0.00312898f $X=6.16 $Y=2.037
+ $X2=0 $Y2=0
cc_671 N_A_1080_47#_M1027_g N_A_857_367#_c_1172_n 0.00284238f $X=6.745 $Y=2.855
+ $X2=0 $Y2=0
cc_672 N_A_1080_47#_c_792_n N_A_857_367#_c_1172_n 0.00687673f $X=5.607 $Y=1.815
+ $X2=0 $Y2=0
cc_673 N_A_1080_47#_c_812_n N_A_857_367#_c_1172_n 0.0247093f $X=6.16 $Y=2.037
+ $X2=0 $Y2=0
cc_674 N_A_1080_47#_c_815_n N_A_857_367#_c_1172_n 0.0181136f $X=6.745 $Y=1.98
+ $X2=0 $Y2=0
cc_675 N_A_1080_47#_c_793_n N_A_857_367#_c_1173_n 0.00413257f $X=6.46 $Y=1.21
+ $X2=0 $Y2=0
cc_676 N_A_1080_47#_c_810_n N_A_857_367#_c_1173_n 9.48461e-19 $X=6.545 $Y=1.98
+ $X2=0 $Y2=0
cc_677 N_A_1080_47#_c_812_n N_A_857_367#_c_1173_n 0.00518753f $X=6.16 $Y=2.037
+ $X2=0 $Y2=0
cc_678 N_A_1080_47#_c_815_n N_A_857_367#_c_1173_n 0.0249314f $X=6.745 $Y=1.98
+ $X2=0 $Y2=0
cc_679 N_A_1080_47#_c_805_n N_A_857_367#_c_1173_n 0.00952309f $X=6.625 $Y=0.525
+ $X2=0 $Y2=0
cc_680 N_A_1080_47#_c_795_n N_A_857_367#_M1008_g 5.64478e-19 $X=6.545 $Y=1.125
+ $X2=0 $Y2=0
cc_681 N_A_1080_47#_c_796_n N_A_857_367#_M1008_g 0.0185221f $X=7.18 $Y=0.382
+ $X2=0 $Y2=0
cc_682 N_A_1080_47#_c_797_n N_A_857_367#_M1008_g 0.00438564f $X=7.265 $Y=0.72
+ $X2=0 $Y2=0
cc_683 N_A_1080_47#_c_831_p N_A_857_367#_M1008_g 0.00332654f $X=7.35 $Y=0.805
+ $X2=0 $Y2=0
cc_684 N_A_1080_47#_c_805_n N_A_857_367#_M1008_g 0.0101149f $X=6.625 $Y=0.525
+ $X2=0 $Y2=0
cc_685 N_A_1080_47#_c_796_n N_A_857_367#_c_1175_n 0.00316552f $X=7.18 $Y=0.382
+ $X2=0 $Y2=0
cc_686 N_A_1080_47#_c_820_n N_A_857_367#_c_1175_n 0.0166672f $X=9.195 $Y=0.805
+ $X2=0 $Y2=0
cc_687 N_A_1080_47#_c_800_n N_A_857_367#_c_1175_n 0.00128489f $X=9.45 $Y=0.355
+ $X2=0 $Y2=0
cc_688 N_A_1080_47#_c_802_n N_A_857_367#_c_1175_n 0.00867237f $X=9.945 $Y=0.36
+ $X2=0 $Y2=0
cc_689 N_A_1080_47#_c_804_n N_A_857_367#_c_1176_n 0.0180755f $X=6.625 $Y=0.36
+ $X2=0 $Y2=0
cc_690 N_A_1080_47#_c_798_n N_A_857_367#_M1016_g 0.00885388f $X=9.322 $Y=0.72
+ $X2=0 $Y2=0
cc_691 N_A_1080_47#_c_799_n N_A_857_367#_M1016_g 0.015339f $X=9.365 $Y=1.755
+ $X2=0 $Y2=0
cc_692 N_A_1080_47#_c_800_n N_A_857_367#_M1016_g 0.00876101f $X=9.45 $Y=0.355
+ $X2=0 $Y2=0
cc_693 N_A_1080_47#_c_889_p N_A_857_367#_M1016_g 0.0113795f $X=9.322 $Y=0.805
+ $X2=0 $Y2=0
cc_694 N_A_1080_47#_c_806_n N_A_857_367#_M1016_g 0.00867589f $X=9.945 $Y=0.525
+ $X2=0 $Y2=0
cc_695 N_A_1080_47#_c_799_n N_A_857_367#_c_1178_n 0.00777861f $X=9.365 $Y=1.755
+ $X2=0 $Y2=0
cc_696 N_A_1080_47#_c_813_n N_A_857_367#_c_1178_n 0.00121249f $X=9.53 $Y=1.92
+ $X2=0 $Y2=0
cc_697 N_A_1080_47#_c_814_n N_A_857_367#_c_1178_n 0.0219808f $X=9.53 $Y=1.92
+ $X2=0 $Y2=0
cc_698 N_A_1080_47#_c_806_n N_A_857_367#_c_1178_n 0.0100252f $X=9.945 $Y=0.525
+ $X2=0 $Y2=0
cc_699 N_A_1080_47#_c_799_n N_A_857_367#_c_1179_n 0.00331033f $X=9.365 $Y=1.755
+ $X2=0 $Y2=0
cc_700 N_A_1080_47#_c_813_n N_A_857_367#_c_1179_n 3.52582e-19 $X=9.53 $Y=1.92
+ $X2=0 $Y2=0
cc_701 N_A_1080_47#_M1006_g N_A_857_367#_M1024_g 0.0283888f $X=9.51 $Y=2.665
+ $X2=0 $Y2=0
cc_702 N_A_1080_47#_c_799_n N_A_857_367#_M1024_g 9.49777e-19 $X=9.365 $Y=1.755
+ $X2=0 $Y2=0
cc_703 N_A_1080_47#_c_813_n N_A_857_367#_M1024_g 2.8557e-19 $X=9.53 $Y=1.92
+ $X2=0 $Y2=0
cc_704 N_A_1080_47#_c_814_n N_A_857_367#_M1024_g 0.0150528f $X=9.53 $Y=1.92
+ $X2=0 $Y2=0
cc_705 N_A_1080_47#_M1027_g N_A_857_367#_c_1189_n 0.0187017f $X=6.745 $Y=2.855
+ $X2=0 $Y2=0
cc_706 N_A_1080_47#_c_810_n N_A_857_367#_c_1189_n 0.00764441f $X=6.545 $Y=1.98
+ $X2=0 $Y2=0
cc_707 N_A_1080_47#_c_812_n N_A_857_367#_c_1189_n 4.14458e-19 $X=6.16 $Y=2.037
+ $X2=0 $Y2=0
cc_708 N_A_1080_47#_c_815_n N_A_857_367#_c_1189_n 5.65657e-19 $X=6.745 $Y=1.98
+ $X2=0 $Y2=0
cc_709 N_A_1080_47#_c_812_n N_A_857_367#_c_1190_n 0.0144661f $X=6.16 $Y=2.037
+ $X2=0 $Y2=0
cc_710 N_A_1080_47#_c_803_n N_A_857_367#_c_1182_n 0.0114684f $X=5.655 $Y=1.06
+ $X2=0 $Y2=0
cc_711 N_A_1080_47#_c_803_n N_A_857_367#_c_1183_n 0.046314f $X=5.655 $Y=1.06
+ $X2=0 $Y2=0
cc_712 N_A_1080_47#_c_812_n N_A_857_367#_c_1183_n 0.00523873f $X=6.16 $Y=2.037
+ $X2=0 $Y2=0
cc_713 N_A_1080_47#_c_792_n N_A_857_367#_c_1184_n 0.00851225f $X=5.607 $Y=1.815
+ $X2=0 $Y2=0
cc_714 N_A_1080_47#_c_802_n N_A_2064_101#_M1029_g 0.0416165f $X=9.945 $Y=0.36
+ $X2=0 $Y2=0
cc_715 N_A_1080_47#_c_798_n N_A_1870_127#_M1016_d 8.08045e-19 $X=9.322 $Y=0.72
+ $X2=-0.19 $Y2=-0.245
cc_716 N_A_1080_47#_c_799_n N_A_1870_127#_M1016_d 0.00374629f $X=9.365 $Y=1.755
+ $X2=-0.19 $Y2=-0.245
cc_717 N_A_1080_47#_c_889_p N_A_1870_127#_M1016_d 0.00168104f $X=9.322 $Y=0.805
+ $X2=-0.19 $Y2=-0.245
cc_718 N_A_1080_47#_c_798_n N_A_1870_127#_c_1419_n 0.00749264f $X=9.322 $Y=0.72
+ $X2=0 $Y2=0
cc_719 N_A_1080_47#_c_799_n N_A_1870_127#_c_1419_n 0.0102762f $X=9.365 $Y=1.755
+ $X2=0 $Y2=0
cc_720 N_A_1080_47#_c_801_n N_A_1870_127#_c_1419_n 0.0268527f $X=9.945 $Y=0.36
+ $X2=0 $Y2=0
cc_721 N_A_1080_47#_c_802_n N_A_1870_127#_c_1419_n 0.00456429f $X=9.945 $Y=0.36
+ $X2=0 $Y2=0
cc_722 N_A_1080_47#_c_889_p N_A_1870_127#_c_1419_n 0.0145233f $X=9.322 $Y=0.805
+ $X2=0 $Y2=0
cc_723 N_A_1080_47#_c_806_n N_A_1870_127#_c_1419_n 0.0131553f $X=9.945 $Y=0.525
+ $X2=0 $Y2=0
cc_724 N_A_1080_47#_M1006_g N_A_1870_127#_c_1420_n 0.00468037f $X=9.51 $Y=2.665
+ $X2=0 $Y2=0
cc_725 N_A_1080_47#_c_799_n N_A_1870_127#_c_1420_n 0.0200476f $X=9.365 $Y=1.755
+ $X2=0 $Y2=0
cc_726 N_A_1080_47#_c_813_n N_A_1870_127#_c_1420_n 0.0248547f $X=9.53 $Y=1.92
+ $X2=0 $Y2=0
cc_727 N_A_1080_47#_c_814_n N_A_1870_127#_c_1420_n 0.00230619f $X=9.53 $Y=1.92
+ $X2=0 $Y2=0
cc_728 N_A_1080_47#_c_801_n N_A_1870_127#_c_1421_n 0.00367878f $X=9.945 $Y=0.36
+ $X2=0 $Y2=0
cc_729 N_A_1080_47#_c_806_n N_A_1870_127#_c_1421_n 0.00766943f $X=9.945 $Y=0.525
+ $X2=0 $Y2=0
cc_730 N_A_1080_47#_c_799_n N_A_1870_127#_c_1423_n 0.0216372f $X=9.365 $Y=1.755
+ $X2=0 $Y2=0
cc_731 N_A_1080_47#_c_806_n N_A_1870_127#_c_1423_n 0.00276914f $X=9.945 $Y=0.525
+ $X2=0 $Y2=0
cc_732 N_A_1080_47#_c_814_n N_A_1870_127#_c_1429_n 0.00203264f $X=9.53 $Y=1.92
+ $X2=0 $Y2=0
cc_733 N_A_1080_47#_M1027_g N_VPWR_c_1602_n 0.00214711f $X=6.745 $Y=2.855 $X2=0
+ $Y2=0
cc_734 N_A_1080_47#_M1006_g N_VPWR_c_1610_n 0.00351226f $X=9.51 $Y=2.665 $X2=0
+ $Y2=0
cc_735 N_A_1080_47#_M1027_g N_VPWR_c_1617_n 0.00522167f $X=6.745 $Y=2.855 $X2=0
+ $Y2=0
cc_736 N_A_1080_47#_M1022_d N_VPWR_c_1597_n 0.00348066f $X=5.4 $Y=1.835 $X2=0
+ $Y2=0
cc_737 N_A_1080_47#_M1027_g N_VPWR_c_1597_n 0.00585499f $X=6.745 $Y=2.855 $X2=0
+ $Y2=0
cc_738 N_A_1080_47#_M1006_g N_VPWR_c_1597_n 0.00557466f $X=9.51 $Y=2.665 $X2=0
+ $Y2=0
cc_739 N_A_1080_47#_c_795_n N_A_229_491#_M1020_s 0.00554459f $X=6.545 $Y=1.125
+ $X2=0 $Y2=0
cc_740 N_A_1080_47#_M1019_d N_A_229_491#_c_1772_n 0.0113352f $X=5.4 $Y=0.235
+ $X2=0 $Y2=0
cc_741 N_A_1080_47#_c_793_n N_A_229_491#_c_1772_n 0.0104678f $X=6.46 $Y=1.21
+ $X2=0 $Y2=0
cc_742 N_A_1080_47#_c_803_n N_A_229_491#_c_1772_n 0.0298154f $X=5.655 $Y=1.06
+ $X2=0 $Y2=0
cc_743 N_A_1080_47#_M1022_d N_A_229_491#_c_1777_n 0.00689834f $X=5.4 $Y=1.835
+ $X2=0 $Y2=0
cc_744 N_A_1080_47#_c_810_n N_A_229_491#_c_1777_n 0.0036704f $X=6.545 $Y=1.98
+ $X2=0 $Y2=0
cc_745 N_A_1080_47#_c_812_n N_A_229_491#_c_1777_n 0.0538404f $X=6.16 $Y=2.037
+ $X2=0 $Y2=0
cc_746 N_A_1080_47#_c_793_n N_A_229_491#_c_1774_n 0.0194195f $X=6.46 $Y=1.21
+ $X2=0 $Y2=0
cc_747 N_A_1080_47#_c_795_n N_A_229_491#_c_1774_n 0.0247093f $X=6.545 $Y=1.125
+ $X2=0 $Y2=0
cc_748 N_A_1080_47#_c_805_n N_A_229_491#_c_1774_n 0.00170198f $X=6.625 $Y=0.525
+ $X2=0 $Y2=0
cc_749 N_A_1080_47#_c_820_n N_VGND_M1009_d 0.0138302f $X=9.195 $Y=0.805 $X2=0
+ $Y2=0
cc_750 N_A_1080_47#_c_820_n N_VGND_c_1946_n 0.0256906f $X=9.195 $Y=0.805 $X2=0
+ $Y2=0
cc_751 N_A_1080_47#_c_801_n N_VGND_c_1947_n 0.00798947f $X=9.945 $Y=0.36 $X2=0
+ $Y2=0
cc_752 N_A_1080_47#_c_802_n N_VGND_c_1947_n 0.00452829f $X=9.945 $Y=0.36 $X2=0
+ $Y2=0
cc_753 N_A_1080_47#_c_794_n N_VGND_c_1951_n 0.0115893f $X=6.545 $Y=0.51 $X2=0
+ $Y2=0
cc_754 N_A_1080_47#_c_796_n N_VGND_c_1951_n 0.0469535f $X=7.18 $Y=0.382 $X2=0
+ $Y2=0
cc_755 N_A_1080_47#_c_820_n N_VGND_c_1951_n 0.00944413f $X=9.195 $Y=0.805 $X2=0
+ $Y2=0
cc_756 N_A_1080_47#_c_804_n N_VGND_c_1951_n 0.00635465f $X=6.625 $Y=0.36 $X2=0
+ $Y2=0
cc_757 N_A_1080_47#_c_820_n N_VGND_c_1952_n 0.00957881f $X=9.195 $Y=0.805 $X2=0
+ $Y2=0
cc_758 N_A_1080_47#_c_800_n N_VGND_c_1952_n 0.0176742f $X=9.45 $Y=0.355 $X2=0
+ $Y2=0
cc_759 N_A_1080_47#_c_801_n N_VGND_c_1952_n 0.0419853f $X=9.945 $Y=0.36 $X2=0
+ $Y2=0
cc_760 N_A_1080_47#_c_802_n N_VGND_c_1952_n 0.00635651f $X=9.945 $Y=0.36 $X2=0
+ $Y2=0
cc_761 N_A_1080_47#_M1019_d N_VGND_c_1955_n 0.00466812f $X=5.4 $Y=0.235 $X2=0
+ $Y2=0
cc_762 N_A_1080_47#_c_794_n N_VGND_c_1955_n 0.00583135f $X=6.545 $Y=0.51 $X2=0
+ $Y2=0
cc_763 N_A_1080_47#_c_796_n N_VGND_c_1955_n 0.0252492f $X=7.18 $Y=0.382 $X2=0
+ $Y2=0
cc_764 N_A_1080_47#_c_820_n N_VGND_c_1955_n 0.0354711f $X=9.195 $Y=0.805 $X2=0
+ $Y2=0
cc_765 N_A_1080_47#_c_800_n N_VGND_c_1955_n 0.00916446f $X=9.45 $Y=0.355 $X2=0
+ $Y2=0
cc_766 N_A_1080_47#_c_801_n N_VGND_c_1955_n 0.0233936f $X=9.945 $Y=0.36 $X2=0
+ $Y2=0
cc_767 N_A_1080_47#_c_802_n N_VGND_c_1955_n 0.00923403f $X=9.945 $Y=0.36 $X2=0
+ $Y2=0
cc_768 N_A_1080_47#_c_804_n N_VGND_c_1955_n 0.00911223f $X=6.625 $Y=0.36 $X2=0
+ $Y2=0
cc_769 N_A_1080_47#_c_831_p A_1437_127# 0.00106014f $X=7.35 $Y=0.805 $X2=-0.19
+ $Y2=-0.245
cc_770 N_A_1080_47#_c_820_n A_1509_127# 0.00251139f $X=9.195 $Y=0.805 $X2=-0.19
+ $Y2=-0.245
cc_771 N_A_1406_399#_c_969_n N_A_1278_529#_M1001_g 0.0140796f $X=8.94 $Y=1.16
+ $X2=0 $Y2=0
cc_772 N_A_1406_399#_c_971_n N_A_1278_529#_M1001_g 0.00617486f $X=9.025 $Y=2.265
+ $X2=0 $Y2=0
cc_773 N_A_1406_399#_c_971_n N_A_1278_529#_c_1058_n 0.0101668f $X=9.025 $Y=2.265
+ $X2=0 $Y2=0
cc_774 N_A_1406_399#_c_971_n N_A_1278_529#_c_1060_n 0.00426677f $X=9.025
+ $Y=2.265 $X2=0 $Y2=0
cc_775 N_A_1406_399#_c_1000_n N_A_1278_529#_c_1060_n 0.00547219f $X=9.11
+ $Y=2.365 $X2=0 $Y2=0
cc_776 N_A_1406_399#_c_1003_n N_A_1278_529#_c_1060_n 0.00313828f $X=9.295
+ $Y=2.37 $X2=0 $Y2=0
cc_777 N_A_1406_399#_M1036_g N_A_1278_529#_c_1061_n 0.00175351f $X=7.105
+ $Y=2.855 $X2=0 $Y2=0
cc_778 N_A_1406_399#_M1007_g N_A_1278_529#_c_1056_n 0.00122807f $X=7.47 $Y=0.845
+ $X2=0 $Y2=0
cc_779 N_A_1406_399#_c_968_n N_A_1278_529#_c_1056_n 0.0567084f $X=7.38 $Y=1.98
+ $X2=0 $Y2=0
cc_780 N_A_1406_399#_c_975_n N_A_1278_529#_c_1056_n 0.00676876f $X=7.38 $Y=1.98
+ $X2=0 $Y2=0
cc_781 N_A_1406_399#_c_970_n N_A_1278_529#_c_1056_n 0.0144602f $X=7.545 $Y=1.16
+ $X2=0 $Y2=0
cc_782 N_A_1406_399#_M1036_g N_A_1278_529#_c_1065_n 8.82443e-19 $X=7.105
+ $Y=2.855 $X2=0 $Y2=0
cc_783 N_A_1406_399#_M1036_g N_A_1278_529#_c_1066_n 0.0116602f $X=7.105 $Y=2.855
+ $X2=0 $Y2=0
cc_784 N_A_1406_399#_c_968_n N_A_1278_529#_c_1066_n 0.0203998f $X=7.38 $Y=1.98
+ $X2=0 $Y2=0
cc_785 N_A_1406_399#_c_975_n N_A_1278_529#_c_1066_n 0.0032127f $X=7.38 $Y=1.98
+ $X2=0 $Y2=0
cc_786 N_A_1406_399#_c_975_n N_A_857_367#_c_1173_n 0.00965412f $X=7.38 $Y=1.98
+ $X2=0 $Y2=0
cc_787 N_A_1406_399#_M1007_g N_A_857_367#_M1008_g 0.0649028f $X=7.47 $Y=0.845
+ $X2=0 $Y2=0
cc_788 N_A_1406_399#_c_968_n N_A_857_367#_M1008_g 0.00262389f $X=7.38 $Y=1.98
+ $X2=0 $Y2=0
cc_789 N_A_1406_399#_c_970_n N_A_857_367#_M1008_g 0.00169562f $X=7.545 $Y=1.16
+ $X2=0 $Y2=0
cc_790 N_A_1406_399#_M1007_g N_A_857_367#_c_1175_n 0.00807149f $X=7.47 $Y=0.845
+ $X2=0 $Y2=0
cc_791 N_A_1406_399#_c_1014_n N_A_857_367#_M1016_g 0.00202048f $X=9.025 $Y=1.26
+ $X2=0 $Y2=0
cc_792 N_A_1406_399#_c_971_n N_A_857_367#_M1016_g 0.0029999f $X=9.025 $Y=2.265
+ $X2=0 $Y2=0
cc_793 N_A_1406_399#_c_1003_n N_A_1870_127#_c_1420_n 0.0063281f $X=9.295 $Y=2.37
+ $X2=0 $Y2=0
cc_794 N_A_1406_399#_c_971_n N_VPWR_M1038_s 2.01365e-19 $X=9.025 $Y=2.265 $X2=0
+ $Y2=0
cc_795 N_A_1406_399#_c_1000_n N_VPWR_M1038_s 0.00223439f $X=9.11 $Y=2.365 $X2=0
+ $Y2=0
cc_796 N_A_1406_399#_M1036_g N_VPWR_c_1602_n 0.010968f $X=7.105 $Y=2.855 $X2=0
+ $Y2=0
cc_797 N_A_1406_399#_M1036_g N_VPWR_c_1617_n 0.00461019f $X=7.105 $Y=2.855 $X2=0
+ $Y2=0
cc_798 N_A_1406_399#_M1038_d N_VPWR_c_1597_n 0.00224374f $X=9.155 $Y=2.245 $X2=0
+ $Y2=0
cc_799 N_A_1406_399#_M1036_g N_VPWR_c_1597_n 0.00427129f $X=7.105 $Y=2.855 $X2=0
+ $Y2=0
cc_800 N_A_1406_399#_c_1000_n N_VPWR_c_1597_n 2.91638e-19 $X=9.11 $Y=2.365 $X2=0
+ $Y2=0
cc_801 N_A_1406_399#_c_969_n N_VGND_M1009_d 0.00960504f $X=8.94 $Y=1.16 $X2=0
+ $Y2=0
cc_802 N_A_1406_399#_M1007_g N_VGND_c_1955_n 9.53055e-19 $X=7.47 $Y=0.845 $X2=0
+ $Y2=0
cc_803 N_A_1278_529#_c_1056_n N_A_857_367#_c_1172_n 0.0035665f $X=6.895 $Y=0.845
+ $X2=0 $Y2=0
cc_804 N_A_1278_529#_c_1056_n N_A_857_367#_c_1173_n 0.0191296f $X=6.895 $Y=0.845
+ $X2=0 $Y2=0
cc_805 N_A_1278_529#_c_1056_n N_A_857_367#_M1008_g 0.00675573f $X=6.895 $Y=0.845
+ $X2=0 $Y2=0
cc_806 N_A_1278_529#_M1001_g N_A_857_367#_c_1175_n 0.00807149f $X=8.615 $Y=0.955
+ $X2=0 $Y2=0
cc_807 N_A_1278_529#_M1001_g N_A_857_367#_M1016_g 0.0191827f $X=8.615 $Y=0.955
+ $X2=0 $Y2=0
cc_808 N_A_1278_529#_c_1061_n N_A_857_367#_c_1189_n 0.00107635f $X=6.53 $Y=2.855
+ $X2=0 $Y2=0
cc_809 N_A_1278_529#_c_1065_n N_A_857_367#_c_1189_n 0.0024308f $X=7 $Y=2.42
+ $X2=0 $Y2=0
cc_810 N_A_1278_529#_c_1061_n N_VPWR_c_1602_n 0.0108528f $X=6.53 $Y=2.855 $X2=0
+ $Y2=0
cc_811 N_A_1278_529#_c_1066_n N_VPWR_c_1602_n 0.0185547f $X=7.625 $Y=2.685 $X2=0
+ $Y2=0
cc_812 N_A_1278_529#_c_1060_n N_VPWR_c_1610_n 0.0038194f $X=9.08 $Y=2.135 $X2=0
+ $Y2=0
cc_813 N_A_1278_529#_c_1061_n N_VPWR_c_1617_n 0.0122081f $X=6.53 $Y=2.855 $X2=0
+ $Y2=0
cc_814 N_A_1278_529#_c_1064_n N_VPWR_c_1618_n 0.00223296f $X=8.28 $Y=2.15 $X2=0
+ $Y2=0
cc_815 N_A_1278_529#_c_1067_n N_VPWR_c_1618_n 0.0382385f $X=8.285 $Y=2.685 $X2=0
+ $Y2=0
cc_816 N_A_1278_529#_c_1060_n N_VPWR_c_1597_n 0.00681349f $X=9.08 $Y=2.135 $X2=0
+ $Y2=0
cc_817 N_A_1278_529#_c_1061_n N_VPWR_c_1597_n 0.0106598f $X=6.53 $Y=2.855 $X2=0
+ $Y2=0
cc_818 N_A_1278_529#_c_1064_n N_VPWR_c_1597_n 0.00194834f $X=8.28 $Y=2.15 $X2=0
+ $Y2=0
cc_819 N_A_1278_529#_c_1065_n N_VPWR_c_1597_n 0.0147292f $X=7 $Y=2.42 $X2=0
+ $Y2=0
cc_820 N_A_1278_529#_c_1066_n N_VPWR_c_1597_n 0.0059121f $X=7.625 $Y=2.685 $X2=0
+ $Y2=0
cc_821 N_A_1278_529#_c_1067_n N_VPWR_c_1597_n 0.0283163f $X=8.285 $Y=2.685 $X2=0
+ $Y2=0
cc_822 N_A_1278_529#_c_1060_n N_VPWR_c_1625_n 0.00658031f $X=9.08 $Y=2.135 $X2=0
+ $Y2=0
cc_823 N_A_1278_529#_c_1067_n N_VPWR_c_1625_n 0.00259155f $X=8.285 $Y=2.685
+ $X2=0 $Y2=0
cc_824 N_A_1278_529#_c_1061_n N_A_229_491#_c_1777_n 0.0069396f $X=6.53 $Y=2.855
+ $X2=0 $Y2=0
cc_825 N_A_1278_529#_c_1065_n N_A_229_491#_c_1777_n 0.0079335f $X=7 $Y=2.42
+ $X2=0 $Y2=0
cc_826 N_A_1278_529#_c_1061_n N_A_229_491#_c_1778_n 0.0035758f $X=6.53 $Y=2.855
+ $X2=0 $Y2=0
cc_827 N_A_1278_529#_M1001_g N_VGND_c_1946_n 0.00133853f $X=8.615 $Y=0.955 $X2=0
+ $Y2=0
cc_828 N_A_1278_529#_M1001_g N_VGND_c_1955_n 9.53055e-19 $X=8.615 $Y=0.955 $X2=0
+ $Y2=0
cc_829 N_A_857_367#_c_1178_n N_A_2064_101#_M1029_g 0.0518916f $X=9.96 $Y=1.47
+ $X2=0 $Y2=0
cc_830 N_A_857_367#_M1024_g N_A_2064_101#_c_1327_n 0.0518916f $X=10.035 $Y=2.875
+ $X2=0 $Y2=0
cc_831 N_A_857_367#_M1016_g N_A_1870_127#_c_1419_n 0.00138099f $X=9.275 $Y=0.955
+ $X2=0 $Y2=0
cc_832 N_A_857_367#_M1016_g N_A_1870_127#_c_1420_n 5.02696e-19 $X=9.275 $Y=0.955
+ $X2=0 $Y2=0
cc_833 N_A_857_367#_c_1178_n N_A_1870_127#_c_1420_n 0.0145101f $X=9.96 $Y=1.47
+ $X2=0 $Y2=0
cc_834 N_A_857_367#_M1024_g N_A_1870_127#_c_1420_n 0.0168826f $X=10.035 $Y=2.875
+ $X2=0 $Y2=0
cc_835 N_A_857_367#_c_1178_n N_A_1870_127#_c_1421_n 0.00298893f $X=9.96 $Y=1.47
+ $X2=0 $Y2=0
cc_836 N_A_857_367#_M1016_g N_A_1870_127#_c_1423_n 0.00126391f $X=9.275 $Y=0.955
+ $X2=0 $Y2=0
cc_837 N_A_857_367#_c_1178_n N_A_1870_127#_c_1423_n 0.00760139f $X=9.96 $Y=1.47
+ $X2=0 $Y2=0
cc_838 N_A_857_367#_M1024_g N_A_1870_127#_c_1429_n 0.00716766f $X=10.035
+ $Y=2.875 $X2=0 $Y2=0
cc_839 N_A_857_367#_c_1190_n N_VPWR_M1022_s 0.00681128f $X=5.045 $Y=2.095 $X2=0
+ $Y2=0
cc_840 N_A_857_367#_c_1183_n N_VPWR_M1022_s 0.00435145f $X=5.13 $Y=1.46 $X2=0
+ $Y2=0
cc_841 N_A_857_367#_M1022_g N_VPWR_c_1601_n 0.015072f $X=5.325 $Y=2.465 $X2=0
+ $Y2=0
cc_842 N_A_857_367#_M1024_g N_VPWR_c_1610_n 0.00351226f $X=10.035 $Y=2.875 $X2=0
+ $Y2=0
cc_843 N_A_857_367#_M1022_g N_VPWR_c_1617_n 0.00364644f $X=5.325 $Y=2.465 $X2=0
+ $Y2=0
cc_844 N_A_857_367#_c_1187_n N_VPWR_c_1617_n 0.00555245f $X=6.315 $Y=2.535 $X2=0
+ $Y2=0
cc_845 N_A_857_367#_M1035_d N_VPWR_c_1597_n 0.00348066f $X=4.285 $Y=1.835 $X2=0
+ $Y2=0
cc_846 N_A_857_367#_M1022_g N_VPWR_c_1597_n 0.00578802f $X=5.325 $Y=2.465 $X2=0
+ $Y2=0
cc_847 N_A_857_367#_c_1187_n N_VPWR_c_1597_n 0.0117713f $X=6.315 $Y=2.535 $X2=0
+ $Y2=0
cc_848 N_A_857_367#_M1024_g N_VPWR_c_1597_n 0.00539338f $X=10.035 $Y=2.875 $X2=0
+ $Y2=0
cc_849 N_A_857_367#_c_1190_n N_A_229_491#_c_1771_n 0.00906358f $X=5.045 $Y=2.095
+ $X2=0 $Y2=0
cc_850 N_A_857_367#_c_1182_n N_A_229_491#_c_1771_n 0.00889803f $X=5.045 $Y=1.065
+ $X2=0 $Y2=0
cc_851 N_A_857_367#_M1023_d N_A_229_491#_c_1772_n 0.00709212f $X=4.41 $Y=0.345
+ $X2=0 $Y2=0
cc_852 N_A_857_367#_M1019_g N_A_229_491#_c_1772_n 0.01997f $X=5.325 $Y=0.655
+ $X2=0 $Y2=0
cc_853 N_A_857_367#_c_1171_n N_A_229_491#_c_1772_n 0.00134281f $X=5.99 $Y=1.5
+ $X2=0 $Y2=0
cc_854 N_A_857_367#_c_1182_n N_A_229_491#_c_1772_n 0.0569176f $X=5.045 $Y=1.065
+ $X2=0 $Y2=0
cc_855 N_A_857_367#_c_1184_n N_A_229_491#_c_1772_n 6.68148e-19 $X=5.4 $Y=1.46
+ $X2=0 $Y2=0
cc_856 N_A_857_367#_M1035_d N_A_229_491#_c_1777_n 0.00689834f $X=4.285 $Y=1.835
+ $X2=0 $Y2=0
cc_857 N_A_857_367#_M1022_g N_A_229_491#_c_1777_n 0.0160842f $X=5.325 $Y=2.465
+ $X2=0 $Y2=0
cc_858 N_A_857_367#_c_1187_n N_A_229_491#_c_1777_n 0.00157638f $X=6.315 $Y=2.535
+ $X2=0 $Y2=0
cc_859 N_A_857_367#_c_1189_n N_A_229_491#_c_1777_n 0.0137412f $X=6.315 $Y=2.46
+ $X2=0 $Y2=0
cc_860 N_A_857_367#_c_1190_n N_A_229_491#_c_1777_n 0.0629193f $X=5.045 $Y=2.095
+ $X2=0 $Y2=0
cc_861 N_A_857_367#_M1022_g N_A_229_491#_c_1778_n 0.00840606f $X=5.325 $Y=2.465
+ $X2=0 $Y2=0
cc_862 N_A_857_367#_c_1187_n N_A_229_491#_c_1778_n 0.00136846f $X=6.315 $Y=2.535
+ $X2=0 $Y2=0
cc_863 N_A_857_367#_M1019_g N_A_229_491#_c_1774_n 0.00386161f $X=5.325 $Y=0.655
+ $X2=0 $Y2=0
cc_864 N_A_857_367#_c_1182_n N_VGND_M1019_s 0.00380435f $X=5.045 $Y=1.065 $X2=0
+ $Y2=0
cc_865 N_A_857_367#_M1019_g N_VGND_c_1945_n 0.0154878f $X=5.325 $Y=0.655 $X2=0
+ $Y2=0
cc_866 N_A_857_367#_c_1175_n N_VGND_c_1946_n 0.0248335f $X=9.2 $Y=0.18 $X2=0
+ $Y2=0
cc_867 N_A_857_367#_M1019_g N_VGND_c_1951_n 0.0035231f $X=5.325 $Y=0.655 $X2=0
+ $Y2=0
cc_868 N_A_857_367#_c_1176_n N_VGND_c_1951_n 0.0267761f $X=7.185 $Y=0.18 $X2=0
+ $Y2=0
cc_869 N_A_857_367#_c_1175_n N_VGND_c_1952_n 0.0229198f $X=9.2 $Y=0.18 $X2=0
+ $Y2=0
cc_870 N_A_857_367#_M1019_g N_VGND_c_1955_n 0.00557134f $X=5.325 $Y=0.655 $X2=0
+ $Y2=0
cc_871 N_A_857_367#_c_1175_n N_VGND_c_1955_n 0.0515628f $X=9.2 $Y=0.18 $X2=0
+ $Y2=0
cc_872 N_A_857_367#_c_1176_n N_VGND_c_1955_n 0.00549737f $X=7.185 $Y=0.18 $X2=0
+ $Y2=0
cc_873 N_A_2064_101#_c_1328_n N_A_1870_127#_M1013_g 0.00458193f $X=11.245
+ $Y=2.875 $X2=0 $Y2=0
cc_874 N_A_2064_101#_c_1329_n N_A_1870_127#_M1013_g 0.00879189f $X=11.305
+ $Y=2.175 $X2=0 $Y2=0
cc_875 N_A_2064_101#_c_1330_n N_A_1870_127#_M1013_g 0.0141851f $X=11.77 $Y=1.88
+ $X2=0 $Y2=0
cc_876 N_A_2064_101#_c_1331_n N_A_1870_127#_M1013_g 0.00139238f $X=11.39 $Y=1.88
+ $X2=0 $Y2=0
cc_877 N_A_2064_101#_c_1323_n N_A_1870_127#_M1013_g 0.00647803f $X=11.855
+ $Y=1.795 $X2=0 $Y2=0
cc_878 N_A_2064_101#_c_1333_n N_A_1870_127#_M1013_g 0.0118896f $X=11.235 $Y=2.34
+ $X2=0 $Y2=0
cc_879 N_A_2064_101#_c_1330_n N_A_1870_127#_c_1413_n 0.00244727f $X=11.77
+ $Y=1.88 $X2=0 $Y2=0
cc_880 N_A_2064_101#_c_1323_n N_A_1870_127#_c_1413_n 0.0142386f $X=11.855
+ $Y=1.795 $X2=0 $Y2=0
cc_881 N_A_2064_101#_c_1330_n N_A_1870_127#_M1004_g 8.16897e-19 $X=11.77 $Y=1.88
+ $X2=0 $Y2=0
cc_882 N_A_2064_101#_c_1323_n N_A_1870_127#_M1004_g 0.00183276f $X=11.855
+ $Y=1.795 $X2=0 $Y2=0
cc_883 N_A_2064_101#_c_1323_n N_A_1870_127#_c_1417_n 0.00124637f $X=11.855
+ $Y=1.795 $X2=0 $Y2=0
cc_884 N_A_2064_101#_M1029_g N_A_1870_127#_c_1419_n 0.00145853f $X=10.395
+ $Y=0.845 $X2=0 $Y2=0
cc_885 N_A_2064_101#_M1029_g N_A_1870_127#_c_1420_n 0.00292054f $X=10.395
+ $Y=0.845 $X2=0 $Y2=0
cc_886 N_A_2064_101#_M1030_d N_A_1870_127#_c_1421_n 8.67508e-19 $X=11.49
+ $Y=0.635 $X2=0 $Y2=0
cc_887 N_A_2064_101#_M1029_g N_A_1870_127#_c_1421_n 0.015939f $X=10.395 $Y=0.845
+ $X2=0 $Y2=0
cc_888 N_A_2064_101#_c_1331_n N_A_1870_127#_c_1421_n 0.00425742f $X=11.39
+ $Y=1.88 $X2=0 $Y2=0
cc_889 N_A_2064_101#_c_1322_n N_A_1870_127#_c_1421_n 0.00618249f $X=11.77
+ $Y=0.725 $X2=0 $Y2=0
cc_890 N_A_2064_101#_c_1323_n N_A_1870_127#_c_1421_n 0.0147776f $X=11.855
+ $Y=1.795 $X2=0 $Y2=0
cc_891 N_A_2064_101#_c_1330_n N_A_1870_127#_c_1422_n 0.0100085f $X=11.77 $Y=1.88
+ $X2=0 $Y2=0
cc_892 N_A_2064_101#_c_1331_n N_A_1870_127#_c_1422_n 0.00275952f $X=11.39
+ $Y=1.88 $X2=0 $Y2=0
cc_893 N_A_2064_101#_c_1323_n N_A_1870_127#_c_1422_n 0.0209558f $X=11.855
+ $Y=1.795 $X2=0 $Y2=0
cc_894 N_A_2064_101#_M1029_g N_A_1870_127#_c_1423_n 0.00276273f $X=10.395
+ $Y=0.845 $X2=0 $Y2=0
cc_895 N_A_2064_101#_c_1330_n N_A_1870_127#_c_1424_n 0.00271849f $X=11.77
+ $Y=1.88 $X2=0 $Y2=0
cc_896 N_A_2064_101#_c_1331_n N_A_1870_127#_c_1424_n 3.21804e-19 $X=11.39
+ $Y=1.88 $X2=0 $Y2=0
cc_897 N_A_2064_101#_c_1322_n N_A_1870_127#_c_1424_n 0.00554605f $X=11.77
+ $Y=0.725 $X2=0 $Y2=0
cc_898 N_A_2064_101#_c_1323_n N_A_1870_127#_c_1424_n 0.00168553f $X=11.855
+ $Y=1.795 $X2=0 $Y2=0
cc_899 N_A_2064_101#_c_1322_n N_A_1870_127#_c_1425_n 0.00615417f $X=11.77
+ $Y=0.725 $X2=0 $Y2=0
cc_900 N_A_2064_101#_c_1323_n N_A_1870_127#_c_1425_n 0.00340935f $X=11.855
+ $Y=1.795 $X2=0 $Y2=0
cc_901 N_A_2064_101#_c_1330_n N_A_2370_351#_M1004_s 0.00327322f $X=11.77 $Y=1.88
+ $X2=0 $Y2=0
cc_902 N_A_2064_101#_c_1323_n N_A_2370_351#_M1004_s 5.10436e-19 $X=11.855
+ $Y=1.795 $X2=0 $Y2=0
cc_903 N_A_2064_101#_c_1329_n N_A_2370_351#_c_1544_n 0.0015384f $X=11.305
+ $Y=2.175 $X2=0 $Y2=0
cc_904 N_A_2064_101#_c_1330_n N_A_2370_351#_c_1544_n 0.0110294f $X=11.77 $Y=1.88
+ $X2=0 $Y2=0
cc_905 N_A_2064_101#_c_1333_n N_A_2370_351#_c_1544_n 0.0104741f $X=11.235
+ $Y=2.34 $X2=0 $Y2=0
cc_906 N_A_2064_101#_c_1322_n N_A_2370_351#_c_1538_n 0.0216869f $X=11.77
+ $Y=0.725 $X2=0 $Y2=0
cc_907 N_A_2064_101#_c_1323_n N_A_2370_351#_c_1538_n 0.0309048f $X=11.855
+ $Y=1.795 $X2=0 $Y2=0
cc_908 N_A_2064_101#_c_1323_n N_A_2370_351#_c_1545_n 0.0133866f $X=11.855
+ $Y=1.795 $X2=0 $Y2=0
cc_909 N_A_2064_101#_c_1323_n N_A_2370_351#_c_1541_n 0.027453f $X=11.855
+ $Y=1.795 $X2=0 $Y2=0
cc_910 N_A_2064_101#_M1012_g N_VPWR_c_1603_n 0.00715047f $X=10.395 $Y=2.875
+ $X2=0 $Y2=0
cc_911 N_A_2064_101#_c_1326_n N_VPWR_c_1603_n 0.0230771f $X=11.08 $Y=2.34 $X2=0
+ $Y2=0
cc_912 N_A_2064_101#_c_1327_n N_VPWR_c_1603_n 0.00466427f $X=10.58 $Y=2.34 $X2=0
+ $Y2=0
cc_913 N_A_2064_101#_c_1328_n N_VPWR_c_1603_n 0.0239156f $X=11.245 $Y=2.875
+ $X2=0 $Y2=0
cc_914 N_A_2064_101#_M1012_g N_VPWR_c_1610_n 0.00575161f $X=10.395 $Y=2.875
+ $X2=0 $Y2=0
cc_915 N_A_2064_101#_c_1328_n N_VPWR_c_1612_n 0.01714f $X=11.245 $Y=2.875 $X2=0
+ $Y2=0
cc_916 N_A_2064_101#_M1033_d N_VPWR_c_1597_n 0.0022756f $X=11.105 $Y=2.665 $X2=0
+ $Y2=0
cc_917 N_A_2064_101#_M1012_g N_VPWR_c_1597_n 0.0110767f $X=10.395 $Y=2.875 $X2=0
+ $Y2=0
cc_918 N_A_2064_101#_c_1326_n N_VPWR_c_1597_n 0.00960911f $X=11.08 $Y=2.34 $X2=0
+ $Y2=0
cc_919 N_A_2064_101#_c_1327_n N_VPWR_c_1597_n 0.00162464f $X=10.58 $Y=2.34 $X2=0
+ $Y2=0
cc_920 N_A_2064_101#_c_1328_n N_VPWR_c_1597_n 0.0114757f $X=11.245 $Y=2.875
+ $X2=0 $Y2=0
cc_921 N_A_2064_101#_c_1333_n N_VPWR_c_1597_n 3.62543e-19 $X=11.235 $Y=2.34
+ $X2=0 $Y2=0
cc_922 N_A_2064_101#_M1029_g N_VGND_c_1947_n 0.0069431f $X=10.395 $Y=0.845 $X2=0
+ $Y2=0
cc_923 N_A_2064_101#_c_1322_n N_VGND_c_1947_n 0.00796204f $X=11.77 $Y=0.725
+ $X2=0 $Y2=0
cc_924 N_A_2064_101#_M1029_g N_VGND_c_1952_n 0.00410092f $X=10.395 $Y=0.845
+ $X2=0 $Y2=0
cc_925 N_A_2064_101#_c_1322_n N_VGND_c_1953_n 0.0099398f $X=11.77 $Y=0.725 $X2=0
+ $Y2=0
cc_926 N_A_2064_101#_M1029_g N_VGND_c_1955_n 0.00466677f $X=10.395 $Y=0.845
+ $X2=0 $Y2=0
cc_927 N_A_2064_101#_c_1322_n N_VGND_c_1955_n 0.0144173f $X=11.77 $Y=0.725 $X2=0
+ $Y2=0
cc_928 N_A_1870_127#_M1004_g N_A_2370_351#_M1025_g 0.017395f $X=12.19 $Y=2.075
+ $X2=0 $Y2=0
cc_929 N_A_1870_127#_M1013_g N_A_2370_351#_c_1544_n 0.00283789f $X=11.46
+ $Y=2.875 $X2=0 $Y2=0
cc_930 N_A_1870_127#_M1004_g N_A_2370_351#_c_1544_n 0.012883f $X=12.19 $Y=2.075
+ $X2=0 $Y2=0
cc_931 N_A_1870_127#_c_1413_n N_A_2370_351#_c_1538_n 0.00140486f $X=12.115
+ $Y=1.24 $X2=0 $Y2=0
cc_932 N_A_1870_127#_c_1414_n N_A_2370_351#_c_1538_n 0.00581294f $X=12.19
+ $Y=1.165 $X2=0 $Y2=0
cc_933 N_A_1870_127#_c_1416_n N_A_2370_351#_c_1538_n 0.00306045f $X=12.44
+ $Y=0.845 $X2=0 $Y2=0
cc_934 N_A_1870_127#_c_1417_n N_A_2370_351#_c_1538_n 0.013503f $X=12.44 $Y=0.92
+ $X2=0 $Y2=0
cc_935 N_A_1870_127#_c_1418_n N_A_2370_351#_c_1538_n 0.0025487f $X=12.19 $Y=1.24
+ $X2=0 $Y2=0
cc_936 N_A_1870_127#_c_1425_n N_A_2370_351#_c_1538_n 0.0023775f $X=11.505
+ $Y=1.165 $X2=0 $Y2=0
cc_937 N_A_1870_127#_M1004_g N_A_2370_351#_c_1545_n 0.0151773f $X=12.19 $Y=2.075
+ $X2=0 $Y2=0
cc_938 N_A_1870_127#_c_1417_n N_A_2370_351#_c_1539_n 0.00629386f $X=12.44
+ $Y=0.92 $X2=0 $Y2=0
cc_939 N_A_1870_127#_c_1418_n N_A_2370_351#_c_1540_n 0.00918211f $X=12.19
+ $Y=1.24 $X2=0 $Y2=0
cc_940 N_A_1870_127#_c_1413_n N_A_2370_351#_c_1541_n 7.24799e-19 $X=12.115
+ $Y=1.24 $X2=0 $Y2=0
cc_941 N_A_1870_127#_M1004_g N_A_2370_351#_c_1541_n 0.0101671f $X=12.19 $Y=2.075
+ $X2=0 $Y2=0
cc_942 N_A_1870_127#_c_1418_n N_A_2370_351#_c_1541_n 0.00149073f $X=12.19
+ $Y=1.24 $X2=0 $Y2=0
cc_943 N_A_1870_127#_c_1414_n N_A_2370_351#_c_1542_n 0.00242909f $X=12.19
+ $Y=1.165 $X2=0 $Y2=0
cc_944 N_A_1870_127#_c_1416_n N_A_2370_351#_c_1542_n 0.0152431f $X=12.44
+ $Y=0.845 $X2=0 $Y2=0
cc_945 N_A_1870_127#_M1013_g N_VPWR_c_1604_n 0.00507981f $X=11.46 $Y=2.875 $X2=0
+ $Y2=0
cc_946 N_A_1870_127#_M1004_g N_VPWR_c_1607_n 0.00509193f $X=12.19 $Y=2.075 $X2=0
+ $Y2=0
cc_947 N_A_1870_127#_M1013_g N_VPWR_c_1612_n 0.00575161f $X=11.46 $Y=2.875 $X2=0
+ $Y2=0
cc_948 N_A_1870_127#_M1006_d N_VPWR_c_1597_n 0.00301588f $X=9.585 $Y=2.245 $X2=0
+ $Y2=0
cc_949 N_A_1870_127#_M1013_g N_VPWR_c_1597_n 0.0118168f $X=11.46 $Y=2.875 $X2=0
+ $Y2=0
cc_950 N_A_1870_127#_M1004_g N_VPWR_c_1597_n 0.00391649f $X=12.19 $Y=2.075 $X2=0
+ $Y2=0
cc_951 N_A_1870_127#_c_1421_n N_VGND_M1029_d 0.00634624f $X=11.34 $Y=1.115 $X2=0
+ $Y2=0
cc_952 N_A_1870_127#_c_1419_n N_VGND_c_1947_n 0.00668622f $X=9.705 $Y=0.79 $X2=0
+ $Y2=0
cc_953 N_A_1870_127#_c_1421_n N_VGND_c_1947_n 0.0267886f $X=11.34 $Y=1.115 $X2=0
+ $Y2=0
cc_954 N_A_1870_127#_c_1414_n N_VGND_c_1948_n 3.60091e-19 $X=12.19 $Y=1.165
+ $X2=0 $Y2=0
cc_955 N_A_1870_127#_c_1416_n N_VGND_c_1948_n 0.00685589f $X=12.44 $Y=0.845
+ $X2=0 $Y2=0
cc_956 N_A_1870_127#_c_1416_n N_VGND_c_1953_n 0.00508422f $X=12.44 $Y=0.845
+ $X2=0 $Y2=0
cc_957 N_A_1870_127#_c_1425_n N_VGND_c_1953_n 0.00394205f $X=11.505 $Y=1.165
+ $X2=0 $Y2=0
cc_958 N_A_1870_127#_c_1416_n N_VGND_c_1955_n 0.0105555f $X=12.44 $Y=0.845 $X2=0
+ $Y2=0
cc_959 N_A_1870_127#_c_1417_n N_VGND_c_1955_n 2.23561e-19 $X=12.44 $Y=0.92 $X2=0
+ $Y2=0
cc_960 N_A_1870_127#_c_1425_n N_VGND_c_1955_n 0.00466677f $X=11.505 $Y=1.165
+ $X2=0 $Y2=0
cc_961 N_A_1870_127#_c_1421_n A_2022_127# 0.00368839f $X=11.34 $Y=1.115
+ $X2=-0.19 $Y2=-0.245
cc_962 N_A_1870_127#_c_1421_n A_2226_127# 0.00368839f $X=11.34 $Y=1.115
+ $X2=-0.19 $Y2=-0.245
cc_963 N_A_2370_351#_c_1544_n N_VPWR_c_1604_n 0.00173188f $X=12.11 $Y=2.275
+ $X2=0 $Y2=0
cc_964 N_A_2370_351#_M1025_g N_VPWR_c_1607_n 0.0217568f $X=12.81 $Y=2.465 $X2=0
+ $Y2=0
cc_965 N_A_2370_351#_c_1544_n N_VPWR_c_1607_n 0.011725f $X=12.11 $Y=2.275 $X2=0
+ $Y2=0
cc_966 N_A_2370_351#_c_1539_n N_VPWR_c_1607_n 0.0223333f $X=12.83 $Y=1.43 $X2=0
+ $Y2=0
cc_967 N_A_2370_351#_c_1540_n N_VPWR_c_1607_n 0.00102501f $X=12.83 $Y=1.43 $X2=0
+ $Y2=0
cc_968 N_A_2370_351#_M1025_g N_VPWR_c_1619_n 0.00579312f $X=12.81 $Y=2.465 $X2=0
+ $Y2=0
cc_969 N_A_2370_351#_M1025_g N_VPWR_c_1597_n 0.0129818f $X=12.81 $Y=2.465 $X2=0
+ $Y2=0
cc_970 N_A_2370_351#_M1025_g Q 0.0127209f $X=12.81 $Y=2.465 $X2=0 $Y2=0
cc_971 N_A_2370_351#_M1025_g N_Q_c_1923_n 0.00695714f $X=12.81 $Y=2.465 $X2=0
+ $Y2=0
cc_972 N_A_2370_351#_c_1539_n N_Q_c_1923_n 0.0270346f $X=12.83 $Y=1.43 $X2=0
+ $Y2=0
cc_973 N_A_2370_351#_c_1542_n N_Q_c_1923_n 0.0163097f $X=12.852 $Y=1.265 $X2=0
+ $Y2=0
cc_974 N_A_2370_351#_M1025_g N_Q_c_1926_n 0.0025085f $X=12.81 $Y=2.465 $X2=0
+ $Y2=0
cc_975 N_A_2370_351#_c_1539_n N_Q_c_1926_n 0.00234559f $X=12.83 $Y=1.43 $X2=0
+ $Y2=0
cc_976 N_A_2370_351#_c_1540_n N_Q_c_1926_n 0.00650555f $X=12.83 $Y=1.43 $X2=0
+ $Y2=0
cc_977 N_A_2370_351#_c_1538_n N_VGND_c_1948_n 0.0290121f $X=12.225 $Y=0.515
+ $X2=0 $Y2=0
cc_978 N_A_2370_351#_c_1539_n N_VGND_c_1948_n 0.0301215f $X=12.83 $Y=1.43 $X2=0
+ $Y2=0
cc_979 N_A_2370_351#_c_1540_n N_VGND_c_1948_n 0.00565946f $X=12.83 $Y=1.43 $X2=0
+ $Y2=0
cc_980 N_A_2370_351#_c_1542_n N_VGND_c_1948_n 0.0210354f $X=12.852 $Y=1.265
+ $X2=0 $Y2=0
cc_981 N_A_2370_351#_c_1538_n N_VGND_c_1953_n 0.00960818f $X=12.225 $Y=0.515
+ $X2=0 $Y2=0
cc_982 N_A_2370_351#_c_1542_n N_VGND_c_1954_n 0.00422142f $X=12.852 $Y=1.265
+ $X2=0 $Y2=0
cc_983 N_A_2370_351#_c_1538_n N_VGND_c_1955_n 0.0089748f $X=12.225 $Y=0.515
+ $X2=0 $Y2=0
cc_984 N_A_2370_351#_c_1542_n N_VGND_c_1955_n 0.00837013f $X=12.852 $Y=1.265
+ $X2=0 $Y2=0
cc_985 N_VPWR_c_1597_n N_A_229_491#_M1032_s 0.00227393f $X=13.2 $Y=3.33 $X2=0
+ $Y2=0
cc_986 N_VPWR_c_1597_n N_A_229_491#_M1018_d 0.00335595f $X=13.2 $Y=3.33 $X2=0
+ $Y2=0
cc_987 N_VPWR_M1037_d N_A_229_491#_c_1781_n 0.0159269f $X=1.92 $Y=2.455 $X2=0
+ $Y2=0
cc_988 N_VPWR_c_1608_n N_A_229_491#_c_1781_n 0.0103265f $X=3.755 $Y=3.33 $X2=0
+ $Y2=0
cc_989 N_VPWR_c_1597_n N_A_229_491#_c_1781_n 0.034005f $X=13.2 $Y=3.33 $X2=0
+ $Y2=0
cc_990 N_VPWR_c_1621_n N_A_229_491#_c_1781_n 0.00951383f $X=1.955 $Y=3.185 $X2=0
+ $Y2=0
cc_991 N_VPWR_c_1622_n N_A_229_491#_c_1781_n 0.0459946f $X=2.625 $Y=3.185 $X2=0
+ $Y2=0
cc_992 N_VPWR_M1000_d N_A_229_491#_c_1775_n 0.00101618f $X=3.71 $Y=2.455 $X2=0
+ $Y2=0
cc_993 N_VPWR_c_1600_n N_A_229_491#_c_1775_n 0.0078049f $X=3.92 $Y=2.88 $X2=0
+ $Y2=0
cc_994 N_VPWR_c_1608_n N_A_229_491#_c_1775_n 0.00263044f $X=3.755 $Y=3.33 $X2=0
+ $Y2=0
cc_995 N_VPWR_c_1597_n N_A_229_491#_c_1775_n 0.00585474f $X=13.2 $Y=3.33 $X2=0
+ $Y2=0
cc_996 N_VPWR_M1000_d N_A_229_491#_c_1771_n 0.00923121f $X=3.71 $Y=2.455 $X2=0
+ $Y2=0
cc_997 N_VPWR_M1000_d N_A_229_491#_c_1777_n 0.00107952f $X=3.71 $Y=2.455 $X2=0
+ $Y2=0
cc_998 N_VPWR_M1022_s N_A_229_491#_c_1777_n 0.00503476f $X=4.985 $Y=1.835 $X2=0
+ $Y2=0
cc_999 N_VPWR_c_1600_n N_A_229_491#_c_1777_n 0.00333414f $X=3.92 $Y=2.88 $X2=0
+ $Y2=0
cc_1000 N_VPWR_c_1601_n N_A_229_491#_c_1777_n 0.0211807f $X=5.11 $Y=2.88 $X2=0
+ $Y2=0
cc_1001 N_VPWR_c_1616_n N_A_229_491#_c_1777_n 0.0117107f $X=4.945 $Y=3.33 $X2=0
+ $Y2=0
cc_1002 N_VPWR_c_1617_n N_A_229_491#_c_1777_n 0.00881392f $X=7.155 $Y=3.33 $X2=0
+ $Y2=0
cc_1003 N_VPWR_c_1597_n N_A_229_491#_c_1777_n 0.0399236f $X=13.2 $Y=3.33 $X2=0
+ $Y2=0
cc_1004 N_VPWR_c_1601_n N_A_229_491#_c_1778_n 0.00721615f $X=5.11 $Y=2.88 $X2=0
+ $Y2=0
cc_1005 N_VPWR_c_1617_n N_A_229_491#_c_1778_n 0.0151227f $X=7.155 $Y=3.33 $X2=0
+ $Y2=0
cc_1006 N_VPWR_c_1597_n N_A_229_491#_c_1778_n 0.0119668f $X=13.2 $Y=3.33 $X2=0
+ $Y2=0
cc_1007 N_VPWR_c_1597_n N_A_229_491#_c_1779_n 0.0116139f $X=13.2 $Y=3.33 $X2=0
+ $Y2=0
cc_1008 N_VPWR_c_1621_n N_A_229_491#_c_1779_n 0.0118206f $X=1.955 $Y=3.185 $X2=0
+ $Y2=0
cc_1009 N_VPWR_c_1608_n N_A_229_491#_c_1780_n 0.0200147f $X=3.755 $Y=3.33 $X2=0
+ $Y2=0
cc_1010 N_VPWR_c_1597_n N_A_229_491#_c_1780_n 0.0127015f $X=13.2 $Y=3.33 $X2=0
+ $Y2=0
cc_1011 N_VPWR_M1000_d N_A_229_491#_c_1834_n 0.0034854f $X=3.71 $Y=2.455 $X2=0
+ $Y2=0
cc_1012 N_VPWR_c_1600_n N_A_229_491#_c_1834_n 0.0146685f $X=3.92 $Y=2.88 $X2=0
+ $Y2=0
cc_1013 N_VPWR_c_1597_n N_A_229_491#_c_1834_n 7.31729e-19 $X=13.2 $Y=3.33 $X2=0
+ $Y2=0
cc_1014 N_VPWR_c_1597_n A_312_491# 0.00218036f $X=13.2 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_1015 N_VPWR_c_1597_n A_562_491# 0.00218036f $X=13.2 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_1016 N_VPWR_c_1597_n A_2022_533# 0.00186271f $X=13.2 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_1017 N_VPWR_c_1597_n N_Q_M1025_d 0.00231914f $X=13.2 $Y=3.33 $X2=0 $Y2=0
cc_1018 N_VPWR_c_1619_n Q 0.0307672f $X=13.2 $Y=3.33 $X2=0 $Y2=0
cc_1019 N_VPWR_c_1597_n Q 0.0179089f $X=13.2 $Y=3.33 $X2=0 $Y2=0
cc_1020 N_VPWR_c_1607_n N_Q_c_1923_n 0.00229217f $X=12.535 $Y=1.96 $X2=0 $Y2=0
cc_1021 N_VPWR_c_1607_n N_Q_c_1926_n 0.0505473f $X=12.535 $Y=1.96 $X2=0 $Y2=0
cc_1022 N_A_229_491#_c_1781_n A_312_491# 0.00245508f $X=3.195 $Y=2.7 $X2=-0.19
+ $Y2=-0.245
cc_1023 N_A_229_491#_c_1781_n A_562_491# 0.00248105f $X=3.195 $Y=2.7 $X2=-0.19
+ $Y2=-0.245
cc_1024 N_A_229_491#_c_1770_n N_VGND_M1034_d 4.0491e-19 $X=3.865 $Y=0.77 $X2=0
+ $Y2=0
cc_1025 N_A_229_491#_c_1771_n N_VGND_M1034_d 0.00472966f $X=3.95 $Y=2.365 $X2=0
+ $Y2=0
cc_1026 N_A_229_491#_c_1772_n N_VGND_M1034_d 0.00698319f $X=6.04 $Y=0.71 $X2=0
+ $Y2=0
cc_1027 N_A_229_491#_c_1826_n N_VGND_M1034_d 0.00439989f $X=3.95 $Y=0.74 $X2=0
+ $Y2=0
cc_1028 N_A_229_491#_c_1772_n N_VGND_M1019_s 0.00544797f $X=6.04 $Y=0.71 $X2=0
+ $Y2=0
cc_1029 N_A_229_491#_c_1772_n N_VGND_c_1944_n 0.012734f $X=6.04 $Y=0.71 $X2=0
+ $Y2=0
cc_1030 N_A_229_491#_c_1826_n N_VGND_c_1944_n 0.0133441f $X=3.95 $Y=0.74 $X2=0
+ $Y2=0
cc_1031 N_A_229_491#_c_1772_n N_VGND_c_1945_n 0.020491f $X=6.04 $Y=0.71 $X2=0
+ $Y2=0
cc_1032 N_A_229_491#_c_1770_n N_VGND_c_1949_n 0.00395912f $X=3.865 $Y=0.77 $X2=0
+ $Y2=0
cc_1033 N_A_229_491#_c_1772_n N_VGND_c_1950_n 0.0123411f $X=6.04 $Y=0.71 $X2=0
+ $Y2=0
cc_1034 N_A_229_491#_c_1772_n N_VGND_c_1951_n 0.013248f $X=6.04 $Y=0.71 $X2=0
+ $Y2=0
cc_1035 N_A_229_491#_c_1774_n N_VGND_c_1951_n 0.00485742f $X=6.165 $Y=0.71 $X2=0
+ $Y2=0
cc_1036 N_A_229_491#_c_1770_n N_VGND_c_1955_n 0.00998677f $X=3.865 $Y=0.77 $X2=0
+ $Y2=0
cc_1037 N_A_229_491#_c_1772_n N_VGND_c_1955_n 0.0443353f $X=6.04 $Y=0.71 $X2=0
+ $Y2=0
cc_1038 N_A_229_491#_c_1826_n N_VGND_c_1955_n 0.00117688f $X=3.95 $Y=0.74 $X2=0
+ $Y2=0
cc_1039 N_A_229_491#_c_1774_n N_VGND_c_1955_n 0.00734198f $X=6.165 $Y=0.71 $X2=0
+ $Y2=0
cc_1040 N_A_229_491#_c_1770_n N_noxref_24_M1015_d 0.00312542f $X=3.865 $Y=0.77
+ $X2=0 $Y2=0
cc_1041 N_A_229_491#_c_1770_n N_noxref_24_c_2074_n 0.0193962f $X=3.865 $Y=0.77
+ $X2=0 $Y2=0
cc_1042 N_A_229_491#_M1028_d N_noxref_24_c_2075_n 0.00552774f $X=2.165 $Y=0.295
+ $X2=0 $Y2=0
cc_1043 N_A_229_491#_c_1770_n N_noxref_24_c_2075_n 0.0217022f $X=3.865 $Y=0.77
+ $X2=0 $Y2=0
cc_1044 N_A_229_491#_c_1773_n N_noxref_24_c_2075_n 0.0232304f $X=2.585 $Y=0.73
+ $X2=0 $Y2=0
cc_1045 N_A_229_491#_c_1770_n noxref_26 0.0018997f $X=3.865 $Y=0.77 $X2=-0.19
+ $Y2=-0.245
cc_1046 N_Q_c_1923_n N_VGND_c_1948_n 0.0315576f $X=13.18 $Y=0.46 $X2=0 $Y2=0
cc_1047 N_Q_c_1923_n N_VGND_c_1954_n 0.0147504f $X=13.18 $Y=0.46 $X2=0 $Y2=0
cc_1048 N_Q_c_1923_n N_VGND_c_1955_n 0.00983143f $X=13.18 $Y=0.46 $X2=0 $Y2=0
cc_1049 N_VGND_c_1949_n N_noxref_24_c_2073_n 0.0206518f $X=3.875 $Y=0 $X2=0
+ $Y2=0
cc_1050 N_VGND_c_1955_n N_noxref_24_c_2073_n 0.0122979f $X=13.2 $Y=0 $X2=0 $Y2=0
cc_1051 N_VGND_c_1944_n N_noxref_24_c_2074_n 0.0100109f $X=4.04 $Y=0.36 $X2=0
+ $Y2=0
cc_1052 N_VGND_c_1949_n N_noxref_24_c_2075_n 0.112255f $X=3.875 $Y=0 $X2=0 $Y2=0
cc_1053 N_VGND_c_1955_n N_noxref_24_c_2075_n 0.0673596f $X=13.2 $Y=0 $X2=0 $Y2=0
cc_1054 N_noxref_24_c_2075_n noxref_25 0.00310834f $X=3.22 $Y=0.39 $X2=-0.19
+ $Y2=-0.245
cc_1055 N_noxref_24_c_2075_n noxref_26 0.00193643f $X=3.22 $Y=0.39 $X2=-0.19
+ $Y2=-0.245
