* File: sky130_fd_sc_lp__a31o_lp.pxi.spice
* Created: Fri Aug 28 09:59:32 2020
* 
x_PM_SKY130_FD_SC_LP__A31O_LP%B1 N_B1_c_73_n N_B1_M1007_g N_B1_c_74_n
+ N_B1_M1003_g N_B1_M1005_g N_B1_c_76_n B1 N_B1_c_78_n
+ PM_SKY130_FD_SC_LP__A31O_LP%B1
x_PM_SKY130_FD_SC_LP__A31O_LP%A1 N_A1_M1008_g N_A1_M1009_g N_A1_c_113_n
+ N_A1_c_114_n A1 N_A1_c_116_n N_A1_c_117_n PM_SKY130_FD_SC_LP__A31O_LP%A1
x_PM_SKY130_FD_SC_LP__A31O_LP%A2 N_A2_M1004_g N_A2_M1010_g A2 A2 A2 N_A2_c_158_n
+ PM_SKY130_FD_SC_LP__A31O_LP%A2
x_PM_SKY130_FD_SC_LP__A31O_LP%A3 N_A3_M1011_g N_A3_M1000_g N_A3_c_201_n
+ N_A3_c_202_n A3 N_A3_c_204_n N_A3_c_205_n PM_SKY130_FD_SC_LP__A31O_LP%A3
x_PM_SKY130_FD_SC_LP__A31O_LP%A_48_409# N_A_48_409#_M1005_d N_A_48_409#_M1003_s
+ N_A_48_409#_c_243_n N_A_48_409#_M1001_g N_A_48_409#_c_244_n
+ N_A_48_409#_c_245_n N_A_48_409#_c_256_n N_A_48_409#_M1006_g
+ N_A_48_409#_c_246_n N_A_48_409#_M1002_g N_A_48_409#_c_247_n
+ N_A_48_409#_c_248_n N_A_48_409#_c_249_n N_A_48_409#_c_250_n
+ N_A_48_409#_c_260_n N_A_48_409#_c_251_n N_A_48_409#_c_252_n
+ N_A_48_409#_c_261_n N_A_48_409#_c_253_n N_A_48_409#_c_254_n
+ N_A_48_409#_c_255_n N_A_48_409#_c_262_n PM_SKY130_FD_SC_LP__A31O_LP%A_48_409#
x_PM_SKY130_FD_SC_LP__A31O_LP%A_155_409# N_A_155_409#_M1003_d
+ N_A_155_409#_M1004_d N_A_155_409#_c_346_n N_A_155_409#_c_347_n
+ N_A_155_409#_c_348_n N_A_155_409#_c_349_n N_A_155_409#_c_350_n
+ PM_SKY130_FD_SC_LP__A31O_LP%A_155_409#
x_PM_SKY130_FD_SC_LP__A31O_LP%VPWR N_VPWR_M1008_d N_VPWR_M1000_d N_VPWR_c_380_n
+ N_VPWR_c_381_n N_VPWR_c_382_n N_VPWR_c_383_n N_VPWR_c_384_n N_VPWR_c_385_n
+ VPWR N_VPWR_c_386_n N_VPWR_c_379_n PM_SKY130_FD_SC_LP__A31O_LP%VPWR
x_PM_SKY130_FD_SC_LP__A31O_LP%X N_X_M1002_d N_X_M1006_d N_X_c_424_n N_X_c_422_n
+ N_X_c_423_n X X PM_SKY130_FD_SC_LP__A31O_LP%X
x_PM_SKY130_FD_SC_LP__A31O_LP%VGND N_VGND_M1007_s N_VGND_M1011_d N_VGND_c_445_n
+ N_VGND_c_446_n N_VGND_c_447_n VGND N_VGND_c_448_n N_VGND_c_449_n
+ N_VGND_c_450_n N_VGND_c_451_n PM_SKY130_FD_SC_LP__A31O_LP%VGND
cc_1 VNB N_B1_c_73_n 0.0316597f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=0.775
cc_2 VNB N_B1_c_74_n 0.0311866f $X=-0.19 $Y=-0.245 $X2=0.602 $Y2=1.323
cc_3 VNB N_B1_M1003_g 0.0112721f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=2.545
cc_4 VNB N_B1_c_76_n 0.0208439f $X=-0.19 $Y=-0.245 $X2=0.685 $Y2=0.925
cc_5 VNB B1 0.00250885f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_6 VNB N_B1_c_78_n 0.0147006f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.33
cc_7 VNB N_A1_M1008_g 0.0104044f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=0.49
cc_8 VNB N_A1_c_113_n 0.0142635f $X=-0.19 $Y=-0.245 $X2=0.865 $Y2=0.775
cc_9 VNB N_A1_c_114_n 0.0121316f $X=-0.19 $Y=-0.245 $X2=0.865 $Y2=0.49
cc_10 VNB A1 0.00422591f $X=-0.19 $Y=-0.245 $X2=0.865 $Y2=0.49
cc_11 VNB N_A1_c_116_n 0.0247914f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_12 VNB N_A1_c_117_n 0.0135787f $X=-0.19 $Y=-0.245 $X2=0.602 $Y2=1.33
cc_13 VNB N_A2_M1004_g 0.0104044f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=0.49
cc_14 VNB N_A2_M1010_g 0.0300601f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=2.545
cc_15 VNB A2 0.00952977f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A2_c_158_n 0.0297569f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A3_M1000_g 0.0101269f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=2.545
cc_18 VNB N_A3_c_201_n 0.0142503f $X=-0.19 $Y=-0.245 $X2=0.865 $Y2=0.775
cc_19 VNB N_A3_c_202_n 0.0132262f $X=-0.19 $Y=-0.245 $X2=0.865 $Y2=0.49
cc_20 VNB A3 0.0047117f $X=-0.19 $Y=-0.245 $X2=0.865 $Y2=0.49
cc_21 VNB N_A3_c_204_n 0.0259984f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_22 VNB N_A3_c_205_n 0.0152708f $X=-0.19 $Y=-0.245 $X2=0.602 $Y2=1.33
cc_23 VNB N_A_48_409#_c_243_n 0.0136814f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=2.545
cc_24 VNB N_A_48_409#_c_244_n 0.00837341f $X=-0.19 $Y=-0.245 $X2=0.865 $Y2=0.775
cc_25 VNB N_A_48_409#_c_245_n 0.0132502f $X=-0.19 $Y=-0.245 $X2=0.865 $Y2=0.49
cc_26 VNB N_A_48_409#_c_246_n 0.0183435f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.33
cc_27 VNB N_A_48_409#_c_247_n 0.016434f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_48_409#_c_248_n 0.0239833f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.33
cc_29 VNB N_A_48_409#_c_249_n 0.00651266f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_48_409#_c_250_n 0.032413f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_48_409#_c_251_n 0.0150687f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_48_409#_c_252_n 0.00977235f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_48_409#_c_253_n 0.00207657f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_48_409#_c_254_n 0.00216019f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_48_409#_c_255_n 0.0146378f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VPWR_c_379_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_X_c_422_n 0.0448728f $X=-0.19 $Y=-0.245 $X2=0.865 $Y2=0.49
cc_38 VNB N_X_c_423_n 0.0266206f $X=-0.19 $Y=-0.245 $X2=0.685 $Y2=0.925
cc_39 VNB N_VGND_c_445_n 0.0116398f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=2.545
cc_40 VNB N_VGND_c_446_n 0.0187263f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_447_n 0.00544811f $X=-0.19 $Y=-0.245 $X2=0.685 $Y2=0.775
cc_42 VNB N_VGND_c_448_n 0.0464048f $X=-0.19 $Y=-0.245 $X2=0.602 $Y2=1.33
cc_43 VNB N_VGND_c_449_n 0.026935f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_450_n 0.215959f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_451_n 0.00494383f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VPB N_B1_M1003_g 0.0462088f $X=-0.19 $Y=1.655 $X2=0.65 $Y2=2.545
cc_47 VPB N_A1_M1008_g 0.0385385f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=0.49
cc_48 VPB N_A2_M1004_g 0.0385646f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=0.49
cc_49 VPB N_A3_M1000_g 0.0382145f $X=-0.19 $Y=1.655 $X2=0.65 $Y2=2.545
cc_50 VPB N_A_48_409#_c_256_n 0.0139187f $X=-0.19 $Y=1.655 $X2=0.865 $Y2=0.49
cc_51 VPB N_A_48_409#_M1006_g 0.0332163f $X=-0.19 $Y=1.655 $X2=0.685 $Y2=0.925
cc_52 VPB N_A_48_409#_c_248_n 0.00177884f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=1.33
cc_53 VPB N_A_48_409#_c_250_n 9.6636e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_54 VPB N_A_48_409#_c_260_n 0.057773f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_55 VPB N_A_48_409#_c_261_n 0.0397953f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_56 VPB N_A_48_409#_c_262_n 0.0158894f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_57 VPB N_A_155_409#_c_346_n 0.0025403f $X=-0.19 $Y=1.655 $X2=0.65 $Y2=2.545
cc_58 VPB N_A_155_409#_c_347_n 0.00207453f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_59 VPB N_A_155_409#_c_348_n 0.00248668f $X=-0.19 $Y=1.655 $X2=0.865 $Y2=0.49
cc_60 VPB N_A_155_409#_c_349_n 0.00254232f $X=-0.19 $Y=1.655 $X2=0.685 $Y2=0.775
cc_61 VPB N_A_155_409#_c_350_n 0.00207453f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_62 VPB N_VPWR_c_380_n 0.00177638f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_63 VPB N_VPWR_c_381_n 0.00426475f $X=-0.19 $Y=1.655 $X2=0.685 $Y2=0.775
cc_64 VPB N_VPWR_c_382_n 0.0349526f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=1.33
cc_65 VPB N_VPWR_c_383_n 0.00497896f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=1.33
cc_66 VPB N_VPWR_c_384_n 0.0187052f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=1.33
cc_67 VPB N_VPWR_c_385_n 0.00497896f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_386_n 0.019711f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_69 VPB N_VPWR_c_379_n 0.0538143f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_70 VPB N_X_c_424_n 0.0154157f $X=-0.19 $Y=1.655 $X2=0.865 $Y2=0.49
cc_71 VPB N_X_c_422_n 0.0177181f $X=-0.19 $Y=1.655 $X2=0.865 $Y2=0.49
cc_72 VPB X 0.0376238f $X=-0.19 $Y=1.655 $X2=0.602 $Y2=1.33
cc_73 N_B1_M1003_g N_A1_M1008_g 0.0340017f $X=0.65 $Y=2.545 $X2=0 $Y2=0
cc_74 N_B1_c_73_n N_A1_c_113_n 0.0111536f $X=0.505 $Y=0.775 $X2=0 $Y2=0
cc_75 N_B1_c_76_n N_A1_c_114_n 0.00894027f $X=0.685 $Y=0.925 $X2=0 $Y2=0
cc_76 N_B1_c_74_n A1 3.86417e-19 $X=0.602 $Y=1.323 $X2=0 $Y2=0
cc_77 B1 A1 0.0252734f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_78 N_B1_c_74_n N_A1_c_116_n 0.0214043f $X=0.602 $Y=1.323 $X2=0 $Y2=0
cc_79 B1 N_A1_c_116_n 0.0011114f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_80 N_B1_c_74_n N_A1_c_117_n 0.00891955f $X=0.602 $Y=1.323 $X2=0 $Y2=0
cc_81 N_B1_c_74_n N_A_48_409#_c_250_n 0.0143743f $X=0.602 $Y=1.323 $X2=0 $Y2=0
cc_82 N_B1_M1003_g N_A_48_409#_c_250_n 0.00590404f $X=0.65 $Y=2.545 $X2=0 $Y2=0
cc_83 B1 N_A_48_409#_c_250_n 0.0238428f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_84 N_B1_M1003_g N_A_48_409#_c_260_n 0.0263184f $X=0.65 $Y=2.545 $X2=0 $Y2=0
cc_85 N_B1_c_74_n N_A_48_409#_c_251_n 0.00924536f $X=0.602 $Y=1.323 $X2=0 $Y2=0
cc_86 N_B1_c_76_n N_A_48_409#_c_251_n 0.0219268f $X=0.685 $Y=0.925 $X2=0 $Y2=0
cc_87 B1 N_A_48_409#_c_251_n 0.0247946f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_88 N_B1_M1003_g N_A_48_409#_c_261_n 0.0178302f $X=0.65 $Y=2.545 $X2=0 $Y2=0
cc_89 B1 N_A_48_409#_c_261_n 0.0176002f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_90 N_B1_c_73_n N_A_48_409#_c_253_n 0.0115883f $X=0.505 $Y=0.775 $X2=0 $Y2=0
cc_91 N_B1_c_76_n N_A_48_409#_c_253_n 0.00221886f $X=0.685 $Y=0.925 $X2=0 $Y2=0
cc_92 N_B1_M1003_g N_A_48_409#_c_262_n 0.00448518f $X=0.65 $Y=2.545 $X2=0 $Y2=0
cc_93 B1 N_A_48_409#_c_262_n 0.00836812f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_94 N_B1_c_78_n N_A_48_409#_c_262_n 0.0028846f $X=0.61 $Y=1.33 $X2=0 $Y2=0
cc_95 N_B1_M1003_g N_A_155_409#_c_346_n 0.0036669f $X=0.65 $Y=2.545 $X2=0 $Y2=0
cc_96 N_B1_M1003_g N_A_155_409#_c_347_n 0.0156243f $X=0.65 $Y=2.545 $X2=0 $Y2=0
cc_97 N_B1_M1003_g N_VPWR_c_380_n 8.49223e-19 $X=0.65 $Y=2.545 $X2=0 $Y2=0
cc_98 N_B1_M1003_g N_VPWR_c_382_n 0.00826654f $X=0.65 $Y=2.545 $X2=0 $Y2=0
cc_99 N_B1_M1003_g N_VPWR_c_379_n 0.0156018f $X=0.65 $Y=2.545 $X2=0 $Y2=0
cc_100 N_B1_c_73_n N_VGND_c_446_n 0.0136008f $X=0.505 $Y=0.775 $X2=0 $Y2=0
cc_101 N_B1_c_73_n N_VGND_c_448_n 0.00956134f $X=0.505 $Y=0.775 $X2=0 $Y2=0
cc_102 N_B1_c_76_n N_VGND_c_448_n 5.88488e-19 $X=0.685 $Y=0.925 $X2=0 $Y2=0
cc_103 N_B1_c_73_n N_VGND_c_450_n 0.00985875f $X=0.505 $Y=0.775 $X2=0 $Y2=0
cc_104 N_B1_c_76_n N_VGND_c_450_n 7.97054e-19 $X=0.685 $Y=0.925 $X2=0 $Y2=0
cc_105 N_A1_M1008_g N_A2_M1004_g 0.0478604f $X=1.18 $Y=2.545 $X2=0 $Y2=0
cc_106 N_A1_c_113_n N_A2_M1010_g 0.0403402f $X=1.267 $Y=0.775 $X2=0 $Y2=0
cc_107 N_A1_c_117_n N_A2_M1010_g 0.00909965f $X=1.15 $Y=1.165 $X2=0 $Y2=0
cc_108 N_A1_c_113_n A2 0.00348756f $X=1.267 $Y=0.775 $X2=0 $Y2=0
cc_109 A1 A2 0.0208755f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_110 N_A1_c_116_n A2 4.14293e-19 $X=1.15 $Y=1.33 $X2=0 $Y2=0
cc_111 N_A1_c_117_n A2 0.0044757f $X=1.15 $Y=1.165 $X2=0 $Y2=0
cc_112 A1 N_A2_c_158_n 0.00114406f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_113 N_A1_c_116_n N_A2_c_158_n 0.0207808f $X=1.15 $Y=1.33 $X2=0 $Y2=0
cc_114 N_A1_M1008_g N_A_48_409#_c_260_n 0.00104556f $X=1.18 $Y=2.545 $X2=0 $Y2=0
cc_115 N_A1_c_114_n N_A_48_409#_c_251_n 0.0030188f $X=1.267 $Y=0.925 $X2=0 $Y2=0
cc_116 A1 N_A_48_409#_c_251_n 0.020736f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_117 N_A1_c_116_n N_A_48_409#_c_251_n 0.00460175f $X=1.15 $Y=1.33 $X2=0 $Y2=0
cc_118 N_A1_c_117_n N_A_48_409#_c_251_n 0.00304073f $X=1.15 $Y=1.165 $X2=0 $Y2=0
cc_119 N_A1_M1008_g N_A_48_409#_c_261_n 0.0149541f $X=1.18 $Y=2.545 $X2=0 $Y2=0
cc_120 A1 N_A_48_409#_c_261_n 0.0228124f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_121 N_A1_c_116_n N_A_48_409#_c_261_n 0.0018211f $X=1.15 $Y=1.33 $X2=0 $Y2=0
cc_122 N_A1_c_113_n N_A_48_409#_c_253_n 0.0088623f $X=1.267 $Y=0.775 $X2=0 $Y2=0
cc_123 N_A1_c_114_n N_A_48_409#_c_253_n 0.00231191f $X=1.267 $Y=0.925 $X2=0
+ $Y2=0
cc_124 N_A1_M1008_g N_A_155_409#_c_346_n 9.82838e-19 $X=1.18 $Y=2.545 $X2=0
+ $Y2=0
cc_125 N_A1_M1008_g N_A_155_409#_c_347_n 0.0155966f $X=1.18 $Y=2.545 $X2=0 $Y2=0
cc_126 N_A1_M1008_g N_A_155_409#_c_348_n 0.0178604f $X=1.18 $Y=2.545 $X2=0 $Y2=0
cc_127 N_A1_M1008_g N_A_155_409#_c_350_n 8.93705e-19 $X=1.18 $Y=2.545 $X2=0
+ $Y2=0
cc_128 N_A1_M1008_g N_VPWR_c_380_n 0.0163548f $X=1.18 $Y=2.545 $X2=0 $Y2=0
cc_129 N_A1_M1008_g N_VPWR_c_382_n 0.00769046f $X=1.18 $Y=2.545 $X2=0 $Y2=0
cc_130 N_A1_M1008_g N_VPWR_c_379_n 0.0134474f $X=1.18 $Y=2.545 $X2=0 $Y2=0
cc_131 N_A1_c_113_n N_VGND_c_448_n 0.0050714f $X=1.267 $Y=0.775 $X2=0 $Y2=0
cc_132 N_A1_c_113_n N_VGND_c_450_n 0.00955779f $X=1.267 $Y=0.775 $X2=0 $Y2=0
cc_133 N_A2_M1004_g N_A3_M1000_g 0.0347392f $X=1.71 $Y=2.545 $X2=0 $Y2=0
cc_134 N_A2_M1010_g N_A3_c_201_n 0.0402302f $X=1.685 $Y=0.49 $X2=0 $Y2=0
cc_135 A2 N_A3_c_201_n 0.00691585f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_136 A2 A3 0.0240992f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_137 N_A2_c_158_n A3 0.00187621f $X=1.69 $Y=1.33 $X2=0 $Y2=0
cc_138 A2 N_A3_c_204_n 3.96006e-19 $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_139 N_A2_c_158_n N_A3_c_204_n 0.0207134f $X=1.69 $Y=1.33 $X2=0 $Y2=0
cc_140 N_A2_M1010_g N_A3_c_205_n 0.00869912f $X=1.685 $Y=0.49 $X2=0 $Y2=0
cc_141 A2 N_A3_c_205_n 0.00543735f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_142 A2 N_A_48_409#_c_251_n 0.00977888f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_143 N_A2_M1004_g N_A_48_409#_c_261_n 0.0149439f $X=1.71 $Y=2.545 $X2=0 $Y2=0
cc_144 A2 N_A_48_409#_c_261_n 0.0241538f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_145 N_A2_c_158_n N_A_48_409#_c_261_n 5.43058e-19 $X=1.69 $Y=1.33 $X2=0 $Y2=0
cc_146 N_A2_M1010_g N_A_48_409#_c_253_n 0.00121905f $X=1.685 $Y=0.49 $X2=0 $Y2=0
cc_147 A2 N_A_48_409#_c_253_n 0.0199941f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_148 N_A2_M1004_g N_A_155_409#_c_347_n 8.93705e-19 $X=1.71 $Y=2.545 $X2=0
+ $Y2=0
cc_149 N_A2_M1004_g N_A_155_409#_c_348_n 0.0178604f $X=1.71 $Y=2.545 $X2=0 $Y2=0
cc_150 N_A2_M1004_g N_A_155_409#_c_349_n 9.82838e-19 $X=1.71 $Y=2.545 $X2=0
+ $Y2=0
cc_151 N_A2_M1004_g N_A_155_409#_c_350_n 0.0155966f $X=1.71 $Y=2.545 $X2=0 $Y2=0
cc_152 N_A2_M1004_g N_VPWR_c_380_n 0.0163548f $X=1.71 $Y=2.545 $X2=0 $Y2=0
cc_153 N_A2_M1004_g N_VPWR_c_381_n 9.45181e-19 $X=1.71 $Y=2.545 $X2=0 $Y2=0
cc_154 N_A2_M1004_g N_VPWR_c_384_n 0.00769046f $X=1.71 $Y=2.545 $X2=0 $Y2=0
cc_155 N_A2_M1004_g N_VPWR_c_379_n 0.0134474f $X=1.71 $Y=2.545 $X2=0 $Y2=0
cc_156 N_A2_M1010_g N_VGND_c_447_n 0.00199711f $X=1.685 $Y=0.49 $X2=0 $Y2=0
cc_157 A2 N_VGND_c_447_n 0.015278f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_158 N_A2_M1010_g N_VGND_c_448_n 0.00360502f $X=1.685 $Y=0.49 $X2=0 $Y2=0
cc_159 A2 N_VGND_c_448_n 0.00846271f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_160 N_A2_M1010_g N_VGND_c_450_n 0.00499696f $X=1.685 $Y=0.49 $X2=0 $Y2=0
cc_161 A2 N_VGND_c_450_n 0.0106888f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_162 A2 A_274_56# 0.00307888f $X=1.595 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_163 A2 A_352_56# 0.00316748f $X=1.595 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_164 N_A3_c_201_n N_A_48_409#_c_243_n 0.0106476f $X=2.107 $Y=0.775 $X2=0 $Y2=0
cc_165 N_A3_c_202_n N_A_48_409#_c_245_n 0.0104671f $X=2.107 $Y=0.925 $X2=0 $Y2=0
cc_166 N_A3_M1000_g N_A_48_409#_M1006_g 0.0166396f $X=2.24 $Y=2.545 $X2=0 $Y2=0
cc_167 N_A3_c_204_n N_A_48_409#_c_247_n 2.7174e-19 $X=2.23 $Y=1.33 $X2=0 $Y2=0
cc_168 N_A3_c_205_n N_A_48_409#_c_247_n 0.0063149f $X=2.23 $Y=1.165 $X2=0 $Y2=0
cc_169 N_A3_M1000_g N_A_48_409#_c_248_n 0.0196833f $X=2.24 $Y=2.545 $X2=0 $Y2=0
cc_170 N_A3_M1000_g N_A_48_409#_c_261_n 0.0207577f $X=2.24 $Y=2.545 $X2=0 $Y2=0
cc_171 A3 N_A_48_409#_c_261_n 0.0243355f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_172 N_A3_c_204_n N_A_48_409#_c_261_n 0.00197701f $X=2.23 $Y=1.33 $X2=0 $Y2=0
cc_173 N_A3_M1000_g N_A_48_409#_c_254_n 0.00121683f $X=2.24 $Y=2.545 $X2=0 $Y2=0
cc_174 A3 N_A_48_409#_c_254_n 0.0202904f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_175 N_A3_c_204_n N_A_48_409#_c_254_n 4.02529e-19 $X=2.23 $Y=1.33 $X2=0 $Y2=0
cc_176 A3 N_A_48_409#_c_255_n 0.00110952f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_177 N_A3_c_204_n N_A_48_409#_c_255_n 0.0201099f $X=2.23 $Y=1.33 $X2=0 $Y2=0
cc_178 N_A3_M1000_g N_A_155_409#_c_349_n 0.00353403f $X=2.24 $Y=2.545 $X2=0
+ $Y2=0
cc_179 N_A3_M1000_g N_A_155_409#_c_350_n 0.0149653f $X=2.24 $Y=2.545 $X2=0 $Y2=0
cc_180 N_A3_M1000_g N_VPWR_c_380_n 8.49223e-19 $X=2.24 $Y=2.545 $X2=0 $Y2=0
cc_181 N_A3_M1000_g N_VPWR_c_381_n 0.0224497f $X=2.24 $Y=2.545 $X2=0 $Y2=0
cc_182 N_A3_M1000_g N_VPWR_c_384_n 0.00769046f $X=2.24 $Y=2.545 $X2=0 $Y2=0
cc_183 N_A3_M1000_g N_VPWR_c_379_n 0.0134474f $X=2.24 $Y=2.545 $X2=0 $Y2=0
cc_184 N_A3_M1000_g N_X_c_424_n 2.7744e-19 $X=2.24 $Y=2.545 $X2=0 $Y2=0
cc_185 N_A3_c_201_n N_VGND_c_447_n 0.0120945f $X=2.107 $Y=0.775 $X2=0 $Y2=0
cc_186 N_A3_c_202_n N_VGND_c_447_n 0.00236517f $X=2.107 $Y=0.925 $X2=0 $Y2=0
cc_187 A3 N_VGND_c_447_n 0.0109499f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_188 N_A3_c_204_n N_VGND_c_447_n 0.0039577f $X=2.23 $Y=1.33 $X2=0 $Y2=0
cc_189 N_A3_c_201_n N_VGND_c_448_n 0.00448994f $X=2.107 $Y=0.775 $X2=0 $Y2=0
cc_190 N_A3_c_201_n N_VGND_c_450_n 0.00806915f $X=2.107 $Y=0.775 $X2=0 $Y2=0
cc_191 N_A_48_409#_c_260_n N_A_155_409#_c_346_n 0.0121893f $X=0.385 $Y=2.19
+ $X2=0 $Y2=0
cc_192 N_A_48_409#_c_261_n N_A_155_409#_c_346_n 0.0263465f $X=2.605 $Y=1.76
+ $X2=0 $Y2=0
cc_193 N_A_48_409#_c_260_n N_A_155_409#_c_347_n 0.0587354f $X=0.385 $Y=2.19
+ $X2=0 $Y2=0
cc_194 N_A_48_409#_c_261_n N_A_155_409#_c_348_n 0.0493217f $X=2.605 $Y=1.76
+ $X2=0 $Y2=0
cc_195 N_A_48_409#_c_261_n N_A_155_409#_c_349_n 0.0263465f $X=2.605 $Y=1.76
+ $X2=0 $Y2=0
cc_196 N_A_48_409#_M1006_g N_A_155_409#_c_350_n 2.28436e-19 $X=2.77 $Y=2.545
+ $X2=0 $Y2=0
cc_197 N_A_48_409#_c_256_n N_VPWR_c_381_n 3.10915e-19 $X=2.77 $Y=1.845 $X2=0
+ $Y2=0
cc_198 N_A_48_409#_M1006_g N_VPWR_c_381_n 0.0237294f $X=2.77 $Y=2.545 $X2=0
+ $Y2=0
cc_199 N_A_48_409#_c_261_n N_VPWR_c_381_n 0.0265231f $X=2.605 $Y=1.76 $X2=0
+ $Y2=0
cc_200 N_A_48_409#_c_260_n N_VPWR_c_382_n 0.0304602f $X=0.385 $Y=2.19 $X2=0
+ $Y2=0
cc_201 N_A_48_409#_M1006_g N_VPWR_c_386_n 0.00769046f $X=2.77 $Y=2.545 $X2=0
+ $Y2=0
cc_202 N_A_48_409#_M1006_g N_VPWR_c_379_n 0.014111f $X=2.77 $Y=2.545 $X2=0 $Y2=0
cc_203 N_A_48_409#_c_260_n N_VPWR_c_379_n 0.0174175f $X=0.385 $Y=2.19 $X2=0
+ $Y2=0
cc_204 N_A_48_409#_c_256_n N_X_c_424_n 9.121e-19 $X=2.77 $Y=1.845 $X2=0 $Y2=0
cc_205 N_A_48_409#_M1006_g N_X_c_424_n 0.00413513f $X=2.77 $Y=2.545 $X2=0 $Y2=0
cc_206 N_A_48_409#_c_261_n N_X_c_424_n 0.00406923f $X=2.605 $Y=1.76 $X2=0 $Y2=0
cc_207 N_A_48_409#_M1006_g N_X_c_422_n 0.00452922f $X=2.77 $Y=2.545 $X2=0 $Y2=0
cc_208 N_A_48_409#_c_246_n N_X_c_422_n 0.00617237f $X=2.865 $Y=0.775 $X2=0 $Y2=0
cc_209 N_A_48_409#_c_247_n N_X_c_422_n 0.0237191f $X=2.77 $Y=1.175 $X2=0 $Y2=0
cc_210 N_A_48_409#_c_261_n N_X_c_422_n 0.0129671f $X=2.605 $Y=1.76 $X2=0 $Y2=0
cc_211 N_A_48_409#_c_254_n N_X_c_422_n 0.035795f $X=2.77 $Y=1.34 $X2=0 $Y2=0
cc_212 N_A_48_409#_c_243_n N_X_c_423_n 0.00123773f $X=2.505 $Y=0.775 $X2=0 $Y2=0
cc_213 N_A_48_409#_c_246_n N_X_c_423_n 0.00993775f $X=2.865 $Y=0.775 $X2=0 $Y2=0
cc_214 N_A_48_409#_M1006_g X 0.0147448f $X=2.77 $Y=2.545 $X2=0 $Y2=0
cc_215 N_A_48_409#_c_251_n N_VGND_c_446_n 0.0119264f $X=0.915 $Y=0.9 $X2=0 $Y2=0
cc_216 N_A_48_409#_c_252_n N_VGND_c_446_n 0.0119494f $X=0.265 $Y=0.9 $X2=0 $Y2=0
cc_217 N_A_48_409#_c_253_n N_VGND_c_446_n 0.0123792f $X=1.08 $Y=0.49 $X2=0 $Y2=0
cc_218 N_A_48_409#_c_243_n N_VGND_c_447_n 0.0133015f $X=2.505 $Y=0.775 $X2=0
+ $Y2=0
cc_219 N_A_48_409#_c_246_n N_VGND_c_447_n 0.0021406f $X=2.865 $Y=0.775 $X2=0
+ $Y2=0
cc_220 N_A_48_409#_c_253_n N_VGND_c_448_n 0.0220438f $X=1.08 $Y=0.49 $X2=0 $Y2=0
cc_221 N_A_48_409#_c_243_n N_VGND_c_449_n 0.00448994f $X=2.505 $Y=0.775 $X2=0
+ $Y2=0
cc_222 N_A_48_409#_c_244_n N_VGND_c_449_n 4.60722e-19 $X=2.785 $Y=0.85 $X2=0
+ $Y2=0
cc_223 N_A_48_409#_c_246_n N_VGND_c_449_n 0.0050714f $X=2.865 $Y=0.775 $X2=0
+ $Y2=0
cc_224 N_A_48_409#_c_243_n N_VGND_c_450_n 0.00798122f $X=2.505 $Y=0.775 $X2=0
+ $Y2=0
cc_225 N_A_48_409#_c_244_n N_VGND_c_450_n 6.34959e-19 $X=2.785 $Y=0.85 $X2=0
+ $Y2=0
cc_226 N_A_48_409#_c_246_n N_VGND_c_450_n 0.0101463f $X=2.865 $Y=0.775 $X2=0
+ $Y2=0
cc_227 N_A_48_409#_c_251_n N_VGND_c_450_n 0.0143823f $X=0.915 $Y=0.9 $X2=0 $Y2=0
cc_228 N_A_48_409#_c_252_n N_VGND_c_450_n 0.00178946f $X=0.265 $Y=0.9 $X2=0
+ $Y2=0
cc_229 N_A_48_409#_c_253_n N_VGND_c_450_n 0.0124902f $X=1.08 $Y=0.49 $X2=0 $Y2=0
cc_230 N_A_155_409#_c_348_n N_VPWR_M1008_d 0.00180746f $X=1.81 $Y=2.11 $X2=-0.19
+ $Y2=1.655
cc_231 N_A_155_409#_c_347_n N_VPWR_c_380_n 0.0454646f $X=0.915 $Y=2.9 $X2=0
+ $Y2=0
cc_232 N_A_155_409#_c_348_n N_VPWR_c_380_n 0.0163515f $X=1.81 $Y=2.11 $X2=0
+ $Y2=0
cc_233 N_A_155_409#_c_350_n N_VPWR_c_380_n 0.0454646f $X=1.975 $Y=2.9 $X2=0
+ $Y2=0
cc_234 N_A_155_409#_c_349_n N_VPWR_c_381_n 0.0119061f $X=1.975 $Y=2.195 $X2=0
+ $Y2=0
cc_235 N_A_155_409#_c_350_n N_VPWR_c_381_n 0.0572919f $X=1.975 $Y=2.9 $X2=0
+ $Y2=0
cc_236 N_A_155_409#_c_347_n N_VPWR_c_382_n 0.021949f $X=0.915 $Y=2.9 $X2=0 $Y2=0
cc_237 N_A_155_409#_c_350_n N_VPWR_c_384_n 0.021949f $X=1.975 $Y=2.9 $X2=0 $Y2=0
cc_238 N_A_155_409#_c_347_n N_VPWR_c_379_n 0.0124703f $X=0.915 $Y=2.9 $X2=0
+ $Y2=0
cc_239 N_A_155_409#_c_350_n N_VPWR_c_379_n 0.0124703f $X=1.975 $Y=2.9 $X2=0
+ $Y2=0
cc_240 N_VPWR_c_381_n N_X_c_424_n 0.0695159f $X=2.505 $Y=2.19 $X2=0 $Y2=0
cc_241 N_VPWR_c_386_n X 0.0267518f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_242 N_VPWR_c_379_n X 0.0152893f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_243 N_X_c_423_n N_VGND_c_447_n 0.0153087f $X=3.08 $Y=0.49 $X2=0 $Y2=0
cc_244 N_X_c_423_n N_VGND_c_449_n 0.0233562f $X=3.08 $Y=0.49 $X2=0 $Y2=0
cc_245 N_X_c_423_n N_VGND_c_450_n 0.0134729f $X=3.08 $Y=0.49 $X2=0 $Y2=0
