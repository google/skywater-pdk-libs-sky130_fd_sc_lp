* File: sky130_fd_sc_lp__nand4_1.pxi.spice
* Created: Wed Sep  2 10:05:28 2020
* 
x_PM_SKY130_FD_SC_LP__NAND4_1%D N_D_M1007_g N_D_M1004_g D D N_D_c_43_n
+ N_D_c_44_n PM_SKY130_FD_SC_LP__NAND4_1%D
x_PM_SKY130_FD_SC_LP__NAND4_1%C N_C_M1003_g N_C_M1001_g C C C N_C_c_68_n
+ N_C_c_69_n PM_SKY130_FD_SC_LP__NAND4_1%C
x_PM_SKY130_FD_SC_LP__NAND4_1%B N_B_M1000_g N_B_M1002_g B B B N_B_c_99_n
+ N_B_c_100_n PM_SKY130_FD_SC_LP__NAND4_1%B
x_PM_SKY130_FD_SC_LP__NAND4_1%A N_A_M1006_g N_A_M1005_g A A A N_A_c_131_n
+ N_A_c_132_n PM_SKY130_FD_SC_LP__NAND4_1%A
x_PM_SKY130_FD_SC_LP__NAND4_1%VPWR N_VPWR_M1004_s N_VPWR_M1001_d N_VPWR_M1005_d
+ N_VPWR_c_161_n N_VPWR_c_162_n N_VPWR_c_163_n N_VPWR_c_164_n N_VPWR_c_165_n
+ N_VPWR_c_166_n VPWR N_VPWR_c_167_n N_VPWR_c_168_n N_VPWR_c_160_n
+ PM_SKY130_FD_SC_LP__NAND4_1%VPWR
x_PM_SKY130_FD_SC_LP__NAND4_1%Y N_Y_M1006_d N_Y_M1004_d N_Y_M1002_d N_Y_c_197_n
+ N_Y_c_196_n Y Y Y Y N_Y_c_201_n N_Y_c_204_n N_Y_c_223_n
+ PM_SKY130_FD_SC_LP__NAND4_1%Y
x_PM_SKY130_FD_SC_LP__NAND4_1%VGND N_VGND_M1007_s N_VGND_c_239_n N_VGND_c_240_n
+ VGND N_VGND_c_241_n N_VGND_c_242_n PM_SKY130_FD_SC_LP__NAND4_1%VGND
cc_1 VNB N_D_M1004_g 0.0114223f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=2.465
cc_2 VNB D 0.026642f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_3 VNB N_D_c_43_n 0.0405089f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=1.35
cc_4 VNB N_D_c_44_n 0.0219223f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=1.185
cc_5 VNB N_C_M1001_g 0.00863754f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=2.465
cc_6 VNB C 0.00515365f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_7 VNB N_C_c_68_n 0.0315099f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=1.185
cc_8 VNB N_C_c_69_n 0.0167966f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.322
cc_9 VNB N_B_M1002_g 0.00863754f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=2.465
cc_10 VNB B 0.00149014f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_11 VNB N_B_c_99_n 0.0342509f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=1.185
cc_12 VNB N_B_c_100_n 0.0182897f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.322
cc_13 VNB N_A_M1005_g 0.00821138f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=2.465
cc_14 VNB A 0.00208946f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_15 VNB N_A_c_131_n 0.0370097f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=1.185
cc_16 VNB N_A_c_132_n 0.0213919f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.322
cc_17 VNB N_VPWR_c_160_n 0.123877f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_Y_c_196_n 0.0291024f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=1.35
cc_19 VNB N_VGND_c_239_n 0.0148529f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.515
cc_20 VNB N_VGND_c_240_n 0.00495479f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=2.465
cc_21 VNB N_VGND_c_241_n 0.072646f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=1.185
cc_22 VNB N_VGND_c_242_n 0.177751f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=1.515
cc_23 VPB N_D_M1004_g 0.0276728f $X=-0.19 $Y=1.655 $X2=0.59 $Y2=2.465
cc_24 VPB N_C_M1001_g 0.0219347f $X=-0.19 $Y=1.655 $X2=0.59 $Y2=2.465
cc_25 VPB N_B_M1002_g 0.0219347f $X=-0.19 $Y=1.655 $X2=0.59 $Y2=2.465
cc_26 VPB N_A_M1005_g 0.0238458f $X=-0.19 $Y=1.655 $X2=0.59 $Y2=2.465
cc_27 VPB N_VPWR_c_161_n 0.0140295f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_28 VPB N_VPWR_c_162_n 0.00444763f $X=-0.19 $Y=1.655 $X2=0.5 $Y2=1.35
cc_29 VPB N_VPWR_c_163_n 0.0198439f $X=-0.19 $Y=1.655 $X2=0.5 $Y2=1.515
cc_30 VPB N_VPWR_c_164_n 0.00443752f $X=-0.19 $Y=1.655 $X2=0.5 $Y2=1.322
cc_31 VPB N_VPWR_c_165_n 0.0140295f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_32 VPB N_VPWR_c_166_n 0.00496839f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_33 VPB N_VPWR_c_167_n 0.0319119f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_34 VPB N_VPWR_c_168_n 0.00401341f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_35 VPB N_VPWR_c_160_n 0.0541716f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_36 VPB N_Y_c_197_n 0.0136692f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_37 VPB N_Y_c_196_n 0.00531653f $X=-0.19 $Y=1.655 $X2=0.5 $Y2=1.35
cc_38 VPB Y 0.00581932f $X=-0.19 $Y=1.655 $X2=0.5 $Y2=1.515
cc_39 VPB Y 0.0101897f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_40 VPB N_Y_c_201_n 0.0112475f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_41 N_D_M1004_g N_C_M1001_g 0.0324001f $X=0.59 $Y=2.465 $X2=0 $Y2=0
cc_42 D C 0.0178279f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_43 N_D_c_43_n C 6.69494e-19 $X=0.5 $Y=1.35 $X2=0 $Y2=0
cc_44 N_D_c_44_n C 0.0030809f $X=0.5 $Y=1.185 $X2=0 $Y2=0
cc_45 D N_C_c_68_n 0.00170116f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_46 N_D_c_43_n N_C_c_68_n 0.0372643f $X=0.5 $Y=1.35 $X2=0 $Y2=0
cc_47 N_D_c_44_n N_C_c_69_n 0.0372643f $X=0.5 $Y=1.185 $X2=0 $Y2=0
cc_48 N_D_M1004_g N_VPWR_c_162_n 0.0077802f $X=0.59 $Y=2.465 $X2=0 $Y2=0
cc_49 D N_VPWR_c_162_n 0.00599389f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_50 N_D_c_43_n N_VPWR_c_162_n 0.00213837f $X=0.5 $Y=1.35 $X2=0 $Y2=0
cc_51 N_D_M1004_g N_VPWR_c_163_n 0.00550419f $X=0.59 $Y=2.465 $X2=0 $Y2=0
cc_52 N_D_M1004_g N_VPWR_c_160_n 0.0108033f $X=0.59 $Y=2.465 $X2=0 $Y2=0
cc_53 N_D_M1004_g Y 0.0183305f $X=0.59 $Y=2.465 $X2=0 $Y2=0
cc_54 D Y 0.00916503f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_55 N_D_M1004_g N_Y_c_204_n 0.00844436f $X=0.59 $Y=2.465 $X2=0 $Y2=0
cc_56 D N_VGND_c_240_n 0.00985004f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_57 N_D_c_43_n N_VGND_c_240_n 0.00306495f $X=0.5 $Y=1.35 $X2=0 $Y2=0
cc_58 N_D_c_44_n N_VGND_c_240_n 0.00460896f $X=0.5 $Y=1.185 $X2=0 $Y2=0
cc_59 N_D_c_44_n N_VGND_c_241_n 0.00585385f $X=0.5 $Y=1.185 $X2=0 $Y2=0
cc_60 N_D_c_44_n N_VGND_c_242_n 0.011642f $X=0.5 $Y=1.185 $X2=0 $Y2=0
cc_61 N_C_M1001_g N_B_M1002_g 0.0304488f $X=1.02 $Y=2.465 $X2=0 $Y2=0
cc_62 C B 0.055344f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_63 N_C_c_68_n B 3.46554e-19 $X=1.07 $Y=1.35 $X2=0 $Y2=0
cc_64 N_C_c_69_n B 6.12644e-19 $X=1.07 $Y=1.185 $X2=0 $Y2=0
cc_65 N_C_c_68_n N_B_c_99_n 0.0174484f $X=1.07 $Y=1.35 $X2=0 $Y2=0
cc_66 C N_B_c_100_n 0.00819668f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_67 N_C_c_69_n N_B_c_100_n 0.0286456f $X=1.07 $Y=1.185 $X2=0 $Y2=0
cc_68 N_C_M1001_g N_VPWR_c_163_n 0.00585385f $X=1.02 $Y=2.465 $X2=0 $Y2=0
cc_69 N_C_M1001_g N_VPWR_c_164_n 0.00192941f $X=1.02 $Y=2.465 $X2=0 $Y2=0
cc_70 N_C_M1001_g N_VPWR_c_160_n 0.0112235f $X=1.02 $Y=2.465 $X2=0 $Y2=0
cc_71 N_C_c_68_n Y 2.24402e-19 $X=1.07 $Y=1.35 $X2=0 $Y2=0
cc_72 N_C_M1001_g N_Y_c_201_n 0.0235573f $X=1.02 $Y=2.465 $X2=0 $Y2=0
cc_73 C N_Y_c_201_n 0.0192072f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_74 N_C_c_68_n N_Y_c_201_n 0.00242458f $X=1.07 $Y=1.35 $X2=0 $Y2=0
cc_75 C N_VGND_c_241_n 0.00774939f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_76 N_C_c_69_n N_VGND_c_241_n 0.00499463f $X=1.07 $Y=1.185 $X2=0 $Y2=0
cc_77 C N_VGND_c_242_n 0.00983356f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_78 N_C_c_69_n N_VGND_c_242_n 0.00880207f $X=1.07 $Y=1.185 $X2=0 $Y2=0
cc_79 C A_211_47# 0.0102108f $X=1.115 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_80 N_B_M1002_g N_A_M1005_g 0.0337732f $X=1.69 $Y=2.465 $X2=0 $Y2=0
cc_81 B A 0.0473044f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_82 N_B_c_99_n A 0.00119094f $X=1.64 $Y=1.35 $X2=0 $Y2=0
cc_83 N_B_c_100_n A 7.29939e-19 $X=1.64 $Y=1.185 $X2=0 $Y2=0
cc_84 B N_A_c_131_n 0.00116585f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_85 N_B_c_99_n N_A_c_131_n 0.0173376f $X=1.64 $Y=1.35 $X2=0 $Y2=0
cc_86 B N_A_c_132_n 0.00506533f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_87 N_B_c_100_n N_A_c_132_n 0.0290479f $X=1.64 $Y=1.185 $X2=0 $Y2=0
cc_88 N_B_M1002_g N_VPWR_c_164_n 0.0110755f $X=1.69 $Y=2.465 $X2=0 $Y2=0
cc_89 N_B_M1002_g N_VPWR_c_167_n 0.00585385f $X=1.69 $Y=2.465 $X2=0 $Y2=0
cc_90 N_B_M1002_g N_VPWR_c_160_n 0.0115441f $X=1.69 $Y=2.465 $X2=0 $Y2=0
cc_91 N_B_c_99_n Y 2.0611e-19 $X=1.64 $Y=1.35 $X2=0 $Y2=0
cc_92 N_B_M1002_g N_Y_c_201_n 0.0222552f $X=1.69 $Y=2.465 $X2=0 $Y2=0
cc_93 B N_Y_c_201_n 0.0129325f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_94 N_B_c_99_n N_Y_c_201_n 0.0050893f $X=1.64 $Y=1.35 $X2=0 $Y2=0
cc_95 B N_VGND_c_241_n 0.00514572f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_96 N_B_c_100_n N_VGND_c_241_n 0.00499463f $X=1.64 $Y=1.185 $X2=0 $Y2=0
cc_97 B N_VGND_c_242_n 0.00675903f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_98 N_B_c_100_n N_VGND_c_242_n 0.00923391f $X=1.64 $Y=1.185 $X2=0 $Y2=0
cc_99 B A_325_47# 0.0080065f $X=1.595 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_100 N_A_M1005_g N_VPWR_c_166_n 0.0165554f $X=2.12 $Y=2.465 $X2=0 $Y2=0
cc_101 N_A_M1005_g N_VPWR_c_167_n 0.00404527f $X=2.12 $Y=2.465 $X2=0 $Y2=0
cc_102 N_A_M1005_g N_VPWR_c_160_n 0.00695434f $X=2.12 $Y=2.465 $X2=0 $Y2=0
cc_103 A N_Y_M1006_d 0.00726786f $X=2.075 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_104 A N_Y_c_197_n 0.00298883f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_105 N_A_c_131_n N_Y_c_197_n 0.00314108f $X=2.21 $Y=1.35 $X2=0 $Y2=0
cc_106 N_A_M1005_g N_Y_c_196_n 0.00745766f $X=2.12 $Y=2.465 $X2=0 $Y2=0
cc_107 A N_Y_c_196_n 0.0752955f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_108 N_A_c_131_n N_Y_c_196_n 0.00812569f $X=2.21 $Y=1.35 $X2=0 $Y2=0
cc_109 N_A_c_132_n N_Y_c_196_n 0.00539828f $X=2.21 $Y=1.185 $X2=0 $Y2=0
cc_110 N_A_M1005_g Y 0.0164738f $X=2.12 $Y=2.465 $X2=0 $Y2=0
cc_111 A Y 0.0110636f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_112 N_A_c_131_n Y 3.79428e-19 $X=2.21 $Y=1.35 $X2=0 $Y2=0
cc_113 N_A_M1005_g N_Y_c_223_n 0.0232165f $X=2.12 $Y=2.465 $X2=0 $Y2=0
cc_114 A N_VGND_c_241_n 0.00535903f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_115 N_A_c_132_n N_VGND_c_241_n 0.00437201f $X=2.21 $Y=1.185 $X2=0 $Y2=0
cc_116 A N_VGND_c_242_n 0.00684951f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_117 N_A_c_132_n N_VGND_c_242_n 0.0083083f $X=2.21 $Y=1.185 $X2=0 $Y2=0
cc_118 N_VPWR_c_160_n N_Y_M1004_d 0.003948f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_119 N_VPWR_c_160_n N_Y_M1002_d 0.003948f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_120 N_VPWR_M1005_d N_Y_c_197_n 0.0112961f $X=2.195 $Y=1.835 $X2=0 $Y2=0
cc_121 N_VPWR_c_166_n N_Y_c_197_n 0.0175169f $X=2.53 $Y=2.27 $X2=0 $Y2=0
cc_122 N_VPWR_c_162_n Y 0.00114446f $X=0.35 $Y=2.27 $X2=0 $Y2=0
cc_123 N_VPWR_M1001_d N_Y_c_201_n 0.0144361f $X=1.095 $Y=1.835 $X2=0 $Y2=0
cc_124 N_VPWR_c_164_n N_Y_c_201_n 0.00994109f $X=1.235 $Y=2.61 $X2=0 $Y2=0
cc_125 N_VPWR_c_162_n N_Y_c_204_n 0.0498626f $X=0.35 $Y=2.27 $X2=0 $Y2=0
cc_126 N_VPWR_c_163_n N_Y_c_204_n 0.00616009f $X=1.13 $Y=3.33 $X2=0 $Y2=0
cc_127 N_VPWR_c_160_n N_Y_c_204_n 0.00894104f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_128 N_VPWR_c_167_n N_Y_c_223_n 0.00984606f $X=2.425 $Y=3.33 $X2=0 $Y2=0
cc_129 N_VPWR_c_160_n N_Y_c_223_n 0.0139961f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_130 N_Y_c_196_n N_VGND_c_241_n 0.00689397f $X=2.58 $Y=0.59 $X2=0 $Y2=0
cc_131 N_Y_M1006_d N_VGND_c_242_n 0.0116079f $X=2.195 $Y=0.235 $X2=0 $Y2=0
cc_132 N_Y_c_196_n N_VGND_c_242_n 0.00732528f $X=2.58 $Y=0.59 $X2=0 $Y2=0
cc_133 N_VGND_c_242_n A_133_47# 0.010279f $X=2.64 $Y=0 $X2=-0.19 $Y2=-0.245
cc_134 N_VGND_c_242_n A_211_47# 0.0103644f $X=2.64 $Y=0 $X2=-0.19 $Y2=-0.245
cc_135 N_VGND_c_242_n A_325_47# 0.0133686f $X=2.64 $Y=0 $X2=-0.19 $Y2=-0.245
