* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__a41o_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
X0 X a_90_53# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X1 VPWR A1 a_453_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X2 a_453_367# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X3 VPWR a_90_53# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X4 a_561_49# A3 a_633_49# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X5 VGND a_90_53# X VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X6 a_633_49# A2 a_741_49# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X7 a_90_53# B1 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X8 VGND A4 a_561_49# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X9 a_741_49# A1 a_90_53# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X10 VPWR A3 a_453_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X11 a_90_53# B1 a_453_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X12 a_453_367# A4 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X13 X a_90_53# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
.ends
