* File: sky130_fd_sc_lp__mux2_2.pex.spice
* Created: Wed Sep  2 10:00:12 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__MUX2_2%A_86_21# 1 2 9 13 17 21 26 27 28 29 30 33 36
+ 37 38 40
r102 45 47 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=0.505 $Y=1.44
+ $X2=0.935 $Y2=1.44
r103 40 43 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=2.25 $Y=2.6 $X2=2.25
+ $Y2=2.68
r104 37 47 13.9889 $w=3.3e-07 $l=8e-08 $layer=POLY_cond $X=1.015 $Y=1.44
+ $X2=0.935 $Y2=1.44
r105 36 39 8.85254 $w=2.43e-07 $l=1.65e-07 $layer=LI1_cond $X=1.052 $Y=1.44
+ $X2=1.052 $Y2=1.605
r106 36 38 8.85254 $w=2.43e-07 $l=1.65e-07 $layer=LI1_cond $X=1.052 $Y=1.44
+ $X2=1.052 $Y2=1.275
r107 36 37 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.015
+ $Y=1.44 $X2=1.015 $Y2=1.44
r108 31 33 5.98384 $w=2.58e-07 $l=1.35e-07 $layer=LI1_cond $X=2.06 $Y=0.595
+ $X2=2.06 $Y2=0.46
r109 29 40 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.085 $Y=2.6
+ $X2=2.25 $Y2=2.6
r110 29 30 59.369 $w=1.68e-07 $l=9.1e-07 $layer=LI1_cond $X=2.085 $Y=2.6
+ $X2=1.175 $Y2=2.6
r111 27 31 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=1.93 $Y=0.68
+ $X2=2.06 $Y2=0.595
r112 27 28 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=1.93 $Y=0.68
+ $X2=1.175 $Y2=0.68
r113 26 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.09 $Y=2.515
+ $X2=1.175 $Y2=2.6
r114 26 39 59.369 $w=1.68e-07 $l=9.1e-07 $layer=LI1_cond $X=1.09 $Y=2.515
+ $X2=1.09 $Y2=1.605
r115 23 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.09 $Y=0.765
+ $X2=1.175 $Y2=0.68
r116 23 38 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=1.09 $Y=0.765
+ $X2=1.09 $Y2=1.275
r117 19 47 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.935 $Y=1.605
+ $X2=0.935 $Y2=1.44
r118 19 21 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=0.935 $Y=1.605
+ $X2=0.935 $Y2=2.465
r119 15 47 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.935 $Y=1.275
+ $X2=0.935 $Y2=1.44
r120 15 17 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=0.935 $Y=1.275
+ $X2=0.935 $Y2=0.655
r121 11 45 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.505 $Y=1.605
+ $X2=0.505 $Y2=1.44
r122 11 13 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=0.505 $Y=1.605
+ $X2=0.505 $Y2=2.465
r123 7 45 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.505 $Y=1.275
+ $X2=0.505 $Y2=1.44
r124 7 9 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=0.505 $Y=1.275
+ $X2=0.505 $Y2=0.655
r125 2 43 600 $w=1.7e-07 $l=5.00125e-07 $layer=licon1_PDIFF $count=1 $X=2.11
+ $Y=2.245 $X2=2.25 $Y2=2.68
r126 1 33 182 $w=1.7e-07 $l=2.85307e-07 $layer=licon1_NDIFF $count=1 $X=1.955
+ $Y=0.24 $X2=2.105 $Y2=0.46
.ends

.subckt PM_SKY130_FD_SC_LP__MUX2_2%A_284_279# 1 2 9 13 17 18 21 22 24 25 28 32
+ 34
r79 30 34 3.351 $w=2.8e-07 $l=9.44722e-08 $layer=LI1_cond $X=3.615 $Y=2.345
+ $X2=3.595 $Y2=2.26
r80 30 32 1.99461 $w=2.58e-07 $l=4.5e-08 $layer=LI1_cond $X=3.615 $Y=2.345
+ $X2=3.615 $Y2=2.39
r81 26 34 3.351 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=3.595 $Y=2.175
+ $X2=3.595 $Y2=2.26
r82 26 28 66.6496 $w=2.98e-07 $l=1.735e-06 $layer=LI1_cond $X=3.595 $Y=2.175
+ $X2=3.595 $Y2=0.44
r83 24 34 3.18746 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=3.445 $Y=2.26
+ $X2=3.595 $Y2=2.26
r84 24 25 110.583 $w=1.68e-07 $l=1.695e-06 $layer=LI1_cond $X=3.445 $Y=2.26
+ $X2=1.75 $Y2=2.26
r85 21 22 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.585
+ $Y=1.56 $X2=1.585 $Y2=1.56
r86 19 25 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.585 $Y=2.175
+ $X2=1.75 $Y2=2.26
r87 19 21 21.4773 $w=3.28e-07 $l=6.15e-07 $layer=LI1_cond $X=1.585 $Y=2.175
+ $X2=1.585 $Y2=1.56
r88 17 22 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.585 $Y=1.9
+ $X2=1.585 $Y2=1.56
r89 17 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.585 $Y=1.9
+ $X2=1.585 $Y2=2.065
r90 16 22 42.4377 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.585 $Y=1.395
+ $X2=1.585 $Y2=1.56
r91 13 18 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=1.675 $Y=2.565
+ $X2=1.675 $Y2=2.065
r92 9 16 484.564 $w=1.5e-07 $l=9.45e-07 $layer=POLY_cond $X=1.52 $Y=0.45
+ $X2=1.52 $Y2=1.395
r93 2 32 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=3.44
+ $Y=2.245 $X2=3.58 $Y2=2.39
r94 1 28 182 $w=1.7e-07 $l=2.60768e-07 $layer=licon1_NDIFF $count=1 $X=3.41
+ $Y=0.24 $X2=3.55 $Y2=0.44
.ends

.subckt PM_SKY130_FD_SC_LP__MUX2_2%A0 3 7 10 12 13 16 23 24 29
c52 23 0 1.04339e-19 $X=2.485 $Y=1.92
c53 12 0 3.86936e-20 $X=1.97 $Y=1.02
r54 27 29 0.657186 $w=4.53e-07 $l=2.5e-08 $layer=LI1_cond $X=2.135 $Y=1.777
+ $X2=2.16 $Y2=1.777
r55 23 26 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.485 $Y=1.92
+ $X2=2.485 $Y2=2.085
r56 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.485
+ $Y=1.92 $X2=2.485 $Y2=1.92
r57 16 27 2.41046 $w=4.55e-07 $l=8.5e-08 $layer=LI1_cond $X=2.05 $Y=1.777
+ $X2=2.135 $Y2=1.777
r58 16 24 7.75479 $w=4.53e-07 $l=2.95e-07 $layer=LI1_cond $X=2.19 $Y=1.777
+ $X2=2.485 $Y2=1.777
r59 16 29 0.788623 $w=4.53e-07 $l=3e-08 $layer=LI1_cond $X=2.19 $Y=1.777
+ $X2=2.16 $Y2=1.777
r60 13 20 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.97 $Y=1.02
+ $X2=1.97 $Y2=0.855
r61 12 15 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=1.97 $Y=1.02
+ $X2=1.97 $Y2=1.185
r62 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.97
+ $Y=1.02 $X2=1.97 $Y2=1.02
r63 10 16 6.43735 $w=1.7e-07 $l=2.27e-07 $layer=LI1_cond $X=2.05 $Y=1.55
+ $X2=2.05 $Y2=1.777
r64 10 15 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=2.05 $Y=1.55
+ $X2=2.05 $Y2=1.185
r65 7 26 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.465 $Y=2.565
+ $X2=2.465 $Y2=2.085
r66 3 20 207.67 $w=1.5e-07 $l=4.05e-07 $layer=POLY_cond $X=1.88 $Y=0.45 $X2=1.88
+ $Y2=0.855
.ends

.subckt PM_SKY130_FD_SC_LP__MUX2_2%A1 3 5 6 9 11 12 13 18
c56 6 0 3.86936e-20 $X=2.11 $Y=1.47
r57 13 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.525
+ $Y=1.295 $X2=2.525 $Y2=1.295
r58 12 13 11.3708 $w=3.73e-07 $l=3.7e-07 $layer=LI1_cond $X=2.547 $Y=0.925
+ $X2=2.547 $Y2=1.295
r59 11 12 11.3708 $w=3.73e-07 $l=3.7e-07 $layer=LI1_cond $X=2.547 $Y=0.555
+ $X2=2.547 $Y2=0.925
r60 7 18 38.5368 $w=3.05e-07 $l=2.07918e-07 $layer=POLY_cond $X=2.42 $Y=1.13
+ $X2=2.517 $Y2=1.295
r61 7 9 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=2.42 $Y=1.13 $X2=2.42
+ $Y2=0.45
r62 5 18 27.6557 $w=3.05e-07 $l=2.46424e-07 $layer=POLY_cond $X=2.345 $Y=1.47
+ $X2=2.517 $Y2=1.295
r63 5 6 120.5 $w=1.5e-07 $l=2.35e-07 $layer=POLY_cond $X=2.345 $Y=1.47 $X2=2.11
+ $Y2=1.47
r64 1 6 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.035 $Y=1.545
+ $X2=2.11 $Y2=1.47
r65 1 3 523.021 $w=1.5e-07 $l=1.02e-06 $layer=POLY_cond $X=2.035 $Y=1.545
+ $X2=2.035 $Y2=2.565
.ends

.subckt PM_SKY130_FD_SC_LP__MUX2_2%S 1 3 6 9 12 15 18 22 25 26 27 28 33
c55 26 0 1.04339e-19 $X=3.12 $Y=0.925
r56 27 28 13.3251 $w=3.18e-07 $l=3.7e-07 $layer=LI1_cond $X=3.115 $Y=1.295
+ $X2=3.115 $Y2=1.665
r57 27 33 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.12
+ $Y=1.345 $X2=3.12 $Y2=1.345
r58 26 27 13.3251 $w=3.18e-07 $l=3.7e-07 $layer=LI1_cond $X=3.115 $Y=0.925
+ $X2=3.115 $Y2=1.295
r59 24 25 58.3064 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=3.35 $Y=0.79
+ $X2=3.35 $Y2=0.94
r60 20 22 99.9894 $w=1.5e-07 $l=1.95e-07 $layer=POLY_cond $X=2.78 $Y=0.845
+ $X2=2.975 $Y2=0.845
r61 16 33 91.0088 $w=2.74e-07 $l=6.02993e-07 $layer=POLY_cond $X=3.365 $Y=1.85
+ $X2=3.15 $Y2=1.345
r62 16 18 366.628 $w=1.5e-07 $l=7.15e-07 $layer=POLY_cond $X=3.365 $Y=1.85
+ $X2=3.365 $Y2=2.565
r63 15 33 31.1986 $w=2.74e-07 $l=2.85832e-07 $layer=POLY_cond $X=3.365 $Y=1.18
+ $X2=3.15 $Y2=1.345
r64 15 25 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=3.365 $Y=1.18
+ $X2=3.365 $Y2=0.94
r65 12 24 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=3.335 $Y=0.45
+ $X2=3.335 $Y2=0.79
r66 9 33 31.1986 $w=2.74e-07 $l=2.43926e-07 $layer=POLY_cond $X=2.975 $Y=1.18
+ $X2=3.15 $Y2=1.345
r67 8 22 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.975 $Y=0.92
+ $X2=2.975 $Y2=0.845
r68 8 9 133.319 $w=1.5e-07 $l=2.6e-07 $layer=POLY_cond $X=2.975 $Y=0.92
+ $X2=2.975 $Y2=1.18
r69 4 33 91.0088 $w=2.74e-07 $l=6.02993e-07 $layer=POLY_cond $X=2.935 $Y=1.85
+ $X2=3.15 $Y2=1.345
r70 4 6 366.628 $w=1.5e-07 $l=7.15e-07 $layer=POLY_cond $X=2.935 $Y=1.85
+ $X2=2.935 $Y2=2.565
r71 1 20 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.78 $Y=0.77 $X2=2.78
+ $Y2=0.845
r72 1 3 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.78 $Y=0.77 $X2=2.78
+ $Y2=0.45
.ends

.subckt PM_SKY130_FD_SC_LP__MUX2_2%VPWR 1 2 3 10 12 18 22 24 26 31 41 42 48 51
r53 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r54 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r55 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r56 42 52 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=3.12 $Y2=3.33
r57 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r58 39 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.315 $Y=3.33
+ $X2=3.15 $Y2=3.33
r59 39 41 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=3.315 $Y=3.33
+ $X2=3.6 $Y2=3.33
r60 38 52 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r61 37 38 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r62 35 49 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r63 34 37 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.68 $Y=3.33 $X2=2.64
+ $Y2=3.33
r64 34 35 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r65 32 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.315 $Y=3.33
+ $X2=1.15 $Y2=3.33
r66 32 34 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=1.315 $Y=3.33
+ $X2=1.68 $Y2=3.33
r67 31 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.985 $Y=3.33
+ $X2=3.15 $Y2=3.33
r68 31 37 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=2.985 $Y=3.33
+ $X2=2.64 $Y2=3.33
r69 30 49 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r70 30 46 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r71 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r72 27 45 4.30888 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=0.41 $Y=3.33
+ $X2=0.205 $Y2=3.33
r73 27 29 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=0.41 $Y=3.33
+ $X2=0.72 $Y2=3.33
r74 26 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.985 $Y=3.33
+ $X2=1.15 $Y2=3.33
r75 26 29 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.985 $Y=3.33
+ $X2=0.72 $Y2=3.33
r76 24 38 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=2.64 $Y2=3.33
r77 24 35 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=1.68 $Y2=3.33
r78 20 51 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.15 $Y=3.245
+ $X2=3.15 $Y2=3.33
r79 20 22 20.7789 $w=3.28e-07 $l=5.95e-07 $layer=LI1_cond $X=3.15 $Y=3.245
+ $X2=3.15 $Y2=2.65
r80 16 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.15 $Y=3.245
+ $X2=1.15 $Y2=3.33
r81 16 18 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=1.15 $Y=3.245
+ $X2=1.15 $Y2=2.97
r82 12 15 39.2235 $w=2.83e-07 $l=9.7e-07 $layer=LI1_cond $X=0.267 $Y=1.98
+ $X2=0.267 $Y2=2.95
r83 10 45 3.08979 $w=2.85e-07 $l=1.11781e-07 $layer=LI1_cond $X=0.267 $Y=3.245
+ $X2=0.205 $Y2=3.33
r84 10 15 11.9288 $w=2.83e-07 $l=2.95e-07 $layer=LI1_cond $X=0.267 $Y=3.245
+ $X2=0.267 $Y2=2.95
r85 3 22 600 $w=1.7e-07 $l=4.69814e-07 $layer=licon1_PDIFF $count=1 $X=3.01
+ $Y=2.245 $X2=3.15 $Y2=2.65
r86 2 18 600 $w=1.7e-07 $l=1.20297e-06 $layer=licon1_PDIFF $count=1 $X=1.01
+ $Y=1.835 $X2=1.15 $Y2=2.97
r87 1 15 400 $w=1.7e-07 $l=1.17584e-06 $layer=licon1_PDIFF $count=1 $X=0.165
+ $Y=1.835 $X2=0.29 $Y2=2.95
r88 1 12 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.165
+ $Y=1.835 $X2=0.29 $Y2=1.98
.ends

.subckt PM_SKY130_FD_SC_LP__MUX2_2%X 1 2 9 13 14 15 16 24 34
r23 21 24 2.71464 $w=2.23e-07 $l=5.3e-08 $layer=LI1_cond $X=0.692 $Y=1.962
+ $X2=0.692 $Y2=2.015
r24 16 31 6.91466 $w=2.23e-07 $l=1.35e-07 $layer=LI1_cond $X=0.692 $Y=2.775
+ $X2=0.692 $Y2=2.91
r25 15 16 18.9513 $w=2.23e-07 $l=3.7e-07 $layer=LI1_cond $X=0.692 $Y=2.405
+ $X2=0.692 $Y2=2.775
r26 14 21 0.307318 $w=2.23e-07 $l=6e-09 $layer=LI1_cond $X=0.692 $Y=1.956
+ $X2=0.692 $Y2=1.962
r27 14 34 6.1449 $w=2.23e-07 $l=1.06e-07 $layer=LI1_cond $X=0.692 $Y=1.956
+ $X2=0.692 $Y2=1.85
r28 14 15 18.644 $w=2.23e-07 $l=3.64e-07 $layer=LI1_cond $X=0.692 $Y=2.041
+ $X2=0.692 $Y2=2.405
r29 14 24 1.33171 $w=2.23e-07 $l=2.6e-08 $layer=LI1_cond $X=0.692 $Y=2.041
+ $X2=0.692 $Y2=2.015
r30 13 34 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=0.665 $Y=1.095
+ $X2=0.665 $Y2=1.85
r31 7 13 7.02311 $w=2.53e-07 $l=1.27e-07 $layer=LI1_cond $X=0.707 $Y=0.968
+ $X2=0.707 $Y2=1.095
r32 7 9 24.7662 $w=2.53e-07 $l=5.48e-07 $layer=LI1_cond $X=0.707 $Y=0.968
+ $X2=0.707 $Y2=0.42
r33 2 31 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=0.58
+ $Y=1.835 $X2=0.72 $Y2=2.91
r34 2 24 400 $w=1.7e-07 $l=2.4e-07 $layer=licon1_PDIFF $count=1 $X=0.58 $Y=1.835
+ $X2=0.72 $Y2=2.015
r35 1 9 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=0.58
+ $Y=0.235 $X2=0.72 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__MUX2_2%VGND 1 2 3 10 12 16 20 22 24 29 39 40 46 49
r60 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r61 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r62 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r63 40 50 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=3.12
+ $Y2=0
r64 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r65 37 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.235 $Y=0 $X2=3.07
+ $Y2=0
r66 37 39 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=3.235 $Y=0 $X2=3.6
+ $Y2=0
r67 36 50 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r68 35 36 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r69 33 47 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r70 32 35 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r71 32 33 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r72 30 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.375 $Y=0 $X2=1.21
+ $Y2=0
r73 30 32 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.375 $Y=0 $X2=1.68
+ $Y2=0
r74 29 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.905 $Y=0 $X2=3.07
+ $Y2=0
r75 29 35 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=2.905 $Y=0 $X2=2.64
+ $Y2=0
r76 28 47 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r77 28 44 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r78 27 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r79 25 43 4.30888 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=0.41 $Y=0 $X2=0.205
+ $Y2=0
r80 25 27 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=0.41 $Y=0 $X2=0.72
+ $Y2=0
r81 24 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.045 $Y=0 $X2=1.21
+ $Y2=0
r82 24 27 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=1.045 $Y=0 $X2=0.72
+ $Y2=0
r83 22 36 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=2.64
+ $Y2=0
r84 22 33 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=1.68
+ $Y2=0
r85 18 49 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.07 $Y=0.085
+ $X2=3.07 $Y2=0
r86 18 20 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=3.07 $Y=0.085
+ $X2=3.07 $Y2=0.45
r87 14 46 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.21 $Y=0.085
+ $X2=1.21 $Y2=0
r88 14 16 8.20679 $w=3.28e-07 $l=2.35e-07 $layer=LI1_cond $X=1.21 $Y=0.085
+ $X2=1.21 $Y2=0.32
r89 10 43 3.08979 $w=2.85e-07 $l=1.11781e-07 $layer=LI1_cond $X=0.267 $Y=0.085
+ $X2=0.205 $Y2=0
r90 10 12 11.9288 $w=2.83e-07 $l=2.95e-07 $layer=LI1_cond $X=0.267 $Y=0.085
+ $X2=0.267 $Y2=0.38
r91 3 20 182 $w=1.7e-07 $l=3.02283e-07 $layer=licon1_NDIFF $count=1 $X=2.855
+ $Y=0.24 $X2=3.07 $Y2=0.45
r92 2 16 182 $w=1.7e-07 $l=2.38747e-07 $layer=licon1_NDIFF $count=1 $X=1.01
+ $Y=0.235 $X2=1.21 $Y2=0.32
r93 1 12 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.165
+ $Y=0.235 $X2=0.29 $Y2=0.38
.ends

