* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__a21bo_4 A1 A2 B1_N VGND VNB VPB VPWR X
X0 a_188_315# a_42_47# a_645_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X1 X a_188_315# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X2 VGND a_188_315# X VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X3 X a_188_315# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X4 a_645_367# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X5 X a_188_315# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X6 VPWR a_188_315# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X7 a_42_47# B1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X8 VGND a_42_47# a_188_315# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X9 a_188_315# A1 a_908_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X10 a_42_47# B1_N VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X11 a_188_315# a_42_47# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X12 a_908_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X13 X a_188_315# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X14 VGND A2 a_908_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X15 a_645_367# a_42_47# a_188_315# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X16 a_908_47# A1 a_188_315# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X17 VPWR a_188_315# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X18 VPWR A2 a_645_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X19 a_645_367# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X20 VPWR A1 a_645_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X21 VGND a_188_315# X VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
.ends
