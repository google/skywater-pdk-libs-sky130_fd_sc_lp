* File: sky130_fd_sc_lp__nor4bb_4.pex.spice
* Created: Wed Sep  2 10:11:46 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__NOR4BB_4%D_N 3 7 9 13 15
c25 7 0 1.55299e-19 $X=0.525 $Y=2.465
r26 12 15 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=0.31 $Y=1.46
+ $X2=0.525 $Y2=1.46
r27 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.31
+ $Y=1.46 $X2=0.31 $Y2=1.46
r28 9 13 6.05771 $w=3.88e-07 $l=2.05e-07 $layer=LI1_cond $X=0.28 $Y=1.665
+ $X2=0.28 $Y2=1.46
r29 5 15 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.525 $Y=1.625
+ $X2=0.525 $Y2=1.46
r30 5 7 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=0.525 $Y=1.625
+ $X2=0.525 $Y2=2.465
r31 1 15 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.525 $Y=1.295
+ $X2=0.525 $Y2=1.46
r32 1 3 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=0.525 $Y=1.295
+ $X2=0.525 $Y2=0.675
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4BB_4%C_N 3 7 9 12 13
r33 12 15 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=1.067 $Y=1.51
+ $X2=1.067 $Y2=1.675
r34 12 14 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=1.067 $Y=1.51
+ $X2=1.067 $Y2=1.345
r35 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.09
+ $Y=1.51 $X2=1.09 $Y2=1.51
r36 9 13 6.15961 $w=2.88e-07 $l=1.55e-07 $layer=LI1_cond $X=1.14 $Y=1.665
+ $X2=1.14 $Y2=1.51
r37 7 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=0.955 $Y=2.465
+ $X2=0.955 $Y2=1.675
r38 3 14 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=0.955 $Y=0.675
+ $X2=0.955 $Y2=1.345
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4BB_4%A_37_51# 1 2 9 13 17 21 25 29 33 37 41 45
+ 47 48 50 51 53 54 57 65 79
c138 33 0 7.76303e-20 $X=3.365 $Y=2.375
r139 78 79 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=3.365 $Y=1.42
+ $X2=3.435 $Y2=1.42
r140 75 76 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=2.935 $Y=1.42
+ $X2=3.005 $Y2=1.42
r141 74 75 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=2.505 $Y=1.42
+ $X2=2.935 $Y2=1.42
r142 73 74 17.4861 $w=3.3e-07 $l=1e-07 $layer=POLY_cond $X=2.405 $Y=1.42
+ $X2=2.505 $Y2=1.42
r143 72 73 57.7042 $w=3.3e-07 $l=3.3e-07 $layer=POLY_cond $X=2.075 $Y=1.42
+ $X2=2.405 $Y2=1.42
r144 68 72 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=1.985 $Y=1.42
+ $X2=2.075 $Y2=1.42
r145 68 69 1.74861 $w=3.3e-07 $l=1e-08 $layer=POLY_cond $X=1.985 $Y=1.42
+ $X2=1.975 $Y2=1.42
r146 67 68 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=1.985
+ $Y=1.42 $X2=1.985 $Y2=1.42
r147 64 65 8.20096 $w=5.48e-07 $l=9e-08 $layer=LI1_cond $X=0.735 $Y=2.205
+ $X2=0.825 $Y2=2.205
r148 63 64 9.24242 $w=5.48e-07 $l=4.25e-07 $layer=LI1_cond $X=0.31 $Y=2.205
+ $X2=0.735 $Y2=2.205
r149 60 63 0.761141 $w=5.48e-07 $l=3.5e-08 $layer=LI1_cond $X=0.275 $Y=2.205
+ $X2=0.31 $Y2=2.205
r150 58 78 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=3.345 $Y=1.42
+ $X2=3.365 $Y2=1.42
r151 58 76 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=3.345 $Y=1.42
+ $X2=3.005 $Y2=1.42
r152 57 58 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=3.345
+ $Y=1.42 $X2=3.345 $Y2=1.42
r153 55 67 3.6578 $w=1.8e-07 $l=1.03e-07 $layer=LI1_cond $X=2.025 $Y=1.425
+ $X2=1.922 $Y2=1.425
r154 55 57 81.3333 $w=1.78e-07 $l=1.32e-06 $layer=LI1_cond $X=2.025 $Y=1.425
+ $X2=3.345 $Y2=1.425
r155 53 67 3.19614 $w=2.05e-07 $l=9e-08 $layer=LI1_cond $X=1.922 $Y=1.515
+ $X2=1.922 $Y2=1.425
r156 53 54 43.0111 $w=2.03e-07 $l=7.95e-07 $layer=LI1_cond $X=1.922 $Y=1.515
+ $X2=1.922 $Y2=2.31
r157 51 54 6.89401 $w=1.7e-07 $l=1.38109e-07 $layer=LI1_cond $X=1.82 $Y=2.395
+ $X2=1.922 $Y2=2.31
r158 51 65 64.9144 $w=1.68e-07 $l=9.95e-07 $layer=LI1_cond $X=1.82 $Y=2.395
+ $X2=0.825 $Y2=2.395
r159 50 64 7.39687 $w=1.8e-07 $l=2.75e-07 $layer=LI1_cond $X=0.735 $Y=1.93
+ $X2=0.735 $Y2=2.205
r160 49 50 45.2879 $w=1.78e-07 $l=7.35e-07 $layer=LI1_cond $X=0.735 $Y=1.195
+ $X2=0.735 $Y2=1.93
r161 47 49 6.82373 $w=1.7e-07 $l=1.25499e-07 $layer=LI1_cond $X=0.645 $Y=1.11
+ $X2=0.735 $Y2=1.195
r162 47 48 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=0.645 $Y=1.11
+ $X2=0.395 $Y2=1.11
r163 43 60 5.13615 $w=2.6e-07 $l=2.75e-07 $layer=LI1_cond $X=0.275 $Y=2.48
+ $X2=0.275 $Y2=2.205
r164 43 45 0.443247 $w=2.58e-07 $l=1e-08 $layer=LI1_cond $X=0.275 $Y=2.48
+ $X2=0.275 $Y2=2.49
r165 39 48 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.27 $Y=1.025
+ $X2=0.395 $Y2=1.11
r166 39 41 27.8891 $w=2.48e-07 $l=6.05e-07 $layer=LI1_cond $X=0.27 $Y=1.025
+ $X2=0.27 $Y2=0.42
r167 35 79 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.435 $Y=1.255
+ $X2=3.435 $Y2=1.42
r168 35 37 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=3.435 $Y=1.255
+ $X2=3.435 $Y2=0.655
r169 31 78 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.365 $Y=1.585
+ $X2=3.365 $Y2=1.42
r170 31 33 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.365 $Y=1.585
+ $X2=3.365 $Y2=2.375
r171 27 76 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.005 $Y=1.255
+ $X2=3.005 $Y2=1.42
r172 27 29 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=3.005 $Y=1.255
+ $X2=3.005 $Y2=0.655
r173 23 75 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.935 $Y=1.585
+ $X2=2.935 $Y2=1.42
r174 23 25 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.935 $Y=1.585
+ $X2=2.935 $Y2=2.375
r175 19 74 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.505 $Y=1.585
+ $X2=2.505 $Y2=1.42
r176 19 21 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.505 $Y=1.585
+ $X2=2.505 $Y2=2.375
r177 15 73 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.405 $Y=1.255
+ $X2=2.405 $Y2=1.42
r178 15 17 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=2.405 $Y=1.255
+ $X2=2.405 $Y2=0.655
r179 11 72 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.075 $Y=1.585
+ $X2=2.075 $Y2=1.42
r180 11 13 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.075 $Y=1.585
+ $X2=2.075 $Y2=2.375
r181 7 69 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.975 $Y=1.255
+ $X2=1.975 $Y2=1.42
r182 7 9 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=1.975 $Y=1.255 $X2=1.975
+ $Y2=0.655
r183 2 63 600 $w=1.7e-07 $l=3.16386e-07 $layer=licon1_PDIFF $count=1 $X=0.185
+ $Y=1.835 $X2=0.31 $Y2=2.095
r184 2 45 300 $w=1.7e-07 $l=7.14773e-07 $layer=licon1_PDIFF $count=2 $X=0.185
+ $Y=1.835 $X2=0.31 $Y2=2.49
r185 1 41 91 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=2 $X=0.185
+ $Y=0.255 $X2=0.31 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4BB_4%A_206_51# 1 2 9 13 17 21 25 29 33 37 39 45
+ 48 49 52 55 61 75
c145 75 0 1.8609e-19 $X=5.225 $Y=1.42
c146 39 0 1.55299e-19 $X=1.455 $Y=2.035
c147 29 0 5.06642e-20 $X=4.795 $Y=0.655
c148 17 0 5.86634e-20 $X=4.225 $Y=2.375
r149 74 75 24.4806 $w=3.3e-07 $l=1.4e-07 $layer=POLY_cond $X=5.085 $Y=1.42
+ $X2=5.225 $Y2=1.42
r150 71 72 24.4806 $w=3.3e-07 $l=1.4e-07 $layer=POLY_cond $X=4.655 $Y=1.42
+ $X2=4.795 $Y2=1.42
r151 70 71 50.7098 $w=3.3e-07 $l=2.9e-07 $layer=POLY_cond $X=4.365 $Y=1.42
+ $X2=4.655 $Y2=1.42
r152 69 70 24.4806 $w=3.3e-07 $l=1.4e-07 $layer=POLY_cond $X=4.225 $Y=1.42
+ $X2=4.365 $Y2=1.42
r153 68 69 50.7098 $w=3.3e-07 $l=2.9e-07 $layer=POLY_cond $X=3.935 $Y=1.42
+ $X2=4.225 $Y2=1.42
r154 64 68 8.74306 $w=3.3e-07 $l=5e-08 $layer=POLY_cond $X=3.885 $Y=1.42
+ $X2=3.935 $Y2=1.42
r155 64 65 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=3.885 $Y=1.42
+ $X2=3.795 $Y2=1.42
r156 63 64 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.885
+ $Y=1.42 $X2=3.885 $Y2=1.42
r157 60 61 5.59224 $w=1.78e-07 $l=9e-08 $layer=LI1_cond $X=1.545 $Y=1.085
+ $X2=1.635 $Y2=1.085
r158 56 74 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=4.905 $Y=1.42
+ $X2=5.085 $Y2=1.42
r159 56 72 19.2347 $w=3.3e-07 $l=1.1e-07 $layer=POLY_cond $X=4.905 $Y=1.42
+ $X2=4.795 $Y2=1.42
r160 55 56 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.905
+ $Y=1.42 $X2=4.905 $Y2=1.42
r161 53 63 3.31438 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=3.89 $Y=1.425
+ $X2=3.805 $Y2=1.425
r162 53 55 62.5404 $w=1.78e-07 $l=1.015e-06 $layer=LI1_cond $X=3.89 $Y=1.425
+ $X2=4.905 $Y2=1.425
r163 52 63 3.50935 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=3.805 $Y=1.335
+ $X2=3.805 $Y2=1.425
r164 51 52 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=3.805 $Y=1.165
+ $X2=3.805 $Y2=1.335
r165 49 51 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.72 $Y=1.08
+ $X2=3.805 $Y2=1.165
r166 49 61 136.027 $w=1.68e-07 $l=2.085e-06 $layer=LI1_cond $X=3.72 $Y=1.08
+ $X2=1.635 $Y2=1.08
r167 47 60 0.716491 $w=1.8e-07 $l=9e-08 $layer=LI1_cond $X=1.545 $Y=1.175
+ $X2=1.545 $Y2=1.085
r168 47 48 46.5202 $w=1.78e-07 $l=7.55e-07 $layer=LI1_cond $X=1.545 $Y=1.175
+ $X2=1.545 $Y2=1.93
r169 43 60 20.9495 $w=1.78e-07 $l=3.4e-07 $layer=LI1_cond $X=1.205 $Y=1.085
+ $X2=1.545 $Y2=1.085
r170 43 45 25.4867 $w=2.58e-07 $l=5.75e-07 $layer=LI1_cond $X=1.205 $Y=0.995
+ $X2=1.205 $Y2=0.42
r171 39 48 6.86909 $w=2.1e-07 $l=1.43091e-07 $layer=LI1_cond $X=1.455 $Y=2.035
+ $X2=1.545 $Y2=1.93
r172 39 41 15.0519 $w=2.08e-07 $l=2.85e-07 $layer=LI1_cond $X=1.455 $Y=2.035
+ $X2=1.17 $Y2=2.035
r173 35 75 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.225 $Y=1.255
+ $X2=5.225 $Y2=1.42
r174 35 37 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=5.225 $Y=1.255
+ $X2=5.225 $Y2=0.655
r175 31 74 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.085 $Y=1.585
+ $X2=5.085 $Y2=1.42
r176 31 33 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=5.085 $Y=1.585
+ $X2=5.085 $Y2=2.375
r177 27 72 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.795 $Y=1.255
+ $X2=4.795 $Y2=1.42
r178 27 29 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=4.795 $Y=1.255
+ $X2=4.795 $Y2=0.655
r179 23 71 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.655 $Y=1.585
+ $X2=4.655 $Y2=1.42
r180 23 25 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=4.655 $Y=1.585
+ $X2=4.655 $Y2=2.375
r181 19 70 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.365 $Y=1.255
+ $X2=4.365 $Y2=1.42
r182 19 21 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=4.365 $Y=1.255
+ $X2=4.365 $Y2=0.655
r183 15 69 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.225 $Y=1.585
+ $X2=4.225 $Y2=1.42
r184 15 17 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=4.225 $Y=1.585
+ $X2=4.225 $Y2=2.375
r185 11 68 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.935 $Y=1.255
+ $X2=3.935 $Y2=1.42
r186 11 13 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=3.935 $Y=1.255
+ $X2=3.935 $Y2=0.655
r187 7 65 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.795 $Y=1.585
+ $X2=3.795 $Y2=1.42
r188 7 9 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.795 $Y=1.585
+ $X2=3.795 $Y2=2.375
r189 2 41 600 $w=1.7e-07 $l=2.60768e-07 $layer=licon1_PDIFF $count=1 $X=1.03
+ $Y=1.835 $X2=1.17 $Y2=2.035
r190 1 45 91 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=2 $X=1.03
+ $Y=0.255 $X2=1.17 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4BB_4%B 3 7 11 15 19 23 27 31 38 41 45 56
c107 45 0 1.8609e-19 $X=5.95 $Y=1.44
r108 55 56 0.874306 $w=3.3e-07 $l=5e-09 $layer=POLY_cond $X=7.325 $Y=1.44
+ $X2=7.33 $Y2=1.44
r109 52 53 0.874306 $w=3.3e-07 $l=5e-09 $layer=POLY_cond $X=6.895 $Y=1.44
+ $X2=6.9 $Y2=1.44
r110 51 52 74.316 $w=3.3e-07 $l=4.25e-07 $layer=POLY_cond $X=6.47 $Y=1.44
+ $X2=6.895 $Y2=1.44
r111 50 51 0.874306 $w=3.3e-07 $l=5e-09 $layer=POLY_cond $X=6.465 $Y=1.44
+ $X2=6.47 $Y2=1.44
r112 47 48 0.874306 $w=3.3e-07 $l=5e-09 $layer=POLY_cond $X=6.035 $Y=1.44
+ $X2=6.04 $Y2=1.44
r113 44 47 14.8632 $w=3.3e-07 $l=8.5e-08 $layer=POLY_cond $X=5.95 $Y=1.44
+ $X2=6.035 $Y2=1.44
r114 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.95
+ $Y=1.44 $X2=5.95 $Y2=1.44
r115 41 45 6.1738 $w=4.18e-07 $l=2.25e-07 $layer=LI1_cond $X=5.995 $Y=1.665
+ $X2=5.995 $Y2=1.44
r116 39 55 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=7.31 $Y=1.44
+ $X2=7.325 $Y2=1.44
r117 39 53 71.6931 $w=3.3e-07 $l=4.1e-07 $layer=POLY_cond $X=7.31 $Y=1.44
+ $X2=6.9 $Y2=1.44
r118 38 39 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.31
+ $Y=1.44 $X2=7.31 $Y2=1.44
r119 36 50 30.6007 $w=3.3e-07 $l=1.75e-07 $layer=POLY_cond $X=6.29 $Y=1.44
+ $X2=6.465 $Y2=1.44
r120 36 48 43.7153 $w=3.3e-07 $l=2.5e-07 $layer=POLY_cond $X=6.29 $Y=1.44
+ $X2=6.04 $Y2=1.44
r121 35 38 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=6.29 $Y=1.44
+ $X2=7.31 $Y2=1.44
r122 35 36 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.29
+ $Y=1.44 $X2=6.29 $Y2=1.44
r123 33 45 6.07598 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=6.205 $Y=1.44
+ $X2=5.995 $Y2=1.44
r124 33 35 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=6.205 $Y=1.44
+ $X2=6.29 $Y2=1.44
r125 29 56 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.33 $Y=1.275
+ $X2=7.33 $Y2=1.44
r126 29 31 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=7.33 $Y=1.275
+ $X2=7.33 $Y2=0.655
r127 25 55 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.325 $Y=1.605
+ $X2=7.325 $Y2=1.44
r128 25 27 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=7.325 $Y=1.605
+ $X2=7.325 $Y2=2.465
r129 21 53 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.9 $Y=1.275
+ $X2=6.9 $Y2=1.44
r130 21 23 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=6.9 $Y=1.275
+ $X2=6.9 $Y2=0.655
r131 17 52 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.895 $Y=1.605
+ $X2=6.895 $Y2=1.44
r132 17 19 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=6.895 $Y=1.605
+ $X2=6.895 $Y2=2.465
r133 13 51 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.47 $Y=1.275
+ $X2=6.47 $Y2=1.44
r134 13 15 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=6.47 $Y=1.275
+ $X2=6.47 $Y2=0.655
r135 9 50 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.465 $Y=1.605
+ $X2=6.465 $Y2=1.44
r136 9 11 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=6.465 $Y=1.605
+ $X2=6.465 $Y2=2.465
r137 5 48 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.04 $Y=1.275
+ $X2=6.04 $Y2=1.44
r138 5 7 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=6.04 $Y=1.275
+ $X2=6.04 $Y2=0.655
r139 1 47 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.035 $Y=1.605
+ $X2=6.035 $Y2=1.44
r140 1 3 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=6.035 $Y=1.605
+ $X2=6.035 $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4BB_4%A 3 7 11 15 19 23 27 31 33 34 35 36 41 43
r77 57 59 10.4917 $w=3.3e-07 $l=6e-08 $layer=POLY_cond $X=8.99 $Y=1.46 $X2=9.05
+ $Y2=1.46
r78 57 58 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=8.99
+ $Y=1.46 $X2=8.99 $Y2=1.46
r79 55 57 64.6987 $w=3.3e-07 $l=3.7e-07 $layer=POLY_cond $X=8.62 $Y=1.46
+ $X2=8.99 $Y2=1.46
r80 53 55 54.207 $w=3.3e-07 $l=3.1e-07 $layer=POLY_cond $X=8.31 $Y=1.46 $X2=8.62
+ $Y2=1.46
r81 53 54 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.31
+ $Y=1.46 $X2=8.31 $Y2=1.46
r82 51 53 20.9834 $w=3.3e-07 $l=1.2e-07 $layer=POLY_cond $X=8.19 $Y=1.46
+ $X2=8.31 $Y2=1.46
r83 50 54 10.1774 $w=3.83e-07 $l=3.4e-07 $layer=LI1_cond $X=7.97 $Y=1.567
+ $X2=8.31 $Y2=1.567
r84 49 51 38.4695 $w=3.3e-07 $l=2.2e-07 $layer=POLY_cond $X=7.97 $Y=1.46
+ $X2=8.19 $Y2=1.46
r85 49 50 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.97
+ $Y=1.46 $X2=7.97 $Y2=1.46
r86 46 49 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=7.76 $Y=1.46
+ $X2=7.97 $Y2=1.46
r87 44 58 10.1774 $w=3.83e-07 $l=3.4e-07 $layer=LI1_cond $X=9.33 $Y=1.567
+ $X2=8.99 $Y2=1.567
r88 43 44 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.33
+ $Y=1.46 $X2=9.33 $Y2=1.46
r89 41 59 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=9.125 $Y=1.46
+ $X2=9.05 $Y2=1.46
r90 41 43 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=9.125 $Y=1.46
+ $X2=9.33 $Y2=1.46
r91 36 44 0.898008 $w=3.83e-07 $l=3e-08 $layer=LI1_cond $X=9.36 $Y=1.567
+ $X2=9.33 $Y2=1.567
r92 35 58 3.29269 $w=3.83e-07 $l=1.1e-07 $layer=LI1_cond $X=8.88 $Y=1.567
+ $X2=8.99 $Y2=1.567
r93 34 35 14.3681 $w=3.83e-07 $l=4.8e-07 $layer=LI1_cond $X=8.4 $Y=1.567
+ $X2=8.88 $Y2=1.567
r94 34 54 2.69402 $w=3.83e-07 $l=9e-08 $layer=LI1_cond $X=8.4 $Y=1.567 $X2=8.31
+ $Y2=1.567
r95 33 50 1.49668 $w=3.83e-07 $l=5e-08 $layer=LI1_cond $X=7.92 $Y=1.567 $X2=7.97
+ $Y2=1.567
r96 29 59 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.05 $Y=1.625
+ $X2=9.05 $Y2=1.46
r97 29 31 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=9.05 $Y=1.625
+ $X2=9.05 $Y2=2.465
r98 25 59 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.05 $Y=1.295
+ $X2=9.05 $Y2=1.46
r99 25 27 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=9.05 $Y=1.295
+ $X2=9.05 $Y2=0.655
r100 21 55 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.62 $Y=1.625
+ $X2=8.62 $Y2=1.46
r101 21 23 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=8.62 $Y=1.625
+ $X2=8.62 $Y2=2.465
r102 17 55 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.62 $Y=1.295
+ $X2=8.62 $Y2=1.46
r103 17 19 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=8.62 $Y=1.295
+ $X2=8.62 $Y2=0.655
r104 13 51 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.19 $Y=1.625
+ $X2=8.19 $Y2=1.46
r105 13 15 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=8.19 $Y=1.625
+ $X2=8.19 $Y2=2.465
r106 9 51 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.19 $Y=1.295
+ $X2=8.19 $Y2=1.46
r107 9 11 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=8.19 $Y=1.295
+ $X2=8.19 $Y2=0.655
r108 5 46 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.76 $Y=1.625
+ $X2=7.76 $Y2=1.46
r109 5 7 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=7.76 $Y=1.625
+ $X2=7.76 $Y2=2.465
r110 1 46 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.76 $Y=1.295
+ $X2=7.76 $Y2=1.46
r111 1 3 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=7.76 $Y=1.295 $X2=7.76
+ $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4BB_4%VPWR 1 2 3 12 16 20 22 24 29 37 44 45 48 51
+ 54
r105 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r106 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r107 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r108 45 55 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=8.88 $Y2=3.33
r109 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r110 42 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9 $Y=3.33 $X2=8.835
+ $Y2=3.33
r111 42 44 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=9 $Y=3.33 $X2=9.36
+ $Y2=3.33
r112 41 55 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=8.88 $Y2=3.33
r113 41 52 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=7.92 $Y2=3.33
r114 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=3.33 $X2=8.4
+ $Y2=3.33
r115 38 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.14 $Y=3.33
+ $X2=7.975 $Y2=3.33
r116 38 40 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=8.14 $Y=3.33
+ $X2=8.4 $Y2=3.33
r117 37 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.67 $Y=3.33
+ $X2=8.835 $Y2=3.33
r118 37 40 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=8.67 $Y=3.33 $X2=8.4
+ $Y2=3.33
r119 36 52 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=7.92 $Y2=3.33
r120 35 36 1.32857 $w=1.7e-07 $l=1.19e-06 $layer=mcon $count=7 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r121 33 49 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r122 32 35 407.102 $w=1.68e-07 $l=6.24e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=7.44 $Y2=3.33
r123 32 33 1.32857 $w=1.7e-07 $l=1.19e-06 $layer=mcon $count=7 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r124 30 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.905 $Y=3.33
+ $X2=0.74 $Y2=3.33
r125 30 32 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.905 $Y=3.33
+ $X2=1.2 $Y2=3.33
r126 29 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.81 $Y=3.33
+ $X2=7.975 $Y2=3.33
r127 29 35 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=7.81 $Y=3.33
+ $X2=7.44 $Y2=3.33
r128 27 49 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r129 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r130 24 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.575 $Y=3.33
+ $X2=0.74 $Y2=3.33
r131 24 26 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=0.575 $Y=3.33
+ $X2=0.24 $Y2=3.33
r132 22 36 0.73586 $w=4.9e-07 $l=2.64e-06 $layer=MET1_cond $X=4.8 $Y=3.33
+ $X2=7.44 $Y2=3.33
r133 22 33 1.00344 $w=4.9e-07 $l=3.6e-06 $layer=MET1_cond $X=4.8 $Y=3.33 $X2=1.2
+ $Y2=3.33
r134 18 54 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.835 $Y=3.245
+ $X2=8.835 $Y2=3.33
r135 18 20 30.208 $w=3.28e-07 $l=8.65e-07 $layer=LI1_cond $X=8.835 $Y=3.245
+ $X2=8.835 $Y2=2.38
r136 14 51 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.975 $Y=3.245
+ $X2=7.975 $Y2=3.33
r137 14 16 30.208 $w=3.28e-07 $l=8.65e-07 $layer=LI1_cond $X=7.975 $Y=3.245
+ $X2=7.975 $Y2=2.38
r138 10 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.74 $Y=3.245
+ $X2=0.74 $Y2=3.33
r139 10 12 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=0.74 $Y=3.245
+ $X2=0.74 $Y2=2.8
r140 3 20 300 $w=1.7e-07 $l=6.11003e-07 $layer=licon1_PDIFF $count=2 $X=8.695
+ $Y=1.835 $X2=8.835 $Y2=2.38
r141 2 16 300 $w=1.7e-07 $l=6.11003e-07 $layer=licon1_PDIFF $count=2 $X=7.835
+ $Y=1.835 $X2=7.975 $Y2=2.38
r142 1 12 600 $w=1.7e-07 $l=1.03263e-06 $layer=licon1_PDIFF $count=1 $X=0.6
+ $Y=1.835 $X2=0.74 $Y2=2.8
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4BB_4%A_347_349# 1 2 3 4 5 16 20 24 26 30 34 36
+ 41 45 49 51
r62 41 43 6.80989 $w=3.28e-07 $l=1.95e-07 $layer=LI1_cond $X=1.86 $Y=2.795
+ $X2=1.86 $Y2=2.99
r63 37 49 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=4.535 $Y=2.12
+ $X2=4.44 $Y2=2.12
r64 36 51 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=5.205 $Y=2.12
+ $X2=5.335 $Y2=2.12
r65 36 37 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.205 $Y=2.12
+ $X2=4.535 $Y2=2.12
r66 32 49 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=4.44 $Y=2.205
+ $X2=4.44 $Y2=2.12
r67 32 34 21.3062 $w=1.88e-07 $l=3.65e-07 $layer=LI1_cond $X=4.44 $Y=2.205
+ $X2=4.44 $Y2=2.57
r68 31 47 3.92798 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=3.675 $Y=2.12
+ $X2=3.565 $Y2=2.12
r69 30 49 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=4.345 $Y=2.12
+ $X2=4.44 $Y2=2.12
r70 30 31 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.345 $Y=2.12
+ $X2=3.675 $Y2=2.12
r71 27 29 1.30959 $w=2.18e-07 $l=2.5e-08 $layer=LI1_cond $X=3.565 $Y=2.905
+ $X2=3.565 $Y2=2.88
r72 26 47 3.03526 $w=2.2e-07 $l=8.5e-08 $layer=LI1_cond $X=3.565 $Y=2.205
+ $X2=3.565 $Y2=2.12
r73 26 29 35.359 $w=2.18e-07 $l=6.75e-07 $layer=LI1_cond $X=3.565 $Y=2.205
+ $X2=3.565 $Y2=2.88
r74 25 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.885 $Y=2.99
+ $X2=2.72 $Y2=2.99
r75 24 27 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=3.455 $Y=2.99
+ $X2=3.565 $Y2=2.905
r76 24 25 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=3.455 $Y=2.99
+ $X2=2.885 $Y2=2.99
r77 20 23 26.8903 $w=3.28e-07 $l=7.7e-07 $layer=LI1_cond $X=2.72 $Y=2.11
+ $X2=2.72 $Y2=2.88
r78 18 45 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.72 $Y=2.905
+ $X2=2.72 $Y2=2.99
r79 18 23 0.873063 $w=3.28e-07 $l=2.5e-08 $layer=LI1_cond $X=2.72 $Y=2.905
+ $X2=2.72 $Y2=2.88
r80 17 43 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.025 $Y=2.99
+ $X2=1.86 $Y2=2.99
r81 16 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.555 $Y=2.99
+ $X2=2.72 $Y2=2.99
r82 16 17 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=2.555 $Y=2.99
+ $X2=2.025 $Y2=2.99
r83 5 51 300 $w=1.7e-07 $l=5.20312e-07 $layer=licon1_PDIFF $count=2 $X=5.16
+ $Y=1.745 $X2=5.3 $Y2=2.2
r84 4 49 600 $w=1.7e-07 $l=4.3946e-07 $layer=licon1_PDIFF $count=1 $X=4.3
+ $Y=1.745 $X2=4.44 $Y2=2.12
r85 4 34 600 $w=1.7e-07 $l=8.92258e-07 $layer=licon1_PDIFF $count=1 $X=4.3
+ $Y=1.745 $X2=4.44 $Y2=2.57
r86 3 47 400 $w=1.7e-07 $l=5.20312e-07 $layer=licon1_PDIFF $count=1 $X=3.44
+ $Y=1.745 $X2=3.58 $Y2=2.2
r87 3 29 400 $w=1.7e-07 $l=1.20297e-06 $layer=licon1_PDIFF $count=1 $X=3.44
+ $Y=1.745 $X2=3.58 $Y2=2.88
r88 2 23 400 $w=1.7e-07 $l=1.20297e-06 $layer=licon1_PDIFF $count=1 $X=2.58
+ $Y=1.745 $X2=2.72 $Y2=2.88
r89 2 20 400 $w=1.7e-07 $l=4.29331e-07 $layer=licon1_PDIFF $count=1 $X=2.58
+ $Y=1.745 $X2=2.72 $Y2=2.11
r90 1 41 600 $w=1.7e-07 $l=1.11074e-06 $layer=licon1_PDIFF $count=1 $X=1.735
+ $Y=1.745 $X2=1.86 $Y2=2.795
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4BB_4%Y 1 2 3 4 5 6 7 8 9 10 33 37 41 42 43 44 47
+ 51 55 57 61 67 68 71 73 74 77 79 83 85 89 91 95 97 98 103 104 105 106 107 111
+ 116
c174 74 0 5.06642e-20 $X=5.615 $Y=1.08
r175 111 116 0.631476 $w=3.63e-07 $l=2e-08 $layer=LI1_cond $X=5.432 $Y=1.685
+ $X2=5.432 $Y2=1.665
r176 107 111 2.61117 $w=3.65e-07 $l=9e-08 $layer=LI1_cond $X=5.432 $Y=1.775
+ $X2=5.432 $Y2=1.685
r177 107 116 1.04193 $w=3.63e-07 $l=3.3e-08 $layer=LI1_cond $X=5.432 $Y=1.632
+ $X2=5.432 $Y2=1.665
r178 106 107 10.6404 $w=3.63e-07 $l=3.37e-07 $layer=LI1_cond $X=5.432 $Y=1.295
+ $X2=5.432 $Y2=1.632
r179 102 106 3.78885 $w=3.63e-07 $l=1.2e-07 $layer=LI1_cond $X=5.432 $Y=1.175
+ $X2=5.432 $Y2=1.295
r180 100 102 27.8292 $w=1.85e-07 $l=4.22e-07 $layer=LI1_cond $X=5.01 $Y=1.08
+ $X2=5.432 $Y2=1.08
r181 93 95 29.9635 $w=2.23e-07 $l=5.85e-07 $layer=LI1_cond $X=8.852 $Y=1.005
+ $X2=8.852 $Y2=0.42
r182 92 105 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=8.07 $Y=1.09
+ $X2=7.975 $Y2=1.09
r183 91 93 6.9898 $w=1.7e-07 $l=1.4854e-07 $layer=LI1_cond $X=8.74 $Y=1.09
+ $X2=8.852 $Y2=1.005
r184 91 92 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=8.74 $Y=1.09
+ $X2=8.07 $Y2=1.09
r185 87 105 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=7.975 $Y=1.005
+ $X2=7.975 $Y2=1.09
r186 87 89 34.1483 $w=1.88e-07 $l=5.85e-07 $layer=LI1_cond $X=7.975 $Y=1.005
+ $X2=7.975 $Y2=0.42
r187 86 104 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=7.21 $Y=1.09
+ $X2=7.115 $Y2=1.09
r188 85 105 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=7.88 $Y=1.09
+ $X2=7.975 $Y2=1.09
r189 85 86 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=7.88 $Y=1.09
+ $X2=7.21 $Y2=1.09
r190 81 104 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=7.115 $Y=1.005
+ $X2=7.115 $Y2=1.09
r191 81 83 34.1483 $w=1.88e-07 $l=5.85e-07 $layer=LI1_cond $X=7.115 $Y=1.005
+ $X2=7.115 $Y2=0.42
r192 80 103 5.40251 $w=1.8e-07 $l=9.98749e-08 $layer=LI1_cond $X=6.35 $Y=1.09
+ $X2=6.255 $Y2=1.08
r193 79 104 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=7.02 $Y=1.09
+ $X2=7.115 $Y2=1.09
r194 79 80 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=7.02 $Y=1.09
+ $X2=6.35 $Y2=1.09
r195 75 103 1.14861 $w=1.9e-07 $l=9.5e-08 $layer=LI1_cond $X=6.255 $Y=0.985
+ $X2=6.255 $Y2=1.08
r196 75 77 32.9809 $w=1.88e-07 $l=5.65e-07 $layer=LI1_cond $X=6.255 $Y=0.985
+ $X2=6.255 $Y2=0.42
r197 74 102 11.7505 $w=1.9e-07 $l=1.83e-07 $layer=LI1_cond $X=5.615 $Y=1.08
+ $X2=5.432 $Y2=1.08
r198 73 103 5.40251 $w=1.8e-07 $l=9.5e-08 $layer=LI1_cond $X=6.16 $Y=1.08
+ $X2=6.255 $Y2=1.08
r199 73 74 31.8134 $w=1.88e-07 $l=5.45e-07 $layer=LI1_cond $X=6.16 $Y=1.08
+ $X2=5.615 $Y2=1.08
r200 69 100 0.553203 $w=1.9e-07 $l=9.5e-08 $layer=LI1_cond $X=5.01 $Y=0.985
+ $X2=5.01 $Y2=1.08
r201 69 71 32.9809 $w=1.88e-07 $l=5.65e-07 $layer=LI1_cond $X=5.01 $Y=0.985
+ $X2=5.01 $Y2=0.42
r202 67 100 6.36665 $w=1.85e-07 $l=9.5e-08 $layer=LI1_cond $X=4.915 $Y=1.08
+ $X2=5.01 $Y2=1.08
r203 67 68 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.915 $Y=1.08
+ $X2=4.245 $Y2=1.08
r204 64 68 6.83233 $w=1.7e-07 $l=1.28662e-07 $layer=LI1_cond $X=4.152 $Y=0.995
+ $X2=4.245 $Y2=1.08
r205 64 66 3.89681 $w=1.83e-07 $l=6.5e-08 $layer=LI1_cond $X=4.152 $Y=0.995
+ $X2=4.152 $Y2=0.93
r206 63 99 4.7579 $w=1.87e-07 $l=8.59942e-08 $layer=LI1_cond $X=4.152 $Y=0.825
+ $X2=4.15 $Y2=0.74
r207 63 66 6.29484 $w=1.83e-07 $l=1.05e-07 $layer=LI1_cond $X=4.152 $Y=0.825
+ $X2=4.152 $Y2=0.93
r208 59 99 4.7579 $w=1.87e-07 $l=8.5e-08 $layer=LI1_cond $X=4.15 $Y=0.655
+ $X2=4.15 $Y2=0.74
r209 59 61 13.7177 $w=1.88e-07 $l=2.35e-07 $layer=LI1_cond $X=4.15 $Y=0.655
+ $X2=4.15 $Y2=0.42
r210 58 97 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.385 $Y=0.74
+ $X2=3.22 $Y2=0.74
r211 57 99 1.69765 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=4.055 $Y=0.74
+ $X2=4.15 $Y2=0.74
r212 57 58 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.055 $Y=0.74
+ $X2=3.385 $Y2=0.74
r213 56 98 6.44382 $w=1.75e-07 $l=1.15e-07 $layer=LI1_cond $X=3.285 $Y=1.775
+ $X2=3.17 $Y2=1.775
r214 55 107 5.28037 $w=1.8e-07 $l=1.82e-07 $layer=LI1_cond $X=5.25 $Y=1.775
+ $X2=5.432 $Y2=1.775
r215 55 56 121.076 $w=1.78e-07 $l=1.965e-06 $layer=LI1_cond $X=5.25 $Y=1.775
+ $X2=3.285 $Y2=1.775
r216 51 53 35.0744 $w=2.28e-07 $l=7e-07 $layer=LI1_cond $X=3.17 $Y=1.87 $X2=3.17
+ $Y2=2.57
r217 49 98 0.379591 $w=2.3e-07 $l=9e-08 $layer=LI1_cond $X=3.17 $Y=1.865
+ $X2=3.17 $Y2=1.775
r218 49 51 0.250531 $w=2.28e-07 $l=5e-09 $layer=LI1_cond $X=3.17 $Y=1.865
+ $X2=3.17 $Y2=1.87
r219 45 97 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.22 $Y=0.655
+ $X2=3.22 $Y2=0.74
r220 45 47 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=3.22 $Y=0.655
+ $X2=3.22 $Y2=0.36
r221 43 98 6.44382 $w=1.75e-07 $l=1.17473e-07 $layer=LI1_cond $X=3.055 $Y=1.77
+ $X2=3.17 $Y2=1.775
r222 43 44 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.055 $Y=1.77
+ $X2=2.385 $Y2=1.77
r223 41 97 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.055 $Y=0.74
+ $X2=3.22 $Y2=0.74
r224 41 42 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.055 $Y=0.74
+ $X2=2.365 $Y2=0.74
r225 37 39 40.8612 $w=1.88e-07 $l=7e-07 $layer=LI1_cond $X=2.29 $Y=1.87 $X2=2.29
+ $Y2=2.57
r226 35 44 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=2.29 $Y=1.855
+ $X2=2.385 $Y2=1.77
r227 35 37 0.875598 $w=1.88e-07 $l=1.5e-08 $layer=LI1_cond $X=2.29 $Y=1.855
+ $X2=2.29 $Y2=1.87
r228 31 42 7.85115 $w=1.7e-07 $l=2.08207e-07 $layer=LI1_cond $X=2.195 $Y=0.655
+ $X2=2.365 $Y2=0.74
r229 31 33 9.99914 $w=3.38e-07 $l=2.95e-07 $layer=LI1_cond $X=2.195 $Y=0.655
+ $X2=2.195 $Y2=0.36
r230 10 53 400 $w=1.7e-07 $l=8.92258e-07 $layer=licon1_PDIFF $count=1 $X=3.01
+ $Y=1.745 $X2=3.15 $Y2=2.57
r231 10 51 400 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=3.01
+ $Y=1.745 $X2=3.15 $Y2=1.87
r232 9 39 400 $w=1.7e-07 $l=8.92258e-07 $layer=licon1_PDIFF $count=1 $X=2.15
+ $Y=1.745 $X2=2.29 $Y2=2.57
r233 9 37 400 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=2.15
+ $Y=1.745 $X2=2.29 $Y2=1.87
r234 8 95 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=8.695
+ $Y=0.235 $X2=8.835 $Y2=0.42
r235 7 89 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=7.835
+ $Y=0.235 $X2=7.975 $Y2=0.42
r236 6 83 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=6.975
+ $Y=0.235 $X2=7.115 $Y2=0.42
r237 5 77 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=6.115
+ $Y=0.235 $X2=6.255 $Y2=0.42
r238 4 71 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=4.87
+ $Y=0.235 $X2=5.01 $Y2=0.42
r239 3 66 182 $w=1.7e-07 $l=7.61791e-07 $layer=licon1_NDIFF $count=1 $X=4.01
+ $Y=0.235 $X2=4.15 $Y2=0.93
r240 3 61 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=4.01
+ $Y=0.235 $X2=4.15 $Y2=0.42
r241 2 47 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=3.08
+ $Y=0.235 $X2=3.22 $Y2=0.36
r242 1 33 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=2.05
+ $Y=0.235 $X2=2.19 $Y2=0.36
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4BB_4%A_774_349# 1 2 3 4 15 17 18 21 23 27 29 31
+ 33 35 36
c65 35 0 5.86634e-20 $X=4.87 $Y=2.98
c66 18 0 7.76303e-20 $X=4.175 $Y=2.99
r67 31 38 2.73294 $w=3.3e-07 $l=9.5e-08 $layer=LI1_cond $X=7.11 $Y=2.885
+ $X2=7.11 $Y2=2.98
r68 31 33 26.0173 $w=3.28e-07 $l=7.45e-07 $layer=LI1_cond $X=7.11 $Y=2.885
+ $X2=7.11 $Y2=2.14
r69 30 36 7.95398 $w=1.9e-07 $l=1.65e-07 $layer=LI1_cond $X=6.415 $Y=2.98
+ $X2=6.25 $Y2=2.98
r70 29 38 4.74669 $w=1.9e-07 $l=1.65e-07 $layer=LI1_cond $X=6.945 $Y=2.98
+ $X2=7.11 $Y2=2.98
r71 29 30 30.9378 $w=1.88e-07 $l=5.3e-07 $layer=LI1_cond $X=6.945 $Y=2.98
+ $X2=6.415 $Y2=2.98
r72 25 36 0.546715 $w=3.3e-07 $l=9.5e-08 $layer=LI1_cond $X=6.25 $Y=2.885
+ $X2=6.25 $Y2=2.98
r73 25 27 13.7944 $w=3.28e-07 $l=3.95e-07 $layer=LI1_cond $X=6.25 $Y=2.885
+ $X2=6.25 $Y2=2.49
r74 24 35 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=5.035 $Y=2.98
+ $X2=4.87 $Y2=2.98
r75 23 36 7.95398 $w=1.9e-07 $l=1.65e-07 $layer=LI1_cond $X=6.085 $Y=2.98
+ $X2=6.25 $Y2=2.98
r76 23 24 61.2919 $w=1.88e-07 $l=1.05e-06 $layer=LI1_cond $X=6.085 $Y=2.98
+ $X2=5.035 $Y2=2.98
r77 19 35 0.718145 $w=3.3e-07 $l=9.5e-08 $layer=LI1_cond $X=4.87 $Y=2.885
+ $X2=4.87 $Y2=2.98
r78 19 21 14.1436 $w=3.28e-07 $l=4.05e-07 $layer=LI1_cond $X=4.87 $Y=2.885
+ $X2=4.87 $Y2=2.48
r79 17 35 8.26956 $w=1.8e-07 $l=1.69926e-07 $layer=LI1_cond $X=4.705 $Y=2.99
+ $X2=4.87 $Y2=2.98
r80 17 18 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=4.705 $Y=2.99
+ $X2=4.175 $Y2=2.99
r81 13 18 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.01 $Y=2.905
+ $X2=4.175 $Y2=2.99
r82 13 15 14.8421 $w=3.28e-07 $l=4.25e-07 $layer=LI1_cond $X=4.01 $Y=2.905
+ $X2=4.01 $Y2=2.48
r83 4 38 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=6.97
+ $Y=1.835 $X2=7.11 $Y2=2.91
r84 4 33 400 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_PDIFF $count=1 $X=6.97
+ $Y=1.835 $X2=7.11 $Y2=2.14
r85 3 27 300 $w=1.7e-07 $l=7.21613e-07 $layer=licon1_PDIFF $count=2 $X=6.11
+ $Y=1.835 $X2=6.25 $Y2=2.49
r86 2 21 300 $w=1.7e-07 $l=8.01951e-07 $layer=licon1_PDIFF $count=2 $X=4.73
+ $Y=1.745 $X2=4.87 $Y2=2.48
r87 1 15 300 $w=1.7e-07 $l=8.01951e-07 $layer=licon1_PDIFF $count=2 $X=3.87
+ $Y=1.745 $X2=4.01 $Y2=2.48
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4BB_4%A_1139_367# 1 2 3 4 5 16 18 20 25 28 30 31
+ 32 34 36 40 42 44 46 50 56
r68 53 54 2.2957 $w=1.86e-07 $l=3.5e-08 $layer=LI1_cond $X=7.542 $Y=1.98
+ $X2=7.542 $Y2=2.015
r69 51 53 12.4624 $w=1.86e-07 $l=1.9e-07 $layer=LI1_cond $X=7.542 $Y=1.79
+ $X2=7.542 $Y2=1.98
r70 44 58 2.85134 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=9.3 $Y=2.1 $X2=9.3
+ $Y2=2.015
r71 44 46 17.2866 $w=2.58e-07 $l=3.9e-07 $layer=LI1_cond $X=9.3 $Y=2.1 $X2=9.3
+ $Y2=2.49
r72 43 56 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=8.5 $Y=2.015
+ $X2=8.405 $Y2=2.015
r73 42 58 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=9.17 $Y=2.015 $X2=9.3
+ $Y2=2.015
r74 42 43 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=9.17 $Y=2.015
+ $X2=8.5 $Y2=2.015
r75 38 56 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=8.405 $Y=2.1
+ $X2=8.405 $Y2=2.015
r76 38 40 22.7656 $w=1.88e-07 $l=3.9e-07 $layer=LI1_cond $X=8.405 $Y=2.1
+ $X2=8.405 $Y2=2.49
r77 37 54 1.25915 $w=1.7e-07 $l=9.8e-08 $layer=LI1_cond $X=7.64 $Y=2.015
+ $X2=7.542 $Y2=2.015
r78 36 56 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=8.31 $Y=2.015
+ $X2=8.405 $Y2=2.015
r79 36 37 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=8.31 $Y=2.015
+ $X2=7.64 $Y2=2.015
r80 32 54 5.31795 $w=1.95e-07 $l=8.5e-08 $layer=LI1_cond $X=7.542 $Y=2.1
+ $X2=7.542 $Y2=2.015
r81 32 34 20.7599 $w=1.93e-07 $l=3.65e-07 $layer=LI1_cond $X=7.542 $Y=2.1
+ $X2=7.542 $Y2=2.465
r82 30 51 1.25915 $w=1.7e-07 $l=9.7e-08 $layer=LI1_cond $X=7.445 $Y=1.79
+ $X2=7.542 $Y2=1.79
r83 30 31 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=7.445 $Y=1.79
+ $X2=6.775 $Y2=1.79
r84 26 50 4.06715 $w=2.25e-07 $l=1.00995e-07 $layer=LI1_cond $X=6.68 $Y=2.205
+ $X2=6.645 $Y2=2.12
r85 26 28 20.1388 $w=1.88e-07 $l=3.45e-07 $layer=LI1_cond $X=6.68 $Y=2.205
+ $X2=6.68 $Y2=2.55
r86 23 50 4.06715 $w=2.25e-07 $l=8.5e-08 $layer=LI1_cond $X=6.645 $Y=2.035
+ $X2=6.645 $Y2=2.12
r87 23 25 2.43786 $w=2.58e-07 $l=5.5e-08 $layer=LI1_cond $X=6.645 $Y=2.035
+ $X2=6.645 $Y2=1.98
r88 22 31 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=6.645 $Y=1.875
+ $X2=6.775 $Y2=1.79
r89 22 25 4.6541 $w=2.58e-07 $l=1.05e-07 $layer=LI1_cond $X=6.645 $Y=1.875
+ $X2=6.645 $Y2=1.98
r90 21 49 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=5.915 $Y=2.12
+ $X2=5.785 $Y2=2.12
r91 20 50 2.36881 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=6.515 $Y=2.12
+ $X2=6.645 $Y2=2.12
r92 20 21 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=6.515 $Y=2.12
+ $X2=5.915 $Y2=2.12
r93 16 49 2.85134 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=5.785 $Y=2.205
+ $X2=5.785 $Y2=2.12
r94 16 18 14.8488 $w=2.58e-07 $l=3.35e-07 $layer=LI1_cond $X=5.785 $Y=2.205
+ $X2=5.785 $Y2=2.54
r95 5 58 600 $w=1.7e-07 $l=2.4e-07 $layer=licon1_PDIFF $count=1 $X=9.125
+ $Y=1.835 $X2=9.265 $Y2=2.015
r96 5 46 300 $w=1.7e-07 $l=7.21613e-07 $layer=licon1_PDIFF $count=2 $X=9.125
+ $Y=1.835 $X2=9.265 $Y2=2.49
r97 4 56 600 $w=1.7e-07 $l=2.4e-07 $layer=licon1_PDIFF $count=1 $X=8.265
+ $Y=1.835 $X2=8.405 $Y2=2.015
r98 4 40 300 $w=1.7e-07 $l=7.21613e-07 $layer=licon1_PDIFF $count=2 $X=8.265
+ $Y=1.835 $X2=8.405 $Y2=2.49
r99 3 53 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=7.4
+ $Y=1.835 $X2=7.54 $Y2=1.98
r100 3 34 300 $w=1.7e-07 $l=6.96491e-07 $layer=licon1_PDIFF $count=2 $X=7.4
+ $Y=1.835 $X2=7.54 $Y2=2.465
r101 2 28 600 $w=1.7e-07 $l=7.81873e-07 $layer=licon1_PDIFF $count=1 $X=6.54
+ $Y=1.835 $X2=6.68 $Y2=2.55
r102 2 25 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=6.54
+ $Y=1.835 $X2=6.68 $Y2=1.98
r103 1 49 600 $w=1.7e-07 $l=3.41833e-07 $layer=licon1_PDIFF $count=1 $X=5.695
+ $Y=1.835 $X2=5.82 $Y2=2.12
r104 1 18 600 $w=1.7e-07 $l=7.64951e-07 $layer=licon1_PDIFF $count=1 $X=5.695
+ $Y=1.835 $X2=5.82 $Y2=2.54
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4BB_4%VGND 1 2 3 4 5 6 7 8 9 10 33 37 41 43 47 51
+ 55 59 61 65 69 71 73 75 76 77 79 84 89 94 99 108 113 119 122 125 128 131 134
+ 137 140 144
r159 143 144 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=0
+ $X2=9.36 $Y2=0
r160 140 141 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r161 137 138 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=0
+ $X2=7.44 $Y2=0
r162 134 135 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0
+ $X2=5.52 $Y2=0
r163 131 132 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=0
+ $X2=4.56 $Y2=0
r164 128 129 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r165 126 129 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0
+ $X2=3.6 $Y2=0
r166 125 126 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0
+ $X2=2.64 $Y2=0
r167 122 123 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0
+ $X2=1.68 $Y2=0
r168 119 120 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0
+ $X2=0.72 $Y2=0
r169 117 144 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=0
+ $X2=9.36 $Y2=0
r170 117 141 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=0
+ $X2=8.4 $Y2=0
r171 116 117 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=0
+ $X2=8.88 $Y2=0
r172 114 140 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.57 $Y=0
+ $X2=8.405 $Y2=0
r173 114 116 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=8.57 $Y=0
+ $X2=8.88 $Y2=0
r174 113 143 4.31539 $w=1.7e-07 $l=2.32e-07 $layer=LI1_cond $X=9.135 $Y=0
+ $X2=9.367 $Y2=0
r175 113 116 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=9.135 $Y=0
+ $X2=8.88 $Y2=0
r176 112 141 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0
+ $X2=8.4 $Y2=0
r177 112 138 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0
+ $X2=7.44 $Y2=0
r178 111 112 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=0
+ $X2=7.92 $Y2=0
r179 109 137 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.71 $Y=0
+ $X2=7.545 $Y2=0
r180 109 111 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=7.71 $Y=0
+ $X2=7.92 $Y2=0
r181 108 140 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.24 $Y=0
+ $X2=8.405 $Y2=0
r182 108 111 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=8.24 $Y=0 $X2=7.92
+ $Y2=0
r183 107 138 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.48 $Y=0
+ $X2=7.44 $Y2=0
r184 107 135 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.48 $Y=0
+ $X2=5.52 $Y2=0
r185 106 107 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=0
+ $X2=6.48 $Y2=0
r186 104 134 13.8148 $w=1.7e-07 $l=3.58e-07 $layer=LI1_cond $X=5.99 $Y=0
+ $X2=5.632 $Y2=0
r187 104 106 31.9679 $w=1.68e-07 $l=4.9e-07 $layer=LI1_cond $X=5.99 $Y=0
+ $X2=6.48 $Y2=0
r188 103 135 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0
+ $X2=5.52 $Y2=0
r189 102 103 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0
+ $X2=5.04 $Y2=0
r190 100 131 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.745 $Y=0
+ $X2=4.58 $Y2=0
r191 100 102 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=4.745 $Y=0
+ $X2=5.04 $Y2=0
r192 99 134 13.8148 $w=1.7e-07 $l=3.57e-07 $layer=LI1_cond $X=5.275 $Y=0
+ $X2=5.632 $Y2=0
r193 99 102 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=5.275 $Y=0
+ $X2=5.04 $Y2=0
r194 98 132 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0
+ $X2=4.56 $Y2=0
r195 98 129 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.6
+ $Y2=0
r196 97 98 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r197 95 128 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.885 $Y=0
+ $X2=3.72 $Y2=0
r198 95 97 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=3.885 $Y=0
+ $X2=4.08 $Y2=0
r199 94 131 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.415 $Y=0
+ $X2=4.58 $Y2=0
r200 94 97 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=4.415 $Y=0
+ $X2=4.08 $Y2=0
r201 93 126 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0
+ $X2=2.64 $Y2=0
r202 93 123 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0
+ $X2=1.68 $Y2=0
r203 92 93 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r204 90 122 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.855 $Y=0
+ $X2=1.69 $Y2=0
r205 90 92 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.855 $Y=0
+ $X2=2.16 $Y2=0
r206 89 125 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.535 $Y=0 $X2=2.7
+ $Y2=0
r207 89 92 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=2.535 $Y=0
+ $X2=2.16 $Y2=0
r208 88 123 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r209 88 120 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r210 87 88 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r211 85 119 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.905 $Y=0
+ $X2=0.74 $Y2=0
r212 85 87 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.905 $Y=0 $X2=1.2
+ $Y2=0
r213 84 122 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.525 $Y=0
+ $X2=1.69 $Y2=0
r214 84 87 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=1.525 $Y=0 $X2=1.2
+ $Y2=0
r215 82 120 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0
+ $X2=0.72 $Y2=0
r216 81 82 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r217 79 119 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.575 $Y=0
+ $X2=0.74 $Y2=0
r218 79 81 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=0.575 $Y=0
+ $X2=0.24 $Y2=0
r219 77 103 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.8 $Y=0
+ $X2=5.04 $Y2=0
r220 77 132 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.8 $Y=0
+ $X2=4.56 $Y2=0
r221 75 106 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=6.52 $Y=0 $X2=6.48
+ $Y2=0
r222 75 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.52 $Y=0 $X2=6.685
+ $Y2=0
r223 71 143 3.16214 $w=2.95e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.282 $Y=0.085
+ $X2=9.367 $Y2=0
r224 71 73 11.5244 $w=2.93e-07 $l=2.95e-07 $layer=LI1_cond $X=9.282 $Y=0.085
+ $X2=9.282 $Y2=0.38
r225 67 140 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.405 $Y=0.085
+ $X2=8.405 $Y2=0
r226 67 69 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=8.405 $Y=0.085
+ $X2=8.405 $Y2=0.38
r227 63 137 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.545 $Y=0.085
+ $X2=7.545 $Y2=0
r228 63 65 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=7.545 $Y=0.085
+ $X2=7.545 $Y2=0.38
r229 62 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.85 $Y=0 $X2=6.685
+ $Y2=0
r230 61 137 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.38 $Y=0
+ $X2=7.545 $Y2=0
r231 61 62 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=7.38 $Y=0 $X2=6.85
+ $Y2=0
r232 57 76 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.685 $Y=0.085
+ $X2=6.685 $Y2=0
r233 57 59 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=6.685 $Y=0.085
+ $X2=6.685 $Y2=0.38
r234 53 134 2.90666 $w=7.15e-07 $l=8.5e-08 $layer=LI1_cond $X=5.632 $Y=0.085
+ $X2=5.632 $Y2=0
r235 53 55 4.6003 $w=7.13e-07 $l=2.75e-07 $layer=LI1_cond $X=5.632 $Y=0.085
+ $X2=5.632 $Y2=0.36
r236 49 131 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.58 $Y=0.085
+ $X2=4.58 $Y2=0
r237 49 51 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=4.58 $Y=0.085
+ $X2=4.58 $Y2=0.36
r238 45 128 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.72 $Y=0.085
+ $X2=3.72 $Y2=0
r239 45 47 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=3.72 $Y=0.085
+ $X2=3.72 $Y2=0.36
r240 44 125 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.865 $Y=0 $X2=2.7
+ $Y2=0
r241 43 128 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.555 $Y=0
+ $X2=3.72 $Y2=0
r242 43 44 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.555 $Y=0 $X2=2.865
+ $Y2=0
r243 39 125 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.7 $Y=0.085
+ $X2=2.7 $Y2=0
r244 39 41 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.7 $Y=0.085
+ $X2=2.7 $Y2=0.36
r245 35 122 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.69 $Y=0.085
+ $X2=1.69 $Y2=0
r246 35 37 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.69 $Y=0.085
+ $X2=1.69 $Y2=0.38
r247 31 119 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.74 $Y=0.085
+ $X2=0.74 $Y2=0
r248 31 33 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=0.74 $Y=0.085
+ $X2=0.74 $Y2=0.4
r249 10 73 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=9.125
+ $Y=0.235 $X2=9.265 $Y2=0.38
r250 9 69 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=8.265
+ $Y=0.235 $X2=8.405 $Y2=0.38
r251 8 65 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=7.405
+ $Y=0.235 $X2=7.545 $Y2=0.38
r252 7 59 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.545
+ $Y=0.235 $X2=6.685 $Y2=0.38
r253 6 55 45.5 $w=1.7e-07 $l=5.84166e-07 $layer=licon1_NDIFF $count=4 $X=5.3
+ $Y=0.235 $X2=5.825 $Y2=0.36
r254 5 51 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=4.44
+ $Y=0.235 $X2=4.58 $Y2=0.36
r255 4 47 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=3.51
+ $Y=0.235 $X2=3.72 $Y2=0.36
r256 3 41 182 $w=1.7e-07 $l=2.755e-07 $layer=licon1_NDIFF $count=1 $X=2.48
+ $Y=0.235 $X2=2.7 $Y2=0.36
r257 2 37 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=1.565
+ $Y=0.235 $X2=1.69 $Y2=0.38
r258 1 33 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=0.6
+ $Y=0.255 $X2=0.74 $Y2=0.4
.ends

