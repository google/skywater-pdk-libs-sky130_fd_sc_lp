* File: sky130_fd_sc_lp__o21ba_0.pex.spice
* Created: Fri Aug 28 11:05:28 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O21BA_0%A_80_225# 1 2 8 11 15 17 20 21 23 24 26 28
+ 31 36 38
c88 38 0 1.3023e-19 $X=2.495 $Y=2.57
r89 35 38 13.3491 $w=2.38e-07 $l=2.78e-07 $layer=LI1_cond $X=2.217 $Y=2.515
+ $X2=2.495 $Y2=2.515
r90 35 36 6.61396 $w=2.38e-07 $l=1.17e-07 $layer=LI1_cond $X=2.217 $Y=2.515
+ $X2=2.1 $Y2=2.515
r91 29 35 0.869974 $w=2.35e-07 $l=1.2e-07 $layer=LI1_cond $X=2.217 $Y=2.395
+ $X2=2.217 $Y2=2.515
r92 29 31 95.6283 $w=2.33e-07 $l=1.95e-06 $layer=LI1_cond $X=2.217 $Y=2.395
+ $X2=2.217 $Y2=0.445
r93 28 36 62.3048 $w=1.68e-07 $l=9.55e-07 $layer=LI1_cond $X=1.145 $Y=2.55
+ $X2=2.1 $Y2=2.55
r94 26 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.06 $Y=2.465
+ $X2=1.145 $Y2=2.55
r95 25 26 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.06 $Y=1.795
+ $X2=1.06 $Y2=2.465
r96 23 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.975 $Y=1.71
+ $X2=1.06 $Y2=1.795
r97 23 24 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=0.975 $Y=1.71
+ $X2=0.755 $Y2=1.71
r98 21 41 46.504 $w=3.55e-07 $l=1.65e-07 $layer=POLY_cond $X=0.577 $Y=1.29
+ $X2=0.577 $Y2=1.125
r99 20 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.59
+ $Y=1.29 $X2=0.59 $Y2=1.29
r100 18 24 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.63 $Y=1.625
+ $X2=0.755 $Y2=1.71
r101 18 20 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=0.63 $Y=1.625
+ $X2=0.63 $Y2=1.29
r102 15 41 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=0.585 $Y=0.445
+ $X2=0.585 $Y2=1.125
r103 11 17 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=0.475 $Y=2.305
+ $X2=0.475 $Y2=1.795
r104 8 17 48.4546 $w=3.55e-07 $l=1.77e-07 $layer=POLY_cond $X=0.577 $Y=1.618
+ $X2=0.577 $Y2=1.795
r105 7 21 1.95057 $w=3.55e-07 $l=1.2e-08 $layer=POLY_cond $X=0.577 $Y=1.302
+ $X2=0.577 $Y2=1.29
r106 7 8 51.3649 $w=3.55e-07 $l=3.16e-07 $layer=POLY_cond $X=0.577 $Y=1.302
+ $X2=0.577 $Y2=1.618
r107 2 38 300 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_PDIFF $count=2 $X=2.355
+ $Y=2.435 $X2=2.495 $Y2=2.57
r108 1 31 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=2.08
+ $Y=0.235 $X2=2.205 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__O21BA_0%B1_N 2 5 9 10 11 12 16 18
r41 16 18 45.5639 $w=3.95e-07 $l=1.65e-07 $layer=POLY_cond $X=1.232 $Y=0.93
+ $X2=1.232 $Y2=0.765
r42 11 12 13.755 $w=3.08e-07 $l=3.7e-07 $layer=LI1_cond $X=1.15 $Y=0.925
+ $X2=1.15 $Y2=1.295
r43 11 16 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.2 $Y=0.93
+ $X2=1.2 $Y2=0.93
r44 9 18 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.355 $Y=0.445
+ $X2=1.355 $Y2=0.765
r45 5 10 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=1.215 $Y=2.195
+ $X2=1.215 $Y2=1.435
r46 2 10 39.7623 $w=3.95e-07 $l=1.97e-07 $layer=POLY_cond $X=1.232 $Y=1.238
+ $X2=1.232 $Y2=1.435
r47 1 16 4.50555 $w=3.95e-07 $l=3.2e-08 $layer=POLY_cond $X=1.232 $Y=0.962
+ $X2=1.232 $Y2=0.93
r48 1 2 38.8604 $w=3.95e-07 $l=2.76e-07 $layer=POLY_cond $X=1.232 $Y=0.962
+ $X2=1.232 $Y2=1.238
.ends

.subckt PM_SKY130_FD_SC_LP__O21BA_0%A_258_397# 1 2 7 9 11 13 16 19 23 26
r49 26 29 15.1331 $w=4.53e-07 $l=5.05e-07 $layer=LI1_cond $X=1.702 $Y=1.03
+ $X2=1.702 $Y2=1.535
r50 26 28 6.51597 $w=4.53e-07 $l=1.65e-07 $layer=LI1_cond $X=1.702 $Y=1.03
+ $X2=1.702 $Y2=0.865
r51 26 27 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.835
+ $Y=1.03 $X2=1.835 $Y2=1.03
r52 21 23 6.3559 $w=3.28e-07 $l=1.82e-07 $layer=LI1_cond $X=1.43 $Y=2.13
+ $X2=1.612 $Y2=2.13
r53 19 23 1.82517 $w=2.75e-07 $l=1.65e-07 $layer=LI1_cond $X=1.612 $Y=1.965
+ $X2=1.612 $Y2=2.13
r54 19 29 18.02 $w=2.73e-07 $l=4.3e-07 $layer=LI1_cond $X=1.612 $Y=1.965
+ $X2=1.612 $Y2=1.535
r55 16 28 18.6164 $w=2.58e-07 $l=4.2e-07 $layer=LI1_cond $X=1.605 $Y=0.445
+ $X2=1.605 $Y2=0.865
r56 11 27 53.2183 $w=6.42e-07 $l=4.51458e-07 $layer=POLY_cond $X=2.42 $Y=0.765
+ $X2=2.082 $Y2=1.03
r57 11 13 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.42 $Y=0.765
+ $X2=2.42 $Y2=0.445
r58 7 27 71.237 $w=6.42e-07 $l=5.95831e-07 $layer=POLY_cond $X=2.28 $Y=1.535
+ $X2=2.082 $Y2=1.03
r59 7 9 625.574 $w=1.5e-07 $l=1.22e-06 $layer=POLY_cond $X=2.28 $Y=1.535
+ $X2=2.28 $Y2=2.755
r60 2 21 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.29
+ $Y=1.985 $X2=1.43 $Y2=2.13
r61 1 16 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.43
+ $Y=0.235 $X2=1.57 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__O21BA_0%A2 3 7 11 12 13 14 15 20
c43 20 0 6.29351e-20 $X=2.76 $Y=1.32
c44 12 0 1.3023e-19 $X=2.76 $Y=1.825
c45 11 0 1.4009e-19 $X=2.76 $Y=1.66
r46 20 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.76
+ $Y=1.32 $X2=2.76 $Y2=1.32
r47 14 15 12.5413 $w=3.38e-07 $l=3.7e-07 $layer=LI1_cond $X=2.675 $Y=1.665
+ $X2=2.675 $Y2=2.035
r48 14 21 11.6939 $w=3.38e-07 $l=3.45e-07 $layer=LI1_cond $X=2.675 $Y=1.665
+ $X2=2.675 $Y2=1.32
r49 13 21 0.847385 $w=3.38e-07 $l=2.5e-08 $layer=LI1_cond $X=2.675 $Y=1.295
+ $X2=2.675 $Y2=1.32
r50 11 20 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.76 $Y=1.66
+ $X2=2.76 $Y2=1.32
r51 11 12 40.8701 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.76 $Y=1.66
+ $X2=2.76 $Y2=1.825
r52 10 20 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.76 $Y=1.155
+ $X2=2.76 $Y2=1.32
r53 7 10 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=2.85 $Y=0.445
+ $X2=2.85 $Y2=1.155
r54 3 12 476.872 $w=1.5e-07 $l=9.3e-07 $layer=POLY_cond $X=2.71 $Y=2.755
+ $X2=2.71 $Y2=1.825
.ends

.subckt PM_SKY130_FD_SC_LP__O21BA_0%A1 3 7 10 11 14 15 16 21
r33 21 22 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.33
+ $Y=1.71 $X2=3.33 $Y2=1.71
r34 16 22 7.40429 $w=5.23e-07 $l=3.25e-07 $layer=LI1_cond $X=3.277 $Y=2.035
+ $X2=3.277 $Y2=1.71
r35 15 22 1.02521 $w=5.23e-07 $l=4.5e-08 $layer=LI1_cond $X=3.277 $Y=1.665
+ $X2=3.277 $Y2=1.71
r36 14 15 8.42951 $w=5.23e-07 $l=3.7e-07 $layer=LI1_cond $X=3.277 $Y=1.295
+ $X2=3.277 $Y2=1.665
r37 13 21 40.8701 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.33 $Y=1.545
+ $X2=3.33 $Y2=1.71
r38 10 21 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=3.33 $Y=2.065
+ $X2=3.33 $Y2=1.71
r39 10 11 43.5886 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=3.26 $Y=2.065
+ $X2=3.26 $Y2=2.215
r40 7 13 564.043 $w=1.5e-07 $l=1.1e-06 $layer=POLY_cond $X=3.28 $Y=0.445
+ $X2=3.28 $Y2=1.545
r41 3 11 276.894 $w=1.5e-07 $l=5.4e-07 $layer=POLY_cond $X=3.1 $Y=2.755 $X2=3.1
+ $Y2=2.215
.ends

.subckt PM_SKY130_FD_SC_LP__O21BA_0%X 1 2 7 8 9 10 11 12 13 47 50
r20 50 51 2.64267 $w=2.68e-07 $l=6e-08 $layer=LI1_cond $X=0.22 $Y=2.035 $X2=0.22
+ $Y2=1.975
r21 24 42 2.36532 $w=2.5e-07 $l=1.65e-07 $layer=LI1_cond $X=0.21 $Y=0.61
+ $X2=0.21 $Y2=0.445
r22 12 13 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.22 $Y=2.405
+ $X2=0.22 $Y2=2.775
r23 11 34 2.90245 $w=2.68e-07 $l=6.8e-08 $layer=LI1_cond $X=0.22 $Y=2.042
+ $X2=0.22 $Y2=2.11
r24 11 50 0.298782 $w=2.68e-07 $l=7e-09 $layer=LI1_cond $X=0.22 $Y=2.042
+ $X2=0.22 $Y2=2.035
r25 11 12 12.3781 $w=2.68e-07 $l=2.9e-07 $layer=LI1_cond $X=0.22 $Y=2.115
+ $X2=0.22 $Y2=2.405
r26 11 34 0.213415 $w=2.68e-07 $l=5e-09 $layer=LI1_cond $X=0.22 $Y=2.115
+ $X2=0.22 $Y2=2.11
r27 11 51 0.59927 $w=2.48e-07 $l=1.3e-08 $layer=LI1_cond $X=0.21 $Y=1.962
+ $X2=0.21 $Y2=1.975
r28 10 11 13.691 $w=2.48e-07 $l=2.97e-07 $layer=LI1_cond $X=0.21 $Y=1.665
+ $X2=0.21 $Y2=1.962
r29 9 10 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=0.21 $Y=1.295
+ $X2=0.21 $Y2=1.665
r30 8 9 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=0.21 $Y=0.925 $X2=0.21
+ $Y2=1.295
r31 7 47 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=0.24 $Y=0.445
+ $X2=0.37 $Y2=0.445
r32 7 42 1.04768 $w=3.28e-07 $l=3e-08 $layer=LI1_cond $X=0.24 $Y=0.445 $X2=0.21
+ $Y2=0.445
r33 7 8 13.8293 $w=2.48e-07 $l=3e-07 $layer=LI1_cond $X=0.21 $Y=0.625 $X2=0.21
+ $Y2=0.925
r34 7 24 0.691466 $w=2.48e-07 $l=1.5e-08 $layer=LI1_cond $X=0.21 $Y=0.625
+ $X2=0.21 $Y2=0.61
r35 2 11 300 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.985 $X2=0.26 $Y2=2.14
r36 1 47 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.245
+ $Y=0.235 $X2=0.37 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__O21BA_0%VPWR 1 2 3 12 16 20 23 24 25 27 32 42 43 46
+ 49
r48 49 50 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r49 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r50 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r51 40 43 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r52 40 50 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.16 $Y2=3.33
r53 39 40 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r54 37 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.21 $Y=3.33
+ $X2=2.045 $Y2=3.33
r55 37 39 59.369 $w=1.68e-07 $l=9.1e-07 $layer=LI1_cond $X=2.21 $Y=3.33 $X2=3.12
+ $Y2=3.33
r56 36 47 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.72 $Y2=3.33
r57 35 36 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r58 33 46 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=0.805 $Y=3.33
+ $X2=0.665 $Y2=3.33
r59 33 35 57.0856 $w=1.68e-07 $l=8.75e-07 $layer=LI1_cond $X=0.805 $Y=3.33
+ $X2=1.68 $Y2=3.33
r60 32 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.88 $Y=3.33
+ $X2=2.045 $Y2=3.33
r61 32 35 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=1.88 $Y=3.33 $X2=1.68
+ $Y2=3.33
r62 30 47 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r63 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r64 27 46 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=0.525 $Y=3.33
+ $X2=0.665 $Y2=3.33
r65 27 29 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.525 $Y=3.33
+ $X2=0.24 $Y2=3.33
r66 25 50 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=2.16 $Y2=3.33
r67 25 36 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=1.68 $Y2=3.33
r68 23 39 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=3.15 $Y=3.33 $X2=3.12
+ $Y2=3.33
r69 23 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.15 $Y=3.33
+ $X2=3.315 $Y2=3.33
r70 22 42 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=3.48 $Y=3.33 $X2=3.6
+ $Y2=3.33
r71 22 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.48 $Y=3.33
+ $X2=3.315 $Y2=3.33
r72 18 24 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.315 $Y=3.245
+ $X2=3.315 $Y2=3.33
r73 18 20 23.2235 $w=3.28e-07 $l=6.65e-07 $layer=LI1_cond $X=3.315 $Y=3.245
+ $X2=3.315 $Y2=2.58
r74 14 49 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.045 $Y=3.245
+ $X2=2.045 $Y2=3.33
r75 14 16 11.5244 $w=3.28e-07 $l=3.3e-07 $layer=LI1_cond $X=2.045 $Y=3.245
+ $X2=2.045 $Y2=2.915
r76 10 46 0.375625 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=0.665 $Y=3.245
+ $X2=0.665 $Y2=3.33
r77 10 12 45.8919 $w=2.78e-07 $l=1.115e-06 $layer=LI1_cond $X=0.665 $Y=3.245
+ $X2=0.665 $Y2=2.13
r78 3 20 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=3.175
+ $Y=2.435 $X2=3.315 $Y2=2.58
r79 2 16 600 $w=1.7e-07 $l=5.38888e-07 $layer=licon1_PDIFF $count=1 $X=1.92
+ $Y=2.435 $X2=2.045 $Y2=2.915
r80 1 12 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=0.55
+ $Y=1.985 $X2=0.69 $Y2=2.13
.ends

.subckt PM_SKY130_FD_SC_LP__O21BA_0%VGND 1 2 9 12 13 14 29 30 35 41
r46 39 41 9.621 $w=6.78e-07 $l=1.05e-07 $layer=LI1_cond $X=1.2 $Y=0.255
+ $X2=1.305 $Y2=0.255
r47 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r48 37 39 1.05536 $w=6.78e-07 $l=6e-08 $layer=LI1_cond $X=1.14 $Y=0.255 $X2=1.2
+ $Y2=0.255
r49 34 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r50 33 37 7.38754 $w=6.78e-07 $l=4.2e-07 $layer=LI1_cond $X=0.72 $Y=0.255
+ $X2=1.14 $Y2=0.255
r51 33 35 9.26921 $w=6.78e-07 $l=8.5e-08 $layer=LI1_cond $X=0.72 $Y=0.255
+ $X2=0.635 $Y2=0.255
r52 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r53 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r54 27 30 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r55 26 27 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r56 24 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r57 23 26 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r58 23 41 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.68 $Y=0 $X2=1.305
+ $Y2=0
r59 23 24 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r60 19 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r61 18 35 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=0.24 $Y=0 $X2=0.635
+ $Y2=0
r62 18 19 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r63 14 27 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=2.64
+ $Y2=0
r64 14 24 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=1.68
+ $Y2=0
r65 12 26 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=2.935 $Y=0 $X2=2.64
+ $Y2=0
r66 12 13 7.34436 $w=1.7e-07 $l=1.32e-07 $layer=LI1_cond $X=2.935 $Y=0 $X2=3.067
+ $Y2=0
r67 11 29 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=3.2 $Y=0 $X2=3.6 $Y2=0
r68 11 13 7.34436 $w=1.7e-07 $l=1.33e-07 $layer=LI1_cond $X=3.2 $Y=0 $X2=3.067
+ $Y2=0
r69 7 13 0.195364 $w=2.65e-07 $l=8.5e-08 $layer=LI1_cond $X=3.067 $Y=0.085
+ $X2=3.067 $Y2=0
r70 7 9 15.6558 $w=2.63e-07 $l=3.6e-07 $layer=LI1_cond $X=3.067 $Y=0.085
+ $X2=3.067 $Y2=0.445
r71 2 9 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.925
+ $Y=0.235 $X2=3.065 $Y2=0.445
r72 1 37 91 $w=1.7e-07 $l=5.755e-07 $layer=licon1_NDIFF $count=2 $X=0.66
+ $Y=0.235 $X2=1.14 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__O21BA_0%A_499_47# 1 2 9 11 12 15
c25 11 0 6.29351e-20 $X=3.37 $Y=0.87
r26 13 15 13.3127 $w=2.88e-07 $l=3.35e-07 $layer=LI1_cond $X=3.515 $Y=0.78
+ $X2=3.515 $Y2=0.445
r27 11 13 7.31368 $w=1.8e-07 $l=1.84594e-07 $layer=LI1_cond $X=3.37 $Y=0.87
+ $X2=3.515 $Y2=0.78
r28 11 12 37.2778 $w=1.78e-07 $l=6.05e-07 $layer=LI1_cond $X=3.37 $Y=0.87
+ $X2=2.765 $Y2=0.87
r29 7 12 7.11373 $w=1.8e-07 $l=1.69115e-07 $layer=LI1_cond $X=2.635 $Y=0.78
+ $X2=2.765 $Y2=0.87
r30 7 9 14.8488 $w=2.58e-07 $l=3.35e-07 $layer=LI1_cond $X=2.635 $Y=0.78
+ $X2=2.635 $Y2=0.445
r31 2 15 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=3.355
+ $Y=0.235 $X2=3.495 $Y2=0.445
r32 1 9 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.495
+ $Y=0.235 $X2=2.635 $Y2=0.445
.ends

