* File: sky130_fd_sc_lp__dlybuf4s18kapwr_1.pex.spice
* Created: Wed Sep  2 09:49:18 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__DLYBUF4S18KAPWR_1%A 3 7 9 10 14
c36 9 0 1.45138e-19 $X=0.24 $Y=1.295
r37 14 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.385 $Y=1.5
+ $X2=0.385 $Y2=1.665
r38 14 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.385 $Y=1.5
+ $X2=0.385 $Y2=1.335
r39 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.385
+ $Y=1.5 $X2=0.385 $Y2=1.5
r40 10 15 4.38562 $w=4.48e-07 $l=1.65e-07 $layer=LI1_cond $X=0.325 $Y=1.665
+ $X2=0.325 $Y2=1.5
r41 9 15 5.4488 $w=4.48e-07 $l=2.05e-07 $layer=LI1_cond $X=0.325 $Y=1.295
+ $X2=0.325 $Y2=1.5
r42 7 17 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=0.475 $Y=2.465
+ $X2=0.475 $Y2=1.665
r43 3 16 443.543 $w=1.5e-07 $l=8.65e-07 $layer=POLY_cond $X=0.475 $Y=0.47
+ $X2=0.475 $Y2=1.335
.ends

.subckt PM_SKY130_FD_SC_LP__DLYBUF4S18KAPWR_1%A_27_52# 1 2 7 9 10 12 16 18 20 22
+ 23 24 27 29
c72 27 0 5.13383e-20 $X=1.087 $Y=1.6
c73 10 0 6.01461e-20 $X=1.32 $Y=1.93
c74 7 0 1.45138e-19 $X=1.32 $Y=1.37
r75 29 30 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.085
+ $Y=1.535 $X2=1.085 $Y2=1.535
r76 27 33 13.9394 $w=4.83e-07 $l=5.7297e-07 $layer=LI1_cond $X=1.087 $Y=1.6
+ $X2=1.205 $Y2=2.117
r77 27 29 2.11011 $w=3.53e-07 $l=6.5e-08 $layer=LI1_cond $X=1.087 $Y=1.6
+ $X2=1.087 $Y2=1.535
r78 26 29 16.7185 $w=3.53e-07 $l=5.15e-07 $layer=LI1_cond $X=1.087 $Y=1.02
+ $X2=1.087 $Y2=1.535
r79 25 32 5.01319 $w=1.75e-07 $l=1.65e-07 $layer=LI1_cond $X=0.425 $Y=2.117
+ $X2=0.26 $Y2=2.117
r80 24 33 6.77202 $w=1.75e-07 $l=2.95e-07 $layer=LI1_cond $X=0.91 $Y=2.117
+ $X2=1.205 $Y2=2.117
r81 24 25 30.7377 $w=1.73e-07 $l=4.85e-07 $layer=LI1_cond $X=0.91 $Y=2.117
+ $X2=0.425 $Y2=2.117
r82 22 26 7.53182 $w=2e-07 $l=2.21425e-07 $layer=LI1_cond $X=0.91 $Y=0.92
+ $X2=1.087 $Y2=1.02
r83 22 23 27.7273 $w=1.98e-07 $l=5e-07 $layer=LI1_cond $X=0.91 $Y=0.92 $X2=0.41
+ $Y2=0.92
r84 18 32 2.6737 $w=3.3e-07 $l=8.8e-08 $layer=LI1_cond $X=0.26 $Y=2.205 $X2=0.26
+ $Y2=2.117
r85 18 20 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=0.26 $Y=2.205
+ $X2=0.26 $Y2=2.915
r86 14 23 7.26812 $w=2e-07 $l=2.01901e-07 $layer=LI1_cond $X=0.252 $Y=0.82
+ $X2=0.41 $Y2=0.92
r87 14 16 12.8049 $w=3.13e-07 $l=3.5e-07 $layer=LI1_cond $X=0.252 $Y=0.82
+ $X2=0.252 $Y2=0.47
r88 10 30 57.7512 $w=6e-07 $l=4.30871e-07 $layer=POLY_cond $X=1.32 $Y=1.93
+ $X2=1.245 $Y2=1.535
r89 10 12 258.492 $w=1.8e-07 $l=6.65e-07 $layer=POLY_cond $X=1.32 $Y=1.93
+ $X2=1.32 $Y2=2.595
r90 7 30 39.2746 $w=6e-07 $l=1.98997e-07 $layer=POLY_cond $X=1.32 $Y=1.37
+ $X2=1.245 $Y2=1.535
r91 7 9 163.344 $w=1.8e-07 $l=6.1e-07 $layer=POLY_cond $X=1.32 $Y=1.37 $X2=1.32
+ $Y2=0.76
r92 2 32 400 $w=1.7e-07 $l=4.17852e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.835 $X2=0.26 $Y2=2.195
r93 2 20 400 $w=1.7e-07 $l=1.14079e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.835 $X2=0.26 $Y2=2.915
r94 1 16 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.26 $X2=0.26 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_LP__DLYBUF4S18KAPWR_1%A_282_52# 1 2 7 9 12 16 18 19 22
+ 23 26
c63 23 0 5.13383e-20 $X=2.52 $Y=1.535
c64 22 0 1.96922e-19 $X=2.52 $Y=1.535
r65 30 31 19.6071 $w=2.52e-07 $l=4.05e-07 $layer=LI1_cond $X=1.67 $Y=1.115
+ $X2=1.67 $Y2=1.52
r66 26 28 9.51376 $w=4.36e-07 $l=3.4e-07 $layer=LI1_cond $X=1.612 $Y=2.265
+ $X2=1.612 $Y2=2.605
r67 23 32 34.0979 $w=3.3e-07 $l=1.95e-07 $layer=POLY_cond $X=2.52 $Y=1.535
+ $X2=2.325 $Y2=1.535
r68 22 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.52
+ $Y=1.535 $X2=2.52 $Y2=1.535
r69 20 31 0.291325 $w=2.7e-07 $l=1.7e-07 $layer=LI1_cond $X=1.84 $Y=1.52
+ $X2=1.67 $Y2=1.52
r70 20 22 29.0245 $w=2.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.84 $Y=1.52
+ $X2=2.52 $Y2=1.52
r71 19 26 9.33164 $w=4.36e-07 $l=2.25433e-07 $layer=LI1_cond $X=1.755 $Y=2.1
+ $X2=1.612 $Y2=2.265
r72 18 31 7.83322 $w=2.52e-07 $l=1.72337e-07 $layer=LI1_cond $X=1.755 $Y=1.655
+ $X2=1.67 $Y2=1.52
r73 18 19 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=1.755 $Y=1.655
+ $X2=1.755 $Y2=2.1
r74 14 30 2.84561 $w=4.05e-07 $l=5.0892e-08 $layer=LI1_cond $X=1.637 $Y=1.078
+ $X2=1.67 $Y2=1.115
r75 14 16 18.2968 $w=4.03e-07 $l=6.43e-07 $layer=LI1_cond $X=1.637 $Y=1.078
+ $X2=1.637 $Y2=0.435
r76 10 32 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.325 $Y=1.7
+ $X2=2.325 $Y2=1.535
r77 10 12 347.895 $w=1.8e-07 $l=8.95e-07 $layer=POLY_cond $X=2.325 $Y=1.7
+ $X2=2.325 $Y2=2.595
r78 7 32 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.325 $Y=1.37
+ $X2=2.325 $Y2=1.535
r79 7 9 163.344 $w=1.8e-07 $l=6.1e-07 $layer=POLY_cond $X=2.325 $Y=1.37
+ $X2=2.325 $Y2=0.76
r80 2 28 300 $w=1.7e-07 $l=5.7576e-07 $layer=licon1_PDIFF $count=2 $X=1.41
+ $Y=2.095 $X2=1.55 $Y2=2.605
r81 2 26 600 $w=1.7e-07 $l=2.29565e-07 $layer=licon1_PDIFF $count=1 $X=1.41
+ $Y=2.095 $X2=1.55 $Y2=2.265
r82 1 30 121.333 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_NDIFF $count=1 $X=1.41
+ $Y=0.26 $X2=1.55 $Y2=1.115
r83 1 16 121.333 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=1 $X=1.41
+ $Y=0.26 $X2=1.55 $Y2=0.435
.ends

.subckt PM_SKY130_FD_SC_LP__DLYBUF4S18KAPWR_1%A_394_52# 1 2 9 13 17 21 22 23 24
+ 25 26 28 32
c77 32 0 1.96922e-19 $X=3.26 $Y=1.46
r78 32 35 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.26 $Y=1.46
+ $X2=3.26 $Y2=1.625
r79 32 34 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.26 $Y=1.46
+ $X2=3.26 $Y2=1.295
r80 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.26
+ $Y=1.46 $X2=3.26 $Y2=1.46
r81 25 31 8.96051 $w=3.33e-07 $l=2.31571e-07 $layer=LI1_cond $X=2.94 $Y=1.625
+ $X2=3.1 $Y2=1.46
r82 25 26 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=2.94 $Y=1.625 $X2=2.94
+ $Y2=1.825
r83 24 28 22.9066 $w=2.51e-07 $l=5.2314e-07 $layer=LI1_cond $X=2.54 $Y=1.91
+ $X2=2.095 $Y2=2.08
r84 23 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.855 $Y=1.91
+ $X2=2.94 $Y2=1.825
r85 23 24 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=2.855 $Y=1.91
+ $X2=2.54 $Y2=1.91
r86 21 31 13.2991 $w=3.33e-07 $l=4.69791e-07 $layer=LI1_cond $X=2.855 $Y=1.097
+ $X2=3.1 $Y2=1.46
r87 21 22 29.1789 $w=2.33e-07 $l=5.95e-07 $layer=LI1_cond $X=2.855 $Y=1.097
+ $X2=2.26 $Y2=1.097
r88 15 22 6.82498 $w=2.35e-07 $l=1.73925e-07 $layer=LI1_cond $X=2.135 $Y=0.98
+ $X2=2.26 $Y2=1.097
r89 15 17 25.1233 $w=2.48e-07 $l=5.45e-07 $layer=LI1_cond $X=2.135 $Y=0.98
+ $X2=2.135 $Y2=0.435
r90 13 35 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=3.17 $Y=2.465
+ $X2=3.17 $Y2=1.625
r91 9 34 423.032 $w=1.5e-07 $l=8.25e-07 $layer=POLY_cond $X=3.17 $Y=0.47
+ $X2=3.17 $Y2=1.295
r92 2 28 300 $w=1.7e-07 $l=2.03101e-07 $layer=licon1_PDIFF $count=2 $X=1.97
+ $Y=2.095 $X2=2.095 $Y2=2.245
r93 1 17 91 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_NDIFF $count=2 $X=1.97
+ $Y=0.26 $X2=2.095 $Y2=0.435
.ends

.subckt PM_SKY130_FD_SC_LP__DLYBUF4S18KAPWR_1%KAPWR 1 2 7 10 17 21
c38 10 0 6.01461e-20 $X=0.76 $Y=2.49
r39 20 21 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.875 $Y=2.81
+ $X2=2.875 $Y2=2.81
r40 17 20 18.8582 $w=3.28e-07 $l=5.4e-07 $layer=LI1_cond $X=2.875 $Y=2.27
+ $X2=2.875 $Y2=2.81
r41 13 14 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.76 $Y=2.81
+ $X2=0.76 $Y2=2.81
r42 10 13 11.1752 $w=3.28e-07 $l=3.2e-07 $layer=LI1_cond $X=0.76 $Y=2.49
+ $X2=0.76 $Y2=2.81
r43 7 21 0.55266 $w=2.55e-07 $l=9.55e-07 $layer=MET1_cond $X=1.92 $Y=2.817
+ $X2=2.875 $Y2=2.817
r44 7 14 0.671294 $w=2.55e-07 $l=1.16e-06 $layer=MET1_cond $X=1.92 $Y=2.817
+ $X2=0.76 $Y2=2.817
r45 2 20 400 $w=1.7e-07 $l=1.06034e-06 $layer=licon1_PDIFF $count=1 $X=2.415
+ $Y=2.095 $X2=2.875 $Y2=2.95
r46 2 17 400 $w=1.7e-07 $l=5.40463e-07 $layer=licon1_PDIFF $count=1 $X=2.415
+ $Y=2.095 $X2=2.875 $Y2=2.27
r47 1 10 300 $w=1.7e-07 $l=7.52712e-07 $layer=licon1_PDIFF $count=2 $X=0.55
+ $Y=1.835 $X2=0.76 $Y2=2.49
.ends

.subckt PM_SKY130_FD_SC_LP__DLYBUF4S18KAPWR_1%X 1 2 7 8 9 10 11 12 13 46 49 53
r26 49 50 7.43121 $w=5.18e-07 $l=1.65e-07 $layer=LI1_cond $X=3.49 $Y=1.98
+ $X2=3.49 $Y2=1.815
r27 32 53 0.92006 $w=5.18e-07 $l=4e-08 $layer=LI1_cond $X=3.49 $Y=2.075 $X2=3.49
+ $Y2=2.035
r28 13 39 3.1052 $w=5.18e-07 $l=1.35e-07 $layer=LI1_cond $X=3.49 $Y=2.775
+ $X2=3.49 $Y2=2.91
r29 12 13 8.51056 $w=5.18e-07 $l=3.7e-07 $layer=LI1_cond $X=3.49 $Y=2.405
+ $X2=3.49 $Y2=2.775
r30 11 53 0.529035 $w=5.18e-07 $l=2.3e-08 $layer=LI1_cond $X=3.49 $Y=2.012
+ $X2=3.49 $Y2=2.035
r31 11 49 0.736048 $w=5.18e-07 $l=3.2e-08 $layer=LI1_cond $X=3.49 $Y=2.012
+ $X2=3.49 $Y2=1.98
r32 11 12 7.08446 $w=5.18e-07 $l=3.08e-07 $layer=LI1_cond $X=3.49 $Y=2.097
+ $X2=3.49 $Y2=2.405
r33 11 32 0.506033 $w=5.18e-07 $l=2.2e-08 $layer=LI1_cond $X=3.49 $Y=2.097
+ $X2=3.49 $Y2=2.075
r34 10 50 7.35602 $w=2.33e-07 $l=1.5e-07 $layer=LI1_cond $X=3.632 $Y=1.665
+ $X2=3.632 $Y2=1.815
r35 9 10 18.1448 $w=2.33e-07 $l=3.7e-07 $layer=LI1_cond $X=3.632 $Y=1.295
+ $X2=3.632 $Y2=1.665
r36 8 9 18.1448 $w=2.33e-07 $l=3.7e-07 $layer=LI1_cond $X=3.632 $Y=0.925
+ $X2=3.632 $Y2=1.295
r37 7 46 1.11752 $w=3.28e-07 $l=3.2e-08 $layer=LI1_cond $X=3.6 $Y=0.475
+ $X2=3.632 $Y2=0.475
r38 7 46 2.74472 $w=2.35e-07 $l=1.65e-07 $layer=LI1_cond $X=3.632 $Y=0.64
+ $X2=3.632 $Y2=0.475
r39 7 42 7.50834 $w=3.28e-07 $l=2.15e-07 $layer=LI1_cond $X=3.6 $Y=0.475
+ $X2=3.385 $Y2=0.475
r40 7 8 10.1233 $w=4.03e-07 $l=2.85e-07 $layer=LI1_cond $X=3.632 $Y=0.64
+ $X2=3.632 $Y2=0.925
r41 2 49 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=3.245
+ $Y=1.835 $X2=3.385 $Y2=1.98
r42 2 39 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=3.245
+ $Y=1.835 $X2=3.385 $Y2=2.91
r43 1 42 182 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_NDIFF $count=1 $X=3.245
+ $Y=0.26 $X2=3.385 $Y2=0.475
.ends

.subckt PM_SKY130_FD_SC_LP__DLYBUF4S18KAPWR_1%VGND 1 2 9 13 16 17 18 20 33 34 37
r37 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r38 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r39 31 34 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r40 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r41 28 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r42 27 30 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.64
+ $Y2=0
r43 27 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r44 25 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.91 $Y=0 $X2=0.745
+ $Y2=0
r45 25 27 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=0.91 $Y=0 $X2=1.2
+ $Y2=0
r46 23 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r47 22 23 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r48 20 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.58 $Y=0 $X2=0.745
+ $Y2=0
r49 20 22 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=0.58 $Y=0 $X2=0.24
+ $Y2=0
r50 18 31 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=2.64
+ $Y2=0
r51 18 28 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=1.2
+ $Y2=0
r52 16 30 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=2.71 $Y=0 $X2=2.64
+ $Y2=0
r53 16 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.71 $Y=0 $X2=2.875
+ $Y2=0
r54 15 33 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=3.04 $Y=0 $X2=3.6
+ $Y2=0
r55 15 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.04 $Y=0 $X2=2.875
+ $Y2=0
r56 11 17 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.875 $Y=0.085
+ $X2=2.875 $Y2=0
r57 11 13 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=2.875 $Y=0.085
+ $X2=2.875 $Y2=0.505
r58 7 37 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.745 $Y=0.085
+ $X2=0.745 $Y2=0
r59 7 9 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=0.745 $Y=0.085
+ $X2=0.745 $Y2=0.47
r60 2 13 182 $w=1.7e-07 $l=5.69473e-07 $layer=licon1_NDIFF $count=1 $X=2.415
+ $Y=0.26 $X2=2.875 $Y2=0.505
r61 1 9 182 $w=1.7e-07 $l=2.91633e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.26 $X2=0.745 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_LP__DLYBUF4S18KAPWR_1%VPWR 1 8 14
r31 5 14 0.00397135 $w=3.84e-06 $l=1.22e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=1.92 $Y2=3.208
r32 5 8 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r33 4 8 219.209 $w=1.68e-07 $l=3.36e-06 $layer=LI1_cond $X=0.24 $Y=3.33 $X2=3.6
+ $Y2=3.33
r34 4 5 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r35 1 14 3.25521e-05 $w=3.84e-06 $l=1e-09 $layer=MET1_cond $X=1.92 $Y=3.207
+ $X2=1.92 $Y2=3.208
.ends

