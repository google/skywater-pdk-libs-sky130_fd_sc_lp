* File: sky130_fd_sc_lp__dfxtp_4.pex.spice
* Created: Wed Sep  2 09:45:21 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__DFXTP_4%CLK 2 5 8 10 11 12 13 14 15 22 24
r29 22 24 45.5639 $w=3.95e-07 $l=1.65e-07 $layer=POLY_cond $X=0.352 $Y=1.045
+ $X2=0.352 $Y2=0.88
r30 22 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.32
+ $Y=1.045 $X2=0.32 $Y2=1.045
r31 14 15 12.5413 $w=3.38e-07 $l=3.7e-07 $layer=LI1_cond $X=0.255 $Y=2.035
+ $X2=0.255 $Y2=2.405
r32 13 14 12.5413 $w=3.38e-07 $l=3.7e-07 $layer=LI1_cond $X=0.255 $Y=1.665
+ $X2=0.255 $Y2=2.035
r33 12 13 12.5413 $w=3.38e-07 $l=3.7e-07 $layer=LI1_cond $X=0.255 $Y=1.295
+ $X2=0.255 $Y2=1.665
r34 12 23 8.47385 $w=3.38e-07 $l=2.5e-07 $layer=LI1_cond $X=0.255 $Y=1.295
+ $X2=0.255 $Y2=1.045
r35 11 23 4.06745 $w=3.38e-07 $l=1.2e-07 $layer=LI1_cond $X=0.255 $Y=0.925
+ $X2=0.255 $Y2=1.045
r36 8 10 569.17 $w=1.5e-07 $l=1.11e-06 $layer=POLY_cond $X=0.475 $Y=2.66
+ $X2=0.475 $Y2=1.55
r37 5 24 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.475 $Y=0.56
+ $X2=0.475 $Y2=0.88
r38 2 10 50.0695 $w=3.95e-07 $l=1.97e-07 $layer=POLY_cond $X=0.352 $Y=1.353
+ $X2=0.352 $Y2=1.55
r39 1 22 4.50555 $w=3.95e-07 $l=3.2e-08 $layer=POLY_cond $X=0.352 $Y=1.077
+ $X2=0.352 $Y2=1.045
r40 1 2 38.8604 $w=3.95e-07 $l=2.76e-07 $layer=POLY_cond $X=0.352 $Y=1.077
+ $X2=0.352 $Y2=1.353
.ends

.subckt PM_SKY130_FD_SC_LP__DFXTP_4%D 3 6 9 11 12 13 14 18 19
r41 18 19 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.99
+ $Y=1.29 $X2=1.99 $Y2=1.29
r42 13 14 8.94038 $w=4.93e-07 $l=3.7e-07 $layer=LI1_cond $X=1.827 $Y=1.295
+ $X2=1.827 $Y2=1.665
r43 13 19 0.120816 $w=4.93e-07 $l=5e-09 $layer=LI1_cond $X=1.827 $Y=1.295
+ $X2=1.827 $Y2=1.29
r44 11 18 42.841 $w=3.3e-07 $l=2.45e-07 $layer=POLY_cond $X=1.99 $Y=1.535
+ $X2=1.99 $Y2=1.29
r45 11 12 62.8233 $w=3.3e-07 $l=2.6e-07 $layer=POLY_cond $X=2.012 $Y=1.535
+ $X2=2.012 $Y2=1.795
r46 9 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.99 $Y=1.125
+ $X2=1.99 $Y2=1.29
r47 6 12 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.125 $Y=2.275
+ $X2=2.125 $Y2=1.795
r48 3 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.08 $Y=0.805 $X2=2.08
+ $Y2=1.125
.ends

.subckt PM_SKY130_FD_SC_LP__DFXTP_4%A_217_413# 1 2 9 11 15 19 22 23 24 27 32 33
+ 36 37 38 41 44 46 49 51 53 56 57 62 63 69
c168 69 0 6.93e-20 $X=2.855 $Y=1.71
c169 49 0 1.30115e-19 $X=4.845 $Y=2.285
c170 46 0 1.17631e-19 $X=4.76 $Y=2.37
r171 63 70 10.0417 $w=2.64e-07 $l=5.5e-08 $layer=POLY_cond $X=4.825 $Y=1.39
+ $X2=4.77 $Y2=1.39
r172 62 65 9.43135 $w=1.98e-07 $l=1.65e-07 $layer=LI1_cond $X=4.83 $Y=1.39
+ $X2=4.83 $Y2=1.555
r173 62 63 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.825
+ $Y=1.39 $X2=4.825 $Y2=1.39
r174 57 59 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=3.41 $Y=2.37
+ $X2=3.41 $Y2=2.62
r175 53 55 7.12573 $w=2.78e-07 $l=1.55e-07 $layer=LI1_cond $X=1.34 $Y=0.805
+ $X2=1.34 $Y2=0.96
r176 49 65 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=4.845 $Y=2.285
+ $X2=4.845 $Y2=1.555
r177 47 57 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.495 $Y=2.37
+ $X2=3.41 $Y2=2.37
r178 46 49 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.76 $Y=2.37
+ $X2=4.845 $Y2=2.285
r179 46 47 82.5294 $w=1.68e-07 $l=1.265e-06 $layer=LI1_cond $X=4.76 $Y=2.37
+ $X2=3.495 $Y2=2.37
r180 45 56 5.41628 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=2.775 $Y=2.62
+ $X2=2.685 $Y2=2.62
r181 44 59 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.325 $Y=2.62
+ $X2=3.41 $Y2=2.62
r182 44 45 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=3.325 $Y=2.62
+ $X2=2.775 $Y2=2.62
r183 42 69 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.69 $Y=1.71
+ $X2=2.855 $Y2=1.71
r184 42 66 23.6063 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=2.69 $Y=1.71
+ $X2=2.555 $Y2=1.71
r185 41 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.69
+ $Y=1.71 $X2=2.69 $Y2=1.71
r186 39 56 1.13756 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.685 $Y=2.535
+ $X2=2.685 $Y2=2.62
r187 39 41 50.8333 $w=1.78e-07 $l=8.25e-07 $layer=LI1_cond $X=2.685 $Y=2.535
+ $X2=2.685 $Y2=1.71
r188 37 56 5.41628 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=2.595 $Y=2.62
+ $X2=2.685 $Y2=2.62
r189 37 38 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=2.595 $Y=2.62
+ $X2=2.075 $Y2=2.62
r190 36 38 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.99 $Y=2.535
+ $X2=2.075 $Y2=2.62
r191 35 36 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=1.99 $Y=2.215
+ $X2=1.99 $Y2=2.535
r192 34 51 2.60907 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=1.41 $Y=2.13
+ $X2=1.227 $Y2=2.13
r193 33 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.905 $Y=2.13
+ $X2=1.99 $Y2=2.215
r194 33 34 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=1.905 $Y=2.13
+ $X2=1.41 $Y2=2.13
r195 32 51 3.84343 $w=2.4e-07 $l=1.17707e-07 $layer=LI1_cond $X=1.305 $Y=2.045
+ $X2=1.227 $Y2=2.13
r196 32 55 57.303 $w=2.08e-07 $l=1.085e-06 $layer=LI1_cond $X=1.305 $Y=2.045
+ $X2=1.305 $Y2=0.96
r197 25 27 225.617 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=5.505 $Y=1.975
+ $X2=5.505 $Y2=2.415
r198 23 25 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.43 $Y=1.9
+ $X2=5.505 $Y2=1.975
r199 23 24 128.191 $w=1.5e-07 $l=2.5e-07 $layer=POLY_cond $X=5.43 $Y=1.9
+ $X2=5.18 $Y2=1.9
r200 22 24 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.105 $Y=1.825
+ $X2=5.18 $Y2=1.9
r201 21 63 51.1212 $w=2.64e-07 $l=3.52987e-07 $layer=POLY_cond $X=5.105 $Y=1.555
+ $X2=4.825 $Y2=1.39
r202 21 22 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=5.105 $Y=1.555
+ $X2=5.105 $Y2=1.825
r203 17 70 15.9823 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.77 $Y=1.225
+ $X2=4.77 $Y2=1.39
r204 17 19 215.362 $w=1.5e-07 $l=4.2e-07 $layer=POLY_cond $X=4.77 $Y=1.225
+ $X2=4.77 $Y2=0.805
r205 13 15 379.447 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=3.135 $Y=1.545
+ $X2=3.135 $Y2=0.805
r206 11 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.06 $Y=1.62
+ $X2=3.135 $Y2=1.545
r207 11 69 105.117 $w=1.5e-07 $l=2.05e-07 $layer=POLY_cond $X=3.06 $Y=1.62
+ $X2=2.855 $Y2=1.62
r208 7 66 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.555 $Y=1.875
+ $X2=2.555 $Y2=1.71
r209 7 9 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=2.555 $Y=1.875
+ $X2=2.555 $Y2=2.275
r210 2 51 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=1.085
+ $Y=2.065 $X2=1.21 $Y2=2.21
r211 1 53 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=1.2
+ $Y=0.595 $X2=1.325 $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_LP__DFXTP_4%A_684_93# 1 2 9 13 17 18 20 21 23 25
c69 18 0 1.17631e-19 $X=3.585 $Y=1.53
r70 25 27 8.61591 $w=2.68e-07 $l=1.65e-07 $layer=LI1_cond $X=4.425 $Y=0.77
+ $X2=4.425 $Y2=0.935
r71 23 29 4.29664 $w=1.7e-07 $l=1.34907e-07 $layer=LI1_cond $X=4.475 $Y=1.855
+ $X2=4.485 $Y2=1.985
r72 23 27 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=4.475 $Y=1.855
+ $X2=4.475 $Y2=0.935
r73 20 29 2.91558 $w=2.6e-07 $l=9.5e-08 $layer=LI1_cond $X=4.39 $Y=1.985
+ $X2=4.485 $Y2=1.985
r74 20 21 28.3678 $w=2.58e-07 $l=6.4e-07 $layer=LI1_cond $X=4.39 $Y=1.985
+ $X2=3.75 $Y2=1.985
r75 18 32 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.585 $Y=1.53
+ $X2=3.585 $Y2=1.695
r76 18 31 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.585 $Y=1.53
+ $X2=3.585 $Y2=1.365
r77 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.585
+ $Y=1.53 $X2=3.585 $Y2=1.53
r78 15 21 6.94204 $w=2.6e-07 $l=2.20624e-07 $layer=LI1_cond $X=3.585 $Y=1.855
+ $X2=3.75 $Y2=1.985
r79 15 17 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=3.585 $Y=1.855
+ $X2=3.585 $Y2=1.53
r80 13 32 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=3.615 $Y=2.275
+ $X2=3.615 $Y2=1.695
r81 9 31 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=3.495 $Y=0.805
+ $X2=3.495 $Y2=1.365
r82 2 29 600 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=4.275
+ $Y=1.895 $X2=4.415 $Y2=2.02
r83 1 25 182 $w=1.7e-07 $l=2.40312e-07 $layer=licon1_NDIFF $count=1 $X=4.3
+ $Y=0.595 $X2=4.455 $Y2=0.77
.ends

.subckt PM_SKY130_FD_SC_LP__DFXTP_4%A_526_413# 1 2 9 13 16 20 22 26 27 29 33
c72 9 0 1.30115e-19 $X=4.2 $Y=2.315
r73 29 31 7.58908 $w=4.23e-07 $l=1.6e-07 $layer=LI1_cond $X=2.932 $Y=1.19
+ $X2=2.932 $Y2=1.35
r74 29 30 2.91128 $w=4.23e-07 $l=8.5e-08 $layer=LI1_cond $X=2.932 $Y=1.19
+ $X2=2.932 $Y2=1.105
r75 27 34 46.3065 $w=3.4e-07 $l=1.65e-07 $layer=POLY_cond $X=4.13 $Y=1.51
+ $X2=4.13 $Y2=1.675
r76 27 33 46.3065 $w=3.4e-07 $l=1.65e-07 $layer=POLY_cond $X=4.13 $Y=1.51
+ $X2=4.13 $Y2=1.345
r77 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.125
+ $Y=1.51 $X2=4.125 $Y2=1.51
r78 24 26 10.4163 $w=2.58e-07 $l=2.35e-07 $layer=LI1_cond $X=4.09 $Y=1.275
+ $X2=4.09 $Y2=1.51
r79 23 29 6.14847 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=3.145 $Y=1.19
+ $X2=2.932 $Y2=1.19
r80 22 24 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=3.96 $Y=1.19
+ $X2=4.09 $Y2=1.275
r81 22 23 53.1711 $w=1.68e-07 $l=8.15e-07 $layer=LI1_cond $X=3.96 $Y=1.19
+ $X2=3.145 $Y2=1.19
r82 20 31 46.5818 $w=1.98e-07 $l=8.4e-07 $layer=LI1_cond $X=3.045 $Y=2.19
+ $X2=3.045 $Y2=1.35
r83 16 30 10.4768 $w=3.28e-07 $l=3e-07 $layer=LI1_cond $X=2.885 $Y=0.805
+ $X2=2.885 $Y2=1.105
r84 13 33 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=4.225 $Y=0.915
+ $X2=4.225 $Y2=1.345
r85 9 34 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=4.2 $Y=2.315 $X2=4.2
+ $Y2=1.675
r86 2 20 600 $w=1.7e-07 $l=4.58258e-07 $layer=licon1_PDIFF $count=1 $X=2.63
+ $Y=2.065 $X2=3.03 $Y2=2.19
r87 1 16 182 $w=1.7e-07 $l=2.93428e-07 $layer=licon1_NDIFF $count=1 $X=2.685
+ $Y=0.595 $X2=2.885 $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_LP__DFXTP_4%A_110_70# 1 2 7 8 12 16 17 18 19 20 23 25 29
+ 31 35 39 43 45 46 49 52 55 58 59 61
c131 61 0 4.11139e-20 $X=0.812 $Y=1.865
r132 58 60 6.22179 $w=4.33e-07 $l=1.65e-07 $layer=LI1_cond $X=0.812 $Y=1.36
+ $X2=0.812 $Y2=1.195
r133 58 59 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.945
+ $Y=1.36 $X2=0.945 $Y2=1.36
r134 55 61 27.4813 $w=2.58e-07 $l=6.2e-07 $layer=LI1_cond $X=0.725 $Y=2.485
+ $X2=0.725 $Y2=1.865
r135 52 61 7.59943 $w=4.33e-07 $l=2.17e-07 $layer=LI1_cond $X=0.812 $Y=1.648
+ $X2=0.812 $Y2=1.865
r136 51 58 1.37763 $w=4.33e-07 $l=5.2e-08 $layer=LI1_cond $X=0.812 $Y=1.412
+ $X2=0.812 $Y2=1.36
r137 51 52 6.25233 $w=4.33e-07 $l=2.36e-07 $layer=LI1_cond $X=0.812 $Y=1.412
+ $X2=0.812 $Y2=1.648
r138 49 60 28.1462 $w=2.58e-07 $l=6.35e-07 $layer=LI1_cond $X=0.725 $Y=0.56
+ $X2=0.725 $Y2=1.195
r139 42 43 58.9681 $w=1.5e-07 $l=1.15e-07 $layer=POLY_cond $X=1.425 $Y=1.27
+ $X2=1.54 $Y2=1.27
r140 41 59 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=0.945 $Y=1.345
+ $X2=0.945 $Y2=1.36
r141 37 39 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=5.275 $Y=0.255
+ $X2=5.275 $Y2=0.805
r142 33 35 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=4.63 $Y=3.075
+ $X2=4.63 $Y2=2.315
r143 32 46 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.33 $Y=3.15
+ $X2=3.255 $Y2=3.15
r144 31 33 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.555 $Y=3.15
+ $X2=4.63 $Y2=3.075
r145 31 32 628.138 $w=1.5e-07 $l=1.225e-06 $layer=POLY_cond $X=4.555 $Y=3.15
+ $X2=3.33 $Y2=3.15
r146 27 46 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.255 $Y=3.075
+ $X2=3.255 $Y2=3.15
r147 27 29 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=3.255 $Y=3.075
+ $X2=3.255 $Y2=2.275
r148 26 45 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.685 $Y=0.18
+ $X2=2.61 $Y2=0.18
r149 25 37 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.2 $Y=0.18
+ $X2=5.275 $Y2=0.255
r150 25 26 1289.61 $w=1.5e-07 $l=2.515e-06 $layer=POLY_cond $X=5.2 $Y=0.18
+ $X2=2.685 $Y2=0.18
r151 21 45 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.61 $Y=0.255
+ $X2=2.61 $Y2=0.18
r152 21 23 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=2.61 $Y=0.255
+ $X2=2.61 $Y2=0.805
r153 19 45 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.535 $Y=0.18
+ $X2=2.61 $Y2=0.18
r154 19 20 471.745 $w=1.5e-07 $l=9.2e-07 $layer=POLY_cond $X=2.535 $Y=0.18
+ $X2=1.615 $Y2=0.18
r155 17 46 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.18 $Y=3.15
+ $X2=3.255 $Y2=3.15
r156 17 18 861.447 $w=1.5e-07 $l=1.68e-06 $layer=POLY_cond $X=3.18 $Y=3.15
+ $X2=1.5 $Y2=3.15
r157 14 43 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.54 $Y=1.195
+ $X2=1.54 $Y2=1.27
r158 14 16 199.979 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=1.54 $Y=1.195
+ $X2=1.54 $Y2=0.805
r159 13 20 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.54 $Y=0.255
+ $X2=1.615 $Y2=0.18
r160 13 16 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=1.54 $Y=0.255
+ $X2=1.54 $Y2=0.805
r161 10 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.425 $Y=3.075
+ $X2=1.5 $Y2=3.15
r162 10 12 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.425 $Y=3.075
+ $X2=1.425 $Y2=2.385
r163 9 42 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.425 $Y=1.345
+ $X2=1.425 $Y2=1.27
r164 9 12 533.277 $w=1.5e-07 $l=1.04e-06 $layer=POLY_cond $X=1.425 $Y=1.345
+ $X2=1.425 $Y2=2.385
r165 8 41 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=1.11 $Y=1.27
+ $X2=0.945 $Y2=1.345
r166 7 42 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.35 $Y=1.27
+ $X2=1.425 $Y2=1.27
r167 7 8 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=1.35 $Y=1.27 $X2=1.11
+ $Y2=1.27
r168 2 55 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=0.55
+ $Y=2.34 $X2=0.69 $Y2=2.485
r169 1 49 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.35 $X2=0.69 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_LP__DFXTP_4%A_1112_93# 1 2 9 13 17 21 25 29 33 37 41 45
+ 49 52 53 54 56 61 67 71 76 82 88
c151 76 0 1.06395e-19 $X=7.265 $Y=1.48
r152 85 86 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=7.77 $Y=1.48
+ $X2=8.2 $Y2=1.48
r153 84 85 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=7.34 $Y=1.48
+ $X2=7.77 $Y2=1.48
r154 76 84 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=7.265 $Y=1.48
+ $X2=7.34 $Y2=1.48
r155 74 75 18.7692 $w=1.95e-07 $l=3e-07 $layer=LI1_cond $X=6.63 $Y=1.48 $X2=6.63
+ $Y2=1.78
r156 71 73 16.8753 $w=4.53e-07 $l=4.55e-07 $layer=LI1_cond $X=6.522 $Y=0.39
+ $X2=6.522 $Y2=0.845
r157 68 88 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=8.45 $Y=1.48
+ $X2=8.63 $Y2=1.48
r158 68 86 43.7153 $w=3.3e-07 $l=2.5e-07 $layer=POLY_cond $X=8.45 $Y=1.48
+ $X2=8.2 $Y2=1.48
r159 67 68 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=8.45
+ $Y=1.48 $X2=8.45 $Y2=1.48
r160 65 76 30.6007 $w=3.3e-07 $l=1.75e-07 $layer=POLY_cond $X=7.09 $Y=1.48
+ $X2=7.265 $Y2=1.48
r161 64 67 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=7.09 $Y=1.48
+ $X2=8.45 $Y2=1.48
r162 64 65 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=7.09
+ $Y=1.48 $X2=7.09 $Y2=1.48
r163 62 74 1.54022 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=6.75 $Y=1.48
+ $X2=6.63 $Y2=1.48
r164 62 64 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=6.75 $Y=1.48
+ $X2=7.09 $Y2=1.48
r165 61 74 5.55076 $w=1.95e-07 $l=1.00995e-07 $layer=LI1_cond $X=6.665 $Y=1.395
+ $X2=6.63 $Y2=1.48
r166 61 73 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=6.665 $Y=1.395
+ $X2=6.665 $Y2=0.845
r167 56 58 46.5779 $w=2.38e-07 $l=9.7e-07 $layer=LI1_cond $X=6.63 $Y=1.87
+ $X2=6.63 $Y2=2.84
r168 54 75 4.78561 $w=2.4e-07 $l=8.5e-08 $layer=LI1_cond $X=6.63 $Y=1.865
+ $X2=6.63 $Y2=1.78
r169 54 56 0.240092 $w=2.38e-07 $l=5e-09 $layer=LI1_cond $X=6.63 $Y=1.865
+ $X2=6.63 $Y2=1.87
r170 52 75 1.54022 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=6.51 $Y=1.78
+ $X2=6.63 $Y2=1.78
r171 52 53 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=6.51 $Y=1.78
+ $X2=5.89 $Y2=1.78
r172 50 82 24.4806 $w=3.3e-07 $l=1.4e-07 $layer=POLY_cond $X=5.725 $Y=1.45
+ $X2=5.865 $Y2=1.45
r173 50 79 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=5.725 $Y=1.45
+ $X2=5.635 $Y2=1.45
r174 49 50 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.725
+ $Y=1.45 $X2=5.725 $Y2=1.45
r175 47 53 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.725 $Y=1.695
+ $X2=5.89 $Y2=1.78
r176 47 49 8.55602 $w=3.28e-07 $l=2.45e-07 $layer=LI1_cond $X=5.725 $Y=1.695
+ $X2=5.725 $Y2=1.45
r177 43 88 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.63 $Y=1.645
+ $X2=8.63 $Y2=1.48
r178 43 45 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=8.63 $Y=1.645
+ $X2=8.63 $Y2=2.465
r179 39 88 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.63 $Y=1.315
+ $X2=8.63 $Y2=1.48
r180 39 41 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=8.63 $Y=1.315
+ $X2=8.63 $Y2=0.655
r181 35 86 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.2 $Y=1.645
+ $X2=8.2 $Y2=1.48
r182 35 37 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=8.2 $Y=1.645
+ $X2=8.2 $Y2=2.465
r183 31 86 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.2 $Y=1.315
+ $X2=8.2 $Y2=1.48
r184 31 33 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=8.2 $Y=1.315
+ $X2=8.2 $Y2=0.655
r185 27 85 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.77 $Y=1.645
+ $X2=7.77 $Y2=1.48
r186 27 29 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=7.77 $Y=1.645
+ $X2=7.77 $Y2=2.465
r187 23 85 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.77 $Y=1.315
+ $X2=7.77 $Y2=1.48
r188 23 25 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=7.77 $Y=1.315
+ $X2=7.77 $Y2=0.655
r189 19 84 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.34 $Y=1.645
+ $X2=7.34 $Y2=1.48
r190 19 21 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=7.34 $Y=1.645
+ $X2=7.34 $Y2=2.465
r191 15 84 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.34 $Y=1.315
+ $X2=7.34 $Y2=1.48
r192 15 17 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=7.34 $Y=1.315
+ $X2=7.34 $Y2=0.655
r193 11 82 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.865 $Y=1.615
+ $X2=5.865 $Y2=1.45
r194 11 13 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=5.865 $Y=1.615
+ $X2=5.865 $Y2=2.415
r195 7 79 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.635 $Y=1.285
+ $X2=5.635 $Y2=1.45
r196 7 9 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=5.635 $Y=1.285
+ $X2=5.635 $Y2=0.805
r197 2 58 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=6.465
+ $Y=1.725 $X2=6.605 $Y2=2.84
r198 2 56 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=6.465
+ $Y=1.725 $X2=6.605 $Y2=1.87
r199 1 71 91 $w=1.7e-07 $l=2.24499e-07 $layer=licon1_NDIFF $count=2 $X=6.3
+ $Y=0.235 $X2=6.46 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_LP__DFXTP_4%A_941_379# 1 2 9 12 14 16 20 24 25 31
c79 24 0 1.06395e-19 $X=6.315 $Y=1.35
r80 28 29 10.7433 $w=3.35e-07 $l=2.95e-07 $layer=LI1_cond $X=5.127 $Y=0.805
+ $X2=5.127 $Y2=1.1
r81 25 32 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.315 $Y=1.35
+ $X2=6.315 $Y2=1.515
r82 25 31 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.315 $Y=1.35
+ $X2=6.315 $Y2=1.185
r83 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.315
+ $Y=1.35 $X2=6.315 $Y2=1.35
r84 22 24 7.31358 $w=2.58e-07 $l=1.65e-07 $layer=LI1_cond $X=6.28 $Y=1.185
+ $X2=6.28 $Y2=1.35
r85 21 29 4.71304 $w=1.7e-07 $l=2.33e-07 $layer=LI1_cond $X=5.36 $Y=1.1
+ $X2=5.127 $Y2=1.1
r86 20 22 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=6.15 $Y=1.1
+ $X2=6.28 $Y2=1.185
r87 20 21 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=6.15 $Y=1.1 $X2=5.36
+ $Y2=1.1
r88 16 18 15.6732 $w=2.48e-07 $l=3.4e-07 $layer=LI1_cond $X=5.235 $Y=2.195
+ $X2=5.235 $Y2=2.535
r89 14 29 3.90748 $w=3.35e-07 $l=1.44375e-07 $layer=LI1_cond $X=5.235 $Y=1.185
+ $X2=5.127 $Y2=1.1
r90 14 16 46.5587 $w=2.48e-07 $l=1.01e-06 $layer=LI1_cond $X=5.235 $Y=1.185
+ $X2=5.235 $Y2=2.195
r91 12 32 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=6.39 $Y=2.355
+ $X2=6.39 $Y2=1.515
r92 9 31 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=6.225 $Y=0.655
+ $X2=6.225 $Y2=1.185
r93 2 18 600 $w=1.7e-07 $l=8.50412e-07 $layer=licon1_PDIFF $count=1 $X=4.705
+ $Y=1.895 $X2=5.195 $Y2=2.535
r94 2 16 600 $w=1.7e-07 $l=6.22174e-07 $layer=licon1_PDIFF $count=1 $X=4.705
+ $Y=1.895 $X2=5.195 $Y2=2.195
r95 1 28 182 $w=1.7e-07 $l=3.02283e-07 $layer=licon1_NDIFF $count=1 $X=4.845
+ $Y=0.595 $X2=5.06 $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_LP__DFXTP_4%VPWR 1 2 3 4 5 6 7 22 24 28 32 36 40 44 50
+ 54 56 58 59 60 62 67 76 81 90 93 96 99 103
r118 102 103 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r119 99 100 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r120 96 97 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r121 93 94 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r122 90 91 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r123 87 88 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r124 85 103 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=8.88 $Y2=3.33
r125 85 100 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=7.92 $Y2=3.33
r126 84 85 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=3.33 $X2=8.4
+ $Y2=3.33
r127 82 99 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.15 $Y=3.33
+ $X2=7.985 $Y2=3.33
r128 82 84 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=8.15 $Y=3.33
+ $X2=8.4 $Y2=3.33
r129 81 102 4.746 $w=1.7e-07 $l=2.2e-07 $layer=LI1_cond $X=8.68 $Y=3.33 $X2=8.9
+ $Y2=3.33
r130 81 84 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=8.68 $Y=3.33
+ $X2=8.4 $Y2=3.33
r131 80 100 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=7.92 $Y2=3.33
r132 80 97 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=6.96 $Y2=3.33
r133 79 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r134 77 96 7.94884 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=7.255 $Y=3.33
+ $X2=7.107 $Y2=3.33
r135 77 79 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=7.255 $Y=3.33
+ $X2=7.44 $Y2=3.33
r136 76 99 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.82 $Y=3.33
+ $X2=7.985 $Y2=3.33
r137 76 79 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=7.82 $Y=3.33
+ $X2=7.44 $Y2=3.33
r138 75 97 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=6.96
+ $Y2=3.33
r139 74 75 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r140 72 93 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.09 $Y=3.33
+ $X2=3.925 $Y2=3.33
r141 72 74 124.61 $w=1.68e-07 $l=1.91e-06 $layer=LI1_cond $X=4.09 $Y=3.33 $X2=6
+ $Y2=3.33
r142 71 94 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r143 71 91 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=1.68 $Y2=3.33
r144 70 71 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r145 68 90 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.725 $Y=3.33
+ $X2=1.63 $Y2=3.33
r146 68 70 122.326 $w=1.68e-07 $l=1.875e-06 $layer=LI1_cond $X=1.725 $Y=3.33
+ $X2=3.6 $Y2=3.33
r147 67 93 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.76 $Y=3.33
+ $X2=3.925 $Y2=3.33
r148 67 70 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=3.76 $Y=3.33
+ $X2=3.6 $Y2=3.33
r149 66 91 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r150 66 88 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.24 $Y2=3.33
r151 65 66 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r152 63 87 4.78091 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=3.33
+ $X2=0.212 $Y2=3.33
r153 63 65 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=0.425 $Y=3.33
+ $X2=1.2 $Y2=3.33
r154 62 90 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.535 $Y=3.33
+ $X2=1.63 $Y2=3.33
r155 62 65 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.535 $Y=3.33
+ $X2=1.2 $Y2=3.33
r156 60 75 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=6 $Y2=3.33
r157 60 94 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=4.08 $Y2=3.33
r158 58 74 0.652406 $w=1.68e-07 $l=1e-08 $layer=LI1_cond $X=6.01 $Y=3.33 $X2=6
+ $Y2=3.33
r159 58 59 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.01 $Y=3.33
+ $X2=6.175 $Y2=3.33
r160 54 102 3.02018 $w=3.3e-07 $l=1.09087e-07 $layer=LI1_cond $X=8.845 $Y=3.245
+ $X2=8.9 $Y2=3.33
r161 54 56 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=8.845 $Y=3.245
+ $X2=8.845 $Y2=2.795
r162 50 53 28.2872 $w=3.28e-07 $l=8.1e-07 $layer=LI1_cond $X=7.985 $Y=2.16
+ $X2=7.985 $Y2=2.97
r163 48 99 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.985 $Y=3.245
+ $X2=7.985 $Y2=3.33
r164 48 53 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=7.985 $Y=3.245
+ $X2=7.985 $Y2=2.97
r165 44 47 37.8939 $w=2.93e-07 $l=9.7e-07 $layer=LI1_cond $X=7.107 $Y=1.98
+ $X2=7.107 $Y2=2.95
r166 42 96 0.543863 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=7.107 $Y=3.245
+ $X2=7.107 $Y2=3.33
r167 42 47 11.5244 $w=2.93e-07 $l=2.95e-07 $layer=LI1_cond $X=7.107 $Y=3.245
+ $X2=7.107 $Y2=2.95
r168 41 59 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.34 $Y=3.33
+ $X2=6.175 $Y2=3.33
r169 40 96 7.94884 $w=1.7e-07 $l=1.47e-07 $layer=LI1_cond $X=6.96 $Y=3.33
+ $X2=7.107 $Y2=3.33
r170 40 41 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=6.96 $Y=3.33
+ $X2=6.34 $Y2=3.33
r171 36 39 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=6.175 $Y=2.16
+ $X2=6.175 $Y2=2.84
r172 34 59 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.175 $Y=3.245
+ $X2=6.175 $Y2=3.33
r173 34 39 14.1436 $w=3.28e-07 $l=4.05e-07 $layer=LI1_cond $X=6.175 $Y=3.245
+ $X2=6.175 $Y2=2.84
r174 30 93 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.925 $Y=3.245
+ $X2=3.925 $Y2=3.33
r175 30 32 18.3343 $w=3.28e-07 $l=5.25e-07 $layer=LI1_cond $X=3.925 $Y=3.245
+ $X2=3.925 $Y2=2.72
r176 26 90 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.63 $Y=3.245
+ $X2=1.63 $Y2=3.33
r177 26 28 39.9856 $w=1.88e-07 $l=6.85e-07 $layer=LI1_cond $X=1.63 $Y=3.245
+ $X2=1.63 $Y2=2.56
r178 22 87 2.98526 $w=3.3e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.26 $Y=3.245
+ $X2=0.212 $Y2=3.33
r179 22 24 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=0.26 $Y=3.245
+ $X2=0.26 $Y2=2.83
r180 7 56 600 $w=1.7e-07 $l=1.02762e-06 $layer=licon1_PDIFF $count=1 $X=8.705
+ $Y=1.835 $X2=8.845 $Y2=2.795
r181 6 53 400 $w=1.7e-07 $l=1.20297e-06 $layer=licon1_PDIFF $count=1 $X=7.845
+ $Y=1.835 $X2=7.985 $Y2=2.97
r182 6 50 400 $w=1.7e-07 $l=3.88748e-07 $layer=licon1_PDIFF $count=1 $X=7.845
+ $Y=1.835 $X2=7.985 $Y2=2.16
r183 5 47 400 $w=1.7e-07 $l=1.17584e-06 $layer=licon1_PDIFF $count=1 $X=7
+ $Y=1.835 $X2=7.125 $Y2=2.95
r184 5 44 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=7
+ $Y=1.835 $X2=7.125 $Y2=1.98
r185 4 39 600 $w=1.7e-07 $l=7.4327e-07 $layer=licon1_PDIFF $count=1 $X=5.94
+ $Y=2.205 $X2=6.175 $Y2=2.84
r186 4 36 300 $w=1.7e-07 $l=2.56515e-07 $layer=licon1_PDIFF $count=2 $X=5.94
+ $Y=2.205 $X2=6.175 $Y2=2.16
r187 3 32 600 $w=1.7e-07 $l=7.63512e-07 $layer=licon1_PDIFF $count=1 $X=3.69
+ $Y=2.065 $X2=3.925 $Y2=2.72
r188 2 28 600 $w=1.7e-07 $l=5.60647e-07 $layer=licon1_PDIFF $count=1 $X=1.5
+ $Y=2.065 $X2=1.64 $Y2=2.56
r189 1 24 600 $w=1.7e-07 $l=5.48954e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.34 $X2=0.26 $Y2=2.83
.ends

.subckt PM_SKY130_FD_SC_LP__DFXTP_4%A_431_119# 1 2 9 11 14 17
c23 14 0 6.93e-20 $X=2.385 $Y=0.79
r24 16 17 63.6096 $w=1.68e-07 $l=9.75e-07 $layer=LI1_cond $X=2.33 $Y=0.955
+ $X2=2.33 $Y2=1.93
r25 14 16 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=2.385 $Y=0.79
+ $X2=2.385 $Y2=0.955
r26 9 17 5.59224 $w=1.78e-07 $l=9e-08 $layer=LI1_cond $X=2.335 $Y=2.02 $X2=2.335
+ $Y2=1.93
r27 9 11 10.4747 $w=1.78e-07 $l=1.7e-07 $layer=LI1_cond $X=2.335 $Y=2.02
+ $X2=2.335 $Y2=2.19
r28 2 11 600 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=2.2
+ $Y=2.065 $X2=2.34 $Y2=2.19
r29 1 14 182 $w=1.7e-07 $l=3.1265e-07 $layer=licon1_NDIFF $count=1 $X=2.155
+ $Y=0.595 $X2=2.385 $Y2=0.79
.ends

.subckt PM_SKY130_FD_SC_LP__DFXTP_4%Q 1 2 3 4 15 19 24 25 26 29 33 38 39 41 42
+ 43 55 59 69 73
r60 53 59 3.36129 $w=2.38e-07 $l=7e-08 $layer=LI1_cond $X=8.915 $Y=1.735
+ $X2=8.915 $Y2=1.665
r61 52 73 3.50224 $w=2.4e-07 $l=1.93e-07 $layer=LI1_cond $X=8.915 $Y=1.225
+ $X2=8.915 $Y2=1.032
r62 52 55 3.36129 $w=2.38e-07 $l=7e-08 $layer=LI1_cond $X=8.915 $Y=1.225
+ $X2=8.915 $Y2=1.295
r63 42 43 17.7668 $w=2.38e-07 $l=3.7e-07 $layer=LI1_cond $X=8.915 $Y=2.035
+ $X2=8.915 $Y2=2.405
r64 42 60 4.32166 $w=2.38e-07 $l=9e-08 $layer=LI1_cond $X=8.915 $Y=2.035
+ $X2=8.915 $Y2=1.945
r65 41 53 4.61626 $w=2.4e-07 $l=1.05e-07 $layer=LI1_cond $X=8.915 $Y=1.84
+ $X2=8.915 $Y2=1.735
r66 41 60 4.61626 $w=2.4e-07 $l=1.05e-07 $layer=LI1_cond $X=8.915 $Y=1.84
+ $X2=8.915 $Y2=1.945
r67 41 59 0.384148 $w=2.38e-07 $l=8e-09 $layer=LI1_cond $X=8.915 $Y=1.657
+ $X2=8.915 $Y2=1.665
r68 39 73 1.04768 $w=3.83e-07 $l=3.5e-08 $layer=LI1_cond $X=8.88 $Y=1.032
+ $X2=8.915 $Y2=1.032
r69 39 41 17.0466 $w=2.38e-07 $l=3.55e-07 $layer=LI1_cond $X=8.915 $Y=1.302
+ $X2=8.915 $Y2=1.657
r70 39 55 0.336129 $w=2.38e-07 $l=7e-09 $layer=LI1_cond $X=8.915 $Y=1.302
+ $X2=8.915 $Y2=1.295
r71 37 41 14.6652 $w=2.23e-07 $l=2.85e-07 $layer=LI1_cond $X=8.51 $Y=1.84
+ $X2=8.795 $Y2=1.84
r72 37 38 5.16603 $w=1.9e-07 $l=9.5e-08 $layer=LI1_cond $X=8.51 $Y=1.84
+ $X2=8.415 $Y2=1.84
r73 33 35 55.4545 $w=1.88e-07 $l=9.5e-07 $layer=LI1_cond $X=8.415 $Y=1.96
+ $X2=8.415 $Y2=2.91
r74 31 38 1.34256 $w=1.9e-07 $l=1.05e-07 $layer=LI1_cond $X=8.415 $Y=1.945
+ $X2=8.415 $Y2=1.84
r75 31 33 0.875598 $w=1.88e-07 $l=1.5e-08 $layer=LI1_cond $X=8.415 $Y=1.945
+ $X2=8.415 $Y2=1.96
r76 27 39 13.9191 $w=3.83e-07 $l=4.65e-07 $layer=LI1_cond $X=8.415 $Y=1.032
+ $X2=8.88 $Y2=1.032
r77 27 69 6.49359 $w=3.83e-07 $l=9.5e-08 $layer=LI1_cond $X=8.415 $Y=1.032
+ $X2=8.32 $Y2=1.032
r78 27 29 24.5167 $w=1.88e-07 $l=4.2e-07 $layer=LI1_cond $X=8.415 $Y=0.84
+ $X2=8.415 $Y2=0.42
r79 25 38 5.16603 $w=1.9e-07 $l=1.04523e-07 $layer=LI1_cond $X=8.32 $Y=1.82
+ $X2=8.415 $Y2=1.84
r80 25 26 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=8.32 $Y=1.82
+ $X2=7.65 $Y2=1.82
r81 24 69 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=7.65 $Y=1.14
+ $X2=8.32 $Y2=1.14
r82 19 21 48.6587 $w=2.23e-07 $l=9.5e-07 $layer=LI1_cond $X=7.537 $Y=1.96
+ $X2=7.537 $Y2=2.91
r83 17 26 6.9898 $w=1.7e-07 $l=1.49579e-07 $layer=LI1_cond $X=7.537 $Y=1.905
+ $X2=7.65 $Y2=1.82
r84 17 19 2.81708 $w=2.23e-07 $l=5.5e-08 $layer=LI1_cond $X=7.537 $Y=1.905
+ $X2=7.537 $Y2=1.96
r85 13 24 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=7.535 $Y=1.055
+ $X2=7.65 $Y2=1.14
r86 13 15 31.8174 $w=2.28e-07 $l=6.35e-07 $layer=LI1_cond $X=7.535 $Y=1.055
+ $X2=7.535 $Y2=0.42
r87 4 35 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=8.275
+ $Y=1.835 $X2=8.415 $Y2=2.91
r88 4 33 400 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=8.275
+ $Y=1.835 $X2=8.415 $Y2=1.96
r89 3 21 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=7.415
+ $Y=1.835 $X2=7.555 $Y2=2.91
r90 3 19 400 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=7.415
+ $Y=1.835 $X2=7.555 $Y2=1.96
r91 2 27 182 $w=1.7e-07 $l=7.81873e-07 $layer=licon1_NDIFF $count=1 $X=8.275
+ $Y=0.235 $X2=8.415 $Y2=0.95
r92 2 29 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=8.275
+ $Y=0.235 $X2=8.415 $Y2=0.42
r93 1 15 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=7.415
+ $Y=0.235 $X2=7.555 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__DFXTP_4%VGND 1 2 3 4 5 6 7 22 24 28 32 36 40 44 48
+ 50 52 55 56 57 59 71 78 83 92 95 98 101 105
r108 104 105 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=0
+ $X2=8.88 $Y2=0
r109 101 102 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=0
+ $X2=7.92 $Y2=0
r110 98 99 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r111 96 99 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.96
+ $Y2=0
r112 95 96 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6 $Y2=0
r113 92 93 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r114 89 90 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r115 87 105 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=0 $X2=8.88
+ $Y2=0
r116 87 102 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=0 $X2=7.92
+ $Y2=0
r117 86 87 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r118 84 101 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.15 $Y=0
+ $X2=7.985 $Y2=0
r119 84 86 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=8.15 $Y=0 $X2=8.4
+ $Y2=0
r120 83 104 4.746 $w=1.7e-07 $l=2.2e-07 $layer=LI1_cond $X=8.68 $Y=0 $X2=8.9
+ $Y2=0
r121 83 86 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=8.68 $Y=0 $X2=8.4
+ $Y2=0
r122 82 102 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0
+ $X2=7.92 $Y2=0
r123 82 99 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0 $X2=6.96
+ $Y2=0
r124 81 82 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r125 79 98 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=7.25 $Y=0 $X2=7.105
+ $Y2=0
r126 79 81 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=7.25 $Y=0 $X2=7.44
+ $Y2=0
r127 78 101 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.82 $Y=0
+ $X2=7.985 $Y2=0
r128 78 81 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=7.82 $Y=0 $X2=7.44
+ $Y2=0
r129 77 96 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=6
+ $Y2=0
r130 76 77 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r131 73 76 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=4.08 $Y=0 $X2=5.52
+ $Y2=0
r132 73 74 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r133 71 95 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.785 $Y=0 $X2=5.95
+ $Y2=0
r134 71 76 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=5.785 $Y=0
+ $X2=5.52 $Y2=0
r135 70 74 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r136 69 70 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r137 67 70 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.6
+ $Y2=0
r138 67 93 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.68
+ $Y2=0
r139 66 69 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=2.16 $Y=0 $X2=3.6
+ $Y2=0
r140 66 67 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r141 64 92 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.98 $Y=0 $X2=1.815
+ $Y2=0
r142 64 66 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=1.98 $Y=0 $X2=2.16
+ $Y2=0
r143 63 93 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r144 63 90 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r145 62 63 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r146 60 89 4.78091 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=0
+ $X2=0.212 $Y2=0
r147 60 62 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.425 $Y=0 $X2=0.72
+ $Y2=0
r148 59 92 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.65 $Y=0 $X2=1.815
+ $Y2=0
r149 59 62 60.6738 $w=1.68e-07 $l=9.3e-07 $layer=LI1_cond $X=1.65 $Y=0 $X2=0.72
+ $Y2=0
r150 57 77 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.52
+ $Y2=0
r151 57 74 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=4.08
+ $Y2=0
r152 55 69 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=3.705 $Y=0 $X2=3.6
+ $Y2=0
r153 55 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.705 $Y=0 $X2=3.87
+ $Y2=0
r154 54 73 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=4.035 $Y=0 $X2=4.08
+ $Y2=0
r155 54 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.035 $Y=0 $X2=3.87
+ $Y2=0
r156 50 104 3.02018 $w=3.3e-07 $l=1.09087e-07 $layer=LI1_cond $X=8.845 $Y=0.085
+ $X2=8.9 $Y2=0
r157 50 52 15.8897 $w=3.28e-07 $l=4.55e-07 $layer=LI1_cond $X=8.845 $Y=0.085
+ $X2=8.845 $Y2=0.54
r158 46 101 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.985 $Y=0.085
+ $X2=7.985 $Y2=0
r159 46 48 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=7.985 $Y=0.085
+ $X2=7.985 $Y2=0.36
r160 42 98 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=7.105 $Y=0.085
+ $X2=7.105 $Y2=0
r161 42 44 11.7231 $w=2.88e-07 $l=2.95e-07 $layer=LI1_cond $X=7.105 $Y=0.085
+ $X2=7.105 $Y2=0.38
r162 41 95 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.115 $Y=0 $X2=5.95
+ $Y2=0
r163 40 98 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=6.96 $Y=0 $X2=7.105
+ $Y2=0
r164 40 41 55.1283 $w=1.68e-07 $l=8.45e-07 $layer=LI1_cond $X=6.96 $Y=0
+ $X2=6.115 $Y2=0
r165 36 38 13.2706 $w=3.28e-07 $l=3.8e-07 $layer=LI1_cond $X=5.95 $Y=0.38
+ $X2=5.95 $Y2=0.76
r166 34 95 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.95 $Y=0.085
+ $X2=5.95 $Y2=0
r167 34 36 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=5.95 $Y=0.085
+ $X2=5.95 $Y2=0.38
r168 30 56 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.87 $Y=0.085
+ $X2=3.87 $Y2=0
r169 30 32 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=3.87 $Y=0.085
+ $X2=3.87 $Y2=0.795
r170 26 92 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.815 $Y=0.085
+ $X2=1.815 $Y2=0
r171 26 28 25.1442 $w=3.28e-07 $l=7.2e-07 $layer=LI1_cond $X=1.815 $Y=0.085
+ $X2=1.815 $Y2=0.805
r172 22 89 2.98526 $w=3.3e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.212 $Y2=0
r173 22 24 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.26 $Y2=0.505
r174 7 52 182 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_NDIFF $count=1 $X=8.705
+ $Y=0.235 $X2=8.845 $Y2=0.54
r175 6 48 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=7.845
+ $Y=0.235 $X2=7.985 $Y2=0.36
r176 5 44 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=7
+ $Y=0.235 $X2=7.125 $Y2=0.38
r177 4 38 182 $w=1.7e-07 $l=3.11769e-07 $layer=licon1_NDIFF $count=1 $X=5.71
+ $Y=0.595 $X2=5.95 $Y2=0.76
r178 4 36 182 $w=1.7e-07 $l=3.30454e-07 $layer=licon1_NDIFF $count=1 $X=5.71
+ $Y=0.595 $X2=5.95 $Y2=0.38
r179 3 32 182 $w=1.7e-07 $l=3.87298e-07 $layer=licon1_NDIFF $count=1 $X=3.57
+ $Y=0.595 $X2=3.87 $Y2=0.795
r180 2 28 182 $w=1.7e-07 $l=2.93428e-07 $layer=licon1_NDIFF $count=1 $X=1.615
+ $Y=0.595 $X2=1.815 $Y2=0.805
r181 1 24 182 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.35 $X2=0.26 $Y2=0.505
.ends

