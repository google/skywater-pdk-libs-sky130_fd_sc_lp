* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__o2bb2ai_lp A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
X0 a_145_419# A2_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X1 a_400_83# B2 VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 VGND B1 a_400_83# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 a_490_419# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X4 Y B2 a_490_419# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X5 VPWR a_145_419# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X6 a_114_57# A2_N a_145_419# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 VGND A1_N a_114_57# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 Y a_145_419# a_400_83# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 VPWR A1_N a_145_419# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
.ends
