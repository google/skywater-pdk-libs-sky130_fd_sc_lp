* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__and3b_lp A_N B C VGND VNB VPB VPWR X
X0 a_248_409# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X1 a_666_57# a_248_409# X VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 a_391_57# B a_469_57# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 a_248_409# a_137_408# a_391_57# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 VPWR a_248_409# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X5 VGND a_248_409# a_666_57# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 VPWR B a_248_409# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X7 VPWR A_N a_137_408# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X8 a_114_57# A_N a_137_408# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 a_248_409# a_137_408# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X10 VGND A_N a_114_57# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X11 a_469_57# C VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
