* File: sky130_fd_sc_lp__a31o_1.pxi.spice
* Created: Wed Sep  2 09:26:18 2020
* 
x_PM_SKY130_FD_SC_LP__A31O_1%A_80_21# N_A_80_21#_M1007_d N_A_80_21#_M1006_d
+ N_A_80_21#_M1004_g N_A_80_21#_M1001_g N_A_80_21#_c_54_n N_A_80_21#_c_55_n
+ N_A_80_21#_c_65_p N_A_80_21#_c_114_p N_A_80_21#_c_121_p N_A_80_21#_c_56_n
+ N_A_80_21#_c_60_n N_A_80_21#_c_81_p N_A_80_21#_c_61_n N_A_80_21#_c_57_n
+ N_A_80_21#_c_58_n PM_SKY130_FD_SC_LP__A31O_1%A_80_21#
x_PM_SKY130_FD_SC_LP__A31O_1%A3 N_A3_M1002_g N_A3_M1005_g A3 A3 A3 A3 A3
+ N_A3_c_129_n N_A3_c_130_n A3 PM_SKY130_FD_SC_LP__A31O_1%A3
x_PM_SKY130_FD_SC_LP__A31O_1%A2 N_A2_M1003_g N_A2_M1009_g A2 N_A2_c_172_n
+ N_A2_c_173_n PM_SKY130_FD_SC_LP__A31O_1%A2
x_PM_SKY130_FD_SC_LP__A31O_1%A1 N_A1_M1007_g N_A1_M1000_g A1 N_A1_c_210_n
+ N_A1_c_211_n PM_SKY130_FD_SC_LP__A31O_1%A1
x_PM_SKY130_FD_SC_LP__A31O_1%B1 N_B1_M1008_g N_B1_M1006_g B1 N_B1_c_244_n
+ N_B1_c_245_n PM_SKY130_FD_SC_LP__A31O_1%B1
x_PM_SKY130_FD_SC_LP__A31O_1%X N_X_M1004_s N_X_M1001_s X X X X X X X N_X_c_271_n
+ X PM_SKY130_FD_SC_LP__A31O_1%X
x_PM_SKY130_FD_SC_LP__A31O_1%VPWR N_VPWR_M1001_d N_VPWR_M1009_d N_VPWR_c_288_n
+ N_VPWR_c_289_n VPWR N_VPWR_c_290_n N_VPWR_c_291_n N_VPWR_c_292_n
+ N_VPWR_c_287_n N_VPWR_c_294_n N_VPWR_c_295_n PM_SKY130_FD_SC_LP__A31O_1%VPWR
x_PM_SKY130_FD_SC_LP__A31O_1%A_269_367# N_A_269_367#_M1005_d
+ N_A_269_367#_M1000_d N_A_269_367#_c_339_n N_A_269_367#_c_332_n
+ N_A_269_367#_c_333_n N_A_269_367#_c_350_n
+ PM_SKY130_FD_SC_LP__A31O_1%A_269_367#
x_PM_SKY130_FD_SC_LP__A31O_1%VGND N_VGND_M1004_d N_VGND_M1008_d N_VGND_c_367_n
+ N_VGND_c_368_n VGND N_VGND_c_369_n N_VGND_c_370_n N_VGND_c_371_n
+ PM_SKY130_FD_SC_LP__A31O_1%VGND
cc_1 VNB N_A_80_21#_M1001_g 0.00904986f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=2.465
cc_2 VNB N_A_80_21#_c_54_n 0.00445611f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.35
cc_3 VNB N_A_80_21#_c_55_n 0.0394763f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.35
cc_4 VNB N_A_80_21#_c_56_n 0.0148526f $X=-0.19 $Y=-0.245 $X2=3.095 $Y2=0.955
cc_5 VNB N_A_80_21#_c_57_n 0.0295944f $X=-0.19 $Y=-0.245 $X2=3.047 $Y2=1.815
cc_6 VNB N_A_80_21#_c_58_n 0.0208967f $X=-0.19 $Y=-0.245 $X2=0.582 $Y2=1.185
cc_7 VNB N_A3_M1002_g 0.0198586f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A3_M1005_g 0.0067552f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.185
cc_9 VNB N_A3_c_129_n 0.032555f $X=-0.19 $Y=-0.245 $X2=2.455 $Y2=0.87
cc_10 VNB N_A3_c_130_n 0.0124759f $X=-0.19 $Y=-0.245 $X2=3.095 $Y2=0.955
cc_11 VNB N_A2_M1009_g 0.00829997f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB A2 0.00172691f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.655
cc_13 VNB N_A2_c_172_n 0.0324803f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=2.465
cc_14 VNB N_A2_c_173_n 0.0172361f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A1_M1007_g 0.0199847f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A1_M1000_g 0.00668834f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.185
cc_17 VNB N_A1_c_210_n 0.0299794f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=2.465
cc_18 VNB N_A1_c_211_n 0.00340285f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_B1_M1008_g 0.0214514f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_B1_M1006_g 0.00673451f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.185
cc_21 VNB N_B1_c_244_n 0.032019f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=2.465
cc_22 VNB N_B1_c_245_n 0.00429971f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_X_c_271_n 0.0617615f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_VPWR_c_287_n 0.143779f $X=-0.19 $Y=-0.245 $X2=3.047 $Y2=1.98
cc_25 VNB N_VGND_c_367_n 0.0149909f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.185
cc_26 VNB N_VGND_c_368_n 0.0209684f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.655
cc_27 VNB N_VGND_c_369_n 0.0284376f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_370_n 0.0447435f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_371_n 0.193611f $X=-0.19 $Y=-0.245 $X2=3.047 $Y2=1.98
cc_30 VPB N_A_80_21#_M1001_g 0.0264898f $X=-0.19 $Y=1.655 $X2=0.515 $Y2=2.465
cc_31 VPB N_A_80_21#_c_60_n 0.0418028f $X=-0.19 $Y=1.655 $X2=2.955 $Y2=2.91
cc_32 VPB N_A_80_21#_c_61_n 0.0195225f $X=-0.19 $Y=1.655 $X2=2.955 $Y2=1.98
cc_33 VPB N_A_80_21#_c_57_n 0.00792896f $X=-0.19 $Y=1.655 $X2=3.047 $Y2=1.815
cc_34 VPB N_A3_M1005_g 0.0229001f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=1.185
cc_35 VPB A3 0.00223428f $X=-0.19 $Y=1.655 $X2=2.975 $Y2=1.985
cc_36 VPB N_A2_M1009_g 0.0210427f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_37 VPB N_A1_M1000_g 0.0204067f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=1.185
cc_38 VPB N_B1_M1006_g 0.0238948f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=1.185
cc_39 VPB X 0.0113483f $X=-0.19 $Y=1.655 $X2=0.515 $Y2=1.515
cc_40 VPB X 0.0499201f $X=-0.19 $Y=1.655 $X2=0.515 $Y2=2.465
cc_41 VPB N_X_c_271_n 0.00215052f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_42 VPB N_VPWR_c_288_n 0.013546f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.655
cc_43 VPB N_VPWR_c_289_n 0.00552886f $X=-0.19 $Y=1.655 $X2=0.64 $Y2=1.35
cc_44 VPB N_VPWR_c_290_n 0.0190404f $X=-0.19 $Y=1.655 $X2=2.455 $Y2=0.87
cc_45 VPB N_VPWR_c_291_n 0.0263291f $X=-0.19 $Y=1.655 $X2=2.62 $Y2=0.955
cc_46 VPB N_VPWR_c_292_n 0.0336276f $X=-0.19 $Y=1.655 $X2=2.455 $Y2=0.955
cc_47 VPB N_VPWR_c_287_n 0.050716f $X=-0.19 $Y=1.655 $X2=3.047 $Y2=1.98
cc_48 VPB N_VPWR_c_294_n 0.00574453f $X=-0.19 $Y=1.655 $X2=3.047 $Y2=1.985
cc_49 VPB N_VPWR_c_295_n 0.00631492f $X=-0.19 $Y=1.655 $X2=0.582 $Y2=1.515
cc_50 VPB N_A_269_367#_c_332_n 0.00944826f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_51 VPB N_A_269_367#_c_333_n 0.00345366f $X=-0.19 $Y=1.655 $X2=0.64 $Y2=1.04
cc_52 N_A_80_21#_c_54_n N_A3_M1002_g 0.00283135f $X=0.6 $Y=1.35 $X2=0 $Y2=0
cc_53 N_A_80_21#_c_55_n N_A3_M1002_g 7.63004e-19 $X=0.6 $Y=1.35 $X2=0 $Y2=0
cc_54 N_A_80_21#_c_65_p N_A3_M1002_g 0.0153845f $X=2.29 $Y=0.955 $X2=0 $Y2=0
cc_55 N_A_80_21#_c_58_n N_A3_M1002_g 0.00924028f $X=0.582 $Y=1.185 $X2=0 $Y2=0
cc_56 N_A_80_21#_M1001_g N_A3_M1005_g 0.0212312f $X=0.515 $Y=2.465 $X2=0 $Y2=0
cc_57 N_A_80_21#_M1001_g N_A3_c_129_n 6.78363e-19 $X=0.515 $Y=2.465 $X2=0 $Y2=0
cc_58 N_A_80_21#_c_54_n N_A3_c_129_n 3.86049e-19 $X=0.6 $Y=1.35 $X2=0 $Y2=0
cc_59 N_A_80_21#_c_55_n N_A3_c_129_n 0.0193397f $X=0.6 $Y=1.35 $X2=0 $Y2=0
cc_60 N_A_80_21#_c_65_p N_A3_c_129_n 0.00142651f $X=2.29 $Y=0.955 $X2=0 $Y2=0
cc_61 N_A_80_21#_M1001_g N_A3_c_130_n 0.00111712f $X=0.515 $Y=2.465 $X2=0 $Y2=0
cc_62 N_A_80_21#_c_54_n N_A3_c_130_n 0.0191781f $X=0.6 $Y=1.35 $X2=0 $Y2=0
cc_63 N_A_80_21#_c_55_n N_A3_c_130_n 0.00108352f $X=0.6 $Y=1.35 $X2=0 $Y2=0
cc_64 N_A_80_21#_c_65_p N_A3_c_130_n 0.0260435f $X=2.29 $Y=0.955 $X2=0 $Y2=0
cc_65 N_A_80_21#_M1001_g A3 0.00399346f $X=0.515 $Y=2.465 $X2=0 $Y2=0
cc_66 N_A_80_21#_c_65_p A2 0.0206931f $X=2.29 $Y=0.955 $X2=0 $Y2=0
cc_67 N_A_80_21#_c_65_p N_A2_c_172_n 0.00372033f $X=2.29 $Y=0.955 $X2=0 $Y2=0
cc_68 N_A_80_21#_c_65_p N_A2_c_173_n 0.0152912f $X=2.29 $Y=0.955 $X2=0 $Y2=0
cc_69 N_A_80_21#_c_65_p N_A1_M1007_g 0.0135135f $X=2.29 $Y=0.955 $X2=0 $Y2=0
cc_70 N_A_80_21#_c_81_p N_A1_c_210_n 0.00464005f $X=2.455 $Y=0.955 $X2=0 $Y2=0
cc_71 N_A_80_21#_c_65_p N_A1_c_211_n 0.0146274f $X=2.29 $Y=0.955 $X2=0 $Y2=0
cc_72 N_A_80_21#_c_81_p N_A1_c_211_n 0.00513439f $X=2.455 $Y=0.955 $X2=0 $Y2=0
cc_73 N_A_80_21#_c_56_n N_B1_M1008_g 0.0165568f $X=3.095 $Y=0.955 $X2=0 $Y2=0
cc_74 N_A_80_21#_c_57_n N_B1_M1008_g 0.00514335f $X=3.047 $Y=1.815 $X2=0 $Y2=0
cc_75 N_A_80_21#_c_61_n N_B1_M1006_g 0.00347437f $X=2.955 $Y=1.98 $X2=0 $Y2=0
cc_76 N_A_80_21#_c_57_n N_B1_M1006_g 0.00716275f $X=3.047 $Y=1.815 $X2=0 $Y2=0
cc_77 N_A_80_21#_c_56_n N_B1_c_244_n 0.00497085f $X=3.095 $Y=0.955 $X2=0 $Y2=0
cc_78 N_A_80_21#_c_61_n N_B1_c_244_n 0.00484439f $X=2.955 $Y=1.98 $X2=0 $Y2=0
cc_79 N_A_80_21#_c_57_n N_B1_c_244_n 0.00806477f $X=3.047 $Y=1.815 $X2=0 $Y2=0
cc_80 N_A_80_21#_c_56_n N_B1_c_245_n 0.0186376f $X=3.095 $Y=0.955 $X2=0 $Y2=0
cc_81 N_A_80_21#_c_81_p N_B1_c_245_n 0.00596323f $X=2.455 $Y=0.955 $X2=0 $Y2=0
cc_82 N_A_80_21#_c_61_n N_B1_c_245_n 0.00554074f $X=2.955 $Y=1.98 $X2=0 $Y2=0
cc_83 N_A_80_21#_c_57_n N_B1_c_245_n 0.0250393f $X=3.047 $Y=1.815 $X2=0 $Y2=0
cc_84 N_A_80_21#_M1001_g X 0.00854845f $X=0.515 $Y=2.465 $X2=0 $Y2=0
cc_85 N_A_80_21#_M1001_g N_X_c_271_n 0.00541643f $X=0.515 $Y=2.465 $X2=0 $Y2=0
cc_86 N_A_80_21#_c_54_n N_X_c_271_n 0.0346263f $X=0.6 $Y=1.35 $X2=0 $Y2=0
cc_87 N_A_80_21#_c_58_n N_X_c_271_n 0.0134745f $X=0.582 $Y=1.185 $X2=0 $Y2=0
cc_88 N_A_80_21#_M1001_g N_VPWR_c_288_n 0.0140797f $X=0.515 $Y=2.465 $X2=0 $Y2=0
cc_89 N_A_80_21#_c_54_n N_VPWR_c_288_n 0.00800468f $X=0.6 $Y=1.35 $X2=0 $Y2=0
cc_90 N_A_80_21#_c_55_n N_VPWR_c_288_n 0.00101857f $X=0.6 $Y=1.35 $X2=0 $Y2=0
cc_91 N_A_80_21#_M1001_g N_VPWR_c_290_n 0.00585385f $X=0.515 $Y=2.465 $X2=0
+ $Y2=0
cc_92 N_A_80_21#_c_60_n N_VPWR_c_292_n 0.0188755f $X=2.955 $Y=2.91 $X2=0 $Y2=0
cc_93 N_A_80_21#_M1006_d N_VPWR_c_287_n 0.0026734f $X=2.815 $Y=1.835 $X2=0 $Y2=0
cc_94 N_A_80_21#_M1001_g N_VPWR_c_287_n 0.0123355f $X=0.515 $Y=2.465 $X2=0 $Y2=0
cc_95 N_A_80_21#_c_60_n N_VPWR_c_287_n 0.0111968f $X=2.955 $Y=2.91 $X2=0 $Y2=0
cc_96 N_A_80_21#_c_65_p N_A_269_367#_c_332_n 0.00468023f $X=2.29 $Y=0.955 $X2=0
+ $Y2=0
cc_97 N_A_80_21#_c_81_p N_A_269_367#_c_332_n 0.00566963f $X=2.455 $Y=0.955 $X2=0
+ $Y2=0
cc_98 N_A_80_21#_c_61_n N_A_269_367#_c_332_n 0.00171339f $X=2.955 $Y=1.98 $X2=0
+ $Y2=0
cc_99 N_A_80_21#_c_57_n N_A_269_367#_c_332_n 0.00457744f $X=3.047 $Y=1.815 $X2=0
+ $Y2=0
cc_100 N_A_80_21#_c_65_p N_A_269_367#_c_333_n 0.00274698f $X=2.29 $Y=0.955 $X2=0
+ $Y2=0
cc_101 N_A_80_21#_c_54_n N_VGND_M1004_d 5.15458e-19 $X=0.6 $Y=1.35 $X2=-0.19
+ $Y2=-0.245
cc_102 N_A_80_21#_c_65_p N_VGND_M1004_d 0.0152352f $X=2.29 $Y=0.955 $X2=-0.19
+ $Y2=-0.245
cc_103 N_A_80_21#_c_114_p N_VGND_M1004_d 0.00199613f $X=0.765 $Y=0.955 $X2=-0.19
+ $Y2=-0.245
cc_104 N_A_80_21#_c_56_n N_VGND_M1008_d 0.00746251f $X=3.095 $Y=0.955 $X2=0
+ $Y2=0
cc_105 N_A_80_21#_c_56_n N_VGND_c_368_n 0.0221865f $X=3.095 $Y=0.955 $X2=0 $Y2=0
cc_106 N_A_80_21#_c_55_n N_VGND_c_369_n 7.65158e-19 $X=0.6 $Y=1.35 $X2=0 $Y2=0
cc_107 N_A_80_21#_c_65_p N_VGND_c_369_n 0.0320963f $X=2.29 $Y=0.955 $X2=0 $Y2=0
cc_108 N_A_80_21#_c_114_p N_VGND_c_369_n 0.0161715f $X=0.765 $Y=0.955 $X2=0
+ $Y2=0
cc_109 N_A_80_21#_c_58_n N_VGND_c_369_n 0.0194953f $X=0.582 $Y=1.185 $X2=0 $Y2=0
cc_110 N_A_80_21#_c_121_p N_VGND_c_370_n 0.0212513f $X=2.455 $Y=0.42 $X2=0 $Y2=0
cc_111 N_A_80_21#_M1007_d N_VGND_c_371_n 0.00526034f $X=2.275 $Y=0.235 $X2=0
+ $Y2=0
cc_112 N_A_80_21#_c_121_p N_VGND_c_371_n 0.0127519f $X=2.455 $Y=0.42 $X2=0 $Y2=0
cc_113 N_A_80_21#_c_58_n N_VGND_c_371_n 0.00917991f $X=0.582 $Y=1.185 $X2=0
+ $Y2=0
cc_114 N_A_80_21#_c_65_p A_269_47# 0.00836926f $X=2.29 $Y=0.955 $X2=-0.19
+ $Y2=-0.245
cc_115 N_A_80_21#_c_65_p A_347_47# 0.0152834f $X=2.29 $Y=0.955 $X2=-0.19
+ $Y2=-0.245
cc_116 N_A3_c_129_n N_A2_M1009_g 0.0211504f $X=1.18 $Y=1.375 $X2=0 $Y2=0
cc_117 N_A3_c_130_n N_A2_M1009_g 7.08578e-19 $X=1.19 $Y=1.645 $X2=0 $Y2=0
cc_118 A3 N_A2_M1009_g 8.3746e-19 $X=1.2 $Y=1.665 $X2=0 $Y2=0
cc_119 N_A3_c_129_n A2 3.84693e-19 $X=1.18 $Y=1.375 $X2=0 $Y2=0
cc_120 N_A3_c_130_n A2 0.0195822f $X=1.19 $Y=1.645 $X2=0 $Y2=0
cc_121 N_A3_M1002_g N_A2_c_172_n 0.0209173f $X=1.27 $Y=0.655 $X2=0 $Y2=0
cc_122 N_A3_c_130_n N_A2_c_172_n 0.00106329f $X=1.19 $Y=1.645 $X2=0 $Y2=0
cc_123 N_A3_M1002_g N_A2_c_173_n 0.0603133f $X=1.27 $Y=0.655 $X2=0 $Y2=0
cc_124 N_A3_c_130_n N_X_c_271_n 0.00411838f $X=1.19 $Y=1.645 $X2=0 $Y2=0
cc_125 A3 N_VPWR_M1001_d 0.0103679f $X=1.2 $Y=1.665 $X2=-0.19 $Y2=-0.245
cc_126 N_A3_M1005_g N_VPWR_c_288_n 0.00838103f $X=1.27 $Y=2.465 $X2=0 $Y2=0
cc_127 A3 N_VPWR_c_288_n 0.0799637f $X=1.2 $Y=1.665 $X2=0 $Y2=0
cc_128 N_A3_M1005_g N_VPWR_c_291_n 0.00474558f $X=1.27 $Y=2.465 $X2=0 $Y2=0
cc_129 A3 N_VPWR_c_291_n 0.00453673f $X=1.2 $Y=1.665 $X2=0 $Y2=0
cc_130 N_A3_M1005_g N_VPWR_c_287_n 0.00853686f $X=1.27 $Y=2.465 $X2=0 $Y2=0
cc_131 A3 N_VPWR_c_287_n 0.00597535f $X=1.2 $Y=1.665 $X2=0 $Y2=0
cc_132 N_A3_M1005_g N_A_269_367#_c_339_n 0.00483201f $X=1.27 $Y=2.465 $X2=0
+ $Y2=0
cc_133 A3 N_A_269_367#_c_339_n 0.0712223f $X=1.2 $Y=1.665 $X2=0 $Y2=0
cc_134 N_A3_M1005_g N_A_269_367#_c_333_n 0.00113639f $X=1.27 $Y=2.465 $X2=0
+ $Y2=0
cc_135 A3 N_A_269_367#_c_333_n 0.0137364f $X=1.2 $Y=1.665 $X2=0 $Y2=0
cc_136 N_A3_M1002_g N_VGND_c_369_n 0.0179901f $X=1.27 $Y=0.655 $X2=0 $Y2=0
cc_137 N_A3_M1002_g N_VGND_c_370_n 0.00487821f $X=1.27 $Y=0.655 $X2=0 $Y2=0
cc_138 N_A3_M1002_g N_VGND_c_371_n 0.00827387f $X=1.27 $Y=0.655 $X2=0 $Y2=0
cc_139 N_A2_c_172_n N_A1_M1007_g 0.0176039f $X=1.72 $Y=1.35 $X2=0 $Y2=0
cc_140 N_A2_c_173_n N_A1_M1007_g 0.0357134f $X=1.72 $Y=1.185 $X2=0 $Y2=0
cc_141 N_A2_M1009_g N_A1_M1000_g 0.040634f $X=1.755 $Y=2.465 $X2=0 $Y2=0
cc_142 N_A2_M1009_g N_A1_c_210_n 9.5668e-19 $X=1.755 $Y=2.465 $X2=0 $Y2=0
cc_143 A2 N_A1_c_210_n 3.3573e-19 $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_144 N_A2_M1009_g N_A1_c_211_n 5.27374e-19 $X=1.755 $Y=2.465 $X2=0 $Y2=0
cc_145 A2 N_A1_c_211_n 0.0241183f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_146 N_A2_c_172_n N_A1_c_211_n 0.00182964f $X=1.72 $Y=1.35 $X2=0 $Y2=0
cc_147 N_A2_M1009_g N_VPWR_c_289_n 0.00948651f $X=1.755 $Y=2.465 $X2=0 $Y2=0
cc_148 N_A2_M1009_g N_VPWR_c_291_n 0.00564131f $X=1.755 $Y=2.465 $X2=0 $Y2=0
cc_149 N_A2_M1009_g N_VPWR_c_287_n 0.0106885f $X=1.755 $Y=2.465 $X2=0 $Y2=0
cc_150 N_A2_M1009_g N_A_269_367#_c_339_n 0.0148278f $X=1.755 $Y=2.465 $X2=0
+ $Y2=0
cc_151 N_A2_M1009_g N_A_269_367#_c_332_n 0.0126032f $X=1.755 $Y=2.465 $X2=0
+ $Y2=0
cc_152 A2 N_A_269_367#_c_332_n 0.0122474f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_153 N_A2_c_172_n N_A_269_367#_c_332_n 3.69604e-19 $X=1.72 $Y=1.35 $X2=0 $Y2=0
cc_154 N_A2_M1009_g N_A_269_367#_c_333_n 0.00174543f $X=1.755 $Y=2.465 $X2=0
+ $Y2=0
cc_155 A2 N_A_269_367#_c_333_n 0.0104945f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_156 N_A2_c_172_n N_A_269_367#_c_333_n 9.56168e-19 $X=1.72 $Y=1.35 $X2=0 $Y2=0
cc_157 N_A2_M1009_g N_A_269_367#_c_350_n 7.37178e-19 $X=1.755 $Y=2.465 $X2=0
+ $Y2=0
cc_158 N_A2_c_173_n N_VGND_c_369_n 0.00343491f $X=1.72 $Y=1.185 $X2=0 $Y2=0
cc_159 N_A2_c_173_n N_VGND_c_370_n 0.00585385f $X=1.72 $Y=1.185 $X2=0 $Y2=0
cc_160 N_A2_c_173_n N_VGND_c_371_n 0.0111877f $X=1.72 $Y=1.185 $X2=0 $Y2=0
cc_161 N_A1_M1007_g N_B1_M1008_g 0.0204145f $X=2.2 $Y=0.655 $X2=0 $Y2=0
cc_162 N_A1_M1000_g N_B1_M1006_g 0.0261021f $X=2.31 $Y=2.465 $X2=0 $Y2=0
cc_163 N_A1_c_210_n N_B1_c_244_n 0.0204448f $X=2.29 $Y=1.375 $X2=0 $Y2=0
cc_164 N_A1_c_211_n N_B1_c_244_n 2.86088e-19 $X=2.29 $Y=1.375 $X2=0 $Y2=0
cc_165 N_A1_c_210_n N_B1_c_245_n 0.00220085f $X=2.29 $Y=1.375 $X2=0 $Y2=0
cc_166 N_A1_c_211_n N_B1_c_245_n 0.0264486f $X=2.29 $Y=1.375 $X2=0 $Y2=0
cc_167 N_A1_M1000_g N_VPWR_c_289_n 0.00939157f $X=2.31 $Y=2.465 $X2=0 $Y2=0
cc_168 N_A1_M1000_g N_VPWR_c_292_n 0.0055654f $X=2.31 $Y=2.465 $X2=0 $Y2=0
cc_169 N_A1_M1000_g N_VPWR_c_287_n 0.0103898f $X=2.31 $Y=2.465 $X2=0 $Y2=0
cc_170 N_A1_M1000_g N_A_269_367#_c_339_n 7.31705e-19 $X=2.31 $Y=2.465 $X2=0
+ $Y2=0
cc_171 N_A1_M1000_g N_A_269_367#_c_332_n 0.0140623f $X=2.31 $Y=2.465 $X2=0 $Y2=0
cc_172 N_A1_c_210_n N_A_269_367#_c_332_n 0.0050112f $X=2.29 $Y=1.375 $X2=0 $Y2=0
cc_173 N_A1_c_211_n N_A_269_367#_c_332_n 0.0238652f $X=2.29 $Y=1.375 $X2=0 $Y2=0
cc_174 N_A1_M1000_g N_A_269_367#_c_350_n 0.0152355f $X=2.31 $Y=2.465 $X2=0 $Y2=0
cc_175 N_A1_M1007_g N_VGND_c_368_n 0.00103262f $X=2.2 $Y=0.655 $X2=0 $Y2=0
cc_176 N_A1_M1007_g N_VGND_c_370_n 0.00585385f $X=2.2 $Y=0.655 $X2=0 $Y2=0
cc_177 N_A1_M1007_g N_VGND_c_371_n 0.0114286f $X=2.2 $Y=0.655 $X2=0 $Y2=0
cc_178 N_B1_M1006_g N_VPWR_c_292_n 0.00585385f $X=2.74 $Y=2.465 $X2=0 $Y2=0
cc_179 N_B1_M1006_g N_VPWR_c_287_n 0.0118344f $X=2.74 $Y=2.465 $X2=0 $Y2=0
cc_180 N_B1_M1006_g N_A_269_367#_c_332_n 0.00168941f $X=2.74 $Y=2.465 $X2=0
+ $Y2=0
cc_181 N_B1_c_245_n N_A_269_367#_c_332_n 0.0101731f $X=2.83 $Y=1.375 $X2=0 $Y2=0
cc_182 N_B1_M1008_g N_VGND_c_368_n 0.0141222f $X=2.74 $Y=0.655 $X2=0 $Y2=0
cc_183 N_B1_M1008_g N_VGND_c_370_n 0.00486043f $X=2.74 $Y=0.655 $X2=0 $Y2=0
cc_184 N_B1_M1008_g N_VGND_c_371_n 0.00864313f $X=2.74 $Y=0.655 $X2=0 $Y2=0
cc_185 X N_VPWR_c_288_n 0.00130678f $X=0.155 $Y=1.58 $X2=0 $Y2=0
cc_186 X N_VPWR_c_290_n 0.0217502f $X=0.155 $Y=1.95 $X2=0 $Y2=0
cc_187 N_X_M1001_s N_VPWR_c_287_n 0.00336915f $X=0.175 $Y=1.835 $X2=0 $Y2=0
cc_188 X N_VPWR_c_287_n 0.0123631f $X=0.155 $Y=1.95 $X2=0 $Y2=0
cc_189 N_X_c_271_n N_VGND_c_369_n 0.0181731f $X=0.26 $Y=0.42 $X2=0 $Y2=0
cc_190 N_X_M1004_s N_VGND_c_371_n 0.0040649f $X=0.135 $Y=0.235 $X2=0 $Y2=0
cc_191 N_X_c_271_n N_VGND_c_371_n 0.0100252f $X=0.26 $Y=0.42 $X2=0 $Y2=0
cc_192 N_VPWR_c_287_n N_A_269_367#_M1005_d 0.00650451f $X=3.12 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_193 N_VPWR_c_287_n N_A_269_367#_M1000_d 0.00240953f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_194 N_VPWR_c_288_n N_A_269_367#_c_339_n 0.00716179f $X=0.81 $Y=1.98 $X2=0
+ $Y2=0
cc_195 N_VPWR_c_291_n N_A_269_367#_c_339_n 0.0146863f $X=1.865 $Y=3.33 $X2=0
+ $Y2=0
cc_196 N_VPWR_c_287_n N_A_269_367#_c_339_n 0.00911565f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_197 N_VPWR_M1009_d N_A_269_367#_c_332_n 0.00320298f $X=1.83 $Y=1.835 $X2=0
+ $Y2=0
cc_198 N_VPWR_c_289_n N_A_269_367#_c_332_n 0.0236753f $X=2.03 $Y=2.135 $X2=0
+ $Y2=0
cc_199 N_VPWR_c_292_n N_A_269_367#_c_350_n 0.0167664f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_200 N_VPWR_c_287_n N_A_269_367#_c_350_n 0.011231f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_201 N_VGND_c_371_n A_269_47# 0.010279f $X=3.12 $Y=0 $X2=-0.19 $Y2=-0.245
cc_202 N_VGND_c_371_n A_347_47# 0.0167135f $X=3.12 $Y=0 $X2=-0.19 $Y2=-0.245
