* File: sky130_fd_sc_lp__inv_8.pex.spice
* Created: Fri Aug 28 10:38:29 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__INV_8%A 3 7 11 15 19 23 27 31 35 39 43 47 51 55 59
+ 63 65 75 78 94
r142 91 92 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=2.88 $Y=1.48
+ $X2=3.31 $Y2=1.48
r143 90 91 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=2.45 $Y=1.48
+ $X2=2.88 $Y2=1.48
r144 88 90 27.9778 $w=3.3e-07 $l=1.6e-07 $layer=POLY_cond $X=2.29 $Y=1.48
+ $X2=2.45 $Y2=1.48
r145 88 89 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=2.29
+ $Y=1.48 $X2=2.29 $Y2=1.48
r146 86 88 47.2125 $w=3.3e-07 $l=2.7e-07 $layer=POLY_cond $X=2.02 $Y=1.48
+ $X2=2.29 $Y2=1.48
r147 83 84 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=1.16 $Y=1.48
+ $X2=1.59 $Y2=1.48
r148 82 83 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=0.73 $Y=1.48
+ $X2=1.16 $Y2=1.48
r149 78 89 6.99023 $w=3.03e-07 $l=1.85e-07 $layer=LI1_cond $X=2.212 $Y=1.295
+ $X2=2.212 $Y2=1.48
r150 76 94 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=3.65 $Y=1.48 $X2=3.74
+ $Y2=1.48
r151 76 92 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=3.65 $Y=1.48
+ $X2=3.31 $Y2=1.48
r152 75 76 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=3.65
+ $Y=1.48 $X2=3.65 $Y2=1.48
r153 73 89 3.20691 $w=2e-07 $l=1.5548e-07 $layer=LI1_cond $X=2.365 $Y=1.485
+ $X2=2.212 $Y2=1.48
r154 73 75 71.2591 $w=1.98e-07 $l=1.285e-06 $layer=LI1_cond $X=2.365 $Y=1.485
+ $X2=3.65 $Y2=1.485
r155 72 86 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=1.95 $Y=1.48 $X2=2.02
+ $Y2=1.48
r156 72 84 62.9501 $w=3.3e-07 $l=3.6e-07 $layer=POLY_cond $X=1.95 $Y=1.48
+ $X2=1.59 $Y2=1.48
r157 71 72 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=1.95
+ $Y=1.48 $X2=1.95 $Y2=1.48
r158 68 82 24.4806 $w=3.3e-07 $l=1.4e-07 $layer=POLY_cond $X=0.59 $Y=1.48
+ $X2=0.73 $Y2=1.48
r159 67 71 79.3876 $w=1.88e-07 $l=1.36e-06 $layer=LI1_cond $X=0.59 $Y=1.49
+ $X2=1.95 $Y2=1.49
r160 67 68 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=0.59
+ $Y=1.48 $X2=0.59 $Y2=1.48
r161 65 89 0.37785 $w=3.03e-07 $l=1e-08 $layer=LI1_cond $X=2.212 $Y=1.49
+ $X2=2.212 $Y2=1.48
r162 65 71 6.42105 $w=1.88e-07 $l=1.1e-07 $layer=LI1_cond $X=2.06 $Y=1.49
+ $X2=1.95 $Y2=1.49
r163 61 94 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.74 $Y=1.645
+ $X2=3.74 $Y2=1.48
r164 61 63 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=3.74 $Y=1.645
+ $X2=3.74 $Y2=2.465
r165 57 94 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.74 $Y=1.315
+ $X2=3.74 $Y2=1.48
r166 57 59 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.74 $Y=1.315
+ $X2=3.74 $Y2=0.655
r167 53 92 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.31 $Y=1.645
+ $X2=3.31 $Y2=1.48
r168 53 55 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=3.31 $Y=1.645
+ $X2=3.31 $Y2=2.465
r169 49 92 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.31 $Y=1.315
+ $X2=3.31 $Y2=1.48
r170 49 51 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.31 $Y=1.315
+ $X2=3.31 $Y2=0.655
r171 45 91 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.88 $Y=1.645
+ $X2=2.88 $Y2=1.48
r172 45 47 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=2.88 $Y=1.645
+ $X2=2.88 $Y2=2.465
r173 41 91 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.88 $Y=1.315
+ $X2=2.88 $Y2=1.48
r174 41 43 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.88 $Y=1.315
+ $X2=2.88 $Y2=0.655
r175 37 90 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.45 $Y=1.645
+ $X2=2.45 $Y2=1.48
r176 37 39 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=2.45 $Y=1.645
+ $X2=2.45 $Y2=2.465
r177 33 90 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.45 $Y=1.315
+ $X2=2.45 $Y2=1.48
r178 33 35 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.45 $Y=1.315
+ $X2=2.45 $Y2=0.655
r179 29 86 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.02 $Y=1.645
+ $X2=2.02 $Y2=1.48
r180 29 31 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=2.02 $Y=1.645
+ $X2=2.02 $Y2=2.465
r181 25 86 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.02 $Y=1.315
+ $X2=2.02 $Y2=1.48
r182 25 27 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.02 $Y=1.315
+ $X2=2.02 $Y2=0.655
r183 21 84 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.59 $Y=1.645
+ $X2=1.59 $Y2=1.48
r184 21 23 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=1.59 $Y=1.645
+ $X2=1.59 $Y2=2.465
r185 17 84 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.59 $Y=1.315
+ $X2=1.59 $Y2=1.48
r186 17 19 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.59 $Y=1.315
+ $X2=1.59 $Y2=0.655
r187 13 83 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.16 $Y=1.645
+ $X2=1.16 $Y2=1.48
r188 13 15 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=1.16 $Y=1.645
+ $X2=1.16 $Y2=2.465
r189 9 83 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.16 $Y=1.315
+ $X2=1.16 $Y2=1.48
r190 9 11 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.16 $Y=1.315
+ $X2=1.16 $Y2=0.655
r191 5 82 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.73 $Y=1.645
+ $X2=0.73 $Y2=1.48
r192 5 7 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=0.73 $Y=1.645
+ $X2=0.73 $Y2=2.465
r193 1 82 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.73 $Y=1.315
+ $X2=0.73 $Y2=1.48
r194 1 3 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.73 $Y=1.315
+ $X2=0.73 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__INV_8%VPWR 1 2 3 4 5 18 24 28 32 38 42 44 49 50 51
+ 52 53 62 67 73 76 80
r63 79 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r64 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r65 71 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r66 71 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=3.12 $Y2=3.33
r67 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r68 68 76 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.225 $Y=3.33
+ $X2=3.095 $Y2=3.33
r69 68 70 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=3.225 $Y=3.33
+ $X2=3.6 $Y2=3.33
r70 67 79 4.27534 $w=1.7e-07 $l=2.47e-07 $layer=LI1_cond $X=3.825 $Y=3.33
+ $X2=4.072 $Y2=3.33
r71 67 70 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=3.825 $Y=3.33
+ $X2=3.6 $Y2=3.33
r72 66 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r73 65 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r74 63 73 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.365 $Y=3.33
+ $X2=2.235 $Y2=3.33
r75 63 65 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=2.365 $Y=3.33
+ $X2=2.64 $Y2=3.33
r76 62 76 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.965 $Y=3.33
+ $X2=3.095 $Y2=3.33
r77 62 65 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=2.965 $Y=3.33
+ $X2=2.64 $Y2=3.33
r78 60 61 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r79 57 61 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.2 $Y2=3.33
r80 56 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r81 53 66 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r82 53 61 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.2 $Y2=3.33
r83 53 73 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r84 51 60 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=1.245 $Y=3.33
+ $X2=1.2 $Y2=3.33
r85 51 52 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.245 $Y=3.33
+ $X2=1.375 $Y2=3.33
r86 49 56 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=0.35 $Y=3.33
+ $X2=0.24 $Y2=3.33
r87 49 50 7.94884 $w=1.7e-07 $l=1.47e-07 $layer=LI1_cond $X=0.35 $Y=3.33
+ $X2=0.497 $Y2=3.33
r88 48 60 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=0.645 $Y=3.33
+ $X2=1.2 $Y2=3.33
r89 48 50 7.94884 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=0.645 $Y=3.33
+ $X2=0.497 $Y2=3.33
r90 44 47 26.5648 $w=2.93e-07 $l=6.8e-07 $layer=LI1_cond $X=3.972 $Y=2.26
+ $X2=3.972 $Y2=2.94
r91 42 79 3.20218 $w=2.95e-07 $l=1.36015e-07 $layer=LI1_cond $X=3.972 $Y=3.245
+ $X2=4.072 $Y2=3.33
r92 42 47 11.9151 $w=2.93e-07 $l=3.05e-07 $layer=LI1_cond $X=3.972 $Y=3.245
+ $X2=3.972 $Y2=2.94
r93 38 41 30.1408 $w=2.58e-07 $l=6.8e-07 $layer=LI1_cond $X=3.095 $Y=2.26
+ $X2=3.095 $Y2=2.94
r94 36 76 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=3.095 $Y=3.245
+ $X2=3.095 $Y2=3.33
r95 36 41 13.519 $w=2.58e-07 $l=3.05e-07 $layer=LI1_cond $X=3.095 $Y=3.245
+ $X2=3.095 $Y2=2.94
r96 32 35 30.1408 $w=2.58e-07 $l=6.8e-07 $layer=LI1_cond $X=2.235 $Y=2.26
+ $X2=2.235 $Y2=2.94
r97 30 73 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=2.235 $Y=3.245
+ $X2=2.235 $Y2=3.33
r98 30 35 13.519 $w=2.58e-07 $l=3.05e-07 $layer=LI1_cond $X=2.235 $Y=3.245
+ $X2=2.235 $Y2=2.94
r99 29 52 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.505 $Y=3.33
+ $X2=1.375 $Y2=3.33
r100 28 73 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.105 $Y=3.33
+ $X2=2.235 $Y2=3.33
r101 28 29 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=2.105 $Y=3.33
+ $X2=1.505 $Y2=3.33
r102 24 27 30.1408 $w=2.58e-07 $l=6.8e-07 $layer=LI1_cond $X=1.375 $Y=2.26
+ $X2=1.375 $Y2=2.94
r103 22 52 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=1.375 $Y=3.245
+ $X2=1.375 $Y2=3.33
r104 22 27 13.519 $w=2.58e-07 $l=3.05e-07 $layer=LI1_cond $X=1.375 $Y=3.245
+ $X2=1.375 $Y2=2.94
r105 18 21 26.5648 $w=2.93e-07 $l=6.8e-07 $layer=LI1_cond $X=0.497 $Y=2.27
+ $X2=0.497 $Y2=2.95
r106 16 50 0.543863 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=0.497 $Y=3.245
+ $X2=0.497 $Y2=3.33
r107 16 21 11.5244 $w=2.93e-07 $l=2.95e-07 $layer=LI1_cond $X=0.497 $Y=3.245
+ $X2=0.497 $Y2=2.95
r108 5 47 400 $w=1.7e-07 $l=1.17291e-06 $layer=licon1_PDIFF $count=1 $X=3.815
+ $Y=1.835 $X2=3.955 $Y2=2.94
r109 5 44 400 $w=1.7e-07 $l=4.90026e-07 $layer=licon1_PDIFF $count=1 $X=3.815
+ $Y=1.835 $X2=3.955 $Y2=2.26
r110 4 41 400 $w=1.7e-07 $l=1.17291e-06 $layer=licon1_PDIFF $count=1 $X=2.955
+ $Y=1.835 $X2=3.095 $Y2=2.94
r111 4 38 400 $w=1.7e-07 $l=4.90026e-07 $layer=licon1_PDIFF $count=1 $X=2.955
+ $Y=1.835 $X2=3.095 $Y2=2.26
r112 3 35 400 $w=1.7e-07 $l=1.17291e-06 $layer=licon1_PDIFF $count=1 $X=2.095
+ $Y=1.835 $X2=2.235 $Y2=2.94
r113 3 32 400 $w=1.7e-07 $l=4.90026e-07 $layer=licon1_PDIFF $count=1 $X=2.095
+ $Y=1.835 $X2=2.235 $Y2=2.26
r114 2 27 400 $w=1.7e-07 $l=1.17291e-06 $layer=licon1_PDIFF $count=1 $X=1.235
+ $Y=1.835 $X2=1.375 $Y2=2.94
r115 2 24 400 $w=1.7e-07 $l=4.90026e-07 $layer=licon1_PDIFF $count=1 $X=1.235
+ $Y=1.835 $X2=1.375 $Y2=2.26
r116 1 21 400 $w=1.7e-07 $l=1.18528e-06 $layer=licon1_PDIFF $count=1 $X=0.37
+ $Y=1.835 $X2=0.515 $Y2=2.95
r117 1 18 400 $w=1.7e-07 $l=5.02295e-07 $layer=licon1_PDIFF $count=1 $X=0.37
+ $Y=1.835 $X2=0.515 $Y2=2.27
.ends

.subckt PM_SKY130_FD_SC_LP__INV_8%Y 1 2 3 4 5 6 7 8 26 27 28 29 30 33 37 41 43
+ 47 51 55 57 61 65 69 71 75 79 83 85 87 88 89 91 92 95 96 97 99 100 104 106
r137 104 106 3.84148 $w=2.38e-07 $l=8e-08 $layer=LI1_cond $X=4.105 $Y=1.215
+ $X2=4.105 $Y2=1.295
r138 99 104 2.93484 $w=2.4e-07 $l=8.5e-08 $layer=LI1_cond $X=4.105 $Y=1.13
+ $X2=4.105 $Y2=1.215
r139 99 100 17.6708 $w=2.38e-07 $l=3.68e-07 $layer=LI1_cond $X=4.105 $Y=1.297
+ $X2=4.105 $Y2=1.665
r140 99 106 0.0960369 $w=2.38e-07 $l=2e-09 $layer=LI1_cond $X=4.105 $Y=1.297
+ $X2=4.105 $Y2=1.295
r141 98 100 4.32166 $w=2.38e-07 $l=9e-08 $layer=LI1_cond $X=4.105 $Y=1.755
+ $X2=4.105 $Y2=1.665
r142 92 93 9.97306 $w=2.58e-07 $l=2.25e-07 $layer=LI1_cond $X=2.665 $Y=0.905
+ $X2=2.665 $Y2=1.13
r143 89 90 11.7308 $w=2.34e-07 $l=2.25e-07 $layer=LI1_cond $X=1.805 $Y=0.905
+ $X2=1.805 $Y2=1.13
r144 86 97 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.655 $Y=1.84
+ $X2=3.525 $Y2=1.84
r145 85 98 7.07814 $w=1.7e-07 $l=1.56844e-07 $layer=LI1_cond $X=3.985 $Y=1.84
+ $X2=4.105 $Y2=1.755
r146 85 86 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=3.985 $Y=1.84
+ $X2=3.655 $Y2=1.84
r147 84 96 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.655 $Y=1.13
+ $X2=3.525 $Y2=1.13
r148 83 99 4.1433 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=3.985 $Y=1.13
+ $X2=4.105 $Y2=1.13
r149 83 84 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=3.985 $Y=1.13
+ $X2=3.655 $Y2=1.13
r150 79 81 35.0165 $w=2.58e-07 $l=7.9e-07 $layer=LI1_cond $X=3.525 $Y=2.07
+ $X2=3.525 $Y2=2.86
r151 77 97 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=3.525 $Y=1.925
+ $X2=3.525 $Y2=1.84
r152 77 79 6.42709 $w=2.58e-07 $l=1.45e-07 $layer=LI1_cond $X=3.525 $Y=1.925
+ $X2=3.525 $Y2=2.07
r153 73 96 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=3.525 $Y=1.045
+ $X2=3.525 $Y2=1.13
r154 73 75 25.7083 $w=2.58e-07 $l=5.8e-07 $layer=LI1_cond $X=3.525 $Y=1.045
+ $X2=3.525 $Y2=0.465
r155 72 95 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.795 $Y=1.84
+ $X2=2.665 $Y2=1.84
r156 71 97 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.395 $Y=1.84
+ $X2=3.525 $Y2=1.84
r157 71 72 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=3.395 $Y=1.84
+ $X2=2.795 $Y2=1.84
r158 70 93 3.22376 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.795 $Y=1.13
+ $X2=2.665 $Y2=1.13
r159 69 96 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.395 $Y=1.13
+ $X2=3.525 $Y2=1.13
r160 69 70 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=3.395 $Y=1.13
+ $X2=2.795 $Y2=1.13
r161 65 67 35.0165 $w=2.58e-07 $l=7.9e-07 $layer=LI1_cond $X=2.665 $Y=2.07
+ $X2=2.665 $Y2=2.86
r162 63 95 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=2.665 $Y=1.925
+ $X2=2.665 $Y2=1.84
r163 63 65 6.42709 $w=2.58e-07 $l=1.45e-07 $layer=LI1_cond $X=2.665 $Y=1.925
+ $X2=2.665 $Y2=2.07
r164 59 92 3.7676 $w=2.58e-07 $l=8.5e-08 $layer=LI1_cond $X=2.665 $Y=0.82
+ $X2=2.665 $Y2=0.905
r165 59 61 15.7353 $w=2.58e-07 $l=3.55e-07 $layer=LI1_cond $X=2.665 $Y=0.82
+ $X2=2.665 $Y2=0.465
r166 58 91 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.935 $Y=1.84
+ $X2=1.805 $Y2=1.84
r167 57 95 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.535 $Y=1.84
+ $X2=2.665 $Y2=1.84
r168 57 58 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=2.535 $Y=1.84
+ $X2=1.935 $Y2=1.84
r169 56 89 2.60974 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.935 $Y=0.905
+ $X2=1.805 $Y2=0.905
r170 55 92 3.22376 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.535 $Y=0.905
+ $X2=2.665 $Y2=0.905
r171 55 56 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=2.535 $Y=0.905
+ $X2=1.935 $Y2=0.905
r172 51 53 35.0165 $w=2.58e-07 $l=7.9e-07 $layer=LI1_cond $X=1.805 $Y=2.07
+ $X2=1.805 $Y2=2.86
r173 49 91 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=1.805 $Y=1.925
+ $X2=1.805 $Y2=1.84
r174 49 51 6.42709 $w=2.58e-07 $l=1.45e-07 $layer=LI1_cond $X=1.805 $Y=1.925
+ $X2=1.805 $Y2=2.07
r175 45 89 4.13705 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=1.805 $Y=0.82
+ $X2=1.805 $Y2=0.905
r176 45 47 15.7353 $w=2.58e-07 $l=3.55e-07 $layer=LI1_cond $X=1.805 $Y=0.82
+ $X2=1.805 $Y2=0.465
r177 44 88 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.075 $Y=1.84
+ $X2=0.945 $Y2=1.84
r178 43 91 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.675 $Y=1.84
+ $X2=1.805 $Y2=1.84
r179 43 44 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=1.675 $Y=1.84
+ $X2=1.075 $Y2=1.84
r180 42 87 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.075 $Y=1.13
+ $X2=0.945 $Y2=1.13
r181 41 90 2.60974 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.675 $Y=1.13
+ $X2=1.805 $Y2=1.13
r182 41 42 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=1.675 $Y=1.13
+ $X2=1.075 $Y2=1.13
r183 37 39 35.0165 $w=2.58e-07 $l=7.9e-07 $layer=LI1_cond $X=0.945 $Y=2.07
+ $X2=0.945 $Y2=2.86
r184 35 88 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=0.945 $Y=1.925
+ $X2=0.945 $Y2=1.84
r185 35 37 6.42709 $w=2.58e-07 $l=1.45e-07 $layer=LI1_cond $X=0.945 $Y=1.925
+ $X2=0.945 $Y2=2.07
r186 31 87 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=0.945 $Y=1.045
+ $X2=0.945 $Y2=1.13
r187 31 33 25.7083 $w=2.58e-07 $l=5.8e-07 $layer=LI1_cond $X=0.945 $Y=1.045
+ $X2=0.945 $Y2=0.465
r188 29 88 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.815 $Y=1.84
+ $X2=0.945 $Y2=1.84
r189 29 30 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=0.815 $Y=1.84
+ $X2=0.255 $Y2=1.84
r190 27 87 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.815 $Y=1.13
+ $X2=0.945 $Y2=1.13
r191 27 28 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=0.815 $Y=1.13
+ $X2=0.255 $Y2=1.13
r192 26 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.17 $Y=1.755
+ $X2=0.255 $Y2=1.84
r193 25 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.17 $Y=1.215
+ $X2=0.255 $Y2=1.13
r194 25 26 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=0.17 $Y=1.215
+ $X2=0.17 $Y2=1.755
r195 8 81 400 $w=1.7e-07 $l=1.09276e-06 $layer=licon1_PDIFF $count=1 $X=3.385
+ $Y=1.835 $X2=3.525 $Y2=2.86
r196 8 79 400 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_PDIFF $count=1 $X=3.385
+ $Y=1.835 $X2=3.525 $Y2=2.07
r197 7 67 400 $w=1.7e-07 $l=1.09276e-06 $layer=licon1_PDIFF $count=1 $X=2.525
+ $Y=1.835 $X2=2.665 $Y2=2.86
r198 7 65 400 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_PDIFF $count=1 $X=2.525
+ $Y=1.835 $X2=2.665 $Y2=2.07
r199 6 53 400 $w=1.7e-07 $l=1.09276e-06 $layer=licon1_PDIFF $count=1 $X=1.665
+ $Y=1.835 $X2=1.805 $Y2=2.86
r200 6 51 400 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_PDIFF $count=1 $X=1.665
+ $Y=1.835 $X2=1.805 $Y2=2.07
r201 5 39 400 $w=1.7e-07 $l=1.09276e-06 $layer=licon1_PDIFF $count=1 $X=0.805
+ $Y=1.835 $X2=0.945 $Y2=2.86
r202 5 37 400 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_PDIFF $count=1 $X=0.805
+ $Y=1.835 $X2=0.945 $Y2=2.07
r203 4 75 91 $w=1.7e-07 $l=2.91719e-07 $layer=licon1_NDIFF $count=2 $X=3.385
+ $Y=0.235 $X2=3.525 $Y2=0.465
r204 3 61 91 $w=1.7e-07 $l=2.91719e-07 $layer=licon1_NDIFF $count=2 $X=2.525
+ $Y=0.235 $X2=2.665 $Y2=0.465
r205 2 47 91 $w=1.7e-07 $l=2.91719e-07 $layer=licon1_NDIFF $count=2 $X=1.665
+ $Y=0.235 $X2=1.805 $Y2=0.465
r206 1 33 91 $w=1.7e-07 $l=2.91719e-07 $layer=licon1_NDIFF $count=2 $X=0.805
+ $Y=0.235 $X2=0.945 $Y2=0.465
.ends

.subckt PM_SKY130_FD_SC_LP__INV_8%VGND 1 2 3 4 5 18 22 24 28 32 34 36 39 40 41
+ 42 43 52 57 63 66 70
r65 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r66 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r67 61 70 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r68 61 67 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=3.12
+ $Y2=0
r69 60 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r70 58 66 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.225 $Y=0 $X2=3.095
+ $Y2=0
r71 58 60 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=3.225 $Y=0 $X2=3.6
+ $Y2=0
r72 57 69 4.27534 $w=1.7e-07 $l=2.47e-07 $layer=LI1_cond $X=3.825 $Y=0 $X2=4.072
+ $Y2=0
r73 57 60 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=3.825 $Y=0 $X2=3.6
+ $Y2=0
r74 56 67 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r75 55 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r76 53 63 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.365 $Y=0 $X2=2.235
+ $Y2=0
r77 53 55 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=2.365 $Y=0 $X2=2.64
+ $Y2=0
r78 52 66 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.965 $Y=0 $X2=3.095
+ $Y2=0
r79 52 55 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=2.965 $Y=0 $X2=2.64
+ $Y2=0
r80 50 51 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r81 47 51 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r82 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r83 43 56 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r84 43 51 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.2
+ $Y2=0
r85 43 63 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r86 41 50 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=1.245 $Y=0 $X2=1.2
+ $Y2=0
r87 41 42 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.245 $Y=0 $X2=1.375
+ $Y2=0
r88 39 46 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=0.35 $Y=0 $X2=0.24
+ $Y2=0
r89 39 40 7.94884 $w=1.7e-07 $l=1.47e-07 $layer=LI1_cond $X=0.35 $Y=0 $X2=0.497
+ $Y2=0
r90 38 50 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=0.645 $Y=0 $X2=1.2
+ $Y2=0
r91 38 40 7.94884 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=0.645 $Y=0 $X2=0.497
+ $Y2=0
r92 34 69 3.20218 $w=2.95e-07 $l=1.36015e-07 $layer=LI1_cond $X=3.972 $Y=0.085
+ $X2=4.072 $Y2=0
r93 34 36 11.1338 $w=2.93e-07 $l=2.85e-07 $layer=LI1_cond $X=3.972 $Y=0.085
+ $X2=3.972 $Y2=0.37
r94 30 66 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=3.095 $Y=0.085
+ $X2=3.095 $Y2=0
r95 30 32 12.6325 $w=2.58e-07 $l=2.85e-07 $layer=LI1_cond $X=3.095 $Y=0.085
+ $X2=3.095 $Y2=0.37
r96 26 63 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=2.235 $Y=0.085
+ $X2=2.235 $Y2=0
r97 26 28 17.7299 $w=2.58e-07 $l=4e-07 $layer=LI1_cond $X=2.235 $Y=0.085
+ $X2=2.235 $Y2=0.485
r98 25 42 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.505 $Y=0 $X2=1.375
+ $Y2=0
r99 24 63 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.105 $Y=0 $X2=2.235
+ $Y2=0
r100 24 25 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=2.105 $Y=0 $X2=1.505
+ $Y2=0
r101 20 42 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=1.375 $Y=0.085
+ $X2=1.375 $Y2=0
r102 20 22 12.6325 $w=2.58e-07 $l=2.85e-07 $layer=LI1_cond $X=1.375 $Y=0.085
+ $X2=1.375 $Y2=0.37
r103 16 40 0.543863 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=0.497 $Y=0.085
+ $X2=0.497 $Y2=0
r104 16 18 11.1338 $w=2.93e-07 $l=2.85e-07 $layer=LI1_cond $X=0.497 $Y=0.085
+ $X2=0.497 $Y2=0.37
r105 5 36 91 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_NDIFF $count=2 $X=3.815
+ $Y=0.235 $X2=3.955 $Y2=0.37
r106 4 32 91 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_NDIFF $count=2 $X=2.955
+ $Y=0.235 $X2=3.095 $Y2=0.37
r107 3 28 182 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=1 $X=2.095
+ $Y=0.235 $X2=2.235 $Y2=0.485
r108 2 22 91 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_NDIFF $count=2 $X=1.235
+ $Y=0.235 $X2=1.375 $Y2=0.37
r109 1 18 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=0.37
+ $Y=0.235 $X2=0.515 $Y2=0.37
.ends

