* NGSPICE file created from sky130_fd_sc_lp__o32a_4.ext - technology: sky130A

.subckt sky130_fd_sc_lp__o32a_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
M1000 X a_547_367# VGND VNB nshort w=840000u l=150000u
+  ad=4.704e+11p pd=4.48e+06u as=1.6884e+12p ps=1.41e+07u
M1001 a_823_367# B1 VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=7.119e+11p pd=6.17e+06u as=1.7262e+12p ps=1.534e+07u
M1002 VPWR A1 a_195_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=7.56e+11p ps=6.24e+06u
M1003 a_44_65# B2 a_547_367# VNB nshort w=840000u l=150000u
+  ad=1.848e+12p pd=1.448e+07u as=5.334e+11p ps=4.63e+06u
M1004 VPWR a_547_367# X VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=7.056e+11p ps=6.16e+06u
M1005 a_547_367# A3 a_112_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=1.0206e+12p pd=9.18e+06u as=1.0206e+12p ps=9.18e+06u
M1006 VGND A1 a_44_65# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND a_547_367# X VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_547_367# B1 a_44_65# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND a_547_367# X VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR B1 a_823_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 X a_547_367# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VGND A2 a_44_65# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_195_367# A2 a_112_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_547_367# B2 a_823_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_112_367# A2 a_195_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 X a_547_367# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VGND A3 a_44_65# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_44_65# A2 VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_44_65# A1 VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 X a_547_367# VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_44_65# B1 a_547_367# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_44_65# A3 VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_547_367# B2 a_44_65# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_195_367# A1 VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_112_367# A3 a_547_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_823_367# B2 a_547_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 VPWR a_547_367# X VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

