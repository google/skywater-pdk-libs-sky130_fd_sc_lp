* NGSPICE file created from sky130_fd_sc_lp__nand2_1.ext - technology: sky130A

.subckt sky130_fd_sc_lp__nand2_1 A B VGND VNB VPB VPWR Y
M1000 a_112_69# B VGND VNB nshort w=840000u l=150000u
+  ad=2.016e+11p pd=2.16e+06u as=2.226e+11p ps=2.21e+06u
M1001 VPWR A Y VPB phighvt w=1.26e+06u l=150000u
+  ad=6.678e+11p pd=6.1e+06u as=3.528e+11p ps=3.08e+06u
M1002 Y A a_112_69# VNB nshort w=840000u l=150000u
+  ad=2.226e+11p pd=2.21e+06u as=0p ps=0u
M1003 Y B VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

