* File: sky130_fd_sc_lp__and4b_lp.pex.spice
* Created: Wed Sep  2 09:33:47 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__AND4B_LP%A_84_21# 1 2 3 10 12 17 19 21 23 24 26 27
+ 28 31 32 34 35 38 42 46 51 52 53 55
c115 51 0 1.28945e-19 $X=2.61 $Y=1.97
r116 55 57 9.16063 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=2.69 $Y=0.445
+ $X2=2.69 $Y2=0.63
r117 51 53 3.351 $w=2.8e-07 $l=1.46458e-07 $layer=LI1_cond $X=2.61 $Y=1.97
+ $X2=2.5 $Y2=2.055
r118 51 57 87.4225 $w=1.68e-07 $l=1.34e-06 $layer=LI1_cond $X=2.61 $Y=1.97
+ $X2=2.61 $Y2=0.63
r119 46 48 20.9804 $w=3.88e-07 $l=7.1e-07 $layer=LI1_cond $X=2.5 $Y=2.19 $X2=2.5
+ $Y2=2.9
r120 44 53 3.351 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.5 $Y=2.14 $X2=2.5
+ $Y2=2.055
r121 44 46 1.47749 $w=3.88e-07 $l=5e-08 $layer=LI1_cond $X=2.5 $Y=2.14 $X2=2.5
+ $Y2=2.19
r122 43 52 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.555 $Y=2.055
+ $X2=1.39 $Y2=2.055
r123 42 53 3.18746 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=2.305 $Y=2.055
+ $X2=2.5 $Y2=2.055
r124 42 43 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=2.305 $Y=2.055
+ $X2=1.555 $Y2=2.055
r125 38 40 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=1.39 $Y=2.19
+ $X2=1.39 $Y2=2.9
r126 36 52 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.39 $Y=2.14
+ $X2=1.39 $Y2=2.055
r127 36 38 1.74613 $w=3.28e-07 $l=5e-08 $layer=LI1_cond $X=1.39 $Y=2.14 $X2=1.39
+ $Y2=2.19
r128 34 52 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.225 $Y=2.055
+ $X2=1.39 $Y2=2.055
r129 34 35 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=1.225 $Y=2.055
+ $X2=0.75 $Y2=2.055
r130 31 32 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.585
+ $Y=1.33 $X2=0.585 $Y2=1.33
r131 29 35 7.59919 $w=1.7e-07 $l=1.92873e-07 $layer=LI1_cond $X=0.595 $Y=1.97
+ $X2=0.75 $Y2=2.055
r132 29 31 23.7924 $w=3.08e-07 $l=6.4e-07 $layer=LI1_cond $X=0.595 $Y=1.97
+ $X2=0.595 $Y2=1.33
r133 27 32 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.585 $Y=1.67
+ $X2=0.585 $Y2=1.33
r134 27 28 30.8683 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.585 $Y=1.67
+ $X2=0.585 $Y2=1.835
r135 26 32 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.585 $Y=1.165
+ $X2=0.585 $Y2=1.33
r136 21 23 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.855 $Y=0.73
+ $X2=0.855 $Y2=0.445
r137 20 24 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.57 $Y=0.805
+ $X2=0.495 $Y2=0.805
r138 19 21 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.78 $Y=0.805
+ $X2=0.855 $Y2=0.73
r139 19 20 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=0.78 $Y=0.805
+ $X2=0.57 $Y2=0.805
r140 17 28 176.402 $w=2.5e-07 $l=7.1e-07 $layer=POLY_cond $X=0.595 $Y=2.545
+ $X2=0.595 $Y2=1.835
r141 13 24 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.495 $Y=0.88
+ $X2=0.495 $Y2=0.805
r142 13 26 146.138 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.495 $Y=0.88
+ $X2=0.495 $Y2=1.165
r143 10 24 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.495 $Y=0.73
+ $X2=0.495 $Y2=0.805
r144 10 12 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.495 $Y=0.73
+ $X2=0.495 $Y2=0.445
r145 3 48 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=2.33
+ $Y=2.045 $X2=2.47 $Y2=2.9
r146 3 46 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.33
+ $Y=2.045 $X2=2.47 $Y2=2.19
r147 2 40 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=1.25
+ $Y=2.045 $X2=1.39 $Y2=2.9
r148 2 38 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.25
+ $Y=2.045 $X2=1.39 $Y2=2.19
r149 1 55 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.55
+ $Y=0.235 $X2=2.69 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__AND4B_LP%D 1 3 7 9 11 12 15 17 18 22
r53 17 18 12.336 $w=3.53e-07 $l=3.8e-07 $layer=LI1_cond $X=1.137 $Y=1.285
+ $X2=1.137 $Y2=1.665
r54 17 22 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.125
+ $Y=1.285 $X2=1.125 $Y2=1.285
r55 13 15 46.1489 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=1.215 $Y=0.805
+ $X2=1.305 $Y2=0.805
r56 12 22 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.125 $Y=1.625
+ $X2=1.125 $Y2=1.285
r57 11 22 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.125 $Y=1.12
+ $X2=1.125 $Y2=1.285
r58 7 15 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.305 $Y=0.73
+ $X2=1.305 $Y2=0.805
r59 7 9 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=1.305 $Y=0.73 $X2=1.305
+ $Y2=0.445
r60 5 13 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.215 $Y=0.88
+ $X2=1.215 $Y2=0.805
r61 5 11 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=1.215 $Y=0.88
+ $X2=1.215 $Y2=1.12
r62 1 12 30.6163 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.125 $Y=1.79
+ $X2=1.125 $Y2=1.625
r63 1 3 187.582 $w=2.5e-07 $l=7.55e-07 $layer=POLY_cond $X=1.125 $Y=1.79
+ $X2=1.125 $Y2=2.545
.ends

.subckt PM_SKY130_FD_SC_LP__AND4B_LP%C 3 7 11 12 13 14 15 16 22
r51 15 16 13.2706 $w=3.28e-07 $l=3.8e-07 $layer=LI1_cond $X=1.665 $Y=1.285
+ $X2=1.665 $Y2=1.665
r52 15 22 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.665
+ $Y=1.285 $X2=1.665 $Y2=1.285
r53 14 15 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=1.665 $Y=0.925
+ $X2=1.665 $Y2=1.285
r54 13 14 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.665 $Y=0.555
+ $X2=1.665 $Y2=0.925
r55 11 22 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.665 $Y=1.625
+ $X2=1.665 $Y2=1.285
r56 11 12 30.8683 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.665 $Y=1.625
+ $X2=1.665 $Y2=1.79
r57 10 22 39.2677 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.665 $Y=1.12
+ $X2=1.665 $Y2=1.285
r58 7 10 346.117 $w=1.5e-07 $l=6.75e-07 $layer=POLY_cond $X=1.695 $Y=0.445
+ $X2=1.695 $Y2=1.12
r59 3 12 187.582 $w=2.5e-07 $l=7.55e-07 $layer=POLY_cond $X=1.655 $Y=2.545
+ $X2=1.655 $Y2=1.79
.ends

.subckt PM_SKY130_FD_SC_LP__AND4B_LP%B 3 6 8 10 11 13 14 15 16 17 18 24
c51 15 0 9.91956e-20 $X=2.16 $Y=0.555
c52 11 0 2.02481e-19 $X=2.1 $Y=0.88
r53 17 18 14.3583 $w=3.03e-07 $l=3.8e-07 $layer=LI1_cond $X=2.192 $Y=1.285
+ $X2=2.192 $Y2=1.665
r54 17 24 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.205
+ $Y=1.285 $X2=2.205 $Y2=1.285
r55 16 17 13.6026 $w=3.03e-07 $l=3.6e-07 $layer=LI1_cond $X=2.192 $Y=0.925
+ $X2=2.192 $Y2=1.285
r56 15 16 13.9805 $w=3.03e-07 $l=3.7e-07 $layer=LI1_cond $X=2.192 $Y=0.555
+ $X2=2.192 $Y2=0.925
r57 14 24 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.205 $Y=1.625
+ $X2=2.205 $Y2=1.285
r58 13 24 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.205 $Y=1.12
+ $X2=2.205 $Y2=1.285
r59 11 13 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=2.115 $Y=0.88
+ $X2=2.115 $Y2=1.12
r60 10 11 58.3064 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=2.1 $Y=0.73 $X2=2.1
+ $Y2=0.88
r61 6 14 30.6163 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.205 $Y=1.79
+ $X2=2.205 $Y2=1.625
r62 6 8 187.582 $w=2.5e-07 $l=7.55e-07 $layer=POLY_cond $X=2.205 $Y=1.79
+ $X2=2.205 $Y2=2.545
r63 3 10 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.085 $Y=0.445
+ $X2=2.085 $Y2=0.73
.ends

.subckt PM_SKY130_FD_SC_LP__AND4B_LP%A_480_21# 1 2 7 9 10 11 12 14 17 18 23 25
+ 30 34
c70 12 0 9.91956e-20 $X=2.735 $Y=1.82
r71 34 36 9.85908 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=4.04 $Y=0.47
+ $X2=4.04 $Y2=0.675
r72 30 32 3.3128 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.12 $Y=1.365
+ $X2=4.12 $Y2=1.53
r73 30 36 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=4.12 $Y=1.365
+ $X2=4.12 $Y2=0.675
r74 25 27 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=3.81 $Y=2.19 $X2=3.81
+ $Y2=2.9
r75 23 32 14.3258 $w=2.64e-07 $l=3.1e-07 $layer=LI1_cond $X=3.81 $Y=1.53
+ $X2=4.12 $Y2=1.53
r76 23 25 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=3.81 $Y=1.695
+ $X2=3.81 $Y2=2.19
r77 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.015
+ $Y=1.53 $X2=3.015 $Y2=1.53
r78 18 23 6.62312 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=3.645 $Y=1.53
+ $X2=3.81 $Y2=1.53
r79 18 20 22.0012 $w=3.28e-07 $l=6.3e-07 $layer=LI1_cond $X=3.645 $Y=1.53
+ $X2=3.015 $Y2=1.53
r80 17 21 8.61411 $w=4.7e-07 $l=9.16515e-08 $layer=POLY_cond $X=2.945 $Y=1.46
+ $X2=2.895 $Y2=1.53
r81 16 17 68.6318 $w=4.7e-07 $l=5.8e-07 $layer=POLY_cond $X=2.945 $Y=0.88
+ $X2=2.945 $Y2=1.46
r82 12 21 41.9244 $w=3.93e-07 $l=3.61248e-07 $layer=POLY_cond $X=2.735 $Y=1.82
+ $X2=2.895 $Y2=1.53
r83 12 14 180.129 $w=2.5e-07 $l=7.25e-07 $layer=POLY_cond $X=2.735 $Y=1.82
+ $X2=2.735 $Y2=2.545
r84 10 16 37.5433 $w=1.5e-07 $l=2.69907e-07 $layer=POLY_cond $X=2.71 $Y=0.805
+ $X2=2.945 $Y2=0.88
r85 10 11 82.0426 $w=1.5e-07 $l=1.6e-07 $layer=POLY_cond $X=2.71 $Y=0.805
+ $X2=2.55 $Y2=0.805
r86 7 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.475 $Y=0.73
+ $X2=2.55 $Y2=0.805
r87 7 9 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.475 $Y=0.73 $X2=2.475
+ $Y2=0.445
r88 2 27 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=3.67
+ $Y=2.045 $X2=3.81 $Y2=2.9
r89 2 25 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=3.67
+ $Y=2.045 $X2=3.81 $Y2=2.19
r90 1 34 182 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=1 $X=3.9
+ $Y=0.235 $X2=4.04 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_LP__AND4B_LP%A_N 3 7 11 15 18 24 29
c42 24 0 1.01448e-20 $X=3.825 $Y=1.02
r43 20 22 13.9889 $w=3.3e-07 $l=8e-08 $layer=POLY_cond $X=3.465 $Y=1.02
+ $X2=3.545 $Y2=1.02
r44 18 29 3.72928 $w=3.73e-07 $l=1.15e-07 $layer=LI1_cond $X=3.12 $Y=0.997
+ $X2=3.235 $Y2=0.997
r45 16 24 24.4806 $w=3.3e-07 $l=1.4e-07 $layer=POLY_cond $X=3.685 $Y=1.02
+ $X2=3.825 $Y2=1.02
r46 16 22 24.4806 $w=3.3e-07 $l=1.4e-07 $layer=POLY_cond $X=3.685 $Y=1.02
+ $X2=3.545 $Y2=1.02
r47 15 29 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=3.685 $Y=1.02
+ $X2=3.235 $Y2=1.02
r48 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.685
+ $Y=1.02 $X2=3.685 $Y2=1.02
r49 9 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.825 $Y=0.855
+ $X2=3.825 $Y2=1.02
r50 9 11 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=3.825 $Y=0.855
+ $X2=3.825 $Y2=0.445
r51 5 22 9.34494 $w=2.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.545 $Y=1.185
+ $X2=3.545 $Y2=1.02
r52 5 7 337.897 $w=2.5e-07 $l=1.36e-06 $layer=POLY_cond $X=3.545 $Y=1.185
+ $X2=3.545 $Y2=2.545
r53 1 20 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.465 $Y=0.855
+ $X2=3.465 $Y2=1.02
r54 1 3 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=3.465 $Y=0.855
+ $X2=3.465 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__AND4B_LP%X 1 2 12 13 14
r20 14 16 1.82704 $w=4.08e-07 $l=6.5e-08 $layer=LI1_cond $X=0.24 $Y=0.47
+ $X2=0.175 $Y2=0.47
r21 12 13 8.6688 $w=4.03e-07 $l=1.65e-07 $layer=LI1_cond $X=0.292 $Y=2.485
+ $X2=0.292 $Y2=2.32
r22 7 16 5.92876 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=0.175 $Y=0.675
+ $X2=0.175 $Y2=0.47
r23 7 13 107.321 $w=1.68e-07 $l=1.645e-06 $layer=LI1_cond $X=0.175 $Y=0.675
+ $X2=0.175 $Y2=2.32
r24 2 12 300 $w=1.7e-07 $l=5.07346e-07 $layer=licon1_PDIFF $count=2 $X=0.185
+ $Y=2.045 $X2=0.33 $Y2=2.485
r25 1 14 182 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.28 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_LP__AND4B_LP%VPWR 1 2 3 14 18 22 27 28 29 35 41 42 45 48
r54 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r55 45 46 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r56 42 49 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.12 $Y2=3.33
r57 41 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r58 39 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.205 $Y=3.33
+ $X2=3.04 $Y2=3.33
r59 39 41 57.0856 $w=1.68e-07 $l=8.75e-07 $layer=LI1_cond $X=3.205 $Y=3.33
+ $X2=4.08 $Y2=3.33
r60 38 49 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r61 37 38 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r62 35 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.875 $Y=3.33
+ $X2=3.04 $Y2=3.33
r63 35 37 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=2.875 $Y=3.33
+ $X2=2.64 $Y2=3.33
r64 34 46 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.72 $Y2=3.33
r65 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r66 31 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.025 $Y=3.33
+ $X2=0.86 $Y2=3.33
r67 31 33 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=1.025 $Y=3.33
+ $X2=1.68 $Y2=3.33
r68 29 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r69 29 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r70 27 33 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=1.755 $Y=3.33
+ $X2=1.68 $Y2=3.33
r71 27 28 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.755 $Y=3.33
+ $X2=1.92 $Y2=3.33
r72 26 37 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=2.085 $Y=3.33
+ $X2=2.64 $Y2=3.33
r73 26 28 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.085 $Y=3.33
+ $X2=1.92 $Y2=3.33
r74 22 25 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=3.04 $Y=2.19 $X2=3.04
+ $Y2=2.9
r75 20 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.04 $Y=3.245
+ $X2=3.04 $Y2=3.33
r76 20 25 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=3.04 $Y=3.245
+ $X2=3.04 $Y2=2.9
r77 16 28 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.92 $Y=3.245
+ $X2=1.92 $Y2=3.33
r78 16 18 26.5411 $w=3.28e-07 $l=7.6e-07 $layer=LI1_cond $X=1.92 $Y=3.245
+ $X2=1.92 $Y2=2.485
r79 12 45 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.86 $Y=3.245
+ $X2=0.86 $Y2=3.33
r80 12 14 26.5411 $w=3.28e-07 $l=7.6e-07 $layer=LI1_cond $X=0.86 $Y=3.245
+ $X2=0.86 $Y2=2.485
r81 3 25 400 $w=1.7e-07 $l=9.40705e-07 $layer=licon1_PDIFF $count=1 $X=2.86
+ $Y=2.045 $X2=3.04 $Y2=2.9
r82 3 22 400 $w=1.7e-07 $l=2.41868e-07 $layer=licon1_PDIFF $count=1 $X=2.86
+ $Y=2.045 $X2=3.04 $Y2=2.19
r83 2 18 300 $w=1.7e-07 $l=5.05173e-07 $layer=licon1_PDIFF $count=2 $X=1.78
+ $Y=2.045 $X2=1.92 $Y2=2.485
r84 1 14 300 $w=1.7e-07 $l=5.05173e-07 $layer=licon1_PDIFF $count=2 $X=0.72
+ $Y=2.045 $X2=0.86 $Y2=2.485
.ends

.subckt PM_SKY130_FD_SC_LP__AND4B_LP%VGND 1 2 9 11 15 17 19 26 27 30 33
c66 11 0 8.36808e-20 $X=3.085 $Y=0
r67 33 34 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r68 30 31 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r69 27 34 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.12
+ $Y2=0
r70 26 27 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r71 24 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.415 $Y=0 $X2=3.25
+ $Y2=0
r72 24 26 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=3.415 $Y=0 $X2=4.08
+ $Y2=0
r73 22 31 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r74 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r75 19 30 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.905 $Y=0 $X2=1.07
+ $Y2=0
r76 19 21 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=0.905 $Y=0 $X2=0.72
+ $Y2=0
r77 17 34 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r78 17 31 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.2
+ $Y2=0
r79 13 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.25 $Y=0.085
+ $X2=3.25 $Y2=0
r80 13 15 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=3.25 $Y=0.085
+ $X2=3.25 $Y2=0.42
r81 12 30 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.235 $Y=0 $X2=1.07
+ $Y2=0
r82 11 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.085 $Y=0 $X2=3.25
+ $Y2=0
r83 11 12 120.695 $w=1.68e-07 $l=1.85e-06 $layer=LI1_cond $X=3.085 $Y=0
+ $X2=1.235 $Y2=0
r84 7 30 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.07 $Y=0.085 $X2=1.07
+ $Y2=0
r85 7 9 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=1.07 $Y=0.085 $X2=1.07
+ $Y2=0.445
r86 2 15 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=3.105
+ $Y=0.235 $X2=3.25 $Y2=0.42
r87 1 9 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.93
+ $Y=0.235 $X2=1.07 $Y2=0.445
.ends

