* File: sky130_fd_sc_lp__o311ai_lp.spice
* Created: Wed Sep  2 10:24:06 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__o311ai_lp.pex.spice"
.subckt sky130_fd_sc_lp__o311ai_lp  VNB VPB A1 A2 A3 B1 C1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* C1	C1
* B1	B1
* A3	A3
* A2	A2
* A1	A1
* VPB	VPB
* VNB	VNB
MM1008 N_A_114_148#_M1008_d N_A1_M1008_g N_VGND_M1008_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0651 AS=0.1197 PD=0.73 PS=1.41 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.3 A=0.063 P=1.14 MULT=1
MM1003 N_VGND_M1003_d N_A2_M1003_g N_A_114_148#_M1008_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1029 AS=0.0651 PD=0.91 PS=0.73 NRD=14.28 NRS=8.568 M=1 R=2.8 SA=75000.7
+ SB=75001.8 A=0.063 P=1.14 MULT=1
MM1004 N_A_114_148#_M1004_d N_A3_M1004_g N_VGND_M1003_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0924 AS=0.1029 PD=0.86 PS=0.91 NRD=22.848 NRS=45.708 M=1 R=2.8 SA=75001.3
+ SB=75001.2 A=0.063 P=1.14 MULT=1
MM1007 A_452_148# N_B1_M1007_g N_A_114_148#_M1004_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0924 PD=0.63 PS=0.86 NRD=14.28 NRS=22.848 M=1 R=2.8 SA=75001.9
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1005 N_Y_M1005_d N_C1_M1005_g A_452_148# VNB NSHORT L=0.15 W=0.42 AD=0.1197
+ AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75002.3 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1009 A_134_419# N_A1_M1009_g N_VPWR_M1009_s VPB PHIGHVT L=0.25 W=1 AD=0.12
+ AS=0.285 PD=1.24 PS=2.57 NRD=12.7853 NRS=0 M=1 R=4 SA=125000 SB=125002 A=0.25
+ P=2.5 MULT=1
MM1000 A_232_419# N_A2_M1000_g A_134_419# VPB PHIGHVT L=0.25 W=1 AD=0.13 AS=0.12
+ PD=1.26 PS=1.24 NRD=14.7553 NRS=12.7853 M=1 R=4 SA=125001 SB=125002 A=0.25
+ P=2.5 MULT=1
MM1001 N_Y_M1001_d N_A3_M1001_g A_232_419# VPB PHIGHVT L=0.25 W=1 AD=0.14
+ AS=0.13 PD=1.28 PS=1.26 NRD=0 NRS=14.7553 M=1 R=4 SA=125001 SB=125001 A=0.25
+ P=2.5 MULT=1
MM1006 N_VPWR_M1006_d N_B1_M1006_g N_Y_M1001_d VPB PHIGHVT L=0.25 W=1 AD=0.15
+ AS=0.14 PD=1.3 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125002 SB=125001 A=0.25 P=2.5
+ MULT=1
MM1002 N_Y_M1002_d N_C1_M1002_g N_VPWR_M1006_d VPB PHIGHVT L=0.25 W=1 AD=0.285
+ AS=0.15 PD=2.57 PS=1.3 NRD=0 NRS=3.9203 M=1 R=4 SA=125002 SB=125000 A=0.25
+ P=2.5 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9751 P=11.21
*
.include "sky130_fd_sc_lp__o311ai_lp.pxi.spice"
*
.ends
*
*
