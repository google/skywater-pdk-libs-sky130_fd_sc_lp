* File: sky130_fd_sc_lp__dlxbn_1.pex.spice
* Created: Fri Aug 28 10:27:45 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__DLXBN_1%D 3 7 9 10 11 12 13 17
r35 17 18 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.54
+ $Y=1.37 $X2=0.54 $Y2=1.37
r36 13 18 7.63979 $w=4.43e-07 $l=2.95e-07 $layer=LI1_cond $X=0.677 $Y=1.665
+ $X2=0.677 $Y2=1.37
r37 12 18 1.94232 $w=4.43e-07 $l=7.5e-08 $layer=LI1_cond $X=0.677 $Y=1.295
+ $X2=0.677 $Y2=1.37
r38 10 17 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.54 $Y=1.71
+ $X2=0.54 $Y2=1.37
r39 10 11 39.2677 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.54 $Y=1.71
+ $X2=0.54 $Y2=1.875
r40 9 17 40.8701 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.54 $Y=1.205
+ $X2=0.54 $Y2=1.37
r41 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.59 $Y=0.885 $X2=0.59
+ $Y2=1.205
r42 3 11 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=0.51 $Y=2.355
+ $X2=0.51 $Y2=1.875
.ends

.subckt PM_SKY130_FD_SC_LP__DLXBN_1%GATE_N 1 3 6 8 11 12 13 14 18
c44 18 0 1.95136e-19 $X=1.6 $Y=0.4
r45 18 21 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.6 $Y=0.4 $X2=1.6
+ $Y2=0.565
r46 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.6 $Y=0.4
+ $X2=1.6 $Y2=0.4
r47 14 19 2.19513 $w=4.18e-07 $l=8e-08 $layer=LI1_cond $X=1.68 $Y=0.465 $X2=1.6
+ $Y2=0.465
r48 13 19 10.9756 $w=4.18e-07 $l=4e-07 $layer=LI1_cond $X=1.2 $Y=0.465 $X2=1.6
+ $Y2=0.465
r49 11 21 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=1.51 $Y=1.205
+ $X2=1.51 $Y2=0.565
r50 9 12 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.095 $Y=1.28
+ $X2=1.02 $Y2=1.28
r51 8 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.435 $Y=1.28
+ $X2=1.51 $Y2=1.205
r52 8 9 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=1.435 $Y=1.28 $X2=1.095
+ $Y2=1.28
r53 4 12 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.02 $Y=1.355
+ $X2=1.02 $Y2=1.28
r54 4 6 512.766 $w=1.5e-07 $l=1e-06 $layer=POLY_cond $X=1.02 $Y=1.355 $X2=1.02
+ $Y2=2.355
r55 1 12 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.02 $Y=1.205
+ $X2=1.02 $Y2=1.28
r56 1 3 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.02 $Y=1.205 $X2=1.02
+ $Y2=0.885
.ends

.subckt PM_SKY130_FD_SC_LP__DLXBN_1%A_219_135# 1 2 9 13 17 19 20 23 27 30 33 34
+ 42 43 47 48
c108 47 0 7.24186e-20 $X=3.145 $Y=1.18
c109 43 0 1.65621e-19 $X=2.035 $Y=1.36
c110 34 0 1.55622e-19 $X=2.98 $Y=1.28
r111 47 48 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.145
+ $Y=1.18 $X2=3.145 $Y2=1.18
r112 42 45 6.55482 $w=9.12e-07 $l=4.9e-07 $layer=LI1_cond $X=1.635 $Y=1.36
+ $X2=1.635 $Y2=1.85
r113 42 43 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.035
+ $Y=1.36 $X2=2.035 $Y2=1.36
r114 40 42 1.07018 $w=9.12e-07 $l=8e-08 $layer=LI1_cond $X=1.635 $Y=1.28
+ $X2=1.635 $Y2=1.36
r115 39 40 4.41447 $w=9.12e-07 $l=5.4037e-07 $layer=LI1_cond $X=1.235 $Y=0.95
+ $X2=1.635 $Y2=1.28
r116 35 40 11.0941 $w=1.7e-07 $l=5.65e-07 $layer=LI1_cond $X=2.2 $Y=1.28
+ $X2=1.635 $Y2=1.28
r117 34 47 4.01693 $w=1.7e-07 $l=1.69115e-07 $layer=LI1_cond $X=2.98 $Y=1.28
+ $X2=3.11 $Y2=1.19
r118 34 35 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=2.98 $Y=1.28
+ $X2=2.2 $Y2=1.28
r119 33 48 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=3.145 $Y=1.535
+ $X2=3.145 $Y2=1.18
r120 32 48 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.145 $Y=1.015
+ $X2=3.145 $Y2=1.18
r121 29 43 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=2.035 $Y=1.715
+ $X2=2.035 $Y2=1.36
r122 29 30 43.5886 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=2.05 $Y=1.715
+ $X2=2.05 $Y2=1.865
r123 27 43 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=2.035 $Y=1.345
+ $X2=2.035 $Y2=1.36
r124 26 27 43.5886 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=2.105 $Y=1.195
+ $X2=2.105 $Y2=1.345
r125 21 23 482 $w=1.5e-07 $l=9.4e-07 $layer=POLY_cond $X=3.745 $Y=1.685
+ $X2=3.745 $Y2=2.625
r126 20 33 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=3.31 $Y=1.61
+ $X2=3.145 $Y2=1.535
r127 19 21 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.67 $Y=1.61
+ $X2=3.745 $Y2=1.685
r128 19 20 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=3.67 $Y=1.61
+ $X2=3.31 $Y2=1.61
r129 17 32 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=3.055 $Y=0.445
+ $X2=3.055 $Y2=1.015
r130 13 26 384.574 $w=1.5e-07 $l=7.5e-07 $layer=POLY_cond $X=2.265 $Y=0.445
+ $X2=2.265 $Y2=1.195
r131 9 30 446.106 $w=1.5e-07 $l=8.7e-07 $layer=POLY_cond $X=2.155 $Y=2.735
+ $X2=2.155 $Y2=1.865
r132 2 45 600 $w=1.7e-07 $l=3.34963e-07 $layer=licon1_PDIFF $count=1 $X=1.095
+ $Y=2.035 $X2=1.35 $Y2=1.85
r133 1 39 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=1.095
+ $Y=0.675 $X2=1.235 $Y2=0.95
.ends

.subckt PM_SKY130_FD_SC_LP__DLXBN_1%A_34_407# 1 2 7 9 13 17 18 20 23 27 33 36
c77 27 0 3.53568e-19 $X=2.605 $Y=1.75
c78 23 0 1.27921e-19 $X=2.44 $Y=2.2
r79 30 33 6.27065 $w=3.38e-07 $l=1.85e-07 $layer=LI1_cond $X=0.19 $Y=0.865
+ $X2=0.375 $Y2=0.865
r80 27 28 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.605
+ $Y=1.75 $X2=2.605 $Y2=1.75
r81 25 27 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=2.605 $Y=2.115
+ $X2=2.605 $Y2=1.75
r82 24 36 2.9446 $w=1.7e-07 $l=1.94715e-07 $layer=LI1_cond $X=0.46 $Y=2.2
+ $X2=0.282 $Y2=2.165
r83 23 25 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.44 $Y=2.2
+ $X2=2.605 $Y2=2.115
r84 23 24 129.176 $w=1.68e-07 $l=1.98e-06 $layer=LI1_cond $X=2.44 $Y=2.2
+ $X2=0.46 $Y2=2.2
r85 20 36 3.55013 $w=2.62e-07 $l=1.59499e-07 $layer=LI1_cond $X=0.19 $Y=2.045
+ $X2=0.282 $Y2=2.165
r86 19 30 4.80115 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=0.19 $Y=1.035
+ $X2=0.19 $Y2=0.865
r87 19 20 65.8931 $w=1.68e-07 $l=1.01e-06 $layer=LI1_cond $X=0.19 $Y=1.035
+ $X2=0.19 $Y2=2.045
r88 17 28 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=2.605 $Y=2.105
+ $X2=2.605 $Y2=1.75
r89 17 18 43.5886 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=2.68 $Y=2.105
+ $X2=2.68 $Y2=2.255
r90 13 18 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.845 $Y=2.735
+ $X2=2.845 $Y2=2.255
r91 7 28 35.1288 $w=2.95e-07 $l=2.56076e-07 $layer=POLY_cond $X=2.695 $Y=1.535
+ $X2=2.605 $Y2=1.75
r92 7 9 558.915 $w=1.5e-07 $l=1.09e-06 $layer=POLY_cond $X=2.695 $Y=1.535
+ $X2=2.695 $Y2=0.445
r93 2 36 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.17
+ $Y=2.035 $X2=0.295 $Y2=2.18
r94 1 33 182 $w=1.7e-07 $l=2.498e-07 $layer=licon1_NDIFF $count=1 $X=0.25
+ $Y=0.675 $X2=0.375 $Y2=0.87
.ends

.subckt PM_SKY130_FD_SC_LP__DLXBN_1%A_363_483# 1 2 9 13 18 20 22 23 25 27 29 34
+ 35 37 41 47
c112 41 0 7.24186e-20 $X=3.685 $Y=0.93
c113 35 0 1.55622e-19 $X=3.495 $Y=2.075
c114 34 0 2.93569e-19 $X=3.295 $Y=2.09
c115 9 0 2.22989e-20 $X=3.205 $Y=2.735
r116 41 47 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.685 $Y=0.93
+ $X2=3.685 $Y2=0.765
r117 40 42 8.53881 $w=3.68e-07 $l=1.65e-07 $layer=LI1_cond $X=3.595 $Y=0.93
+ $X2=3.595 $Y2=1.095
r118 40 41 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.685
+ $Y=0.93 $X2=3.685 $Y2=0.93
r119 37 40 5.29501 $w=3.68e-07 $l=1.7e-07 $layer=LI1_cond $X=3.595 $Y=0.76
+ $X2=3.595 $Y2=0.93
r120 34 45 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.295 $Y=2.09
+ $X2=3.295 $Y2=2.255
r121 33 35 7.68295 $w=2.98e-07 $l=2e-07 $layer=LI1_cond $X=3.295 $Y=2.075
+ $X2=3.495 $Y2=2.075
r122 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.295
+ $Y=2.09 $X2=3.295 $Y2=2.09
r123 30 33 9.02747 $w=2.98e-07 $l=2.35e-07 $layer=LI1_cond $X=3.06 $Y=2.075
+ $X2=3.295 $Y2=2.075
r124 27 35 4.061 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=3.495 $Y=1.925
+ $X2=3.495 $Y2=2.075
r125 27 42 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=3.495 $Y=1.925
+ $X2=3.495 $Y2=1.095
r126 24 30 4.061 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=3.06 $Y=2.225 $X2=3.06
+ $Y2=2.075
r127 24 25 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=3.06 $Y=2.225
+ $X2=3.06 $Y2=2.455
r128 22 37 5.30706 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=3.41 $Y=0.76
+ $X2=3.595 $Y2=0.76
r129 22 23 83.1818 $w=1.68e-07 $l=1.275e-06 $layer=LI1_cond $X=3.41 $Y=0.76
+ $X2=2.135 $Y2=0.76
r130 21 29 4.92601 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=2.105 $Y=2.545
+ $X2=1.94 $Y2=2.545
r131 20 25 6.82373 $w=1.8e-07 $l=1.25499e-07 $layer=LI1_cond $X=2.975 $Y=2.545
+ $X2=3.06 $Y2=2.455
r132 20 21 53.6061 $w=1.78e-07 $l=8.7e-07 $layer=LI1_cond $X=2.975 $Y=2.545
+ $X2=2.105 $Y2=2.545
r133 16 23 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=2.04 $Y=0.675
+ $X2=2.135 $Y2=0.76
r134 16 18 13.134 $w=1.88e-07 $l=2.25e-07 $layer=LI1_cond $X=2.04 $Y=0.675
+ $X2=2.04 $Y2=0.45
r135 13 47 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=3.595 $Y=0.445
+ $X2=3.595 $Y2=0.765
r136 9 45 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=3.205 $Y=2.735
+ $X2=3.205 $Y2=2.255
r137 2 29 300 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_PDIFF $count=2 $X=1.815
+ $Y=2.415 $X2=1.94 $Y2=2.57
r138 1 18 182 $w=1.7e-07 $l=2.7037e-07 $layer=licon1_NDIFF $count=1 $X=1.925
+ $Y=0.235 $X2=2.05 $Y2=0.45
.ends

.subckt PM_SKY130_FD_SC_LP__DLXBN_1%A_806_385# 1 2 9 13 18 21 23 25 28 32 34 37
+ 41 44 45 47 48 49 50 52 53 54 57 61 66 69 78
r146 69 75 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.74 $Y=0.51
+ $X2=5.74 $Y2=0.675
r147 68 69 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.74
+ $Y=0.51 $X2=5.74 $Y2=0.51
r148 63 64 20.9993 $w=4.23e-07 $l=6.3e-07 $layer=LI1_cond $X=4.982 $Y=0.465
+ $X2=4.982 $Y2=1.095
r149 61 63 1.22023 $w=4.23e-07 $l=4.5e-08 $layer=LI1_cond $X=4.982 $Y=0.42
+ $X2=4.982 $Y2=0.465
r150 58 78 39.3438 $w=3.3e-07 $l=2.25e-07 $layer=POLY_cond $X=7.46 $Y=1.35
+ $X2=7.685 $Y2=1.35
r151 57 58 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.46
+ $Y=1.35 $X2=7.46 $Y2=1.35
r152 55 57 18.3343 $w=3.28e-07 $l=5.25e-07 $layer=LI1_cond $X=7.46 $Y=0.825
+ $X2=7.46 $Y2=1.35
r153 53 55 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=7.295 $Y=0.74
+ $X2=7.46 $Y2=0.825
r154 53 54 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=7.295 $Y=0.74
+ $X2=6.615 $Y2=0.74
r155 51 54 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.53 $Y=0.825
+ $X2=6.615 $Y2=0.74
r156 51 52 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=6.53 $Y=0.825
+ $X2=6.53 $Y2=1.075
r157 49 52 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.445 $Y=1.16
+ $X2=6.53 $Y2=1.075
r158 49 50 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=6.445 $Y=1.16
+ $X2=5.895 $Y2=1.16
r159 48 50 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.81 $Y=1.075
+ $X2=5.895 $Y2=1.16
r160 47 68 6.0829 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=5.81 $Y=0.675
+ $X2=5.81 $Y2=0.465
r161 47 48 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=5.81 $Y=0.675
+ $X2=5.81 $Y2=1.075
r162 46 63 0.788567 $w=4.2e-07 $l=2.13e-07 $layer=LI1_cond $X=5.195 $Y=0.465
+ $X2=4.982 $Y2=0.465
r163 45 68 2.46213 $w=4.2e-07 $l=8.5e-08 $layer=LI1_cond $X=5.725 $Y=0.465
+ $X2=5.81 $Y2=0.465
r164 45 46 14.5427 $w=4.18e-07 $l=5.3e-07 $layer=LI1_cond $X=5.725 $Y=0.465
+ $X2=5.195 $Y2=0.465
r165 44 66 6.51676 $w=2.47e-07 $l=1.76125e-07 $layer=LI1_cond $X=5.105 $Y=1.925
+ $X2=5.082 $Y2=2.09
r166 44 64 51.1414 $w=1.78e-07 $l=8.3e-07 $layer=LI1_cond $X=5.105 $Y=1.925
+ $X2=5.105 $Y2=1.095
r167 39 66 6.51676 $w=2.47e-07 $l=1.65e-07 $layer=LI1_cond $X=5.082 $Y=2.255
+ $X2=5.082 $Y2=2.09
r168 39 41 23.9635 $w=3.13e-07 $l=6.55e-07 $layer=LI1_cond $X=5.082 $Y=2.255
+ $X2=5.082 $Y2=2.91
r169 37 72 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.195 $Y=2.09
+ $X2=4.195 $Y2=2.255
r170 37 71 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.195 $Y=2.09
+ $X2=4.195 $Y2=1.925
r171 36 37 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.195
+ $Y=2.09 $X2=4.195 $Y2=2.09
r172 34 66 0.330231 $w=3.3e-07 $l=1.57e-07 $layer=LI1_cond $X=4.925 $Y=2.09
+ $X2=5.082 $Y2=2.09
r173 34 36 25.4934 $w=3.28e-07 $l=7.3e-07 $layer=LI1_cond $X=4.925 $Y=2.09
+ $X2=4.195 $Y2=2.09
r174 30 32 146.138 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=5.685 $Y=1.41
+ $X2=5.97 $Y2=1.41
r175 26 78 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.685 $Y=1.515
+ $X2=7.685 $Y2=1.35
r176 26 28 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=7.685 $Y=1.515
+ $X2=7.685 $Y2=2.465
r177 23 78 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.685 $Y=1.185
+ $X2=7.685 $Y2=1.35
r178 23 25 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=7.685 $Y=1.185
+ $X2=7.685 $Y2=0.655
r179 19 32 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.97 $Y=1.485
+ $X2=5.97 $Y2=1.41
r180 19 21 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.97 $Y=1.485
+ $X2=5.97 $Y2=2.145
r181 18 75 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=5.685 $Y=1.015
+ $X2=5.685 $Y2=0.675
r182 16 30 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.685 $Y=1.335
+ $X2=5.685 $Y2=1.41
r183 16 18 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=5.685 $Y=1.335
+ $X2=5.685 $Y2=1.015
r184 13 71 758.894 $w=1.5e-07 $l=1.48e-06 $layer=POLY_cond $X=4.135 $Y=0.445
+ $X2=4.135 $Y2=1.925
r185 9 72 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=4.105 $Y=2.625
+ $X2=4.105 $Y2=2.255
r186 2 66 400 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_PDIFF $count=1 $X=4.95
+ $Y=1.815 $X2=5.09 $Y2=2.03
r187 2 41 400 $w=1.7e-07 $l=1.1629e-06 $layer=licon1_PDIFF $count=1 $X=4.95
+ $Y=1.815 $X2=5.09 $Y2=2.91
r188 1 61 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=4.735
+ $Y=0.235 $X2=4.875 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__DLXBN_1%A_626_47# 1 2 9 13 15 21 24 25 28 29 32 41
r85 36 41 21.8577 $w=3.3e-07 $l=1.25e-07 $layer=POLY_cond $X=4.75 $Y=1.44
+ $X2=4.875 $Y2=1.44
r86 36 38 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=4.75 $Y=1.44 $X2=4.66
+ $Y2=1.44
r87 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.75
+ $Y=1.44 $X2=4.75 $Y2=1.44
r88 32 35 3.54598 $w=2.58e-07 $l=8e-08 $layer=LI1_cond $X=4.715 $Y=1.36
+ $X2=4.715 $Y2=1.44
r89 28 29 10.2539 $w=6.13e-07 $l=1.65e-07 $layer=LI1_cond $X=3.622 $Y=2.56
+ $X2=3.622 $Y2=2.395
r90 26 31 2.70854 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=4.12 $Y=1.36 $X2=3.95
+ $Y2=1.36
r91 25 32 3.22376 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=4.585 $Y=1.36
+ $X2=4.715 $Y2=1.36
r92 25 26 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=4.585 $Y=1.36
+ $X2=4.12 $Y2=1.36
r93 24 31 5.37115 $w=2.38e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.035 $Y=1.275
+ $X2=3.95 $Y2=1.36
r94 23 24 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=4.035 $Y=0.485
+ $X2=4.035 $Y2=1.275
r95 21 31 20.7493 $w=2.38e-07 $l=4.34339e-07 $layer=LI1_cond $X=3.845 $Y=1.745
+ $X2=3.95 $Y2=1.36
r96 21 29 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=3.845 $Y=1.745
+ $X2=3.845 $Y2=2.395
r97 15 23 6.91519 $w=2.1e-07 $l=1.41244e-07 $layer=LI1_cond $X=3.95 $Y=0.38
+ $X2=4.035 $Y2=0.485
r98 15 17 32.7446 $w=2.08e-07 $l=6.2e-07 $layer=LI1_cond $X=3.95 $Y=0.38
+ $X2=3.33 $Y2=0.38
r99 11 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.875 $Y=1.605
+ $X2=4.875 $Y2=1.44
r100 11 13 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=4.875 $Y=1.605
+ $X2=4.875 $Y2=2.445
r101 7 38 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.66 $Y=1.275
+ $X2=4.66 $Y2=1.44
r102 7 9 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=4.66 $Y=1.275
+ $X2=4.66 $Y2=0.655
r103 2 28 300 $w=1.7e-07 $l=3.14245e-07 $layer=licon1_PDIFF $count=2 $X=3.28
+ $Y=2.415 $X2=3.53 $Y2=2.56
r104 1 17 182 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_NDIFF $count=1 $X=3.13
+ $Y=0.235 $X2=3.33 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_LP__DLXBN_1%A_1069_161# 1 2 9 11 13 16 20 22 24 32
r50 31 32 48.0869 $w=3.3e-07 $l=2.75e-07 $layer=POLY_cond $X=6.46 $Y=1.5
+ $X2=6.735 $Y2=1.5
r51 25 31 1.74861 $w=3.3e-07 $l=1e-08 $layer=POLY_cond $X=6.45 $Y=1.5 $X2=6.46
+ $Y2=1.5
r52 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.45
+ $Y=1.5 $X2=6.45 $Y2=1.5
r53 22 24 27.7634 $w=2.18e-07 $l=5.3e-07 $layer=LI1_cond $X=5.92 $Y=1.525
+ $X2=6.45 $Y2=1.525
r54 18 22 9.28663 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=5.755 $Y=1.525
+ $X2=5.92 $Y2=1.525
r55 18 27 18.0854 $w=1.99e-07 $l=2.95e-07 $layer=LI1_cond $X=5.755 $Y=1.525
+ $X2=5.46 $Y2=1.525
r56 18 20 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=5.755 $Y=1.635
+ $X2=5.755 $Y2=1.97
r57 14 27 0.997118 $w=1.9e-07 $l=1.1e-07 $layer=LI1_cond $X=5.46 $Y=1.415
+ $X2=5.46 $Y2=1.525
r58 14 16 23.0574 $w=1.88e-07 $l=3.95e-07 $layer=LI1_cond $X=5.46 $Y=1.415
+ $X2=5.46 $Y2=1.02
r59 11 32 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.735 $Y=1.335
+ $X2=6.735 $Y2=1.5
r60 11 13 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=6.735 $Y=1.335
+ $X2=6.735 $Y2=0.805
r61 7 31 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.46 $Y=1.665
+ $X2=6.46 $Y2=1.5
r62 7 9 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=6.46 $Y=1.665 $X2=6.46
+ $Y2=2.455
r63 2 20 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=5.63
+ $Y=1.825 $X2=5.755 $Y2=1.97
r64 1 16 182 $w=1.7e-07 $l=2.7037e-07 $layer=licon1_NDIFF $count=1 $X=5.345
+ $Y=0.805 $X2=5.47 $Y2=1.02
.ends

.subckt PM_SKY130_FD_SC_LP__DLXBN_1%VPWR 1 2 3 4 5 20 24 28 32 38 43 44 45 47 55
+ 67 73 74 77 80 83 86
r86 86 87 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r87 83 84 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r88 80 81 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r89 77 78 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r90 74 87 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=7.44 $Y2=3.33
r91 73 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r92 71 86 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.635 $Y=3.33
+ $X2=7.47 $Y2=3.33
r93 71 73 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=7.635 $Y=3.33
+ $X2=7.92 $Y2=3.33
r94 70 87 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=7.44 $Y2=3.33
r95 69 70 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r96 67 86 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.305 $Y=3.33
+ $X2=7.47 $Y2=3.33
r97 67 69 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=7.305 $Y=3.33
+ $X2=6.96 $Y2=3.33
r98 66 70 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=6.96
+ $Y2=3.33
r99 65 66 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r100 63 66 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=3.33 $X2=6
+ $Y2=3.33
r101 63 84 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=4.56 $Y2=3.33
r102 62 65 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=5.04 $Y=3.33 $X2=6
+ $Y2=3.33
r103 62 63 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r104 60 83 12.559 $w=1.7e-07 $l=3e-07 $layer=LI1_cond $X=4.755 $Y=3.33 $X2=4.455
+ $Y2=3.33
r105 60 62 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=4.755 $Y=3.33
+ $X2=5.04 $Y2=3.33
r106 56 80 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.68 $Y=3.33
+ $X2=2.515 $Y2=3.33
r107 56 58 91.3369 $w=1.68e-07 $l=1.4e-06 $layer=LI1_cond $X=2.68 $Y=3.33
+ $X2=4.08 $Y2=3.33
r108 55 83 12.559 $w=1.7e-07 $l=3e-07 $layer=LI1_cond $X=4.155 $Y=3.33 $X2=4.455
+ $Y2=3.33
r109 55 58 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=4.155 $Y=3.33
+ $X2=4.08 $Y2=3.33
r110 54 81 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r111 53 54 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r112 51 54 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r113 51 78 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r114 50 53 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=3.33 $X2=2.16
+ $Y2=3.33
r115 50 51 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r116 48 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.97 $Y=3.33
+ $X2=0.805 $Y2=3.33
r117 48 50 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=0.97 $Y=3.33
+ $X2=1.2 $Y2=3.33
r118 47 80 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.35 $Y=3.33
+ $X2=2.515 $Y2=3.33
r119 47 53 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=2.35 $Y=3.33
+ $X2=2.16 $Y2=3.33
r120 45 84 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r121 45 81 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=2.64 $Y2=3.33
r122 45 58 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r123 43 65 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=6.09 $Y=3.33 $X2=6
+ $Y2=3.33
r124 43 44 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=6.09 $Y=3.33
+ $X2=6.22 $Y2=3.33
r125 42 69 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=6.35 $Y=3.33
+ $X2=6.96 $Y2=3.33
r126 42 44 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=6.35 $Y=3.33
+ $X2=6.22 $Y2=3.33
r127 38 41 33.8748 $w=3.28e-07 $l=9.7e-07 $layer=LI1_cond $X=7.47 $Y=1.98
+ $X2=7.47 $Y2=2.95
r128 36 86 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.47 $Y=3.245
+ $X2=7.47 $Y2=3.33
r129 36 41 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=7.47 $Y=3.245
+ $X2=7.47 $Y2=2.95
r130 32 35 20.8326 $w=2.58e-07 $l=4.7e-07 $layer=LI1_cond $X=6.22 $Y=1.97
+ $X2=6.22 $Y2=2.44
r131 30 44 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=6.22 $Y=3.245
+ $X2=6.22 $Y2=3.33
r132 30 35 35.6814 $w=2.58e-07 $l=8.05e-07 $layer=LI1_cond $X=6.22 $Y=3.245
+ $X2=6.22 $Y2=2.44
r133 26 83 2.52064 $w=6e-07 $l=8.5e-08 $layer=LI1_cond $X=4.455 $Y=3.245
+ $X2=4.455 $Y2=3.33
r134 26 28 13.0572 $w=5.98e-07 $l=6.55e-07 $layer=LI1_cond $X=4.455 $Y=3.245
+ $X2=4.455 $Y2=2.59
r135 22 80 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.515 $Y=3.245
+ $X2=2.515 $Y2=3.33
r136 22 24 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=2.515 $Y=3.245
+ $X2=2.515 $Y2=2.93
r137 18 77 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.805 $Y=3.245
+ $X2=0.805 $Y2=3.33
r138 18 20 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=0.805 $Y=3.245
+ $X2=0.805 $Y2=2.55
r139 5 41 400 $w=1.7e-07 $l=1.17584e-06 $layer=licon1_PDIFF $count=1 $X=7.345
+ $Y=1.835 $X2=7.47 $Y2=2.95
r140 5 38 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=7.345
+ $Y=1.835 $X2=7.47 $Y2=1.98
r141 4 35 300 $w=1.7e-07 $l=7.07972e-07 $layer=licon1_PDIFF $count=2 $X=6.045
+ $Y=1.825 $X2=6.245 $Y2=2.44
r142 4 32 600 $w=1.7e-07 $l=2.26164e-07 $layer=licon1_PDIFF $count=1 $X=6.045
+ $Y=1.825 $X2=6.21 $Y2=1.97
r143 3 28 200 $w=1.7e-07 $l=5.60714e-07 $layer=licon1_PDIFF $count=3 $X=4.18
+ $Y=2.415 $X2=4.66 $Y2=2.59
r144 2 24 600 $w=1.7e-07 $l=6.41872e-07 $layer=licon1_PDIFF $count=1 $X=2.23
+ $Y=2.415 $X2=2.515 $Y2=2.93
r145 1 20 600 $w=1.7e-07 $l=6.15244e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=2.035 $X2=0.805 $Y2=2.55
.ends

.subckt PM_SKY130_FD_SC_LP__DLXBN_1%Q_N 1 2 7 8 9 10 18 32 36
r24 32 33 5.27152 $w=5.33e-07 $l=1.65e-07 $layer=LI1_cond $X=6.857 $Y=1.97
+ $X2=6.857 $Y2=1.805
r25 22 36 0.827194 $w=5.33e-07 $l=3.7e-08 $layer=LI1_cond $X=6.857 $Y=2.072
+ $X2=6.857 $Y2=2.035
r26 10 29 3.01814 $w=5.33e-07 $l=1.35e-07 $layer=LI1_cond $X=6.857 $Y=2.775
+ $X2=6.857 $Y2=2.91
r27 9 10 8.27194 $w=5.33e-07 $l=3.7e-07 $layer=LI1_cond $X=6.857 $Y=2.405
+ $X2=6.857 $Y2=2.775
r28 8 36 0.536559 $w=5.33e-07 $l=2.4e-08 $layer=LI1_cond $X=6.857 $Y=2.011
+ $X2=6.857 $Y2=2.035
r29 8 32 0.916621 $w=5.33e-07 $l=4.1e-08 $layer=LI1_cond $X=6.857 $Y=2.011
+ $X2=6.857 $Y2=1.97
r30 8 9 6.90819 $w=5.33e-07 $l=3.09e-07 $layer=LI1_cond $X=6.857 $Y=2.096
+ $X2=6.857 $Y2=2.405
r31 8 22 0.536559 $w=5.33e-07 $l=2.4e-08 $layer=LI1_cond $X=6.857 $Y=2.096
+ $X2=6.857 $Y2=2.072
r32 7 33 4.74535 $w=3.38e-07 $l=1.4e-07 $layer=LI1_cond $X=6.955 $Y=1.665
+ $X2=6.955 $Y2=1.805
r33 7 18 19.8288 $w=3.38e-07 $l=5.85e-07 $layer=LI1_cond $X=6.955 $Y=1.665
+ $X2=6.955 $Y2=1.08
r34 2 32 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=6.535
+ $Y=1.825 $X2=6.675 $Y2=1.97
r35 2 29 400 $w=1.7e-07 $l=1.15288e-06 $layer=licon1_PDIFF $count=1 $X=6.535
+ $Y=1.825 $X2=6.675 $Y2=2.91
r36 1 18 182 $w=1.7e-07 $l=7.61791e-07 $layer=licon1_NDIFF $count=1 $X=6.81
+ $Y=0.385 $X2=6.95 $Y2=1.08
.ends

.subckt PM_SKY130_FD_SC_LP__DLXBN_1%Q 1 2 7 8 9 10 11 12 13 22
r11 13 40 5.98384 $w=2.58e-07 $l=1.35e-07 $layer=LI1_cond $X=7.935 $Y=2.775
+ $X2=7.935 $Y2=2.91
r12 12 13 16.4002 $w=2.58e-07 $l=3.7e-07 $layer=LI1_cond $X=7.935 $Y=2.405
+ $X2=7.935 $Y2=2.775
r13 11 12 18.838 $w=2.58e-07 $l=4.25e-07 $layer=LI1_cond $X=7.935 $Y=1.98
+ $X2=7.935 $Y2=2.405
r14 10 11 13.9623 $w=2.58e-07 $l=3.15e-07 $layer=LI1_cond $X=7.935 $Y=1.665
+ $X2=7.935 $Y2=1.98
r15 9 10 16.4002 $w=2.58e-07 $l=3.7e-07 $layer=LI1_cond $X=7.935 $Y=1.295
+ $X2=7.935 $Y2=1.665
r16 8 9 16.4002 $w=2.58e-07 $l=3.7e-07 $layer=LI1_cond $X=7.935 $Y=0.925
+ $X2=7.935 $Y2=1.295
r17 7 8 16.4002 $w=2.58e-07 $l=3.7e-07 $layer=LI1_cond $X=7.935 $Y=0.555
+ $X2=7.935 $Y2=0.925
r18 7 22 5.98384 $w=2.58e-07 $l=1.35e-07 $layer=LI1_cond $X=7.935 $Y=0.555
+ $X2=7.935 $Y2=0.42
r19 2 40 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=7.76
+ $Y=1.835 $X2=7.9 $Y2=2.91
r20 2 11 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=7.76
+ $Y=1.835 $X2=7.9 $Y2=1.98
r21 1 22 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=7.76
+ $Y=0.235 $X2=7.9 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__DLXBN_1%VGND 1 2 3 4 5 20 24 28 34 38 41 42 43 45 53
+ 62 68 69 72 75 78 81
c104 24 0 1.95136e-19 $X=2.48 $Y=0.4
r105 81 82 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r106 78 79 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r107 75 76 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r108 72 73 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r109 69 82 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=7.44
+ $Y2=0
r110 68 69 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r111 66 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.635 $Y=0 $X2=7.47
+ $Y2=0
r112 66 68 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=7.635 $Y=0
+ $X2=7.92 $Y2=0
r113 65 82 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=7.44
+ $Y2=0
r114 64 65 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r115 62 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.305 $Y=0 $X2=7.47
+ $Y2=0
r116 62 64 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=7.305 $Y=0 $X2=6.96
+ $Y2=0
r117 61 65 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.96
+ $Y2=0
r118 61 79 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=6 $Y=0 $X2=4.56
+ $Y2=0
r119 60 61 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=0 $X2=6 $Y2=0
r120 58 78 8.23795 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=4.6 $Y=0 $X2=4.445
+ $Y2=0
r121 58 60 91.3369 $w=1.68e-07 $l=1.4e-06 $layer=LI1_cond $X=4.6 $Y=0 $X2=6
+ $Y2=0
r122 54 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.645 $Y=0 $X2=2.48
+ $Y2=0
r123 54 56 93.6203 $w=1.68e-07 $l=1.435e-06 $layer=LI1_cond $X=2.645 $Y=0
+ $X2=4.08 $Y2=0
r124 53 78 8.23795 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=4.29 $Y=0 $X2=4.445
+ $Y2=0
r125 53 56 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=4.29 $Y=0 $X2=4.08
+ $Y2=0
r126 52 76 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r127 51 52 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r128 49 52 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r129 49 73 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r130 48 51 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r131 48 49 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r132 46 72 6.25164 $w=1.7e-07 $l=1.08e-07 $layer=LI1_cond $X=0.89 $Y=0 $X2=0.782
+ $Y2=0
r133 46 48 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=0.89 $Y=0 $X2=1.2
+ $Y2=0
r134 45 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.315 $Y=0 $X2=2.48
+ $Y2=0
r135 45 51 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=2.315 $Y=0
+ $X2=2.16 $Y2=0
r136 43 79 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=4.56
+ $Y2=0
r137 43 76 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=4.08 $Y=0
+ $X2=2.64 $Y2=0
r138 43 56 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r139 41 60 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=6.065 $Y=0 $X2=6
+ $Y2=0
r140 41 42 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=6.065 $Y=0 $X2=6.17
+ $Y2=0
r141 40 64 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=6.275 $Y=0
+ $X2=6.96 $Y2=0
r142 40 42 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=6.275 $Y=0 $X2=6.17
+ $Y2=0
r143 36 81 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.47 $Y=0.085
+ $X2=7.47 $Y2=0
r144 36 38 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=7.47 $Y=0.085
+ $X2=7.47 $Y2=0.38
r145 32 42 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=6.17 $Y=0.085
+ $X2=6.17 $Y2=0
r146 32 34 34.5931 $w=2.08e-07 $l=6.55e-07 $layer=LI1_cond $X=6.17 $Y=0.085
+ $X2=6.17 $Y2=0.74
r147 28 30 20.4466 $w=3.08e-07 $l=5.5e-07 $layer=LI1_cond $X=4.445 $Y=0.38
+ $X2=4.445 $Y2=0.93
r148 26 78 0.701276 $w=3.1e-07 $l=8.5e-08 $layer=LI1_cond $X=4.445 $Y=0.085
+ $X2=4.445 $Y2=0
r149 26 28 10.9668 $w=3.08e-07 $l=2.95e-07 $layer=LI1_cond $X=4.445 $Y=0.085
+ $X2=4.445 $Y2=0.38
r150 22 75 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.48 $Y=0.085
+ $X2=2.48 $Y2=0
r151 22 24 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=2.48 $Y=0.085
+ $X2=2.48 $Y2=0.4
r152 18 72 0.512231 $w=2.15e-07 $l=8.5e-08 $layer=LI1_cond $X=0.782 $Y=0.085
+ $X2=0.782 $Y2=0
r153 18 20 42.0776 $w=2.13e-07 $l=7.85e-07 $layer=LI1_cond $X=0.782 $Y=0.085
+ $X2=0.782 $Y2=0.87
r154 5 38 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=7.345
+ $Y=0.235 $X2=7.47 $Y2=0.38
r155 4 34 182 $w=1.7e-07 $l=4.41305e-07 $layer=licon1_NDIFF $count=1 $X=5.76
+ $Y=0.805 $X2=6.17 $Y2=0.74
r156 3 30 182 $w=1.7e-07 $l=8.03959e-07 $layer=licon1_NDIFF $count=1 $X=4.21
+ $Y=0.235 $X2=4.445 $Y2=0.93
r157 3 28 182 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_NDIFF $count=1 $X=4.21
+ $Y=0.235 $X2=4.405 $Y2=0.38
r158 2 24 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=2.34
+ $Y=0.235 $X2=2.48 $Y2=0.4
r159 1 20 182 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_NDIFF $count=1 $X=0.665
+ $Y=0.675 $X2=0.805 $Y2=0.87
.ends

