* File: sky130_fd_sc_lp__and3_2.spice
* Created: Wed Sep  2 09:31:40 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__and3_2.pex.spice"
.subckt sky130_fd_sc_lp__and3_2  VNB VPB A B C VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* C	C
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1008 A_124_47# N_A_M1008_g N_A_27_385#_M1008_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1113 PD=0.63 PS=1.37 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002 A=0.063 P=1.14 MULT=1
MM1004 A_196_47# N_B_M1004_g A_124_47# VNB NSHORT L=0.15 W=0.42 AD=0.0441
+ AS=0.0441 PD=0.63 PS=0.63 NRD=14.28 NRS=14.28 M=1 R=2.8 SA=75000.6 SB=75001.7
+ A=0.063 P=1.14 MULT=1
MM1005 N_VGND_M1005_d N_C_M1005_g A_196_47# VNB NSHORT L=0.15 W=0.42 AD=0.1099
+ AS=0.0441 PD=0.906667 PS=0.63 NRD=37.14 NRS=14.28 M=1 R=2.8 SA=75000.9
+ SB=75001.3 A=0.063 P=1.14 MULT=1
MM1002 N_X_M1002_d N_A_27_385#_M1002_g N_VGND_M1005_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2198 PD=1.12 PS=1.81333 NRD=0 NRS=15.708 M=1 R=5.6 SA=75000.9
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1009 N_X_M1002_d N_A_27_385#_M1009_g N_VGND_M1009_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2352 PD=1.12 PS=2.24 NRD=0 NRS=2.136 M=1 R=5.6 SA=75001.3
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1000 N_VPWR_M1000_d N_A_M1000_g N_A_27_385#_M1000_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75002.1
+ A=0.063 P=1.14 MULT=1
MM1003 N_A_27_385#_M1003_d N_B_M1003_g N_VPWR_M1000_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.07455 AS=0.0588 PD=0.775 PS=0.7 NRD=16.4101 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75001.7 A=0.063 P=1.14 MULT=1
MM1006 N_VPWR_M1006_d N_C_M1006_g N_A_27_385#_M1003_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.095025 AS=0.07455 PD=0.8175 PS=0.775 NRD=0 NRS=18.7544 M=1 R=2.8
+ SA=75001.1 SB=75001.2 A=0.063 P=1.14 MULT=1
MM1001 N_X_M1001_d N_A_27_385#_M1001_g N_VPWR_M1006_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.285075 PD=1.54 PS=2.4525 NRD=0 NRS=4.9447 M=1 R=8.4 SA=75000.7
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1007 N_X_M1001_d N_A_27_385#_M1007_g N_VPWR_M1007_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.3528 PD=1.54 PS=3.08 NRD=0 NRS=2.3443 M=1 R=8.4 SA=75001.1
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.0799 P=10.25
*
.include "sky130_fd_sc_lp__and3_2.pxi.spice"
*
.ends
*
*
