* File: sky130_fd_sc_lp__nand4bb_lp.spice
* Created: Fri Aug 28 10:52:44 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__nand4bb_lp.pex.spice"
.subckt sky130_fd_sc_lp__nand4bb_lp  VNB VPB A_N C D B_N VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B_N	B_N
* D	D
* C	C
* A_N	A_N
* VPB	VPB
* VNB	VNB
MM1002 A_114_47# N_A_N_M1002_g N_A_27_47#_M1002_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1197 PD=0.63 PS=1.41 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1011 N_VGND_M1011_d N_A_N_M1011_g A_114_47# VNB NSHORT L=0.15 W=0.42 AD=0.1197
+ AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1003 A_384_47# N_A_27_47#_M1003_g N_Y_M1003_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1197 PD=0.63 PS=1.41 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.2 A=0.063 P=1.14 MULT=1
MM1005 A_456_47# N_A_332_352#_M1005_g A_384_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.0441 PD=0.66 PS=0.63 NRD=18.564 NRS=14.28 M=1 R=2.8 SA=75000.6
+ SB=75001.8 A=0.063 P=1.14 MULT=1
MM1006 A_534_47# N_C_M1006_g A_456_47# VNB NSHORT L=0.15 W=0.42 AD=0.0504
+ AS=0.0504 PD=0.66 PS=0.66 NRD=18.564 NRS=18.564 M=1 R=2.8 SA=75001 SB=75001.4
+ A=0.063 P=1.14 MULT=1
MM1013 N_VGND_M1013_d N_D_M1013_g A_534_47# VNB NSHORT L=0.15 W=0.42 AD=0.0693
+ AS=0.0504 PD=0.75 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75001.3 SB=75001.1
+ A=0.063 P=1.14 MULT=1
MM1007 A_708_47# N_B_N_M1007_g N_VGND_M1013_d VNB NSHORT L=0.15 W=0.42 AD=0.0441
+ AS=0.0693 PD=0.63 PS=0.75 NRD=14.28 NRS=14.28 M=1 R=2.8 SA=75001.8 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1001 N_A_332_352#_M1001_d N_B_N_M1001_g A_708_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75002.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1008 N_VPWR_M1008_d N_A_N_M1008_g N_A_27_47#_M1008_s VPB PHIGHVT L=0.25 W=1
+ AD=0.14 AS=0.285 PD=1.28 PS=2.57 NRD=0 NRS=0 M=1 R=4 SA=125000 SB=125003
+ A=0.25 P=2.5 MULT=1
MM1000 N_Y_M1000_d N_A_27_47#_M1000_g N_VPWR_M1008_d VPB PHIGHVT L=0.25 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125001 SB=125003 A=0.25
+ P=2.5 MULT=1
MM1009 N_VPWR_M1009_d N_A_332_352#_M1009_g N_Y_M1000_d VPB PHIGHVT L=0.25 W=1
+ AD=0.295 AS=0.14 PD=1.59 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125001 SB=125002
+ A=0.25 P=2.5 MULT=1
MM1004 N_Y_M1004_d N_C_M1004_g N_VPWR_M1009_d VPB PHIGHVT L=0.25 W=1 AD=0.14
+ AS=0.295 PD=1.28 PS=1.59 NRD=0 NRS=61.0503 M=1 R=4 SA=125002 SB=125001 A=0.25
+ P=2.5 MULT=1
MM1012 N_VPWR_M1012_d N_D_M1012_g N_Y_M1004_d VPB PHIGHVT L=0.25 W=1 AD=0.16
+ AS=0.14 PD=1.32 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125003 SB=125001 A=0.25 P=2.5
+ MULT=1
MM1010 N_A_332_352#_M1010_d N_B_N_M1010_g N_VPWR_M1012_d VPB PHIGHVT L=0.25 W=1
+ AD=0.285 AS=0.16 PD=2.57 PS=1.32 NRD=0 NRS=7.8603 M=1 R=4 SA=125003 SB=125000
+ A=0.25 P=2.5 MULT=1
DX14_noxref VNB VPB NWDIODE A=8.7655 P=13.13
c_47 VNB 0 1.06129e-19 $X=0 $Y=0
*
.include "sky130_fd_sc_lp__nand4bb_lp.pxi.spice"
*
.ends
*
*
