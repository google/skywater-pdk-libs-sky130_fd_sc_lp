* File: sky130_fd_sc_lp__inputisolatch_lp.spice
* Created: Fri Aug 28 10:37:39 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__inputisolatch_lp.pex.spice"
.subckt sky130_fd_sc_lp__inputisolatch_lp  VNB VPB D SLEEP_B VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* SLEEP_B	SLEEP_B
* D	D
* VPB	VPB
* VNB	VNB
MM1018 N_VGND_M1018_d N_A_21_179#_M1018_g N_A_36_73#_M1018_s VNB NSHORT L=0.15
+ W=0.42 AD=0.10115 AS=0.1197 PD=1.075 PS=1.41 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1010 A_232_125# N_D_M1010_g N_VGND_M1018_d VNB NSHORT L=0.15 W=0.42 AD=0.0504
+ AS=0.10115 PD=0.66 PS=1.075 NRD=18.564 NRS=53.088 M=1 R=2.8 SA=75000.4
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1008 N_A_281_535#_M1008_d N_A_36_73#_M1008_g A_232_125# VNB NSHORT L=0.15
+ W=0.42 AD=0.10115 AS=0.0504 PD=1.075 PS=0.66 NRD=53.088 NRS=18.564 M=1 R=2.8
+ SA=75000.8 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1013 A_419_73# N_A_21_179#_M1013_g N_A_281_535#_M1008_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0756 AS=0.10115 PD=0.78 PS=1.075 NRD=35.712 NRS=0 M=1 R=2.8
+ SA=75000.8 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1015 A_521_73# N_A_458_293#_M1015_g A_419_73# VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.0756 PD=0.66 PS=0.78 NRD=18.564 NRS=35.712 M=1 R=2.8 SA=75001.3
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1000 N_VGND_M1000_d N_A_458_293#_M1000_g A_521_73# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0504 PD=1.41 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75001.7
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1002 A_837_93# N_SLEEP_B_M1002_g N_A_21_179#_M1002_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1197 PD=0.63 PS=1.41 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1017 N_VGND_M1017_d N_SLEEP_B_M1017_g A_837_93# VNB NSHORT L=0.15 W=0.42
+ AD=0.0735 AS=0.0441 PD=0.77 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1016 A_1009_93# N_A_281_535#_M1016_g N_VGND_M1017_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0735 PD=0.63 PS=0.77 NRD=14.28 NRS=19.992 M=1 R=2.8 SA=75001.1
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1007 N_A_458_293#_M1007_d N_A_281_535#_M1007_g A_1009_93# VNB NSHORT L=0.15
+ W=0.42 AD=0.1113 AS=0.0441 PD=1.37 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8
+ SA=75001.4 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1009 A_1284_177# N_A_281_535#_M1009_g N_VGND_M1009_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.126 PD=0.63 PS=1.44 NRD=14.28 NRS=4.284 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1005 N_Q_M1005_d N_A_281_535#_M1005_g A_1284_177# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1001 A_117_535# N_D_M1001_g N_VPWR_M1001_s VPB PHIGHVT L=0.15 W=0.42 AD=0.1407
+ AS=0.1197 PD=1.09 PS=1.41 NRD=131.32 NRS=0 M=1 R=2.8 SA=75000.2 SB=75002.7
+ A=0.063 P=1.14 MULT=1
MM1019 N_A_281_535#_M1019_d N_A_21_179#_M1019_g A_117_535# VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0979606 AS=0.1407 PD=0.825211 PS=1.09 NRD=83.5871 NRS=131.32 M=1
+ R=2.8 SA=75001 SB=75001.9 A=0.063 P=1.14 MULT=1
MM1011 A_410_419# N_A_36_73#_M1011_g N_A_281_535#_M1019_d VPB PHIGHVT L=0.25 W=1
+ AD=0.12 AS=0.233239 PD=1.24 PS=1.96479 NRD=12.7853 NRS=0 M=1 R=4 SA=125001
+ SB=125001 A=0.25 P=2.5 MULT=1
MM1003 N_VPWR_M1003_d N_A_458_293#_M1003_g A_410_419# VPB PHIGHVT L=0.25 W=1
+ AD=0.14 AS=0.12 PD=1.28 PS=1.24 NRD=0 NRS=12.7853 M=1 R=4 SA=125001 SB=125001
+ A=0.25 P=2.5 MULT=1
MM1014 N_A_36_73#_M1014_d N_A_21_179#_M1014_g N_VPWR_M1003_d VPB PHIGHVT L=0.25
+ W=1 AD=0.285 AS=0.14 PD=2.57 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125002 SB=125000
+ A=0.25 P=2.5 MULT=1
MM1006 N_VPWR_M1006_d N_SLEEP_B_M1006_g N_A_21_179#_M1006_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.32 AS=0.256 PD=2.28 PS=2.08 NRD=66.1723 NRS=35.3812 M=1 R=4.26667
+ SA=75000.3 SB=75000.4 A=0.096 P=1.58 MULT=1
MM1012 N_VPWR_M1012_d N_A_281_535#_M1012_g N_A_458_293#_M1012_s VPB PHIGHVT
+ L=0.25 W=1 AD=0.14 AS=0.285 PD=1.28 PS=2.57 NRD=0 NRS=0 M=1 R=4 SA=125000
+ SB=125001 A=0.25 P=2.5 MULT=1
MM1004 N_Q_M1004_d N_A_281_535#_M1004_g N_VPWR_M1012_d VPB PHIGHVT L=0.25 W=1
+ AD=0.34 AS=0.14 PD=2.68 PS=1.28 NRD=10.8153 NRS=0 M=1 R=4 SA=125001 SB=125000
+ A=0.25 P=2.5 MULT=1
DX20_noxref VNB VPB NWDIODE A=14.1367 P=18.89
*
.include "sky130_fd_sc_lp__inputisolatch_lp.pxi.spice"
*
.ends
*
*
