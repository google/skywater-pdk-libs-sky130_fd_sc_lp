* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_lp__and3b_2 A_N B C VGND VNB VPB VPWR X
*.PININFO A_N:I B:I C:I VGND:I VNB:I VPB:I VPWR:I X:O
MMP0 y A VPB phighvt m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 y B VPB phighvt m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 y C VPB phighvt m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIP0 A A_N VPB phighvt m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIP1 X y VPB phighvt m=2 w=1.26 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A VNB nshort m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265 sd=0.28
+ topography=normal area=0.063 perim=1.14
MMN1 sndA B VNB nshort m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 sndB C VNB nshort m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN0 A A_N VNB nshort m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN1 X y VNB nshort m=2 w=0.84 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_sc_lp__and3b_2
