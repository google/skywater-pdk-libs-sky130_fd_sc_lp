# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__a31o_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_lp__a31o_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.720000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.915000 1.415000 6.565000 1.760000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.955000 1.415000 5.605000 1.760000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.515000 1.415000 4.645000 1.750000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.155000 1.210000 0.425000 1.760000 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  1.593200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.025000 0.975000 2.900000 1.185000 ;
        RECT 1.025000 1.185000 1.690000 1.760000 ;
        RECT 1.405000 1.760000 1.690000 1.930000 ;
        RECT 1.405000 1.930000 3.575000 2.260000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 6.720000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 6.720000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.720000 0.085000 ;
      RECT 0.000000  3.245000 6.720000 3.415000 ;
      RECT 0.095000  0.085000 0.425000 1.040000 ;
      RECT 0.095000  1.930000 0.425000 2.905000 ;
      RECT 0.095000  2.905000 1.285000 3.075000 ;
      RECT 0.595000  0.255000 0.785000 0.635000 ;
      RECT 0.595000  0.635000 3.250000 0.805000 ;
      RECT 0.595000  0.805000 0.855000 2.735000 ;
      RECT 0.955000  0.085000 1.285000 0.465000 ;
      RECT 1.025000  1.930000 1.235000 2.440000 ;
      RECT 1.025000  2.440000 4.385000 2.610000 ;
      RECT 1.025000  2.610000 1.285000 2.905000 ;
      RECT 1.890000  1.355000 3.250000 1.645000 ;
      RECT 1.955000  2.780000 2.285000 3.245000 ;
      RECT 2.045000  0.085000 2.375000 0.465000 ;
      RECT 2.815000  2.780000 3.145000 3.245000 ;
      RECT 3.080000  0.805000 3.250000 1.075000 ;
      RECT 3.080000  1.075000 6.195000 1.245000 ;
      RECT 3.080000  1.245000 3.250000 1.355000 ;
      RECT 3.095000  0.085000 3.425000 0.465000 ;
      RECT 3.605000  0.345000 3.935000 0.725000 ;
      RECT 3.605000  0.725000 5.335000 0.905000 ;
      RECT 3.675000  2.780000 4.005000 3.245000 ;
      RECT 4.105000  0.085000 4.305000 0.545000 ;
      RECT 4.105000  1.930000 6.125000 2.100000 ;
      RECT 4.105000  2.100000 4.385000 2.440000 ;
      RECT 4.175000  2.610000 4.385000 3.075000 ;
      RECT 4.555000  2.270000 4.885000 3.245000 ;
      RECT 4.575000  0.275000 6.625000 0.445000 ;
      RECT 4.575000  0.445000 5.695000 0.555000 ;
      RECT 5.055000  2.100000 5.265000 3.075000 ;
      RECT 5.435000  2.270000 5.765000 3.245000 ;
      RECT 5.515000  0.555000 5.695000 0.645000 ;
      RECT 5.865000  0.615000 6.195000 1.075000 ;
      RECT 5.935000  2.100000 6.125000 3.075000 ;
      RECT 6.295000  1.930000 6.625000 3.245000 ;
      RECT 6.365000  0.445000 6.625000 1.195000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
  END
END sky130_fd_sc_lp__a31o_4
END LIBRARY
