* File: sky130_fd_sc_lp__buflp_1.pex.spice
* Created: Wed Sep  2 09:36:27 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__BUFLP_1%A_86_21# 1 2 9 13 15 19 22 24 27 28 30 31 34
+ 37 42
r64 43 44 30.474 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=0.985 $Y=1.44
+ $X2=0.985 $Y2=1.515
r65 39 40 3.67308 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=2.07 $Y=0.93
+ $X2=2.07 $Y2=1.015
r66 37 39 3.66686 $w=3.28e-07 $l=1.05e-07 $layer=LI1_cond $X=2.07 $Y=0.825
+ $X2=2.07 $Y2=0.93
r67 34 40 52.7819 $w=2.48e-07 $l=1.145e-06 $layer=LI1_cond $X=2.11 $Y=2.16
+ $X2=2.11 $Y2=1.015
r68 30 39 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.905 $Y=0.93
+ $X2=2.07 $Y2=0.93
r69 30 31 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=1.905 $Y=0.93
+ $X2=1.15 $Y2=0.93
r70 28 43 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=0.985 $Y=1.35
+ $X2=0.985 $Y2=1.44
r71 28 42 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.985 $Y=1.35
+ $X2=0.985 $Y2=1.185
r72 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.985
+ $Y=1.35 $X2=0.985 $Y2=1.35
r73 25 31 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.985 $Y=1.015
+ $X2=1.15 $Y2=0.93
r74 25 27 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=0.985 $Y=1.015
+ $X2=0.985 $Y2=1.35
r75 22 44 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=0.895 $Y=2.465
+ $X2=0.895 $Y2=1.515
r76 19 42 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.895 $Y=0.655
+ $X2=0.895 $Y2=1.185
r77 16 24 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.58 $Y=1.44
+ $X2=0.505 $Y2=1.44
r78 15 43 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.82 $Y=1.44
+ $X2=0.985 $Y2=1.44
r79 15 16 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=0.82 $Y=1.44
+ $X2=0.58 $Y2=1.44
r80 11 24 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.505 $Y=1.515
+ $X2=0.505 $Y2=1.44
r81 11 13 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=0.505 $Y=1.515
+ $X2=0.505 $Y2=2.465
r82 7 24 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.505 $Y=1.365
+ $X2=0.505 $Y2=1.44
r83 7 9 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=0.505 $Y=1.365
+ $X2=0.505 $Y2=0.655
r84 2 34 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=1.93
+ $Y=2.015 $X2=2.07 $Y2=2.16
r85 1 37 182 $w=1.7e-07 $l=2.29565e-07 $layer=licon1_NDIFF $count=1 $X=1.93
+ $Y=0.655 $X2=2.07 $Y2=0.825
.ends

.subckt PM_SKY130_FD_SC_LP__BUFLP_1%A 1 3 6 8 10 13 15 16 17 18 27 28
r38 26 28 42.841 $w=3.3e-07 $l=2.45e-07 $layer=POLY_cond $X=1.61 $Y=1.35
+ $X2=1.855 $Y2=1.35
r39 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.61
+ $Y=1.35 $X2=1.61 $Y2=1.35
r40 23 26 25.3549 $w=3.3e-07 $l=1.45e-07 $layer=POLY_cond $X=1.465 $Y=1.35
+ $X2=1.61 $Y2=1.35
r41 17 18 12.183 $w=3.48e-07 $l=3.7e-07 $layer=LI1_cond $X=1.62 $Y=2.405
+ $X2=1.62 $Y2=2.775
r42 16 17 12.183 $w=3.48e-07 $l=3.7e-07 $layer=LI1_cond $X=1.62 $Y=2.035
+ $X2=1.62 $Y2=2.405
r43 15 16 12.183 $w=3.48e-07 $l=3.7e-07 $layer=LI1_cond $X=1.62 $Y=1.665
+ $X2=1.62 $Y2=2.035
r44 15 27 10.372 $w=3.48e-07 $l=3.15e-07 $layer=LI1_cond $X=1.62 $Y=1.665
+ $X2=1.62 $Y2=1.35
r45 11 28 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.855 $Y=1.515
+ $X2=1.855 $Y2=1.35
r46 11 13 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=1.855 $Y=1.515
+ $X2=1.855 $Y2=2.335
r47 8 28 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.855 $Y=1.185
+ $X2=1.855 $Y2=1.35
r48 8 10 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.855 $Y=1.185
+ $X2=1.855 $Y2=0.865
r49 4 23 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.465 $Y=1.515
+ $X2=1.465 $Y2=1.35
r50 4 6 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=1.465 $Y=1.515
+ $X2=1.465 $Y2=2.335
r51 1 23 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.465 $Y=1.185
+ $X2=1.465 $Y2=1.35
r52 1 3 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.465 $Y=1.185
+ $X2=1.465 $Y2=0.865
.ends

.subckt PM_SKY130_FD_SC_LP__BUFLP_1%X 1 2 7 8 9 10 11 12 13 22
r17 13 40 4.71454 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=0.29 $Y=2.775
+ $X2=0.29 $Y2=2.91
r18 12 13 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.29 $Y=2.405
+ $X2=0.29 $Y2=2.775
r19 11 12 14.8421 $w=3.28e-07 $l=4.25e-07 $layer=LI1_cond $X=0.29 $Y=1.98
+ $X2=0.29 $Y2=2.405
r20 10 11 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=0.29 $Y=1.665
+ $X2=0.29 $Y2=1.98
r21 9 10 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.29 $Y=1.295
+ $X2=0.29 $Y2=1.665
r22 8 9 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.29 $Y=0.925 $X2=0.29
+ $Y2=1.295
r23 7 8 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.29 $Y=0.555 $X2=0.29
+ $Y2=0.925
r24 7 22 4.71454 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=0.29 $Y=0.555
+ $X2=0.29 $Y2=0.42
r25 2 40 400 $w=1.7e-07 $l=1.14521e-06 $layer=licon1_PDIFF $count=1 $X=0.145
+ $Y=1.835 $X2=0.29 $Y2=2.91
r26 2 11 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.145
+ $Y=1.835 $X2=0.29 $Y2=1.98
r27 1 22 91 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=2 $X=0.145
+ $Y=0.235 $X2=0.29 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__BUFLP_1%VPWR 1 6 12 14 21 22 25
r29 21 22 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r30 19 25 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.275 $Y=3.33
+ $X2=1.11 $Y2=3.33
r31 19 21 57.738 $w=1.68e-07 $l=8.85e-07 $layer=LI1_cond $X=1.275 $Y=3.33
+ $X2=2.16 $Y2=3.33
r32 16 17 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r33 14 25 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.945 $Y=3.33
+ $X2=1.11 $Y2=3.33
r34 14 16 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=0.945 $Y=3.33
+ $X2=0.72 $Y2=3.33
r35 12 22 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r36 12 17 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r37 12 25 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r38 9 11 16.9374 $w=3.28e-07 $l=4.85e-07 $layer=LI1_cond $X=1.11 $Y=2.465
+ $X2=1.11 $Y2=2.95
r39 6 9 16.9374 $w=3.28e-07 $l=4.85e-07 $layer=LI1_cond $X=1.11 $Y=1.98 $X2=1.11
+ $Y2=2.465
r40 4 25 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.11 $Y=3.245 $X2=1.11
+ $Y2=3.33
r41 4 11 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.11 $Y=3.245
+ $X2=1.11 $Y2=2.95
r42 1 11 600 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=0.97
+ $Y=1.835 $X2=1.11 $Y2=2.95
r43 1 9 600 $w=1.7e-07 $l=6.96491e-07 $layer=licon1_PDIFF $count=1 $X=0.97
+ $Y=1.835 $X2=1.11 $Y2=2.465
r44 1 6 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.97
+ $Y=1.835 $X2=1.11 $Y2=1.98
.ends

.subckt PM_SKY130_FD_SC_LP__BUFLP_1%VGND 1 6 8 10 17 18 21
r32 17 18 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r33 15 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.275 $Y=0 $X2=1.11
+ $Y2=0
r34 15 17 57.738 $w=1.68e-07 $l=8.85e-07 $layer=LI1_cond $X=1.275 $Y=0 $X2=2.16
+ $Y2=0
r35 12 13 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r36 10 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.945 $Y=0 $X2=1.11
+ $Y2=0
r37 10 12 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=0.945 $Y=0 $X2=0.72
+ $Y2=0
r38 8 18 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r39 8 13 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r40 8 21 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r41 4 21 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.11 $Y=0.085 $X2=1.11
+ $Y2=0
r42 4 6 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=1.11 $Y=0.085 $X2=1.11
+ $Y2=0.445
r43 1 6 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.97
+ $Y=0.235 $X2=1.11 $Y2=0.445
.ends

