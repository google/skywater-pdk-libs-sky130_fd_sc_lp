* File: sky130_fd_sc_lp__clkbuf_16.pxi.spice
* Created: Wed Sep  2 09:38:14 2020
* 
x_PM_SKY130_FD_SC_LP__CLKBUF_16%A N_A_M1011_g N_A_M1004_g N_A_M1026_g
+ N_A_M1021_g N_A_M1029_g N_A_M1025_g N_A_M1030_g N_A_M1035_g A A A N_A_c_177_n
+ PM_SKY130_FD_SC_LP__CLKBUF_16%A
x_PM_SKY130_FD_SC_LP__CLKBUF_16%A_116_47# N_A_116_47#_M1011_d
+ N_A_116_47#_M1029_d N_A_116_47#_M1004_s N_A_116_47#_M1025_s
+ N_A_116_47#_M1001_g N_A_116_47#_M1000_g N_A_116_47#_M1003_g
+ N_A_116_47#_M1002_g N_A_116_47#_M1005_g N_A_116_47#_M1010_g
+ N_A_116_47#_M1006_g N_A_116_47#_M1013_g N_A_116_47#_M1007_g
+ N_A_116_47#_M1014_g N_A_116_47#_M1008_g N_A_116_47#_M1015_g
+ N_A_116_47#_M1009_g N_A_116_47#_M1016_g N_A_116_47#_M1012_g
+ N_A_116_47#_M1017_g N_A_116_47#_M1018_g N_A_116_47#_M1019_g
+ N_A_116_47#_M1020_g N_A_116_47#_M1022_g N_A_116_47#_M1023_g
+ N_A_116_47#_M1028_g N_A_116_47#_M1024_g N_A_116_47#_M1032_g
+ N_A_116_47#_M1027_g N_A_116_47#_M1034_g N_A_116_47#_M1031_g
+ N_A_116_47#_M1037_g N_A_116_47#_M1033_g N_A_116_47#_M1038_g
+ N_A_116_47#_c_272_n N_A_116_47#_M1036_g N_A_116_47#_M1039_g
+ N_A_116_47#_c_275_n N_A_116_47#_c_417_p N_A_116_47#_c_276_n
+ N_A_116_47#_c_277_n N_A_116_47#_c_308_n N_A_116_47#_c_309_n
+ N_A_116_47#_c_278_n N_A_116_47#_c_418_p N_A_116_47#_c_279_n
+ N_A_116_47#_c_310_n N_A_116_47#_c_280_n N_A_116_47#_c_281_n
+ N_A_116_47#_c_282_n N_A_116_47#_c_312_n N_A_116_47#_c_283_n
+ N_A_116_47#_c_284_n N_A_116_47#_c_285_n N_A_116_47#_c_286_n
+ N_A_116_47#_c_287_n N_A_116_47#_c_288_n N_A_116_47#_c_289_n
+ N_A_116_47#_c_290_n N_A_116_47#_c_291_n
+ PM_SKY130_FD_SC_LP__CLKBUF_16%A_116_47#
x_PM_SKY130_FD_SC_LP__CLKBUF_16%VPWR N_VPWR_M1004_d N_VPWR_M1021_d
+ N_VPWR_M1035_d N_VPWR_M1002_d N_VPWR_M1013_d N_VPWR_M1015_d N_VPWR_M1017_d
+ N_VPWR_M1022_d N_VPWR_M1032_d N_VPWR_M1037_d N_VPWR_M1039_d N_VPWR_c_635_n
+ N_VPWR_c_636_n N_VPWR_c_637_n N_VPWR_c_638_n N_VPWR_c_639_n N_VPWR_c_640_n
+ N_VPWR_c_641_n N_VPWR_c_642_n N_VPWR_c_643_n N_VPWR_c_644_n N_VPWR_c_645_n
+ N_VPWR_c_646_n N_VPWR_c_647_n N_VPWR_c_648_n N_VPWR_c_649_n N_VPWR_c_650_n
+ N_VPWR_c_651_n N_VPWR_c_652_n N_VPWR_c_653_n VPWR N_VPWR_c_654_n
+ N_VPWR_c_655_n N_VPWR_c_656_n N_VPWR_c_657_n N_VPWR_c_658_n N_VPWR_c_659_n
+ N_VPWR_c_660_n N_VPWR_c_661_n N_VPWR_c_662_n N_VPWR_c_663_n N_VPWR_c_664_n
+ N_VPWR_c_665_n N_VPWR_c_666_n N_VPWR_c_634_n VPWR
+ PM_SKY130_FD_SC_LP__CLKBUF_16%VPWR
x_PM_SKY130_FD_SC_LP__CLKBUF_16%X N_X_M1001_s N_X_M1005_s N_X_M1007_s
+ N_X_M1009_s N_X_M1018_s N_X_M1023_s N_X_M1027_s N_X_M1033_s N_X_M1000_s
+ N_X_M1010_s N_X_M1014_s N_X_M1016_s N_X_M1019_s N_X_M1028_s N_X_M1034_s
+ N_X_M1038_s X N_X_c_827_n N_X_c_828_n N_X_c_829_n N_X_c_830_n N_X_c_831_n
+ N_X_c_832_n N_X_c_833_n N_X_c_834_n N_X_c_909_n
+ PM_SKY130_FD_SC_LP__CLKBUF_16%X
x_PM_SKY130_FD_SC_LP__CLKBUF_16%VGND N_VGND_M1011_s N_VGND_M1026_s
+ N_VGND_M1030_s N_VGND_M1003_d N_VGND_M1006_d N_VGND_M1008_d N_VGND_M1012_d
+ N_VGND_M1020_d N_VGND_M1024_d N_VGND_M1031_d N_VGND_M1036_d N_VGND_c_1006_n
+ N_VGND_c_1007_n N_VGND_c_1008_n N_VGND_c_1009_n N_VGND_c_1010_n
+ N_VGND_c_1011_n N_VGND_c_1012_n N_VGND_c_1013_n N_VGND_c_1014_n
+ N_VGND_c_1015_n N_VGND_c_1016_n N_VGND_c_1017_n N_VGND_c_1018_n
+ N_VGND_c_1019_n N_VGND_c_1020_n N_VGND_c_1021_n N_VGND_c_1022_n
+ N_VGND_c_1023_n VGND N_VGND_c_1024_n N_VGND_c_1025_n N_VGND_c_1026_n
+ N_VGND_c_1027_n N_VGND_c_1028_n N_VGND_c_1029_n N_VGND_c_1030_n
+ N_VGND_c_1031_n N_VGND_c_1032_n N_VGND_c_1033_n N_VGND_c_1034_n
+ N_VGND_c_1035_n N_VGND_c_1036_n N_VGND_c_1037_n VGND
+ PM_SKY130_FD_SC_LP__CLKBUF_16%VGND
cc_1 VNB N_A_M1011_g 0.0509575f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=0.445
cc_2 VNB N_A_M1004_g 0.0160144f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.465
cc_3 VNB N_A_M1026_g 0.0330149f $X=-0.19 $Y=-0.245 $X2=0.935 $Y2=0.445
cc_4 VNB N_A_M1021_g 0.0101204f $X=-0.19 $Y=-0.245 $X2=0.935 $Y2=2.465
cc_5 VNB N_A_M1029_g 0.0329924f $X=-0.19 $Y=-0.245 $X2=1.365 $Y2=0.445
cc_6 VNB N_A_M1025_g 0.0101148f $X=-0.19 $Y=-0.245 $X2=1.365 $Y2=2.465
cc_7 VNB N_A_M1030_g 0.0369246f $X=-0.19 $Y=-0.245 $X2=1.795 $Y2=0.445
cc_8 VNB N_A_M1035_g 0.0115107f $X=-0.19 $Y=-0.245 $X2=1.795 $Y2=2.465
cc_9 VNB A 0.0133586f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.21
cc_10 VNB N_A_c_177_n 0.0806664f $X=-0.19 $Y=-0.245 $X2=1.795 $Y2=1.29
cc_11 VNB N_A_116_47#_M1001_g 0.0245706f $X=-0.19 $Y=-0.245 $X2=0.935 $Y2=2.465
cc_12 VNB N_A_116_47#_M1000_g 0.0074914f $X=-0.19 $Y=-0.245 $X2=1.365 $Y2=0.445
cc_13 VNB N_A_116_47#_M1003_g 0.0380497f $X=-0.19 $Y=-0.245 $X2=1.365 $Y2=2.465
cc_14 VNB N_A_116_47#_M1002_g 0.00600768f $X=-0.19 $Y=-0.245 $X2=1.795 $Y2=0.445
cc_15 VNB N_A_116_47#_M1005_g 0.0380497f $X=-0.19 $Y=-0.245 $X2=1.795 $Y2=2.465
cc_16 VNB N_A_116_47#_M1010_g 0.00600768f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.21
cc_17 VNB N_A_116_47#_M1006_g 0.0380497f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.29
cc_18 VNB N_A_116_47#_M1013_g 0.00600768f $X=-0.19 $Y=-0.245 $X2=0.675 $Y2=1.29
cc_19 VNB N_A_116_47#_M1007_g 0.0380497f $X=-0.19 $Y=-0.245 $X2=1.695 $Y2=1.29
cc_20 VNB N_A_116_47#_M1014_g 0.00600768f $X=-0.19 $Y=-0.245 $X2=0.675 $Y2=1.29
cc_21 VNB N_A_116_47#_M1008_g 0.0380497f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_116_47#_M1015_g 0.00600768f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_116_47#_M1009_g 0.0380497f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_116_47#_M1016_g 0.00600768f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_116_47#_M1012_g 0.0380497f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_116_47#_M1017_g 0.00600768f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_116_47#_M1018_g 0.0380497f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_116_47#_M1019_g 0.00600768f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_116_47#_M1020_g 0.0380488f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_116_47#_M1022_g 0.00600748f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_116_47#_M1023_g 0.038077f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_116_47#_M1028_g 0.00600754f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_116_47#_M1024_g 0.0380497f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_116_47#_M1032_g 0.00600768f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_116_47#_M1027_g 0.0380497f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_116_47#_M1034_g 0.00600768f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_116_47#_M1031_g 0.0380497f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_116_47#_M1037_g 0.00600768f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_116_47#_M1033_g 0.0381391f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_116_47#_M1038_g 0.00600768f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_116_47#_c_272_n 0.408604f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_116_47#_M1036_g 0.0565027f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_116_47#_M1039_g 0.00953809f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_116_47#_c_275_n 0.00247758f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_116_47#_c_276_n 0.00566142f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_116_47#_c_277_n 0.00442754f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_116_47#_c_278_n 0.00208514f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_116_47#_c_279_n 0.00963554f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_116_47#_c_280_n 0.00249619f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_116_47#_c_281_n 0.00232292f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_116_47#_c_282_n 0.00199612f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_116_47#_c_283_n 0.00667702f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_116_47#_c_284_n 0.00194335f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_116_47#_c_285_n 0.00194335f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_116_47#_c_286_n 0.00194335f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_116_47#_c_287_n 0.00194335f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_116_47#_c_288_n 0.00194335f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_116_47#_c_289_n 0.00194335f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_116_47#_c_290_n 0.0434608f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_116_47#_c_291_n 0.00194335f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_VPWR_c_634_n 0.40251f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_X_c_827_n 0.0130638f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_X_c_828_n 0.0141044f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_X_c_829_n 0.0141044f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_X_c_830_n 0.0141044f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_X_c_831_n 0.0140824f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_X_c_832_n 0.0141475f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_X_c_833_n 0.0141044f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_X_c_834_n 0.0145687f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_VGND_c_1006_n 0.0118373f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.21
cc_71 VNB N_VGND_c_1007_n 0.0188511f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_VGND_c_1008_n 0.00408721f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_VGND_c_1009_n 0.0135711f $X=-0.19 $Y=-0.245 $X2=0.675 $Y2=1.29
cc_74 VNB N_VGND_c_1010_n 3.16879e-19 $X=-0.19 $Y=-0.245 $X2=1.695 $Y2=1.29
cc_75 VNB N_VGND_c_1011_n 3.16188e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_VGND_c_1012_n 3.16188e-19 $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=1.29
cc_77 VNB N_VGND_c_1013_n 3.16188e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_VGND_c_1014_n 3.17051e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_VGND_c_1015_n 0.0135769f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_VGND_c_1016_n 3.17051e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_VGND_c_1017_n 3.16188e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_VGND_c_1018_n 0.012121f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_VGND_c_1019_n 0.0183788f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_VGND_c_1020_n 0.0134631f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_VGND_c_1021_n 0.00410281f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_VGND_c_1022_n 0.0134631f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_VGND_c_1023_n 0.00403622f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_VGND_c_1024_n 0.0164895f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_VGND_c_1025_n 0.0134631f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_VGND_c_1026_n 0.0134631f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_VGND_c_1027_n 0.0134631f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_VGND_c_1028_n 0.0134631f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_93 VNB N_VGND_c_1029_n 0.00536026f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_94 VNB N_VGND_c_1030_n 0.0163239f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_95 VNB N_VGND_c_1031_n 0.0159754f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_96 VNB N_VGND_c_1032_n 0.00410281f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_97 VNB N_VGND_c_1033_n 0.00410281f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_98 VNB N_VGND_c_1034_n 0.00410281f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_99 VNB N_VGND_c_1035_n 0.00410281f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_100 VNB N_VGND_c_1036_n 0.00410281f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_101 VNB N_VGND_c_1037_n 0.450575f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_102 VPB N_A_M1004_g 0.0277461f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=2.465
cc_103 VPB N_A_M1021_g 0.0185278f $X=-0.19 $Y=1.655 $X2=0.935 $Y2=2.465
cc_104 VPB N_A_M1025_g 0.018496f $X=-0.19 $Y=1.655 $X2=1.365 $Y2=2.465
cc_105 VPB N_A_M1035_g 0.0218179f $X=-0.19 $Y=1.655 $X2=1.795 $Y2=2.465
cc_106 VPB N_A_116_47#_M1000_g 0.0231789f $X=-0.19 $Y=1.655 $X2=1.365 $Y2=0.445
cc_107 VPB N_A_116_47#_M1002_g 0.0196061f $X=-0.19 $Y=1.655 $X2=1.795 $Y2=0.445
cc_108 VPB N_A_116_47#_M1010_g 0.0196061f $X=-0.19 $Y=1.655 $X2=1.595 $Y2=1.21
cc_109 VPB N_A_116_47#_M1013_g 0.0196061f $X=-0.19 $Y=1.655 $X2=0.675 $Y2=1.29
cc_110 VPB N_A_116_47#_M1014_g 0.0196061f $X=-0.19 $Y=1.655 $X2=0.675 $Y2=1.29
cc_111 VPB N_A_116_47#_M1015_g 0.0196061f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_112 VPB N_A_116_47#_M1016_g 0.0196061f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_113 VPB N_A_116_47#_M1017_g 0.0196061f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_114 VPB N_A_116_47#_M1019_g 0.0196061f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_115 VPB N_A_116_47#_M1022_g 0.0196058f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_116 VPB N_A_116_47#_M1028_g 0.0196338f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_117 VPB N_A_116_47#_M1032_g 0.0196061f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_118 VPB N_A_116_47#_M1034_g 0.0196061f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_119 VPB N_A_116_47#_M1037_g 0.0196061f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_120 VPB N_A_116_47#_M1038_g 0.0196061f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_121 VPB N_A_116_47#_M1039_g 0.0269266f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_122 VPB N_A_116_47#_c_308_n 0.00271941f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_123 VPB N_A_116_47#_c_309_n 0.00451764f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_124 VPB N_A_116_47#_c_310_n 0.00567517f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_125 VPB N_A_116_47#_c_281_n 5.66089e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_126 VPB N_A_116_47#_c_312_n 0.00226968f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_127 VPB N_VPWR_c_635_n 0.0118367f $X=-0.19 $Y=1.655 $X2=1.115 $Y2=1.21
cc_128 VPB N_VPWR_c_636_n 0.0502122f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_129 VPB N_VPWR_c_637_n 0.00403106f $X=-0.19 $Y=1.655 $X2=0.675 $Y2=1.29
cc_130 VPB N_VPWR_c_638_n 0.00408044f $X=-0.19 $Y=1.655 $X2=1.695 $Y2=1.29
cc_131 VPB N_VPWR_c_639_n 0.0135769f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_132 VPB N_VPWR_c_640_n 3.17051e-19 $X=-0.19 $Y=1.655 $X2=1.68 $Y2=1.29
cc_133 VPB N_VPWR_c_641_n 3.16188e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_134 VPB N_VPWR_c_642_n 3.16188e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_135 VPB N_VPWR_c_643_n 3.16188e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_136 VPB N_VPWR_c_644_n 3.17051e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_137 VPB N_VPWR_c_645_n 0.0135769f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_138 VPB N_VPWR_c_646_n 3.17051e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_139 VPB N_VPWR_c_647_n 3.16188e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_140 VPB N_VPWR_c_648_n 0.0121205f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_141 VPB N_VPWR_c_649_n 0.0511612f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_142 VPB N_VPWR_c_650_n 0.0134631f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_143 VPB N_VPWR_c_651_n 0.00410235f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_144 VPB N_VPWR_c_652_n 0.0134631f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_145 VPB N_VPWR_c_653_n 0.00403576f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_146 VPB N_VPWR_c_654_n 0.0167145f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_147 VPB N_VPWR_c_655_n 0.0163782f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_148 VPB N_VPWR_c_656_n 0.0134631f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_149 VPB N_VPWR_c_657_n 0.0134631f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_150 VPB N_VPWR_c_658_n 0.0134631f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_151 VPB N_VPWR_c_659_n 0.0134631f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_152 VPB N_VPWR_c_660_n 0.00507132f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_153 VPB N_VPWR_c_661_n 0.011737f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_154 VPB N_VPWR_c_662_n 0.00410235f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_155 VPB N_VPWR_c_663_n 0.00410235f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_156 VPB N_VPWR_c_664_n 0.00410235f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_157 VPB N_VPWR_c_665_n 0.00410235f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_158 VPB N_VPWR_c_666_n 0.00410235f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_159 VPB N_VPWR_c_634_n 0.0480432f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_160 VPB N_X_c_827_n 0.00396599f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_161 VPB N_X_c_828_n 0.00387487f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_162 VPB N_X_c_829_n 0.00387487f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_163 VPB N_X_c_830_n 0.00387487f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_164 VPB N_X_c_831_n 0.003869f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_165 VPB N_X_c_832_n 0.00389014f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_166 VPB N_X_c_833_n 0.00387487f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_167 VPB N_X_c_834_n 0.0040245f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_168 N_A_M1030_g N_A_116_47#_M1001_g 0.00600458f $X=1.795 $Y=0.445 $X2=0 $Y2=0
cc_169 N_A_M1035_g N_A_116_47#_M1000_g 0.00815828f $X=1.795 $Y=2.465 $X2=0 $Y2=0
cc_170 N_A_M1030_g N_A_116_47#_c_272_n 0.0346721f $X=1.795 $Y=0.445 $X2=0 $Y2=0
cc_171 A N_A_116_47#_c_272_n 2.98227e-19 $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_172 N_A_M1011_g N_A_116_47#_c_275_n 0.00328851f $X=0.505 $Y=0.445 $X2=0 $Y2=0
cc_173 N_A_M1026_g N_A_116_47#_c_275_n 0.00176083f $X=0.935 $Y=0.445 $X2=0 $Y2=0
cc_174 N_A_M1026_g N_A_116_47#_c_276_n 0.0114646f $X=0.935 $Y=0.445 $X2=0 $Y2=0
cc_175 N_A_M1029_g N_A_116_47#_c_276_n 0.0117609f $X=1.365 $Y=0.445 $X2=0 $Y2=0
cc_176 A N_A_116_47#_c_276_n 0.0434316f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_177 N_A_c_177_n N_A_116_47#_c_276_n 0.00222766f $X=1.795 $Y=1.29 $X2=0 $Y2=0
cc_178 N_A_M1011_g N_A_116_47#_c_277_n 0.00568793f $X=0.505 $Y=0.445 $X2=0 $Y2=0
cc_179 A N_A_116_47#_c_277_n 0.020161f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_180 N_A_c_177_n N_A_116_47#_c_277_n 0.00231242f $X=1.795 $Y=1.29 $X2=0 $Y2=0
cc_181 N_A_M1021_g N_A_116_47#_c_308_n 0.0149533f $X=0.935 $Y=2.465 $X2=0 $Y2=0
cc_182 N_A_M1025_g N_A_116_47#_c_308_n 0.0152312f $X=1.365 $Y=2.465 $X2=0 $Y2=0
cc_183 A N_A_116_47#_c_308_n 0.0350488f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_184 N_A_c_177_n N_A_116_47#_c_308_n 0.0021537f $X=1.795 $Y=1.29 $X2=0 $Y2=0
cc_185 N_A_M1004_g N_A_116_47#_c_309_n 0.00503628f $X=0.505 $Y=2.465 $X2=0 $Y2=0
cc_186 A N_A_116_47#_c_309_n 0.0178325f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_187 N_A_c_177_n N_A_116_47#_c_309_n 0.00225633f $X=1.795 $Y=1.29 $X2=0 $Y2=0
cc_188 N_A_M1029_g N_A_116_47#_c_278_n 0.0017555f $X=1.365 $Y=0.445 $X2=0 $Y2=0
cc_189 N_A_M1030_g N_A_116_47#_c_278_n 0.00325493f $X=1.795 $Y=0.445 $X2=0 $Y2=0
cc_190 N_A_M1030_g N_A_116_47#_c_279_n 0.0140837f $X=1.795 $Y=0.445 $X2=0 $Y2=0
cc_191 A N_A_116_47#_c_279_n 0.00752417f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_192 N_A_M1035_g N_A_116_47#_c_310_n 0.0176848f $X=1.795 $Y=2.465 $X2=0 $Y2=0
cc_193 A N_A_116_47#_c_310_n 0.00589724f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_194 N_A_M1030_g N_A_116_47#_c_280_n 0.00453701f $X=1.795 $Y=0.445 $X2=0 $Y2=0
cc_195 A N_A_116_47#_c_280_n 0.0247902f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_196 N_A_M1035_g N_A_116_47#_c_281_n 0.00453701f $X=1.795 $Y=2.465 $X2=0 $Y2=0
cc_197 A N_A_116_47#_c_282_n 0.0197577f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_198 N_A_c_177_n N_A_116_47#_c_282_n 0.00231242f $X=1.795 $Y=1.29 $X2=0 $Y2=0
cc_199 A N_A_116_47#_c_312_n 0.016823f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_200 N_A_c_177_n N_A_116_47#_c_312_n 0.00225633f $X=1.795 $Y=1.29 $X2=0 $Y2=0
cc_201 N_A_c_177_n N_A_116_47#_c_283_n 0.00453701f $X=1.795 $Y=1.29 $X2=0 $Y2=0
cc_202 A N_A_116_47#_c_290_n 0.00796421f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_203 N_A_c_177_n N_A_116_47#_c_290_n 0.00498172f $X=1.795 $Y=1.29 $X2=0 $Y2=0
cc_204 N_A_M1004_g N_VPWR_c_636_n 0.0050322f $X=0.505 $Y=2.465 $X2=0 $Y2=0
cc_205 N_A_M1021_g N_VPWR_c_637_n 0.00162181f $X=0.935 $Y=2.465 $X2=0 $Y2=0
cc_206 N_A_M1025_g N_VPWR_c_637_n 0.00162973f $X=1.365 $Y=2.465 $X2=0 $Y2=0
cc_207 N_A_M1035_g N_VPWR_c_638_n 0.00229987f $X=1.795 $Y=2.465 $X2=0 $Y2=0
cc_208 N_A_M1004_g N_VPWR_c_654_n 0.00585385f $X=0.505 $Y=2.465 $X2=0 $Y2=0
cc_209 N_A_M1021_g N_VPWR_c_654_n 0.00585385f $X=0.935 $Y=2.465 $X2=0 $Y2=0
cc_210 N_A_M1025_g N_VPWR_c_655_n 0.00583607f $X=1.365 $Y=2.465 $X2=0 $Y2=0
cc_211 N_A_M1035_g N_VPWR_c_655_n 0.00585385f $X=1.795 $Y=2.465 $X2=0 $Y2=0
cc_212 N_A_M1004_g N_VPWR_c_634_n 0.0116789f $X=0.505 $Y=2.465 $X2=0 $Y2=0
cc_213 N_A_M1021_g N_VPWR_c_634_n 0.0105977f $X=0.935 $Y=2.465 $X2=0 $Y2=0
cc_214 N_A_M1025_g N_VPWR_c_634_n 0.0105506f $X=1.365 $Y=2.465 $X2=0 $Y2=0
cc_215 N_A_M1035_g N_VPWR_c_634_n 0.0112877f $X=1.795 $Y=2.465 $X2=0 $Y2=0
cc_216 N_A_M1011_g N_VGND_c_1007_n 0.00370285f $X=0.505 $Y=0.445 $X2=0 $Y2=0
cc_217 N_A_M1026_g N_VGND_c_1008_n 0.00171697f $X=0.935 $Y=0.445 $X2=0 $Y2=0
cc_218 N_A_M1029_g N_VGND_c_1008_n 0.00170842f $X=1.365 $Y=0.445 $X2=0 $Y2=0
cc_219 N_A_M1011_g N_VGND_c_1024_n 0.00585385f $X=0.505 $Y=0.445 $X2=0 $Y2=0
cc_220 N_A_M1026_g N_VGND_c_1024_n 0.00583607f $X=0.935 $Y=0.445 $X2=0 $Y2=0
cc_221 N_A_M1029_g N_VGND_c_1030_n 0.00583607f $X=1.365 $Y=0.445 $X2=0 $Y2=0
cc_222 N_A_M1030_g N_VGND_c_1030_n 0.00585385f $X=1.795 $Y=0.445 $X2=0 $Y2=0
cc_223 N_A_M1030_g N_VGND_c_1031_n 0.00241256f $X=1.795 $Y=0.445 $X2=0 $Y2=0
cc_224 N_A_M1011_g N_VGND_c_1037_n 0.0117712f $X=0.505 $Y=0.445 $X2=0 $Y2=0
cc_225 N_A_M1026_g N_VGND_c_1037_n 0.00608505f $X=0.935 $Y=0.445 $X2=0 $Y2=0
cc_226 N_A_M1029_g N_VGND_c_1037_n 0.00608505f $X=1.365 $Y=0.445 $X2=0 $Y2=0
cc_227 N_A_M1030_g N_VGND_c_1037_n 0.00685381f $X=1.795 $Y=0.445 $X2=0 $Y2=0
cc_228 N_A_116_47#_c_308_n N_VPWR_M1021_d 0.00176461f $X=1.46 $Y=1.77 $X2=0
+ $Y2=0
cc_229 N_A_116_47#_c_310_n N_VPWR_M1035_d 0.00345375f $X=1.985 $Y=1.77 $X2=0
+ $Y2=0
cc_230 N_A_116_47#_c_308_n N_VPWR_c_637_n 0.0135055f $X=1.46 $Y=1.77 $X2=0 $Y2=0
cc_231 N_A_116_47#_M1000_g N_VPWR_c_638_n 0.0145089f $X=2.615 $Y=2.465 $X2=0
+ $Y2=0
cc_232 N_A_116_47#_M1002_g N_VPWR_c_638_n 7.6476e-19 $X=3.045 $Y=2.465 $X2=0
+ $Y2=0
cc_233 N_A_116_47#_c_272_n N_VPWR_c_638_n 0.00235812f $X=9.065 $Y=1.205 $X2=0
+ $Y2=0
cc_234 N_A_116_47#_c_310_n N_VPWR_c_638_n 0.0235837f $X=1.985 $Y=1.77 $X2=0
+ $Y2=0
cc_235 N_A_116_47#_c_283_n N_VPWR_c_638_n 0.0101191f $X=2.465 $Y=1.295 $X2=0
+ $Y2=0
cc_236 N_A_116_47#_c_290_n N_VPWR_c_638_n 0.0031131f $X=8.425 $Y=1.295 $X2=0
+ $Y2=0
cc_237 N_A_116_47#_M1000_g N_VPWR_c_639_n 0.00544582f $X=2.615 $Y=2.465 $X2=0
+ $Y2=0
cc_238 N_A_116_47#_M1002_g N_VPWR_c_639_n 0.00525069f $X=3.045 $Y=2.465 $X2=0
+ $Y2=0
cc_239 N_A_116_47#_M1000_g N_VPWR_c_640_n 8.84817e-19 $X=2.615 $Y=2.465 $X2=0
+ $Y2=0
cc_240 N_A_116_47#_M1002_g N_VPWR_c_640_n 0.0157287f $X=3.045 $Y=2.465 $X2=0
+ $Y2=0
cc_241 N_A_116_47#_M1010_g N_VPWR_c_640_n 0.0157158f $X=3.475 $Y=2.465 $X2=0
+ $Y2=0
cc_242 N_A_116_47#_M1013_g N_VPWR_c_640_n 8.8273e-19 $X=3.905 $Y=2.465 $X2=0
+ $Y2=0
cc_243 N_A_116_47#_c_272_n N_VPWR_c_640_n 7.24868e-19 $X=9.065 $Y=1.205 $X2=0
+ $Y2=0
cc_244 N_A_116_47#_c_284_n N_VPWR_c_640_n 0.00820577f $X=3.265 $Y=1.295 $X2=0
+ $Y2=0
cc_245 N_A_116_47#_c_290_n N_VPWR_c_640_n 0.00147571f $X=8.425 $Y=1.295 $X2=0
+ $Y2=0
cc_246 N_A_116_47#_M1010_g N_VPWR_c_641_n 8.8273e-19 $X=3.475 $Y=2.465 $X2=0
+ $Y2=0
cc_247 N_A_116_47#_M1013_g N_VPWR_c_641_n 0.0157158f $X=3.905 $Y=2.465 $X2=0
+ $Y2=0
cc_248 N_A_116_47#_M1014_g N_VPWR_c_641_n 0.0157158f $X=4.335 $Y=2.465 $X2=0
+ $Y2=0
cc_249 N_A_116_47#_M1015_g N_VPWR_c_641_n 8.8273e-19 $X=4.765 $Y=2.465 $X2=0
+ $Y2=0
cc_250 N_A_116_47#_c_272_n N_VPWR_c_641_n 7.24868e-19 $X=9.065 $Y=1.205 $X2=0
+ $Y2=0
cc_251 N_A_116_47#_c_285_n N_VPWR_c_641_n 0.00820577f $X=4.125 $Y=1.295 $X2=0
+ $Y2=0
cc_252 N_A_116_47#_c_290_n N_VPWR_c_641_n 0.00147571f $X=8.425 $Y=1.295 $X2=0
+ $Y2=0
cc_253 N_A_116_47#_M1014_g N_VPWR_c_642_n 8.8273e-19 $X=4.335 $Y=2.465 $X2=0
+ $Y2=0
cc_254 N_A_116_47#_M1015_g N_VPWR_c_642_n 0.0157158f $X=4.765 $Y=2.465 $X2=0
+ $Y2=0
cc_255 N_A_116_47#_M1016_g N_VPWR_c_642_n 0.0157158f $X=5.195 $Y=2.465 $X2=0
+ $Y2=0
cc_256 N_A_116_47#_M1017_g N_VPWR_c_642_n 8.8273e-19 $X=5.625 $Y=2.465 $X2=0
+ $Y2=0
cc_257 N_A_116_47#_c_272_n N_VPWR_c_642_n 7.24868e-19 $X=9.065 $Y=1.205 $X2=0
+ $Y2=0
cc_258 N_A_116_47#_c_286_n N_VPWR_c_642_n 0.00820577f $X=4.985 $Y=1.295 $X2=0
+ $Y2=0
cc_259 N_A_116_47#_c_290_n N_VPWR_c_642_n 0.00147571f $X=8.425 $Y=1.295 $X2=0
+ $Y2=0
cc_260 N_A_116_47#_M1016_g N_VPWR_c_643_n 8.8273e-19 $X=5.195 $Y=2.465 $X2=0
+ $Y2=0
cc_261 N_A_116_47#_M1017_g N_VPWR_c_643_n 0.0157158f $X=5.625 $Y=2.465 $X2=0
+ $Y2=0
cc_262 N_A_116_47#_M1019_g N_VPWR_c_643_n 0.0157158f $X=6.055 $Y=2.465 $X2=0
+ $Y2=0
cc_263 N_A_116_47#_M1022_g N_VPWR_c_643_n 8.8273e-19 $X=6.485 $Y=2.465 $X2=0
+ $Y2=0
cc_264 N_A_116_47#_c_272_n N_VPWR_c_643_n 7.24868e-19 $X=9.065 $Y=1.205 $X2=0
+ $Y2=0
cc_265 N_A_116_47#_c_287_n N_VPWR_c_643_n 0.00820577f $X=5.845 $Y=1.295 $X2=0
+ $Y2=0
cc_266 N_A_116_47#_c_290_n N_VPWR_c_643_n 0.00147571f $X=8.425 $Y=1.295 $X2=0
+ $Y2=0
cc_267 N_A_116_47#_M1019_g N_VPWR_c_644_n 8.82258e-19 $X=6.055 $Y=2.465 $X2=0
+ $Y2=0
cc_268 N_A_116_47#_M1022_g N_VPWR_c_644_n 0.0157158f $X=6.485 $Y=2.465 $X2=0
+ $Y2=0
cc_269 N_A_116_47#_M1028_g N_VPWR_c_644_n 0.0150735f $X=6.915 $Y=2.465 $X2=0
+ $Y2=0
cc_270 N_A_116_47#_M1032_g N_VPWR_c_644_n 8.7318e-19 $X=7.345 $Y=2.465 $X2=0
+ $Y2=0
cc_271 N_A_116_47#_c_272_n N_VPWR_c_644_n 7.24868e-19 $X=9.065 $Y=1.205 $X2=0
+ $Y2=0
cc_272 N_A_116_47#_c_288_n N_VPWR_c_644_n 0.00804519f $X=6.7 $Y=1.295 $X2=0
+ $Y2=0
cc_273 N_A_116_47#_c_290_n N_VPWR_c_644_n 0.00145491f $X=8.425 $Y=1.295 $X2=0
+ $Y2=0
cc_274 N_A_116_47#_M1028_g N_VPWR_c_645_n 0.00544582f $X=6.915 $Y=2.465 $X2=0
+ $Y2=0
cc_275 N_A_116_47#_M1032_g N_VPWR_c_645_n 0.00525069f $X=7.345 $Y=2.465 $X2=0
+ $Y2=0
cc_276 N_A_116_47#_M1028_g N_VPWR_c_646_n 8.84817e-19 $X=6.915 $Y=2.465 $X2=0
+ $Y2=0
cc_277 N_A_116_47#_M1032_g N_VPWR_c_646_n 0.0157287f $X=7.345 $Y=2.465 $X2=0
+ $Y2=0
cc_278 N_A_116_47#_M1034_g N_VPWR_c_646_n 0.0157158f $X=7.775 $Y=2.465 $X2=0
+ $Y2=0
cc_279 N_A_116_47#_M1037_g N_VPWR_c_646_n 8.8273e-19 $X=8.205 $Y=2.465 $X2=0
+ $Y2=0
cc_280 N_A_116_47#_c_272_n N_VPWR_c_646_n 7.24868e-19 $X=9.065 $Y=1.205 $X2=0
+ $Y2=0
cc_281 N_A_116_47#_c_289_n N_VPWR_c_646_n 0.00820577f $X=7.565 $Y=1.295 $X2=0
+ $Y2=0
cc_282 N_A_116_47#_c_290_n N_VPWR_c_646_n 0.00147571f $X=8.425 $Y=1.295 $X2=0
+ $Y2=0
cc_283 N_A_116_47#_M1034_g N_VPWR_c_647_n 8.8273e-19 $X=7.775 $Y=2.465 $X2=0
+ $Y2=0
cc_284 N_A_116_47#_M1037_g N_VPWR_c_647_n 0.0157158f $X=8.205 $Y=2.465 $X2=0
+ $Y2=0
cc_285 N_A_116_47#_M1038_g N_VPWR_c_647_n 0.0157158f $X=8.635 $Y=2.465 $X2=0
+ $Y2=0
cc_286 N_A_116_47#_c_272_n N_VPWR_c_647_n 7.24868e-19 $X=9.065 $Y=1.205 $X2=0
+ $Y2=0
cc_287 N_A_116_47#_M1039_g N_VPWR_c_647_n 8.8273e-19 $X=9.065 $Y=2.465 $X2=0
+ $Y2=0
cc_288 N_A_116_47#_c_290_n N_VPWR_c_647_n 0.00147571f $X=8.425 $Y=1.295 $X2=0
+ $Y2=0
cc_289 N_A_116_47#_c_291_n N_VPWR_c_647_n 0.00820577f $X=8.425 $Y=1.295 $X2=0
+ $Y2=0
cc_290 N_A_116_47#_M1038_g N_VPWR_c_649_n 8.01391e-19 $X=8.635 $Y=2.465 $X2=0
+ $Y2=0
cc_291 N_A_116_47#_M1039_g N_VPWR_c_649_n 0.0184839f $X=9.065 $Y=2.465 $X2=0
+ $Y2=0
cc_292 N_A_116_47#_M1016_g N_VPWR_c_650_n 0.00525069f $X=5.195 $Y=2.465 $X2=0
+ $Y2=0
cc_293 N_A_116_47#_M1017_g N_VPWR_c_650_n 0.00525069f $X=5.625 $Y=2.465 $X2=0
+ $Y2=0
cc_294 N_A_116_47#_M1019_g N_VPWR_c_652_n 0.00525069f $X=6.055 $Y=2.465 $X2=0
+ $Y2=0
cc_295 N_A_116_47#_M1022_g N_VPWR_c_652_n 0.00525069f $X=6.485 $Y=2.465 $X2=0
+ $Y2=0
cc_296 N_A_116_47#_c_417_p N_VPWR_c_654_n 0.0151136f $X=0.72 $Y=2.04 $X2=0 $Y2=0
cc_297 N_A_116_47#_c_418_p N_VPWR_c_655_n 0.0145813f $X=1.58 $Y=2.04 $X2=0 $Y2=0
cc_298 N_A_116_47#_M1010_g N_VPWR_c_656_n 0.00525069f $X=3.475 $Y=2.465 $X2=0
+ $Y2=0
cc_299 N_A_116_47#_M1013_g N_VPWR_c_656_n 0.00525069f $X=3.905 $Y=2.465 $X2=0
+ $Y2=0
cc_300 N_A_116_47#_M1014_g N_VPWR_c_657_n 0.00525069f $X=4.335 $Y=2.465 $X2=0
+ $Y2=0
cc_301 N_A_116_47#_M1015_g N_VPWR_c_657_n 0.00525069f $X=4.765 $Y=2.465 $X2=0
+ $Y2=0
cc_302 N_A_116_47#_M1034_g N_VPWR_c_658_n 0.00525069f $X=7.775 $Y=2.465 $X2=0
+ $Y2=0
cc_303 N_A_116_47#_M1037_g N_VPWR_c_658_n 0.00525069f $X=8.205 $Y=2.465 $X2=0
+ $Y2=0
cc_304 N_A_116_47#_M1038_g N_VPWR_c_659_n 0.00525069f $X=8.635 $Y=2.465 $X2=0
+ $Y2=0
cc_305 N_A_116_47#_M1039_g N_VPWR_c_659_n 0.00525069f $X=9.065 $Y=2.465 $X2=0
+ $Y2=0
cc_306 N_A_116_47#_M1004_s N_VPWR_c_634_n 0.0027574f $X=0.58 $Y=1.835 $X2=0
+ $Y2=0
cc_307 N_A_116_47#_M1025_s N_VPWR_c_634_n 0.00327921f $X=1.44 $Y=1.835 $X2=0
+ $Y2=0
cc_308 N_A_116_47#_M1000_g N_VPWR_c_634_n 0.00923564f $X=2.615 $Y=2.465 $X2=0
+ $Y2=0
cc_309 N_A_116_47#_M1002_g N_VPWR_c_634_n 0.00892673f $X=3.045 $Y=2.465 $X2=0
+ $Y2=0
cc_310 N_A_116_47#_M1010_g N_VPWR_c_634_n 0.00892673f $X=3.475 $Y=2.465 $X2=0
+ $Y2=0
cc_311 N_A_116_47#_M1013_g N_VPWR_c_634_n 0.00892673f $X=3.905 $Y=2.465 $X2=0
+ $Y2=0
cc_312 N_A_116_47#_M1014_g N_VPWR_c_634_n 0.00892673f $X=4.335 $Y=2.465 $X2=0
+ $Y2=0
cc_313 N_A_116_47#_M1015_g N_VPWR_c_634_n 0.00892673f $X=4.765 $Y=2.465 $X2=0
+ $Y2=0
cc_314 N_A_116_47#_M1016_g N_VPWR_c_634_n 0.00892673f $X=5.195 $Y=2.465 $X2=0
+ $Y2=0
cc_315 N_A_116_47#_M1017_g N_VPWR_c_634_n 0.00892673f $X=5.625 $Y=2.465 $X2=0
+ $Y2=0
cc_316 N_A_116_47#_M1019_g N_VPWR_c_634_n 0.00892673f $X=6.055 $Y=2.465 $X2=0
+ $Y2=0
cc_317 N_A_116_47#_M1022_g N_VPWR_c_634_n 0.00892673f $X=6.485 $Y=2.465 $X2=0
+ $Y2=0
cc_318 N_A_116_47#_M1028_g N_VPWR_c_634_n 0.00923564f $X=6.915 $Y=2.465 $X2=0
+ $Y2=0
cc_319 N_A_116_47#_M1032_g N_VPWR_c_634_n 0.00892673f $X=7.345 $Y=2.465 $X2=0
+ $Y2=0
cc_320 N_A_116_47#_M1034_g N_VPWR_c_634_n 0.00892673f $X=7.775 $Y=2.465 $X2=0
+ $Y2=0
cc_321 N_A_116_47#_M1037_g N_VPWR_c_634_n 0.00892673f $X=8.205 $Y=2.465 $X2=0
+ $Y2=0
cc_322 N_A_116_47#_M1038_g N_VPWR_c_634_n 0.00892673f $X=8.635 $Y=2.465 $X2=0
+ $Y2=0
cc_323 N_A_116_47#_M1039_g N_VPWR_c_634_n 0.00892673f $X=9.065 $Y=2.465 $X2=0
+ $Y2=0
cc_324 N_A_116_47#_c_417_p N_VPWR_c_634_n 0.0102248f $X=0.72 $Y=2.04 $X2=0 $Y2=0
cc_325 N_A_116_47#_c_418_p N_VPWR_c_634_n 0.00964167f $X=1.58 $Y=2.04 $X2=0
+ $Y2=0
cc_326 N_A_116_47#_M1001_g N_X_c_827_n 0.00691693f $X=2.615 $Y=0.445 $X2=0 $Y2=0
cc_327 N_A_116_47#_M1000_g N_X_c_827_n 0.00519941f $X=2.615 $Y=2.465 $X2=0 $Y2=0
cc_328 N_A_116_47#_M1003_g N_X_c_827_n 0.00767605f $X=3.045 $Y=0.445 $X2=0 $Y2=0
cc_329 N_A_116_47#_M1002_g N_X_c_827_n 0.00478785f $X=3.045 $Y=2.465 $X2=0 $Y2=0
cc_330 N_A_116_47#_c_272_n N_X_c_827_n 0.0179156f $X=9.065 $Y=1.205 $X2=0 $Y2=0
cc_331 N_A_116_47#_c_279_n N_X_c_827_n 0.013775f $X=1.985 $Y=0.86 $X2=0 $Y2=0
cc_332 N_A_116_47#_c_310_n N_X_c_827_n 0.0062498f $X=1.985 $Y=1.77 $X2=0 $Y2=0
cc_333 N_A_116_47#_c_280_n N_X_c_827_n 0.0432521f $X=2.28 $Y=1.03 $X2=0 $Y2=0
cc_334 N_A_116_47#_c_281_n N_X_c_827_n 0.00532075f $X=2.092 $Y=1.685 $X2=0 $Y2=0
cc_335 N_A_116_47#_c_284_n N_X_c_827_n 0.0224022f $X=3.265 $Y=1.295 $X2=0 $Y2=0
cc_336 N_A_116_47#_c_290_n N_X_c_827_n 0.027968f $X=8.425 $Y=1.295 $X2=0 $Y2=0
cc_337 N_A_116_47#_M1005_g N_X_c_828_n 0.00761263f $X=3.475 $Y=0.445 $X2=0 $Y2=0
cc_338 N_A_116_47#_M1010_g N_X_c_828_n 0.0047717f $X=3.475 $Y=2.465 $X2=0 $Y2=0
cc_339 N_A_116_47#_M1006_g N_X_c_828_n 0.00761263f $X=3.905 $Y=0.445 $X2=0 $Y2=0
cc_340 N_A_116_47#_M1013_g N_X_c_828_n 0.0047717f $X=3.905 $Y=2.465 $X2=0 $Y2=0
cc_341 N_A_116_47#_c_272_n N_X_c_828_n 0.0179348f $X=9.065 $Y=1.205 $X2=0 $Y2=0
cc_342 N_A_116_47#_c_284_n N_X_c_828_n 0.0223699f $X=3.265 $Y=1.295 $X2=0 $Y2=0
cc_343 N_A_116_47#_c_285_n N_X_c_828_n 0.0223699f $X=4.125 $Y=1.295 $X2=0 $Y2=0
cc_344 N_A_116_47#_c_290_n N_X_c_828_n 0.0277981f $X=8.425 $Y=1.295 $X2=0 $Y2=0
cc_345 N_A_116_47#_M1007_g N_X_c_829_n 0.00761263f $X=4.335 $Y=0.445 $X2=0 $Y2=0
cc_346 N_A_116_47#_M1014_g N_X_c_829_n 0.0047717f $X=4.335 $Y=2.465 $X2=0 $Y2=0
cc_347 N_A_116_47#_M1008_g N_X_c_829_n 0.00761263f $X=4.765 $Y=0.445 $X2=0 $Y2=0
cc_348 N_A_116_47#_M1015_g N_X_c_829_n 0.0047717f $X=4.765 $Y=2.465 $X2=0 $Y2=0
cc_349 N_A_116_47#_c_272_n N_X_c_829_n 0.0179348f $X=9.065 $Y=1.205 $X2=0 $Y2=0
cc_350 N_A_116_47#_c_285_n N_X_c_829_n 0.0223699f $X=4.125 $Y=1.295 $X2=0 $Y2=0
cc_351 N_A_116_47#_c_286_n N_X_c_829_n 0.0223699f $X=4.985 $Y=1.295 $X2=0 $Y2=0
cc_352 N_A_116_47#_c_290_n N_X_c_829_n 0.0277981f $X=8.425 $Y=1.295 $X2=0 $Y2=0
cc_353 N_A_116_47#_M1009_g N_X_c_830_n 0.00761263f $X=5.195 $Y=0.445 $X2=0 $Y2=0
cc_354 N_A_116_47#_M1016_g N_X_c_830_n 0.0047717f $X=5.195 $Y=2.465 $X2=0 $Y2=0
cc_355 N_A_116_47#_M1012_g N_X_c_830_n 0.00761263f $X=5.625 $Y=0.445 $X2=0 $Y2=0
cc_356 N_A_116_47#_M1017_g N_X_c_830_n 0.0047717f $X=5.625 $Y=2.465 $X2=0 $Y2=0
cc_357 N_A_116_47#_c_272_n N_X_c_830_n 0.0179348f $X=9.065 $Y=1.205 $X2=0 $Y2=0
cc_358 N_A_116_47#_c_286_n N_X_c_830_n 0.0223699f $X=4.985 $Y=1.295 $X2=0 $Y2=0
cc_359 N_A_116_47#_c_287_n N_X_c_830_n 0.0223699f $X=5.845 $Y=1.295 $X2=0 $Y2=0
cc_360 N_A_116_47#_c_290_n N_X_c_830_n 0.0277981f $X=8.425 $Y=1.295 $X2=0 $Y2=0
cc_361 N_A_116_47#_M1018_g N_X_c_831_n 0.00761263f $X=6.055 $Y=0.445 $X2=0 $Y2=0
cc_362 N_A_116_47#_M1019_g N_X_c_831_n 0.0047717f $X=6.055 $Y=2.465 $X2=0 $Y2=0
cc_363 N_A_116_47#_M1020_g N_X_c_831_n 0.00758371f $X=6.485 $Y=0.445 $X2=0 $Y2=0
cc_364 N_A_116_47#_M1022_g N_X_c_831_n 0.00475583f $X=6.485 $Y=2.465 $X2=0 $Y2=0
cc_365 N_A_116_47#_c_272_n N_X_c_831_n 0.0179348f $X=9.065 $Y=1.205 $X2=0 $Y2=0
cc_366 N_A_116_47#_c_287_n N_X_c_831_n 0.0223699f $X=5.845 $Y=1.295 $X2=0 $Y2=0
cc_367 N_A_116_47#_c_288_n N_X_c_831_n 0.0223575f $X=6.7 $Y=1.295 $X2=0 $Y2=0
cc_368 N_A_116_47#_c_290_n N_X_c_831_n 0.0277956f $X=8.425 $Y=1.295 $X2=0 $Y2=0
cc_369 N_A_116_47#_M1023_g N_X_c_832_n 0.00768787f $X=6.915 $Y=0.445 $X2=0 $Y2=0
cc_370 N_A_116_47#_M1028_g N_X_c_832_n 0.00482092f $X=6.915 $Y=2.465 $X2=0 $Y2=0
cc_371 N_A_116_47#_M1024_g N_X_c_832_n 0.00764f $X=7.345 $Y=0.445 $X2=0 $Y2=0
cc_372 N_A_116_47#_M1032_g N_X_c_832_n 0.00478785f $X=7.345 $Y=2.465 $X2=0 $Y2=0
cc_373 N_A_116_47#_c_272_n N_X_c_832_n 0.0180935f $X=9.065 $Y=1.205 $X2=0 $Y2=0
cc_374 N_A_116_47#_c_288_n N_X_c_832_n 0.0223746f $X=6.7 $Y=1.295 $X2=0 $Y2=0
cc_375 N_A_116_47#_c_289_n N_X_c_832_n 0.0223871f $X=7.565 $Y=1.295 $X2=0 $Y2=0
cc_376 N_A_116_47#_c_290_n N_X_c_832_n 0.0283445f $X=8.425 $Y=1.295 $X2=0 $Y2=0
cc_377 N_A_116_47#_M1027_g N_X_c_833_n 0.00761263f $X=7.775 $Y=0.445 $X2=0 $Y2=0
cc_378 N_A_116_47#_M1034_g N_X_c_833_n 0.0047717f $X=7.775 $Y=2.465 $X2=0 $Y2=0
cc_379 N_A_116_47#_M1031_g N_X_c_833_n 0.00761263f $X=8.205 $Y=0.445 $X2=0 $Y2=0
cc_380 N_A_116_47#_M1037_g N_X_c_833_n 0.0047717f $X=8.205 $Y=2.465 $X2=0 $Y2=0
cc_381 N_A_116_47#_c_272_n N_X_c_833_n 0.0179348f $X=9.065 $Y=1.205 $X2=0 $Y2=0
cc_382 N_A_116_47#_c_289_n N_X_c_833_n 0.0223699f $X=7.565 $Y=1.295 $X2=0 $Y2=0
cc_383 N_A_116_47#_c_290_n N_X_c_833_n 0.0277707f $X=8.425 $Y=1.295 $X2=0 $Y2=0
cc_384 N_A_116_47#_c_291_n N_X_c_833_n 0.0223699f $X=8.425 $Y=1.295 $X2=0 $Y2=0
cc_385 N_A_116_47#_M1033_g N_X_c_834_n 0.00766326f $X=8.635 $Y=0.445 $X2=0 $Y2=0
cc_386 N_A_116_47#_M1038_g N_X_c_834_n 0.0047717f $X=8.635 $Y=2.465 $X2=0 $Y2=0
cc_387 N_A_116_47#_c_272_n N_X_c_834_n 0.0289495f $X=9.065 $Y=1.205 $X2=0 $Y2=0
cc_388 N_A_116_47#_M1036_g N_X_c_834_n 0.0140794f $X=9.065 $Y=0.445 $X2=0 $Y2=0
cc_389 N_A_116_47#_M1039_g N_X_c_834_n 0.00826608f $X=9.065 $Y=2.465 $X2=0 $Y2=0
cc_390 N_A_116_47#_c_290_n N_X_c_834_n 0.00708764f $X=8.425 $Y=1.295 $X2=0 $Y2=0
cc_391 N_A_116_47#_c_291_n N_X_c_834_n 0.021437f $X=8.425 $Y=1.295 $X2=0 $Y2=0
cc_392 N_A_116_47#_M1000_g N_X_c_909_n 0.00525656f $X=2.615 $Y=2.465 $X2=0 $Y2=0
cc_393 N_A_116_47#_M1002_g N_X_c_909_n 0.00798792f $X=3.045 $Y=2.465 $X2=0 $Y2=0
cc_394 N_A_116_47#_M1010_g N_X_c_909_n 0.00798792f $X=3.475 $Y=2.465 $X2=0 $Y2=0
cc_395 N_A_116_47#_M1013_g N_X_c_909_n 0.00798792f $X=3.905 $Y=2.465 $X2=0 $Y2=0
cc_396 N_A_116_47#_M1014_g N_X_c_909_n 0.00798792f $X=4.335 $Y=2.465 $X2=0 $Y2=0
cc_397 N_A_116_47#_M1015_g N_X_c_909_n 0.00798792f $X=4.765 $Y=2.465 $X2=0 $Y2=0
cc_398 N_A_116_47#_M1016_g N_X_c_909_n 0.00798792f $X=5.195 $Y=2.465 $X2=0 $Y2=0
cc_399 N_A_116_47#_M1017_g N_X_c_909_n 0.00798792f $X=5.625 $Y=2.465 $X2=0 $Y2=0
cc_400 N_A_116_47#_M1019_g N_X_c_909_n 0.00798792f $X=6.055 $Y=2.465 $X2=0 $Y2=0
cc_401 N_A_116_47#_M1022_g N_X_c_909_n 0.00798792f $X=6.485 $Y=2.465 $X2=0 $Y2=0
cc_402 N_A_116_47#_M1028_g N_X_c_909_n 0.00828377f $X=6.915 $Y=2.465 $X2=0 $Y2=0
cc_403 N_A_116_47#_M1032_g N_X_c_909_n 0.00798792f $X=7.345 $Y=2.465 $X2=0 $Y2=0
cc_404 N_A_116_47#_M1034_g N_X_c_909_n 0.00798792f $X=7.775 $Y=2.465 $X2=0 $Y2=0
cc_405 N_A_116_47#_M1037_g N_X_c_909_n 0.00798792f $X=8.205 $Y=2.465 $X2=0 $Y2=0
cc_406 N_A_116_47#_M1038_g N_X_c_909_n 0.0106488f $X=8.635 $Y=2.465 $X2=0 $Y2=0
cc_407 N_A_116_47#_M1039_g N_X_c_909_n 0.00564645f $X=9.065 $Y=2.465 $X2=0 $Y2=0
cc_408 N_A_116_47#_c_284_n N_X_c_909_n 0.00130876f $X=3.265 $Y=1.295 $X2=0 $Y2=0
cc_409 N_A_116_47#_c_285_n N_X_c_909_n 0.00130876f $X=4.125 $Y=1.295 $X2=0 $Y2=0
cc_410 N_A_116_47#_c_286_n N_X_c_909_n 0.00130876f $X=4.985 $Y=1.295 $X2=0 $Y2=0
cc_411 N_A_116_47#_c_287_n N_X_c_909_n 0.00130876f $X=5.845 $Y=1.295 $X2=0 $Y2=0
cc_412 N_A_116_47#_c_288_n N_X_c_909_n 0.00128751f $X=6.7 $Y=1.295 $X2=0 $Y2=0
cc_413 N_A_116_47#_c_289_n N_X_c_909_n 0.00130876f $X=7.565 $Y=1.295 $X2=0 $Y2=0
cc_414 N_A_116_47#_c_290_n N_X_c_909_n 0.269372f $X=8.425 $Y=1.295 $X2=0 $Y2=0
cc_415 N_A_116_47#_c_291_n N_X_c_909_n 0.00130876f $X=8.425 $Y=1.295 $X2=0 $Y2=0
cc_416 N_A_116_47#_c_276_n N_VGND_c_1008_n 0.017321f $X=1.46 $Y=0.86 $X2=0 $Y2=0
cc_417 N_A_116_47#_M1001_g N_VGND_c_1009_n 0.00544582f $X=2.615 $Y=0.445 $X2=0
+ $Y2=0
cc_418 N_A_116_47#_M1003_g N_VGND_c_1009_n 0.00525069f $X=3.045 $Y=0.445 $X2=0
+ $Y2=0
cc_419 N_A_116_47#_M1001_g N_VGND_c_1010_n 5.68147e-19 $X=2.615 $Y=0.445 $X2=0
+ $Y2=0
cc_420 N_A_116_47#_M1003_g N_VGND_c_1010_n 0.00769543f $X=3.045 $Y=0.445 $X2=0
+ $Y2=0
cc_421 N_A_116_47#_M1005_g N_VGND_c_1010_n 0.00769334f $X=3.475 $Y=0.445 $X2=0
+ $Y2=0
cc_422 N_A_116_47#_M1006_g N_VGND_c_1010_n 5.66477e-19 $X=3.905 $Y=0.445 $X2=0
+ $Y2=0
cc_423 N_A_116_47#_c_272_n N_VGND_c_1010_n 6.26773e-19 $X=9.065 $Y=1.205 $X2=0
+ $Y2=0
cc_424 N_A_116_47#_c_284_n N_VGND_c_1010_n 0.00353566f $X=3.265 $Y=1.295 $X2=0
+ $Y2=0
cc_425 N_A_116_47#_c_290_n N_VGND_c_1010_n 0.00684837f $X=8.425 $Y=1.295 $X2=0
+ $Y2=0
cc_426 N_A_116_47#_M1005_g N_VGND_c_1011_n 5.66477e-19 $X=3.475 $Y=0.445 $X2=0
+ $Y2=0
cc_427 N_A_116_47#_M1006_g N_VGND_c_1011_n 0.00769334f $X=3.905 $Y=0.445 $X2=0
+ $Y2=0
cc_428 N_A_116_47#_M1007_g N_VGND_c_1011_n 0.00769334f $X=4.335 $Y=0.445 $X2=0
+ $Y2=0
cc_429 N_A_116_47#_M1008_g N_VGND_c_1011_n 5.66477e-19 $X=4.765 $Y=0.445 $X2=0
+ $Y2=0
cc_430 N_A_116_47#_c_272_n N_VGND_c_1011_n 6.26773e-19 $X=9.065 $Y=1.205 $X2=0
+ $Y2=0
cc_431 N_A_116_47#_c_285_n N_VGND_c_1011_n 0.00353566f $X=4.125 $Y=1.295 $X2=0
+ $Y2=0
cc_432 N_A_116_47#_c_290_n N_VGND_c_1011_n 0.00684837f $X=8.425 $Y=1.295 $X2=0
+ $Y2=0
cc_433 N_A_116_47#_M1007_g N_VGND_c_1012_n 5.66477e-19 $X=4.335 $Y=0.445 $X2=0
+ $Y2=0
cc_434 N_A_116_47#_M1008_g N_VGND_c_1012_n 0.00769334f $X=4.765 $Y=0.445 $X2=0
+ $Y2=0
cc_435 N_A_116_47#_M1009_g N_VGND_c_1012_n 0.00769334f $X=5.195 $Y=0.445 $X2=0
+ $Y2=0
cc_436 N_A_116_47#_M1012_g N_VGND_c_1012_n 5.66477e-19 $X=5.625 $Y=0.445 $X2=0
+ $Y2=0
cc_437 N_A_116_47#_c_272_n N_VGND_c_1012_n 6.26773e-19 $X=9.065 $Y=1.205 $X2=0
+ $Y2=0
cc_438 N_A_116_47#_c_286_n N_VGND_c_1012_n 0.00353566f $X=4.985 $Y=1.295 $X2=0
+ $Y2=0
cc_439 N_A_116_47#_c_290_n N_VGND_c_1012_n 0.00684837f $X=8.425 $Y=1.295 $X2=0
+ $Y2=0
cc_440 N_A_116_47#_M1009_g N_VGND_c_1013_n 5.66477e-19 $X=5.195 $Y=0.445 $X2=0
+ $Y2=0
cc_441 N_A_116_47#_M1012_g N_VGND_c_1013_n 0.00769334f $X=5.625 $Y=0.445 $X2=0
+ $Y2=0
cc_442 N_A_116_47#_M1018_g N_VGND_c_1013_n 0.00769334f $X=6.055 $Y=0.445 $X2=0
+ $Y2=0
cc_443 N_A_116_47#_M1020_g N_VGND_c_1013_n 5.66477e-19 $X=6.485 $Y=0.445 $X2=0
+ $Y2=0
cc_444 N_A_116_47#_c_272_n N_VGND_c_1013_n 6.26773e-19 $X=9.065 $Y=1.205 $X2=0
+ $Y2=0
cc_445 N_A_116_47#_c_287_n N_VGND_c_1013_n 0.00353566f $X=5.845 $Y=1.295 $X2=0
+ $Y2=0
cc_446 N_A_116_47#_c_290_n N_VGND_c_1013_n 0.00684837f $X=8.425 $Y=1.295 $X2=0
+ $Y2=0
cc_447 N_A_116_47#_M1018_g N_VGND_c_1014_n 5.6615e-19 $X=6.055 $Y=0.445 $X2=0
+ $Y2=0
cc_448 N_A_116_47#_M1020_g N_VGND_c_1014_n 0.00769334f $X=6.485 $Y=0.445 $X2=0
+ $Y2=0
cc_449 N_A_116_47#_M1023_g N_VGND_c_1014_n 0.00729875f $X=6.915 $Y=0.445 $X2=0
+ $Y2=0
cc_450 N_A_116_47#_M1024_g N_VGND_c_1014_n 5.61169e-19 $X=7.345 $Y=0.445 $X2=0
+ $Y2=0
cc_451 N_A_116_47#_c_272_n N_VGND_c_1014_n 6.26773e-19 $X=9.065 $Y=1.205 $X2=0
+ $Y2=0
cc_452 N_A_116_47#_c_288_n N_VGND_c_1014_n 0.00346643f $X=6.7 $Y=1.295 $X2=0
+ $Y2=0
cc_453 N_A_116_47#_c_290_n N_VGND_c_1014_n 0.00675797f $X=8.425 $Y=1.295 $X2=0
+ $Y2=0
cc_454 N_A_116_47#_M1023_g N_VGND_c_1015_n 0.00544582f $X=6.915 $Y=0.445 $X2=0
+ $Y2=0
cc_455 N_A_116_47#_M1024_g N_VGND_c_1015_n 0.00525069f $X=7.345 $Y=0.445 $X2=0
+ $Y2=0
cc_456 N_A_116_47#_M1023_g N_VGND_c_1016_n 5.68564e-19 $X=6.915 $Y=0.445 $X2=0
+ $Y2=0
cc_457 N_A_116_47#_M1024_g N_VGND_c_1016_n 0.00770619f $X=7.345 $Y=0.445 $X2=0
+ $Y2=0
cc_458 N_A_116_47#_M1027_g N_VGND_c_1016_n 0.00769334f $X=7.775 $Y=0.445 $X2=0
+ $Y2=0
cc_459 N_A_116_47#_M1031_g N_VGND_c_1016_n 5.66477e-19 $X=8.205 $Y=0.445 $X2=0
+ $Y2=0
cc_460 N_A_116_47#_c_272_n N_VGND_c_1016_n 6.26773e-19 $X=9.065 $Y=1.205 $X2=0
+ $Y2=0
cc_461 N_A_116_47#_c_289_n N_VGND_c_1016_n 0.00353566f $X=7.565 $Y=1.295 $X2=0
+ $Y2=0
cc_462 N_A_116_47#_c_290_n N_VGND_c_1016_n 0.00684837f $X=8.425 $Y=1.295 $X2=0
+ $Y2=0
cc_463 N_A_116_47#_M1027_g N_VGND_c_1017_n 5.66477e-19 $X=7.775 $Y=0.445 $X2=0
+ $Y2=0
cc_464 N_A_116_47#_M1031_g N_VGND_c_1017_n 0.00769334f $X=8.205 $Y=0.445 $X2=0
+ $Y2=0
cc_465 N_A_116_47#_M1033_g N_VGND_c_1017_n 0.00769334f $X=8.635 $Y=0.445 $X2=0
+ $Y2=0
cc_466 N_A_116_47#_c_272_n N_VGND_c_1017_n 6.26773e-19 $X=9.065 $Y=1.205 $X2=0
+ $Y2=0
cc_467 N_A_116_47#_M1036_g N_VGND_c_1017_n 5.66477e-19 $X=9.065 $Y=0.445 $X2=0
+ $Y2=0
cc_468 N_A_116_47#_c_290_n N_VGND_c_1017_n 0.00684837f $X=8.425 $Y=1.295 $X2=0
+ $Y2=0
cc_469 N_A_116_47#_c_291_n N_VGND_c_1017_n 0.00353566f $X=8.425 $Y=1.295 $X2=0
+ $Y2=0
cc_470 N_A_116_47#_M1033_g N_VGND_c_1019_n 5.67119e-19 $X=8.635 $Y=0.445 $X2=0
+ $Y2=0
cc_471 N_A_116_47#_M1036_g N_VGND_c_1019_n 0.00915342f $X=9.065 $Y=0.445 $X2=0
+ $Y2=0
cc_472 N_A_116_47#_M1009_g N_VGND_c_1020_n 0.00525069f $X=5.195 $Y=0.445 $X2=0
+ $Y2=0
cc_473 N_A_116_47#_M1012_g N_VGND_c_1020_n 0.00525069f $X=5.625 $Y=0.445 $X2=0
+ $Y2=0
cc_474 N_A_116_47#_M1018_g N_VGND_c_1022_n 0.00525069f $X=6.055 $Y=0.445 $X2=0
+ $Y2=0
cc_475 N_A_116_47#_M1020_g N_VGND_c_1022_n 0.00525069f $X=6.485 $Y=0.445 $X2=0
+ $Y2=0
cc_476 N_A_116_47#_c_275_n N_VGND_c_1024_n 0.0125732f $X=0.72 $Y=0.445 $X2=0
+ $Y2=0
cc_477 N_A_116_47#_M1005_g N_VGND_c_1025_n 0.00525069f $X=3.475 $Y=0.445 $X2=0
+ $Y2=0
cc_478 N_A_116_47#_M1006_g N_VGND_c_1025_n 0.00525069f $X=3.905 $Y=0.445 $X2=0
+ $Y2=0
cc_479 N_A_116_47#_M1007_g N_VGND_c_1026_n 0.00525069f $X=4.335 $Y=0.445 $X2=0
+ $Y2=0
cc_480 N_A_116_47#_M1008_g N_VGND_c_1026_n 0.00525069f $X=4.765 $Y=0.445 $X2=0
+ $Y2=0
cc_481 N_A_116_47#_M1027_g N_VGND_c_1027_n 0.00525069f $X=7.775 $Y=0.445 $X2=0
+ $Y2=0
cc_482 N_A_116_47#_M1031_g N_VGND_c_1027_n 0.00525069f $X=8.205 $Y=0.445 $X2=0
+ $Y2=0
cc_483 N_A_116_47#_M1033_g N_VGND_c_1028_n 0.00525069f $X=8.635 $Y=0.445 $X2=0
+ $Y2=0
cc_484 N_A_116_47#_M1036_g N_VGND_c_1028_n 0.00525069f $X=9.065 $Y=0.445 $X2=0
+ $Y2=0
cc_485 N_A_116_47#_c_278_n N_VGND_c_1030_n 0.0124184f $X=1.58 $Y=0.445 $X2=0
+ $Y2=0
cc_486 N_A_116_47#_M1001_g N_VGND_c_1031_n 0.00837538f $X=2.615 $Y=0.445 $X2=0
+ $Y2=0
cc_487 N_A_116_47#_M1003_g N_VGND_c_1031_n 5.78376e-19 $X=3.045 $Y=0.445 $X2=0
+ $Y2=0
cc_488 N_A_116_47#_c_272_n N_VGND_c_1031_n 0.00249081f $X=9.065 $Y=1.205 $X2=0
+ $Y2=0
cc_489 N_A_116_47#_c_279_n N_VGND_c_1031_n 0.0526157f $X=1.985 $Y=0.86 $X2=0
+ $Y2=0
cc_490 N_A_116_47#_c_290_n N_VGND_c_1031_n 0.00223347f $X=8.425 $Y=1.295 $X2=0
+ $Y2=0
cc_491 N_A_116_47#_M1011_d N_VGND_c_1037_n 0.00274817f $X=0.58 $Y=0.235 $X2=0
+ $Y2=0
cc_492 N_A_116_47#_M1029_d N_VGND_c_1037_n 0.00244217f $X=1.44 $Y=0.235 $X2=0
+ $Y2=0
cc_493 N_A_116_47#_M1001_g N_VGND_c_1037_n 0.00918681f $X=2.615 $Y=0.445 $X2=0
+ $Y2=0
cc_494 N_A_116_47#_M1003_g N_VGND_c_1037_n 0.00892673f $X=3.045 $Y=0.445 $X2=0
+ $Y2=0
cc_495 N_A_116_47#_M1005_g N_VGND_c_1037_n 0.00892673f $X=3.475 $Y=0.445 $X2=0
+ $Y2=0
cc_496 N_A_116_47#_M1006_g N_VGND_c_1037_n 0.00892673f $X=3.905 $Y=0.445 $X2=0
+ $Y2=0
cc_497 N_A_116_47#_M1007_g N_VGND_c_1037_n 0.00892673f $X=4.335 $Y=0.445 $X2=0
+ $Y2=0
cc_498 N_A_116_47#_M1008_g N_VGND_c_1037_n 0.00892673f $X=4.765 $Y=0.445 $X2=0
+ $Y2=0
cc_499 N_A_116_47#_M1009_g N_VGND_c_1037_n 0.00892673f $X=5.195 $Y=0.445 $X2=0
+ $Y2=0
cc_500 N_A_116_47#_M1012_g N_VGND_c_1037_n 0.00892673f $X=5.625 $Y=0.445 $X2=0
+ $Y2=0
cc_501 N_A_116_47#_M1018_g N_VGND_c_1037_n 0.00892673f $X=6.055 $Y=0.445 $X2=0
+ $Y2=0
cc_502 N_A_116_47#_M1020_g N_VGND_c_1037_n 0.00892673f $X=6.485 $Y=0.445 $X2=0
+ $Y2=0
cc_503 N_A_116_47#_M1023_g N_VGND_c_1037_n 0.00923564f $X=6.915 $Y=0.445 $X2=0
+ $Y2=0
cc_504 N_A_116_47#_M1024_g N_VGND_c_1037_n 0.00892673f $X=7.345 $Y=0.445 $X2=0
+ $Y2=0
cc_505 N_A_116_47#_M1027_g N_VGND_c_1037_n 0.00892673f $X=7.775 $Y=0.445 $X2=0
+ $Y2=0
cc_506 N_A_116_47#_M1031_g N_VGND_c_1037_n 0.00892673f $X=8.205 $Y=0.445 $X2=0
+ $Y2=0
cc_507 N_A_116_47#_M1033_g N_VGND_c_1037_n 0.00892673f $X=8.635 $Y=0.445 $X2=0
+ $Y2=0
cc_508 N_A_116_47#_M1036_g N_VGND_c_1037_n 0.00892673f $X=9.065 $Y=0.445 $X2=0
+ $Y2=0
cc_509 N_A_116_47#_c_275_n N_VGND_c_1037_n 0.00951847f $X=0.72 $Y=0.445 $X2=0
+ $Y2=0
cc_510 N_A_116_47#_c_276_n N_VGND_c_1037_n 0.0112116f $X=1.46 $Y=0.86 $X2=0
+ $Y2=0
cc_511 N_A_116_47#_c_278_n N_VGND_c_1037_n 0.00932657f $X=1.58 $Y=0.445 $X2=0
+ $Y2=0
cc_512 N_A_116_47#_c_279_n N_VGND_c_1037_n 0.00771845f $X=1.985 $Y=0.86 $X2=0
+ $Y2=0
cc_513 N_VPWR_c_634_n N_X_M1000_s 0.00450209f $X=9.36 $Y=3.33 $X2=0 $Y2=0
cc_514 N_VPWR_c_634_n N_X_M1010_s 0.00467591f $X=9.36 $Y=3.33 $X2=0 $Y2=0
cc_515 N_VPWR_c_634_n N_X_M1014_s 0.00467591f $X=9.36 $Y=3.33 $X2=0 $Y2=0
cc_516 N_VPWR_c_634_n N_X_M1016_s 0.00467591f $X=9.36 $Y=3.33 $X2=0 $Y2=0
cc_517 N_VPWR_c_634_n N_X_M1019_s 0.00467591f $X=9.36 $Y=3.33 $X2=0 $Y2=0
cc_518 N_VPWR_c_634_n N_X_M1028_s 0.00450209f $X=9.36 $Y=3.33 $X2=0 $Y2=0
cc_519 N_VPWR_c_634_n N_X_M1034_s 0.00467591f $X=9.36 $Y=3.33 $X2=0 $Y2=0
cc_520 N_VPWR_c_634_n N_X_M1038_s 0.00467591f $X=9.36 $Y=3.33 $X2=0 $Y2=0
cc_521 N_VPWR_c_638_n N_X_c_827_n 0.0442334f $X=2.01 $Y=2.19 $X2=0 $Y2=0
cc_522 N_VPWR_c_639_n N_X_c_827_n 0.0118321f $X=3.105 $Y=3.33 $X2=0 $Y2=0
cc_523 N_VPWR_c_640_n N_X_c_827_n 0.0468931f $X=3.26 $Y=2.04 $X2=0 $Y2=0
cc_524 N_VPWR_c_634_n N_X_c_827_n 0.00820109f $X=9.36 $Y=3.33 $X2=0 $Y2=0
cc_525 N_VPWR_c_640_n N_X_c_828_n 0.04689f $X=3.26 $Y=2.04 $X2=0 $Y2=0
cc_526 N_VPWR_c_641_n N_X_c_828_n 0.04689f $X=4.12 $Y=2.04 $X2=0 $Y2=0
cc_527 N_VPWR_c_656_n N_X_c_828_n 0.0116733f $X=3.965 $Y=3.33 $X2=0 $Y2=0
cc_528 N_VPWR_c_634_n N_X_c_828_n 0.00800858f $X=9.36 $Y=3.33 $X2=0 $Y2=0
cc_529 N_VPWR_c_641_n N_X_c_829_n 0.04689f $X=4.12 $Y=2.04 $X2=0 $Y2=0
cc_530 N_VPWR_c_642_n N_X_c_829_n 0.04689f $X=4.98 $Y=2.04 $X2=0 $Y2=0
cc_531 N_VPWR_c_657_n N_X_c_829_n 0.0116733f $X=4.825 $Y=3.33 $X2=0 $Y2=0
cc_532 N_VPWR_c_634_n N_X_c_829_n 0.00800858f $X=9.36 $Y=3.33 $X2=0 $Y2=0
cc_533 N_VPWR_c_642_n N_X_c_830_n 0.04689f $X=4.98 $Y=2.04 $X2=0 $Y2=0
cc_534 N_VPWR_c_643_n N_X_c_830_n 0.04689f $X=5.84 $Y=2.04 $X2=0 $Y2=0
cc_535 N_VPWR_c_650_n N_X_c_830_n 0.0116733f $X=5.685 $Y=3.33 $X2=0 $Y2=0
cc_536 N_VPWR_c_634_n N_X_c_830_n 0.00800858f $X=9.36 $Y=3.33 $X2=0 $Y2=0
cc_537 N_VPWR_c_643_n N_X_c_831_n 0.04689f $X=5.84 $Y=2.04 $X2=0 $Y2=0
cc_538 N_VPWR_c_644_n N_X_c_831_n 0.0468012f $X=6.7 $Y=2.04 $X2=0 $Y2=0
cc_539 N_VPWR_c_652_n N_X_c_831_n 0.0116733f $X=6.545 $Y=3.33 $X2=0 $Y2=0
cc_540 N_VPWR_c_634_n N_X_c_831_n 0.00800858f $X=9.36 $Y=3.33 $X2=0 $Y2=0
cc_541 N_VPWR_c_644_n N_X_c_832_n 0.0468042f $X=6.7 $Y=2.04 $X2=0 $Y2=0
cc_542 N_VPWR_c_645_n N_X_c_832_n 0.0118321f $X=7.405 $Y=3.33 $X2=0 $Y2=0
cc_543 N_VPWR_c_646_n N_X_c_832_n 0.0468931f $X=7.56 $Y=2.04 $X2=0 $Y2=0
cc_544 N_VPWR_c_634_n N_X_c_832_n 0.00820109f $X=9.36 $Y=3.33 $X2=0 $Y2=0
cc_545 N_VPWR_c_646_n N_X_c_833_n 0.04689f $X=7.56 $Y=2.04 $X2=0 $Y2=0
cc_546 N_VPWR_c_647_n N_X_c_833_n 0.04689f $X=8.42 $Y=2.04 $X2=0 $Y2=0
cc_547 N_VPWR_c_658_n N_X_c_833_n 0.0116733f $X=8.265 $Y=3.33 $X2=0 $Y2=0
cc_548 N_VPWR_c_634_n N_X_c_833_n 0.00800858f $X=9.36 $Y=3.33 $X2=0 $Y2=0
cc_549 N_VPWR_c_647_n N_X_c_834_n 0.04689f $X=8.42 $Y=2.04 $X2=0 $Y2=0
cc_550 N_VPWR_c_649_n N_X_c_834_n 0.0463091f $X=9.28 $Y=2.04 $X2=0 $Y2=0
cc_551 N_VPWR_c_659_n N_X_c_834_n 0.0116733f $X=9.125 $Y=3.33 $X2=0 $Y2=0
cc_552 N_VPWR_c_634_n N_X_c_834_n 0.00800858f $X=9.36 $Y=3.33 $X2=0 $Y2=0
cc_553 N_VPWR_c_638_n N_X_c_909_n 0.00386445f $X=2.01 $Y=2.19 $X2=0 $Y2=0
cc_554 N_VPWR_c_640_n N_X_c_909_n 0.0339375f $X=3.26 $Y=2.04 $X2=0 $Y2=0
cc_555 N_VPWR_c_641_n N_X_c_909_n 0.0339375f $X=4.12 $Y=2.04 $X2=0 $Y2=0
cc_556 N_VPWR_c_642_n N_X_c_909_n 0.0339375f $X=4.98 $Y=2.04 $X2=0 $Y2=0
cc_557 N_VPWR_c_643_n N_X_c_909_n 0.0339375f $X=5.84 $Y=2.04 $X2=0 $Y2=0
cc_558 N_VPWR_c_644_n N_X_c_909_n 0.0334539f $X=6.7 $Y=2.04 $X2=0 $Y2=0
cc_559 N_VPWR_c_646_n N_X_c_909_n 0.0339375f $X=7.56 $Y=2.04 $X2=0 $Y2=0
cc_560 N_VPWR_c_647_n N_X_c_909_n 0.0339375f $X=8.42 $Y=2.04 $X2=0 $Y2=0
cc_561 N_VPWR_c_649_n N_X_c_909_n 0.0074036f $X=9.28 $Y=2.04 $X2=0 $Y2=0
cc_562 N_X_c_827_n N_VGND_c_1009_n 0.0118321f $X=2.83 $Y=0.44 $X2=0 $Y2=0
cc_563 N_X_c_832_n N_VGND_c_1015_n 0.0118321f $X=7.13 $Y=0.44 $X2=0 $Y2=0
cc_564 N_X_c_830_n N_VGND_c_1020_n 0.0116733f $X=5.41 $Y=0.44 $X2=0 $Y2=0
cc_565 N_X_c_831_n N_VGND_c_1022_n 0.0116733f $X=6.27 $Y=0.44 $X2=0 $Y2=0
cc_566 N_X_c_828_n N_VGND_c_1025_n 0.0116733f $X=3.69 $Y=0.44 $X2=0 $Y2=0
cc_567 N_X_c_829_n N_VGND_c_1026_n 0.0116733f $X=4.55 $Y=0.44 $X2=0 $Y2=0
cc_568 N_X_c_833_n N_VGND_c_1027_n 0.0116733f $X=7.99 $Y=0.44 $X2=0 $Y2=0
cc_569 N_X_c_834_n N_VGND_c_1028_n 0.0116733f $X=8.85 $Y=0.44 $X2=0 $Y2=0
cc_570 N_X_M1001_s N_VGND_c_1037_n 0.00450209f $X=2.69 $Y=0.235 $X2=0 $Y2=0
cc_571 N_X_M1005_s N_VGND_c_1037_n 0.00467591f $X=3.55 $Y=0.235 $X2=0 $Y2=0
cc_572 N_X_M1007_s N_VGND_c_1037_n 0.00467591f $X=4.41 $Y=0.235 $X2=0 $Y2=0
cc_573 N_X_M1009_s N_VGND_c_1037_n 0.00467591f $X=5.27 $Y=0.235 $X2=0 $Y2=0
cc_574 N_X_M1018_s N_VGND_c_1037_n 0.00467591f $X=6.13 $Y=0.235 $X2=0 $Y2=0
cc_575 N_X_M1023_s N_VGND_c_1037_n 0.00450209f $X=6.99 $Y=0.235 $X2=0 $Y2=0
cc_576 N_X_M1027_s N_VGND_c_1037_n 0.00467591f $X=7.85 $Y=0.235 $X2=0 $Y2=0
cc_577 N_X_M1033_s N_VGND_c_1037_n 0.00467591f $X=8.71 $Y=0.235 $X2=0 $Y2=0
cc_578 N_X_c_827_n N_VGND_c_1037_n 0.00820109f $X=2.83 $Y=0.44 $X2=0 $Y2=0
cc_579 N_X_c_828_n N_VGND_c_1037_n 0.00800858f $X=3.69 $Y=0.44 $X2=0 $Y2=0
cc_580 N_X_c_829_n N_VGND_c_1037_n 0.00800858f $X=4.55 $Y=0.44 $X2=0 $Y2=0
cc_581 N_X_c_830_n N_VGND_c_1037_n 0.00800858f $X=5.41 $Y=0.44 $X2=0 $Y2=0
cc_582 N_X_c_831_n N_VGND_c_1037_n 0.00800858f $X=6.27 $Y=0.44 $X2=0 $Y2=0
cc_583 N_X_c_832_n N_VGND_c_1037_n 0.00820109f $X=7.13 $Y=0.44 $X2=0 $Y2=0
cc_584 N_X_c_833_n N_VGND_c_1037_n 0.00800858f $X=7.99 $Y=0.44 $X2=0 $Y2=0
cc_585 N_X_c_834_n N_VGND_c_1037_n 0.00800858f $X=8.85 $Y=0.44 $X2=0 $Y2=0
