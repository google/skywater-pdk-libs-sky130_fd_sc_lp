* File: sky130_fd_sc_lp__dlclkp_lp.pxi.spice
* Created: Wed Sep  2 09:46:01 2020
* 
x_PM_SKY130_FD_SC_LP__DLCLKP_LP%A_80_21# N_A_80_21#_M1016_s N_A_80_21#_M1020_s
+ N_A_80_21#_M1013_g N_A_80_21#_M1003_g N_A_80_21#_M1000_g N_A_80_21#_M1010_g
+ N_A_80_21#_M1012_g N_A_80_21#_c_139_n N_A_80_21#_c_140_n N_A_80_21#_c_141_n
+ N_A_80_21#_c_150_n N_A_80_21#_c_142_n N_A_80_21#_c_143_n N_A_80_21#_c_158_p
+ N_A_80_21#_c_144_n N_A_80_21#_c_145_n N_A_80_21#_c_146_n N_A_80_21#_c_154_n
+ N_A_80_21#_c_155_n PM_SKY130_FD_SC_LP__DLCLKP_LP%A_80_21#
x_PM_SKY130_FD_SC_LP__DLCLKP_LP%GATE N_GATE_M1007_g N_GATE_c_285_n
+ N_GATE_M1009_g N_GATE_c_286_n GATE N_GATE_c_287_n N_GATE_c_288_n
+ N_GATE_c_289_n PM_SKY130_FD_SC_LP__DLCLKP_LP%GATE
x_PM_SKY130_FD_SC_LP__DLCLKP_LP%A_27_47# N_A_27_47#_M1013_s N_A_27_47#_M1003_s
+ N_A_27_47#_M1018_g N_A_27_47#_c_342_n N_A_27_47#_c_343_n N_A_27_47#_c_333_n
+ N_A_27_47#_c_334_n N_A_27_47#_c_335_n N_A_27_47#_M1022_g N_A_27_47#_c_336_n
+ N_A_27_47#_c_337_n N_A_27_47#_c_338_n N_A_27_47#_c_345_n N_A_27_47#_c_339_n
+ N_A_27_47#_c_340_n PM_SKY130_FD_SC_LP__DLCLKP_LP%A_27_47#
x_PM_SKY130_FD_SC_LP__DLCLKP_LP%A_584_21# N_A_584_21#_M1023_d
+ N_A_584_21#_M1015_d N_A_584_21#_M1011_g N_A_584_21#_M1001_g
+ N_A_584_21#_c_423_n N_A_584_21#_M1005_g N_A_584_21#_M1004_g
+ N_A_584_21#_c_424_n N_A_584_21#_c_425_n N_A_584_21#_c_426_n
+ N_A_584_21#_c_427_n N_A_584_21#_c_428_n N_A_584_21#_c_438_n
+ N_A_584_21#_c_439_n N_A_584_21#_c_440_n N_A_584_21#_c_429_n
+ N_A_584_21#_c_430_n N_A_584_21#_c_431_n N_A_584_21#_c_444_n
+ N_A_584_21#_c_432_n N_A_584_21#_c_433_n
+ PM_SKY130_FD_SC_LP__DLCLKP_LP%A_584_21#
x_PM_SKY130_FD_SC_LP__DLCLKP_LP%A_352_419# N_A_352_419#_M1010_d
+ N_A_352_419#_M1018_d N_A_352_419#_M1019_g N_A_352_419#_M1015_g
+ N_A_352_419#_M1023_g N_A_352_419#_c_598_n N_A_352_419#_c_591_n
+ N_A_352_419#_c_584_n N_A_352_419#_c_585_n N_A_352_419#_c_586_n
+ N_A_352_419#_c_592_n N_A_352_419#_c_593_n N_A_352_419#_c_587_n
+ N_A_352_419#_c_588_n N_A_352_419#_c_589_n
+ PM_SKY130_FD_SC_LP__DLCLKP_LP%A_352_419#
x_PM_SKY130_FD_SC_LP__DLCLKP_LP%CLK N_CLK_c_688_n N_CLK_M1016_g N_CLK_c_689_n
+ N_CLK_c_690_n N_CLK_c_691_n N_CLK_M1014_g N_CLK_M1020_g N_CLK_c_692_n
+ N_CLK_M1017_g N_CLK_M1008_g CLK N_CLK_c_694_n
+ PM_SKY130_FD_SC_LP__DLCLKP_LP%CLK
x_PM_SKY130_FD_SC_LP__DLCLKP_LP%A_1147_419# N_A_1147_419#_M1005_d
+ N_A_1147_419#_M1008_d N_A_1147_419#_M1002_g N_A_1147_419#_M1021_g
+ N_A_1147_419#_M1006_g N_A_1147_419#_c_743_n N_A_1147_419#_c_744_n
+ N_A_1147_419#_c_759_n N_A_1147_419#_c_745_n N_A_1147_419#_c_746_n
+ N_A_1147_419#_c_763_n N_A_1147_419#_c_747_n N_A_1147_419#_c_768_n
+ N_A_1147_419#_c_748_n N_A_1147_419#_c_749_n N_A_1147_419#_c_775_n
+ PM_SKY130_FD_SC_LP__DLCLKP_LP%A_1147_419#
x_PM_SKY130_FD_SC_LP__DLCLKP_LP%VPWR N_VPWR_M1003_d N_VPWR_M1001_d
+ N_VPWR_M1020_d N_VPWR_M1004_d N_VPWR_c_811_n N_VPWR_c_812_n N_VPWR_c_813_n
+ N_VPWR_c_814_n N_VPWR_c_815_n N_VPWR_c_816_n N_VPWR_c_817_n N_VPWR_c_818_n
+ VPWR N_VPWR_c_819_n N_VPWR_c_820_n N_VPWR_c_810_n N_VPWR_c_822_n
+ N_VPWR_c_823_n PM_SKY130_FD_SC_LP__DLCLKP_LP%VPWR
x_PM_SKY130_FD_SC_LP__DLCLKP_LP%GCLK N_GCLK_M1006_d N_GCLK_M1021_d
+ N_GCLK_c_896_n GCLK GCLK GCLK N_GCLK_c_897_n GCLK
+ PM_SKY130_FD_SC_LP__DLCLKP_LP%GCLK
x_PM_SKY130_FD_SC_LP__DLCLKP_LP%VGND N_VGND_M1000_d N_VGND_M1011_d
+ N_VGND_M1014_d N_VGND_M1002_s N_VGND_c_919_n N_VGND_c_920_n N_VGND_c_921_n
+ N_VGND_c_922_n N_VGND_c_923_n N_VGND_c_924_n N_VGND_c_925_n N_VGND_c_926_n
+ VGND N_VGND_c_927_n N_VGND_c_928_n N_VGND_c_929_n N_VGND_c_930_n
+ N_VGND_c_931_n N_VGND_c_932_n PM_SKY130_FD_SC_LP__DLCLKP_LP%VGND
cc_1 VNB N_A_80_21#_M1013_g 0.036286f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.445
cc_2 VNB N_A_80_21#_M1003_g 0.0186852f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=2.595
cc_3 VNB N_A_80_21#_M1000_g 0.0281975f $X=-0.19 $Y=-0.245 $X2=0.835 $Y2=0.445
cc_4 VNB N_A_80_21#_M1010_g 0.0331082f $X=-0.19 $Y=-0.245 $X2=1.735 $Y2=0.445
cc_5 VNB N_A_80_21#_c_139_n 0.0141149f $X=-0.19 $Y=-0.245 $X2=1.48 $Y2=1.23
cc_6 VNB N_A_80_21#_c_140_n 0.0370858f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.23
cc_7 VNB N_A_80_21#_c_141_n 0.0117478f $X=-0.19 $Y=-0.245 $X2=1.725 $Y2=1.78
cc_8 VNB N_A_80_21#_c_142_n 0.00645722f $X=-0.19 $Y=-0.245 $X2=2.545 $Y2=1.615
cc_9 VNB N_A_80_21#_c_143_n 0.0251433f $X=-0.19 $Y=-0.245 $X2=2.545 $Y2=1.615
cc_10 VNB N_A_80_21#_c_144_n 0.0073279f $X=-0.19 $Y=-0.245 $X2=4.405 $Y2=2.315
cc_11 VNB N_A_80_21#_c_145_n 0.0277522f $X=-0.19 $Y=-0.245 $X2=1.645 $Y2=1.285
cc_12 VNB N_A_80_21#_c_146_n 0.00588765f $X=-0.19 $Y=-0.245 $X2=4.325 $Y2=1.06
cc_13 VNB N_GATE_c_285_n 0.0148981f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.065
cc_14 VNB N_GATE_c_286_n 0.0165759f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=2.595
cc_15 VNB N_GATE_c_287_n 0.00838345f $X=-0.19 $Y=-0.245 $X2=0.835 $Y2=0.445
cc_16 VNB N_GATE_c_288_n 0.00243064f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_GATE_c_289_n 0.036624f $X=-0.19 $Y=-0.245 $X2=1.735 $Y2=1.12
cc_18 VNB N_A_27_47#_c_333_n 0.0400976f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=2.595
cc_19 VNB N_A_27_47#_c_334_n 0.0382449f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_27_47#_c_335_n 0.0187157f $X=-0.19 $Y=-0.245 $X2=0.835 $Y2=1.065
cc_21 VNB N_A_27_47#_c_336_n 0.0178557f $X=-0.19 $Y=-0.245 $X2=1.735 $Y2=0.445
cc_22 VNB N_A_27_47#_c_337_n 0.0229559f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_27_47#_c_338_n 0.0131464f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.23
cc_24 VNB N_A_27_47#_c_339_n 0.0368319f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_27_47#_c_340_n 0.00489305f $X=-0.19 $Y=-0.245 $X2=1.725 $Y2=1.78
cc_26 VNB N_A_584_21#_M1011_g 0.0585295f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.445
cc_27 VNB N_A_584_21#_c_423_n 0.0177893f $X=-0.19 $Y=-0.245 $X2=0.835 $Y2=1.065
cc_28 VNB N_A_584_21#_c_424_n 0.0079402f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_584_21#_c_425_n 0.0134323f $X=-0.19 $Y=-0.245 $X2=2.505 $Y2=2.595
cc_30 VNB N_A_584_21#_c_426_n 0.0100624f $X=-0.19 $Y=-0.245 $X2=1.48 $Y2=1.23
cc_31 VNB N_A_584_21#_c_427_n 0.0186155f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.23
cc_32 VNB N_A_584_21#_c_428_n 0.0160906f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_584_21#_c_429_n 0.0370501f $X=-0.19 $Y=-0.245 $X2=2.545 $Y2=1.615
cc_34 VNB N_A_584_21#_c_430_n 0.0018159f $X=-0.19 $Y=-0.245 $X2=4.32 $Y2=2.6
cc_35 VNB N_A_584_21#_c_431_n 0.0253693f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_584_21#_c_432_n 0.013384f $X=-0.19 $Y=-0.245 $X2=4.405 $Y2=2.5
cc_37 VNB N_A_584_21#_c_433_n 0.00885582f $X=-0.19 $Y=-0.245 $X2=4.815 $Y2=2.5
cc_38 VNB N_A_352_419#_M1019_g 0.0182992f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.445
cc_39 VNB N_A_352_419#_M1023_g 0.0224802f $X=-0.19 $Y=-0.245 $X2=1.735 $Y2=1.12
cc_40 VNB N_A_352_419#_c_584_n 0.00363255f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.23
cc_41 VNB N_A_352_419#_c_585_n 0.00750859f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_352_419#_c_586_n 0.0119505f $X=-0.19 $Y=-0.245 $X2=1.725 $Y2=2.515
cc_43 VNB N_A_352_419#_c_587_n 0.00913096f $X=-0.19 $Y=-0.245 $X2=4.405
+ $Y2=2.315
cc_44 VNB N_A_352_419#_c_588_n 0.0427738f $X=-0.19 $Y=-0.245 $X2=1.645 $Y2=1.285
cc_45 VNB N_A_352_419#_c_589_n 0.0273979f $X=-0.19 $Y=-0.245 $X2=1.645 $Y2=1.615
cc_46 VNB N_CLK_c_688_n 0.0186823f $X=-0.19 $Y=-0.245 $X2=4.18 $Y2=0.925
cc_47 VNB N_CLK_c_689_n 0.0202608f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_CLK_c_690_n 0.0142894f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_CLK_c_691_n 0.0179093f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_CLK_c_692_n 0.01758f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=2.595
cc_51 VNB CLK 0.00637682f $X=-0.19 $Y=-0.245 $X2=1.735 $Y2=0.445
cc_52 VNB N_CLK_c_694_n 0.0344081f $X=-0.19 $Y=-0.245 $X2=1.48 $Y2=1.23
cc_53 VNB N_A_1147_419#_M1002_g 0.0281873f $X=-0.19 $Y=-0.245 $X2=0.475
+ $Y2=0.445
cc_54 VNB N_A_1147_419#_M1021_g 0.004948f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=2.595
cc_55 VNB N_A_1147_419#_M1006_g 0.0260781f $X=-0.19 $Y=-0.245 $X2=0.835
+ $Y2=0.445
cc_56 VNB N_A_1147_419#_c_743_n 0.0226787f $X=-0.19 $Y=-0.245 $X2=2.505 $Y2=1.78
cc_57 VNB N_A_1147_419#_c_744_n 0.0153384f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_1147_419#_c_745_n 0.0086528f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_1147_419#_c_746_n 0.00122182f $X=-0.19 $Y=-0.245 $X2=1.725
+ $Y2=2.515
cc_60 VNB N_A_1147_419#_c_747_n 7.1295e-19 $X=-0.19 $Y=-0.245 $X2=2.545
+ $Y2=1.615
cc_61 VNB N_A_1147_419#_c_748_n 0.00883638f $X=-0.19 $Y=-0.245 $X2=4.32 $Y2=2.6
cc_62 VNB N_A_1147_419#_c_749_n 0.0305946f $X=-0.19 $Y=-0.245 $X2=1.645
+ $Y2=1.285
cc_63 VNB N_VPWR_c_810_n 0.302998f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.23
cc_64 VNB N_GCLK_c_896_n 0.0216665f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_GCLK_c_897_n 0.0463558f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.23
cc_66 VNB N_VGND_c_919_n 0.002833f $X=-0.19 $Y=-0.245 $X2=0.835 $Y2=1.065
cc_67 VNB N_VGND_c_920_n 0.0458922f $X=-0.19 $Y=-0.245 $X2=0.835 $Y2=0.445
cc_68 VNB N_VGND_c_921_n 4.89148e-19 $X=-0.19 $Y=-0.245 $X2=1.735 $Y2=0.445
cc_69 VNB N_VGND_c_922_n 0.0328503f $X=-0.19 $Y=-0.245 $X2=2.505 $Y2=2.595
cc_70 VNB N_VGND_c_923_n 0.0180749f $X=-0.19 $Y=-0.245 $X2=1.48 $Y2=1.23
cc_71 VNB N_VGND_c_924_n 0.0117334f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_VGND_c_925_n 0.0454109f $X=-0.19 $Y=-0.245 $X2=1.725 $Y2=2.515
cc_73 VNB N_VGND_c_926_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=1.81 $Y2=1.615
cc_74 VNB N_VGND_c_927_n 0.0244814f $X=-0.19 $Y=-0.245 $X2=2.545 $Y2=1.615
cc_75 VNB N_VGND_c_928_n 0.0266387f $X=-0.19 $Y=-0.245 $X2=4.325 $Y2=1.06
cc_76 VNB N_VGND_c_929_n 0.379127f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_VGND_c_930_n 0.0051053f $X=-0.19 $Y=-0.245 $X2=4.32 $Y2=2.5
cc_78 VNB N_VGND_c_931_n 0.00437061f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_VGND_c_932_n 0.00513431f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.23
cc_80 VPB N_A_80_21#_M1003_g 0.0458207f $X=-0.19 $Y=1.655 $X2=0.575 $Y2=2.595
cc_81 VPB N_A_80_21#_M1012_g 0.0402315f $X=-0.19 $Y=1.655 $X2=2.505 $Y2=2.595
cc_82 VPB N_A_80_21#_c_141_n 3.15809e-19 $X=-0.19 $Y=1.655 $X2=1.725 $Y2=1.78
cc_83 VPB N_A_80_21#_c_150_n 0.003375f $X=-0.19 $Y=1.655 $X2=1.725 $Y2=2.515
cc_84 VPB N_A_80_21#_c_142_n 0.00357971f $X=-0.19 $Y=1.655 $X2=2.545 $Y2=1.615
cc_85 VPB N_A_80_21#_c_143_n 0.0090953f $X=-0.19 $Y=1.655 $X2=2.545 $Y2=1.615
cc_86 VPB N_A_80_21#_c_144_n 0.00968892f $X=-0.19 $Y=1.655 $X2=4.405 $Y2=2.315
cc_87 VPB N_A_80_21#_c_154_n 0.0110109f $X=-0.19 $Y=1.655 $X2=4.32 $Y2=2.5
cc_88 VPB N_A_80_21#_c_155_n 0.034039f $X=-0.19 $Y=1.655 $X2=4.815 $Y2=2.48
cc_89 VPB N_GATE_M1007_g 0.0239114f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_90 VPB N_GATE_c_287_n 0.0191834f $X=-0.19 $Y=1.655 $X2=0.835 $Y2=0.445
cc_91 VPB N_GATE_c_288_n 0.00382f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_92 VPB N_A_27_47#_M1018_g 0.0335546f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.445
cc_93 VPB N_A_27_47#_c_342_n 0.0275712f $X=-0.19 $Y=1.655 $X2=0.575 $Y2=1.395
cc_94 VPB N_A_27_47#_c_343_n 0.0104708f $X=-0.19 $Y=1.655 $X2=0.575 $Y2=2.595
cc_95 VPB N_A_27_47#_c_334_n 0.00186175f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_96 VPB N_A_27_47#_c_345_n 0.0302161f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=1.23
cc_97 VPB N_A_27_47#_c_339_n 0.0301675f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_98 VPB N_A_584_21#_M1001_g 0.0408934f $X=-0.19 $Y=1.655 $X2=0.575 $Y2=2.595
cc_99 VPB N_A_584_21#_M1004_g 0.0268772f $X=-0.19 $Y=1.655 $X2=1.735 $Y2=0.445
cc_100 VPB N_A_584_21#_c_426_n 0.00492808f $X=-0.19 $Y=1.655 $X2=1.48 $Y2=1.23
cc_101 VPB N_A_584_21#_c_428_n 0.00106255f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_102 VPB N_A_584_21#_c_438_n 0.00736909f $X=-0.19 $Y=1.655 $X2=1.725 $Y2=1.78
cc_103 VPB N_A_584_21#_c_439_n 0.00213271f $X=-0.19 $Y=1.655 $X2=1.725 $Y2=2.515
cc_104 VPB N_A_584_21#_c_440_n 0.00156239f $X=-0.19 $Y=1.655 $X2=2.545 $Y2=1.615
cc_105 VPB N_A_584_21#_c_429_n 0.0166419f $X=-0.19 $Y=1.655 $X2=2.545 $Y2=1.615
cc_106 VPB N_A_584_21#_c_430_n 9.80967e-19 $X=-0.19 $Y=1.655 $X2=4.32 $Y2=2.6
cc_107 VPB N_A_584_21#_c_431_n 0.00632394f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_108 VPB N_A_584_21#_c_444_n 0.00260452f $X=-0.19 $Y=1.655 $X2=1.645 $Y2=1.285
cc_109 VPB N_A_352_419#_M1015_g 0.0289865f $X=-0.19 $Y=1.655 $X2=0.835 $Y2=1.065
cc_110 VPB N_A_352_419#_c_591_n 0.0151101f $X=-0.19 $Y=1.655 $X2=2.505 $Y2=2.595
cc_111 VPB N_A_352_419#_c_592_n 0.00147816f $X=-0.19 $Y=1.655 $X2=2.545
+ $Y2=1.615
cc_112 VPB N_A_352_419#_c_593_n 0.00295875f $X=-0.19 $Y=1.655 $X2=4.405
+ $Y2=1.145
cc_113 VPB N_A_352_419#_c_587_n 0.0232233f $X=-0.19 $Y=1.655 $X2=4.405 $Y2=2.315
cc_114 VPB N_CLK_M1020_g 0.0268804f $X=-0.19 $Y=1.655 $X2=0.575 $Y2=1.395
cc_115 VPB N_CLK_M1008_g 0.0222335f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_116 VPB CLK 0.00148588f $X=-0.19 $Y=1.655 $X2=1.735 $Y2=0.445
cc_117 VPB N_CLK_c_694_n 0.031505f $X=-0.19 $Y=1.655 $X2=1.48 $Y2=1.23
cc_118 VPB N_A_1147_419#_M1021_g 0.0453963f $X=-0.19 $Y=1.655 $X2=0.575
+ $Y2=2.595
cc_119 VPB N_A_1147_419#_c_747_n 0.00268785f $X=-0.19 $Y=1.655 $X2=2.545
+ $Y2=1.615
cc_120 VPB N_VPWR_c_811_n 0.00283153f $X=-0.19 $Y=1.655 $X2=0.835 $Y2=0.445
cc_121 VPB N_VPWR_c_812_n 0.00286019f $X=-0.19 $Y=1.655 $X2=1.735 $Y2=0.445
cc_122 VPB N_VPWR_c_813_n 4.89148e-19 $X=-0.19 $Y=1.655 $X2=2.505 $Y2=2.595
cc_123 VPB N_VPWR_c_814_n 4.89148e-19 $X=-0.19 $Y=1.655 $X2=0.61 $Y2=1.23
cc_124 VPB N_VPWR_c_815_n 0.0613979f $X=-0.19 $Y=1.655 $X2=1.725 $Y2=1.78
cc_125 VPB N_VPWR_c_816_n 0.00513086f $X=-0.19 $Y=1.655 $X2=1.725 $Y2=2.515
cc_126 VPB N_VPWR_c_817_n 0.0440282f $X=-0.19 $Y=1.655 $X2=2.545 $Y2=1.615
cc_127 VPB N_VPWR_c_818_n 0.00436868f $X=-0.19 $Y=1.655 $X2=2.545 $Y2=1.615
cc_128 VPB N_VPWR_c_819_n 0.0180468f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_129 VPB N_VPWR_c_820_n 0.018718f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_130 VPB N_VPWR_c_810_n 0.0527941f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=1.23
cc_131 VPB N_VPWR_c_822_n 0.0241975f $X=-0.19 $Y=1.655 $X2=0.835 $Y2=1.065
cc_132 VPB N_VPWR_c_823_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_133 VPB GCLK 0.0499724f $X=-0.19 $Y=1.655 $X2=0.575 $Y2=2.595
cc_134 VPB N_GCLK_c_897_n 0.0125713f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=1.23
cc_135 N_A_80_21#_M1003_g N_GATE_M1007_g 0.0230569f $X=0.575 $Y=2.595 $X2=0
+ $Y2=0
cc_136 N_A_80_21#_c_150_n N_GATE_M1007_g 0.00154348f $X=1.725 $Y=2.515 $X2=0
+ $Y2=0
cc_137 N_A_80_21#_c_158_p N_GATE_M1007_g 5.48377e-19 $X=1.81 $Y=2.6 $X2=0 $Y2=0
cc_138 N_A_80_21#_M1000_g N_GATE_c_285_n 0.0144921f $X=0.835 $Y=0.445 $X2=0
+ $Y2=0
cc_139 N_A_80_21#_M1010_g N_GATE_c_285_n 0.0422575f $X=1.735 $Y=0.445 $X2=0
+ $Y2=0
cc_140 N_A_80_21#_M1000_g N_GATE_c_286_n 0.0157712f $X=0.835 $Y=0.445 $X2=0
+ $Y2=0
cc_141 N_A_80_21#_c_139_n N_GATE_c_286_n 0.00107342f $X=1.48 $Y=1.23 $X2=0 $Y2=0
cc_142 N_A_80_21#_M1003_g N_GATE_c_287_n 0.0181349f $X=0.575 $Y=2.595 $X2=0
+ $Y2=0
cc_143 N_A_80_21#_c_139_n N_GATE_c_287_n 0.00438096f $X=1.48 $Y=1.23 $X2=0 $Y2=0
cc_144 N_A_80_21#_c_141_n N_GATE_c_287_n 6.94548e-19 $X=1.725 $Y=1.78 $X2=0
+ $Y2=0
cc_145 N_A_80_21#_c_150_n N_GATE_c_287_n 3.92605e-19 $X=1.725 $Y=2.515 $X2=0
+ $Y2=0
cc_146 N_A_80_21#_M1003_g N_GATE_c_288_n 0.0238757f $X=0.575 $Y=2.595 $X2=0
+ $Y2=0
cc_147 N_A_80_21#_c_139_n N_GATE_c_288_n 0.0463577f $X=1.48 $Y=1.23 $X2=0 $Y2=0
cc_148 N_A_80_21#_c_140_n N_GATE_c_288_n 0.00265838f $X=0.61 $Y=1.23 $X2=0 $Y2=0
cc_149 N_A_80_21#_c_141_n N_GATE_c_288_n 0.00822456f $X=1.725 $Y=1.78 $X2=0
+ $Y2=0
cc_150 N_A_80_21#_c_150_n N_GATE_c_288_n 0.0149214f $X=1.725 $Y=2.515 $X2=0
+ $Y2=0
cc_151 N_A_80_21#_M1003_g N_GATE_c_289_n 0.00764736f $X=0.575 $Y=2.595 $X2=0
+ $Y2=0
cc_152 N_A_80_21#_M1010_g N_GATE_c_289_n 0.00848293f $X=1.735 $Y=0.445 $X2=0
+ $Y2=0
cc_153 N_A_80_21#_c_139_n N_GATE_c_289_n 0.0162381f $X=1.48 $Y=1.23 $X2=0 $Y2=0
cc_154 N_A_80_21#_c_140_n N_GATE_c_289_n 0.0219693f $X=0.61 $Y=1.23 $X2=0 $Y2=0
cc_155 N_A_80_21#_c_141_n N_GATE_c_289_n 0.00554248f $X=1.725 $Y=1.78 $X2=0
+ $Y2=0
cc_156 N_A_80_21#_c_145_n N_GATE_c_289_n 0.0210439f $X=1.645 $Y=1.285 $X2=0
+ $Y2=0
cc_157 N_A_80_21#_M1012_g N_A_27_47#_M1018_g 0.0221254f $X=2.505 $Y=2.595 $X2=0
+ $Y2=0
cc_158 N_A_80_21#_c_150_n N_A_27_47#_M1018_g 0.0240019f $X=1.725 $Y=2.515 $X2=0
+ $Y2=0
cc_159 N_A_80_21#_c_158_p N_A_27_47#_M1018_g 0.0108801f $X=1.81 $Y=2.6 $X2=0
+ $Y2=0
cc_160 N_A_80_21#_M1012_g N_A_27_47#_c_342_n 0.0128861f $X=2.505 $Y=2.595 $X2=0
+ $Y2=0
cc_161 N_A_80_21#_c_141_n N_A_27_47#_c_342_n 9.14057e-19 $X=1.725 $Y=1.78 $X2=0
+ $Y2=0
cc_162 N_A_80_21#_c_150_n N_A_27_47#_c_342_n 0.00250374f $X=1.725 $Y=2.515 $X2=0
+ $Y2=0
cc_163 N_A_80_21#_c_142_n N_A_27_47#_c_342_n 0.0193336f $X=2.545 $Y=1.615 $X2=0
+ $Y2=0
cc_164 N_A_80_21#_c_154_n N_A_27_47#_c_342_n 0.00563835f $X=4.32 $Y=2.5 $X2=0
+ $Y2=0
cc_165 N_A_80_21#_c_141_n N_A_27_47#_c_343_n 0.00435739f $X=1.725 $Y=1.78 $X2=0
+ $Y2=0
cc_166 N_A_80_21#_c_150_n N_A_27_47#_c_343_n 0.00138759f $X=1.725 $Y=2.515 $X2=0
+ $Y2=0
cc_167 N_A_80_21#_c_145_n N_A_27_47#_c_343_n 0.0167319f $X=1.645 $Y=1.285 $X2=0
+ $Y2=0
cc_168 N_A_80_21#_M1010_g N_A_27_47#_c_333_n 0.0154372f $X=1.735 $Y=0.445 $X2=0
+ $Y2=0
cc_169 N_A_80_21#_c_141_n N_A_27_47#_c_333_n 0.00245476f $X=1.725 $Y=1.78 $X2=0
+ $Y2=0
cc_170 N_A_80_21#_c_142_n N_A_27_47#_c_333_n 0.00141188f $X=2.545 $Y=1.615 $X2=0
+ $Y2=0
cc_171 N_A_80_21#_c_143_n N_A_27_47#_c_333_n 0.00139789f $X=2.545 $Y=1.615 $X2=0
+ $Y2=0
cc_172 N_A_80_21#_c_142_n N_A_27_47#_c_334_n 0.013893f $X=2.545 $Y=1.615 $X2=0
+ $Y2=0
cc_173 N_A_80_21#_c_143_n N_A_27_47#_c_334_n 0.0128861f $X=2.545 $Y=1.615 $X2=0
+ $Y2=0
cc_174 N_A_80_21#_c_145_n N_A_27_47#_c_334_n 0.0154372f $X=1.645 $Y=1.285 $X2=0
+ $Y2=0
cc_175 N_A_80_21#_M1010_g N_A_27_47#_c_335_n 0.0216275f $X=1.735 $Y=0.445 $X2=0
+ $Y2=0
cc_176 N_A_80_21#_M1013_g N_A_27_47#_c_336_n 0.00898882f $X=0.475 $Y=0.445 $X2=0
+ $Y2=0
cc_177 N_A_80_21#_M1000_g N_A_27_47#_c_336_n 0.00163457f $X=0.835 $Y=0.445 $X2=0
+ $Y2=0
cc_178 N_A_80_21#_M1013_g N_A_27_47#_c_337_n 0.00887731f $X=0.475 $Y=0.445 $X2=0
+ $Y2=0
cc_179 N_A_80_21#_M1000_g N_A_27_47#_c_337_n 0.0110391f $X=0.835 $Y=0.445 $X2=0
+ $Y2=0
cc_180 N_A_80_21#_M1010_g N_A_27_47#_c_337_n 0.0115942f $X=1.735 $Y=0.445 $X2=0
+ $Y2=0
cc_181 N_A_80_21#_c_139_n N_A_27_47#_c_337_n 0.0746893f $X=1.48 $Y=1.23 $X2=0
+ $Y2=0
cc_182 N_A_80_21#_c_140_n N_A_27_47#_c_337_n 7.85225e-19 $X=0.61 $Y=1.23 $X2=0
+ $Y2=0
cc_183 N_A_80_21#_c_141_n N_A_27_47#_c_337_n 0.0249207f $X=1.725 $Y=1.78 $X2=0
+ $Y2=0
cc_184 N_A_80_21#_c_142_n N_A_27_47#_c_337_n 0.00932518f $X=2.545 $Y=1.615 $X2=0
+ $Y2=0
cc_185 N_A_80_21#_c_145_n N_A_27_47#_c_337_n 0.00108366f $X=1.645 $Y=1.285 $X2=0
+ $Y2=0
cc_186 N_A_80_21#_M1013_g N_A_27_47#_c_338_n 0.00499595f $X=0.475 $Y=0.445 $X2=0
+ $Y2=0
cc_187 N_A_80_21#_M1003_g N_A_27_47#_c_345_n 0.0141471f $X=0.575 $Y=2.595 $X2=0
+ $Y2=0
cc_188 N_A_80_21#_M1013_g N_A_27_47#_c_339_n 0.0128246f $X=0.475 $Y=0.445 $X2=0
+ $Y2=0
cc_189 N_A_80_21#_M1003_g N_A_27_47#_c_339_n 0.0245003f $X=0.575 $Y=2.595 $X2=0
+ $Y2=0
cc_190 N_A_80_21#_c_139_n N_A_27_47#_c_339_n 0.0250954f $X=1.48 $Y=1.23 $X2=0
+ $Y2=0
cc_191 N_A_80_21#_M1010_g N_A_27_47#_c_340_n 0.00120383f $X=1.735 $Y=0.445 $X2=0
+ $Y2=0
cc_192 N_A_80_21#_c_141_n N_A_27_47#_c_340_n 0.00160415f $X=1.725 $Y=1.78 $X2=0
+ $Y2=0
cc_193 N_A_80_21#_c_142_n N_A_27_47#_c_340_n 0.0147059f $X=2.545 $Y=1.615 $X2=0
+ $Y2=0
cc_194 N_A_80_21#_c_154_n N_A_584_21#_M1015_d 0.00748071f $X=4.32 $Y=2.5 $X2=0
+ $Y2=0
cc_195 N_A_80_21#_M1012_g N_A_584_21#_M1001_g 0.064089f $X=2.505 $Y=2.595 $X2=0
+ $Y2=0
cc_196 N_A_80_21#_c_142_n N_A_584_21#_M1001_g 4.28013e-19 $X=2.545 $Y=1.615
+ $X2=0 $Y2=0
cc_197 N_A_80_21#_c_143_n N_A_584_21#_M1001_g 0.00338753f $X=2.545 $Y=1.615
+ $X2=0 $Y2=0
cc_198 N_A_80_21#_c_154_n N_A_584_21#_M1001_g 0.0176535f $X=4.32 $Y=2.5 $X2=0
+ $Y2=0
cc_199 N_A_80_21#_c_144_n N_A_584_21#_c_425_n 0.0081224f $X=4.405 $Y=2.315 $X2=0
+ $Y2=0
cc_200 N_A_80_21#_c_146_n N_A_584_21#_c_425_n 0.0189687f $X=4.325 $Y=1.06 $X2=0
+ $Y2=0
cc_201 N_A_80_21#_c_144_n N_A_584_21#_c_426_n 0.0477354f $X=4.405 $Y=2.315 $X2=0
+ $Y2=0
cc_202 N_A_80_21#_c_144_n N_A_584_21#_c_428_n 0.0496545f $X=4.405 $Y=2.315 $X2=0
+ $Y2=0
cc_203 N_A_80_21#_c_146_n N_A_584_21#_c_428_n 0.00995243f $X=4.325 $Y=1.06 $X2=0
+ $Y2=0
cc_204 N_A_80_21#_M1020_s N_A_584_21#_c_438_n 6.22097e-19 $X=4.67 $Y=2.095 $X2=0
+ $Y2=0
cc_205 N_A_80_21#_c_155_n N_A_584_21#_c_438_n 0.00593632f $X=4.815 $Y=2.48 $X2=0
+ $Y2=0
cc_206 N_A_80_21#_M1020_s N_A_584_21#_c_439_n 0.00261901f $X=4.67 $Y=2.095 $X2=0
+ $Y2=0
cc_207 N_A_80_21#_c_144_n N_A_584_21#_c_439_n 0.0137159f $X=4.405 $Y=2.315 $X2=0
+ $Y2=0
cc_208 N_A_80_21#_c_155_n N_A_584_21#_c_439_n 0.0139849f $X=4.815 $Y=2.48 $X2=0
+ $Y2=0
cc_209 N_A_80_21#_c_142_n N_A_584_21#_c_430_n 0.0177797f $X=2.545 $Y=1.615 $X2=0
+ $Y2=0
cc_210 N_A_80_21#_c_143_n N_A_584_21#_c_430_n 3.33456e-19 $X=2.545 $Y=1.615
+ $X2=0 $Y2=0
cc_211 N_A_80_21#_c_142_n N_A_584_21#_c_431_n 9.17588e-19 $X=2.545 $Y=1.615
+ $X2=0 $Y2=0
cc_212 N_A_80_21#_c_143_n N_A_584_21#_c_431_n 0.0166807f $X=2.545 $Y=1.615 $X2=0
+ $Y2=0
cc_213 N_A_80_21#_c_144_n N_A_584_21#_c_444_n 0.0122461f $X=4.405 $Y=2.315 $X2=0
+ $Y2=0
cc_214 N_A_80_21#_c_154_n N_A_584_21#_c_444_n 0.0211286f $X=4.32 $Y=2.5 $X2=0
+ $Y2=0
cc_215 N_A_80_21#_c_155_n N_A_584_21#_c_444_n 0.00154168f $X=4.815 $Y=2.48 $X2=0
+ $Y2=0
cc_216 N_A_80_21#_c_146_n N_A_584_21#_c_432_n 0.021397f $X=4.325 $Y=1.06 $X2=0
+ $Y2=0
cc_217 N_A_80_21#_c_144_n N_A_584_21#_c_433_n 0.0135989f $X=4.405 $Y=2.315 $X2=0
+ $Y2=0
cc_218 N_A_80_21#_c_154_n N_A_352_419#_M1018_d 0.0185516f $X=4.32 $Y=2.5 $X2=0
+ $Y2=0
cc_219 N_A_80_21#_c_154_n N_A_352_419#_M1015_g 0.0220262f $X=4.32 $Y=2.5 $X2=0
+ $Y2=0
cc_220 N_A_80_21#_c_155_n N_A_352_419#_M1015_g 0.00398439f $X=4.815 $Y=2.48
+ $X2=0 $Y2=0
cc_221 N_A_80_21#_M1010_g N_A_352_419#_c_598_n 0.00536545f $X=1.735 $Y=0.445
+ $X2=0 $Y2=0
cc_222 N_A_80_21#_M1012_g N_A_352_419#_c_591_n 0.017999f $X=2.505 $Y=2.595 $X2=0
+ $Y2=0
cc_223 N_A_80_21#_c_150_n N_A_352_419#_c_591_n 0.00887143f $X=1.725 $Y=2.515
+ $X2=0 $Y2=0
cc_224 N_A_80_21#_c_142_n N_A_352_419#_c_591_n 0.0325942f $X=2.545 $Y=1.615
+ $X2=0 $Y2=0
cc_225 N_A_80_21#_c_143_n N_A_352_419#_c_591_n 0.00166727f $X=2.545 $Y=1.615
+ $X2=0 $Y2=0
cc_226 N_A_80_21#_c_154_n N_A_352_419#_c_591_n 0.0866509f $X=4.32 $Y=2.5 $X2=0
+ $Y2=0
cc_227 N_A_80_21#_c_142_n N_A_352_419#_c_585_n 0.00600601f $X=2.545 $Y=1.615
+ $X2=0 $Y2=0
cc_228 N_A_80_21#_c_143_n N_A_352_419#_c_585_n 0.00247228f $X=2.545 $Y=1.615
+ $X2=0 $Y2=0
cc_229 N_A_80_21#_c_154_n N_A_352_419#_c_593_n 0.00461473f $X=4.32 $Y=2.5 $X2=0
+ $Y2=0
cc_230 N_A_80_21#_c_154_n N_A_352_419#_c_587_n 2.28234e-19 $X=4.32 $Y=2.5 $X2=0
+ $Y2=0
cc_231 N_A_80_21#_c_146_n N_A_352_419#_c_588_n 2.36794e-19 $X=4.325 $Y=1.06
+ $X2=0 $Y2=0
cc_232 N_A_80_21#_c_144_n N_A_352_419#_c_589_n 8.94466e-19 $X=4.405 $Y=2.315
+ $X2=0 $Y2=0
cc_233 N_A_80_21#_c_144_n N_CLK_c_688_n 0.00679063f $X=4.405 $Y=2.315 $X2=-0.19
+ $Y2=-0.245
cc_234 N_A_80_21#_c_146_n N_CLK_c_688_n 0.00333432f $X=4.325 $Y=1.06 $X2=-0.19
+ $Y2=-0.245
cc_235 N_A_80_21#_c_144_n N_CLK_c_690_n 0.00557936f $X=4.405 $Y=2.315 $X2=0
+ $Y2=0
cc_236 N_A_80_21#_c_144_n N_CLK_M1020_g 0.00504717f $X=4.405 $Y=2.315 $X2=0
+ $Y2=0
cc_237 N_A_80_21#_c_155_n N_CLK_M1020_g 0.014117f $X=4.815 $Y=2.48 $X2=0 $Y2=0
cc_238 N_A_80_21#_c_154_n N_VPWR_M1001_d 0.00511493f $X=4.32 $Y=2.5 $X2=0 $Y2=0
cc_239 N_A_80_21#_M1003_g N_VPWR_c_811_n 0.0199704f $X=0.575 $Y=2.595 $X2=0
+ $Y2=0
cc_240 N_A_80_21#_M1012_g N_VPWR_c_812_n 0.001781f $X=2.505 $Y=2.595 $X2=0 $Y2=0
cc_241 N_A_80_21#_c_154_n N_VPWR_c_812_n 0.0187678f $X=4.32 $Y=2.5 $X2=0 $Y2=0
cc_242 N_A_80_21#_c_155_n N_VPWR_c_813_n 0.0507784f $X=4.815 $Y=2.48 $X2=0 $Y2=0
cc_243 N_A_80_21#_M1012_g N_VPWR_c_815_n 0.00710941f $X=2.505 $Y=2.595 $X2=0
+ $Y2=0
cc_244 N_A_80_21#_c_158_p N_VPWR_c_815_n 0.0025723f $X=1.81 $Y=2.6 $X2=0 $Y2=0
cc_245 N_A_80_21#_c_154_n N_VPWR_c_815_n 0.0215114f $X=4.32 $Y=2.5 $X2=0 $Y2=0
cc_246 N_A_80_21#_c_154_n N_VPWR_c_817_n 0.0192064f $X=4.32 $Y=2.5 $X2=0 $Y2=0
cc_247 N_A_80_21#_c_155_n N_VPWR_c_817_n 0.0190308f $X=4.815 $Y=2.48 $X2=0 $Y2=0
cc_248 N_A_80_21#_M1020_s N_VPWR_c_810_n 0.0023218f $X=4.67 $Y=2.095 $X2=0 $Y2=0
cc_249 N_A_80_21#_M1003_g N_VPWR_c_810_n 0.01455f $X=0.575 $Y=2.595 $X2=0 $Y2=0
cc_250 N_A_80_21#_M1012_g N_VPWR_c_810_n 0.00977333f $X=2.505 $Y=2.595 $X2=0
+ $Y2=0
cc_251 N_A_80_21#_c_158_p N_VPWR_c_810_n 0.00448973f $X=1.81 $Y=2.6 $X2=0 $Y2=0
cc_252 N_A_80_21#_c_154_n N_VPWR_c_810_n 0.0693537f $X=4.32 $Y=2.5 $X2=0 $Y2=0
cc_253 N_A_80_21#_c_155_n N_VPWR_c_810_n 0.0123181f $X=4.815 $Y=2.48 $X2=0 $Y2=0
cc_254 N_A_80_21#_M1003_g N_VPWR_c_822_n 0.00840199f $X=0.575 $Y=2.595 $X2=0
+ $Y2=0
cc_255 N_A_80_21#_c_154_n A_526_419# 0.00587672f $X=4.32 $Y=2.5 $X2=-0.19
+ $Y2=-0.245
cc_256 N_A_80_21#_M1013_g N_VGND_c_919_n 0.00201689f $X=0.475 $Y=0.445 $X2=0
+ $Y2=0
cc_257 N_A_80_21#_M1000_g N_VGND_c_919_n 0.0100125f $X=0.835 $Y=0.445 $X2=0
+ $Y2=0
cc_258 N_A_80_21#_M1010_g N_VGND_c_920_n 0.00423733f $X=1.735 $Y=0.445 $X2=0
+ $Y2=0
cc_259 N_A_80_21#_M1013_g N_VGND_c_927_n 0.00425202f $X=0.475 $Y=0.445 $X2=0
+ $Y2=0
cc_260 N_A_80_21#_M1000_g N_VGND_c_927_n 0.00362954f $X=0.835 $Y=0.445 $X2=0
+ $Y2=0
cc_261 N_A_80_21#_M1013_g N_VGND_c_929_n 0.00687266f $X=0.475 $Y=0.445 $X2=0
+ $Y2=0
cc_262 N_A_80_21#_M1000_g N_VGND_c_929_n 0.00414614f $X=0.835 $Y=0.445 $X2=0
+ $Y2=0
cc_263 N_A_80_21#_M1010_g N_VGND_c_929_n 0.00602521f $X=1.735 $Y=0.445 $X2=0
+ $Y2=0
cc_264 N_GATE_M1007_g N_A_27_47#_M1018_g 0.043123f $X=1.145 $Y=2.595 $X2=0 $Y2=0
cc_265 N_GATE_c_287_n N_A_27_47#_c_343_n 0.043123f $X=1.105 $Y=1.77 $X2=0 $Y2=0
cc_266 N_GATE_c_288_n N_A_27_47#_c_343_n 0.00184002f $X=1.105 $Y=1.77 $X2=0
+ $Y2=0
cc_267 N_GATE_c_285_n N_A_27_47#_c_337_n 0.00426087f $X=1.345 $Y=0.73 $X2=0
+ $Y2=0
cc_268 N_GATE_c_286_n N_A_27_47#_c_337_n 0.0113137f $X=1.345 $Y=0.805 $X2=0
+ $Y2=0
cc_269 N_GATE_c_289_n N_A_27_47#_c_337_n 0.00215693f $X=1.105 $Y=1.605 $X2=0
+ $Y2=0
cc_270 N_GATE_c_288_n N_A_27_47#_c_339_n 0.0256226f $X=1.105 $Y=1.77 $X2=0 $Y2=0
cc_271 N_GATE_c_285_n N_A_352_419#_c_598_n 7.8437e-19 $X=1.345 $Y=0.73 $X2=0
+ $Y2=0
cc_272 N_GATE_c_288_n N_VPWR_M1003_d 0.00232502f $X=1.105 $Y=1.77 $X2=-0.19
+ $Y2=-0.245
cc_273 N_GATE_M1007_g N_VPWR_c_811_n 0.00362166f $X=1.145 $Y=2.595 $X2=0 $Y2=0
cc_274 N_GATE_c_287_n N_VPWR_c_811_n 2.25906e-19 $X=1.105 $Y=1.77 $X2=0 $Y2=0
cc_275 N_GATE_c_288_n N_VPWR_c_811_n 0.0192848f $X=1.105 $Y=1.77 $X2=0 $Y2=0
cc_276 N_GATE_M1007_g N_VPWR_c_815_n 0.00975641f $X=1.145 $Y=2.595 $X2=0 $Y2=0
cc_277 N_GATE_M1007_g N_VPWR_c_810_n 0.0168693f $X=1.145 $Y=2.595 $X2=0 $Y2=0
cc_278 N_GATE_c_285_n N_VGND_c_919_n 0.00458721f $X=1.345 $Y=0.73 $X2=0 $Y2=0
cc_279 N_GATE_c_286_n N_VGND_c_919_n 6.89717e-19 $X=1.345 $Y=0.805 $X2=0 $Y2=0
cc_280 N_GATE_c_285_n N_VGND_c_920_n 0.00436487f $X=1.345 $Y=0.73 $X2=0 $Y2=0
cc_281 N_GATE_c_285_n N_VGND_c_929_n 0.00624169f $X=1.345 $Y=0.73 $X2=0 $Y2=0
cc_282 N_A_27_47#_c_333_n N_A_584_21#_M1011_g 0.00590588f $X=2.095 $Y=1.095
+ $X2=0 $Y2=0
cc_283 N_A_27_47#_c_335_n N_A_584_21#_M1011_g 0.00743726f $X=2.165 $Y=0.765
+ $X2=0 $Y2=0
cc_284 N_A_27_47#_c_340_n N_A_584_21#_M1011_g 2.46693e-19 $X=2.255 $Y=0.8 $X2=0
+ $Y2=0
cc_285 N_A_27_47#_c_333_n N_A_352_419#_c_598_n 0.00100251f $X=2.095 $Y=1.095
+ $X2=0 $Y2=0
cc_286 N_A_27_47#_c_335_n N_A_352_419#_c_598_n 0.0124321f $X=2.165 $Y=0.765
+ $X2=0 $Y2=0
cc_287 N_A_27_47#_c_337_n N_A_352_419#_c_598_n 0.0169705f $X=2.09 $Y=0.8 $X2=0
+ $Y2=0
cc_288 N_A_27_47#_c_340_n N_A_352_419#_c_598_n 0.0214529f $X=2.255 $Y=0.8 $X2=0
+ $Y2=0
cc_289 N_A_27_47#_M1018_g N_A_352_419#_c_591_n 0.00119285f $X=1.635 $Y=2.595
+ $X2=0 $Y2=0
cc_290 N_A_27_47#_c_342_n N_A_352_419#_c_591_n 0.00247499f $X=2.02 $Y=1.765
+ $X2=0 $Y2=0
cc_291 N_A_27_47#_c_333_n N_A_352_419#_c_584_n 4.33799e-19 $X=2.095 $Y=1.095
+ $X2=0 $Y2=0
cc_292 N_A_27_47#_c_335_n N_A_352_419#_c_584_n 0.00357318f $X=2.165 $Y=0.765
+ $X2=0 $Y2=0
cc_293 N_A_27_47#_c_340_n N_A_352_419#_c_584_n 0.00737081f $X=2.255 $Y=0.8 $X2=0
+ $Y2=0
cc_294 N_A_27_47#_c_333_n N_A_352_419#_c_585_n 0.00273601f $X=2.095 $Y=1.095
+ $X2=0 $Y2=0
cc_295 N_A_27_47#_c_334_n N_A_352_419#_c_585_n 0.00154911f $X=2.095 $Y=1.69
+ $X2=0 $Y2=0
cc_296 N_A_27_47#_c_340_n N_A_352_419#_c_585_n 0.0226185f $X=2.255 $Y=0.8 $X2=0
+ $Y2=0
cc_297 N_A_27_47#_c_345_n N_VPWR_c_811_n 0.0489245f $X=0.31 $Y=2.495 $X2=0 $Y2=0
cc_298 N_A_27_47#_M1018_g N_VPWR_c_815_n 0.00848468f $X=1.635 $Y=2.595 $X2=0
+ $Y2=0
cc_299 N_A_27_47#_M1003_s N_VPWR_c_810_n 0.0023218f $X=0.165 $Y=2.095 $X2=0
+ $Y2=0
cc_300 N_A_27_47#_M1018_g N_VPWR_c_810_n 0.013835f $X=1.635 $Y=2.595 $X2=0 $Y2=0
cc_301 N_A_27_47#_c_345_n N_VPWR_c_810_n 0.0144427f $X=0.31 $Y=2.495 $X2=0 $Y2=0
cc_302 N_A_27_47#_c_345_n N_VPWR_c_822_n 0.0231292f $X=0.31 $Y=2.495 $X2=0 $Y2=0
cc_303 N_A_27_47#_c_336_n N_VGND_c_919_n 0.00903348f $X=0.26 $Y=0.47 $X2=0 $Y2=0
cc_304 N_A_27_47#_c_337_n N_VGND_c_919_n 0.0221076f $X=2.09 $Y=0.8 $X2=0 $Y2=0
cc_305 N_A_27_47#_c_335_n N_VGND_c_920_n 0.00359964f $X=2.165 $Y=0.765 $X2=0
+ $Y2=0
cc_306 N_A_27_47#_c_337_n N_VGND_c_920_n 0.00831946f $X=2.09 $Y=0.8 $X2=0 $Y2=0
cc_307 N_A_27_47#_c_336_n N_VGND_c_927_n 0.0197709f $X=0.26 $Y=0.47 $X2=0 $Y2=0
cc_308 N_A_27_47#_c_337_n N_VGND_c_927_n 0.00665482f $X=2.09 $Y=0.8 $X2=0 $Y2=0
cc_309 N_A_27_47#_M1013_s N_VGND_c_929_n 0.00216211f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_310 N_A_27_47#_c_335_n N_VGND_c_929_n 0.00621233f $X=2.165 $Y=0.765 $X2=0
+ $Y2=0
cc_311 N_A_27_47#_c_336_n N_VGND_c_929_n 0.0125654f $X=0.26 $Y=0.47 $X2=0 $Y2=0
cc_312 N_A_27_47#_c_337_n N_VGND_c_929_n 0.0269021f $X=2.09 $Y=0.8 $X2=0 $Y2=0
cc_313 N_A_584_21#_M1011_g N_A_352_419#_M1019_g 0.0149944f $X=2.995 $Y=0.445
+ $X2=0 $Y2=0
cc_314 N_A_584_21#_c_425_n N_A_352_419#_M1019_g 7.78171e-19 $X=3.895 $Y=1.325
+ $X2=0 $Y2=0
cc_315 N_A_584_21#_c_432_n N_A_352_419#_M1019_g 0.00135363f $X=4.195 $Y=0.47
+ $X2=0 $Y2=0
cc_316 N_A_584_21#_M1001_g N_A_352_419#_M1015_g 0.0398677f $X=3.075 $Y=2.595
+ $X2=0 $Y2=0
cc_317 N_A_584_21#_c_444_n N_A_352_419#_M1015_g 0.00375038f $X=4.055 $Y=2.245
+ $X2=0 $Y2=0
cc_318 N_A_584_21#_c_425_n N_A_352_419#_M1023_g 0.00551413f $X=3.895 $Y=1.325
+ $X2=0 $Y2=0
cc_319 N_A_584_21#_c_432_n N_A_352_419#_M1023_g 0.00963098f $X=4.195 $Y=0.47
+ $X2=0 $Y2=0
cc_320 N_A_584_21#_M1011_g N_A_352_419#_c_598_n 0.00329049f $X=2.995 $Y=0.445
+ $X2=0 $Y2=0
cc_321 N_A_584_21#_M1001_g N_A_352_419#_c_591_n 0.0219547f $X=3.075 $Y=2.595
+ $X2=0 $Y2=0
cc_322 N_A_584_21#_c_424_n N_A_352_419#_c_591_n 0.00595601f $X=3.81 $Y=1.41
+ $X2=0 $Y2=0
cc_323 N_A_584_21#_c_426_n N_A_352_419#_c_591_n 0.00347008f $X=4.055 $Y=2.155
+ $X2=0 $Y2=0
cc_324 N_A_584_21#_c_430_n N_A_352_419#_c_591_n 0.0137648f $X=3.085 $Y=1.41
+ $X2=0 $Y2=0
cc_325 N_A_584_21#_c_431_n N_A_352_419#_c_591_n 4.89801e-19 $X=3.085 $Y=1.55
+ $X2=0 $Y2=0
cc_326 N_A_584_21#_c_444_n N_A_352_419#_c_591_n 0.0137214f $X=4.055 $Y=2.245
+ $X2=0 $Y2=0
cc_327 N_A_584_21#_M1011_g N_A_352_419#_c_584_n 0.00547614f $X=2.995 $Y=0.445
+ $X2=0 $Y2=0
cc_328 N_A_584_21#_M1011_g N_A_352_419#_c_586_n 0.018689f $X=2.995 $Y=0.445
+ $X2=0 $Y2=0
cc_329 N_A_584_21#_c_424_n N_A_352_419#_c_586_n 0.0270354f $X=3.81 $Y=1.41 $X2=0
+ $Y2=0
cc_330 N_A_584_21#_c_425_n N_A_352_419#_c_586_n 0.0245347f $X=3.895 $Y=1.325
+ $X2=0 $Y2=0
cc_331 N_A_584_21#_c_430_n N_A_352_419#_c_586_n 0.0254321f $X=3.085 $Y=1.41
+ $X2=0 $Y2=0
cc_332 N_A_584_21#_c_431_n N_A_352_419#_c_586_n 0.00111385f $X=3.085 $Y=1.55
+ $X2=0 $Y2=0
cc_333 N_A_584_21#_M1001_g N_A_352_419#_c_592_n 0.00283734f $X=3.075 $Y=2.595
+ $X2=0 $Y2=0
cc_334 N_A_584_21#_c_426_n N_A_352_419#_c_592_n 0.00557292f $X=4.055 $Y=2.155
+ $X2=0 $Y2=0
cc_335 N_A_584_21#_M1001_g N_A_352_419#_c_593_n 0.0049236f $X=3.075 $Y=2.595
+ $X2=0 $Y2=0
cc_336 N_A_584_21#_c_424_n N_A_352_419#_c_593_n 0.0250064f $X=3.81 $Y=1.41 $X2=0
+ $Y2=0
cc_337 N_A_584_21#_c_426_n N_A_352_419#_c_593_n 0.0187832f $X=4.055 $Y=2.155
+ $X2=0 $Y2=0
cc_338 N_A_584_21#_c_430_n N_A_352_419#_c_593_n 0.00299117f $X=3.085 $Y=1.41
+ $X2=0 $Y2=0
cc_339 N_A_584_21#_c_431_n N_A_352_419#_c_593_n 2.22854e-19 $X=3.085 $Y=1.55
+ $X2=0 $Y2=0
cc_340 N_A_584_21#_c_444_n N_A_352_419#_c_593_n 5.72585e-19 $X=4.055 $Y=2.245
+ $X2=0 $Y2=0
cc_341 N_A_584_21#_M1001_g N_A_352_419#_c_587_n 0.0103528f $X=3.075 $Y=2.595
+ $X2=0 $Y2=0
cc_342 N_A_584_21#_c_424_n N_A_352_419#_c_587_n 0.0025571f $X=3.81 $Y=1.41 $X2=0
+ $Y2=0
cc_343 N_A_584_21#_c_426_n N_A_352_419#_c_587_n 0.0126453f $X=4.055 $Y=2.155
+ $X2=0 $Y2=0
cc_344 N_A_584_21#_c_430_n N_A_352_419#_c_587_n 5.5464e-19 $X=3.085 $Y=1.41
+ $X2=0 $Y2=0
cc_345 N_A_584_21#_c_431_n N_A_352_419#_c_587_n 0.0072578f $X=3.085 $Y=1.55
+ $X2=0 $Y2=0
cc_346 N_A_584_21#_M1011_g N_A_352_419#_c_588_n 0.0190979f $X=2.995 $Y=0.445
+ $X2=0 $Y2=0
cc_347 N_A_584_21#_c_424_n N_A_352_419#_c_588_n 0.00790171f $X=3.81 $Y=1.41
+ $X2=0 $Y2=0
cc_348 N_A_584_21#_c_425_n N_A_352_419#_c_588_n 0.016758f $X=3.895 $Y=1.325
+ $X2=0 $Y2=0
cc_349 N_A_584_21#_c_433_n N_A_352_419#_c_588_n 2.31092e-19 $X=4.055 $Y=1.41
+ $X2=0 $Y2=0
cc_350 N_A_584_21#_M1011_g N_A_352_419#_c_589_n 0.00784646f $X=2.995 $Y=0.445
+ $X2=0 $Y2=0
cc_351 N_A_584_21#_c_424_n N_A_352_419#_c_589_n 0.0124929f $X=3.81 $Y=1.41 $X2=0
+ $Y2=0
cc_352 N_A_584_21#_c_426_n N_A_352_419#_c_589_n 0.00316148f $X=4.055 $Y=2.155
+ $X2=0 $Y2=0
cc_353 N_A_584_21#_c_430_n N_A_352_419#_c_589_n 8.51848e-19 $X=3.085 $Y=1.41
+ $X2=0 $Y2=0
cc_354 N_A_584_21#_c_431_n N_A_352_419#_c_589_n 0.0121506f $X=3.085 $Y=1.55
+ $X2=0 $Y2=0
cc_355 N_A_584_21#_c_425_n N_CLK_c_688_n 0.00253914f $X=3.895 $Y=1.325 $X2=-0.19
+ $Y2=-0.245
cc_356 N_A_584_21#_c_427_n N_CLK_c_688_n 0.00619211f $X=4.67 $Y=0.59 $X2=-0.19
+ $Y2=-0.245
cc_357 N_A_584_21#_c_428_n N_CLK_c_688_n 0.00554447f $X=4.755 $Y=1.965 $X2=-0.19
+ $Y2=-0.245
cc_358 N_A_584_21#_c_433_n N_CLK_c_688_n 9.43282e-19 $X=4.055 $Y=1.41 $X2=-0.19
+ $Y2=-0.245
cc_359 N_A_584_21#_c_428_n N_CLK_c_689_n 0.0136217f $X=4.755 $Y=1.965 $X2=0
+ $Y2=0
cc_360 N_A_584_21#_c_438_n N_CLK_c_689_n 0.00329847f $X=5.945 $Y=2.05 $X2=0
+ $Y2=0
cc_361 N_A_584_21#_c_426_n N_CLK_c_690_n 5.34804e-19 $X=4.055 $Y=2.155 $X2=0
+ $Y2=0
cc_362 N_A_584_21#_c_428_n N_CLK_c_691_n 0.00781715f $X=4.755 $Y=1.965 $X2=0
+ $Y2=0
cc_363 N_A_584_21#_c_438_n N_CLK_M1020_g 0.0243517f $X=5.945 $Y=2.05 $X2=0 $Y2=0
cc_364 N_A_584_21#_c_423_n N_CLK_c_692_n 0.0201417f $X=5.835 $Y=1.42 $X2=0 $Y2=0
cc_365 N_A_584_21#_c_438_n N_CLK_M1008_g 0.0229471f $X=5.945 $Y=2.05 $X2=0 $Y2=0
cc_366 N_A_584_21#_c_428_n CLK 0.0243332f $X=4.755 $Y=1.965 $X2=0 $Y2=0
cc_367 N_A_584_21#_c_438_n CLK 0.0434832f $X=5.945 $Y=2.05 $X2=0 $Y2=0
cc_368 N_A_584_21#_c_440_n CLK 0.0127821f $X=6.11 $Y=1.71 $X2=0 $Y2=0
cc_369 N_A_584_21#_c_429_n CLK 0.0045851f $X=6.11 $Y=1.71 $X2=0 $Y2=0
cc_370 N_A_584_21#_M1004_g N_CLK_c_694_n 0.0280173f $X=6.14 $Y=2.595 $X2=0 $Y2=0
cc_371 N_A_584_21#_c_428_n N_CLK_c_694_n 0.0127675f $X=4.755 $Y=1.965 $X2=0
+ $Y2=0
cc_372 N_A_584_21#_c_438_n N_CLK_c_694_n 0.00396695f $X=5.945 $Y=2.05 $X2=0
+ $Y2=0
cc_373 N_A_584_21#_c_440_n N_CLK_c_694_n 0.00303593f $X=6.11 $Y=1.71 $X2=0 $Y2=0
cc_374 N_A_584_21#_c_429_n N_CLK_c_694_n 0.030948f $X=6.11 $Y=1.71 $X2=0 $Y2=0
cc_375 N_A_584_21#_c_438_n N_A_1147_419#_M1008_d 0.00179048f $X=5.945 $Y=2.05
+ $X2=0 $Y2=0
cc_376 N_A_584_21#_c_423_n N_A_1147_419#_M1002_g 0.0074551f $X=5.835 $Y=1.42
+ $X2=0 $Y2=0
cc_377 N_A_584_21#_M1004_g N_A_1147_419#_M1021_g 0.0431392f $X=6.14 $Y=2.595
+ $X2=0 $Y2=0
cc_378 N_A_584_21#_c_438_n N_A_1147_419#_M1021_g 5.07547e-19 $X=5.945 $Y=2.05
+ $X2=0 $Y2=0
cc_379 N_A_584_21#_c_440_n N_A_1147_419#_M1021_g 6.34981e-19 $X=6.11 $Y=1.71
+ $X2=0 $Y2=0
cc_380 N_A_584_21#_c_429_n N_A_1147_419#_M1021_g 0.0136187f $X=6.11 $Y=1.71
+ $X2=0 $Y2=0
cc_381 N_A_584_21#_c_429_n N_A_1147_419#_c_744_n 0.0105993f $X=6.11 $Y=1.71
+ $X2=0 $Y2=0
cc_382 N_A_584_21#_M1004_g N_A_1147_419#_c_759_n 0.0138364f $X=6.14 $Y=2.595
+ $X2=0 $Y2=0
cc_383 N_A_584_21#_c_438_n N_A_1147_419#_c_759_n 0.0161411f $X=5.945 $Y=2.05
+ $X2=0 $Y2=0
cc_384 N_A_584_21#_c_440_n N_A_1147_419#_c_745_n 0.00216063f $X=6.11 $Y=1.71
+ $X2=0 $Y2=0
cc_385 N_A_584_21#_c_429_n N_A_1147_419#_c_745_n 0.00135769f $X=6.11 $Y=1.71
+ $X2=0 $Y2=0
cc_386 N_A_584_21#_c_423_n N_A_1147_419#_c_763_n 3.77262e-19 $X=5.835 $Y=1.42
+ $X2=0 $Y2=0
cc_387 N_A_584_21#_c_429_n N_A_1147_419#_c_763_n 0.00104031f $X=6.11 $Y=1.71
+ $X2=0 $Y2=0
cc_388 N_A_584_21#_M1004_g N_A_1147_419#_c_747_n 0.00438896f $X=6.14 $Y=2.595
+ $X2=0 $Y2=0
cc_389 N_A_584_21#_c_438_n N_A_1147_419#_c_747_n 0.0106632f $X=5.945 $Y=2.05
+ $X2=0 $Y2=0
cc_390 N_A_584_21#_c_429_n N_A_1147_419#_c_747_n 0.00181047f $X=6.11 $Y=1.71
+ $X2=0 $Y2=0
cc_391 N_A_584_21#_M1004_g N_A_1147_419#_c_768_n 0.0116315f $X=6.14 $Y=2.595
+ $X2=0 $Y2=0
cc_392 N_A_584_21#_c_438_n N_A_1147_419#_c_768_n 0.0167406f $X=5.945 $Y=2.05
+ $X2=0 $Y2=0
cc_393 N_A_584_21#_c_423_n N_A_1147_419#_c_748_n 0.0102092f $X=5.835 $Y=1.42
+ $X2=0 $Y2=0
cc_394 N_A_584_21#_c_438_n N_A_1147_419#_c_748_n 0.00186922f $X=5.945 $Y=2.05
+ $X2=0 $Y2=0
cc_395 N_A_584_21#_c_440_n N_A_1147_419#_c_748_n 0.0219545f $X=6.11 $Y=1.71
+ $X2=0 $Y2=0
cc_396 N_A_584_21#_c_429_n N_A_1147_419#_c_748_n 0.00922015f $X=6.11 $Y=1.71
+ $X2=0 $Y2=0
cc_397 N_A_584_21#_c_423_n N_A_1147_419#_c_749_n 0.00371424f $X=5.835 $Y=1.42
+ $X2=0 $Y2=0
cc_398 N_A_584_21#_c_440_n N_A_1147_419#_c_775_n 0.027199f $X=6.11 $Y=1.71 $X2=0
+ $Y2=0
cc_399 N_A_584_21#_c_438_n N_VPWR_M1020_d 0.00180746f $X=5.945 $Y=2.05 $X2=0
+ $Y2=0
cc_400 N_A_584_21#_M1001_g N_VPWR_c_812_n 0.00986369f $X=3.075 $Y=2.595 $X2=0
+ $Y2=0
cc_401 N_A_584_21#_M1004_g N_VPWR_c_813_n 0.00113722f $X=6.14 $Y=2.595 $X2=0
+ $Y2=0
cc_402 N_A_584_21#_c_438_n N_VPWR_c_813_n 0.0163514f $X=5.945 $Y=2.05 $X2=0
+ $Y2=0
cc_403 N_A_584_21#_M1004_g N_VPWR_c_814_n 0.0131232f $X=6.14 $Y=2.595 $X2=0
+ $Y2=0
cc_404 N_A_584_21#_M1001_g N_VPWR_c_815_n 0.00653347f $X=3.075 $Y=2.595 $X2=0
+ $Y2=0
cc_405 N_A_584_21#_M1004_g N_VPWR_c_819_n 0.00840199f $X=6.14 $Y=2.595 $X2=0
+ $Y2=0
cc_406 N_A_584_21#_M1015_d N_VPWR_c_810_n 0.00339068f $X=3.805 $Y=2.095 $X2=0
+ $Y2=0
cc_407 N_A_584_21#_M1001_g N_VPWR_c_810_n 0.00738073f $X=3.075 $Y=2.595 $X2=0
+ $Y2=0
cc_408 N_A_584_21#_M1004_g N_VPWR_c_810_n 0.00761444f $X=6.14 $Y=2.595 $X2=0
+ $Y2=0
cc_409 N_A_584_21#_M1011_g N_VGND_c_920_n 0.00486043f $X=2.995 $Y=0.445 $X2=0
+ $Y2=0
cc_410 N_A_584_21#_M1011_g N_VGND_c_921_n 0.0113055f $X=2.995 $Y=0.445 $X2=0
+ $Y2=0
cc_411 N_A_584_21#_c_432_n N_VGND_c_921_n 0.0133459f $X=4.195 $Y=0.47 $X2=0
+ $Y2=0
cc_412 N_A_584_21#_c_423_n N_VGND_c_922_n 0.00159256f $X=5.835 $Y=1.42 $X2=0
+ $Y2=0
cc_413 N_A_584_21#_c_427_n N_VGND_c_922_n 0.0123493f $X=4.67 $Y=0.59 $X2=0 $Y2=0
cc_414 N_A_584_21#_c_428_n N_VGND_c_922_n 0.0365362f $X=4.755 $Y=1.965 $X2=0
+ $Y2=0
cc_415 N_A_584_21#_c_427_n N_VGND_c_925_n 0.016357f $X=4.67 $Y=0.59 $X2=0 $Y2=0
cc_416 N_A_584_21#_c_432_n N_VGND_c_925_n 0.0225281f $X=4.195 $Y=0.47 $X2=0
+ $Y2=0
cc_417 N_A_584_21#_M1023_d N_VGND_c_929_n 0.00233022f $X=3.89 $Y=0.235 $X2=0
+ $Y2=0
cc_418 N_A_584_21#_M1011_g N_VGND_c_929_n 0.00533746f $X=2.995 $Y=0.445 $X2=0
+ $Y2=0
cc_419 N_A_584_21#_c_423_n N_VGND_c_929_n 0.00393927f $X=5.835 $Y=1.42 $X2=0
+ $Y2=0
cc_420 N_A_584_21#_c_427_n N_VGND_c_929_n 0.0206562f $X=4.67 $Y=0.59 $X2=0 $Y2=0
cc_421 N_A_584_21#_c_432_n N_VGND_c_929_n 0.0143225f $X=4.195 $Y=0.47 $X2=0
+ $Y2=0
cc_422 N_A_584_21#_c_428_n A_923_185# 0.00721863f $X=4.755 $Y=1.965 $X2=-0.19
+ $Y2=-0.245
cc_423 N_A_352_419#_M1023_g N_CLK_c_688_n 0.0022372f $X=3.815 $Y=0.445 $X2=-0.19
+ $Y2=-0.245
cc_424 N_A_352_419#_c_591_n N_VPWR_M1001_d 0.00265118f $X=3.43 $Y=2.205 $X2=0
+ $Y2=0
cc_425 N_A_352_419#_M1015_g N_VPWR_c_812_n 0.00446878f $X=3.68 $Y=2.595 $X2=0
+ $Y2=0
cc_426 N_A_352_419#_M1015_g N_VPWR_c_817_n 0.00710941f $X=3.68 $Y=2.595 $X2=0
+ $Y2=0
cc_427 N_A_352_419#_M1018_d N_VPWR_c_810_n 0.00738611f $X=1.76 $Y=2.095 $X2=0
+ $Y2=0
cc_428 N_A_352_419#_M1015_g N_VPWR_c_810_n 0.0104338f $X=3.68 $Y=2.595 $X2=0
+ $Y2=0
cc_429 N_A_352_419#_c_591_n A_526_419# 0.00227802f $X=3.43 $Y=2.205 $X2=-0.19
+ $Y2=-0.245
cc_430 N_A_352_419#_c_598_n N_VGND_c_920_n 0.0561134f $X=2.6 $Y=0.4 $X2=0 $Y2=0
cc_431 N_A_352_419#_M1019_g N_VGND_c_921_n 0.0116168f $X=3.425 $Y=0.445 $X2=0
+ $Y2=0
cc_432 N_A_352_419#_M1023_g N_VGND_c_921_n 0.00225635f $X=3.815 $Y=0.445 $X2=0
+ $Y2=0
cc_433 N_A_352_419#_c_598_n N_VGND_c_921_n 0.0154068f $X=2.6 $Y=0.4 $X2=0 $Y2=0
cc_434 N_A_352_419#_c_584_n N_VGND_c_921_n 0.0050777f $X=2.685 $Y=0.815 $X2=0
+ $Y2=0
cc_435 N_A_352_419#_c_586_n N_VGND_c_921_n 0.0211032f $X=3.465 $Y=0.98 $X2=0
+ $Y2=0
cc_436 N_A_352_419#_M1019_g N_VGND_c_925_n 0.00486043f $X=3.425 $Y=0.445 $X2=0
+ $Y2=0
cc_437 N_A_352_419#_M1023_g N_VGND_c_925_n 0.00465161f $X=3.815 $Y=0.445 $X2=0
+ $Y2=0
cc_438 N_A_352_419#_M1010_d N_VGND_c_929_n 0.00223855f $X=1.81 $Y=0.235 $X2=0
+ $Y2=0
cc_439 N_A_352_419#_M1019_g N_VGND_c_929_n 0.00444995f $X=3.425 $Y=0.445 $X2=0
+ $Y2=0
cc_440 N_A_352_419#_M1023_g N_VGND_c_929_n 0.00929057f $X=3.815 $Y=0.445 $X2=0
+ $Y2=0
cc_441 N_A_352_419#_c_598_n N_VGND_c_929_n 0.0364096f $X=2.6 $Y=0.4 $X2=0 $Y2=0
cc_442 N_A_352_419#_c_586_n N_VGND_c_929_n 0.0187417f $X=3.465 $Y=0.98 $X2=0
+ $Y2=0
cc_443 N_A_352_419#_c_588_n N_VGND_c_929_n 0.00150475f $X=3.565 $Y=0.98 $X2=0
+ $Y2=0
cc_444 N_A_352_419#_c_598_n A_448_47# 0.0210199f $X=2.6 $Y=0.4 $X2=-0.19
+ $Y2=-0.245
cc_445 N_A_352_419#_c_584_n A_448_47# 0.00391905f $X=2.685 $Y=0.815 $X2=-0.19
+ $Y2=-0.245
cc_446 N_CLK_M1008_g N_A_1147_419#_c_768_n 0.0135525f $X=5.61 $Y=2.595 $X2=0
+ $Y2=0
cc_447 N_CLK_c_692_n N_A_1147_419#_c_748_n 0.00149342f $X=5.445 $Y=1.455 $X2=0
+ $Y2=0
cc_448 N_CLK_M1020_g N_VPWR_c_813_n 0.0204786f $X=5.08 $Y=2.595 $X2=0 $Y2=0
cc_449 N_CLK_M1008_g N_VPWR_c_813_n 0.0194516f $X=5.61 $Y=2.595 $X2=0 $Y2=0
cc_450 N_CLK_M1008_g N_VPWR_c_814_n 0.00104821f $X=5.61 $Y=2.595 $X2=0 $Y2=0
cc_451 N_CLK_M1020_g N_VPWR_c_817_n 0.0083914f $X=5.08 $Y=2.595 $X2=0 $Y2=0
cc_452 N_CLK_M1008_g N_VPWR_c_819_n 0.00840199f $X=5.61 $Y=2.595 $X2=0 $Y2=0
cc_453 N_CLK_M1020_g N_VPWR_c_810_n 0.0148509f $X=5.08 $Y=2.595 $X2=0 $Y2=0
cc_454 N_CLK_M1008_g N_VPWR_c_810_n 0.0136033f $X=5.61 $Y=2.595 $X2=0 $Y2=0
cc_455 N_CLK_c_691_n N_VGND_c_922_n 0.00799283f $X=5.015 $Y=1.455 $X2=0 $Y2=0
cc_456 N_CLK_c_692_n N_VGND_c_922_n 0.010581f $X=5.445 $Y=1.455 $X2=0 $Y2=0
cc_457 CLK N_VGND_c_922_n 0.0207973f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_458 N_CLK_c_694_n N_VGND_c_922_n 0.00270827f $X=5.445 $Y=1.707 $X2=0 $Y2=0
cc_459 N_CLK_c_691_n N_VGND_c_929_n 0.00330899f $X=5.015 $Y=1.455 $X2=0 $Y2=0
cc_460 N_CLK_c_692_n N_VGND_c_929_n 0.00330899f $X=5.445 $Y=1.455 $X2=0 $Y2=0
cc_461 N_A_1147_419#_c_759_n N_VPWR_M1004_d 0.00792101f $X=6.485 $Y=2.4 $X2=0
+ $Y2=0
cc_462 N_A_1147_419#_c_747_n N_VPWR_M1004_d 0.00252199f $X=6.57 $Y=2.315 $X2=0
+ $Y2=0
cc_463 N_A_1147_419#_c_768_n N_VPWR_c_813_n 0.0500898f $X=5.875 $Y=2.48 $X2=0
+ $Y2=0
cc_464 N_A_1147_419#_M1021_g N_VPWR_c_814_n 0.0131682f $X=6.67 $Y=2.595 $X2=0
+ $Y2=0
cc_465 N_A_1147_419#_c_759_n N_VPWR_c_814_n 0.0159804f $X=6.485 $Y=2.4 $X2=0
+ $Y2=0
cc_466 N_A_1147_419#_c_768_n N_VPWR_c_814_n 0.0263563f $X=5.875 $Y=2.48 $X2=0
+ $Y2=0
cc_467 N_A_1147_419#_c_768_n N_VPWR_c_819_n 0.0177952f $X=5.875 $Y=2.48 $X2=0
+ $Y2=0
cc_468 N_A_1147_419#_M1021_g N_VPWR_c_820_n 0.008763f $X=6.67 $Y=2.595 $X2=0
+ $Y2=0
cc_469 N_A_1147_419#_M1008_d N_VPWR_c_810_n 0.00223819f $X=5.735 $Y=2.095 $X2=0
+ $Y2=0
cc_470 N_A_1147_419#_M1021_g N_VPWR_c_810_n 0.0128187f $X=6.67 $Y=2.595 $X2=0
+ $Y2=0
cc_471 N_A_1147_419#_c_759_n N_VPWR_c_810_n 0.00926284f $X=6.485 $Y=2.4 $X2=0
+ $Y2=0
cc_472 N_A_1147_419#_c_768_n N_VPWR_c_810_n 0.0123247f $X=5.875 $Y=2.48 $X2=0
+ $Y2=0
cc_473 N_A_1147_419#_M1002_g N_GCLK_c_896_n 0.00111532f $X=6.345 $Y=0.445 $X2=0
+ $Y2=0
cc_474 N_A_1147_419#_M1006_g N_GCLK_c_896_n 0.00851821f $X=6.705 $Y=0.445 $X2=0
+ $Y2=0
cc_475 N_A_1147_419#_c_743_n N_GCLK_c_896_n 0.00148461f $X=6.705 $Y=0.98 $X2=0
+ $Y2=0
cc_476 N_A_1147_419#_M1021_g GCLK 0.0102259f $X=6.67 $Y=2.595 $X2=0 $Y2=0
cc_477 N_A_1147_419#_c_747_n GCLK 0.0186519f $X=6.57 $Y=2.315 $X2=0 $Y2=0
cc_478 N_A_1147_419#_M1021_g N_GCLK_c_897_n 0.00797605f $X=6.67 $Y=2.595 $X2=0
+ $Y2=0
cc_479 N_A_1147_419#_M1006_g N_GCLK_c_897_n 0.00792544f $X=6.705 $Y=0.445 $X2=0
+ $Y2=0
cc_480 N_A_1147_419#_c_743_n N_GCLK_c_897_n 0.0162675f $X=6.705 $Y=0.98 $X2=0
+ $Y2=0
cc_481 N_A_1147_419#_c_746_n N_GCLK_c_897_n 0.0127439f $X=6.622 $Y=1.075 $X2=0
+ $Y2=0
cc_482 N_A_1147_419#_c_763_n N_GCLK_c_897_n 0.0353931f $X=6.622 $Y=1.438 $X2=0
+ $Y2=0
cc_483 N_A_1147_419#_c_747_n N_GCLK_c_897_n 0.0167459f $X=6.57 $Y=2.315 $X2=0
+ $Y2=0
cc_484 N_A_1147_419#_c_748_n N_VGND_c_922_n 0.0117218f $X=6.05 $Y=0.99 $X2=0
+ $Y2=0
cc_485 N_A_1147_419#_M1002_g N_VGND_c_924_n 0.014372f $X=6.345 $Y=0.445 $X2=0
+ $Y2=0
cc_486 N_A_1147_419#_M1006_g N_VGND_c_924_n 0.00239794f $X=6.705 $Y=0.445 $X2=0
+ $Y2=0
cc_487 N_A_1147_419#_c_745_n N_VGND_c_924_n 0.00519083f $X=6.485 $Y=0.99 $X2=0
+ $Y2=0
cc_488 N_A_1147_419#_c_748_n N_VGND_c_924_n 0.0182348f $X=6.05 $Y=0.99 $X2=0
+ $Y2=0
cc_489 N_A_1147_419#_M1002_g N_VGND_c_928_n 0.00486043f $X=6.345 $Y=0.445 $X2=0
+ $Y2=0
cc_490 N_A_1147_419#_M1006_g N_VGND_c_928_n 0.00549284f $X=6.705 $Y=0.445 $X2=0
+ $Y2=0
cc_491 N_A_1147_419#_M1002_g N_VGND_c_929_n 0.00814425f $X=6.345 $Y=0.445 $X2=0
+ $Y2=0
cc_492 N_A_1147_419#_M1006_g N_VGND_c_929_n 0.010905f $X=6.705 $Y=0.445 $X2=0
+ $Y2=0
cc_493 N_VPWR_c_810_n A_254_419# 0.010279f $X=6.96 $Y=3.33 $X2=-0.19 $Y2=-0.245
cc_494 N_VPWR_c_810_n A_526_419# 0.00376744f $X=6.96 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_495 N_VPWR_c_810_n N_GCLK_M1021_d 0.0039349f $X=6.96 $Y=3.33 $X2=0 $Y2=0
cc_496 N_VPWR_c_820_n GCLK 0.0172394f $X=6.96 $Y=3.33 $X2=0 $Y2=0
cc_497 N_VPWR_c_810_n GCLK 0.0101763f $X=6.96 $Y=3.33 $X2=0 $Y2=0
cc_498 N_GCLK_c_896_n N_VGND_c_924_n 0.0137946f $X=6.92 $Y=0.47 $X2=0 $Y2=0
cc_499 N_GCLK_c_896_n N_VGND_c_928_n 0.0211775f $X=6.92 $Y=0.47 $X2=0 $Y2=0
cc_500 N_GCLK_M1006_d N_VGND_c_929_n 0.00232985f $X=6.78 $Y=0.235 $X2=0 $Y2=0
cc_501 N_GCLK_c_896_n N_VGND_c_929_n 0.0134544f $X=6.92 $Y=0.47 $X2=0 $Y2=0
cc_502 A_110_47# N_VGND_c_929_n 0.00268865f $X=0.55 $Y=0.235 $X2=6.96 $Y2=0
cc_503 N_VGND_c_929_n A_284_47# 0.00307274f $X=6.96 $Y=0 $X2=-0.19 $Y2=-0.245
cc_504 N_VGND_c_929_n A_448_47# 0.00651211f $X=6.96 $Y=0 $X2=-0.19 $Y2=-0.245
cc_505 N_VGND_c_929_n A_700_47# 0.00611671f $X=6.96 $Y=0 $X2=-0.19 $Y2=-0.245
cc_506 N_VGND_c_929_n A_1284_47# 0.00899413f $X=6.96 $Y=0 $X2=-0.19 $Y2=-0.245
