# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_sc_lp__ebufn_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_lp__ebufn_8 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.600000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.705000 1.180000 9.035000 1.515000 ;
    END
  END A
  PIN TE_B
    ANTENNAGATEAREA  1.827000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.805000 1.180000 8.195000 1.515000 ;
    END
  END TE_B
  PIN Z
    ANTENNADIFFAREA  2.352000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.180000 0.835000 1.410000 ;
        RECT 0.545000 0.595000 0.875000 0.975000 ;
        RECT 0.545000 0.975000 3.455000 1.145000 ;
        RECT 0.545000 1.145000 0.835000 1.180000 ;
        RECT 0.625000 1.410000 0.795000 1.815000 ;
        RECT 0.625000 1.815000 3.455000 1.985000 ;
        RECT 0.625000 1.985000 0.795000 2.735000 ;
        RECT 1.405000 0.595000 1.735000 0.975000 ;
        RECT 1.405000 1.985000 1.735000 2.735000 ;
        RECT 2.265000 0.595000 2.595000 0.975000 ;
        RECT 2.265000 1.985000 2.595000 2.735000 ;
        RECT 3.125000 0.595000 3.455000 0.975000 ;
        RECT 3.125000 1.985000 3.455000 2.735000 ;
    END
  END Z
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 9.600000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.000000 0.000000 9.600000 0.245000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.655000 9.790000 3.520000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 9.600000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 9.600000 0.085000 ;
      RECT 0.000000  3.245000 9.600000 3.415000 ;
      RECT 0.115000  0.255000 3.805000 0.425000 ;
      RECT 0.115000  0.425000 0.365000 1.010000 ;
      RECT 0.115000  1.815000 0.445000 2.905000 ;
      RECT 0.115000  2.905000 3.805000 3.075000 ;
      RECT 0.975000  2.155000 1.225000 2.905000 ;
      RECT 1.055000  0.425000 1.225000 0.805000 ;
      RECT 1.095000  1.315000 3.465000 1.475000 ;
      RECT 1.095000  1.475000 6.725000 1.645000 ;
      RECT 1.915000  0.425000 2.085000 0.805000 ;
      RECT 1.915000  2.155000 2.085000 2.905000 ;
      RECT 2.775000  0.425000 2.945000 0.805000 ;
      RECT 2.775000  2.155000 2.945000 2.905000 ;
      RECT 3.635000  0.425000 3.805000 1.135000 ;
      RECT 3.635000  1.135000 7.245000 1.305000 ;
      RECT 3.635000  1.815000 6.385000 1.985000 ;
      RECT 3.635000  1.985000 3.805000 2.905000 ;
      RECT 3.985000  0.085000 4.235000 0.965000 ;
      RECT 3.985000  2.155000 4.235000 3.245000 ;
      RECT 4.415000  0.255000 4.745000 1.135000 ;
      RECT 4.415000  1.985000 4.745000 3.075000 ;
      RECT 4.925000  0.085000 5.095000 0.965000 ;
      RECT 4.925000  2.155000 5.095000 3.245000 ;
      RECT 5.275000  0.295000 5.605000 1.135000 ;
      RECT 5.275000  1.985000 5.605000 3.075000 ;
      RECT 5.785000  0.085000 5.955000 0.965000 ;
      RECT 5.785000  2.155000 5.955000 3.245000 ;
      RECT 6.135000  0.255000 6.465000 1.135000 ;
      RECT 6.135000  1.985000 6.385000 2.365000 ;
      RECT 6.135000  2.365000 7.325000 2.535000 ;
      RECT 6.135000  2.535000 6.385000 3.075000 ;
      RECT 6.555000  1.645000 6.725000 2.025000 ;
      RECT 6.555000  2.025000 7.665000 2.195000 ;
      RECT 6.565000  2.705000 6.815000 3.245000 ;
      RECT 6.645000  0.085000 6.815000 0.965000 ;
      RECT 6.995000  0.255000 7.245000 1.135000 ;
      RECT 6.995000  2.535000 7.325000 3.075000 ;
      RECT 7.415000  0.255000 8.165000 1.010000 ;
      RECT 7.415000  1.010000 7.635000 1.685000 ;
      RECT 7.415000  1.685000 8.165000 1.855000 ;
      RECT 7.495000  2.195000 7.665000 2.315000 ;
      RECT 7.495000  2.315000 9.025000 2.485000 ;
      RECT 7.835000  1.855000 8.165000 2.145000 ;
      RECT 8.265000  2.655000 8.515000 3.245000 ;
      RECT 8.345000  0.085000 8.515000 0.670000 ;
      RECT 8.365000  0.840000 9.025000 1.010000 ;
      RECT 8.365000  1.010000 8.535000 1.815000 ;
      RECT 8.365000  1.815000 9.025000 2.315000 ;
      RECT 8.695000  0.255000 9.025000 0.840000 ;
      RECT 8.695000  2.485000 9.025000 3.075000 ;
      RECT 9.205000  0.085000 9.455000 1.095000 ;
      RECT 9.205000  1.815000 9.455000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
      RECT 8.315000 -0.085000 8.485000 0.085000 ;
      RECT 8.315000  3.245000 8.485000 3.415000 ;
      RECT 8.795000 -0.085000 8.965000 0.085000 ;
      RECT 8.795000  3.245000 8.965000 3.415000 ;
      RECT 9.275000 -0.085000 9.445000 0.085000 ;
      RECT 9.275000  3.245000 9.445000 3.415000 ;
  END
END sky130_fd_sc_lp__ebufn_8
END LIBRARY
