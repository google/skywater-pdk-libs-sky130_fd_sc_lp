# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__bufinv_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_lp__bufinv_8 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.240000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.315000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.750000 1.210000 6.155000 1.800000 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  2.352000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.095000 1.160000 3.410000 1.225000 ;
        RECT 0.095000 1.225000 0.815000 1.755000 ;
        RECT 0.095000 1.755000 3.410000 1.925000 ;
        RECT 0.570000 0.255000 0.830000 1.055000 ;
        RECT 0.570000 1.055000 3.410000 1.160000 ;
        RECT 0.570000 1.925000 0.830000 3.055000 ;
        RECT 1.430000 0.255000 1.690000 1.055000 ;
        RECT 1.430000 1.925000 1.690000 3.055000 ;
        RECT 2.290000 0.255000 2.550000 1.055000 ;
        RECT 2.290000 1.925000 2.550000 3.055000 ;
        RECT 3.150000 0.255000 3.410000 1.055000 ;
        RECT 3.150000 1.925000 3.410000 3.055000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 6.240000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 6.240000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.240000 0.085000 ;
      RECT 0.000000  3.245000 6.240000 3.415000 ;
      RECT 0.105000  0.085000 0.400000 0.990000 ;
      RECT 0.105000  2.095000 0.400000 3.245000 ;
      RECT 0.985000  1.395000 4.210000 1.585000 ;
      RECT 1.000000  0.085000 1.260000 0.885000 ;
      RECT 1.000000  2.095000 1.260000 3.245000 ;
      RECT 1.860000  0.085000 2.120000 0.885000 ;
      RECT 1.860000  2.095000 2.120000 3.245000 ;
      RECT 2.720000  0.085000 2.980000 0.885000 ;
      RECT 2.720000  2.095000 2.980000 3.245000 ;
      RECT 3.580000  0.085000 3.860000 1.070000 ;
      RECT 3.580000  1.840000 3.870000 3.245000 ;
      RECT 4.030000  0.255000 4.335000 1.055000 ;
      RECT 4.030000  1.055000 5.195000 1.225000 ;
      RECT 4.030000  1.225000 4.210000 1.395000 ;
      RECT 4.040000  1.585000 4.210000 1.755000 ;
      RECT 4.040000  1.755000 5.195000 1.925000 ;
      RECT 4.040000  1.925000 4.375000 3.055000 ;
      RECT 4.380000  1.395000 5.555000 1.585000 ;
      RECT 4.505000  0.085000 4.835000 0.885000 ;
      RECT 4.545000  2.095000 4.800000 3.245000 ;
      RECT 4.970000  1.925000 5.195000 3.055000 ;
      RECT 5.005000  0.255000 5.195000 1.055000 ;
      RECT 5.365000  0.085000 5.695000 0.700000 ;
      RECT 5.365000  2.310000 5.695000 3.245000 ;
      RECT 5.385000  0.870000 6.145000 1.040000 ;
      RECT 5.385000  1.040000 5.555000 1.395000 ;
      RECT 5.385000  1.585000 5.555000 1.970000 ;
      RECT 5.385000  1.970000 6.125000 2.140000 ;
      RECT 5.865000  0.255000 6.145000 0.870000 ;
      RECT 5.865000  2.140000 6.125000 3.055000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
  END
END sky130_fd_sc_lp__bufinv_8
END LIBRARY
