* File: sky130_fd_sc_lp__edfxbp_1.spice
* Created: Fri Aug 28 10:32:25 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__edfxbp_1.pex.spice"
.subckt sky130_fd_sc_lp__edfxbp_1  VNB VPB DE D CLK VPWR Q_N Q VGND
* 
* VGND	VGND
* Q	Q
* Q_N	Q_N
* VPWR	VPWR
* CLK	CLK
* D	D
* DE	DE
* VPB	VPB
* VNB	VNB
MM1007 N_A_120_179#_M1007_d N_DE_M1007_g N_VGND_M1007_s VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.1197 PD=1.41 PS=1.41 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1022 N_VGND_M1022_d N_DE_M1022_g N_A_231_53#_M1022_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.1197 PD=0.7 PS=1.41 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1002 N_A_404_53#_M1002_d N_A_120_179#_M1002_g N_VGND_M1022_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1197 AS=0.0588 PD=1.41 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1029 N_A_531_423#_M1029_d N_D_M1029_g N_A_231_53#_M1029_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0588 AS=0.1197 PD=0.7 PS=1.41 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1017 N_A_404_53#_M1017_d N_A_587_350#_M1017_g N_A_531_423#_M1029_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.1533 AS=0.0588 PD=1.57 PS=0.7 NRD=22.848 NRS=0 M=1 R=2.8
+ SA=75000.6 SB=75000.3 A=0.063 P=1.14 MULT=1
MM1013 N_A_902_396#_M1013_d N_A_872_324#_M1013_g N_A_531_423#_M1013_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.0672 AS=0.1365 PD=0.74 PS=1.49 NRD=11.424 NRS=11.424 M=1
+ R=2.8 SA=75000.2 SB=75001.8 A=0.063 P=1.14 MULT=1
MM1011 A_1004_91# N_A_958_290#_M1011_g N_A_902_396#_M1013_d VNB NSHORT L=0.15
+ W=0.42 AD=0.06615 AS=0.0672 PD=0.735 PS=0.74 NRD=29.28 NRS=0 M=1 R=2.8
+ SA=75000.7 SB=75001.3 A=0.063 P=1.14 MULT=1
MM1014 N_VGND_M1014_d N_A_1067_65#_M1014_g A_1004_91# VNB NSHORT L=0.15 W=0.42
+ AD=0.10084 AS=0.06615 PD=0.883585 PS=0.735 NRD=0 NRS=29.28 M=1 R=2.8
+ SA=75001.2 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1035 N_A_1067_65#_M1035_d N_A_902_396#_M1035_g N_VGND_M1014_d VNB NSHORT
+ L=0.15 W=0.64 AD=0.1824 AS=0.15366 PD=1.85 PS=1.34642 NRD=0 NRS=36.552 M=1
+ R=4.26667 SA=75001.2 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1018 N_VGND_M1018_d N_CLK_M1018_g N_A_872_324#_M1018_s VNB NSHORT L=0.15
+ W=0.42 AD=0.1155 AS=0.168 PD=0.97 PS=1.64 NRD=54.276 NRS=32.856 M=1 R=2.8
+ SA=75000.3 SB=75000.9 A=0.063 P=1.14 MULT=1
MM1032 N_A_958_290#_M1032_d N_A_872_324#_M1032_g N_VGND_M1018_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.1197 AS=0.1155 PD=1.41 PS=0.97 NRD=0 NRS=22.848 M=1 R=2.8
+ SA=75001 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1020 N_A_1865_367#_M1020_d N_A_872_324#_M1020_g N_A_1789_141#_M1020_s VNB
+ NSHORT L=0.15 W=0.42 AD=0.0966 AS=0.1197 PD=0.826667 PS=1.41 NRD=49.992 NRS=0
+ M=1 R=2.8 SA=75000.2 SB=75002.1 A=0.063 P=1.14 MULT=1
MM1006 A_1986_57# N_A_958_290#_M1006_g N_A_1865_367#_M1020_d VNB NSHORT L=0.15
+ W=0.84 AD=0.1092 AS=0.1932 PD=1.1 PS=1.65333 NRD=10.704 NRS=0.708 M=1 R=5.6
+ SA=75000.5 SB=75001.2 A=0.126 P=1.98 MULT=1
MM1028 N_VGND_M1028_d N_A_1067_65#_M1028_g A_1986_57# VNB NSHORT L=0.15 W=0.84
+ AD=0.3412 AS=0.1092 PD=2.27333 PS=1.1 NRD=17.136 NRS=10.704 M=1 R=5.6
+ SA=75000.9 SB=75000.7 A=0.126 P=1.98 MULT=1
MM1016 N_A_1789_141#_M1016_d N_A_587_350#_M1016_g N_VGND_M1028_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.1617 AS=0.1706 PD=1.61 PS=1.13667 NRD=31.428 NRS=100.332
+ M=1 R=2.8 SA=75002 SB=75000.3 A=0.063 P=1.14 MULT=1
MM1024 N_VGND_M1024_d N_A_1865_367#_M1024_g N_A_587_350#_M1024_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.1272 AS=0.1155 PD=0.953333 PS=1.39 NRD=70.812 NRS=0 M=1
+ R=2.8 SA=75000.2 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1000 N_Q_N_M1000_d N_A_587_350#_M1000_g N_VGND_M1024_d VNB NSHORT L=0.15
+ W=0.84 AD=0.231 AS=0.2544 PD=2.23 PS=1.90667 NRD=0 NRS=12.132 M=1 R=5.6
+ SA=75000.5 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1012 N_Q_M1012_d N_A_1865_367#_M1012_g N_VGND_M1012_s VNB NSHORT L=0.15 W=0.84
+ AD=0.231 AS=0.3556 PD=2.23 PS=2.66 NRD=0 NRS=17.136 M=1 R=5.6 SA=75000.3
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1001 N_A_120_179#_M1001_d N_DE_M1001_g N_VPWR_M1001_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1824 AS=0.1824 PD=1.85 PS=1.85 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1005 N_VPWR_M1005_d N_DE_M1005_g N_A_286_423#_M1005_s VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0588 AS=0.1197 PD=0.7 PS=1.41 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1026 A_459_423# N_A_120_179#_M1026_g N_VPWR_M1005_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=23.443 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1025 N_A_531_423#_M1025_d N_D_M1025_g A_459_423# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=23.443 M=1 R=2.8 SA=75001
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1003 N_A_286_423#_M1003_d N_A_587_350#_M1003_g N_A_531_423#_M1025_d VPB
+ PHIGHVT L=0.15 W=0.42 AD=0.1197 AS=0.0588 PD=1.41 PS=0.7 NRD=0 NRS=0 M=1 R=2.8
+ SA=75001.4 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1008 N_A_902_396#_M1008_d N_A_872_324#_M1008_g N_A_761_396#_M1008_s VPB
+ PHIGHVT L=0.15 W=0.42 AD=0.0588 AS=0.2331 PD=0.7 PS=1.95 NRD=0 NRS=126.632 M=1
+ R=2.8 SA=75000.5 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1033 N_A_531_423#_M1033_d N_A_958_290#_M1033_g N_A_902_396#_M1008_d VPB
+ PHIGHVT L=0.15 W=0.42 AD=0.1134 AS=0.0588 PD=1.38 PS=0.7 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.9 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1027 N_VPWR_M1027_d N_A_1067_65#_M1027_g N_A_761_396#_M1027_s VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.0924 AS=0.1134 PD=0.816667 PS=1.38 NRD=49.25 NRS=0 M=1
+ R=2.8 SA=75000.2 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1015 N_A_1067_65#_M1015_d N_A_902_396#_M1015_g N_VPWR_M1027_d VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.2268 AS=0.1848 PD=2.22 PS=1.63333 NRD=0 NRS=0 M=1 R=5.6
+ SA=75000.5 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1023 N_VPWR_M1023_d N_CLK_M1023_g N_A_872_324#_M1023_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.2624 AS=0.1728 PD=1.46 PS=1.82 NRD=83.0946 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75001.2 A=0.096 P=1.58 MULT=1
MM1021 N_A_958_290#_M1021_d N_A_872_324#_M1021_g N_VPWR_M1023_d VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.1728 AS=0.2624 PD=1.82 PS=1.46 NRD=0 NRS=83.0946 M=1
+ R=4.26667 SA=75001.2 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1030 N_A_1865_367#_M1030_d N_A_872_324#_M1030_g N_A_1781_367#_M1030_s VPB
+ PHIGHVT L=0.15 W=1.26 AD=0.2898 AS=0.3402 PD=2.46 PS=3.06 NRD=0 NRS=0 M=1
+ R=8.4 SA=75000.2 SB=75000.4 A=0.189 P=2.82 MULT=1
MM1004 N_A_1971_388#_M1004_d N_A_958_290#_M1004_g N_A_1865_367#_M1030_d VPB
+ PHIGHVT L=0.15 W=0.42 AD=0.1134 AS=0.0966 PD=1.38 PS=0.82 NRD=0 NRS=82.0702
+ M=1 R=2.8 SA=75000.7 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1009 N_VPWR_M1009_d N_A_1067_65#_M1009_g N_A_1781_367#_M1009_s VPB PHIGHVT
+ L=0.15 W=1.26 AD=0.29925 AS=0.3402 PD=2.475 PS=3.06 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.2 SB=75000.4 A=0.189 P=2.82 MULT=1
MM1019 N_A_1971_388#_M1019_d N_A_587_350#_M1019_g N_VPWR_M1009_d VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.1806 AS=0.09975 PD=1.7 PS=0.825 NRD=75.0373 NRS=85.5965 M=1
+ R=2.8 SA=75000.7 SB=75000.4 A=0.063 P=1.14 MULT=1
MM1034 N_VPWR_M1034_d N_A_1865_367#_M1034_g N_A_587_350#_M1034_s VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.142552 AS=0.1728 PD=1.11158 PS=1.82 NRD=51.614 NRS=0 M=1
+ R=4.26667 SA=75000.2 SB=75000.7 A=0.096 P=1.58 MULT=1
MM1010 N_Q_N_M1010_d N_A_587_350#_M1010_g N_VPWR_M1034_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3528 AS=0.280648 PD=3.08 PS=2.18842 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.5 SB=75000.2 A=0.189 P=2.82 MULT=1
MM1031 N_Q_M1031_d N_A_1865_367#_M1031_g N_VPWR_M1031_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3402 AS=0.3528 PD=3.06 PS=3.08 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX36_noxref VNB VPB NWDIODE A=27.5967 P=33.33
c_135 VNB 0 1.25302e-19 $X=0 $Y=0
*
.include "sky130_fd_sc_lp__edfxbp_1.pxi.spice"
*
.ends
*
*
