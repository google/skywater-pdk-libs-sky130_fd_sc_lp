* File: sky130_fd_sc_lp__dfsbp_1.pxi.spice
* Created: Wed Sep  2 09:44:01 2020
* 
x_PM_SKY130_FD_SC_LP__DFSBP_1%CLK N_CLK_c_259_n N_CLK_M1025_g N_CLK_M1021_g
+ N_CLK_c_265_n CLK CLK CLK CLK N_CLK_c_261_n N_CLK_c_262_n CLK
+ PM_SKY130_FD_SC_LP__DFSBP_1%CLK
x_PM_SKY130_FD_SC_LP__DFSBP_1%A_111_156# N_A_111_156#_M1025_d
+ N_A_111_156#_M1021_d N_A_111_156#_c_322_n N_A_111_156#_c_293_n
+ N_A_111_156#_M1011_g N_A_111_156#_c_323_n N_A_111_156#_M1002_g
+ N_A_111_156#_M1010_g N_A_111_156#_c_295_n N_A_111_156#_c_296_n
+ N_A_111_156#_M1028_g N_A_111_156#_M1019_g N_A_111_156#_M1007_g
+ N_A_111_156#_c_326_n N_A_111_156#_c_298_n N_A_111_156#_c_328_n
+ N_A_111_156#_c_299_n N_A_111_156#_c_300_n N_A_111_156#_c_301_n
+ N_A_111_156#_c_302_n N_A_111_156#_c_303_n N_A_111_156#_c_304_n
+ N_A_111_156#_c_305_n N_A_111_156#_c_306_n N_A_111_156#_c_307_n
+ N_A_111_156#_c_308_n N_A_111_156#_c_309_n N_A_111_156#_c_310_n
+ N_A_111_156#_c_311_n N_A_111_156#_c_312_n N_A_111_156#_c_313_n
+ N_A_111_156#_c_314_n N_A_111_156#_c_315_n N_A_111_156#_c_333_n
+ N_A_111_156#_c_334_n N_A_111_156#_c_316_n N_A_111_156#_c_317_n
+ N_A_111_156#_c_318_n N_A_111_156#_c_319_n N_A_111_156#_c_320_n
+ N_A_111_156#_c_321_n PM_SKY130_FD_SC_LP__DFSBP_1%A_111_156#
x_PM_SKY130_FD_SC_LP__DFSBP_1%D N_D_M1008_g N_D_M1018_g D D D N_D_c_559_n
+ N_D_c_560_n N_D_c_563_n N_D_c_564_n PM_SKY130_FD_SC_LP__DFSBP_1%D
x_PM_SKY130_FD_SC_LP__DFSBP_1%A_708_93# N_A_708_93#_M1012_s N_A_708_93#_M1029_d
+ N_A_708_93#_c_615_n N_A_708_93#_M1023_g N_A_708_93#_c_622_n
+ N_A_708_93#_M1031_g N_A_708_93#_c_616_n N_A_708_93#_c_617_n
+ N_A_708_93#_c_623_n N_A_708_93#_c_624_n N_A_708_93#_c_618_n
+ N_A_708_93#_c_619_n N_A_708_93#_c_625_n N_A_708_93#_c_620_n
+ N_A_708_93#_c_700_p N_A_708_93#_c_662_p N_A_708_93#_c_626_n
+ N_A_708_93#_c_627_n N_A_708_93#_c_621_n N_A_708_93#_c_629_n
+ PM_SKY130_FD_SC_LP__DFSBP_1%A_708_93#
x_PM_SKY130_FD_SC_LP__DFSBP_1%A_580_119# N_A_580_119#_M1010_d
+ N_A_580_119#_M1003_d N_A_580_119#_M1012_g N_A_580_119#_c_730_n
+ N_A_580_119#_c_731_n N_A_580_119#_c_732_n N_A_580_119#_M1029_g
+ N_A_580_119#_M1026_g N_A_580_119#_c_720_n N_A_580_119#_c_721_n
+ N_A_580_119#_M1032_g N_A_580_119#_c_734_n N_A_580_119#_c_722_n
+ N_A_580_119#_c_723_n N_A_580_119#_c_767_n N_A_580_119#_c_736_n
+ N_A_580_119#_c_737_n N_A_580_119#_c_738_n N_A_580_119#_c_739_n
+ N_A_580_119#_c_724_n N_A_580_119#_c_741_n N_A_580_119#_c_742_n
+ N_A_580_119#_c_743_n N_A_580_119#_c_725_n N_A_580_119#_c_726_n
+ N_A_580_119#_c_745_n N_A_580_119#_c_727_n N_A_580_119#_c_728_n
+ N_A_580_119#_c_748_n PM_SKY130_FD_SC_LP__DFSBP_1%A_580_119#
x_PM_SKY130_FD_SC_LP__DFSBP_1%SET_B N_SET_B_M1009_g N_SET_B_c_892_n
+ N_SET_B_M1013_g N_SET_B_M1015_g N_SET_B_M1005_g N_SET_B_c_894_n
+ N_SET_B_c_911_n N_SET_B_c_899_n N_SET_B_c_1002_p N_SET_B_c_900_n
+ N_SET_B_c_901_n N_SET_B_c_902_n N_SET_B_c_903_n N_SET_B_c_904_n
+ N_SET_B_c_905_n SET_B N_SET_B_c_906_n PM_SKY130_FD_SC_LP__DFSBP_1%SET_B
x_PM_SKY130_FD_SC_LP__DFSBP_1%A_161_21# N_A_161_21#_M1011_s N_A_161_21#_M1002_s
+ N_A_161_21#_c_1018_n N_A_161_21#_c_1019_n N_A_161_21#_c_1030_n
+ N_A_161_21#_M1003_g N_A_161_21#_M1000_g N_A_161_21#_c_1021_n
+ N_A_161_21#_M1020_g N_A_161_21#_M1033_g N_A_161_21#_c_1024_n
+ N_A_161_21#_c_1025_n N_A_161_21#_c_1026_n N_A_161_21#_c_1033_n
+ N_A_161_21#_c_1027_n N_A_161_21#_c_1034_n N_A_161_21#_c_1028_n
+ N_A_161_21#_c_1035_n PM_SKY130_FD_SC_LP__DFSBP_1%A_161_21#
x_PM_SKY130_FD_SC_LP__DFSBP_1%A_1535_177# N_A_1535_177#_M1024_s
+ N_A_1535_177#_M1006_s N_A_1535_177#_M1030_g N_A_1535_177#_c_1169_n
+ N_A_1535_177#_c_1170_n N_A_1535_177#_c_1164_n N_A_1535_177#_M1016_g
+ N_A_1535_177#_c_1165_n N_A_1535_177#_c_1171_n N_A_1535_177#_c_1172_n
+ N_A_1535_177#_c_1166_n N_A_1535_177#_c_1173_n N_A_1535_177#_c_1167_n
+ PM_SKY130_FD_SC_LP__DFSBP_1%A_1535_177#
x_PM_SKY130_FD_SC_LP__DFSBP_1%A_1331_151# N_A_1331_151#_M1019_d
+ N_A_1331_151#_M1007_d N_A_1331_151#_M1015_d N_A_1331_151#_c_1256_n
+ N_A_1331_151#_M1006_g N_A_1331_151#_c_1237_n N_A_1331_151#_M1024_g
+ N_A_1331_151#_c_1238_n N_A_1331_151#_c_1257_n N_A_1331_151#_c_1239_n
+ N_A_1331_151#_M1027_g N_A_1331_151#_c_1258_n N_A_1331_151#_M1017_g
+ N_A_1331_151#_M1004_g N_A_1331_151#_c_1241_n N_A_1331_151#_M1001_g
+ N_A_1331_151#_c_1242_n N_A_1331_151#_c_1260_n N_A_1331_151#_c_1243_n
+ N_A_1331_151#_c_1244_n N_A_1331_151#_c_1245_n N_A_1331_151#_c_1246_n
+ N_A_1331_151#_c_1247_n N_A_1331_151#_c_1248_n N_A_1331_151#_c_1263_n
+ N_A_1331_151#_c_1264_n N_A_1331_151#_c_1249_n N_A_1331_151#_c_1273_n
+ N_A_1331_151#_c_1266_n N_A_1331_151#_c_1250_n N_A_1331_151#_c_1251_n
+ N_A_1331_151#_c_1268_n N_A_1331_151#_c_1252_n N_A_1331_151#_c_1269_n
+ N_A_1331_151#_c_1253_n N_A_1331_151#_c_1254_n N_A_1331_151#_c_1255_n
+ PM_SKY130_FD_SC_LP__DFSBP_1%A_1331_151#
x_PM_SKY130_FD_SC_LP__DFSBP_1%A_2005_119# N_A_2005_119#_M1027_d
+ N_A_2005_119#_M1017_d N_A_2005_119#_c_1416_n N_A_2005_119#_M1014_g
+ N_A_2005_119#_M1022_g N_A_2005_119#_c_1419_n N_A_2005_119#_c_1420_n
+ N_A_2005_119#_c_1421_n N_A_2005_119#_c_1424_n N_A_2005_119#_c_1425_n
+ N_A_2005_119#_c_1426_n N_A_2005_119#_c_1422_n
+ PM_SKY130_FD_SC_LP__DFSBP_1%A_2005_119#
x_PM_SKY130_FD_SC_LP__DFSBP_1%VPWR N_VPWR_M1021_s N_VPWR_M1002_d N_VPWR_M1031_d
+ N_VPWR_M1013_d N_VPWR_M1030_d N_VPWR_M1006_d N_VPWR_M1014_d N_VPWR_c_1480_n
+ N_VPWR_c_1481_n N_VPWR_c_1482_n N_VPWR_c_1483_n N_VPWR_c_1484_n
+ N_VPWR_c_1485_n N_VPWR_c_1486_n N_VPWR_c_1487_n N_VPWR_c_1488_n
+ N_VPWR_c_1489_n VPWR N_VPWR_c_1490_n N_VPWR_c_1491_n N_VPWR_c_1492_n
+ N_VPWR_c_1493_n N_VPWR_c_1494_n N_VPWR_c_1495_n N_VPWR_c_1479_n
+ N_VPWR_c_1497_n N_VPWR_c_1498_n N_VPWR_c_1499_n N_VPWR_c_1500_n
+ N_VPWR_c_1501_n PM_SKY130_FD_SC_LP__DFSBP_1%VPWR
x_PM_SKY130_FD_SC_LP__DFSBP_1%A_494_119# N_A_494_119#_M1008_d
+ N_A_494_119#_M1018_d N_A_494_119#_c_1626_n N_A_494_119#_c_1628_n
+ N_A_494_119#_c_1634_n N_A_494_119#_c_1644_n N_A_494_119#_c_1629_n
+ PM_SKY130_FD_SC_LP__DFSBP_1%A_494_119#
x_PM_SKY130_FD_SC_LP__DFSBP_1%Q N_Q_M1022_s N_Q_M1014_s Q Q Q Q Q
+ PM_SKY130_FD_SC_LP__DFSBP_1%Q
x_PM_SKY130_FD_SC_LP__DFSBP_1%Q_N N_Q_N_M1001_d N_Q_N_M1004_d Q_N Q_N Q_N Q_N
+ Q_N Q_N Q_N N_Q_N_c_1693_n Q_N N_Q_N_c_1696_n Q_N
+ PM_SKY130_FD_SC_LP__DFSBP_1%Q_N
x_PM_SKY130_FD_SC_LP__DFSBP_1%VGND N_VGND_M1025_s N_VGND_M1011_d N_VGND_M1023_d
+ N_VGND_M1009_d N_VGND_M1005_d N_VGND_M1024_d N_VGND_M1022_d N_VGND_c_1711_n
+ N_VGND_c_1712_n N_VGND_c_1713_n N_VGND_c_1714_n N_VGND_c_1715_n
+ N_VGND_c_1716_n N_VGND_c_1717_n N_VGND_c_1718_n N_VGND_c_1719_n
+ N_VGND_c_1720_n N_VGND_c_1721_n N_VGND_c_1722_n N_VGND_c_1723_n
+ N_VGND_c_1724_n VGND N_VGND_c_1725_n N_VGND_c_1726_n N_VGND_c_1727_n
+ N_VGND_c_1728_n N_VGND_c_1729_n N_VGND_c_1730_n N_VGND_c_1731_n
+ N_VGND_c_1732_n PM_SKY130_FD_SC_LP__DFSBP_1%VGND
x_PM_SKY130_FD_SC_LP__DFSBP_1%A_1141_125# N_A_1141_125#_M1026_d
+ N_A_1141_125#_M1020_d N_A_1141_125#_c_1841_n N_A_1141_125#_c_1842_n
+ N_A_1141_125#_c_1843_n PM_SKY130_FD_SC_LP__DFSBP_1%A_1141_125#
x_PM_SKY130_FD_SC_LP__DFSBP_1%A_1248_151# N_A_1248_151#_M1019_s
+ N_A_1248_151#_M1016_s N_A_1248_151#_c_1865_n N_A_1248_151#_c_1866_n
+ N_A_1248_151#_c_1867_n PM_SKY130_FD_SC_LP__DFSBP_1%A_1248_151#
cc_1 VNB N_CLK_c_259_n 0.0156313f $X=-0.19 $Y=-0.245 $X2=0.387 $Y2=1.813
cc_2 VNB CLK 0.0203604f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_3 VNB N_CLK_c_261_n 0.0200286f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.475
cc_4 VNB N_CLK_c_262_n 0.0215525f $X=-0.19 $Y=-0.245 $X2=0.387 $Y2=1.31
cc_5 VNB N_A_111_156#_c_293_n 0.0170642f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_6 VNB N_A_111_156#_M1010_g 0.031203f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_A_111_156#_c_295_n 0.0416966f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_111_156#_c_296_n 0.00674607f $X=-0.19 $Y=-0.245 $X2=0.387 $Y2=1.475
cc_9 VNB N_A_111_156#_M1019_g 0.0224862f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_111_156#_c_298_n 0.0113724f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=2.035
cc_11 VNB N_A_111_156#_c_299_n 0.00580853f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_111_156#_c_300_n 0.00425495f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_111_156#_c_301_n 0.0136902f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_111_156#_c_302_n 0.00199113f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_111_156#_c_303_n 0.0146334f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_111_156#_c_304_n 0.00241947f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_111_156#_c_305_n 0.00125285f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_111_156#_c_306_n 0.0039119f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_111_156#_c_307_n 0.00460341f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_111_156#_c_308_n 0.0104264f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_111_156#_c_309_n 0.00612881f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_111_156#_c_310_n 0.0147335f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_111_156#_c_311_n 0.0037109f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_111_156#_c_312_n 4.53895e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_111_156#_c_313_n 0.0159473f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_111_156#_c_314_n 0.00132304f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_111_156#_c_315_n 0.0121108f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_111_156#_c_316_n 0.00437164f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_111_156#_c_317_n 0.0021934f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_111_156#_c_318_n 0.0162393f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_111_156#_c_319_n 0.0397508f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_111_156#_c_320_n 0.00344821f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_111_156#_c_321_n 0.0181458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_D_M1008_g 0.0253393f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=1.31
cc_35 VNB N_D_c_559_n 0.00963786f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_D_c_560_n 0.0356483f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_708_93#_c_615_n 0.0161913f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=2.6
cc_38 VNB N_A_708_93#_c_616_n 0.0345737f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.95
cc_39 VNB N_A_708_93#_c_617_n 0.008862f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=2.32
cc_40 VNB N_A_708_93#_c_618_n 0.0112963f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.475
cc_41 VNB N_A_708_93#_c_619_n 0.0175407f $X=-0.19 $Y=-0.245 $X2=0.277 $Y2=1.898
cc_42 VNB N_A_708_93#_c_620_n 0.00340272f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_708_93#_c_621_n 0.0110321f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_580_119#_M1012_g 0.0307418f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_580_119#_M1026_g 0.0233217f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_580_119#_c_720_n 0.0314598f $X=-0.19 $Y=-0.245 $X2=0.387 $Y2=1.475
cc_47 VNB N_A_580_119#_c_721_n 0.00764755f $X=-0.19 $Y=-0.245 $X2=0.385
+ $Y2=1.475
cc_48 VNB N_A_580_119#_c_722_n 0.00723952f $X=-0.19 $Y=-0.245 $X2=0.257
+ $Y2=2.405
cc_49 VNB N_A_580_119#_c_723_n 5.5861e-19 $X=-0.19 $Y=-0.245 $X2=0.277 $Y2=2.02
cc_50 VNB N_A_580_119#_c_724_n 0.00157692f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_580_119#_c_725_n 0.00234902f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_580_119#_c_726_n 0.00215745f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_580_119#_c_727_n 0.00346148f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_580_119#_c_728_n 2.98278e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_SET_B_M1009_g 0.0189784f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=1.31
cc_56 VNB N_SET_B_c_892_n 0.00290174f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=1.98
cc_57 VNB N_SET_B_M1005_g 0.0719924f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_SET_B_c_894_n 0.0164262f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.475
cc_59 VNB N_A_161_21#_c_1018_n 0.0743332f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=2.6
cc_60 VNB N_A_161_21#_c_1019_n 0.144987f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_A_161_21#_M1000_g 0.0307691f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_A_161_21#_c_1021_n 0.287941f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.475
cc_63 VNB N_A_161_21#_M1020_g 0.0290823f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_A_161_21#_M1033_g 0.0122394f $X=-0.19 $Y=-0.245 $X2=0.277 $Y2=1.665
cc_65 VNB N_A_161_21#_c_1024_n 0.00749069f $X=-0.19 $Y=-0.245 $X2=0.257 $Y2=2.09
cc_66 VNB N_A_161_21#_c_1025_n 0.0190211f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_A_161_21#_c_1026_n 0.0110358f $X=-0.19 $Y=-0.245 $X2=0.277 $Y2=2.02
cc_68 VNB N_A_161_21#_c_1027_n 0.00557728f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_161_21#_c_1028_n 0.0493572f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_A_1535_177#_M1030_g 0.0249681f $X=-0.19 $Y=-0.245 $X2=0.387 $Y2=1.98
cc_71 VNB N_A_1535_177#_c_1164_n 0.0217556f $X=-0.19 $Y=-0.245 $X2=0.155
+ $Y2=1.95
cc_72 VNB N_A_1535_177#_c_1165_n 0.030063f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_A_1535_177#_c_1166_n 0.00470284f $X=-0.19 $Y=-0.245 $X2=0.277
+ $Y2=1.475
cc_74 VNB N_A_1535_177#_c_1167_n 0.0574283f $X=-0.19 $Y=-0.245 $X2=0.24
+ $Y2=2.035
cc_75 VNB N_A_1331_151#_c_1237_n 0.0184462f $X=-0.19 $Y=-0.245 $X2=0.155
+ $Y2=1.95
cc_76 VNB N_A_1331_151#_c_1238_n 0.0241336f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_A_1331_151#_c_1239_n 0.0209974f $X=-0.19 $Y=-0.245 $X2=0.387
+ $Y2=1.475
cc_78 VNB N_A_1331_151#_M1004_g 0.00483366f $X=-0.19 $Y=-0.245 $X2=0.277
+ $Y2=1.475
cc_79 VNB N_A_1331_151#_c_1241_n 0.0208735f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_A_1331_151#_c_1242_n 0.0267938f $X=-0.19 $Y=-0.245 $X2=0.257
+ $Y2=2.405
cc_81 VNB N_A_1331_151#_c_1243_n 0.0013291f $X=-0.19 $Y=-0.245 $X2=0.24
+ $Y2=2.035
cc_82 VNB N_A_1331_151#_c_1244_n 0.0263034f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_A_1331_151#_c_1245_n 0.0017313f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_A_1331_151#_c_1246_n 0.0259087f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_A_1331_151#_c_1247_n 0.0258866f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_A_1331_151#_c_1248_n 3.23103e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_A_1331_151#_c_1249_n 9.08564e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_A_1331_151#_c_1250_n 0.00269488f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_A_1331_151#_c_1251_n 0.0010728f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_A_1331_151#_c_1252_n 5.6343e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_A_1331_151#_c_1253_n 0.0232426f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_A_1331_151#_c_1254_n 0.00343755f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_93 VNB N_A_1331_151#_c_1255_n 0.0376583f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_94 VNB N_A_2005_119#_c_1416_n 0.0422023f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=2.6
cc_95 VNB N_A_2005_119#_M1014_g 0.00111396f $X=-0.19 $Y=-0.245 $X2=0.155
+ $Y2=1.21
cc_96 VNB N_A_2005_119#_M1022_g 0.0354228f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_97 VNB N_A_2005_119#_c_1419_n 0.00716485f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_98 VNB N_A_2005_119#_c_1420_n 0.0175356f $X=-0.19 $Y=-0.245 $X2=0.385
+ $Y2=1.475
cc_99 VNB N_A_2005_119#_c_1421_n 0.0577265f $X=-0.19 $Y=-0.245 $X2=0.387
+ $Y2=1.31
cc_100 VNB N_A_2005_119#_c_1422_n 0.0161277f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_101 VNB N_VPWR_c_1479_n 0.521925f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_102 VNB N_A_494_119#_c_1626_n 0.00518463f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=2.6
cc_103 VNB Q 0.0169702f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=2.6
cc_104 VNB N_Q_N_c_1693_n 0.0634031f $X=-0.19 $Y=-0.245 $X2=0.277 $Y2=1.295
cc_105 VNB N_VGND_c_1711_n 0.0117383f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.475
cc_106 VNB N_VGND_c_1712_n 0.0450037f $X=-0.19 $Y=-0.245 $X2=0.277 $Y2=1.898
cc_107 VNB N_VGND_c_1713_n 0.00737785f $X=-0.19 $Y=-0.245 $X2=0.277 $Y2=1.475
cc_108 VNB N_VGND_c_1714_n 0.0161662f $X=-0.19 $Y=-0.245 $X2=0.257 $Y2=2.105
cc_109 VNB N_VGND_c_1715_n 0.021004f $X=-0.19 $Y=-0.245 $X2=0.277 $Y2=2.02
cc_110 VNB N_VGND_c_1716_n 0.0112861f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_111 VNB N_VGND_c_1717_n 0.0219344f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_112 VNB N_VGND_c_1718_n 0.00705983f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_113 VNB N_VGND_c_1719_n 0.0419174f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_114 VNB N_VGND_c_1720_n 0.00266338f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_115 VNB N_VGND_c_1721_n 0.0358067f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_116 VNB N_VGND_c_1722_n 0.00359556f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_117 VNB N_VGND_c_1723_n 0.0770805f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_118 VNB N_VGND_c_1724_n 0.00604418f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_119 VNB N_VGND_c_1725_n 0.0314716f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_120 VNB N_VGND_c_1726_n 0.0194883f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_121 VNB N_VGND_c_1727_n 0.0491829f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_122 VNB N_VGND_c_1728_n 0.0177851f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_123 VNB N_VGND_c_1729_n 0.639426f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_124 VNB N_VGND_c_1730_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_125 VNB N_VGND_c_1731_n 0.00500104f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_126 VNB N_VGND_c_1732_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_127 VNB N_A_1141_125#_c_1841_n 0.0135945f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_128 VNB N_A_1141_125#_c_1842_n 0.0049042f $X=-0.19 $Y=-0.245 $X2=0.155
+ $Y2=1.21
cc_129 VNB N_A_1141_125#_c_1843_n 0.0291912f $X=-0.19 $Y=-0.245 $X2=0.155
+ $Y2=1.95
cc_130 VNB N_A_1248_151#_c_1865_n 0.00833653f $X=-0.19 $Y=-0.245 $X2=0.48
+ $Y2=2.6
cc_131 VNB N_A_1248_151#_c_1866_n 0.00680851f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_132 VNB N_A_1248_151#_c_1867_n 0.0059619f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_133 VPB N_CLK_c_259_n 0.0138651f $X=-0.19 $Y=1.655 $X2=0.387 $Y2=1.813
cc_134 VPB N_CLK_M1021_g 0.0329246f $X=-0.19 $Y=1.655 $X2=0.48 $Y2=2.6
cc_135 VPB N_CLK_c_265_n 0.0199276f $X=-0.19 $Y=1.655 $X2=0.387 $Y2=1.98
cc_136 VPB CLK 0.00919081f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_137 VPB CLK 0.0239333f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.95
cc_138 VPB N_A_111_156#_c_322_n 0.0393608f $X=-0.19 $Y=1.655 $X2=0.48 $Y2=2.6
cc_139 VPB N_A_111_156#_c_323_n 0.0183034f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_140 VPB N_A_111_156#_M1028_g 0.0368072f $X=-0.19 $Y=1.655 $X2=0.387 $Y2=1.31
cc_141 VPB N_A_111_156#_M1007_g 0.028459f $X=-0.19 $Y=1.655 $X2=0.257 $Y2=2.09
cc_142 VPB N_A_111_156#_c_326_n 0.0262003f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_143 VPB N_A_111_156#_c_298_n 0.0136377f $X=-0.19 $Y=1.655 $X2=0.24 $Y2=2.035
cc_144 VPB N_A_111_156#_c_328_n 0.0173508f $X=-0.19 $Y=1.655 $X2=0.277 $Y2=2.09
cc_145 VPB N_A_111_156#_c_300_n 0.0134622f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_146 VPB N_A_111_156#_c_306_n 0.00215648f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_147 VPB N_A_111_156#_c_307_n 0.0261001f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_148 VPB N_A_111_156#_c_315_n 0.00727884f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_149 VPB N_A_111_156#_c_333_n 0.0275672f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_150 VPB N_A_111_156#_c_334_n 0.0508381f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_151 VPB N_D_M1018_g 0.0216947f $X=-0.19 $Y=1.655 $X2=0.48 $Y2=2.6
cc_152 VPB N_D_c_559_n 0.0114196f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_153 VPB N_D_c_563_n 0.0330878f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.475
cc_154 VPB N_D_c_564_n 0.00667677f $X=-0.19 $Y=1.655 $X2=0.387 $Y2=1.31
cc_155 VPB N_A_708_93#_c_622_n 0.0181196f $X=-0.19 $Y=1.655 $X2=0.387 $Y2=1.98
cc_156 VPB N_A_708_93#_c_623_n 0.0182778f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_157 VPB N_A_708_93#_c_624_n 0.0119505f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_158 VPB N_A_708_93#_c_625_n 0.00545185f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_159 VPB N_A_708_93#_c_626_n 0.0391492f $X=-0.19 $Y=1.655 $X2=0.24 $Y2=2.035
cc_160 VPB N_A_708_93#_c_627_n 0.00301053f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_161 VPB N_A_708_93#_c_621_n 0.00519814f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_162 VPB N_A_708_93#_c_629_n 0.0298285f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_163 VPB N_A_580_119#_M1012_g 0.00981672f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_164 VPB N_A_580_119#_c_730_n 0.0235032f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_165 VPB N_A_580_119#_c_731_n 0.0162348f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_166 VPB N_A_580_119#_c_732_n 0.0223196f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.95
cc_167 VPB N_A_580_119#_M1032_g 0.0259422f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_168 VPB N_A_580_119#_c_734_n 0.029139f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_169 VPB N_A_580_119#_c_723_n 0.00821981f $X=-0.19 $Y=1.655 $X2=0.277 $Y2=2.02
cc_170 VPB N_A_580_119#_c_736_n 0.00719111f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_171 VPB N_A_580_119#_c_737_n 0.00828312f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_172 VPB N_A_580_119#_c_738_n 0.014051f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_173 VPB N_A_580_119#_c_739_n 0.00314372f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_174 VPB N_A_580_119#_c_724_n 0.00194635f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_175 VPB N_A_580_119#_c_741_n 0.00327496f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_176 VPB N_A_580_119#_c_742_n 0.0160594f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_177 VPB N_A_580_119#_c_743_n 0.00204504f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_178 VPB N_A_580_119#_c_725_n 0.0146517f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_179 VPB N_A_580_119#_c_745_n 0.00191969f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_180 VPB N_A_580_119#_c_727_n 0.00414615f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_181 VPB N_A_580_119#_c_728_n 0.00524104f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_182 VPB N_A_580_119#_c_748_n 0.0165848f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_183 VPB N_SET_B_c_892_n 0.0124783f $X=-0.19 $Y=1.655 $X2=0.48 $Y2=1.98
cc_184 VPB N_SET_B_M1013_g 0.0379007f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_185 VPB N_SET_B_M1015_g 0.0227367f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.95
cc_186 VPB N_SET_B_M1005_g 0.00409284f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_187 VPB N_SET_B_c_899_n 0.0170752f $X=-0.19 $Y=1.655 $X2=0.277 $Y2=1.295
cc_188 VPB N_SET_B_c_900_n 0.00349417f $X=-0.19 $Y=1.655 $X2=0.277 $Y2=1.475
cc_189 VPB N_SET_B_c_901_n 0.004369f $X=-0.19 $Y=1.655 $X2=0.277 $Y2=1.665
cc_190 VPB N_SET_B_c_902_n 0.00629059f $X=-0.19 $Y=1.655 $X2=0.257 $Y2=2.09
cc_191 VPB N_SET_B_c_903_n 0.00393528f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_192 VPB N_SET_B_c_904_n 0.0490389f $X=-0.19 $Y=1.655 $X2=0.277 $Y2=2.02
cc_193 VPB N_SET_B_c_905_n 0.0112725f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_194 VPB N_SET_B_c_906_n 0.0521473f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_195 VPB N_A_161_21#_c_1018_n 0.00969484f $X=-0.19 $Y=1.655 $X2=0.48 $Y2=2.6
cc_196 VPB N_A_161_21#_c_1030_n 0.103527f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_197 VPB N_A_161_21#_M1003_g 0.0459945f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_198 VPB N_A_161_21#_M1033_g 0.0456108f $X=-0.19 $Y=1.655 $X2=0.277 $Y2=1.665
cc_199 VPB N_A_161_21#_c_1033_n 0.00877774f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_200 VPB N_A_161_21#_c_1034_n 0.00611977f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_201 VPB N_A_161_21#_c_1035_n 0.0431413f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_202 VPB N_A_1535_177#_M1030_g 0.0486866f $X=-0.19 $Y=1.655 $X2=0.387 $Y2=1.98
cc_203 VPB N_A_1535_177#_c_1169_n 0.0693887f $X=-0.19 $Y=1.655 $X2=0.155
+ $Y2=1.21
cc_204 VPB N_A_1535_177#_c_1170_n 0.0125868f $X=-0.19 $Y=1.655 $X2=0.155
+ $Y2=1.58
cc_205 VPB N_A_1535_177#_c_1171_n 0.00533367f $X=-0.19 $Y=1.655 $X2=0.387
+ $Y2=1.31
cc_206 VPB N_A_1535_177#_c_1172_n 0.0657908f $X=-0.19 $Y=1.655 $X2=0.277
+ $Y2=1.898
cc_207 VPB N_A_1535_177#_c_1173_n 0.014562f $X=-0.19 $Y=1.655 $X2=0.257
+ $Y2=2.405
cc_208 VPB N_A_1331_151#_c_1256_n 0.0205026f $X=-0.19 $Y=1.655 $X2=0.387
+ $Y2=1.98
cc_209 VPB N_A_1331_151#_c_1257_n 0.0286753f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_210 VPB N_A_1331_151#_c_1258_n 0.0222939f $X=-0.19 $Y=1.655 $X2=0.387
+ $Y2=1.31
cc_211 VPB N_A_1331_151#_M1004_g 0.0223614f $X=-0.19 $Y=1.655 $X2=0.277
+ $Y2=1.475
cc_212 VPB N_A_1331_151#_c_1260_n 0.0126523f $X=-0.19 $Y=1.655 $X2=0.277
+ $Y2=2.02
cc_213 VPB N_A_1331_151#_c_1245_n 0.00913082f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_214 VPB N_A_1331_151#_c_1248_n 0.0151092f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_215 VPB N_A_1331_151#_c_1263_n 0.00991418f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_216 VPB N_A_1331_151#_c_1264_n 0.00600797f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_217 VPB N_A_1331_151#_c_1249_n 0.00105813f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_218 VPB N_A_1331_151#_c_1266_n 4.22143e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_219 VPB N_A_1331_151#_c_1250_n 0.0127631f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_220 VPB N_A_1331_151#_c_1268_n 0.00895171f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_221 VPB N_A_1331_151#_c_1269_n 0.00111305f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_222 VPB N_A_1331_151#_c_1253_n 0.020598f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_223 VPB N_A_2005_119#_M1014_g 0.0236393f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_224 VPB N_A_2005_119#_c_1424_n 0.0176362f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_225 VPB N_A_2005_119#_c_1425_n 0.0116642f $X=-0.19 $Y=1.655 $X2=0.277
+ $Y2=1.665
cc_226 VPB N_A_2005_119#_c_1426_n 0.00110315f $X=-0.19 $Y=1.655 $X2=0.257
+ $Y2=2.09
cc_227 VPB N_A_2005_119#_c_1422_n 0.046173f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_228 VPB N_VPWR_c_1480_n 0.0117124f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.475
cc_229 VPB N_VPWR_c_1481_n 0.0226984f $X=-0.19 $Y=1.655 $X2=0.277 $Y2=1.898
cc_230 VPB N_VPWR_c_1482_n 0.00765578f $X=-0.19 $Y=1.655 $X2=0.277 $Y2=1.475
cc_231 VPB N_VPWR_c_1483_n 0.00314922f $X=-0.19 $Y=1.655 $X2=0.257 $Y2=2.105
cc_232 VPB N_VPWR_c_1484_n 0.00368255f $X=-0.19 $Y=1.655 $X2=0.277 $Y2=2.02
cc_233 VPB N_VPWR_c_1485_n 0.0153857f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_234 VPB N_VPWR_c_1486_n 0.0250215f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_235 VPB N_VPWR_c_1487_n 4.89148e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_236 VPB N_VPWR_c_1488_n 0.046806f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_237 VPB N_VPWR_c_1489_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_238 VPB N_VPWR_c_1490_n 0.0416391f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_239 VPB N_VPWR_c_1491_n 0.0376044f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_240 VPB N_VPWR_c_1492_n 0.0439334f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_241 VPB N_VPWR_c_1493_n 0.0393781f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_242 VPB N_VPWR_c_1494_n 0.0439154f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_243 VPB N_VPWR_c_1495_n 0.0194284f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_244 VPB N_VPWR_c_1479_n 0.0979985f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_245 VPB N_VPWR_c_1497_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_246 VPB N_VPWR_c_1498_n 0.00517946f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_247 VPB N_VPWR_c_1499_n 0.0052952f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_248 VPB N_VPWR_c_1500_n 0.00352523f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_249 VPB N_VPWR_c_1501_n 0.00603306f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_250 VPB N_A_494_119#_c_1626_n 0.00225539f $X=-0.19 $Y=1.655 $X2=0.48 $Y2=2.6
cc_251 VPB N_A_494_119#_c_1628_n 0.00581012f $X=-0.19 $Y=1.655 $X2=0.387
+ $Y2=1.98
cc_252 VPB N_A_494_119#_c_1629_n 0.00234741f $X=-0.19 $Y=1.655 $X2=0.385
+ $Y2=1.475
cc_253 VPB Q 0.00480048f $X=-0.19 $Y=1.655 $X2=0.48 $Y2=2.6
cc_254 VPB Q_N 0.0154561f $X=-0.19 $Y=1.655 $X2=0.387 $Y2=1.98
cc_255 VPB N_Q_N_c_1693_n 0.00455019f $X=-0.19 $Y=1.655 $X2=0.277 $Y2=1.295
cc_256 VPB N_Q_N_c_1696_n 0.0541945f $X=-0.19 $Y=1.655 $X2=0.24 $Y2=2.035
cc_257 CLK N_A_111_156#_c_299_n 0.0058512f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_258 N_CLK_c_262_n N_A_111_156#_c_299_n 0.00505414f $X=0.387 $Y=1.31 $X2=0
+ $Y2=0
cc_259 CLK N_A_111_156#_c_300_n 0.0486934f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_260 CLK N_A_111_156#_c_300_n 0.0110102f $X=0.155 $Y=1.95 $X2=0 $Y2=0
cc_261 N_CLK_c_261_n N_A_111_156#_c_300_n 0.00893244f $X=0.385 $Y=1.475 $X2=0
+ $Y2=0
cc_262 N_CLK_M1021_g N_A_111_156#_c_333_n 0.00149065f $X=0.48 $Y=2.6 $X2=0 $Y2=0
cc_263 CLK N_A_111_156#_c_333_n 0.00962282f $X=0.155 $Y=1.95 $X2=0 $Y2=0
cc_264 N_CLK_M1021_g N_A_111_156#_c_334_n 0.00485563f $X=0.48 $Y=2.6 $X2=0 $Y2=0
cc_265 CLK N_A_111_156#_c_316_n 0.0144494f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_266 N_CLK_c_262_n N_A_111_156#_c_316_n 0.00175122f $X=0.387 $Y=1.31 $X2=0
+ $Y2=0
cc_267 CLK N_A_161_21#_c_1018_n 2.76313e-19 $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_268 N_CLK_c_262_n N_A_161_21#_c_1018_n 0.0136619f $X=0.387 $Y=1.31 $X2=0
+ $Y2=0
cc_269 N_CLK_c_259_n N_A_161_21#_c_1035_n 0.0136619f $X=0.387 $Y=1.813 $X2=0
+ $Y2=0
cc_270 CLK N_VPWR_M1021_s 0.00325852f $X=0.155 $Y=1.95 $X2=-0.19 $Y2=-0.245
cc_271 N_CLK_M1021_g N_VPWR_c_1481_n 0.00845652f $X=0.48 $Y=2.6 $X2=0 $Y2=0
cc_272 N_CLK_c_265_n N_VPWR_c_1481_n 4.66209e-19 $X=0.387 $Y=1.98 $X2=0 $Y2=0
cc_273 CLK N_VPWR_c_1481_n 0.0238082f $X=0.155 $Y=1.95 $X2=0 $Y2=0
cc_274 N_CLK_M1021_g N_VPWR_c_1490_n 0.00455951f $X=0.48 $Y=2.6 $X2=0 $Y2=0
cc_275 N_CLK_M1021_g N_VPWR_c_1479_n 0.00447788f $X=0.48 $Y=2.6 $X2=0 $Y2=0
cc_276 CLK N_VPWR_c_1479_n 0.00177675f $X=0.155 $Y=1.95 $X2=0 $Y2=0
cc_277 CLK N_VGND_c_1712_n 0.0274352f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_278 N_CLK_c_261_n N_VGND_c_1712_n 9.83752e-19 $X=0.385 $Y=1.475 $X2=0 $Y2=0
cc_279 N_CLK_c_262_n N_VGND_c_1712_n 0.00961427f $X=0.387 $Y=1.31 $X2=0 $Y2=0
cc_280 N_CLK_c_262_n N_VGND_c_1725_n 0.00284536f $X=0.387 $Y=1.31 $X2=0 $Y2=0
cc_281 N_CLK_c_262_n N_VGND_c_1729_n 0.00360052f $X=0.387 $Y=1.31 $X2=0 $Y2=0
cc_282 N_A_111_156#_c_293_n N_D_M1008_g 0.00477349f $X=1.585 $Y=1.125 $X2=0
+ $Y2=0
cc_283 N_A_111_156#_M1010_g N_D_M1008_g 0.015991f $X=2.825 $Y=0.805 $X2=0 $Y2=0
cc_284 N_A_111_156#_c_301_n N_D_M1008_g 0.00250774f $X=2.145 $Y=1.1 $X2=0 $Y2=0
cc_285 N_A_111_156#_c_302_n N_D_M1008_g 0.00764588f $X=2.23 $Y=1.015 $X2=0 $Y2=0
cc_286 N_A_111_156#_c_303_n N_D_M1008_g 0.00758946f $X=3.325 $Y=0.385 $X2=0
+ $Y2=0
cc_287 N_A_111_156#_c_317_n N_D_M1008_g 4.60587e-19 $X=1.732 $Y=1.1 $X2=0 $Y2=0
cc_288 N_A_111_156#_c_319_n N_D_M1008_g 0.00406518f $X=1.72 $Y=1.29 $X2=0 $Y2=0
cc_289 N_A_111_156#_c_323_n N_D_M1018_g 0.0123739f $X=1.815 $Y=3.075 $X2=0 $Y2=0
cc_290 N_A_111_156#_M1010_g N_D_c_559_n 2.31615e-19 $X=2.825 $Y=0.805 $X2=0
+ $Y2=0
cc_291 N_A_111_156#_c_301_n N_D_c_559_n 0.0270516f $X=2.145 $Y=1.1 $X2=0 $Y2=0
cc_292 N_A_111_156#_c_317_n N_D_c_559_n 0.00778464f $X=1.732 $Y=1.1 $X2=0 $Y2=0
cc_293 N_A_111_156#_c_319_n N_D_c_559_n 6.5673e-19 $X=1.72 $Y=1.29 $X2=0 $Y2=0
cc_294 N_A_111_156#_c_296_n N_D_c_560_n 0.015991f $X=2.9 $Y=1.53 $X2=0 $Y2=0
cc_295 N_A_111_156#_c_301_n N_D_c_560_n 0.00559069f $X=2.145 $Y=1.1 $X2=0 $Y2=0
cc_296 N_A_111_156#_c_317_n N_D_c_560_n 6.05682e-19 $X=1.732 $Y=1.1 $X2=0 $Y2=0
cc_297 N_A_111_156#_c_319_n N_D_c_560_n 0.011833f $X=1.72 $Y=1.29 $X2=0 $Y2=0
cc_298 N_A_111_156#_c_323_n N_D_c_563_n 0.00727076f $X=1.815 $Y=3.075 $X2=0
+ $Y2=0
cc_299 N_A_111_156#_c_323_n N_D_c_564_n 0.00297115f $X=1.815 $Y=3.075 $X2=0
+ $Y2=0
cc_300 N_A_111_156#_c_305_n N_A_708_93#_c_615_n 0.00294884f $X=3.41 $Y=1.075
+ $X2=0 $Y2=0
cc_301 N_A_111_156#_c_308_n N_A_708_93#_c_615_n 0.00489135f $X=4.095 $Y=1.16
+ $X2=0 $Y2=0
cc_302 N_A_111_156#_c_309_n N_A_708_93#_c_615_n 0.00275679f $X=4.18 $Y=1.075
+ $X2=0 $Y2=0
cc_303 N_A_111_156#_c_320_n N_A_708_93#_c_615_n 0.00466565f $X=3.325 $Y=1.075
+ $X2=0 $Y2=0
cc_304 N_A_111_156#_c_308_n N_A_708_93#_c_616_n 0.0253012f $X=4.095 $Y=1.16
+ $X2=0 $Y2=0
cc_305 N_A_111_156#_M1010_g N_A_708_93#_c_617_n 0.00150216f $X=2.825 $Y=0.805
+ $X2=0 $Y2=0
cc_306 N_A_111_156#_c_295_n N_A_708_93#_c_617_n 0.00835095f $X=3.215 $Y=1.53
+ $X2=0 $Y2=0
cc_307 N_A_111_156#_c_306_n N_A_708_93#_c_617_n 0.00316595f $X=3.495 $Y=1.66
+ $X2=0 $Y2=0
cc_308 N_A_111_156#_c_308_n N_A_708_93#_c_617_n 0.00242507f $X=4.095 $Y=1.16
+ $X2=0 $Y2=0
cc_309 N_A_111_156#_c_320_n N_A_708_93#_c_617_n 0.00233189f $X=3.325 $Y=1.075
+ $X2=0 $Y2=0
cc_310 N_A_111_156#_M1028_g N_A_708_93#_c_624_n 0.0504846f $X=3.36 $Y=2.875
+ $X2=0 $Y2=0
cc_311 N_A_111_156#_c_326_n N_A_708_93#_c_624_n 0.00100247f $X=3.437 $Y=2.165
+ $X2=0 $Y2=0
cc_312 N_A_111_156#_c_295_n N_A_708_93#_c_618_n 3.88491e-19 $X=3.215 $Y=1.53
+ $X2=0 $Y2=0
cc_313 N_A_111_156#_c_306_n N_A_708_93#_c_618_n 0.00887771f $X=3.495 $Y=1.66
+ $X2=0 $Y2=0
cc_314 N_A_111_156#_c_308_n N_A_708_93#_c_618_n 0.026356f $X=4.095 $Y=1.16 $X2=0
+ $Y2=0
cc_315 N_A_111_156#_c_310_n N_A_708_93#_c_618_n 0.00534994f $X=4.815 $Y=0.69
+ $X2=0 $Y2=0
cc_316 N_A_111_156#_c_295_n N_A_708_93#_c_619_n 0.00563733f $X=3.215 $Y=1.53
+ $X2=0 $Y2=0
cc_317 N_A_111_156#_c_306_n N_A_708_93#_c_619_n 0.004967f $X=3.495 $Y=1.66 $X2=0
+ $Y2=0
cc_318 N_A_111_156#_c_308_n N_A_708_93#_c_620_n 0.0136568f $X=4.095 $Y=1.16
+ $X2=0 $Y2=0
cc_319 N_A_111_156#_c_309_n N_A_708_93#_c_620_n 0.0085502f $X=4.18 $Y=1.075
+ $X2=0 $Y2=0
cc_320 N_A_111_156#_c_310_n N_A_708_93#_c_620_n 0.0139262f $X=4.815 $Y=0.69
+ $X2=0 $Y2=0
cc_321 N_A_111_156#_c_314_n N_A_708_93#_c_620_n 0.0122989f $X=4.985 $Y=1.33
+ $X2=0 $Y2=0
cc_322 N_A_111_156#_c_306_n N_A_708_93#_c_621_n 5.10435e-19 $X=3.495 $Y=1.66
+ $X2=0 $Y2=0
cc_323 N_A_111_156#_c_307_n N_A_708_93#_c_621_n 0.00497831f $X=3.495 $Y=1.66
+ $X2=0 $Y2=0
cc_324 N_A_111_156#_M1028_g N_A_708_93#_c_629_n 0.00278895f $X=3.36 $Y=2.875
+ $X2=0 $Y2=0
cc_325 N_A_111_156#_c_306_n N_A_708_93#_c_629_n 7.35108e-19 $X=3.495 $Y=1.66
+ $X2=0 $Y2=0
cc_326 N_A_111_156#_c_307_n N_A_708_93#_c_629_n 0.0133114f $X=3.495 $Y=1.66
+ $X2=0 $Y2=0
cc_327 N_A_111_156#_c_309_n N_A_580_119#_M1012_g 0.00287335f $X=4.18 $Y=1.075
+ $X2=0 $Y2=0
cc_328 N_A_111_156#_c_310_n N_A_580_119#_M1012_g 0.0103927f $X=4.815 $Y=0.69
+ $X2=0 $Y2=0
cc_329 N_A_111_156#_c_312_n N_A_580_119#_M1012_g 0.00887655f $X=4.9 $Y=1.245
+ $X2=0 $Y2=0
cc_330 N_A_111_156#_c_314_n N_A_580_119#_M1012_g 0.00318488f $X=4.985 $Y=1.33
+ $X2=0 $Y2=0
cc_331 N_A_111_156#_c_313_n N_A_580_119#_M1026_g 0.0175645f $X=6.27 $Y=1.33
+ $X2=0 $Y2=0
cc_332 N_A_111_156#_c_315_n N_A_580_119#_M1026_g 0.00154431f $X=6.635 $Y=1.505
+ $X2=0 $Y2=0
cc_333 N_A_111_156#_c_313_n N_A_580_119#_c_720_n 0.0159161f $X=6.27 $Y=1.33
+ $X2=0 $Y2=0
cc_334 N_A_111_156#_c_315_n N_A_580_119#_c_720_n 0.00578335f $X=6.635 $Y=1.505
+ $X2=0 $Y2=0
cc_335 N_A_111_156#_c_321_n N_A_580_119#_c_720_n 0.011351f $X=6.67 $Y=1.5 $X2=0
+ $Y2=0
cc_336 N_A_111_156#_M1010_g N_A_580_119#_c_722_n 0.00637176f $X=2.825 $Y=0.805
+ $X2=0 $Y2=0
cc_337 N_A_111_156#_c_303_n N_A_580_119#_c_722_n 0.0142211f $X=3.325 $Y=0.385
+ $X2=0 $Y2=0
cc_338 N_A_111_156#_c_305_n N_A_580_119#_c_722_n 0.0168311f $X=3.41 $Y=1.075
+ $X2=0 $Y2=0
cc_339 N_A_111_156#_c_306_n N_A_580_119#_c_722_n 0.0102035f $X=3.495 $Y=1.66
+ $X2=0 $Y2=0
cc_340 N_A_111_156#_c_320_n N_A_580_119#_c_722_n 0.014055f $X=3.325 $Y=1.075
+ $X2=0 $Y2=0
cc_341 N_A_111_156#_c_295_n N_A_580_119#_c_723_n 0.00456652f $X=3.215 $Y=1.53
+ $X2=0 $Y2=0
cc_342 N_A_111_156#_M1028_g N_A_580_119#_c_723_n 0.00378512f $X=3.36 $Y=2.875
+ $X2=0 $Y2=0
cc_343 N_A_111_156#_c_326_n N_A_580_119#_c_723_n 0.00496052f $X=3.437 $Y=2.165
+ $X2=0 $Y2=0
cc_344 N_A_111_156#_c_307_n N_A_580_119#_c_723_n 0.00937621f $X=3.495 $Y=1.66
+ $X2=0 $Y2=0
cc_345 N_A_111_156#_M1028_g N_A_580_119#_c_767_n 0.0069512f $X=3.36 $Y=2.875
+ $X2=0 $Y2=0
cc_346 N_A_111_156#_M1028_g N_A_580_119#_c_736_n 0.0110691f $X=3.36 $Y=2.875
+ $X2=0 $Y2=0
cc_347 N_A_111_156#_c_326_n N_A_580_119#_c_736_n 0.00227442f $X=3.437 $Y=2.165
+ $X2=0 $Y2=0
cc_348 N_A_111_156#_c_306_n N_A_580_119#_c_736_n 0.0104471f $X=3.495 $Y=1.66
+ $X2=0 $Y2=0
cc_349 N_A_111_156#_M1028_g N_A_580_119#_c_737_n 0.0024229f $X=3.36 $Y=2.875
+ $X2=0 $Y2=0
cc_350 N_A_111_156#_c_306_n N_A_580_119#_c_737_n 0.0166635f $X=3.495 $Y=1.66
+ $X2=0 $Y2=0
cc_351 N_A_111_156#_c_307_n N_A_580_119#_c_737_n 0.00199468f $X=3.495 $Y=1.66
+ $X2=0 $Y2=0
cc_352 N_A_111_156#_c_306_n N_A_580_119#_c_739_n 0.0139282f $X=3.495 $Y=1.66
+ $X2=0 $Y2=0
cc_353 N_A_111_156#_c_307_n N_A_580_119#_c_739_n 0.00164173f $X=3.495 $Y=1.66
+ $X2=0 $Y2=0
cc_354 N_A_111_156#_c_308_n N_A_580_119#_c_739_n 0.0040153f $X=4.095 $Y=1.16
+ $X2=0 $Y2=0
cc_355 N_A_111_156#_c_314_n N_A_580_119#_c_724_n 0.015246f $X=4.985 $Y=1.33
+ $X2=0 $Y2=0
cc_356 N_A_111_156#_c_314_n N_A_580_119#_c_742_n 4.82014e-19 $X=4.985 $Y=1.33
+ $X2=0 $Y2=0
cc_357 N_A_111_156#_c_298_n N_A_580_119#_c_743_n 9.81271e-19 $X=6.67 $Y=1.84
+ $X2=0 $Y2=0
cc_358 N_A_111_156#_c_313_n N_A_580_119#_c_743_n 0.0201453f $X=6.27 $Y=1.33
+ $X2=0 $Y2=0
cc_359 N_A_111_156#_c_315_n N_A_580_119#_c_743_n 0.016024f $X=6.635 $Y=1.505
+ $X2=0 $Y2=0
cc_360 N_A_111_156#_c_298_n N_A_580_119#_c_725_n 0.011351f $X=6.67 $Y=1.84 $X2=0
+ $Y2=0
cc_361 N_A_111_156#_c_295_n N_A_580_119#_c_726_n 0.0156111f $X=3.215 $Y=1.53
+ $X2=0 $Y2=0
cc_362 N_A_111_156#_c_306_n N_A_580_119#_c_726_n 0.0525446f $X=3.495 $Y=1.66
+ $X2=0 $Y2=0
cc_363 N_A_111_156#_M1028_g N_A_580_119#_c_745_n 0.00316256f $X=3.36 $Y=2.875
+ $X2=0 $Y2=0
cc_364 N_A_111_156#_c_326_n N_A_580_119#_c_745_n 0.0022031f $X=3.437 $Y=2.165
+ $X2=0 $Y2=0
cc_365 N_A_111_156#_c_313_n N_A_580_119#_c_727_n 0.0608509f $X=6.27 $Y=1.33
+ $X2=0 $Y2=0
cc_366 N_A_111_156#_c_315_n N_A_580_119#_c_728_n 0.00248961f $X=6.635 $Y=1.505
+ $X2=0 $Y2=0
cc_367 N_A_111_156#_M1007_g N_A_580_119#_c_748_n 0.0325237f $X=6.76 $Y=2.665
+ $X2=0 $Y2=0
cc_368 N_A_111_156#_c_328_n N_A_580_119#_c_748_n 0.011351f $X=6.67 $Y=2.005
+ $X2=0 $Y2=0
cc_369 N_A_111_156#_c_310_n N_SET_B_M1009_g 5.52862e-19 $X=4.815 $Y=0.69 $X2=0
+ $Y2=0
cc_370 N_A_111_156#_c_312_n N_SET_B_M1009_g 0.00184865f $X=4.9 $Y=1.245 $X2=0
+ $Y2=0
cc_371 N_A_111_156#_c_313_n N_SET_B_M1009_g 0.0141906f $X=6.27 $Y=1.33 $X2=0
+ $Y2=0
cc_372 N_A_111_156#_c_313_n N_SET_B_c_894_n 0.00421866f $X=6.27 $Y=1.33 $X2=0
+ $Y2=0
cc_373 N_A_111_156#_M1007_g N_SET_B_c_911_n 0.00509745f $X=6.76 $Y=2.665 $X2=0
+ $Y2=0
cc_374 N_A_111_156#_M1007_g N_SET_B_c_899_n 0.019159f $X=6.76 $Y=2.665 $X2=0
+ $Y2=0
cc_375 N_A_111_156#_M1007_g N_SET_B_c_900_n 0.00116931f $X=6.76 $Y=2.665 $X2=0
+ $Y2=0
cc_376 N_A_111_156#_M1007_g N_SET_B_c_905_n 0.00238413f $X=6.76 $Y=2.665 $X2=0
+ $Y2=0
cc_377 N_A_111_156#_c_299_n N_A_161_21#_c_1018_n 0.0102702f $X=0.735 $Y=0.995
+ $X2=0 $Y2=0
cc_378 N_A_111_156#_c_300_n N_A_161_21#_c_1018_n 0.0120089f $X=0.74 $Y=2.26
+ $X2=0 $Y2=0
cc_379 N_A_111_156#_c_317_n N_A_161_21#_c_1018_n 0.00134951f $X=1.732 $Y=1.1
+ $X2=0 $Y2=0
cc_380 N_A_111_156#_c_318_n N_A_161_21#_c_1018_n 0.0177561f $X=1.72 $Y=1.29
+ $X2=0 $Y2=0
cc_381 N_A_111_156#_c_319_n N_A_161_21#_c_1018_n 0.0112983f $X=1.72 $Y=1.29
+ $X2=0 $Y2=0
cc_382 N_A_111_156#_c_293_n N_A_161_21#_c_1019_n 0.0103562f $X=1.585 $Y=1.125
+ $X2=0 $Y2=0
cc_383 N_A_111_156#_M1010_g N_A_161_21#_c_1019_n 0.00880114f $X=2.825 $Y=0.805
+ $X2=0 $Y2=0
cc_384 N_A_111_156#_c_303_n N_A_161_21#_c_1019_n 0.0129137f $X=3.325 $Y=0.385
+ $X2=0 $Y2=0
cc_385 N_A_111_156#_c_304_n N_A_161_21#_c_1019_n 0.00412631f $X=2.315 $Y=0.385
+ $X2=0 $Y2=0
cc_386 N_A_111_156#_c_323_n N_A_161_21#_c_1030_n 0.0100632f $X=1.815 $Y=3.075
+ $X2=0 $Y2=0
cc_387 N_A_111_156#_c_296_n N_A_161_21#_c_1030_n 0.0174145f $X=2.9 $Y=1.53 $X2=0
+ $Y2=0
cc_388 N_A_111_156#_c_301_n N_A_161_21#_c_1030_n 0.00294862f $X=2.145 $Y=1.1
+ $X2=0 $Y2=0
cc_389 N_A_111_156#_c_307_n N_A_161_21#_c_1030_n 0.0107376f $X=3.495 $Y=1.66
+ $X2=0 $Y2=0
cc_390 N_A_111_156#_c_317_n N_A_161_21#_c_1030_n 5.41831e-19 $X=1.732 $Y=1.1
+ $X2=0 $Y2=0
cc_391 N_A_111_156#_c_318_n N_A_161_21#_c_1030_n 3.12266e-19 $X=1.72 $Y=1.29
+ $X2=0 $Y2=0
cc_392 N_A_111_156#_c_319_n N_A_161_21#_c_1030_n 0.0125601f $X=1.72 $Y=1.29
+ $X2=0 $Y2=0
cc_393 N_A_111_156#_M1028_g N_A_161_21#_M1003_g 0.0261571f $X=3.36 $Y=2.875
+ $X2=0 $Y2=0
cc_394 N_A_111_156#_c_326_n N_A_161_21#_M1003_g 0.0107376f $X=3.437 $Y=2.165
+ $X2=0 $Y2=0
cc_395 N_A_111_156#_M1010_g N_A_161_21#_M1000_g 0.011754f $X=2.825 $Y=0.805
+ $X2=0 $Y2=0
cc_396 N_A_111_156#_c_295_n N_A_161_21#_M1000_g 0.00780919f $X=3.215 $Y=1.53
+ $X2=0 $Y2=0
cc_397 N_A_111_156#_c_303_n N_A_161_21#_M1000_g 0.0170187f $X=3.325 $Y=0.385
+ $X2=0 $Y2=0
cc_398 N_A_111_156#_c_305_n N_A_161_21#_M1000_g 0.0101175f $X=3.41 $Y=1.075
+ $X2=0 $Y2=0
cc_399 N_A_111_156#_c_320_n N_A_161_21#_M1000_g 0.00128001f $X=3.325 $Y=1.075
+ $X2=0 $Y2=0
cc_400 N_A_111_156#_M1019_g N_A_161_21#_c_1021_n 0.00409527f $X=6.58 $Y=0.965
+ $X2=0 $Y2=0
cc_401 N_A_111_156#_c_303_n N_A_161_21#_c_1021_n 0.00182043f $X=3.325 $Y=0.385
+ $X2=0 $Y2=0
cc_402 N_A_111_156#_c_310_n N_A_161_21#_c_1021_n 0.0118222f $X=4.815 $Y=0.69
+ $X2=0 $Y2=0
cc_403 N_A_111_156#_c_311_n N_A_161_21#_c_1021_n 0.00334788f $X=4.265 $Y=0.69
+ $X2=0 $Y2=0
cc_404 N_A_111_156#_M1019_g N_A_161_21#_M1020_g 0.0150342f $X=6.58 $Y=0.965
+ $X2=0 $Y2=0
cc_405 N_A_111_156#_c_321_n N_A_161_21#_M1033_g 0.0289994f $X=6.67 $Y=1.5 $X2=0
+ $Y2=0
cc_406 N_A_111_156#_c_321_n N_A_161_21#_c_1025_n 0.00600905f $X=6.67 $Y=1.5
+ $X2=0 $Y2=0
cc_407 N_A_111_156#_c_293_n N_A_161_21#_c_1026_n 4.80654e-19 $X=1.585 $Y=1.125
+ $X2=0 $Y2=0
cc_408 N_A_111_156#_c_299_n N_A_161_21#_c_1026_n 0.00425091f $X=0.735 $Y=0.995
+ $X2=0 $Y2=0
cc_409 N_A_111_156#_c_300_n N_A_161_21#_c_1033_n 0.0211354f $X=0.74 $Y=2.26
+ $X2=0 $Y2=0
cc_410 N_A_111_156#_c_333_n N_A_161_21#_c_1033_n 0.02457f $X=0.695 $Y=2.425
+ $X2=0 $Y2=0
cc_411 N_A_111_156#_c_317_n N_A_161_21#_c_1033_n 0.00575883f $X=1.732 $Y=1.1
+ $X2=0 $Y2=0
cc_412 N_A_111_156#_c_318_n N_A_161_21#_c_1033_n 0.0255594f $X=1.72 $Y=1.29
+ $X2=0 $Y2=0
cc_413 N_A_111_156#_c_319_n N_A_161_21#_c_1033_n 7.71804e-19 $X=1.72 $Y=1.29
+ $X2=0 $Y2=0
cc_414 N_A_111_156#_c_293_n N_A_161_21#_c_1027_n 6.9934e-19 $X=1.585 $Y=1.125
+ $X2=0 $Y2=0
cc_415 N_A_111_156#_c_299_n N_A_161_21#_c_1027_n 0.00614305f $X=0.735 $Y=0.995
+ $X2=0 $Y2=0
cc_416 N_A_111_156#_c_318_n N_A_161_21#_c_1027_n 0.0127466f $X=1.72 $Y=1.29
+ $X2=0 $Y2=0
cc_417 N_A_111_156#_c_322_n N_A_161_21#_c_1034_n 0.00386976f $X=1.74 $Y=3.15
+ $X2=0 $Y2=0
cc_418 N_A_111_156#_c_323_n N_A_161_21#_c_1034_n 0.0141521f $X=1.815 $Y=3.075
+ $X2=0 $Y2=0
cc_419 N_A_111_156#_c_300_n N_A_161_21#_c_1034_n 0.00525431f $X=0.74 $Y=2.26
+ $X2=0 $Y2=0
cc_420 N_A_111_156#_c_333_n N_A_161_21#_c_1034_n 0.0607137f $X=0.695 $Y=2.425
+ $X2=0 $Y2=0
cc_421 N_A_111_156#_c_334_n N_A_161_21#_c_1034_n 7.66122e-19 $X=1.15 $Y=2.94
+ $X2=0 $Y2=0
cc_422 N_A_111_156#_c_293_n N_A_161_21#_c_1028_n 0.0112983f $X=1.585 $Y=1.125
+ $X2=0 $Y2=0
cc_423 N_A_111_156#_c_299_n N_A_161_21#_c_1028_n 0.00208703f $X=0.735 $Y=0.995
+ $X2=0 $Y2=0
cc_424 N_A_111_156#_c_333_n N_A_161_21#_c_1035_n 0.0050534f $X=0.695 $Y=2.425
+ $X2=0 $Y2=0
cc_425 N_A_111_156#_c_334_n N_A_161_21#_c_1035_n 0.0039883f $X=1.15 $Y=2.94
+ $X2=0 $Y2=0
cc_426 N_A_111_156#_c_318_n N_A_161_21#_c_1035_n 0.00646261f $X=1.72 $Y=1.29
+ $X2=0 $Y2=0
cc_427 N_A_111_156#_M1019_g N_A_1331_151#_c_1243_n 0.00205058f $X=6.58 $Y=0.965
+ $X2=0 $Y2=0
cc_428 N_A_111_156#_c_315_n N_A_1331_151#_c_1243_n 0.00288606f $X=6.635 $Y=1.505
+ $X2=0 $Y2=0
cc_429 N_A_111_156#_c_315_n N_A_1331_151#_c_1273_n 0.0047274f $X=6.635 $Y=1.505
+ $X2=0 $Y2=0
cc_430 N_A_111_156#_c_321_n N_A_1331_151#_c_1273_n 0.00339772f $X=6.67 $Y=1.5
+ $X2=0 $Y2=0
cc_431 N_A_111_156#_M1007_g N_A_1331_151#_c_1266_n 0.00713829f $X=6.76 $Y=2.665
+ $X2=0 $Y2=0
cc_432 N_A_111_156#_c_315_n N_A_1331_151#_c_1250_n 0.0388738f $X=6.635 $Y=1.505
+ $X2=0 $Y2=0
cc_433 N_A_111_156#_c_321_n N_A_1331_151#_c_1250_n 0.0107416f $X=6.67 $Y=1.5
+ $X2=0 $Y2=0
cc_434 N_A_111_156#_c_315_n N_A_1331_151#_c_1251_n 0.0141401f $X=6.635 $Y=1.505
+ $X2=0 $Y2=0
cc_435 N_A_111_156#_c_321_n N_A_1331_151#_c_1251_n 0.00118378f $X=6.67 $Y=1.5
+ $X2=0 $Y2=0
cc_436 N_A_111_156#_c_333_n N_VPWR_c_1481_n 0.0155886f $X=0.695 $Y=2.425 $X2=0
+ $Y2=0
cc_437 N_A_111_156#_c_334_n N_VPWR_c_1481_n 0.00286963f $X=1.15 $Y=2.94 $X2=0
+ $Y2=0
cc_438 N_A_111_156#_c_323_n N_VPWR_c_1482_n 0.00955628f $X=1.815 $Y=3.075 $X2=0
+ $Y2=0
cc_439 N_A_111_156#_M1028_g N_VPWR_c_1483_n 0.00188523f $X=3.36 $Y=2.875 $X2=0
+ $Y2=0
cc_440 N_A_111_156#_M1007_g N_VPWR_c_1484_n 0.00107108f $X=6.76 $Y=2.665 $X2=0
+ $Y2=0
cc_441 N_A_111_156#_c_333_n N_VPWR_c_1490_n 0.0374786f $X=0.695 $Y=2.425 $X2=0
+ $Y2=0
cc_442 N_A_111_156#_c_334_n N_VPWR_c_1490_n 0.0251103f $X=1.15 $Y=2.94 $X2=0
+ $Y2=0
cc_443 N_A_111_156#_M1028_g N_VPWR_c_1491_n 0.0041283f $X=3.36 $Y=2.875 $X2=0
+ $Y2=0
cc_444 N_A_111_156#_M1007_g N_VPWR_c_1493_n 0.00351226f $X=6.76 $Y=2.665 $X2=0
+ $Y2=0
cc_445 N_A_111_156#_c_322_n N_VPWR_c_1479_n 0.0259298f $X=1.74 $Y=3.15 $X2=0
+ $Y2=0
cc_446 N_A_111_156#_M1028_g N_VPWR_c_1479_n 0.00575681f $X=3.36 $Y=2.875 $X2=0
+ $Y2=0
cc_447 N_A_111_156#_M1007_g N_VPWR_c_1479_n 0.00687926f $X=6.76 $Y=2.665 $X2=0
+ $Y2=0
cc_448 N_A_111_156#_c_333_n N_VPWR_c_1479_n 0.0251605f $X=0.695 $Y=2.425 $X2=0
+ $Y2=0
cc_449 N_A_111_156#_c_334_n N_VPWR_c_1479_n 0.0101216f $X=1.15 $Y=2.94 $X2=0
+ $Y2=0
cc_450 N_A_111_156#_M1010_g N_A_494_119#_c_1626_n 0.00830006f $X=2.825 $Y=0.805
+ $X2=0 $Y2=0
cc_451 N_A_111_156#_c_296_n N_A_494_119#_c_1626_n 0.00371273f $X=2.9 $Y=1.53
+ $X2=0 $Y2=0
cc_452 N_A_111_156#_c_301_n N_A_494_119#_c_1626_n 0.00957223f $X=2.145 $Y=1.1
+ $X2=0 $Y2=0
cc_453 N_A_111_156#_c_307_n N_A_494_119#_c_1626_n 7.42124e-19 $X=3.495 $Y=1.66
+ $X2=0 $Y2=0
cc_454 N_A_111_156#_M1010_g N_A_494_119#_c_1634_n 0.00364626f $X=2.825 $Y=0.805
+ $X2=0 $Y2=0
cc_455 N_A_111_156#_c_303_n N_A_494_119#_c_1634_n 0.0176282f $X=3.325 $Y=0.385
+ $X2=0 $Y2=0
cc_456 N_A_111_156#_c_296_n N_A_494_119#_c_1629_n 0.00248716f $X=2.9 $Y=1.53
+ $X2=0 $Y2=0
cc_457 N_A_111_156#_c_307_n N_A_494_119#_c_1629_n 3.39066e-19 $X=3.495 $Y=1.66
+ $X2=0 $Y2=0
cc_458 N_A_111_156#_c_302_n N_VGND_M1011_d 0.00728913f $X=2.23 $Y=1.015 $X2=0
+ $Y2=0
cc_459 N_A_111_156#_c_317_n N_VGND_M1011_d 0.00184553f $X=1.732 $Y=1.1 $X2=0
+ $Y2=0
cc_460 N_A_111_156#_c_313_n N_VGND_M1009_d 0.00317561f $X=6.27 $Y=1.33 $X2=0
+ $Y2=0
cc_461 N_A_111_156#_c_299_n N_VGND_c_1712_n 0.0136042f $X=0.735 $Y=0.995 $X2=0
+ $Y2=0
cc_462 N_A_111_156#_c_293_n N_VGND_c_1713_n 0.00620105f $X=1.585 $Y=1.125 $X2=0
+ $Y2=0
cc_463 N_A_111_156#_c_301_n N_VGND_c_1713_n 0.0119073f $X=2.145 $Y=1.1 $X2=0
+ $Y2=0
cc_464 N_A_111_156#_c_302_n N_VGND_c_1713_n 0.0289778f $X=2.23 $Y=1.015 $X2=0
+ $Y2=0
cc_465 N_A_111_156#_c_304_n N_VGND_c_1713_n 0.0150385f $X=2.315 $Y=0.385 $X2=0
+ $Y2=0
cc_466 N_A_111_156#_c_317_n N_VGND_c_1713_n 0.0132961f $X=1.732 $Y=1.1 $X2=0
+ $Y2=0
cc_467 N_A_111_156#_c_319_n N_VGND_c_1713_n 0.00120849f $X=1.72 $Y=1.29 $X2=0
+ $Y2=0
cc_468 N_A_111_156#_c_303_n N_VGND_c_1714_n 0.0117407f $X=3.325 $Y=0.385 $X2=0
+ $Y2=0
cc_469 N_A_111_156#_c_305_n N_VGND_c_1714_n 0.00761308f $X=3.41 $Y=1.075 $X2=0
+ $Y2=0
cc_470 N_A_111_156#_c_308_n N_VGND_c_1714_n 0.0154298f $X=4.095 $Y=1.16 $X2=0
+ $Y2=0
cc_471 N_A_111_156#_c_309_n N_VGND_c_1714_n 0.0096943f $X=4.18 $Y=1.075 $X2=0
+ $Y2=0
cc_472 N_A_111_156#_c_311_n N_VGND_c_1714_n 0.0142846f $X=4.265 $Y=0.69 $X2=0
+ $Y2=0
cc_473 N_A_111_156#_c_310_n N_VGND_c_1715_n 0.0108629f $X=4.815 $Y=0.69 $X2=0
+ $Y2=0
cc_474 N_A_111_156#_c_312_n N_VGND_c_1715_n 0.0104018f $X=4.9 $Y=1.245 $X2=0
+ $Y2=0
cc_475 N_A_111_156#_c_313_n N_VGND_c_1715_n 0.0200956f $X=6.27 $Y=1.33 $X2=0
+ $Y2=0
cc_476 N_A_111_156#_c_303_n N_VGND_c_1719_n 0.0597772f $X=3.325 $Y=0.385 $X2=0
+ $Y2=0
cc_477 N_A_111_156#_c_304_n N_VGND_c_1719_n 0.00947234f $X=2.315 $Y=0.385 $X2=0
+ $Y2=0
cc_478 N_A_111_156#_c_310_n N_VGND_c_1721_n 0.014331f $X=4.815 $Y=0.69 $X2=0
+ $Y2=0
cc_479 N_A_111_156#_c_311_n N_VGND_c_1721_n 0.00364552f $X=4.265 $Y=0.69 $X2=0
+ $Y2=0
cc_480 N_A_111_156#_c_293_n N_VGND_c_1729_n 8.51577e-19 $X=1.585 $Y=1.125 $X2=0
+ $Y2=0
cc_481 N_A_111_156#_c_299_n N_VGND_c_1729_n 0.00683311f $X=0.735 $Y=0.995 $X2=0
+ $Y2=0
cc_482 N_A_111_156#_c_303_n N_VGND_c_1729_n 0.038504f $X=3.325 $Y=0.385 $X2=0
+ $Y2=0
cc_483 N_A_111_156#_c_304_n N_VGND_c_1729_n 0.00578067f $X=2.315 $Y=0.385 $X2=0
+ $Y2=0
cc_484 N_A_111_156#_c_310_n N_VGND_c_1729_n 0.0185041f $X=4.815 $Y=0.69 $X2=0
+ $Y2=0
cc_485 N_A_111_156#_c_311_n N_VGND_c_1729_n 0.00458776f $X=4.265 $Y=0.69 $X2=0
+ $Y2=0
cc_486 N_A_111_156#_c_313_n N_A_1141_125#_M1026_d 0.00230047f $X=6.27 $Y=1.33
+ $X2=-0.19 $Y2=-0.245
cc_487 N_A_111_156#_M1019_g N_A_1141_125#_c_1841_n 9.96624e-19 $X=6.58 $Y=0.965
+ $X2=0 $Y2=0
cc_488 N_A_111_156#_c_313_n N_A_1141_125#_c_1841_n 0.0202164f $X=6.27 $Y=1.33
+ $X2=0 $Y2=0
cc_489 N_A_111_156#_M1019_g N_A_1141_125#_c_1843_n 4.96616e-19 $X=6.58 $Y=0.965
+ $X2=0 $Y2=0
cc_490 N_A_111_156#_M1019_g N_A_1248_151#_c_1865_n 0.00867354f $X=6.58 $Y=0.965
+ $X2=0 $Y2=0
cc_491 N_A_111_156#_c_315_n N_A_1248_151#_c_1865_n 0.00433468f $X=6.635 $Y=1.505
+ $X2=0 $Y2=0
cc_492 N_A_111_156#_M1019_g N_A_1248_151#_c_1866_n 0.00877782f $X=6.58 $Y=0.965
+ $X2=0 $Y2=0
cc_493 N_A_111_156#_c_313_n N_A_1248_151#_c_1866_n 0.00555706f $X=6.27 $Y=1.33
+ $X2=0 $Y2=0
cc_494 N_A_111_156#_c_315_n N_A_1248_151#_c_1866_n 0.0190332f $X=6.635 $Y=1.505
+ $X2=0 $Y2=0
cc_495 N_D_M1008_g N_A_161_21#_c_1019_n 0.00880114f $X=2.395 $Y=0.805 $X2=0
+ $Y2=0
cc_496 N_D_c_559_n N_A_161_21#_c_1030_n 0.0237962f $X=2.26 $Y=1.44 $X2=0 $Y2=0
cc_497 N_D_c_560_n N_A_161_21#_c_1030_n 0.0245828f $X=2.395 $Y=1.44 $X2=0 $Y2=0
cc_498 N_D_c_563_n N_A_161_21#_c_1030_n 0.0220859f $X=2.465 $Y=2.34 $X2=0 $Y2=0
cc_499 N_D_c_564_n N_A_161_21#_c_1030_n 8.28749e-19 $X=2.465 $Y=2.34 $X2=0 $Y2=0
cc_500 N_D_M1018_g N_A_161_21#_M1003_g 0.0142331f $X=2.5 $Y=2.875 $X2=0 $Y2=0
cc_501 N_D_c_559_n N_A_161_21#_M1003_g 0.00112944f $X=2.26 $Y=1.44 $X2=0 $Y2=0
cc_502 N_D_c_563_n N_A_161_21#_M1003_g 0.0203793f $X=2.465 $Y=2.34 $X2=0 $Y2=0
cc_503 N_D_c_564_n N_A_161_21#_M1003_g 2.76356e-19 $X=2.465 $Y=2.34 $X2=0 $Y2=0
cc_504 N_D_c_559_n N_A_161_21#_c_1033_n 0.0183762f $X=2.26 $Y=1.44 $X2=0 $Y2=0
cc_505 N_D_M1018_g N_A_161_21#_c_1034_n 7.88709e-19 $X=2.5 $Y=2.875 $X2=0 $Y2=0
cc_506 N_D_c_559_n N_A_161_21#_c_1034_n 0.0265335f $X=2.26 $Y=1.44 $X2=0 $Y2=0
cc_507 N_D_c_563_n N_A_161_21#_c_1034_n 3.03283e-19 $X=2.465 $Y=2.34 $X2=0 $Y2=0
cc_508 N_D_c_559_n N_A_161_21#_c_1035_n 5.11906e-19 $X=2.26 $Y=1.44 $X2=0 $Y2=0
cc_509 N_D_c_564_n N_VPWR_M1002_d 0.00444485f $X=2.465 $Y=2.34 $X2=0 $Y2=0
cc_510 N_D_M1018_g N_VPWR_c_1482_n 0.00798875f $X=2.5 $Y=2.875 $X2=0 $Y2=0
cc_511 N_D_c_563_n N_VPWR_c_1482_n 2.29527e-19 $X=2.465 $Y=2.34 $X2=0 $Y2=0
cc_512 N_D_c_564_n N_VPWR_c_1482_n 0.0290109f $X=2.465 $Y=2.34 $X2=0 $Y2=0
cc_513 N_D_M1018_g N_VPWR_c_1491_n 0.00538679f $X=2.5 $Y=2.875 $X2=0 $Y2=0
cc_514 N_D_M1018_g N_VPWR_c_1479_n 0.00672525f $X=2.5 $Y=2.875 $X2=0 $Y2=0
cc_515 N_D_c_564_n N_VPWR_c_1479_n 0.00836374f $X=2.465 $Y=2.34 $X2=0 $Y2=0
cc_516 N_D_M1008_g N_A_494_119#_c_1626_n 0.00689438f $X=2.395 $Y=0.805 $X2=0
+ $Y2=0
cc_517 N_D_c_559_n N_A_494_119#_c_1626_n 0.0307837f $X=2.26 $Y=1.44 $X2=0 $Y2=0
cc_518 N_D_M1018_g N_A_494_119#_c_1628_n 0.00389131f $X=2.5 $Y=2.875 $X2=0 $Y2=0
cc_519 N_D_c_559_n N_A_494_119#_c_1628_n 0.0129693f $X=2.26 $Y=1.44 $X2=0 $Y2=0
cc_520 N_D_c_563_n N_A_494_119#_c_1628_n 0.00212376f $X=2.465 $Y=2.34 $X2=0
+ $Y2=0
cc_521 N_D_c_564_n N_A_494_119#_c_1628_n 0.0258047f $X=2.465 $Y=2.34 $X2=0 $Y2=0
cc_522 N_D_M1018_g N_A_494_119#_c_1644_n 0.00515634f $X=2.5 $Y=2.875 $X2=0 $Y2=0
cc_523 N_D_c_563_n N_A_494_119#_c_1644_n 0.00159909f $X=2.465 $Y=2.34 $X2=0
+ $Y2=0
cc_524 N_D_c_559_n N_A_494_119#_c_1629_n 0.0126169f $X=2.26 $Y=1.44 $X2=0 $Y2=0
cc_525 N_D_c_563_n N_A_494_119#_c_1629_n 2.67811e-19 $X=2.465 $Y=2.34 $X2=0
+ $Y2=0
cc_526 N_D_M1008_g N_VGND_c_1713_n 6.92788e-19 $X=2.395 $Y=0.805 $X2=0 $Y2=0
cc_527 N_A_708_93#_c_616_n N_A_580_119#_M1012_g 0.0105245f $X=3.9 $Y=1.21 $X2=0
+ $Y2=0
cc_528 N_A_708_93#_c_618_n N_A_580_119#_M1012_g 0.00586305f $X=4.445 $Y=1.5
+ $X2=0 $Y2=0
cc_529 N_A_708_93#_c_620_n N_A_580_119#_M1012_g 0.0014272f $X=4.53 $Y=1.12 $X2=0
+ $Y2=0
cc_530 N_A_708_93#_c_629_n N_A_580_119#_M1012_g 0.00423741f $X=4.22 $Y=2.175
+ $X2=0 $Y2=0
cc_531 N_A_708_93#_c_625_n N_A_580_119#_c_731_n 0.00108412f $X=4.365 $Y=2.685
+ $X2=0 $Y2=0
cc_532 N_A_708_93#_c_662_p N_A_580_119#_c_731_n 0.0179406f $X=5.46 $Y=2.85 $X2=0
+ $Y2=0
cc_533 N_A_708_93#_c_662_p N_A_580_119#_c_732_n 0.0162869f $X=5.46 $Y=2.85 $X2=0
+ $Y2=0
cc_534 N_A_708_93#_c_626_n N_A_580_119#_c_734_n 0.0242619f $X=4.22 $Y=2.34 $X2=0
+ $Y2=0
cc_535 N_A_708_93#_c_627_n N_A_580_119#_c_734_n 0.00224863f $X=4.365 $Y=2.34
+ $X2=0 $Y2=0
cc_536 N_A_708_93#_c_615_n N_A_580_119#_c_722_n 4.07506e-19 $X=3.615 $Y=1.135
+ $X2=0 $Y2=0
cc_537 N_A_708_93#_c_622_n N_A_580_119#_c_767_n 0.00146699f $X=3.72 $Y=2.555
+ $X2=0 $Y2=0
cc_538 N_A_708_93#_c_622_n N_A_580_119#_c_736_n 0.00730336f $X=3.72 $Y=2.555
+ $X2=0 $Y2=0
cc_539 N_A_708_93#_c_623_n N_A_580_119#_c_736_n 0.00489694f $X=4.055 $Y=2.48
+ $X2=0 $Y2=0
cc_540 N_A_708_93#_c_624_n N_A_580_119#_c_736_n 0.00646013f $X=3.795 $Y=2.48
+ $X2=0 $Y2=0
cc_541 N_A_708_93#_c_625_n N_A_580_119#_c_736_n 0.00764331f $X=4.365 $Y=2.685
+ $X2=0 $Y2=0
cc_542 N_A_708_93#_c_627_n N_A_580_119#_c_736_n 0.00145062f $X=4.365 $Y=2.34
+ $X2=0 $Y2=0
cc_543 N_A_708_93#_c_623_n N_A_580_119#_c_737_n 0.00596752f $X=4.055 $Y=2.48
+ $X2=0 $Y2=0
cc_544 N_A_708_93#_c_624_n N_A_580_119#_c_737_n 0.00151832f $X=3.795 $Y=2.48
+ $X2=0 $Y2=0
cc_545 N_A_708_93#_c_627_n N_A_580_119#_c_737_n 0.0219334f $X=4.365 $Y=2.34
+ $X2=0 $Y2=0
cc_546 N_A_708_93#_c_629_n N_A_580_119#_c_737_n 0.00839922f $X=4.22 $Y=2.175
+ $X2=0 $Y2=0
cc_547 N_A_708_93#_c_623_n N_A_580_119#_c_738_n 0.00247236f $X=4.055 $Y=2.48
+ $X2=0 $Y2=0
cc_548 N_A_708_93#_c_618_n N_A_580_119#_c_738_n 0.0490668f $X=4.445 $Y=1.5 $X2=0
+ $Y2=0
cc_549 N_A_708_93#_c_626_n N_A_580_119#_c_738_n 0.00362719f $X=4.22 $Y=2.34
+ $X2=0 $Y2=0
cc_550 N_A_708_93#_c_627_n N_A_580_119#_c_738_n 0.018299f $X=4.365 $Y=2.34 $X2=0
+ $Y2=0
cc_551 N_A_708_93#_c_621_n N_A_580_119#_c_738_n 0.00297477f $X=4.065 $Y=1.665
+ $X2=0 $Y2=0
cc_552 N_A_708_93#_c_629_n N_A_580_119#_c_738_n 0.0137645f $X=4.22 $Y=2.175
+ $X2=0 $Y2=0
cc_553 N_A_708_93#_c_616_n N_A_580_119#_c_739_n 0.0019346f $X=3.9 $Y=1.21 $X2=0
+ $Y2=0
cc_554 N_A_708_93#_c_618_n N_A_580_119#_c_739_n 0.00425068f $X=4.445 $Y=1.5
+ $X2=0 $Y2=0
cc_555 N_A_708_93#_c_621_n N_A_580_119#_c_739_n 0.00154252f $X=4.065 $Y=1.665
+ $X2=0 $Y2=0
cc_556 N_A_708_93#_c_621_n N_A_580_119#_c_724_n 3.36841e-19 $X=4.065 $Y=1.665
+ $X2=0 $Y2=0
cc_557 N_A_708_93#_c_629_n N_A_580_119#_c_724_n 4.25934e-19 $X=4.22 $Y=2.175
+ $X2=0 $Y2=0
cc_558 N_A_708_93#_c_662_p N_A_580_119#_c_741_n 0.0234808f $X=5.46 $Y=2.85 $X2=0
+ $Y2=0
cc_559 N_A_708_93#_c_626_n N_A_580_119#_c_741_n 3.23013e-19 $X=4.22 $Y=2.34
+ $X2=0 $Y2=0
cc_560 N_A_708_93#_c_627_n N_A_580_119#_c_741_n 0.0209299f $X=4.365 $Y=2.34
+ $X2=0 $Y2=0
cc_561 N_A_708_93#_c_629_n N_A_580_119#_c_741_n 0.00119508f $X=4.22 $Y=2.175
+ $X2=0 $Y2=0
cc_562 N_A_708_93#_c_618_n N_A_580_119#_c_742_n 2.57655e-19 $X=4.445 $Y=1.5
+ $X2=0 $Y2=0
cc_563 N_A_708_93#_c_629_n N_A_580_119#_c_742_n 0.0100022f $X=4.22 $Y=2.175
+ $X2=0 $Y2=0
cc_564 N_A_708_93#_c_662_p N_SET_B_c_903_n 0.0210746f $X=5.46 $Y=2.85 $X2=0
+ $Y2=0
cc_565 N_A_708_93#_c_662_p N_SET_B_c_904_n 7.75395e-19 $X=5.46 $Y=2.85 $X2=0
+ $Y2=0
cc_566 N_A_708_93#_c_662_p N_SET_B_c_905_n 0.00408458f $X=5.46 $Y=2.85 $X2=0
+ $Y2=0
cc_567 N_A_708_93#_c_615_n N_A_161_21#_M1000_g 0.0399478f $X=3.615 $Y=1.135
+ $X2=0 $Y2=0
cc_568 N_A_708_93#_c_615_n N_A_161_21#_c_1021_n 0.0104164f $X=3.615 $Y=1.135
+ $X2=0 $Y2=0
cc_569 N_A_708_93#_c_625_n N_VPWR_M1031_d 0.00101379f $X=4.365 $Y=2.685 $X2=0
+ $Y2=0
cc_570 N_A_708_93#_c_700_p N_VPWR_M1031_d 0.00890198f $X=4.45 $Y=2.85 $X2=0
+ $Y2=0
cc_571 N_A_708_93#_c_662_p N_VPWR_M1031_d 0.0278467f $X=5.46 $Y=2.85 $X2=0 $Y2=0
cc_572 N_A_708_93#_c_622_n N_VPWR_c_1483_n 0.01035f $X=3.72 $Y=2.555 $X2=0 $Y2=0
cc_573 N_A_708_93#_c_623_n N_VPWR_c_1483_n 0.00628999f $X=4.055 $Y=2.48 $X2=0
+ $Y2=0
cc_574 N_A_708_93#_c_700_p N_VPWR_c_1483_n 0.0155039f $X=4.45 $Y=2.85 $X2=0
+ $Y2=0
cc_575 N_A_708_93#_c_622_n N_VPWR_c_1491_n 0.00351296f $X=3.72 $Y=2.555 $X2=0
+ $Y2=0
cc_576 N_A_708_93#_c_700_p N_VPWR_c_1492_n 0.00838606f $X=4.45 $Y=2.85 $X2=0
+ $Y2=0
cc_577 N_A_708_93#_c_662_p N_VPWR_c_1492_n 0.0501585f $X=5.46 $Y=2.85 $X2=0
+ $Y2=0
cc_578 N_A_708_93#_c_626_n N_VPWR_c_1492_n 0.0036324f $X=4.22 $Y=2.34 $X2=0
+ $Y2=0
cc_579 N_A_708_93#_M1029_d N_VPWR_c_1479_n 0.002513f $X=5.32 $Y=2.665 $X2=0
+ $Y2=0
cc_580 N_A_708_93#_c_622_n N_VPWR_c_1479_n 0.00406706f $X=3.72 $Y=2.555 $X2=0
+ $Y2=0
cc_581 N_A_708_93#_c_700_p N_VPWR_c_1479_n 0.00633924f $X=4.45 $Y=2.85 $X2=0
+ $Y2=0
cc_582 N_A_708_93#_c_662_p N_VPWR_c_1479_n 0.0403723f $X=5.46 $Y=2.85 $X2=0
+ $Y2=0
cc_583 N_A_708_93#_c_626_n N_VPWR_c_1479_n 0.00463141f $X=4.22 $Y=2.34 $X2=0
+ $Y2=0
cc_584 N_A_708_93#_c_627_n N_VPWR_c_1479_n 0.00489801f $X=4.365 $Y=2.34 $X2=0
+ $Y2=0
cc_585 N_A_708_93#_c_615_n N_VGND_c_1714_n 0.00305576f $X=3.615 $Y=1.135 $X2=0
+ $Y2=0
cc_586 N_A_708_93#_c_616_n N_VGND_c_1714_n 0.00129224f $X=3.9 $Y=1.21 $X2=0
+ $Y2=0
cc_587 N_A_708_93#_c_615_n N_VGND_c_1729_n 9.39239e-19 $X=3.615 $Y=1.135 $X2=0
+ $Y2=0
cc_588 N_A_580_119#_M1012_g N_SET_B_M1009_g 0.0533533f $X=4.745 $Y=1.055 $X2=0
+ $Y2=0
cc_589 N_A_580_119#_M1026_g N_SET_B_M1009_g 0.0158251f $X=5.63 $Y=0.945 $X2=0
+ $Y2=0
cc_590 N_A_580_119#_M1012_g N_SET_B_c_892_n 0.00792255f $X=4.745 $Y=1.055 $X2=0
+ $Y2=0
cc_591 N_A_580_119#_c_721_n N_SET_B_c_892_n 0.00587455f $X=5.705 $Y=1.55 $X2=0
+ $Y2=0
cc_592 N_A_580_119#_c_724_n N_SET_B_c_892_n 0.00466693f $X=4.83 $Y=1.935 $X2=0
+ $Y2=0
cc_593 N_A_580_119#_c_742_n N_SET_B_c_892_n 0.00960646f $X=4.76 $Y=2 $X2=0 $Y2=0
cc_594 N_A_580_119#_c_725_n N_SET_B_c_892_n 0.0027072f $X=6.13 $Y=1.85 $X2=0
+ $Y2=0
cc_595 N_A_580_119#_c_727_n N_SET_B_c_892_n 0.0112183f $X=5.675 $Y=1.805 $X2=0
+ $Y2=0
cc_596 N_A_580_119#_c_728_n N_SET_B_c_892_n 0.00233093f $X=5.845 $Y=1.805 $X2=0
+ $Y2=0
cc_597 N_A_580_119#_c_730_n N_SET_B_M1013_g 0.0214933f $X=5.17 $Y=2.48 $X2=0
+ $Y2=0
cc_598 N_A_580_119#_c_734_n N_SET_B_M1013_g 0.0021575f $X=4.76 $Y=2.405 $X2=0
+ $Y2=0
cc_599 N_A_580_119#_M1026_g N_SET_B_c_894_n 0.00587455f $X=5.63 $Y=0.945 $X2=0
+ $Y2=0
cc_600 N_A_580_119#_c_727_n N_SET_B_c_894_n 0.00438151f $X=5.675 $Y=1.805 $X2=0
+ $Y2=0
cc_601 N_A_580_119#_c_730_n N_SET_B_c_903_n 0.00681257f $X=5.17 $Y=2.48 $X2=0
+ $Y2=0
cc_602 N_A_580_119#_M1032_g N_SET_B_c_903_n 7.02785e-19 $X=6.22 $Y=2.665 $X2=0
+ $Y2=0
cc_603 N_A_580_119#_c_734_n N_SET_B_c_903_n 8.15853e-19 $X=4.76 $Y=2.405 $X2=0
+ $Y2=0
cc_604 N_A_580_119#_c_741_n N_SET_B_c_903_n 0.041638f $X=4.76 $Y=2 $X2=0 $Y2=0
cc_605 N_A_580_119#_c_742_n N_SET_B_c_903_n 2.82462e-19 $X=4.76 $Y=2 $X2=0 $Y2=0
cc_606 N_A_580_119#_c_727_n N_SET_B_c_903_n 0.0240964f $X=5.675 $Y=1.805 $X2=0
+ $Y2=0
cc_607 N_A_580_119#_c_728_n N_SET_B_c_903_n 0.00546859f $X=5.845 $Y=1.805 $X2=0
+ $Y2=0
cc_608 N_A_580_119#_c_730_n N_SET_B_c_904_n 0.0101122f $X=5.17 $Y=2.48 $X2=0
+ $Y2=0
cc_609 N_A_580_119#_c_721_n N_SET_B_c_904_n 0.00506641f $X=5.705 $Y=1.55 $X2=0
+ $Y2=0
cc_610 N_A_580_119#_M1032_g N_SET_B_c_904_n 0.0291165f $X=6.22 $Y=2.665 $X2=0
+ $Y2=0
cc_611 N_A_580_119#_c_734_n N_SET_B_c_904_n 0.00960646f $X=4.76 $Y=2.405 $X2=0
+ $Y2=0
cc_612 N_A_580_119#_c_741_n N_SET_B_c_904_n 0.00178648f $X=4.76 $Y=2 $X2=0 $Y2=0
cc_613 N_A_580_119#_c_727_n N_SET_B_c_904_n 0.00621671f $X=5.675 $Y=1.805 $X2=0
+ $Y2=0
cc_614 N_A_580_119#_c_728_n N_SET_B_c_904_n 0.00393927f $X=5.845 $Y=1.805 $X2=0
+ $Y2=0
cc_615 N_A_580_119#_c_748_n N_SET_B_c_904_n 0.00304207f $X=6.13 $Y=2.015 $X2=0
+ $Y2=0
cc_616 N_A_580_119#_c_720_n N_SET_B_c_905_n 3.1477e-19 $X=5.965 $Y=1.55 $X2=0
+ $Y2=0
cc_617 N_A_580_119#_M1032_g N_SET_B_c_905_n 0.018283f $X=6.22 $Y=2.665 $X2=0
+ $Y2=0
cc_618 N_A_580_119#_c_727_n N_SET_B_c_905_n 0.00478359f $X=5.675 $Y=1.805 $X2=0
+ $Y2=0
cc_619 N_A_580_119#_c_728_n N_SET_B_c_905_n 0.0319418f $X=5.845 $Y=1.805 $X2=0
+ $Y2=0
cc_620 N_A_580_119#_c_748_n N_SET_B_c_905_n 0.0041636f $X=6.13 $Y=2.015 $X2=0
+ $Y2=0
cc_621 N_A_580_119#_c_723_n N_A_161_21#_c_1030_n 0.00455448f $X=3.145 $Y=2.485
+ $X2=0 $Y2=0
cc_622 N_A_580_119#_c_726_n N_A_161_21#_c_1030_n 4.28437e-19 $X=3.087 $Y=1.585
+ $X2=0 $Y2=0
cc_623 N_A_580_119#_c_745_n N_A_161_21#_M1003_g 0.00137314f $X=3.185 $Y=2.57
+ $X2=0 $Y2=0
cc_624 N_A_580_119#_c_722_n N_A_161_21#_M1000_g 0.00102738f $X=3.04 $Y=0.81
+ $X2=0 $Y2=0
cc_625 N_A_580_119#_c_726_n N_A_161_21#_M1000_g 0.00127728f $X=3.087 $Y=1.585
+ $X2=0 $Y2=0
cc_626 N_A_580_119#_M1012_g N_A_161_21#_c_1021_n 0.00314123f $X=4.745 $Y=1.055
+ $X2=0 $Y2=0
cc_627 N_A_580_119#_M1026_g N_A_161_21#_c_1021_n 0.00907339f $X=5.63 $Y=0.945
+ $X2=0 $Y2=0
cc_628 N_A_580_119#_M1032_g N_A_1331_151#_c_1266_n 2.42085e-19 $X=6.22 $Y=2.665
+ $X2=0 $Y2=0
cc_629 N_A_580_119#_c_767_n N_VPWR_c_1483_n 0.00737112f $X=3.145 $Y=2.885 $X2=0
+ $Y2=0
cc_630 N_A_580_119#_c_736_n N_VPWR_c_1483_n 0.0131185f $X=3.785 $Y=2.57 $X2=0
+ $Y2=0
cc_631 N_A_580_119#_M1032_g N_VPWR_c_1484_n 0.0091284f $X=6.22 $Y=2.665 $X2=0
+ $Y2=0
cc_632 N_A_580_119#_c_767_n N_VPWR_c_1491_n 0.0132057f $X=3.145 $Y=2.885 $X2=0
+ $Y2=0
cc_633 N_A_580_119#_c_736_n N_VPWR_c_1491_n 0.00723599f $X=3.785 $Y=2.57 $X2=0
+ $Y2=0
cc_634 N_A_580_119#_c_732_n N_VPWR_c_1492_n 0.00363139f $X=5.245 $Y=2.555 $X2=0
+ $Y2=0
cc_635 N_A_580_119#_M1032_g N_VPWR_c_1493_n 0.00554242f $X=6.22 $Y=2.665 $X2=0
+ $Y2=0
cc_636 N_A_580_119#_M1003_d N_VPWR_c_1479_n 0.00420763f $X=3.005 $Y=2.665 $X2=0
+ $Y2=0
cc_637 N_A_580_119#_c_732_n N_VPWR_c_1479_n 0.00666269f $X=5.245 $Y=2.555 $X2=0
+ $Y2=0
cc_638 N_A_580_119#_M1032_g N_VPWR_c_1479_n 0.00548042f $X=6.22 $Y=2.665 $X2=0
+ $Y2=0
cc_639 N_A_580_119#_c_767_n N_VPWR_c_1479_n 0.00938117f $X=3.145 $Y=2.885 $X2=0
+ $Y2=0
cc_640 N_A_580_119#_c_736_n N_VPWR_c_1479_n 0.0123717f $X=3.785 $Y=2.57 $X2=0
+ $Y2=0
cc_641 N_A_580_119#_c_723_n N_A_494_119#_c_1626_n 0.00929078f $X=3.145 $Y=2.485
+ $X2=0 $Y2=0
cc_642 N_A_580_119#_c_726_n N_A_494_119#_c_1626_n 0.0273025f $X=3.087 $Y=1.585
+ $X2=0 $Y2=0
cc_643 N_A_580_119#_c_723_n N_A_494_119#_c_1628_n 0.0392613f $X=3.145 $Y=2.485
+ $X2=0 $Y2=0
cc_644 N_A_580_119#_c_767_n N_A_494_119#_c_1628_n 0.00252201f $X=3.145 $Y=2.885
+ $X2=0 $Y2=0
cc_645 N_A_580_119#_c_745_n N_A_494_119#_c_1628_n 0.0137141f $X=3.185 $Y=2.57
+ $X2=0 $Y2=0
cc_646 N_A_580_119#_c_722_n N_A_494_119#_c_1634_n 0.0273025f $X=3.04 $Y=0.81
+ $X2=0 $Y2=0
cc_647 N_A_580_119#_c_723_n N_A_494_119#_c_1629_n 0.0127456f $X=3.145 $Y=2.485
+ $X2=0 $Y2=0
cc_648 N_A_580_119#_M1026_g N_VGND_c_1715_n 0.00483343f $X=5.63 $Y=0.945 $X2=0
+ $Y2=0
cc_649 N_A_580_119#_M1026_g N_VGND_c_1729_n 9.49986e-19 $X=5.63 $Y=0.945 $X2=0
+ $Y2=0
cc_650 N_A_580_119#_M1026_g N_A_1141_125#_c_1841_n 0.00483343f $X=5.63 $Y=0.945
+ $X2=0 $Y2=0
cc_651 N_SET_B_M1009_g N_A_161_21#_c_1021_n 0.00462072f $X=5.105 $Y=1.055 $X2=0
+ $Y2=0
cc_652 N_SET_B_c_899_n N_A_161_21#_M1033_g 0.00731076f $X=7.51 $Y=2.96 $X2=0
+ $Y2=0
cc_653 N_SET_B_c_900_n N_A_161_21#_M1033_g 0.00789327f $X=7.595 $Y=2.845 $X2=0
+ $Y2=0
cc_654 N_SET_B_c_901_n N_A_161_21#_M1033_g 0.00337654f $X=7.68 $Y=1.88 $X2=0
+ $Y2=0
cc_655 N_SET_B_M1005_g N_A_1535_177#_M1030_g 0.00726237f $X=8.57 $Y=0.565 $X2=0
+ $Y2=0
cc_656 N_SET_B_c_899_n N_A_1535_177#_M1030_g 0.00691892f $X=7.51 $Y=2.96 $X2=0
+ $Y2=0
cc_657 N_SET_B_c_900_n N_A_1535_177#_M1030_g 0.0160245f $X=7.595 $Y=2.845 $X2=0
+ $Y2=0
cc_658 N_SET_B_c_901_n N_A_1535_177#_M1030_g 0.00306915f $X=7.68 $Y=1.88 $X2=0
+ $Y2=0
cc_659 N_SET_B_c_902_n N_A_1535_177#_M1030_g 0.0175327f $X=8.27 $Y=1.88 $X2=0
+ $Y2=0
cc_660 N_SET_B_c_906_n N_A_1535_177#_M1030_g 0.0296319f $X=8.57 $Y=1.88 $X2=0
+ $Y2=0
cc_661 N_SET_B_M1015_g N_A_1535_177#_c_1169_n 0.00914649f $X=8.18 $Y=2.455 $X2=0
+ $Y2=0
cc_662 N_SET_B_c_899_n N_A_1535_177#_c_1170_n 0.00162339f $X=7.51 $Y=2.96 $X2=0
+ $Y2=0
cc_663 N_SET_B_M1005_g N_A_1535_177#_c_1164_n 0.0623931f $X=8.57 $Y=0.565 $X2=0
+ $Y2=0
cc_664 N_SET_B_M1005_g N_A_1535_177#_c_1165_n 0.0169542f $X=8.57 $Y=0.565 $X2=0
+ $Y2=0
cc_665 N_SET_B_M1015_g N_A_1535_177#_c_1171_n 0.00405554f $X=8.18 $Y=2.455 $X2=0
+ $Y2=0
cc_666 N_SET_B_M1015_g N_A_1535_177#_c_1172_n 0.00145495f $X=8.18 $Y=2.455 $X2=0
+ $Y2=0
cc_667 N_SET_B_M1005_g N_A_1535_177#_c_1166_n 0.00547862f $X=8.57 $Y=0.565 $X2=0
+ $Y2=0
cc_668 N_SET_B_M1015_g N_A_1535_177#_c_1173_n 4.34705e-19 $X=8.18 $Y=2.455 $X2=0
+ $Y2=0
cc_669 N_SET_B_c_906_n N_A_1535_177#_c_1167_n 0.00337248f $X=8.57 $Y=1.88 $X2=0
+ $Y2=0
cc_670 N_SET_B_c_899_n N_A_1331_151#_M1007_d 0.00527599f $X=7.51 $Y=2.96 $X2=0
+ $Y2=0
cc_671 N_SET_B_M1005_g N_A_1331_151#_c_1242_n 0.00528014f $X=8.57 $Y=0.565 $X2=0
+ $Y2=0
cc_672 N_SET_B_M1005_g N_A_1331_151#_c_1244_n 0.00620571f $X=8.57 $Y=0.565 $X2=0
+ $Y2=0
cc_673 N_SET_B_c_901_n N_A_1331_151#_c_1244_n 0.0115691f $X=7.68 $Y=1.88 $X2=0
+ $Y2=0
cc_674 N_SET_B_c_902_n N_A_1331_151#_c_1244_n 0.04166f $X=8.27 $Y=1.88 $X2=0
+ $Y2=0
cc_675 N_SET_B_c_906_n N_A_1331_151#_c_1244_n 0.00799579f $X=8.57 $Y=1.88 $X2=0
+ $Y2=0
cc_676 N_SET_B_M1015_g N_A_1331_151#_c_1245_n 0.00546311f $X=8.18 $Y=2.455 $X2=0
+ $Y2=0
cc_677 N_SET_B_M1005_g N_A_1331_151#_c_1245_n 0.0132061f $X=8.57 $Y=0.565 $X2=0
+ $Y2=0
cc_678 N_SET_B_c_902_n N_A_1331_151#_c_1245_n 0.0249855f $X=8.27 $Y=1.88 $X2=0
+ $Y2=0
cc_679 N_SET_B_c_906_n N_A_1331_151#_c_1245_n 0.0136182f $X=8.57 $Y=1.88 $X2=0
+ $Y2=0
cc_680 N_SET_B_c_911_n N_A_1331_151#_c_1266_n 0.00858734f $X=6.415 $Y=2.845
+ $X2=0 $Y2=0
cc_681 N_SET_B_c_899_n N_A_1331_151#_c_1266_n 0.0210891f $X=7.51 $Y=2.96 $X2=0
+ $Y2=0
cc_682 N_SET_B_c_905_n N_A_1331_151#_c_1266_n 0.0106706f $X=6.33 $Y=2.367 $X2=0
+ $Y2=0
cc_683 N_SET_B_c_900_n N_A_1331_151#_c_1250_n 0.0273392f $X=7.595 $Y=2.845 $X2=0
+ $Y2=0
cc_684 N_SET_B_c_901_n N_A_1331_151#_c_1250_n 0.0163896f $X=7.68 $Y=1.88 $X2=0
+ $Y2=0
cc_685 N_SET_B_c_905_n N_A_1331_151#_c_1250_n 0.00162207f $X=6.33 $Y=2.367 $X2=0
+ $Y2=0
cc_686 N_SET_B_M1015_g N_A_1331_151#_c_1268_n 5.61829e-19 $X=8.18 $Y=2.455 $X2=0
+ $Y2=0
cc_687 N_SET_B_c_900_n N_A_1331_151#_c_1268_n 9.49668e-19 $X=7.595 $Y=2.845
+ $X2=0 $Y2=0
cc_688 N_SET_B_c_902_n N_A_1331_151#_c_1268_n 0.00568604f $X=8.27 $Y=1.88 $X2=0
+ $Y2=0
cc_689 N_SET_B_c_906_n N_A_1331_151#_c_1268_n 0.0092019f $X=8.57 $Y=1.88 $X2=0
+ $Y2=0
cc_690 N_SET_B_M1005_g N_A_1331_151#_c_1252_n 0.00668968f $X=8.57 $Y=0.565 $X2=0
+ $Y2=0
cc_691 N_SET_B_M1005_g N_A_1331_151#_c_1269_n 5.03855e-19 $X=8.57 $Y=0.565 $X2=0
+ $Y2=0
cc_692 N_SET_B_c_906_n N_A_1331_151#_c_1253_n 0.00528014f $X=8.57 $Y=1.88 $X2=0
+ $Y2=0
cc_693 N_SET_B_c_905_n N_VPWR_M1013_d 0.00526696f $X=6.33 $Y=2.367 $X2=0 $Y2=0
cc_694 N_SET_B_M1013_g N_VPWR_c_1484_n 0.00889946f $X=5.675 $Y=2.875 $X2=0 $Y2=0
cc_695 N_SET_B_c_905_n N_VPWR_c_1484_n 0.0221538f $X=6.33 $Y=2.367 $X2=0 $Y2=0
cc_696 N_SET_B_M1015_g N_VPWR_c_1485_n 0.00357865f $X=8.18 $Y=2.455 $X2=0 $Y2=0
cc_697 N_SET_B_c_899_n N_VPWR_c_1485_n 0.0186494f $X=7.51 $Y=2.96 $X2=0 $Y2=0
cc_698 N_SET_B_c_900_n N_VPWR_c_1485_n 0.0262106f $X=7.595 $Y=2.845 $X2=0 $Y2=0
cc_699 N_SET_B_c_902_n N_VPWR_c_1485_n 0.0137875f $X=8.27 $Y=1.88 $X2=0 $Y2=0
cc_700 N_SET_B_M1013_g N_VPWR_c_1492_n 0.00575161f $X=5.675 $Y=2.875 $X2=0 $Y2=0
cc_701 N_SET_B_c_899_n N_VPWR_c_1493_n 0.0742518f $X=7.51 $Y=2.96 $X2=0 $Y2=0
cc_702 N_SET_B_c_1002_p N_VPWR_c_1493_n 0.0111868f $X=6.5 $Y=2.96 $X2=0 $Y2=0
cc_703 N_SET_B_M1013_g N_VPWR_c_1479_n 0.0066471f $X=5.675 $Y=2.875 $X2=0 $Y2=0
cc_704 N_SET_B_M1015_g N_VPWR_c_1479_n 9.03821e-19 $X=8.18 $Y=2.455 $X2=0 $Y2=0
cc_705 N_SET_B_c_899_n N_VPWR_c_1479_n 0.0441172f $X=7.51 $Y=2.96 $X2=0 $Y2=0
cc_706 N_SET_B_c_1002_p N_VPWR_c_1479_n 0.00660921f $X=6.5 $Y=2.96 $X2=0 $Y2=0
cc_707 N_SET_B_c_905_n N_VPWR_c_1479_n 0.0146307f $X=6.33 $Y=2.367 $X2=0 $Y2=0
cc_708 N_SET_B_c_911_n A_1259_449# 0.0056188f $X=6.415 $Y=2.845 $X2=-0.19
+ $Y2=-0.245
cc_709 N_SET_B_c_899_n A_1259_449# 0.00628051f $X=7.51 $Y=2.96 $X2=-0.19
+ $Y2=-0.245
cc_710 N_SET_B_c_1002_p A_1259_449# 0.00333126f $X=6.5 $Y=2.96 $X2=-0.19
+ $Y2=-0.245
cc_711 N_SET_B_c_905_n A_1259_449# 0.00983723f $X=6.33 $Y=2.367 $X2=-0.19
+ $Y2=-0.245
cc_712 N_SET_B_c_900_n A_1472_449# 0.00481456f $X=7.595 $Y=2.845 $X2=-0.19
+ $Y2=-0.245
cc_713 N_SET_B_M1009_g N_VGND_c_1715_n 0.00349814f $X=5.105 $Y=1.055 $X2=0 $Y2=0
cc_714 N_SET_B_M1005_g N_VGND_c_1716_n 0.0125082f $X=8.57 $Y=0.565 $X2=0 $Y2=0
cc_715 N_SET_B_M1005_g N_VGND_c_1723_n 0.00393414f $X=8.57 $Y=0.565 $X2=0 $Y2=0
cc_716 N_SET_B_M1009_g N_VGND_c_1729_n 9.7053e-19 $X=5.105 $Y=1.055 $X2=0 $Y2=0
cc_717 N_SET_B_M1005_g N_VGND_c_1729_n 0.00765569f $X=8.57 $Y=0.565 $X2=0 $Y2=0
cc_718 N_A_161_21#_c_1025_n N_A_1535_177#_M1030_g 0.0547368f $X=7.285 $Y=1.36
+ $X2=0 $Y2=0
cc_719 N_A_161_21#_M1020_g N_A_1535_177#_c_1165_n 8.20375e-19 $X=7.125 $Y=0.855
+ $X2=0 $Y2=0
cc_720 N_A_161_21#_M1020_g N_A_1535_177#_c_1167_n 0.0110772f $X=7.125 $Y=0.855
+ $X2=0 $Y2=0
cc_721 N_A_161_21#_M1020_g N_A_1331_151#_c_1243_n 0.00375521f $X=7.125 $Y=0.855
+ $X2=0 $Y2=0
cc_722 N_A_161_21#_c_1025_n N_A_1331_151#_c_1243_n 9.22829e-19 $X=7.285 $Y=1.36
+ $X2=0 $Y2=0
cc_723 N_A_161_21#_M1033_g N_A_1331_151#_c_1244_n 0.00850597f $X=7.285 $Y=2.455
+ $X2=0 $Y2=0
cc_724 N_A_161_21#_c_1025_n N_A_1331_151#_c_1244_n 0.00890136f $X=7.285 $Y=1.36
+ $X2=0 $Y2=0
cc_725 N_A_161_21#_M1020_g N_A_1331_151#_c_1273_n 0.0058868f $X=7.125 $Y=0.855
+ $X2=0 $Y2=0
cc_726 N_A_161_21#_M1033_g N_A_1331_151#_c_1250_n 0.0164844f $X=7.285 $Y=2.455
+ $X2=0 $Y2=0
cc_727 N_A_161_21#_c_1025_n N_A_1331_151#_c_1251_n 0.00489927f $X=7.285 $Y=1.36
+ $X2=0 $Y2=0
cc_728 N_A_161_21#_c_1034_n N_VPWR_c_1482_n 0.0179627f $X=1.6 $Y=2.47 $X2=0
+ $Y2=0
cc_729 N_A_161_21#_c_1034_n N_VPWR_c_1490_n 0.0120829f $X=1.6 $Y=2.47 $X2=0
+ $Y2=0
cc_730 N_A_161_21#_M1003_g N_VPWR_c_1491_n 0.00524086f $X=2.93 $Y=2.875 $X2=0
+ $Y2=0
cc_731 N_A_161_21#_M1003_g N_VPWR_c_1479_n 0.00961687f $X=2.93 $Y=2.875 $X2=0
+ $Y2=0
cc_732 N_A_161_21#_c_1034_n N_VPWR_c_1479_n 0.0090757f $X=1.6 $Y=2.47 $X2=0
+ $Y2=0
cc_733 N_A_161_21#_c_1030_n N_A_494_119#_c_1626_n 0.00140227f $X=2.855 $Y=1.89
+ $X2=0 $Y2=0
cc_734 N_A_161_21#_c_1030_n N_A_494_119#_c_1628_n 0.00495804f $X=2.855 $Y=1.89
+ $X2=0 $Y2=0
cc_735 N_A_161_21#_M1003_g N_A_494_119#_c_1628_n 0.0149657f $X=2.93 $Y=2.875
+ $X2=0 $Y2=0
cc_736 N_A_161_21#_M1003_g N_A_494_119#_c_1644_n 0.00397142f $X=2.93 $Y=2.875
+ $X2=0 $Y2=0
cc_737 N_A_161_21#_c_1030_n N_A_494_119#_c_1629_n 0.0121617f $X=2.855 $Y=1.89
+ $X2=0 $Y2=0
cc_738 N_A_161_21#_c_1018_n N_VGND_c_1712_n 0.00420742f $X=1.06 $Y=1.815 $X2=0
+ $Y2=0
cc_739 N_A_161_21#_c_1026_n N_VGND_c_1712_n 0.011475f $X=1.205 $Y=0.39 $X2=0
+ $Y2=0
cc_740 N_A_161_21#_c_1028_n N_VGND_c_1712_n 0.00537711f $X=0.97 $Y=0.18 $X2=0
+ $Y2=0
cc_741 N_A_161_21#_c_1019_n N_VGND_c_1713_n 0.0256696f $X=3.18 $Y=0.18 $X2=0
+ $Y2=0
cc_742 N_A_161_21#_c_1026_n N_VGND_c_1713_n 0.0209779f $X=1.205 $Y=0.39 $X2=0
+ $Y2=0
cc_743 N_A_161_21#_c_1027_n N_VGND_c_1713_n 0.0148339f $X=1.37 $Y=0.78 $X2=0
+ $Y2=0
cc_744 N_A_161_21#_c_1028_n N_VGND_c_1713_n 5.52035e-19 $X=0.97 $Y=0.18 $X2=0
+ $Y2=0
cc_745 N_A_161_21#_M1000_g N_VGND_c_1714_n 0.0021727f $X=3.255 $Y=0.805 $X2=0
+ $Y2=0
cc_746 N_A_161_21#_c_1021_n N_VGND_c_1714_n 0.0186898f $X=7.05 $Y=0.18 $X2=0
+ $Y2=0
cc_747 N_A_161_21#_c_1021_n N_VGND_c_1715_n 0.022762f $X=7.05 $Y=0.18 $X2=0
+ $Y2=0
cc_748 N_A_161_21#_c_1019_n N_VGND_c_1719_n 0.0432762f $X=3.18 $Y=0.18 $X2=0
+ $Y2=0
cc_749 N_A_161_21#_c_1021_n N_VGND_c_1721_n 0.0369547f $X=7.05 $Y=0.18 $X2=0
+ $Y2=0
cc_750 N_A_161_21#_c_1021_n N_VGND_c_1723_n 0.0382127f $X=7.05 $Y=0.18 $X2=0
+ $Y2=0
cc_751 N_A_161_21#_c_1026_n N_VGND_c_1725_n 0.0414112f $X=1.205 $Y=0.39 $X2=0
+ $Y2=0
cc_752 N_A_161_21#_c_1028_n N_VGND_c_1725_n 0.0209993f $X=0.97 $Y=0.18 $X2=0
+ $Y2=0
cc_753 N_A_161_21#_c_1019_n N_VGND_c_1729_n 0.0477761f $X=3.18 $Y=0.18 $X2=0
+ $Y2=0
cc_754 N_A_161_21#_c_1021_n N_VGND_c_1729_n 0.101784f $X=7.05 $Y=0.18 $X2=0
+ $Y2=0
cc_755 N_A_161_21#_c_1024_n N_VGND_c_1729_n 0.0037242f $X=3.255 $Y=0.18 $X2=0
+ $Y2=0
cc_756 N_A_161_21#_c_1026_n N_VGND_c_1729_n 0.0222759f $X=1.205 $Y=0.39 $X2=0
+ $Y2=0
cc_757 N_A_161_21#_c_1028_n N_VGND_c_1729_n 0.0102885f $X=0.97 $Y=0.18 $X2=0
+ $Y2=0
cc_758 N_A_161_21#_c_1021_n N_A_1141_125#_c_1842_n 0.00665102f $X=7.05 $Y=0.18
+ $X2=0 $Y2=0
cc_759 N_A_161_21#_c_1021_n N_A_1141_125#_c_1843_n 0.0200857f $X=7.05 $Y=0.18
+ $X2=0 $Y2=0
cc_760 N_A_161_21#_M1020_g N_A_1141_125#_c_1843_n 0.0140871f $X=7.125 $Y=0.855
+ $X2=0 $Y2=0
cc_761 N_A_161_21#_M1020_g N_A_1248_151#_c_1865_n 0.0141204f $X=7.125 $Y=0.855
+ $X2=0 $Y2=0
cc_762 N_A_161_21#_c_1025_n N_A_1248_151#_c_1865_n 0.00302692f $X=7.285 $Y=1.36
+ $X2=0 $Y2=0
cc_763 N_A_161_21#_M1020_g N_A_1248_151#_c_1866_n 6.44814e-19 $X=7.125 $Y=0.855
+ $X2=0 $Y2=0
cc_764 N_A_161_21#_M1020_g N_A_1248_151#_c_1867_n 0.0043223f $X=7.125 $Y=0.855
+ $X2=0 $Y2=0
cc_765 N_A_1535_177#_c_1171_n N_A_1331_151#_c_1256_n 0.00311093f $X=8.97 $Y=2.9
+ $X2=0 $Y2=0
cc_766 N_A_1535_177#_c_1173_n N_A_1331_151#_c_1256_n 0.00429613f $X=9.235
+ $Y=2.365 $X2=0 $Y2=0
cc_767 N_A_1535_177#_c_1165_n N_A_1331_151#_c_1237_n 0.00464207f $X=9.14 $Y=1.05
+ $X2=0 $Y2=0
cc_768 N_A_1535_177#_c_1165_n N_A_1331_151#_c_1242_n 0.00480149f $X=9.14 $Y=1.05
+ $X2=0 $Y2=0
cc_769 N_A_1535_177#_c_1173_n N_A_1331_151#_c_1260_n 6.02103e-19 $X=9.235
+ $Y=2.365 $X2=0 $Y2=0
cc_770 N_A_1535_177#_c_1167_n N_A_1331_151#_c_1243_n 8.14515e-19 $X=8.21 $Y=1.05
+ $X2=0 $Y2=0
cc_771 N_A_1535_177#_M1030_g N_A_1331_151#_c_1244_n 0.0135528f $X=7.75 $Y=2.455
+ $X2=0 $Y2=0
cc_772 N_A_1535_177#_c_1165_n N_A_1331_151#_c_1244_n 0.0531833f $X=9.14 $Y=1.05
+ $X2=0 $Y2=0
cc_773 N_A_1535_177#_c_1167_n N_A_1331_151#_c_1244_n 0.00884672f $X=8.21 $Y=1.05
+ $X2=0 $Y2=0
cc_774 N_A_1535_177#_c_1173_n N_A_1331_151#_c_1245_n 0.00198433f $X=9.235
+ $Y=2.365 $X2=0 $Y2=0
cc_775 N_A_1535_177#_c_1165_n N_A_1331_151#_c_1246_n 0.043226f $X=9.14 $Y=1.05
+ $X2=0 $Y2=0
cc_776 N_A_1535_177#_c_1167_n N_A_1331_151#_c_1273_n 0.00117246f $X=8.21 $Y=1.05
+ $X2=0 $Y2=0
cc_777 N_A_1535_177#_c_1169_n N_A_1331_151#_c_1268_n 0.01078f $X=8.805 $Y=3.11
+ $X2=0 $Y2=0
cc_778 N_A_1535_177#_c_1171_n N_A_1331_151#_c_1268_n 0.00200454f $X=8.97 $Y=2.9
+ $X2=0 $Y2=0
cc_779 N_A_1535_177#_c_1173_n N_A_1331_151#_c_1268_n 0.026833f $X=9.235 $Y=2.365
+ $X2=0 $Y2=0
cc_780 N_A_1535_177#_c_1165_n N_A_1331_151#_c_1252_n 0.0135503f $X=9.14 $Y=1.05
+ $X2=0 $Y2=0
cc_781 N_A_1535_177#_c_1165_n N_A_1331_151#_c_1269_n 0.0147931f $X=9.14 $Y=1.05
+ $X2=0 $Y2=0
cc_782 N_A_1535_177#_c_1173_n N_A_1331_151#_c_1269_n 0.00717088f $X=9.235
+ $Y=2.365 $X2=0 $Y2=0
cc_783 N_A_1535_177#_c_1165_n N_A_2005_119#_c_1420_n 0.00492391f $X=9.14 $Y=1.05
+ $X2=0 $Y2=0
cc_784 N_A_1535_177#_M1030_g N_VPWR_c_1485_n 0.00455764f $X=7.75 $Y=2.455 $X2=0
+ $Y2=0
cc_785 N_A_1535_177#_c_1169_n N_VPWR_c_1485_n 0.0197287f $X=8.805 $Y=3.11 $X2=0
+ $Y2=0
cc_786 N_A_1535_177#_c_1171_n N_VPWR_c_1486_n 0.0201375f $X=8.97 $Y=2.9 $X2=0
+ $Y2=0
cc_787 N_A_1535_177#_c_1172_n N_VPWR_c_1486_n 0.00895302f $X=8.97 $Y=2.9 $X2=0
+ $Y2=0
cc_788 N_A_1535_177#_c_1170_n N_VPWR_c_1493_n 0.00625713f $X=7.825 $Y=3.11 $X2=0
+ $Y2=0
cc_789 N_A_1535_177#_c_1169_n N_VPWR_c_1494_n 0.0318598f $X=8.805 $Y=3.11 $X2=0
+ $Y2=0
cc_790 N_A_1535_177#_c_1171_n N_VPWR_c_1494_n 0.0159061f $X=8.97 $Y=2.9 $X2=0
+ $Y2=0
cc_791 N_A_1535_177#_c_1169_n N_VPWR_c_1479_n 0.0271328f $X=8.805 $Y=3.11 $X2=0
+ $Y2=0
cc_792 N_A_1535_177#_c_1170_n N_VPWR_c_1479_n 0.0105968f $X=7.825 $Y=3.11 $X2=0
+ $Y2=0
cc_793 N_A_1535_177#_c_1171_n N_VPWR_c_1479_n 0.0085619f $X=8.97 $Y=2.9 $X2=0
+ $Y2=0
cc_794 N_A_1535_177#_c_1172_n N_VPWR_c_1479_n 0.0118827f $X=8.97 $Y=2.9 $X2=0
+ $Y2=0
cc_795 N_A_1535_177#_c_1173_n N_VPWR_c_1479_n 0.0101942f $X=9.235 $Y=2.365 $X2=0
+ $Y2=0
cc_796 N_A_1535_177#_c_1164_n N_VGND_c_1716_n 0.00187458f $X=8.21 $Y=0.885 $X2=0
+ $Y2=0
cc_797 N_A_1535_177#_c_1165_n N_VGND_c_1716_n 0.0201114f $X=9.14 $Y=1.05 $X2=0
+ $Y2=0
cc_798 N_A_1535_177#_c_1166_n N_VGND_c_1716_n 0.00687192f $X=9.305 $Y=0.805
+ $X2=0 $Y2=0
cc_799 N_A_1535_177#_c_1164_n N_VGND_c_1723_n 0.00473823f $X=8.21 $Y=0.885 $X2=0
+ $Y2=0
cc_800 N_A_1535_177#_c_1166_n N_VGND_c_1726_n 0.00509161f $X=9.305 $Y=0.805
+ $X2=0 $Y2=0
cc_801 N_A_1535_177#_c_1164_n N_VGND_c_1729_n 0.00954057f $X=8.21 $Y=0.885 $X2=0
+ $Y2=0
cc_802 N_A_1535_177#_c_1166_n N_VGND_c_1729_n 0.00873769f $X=9.305 $Y=0.805
+ $X2=0 $Y2=0
cc_803 N_A_1535_177#_c_1167_n N_VGND_c_1729_n 8.17771e-19 $X=8.21 $Y=1.05 $X2=0
+ $Y2=0
cc_804 N_A_1535_177#_c_1164_n N_A_1141_125#_c_1843_n 0.00357125f $X=8.21
+ $Y=0.885 $X2=0 $Y2=0
cc_805 N_A_1535_177#_c_1165_n N_A_1248_151#_c_1865_n 0.00180257f $X=9.14 $Y=1.05
+ $X2=0 $Y2=0
cc_806 N_A_1535_177#_c_1167_n N_A_1248_151#_c_1865_n 0.00496391f $X=8.21 $Y=1.05
+ $X2=0 $Y2=0
cc_807 N_A_1535_177#_c_1164_n N_A_1248_151#_c_1867_n 6.90734e-19 $X=8.21
+ $Y=0.885 $X2=0 $Y2=0
cc_808 N_A_1535_177#_c_1165_n N_A_1248_151#_c_1867_n 0.0207543f $X=9.14 $Y=1.05
+ $X2=0 $Y2=0
cc_809 N_A_1535_177#_c_1167_n N_A_1248_151#_c_1867_n 0.00667172f $X=8.21 $Y=1.05
+ $X2=0 $Y2=0
cc_810 N_A_1331_151#_c_1247_n N_A_2005_119#_c_1416_n 0.00115459f $X=10.7 $Y=1.41
+ $X2=0 $Y2=0
cc_811 N_A_1331_151#_c_1248_n N_A_2005_119#_c_1416_n 0.00712657f $X=10.785
+ $Y=2.395 $X2=0 $Y2=0
cc_812 N_A_1331_151#_M1004_g N_A_2005_119#_M1014_g 0.0505406f $X=11.82 $Y=2.465
+ $X2=0 $Y2=0
cc_813 N_A_1331_151#_c_1248_n N_A_2005_119#_M1014_g 0.00494553f $X=10.785
+ $Y=2.395 $X2=0 $Y2=0
cc_814 N_A_1331_151#_c_1263_n N_A_2005_119#_M1014_g 0.0150919f $X=11.58 $Y=2.48
+ $X2=0 $Y2=0
cc_815 N_A_1331_151#_c_1249_n N_A_2005_119#_M1014_g 0.00738386f $X=11.665
+ $Y=2.395 $X2=0 $Y2=0
cc_816 N_A_1331_151#_c_1241_n N_A_2005_119#_M1022_g 0.0152118f $X=12.005 $Y=1.23
+ $X2=0 $Y2=0
cc_817 N_A_1331_151#_c_1247_n N_A_2005_119#_M1022_g 3.9712e-19 $X=10.7 $Y=1.41
+ $X2=0 $Y2=0
cc_818 N_A_1331_151#_c_1254_n N_A_2005_119#_M1022_g 0.00212281f $X=11.87
+ $Y=1.395 $X2=0 $Y2=0
cc_819 N_A_1331_151#_c_1255_n N_A_2005_119#_M1022_g 0.0198581f $X=12.005
+ $Y=1.395 $X2=0 $Y2=0
cc_820 N_A_1331_151#_M1004_g N_A_2005_119#_c_1419_n 0.00387977f $X=11.82
+ $Y=2.465 $X2=0 $Y2=0
cc_821 N_A_1331_151#_c_1249_n N_A_2005_119#_c_1419_n 5.79366e-19 $X=11.665
+ $Y=2.395 $X2=0 $Y2=0
cc_822 N_A_1331_151#_c_1239_n N_A_2005_119#_c_1420_n 0.00281181f $X=9.95
+ $Y=1.125 $X2=0 $Y2=0
cc_823 N_A_1331_151#_c_1247_n N_A_2005_119#_c_1420_n 0.0546533f $X=10.7 $Y=1.41
+ $X2=0 $Y2=0
cc_824 N_A_1331_151#_c_1239_n N_A_2005_119#_c_1421_n 0.0111704f $X=9.95 $Y=1.125
+ $X2=0 $Y2=0
cc_825 N_A_1331_151#_c_1247_n N_A_2005_119#_c_1421_n 0.0153575f $X=10.7 $Y=1.41
+ $X2=0 $Y2=0
cc_826 N_A_1331_151#_c_1258_n N_A_2005_119#_c_1424_n 0.00673128f $X=9.995
+ $Y=2.045 $X2=0 $Y2=0
cc_827 N_A_1331_151#_c_1248_n N_A_2005_119#_c_1424_n 0.0111747f $X=10.785
+ $Y=2.395 $X2=0 $Y2=0
cc_828 N_A_1331_151#_c_1264_n N_A_2005_119#_c_1424_n 0.00883952f $X=10.87
+ $Y=2.48 $X2=0 $Y2=0
cc_829 N_A_1331_151#_c_1256_n N_A_2005_119#_c_1425_n 4.89574e-19 $X=9.45
+ $Y=2.045 $X2=0 $Y2=0
cc_830 N_A_1331_151#_c_1257_n N_A_2005_119#_c_1425_n 0.00444596f $X=9.92 $Y=1.97
+ $X2=0 $Y2=0
cc_831 N_A_1331_151#_c_1258_n N_A_2005_119#_c_1425_n 0.00461799f $X=9.995
+ $Y=2.045 $X2=0 $Y2=0
cc_832 N_A_1331_151#_c_1247_n N_A_2005_119#_c_1425_n 0.00815092f $X=10.7 $Y=1.41
+ $X2=0 $Y2=0
cc_833 N_A_1331_151#_c_1248_n N_A_2005_119#_c_1425_n 0.0137387f $X=10.785
+ $Y=2.395 $X2=0 $Y2=0
cc_834 N_A_1331_151#_c_1257_n N_A_2005_119#_c_1426_n 6.9482e-19 $X=9.92 $Y=1.97
+ $X2=0 $Y2=0
cc_835 N_A_1331_151#_c_1247_n N_A_2005_119#_c_1426_n 0.0182045f $X=10.7 $Y=1.41
+ $X2=0 $Y2=0
cc_836 N_A_1331_151#_c_1248_n N_A_2005_119#_c_1426_n 0.0235475f $X=10.785
+ $Y=2.395 $X2=0 $Y2=0
cc_837 N_A_1331_151#_c_1253_n N_A_2005_119#_c_1426_n 7.40229e-19 $X=9.43 $Y=1.48
+ $X2=0 $Y2=0
cc_838 N_A_1331_151#_c_1257_n N_A_2005_119#_c_1422_n 0.00690777f $X=9.92 $Y=1.97
+ $X2=0 $Y2=0
cc_839 N_A_1331_151#_c_1247_n N_A_2005_119#_c_1422_n 0.0103854f $X=10.7 $Y=1.41
+ $X2=0 $Y2=0
cc_840 N_A_1331_151#_c_1248_n N_A_2005_119#_c_1422_n 0.0116719f $X=10.785
+ $Y=2.395 $X2=0 $Y2=0
cc_841 N_A_1331_151#_c_1269_n N_A_2005_119#_c_1422_n 0.00222409f $X=9.43 $Y=1.48
+ $X2=0 $Y2=0
cc_842 N_A_1331_151#_c_1253_n N_A_2005_119#_c_1422_n 0.00205889f $X=9.43 $Y=1.48
+ $X2=0 $Y2=0
cc_843 N_A_1331_151#_c_1263_n N_VPWR_M1014_d 0.00392858f $X=11.58 $Y=2.48 $X2=0
+ $Y2=0
cc_844 N_A_1331_151#_c_1249_n N_VPWR_M1014_d 0.00510945f $X=11.665 $Y=2.395
+ $X2=0 $Y2=0
cc_845 N_A_1331_151#_c_1256_n N_VPWR_c_1486_n 0.00206293f $X=9.45 $Y=2.045 $X2=0
+ $Y2=0
cc_846 N_A_1331_151#_c_1257_n N_VPWR_c_1486_n 0.00623931f $X=9.92 $Y=1.97 $X2=0
+ $Y2=0
cc_847 N_A_1331_151#_c_1258_n N_VPWR_c_1486_n 0.00724f $X=9.995 $Y=2.045 $X2=0
+ $Y2=0
cc_848 N_A_1331_151#_c_1247_n N_VPWR_c_1486_n 0.00847365f $X=10.7 $Y=1.41 $X2=0
+ $Y2=0
cc_849 N_A_1331_151#_c_1269_n N_VPWR_c_1486_n 0.00151226f $X=9.43 $Y=1.48 $X2=0
+ $Y2=0
cc_850 N_A_1331_151#_M1004_g N_VPWR_c_1487_n 0.0099987f $X=11.82 $Y=2.465 $X2=0
+ $Y2=0
cc_851 N_A_1331_151#_c_1263_n N_VPWR_c_1487_n 0.0159924f $X=11.58 $Y=2.48 $X2=0
+ $Y2=0
cc_852 N_A_1331_151#_c_1258_n N_VPWR_c_1488_n 0.00455206f $X=9.995 $Y=2.045
+ $X2=0 $Y2=0
cc_853 N_A_1331_151#_c_1256_n N_VPWR_c_1494_n 0.00352953f $X=9.45 $Y=2.045 $X2=0
+ $Y2=0
cc_854 N_A_1331_151#_M1004_g N_VPWR_c_1495_n 0.00486043f $X=11.82 $Y=2.465 $X2=0
+ $Y2=0
cc_855 N_A_1331_151#_M1007_d N_VPWR_c_1479_n 0.00213122f $X=6.835 $Y=2.245 $X2=0
+ $Y2=0
cc_856 N_A_1331_151#_c_1256_n N_VPWR_c_1479_n 0.00434946f $X=9.45 $Y=2.045 $X2=0
+ $Y2=0
cc_857 N_A_1331_151#_c_1258_n N_VPWR_c_1479_n 0.00495025f $X=9.995 $Y=2.045
+ $X2=0 $Y2=0
cc_858 N_A_1331_151#_M1004_g N_VPWR_c_1479_n 0.00931409f $X=11.82 $Y=2.465 $X2=0
+ $Y2=0
cc_859 N_A_1331_151#_c_1263_n N_VPWR_c_1479_n 0.0213307f $X=11.58 $Y=2.48 $X2=0
+ $Y2=0
cc_860 N_A_1331_151#_c_1264_n N_VPWR_c_1479_n 0.0071207f $X=10.87 $Y=2.48 $X2=0
+ $Y2=0
cc_861 N_A_1331_151#_c_1268_n N_VPWR_c_1479_n 0.0145241f $X=8.62 $Y=2.39 $X2=0
+ $Y2=0
cc_862 N_A_1331_151#_c_1263_n N_Q_M1014_s 0.00691167f $X=11.58 $Y=2.48 $X2=0
+ $Y2=0
cc_863 N_A_1331_151#_M1004_g Q 5.91204e-19 $X=11.82 $Y=2.465 $X2=0 $Y2=0
cc_864 N_A_1331_151#_c_1241_n Q 7.84735e-19 $X=12.005 $Y=1.23 $X2=0 $Y2=0
cc_865 N_A_1331_151#_c_1247_n Q 0.0150744f $X=10.7 $Y=1.41 $X2=0 $Y2=0
cc_866 N_A_1331_151#_c_1248_n Q 0.0572625f $X=10.785 $Y=2.395 $X2=0 $Y2=0
cc_867 N_A_1331_151#_c_1263_n Q 0.0248011f $X=11.58 $Y=2.48 $X2=0 $Y2=0
cc_868 N_A_1331_151#_c_1249_n Q 0.0498653f $X=11.665 $Y=2.395 $X2=0 $Y2=0
cc_869 N_A_1331_151#_c_1254_n Q 0.0265291f $X=11.87 $Y=1.395 $X2=0 $Y2=0
cc_870 N_A_1331_151#_c_1255_n Q 2.80053e-19 $X=12.005 $Y=1.395 $X2=0 $Y2=0
cc_871 N_A_1331_151#_M1004_g Q_N 0.00511517f $X=11.82 $Y=2.465 $X2=0 $Y2=0
cc_872 N_A_1331_151#_c_1249_n Q_N 0.0240704f $X=11.665 $Y=2.395 $X2=0 $Y2=0
cc_873 N_A_1331_151#_c_1254_n Q_N 0.00113093f $X=11.87 $Y=1.395 $X2=0 $Y2=0
cc_874 N_A_1331_151#_c_1255_n Q_N 0.00636238f $X=12.005 $Y=1.395 $X2=0 $Y2=0
cc_875 N_A_1331_151#_M1004_g N_Q_N_c_1693_n 0.00362638f $X=11.82 $Y=2.465 $X2=0
+ $Y2=0
cc_876 N_A_1331_151#_c_1241_n N_Q_N_c_1693_n 0.0170324f $X=12.005 $Y=1.23 $X2=0
+ $Y2=0
cc_877 N_A_1331_151#_c_1249_n N_Q_N_c_1693_n 0.00738648f $X=11.665 $Y=2.395
+ $X2=0 $Y2=0
cc_878 N_A_1331_151#_c_1254_n N_Q_N_c_1693_n 0.025914f $X=11.87 $Y=1.395 $X2=0
+ $Y2=0
cc_879 N_A_1331_151#_c_1237_n N_VGND_c_1716_n 0.00269764f $X=9.52 $Y=1.125 $X2=0
+ $Y2=0
cc_880 N_A_1331_151#_c_1237_n N_VGND_c_1717_n 0.00201661f $X=9.52 $Y=1.125 $X2=0
+ $Y2=0
cc_881 N_A_1331_151#_c_1238_n N_VGND_c_1717_n 0.00232793f $X=9.875 $Y=1.2 $X2=0
+ $Y2=0
cc_882 N_A_1331_151#_c_1239_n N_VGND_c_1717_n 0.00360949f $X=9.95 $Y=1.125 $X2=0
+ $Y2=0
cc_883 N_A_1331_151#_c_1247_n N_VGND_c_1717_n 0.0101489f $X=10.7 $Y=1.41 $X2=0
+ $Y2=0
cc_884 N_A_1331_151#_c_1241_n N_VGND_c_1718_n 0.00397264f $X=12.005 $Y=1.23
+ $X2=0 $Y2=0
cc_885 N_A_1331_151#_c_1254_n N_VGND_c_1718_n 0.0259804f $X=11.87 $Y=1.395 $X2=0
+ $Y2=0
cc_886 N_A_1331_151#_c_1255_n N_VGND_c_1718_n 0.00523425f $X=12.005 $Y=1.395
+ $X2=0 $Y2=0
cc_887 N_A_1331_151#_c_1237_n N_VGND_c_1726_n 0.00431487f $X=9.52 $Y=1.125 $X2=0
+ $Y2=0
cc_888 N_A_1331_151#_c_1239_n N_VGND_c_1727_n 0.00431487f $X=9.95 $Y=1.125 $X2=0
+ $Y2=0
cc_889 N_A_1331_151#_c_1241_n N_VGND_c_1728_n 0.00540763f $X=12.005 $Y=1.23
+ $X2=0 $Y2=0
cc_890 N_A_1331_151#_c_1237_n N_VGND_c_1729_n 0.00477801f $X=9.52 $Y=1.125 $X2=0
+ $Y2=0
cc_891 N_A_1331_151#_c_1239_n N_VGND_c_1729_n 0.00477801f $X=9.95 $Y=1.125 $X2=0
+ $Y2=0
cc_892 N_A_1331_151#_c_1241_n N_VGND_c_1729_n 0.0112074f $X=12.005 $Y=1.23 $X2=0
+ $Y2=0
cc_893 N_A_1331_151#_M1019_d N_A_1248_151#_c_1865_n 0.00520986f $X=6.655
+ $Y=0.755 $X2=0 $Y2=0
cc_894 N_A_1331_151#_c_1244_n N_A_1248_151#_c_1865_n 0.0197002f $X=8.535 $Y=1.4
+ $X2=0 $Y2=0
cc_895 N_A_1331_151#_c_1273_n N_A_1248_151#_c_1865_n 0.0244929f $X=7.02 $Y=1.06
+ $X2=0 $Y2=0
cc_896 N_A_1331_151#_c_1251_n N_A_1248_151#_c_1865_n 0.00104774f $X=7.037 $Y=1.4
+ $X2=0 $Y2=0
cc_897 N_A_2005_119#_c_1424_n N_VPWR_c_1486_n 0.0242198f $X=10.21 $Y=2.3 $X2=0
+ $Y2=0
cc_898 N_A_2005_119#_M1014_g N_VPWR_c_1487_n 0.0204595f $X=11.39 $Y=2.465 $X2=0
+ $Y2=0
cc_899 N_A_2005_119#_M1014_g N_VPWR_c_1488_n 0.00486043f $X=11.39 $Y=2.465 $X2=0
+ $Y2=0
cc_900 N_A_2005_119#_c_1424_n N_VPWR_c_1488_n 0.00728674f $X=10.21 $Y=2.3 $X2=0
+ $Y2=0
cc_901 N_A_2005_119#_M1014_g N_VPWR_c_1479_n 0.00586151f $X=11.39 $Y=2.465 $X2=0
+ $Y2=0
cc_902 N_A_2005_119#_c_1424_n N_VPWR_c_1479_n 0.00926863f $X=10.21 $Y=2.3 $X2=0
+ $Y2=0
cc_903 N_A_2005_119#_c_1416_n Q 0.015422f $X=11.315 $Y=1.56 $X2=0 $Y2=0
cc_904 N_A_2005_119#_M1014_g Q 0.0138594f $X=11.39 $Y=2.465 $X2=0 $Y2=0
cc_905 N_A_2005_119#_M1022_g Q 0.0218573f $X=11.42 $Y=0.7 $X2=0 $Y2=0
cc_906 N_A_2005_119#_c_1419_n Q 0.00233759f $X=11.405 $Y=1.56 $X2=0 $Y2=0
cc_907 N_A_2005_119#_c_1420_n Q 0.0289856f $X=10.565 $Y=1.07 $X2=0 $Y2=0
cc_908 N_A_2005_119#_c_1421_n Q 0.0057342f $X=10.565 $Y=1.07 $X2=0 $Y2=0
cc_909 N_A_2005_119#_M1022_g N_VGND_c_1718_n 0.0135792f $X=11.42 $Y=0.7 $X2=0
+ $Y2=0
cc_910 N_A_2005_119#_M1022_g N_VGND_c_1727_n 0.00465848f $X=11.42 $Y=0.7 $X2=0
+ $Y2=0
cc_911 N_A_2005_119#_c_1420_n N_VGND_c_1727_n 0.0129444f $X=10.565 $Y=1.07 $X2=0
+ $Y2=0
cc_912 N_A_2005_119#_M1022_g N_VGND_c_1729_n 0.00938259f $X=11.42 $Y=0.7 $X2=0
+ $Y2=0
cc_913 N_A_2005_119#_c_1420_n N_VGND_c_1729_n 0.0207252f $X=10.565 $Y=1.07 $X2=0
+ $Y2=0
cc_914 N_VPWR_c_1479_n N_A_494_119#_M1018_d 0.00226211f $X=12.24 $Y=3.33 $X2=0
+ $Y2=0
cc_915 N_VPWR_c_1482_n N_A_494_119#_c_1628_n 0.00186388f $X=2.165 $Y=2.84 $X2=0
+ $Y2=0
cc_916 N_VPWR_c_1482_n N_A_494_119#_c_1644_n 0.0210129f $X=2.165 $Y=2.84 $X2=0
+ $Y2=0
cc_917 N_VPWR_c_1491_n N_A_494_119#_c_1644_n 0.0162502f $X=3.77 $Y=3.33 $X2=0
+ $Y2=0
cc_918 N_VPWR_c_1479_n N_A_494_119#_c_1644_n 0.0124941f $X=12.24 $Y=3.33 $X2=0
+ $Y2=0
cc_919 N_VPWR_c_1479_n A_687_533# 0.00256433f $X=12.24 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_920 N_VPWR_c_1479_n A_1259_449# 0.00336853f $X=12.24 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_921 N_VPWR_c_1479_n N_Q_M1014_s 0.00361946f $X=12.24 $Y=3.33 $X2=0 $Y2=0
cc_922 N_VPWR_c_1479_n N_Q_N_M1004_d 0.00371702f $X=12.24 $Y=3.33 $X2=0 $Y2=0
cc_923 N_VPWR_c_1495_n N_Q_N_c_1696_n 0.03179f $X=12.24 $Y=3.33 $X2=0 $Y2=0
cc_924 N_VPWR_c_1479_n N_Q_N_c_1696_n 0.0176116f $X=12.24 $Y=3.33 $X2=0 $Y2=0
cc_925 Q N_VGND_c_1718_n 0.0461897f $X=11.195 $Y=0.47 $X2=0 $Y2=0
cc_926 Q N_VGND_c_1727_n 0.00981119f $X=11.195 $Y=0.47 $X2=0 $Y2=0
cc_927 Q N_VGND_c_1729_n 0.0122366f $X=11.195 $Y=0.47 $X2=0 $Y2=0
cc_928 N_Q_N_c_1693_n N_VGND_c_1718_n 0.00132054f $X=12.22 $Y=0.425 $X2=0 $Y2=0
cc_929 N_Q_N_c_1693_n N_VGND_c_1728_n 0.0186238f $X=12.22 $Y=0.425 $X2=0 $Y2=0
cc_930 N_Q_N_c_1693_n N_VGND_c_1729_n 0.0103947f $X=12.22 $Y=0.425 $X2=0 $Y2=0
cc_931 N_VGND_c_1729_n N_A_1141_125#_M1020_d 0.00248311f $X=12.24 $Y=0 $X2=0
+ $Y2=0
cc_932 N_VGND_c_1715_n N_A_1141_125#_c_1841_n 0.012028f $X=5.415 $Y=0.91 $X2=0
+ $Y2=0
cc_933 N_VGND_c_1715_n N_A_1141_125#_c_1842_n 0.013094f $X=5.415 $Y=0.91 $X2=0
+ $Y2=0
cc_934 N_VGND_c_1723_n N_A_1141_125#_c_1842_n 0.018197f $X=8.62 $Y=0 $X2=0 $Y2=0
cc_935 N_VGND_c_1729_n N_A_1141_125#_c_1842_n 0.00937024f $X=12.24 $Y=0 $X2=0
+ $Y2=0
cc_936 N_VGND_c_1723_n N_A_1141_125#_c_1843_n 0.0972221f $X=8.62 $Y=0 $X2=0
+ $Y2=0
cc_937 N_VGND_c_1729_n N_A_1141_125#_c_1843_n 0.0553776f $X=12.24 $Y=0 $X2=0
+ $Y2=0
cc_938 N_VGND_c_1723_n N_A_1248_151#_c_1865_n 0.00399754f $X=8.62 $Y=0 $X2=0
+ $Y2=0
cc_939 N_VGND_c_1729_n N_A_1248_151#_c_1865_n 0.0082531f $X=12.24 $Y=0 $X2=0
+ $Y2=0
cc_940 N_VGND_c_1723_n N_A_1248_151#_c_1867_n 0.00900326f $X=8.62 $Y=0 $X2=0
+ $Y2=0
cc_941 N_VGND_c_1729_n N_A_1248_151#_c_1867_n 0.00940099f $X=12.24 $Y=0 $X2=0
+ $Y2=0
cc_942 N_A_1141_125#_M1020_d N_A_1248_151#_c_1865_n 0.0116276f $X=7.2 $Y=0.535
+ $X2=0 $Y2=0
cc_943 N_A_1141_125#_c_1843_n N_A_1248_151#_c_1865_n 0.0719352f $X=7.455 $Y=0.35
+ $X2=0 $Y2=0
cc_944 N_A_1141_125#_c_1841_n N_A_1248_151#_c_1866_n 0.0348912f $X=5.845 $Y=0.91
+ $X2=0 $Y2=0
cc_945 N_A_1141_125#_c_1843_n N_A_1248_151#_c_1866_n 0.0253546f $X=7.455 $Y=0.35
+ $X2=0 $Y2=0
cc_946 N_A_1141_125#_c_1843_n N_A_1248_151#_c_1867_n 0.00330631f $X=7.455
+ $Y=0.35 $X2=0 $Y2=0
