* File: sky130_fd_sc_lp__o2bb2ai_lp.spice
* Created: Wed Sep  2 10:22:31 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__o2bb2ai_lp.pex.spice"
.subckt sky130_fd_sc_lp__o2bb2ai_lp  VNB VPB A1_N A2_N B2 B1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B1	B1
* B2	B2
* A2_N	A2_N
* A1_N	A1_N
* VPB	VPB
* VNB	VNB
MM1001 A_114_57# N_A1_N_M1001_g N_VGND_M1001_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.1197 PD=0.66 PS=1.41 NRD=18.564 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1009 N_A_145_419#_M1009_d N_A2_N_M1009_g A_114_57# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0504 PD=1.41 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1007 N_A_400_83#_M1007_d N_A_145_419#_M1007_g N_Y_M1007_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0588 AS=0.1197 PD=0.7 PS=1.41 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1003 N_VGND_M1003_d N_B2_M1003_g N_A_400_83#_M1007_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0651 AS=0.0588 PD=0.73 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1000 N_A_400_83#_M1000_d N_B1_M1000_g N_VGND_M1003_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.0651 PD=1.37 PS=0.73 NRD=0 NRS=8.568 M=1 R=2.8 SA=75001.1
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1006 N_A_145_419#_M1006_d N_A1_N_M1006_g N_VPWR_M1006_s VPB PHIGHVT L=0.25 W=1
+ AD=0.14 AS=0.295 PD=1.28 PS=2.59 NRD=0 NRS=1.9503 M=1 R=4 SA=125000 SB=125002
+ A=0.25 P=2.5 MULT=1
MM1005 N_VPWR_M1005_d N_A2_N_M1005_g N_A_145_419#_M1006_d VPB PHIGHVT L=0.25 W=1
+ AD=0.2075 AS=0.14 PD=1.415 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125001 SB=125002
+ A=0.25 P=2.5 MULT=1
MM1002 N_Y_M1002_d N_A_145_419#_M1002_g N_VPWR_M1005_d VPB PHIGHVT L=0.25 W=1
+ AD=0.14 AS=0.2075 PD=1.28 PS=1.415 NRD=0 NRS=26.5753 M=1 R=4 SA=125001
+ SB=125001 A=0.25 P=2.5 MULT=1
MM1008 A_490_419# N_B2_M1008_g N_Y_M1002_d VPB PHIGHVT L=0.25 W=1 AD=0.12
+ AS=0.14 PD=1.24 PS=1.28 NRD=12.7853 NRS=0 M=1 R=4 SA=125002 SB=125001 A=0.25
+ P=2.5 MULT=1
MM1004 N_VPWR_M1004_d N_B1_M1004_g A_490_419# VPB PHIGHVT L=0.25 W=1 AD=0.265
+ AS=0.12 PD=2.53 PS=1.24 NRD=0 NRS=12.7853 M=1 R=4 SA=125002 SB=125000 A=0.25
+ P=2.5 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9751 P=11.21
c_37 VNB 0 1.34366e-19 $X=0 $Y=0
*
.include "sky130_fd_sc_lp__o2bb2ai_lp.pxi.spice"
*
.ends
*
*
