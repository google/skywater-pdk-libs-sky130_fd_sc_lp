* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__srsdfrtn_1 CLK_N D RESET_B SCD SCE SLEEP_B KAPWR VGND VNB
+ VPB VPWR Q
X0 VPWR SCE a_247_491# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X1 a_411_491# SCD VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X2 a_1373_77# a_1343_51# a_1453_77# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 VPWR a_3368_57# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X4 KAPWR CLK_N a_742_63# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X5 a_2562_427# a_742_63# a_2645_427# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X6 a_2562_427# a_2999_73# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X7 VGND SLEEP_B a_2480_97# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 a_247_491# D a_305_97# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X9 a_2198_97# SLEEP_B a_2276_97# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 a_3115_99# a_2717_427# a_2999_73# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X11 VGND a_3368_57# Q VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X12 a_1682_341# a_1724_21# KAPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X13 a_2717_427# a_666_89# a_1343_51# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X14 a_391_97# a_27_55# a_469_97# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X15 a_2717_427# a_666_89# a_2879_99# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X16 VGND RESET_B a_469_97# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X17 a_469_97# SCD a_220_97# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X18 a_2999_73# a_2717_427# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X19 a_666_89# a_742_63# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X20 a_220_97# SCE a_305_97# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X21 a_742_63# SLEEP_B KAPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X22 VPWR RESET_B a_2999_73# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X23 a_305_97# a_27_55# a_411_491# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X24 a_305_97# a_742_63# a_1041_419# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X25 a_305_97# D a_391_97# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X26 a_666_89# a_742_63# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X27 a_3368_57# a_2717_427# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X28 KAPWR a_1113_419# a_1343_51# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X29 a_27_55# SCE VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X30 a_742_63# CLK_N a_2198_97# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X31 VGND RESET_B a_1453_77# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X32 VGND RESET_B a_3115_99# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X33 a_3368_57# a_2717_427# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X34 a_1453_77# a_1724_21# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X35 a_1242_419# a_1343_51# KAPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X36 a_2645_427# a_742_63# a_2717_427# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X37 VGND a_1113_419# a_1840_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X38 a_1009_107# a_742_63# a_1113_419# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X39 a_1113_419# RESET_B a_1682_341# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X40 a_1343_51# a_742_63# a_2717_427# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X41 a_2879_99# a_666_89# a_2951_99# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X42 a_1840_47# a_1113_419# a_1343_51# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X43 VPWR RESET_B a_305_97# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X44 a_1201_215# a_666_89# a_305_97# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X45 a_2276_97# SLEEP_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X46 a_27_55# SCE VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X47 a_1113_419# a_666_89# a_1242_419# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X48 a_1041_419# a_742_63# a_1113_419# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X49 a_1113_419# a_666_89# a_1201_215# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X50 a_2480_97# SLEEP_B a_1724_21# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X51 KAPWR SLEEP_B a_1724_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X52 a_2951_99# a_2999_73# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X53 a_1009_107# a_1343_51# a_1373_77# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
