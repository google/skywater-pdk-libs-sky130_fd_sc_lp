* File: sky130_fd_sc_lp__and4_m.pex.spice
* Created: Wed Sep  2 09:33:19 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__AND4_M%A 1 5 9 14 16 18 19 20 25
c33 18 0 8.08206e-20 $X=0.24 $Y=0.925
c34 14 0 2.96048e-20 $X=0.605 $Y=1.03
r35 25 26 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.27
+ $Y=1.12 $X2=0.27 $Y2=1.12
r36 19 20 20.5182 $w=1.98e-07 $l=3.7e-07 $layer=LI1_cond $X=0.255 $Y=1.295
+ $X2=0.255 $Y2=1.665
r37 19 26 9.70455 $w=1.98e-07 $l=1.75e-07 $layer=LI1_cond $X=0.255 $Y=1.295
+ $X2=0.255 $Y2=1.12
r38 18 26 10.8136 $w=1.98e-07 $l=1.95e-07 $layer=LI1_cond $X=0.255 $Y=0.925
+ $X2=0.255 $Y2=1.12
r39 16 25 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.27 $Y=1.46
+ $X2=0.27 $Y2=1.12
r40 16 17 46.7501 $w=3.3e-07 $l=2.97405e-07 $layer=POLY_cond $X=0.27 $Y=1.46
+ $X2=0.285 $Y2=1.75
r41 12 25 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=0.27 $Y=1.105
+ $X2=0.27 $Y2=1.12
r42 12 14 171.777 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=0.27 $Y=1.03
+ $X2=0.605 $Y2=1.03
r43 7 9 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=0.685 $Y=1.825
+ $X2=0.685 $Y2=2.165
r44 3 14 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.605 $Y=0.955
+ $X2=0.605 $Y2=1.03
r45 3 5 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=0.605 $Y=0.955
+ $X2=0.605 $Y2=0.445
r46 2 17 12.8954 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=0.435 $Y=1.75
+ $X2=0.285 $Y2=1.75
r47 1 7 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.61 $Y=1.75
+ $X2=0.685 $Y2=1.825
r48 1 2 89.734 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=0.61 $Y=1.75 $X2=0.435
+ $Y2=1.75
.ends

.subckt PM_SKY130_FD_SC_LP__AND4_M%B 3 6 9 10 11 12 13 14 19
c40 11 0 1.88521e-19 $X=1.055 $Y=1.435
c41 6 0 8.08206e-20 $X=1.115 $Y=2.165
r42 19 20 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.055
+ $Y=0.93 $X2=1.055 $Y2=0.93
r43 14 20 13.3537 $w=3.13e-07 $l=3.65e-07 $layer=LI1_cond $X=1.127 $Y=1.295
+ $X2=1.127 $Y2=0.93
r44 13 20 0.182927 $w=3.13e-07 $l=5e-09 $layer=LI1_cond $X=1.127 $Y=0.925
+ $X2=1.127 $Y2=0.93
r45 12 13 13.5366 $w=3.13e-07 $l=3.7e-07 $layer=LI1_cond $X=1.127 $Y=0.555
+ $X2=1.127 $Y2=0.925
r46 10 19 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.055 $Y=1.27
+ $X2=1.055 $Y2=0.93
r47 10 11 41.8716 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.055 $Y=1.27
+ $X2=1.055 $Y2=1.435
r48 9 19 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.055 $Y=0.765
+ $X2=1.055 $Y2=0.93
r49 6 11 374.319 $w=1.5e-07 $l=7.3e-07 $layer=POLY_cond $X=1.115 $Y=2.165
+ $X2=1.115 $Y2=1.435
r50 3 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.965 $Y=0.445
+ $X2=0.965 $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_LP__AND4_M%C 3 7 9 10 11 16
r38 16 19 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.595 $Y=1.32
+ $X2=1.595 $Y2=1.485
r39 16 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.595 $Y=1.32
+ $X2=1.595 $Y2=1.155
r40 11 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.595
+ $Y=1.32 $X2=1.595 $Y2=1.32
r41 10 11 16.7217 $w=2.53e-07 $l=3.7e-07 $layer=LI1_cond $X=1.637 $Y=0.925
+ $X2=1.637 $Y2=1.295
r42 9 10 16.7217 $w=2.53e-07 $l=3.7e-07 $layer=LI1_cond $X=1.637 $Y=0.555
+ $X2=1.637 $Y2=0.925
r43 7 19 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=1.545 $Y=2.165
+ $X2=1.545 $Y2=1.485
r44 3 18 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=1.505 $Y=0.445
+ $X2=1.505 $Y2=1.155
.ends

.subckt PM_SKY130_FD_SC_LP__AND4_M%D 1 3 6 13 15 16 17 18 19 24 26
c51 13 0 1.62226e-19 $X=2.045 $Y=0.84
r52 24 27 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.135 $Y=1.29
+ $X2=2.135 $Y2=1.455
r53 24 26 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.135 $Y=1.29
+ $X2=2.135 $Y2=1.125
r54 18 19 21.3287 $w=1.93e-07 $l=3.75e-07 $layer=LI1_cond $X=2.147 $Y=1.29
+ $X2=2.147 $Y2=1.665
r55 18 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.135
+ $Y=1.29 $X2=2.135 $Y2=1.29
r56 17 18 20.7599 $w=1.93e-07 $l=3.65e-07 $layer=LI1_cond $X=2.147 $Y=0.925
+ $X2=2.147 $Y2=1.29
r57 15 16 43.7534 $w=2.2e-07 $l=1.5e-07 $layer=POLY_cond $X=2.01 $Y=1.695
+ $X2=2.01 $Y2=1.845
r58 15 27 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=2.045 $Y=1.695
+ $X2=2.045 $Y2=1.455
r59 11 13 92.2979 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=1.865 $Y=0.84
+ $X2=2.045 $Y2=0.84
r60 7 13 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.045 $Y=0.915
+ $X2=2.045 $Y2=0.84
r61 7 26 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=2.045 $Y=0.915
+ $X2=2.045 $Y2=1.125
r62 6 16 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.975 $Y=2.165
+ $X2=1.975 $Y2=1.845
r63 1 11 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.865 $Y=0.765
+ $X2=1.865 $Y2=0.84
r64 1 3 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.865 $Y=0.765
+ $X2=1.865 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__AND4_M%A_53_47# 1 2 3 10 12 14 18 20 23 27 29 34 37
+ 39 40 43 46
c84 40 0 2.96048e-20 $X=1.005 $Y=1.8
c85 39 0 1.88521e-19 $X=1.655 $Y=1.8
r86 46 53 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=1.78 $Y=2.88 $X2=1.78
+ $Y2=2.97
r87 45 46 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.78
+ $Y=2.88 $X2=1.78 $Y2=2.88
r88 43 45 34.329 $w=2.08e-07 $l=6.5e-07 $layer=LI1_cond $X=1.76 $Y=2.23 $X2=1.76
+ $Y2=2.88
r89 41 43 18.2208 $w=2.08e-07 $l=3.45e-07 $layer=LI1_cond $X=1.76 $Y=1.885
+ $X2=1.76 $Y2=2.23
r90 39 41 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=1.655 $Y=1.8
+ $X2=1.76 $Y2=1.885
r91 39 40 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=1.655 $Y=1.8
+ $X2=1.005 $Y2=1.8
r92 35 40 7.04599 $w=1.68e-07 $l=1.08e-07 $layer=LI1_cond $X=0.897 $Y=1.8
+ $X2=1.005 $Y2=1.8
r93 35 48 12.5262 $w=1.68e-07 $l=1.92e-07 $layer=LI1_cond $X=0.897 $Y=1.8
+ $X2=0.705 $Y2=1.8
r94 35 37 11.5244 $w=2.13e-07 $l=2.15e-07 $layer=LI1_cond $X=0.897 $Y=1.885
+ $X2=0.897 $Y2=2.1
r95 34 48 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.705 $Y=1.715
+ $X2=0.705 $Y2=1.8
r96 33 34 68.8289 $w=1.68e-07 $l=1.055e-06 $layer=LI1_cond $X=0.705 $Y=0.66
+ $X2=0.705 $Y2=1.715
r97 29 33 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.62 $Y=0.495
+ $X2=0.705 $Y2=0.66
r98 29 31 8.03218 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=0.62 $Y=0.495
+ $X2=0.39 $Y2=0.495
r99 25 27 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=2.405 $Y=1.77
+ $X2=2.615 $Y2=1.77
r100 21 23 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=2.405 $Y=0.84
+ $X2=2.615 $Y2=0.84
r101 20 27 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.615 $Y=1.695
+ $X2=2.615 $Y2=1.77
r102 19 23 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.615 $Y=0.915
+ $X2=2.615 $Y2=0.84
r103 19 20 399.957 $w=1.5e-07 $l=7.8e-07 $layer=POLY_cond $X=2.615 $Y=0.915
+ $X2=2.615 $Y2=1.695
r104 16 18 374.319 $w=1.5e-07 $l=7.3e-07 $layer=POLY_cond $X=2.405 $Y=2.895
+ $X2=2.405 $Y2=2.165
r105 15 25 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.405 $Y=1.845
+ $X2=2.405 $Y2=1.77
r106 15 18 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.405 $Y=1.845
+ $X2=2.405 $Y2=2.165
r107 12 21 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.405 $Y=0.765
+ $X2=2.405 $Y2=0.84
r108 12 14 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.405 $Y=0.765
+ $X2=2.405 $Y2=0.445
r109 11 53 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.945 $Y=2.97
+ $X2=1.78 $Y2=2.97
r110 10 16 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.33 $Y=2.97
+ $X2=2.405 $Y2=2.895
r111 10 11 197.415 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=2.33 $Y=2.97
+ $X2=1.945 $Y2=2.97
r112 3 43 600 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=1 $X=1.62
+ $Y=1.955 $X2=1.76 $Y2=2.23
r113 2 37 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.76
+ $Y=1.955 $X2=0.9 $Y2=2.1
r114 1 31 182 $w=1.7e-07 $l=3.16386e-07 $layer=licon1_NDIFF $count=1 $X=0.265
+ $Y=0.235 $X2=0.39 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__AND4_M%VPWR 1 2 3 12 16 18 22 25 26 27 28 29 40 41
+ 44
r37 44 45 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r38 41 45 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r39 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r40 38 44 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=2.295 $Y=3.33
+ $X2=2.19 $Y2=3.33
r41 38 40 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=2.295 $Y=3.33
+ $X2=2.64 $Y2=3.33
r42 36 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r43 33 37 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.2 $Y2=3.33
r44 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r45 29 45 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=2.16 $Y2=3.33
r46 29 37 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=1.2 $Y2=3.33
r47 27 36 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=1.225 $Y=3.33
+ $X2=1.2 $Y2=3.33
r48 27 28 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.225 $Y=3.33
+ $X2=1.33 $Y2=3.33
r49 25 32 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=0.365 $Y=3.33
+ $X2=0.24 $Y2=3.33
r50 25 26 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=0.365 $Y=3.33
+ $X2=0.47 $Y2=3.33
r51 24 36 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=0.575 $Y=3.33
+ $X2=1.2 $Y2=3.33
r52 24 26 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=0.575 $Y=3.33
+ $X2=0.47 $Y2=3.33
r53 20 44 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=2.19 $Y=3.245
+ $X2=2.19 $Y2=3.33
r54 20 22 53.6061 $w=2.08e-07 $l=1.015e-06 $layer=LI1_cond $X=2.19 $Y=3.245
+ $X2=2.19 $Y2=2.23
r55 19 28 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.435 $Y=3.33
+ $X2=1.33 $Y2=3.33
r56 18 44 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=2.085 $Y=3.33
+ $X2=2.19 $Y2=3.33
r57 18 19 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=2.085 $Y=3.33
+ $X2=1.435 $Y2=3.33
r58 14 28 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=1.33 $Y=3.245
+ $X2=1.33 $Y2=3.33
r59 14 16 53.6061 $w=2.08e-07 $l=1.015e-06 $layer=LI1_cond $X=1.33 $Y=3.245
+ $X2=1.33 $Y2=2.23
r60 10 26 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=0.47 $Y=3.245
+ $X2=0.47 $Y2=3.33
r61 10 12 53.6061 $w=2.08e-07 $l=1.015e-06 $layer=LI1_cond $X=0.47 $Y=3.245
+ $X2=0.47 $Y2=2.23
r62 3 22 600 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=1 $X=2.05
+ $Y=1.955 $X2=2.19 $Y2=2.23
r63 2 16 600 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=1 $X=1.19
+ $Y=1.955 $X2=1.33 $Y2=2.23
r64 1 12 600 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_PDIFF $count=1 $X=0.345
+ $Y=1.955 $X2=0.47 $Y2=2.23
.ends

.subckt PM_SKY130_FD_SC_LP__AND4_M%X 1 2 7 8 9 10 11 12 13
r21 12 13 19.5411 $w=2.08e-07 $l=3.7e-07 $layer=LI1_cond $X=2.62 $Y=2.405
+ $X2=2.62 $Y2=2.775
r22 11 12 19.5411 $w=2.08e-07 $l=3.7e-07 $layer=LI1_cond $X=2.62 $Y=2.035
+ $X2=2.62 $Y2=2.405
r23 10 11 19.5411 $w=2.08e-07 $l=3.7e-07 $layer=LI1_cond $X=2.62 $Y=1.665
+ $X2=2.62 $Y2=2.035
r24 9 10 19.5411 $w=2.08e-07 $l=3.7e-07 $layer=LI1_cond $X=2.62 $Y=1.295
+ $X2=2.62 $Y2=1.665
r25 8 9 19.5411 $w=2.08e-07 $l=3.7e-07 $layer=LI1_cond $X=2.62 $Y=0.925 $X2=2.62
+ $Y2=1.295
r26 7 8 21.9177 $w=2.08e-07 $l=4.15e-07 $layer=LI1_cond $X=2.62 $Y=0.51 $X2=2.62
+ $Y2=0.925
r27 2 11 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.48
+ $Y=1.955 $X2=2.62 $Y2=2.1
r28 1 7 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=2.48
+ $Y=0.235 $X2=2.62 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_LP__AND4_M%VGND 1 6 8 10 20 21 24
c38 21 0 9.0026e-20 $X=2.64 $Y=0
c39 10 0 7.22003e-20 $X=1.945 $Y=0
r40 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r41 21 25 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=2.16
+ $Y2=0
r42 20 21 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r43 18 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.275 $Y=0 $X2=2.11
+ $Y2=0
r44 18 20 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=2.275 $Y=0 $X2=2.64
+ $Y2=0
r45 17 25 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r46 16 17 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r47 12 16 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=0.24 $Y=0 $X2=1.68
+ $Y2=0
r48 12 13 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r49 10 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.945 $Y=0 $X2=2.11
+ $Y2=0
r50 10 16 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=1.945 $Y=0 $X2=1.68
+ $Y2=0
r51 8 17 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=1.68
+ $Y2=0
r52 8 13 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=1.44 $Y=0 $X2=0.24
+ $Y2=0
r53 4 24 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.11 $Y=0.085 $X2=2.11
+ $Y2=0
r54 4 6 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.11 $Y=0.085
+ $X2=2.11 $Y2=0.38
r55 1 6 182 $w=1.7e-07 $l=2.31409e-07 $layer=licon1_NDIFF $count=1 $X=1.94
+ $Y=0.235 $X2=2.11 $Y2=0.38
.ends

