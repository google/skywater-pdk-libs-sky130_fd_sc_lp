* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__o311ai_0 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
M1000 VGND A2 a_193_48# VNB nshort w=420000u l=150000u
+  ad=2.541e+11p pd=2.89e+06u as=2.352e+11p ps=2.8e+06u
M1001 a_193_466# A1 VPWR VPB phighvt w=640000u l=150000u
+  ad=1.344e+11p pd=1.7e+06u as=4.128e+11p ps=3.85e+06u
M1002 a_265_466# A2 a_193_466# VPB phighvt w=640000u l=150000u
+  ad=1.344e+11p pd=1.7e+06u as=0p ps=0u
M1003 Y C1 VPWR VPB phighvt w=640000u l=150000u
+  ad=3.872e+11p pd=3.77e+06u as=0p ps=0u
M1004 Y A3 a_265_466# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_193_48# A1 VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_193_48# A3 VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR B1 Y VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 Y C1 a_463_48# VNB nshort w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=1.008e+11p ps=1.32e+06u
M1009 a_463_48# B1 a_193_48# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
