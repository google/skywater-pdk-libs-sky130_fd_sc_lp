* File: sky130_fd_sc_lp__a41o_lp.spice
* Created: Wed Sep  2 09:29:15 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__a41o_lp.pex.spice"
.subckt sky130_fd_sc_lp__a41o_lp  VNB VPB A4 A3 A2 A1 B1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* B1	B1
* A1	A1
* A2	A2
* A3	A3
* A4	A4
* VPB	VPB
* VNB	VNB
MM1010 A_128_47# N_A4_M1010_g N_VGND_M1010_s VNB NSHORT L=0.15 W=0.42 AD=0.0504
+ AS=0.1197 PD=0.66 PS=1.41 NRD=18.564 NRS=0 M=1 R=2.8 SA=75000.2 SB=75003.4
+ A=0.063 P=1.14 MULT=1
MM1005 A_206_47# N_A3_M1005_g A_128_47# VNB NSHORT L=0.15 W=0.42 AD=0.0819
+ AS=0.0504 PD=0.81 PS=0.66 NRD=39.996 NRS=18.564 M=1 R=2.8 SA=75000.6 SB=75003
+ A=0.063 P=1.14 MULT=1
MM1007 A_314_47# N_A2_M1007_g A_206_47# VNB NSHORT L=0.15 W=0.42 AD=0.0882
+ AS=0.0819 PD=0.84 PS=0.81 NRD=44.28 NRS=39.996 M=1 R=2.8 SA=75001.1 SB=75002.5
+ A=0.063 P=1.14 MULT=1
MM1000 N_A_428_47#_M1000_d N_A1_M1000_g A_314_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.0882 AS=0.0882 PD=0.84 PS=0.84 NRD=39.996 NRS=44.28 M=1 R=2.8 SA=75001.7
+ SB=75001.9 A=0.063 P=1.14 MULT=1
MM1008 A_542_47# N_B1_M1008_g N_A_428_47#_M1000_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0882 PD=0.63 PS=0.84 NRD=14.28 NRS=0 M=1 R=2.8 SA=75002.3
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1004 N_VGND_M1004_d N_B1_M1004_g A_542_47# VNB NSHORT L=0.15 W=0.42 AD=0.0588
+ AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75002.6 SB=75001 A=0.063
+ P=1.14 MULT=1
MM1009 A_700_47# N_A_428_47#_M1009_g N_VGND_M1004_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75003.1
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1011 N_X_M1011_d N_A_428_47#_M1011_g A_700_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75003.4
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1002 N_VPWR_M1002_d N_A4_M1002_g N_A_27_409#_M1002_s VPB PHIGHVT L=0.25 W=1
+ AD=0.14 AS=0.285 PD=1.28 PS=2.57 NRD=0 NRS=0 M=1 R=4 SA=125000 SB=125002
+ A=0.25 P=2.5 MULT=1
MM1006 N_A_27_409#_M1006_d N_A3_M1006_g N_VPWR_M1002_d VPB PHIGHVT L=0.25 W=1
+ AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125001 SB=125002 A=0.25
+ P=2.5 MULT=1
MM1001 N_VPWR_M1001_d N_A2_M1001_g N_A_27_409#_M1006_d VPB PHIGHVT L=0.25 W=1
+ AD=0.15 AS=0.14 PD=1.3 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125001 SB=125001 A=0.25
+ P=2.5 MULT=1
MM1012 N_A_27_409#_M1012_d N_A1_M1012_g N_VPWR_M1001_d VPB PHIGHVT L=0.25 W=1
+ AD=0.14 AS=0.15 PD=1.28 PS=1.3 NRD=0 NRS=3.9203 M=1 R=4 SA=125002 SB=125001
+ A=0.25 P=2.5 MULT=1
MM1003 N_A_428_47#_M1003_d N_B1_M1003_g N_A_27_409#_M1012_d VPB PHIGHVT L=0.25
+ W=1 AD=0.285 AS=0.14 PD=2.57 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125002 SB=125000
+ A=0.25 P=2.5 MULT=1
MM1013 N_X_M1013_d N_A_428_47#_M1013_g N_VPWR_M1013_s VPB PHIGHVT L=0.25 W=1
+ AD=0.285 AS=0.285 PD=2.57 PS=2.57 NRD=0 NRS=0 M=1 R=4 SA=125000 SB=125000
+ A=0.25 P=2.5 MULT=1
DX14_noxref VNB VPB NWDIODE A=8.7655 P=13.13
*
.include "sky130_fd_sc_lp__a41o_lp.pxi.spice"
*
.ends
*
*
