# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__o32a_m
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__o32a_m ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.840000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.635000 0.840000 1.120000 1.750000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.535000 1.185000 1.765000 2.490000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.075000 1.185000 2.245000 2.490000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.395000 0.840000 3.685000 1.750000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.535000 1.185000 2.865000 1.695000 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  0.222600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.155000 0.470000 0.395000 0.800000 ;
        RECT 0.155000 0.800000 0.325000 2.125000 ;
        RECT 0.155000 2.125000 0.395000 2.860000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 3.840000 0.085000 ;
        RECT 0.575000  0.085000 0.905000 0.655000 ;
        RECT 1.670000  0.085000 2.000000 0.655000 ;
      LAYER mcon ;
        RECT 0.155000 -0.085000 0.325000 0.085000 ;
        RECT 0.635000 -0.085000 0.805000 0.085000 ;
        RECT 1.115000 -0.085000 1.285000 0.085000 ;
        RECT 1.595000 -0.085000 1.765000 0.085000 ;
        RECT 2.075000 -0.085000 2.245000 0.085000 ;
        RECT 2.555000 -0.085000 2.725000 0.085000 ;
        RECT 3.035000 -0.085000 3.205000 0.085000 ;
        RECT 3.515000 -0.085000 3.685000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.840000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.245000 3.840000 3.415000 ;
        RECT 0.575000 2.185000 0.905000 3.245000 ;
        RECT 3.200000 2.225000 3.530000 3.245000 ;
      LAYER mcon ;
        RECT 0.155000 3.245000 0.325000 3.415000 ;
        RECT 0.635000 3.245000 0.805000 3.415000 ;
        RECT 1.115000 3.245000 1.285000 3.415000 ;
        RECT 1.595000 3.245000 1.765000 3.415000 ;
        RECT 2.075000 3.245000 2.245000 3.415000 ;
        RECT 2.555000 3.245000 2.725000 3.415000 ;
        RECT 3.035000 3.245000 3.205000 3.415000 ;
        RECT 3.515000 3.245000 3.685000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 3.840000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 1.300000 0.515000 1.490000 0.835000 ;
      RECT 1.300000 0.835000 2.550000 1.005000 ;
      RECT 2.110000 2.855000 2.635000 3.025000 ;
      RECT 2.360000 0.265000 3.570000 0.435000 ;
      RECT 2.360000 0.435000 2.550000 0.835000 ;
      RECT 2.425000 2.125000 2.635000 2.855000 ;
      RECT 2.465000 1.875000 3.215000 2.045000 ;
      RECT 2.465000 2.045000 2.635000 2.125000 ;
      RECT 2.730000 0.615000 3.060000 0.835000 ;
      RECT 2.730000 0.835000 3.215000 1.005000 ;
      RECT 3.045000 1.005000 3.215000 1.875000 ;
      RECT 3.240000 0.435000 3.570000 0.655000 ;
  END
END sky130_fd_sc_lp__o32a_m
