* File: sky130_fd_sc_lp__decap_12.pxi.spice
* Created: Wed Sep  2 09:41:46 2020
* 
x_PM_SKY130_FD_SC_LP__DECAP_12%VGND N_VGND_M1000_s N_VGND_c_28_n N_VGND_M1001_g
+ N_VGND_c_29_n N_VGND_c_30_n N_VGND_c_31_n N_VGND_c_32_n VGND N_VGND_c_33_n
+ N_VGND_c_34_n N_VGND_c_35_n N_VGND_c_36_n N_VGND_c_37_n
+ PM_SKY130_FD_SC_LP__DECAP_12%VGND
x_PM_SKY130_FD_SC_LP__DECAP_12%VPWR N_VPWR_M1001_s N_VPWR_c_61_n N_VPWR_c_57_n
+ N_VPWR_c_58_n N_VPWR_c_64_n VPWR N_VPWR_M1000_g N_VPWR_c_65_n N_VPWR_c_66_n
+ N_VPWR_c_67_n N_VPWR_c_60_n N_VPWR_c_69_n N_VPWR_c_70_n
+ PM_SKY130_FD_SC_LP__DECAP_12%VPWR
cc_1 VNB N_VGND_c_28_n 0.0434284f $X=-0.19 $Y=-0.245 $X2=2.58 $Y2=2.555
cc_2 VNB N_VGND_c_29_n 0.0651019f $X=-0.19 $Y=-0.245 $X2=0.815 $Y2=0.38
cc_3 VNB N_VGND_c_30_n 0.00211035f $X=-0.19 $Y=-0.245 $X2=0.98 $Y2=1.77
cc_4 VNB N_VGND_c_31_n 4.23625e-19 $X=-0.19 $Y=-0.245 $X2=2.415 $Y2=1.77
cc_5 VNB N_VGND_c_32_n 0.0371702f $X=-0.19 $Y=-0.245 $X2=5.095 $Y2=0.36
cc_6 VNB N_VGND_c_33_n 0.12354f $X=-0.19 $Y=-0.245 $X2=4.93 $Y2=0
cc_7 VNB N_VGND_c_34_n 0.0180543f $X=-0.19 $Y=-0.245 $X2=5.52 $Y2=0
cc_8 VNB N_VGND_c_35_n 0.327077f $X=-0.19 $Y=-0.245 $X2=5.52 $Y2=0
cc_9 VNB N_VGND_c_36_n 0.0279619f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=0
cc_10 VNB N_VGND_c_37_n 0.00513431f $X=-0.19 $Y=-0.245 $X2=5.04 $Y2=0
cc_11 VNB N_VPWR_c_57_n 0.0262142f $X=-0.19 $Y=-0.245 $X2=0.815 $Y2=0.38
cc_12 VNB N_VPWR_c_58_n 0.213478f $X=-0.19 $Y=-0.245 $X2=2.415 $Y2=1.77
cc_13 VNB N_VPWR_M1000_g 0.167743f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_VPWR_c_60_n 0.243291f $X=-0.19 $Y=-0.245 $X2=5.04 $Y2=0
cc_15 VPB N_VGND_c_28_n 0.401857f $X=-0.19 $Y=1.655 $X2=2.58 $Y2=2.555
cc_16 VPB N_VGND_c_30_n 0.0140672f $X=-0.19 $Y=1.655 $X2=0.98 $Y2=1.77
cc_17 VPB N_VGND_c_31_n 0.00875776f $X=-0.19 $Y=1.655 $X2=2.415 $Y2=1.77
cc_18 VPB N_VPWR_c_61_n 0.0425694f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_19 VPB N_VPWR_c_57_n 0.0010232f $X=-0.19 $Y=1.655 $X2=0.815 $Y2=0.38
cc_20 VPB N_VPWR_c_58_n 0.0404704f $X=-0.19 $Y=1.655 $X2=2.415 $Y2=1.77
cc_21 VPB N_VPWR_c_64_n 0.0654693f $X=-0.19 $Y=1.655 $X2=5.095 $Y2=0.085
cc_22 VPB N_VPWR_c_65_n 0.0204409f $X=-0.19 $Y=1.655 $X2=0.98 $Y2=0
cc_23 VPB N_VPWR_c_66_n 0.123858f $X=-0.19 $Y=1.655 $X2=4.56 $Y2=0
cc_24 VPB N_VPWR_c_67_n 0.0201227f $X=-0.19 $Y=1.655 $X2=5.095 $Y2=0
cc_25 VPB N_VPWR_c_60_n 0.08337f $X=-0.19 $Y=1.655 $X2=5.04 $Y2=0
cc_26 VPB N_VPWR_c_69_n 0.00516759f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_27 VPB N_VPWR_c_70_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_28 N_VGND_c_28_n N_VPWR_c_61_n 0.0546006f $X=2.58 $Y=2.555 $X2=0 $Y2=0
cc_29 N_VGND_c_30_n N_VPWR_c_61_n 0.0205458f $X=0.98 $Y=1.77 $X2=0 $Y2=0
cc_30 N_VGND_c_28_n N_VPWR_c_57_n 0.0149963f $X=2.58 $Y=2.555 $X2=0 $Y2=0
cc_31 N_VGND_c_31_n N_VPWR_c_57_n 0.00324791f $X=2.415 $Y=1.77 $X2=0 $Y2=0
cc_32 N_VGND_c_32_n N_VPWR_c_57_n 0.0180876f $X=5.095 $Y=0.36 $X2=0 $Y2=0
cc_33 N_VGND_c_28_n N_VPWR_c_58_n 0.151712f $X=2.58 $Y=2.555 $X2=0 $Y2=0
cc_34 N_VGND_c_32_n N_VPWR_c_58_n 0.0510144f $X=5.095 $Y=0.36 $X2=0 $Y2=0
cc_35 N_VGND_c_35_n N_VPWR_c_58_n 0.123649f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_36 N_VGND_c_28_n N_VPWR_c_64_n 0.0710714f $X=2.58 $Y=2.555 $X2=0 $Y2=0
cc_37 N_VGND_c_28_n N_VPWR_M1000_g 0.119822f $X=2.58 $Y=2.555 $X2=0 $Y2=0
cc_38 N_VGND_c_29_n N_VPWR_M1000_g 0.0654854f $X=0.815 $Y=0.38 $X2=0 $Y2=0
cc_39 N_VGND_c_31_n N_VPWR_M1000_g 0.0121106f $X=2.415 $Y=1.77 $X2=0 $Y2=0
cc_40 N_VGND_c_33_n N_VPWR_M1000_g 0.154094f $X=4.93 $Y=0 $X2=0 $Y2=0
cc_41 N_VGND_c_35_n N_VPWR_M1000_g 0.11988f $X=5.52 $Y=0 $X2=0 $Y2=0
cc_42 N_VGND_c_28_n N_VPWR_c_66_n 0.154485f $X=2.58 $Y=2.555 $X2=0 $Y2=0
cc_43 N_VGND_c_28_n N_VPWR_c_60_n 0.244147f $X=2.58 $Y=2.555 $X2=0 $Y2=0
