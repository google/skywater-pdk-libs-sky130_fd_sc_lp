* File: sky130_fd_sc_lp__dfrtp_2.pxi.spice
* Created: Wed Sep  2 09:43:47 2020
* 
x_PM_SKY130_FD_SC_LP__DFRTP_2%CLK N_CLK_M1009_g N_CLK_M1003_g N_CLK_c_261_n
+ N_CLK_c_266_n CLK CLK N_CLK_c_262_n N_CLK_c_263_n
+ PM_SKY130_FD_SC_LP__DFRTP_2%CLK
x_PM_SKY130_FD_SC_LP__DFRTP_2%A_27_101# N_A_27_101#_M1009_s N_A_27_101#_M1003_s
+ N_A_27_101#_c_296_n N_A_27_101#_M1019_g N_A_27_101#_M1021_g
+ N_A_27_101#_M1006_g N_A_27_101#_M1004_g N_A_27_101#_M1030_g
+ N_A_27_101#_M1012_g N_A_27_101#_c_298_n N_A_27_101#_c_299_n
+ N_A_27_101#_c_329_n N_A_27_101#_c_300_n N_A_27_101#_c_301_n
+ N_A_27_101#_c_330_n N_A_27_101#_c_302_n N_A_27_101#_c_303_n
+ N_A_27_101#_c_304_n N_A_27_101#_c_305_n N_A_27_101#_c_306_n
+ N_A_27_101#_c_360_p N_A_27_101#_c_307_n N_A_27_101#_c_447_p
+ N_A_27_101#_c_308_n N_A_27_101#_c_309_n N_A_27_101#_c_310_n
+ N_A_27_101#_c_311_n N_A_27_101#_c_373_p N_A_27_101#_c_376_p
+ N_A_27_101#_c_312_n N_A_27_101#_c_313_n N_A_27_101#_c_314_n
+ N_A_27_101#_c_332_n N_A_27_101#_c_315_n N_A_27_101#_c_316_n
+ N_A_27_101#_c_333_n N_A_27_101#_c_317_n N_A_27_101#_c_318_n
+ N_A_27_101#_c_319_n N_A_27_101#_c_320_n N_A_27_101#_c_452_p
+ N_A_27_101#_c_321_n N_A_27_101#_c_322_n N_A_27_101#_c_323_n
+ N_A_27_101#_c_324_n PM_SKY130_FD_SC_LP__DFRTP_2%A_27_101#
x_PM_SKY130_FD_SC_LP__DFRTP_2%D N_D_M1026_g N_D_c_573_n N_D_c_574_n N_D_M1002_g
+ N_D_c_579_n D N_D_c_577_n PM_SKY130_FD_SC_LP__DFRTP_2%D
x_PM_SKY130_FD_SC_LP__DFRTP_2%A_196_464# N_A_196_464#_M1021_d
+ N_A_196_464#_M1019_d N_A_196_464#_M1010_g N_A_196_464#_c_630_n
+ N_A_196_464#_M1023_g N_A_196_464#_M1020_g N_A_196_464#_c_633_n
+ N_A_196_464#_c_634_n N_A_196_464#_M1015_g N_A_196_464#_c_647_n
+ N_A_196_464#_c_648_n N_A_196_464#_c_635_n N_A_196_464#_c_649_n
+ N_A_196_464#_c_650_n N_A_196_464#_c_651_n N_A_196_464#_c_652_n
+ N_A_196_464#_c_653_n N_A_196_464#_c_636_n N_A_196_464#_c_637_n
+ N_A_196_464#_c_638_n N_A_196_464#_c_639_n N_A_196_464#_c_640_n
+ N_A_196_464#_c_768_p N_A_196_464#_c_641_n N_A_196_464#_c_642_n
+ N_A_196_464#_c_643_n PM_SKY130_FD_SC_LP__DFRTP_2%A_196_464#
x_PM_SKY130_FD_SC_LP__DFRTP_2%A_709_411# N_A_709_411#_M1017_d
+ N_A_709_411#_M1007_d N_A_709_411#_M1008_g N_A_709_411#_c_863_n
+ N_A_709_411#_c_864_n N_A_709_411#_c_857_n N_A_709_411#_c_866_n
+ N_A_709_411#_M1014_g N_A_709_411#_c_859_n N_A_709_411#_c_860_n
+ N_A_709_411#_c_861_n N_A_709_411#_c_909_p N_A_709_411#_c_869_n
+ PM_SKY130_FD_SC_LP__DFRTP_2%A_709_411#
x_PM_SKY130_FD_SC_LP__DFRTP_2%RESET_B N_RESET_B_c_944_n N_RESET_B_c_945_n
+ N_RESET_B_c_946_n N_RESET_B_M1001_g N_RESET_B_M1032_g N_RESET_B_c_948_n
+ N_RESET_B_c_956_n N_RESET_B_M1011_g N_RESET_B_c_957_n N_RESET_B_M1027_g
+ N_RESET_B_c_950_n N_RESET_B_M1028_g N_RESET_B_M1031_g N_RESET_B_c_961_n
+ N_RESET_B_c_952_n N_RESET_B_c_953_n N_RESET_B_c_962_n N_RESET_B_c_963_n
+ N_RESET_B_c_964_n N_RESET_B_c_1125_p N_RESET_B_c_997_n N_RESET_B_c_1126_p
+ N_RESET_B_c_965_n N_RESET_B_c_966_n N_RESET_B_c_967_n N_RESET_B_c_968_n
+ N_RESET_B_c_969_n RESET_B N_RESET_B_c_970_n N_RESET_B_c_971_n
+ N_RESET_B_c_972_n N_RESET_B_c_973_n PM_SKY130_FD_SC_LP__DFRTP_2%RESET_B
x_PM_SKY130_FD_SC_LP__DFRTP_2%A_573_535# N_A_573_535#_M1004_d
+ N_A_573_535#_M1010_d N_A_573_535#_M1011_d N_A_573_535#_c_1172_n
+ N_A_573_535#_c_1173_n N_A_573_535#_M1017_g N_A_573_535#_M1007_g
+ N_A_573_535#_c_1194_n N_A_573_535#_c_1180_n N_A_573_535#_c_1181_n
+ N_A_573_535#_c_1182_n N_A_573_535#_c_1174_n N_A_573_535#_c_1175_n
+ N_A_573_535#_c_1176_n N_A_573_535#_c_1183_n N_A_573_535#_c_1184_n
+ N_A_573_535#_c_1185_n N_A_573_535#_c_1186_n N_A_573_535#_c_1177_n
+ PM_SKY130_FD_SC_LP__DFRTP_2%A_573_535#
x_PM_SKY130_FD_SC_LP__DFRTP_2%A_1399_473# N_A_1399_473#_M1018_d
+ N_A_1399_473#_M1031_d N_A_1399_473#_M1005_g N_A_1399_473#_c_1303_n
+ N_A_1399_473#_M1024_g N_A_1399_473#_c_1305_n N_A_1399_473#_c_1306_n
+ N_A_1399_473#_c_1299_n N_A_1399_473#_c_1307_n N_A_1399_473#_c_1308_n
+ N_A_1399_473#_c_1300_n N_A_1399_473#_c_1310_n N_A_1399_473#_c_1311_n
+ N_A_1399_473#_c_1301_n N_A_1399_473#_c_1312_n
+ PM_SKY130_FD_SC_LP__DFRTP_2%A_1399_473#
x_PM_SKY130_FD_SC_LP__DFRTP_2%A_1252_451# N_A_1252_451#_M1020_d
+ N_A_1252_451#_M1030_d N_A_1252_451#_M1018_g N_A_1252_451#_c_1416_n
+ N_A_1252_451#_c_1417_n N_A_1252_451#_M1016_g N_A_1252_451#_c_1418_n
+ N_A_1252_451#_M1013_g N_A_1252_451#_c_1420_n N_A_1252_451#_M1000_g
+ N_A_1252_451#_c_1433_n N_A_1252_451#_c_1421_n N_A_1252_451#_c_1422_n
+ N_A_1252_451#_c_1434_n N_A_1252_451#_c_1423_n N_A_1252_451#_c_1424_n
+ N_A_1252_451#_c_1425_n N_A_1252_451#_c_1426_n N_A_1252_451#_c_1436_n
+ N_A_1252_451#_c_1427_n N_A_1252_451#_c_1428_n N_A_1252_451#_c_1437_n
+ N_A_1252_451#_c_1429_n PM_SKY130_FD_SC_LP__DFRTP_2%A_1252_451#
x_PM_SKY130_FD_SC_LP__DFRTP_2%A_1836_47# N_A_1836_47#_M1013_s
+ N_A_1836_47#_M1000_s N_A_1836_47#_M1022_g N_A_1836_47#_M1029_g
+ N_A_1836_47#_c_1564_n N_A_1836_47#_c_1565_n N_A_1836_47#_M1025_g
+ N_A_1836_47#_M1033_g N_A_1836_47#_c_1567_n N_A_1836_47#_c_1568_n
+ N_A_1836_47#_c_1569_n N_A_1836_47#_c_1570_n N_A_1836_47#_c_1571_n
+ N_A_1836_47#_c_1578_n N_A_1836_47#_c_1572_n N_A_1836_47#_c_1573_n
+ N_A_1836_47#_c_1574_n N_A_1836_47#_c_1575_n
+ PM_SKY130_FD_SC_LP__DFRTP_2%A_1836_47#
x_PM_SKY130_FD_SC_LP__DFRTP_2%VPWR N_VPWR_M1003_d N_VPWR_M1001_d N_VPWR_M1008_d
+ N_VPWR_M1007_s N_VPWR_M1005_d N_VPWR_M1016_d N_VPWR_M1000_d N_VPWR_M1033_s
+ N_VPWR_c_1649_n N_VPWR_c_1650_n N_VPWR_c_1651_n N_VPWR_c_1652_n
+ N_VPWR_c_1653_n N_VPWR_c_1654_n N_VPWR_c_1655_n N_VPWR_c_1656_n
+ N_VPWR_c_1657_n N_VPWR_c_1658_n N_VPWR_c_1659_n N_VPWR_c_1660_n VPWR
+ N_VPWR_c_1661_n N_VPWR_c_1662_n N_VPWR_c_1663_n N_VPWR_c_1664_n
+ N_VPWR_c_1665_n N_VPWR_c_1666_n N_VPWR_c_1667_n N_VPWR_c_1668_n
+ N_VPWR_c_1669_n N_VPWR_c_1670_n N_VPWR_c_1671_n N_VPWR_c_1648_n
+ PM_SKY130_FD_SC_LP__DFRTP_2%VPWR
x_PM_SKY130_FD_SC_LP__DFRTP_2%A_318_535# N_A_318_535#_M1002_d
+ N_A_318_535#_M1001_s N_A_318_535#_M1026_d N_A_318_535#_c_1807_n
+ N_A_318_535#_c_1808_n N_A_318_535#_c_1809_n N_A_318_535#_c_1810_n
+ N_A_318_535#_c_1811_n N_A_318_535#_c_1805_n N_A_318_535#_c_1812_n
+ N_A_318_535#_c_1813_n N_A_318_535#_c_1823_n N_A_318_535#_c_1806_n
+ PM_SKY130_FD_SC_LP__DFRTP_2%A_318_535#
x_PM_SKY130_FD_SC_LP__DFRTP_2%Q N_Q_M1022_d N_Q_M1029_d Q Q Q Q Q Q Q
+ N_Q_c_1895_n PM_SKY130_FD_SC_LP__DFRTP_2%Q
x_PM_SKY130_FD_SC_LP__DFRTP_2%VGND N_VGND_M1009_d N_VGND_M1032_s N_VGND_M1027_d
+ N_VGND_M1024_d N_VGND_M1013_d N_VGND_M1025_s N_VGND_c_1913_n N_VGND_c_1914_n
+ N_VGND_c_1915_n N_VGND_c_1916_n N_VGND_c_1917_n N_VGND_c_1918_n
+ N_VGND_c_1919_n N_VGND_c_1920_n N_VGND_c_1921_n N_VGND_c_1922_n
+ N_VGND_c_1923_n VGND N_VGND_c_1924_n N_VGND_c_1925_n N_VGND_c_1926_n
+ N_VGND_c_1927_n N_VGND_c_1928_n N_VGND_c_1929_n N_VGND_c_1930_n
+ N_VGND_c_1931_n PM_SKY130_FD_SC_LP__DFRTP_2%VGND
cc_1 VNB N_CLK_M1009_g 0.0498794f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.715
cc_2 VNB N_CLK_c_261_n 0.00317347f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.955
cc_3 VNB N_CLK_c_262_n 0.018564f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.615
cc_4 VNB N_CLK_c_263_n 0.00992817f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.615
cc_5 VNB N_A_27_101#_c_296_n 0.0228415f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_6 VNB N_A_27_101#_M1006_g 0.0116615f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.615
cc_7 VNB N_A_27_101#_c_298_n 0.00992859f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_27_101#_c_299_n 0.023525f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_27_101#_c_300_n 0.00605812f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_27_101#_c_301_n 0.0116439f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_27_101#_c_302_n 0.0159014f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_27_101#_c_303_n 0.00271285f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_27_101#_c_304_n 0.00356352f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_27_101#_c_305_n 0.0126784f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_27_101#_c_306_n 9.02063e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_27_101#_c_307_n 0.0106953f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_27_101#_c_308_n 0.00599719f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_27_101#_c_309_n 0.0163675f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_27_101#_c_310_n 0.00111447f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_27_101#_c_311_n 0.00637231f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_27_101#_c_312_n 0.00308383f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_27_101#_c_313_n 0.00142946f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_27_101#_c_314_n 0.00560177f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_27_101#_c_315_n 0.00726879f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_27_101#_c_316_n 0.0448783f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_27_101#_c_317_n 0.0049558f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_27_101#_c_318_n 0.0015602f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_27_101#_c_319_n 0.0246512f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_27_101#_c_320_n 0.0333628f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_27_101#_c_321_n 3.63984e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_27_101#_c_322_n 0.0181041f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_27_101#_c_323_n 0.0153635f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_27_101#_c_324_n 0.0159403f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_D_c_573_n 0.0378718f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.12
cc_35 VNB N_D_c_574_n 0.0189387f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.64
cc_36 VNB N_D_M1002_g 0.0226173f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.615
cc_37 VNB D 0.00290651f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_D_c_577_n 0.0261483f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.615
cc_39 VNB N_A_196_464#_c_630_n 0.0339787f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.955
cc_40 VNB N_A_196_464#_M1023_g 0.0184449f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_41 VNB N_A_196_464#_M1020_g 0.0374049f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.615
cc_42 VNB N_A_196_464#_c_633_n 0.0417303f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.615
cc_43 VNB N_A_196_464#_c_634_n 0.00824362f $X=-0.19 $Y=-0.245 $X2=0.312
+ $Y2=1.615
cc_44 VNB N_A_196_464#_c_635_n 0.0121119f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_196_464#_c_636_n 0.00744561f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_196_464#_c_637_n 3.31215e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_196_464#_c_638_n 0.0105376f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_196_464#_c_639_n 0.00674616f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_196_464#_c_640_n 0.00830966f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_196_464#_c_641_n 0.0118515f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_196_464#_c_642_n 0.0014378f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_196_464#_c_643_n 0.00385617f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_709_411#_c_857_n 0.0213261f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_54 VNB N_A_709_411#_M1014_g 0.0299691f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.615
cc_55 VNB N_A_709_411#_c_859_n 0.0111938f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.615
cc_56 VNB N_A_709_411#_c_860_n 0.0112971f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_709_411#_c_861_n 0.0019574f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_RESET_B_c_944_n 0.0855113f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.715
cc_59 VNB N_RESET_B_c_945_n 0.0336798f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.715
cc_60 VNB N_RESET_B_c_946_n 0.012806f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_RESET_B_M1032_g 0.0179426f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.955
cc_62 VNB N_RESET_B_c_948_n 0.179994f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_63 VNB N_RESET_B_M1027_g 0.0276392f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_RESET_B_c_950_n 0.0221122f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_RESET_B_M1028_g 0.0428935f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_RESET_B_c_952_n 0.00749069f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_RESET_B_c_953_n 0.0103168f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_A_573_535#_c_1172_n 0.0157306f $X=-0.19 $Y=-0.245 $X2=0.385
+ $Y2=1.955
cc_69 VNB N_A_573_535#_c_1173_n 0.0204288f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=2.12
cc_70 VNB N_A_573_535#_c_1174_n 0.00203566f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_A_573_535#_c_1175_n 0.00216664f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_A_573_535#_c_1176_n 0.0165669f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_A_573_535#_c_1177_n 0.0444957f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_A_1399_473#_M1024_g 0.0449072f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_A_1399_473#_c_1299_n 0.0257214f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_A_1399_473#_c_1300_n 0.00789141f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_A_1399_473#_c_1301_n 0.0126007f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_A_1252_451#_M1018_g 0.0310529f $X=-0.19 $Y=-0.245 $X2=0.385
+ $Y2=1.615
cc_79 VNB N_A_1252_451#_c_1416_n 0.0155198f $X=-0.19 $Y=-0.245 $X2=0.385
+ $Y2=1.955
cc_80 VNB N_A_1252_451#_c_1417_n 0.00600108f $X=-0.19 $Y=-0.245 $X2=0.385
+ $Y2=2.12
cc_81 VNB N_A_1252_451#_c_1418_n 0.0319508f $X=-0.19 $Y=-0.245 $X2=0.385
+ $Y2=1.615
cc_82 VNB N_A_1252_451#_M1013_g 0.0549897f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_A_1252_451#_c_1420_n 0.0126556f $X=-0.19 $Y=-0.245 $X2=0.312
+ $Y2=2.035
cc_84 VNB N_A_1252_451#_c_1421_n 0.0136482f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_A_1252_451#_c_1422_n 0.00391059f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_A_1252_451#_c_1423_n 7.14815e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_A_1252_451#_c_1424_n 0.00337964f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_A_1252_451#_c_1425_n 0.0105655f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_A_1252_451#_c_1426_n 0.0206938f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_A_1252_451#_c_1427_n 0.00210256f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_A_1252_451#_c_1428_n 0.0112078f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_A_1252_451#_c_1429_n 0.0201888f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_93 VNB N_A_1836_47#_M1029_g 0.00800597f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=2.12
cc_94 VNB N_A_1836_47#_c_1564_n 0.0101534f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.95
cc_95 VNB N_A_1836_47#_c_1565_n 0.0215271f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_96 VNB N_A_1836_47#_M1033_g 0.0255672f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_97 VNB N_A_1836_47#_c_1567_n 0.0106787f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_98 VNB N_A_1836_47#_c_1568_n 0.0150542f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_99 VNB N_A_1836_47#_c_1569_n 0.00788177f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_100 VNB N_A_1836_47#_c_1570_n 0.00874635f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_101 VNB N_A_1836_47#_c_1571_n 0.00687201f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_102 VNB N_A_1836_47#_c_1572_n 9.62749e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_103 VNB N_A_1836_47#_c_1573_n 0.00146498f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_104 VNB N_A_1836_47#_c_1574_n 0.0313477f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_105 VNB N_A_1836_47#_c_1575_n 0.0174449f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_106 VNB N_VPWR_c_1648_n 0.462217f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_107 VNB N_A_318_535#_c_1805_n 0.00668304f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_108 VNB N_A_318_535#_c_1806_n 0.00466783f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_109 VNB N_Q_c_1895_n 0.00844637f $X=-0.19 $Y=-0.245 $X2=0.312 $Y2=1.665
cc_110 VNB N_VGND_c_1913_n 0.0156267f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_111 VNB N_VGND_c_1914_n 0.00237577f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_112 VNB N_VGND_c_1915_n 0.00983419f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_113 VNB N_VGND_c_1916_n 0.0185424f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_114 VNB N_VGND_c_1917_n 0.00344689f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_115 VNB N_VGND_c_1918_n 0.0117031f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_116 VNB N_VGND_c_1919_n 0.0496202f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_117 VNB N_VGND_c_1920_n 0.0710942f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_118 VNB N_VGND_c_1921_n 0.00516907f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_119 VNB N_VGND_c_1922_n 0.0533726f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_120 VNB N_VGND_c_1923_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_121 VNB N_VGND_c_1924_n 0.0184044f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_122 VNB N_VGND_c_1925_n 0.0291036f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_123 VNB N_VGND_c_1926_n 0.0495733f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_124 VNB N_VGND_c_1927_n 0.014797f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_125 VNB N_VGND_c_1928_n 0.00432782f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_126 VNB N_VGND_c_1929_n 0.00326264f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_127 VNB N_VGND_c_1930_n 0.00785353f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_128 VNB N_VGND_c_1931_n 0.586985f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_129 VPB N_CLK_M1003_g 0.0302639f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.64
cc_130 VPB N_CLK_c_261_n 0.0247109f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.955
cc_131 VPB N_CLK_c_266_n 0.0188165f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=2.12
cc_132 VPB N_CLK_c_263_n 0.0195636f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.615
cc_133 VPB N_A_27_101#_M1019_g 0.0481866f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.955
cc_134 VPB N_A_27_101#_M1006_g 0.0654305f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.615
cc_135 VPB N_A_27_101#_M1030_g 0.0214243f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_136 VPB N_A_27_101#_c_298_n 0.0099246f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_137 VPB N_A_27_101#_c_329_n 0.004186f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_138 VPB N_A_27_101#_c_330_n 0.00420065f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_139 VPB N_A_27_101#_c_314_n 0.00198741f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_140 VPB N_A_27_101#_c_332_n 0.0368368f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_141 VPB N_A_27_101#_c_333_n 0.0322901f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_142 VPB N_A_27_101#_c_317_n 0.00342268f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_143 VPB N_D_M1026_g 0.0524042f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.715
cc_144 VPB N_D_c_579_n 0.0236052f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.95
cc_145 VPB D 0.00286922f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_146 VPB N_D_c_577_n 0.00655157f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.615
cc_147 VPB N_A_196_464#_M1010_g 0.0322635f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.615
cc_148 VPB N_A_196_464#_c_630_n 0.0162902f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.955
cc_149 VPB N_A_196_464#_M1015_g 0.0405081f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_150 VPB N_A_196_464#_c_647_n 0.0303142f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_151 VPB N_A_196_464#_c_648_n 0.0121003f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_152 VPB N_A_196_464#_c_649_n 0.00696269f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_153 VPB N_A_196_464#_c_650_n 0.0157762f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_154 VPB N_A_196_464#_c_651_n 0.0173691f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_155 VPB N_A_196_464#_c_652_n 0.00241298f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_156 VPB N_A_196_464#_c_653_n 0.0335666f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_157 VPB N_A_196_464#_c_636_n 0.0126075f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_158 VPB N_A_196_464#_c_637_n 3.31215e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_159 VPB N_A_196_464#_c_638_n 0.0180796f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_160 VPB N_A_196_464#_c_639_n 0.00177431f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_161 VPB N_A_196_464#_c_640_n 0.00497027f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_162 VPB N_A_196_464#_c_641_n 0.0198035f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_163 VPB N_A_196_464#_c_642_n 0.00152246f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_164 VPB N_A_196_464#_c_643_n 0.00275523f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_165 VPB N_A_709_411#_M1008_g 0.0337036f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.615
cc_166 VPB N_A_709_411#_c_863_n 0.0352582f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.955
cc_167 VPB N_A_709_411#_c_864_n 0.00782356f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=2.12
cc_168 VPB N_A_709_411#_c_857_n 0.0126691f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_169 VPB N_A_709_411#_c_866_n 0.0199932f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.95
cc_170 VPB N_A_709_411#_c_859_n 0.00484021f $X=-0.19 $Y=1.655 $X2=0.385
+ $Y2=1.615
cc_171 VPB N_A_709_411#_c_861_n 3.24298e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_172 VPB N_A_709_411#_c_869_n 0.0120646f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_173 VPB N_RESET_B_c_944_n 0.026181f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.715
cc_174 VPB N_RESET_B_M1001_g 0.0373959f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.64
cc_175 VPB N_RESET_B_c_956_n 0.0197123f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_176 VPB N_RESET_B_c_957_n 0.0080737f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.615
cc_177 VPB N_RESET_B_c_950_n 0.0334177f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_178 VPB N_RESET_B_M1028_g 5.87215e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_179 VPB N_RESET_B_M1031_g 0.0325455f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_180 VPB N_RESET_B_c_961_n 0.0249941f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_181 VPB N_RESET_B_c_962_n 0.0283571f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_182 VPB N_RESET_B_c_963_n 0.0153767f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_183 VPB N_RESET_B_c_964_n 0.00675311f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_184 VPB N_RESET_B_c_965_n 6.99208e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_185 VPB N_RESET_B_c_966_n 0.00480896f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_186 VPB N_RESET_B_c_967_n 0.00777951f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_187 VPB N_RESET_B_c_968_n 0.00340604f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_188 VPB N_RESET_B_c_969_n 0.010793f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_189 VPB N_RESET_B_c_970_n 0.0241575f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_190 VPB N_RESET_B_c_971_n 0.00581296f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_191 VPB N_RESET_B_c_972_n 0.0287064f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_192 VPB N_RESET_B_c_973_n 0.0453962f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_193 VPB N_A_573_535#_c_1172_n 0.00697732f $X=-0.19 $Y=1.655 $X2=0.385
+ $Y2=1.955
cc_194 VPB N_A_573_535#_M1007_g 0.0238374f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.615
cc_195 VPB N_A_573_535#_c_1180_n 0.00289503f $X=-0.19 $Y=1.655 $X2=0.312
+ $Y2=2.035
cc_196 VPB N_A_573_535#_c_1181_n 0.0114661f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_197 VPB N_A_573_535#_c_1182_n 0.00297798f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_198 VPB N_A_573_535#_c_1183_n 0.0161176f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_199 VPB N_A_573_535#_c_1184_n 0.0125379f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_200 VPB N_A_573_535#_c_1185_n 0.0448928f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_201 VPB N_A_573_535#_c_1186_n 0.00608073f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_202 VPB N_A_1399_473#_M1005_g 0.022965f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.615
cc_203 VPB N_A_1399_473#_c_1303_n 0.00597564f $X=-0.19 $Y=1.655 $X2=0.385
+ $Y2=2.12
cc_204 VPB N_A_1399_473#_M1024_g 0.0281924f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_205 VPB N_A_1399_473#_c_1305_n 0.00649178f $X=-0.19 $Y=1.655 $X2=0.385
+ $Y2=1.615
cc_206 VPB N_A_1399_473#_c_1306_n 0.00125597f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_207 VPB N_A_1399_473#_c_1307_n 0.016261f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_208 VPB N_A_1399_473#_c_1308_n 0.00970623f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_209 VPB N_A_1399_473#_c_1300_n 0.01012f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_210 VPB N_A_1399_473#_c_1310_n 0.005248f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_211 VPB N_A_1399_473#_c_1311_n 0.0462195f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_212 VPB N_A_1399_473#_c_1312_n 0.0174211f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_213 VPB N_A_1252_451#_M1016_g 0.0529498f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_214 VPB N_A_1252_451#_c_1420_n 0.0060397f $X=-0.19 $Y=1.655 $X2=0.312
+ $Y2=2.035
cc_215 VPB N_A_1252_451#_M1000_g 0.0493991f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_216 VPB N_A_1252_451#_c_1433_n 0.0185692f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_217 VPB N_A_1252_451#_c_1434_n 0.0144999f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_218 VPB N_A_1252_451#_c_1424_n 0.0057291f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_219 VPB N_A_1252_451#_c_1436_n 3.11212e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_220 VPB N_A_1252_451#_c_1437_n 0.0012329f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_221 VPB N_A_1252_451#_c_1429_n 0.0147588f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_222 VPB N_A_1836_47#_M1029_g 0.0208864f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=2.12
cc_223 VPB N_A_1836_47#_M1033_g 0.0272176f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_224 VPB N_A_1836_47#_c_1578_n 0.008108f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_225 VPB N_A_1836_47#_c_1572_n 0.00632237f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_226 VPB N_VPWR_c_1649_n 0.00396467f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_227 VPB N_VPWR_c_1650_n 4.89148e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_228 VPB N_VPWR_c_1651_n 0.00507815f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_229 VPB N_VPWR_c_1652_n 0.0121651f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_230 VPB N_VPWR_c_1653_n 0.00621655f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_231 VPB N_VPWR_c_1654_n 0.0101483f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_232 VPB N_VPWR_c_1655_n 0.0116772f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_233 VPB N_VPWR_c_1656_n 0.0656709f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_234 VPB N_VPWR_c_1657_n 0.0352636f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_235 VPB N_VPWR_c_1658_n 0.00459098f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_236 VPB N_VPWR_c_1659_n 0.0313545f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_237 VPB N_VPWR_c_1660_n 0.00497514f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_238 VPB N_VPWR_c_1661_n 0.0167155f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_239 VPB N_VPWR_c_1662_n 0.0296156f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_240 VPB N_VPWR_c_1663_n 0.011965f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_241 VPB N_VPWR_c_1664_n 0.0187941f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_242 VPB N_VPWR_c_1665_n 0.0147711f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_243 VPB N_VPWR_c_1666_n 0.00601644f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_244 VPB N_VPWR_c_1667_n 0.00436716f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_245 VPB N_VPWR_c_1668_n 0.0441543f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_246 VPB N_VPWR_c_1669_n 0.0234374f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_247 VPB N_VPWR_c_1670_n 0.00506755f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_248 VPB N_VPWR_c_1671_n 0.00520126f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_249 VPB N_VPWR_c_1648_n 0.0818225f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_250 VPB N_A_318_535#_c_1807_n 0.00626478f $X=-0.19 $Y=1.655 $X2=0.385
+ $Y2=2.12
cc_251 VPB N_A_318_535#_c_1808_n 0.00636642f $X=-0.19 $Y=1.655 $X2=0.155
+ $Y2=1.95
cc_252 VPB N_A_318_535#_c_1809_n 0.00399218f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_253 VPB N_A_318_535#_c_1810_n 0.00139619f $X=-0.19 $Y=1.655 $X2=0.385
+ $Y2=1.615
cc_254 VPB N_A_318_535#_c_1811_n 0.00736942f $X=-0.19 $Y=1.655 $X2=0.312
+ $Y2=1.615
cc_255 VPB N_A_318_535#_c_1812_n 0.00634309f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_256 VPB N_A_318_535#_c_1813_n 0.00186219f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_257 VPB N_A_318_535#_c_1806_n 0.00385634f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_258 VPB N_Q_c_1895_n 0.00467442f $X=-0.19 $Y=1.655 $X2=0.312 $Y2=1.665
cc_259 N_CLK_c_262_n N_A_27_101#_c_296_n 0.0116281f $X=0.385 $Y=1.615 $X2=0
+ $Y2=0
cc_260 N_CLK_c_263_n N_A_27_101#_c_296_n 2.28868e-19 $X=0.385 $Y=1.615 $X2=0
+ $Y2=0
cc_261 N_CLK_c_261_n N_A_27_101#_M1019_g 0.0424871f $X=0.385 $Y=1.955 $X2=0
+ $Y2=0
cc_262 N_CLK_c_263_n N_A_27_101#_M1019_g 3.63795e-19 $X=0.385 $Y=1.615 $X2=0
+ $Y2=0
cc_263 N_CLK_c_261_n N_A_27_101#_c_298_n 0.0116281f $X=0.385 $Y=1.955 $X2=0
+ $Y2=0
cc_264 N_CLK_M1009_g N_A_27_101#_c_299_n 0.00549066f $X=0.475 $Y=0.715 $X2=0
+ $Y2=0
cc_265 N_CLK_M1003_g N_A_27_101#_c_329_n 0.0125058f $X=0.475 $Y=2.64 $X2=0 $Y2=0
cc_266 N_CLK_c_266_n N_A_27_101#_c_329_n 3.07325e-19 $X=0.385 $Y=2.12 $X2=0
+ $Y2=0
cc_267 N_CLK_c_263_n N_A_27_101#_c_329_n 0.0084158f $X=0.385 $Y=1.615 $X2=0
+ $Y2=0
cc_268 N_CLK_M1009_g N_A_27_101#_c_300_n 0.0178855f $X=0.475 $Y=0.715 $X2=0
+ $Y2=0
cc_269 N_CLK_c_263_n N_A_27_101#_c_300_n 0.00574094f $X=0.385 $Y=1.615 $X2=0
+ $Y2=0
cc_270 N_CLK_c_262_n N_A_27_101#_c_301_n 0.00132139f $X=0.385 $Y=1.615 $X2=0
+ $Y2=0
cc_271 N_CLK_c_263_n N_A_27_101#_c_301_n 0.0202468f $X=0.385 $Y=1.615 $X2=0
+ $Y2=0
cc_272 N_CLK_c_261_n N_A_27_101#_c_330_n 0.00680351f $X=0.385 $Y=1.955 $X2=0
+ $Y2=0
cc_273 N_CLK_M1003_g N_A_27_101#_c_333_n 2.21843e-19 $X=0.475 $Y=2.64 $X2=0
+ $Y2=0
cc_274 N_CLK_c_266_n N_A_27_101#_c_333_n 0.0010425f $X=0.385 $Y=2.12 $X2=0 $Y2=0
cc_275 N_CLK_c_263_n N_A_27_101#_c_333_n 0.0172425f $X=0.385 $Y=1.615 $X2=0
+ $Y2=0
cc_276 N_CLK_M1009_g N_A_27_101#_c_317_n 0.00699423f $X=0.475 $Y=0.715 $X2=0
+ $Y2=0
cc_277 N_CLK_c_263_n N_A_27_101#_c_317_n 0.0465708f $X=0.385 $Y=1.615 $X2=0
+ $Y2=0
cc_278 N_CLK_M1009_g N_A_27_101#_c_318_n 0.00114972f $X=0.475 $Y=0.715 $X2=0
+ $Y2=0
cc_279 N_CLK_M1009_g N_A_27_101#_c_319_n 0.0116281f $X=0.475 $Y=0.715 $X2=0
+ $Y2=0
cc_280 N_CLK_M1009_g N_A_27_101#_c_322_n 0.0099183f $X=0.475 $Y=0.715 $X2=0
+ $Y2=0
cc_281 N_CLK_M1003_g N_VPWR_c_1649_n 0.0109495f $X=0.475 $Y=2.64 $X2=0 $Y2=0
cc_282 N_CLK_M1003_g N_VPWR_c_1661_n 0.00383152f $X=0.475 $Y=2.64 $X2=0 $Y2=0
cc_283 N_CLK_M1003_g N_VPWR_c_1648_n 0.00391732f $X=0.475 $Y=2.64 $X2=0 $Y2=0
cc_284 N_CLK_M1009_g N_VGND_c_1913_n 0.00385181f $X=0.475 $Y=0.715 $X2=0 $Y2=0
cc_285 N_CLK_M1009_g N_VGND_c_1924_n 0.00484506f $X=0.475 $Y=0.715 $X2=0 $Y2=0
cc_286 N_CLK_M1009_g N_VGND_c_1931_n 0.00503886f $X=0.475 $Y=0.715 $X2=0 $Y2=0
cc_287 N_A_27_101#_c_305_n N_D_c_573_n 0.00691999f $X=2.41 $Y=0.955 $X2=0 $Y2=0
cc_288 N_A_27_101#_c_305_n N_D_c_574_n 0.00390334f $X=2.41 $Y=0.955 $X2=0 $Y2=0
cc_289 N_A_27_101#_c_305_n N_D_M1002_g 0.00252978f $X=2.41 $Y=0.955 $X2=0 $Y2=0
cc_290 N_A_27_101#_c_360_p N_D_M1002_g 0.00502094f $X=2.495 $Y=0.87 $X2=0 $Y2=0
cc_291 N_A_27_101#_c_307_n N_D_M1002_g 0.00347885f $X=3.33 $Y=0.362 $X2=0 $Y2=0
cc_292 N_A_27_101#_c_308_n N_D_M1002_g 0.00119227f $X=3.415 $Y=1.14 $X2=0 $Y2=0
cc_293 N_A_27_101#_c_320_n N_D_M1002_g 0.0145731f $X=3.3 $Y=1.3 $X2=0 $Y2=0
cc_294 N_A_27_101#_c_323_n N_D_M1002_g 0.0117037f $X=3.3 $Y=1.135 $X2=0 $Y2=0
cc_295 N_A_27_101#_c_305_n D 0.0254764f $X=2.41 $Y=0.955 $X2=0 $Y2=0
cc_296 N_A_27_101#_M1006_g N_A_196_464#_M1010_g 0.0219289f $X=3.26 $Y=2.885
+ $X2=0 $Y2=0
cc_297 N_A_27_101#_M1006_g N_A_196_464#_c_630_n 0.0132527f $X=3.26 $Y=2.885
+ $X2=0 $Y2=0
cc_298 N_A_27_101#_c_308_n N_A_196_464#_c_630_n 0.00150088f $X=3.415 $Y=1.14
+ $X2=0 $Y2=0
cc_299 N_A_27_101#_c_320_n N_A_196_464#_c_630_n 0.00830992f $X=3.3 $Y=1.3 $X2=0
+ $Y2=0
cc_300 N_A_27_101#_c_308_n N_A_196_464#_M1023_g 0.00213851f $X=3.415 $Y=1.14
+ $X2=0 $Y2=0
cc_301 N_A_27_101#_c_309_n N_A_196_464#_M1023_g 0.00535437f $X=4.05 $Y=0.362
+ $X2=0 $Y2=0
cc_302 N_A_27_101#_c_310_n N_A_196_464#_M1023_g 0.00647446f $X=4.135 $Y=0.805
+ $X2=0 $Y2=0
cc_303 N_A_27_101#_c_373_p N_A_196_464#_M1023_g 0.00315998f $X=4.22 $Y=0.89
+ $X2=0 $Y2=0
cc_304 N_A_27_101#_c_320_n N_A_196_464#_M1023_g 0.00163858f $X=3.3 $Y=1.3 $X2=0
+ $Y2=0
cc_305 N_A_27_101#_c_323_n N_A_196_464#_M1023_g 0.00732488f $X=3.3 $Y=1.135
+ $X2=0 $Y2=0
cc_306 N_A_27_101#_c_376_p N_A_196_464#_M1020_g 2.10461e-19 $X=5.57 $Y=0.805
+ $X2=0 $Y2=0
cc_307 N_A_27_101#_c_314_n N_A_196_464#_M1020_g 0.0258025f $X=6.26 $Y=1.91 $X2=0
+ $Y2=0
cc_308 N_A_27_101#_c_315_n N_A_196_464#_M1020_g 0.00430702f $X=7.01 $Y=0.35
+ $X2=0 $Y2=0
cc_309 N_A_27_101#_c_316_n N_A_196_464#_M1020_g 0.0199719f $X=7.01 $Y=0.35 $X2=0
+ $Y2=0
cc_310 N_A_27_101#_c_321_n N_A_196_464#_M1020_g 0.00596145f $X=6.265 $Y=0.345
+ $X2=0 $Y2=0
cc_311 N_A_27_101#_c_324_n N_A_196_464#_c_633_n 0.00686857f $X=7.01 $Y=0.515
+ $X2=0 $Y2=0
cc_312 N_A_27_101#_c_314_n N_A_196_464#_c_634_n 0.00724468f $X=6.26 $Y=1.91
+ $X2=0 $Y2=0
cc_313 N_A_27_101#_c_332_n N_A_196_464#_c_634_n 0.0133183f $X=6.26 $Y=1.91 $X2=0
+ $Y2=0
cc_314 N_A_27_101#_M1030_g N_A_196_464#_c_647_n 0.0298296f $X=6.185 $Y=2.675
+ $X2=0 $Y2=0
cc_315 N_A_27_101#_M1019_g N_A_196_464#_c_648_n 0.00153613f $X=0.905 $Y=2.64
+ $X2=0 $Y2=0
cc_316 N_A_27_101#_c_329_n N_A_196_464#_c_648_n 0.00725482f $X=0.665 $Y=2.385
+ $X2=0 $Y2=0
cc_317 N_A_27_101#_c_330_n N_A_196_464#_c_648_n 0.00303369f $X=0.75 $Y=2.3 $X2=0
+ $Y2=0
cc_318 N_A_27_101#_c_302_n N_A_196_464#_c_635_n 0.0145595f $X=1.655 $Y=0.34
+ $X2=0 $Y2=0
cc_319 N_A_27_101#_c_304_n N_A_196_464#_c_635_n 0.0194404f $X=1.74 $Y=0.87 $X2=0
+ $Y2=0
cc_320 N_A_27_101#_c_306_n N_A_196_464#_c_635_n 0.0136205f $X=1.825 $Y=0.955
+ $X2=0 $Y2=0
cc_321 N_A_27_101#_c_318_n N_A_196_464#_c_635_n 0.0669909f $X=0.895 $Y=1.1 $X2=0
+ $Y2=0
cc_322 N_A_27_101#_c_322_n N_A_196_464#_c_635_n 0.00753584f $X=0.972 $Y=1.035
+ $X2=0 $Y2=0
cc_323 N_A_27_101#_M1019_g N_A_196_464#_c_649_n 0.00233752f $X=0.905 $Y=2.64
+ $X2=0 $Y2=0
cc_324 N_A_27_101#_c_330_n N_A_196_464#_c_649_n 0.00870842f $X=0.75 $Y=2.3 $X2=0
+ $Y2=0
cc_325 N_A_27_101#_M1019_g N_A_196_464#_c_651_n 0.00213121f $X=0.905 $Y=2.64
+ $X2=0 $Y2=0
cc_326 N_A_27_101#_c_298_n N_A_196_464#_c_651_n 0.00160924f $X=0.972 $Y=1.705
+ $X2=0 $Y2=0
cc_327 N_A_27_101#_c_330_n N_A_196_464#_c_651_n 0.0124681f $X=0.75 $Y=2.3 $X2=0
+ $Y2=0
cc_328 N_A_27_101#_c_317_n N_A_196_464#_c_651_n 0.00431851f $X=0.895 $Y=1.185
+ $X2=0 $Y2=0
cc_329 N_A_27_101#_M1006_g N_A_196_464#_c_652_n 3.01767e-19 $X=3.26 $Y=2.885
+ $X2=0 $Y2=0
cc_330 N_A_27_101#_M1006_g N_A_196_464#_c_653_n 0.0203599f $X=3.26 $Y=2.885
+ $X2=0 $Y2=0
cc_331 N_A_27_101#_M1006_g N_A_196_464#_c_636_n 0.00557535f $X=3.26 $Y=2.885
+ $X2=0 $Y2=0
cc_332 N_A_27_101#_c_305_n N_A_196_464#_c_636_n 0.0151921f $X=2.41 $Y=0.955
+ $X2=0 $Y2=0
cc_333 N_A_27_101#_c_308_n N_A_196_464#_c_636_n 0.00773838f $X=3.415 $Y=1.14
+ $X2=0 $Y2=0
cc_334 N_A_27_101#_c_320_n N_A_196_464#_c_636_n 0.00205331f $X=3.3 $Y=1.3 $X2=0
+ $Y2=0
cc_335 N_A_27_101#_c_306_n N_A_196_464#_c_637_n 0.00116209f $X=1.825 $Y=0.955
+ $X2=0 $Y2=0
cc_336 N_A_27_101#_c_317_n N_A_196_464#_c_637_n 6.68146e-19 $X=0.895 $Y=1.185
+ $X2=0 $Y2=0
cc_337 N_A_27_101#_c_311_n N_A_196_464#_c_638_n 3.37845e-19 $X=5.485 $Y=0.89
+ $X2=0 $Y2=0
cc_338 N_A_27_101#_c_314_n N_A_196_464#_c_638_n 0.0156358f $X=6.26 $Y=1.91 $X2=0
+ $Y2=0
cc_339 N_A_27_101#_c_332_n N_A_196_464#_c_638_n 0.00342731f $X=6.26 $Y=1.91
+ $X2=0 $Y2=0
cc_340 N_A_27_101#_M1006_g N_A_196_464#_c_639_n 6.0018e-19 $X=3.26 $Y=2.885
+ $X2=0 $Y2=0
cc_341 N_A_27_101#_c_308_n N_A_196_464#_c_639_n 0.00124885f $X=3.415 $Y=1.14
+ $X2=0 $Y2=0
cc_342 N_A_27_101#_c_320_n N_A_196_464#_c_639_n 2.72074e-19 $X=3.3 $Y=1.3 $X2=0
+ $Y2=0
cc_343 N_A_27_101#_c_296_n N_A_196_464#_c_640_n 0.00194431f $X=0.972 $Y=1.523
+ $X2=0 $Y2=0
cc_344 N_A_27_101#_M1019_g N_A_196_464#_c_640_n 0.00127644f $X=0.905 $Y=2.64
+ $X2=0 $Y2=0
cc_345 N_A_27_101#_c_330_n N_A_196_464#_c_640_n 0.00464808f $X=0.75 $Y=2.3 $X2=0
+ $Y2=0
cc_346 N_A_27_101#_c_306_n N_A_196_464#_c_640_n 0.00536286f $X=1.825 $Y=0.955
+ $X2=0 $Y2=0
cc_347 N_A_27_101#_c_317_n N_A_196_464#_c_640_n 0.0166262f $X=0.895 $Y=1.185
+ $X2=0 $Y2=0
cc_348 N_A_27_101#_c_314_n N_A_196_464#_c_641_n 0.00134199f $X=6.26 $Y=1.91
+ $X2=0 $Y2=0
cc_349 N_A_27_101#_c_332_n N_A_196_464#_c_641_n 0.0204574f $X=6.26 $Y=1.91 $X2=0
+ $Y2=0
cc_350 N_A_27_101#_M1006_g N_A_196_464#_c_643_n 0.00143807f $X=3.26 $Y=2.885
+ $X2=0 $Y2=0
cc_351 N_A_27_101#_c_308_n N_A_196_464#_c_643_n 0.00573238f $X=3.415 $Y=1.14
+ $X2=0 $Y2=0
cc_352 N_A_27_101#_c_320_n N_A_196_464#_c_643_n 0.00123167f $X=3.3 $Y=1.3 $X2=0
+ $Y2=0
cc_353 N_A_27_101#_c_312_n N_A_709_411#_M1017_d 0.00871221f $X=6.175 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_354 N_A_27_101#_M1006_g N_A_709_411#_c_864_n 0.0716219f $X=3.26 $Y=2.885
+ $X2=0 $Y2=0
cc_355 N_A_27_101#_c_310_n N_A_709_411#_M1014_g 0.00355727f $X=4.135 $Y=0.805
+ $X2=0 $Y2=0
cc_356 N_A_27_101#_c_311_n N_A_709_411#_M1014_g 0.00987813f $X=5.485 $Y=0.89
+ $X2=0 $Y2=0
cc_357 N_A_27_101#_c_311_n N_A_709_411#_c_859_n 2.82186e-19 $X=5.485 $Y=0.89
+ $X2=0 $Y2=0
cc_358 N_A_27_101#_c_311_n N_A_709_411#_c_860_n 0.00788523f $X=5.485 $Y=0.89
+ $X2=0 $Y2=0
cc_359 N_A_27_101#_c_312_n N_A_709_411#_c_860_n 0.013472f $X=6.175 $Y=0.34 $X2=0
+ $Y2=0
cc_360 N_A_27_101#_c_314_n N_A_709_411#_c_860_n 0.0541208f $X=6.26 $Y=1.91 $X2=0
+ $Y2=0
cc_361 N_A_27_101#_c_314_n N_A_709_411#_c_861_n 0.0142872f $X=6.26 $Y=1.91 $X2=0
+ $Y2=0
cc_362 N_A_27_101#_M1030_g N_A_709_411#_c_869_n 0.00330902f $X=6.185 $Y=2.675
+ $X2=0 $Y2=0
cc_363 N_A_27_101#_c_314_n N_A_709_411#_c_869_n 0.0286568f $X=6.26 $Y=1.91 $X2=0
+ $Y2=0
cc_364 N_A_27_101#_c_332_n N_A_709_411#_c_869_n 0.00288222f $X=6.26 $Y=1.91
+ $X2=0 $Y2=0
cc_365 N_A_27_101#_M1019_g N_RESET_B_c_944_n 0.00643547f $X=0.905 $Y=2.64 $X2=0
+ $Y2=0
cc_366 N_A_27_101#_c_302_n N_RESET_B_c_944_n 0.00932968f $X=1.655 $Y=0.34 $X2=0
+ $Y2=0
cc_367 N_A_27_101#_c_304_n N_RESET_B_c_944_n 0.0123559f $X=1.74 $Y=0.87 $X2=0
+ $Y2=0
cc_368 N_A_27_101#_c_306_n N_RESET_B_c_944_n 0.00878148f $X=1.825 $Y=0.955 $X2=0
+ $Y2=0
cc_369 N_A_27_101#_c_318_n N_RESET_B_c_944_n 8.21274e-19 $X=0.895 $Y=1.1 $X2=0
+ $Y2=0
cc_370 N_A_27_101#_c_322_n N_RESET_B_c_944_n 0.0256517f $X=0.972 $Y=1.035 $X2=0
+ $Y2=0
cc_371 N_A_27_101#_c_302_n N_RESET_B_c_945_n 5.91049e-19 $X=1.655 $Y=0.34 $X2=0
+ $Y2=0
cc_372 N_A_27_101#_c_305_n N_RESET_B_c_945_n 0.00377837f $X=2.41 $Y=0.955 $X2=0
+ $Y2=0
cc_373 N_A_27_101#_c_302_n N_RESET_B_c_946_n 8.56593e-19 $X=1.655 $Y=0.34 $X2=0
+ $Y2=0
cc_374 N_A_27_101#_c_304_n N_RESET_B_M1032_g 0.00152111f $X=1.74 $Y=0.87 $X2=0
+ $Y2=0
cc_375 N_A_27_101#_c_305_n N_RESET_B_M1032_g 0.0101313f $X=2.41 $Y=0.955 $X2=0
+ $Y2=0
cc_376 N_A_27_101#_c_360_p N_RESET_B_M1032_g 0.00892444f $X=2.495 $Y=0.87 $X2=0
+ $Y2=0
cc_377 N_A_27_101#_c_447_p N_RESET_B_M1032_g 0.00708932f $X=2.58 $Y=0.362 $X2=0
+ $Y2=0
cc_378 N_A_27_101#_c_307_n N_RESET_B_c_948_n 0.0131446f $X=3.33 $Y=0.362 $X2=0
+ $Y2=0
cc_379 N_A_27_101#_c_447_p N_RESET_B_c_948_n 0.00321157f $X=2.58 $Y=0.362 $X2=0
+ $Y2=0
cc_380 N_A_27_101#_c_309_n N_RESET_B_c_948_n 0.0147033f $X=4.05 $Y=0.362 $X2=0
+ $Y2=0
cc_381 N_A_27_101#_c_311_n N_RESET_B_c_948_n 0.00675701f $X=5.485 $Y=0.89 $X2=0
+ $Y2=0
cc_382 N_A_27_101#_c_452_p N_RESET_B_c_948_n 0.00378523f $X=3.415 $Y=0.362 $X2=0
+ $Y2=0
cc_383 N_A_27_101#_c_323_n N_RESET_B_c_948_n 0.00895246f $X=3.3 $Y=1.135 $X2=0
+ $Y2=0
cc_384 N_A_27_101#_c_309_n N_RESET_B_M1027_g 0.00560683f $X=4.05 $Y=0.362 $X2=0
+ $Y2=0
cc_385 N_A_27_101#_c_311_n N_RESET_B_M1027_g 0.0138538f $X=5.485 $Y=0.89 $X2=0
+ $Y2=0
cc_386 N_A_27_101#_c_376_p N_RESET_B_M1027_g 0.00288071f $X=5.57 $Y=0.805 $X2=0
+ $Y2=0
cc_387 N_A_27_101#_c_311_n N_RESET_B_c_953_n 8.68359e-19 $X=5.485 $Y=0.89 $X2=0
+ $Y2=0
cc_388 N_A_27_101#_M1030_g N_RESET_B_c_997_n 0.0147178f $X=6.185 $Y=2.675 $X2=0
+ $Y2=0
cc_389 N_A_27_101#_c_308_n N_A_573_535#_M1004_d 0.00407654f $X=3.415 $Y=1.14
+ $X2=-0.19 $Y2=-0.245
cc_390 N_A_27_101#_c_332_n N_A_573_535#_c_1172_n 2.23154e-19 $X=6.26 $Y=1.91
+ $X2=0 $Y2=0
cc_391 N_A_27_101#_c_311_n N_A_573_535#_c_1173_n 0.00591979f $X=5.485 $Y=0.89
+ $X2=0 $Y2=0
cc_392 N_A_27_101#_c_376_p N_A_573_535#_c_1173_n 0.0105231f $X=5.57 $Y=0.805
+ $X2=0 $Y2=0
cc_393 N_A_27_101#_c_312_n N_A_573_535#_c_1173_n 0.010391f $X=6.175 $Y=0.34
+ $X2=0 $Y2=0
cc_394 N_A_27_101#_c_313_n N_A_573_535#_c_1173_n 0.00305089f $X=5.655 $Y=0.34
+ $X2=0 $Y2=0
cc_395 N_A_27_101#_c_314_n N_A_573_535#_c_1173_n 0.00105914f $X=6.26 $Y=1.91
+ $X2=0 $Y2=0
cc_396 N_A_27_101#_M1006_g N_A_573_535#_c_1194_n 0.0130061f $X=3.26 $Y=2.885
+ $X2=0 $Y2=0
cc_397 N_A_27_101#_M1006_g N_A_573_535#_c_1180_n 0.00589784f $X=3.26 $Y=2.885
+ $X2=0 $Y2=0
cc_398 N_A_27_101#_M1006_g N_A_573_535#_c_1182_n 0.0041276f $X=3.26 $Y=2.885
+ $X2=0 $Y2=0
cc_399 N_A_27_101#_c_308_n N_A_573_535#_c_1174_n 0.0372409f $X=3.415 $Y=1.14
+ $X2=0 $Y2=0
cc_400 N_A_27_101#_c_309_n N_A_573_535#_c_1174_n 0.0152993f $X=4.05 $Y=0.362
+ $X2=0 $Y2=0
cc_401 N_A_27_101#_c_323_n N_A_573_535#_c_1174_n 0.00138349f $X=3.3 $Y=1.135
+ $X2=0 $Y2=0
cc_402 N_A_27_101#_c_308_n N_A_573_535#_c_1175_n 0.0161091f $X=3.415 $Y=1.14
+ $X2=0 $Y2=0
cc_403 N_A_27_101#_c_320_n N_A_573_535#_c_1175_n 7.18081e-19 $X=3.3 $Y=1.3 $X2=0
+ $Y2=0
cc_404 N_A_27_101#_c_309_n N_A_573_535#_c_1176_n 0.00388046f $X=4.05 $Y=0.362
+ $X2=0 $Y2=0
cc_405 N_A_27_101#_c_311_n N_A_573_535#_c_1176_n 0.101085f $X=5.485 $Y=0.89
+ $X2=0 $Y2=0
cc_406 N_A_27_101#_c_373_p N_A_573_535#_c_1176_n 0.0108192f $X=4.22 $Y=0.89
+ $X2=0 $Y2=0
cc_407 N_A_27_101#_M1030_g N_A_573_535#_c_1185_n 0.0322139f $X=6.185 $Y=2.675
+ $X2=0 $Y2=0
cc_408 N_A_27_101#_c_332_n N_A_573_535#_c_1185_n 0.00944521f $X=6.26 $Y=1.91
+ $X2=0 $Y2=0
cc_409 N_A_27_101#_c_311_n N_A_573_535#_c_1177_n 0.0082984f $X=5.485 $Y=0.89
+ $X2=0 $Y2=0
cc_410 N_A_27_101#_c_316_n N_A_1399_473#_M1024_g 0.00129738f $X=7.01 $Y=0.35
+ $X2=0 $Y2=0
cc_411 N_A_27_101#_c_324_n N_A_1399_473#_M1024_g 0.0198517f $X=7.01 $Y=0.515
+ $X2=0 $Y2=0
cc_412 N_A_27_101#_c_315_n N_A_1252_451#_M1020_d 0.00656171f $X=7.01 $Y=0.35
+ $X2=-0.19 $Y2=-0.245
cc_413 N_A_27_101#_c_314_n N_A_1252_451#_c_1423_n 0.0326732f $X=6.26 $Y=1.91
+ $X2=0 $Y2=0
cc_414 N_A_27_101#_c_315_n N_A_1252_451#_c_1423_n 0.0190645f $X=7.01 $Y=0.35
+ $X2=0 $Y2=0
cc_415 N_A_27_101#_c_324_n N_A_1252_451#_c_1423_n 0.0123382f $X=7.01 $Y=0.515
+ $X2=0 $Y2=0
cc_416 N_A_27_101#_M1030_g N_A_1252_451#_c_1424_n 0.0026978f $X=6.185 $Y=2.675
+ $X2=0 $Y2=0
cc_417 N_A_27_101#_c_314_n N_A_1252_451#_c_1424_n 0.0602416f $X=6.26 $Y=1.91
+ $X2=0 $Y2=0
cc_418 N_A_27_101#_c_332_n N_A_1252_451#_c_1424_n 0.00200461f $X=6.26 $Y=1.91
+ $X2=0 $Y2=0
cc_419 N_A_27_101#_c_315_n N_A_1252_451#_c_1425_n 0.0104794f $X=7.01 $Y=0.35
+ $X2=0 $Y2=0
cc_420 N_A_27_101#_c_316_n N_A_1252_451#_c_1425_n 0.00311395f $X=7.01 $Y=0.35
+ $X2=0 $Y2=0
cc_421 N_A_27_101#_c_324_n N_A_1252_451#_c_1425_n 0.00960376f $X=7.01 $Y=0.515
+ $X2=0 $Y2=0
cc_422 N_A_27_101#_c_314_n N_A_1252_451#_c_1436_n 0.00311214f $X=6.26 $Y=1.91
+ $X2=0 $Y2=0
cc_423 N_A_27_101#_c_332_n N_A_1252_451#_c_1436_n 0.00282952f $X=6.26 $Y=1.91
+ $X2=0 $Y2=0
cc_424 N_A_27_101#_c_314_n N_A_1252_451#_c_1427_n 0.0138012f $X=6.26 $Y=1.91
+ $X2=0 $Y2=0
cc_425 N_A_27_101#_c_329_n N_VPWR_M1003_d 0.00177916f $X=0.665 $Y=2.385
+ $X2=-0.19 $Y2=-0.245
cc_426 N_A_27_101#_M1019_g N_VPWR_c_1649_n 0.0116025f $X=0.905 $Y=2.64 $X2=0
+ $Y2=0
cc_427 N_A_27_101#_c_329_n N_VPWR_c_1649_n 0.0162291f $X=0.665 $Y=2.385 $X2=0
+ $Y2=0
cc_428 N_A_27_101#_c_333_n N_VPWR_c_1649_n 0.0127436f $X=0.26 $Y=2.465 $X2=0
+ $Y2=0
cc_429 N_A_27_101#_M1006_g N_VPWR_c_1657_n 0.00363059f $X=3.26 $Y=2.885 $X2=0
+ $Y2=0
cc_430 N_A_27_101#_c_333_n N_VPWR_c_1661_n 0.0110559f $X=0.26 $Y=2.465 $X2=0
+ $Y2=0
cc_431 N_A_27_101#_M1019_g N_VPWR_c_1662_n 0.00383152f $X=0.905 $Y=2.64 $X2=0
+ $Y2=0
cc_432 N_A_27_101#_M1030_g N_VPWR_c_1668_n 0.00357877f $X=6.185 $Y=2.675 $X2=0
+ $Y2=0
cc_433 N_A_27_101#_M1019_g N_VPWR_c_1648_n 0.00762539f $X=0.905 $Y=2.64 $X2=0
+ $Y2=0
cc_434 N_A_27_101#_M1006_g N_VPWR_c_1648_n 0.00538836f $X=3.26 $Y=2.885 $X2=0
+ $Y2=0
cc_435 N_A_27_101#_M1030_g N_VPWR_c_1648_n 0.00570473f $X=6.185 $Y=2.675 $X2=0
+ $Y2=0
cc_436 N_A_27_101#_c_329_n N_VPWR_c_1648_n 0.00588972f $X=0.665 $Y=2.385 $X2=0
+ $Y2=0
cc_437 N_A_27_101#_c_333_n N_VPWR_c_1648_n 0.00946638f $X=0.26 $Y=2.465 $X2=0
+ $Y2=0
cc_438 N_A_27_101#_M1019_g N_A_318_535#_c_1807_n 0.00256076f $X=0.905 $Y=2.64
+ $X2=0 $Y2=0
cc_439 N_A_27_101#_M1006_g N_A_318_535#_c_1811_n 0.0051991f $X=3.26 $Y=2.885
+ $X2=0 $Y2=0
cc_440 N_A_27_101#_M1006_g N_A_318_535#_c_1805_n 0.00309009f $X=3.26 $Y=2.885
+ $X2=0 $Y2=0
cc_441 N_A_27_101#_c_305_n N_A_318_535#_c_1805_n 0.00482842f $X=2.41 $Y=0.955
+ $X2=0 $Y2=0
cc_442 N_A_27_101#_c_308_n N_A_318_535#_c_1805_n 0.0234389f $X=3.415 $Y=1.14
+ $X2=0 $Y2=0
cc_443 N_A_27_101#_c_320_n N_A_318_535#_c_1805_n 0.00388386f $X=3.3 $Y=1.3 $X2=0
+ $Y2=0
cc_444 N_A_27_101#_c_323_n N_A_318_535#_c_1805_n 8.39165e-19 $X=3.3 $Y=1.135
+ $X2=0 $Y2=0
cc_445 N_A_27_101#_M1006_g N_A_318_535#_c_1812_n 0.017995f $X=3.26 $Y=2.885
+ $X2=0 $Y2=0
cc_446 N_A_27_101#_c_305_n N_A_318_535#_c_1823_n 0.0071682f $X=2.41 $Y=0.955
+ $X2=0 $Y2=0
cc_447 N_A_27_101#_c_360_p N_A_318_535#_c_1823_n 0.0148128f $X=2.495 $Y=0.87
+ $X2=0 $Y2=0
cc_448 N_A_27_101#_c_307_n N_A_318_535#_c_1823_n 0.0247504f $X=3.33 $Y=0.362
+ $X2=0 $Y2=0
cc_449 N_A_27_101#_c_308_n N_A_318_535#_c_1823_n 0.00141755f $X=3.415 $Y=1.14
+ $X2=0 $Y2=0
cc_450 N_A_27_101#_c_320_n N_A_318_535#_c_1823_n 5.41963e-19 $X=3.3 $Y=1.3 $X2=0
+ $Y2=0
cc_451 N_A_27_101#_M1006_g N_A_318_535#_c_1806_n 0.00608881f $X=3.26 $Y=2.885
+ $X2=0 $Y2=0
cc_452 N_A_27_101#_c_308_n N_A_318_535#_c_1806_n 0.00679537f $X=3.415 $Y=1.14
+ $X2=0 $Y2=0
cc_453 N_A_27_101#_c_320_n N_A_318_535#_c_1806_n 0.00122451f $X=3.3 $Y=1.3 $X2=0
+ $Y2=0
cc_454 N_A_27_101#_c_311_n N_VGND_M1027_d 0.00929582f $X=5.485 $Y=0.89 $X2=0
+ $Y2=0
cc_455 N_A_27_101#_c_376_p N_VGND_M1027_d 0.00466975f $X=5.57 $Y=0.805 $X2=0
+ $Y2=0
cc_456 N_A_27_101#_c_313_n N_VGND_M1027_d 0.00109436f $X=5.655 $Y=0.34 $X2=0
+ $Y2=0
cc_457 N_A_27_101#_c_300_n N_VGND_c_1913_n 0.00542902f $X=0.665 $Y=1.185 $X2=0
+ $Y2=0
cc_458 N_A_27_101#_c_303_n N_VGND_c_1913_n 0.0146372f $X=1.125 $Y=0.34 $X2=0
+ $Y2=0
cc_459 N_A_27_101#_c_317_n N_VGND_c_1913_n 0.00899376f $X=0.895 $Y=1.185 $X2=0
+ $Y2=0
cc_460 N_A_27_101#_c_318_n N_VGND_c_1913_n 0.0202813f $X=0.895 $Y=1.1 $X2=0
+ $Y2=0
cc_461 N_A_27_101#_c_322_n N_VGND_c_1913_n 0.00169404f $X=0.972 $Y=1.035 $X2=0
+ $Y2=0
cc_462 N_A_27_101#_c_302_n N_VGND_c_1914_n 0.014674f $X=1.655 $Y=0.34 $X2=0
+ $Y2=0
cc_463 N_A_27_101#_c_304_n N_VGND_c_1914_n 0.0208647f $X=1.74 $Y=0.87 $X2=0
+ $Y2=0
cc_464 N_A_27_101#_c_305_n N_VGND_c_1914_n 0.0187022f $X=2.41 $Y=0.955 $X2=0
+ $Y2=0
cc_465 N_A_27_101#_c_447_p N_VGND_c_1914_n 0.014366f $X=2.58 $Y=0.362 $X2=0
+ $Y2=0
cc_466 N_A_27_101#_c_311_n N_VGND_c_1915_n 0.021361f $X=5.485 $Y=0.89 $X2=0
+ $Y2=0
cc_467 N_A_27_101#_c_376_p N_VGND_c_1915_n 0.0157636f $X=5.57 $Y=0.805 $X2=0
+ $Y2=0
cc_468 N_A_27_101#_c_313_n N_VGND_c_1915_n 0.0144694f $X=5.655 $Y=0.34 $X2=0
+ $Y2=0
cc_469 N_A_27_101#_c_315_n N_VGND_c_1916_n 0.00898475f $X=7.01 $Y=0.35 $X2=0
+ $Y2=0
cc_470 N_A_27_101#_c_316_n N_VGND_c_1916_n 0.00505103f $X=7.01 $Y=0.35 $X2=0
+ $Y2=0
cc_471 N_A_27_101#_c_324_n N_VGND_c_1916_n 0.00171223f $X=7.01 $Y=0.515 $X2=0
+ $Y2=0
cc_472 N_A_27_101#_c_307_n N_VGND_c_1920_n 0.0490306f $X=3.33 $Y=0.362 $X2=0
+ $Y2=0
cc_473 N_A_27_101#_c_447_p N_VGND_c_1920_n 0.0115566f $X=2.58 $Y=0.362 $X2=0
+ $Y2=0
cc_474 N_A_27_101#_c_309_n N_VGND_c_1920_n 0.0475775f $X=4.05 $Y=0.362 $X2=0
+ $Y2=0
cc_475 N_A_27_101#_c_452_p N_VGND_c_1920_n 0.0115893f $X=3.415 $Y=0.362 $X2=0
+ $Y2=0
cc_476 N_A_27_101#_c_312_n N_VGND_c_1922_n 0.0331074f $X=6.175 $Y=0.34 $X2=0
+ $Y2=0
cc_477 N_A_27_101#_c_313_n N_VGND_c_1922_n 0.0121159f $X=5.655 $Y=0.34 $X2=0
+ $Y2=0
cc_478 N_A_27_101#_c_315_n N_VGND_c_1922_n 0.0519785f $X=7.01 $Y=0.35 $X2=0
+ $Y2=0
cc_479 N_A_27_101#_c_316_n N_VGND_c_1922_n 0.00647615f $X=7.01 $Y=0.35 $X2=0
+ $Y2=0
cc_480 N_A_27_101#_c_321_n N_VGND_c_1922_n 0.0124467f $X=6.265 $Y=0.345 $X2=0
+ $Y2=0
cc_481 N_A_27_101#_c_299_n N_VGND_c_1924_n 0.00647246f $X=0.26 $Y=0.715 $X2=0
+ $Y2=0
cc_482 N_A_27_101#_c_302_n N_VGND_c_1925_n 0.0454974f $X=1.655 $Y=0.34 $X2=0
+ $Y2=0
cc_483 N_A_27_101#_c_303_n N_VGND_c_1925_n 0.0121867f $X=1.125 $Y=0.34 $X2=0
+ $Y2=0
cc_484 N_A_27_101#_c_322_n N_VGND_c_1925_n 7.16913e-19 $X=0.972 $Y=1.035 $X2=0
+ $Y2=0
cc_485 N_A_27_101#_c_299_n N_VGND_c_1931_n 0.00949401f $X=0.26 $Y=0.715 $X2=0
+ $Y2=0
cc_486 N_A_27_101#_c_302_n N_VGND_c_1931_n 0.0254889f $X=1.655 $Y=0.34 $X2=0
+ $Y2=0
cc_487 N_A_27_101#_c_303_n N_VGND_c_1931_n 0.00660921f $X=1.125 $Y=0.34 $X2=0
+ $Y2=0
cc_488 N_A_27_101#_c_307_n N_VGND_c_1931_n 0.0253444f $X=3.33 $Y=0.362 $X2=0
+ $Y2=0
cc_489 N_A_27_101#_c_447_p N_VGND_c_1931_n 0.00579705f $X=2.58 $Y=0.362 $X2=0
+ $Y2=0
cc_490 N_A_27_101#_c_309_n N_VGND_c_1931_n 0.0244249f $X=4.05 $Y=0.362 $X2=0
+ $Y2=0
cc_491 N_A_27_101#_c_311_n N_VGND_c_1931_n 0.0325597f $X=5.485 $Y=0.89 $X2=0
+ $Y2=0
cc_492 N_A_27_101#_c_312_n N_VGND_c_1931_n 0.01902f $X=6.175 $Y=0.34 $X2=0 $Y2=0
cc_493 N_A_27_101#_c_313_n N_VGND_c_1931_n 0.00645908f $X=5.655 $Y=0.34 $X2=0
+ $Y2=0
cc_494 N_A_27_101#_c_315_n N_VGND_c_1931_n 0.0292708f $X=7.01 $Y=0.35 $X2=0
+ $Y2=0
cc_495 N_A_27_101#_c_316_n N_VGND_c_1931_n 0.00968077f $X=7.01 $Y=0.35 $X2=0
+ $Y2=0
cc_496 N_A_27_101#_c_452_p N_VGND_c_1931_n 0.00583135f $X=3.415 $Y=0.362 $X2=0
+ $Y2=0
cc_497 N_A_27_101#_c_321_n N_VGND_c_1931_n 0.00640315f $X=6.265 $Y=0.345 $X2=0
+ $Y2=0
cc_498 N_A_27_101#_c_305_n A_483_78# 0.00135969f $X=2.41 $Y=0.955 $X2=-0.19
+ $Y2=-0.245
cc_499 N_A_27_101#_c_360_p A_483_78# 0.00407171f $X=2.495 $Y=0.87 $X2=-0.19
+ $Y2=-0.245
cc_500 N_A_27_101#_c_307_n A_483_78# 0.00329747f $X=3.33 $Y=0.362 $X2=-0.19
+ $Y2=-0.245
cc_501 N_A_27_101#_c_373_p A_811_119# 0.00105415f $X=4.22 $Y=0.89 $X2=-0.19
+ $Y2=-0.245
cc_502 N_A_27_101#_c_311_n A_883_119# 0.00480767f $X=5.485 $Y=0.89 $X2=-0.19
+ $Y2=-0.245
cc_503 N_D_M1026_g N_A_196_464#_M1010_g 0.026317f $X=2.36 $Y=2.885 $X2=0 $Y2=0
cc_504 D N_A_196_464#_c_635_n 0.00955906f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_505 D N_A_196_464#_c_649_n 0.00161826f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_506 N_D_M1026_g N_A_196_464#_c_650_n 0.0109305f $X=2.36 $Y=2.885 $X2=0 $Y2=0
cc_507 N_D_c_579_n N_A_196_464#_c_650_n 0.00190326f $X=2.215 $Y=1.88 $X2=0 $Y2=0
cc_508 D N_A_196_464#_c_650_n 0.0207715f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_509 N_D_M1026_g N_A_196_464#_c_652_n 0.00118604f $X=2.36 $Y=2.885 $X2=0 $Y2=0
cc_510 N_D_c_573_n N_A_196_464#_c_652_n 7.26496e-19 $X=2.775 $Y=1.285 $X2=0
+ $Y2=0
cc_511 N_D_M1026_g N_A_196_464#_c_653_n 0.021261f $X=2.36 $Y=2.885 $X2=0 $Y2=0
cc_512 N_D_c_573_n N_A_196_464#_c_653_n 0.00440472f $X=2.775 $Y=1.285 $X2=0
+ $Y2=0
cc_513 N_D_c_573_n N_A_196_464#_c_636_n 0.00671022f $X=2.775 $Y=1.285 $X2=0
+ $Y2=0
cc_514 N_D_c_579_n N_A_196_464#_c_636_n 0.00145109f $X=2.215 $Y=1.88 $X2=0 $Y2=0
cc_515 D N_A_196_464#_c_636_n 0.0197298f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_516 N_D_c_577_n N_A_196_464#_c_636_n 0.00385571f $X=2.16 $Y=1.375 $X2=0 $Y2=0
cc_517 D N_A_196_464#_c_637_n 6.74348e-19 $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_518 D N_A_196_464#_c_640_n 0.0239134f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_519 N_D_c_577_n N_A_196_464#_c_640_n 0.00179085f $X=2.16 $Y=1.375 $X2=0 $Y2=0
cc_520 N_D_M1026_g N_RESET_B_c_944_n 0.00424012f $X=2.36 $Y=2.885 $X2=0 $Y2=0
cc_521 N_D_c_574_n N_RESET_B_c_944_n 0.0365612f $X=2.395 $Y=1.285 $X2=0 $Y2=0
cc_522 D N_RESET_B_c_944_n 0.00173923f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_523 N_D_c_574_n N_RESET_B_M1032_g 0.00708704f $X=2.395 $Y=1.285 $X2=0 $Y2=0
cc_524 N_D_M1002_g N_RESET_B_M1032_g 0.013707f $X=2.85 $Y=0.805 $X2=0 $Y2=0
cc_525 N_D_M1002_g N_RESET_B_c_948_n 0.00879187f $X=2.85 $Y=0.805 $X2=0 $Y2=0
cc_526 N_D_M1026_g N_RESET_B_c_961_n 0.0329467f $X=2.36 $Y=2.885 $X2=0 $Y2=0
cc_527 N_D_c_579_n N_RESET_B_c_961_n 5.63184e-19 $X=2.215 $Y=1.88 $X2=0 $Y2=0
cc_528 N_D_M1026_g N_VPWR_c_1650_n 0.00898125f $X=2.36 $Y=2.885 $X2=0 $Y2=0
cc_529 N_D_M1026_g N_VPWR_c_1657_n 0.00365202f $X=2.36 $Y=2.885 $X2=0 $Y2=0
cc_530 N_D_M1026_g N_VPWR_c_1648_n 0.00442612f $X=2.36 $Y=2.885 $X2=0 $Y2=0
cc_531 N_D_M1026_g N_A_318_535#_c_1808_n 0.011869f $X=2.36 $Y=2.885 $X2=0 $Y2=0
cc_532 N_D_M1026_g N_A_318_535#_c_1810_n 0.00115233f $X=2.36 $Y=2.885 $X2=0
+ $Y2=0
cc_533 N_D_c_573_n N_A_318_535#_c_1805_n 0.00773242f $X=2.775 $Y=1.285 $X2=0
+ $Y2=0
cc_534 N_D_M1002_g N_A_318_535#_c_1805_n 0.0108365f $X=2.85 $Y=0.805 $X2=0 $Y2=0
cc_535 D N_A_318_535#_c_1805_n 0.0120641f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_536 N_D_c_577_n N_A_318_535#_c_1805_n 0.00414256f $X=2.16 $Y=1.375 $X2=0
+ $Y2=0
cc_537 N_D_c_579_n N_A_318_535#_c_1812_n 0.00441067f $X=2.215 $Y=1.88 $X2=0
+ $Y2=0
cc_538 N_D_M1002_g N_A_318_535#_c_1823_n 0.00834552f $X=2.85 $Y=0.805 $X2=0
+ $Y2=0
cc_539 N_D_c_573_n N_A_318_535#_c_1806_n 2.08955e-19 $X=2.775 $Y=1.285 $X2=0
+ $Y2=0
cc_540 D N_A_318_535#_c_1806_n 0.00418027f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_541 N_D_c_577_n N_A_318_535#_c_1806_n 0.00236432f $X=2.16 $Y=1.375 $X2=0
+ $Y2=0
cc_542 N_A_196_464#_c_630_n N_A_709_411#_c_863_n 6.08083e-19 $X=3.98 $Y=1.205
+ $X2=0 $Y2=0
cc_543 N_A_196_464#_c_630_n N_A_709_411#_c_864_n 0.0175611f $X=3.98 $Y=1.205
+ $X2=0 $Y2=0
cc_544 N_A_196_464#_c_643_n N_A_709_411#_c_864_n 9.33695e-19 $X=3.84 $Y=1.65
+ $X2=0 $Y2=0
cc_545 N_A_196_464#_c_630_n N_A_709_411#_c_857_n 0.0149732f $X=3.98 $Y=1.205
+ $X2=0 $Y2=0
cc_546 N_A_196_464#_c_638_n N_A_709_411#_c_857_n 0.0039633f $X=6.815 $Y=1.665
+ $X2=0 $Y2=0
cc_547 N_A_196_464#_c_643_n N_A_709_411#_c_857_n 0.0011533f $X=3.84 $Y=1.65
+ $X2=0 $Y2=0
cc_548 N_A_196_464#_c_630_n N_A_709_411#_M1014_g 0.0127927f $X=3.98 $Y=1.205
+ $X2=0 $Y2=0
cc_549 N_A_196_464#_M1023_g N_A_709_411#_M1014_g 0.0548041f $X=3.98 $Y=0.805
+ $X2=0 $Y2=0
cc_550 N_A_196_464#_c_630_n N_A_709_411#_c_859_n 6.20601e-19 $X=3.98 $Y=1.205
+ $X2=0 $Y2=0
cc_551 N_A_196_464#_c_638_n N_A_709_411#_c_859_n 0.0453997f $X=6.815 $Y=1.665
+ $X2=0 $Y2=0
cc_552 N_A_196_464#_c_639_n N_A_709_411#_c_859_n 3.74974e-19 $X=3.745 $Y=1.665
+ $X2=0 $Y2=0
cc_553 N_A_196_464#_c_643_n N_A_709_411#_c_859_n 0.00536445f $X=3.84 $Y=1.65
+ $X2=0 $Y2=0
cc_554 N_A_196_464#_M1020_g N_A_709_411#_c_860_n 0.00320195f $X=6.3 $Y=0.635
+ $X2=0 $Y2=0
cc_555 N_A_196_464#_c_634_n N_A_709_411#_c_861_n 2.74305e-19 $X=6.375 $Y=1.46
+ $X2=0 $Y2=0
cc_556 N_A_196_464#_c_638_n N_A_709_411#_c_861_n 0.0122773f $X=6.815 $Y=1.665
+ $X2=0 $Y2=0
cc_557 N_A_196_464#_c_638_n N_A_709_411#_c_869_n 0.0126928f $X=6.815 $Y=1.665
+ $X2=0 $Y2=0
cc_558 N_A_196_464#_c_635_n N_RESET_B_c_944_n 0.0111949f $X=1.39 $Y=0.76 $X2=0
+ $Y2=0
cc_559 N_A_196_464#_c_649_n N_RESET_B_c_944_n 0.00604944f $X=1.385 $Y=2.085
+ $X2=0 $Y2=0
cc_560 N_A_196_464#_c_650_n N_RESET_B_c_944_n 0.0033546f $X=2.645 $Y=2.17 $X2=0
+ $Y2=0
cc_561 N_A_196_464#_c_640_n N_RESET_B_c_944_n 0.0183308f $X=1.68 $Y=1.665 $X2=0
+ $Y2=0
cc_562 N_A_196_464#_c_648_n N_RESET_B_M1001_g 0.00500104f $X=1.12 $Y=2.465 $X2=0
+ $Y2=0
cc_563 N_A_196_464#_M1023_g N_RESET_B_c_948_n 0.00882699f $X=3.98 $Y=0.805 $X2=0
+ $Y2=0
cc_564 N_A_196_464#_c_638_n N_RESET_B_c_950_n 0.00204699f $X=6.815 $Y=1.665
+ $X2=0 $Y2=0
cc_565 N_A_196_464#_c_648_n N_RESET_B_c_961_n 3.38616e-19 $X=1.12 $Y=2.465 $X2=0
+ $Y2=0
cc_566 N_A_196_464#_c_650_n N_RESET_B_c_961_n 0.0161089f $X=2.645 $Y=2.17 $X2=0
+ $Y2=0
cc_567 N_A_196_464#_c_640_n N_RESET_B_c_961_n 4.53814e-19 $X=1.68 $Y=1.665 $X2=0
+ $Y2=0
cc_568 N_A_196_464#_c_638_n N_RESET_B_c_964_n 7.72593e-19 $X=6.815 $Y=1.665
+ $X2=0 $Y2=0
cc_569 N_A_196_464#_M1015_g N_RESET_B_c_997_n 0.0124164f $X=6.71 $Y=2.885 $X2=0
+ $Y2=0
cc_570 N_A_196_464#_M1015_g N_RESET_B_c_965_n 0.00451541f $X=6.71 $Y=2.885 $X2=0
+ $Y2=0
cc_571 N_A_196_464#_M1015_g N_RESET_B_c_966_n 0.00130596f $X=6.71 $Y=2.885 $X2=0
+ $Y2=0
cc_572 N_A_196_464#_c_647_n N_RESET_B_c_966_n 8.09863e-19 $X=6.88 $Y=2.125 $X2=0
+ $Y2=0
cc_573 N_A_196_464#_c_642_n N_RESET_B_c_966_n 0.00786216f $X=6.96 $Y=1.62 $X2=0
+ $Y2=0
cc_574 N_A_196_464#_c_768_p N_RESET_B_c_968_n 9.70772e-19 $X=6.96 $Y=1.665 $X2=0
+ $Y2=0
cc_575 N_A_196_464#_c_641_n N_RESET_B_c_968_n 0.00226324f $X=6.96 $Y=1.62 $X2=0
+ $Y2=0
cc_576 N_A_196_464#_c_642_n N_RESET_B_c_968_n 0.0214316f $X=6.96 $Y=1.62 $X2=0
+ $Y2=0
cc_577 N_A_196_464#_M1015_g N_RESET_B_c_969_n 0.00232458f $X=6.71 $Y=2.885 $X2=0
+ $Y2=0
cc_578 N_A_196_464#_c_647_n N_RESET_B_c_969_n 0.00304716f $X=6.88 $Y=2.125 $X2=0
+ $Y2=0
cc_579 N_A_196_464#_c_768_p N_RESET_B_c_969_n 0.00270119f $X=6.96 $Y=1.665 $X2=0
+ $Y2=0
cc_580 N_A_196_464#_c_642_n N_RESET_B_c_969_n 0.0143639f $X=6.96 $Y=1.62 $X2=0
+ $Y2=0
cc_581 N_A_196_464#_c_638_n N_A_573_535#_c_1172_n 0.00254269f $X=6.815 $Y=1.665
+ $X2=0 $Y2=0
cc_582 N_A_196_464#_M1020_g N_A_573_535#_c_1173_n 0.0112151f $X=6.3 $Y=0.635
+ $X2=0 $Y2=0
cc_583 N_A_196_464#_c_630_n N_A_573_535#_c_1181_n 0.00280649f $X=3.98 $Y=1.205
+ $X2=0 $Y2=0
cc_584 N_A_196_464#_c_638_n N_A_573_535#_c_1181_n 0.00704531f $X=6.815 $Y=1.665
+ $X2=0 $Y2=0
cc_585 N_A_196_464#_c_639_n N_A_573_535#_c_1181_n 0.00433358f $X=3.745 $Y=1.665
+ $X2=0 $Y2=0
cc_586 N_A_196_464#_c_643_n N_A_573_535#_c_1181_n 0.0283867f $X=3.84 $Y=1.65
+ $X2=0 $Y2=0
cc_587 N_A_196_464#_c_636_n N_A_573_535#_c_1182_n 3.30792e-19 $X=3.455 $Y=1.665
+ $X2=0 $Y2=0
cc_588 N_A_196_464#_c_639_n N_A_573_535#_c_1182_n 0.00382208f $X=3.745 $Y=1.665
+ $X2=0 $Y2=0
cc_589 N_A_196_464#_c_643_n N_A_573_535#_c_1182_n 0.0125646f $X=3.84 $Y=1.65
+ $X2=0 $Y2=0
cc_590 N_A_196_464#_M1023_g N_A_573_535#_c_1174_n 0.0038544f $X=3.98 $Y=0.805
+ $X2=0 $Y2=0
cc_591 N_A_196_464#_c_630_n N_A_573_535#_c_1175_n 0.00691092f $X=3.98 $Y=1.205
+ $X2=0 $Y2=0
cc_592 N_A_196_464#_c_638_n N_A_573_535#_c_1175_n 0.00103545f $X=6.815 $Y=1.665
+ $X2=0 $Y2=0
cc_593 N_A_196_464#_c_639_n N_A_573_535#_c_1175_n 0.00182203f $X=3.745 $Y=1.665
+ $X2=0 $Y2=0
cc_594 N_A_196_464#_c_643_n N_A_573_535#_c_1175_n 0.0112939f $X=3.84 $Y=1.65
+ $X2=0 $Y2=0
cc_595 N_A_196_464#_c_630_n N_A_573_535#_c_1176_n 0.00606564f $X=3.98 $Y=1.205
+ $X2=0 $Y2=0
cc_596 N_A_196_464#_M1023_g N_A_573_535#_c_1176_n 0.00634378f $X=3.98 $Y=0.805
+ $X2=0 $Y2=0
cc_597 N_A_196_464#_c_638_n N_A_573_535#_c_1176_n 0.0157258f $X=6.815 $Y=1.665
+ $X2=0 $Y2=0
cc_598 N_A_196_464#_c_643_n N_A_573_535#_c_1176_n 0.00591468f $X=3.84 $Y=1.65
+ $X2=0 $Y2=0
cc_599 N_A_196_464#_c_638_n N_A_573_535#_c_1184_n 0.0304364f $X=6.815 $Y=1.665
+ $X2=0 $Y2=0
cc_600 N_A_196_464#_c_638_n N_A_573_535#_c_1185_n 0.00637153f $X=6.815 $Y=1.665
+ $X2=0 $Y2=0
cc_601 N_A_196_464#_c_638_n N_A_573_535#_c_1186_n 0.0077771f $X=6.815 $Y=1.665
+ $X2=0 $Y2=0
cc_602 N_A_196_464#_c_634_n N_A_573_535#_c_1177_n 0.0112151f $X=6.375 $Y=1.46
+ $X2=0 $Y2=0
cc_603 N_A_196_464#_M1015_g N_A_1399_473#_c_1303_n 0.0527711f $X=6.71 $Y=2.885
+ $X2=0 $Y2=0
cc_604 N_A_196_464#_c_647_n N_A_1399_473#_c_1303_n 0.00723221f $X=6.88 $Y=2.125
+ $X2=0 $Y2=0
cc_605 N_A_196_464#_c_633_n N_A_1399_473#_M1024_g 0.0342592f $X=6.635 $Y=1.46
+ $X2=0 $Y2=0
cc_606 N_A_196_464#_M1015_g N_A_1399_473#_M1024_g 0.00298907f $X=6.71 $Y=2.885
+ $X2=0 $Y2=0
cc_607 N_A_196_464#_c_768_p N_A_1399_473#_M1024_g 0.0010269f $X=6.96 $Y=1.665
+ $X2=0 $Y2=0
cc_608 N_A_196_464#_c_642_n N_A_1399_473#_M1024_g 0.00231326f $X=6.96 $Y=1.62
+ $X2=0 $Y2=0
cc_609 N_A_196_464#_M1020_g N_A_1252_451#_c_1423_n 0.0035611f $X=6.3 $Y=0.635
+ $X2=0 $Y2=0
cc_610 N_A_196_464#_M1020_g N_A_1252_451#_c_1424_n 0.00310851f $X=6.3 $Y=0.635
+ $X2=0 $Y2=0
cc_611 N_A_196_464#_c_633_n N_A_1252_451#_c_1424_n 0.0132584f $X=6.635 $Y=1.46
+ $X2=0 $Y2=0
cc_612 N_A_196_464#_M1015_g N_A_1252_451#_c_1424_n 0.00745171f $X=6.71 $Y=2.885
+ $X2=0 $Y2=0
cc_613 N_A_196_464#_c_647_n N_A_1252_451#_c_1424_n 0.0059388f $X=6.88 $Y=2.125
+ $X2=0 $Y2=0
cc_614 N_A_196_464#_c_638_n N_A_1252_451#_c_1424_n 0.020285f $X=6.815 $Y=1.665
+ $X2=0 $Y2=0
cc_615 N_A_196_464#_c_768_p N_A_1252_451#_c_1424_n 0.00232708f $X=6.96 $Y=1.665
+ $X2=0 $Y2=0
cc_616 N_A_196_464#_c_641_n N_A_1252_451#_c_1424_n 0.00966503f $X=6.96 $Y=1.62
+ $X2=0 $Y2=0
cc_617 N_A_196_464#_c_642_n N_A_1252_451#_c_1424_n 0.0442487f $X=6.96 $Y=1.62
+ $X2=0 $Y2=0
cc_618 N_A_196_464#_c_633_n N_A_1252_451#_c_1425_n 0.00701378f $X=6.635 $Y=1.46
+ $X2=0 $Y2=0
cc_619 N_A_196_464#_c_638_n N_A_1252_451#_c_1425_n 0.00131932f $X=6.815 $Y=1.665
+ $X2=0 $Y2=0
cc_620 N_A_196_464#_c_768_p N_A_1252_451#_c_1425_n 0.00522434f $X=6.96 $Y=1.665
+ $X2=0 $Y2=0
cc_621 N_A_196_464#_c_642_n N_A_1252_451#_c_1425_n 0.0101343f $X=6.96 $Y=1.62
+ $X2=0 $Y2=0
cc_622 N_A_196_464#_M1015_g N_A_1252_451#_c_1436_n 0.00950181f $X=6.71 $Y=2.885
+ $X2=0 $Y2=0
cc_623 N_A_196_464#_M1020_g N_A_1252_451#_c_1427_n 0.00205211f $X=6.3 $Y=0.635
+ $X2=0 $Y2=0
cc_624 N_A_196_464#_c_633_n N_A_1252_451#_c_1427_n 0.00384814f $X=6.635 $Y=1.46
+ $X2=0 $Y2=0
cc_625 N_A_196_464#_c_638_n N_A_1252_451#_c_1427_n 0.00314954f $X=6.815 $Y=1.665
+ $X2=0 $Y2=0
cc_626 N_A_196_464#_c_633_n N_A_1252_451#_c_1428_n 9.43869e-19 $X=6.635 $Y=1.46
+ $X2=0 $Y2=0
cc_627 N_A_196_464#_c_642_n N_A_1252_451#_c_1428_n 0.00275186f $X=6.96 $Y=1.62
+ $X2=0 $Y2=0
cc_628 N_A_196_464#_c_648_n N_VPWR_c_1649_n 0.0127436f $X=1.12 $Y=2.465 $X2=0
+ $Y2=0
cc_629 N_A_196_464#_M1010_g N_VPWR_c_1650_n 0.00126615f $X=2.79 $Y=2.885 $X2=0
+ $Y2=0
cc_630 N_A_196_464#_M1010_g N_VPWR_c_1657_n 0.00439206f $X=2.79 $Y=2.885 $X2=0
+ $Y2=0
cc_631 N_A_196_464#_c_648_n N_VPWR_c_1662_n 0.0111085f $X=1.12 $Y=2.465 $X2=0
+ $Y2=0
cc_632 N_A_196_464#_M1015_g N_VPWR_c_1668_n 0.00357877f $X=6.71 $Y=2.885 $X2=0
+ $Y2=0
cc_633 N_A_196_464#_M1010_g N_VPWR_c_1648_n 0.00642652f $X=2.79 $Y=2.885 $X2=0
+ $Y2=0
cc_634 N_A_196_464#_M1015_g N_VPWR_c_1648_n 0.0055095f $X=6.71 $Y=2.885 $X2=0
+ $Y2=0
cc_635 N_A_196_464#_c_648_n N_VPWR_c_1648_n 0.00948794f $X=1.12 $Y=2.465 $X2=0
+ $Y2=0
cc_636 N_A_196_464#_c_648_n N_A_318_535#_c_1807_n 0.0220886f $X=1.12 $Y=2.465
+ $X2=0 $Y2=0
cc_637 N_A_196_464#_c_650_n N_A_318_535#_c_1808_n 0.0479501f $X=2.645 $Y=2.17
+ $X2=0 $Y2=0
cc_638 N_A_196_464#_c_648_n N_A_318_535#_c_1809_n 0.0108414f $X=1.12 $Y=2.465
+ $X2=0 $Y2=0
cc_639 N_A_196_464#_c_650_n N_A_318_535#_c_1809_n 0.0210335f $X=2.645 $Y=2.17
+ $X2=0 $Y2=0
cc_640 N_A_196_464#_M1010_g N_A_318_535#_c_1810_n 0.0021353f $X=2.79 $Y=2.885
+ $X2=0 $Y2=0
cc_641 N_A_196_464#_M1010_g N_A_318_535#_c_1811_n 0.0124018f $X=2.79 $Y=2.885
+ $X2=0 $Y2=0
cc_642 N_A_196_464#_c_652_n N_A_318_535#_c_1811_n 0.0148087f $X=2.81 $Y=2.09
+ $X2=0 $Y2=0
cc_643 N_A_196_464#_c_653_n N_A_318_535#_c_1811_n 0.0030457f $X=2.81 $Y=2.09
+ $X2=0 $Y2=0
cc_644 N_A_196_464#_c_636_n N_A_318_535#_c_1805_n 0.00242771f $X=3.455 $Y=1.665
+ $X2=0 $Y2=0
cc_645 N_A_196_464#_c_639_n N_A_318_535#_c_1805_n 2.69345e-19 $X=3.745 $Y=1.665
+ $X2=0 $Y2=0
cc_646 N_A_196_464#_c_643_n N_A_318_535#_c_1805_n 3.10974e-19 $X=3.84 $Y=1.65
+ $X2=0 $Y2=0
cc_647 N_A_196_464#_M1010_g N_A_318_535#_c_1812_n 0.00339521f $X=2.79 $Y=2.885
+ $X2=0 $Y2=0
cc_648 N_A_196_464#_c_630_n N_A_318_535#_c_1812_n 3.43548e-19 $X=3.98 $Y=1.205
+ $X2=0 $Y2=0
cc_649 N_A_196_464#_c_652_n N_A_318_535#_c_1812_n 0.0243553f $X=2.81 $Y=2.09
+ $X2=0 $Y2=0
cc_650 N_A_196_464#_c_653_n N_A_318_535#_c_1812_n 0.00200461f $X=2.81 $Y=2.09
+ $X2=0 $Y2=0
cc_651 N_A_196_464#_c_636_n N_A_318_535#_c_1812_n 0.00447606f $X=3.455 $Y=1.665
+ $X2=0 $Y2=0
cc_652 N_A_196_464#_c_639_n N_A_318_535#_c_1812_n 0.00142684f $X=3.745 $Y=1.665
+ $X2=0 $Y2=0
cc_653 N_A_196_464#_c_643_n N_A_318_535#_c_1812_n 0.00103366f $X=3.84 $Y=1.65
+ $X2=0 $Y2=0
cc_654 N_A_196_464#_c_650_n N_A_318_535#_c_1813_n 0.0138396f $X=2.645 $Y=2.17
+ $X2=0 $Y2=0
cc_655 N_A_196_464#_c_652_n N_A_318_535#_c_1813_n 0.00454495f $X=2.81 $Y=2.09
+ $X2=0 $Y2=0
cc_656 N_A_196_464#_c_653_n N_A_318_535#_c_1813_n 4.22294e-19 $X=2.81 $Y=2.09
+ $X2=0 $Y2=0
cc_657 N_A_196_464#_c_652_n N_A_318_535#_c_1806_n 0.00699853f $X=2.81 $Y=2.09
+ $X2=0 $Y2=0
cc_658 N_A_196_464#_c_653_n N_A_318_535#_c_1806_n 0.00247568f $X=2.81 $Y=2.09
+ $X2=0 $Y2=0
cc_659 N_A_196_464#_c_636_n N_A_318_535#_c_1806_n 0.0249352f $X=3.455 $Y=1.665
+ $X2=0 $Y2=0
cc_660 N_A_196_464#_c_643_n N_A_318_535#_c_1806_n 0.0120563f $X=3.84 $Y=1.65
+ $X2=0 $Y2=0
cc_661 N_A_196_464#_M1020_g N_VGND_c_1922_n 0.00308034f $X=6.3 $Y=0.635 $X2=0
+ $Y2=0
cc_662 N_A_196_464#_M1020_g N_VGND_c_1931_n 0.00489791f $X=6.3 $Y=0.635 $X2=0
+ $Y2=0
cc_663 N_A_709_411#_M1014_g N_RESET_B_c_948_n 0.0100117f $X=4.34 $Y=0.805 $X2=0
+ $Y2=0
cc_664 N_A_709_411#_M1008_g N_RESET_B_c_957_n 0.0173854f $X=3.62 $Y=2.885 $X2=0
+ $Y2=0
cc_665 N_A_709_411#_c_863_n N_RESET_B_c_957_n 0.0237208f $X=4.215 $Y=2.13 $X2=0
+ $Y2=0
cc_666 N_A_709_411#_M1014_g N_RESET_B_M1027_g 0.023833f $X=4.34 $Y=0.805 $X2=0
+ $Y2=0
cc_667 N_A_709_411#_c_857_n N_RESET_B_c_950_n 0.0191032f $X=4.29 $Y=1.745 $X2=0
+ $Y2=0
cc_668 N_A_709_411#_c_866_n N_RESET_B_c_950_n 0.0107195f $X=4.29 $Y=2.055 $X2=0
+ $Y2=0
cc_669 N_A_709_411#_M1014_g N_RESET_B_c_950_n 0.00596865f $X=4.34 $Y=0.805 $X2=0
+ $Y2=0
cc_670 N_A_709_411#_c_859_n N_RESET_B_c_950_n 0.00988873f $X=5.825 $Y=1.585
+ $X2=0 $Y2=0
cc_671 N_A_709_411#_c_859_n N_RESET_B_c_964_n 4.14947e-19 $X=5.825 $Y=1.585
+ $X2=0 $Y2=0
cc_672 N_A_709_411#_c_869_n N_RESET_B_c_964_n 0.00160357f $X=5.965 $Y=2.405
+ $X2=0 $Y2=0
cc_673 N_A_709_411#_M1007_d N_RESET_B_c_997_n 0.00332344f $X=5.83 $Y=2.255 $X2=0
+ $Y2=0
cc_674 N_A_709_411#_c_909_p N_RESET_B_c_997_n 0.0124413f $X=5.97 $Y=2.57 $X2=0
+ $Y2=0
cc_675 N_A_709_411#_c_857_n N_RESET_B_c_972_n 0.00239442f $X=4.29 $Y=1.745 $X2=0
+ $Y2=0
cc_676 N_A_709_411#_c_859_n N_A_573_535#_c_1172_n 0.0121443f $X=5.825 $Y=1.585
+ $X2=0 $Y2=0
cc_677 N_A_709_411#_c_860_n N_A_573_535#_c_1172_n 0.00278839f $X=5.91 $Y=0.76
+ $X2=0 $Y2=0
cc_678 N_A_709_411#_c_869_n N_A_573_535#_c_1172_n 0.00177893f $X=5.965 $Y=2.405
+ $X2=0 $Y2=0
cc_679 N_A_709_411#_c_860_n N_A_573_535#_c_1173_n 0.00879282f $X=5.91 $Y=0.76
+ $X2=0 $Y2=0
cc_680 N_A_709_411#_M1008_g N_A_573_535#_c_1194_n 0.0061303f $X=3.62 $Y=2.885
+ $X2=0 $Y2=0
cc_681 N_A_709_411#_M1008_g N_A_573_535#_c_1180_n 0.0134312f $X=3.62 $Y=2.885
+ $X2=0 $Y2=0
cc_682 N_A_709_411#_M1008_g N_A_573_535#_c_1181_n 0.00559489f $X=3.62 $Y=2.885
+ $X2=0 $Y2=0
cc_683 N_A_709_411#_c_863_n N_A_573_535#_c_1181_n 0.0155591f $X=4.215 $Y=2.13
+ $X2=0 $Y2=0
cc_684 N_A_709_411#_c_864_n N_A_573_535#_c_1181_n 0.00317485f $X=3.695 $Y=2.13
+ $X2=0 $Y2=0
cc_685 N_A_709_411#_c_864_n N_A_573_535#_c_1182_n 0.00201983f $X=3.695 $Y=2.13
+ $X2=0 $Y2=0
cc_686 N_A_709_411#_c_857_n N_A_573_535#_c_1176_n 0.0053588f $X=4.29 $Y=1.745
+ $X2=0 $Y2=0
cc_687 N_A_709_411#_M1014_g N_A_573_535#_c_1176_n 0.0109358f $X=4.34 $Y=0.805
+ $X2=0 $Y2=0
cc_688 N_A_709_411#_c_859_n N_A_573_535#_c_1176_n 0.09257f $X=5.825 $Y=1.585
+ $X2=0 $Y2=0
cc_689 N_A_709_411#_c_860_n N_A_573_535#_c_1176_n 0.013674f $X=5.91 $Y=0.76
+ $X2=0 $Y2=0
cc_690 N_A_709_411#_M1008_g N_A_573_535#_c_1183_n 0.00365143f $X=3.62 $Y=2.885
+ $X2=0 $Y2=0
cc_691 N_A_709_411#_c_857_n N_A_573_535#_c_1184_n 0.00169303f $X=4.29 $Y=1.745
+ $X2=0 $Y2=0
cc_692 N_A_709_411#_c_859_n N_A_573_535#_c_1184_n 0.0761182f $X=5.825 $Y=1.585
+ $X2=0 $Y2=0
cc_693 N_A_709_411#_c_869_n N_A_573_535#_c_1184_n 0.0160086f $X=5.965 $Y=2.405
+ $X2=0 $Y2=0
cc_694 N_A_709_411#_c_859_n N_A_573_535#_c_1185_n 0.00537573f $X=5.825 $Y=1.585
+ $X2=0 $Y2=0
cc_695 N_A_709_411#_c_869_n N_A_573_535#_c_1185_n 0.00841839f $X=5.965 $Y=2.405
+ $X2=0 $Y2=0
cc_696 N_A_709_411#_c_863_n N_A_573_535#_c_1186_n 0.00700853f $X=4.215 $Y=2.13
+ $X2=0 $Y2=0
cc_697 N_A_709_411#_c_857_n N_A_573_535#_c_1186_n 0.0012583f $X=4.29 $Y=1.745
+ $X2=0 $Y2=0
cc_698 N_A_709_411#_c_866_n N_A_573_535#_c_1186_n 0.0130687f $X=4.29 $Y=2.055
+ $X2=0 $Y2=0
cc_699 N_A_709_411#_c_859_n N_A_573_535#_c_1186_n 0.0128715f $X=5.825 $Y=1.585
+ $X2=0 $Y2=0
cc_700 N_A_709_411#_c_859_n N_A_573_535#_c_1177_n 0.00500217f $X=5.825 $Y=1.585
+ $X2=0 $Y2=0
cc_701 N_A_709_411#_c_869_n N_A_1252_451#_c_1424_n 0.0111402f $X=5.965 $Y=2.405
+ $X2=0 $Y2=0
cc_702 N_A_709_411#_M1008_g N_VPWR_c_1651_n 0.00470014f $X=3.62 $Y=2.885 $X2=0
+ $Y2=0
cc_703 N_A_709_411#_c_863_n N_VPWR_c_1651_n 0.00133849f $X=4.215 $Y=2.13 $X2=0
+ $Y2=0
cc_704 N_A_709_411#_M1008_g N_VPWR_c_1657_n 0.00526043f $X=3.62 $Y=2.885 $X2=0
+ $Y2=0
cc_705 N_A_709_411#_M1007_d N_VPWR_c_1648_n 0.00225186f $X=5.83 $Y=2.255 $X2=0
+ $Y2=0
cc_706 N_A_709_411#_M1008_g N_VPWR_c_1648_n 0.00931664f $X=3.62 $Y=2.885 $X2=0
+ $Y2=0
cc_707 N_A_709_411#_c_864_n N_A_318_535#_c_1812_n 3.16537e-19 $X=3.695 $Y=2.13
+ $X2=0 $Y2=0
cc_708 N_A_709_411#_M1014_g N_VGND_c_1931_n 9.39239e-19 $X=4.34 $Y=0.805 $X2=0
+ $Y2=0
cc_709 N_RESET_B_c_950_n N_A_573_535#_c_1172_n 0.0208795f $X=4.91 $Y=2.235 $X2=0
+ $Y2=0
cc_710 N_RESET_B_c_948_n N_A_573_535#_c_1173_n 0.0107241f $X=4.805 $Y=0.18 $X2=0
+ $Y2=0
cc_711 N_RESET_B_c_950_n N_A_573_535#_M1007_g 0.00603288f $X=4.91 $Y=2.235 $X2=0
+ $Y2=0
cc_712 N_RESET_B_c_964_n N_A_573_535#_M1007_g 0.00322344f $X=5.495 $Y=2.4 $X2=0
+ $Y2=0
cc_713 N_RESET_B_c_997_n N_A_573_535#_M1007_g 0.0152979f $X=6.865 $Y=2.99 $X2=0
+ $Y2=0
cc_714 N_RESET_B_c_957_n N_A_573_535#_c_1180_n 0.00104427f $X=4.15 $Y=2.49 $X2=0
+ $Y2=0
cc_715 N_RESET_B_c_957_n N_A_573_535#_c_1181_n 0.00371437f $X=4.15 $Y=2.49 $X2=0
+ $Y2=0
cc_716 N_RESET_B_c_950_n N_A_573_535#_c_1176_n 0.00667941f $X=4.91 $Y=2.235
+ $X2=0 $Y2=0
cc_717 N_RESET_B_c_953_n N_A_573_535#_c_1176_n 0.00590214f $X=4.895 $Y=1.215
+ $X2=0 $Y2=0
cc_718 N_RESET_B_c_956_n N_A_573_535#_c_1183_n 0.00353822f $X=4.075 $Y=2.565
+ $X2=0 $Y2=0
cc_719 N_RESET_B_c_950_n N_A_573_535#_c_1183_n 4.09025e-19 $X=4.91 $Y=2.235
+ $X2=0 $Y2=0
cc_720 N_RESET_B_c_964_n N_A_573_535#_c_1183_n 0.0266592f $X=5.495 $Y=2.4 $X2=0
+ $Y2=0
cc_721 N_RESET_B_c_972_n N_A_573_535#_c_1183_n 0.0187064f $X=4.595 $Y=2.4 $X2=0
+ $Y2=0
cc_722 N_RESET_B_c_973_n N_A_573_535#_c_1183_n 0.00439651f $X=4.91 $Y=2.4 $X2=0
+ $Y2=0
cc_723 N_RESET_B_c_950_n N_A_573_535#_c_1184_n 0.0137339f $X=4.91 $Y=2.235 $X2=0
+ $Y2=0
cc_724 N_RESET_B_c_964_n N_A_573_535#_c_1184_n 0.076836f $X=5.495 $Y=2.4 $X2=0
+ $Y2=0
cc_725 N_RESET_B_c_972_n N_A_573_535#_c_1184_n 0.0028126f $X=4.595 $Y=2.4 $X2=0
+ $Y2=0
cc_726 N_RESET_B_c_973_n N_A_573_535#_c_1184_n 0.00589537f $X=4.91 $Y=2.4 $X2=0
+ $Y2=0
cc_727 N_RESET_B_c_964_n N_A_573_535#_c_1185_n 0.00901273f $X=5.495 $Y=2.4 $X2=0
+ $Y2=0
cc_728 N_RESET_B_c_950_n N_A_573_535#_c_1186_n 0.00370498f $X=4.91 $Y=2.235
+ $X2=0 $Y2=0
cc_729 N_RESET_B_c_953_n N_A_573_535#_c_1177_n 0.0208795f $X=4.895 $Y=1.215
+ $X2=0 $Y2=0
cc_730 N_RESET_B_c_997_n N_A_1399_473#_M1005_g 0.00386032f $X=6.865 $Y=2.99
+ $X2=0 $Y2=0
cc_731 N_RESET_B_c_965_n N_A_1399_473#_M1005_g 0.0102675f $X=6.95 $Y=2.905 $X2=0
+ $Y2=0
cc_732 N_RESET_B_c_969_n N_A_1399_473#_M1005_g 0.00642348f $X=7.3 $Y=2.45 $X2=0
+ $Y2=0
cc_733 N_RESET_B_c_969_n N_A_1399_473#_c_1303_n 0.00374412f $X=7.3 $Y=2.45 $X2=0
+ $Y2=0
cc_734 N_RESET_B_M1028_g N_A_1399_473#_M1024_g 0.0459766f $X=7.89 $Y=0.835 $X2=0
+ $Y2=0
cc_735 N_RESET_B_c_966_n N_A_1399_473#_M1024_g 0.00424489f $X=7.3 $Y=2.295 $X2=0
+ $Y2=0
cc_736 N_RESET_B_c_967_n N_A_1399_473#_M1024_g 0.0171554f $X=8.035 $Y=1.88 $X2=0
+ $Y2=0
cc_737 N_RESET_B_c_968_n N_A_1399_473#_M1024_g 0.0019885f $X=7.385 $Y=1.88 $X2=0
+ $Y2=0
cc_738 N_RESET_B_c_970_n N_A_1399_473#_M1024_g 0.00741962f $X=8.2 $Y=1.83 $X2=0
+ $Y2=0
cc_739 N_RESET_B_c_971_n N_A_1399_473#_M1024_g 7.91702e-19 $X=8.2 $Y=1.83 $X2=0
+ $Y2=0
cc_740 N_RESET_B_M1031_g N_A_1399_473#_c_1305_n 0.0129099f $X=8.22 $Y=2.885
+ $X2=0 $Y2=0
cc_741 N_RESET_B_c_962_n N_A_1399_473#_c_1305_n 8.6007e-19 $X=8.2 $Y=1.815 $X2=0
+ $Y2=0
cc_742 N_RESET_B_c_963_n N_A_1399_473#_c_1305_n 0.0041174f $X=8.2 $Y=2.335 $X2=0
+ $Y2=0
cc_743 N_RESET_B_c_967_n N_A_1399_473#_c_1305_n 0.0087735f $X=8.035 $Y=1.88
+ $X2=0 $Y2=0
cc_744 N_RESET_B_c_971_n N_A_1399_473#_c_1305_n 0.0213855f $X=8.2 $Y=1.83 $X2=0
+ $Y2=0
cc_745 N_RESET_B_M1031_g N_A_1399_473#_c_1306_n 0.00179158f $X=8.22 $Y=2.885
+ $X2=0 $Y2=0
cc_746 N_RESET_B_M1031_g N_A_1399_473#_c_1308_n 5.23894e-19 $X=8.22 $Y=2.885
+ $X2=0 $Y2=0
cc_747 N_RESET_B_c_963_n N_A_1399_473#_c_1308_n 0.00155188f $X=8.2 $Y=2.335
+ $X2=0 $Y2=0
cc_748 N_RESET_B_c_971_n N_A_1399_473#_c_1308_n 0.0209343f $X=8.2 $Y=1.83 $X2=0
+ $Y2=0
cc_749 N_RESET_B_c_971_n N_A_1399_473#_c_1300_n 0.00659505f $X=8.2 $Y=1.83 $X2=0
+ $Y2=0
cc_750 N_RESET_B_M1031_g N_A_1399_473#_c_1310_n 9.60413e-19 $X=8.22 $Y=2.885
+ $X2=0 $Y2=0
cc_751 N_RESET_B_c_963_n N_A_1399_473#_c_1310_n 8.17366e-19 $X=8.2 $Y=2.335
+ $X2=0 $Y2=0
cc_752 N_RESET_B_c_966_n N_A_1399_473#_c_1310_n 0.0074446f $X=7.3 $Y=2.295 $X2=0
+ $Y2=0
cc_753 N_RESET_B_c_967_n N_A_1399_473#_c_1310_n 0.0197623f $X=8.035 $Y=1.88
+ $X2=0 $Y2=0
cc_754 N_RESET_B_c_969_n N_A_1399_473#_c_1310_n 0.022315f $X=7.3 $Y=2.45 $X2=0
+ $Y2=0
cc_755 N_RESET_B_c_971_n N_A_1399_473#_c_1310_n 0.00445935f $X=8.2 $Y=1.83 $X2=0
+ $Y2=0
cc_756 N_RESET_B_M1031_g N_A_1399_473#_c_1311_n 0.00745113f $X=8.22 $Y=2.885
+ $X2=0 $Y2=0
cc_757 N_RESET_B_c_962_n N_A_1399_473#_c_1311_n 3.20503e-19 $X=8.2 $Y=1.815
+ $X2=0 $Y2=0
cc_758 N_RESET_B_c_963_n N_A_1399_473#_c_1311_n 0.00990269f $X=8.2 $Y=2.335
+ $X2=0 $Y2=0
cc_759 N_RESET_B_c_967_n N_A_1399_473#_c_1311_n 0.00339649f $X=8.035 $Y=1.88
+ $X2=0 $Y2=0
cc_760 N_RESET_B_c_969_n N_A_1399_473#_c_1311_n 0.00336337f $X=7.3 $Y=2.45 $X2=0
+ $Y2=0
cc_761 N_RESET_B_c_971_n N_A_1399_473#_c_1311_n 2.56951e-19 $X=8.2 $Y=1.83 $X2=0
+ $Y2=0
cc_762 N_RESET_B_M1028_g N_A_1399_473#_c_1301_n 0.00193941f $X=7.89 $Y=0.835
+ $X2=0 $Y2=0
cc_763 N_RESET_B_c_966_n N_A_1399_473#_c_1312_n 0.00134937f $X=7.3 $Y=2.295
+ $X2=0 $Y2=0
cc_764 N_RESET_B_c_969_n N_A_1399_473#_c_1312_n 0.0108549f $X=7.3 $Y=2.45 $X2=0
+ $Y2=0
cc_765 N_RESET_B_c_997_n N_A_1252_451#_M1030_d 0.005361f $X=6.865 $Y=2.99 $X2=0
+ $Y2=0
cc_766 N_RESET_B_M1028_g N_A_1252_451#_M1018_g 0.0575628f $X=7.89 $Y=0.835 $X2=0
+ $Y2=0
cc_767 N_RESET_B_c_971_n N_A_1252_451#_c_1416_n 8.1018e-19 $X=8.2 $Y=1.83 $X2=0
+ $Y2=0
cc_768 N_RESET_B_c_962_n N_A_1252_451#_c_1417_n 0.0106029f $X=8.2 $Y=1.815 $X2=0
+ $Y2=0
cc_769 N_RESET_B_M1031_g N_A_1252_451#_M1016_g 0.0223782f $X=8.22 $Y=2.885 $X2=0
+ $Y2=0
cc_770 N_RESET_B_c_963_n N_A_1252_451#_M1016_g 0.0148265f $X=8.2 $Y=2.335 $X2=0
+ $Y2=0
cc_771 N_RESET_B_c_970_n N_A_1252_451#_c_1433_n 0.0148265f $X=8.2 $Y=1.83 $X2=0
+ $Y2=0
cc_772 N_RESET_B_c_971_n N_A_1252_451#_c_1433_n 0.00377092f $X=8.2 $Y=1.83 $X2=0
+ $Y2=0
cc_773 N_RESET_B_c_966_n N_A_1252_451#_c_1424_n 0.00524194f $X=7.3 $Y=2.295
+ $X2=0 $Y2=0
cc_774 N_RESET_B_c_969_n N_A_1252_451#_c_1424_n 0.00859251f $X=7.3 $Y=2.45 $X2=0
+ $Y2=0
cc_775 N_RESET_B_c_968_n N_A_1252_451#_c_1425_n 3.82315e-19 $X=7.385 $Y=1.88
+ $X2=0 $Y2=0
cc_776 N_RESET_B_M1028_g N_A_1252_451#_c_1426_n 0.015237f $X=7.89 $Y=0.835 $X2=0
+ $Y2=0
cc_777 N_RESET_B_c_962_n N_A_1252_451#_c_1426_n 0.00656542f $X=8.2 $Y=1.815
+ $X2=0 $Y2=0
cc_778 N_RESET_B_c_967_n N_A_1252_451#_c_1426_n 0.0355629f $X=8.035 $Y=1.88
+ $X2=0 $Y2=0
cc_779 N_RESET_B_c_971_n N_A_1252_451#_c_1426_n 0.0273374f $X=8.2 $Y=1.83 $X2=0
+ $Y2=0
cc_780 N_RESET_B_c_997_n N_A_1252_451#_c_1436_n 0.0226973f $X=6.865 $Y=2.99
+ $X2=0 $Y2=0
cc_781 N_RESET_B_c_965_n N_A_1252_451#_c_1436_n 0.00986474f $X=6.95 $Y=2.905
+ $X2=0 $Y2=0
cc_782 N_RESET_B_c_969_n N_A_1252_451#_c_1436_n 0.0167195f $X=7.3 $Y=2.45 $X2=0
+ $Y2=0
cc_783 N_RESET_B_M1028_g N_A_1252_451#_c_1428_n 0.00137088f $X=7.89 $Y=0.835
+ $X2=0 $Y2=0
cc_784 N_RESET_B_c_967_n N_A_1252_451#_c_1428_n 4.74919e-19 $X=8.035 $Y=1.88
+ $X2=0 $Y2=0
cc_785 N_RESET_B_c_968_n N_A_1252_451#_c_1428_n 0.0108189f $X=7.385 $Y=1.88
+ $X2=0 $Y2=0
cc_786 N_RESET_B_c_962_n N_A_1252_451#_c_1437_n 7.13715e-19 $X=8.2 $Y=1.815
+ $X2=0 $Y2=0
cc_787 N_RESET_B_c_971_n N_A_1252_451#_c_1437_n 0.0178321f $X=8.2 $Y=1.83 $X2=0
+ $Y2=0
cc_788 N_RESET_B_M1028_g N_A_1252_451#_c_1429_n 0.00510792f $X=7.89 $Y=0.835
+ $X2=0 $Y2=0
cc_789 N_RESET_B_c_962_n N_A_1252_451#_c_1429_n 0.0101271f $X=8.2 $Y=1.815 $X2=0
+ $Y2=0
cc_790 N_RESET_B_c_971_n N_A_1252_451#_c_1429_n 7.33102e-19 $X=8.2 $Y=1.83 $X2=0
+ $Y2=0
cc_791 N_RESET_B_c_964_n N_VPWR_M1007_s 0.0138262f $X=5.495 $Y=2.4 $X2=0 $Y2=0
cc_792 N_RESET_B_c_1125_p N_VPWR_M1007_s 0.0094133f $X=5.58 $Y=2.905 $X2=0 $Y2=0
cc_793 N_RESET_B_c_1126_p N_VPWR_M1007_s 0.00318452f $X=5.665 $Y=2.99 $X2=0
+ $Y2=0
cc_794 N_RESET_B_M1001_g N_VPWR_c_1650_n 0.0100308f $X=1.93 $Y=2.885 $X2=0 $Y2=0
cc_795 N_RESET_B_c_956_n N_VPWR_c_1651_n 0.00321358f $X=4.075 $Y=2.565 $X2=0
+ $Y2=0
cc_796 N_RESET_B_c_964_n N_VPWR_c_1652_n 0.0213599f $X=5.495 $Y=2.4 $X2=0 $Y2=0
cc_797 N_RESET_B_c_1125_p N_VPWR_c_1652_n 0.0127169f $X=5.58 $Y=2.905 $X2=0
+ $Y2=0
cc_798 N_RESET_B_c_1126_p N_VPWR_c_1652_n 0.0142383f $X=5.665 $Y=2.99 $X2=0
+ $Y2=0
cc_799 N_RESET_B_M1031_g N_VPWR_c_1653_n 5.76653e-19 $X=8.22 $Y=2.885 $X2=0
+ $Y2=0
cc_800 N_RESET_B_c_956_n N_VPWR_c_1659_n 0.00585385f $X=4.075 $Y=2.565 $X2=0
+ $Y2=0
cc_801 N_RESET_B_c_972_n N_VPWR_c_1659_n 0.0102605f $X=4.595 $Y=2.4 $X2=0 $Y2=0
cc_802 N_RESET_B_M1001_g N_VPWR_c_1662_n 0.00365202f $X=1.93 $Y=2.885 $X2=0
+ $Y2=0
cc_803 N_RESET_B_M1031_g N_VPWR_c_1663_n 0.00393274f $X=8.22 $Y=2.885 $X2=0
+ $Y2=0
cc_804 N_RESET_B_c_997_n N_VPWR_c_1668_n 0.0763992f $X=6.865 $Y=2.99 $X2=0 $Y2=0
cc_805 N_RESET_B_c_1126_p N_VPWR_c_1668_n 0.0104902f $X=5.665 $Y=2.99 $X2=0
+ $Y2=0
cc_806 N_RESET_B_c_969_n N_VPWR_c_1668_n 0.00249091f $X=7.3 $Y=2.45 $X2=0 $Y2=0
cc_807 N_RESET_B_M1031_g N_VPWR_c_1669_n 0.00891905f $X=8.22 $Y=2.885 $X2=0
+ $Y2=0
cc_808 N_RESET_B_c_997_n N_VPWR_c_1669_n 0.0148585f $X=6.865 $Y=2.99 $X2=0 $Y2=0
cc_809 N_RESET_B_c_965_n N_VPWR_c_1669_n 0.0101479f $X=6.95 $Y=2.905 $X2=0 $Y2=0
cc_810 N_RESET_B_c_969_n N_VPWR_c_1669_n 0.0148266f $X=7.3 $Y=2.45 $X2=0 $Y2=0
cc_811 N_RESET_B_M1001_g N_VPWR_c_1648_n 0.0057985f $X=1.93 $Y=2.885 $X2=0 $Y2=0
cc_812 N_RESET_B_c_956_n N_VPWR_c_1648_n 0.0122148f $X=4.075 $Y=2.565 $X2=0
+ $Y2=0
cc_813 N_RESET_B_M1031_g N_VPWR_c_1648_n 0.00469006f $X=8.22 $Y=2.885 $X2=0
+ $Y2=0
cc_814 N_RESET_B_c_964_n N_VPWR_c_1648_n 0.0236437f $X=5.495 $Y=2.4 $X2=0 $Y2=0
cc_815 N_RESET_B_c_997_n N_VPWR_c_1648_n 0.0494211f $X=6.865 $Y=2.99 $X2=0 $Y2=0
cc_816 N_RESET_B_c_1126_p N_VPWR_c_1648_n 0.00660921f $X=5.665 $Y=2.99 $X2=0
+ $Y2=0
cc_817 N_RESET_B_c_969_n N_VPWR_c_1648_n 0.00483237f $X=7.3 $Y=2.45 $X2=0 $Y2=0
cc_818 N_RESET_B_c_972_n N_VPWR_c_1648_n 0.0130196f $X=4.595 $Y=2.4 $X2=0 $Y2=0
cc_819 N_RESET_B_M1001_g N_A_318_535#_c_1807_n 0.00261315f $X=1.93 $Y=2.885
+ $X2=0 $Y2=0
cc_820 N_RESET_B_M1001_g N_A_318_535#_c_1808_n 0.0132982f $X=1.93 $Y=2.885 $X2=0
+ $Y2=0
cc_821 N_RESET_B_c_961_n N_A_318_535#_c_1808_n 8.72279e-19 $X=1.93 $Y=2.195
+ $X2=0 $Y2=0
cc_822 N_RESET_B_c_961_n N_A_318_535#_c_1809_n 0.00525721f $X=1.93 $Y=2.195
+ $X2=0 $Y2=0
cc_823 N_RESET_B_M1032_g N_A_318_535#_c_1823_n 3.0029e-19 $X=2.34 $Y=0.6 $X2=0
+ $Y2=0
cc_824 N_RESET_B_c_997_n A_1357_535# 0.00174214f $X=6.865 $Y=2.99 $X2=-0.19
+ $Y2=-0.245
cc_825 N_RESET_B_c_965_n A_1357_535# 0.00236267f $X=6.95 $Y=2.905 $X2=-0.19
+ $Y2=-0.245
cc_826 N_RESET_B_c_944_n N_VGND_c_1914_n 0.00118804f $X=1.68 $Y=2.12 $X2=0 $Y2=0
cc_827 N_RESET_B_c_945_n N_VGND_c_1914_n 0.0191562f $X=2.265 $Y=0.18 $X2=0 $Y2=0
cc_828 N_RESET_B_M1032_g N_VGND_c_1914_n 0.00252433f $X=2.34 $Y=0.6 $X2=0 $Y2=0
cc_829 N_RESET_B_c_948_n N_VGND_c_1915_n 0.015666f $X=4.805 $Y=0.18 $X2=0 $Y2=0
cc_830 N_RESET_B_M1028_g N_VGND_c_1916_n 0.00908555f $X=7.89 $Y=0.835 $X2=0
+ $Y2=0
cc_831 N_RESET_B_c_945_n N_VGND_c_1920_n 0.070177f $X=2.265 $Y=0.18 $X2=0 $Y2=0
cc_832 N_RESET_B_c_946_n N_VGND_c_1925_n 0.0112828f $X=1.755 $Y=0.18 $X2=0 $Y2=0
cc_833 N_RESET_B_M1028_g N_VGND_c_1926_n 0.00345209f $X=7.89 $Y=0.835 $X2=0
+ $Y2=0
cc_834 N_RESET_B_c_945_n N_VGND_c_1931_n 0.0123585f $X=2.265 $Y=0.18 $X2=0 $Y2=0
cc_835 N_RESET_B_c_946_n N_VGND_c_1931_n 0.00604509f $X=1.755 $Y=0.18 $X2=0
+ $Y2=0
cc_836 N_RESET_B_c_948_n N_VGND_c_1931_n 0.066104f $X=4.805 $Y=0.18 $X2=0 $Y2=0
cc_837 N_RESET_B_M1028_g N_VGND_c_1931_n 0.00394323f $X=7.89 $Y=0.835 $X2=0
+ $Y2=0
cc_838 N_RESET_B_c_952_n N_VGND_c_1931_n 0.00887976f $X=2.34 $Y=0.18 $X2=0 $Y2=0
cc_839 N_A_573_535#_c_1194_n N_VPWR_c_1651_n 0.0230429f $X=3.415 $Y=2.907 $X2=0
+ $Y2=0
cc_840 N_A_573_535#_c_1180_n N_VPWR_c_1651_n 0.00321192f $X=3.5 $Y=2.765 $X2=0
+ $Y2=0
cc_841 N_A_573_535#_c_1181_n N_VPWR_c_1651_n 0.00841261f $X=4.165 $Y=2.07 $X2=0
+ $Y2=0
cc_842 N_A_573_535#_M1007_g N_VPWR_c_1652_n 0.00422835f $X=5.755 $Y=2.675 $X2=0
+ $Y2=0
cc_843 N_A_573_535#_c_1183_n N_VPWR_c_1652_n 0.0104888f $X=4.29 $Y=2.885 $X2=0
+ $Y2=0
cc_844 N_A_573_535#_c_1194_n N_VPWR_c_1657_n 0.0347383f $X=3.415 $Y=2.907 $X2=0
+ $Y2=0
cc_845 N_A_573_535#_c_1183_n N_VPWR_c_1659_n 0.0162773f $X=4.29 $Y=2.885 $X2=0
+ $Y2=0
cc_846 N_A_573_535#_M1007_g N_VPWR_c_1668_n 0.00357877f $X=5.755 $Y=2.675 $X2=0
+ $Y2=0
cc_847 N_A_573_535#_M1010_d N_VPWR_c_1648_n 0.00261038f $X=2.865 $Y=2.675 $X2=0
+ $Y2=0
cc_848 N_A_573_535#_M1011_d N_VPWR_c_1648_n 0.00235618f $X=4.15 $Y=2.675 $X2=0
+ $Y2=0
cc_849 N_A_573_535#_M1007_g N_VPWR_c_1648_n 0.00684889f $X=5.755 $Y=2.675 $X2=0
+ $Y2=0
cc_850 N_A_573_535#_c_1194_n N_VPWR_c_1648_n 0.0260621f $X=3.415 $Y=2.907 $X2=0
+ $Y2=0
cc_851 N_A_573_535#_c_1183_n N_VPWR_c_1648_n 0.0110608f $X=4.29 $Y=2.885 $X2=0
+ $Y2=0
cc_852 N_A_573_535#_c_1194_n N_A_318_535#_c_1811_n 0.0244877f $X=3.415 $Y=2.907
+ $X2=0 $Y2=0
cc_853 N_A_573_535#_c_1180_n N_A_318_535#_c_1811_n 0.0135843f $X=3.5 $Y=2.765
+ $X2=0 $Y2=0
cc_854 N_A_573_535#_c_1180_n N_A_318_535#_c_1812_n 0.0145893f $X=3.5 $Y=2.765
+ $X2=0 $Y2=0
cc_855 N_A_573_535#_c_1182_n N_A_318_535#_c_1812_n 0.024202f $X=3.585 $Y=2.07
+ $X2=0 $Y2=0
cc_856 N_A_573_535#_c_1194_n A_667_535# 0.00185853f $X=3.415 $Y=2.907 $X2=-0.19
+ $Y2=-0.245
cc_857 N_A_573_535#_c_1180_n A_667_535# 9.85144e-19 $X=3.5 $Y=2.765 $X2=-0.19
+ $Y2=-0.245
cc_858 N_A_573_535#_c_1173_n N_VGND_c_1915_n 0.00233827f $X=5.695 $Y=1.065 $X2=0
+ $Y2=0
cc_859 N_A_573_535#_c_1173_n N_VGND_c_1922_n 0.00308141f $X=5.695 $Y=1.065 $X2=0
+ $Y2=0
cc_860 N_A_573_535#_c_1173_n N_VGND_c_1931_n 0.00502818f $X=5.695 $Y=1.065 $X2=0
+ $Y2=0
cc_861 N_A_1399_473#_c_1299_n N_A_1252_451#_M1018_g 4.27466e-19 $X=9.025 $Y=1.07
+ $X2=0 $Y2=0
cc_862 N_A_1399_473#_c_1301_n N_A_1252_451#_M1018_g 0.0113648f $X=8.465 $Y=0.835
+ $X2=0 $Y2=0
cc_863 N_A_1399_473#_c_1301_n N_A_1252_451#_c_1416_n 0.00464748f $X=8.465
+ $Y=0.835 $X2=0 $Y2=0
cc_864 N_A_1399_473#_c_1306_n N_A_1252_451#_M1016_g 0.00176831f $X=8.435
+ $Y=2.885 $X2=0 $Y2=0
cc_865 N_A_1399_473#_c_1308_n N_A_1252_451#_M1016_g 0.0261737f $X=8.835 $Y=2.26
+ $X2=0 $Y2=0
cc_866 N_A_1399_473#_c_1300_n N_A_1252_451#_M1016_g 0.00347008f $X=9.11 $Y=2.175
+ $X2=0 $Y2=0
cc_867 N_A_1399_473#_c_1300_n N_A_1252_451#_c_1418_n 0.0153142f $X=9.11 $Y=2.175
+ $X2=0 $Y2=0
cc_868 N_A_1399_473#_c_1299_n N_A_1252_451#_M1013_g 0.0010866f $X=9.025 $Y=1.07
+ $X2=0 $Y2=0
cc_869 N_A_1399_473#_c_1300_n N_A_1252_451#_M1013_g 6.99751e-19 $X=9.11 $Y=2.175
+ $X2=0 $Y2=0
cc_870 N_A_1399_473#_c_1300_n N_A_1252_451#_c_1420_n 0.00148264f $X=9.11
+ $Y=2.175 $X2=0 $Y2=0
cc_871 N_A_1399_473#_c_1307_n N_A_1252_451#_M1000_g 9.06288e-19 $X=9.025 $Y=2.26
+ $X2=0 $Y2=0
cc_872 N_A_1399_473#_c_1308_n N_A_1252_451#_M1000_g 9.17467e-19 $X=8.835 $Y=2.26
+ $X2=0 $Y2=0
cc_873 N_A_1399_473#_c_1300_n N_A_1252_451#_M1000_g 0.00111142f $X=9.11 $Y=2.175
+ $X2=0 $Y2=0
cc_874 N_A_1399_473#_c_1307_n N_A_1252_451#_c_1433_n 0.0034542f $X=9.025 $Y=2.26
+ $X2=0 $Y2=0
cc_875 N_A_1399_473#_c_1308_n N_A_1252_451#_c_1433_n 8.15859e-19 $X=8.835
+ $Y=2.26 $X2=0 $Y2=0
cc_876 N_A_1399_473#_c_1299_n N_A_1252_451#_c_1421_n 0.01369f $X=9.025 $Y=1.07
+ $X2=0 $Y2=0
cc_877 N_A_1399_473#_M1024_g N_A_1252_451#_c_1424_n 7.31742e-19 $X=7.46 $Y=0.835
+ $X2=0 $Y2=0
cc_878 N_A_1399_473#_M1024_g N_A_1252_451#_c_1425_n 4.19809e-19 $X=7.46 $Y=0.835
+ $X2=0 $Y2=0
cc_879 N_A_1399_473#_M1024_g N_A_1252_451#_c_1426_n 0.0127305f $X=7.46 $Y=0.835
+ $X2=0 $Y2=0
cc_880 N_A_1399_473#_c_1299_n N_A_1252_451#_c_1426_n 0.00389968f $X=9.025
+ $Y=1.07 $X2=0 $Y2=0
cc_881 N_A_1399_473#_c_1301_n N_A_1252_451#_c_1426_n 0.0255354f $X=8.465
+ $Y=0.835 $X2=0 $Y2=0
cc_882 N_A_1399_473#_M1024_g N_A_1252_451#_c_1428_n 0.0116307f $X=7.46 $Y=0.835
+ $X2=0 $Y2=0
cc_883 N_A_1399_473#_c_1299_n N_A_1252_451#_c_1437_n 0.0135689f $X=9.025 $Y=1.07
+ $X2=0 $Y2=0
cc_884 N_A_1399_473#_c_1307_n N_A_1252_451#_c_1437_n 0.00141578f $X=9.025
+ $Y=2.26 $X2=0 $Y2=0
cc_885 N_A_1399_473#_c_1308_n N_A_1252_451#_c_1437_n 0.0120926f $X=8.835 $Y=2.26
+ $X2=0 $Y2=0
cc_886 N_A_1399_473#_c_1300_n N_A_1252_451#_c_1437_n 0.0488596f $X=9.11 $Y=2.175
+ $X2=0 $Y2=0
cc_887 N_A_1399_473#_c_1300_n N_A_1252_451#_c_1429_n 0.00600241f $X=9.11
+ $Y=2.175 $X2=0 $Y2=0
cc_888 N_A_1399_473#_c_1299_n N_A_1836_47#_c_1569_n 0.0141411f $X=9.025 $Y=1.07
+ $X2=0 $Y2=0
cc_889 N_A_1399_473#_c_1300_n N_A_1836_47#_c_1569_n 0.00218347f $X=9.11 $Y=2.175
+ $X2=0 $Y2=0
cc_890 N_A_1399_473#_c_1299_n N_A_1836_47#_c_1571_n 0.00464527f $X=9.025 $Y=1.07
+ $X2=0 $Y2=0
cc_891 N_A_1399_473#_c_1301_n N_A_1836_47#_c_1571_n 0.00569312f $X=8.465
+ $Y=0.835 $X2=0 $Y2=0
cc_892 N_A_1399_473#_c_1308_n N_A_1836_47#_c_1578_n 0.00451933f $X=8.835 $Y=2.26
+ $X2=0 $Y2=0
cc_893 N_A_1399_473#_c_1307_n N_A_1836_47#_c_1572_n 0.0141753f $X=9.025 $Y=2.26
+ $X2=0 $Y2=0
cc_894 N_A_1399_473#_c_1308_n N_A_1836_47#_c_1572_n 0.00609466f $X=8.835 $Y=2.26
+ $X2=0 $Y2=0
cc_895 N_A_1399_473#_c_1300_n N_A_1836_47#_c_1572_n 0.0500412f $X=9.11 $Y=2.175
+ $X2=0 $Y2=0
cc_896 N_A_1399_473#_c_1300_n N_A_1836_47#_c_1573_n 0.0266757f $X=9.11 $Y=2.175
+ $X2=0 $Y2=0
cc_897 N_A_1399_473#_c_1307_n N_VPWR_c_1653_n 0.00805426f $X=9.025 $Y=2.26 $X2=0
+ $Y2=0
cc_898 N_A_1399_473#_c_1308_n N_VPWR_c_1653_n 0.00866367f $X=8.835 $Y=2.26 $X2=0
+ $Y2=0
cc_899 N_A_1399_473#_c_1305_n N_VPWR_c_1663_n 0.00232082f $X=8.33 $Y=2.52 $X2=0
+ $Y2=0
cc_900 N_A_1399_473#_c_1306_n N_VPWR_c_1663_n 0.0109693f $X=8.435 $Y=2.885 $X2=0
+ $Y2=0
cc_901 N_A_1399_473#_c_1308_n N_VPWR_c_1663_n 0.00238332f $X=8.835 $Y=2.26 $X2=0
+ $Y2=0
cc_902 N_A_1399_473#_M1005_g N_VPWR_c_1668_n 0.0041647f $X=7.07 $Y=2.885 $X2=0
+ $Y2=0
cc_903 N_A_1399_473#_M1005_g N_VPWR_c_1669_n 0.0123727f $X=7.07 $Y=2.885 $X2=0
+ $Y2=0
cc_904 N_A_1399_473#_c_1305_n N_VPWR_c_1669_n 0.0238243f $X=8.33 $Y=2.52 $X2=0
+ $Y2=0
cc_905 N_A_1399_473#_c_1310_n N_VPWR_c_1669_n 0.0209779f $X=7.66 $Y=2.35 $X2=0
+ $Y2=0
cc_906 N_A_1399_473#_c_1311_n N_VPWR_c_1669_n 0.00966479f $X=7.66 $Y=2.35 $X2=0
+ $Y2=0
cc_907 N_A_1399_473#_c_1312_n N_VPWR_c_1669_n 0.00113203f $X=7.385 $Y=2.35 $X2=0
+ $Y2=0
cc_908 N_A_1399_473#_M1031_d N_VPWR_c_1648_n 0.00263469f $X=8.295 $Y=2.675 $X2=0
+ $Y2=0
cc_909 N_A_1399_473#_M1005_g N_VPWR_c_1648_n 0.00714868f $X=7.07 $Y=2.885 $X2=0
+ $Y2=0
cc_910 N_A_1399_473#_c_1305_n N_VPWR_c_1648_n 0.00513151f $X=8.33 $Y=2.52 $X2=0
+ $Y2=0
cc_911 N_A_1399_473#_c_1306_n N_VPWR_c_1648_n 0.00758253f $X=8.435 $Y=2.885
+ $X2=0 $Y2=0
cc_912 N_A_1399_473#_c_1308_n N_VPWR_c_1648_n 0.00452851f $X=8.835 $Y=2.26 $X2=0
+ $Y2=0
cc_913 N_A_1399_473#_c_1310_n N_VPWR_c_1648_n 0.00103341f $X=7.66 $Y=2.35 $X2=0
+ $Y2=0
cc_914 N_A_1399_473#_M1024_g N_VGND_c_1916_n 0.0103471f $X=7.46 $Y=0.835 $X2=0
+ $Y2=0
cc_915 N_A_1399_473#_c_1301_n N_VGND_c_1916_n 0.00719333f $X=8.465 $Y=0.835
+ $X2=0 $Y2=0
cc_916 N_A_1399_473#_M1024_g N_VGND_c_1922_n 0.00345209f $X=7.46 $Y=0.835 $X2=0
+ $Y2=0
cc_917 N_A_1399_473#_c_1301_n N_VGND_c_1926_n 0.00524028f $X=8.465 $Y=0.835
+ $X2=0 $Y2=0
cc_918 N_A_1399_473#_M1024_g N_VGND_c_1931_n 0.00394323f $X=7.46 $Y=0.835 $X2=0
+ $Y2=0
cc_919 N_A_1399_473#_c_1301_n N_VGND_c_1931_n 0.00950543f $X=8.465 $Y=0.835
+ $X2=0 $Y2=0
cc_920 N_A_1252_451#_c_1420_n N_A_1836_47#_M1029_g 0.00563542f $X=9.52 $Y=1.755
+ $X2=0 $Y2=0
cc_921 N_A_1252_451#_c_1434_n N_A_1836_47#_M1029_g 0.0267099f $X=9.6 $Y=1.83
+ $X2=0 $Y2=0
cc_922 N_A_1252_451#_M1013_g N_A_1836_47#_c_1569_n 0.0131358f $X=9.52 $Y=0.445
+ $X2=0 $Y2=0
cc_923 N_A_1252_451#_M1013_g N_A_1836_47#_c_1570_n 0.00297383f $X=9.52 $Y=0.445
+ $X2=0 $Y2=0
cc_924 N_A_1252_451#_c_1420_n N_A_1836_47#_c_1570_n 0.00297383f $X=9.52 $Y=1.755
+ $X2=0 $Y2=0
cc_925 N_A_1252_451#_c_1422_n N_A_1836_47#_c_1570_n 0.00192766f $X=9.52 $Y=1.35
+ $X2=0 $Y2=0
cc_926 N_A_1252_451#_c_1434_n N_A_1836_47#_c_1570_n 0.00329215f $X=9.6 $Y=1.83
+ $X2=0 $Y2=0
cc_927 N_A_1252_451#_c_1418_n N_A_1836_47#_c_1571_n 0.00425397f $X=9.445 $Y=1.35
+ $X2=0 $Y2=0
cc_928 N_A_1252_451#_M1013_g N_A_1836_47#_c_1571_n 0.00824423f $X=9.52 $Y=0.445
+ $X2=0 $Y2=0
cc_929 N_A_1252_451#_M1016_g N_A_1836_47#_c_1578_n 0.00393506f $X=8.65 $Y=2.885
+ $X2=0 $Y2=0
cc_930 N_A_1252_451#_M1000_g N_A_1836_47#_c_1578_n 0.00615098f $X=9.6 $Y=2.775
+ $X2=0 $Y2=0
cc_931 N_A_1252_451#_M1016_g N_A_1836_47#_c_1572_n 0.00125167f $X=8.65 $Y=2.885
+ $X2=0 $Y2=0
cc_932 N_A_1252_451#_c_1420_n N_A_1836_47#_c_1572_n 0.00857282f $X=9.52 $Y=1.755
+ $X2=0 $Y2=0
cc_933 N_A_1252_451#_M1000_g N_A_1836_47#_c_1572_n 0.0156955f $X=9.6 $Y=2.775
+ $X2=0 $Y2=0
cc_934 N_A_1252_451#_c_1434_n N_A_1836_47#_c_1572_n 0.0068023f $X=9.6 $Y=1.83
+ $X2=0 $Y2=0
cc_935 N_A_1252_451#_c_1418_n N_A_1836_47#_c_1573_n 0.00329229f $X=9.445 $Y=1.35
+ $X2=0 $Y2=0
cc_936 N_A_1252_451#_M1013_g N_A_1836_47#_c_1573_n 0.00336353f $X=9.52 $Y=0.445
+ $X2=0 $Y2=0
cc_937 N_A_1252_451#_c_1420_n N_A_1836_47#_c_1573_n 0.00179612f $X=9.52 $Y=1.755
+ $X2=0 $Y2=0
cc_938 N_A_1252_451#_c_1422_n N_A_1836_47#_c_1573_n 0.00155371f $X=9.52 $Y=1.35
+ $X2=0 $Y2=0
cc_939 N_A_1252_451#_M1013_g N_A_1836_47#_c_1574_n 0.0214019f $X=9.52 $Y=0.445
+ $X2=0 $Y2=0
cc_940 N_A_1252_451#_M1013_g N_A_1836_47#_c_1575_n 0.0162256f $X=9.52 $Y=0.445
+ $X2=0 $Y2=0
cc_941 N_A_1252_451#_M1016_g N_VPWR_c_1653_n 0.00893402f $X=8.65 $Y=2.885 $X2=0
+ $Y2=0
cc_942 N_A_1252_451#_M1000_g N_VPWR_c_1653_n 0.00230008f $X=9.6 $Y=2.775 $X2=0
+ $Y2=0
cc_943 N_A_1252_451#_c_1434_n N_VPWR_c_1654_n 0.0101681f $X=9.6 $Y=1.83 $X2=0
+ $Y2=0
cc_944 N_A_1252_451#_M1016_g N_VPWR_c_1663_n 0.00363971f $X=8.65 $Y=2.885 $X2=0
+ $Y2=0
cc_945 N_A_1252_451#_M1000_g N_VPWR_c_1664_n 0.00541359f $X=9.6 $Y=2.775 $X2=0
+ $Y2=0
cc_946 N_A_1252_451#_M1016_g N_VPWR_c_1669_n 5.8e-19 $X=8.65 $Y=2.885 $X2=0
+ $Y2=0
cc_947 N_A_1252_451#_M1030_d N_VPWR_c_1648_n 0.00301588f $X=6.26 $Y=2.255 $X2=0
+ $Y2=0
cc_948 N_A_1252_451#_M1016_g N_VPWR_c_1648_n 0.00440307f $X=8.65 $Y=2.885 $X2=0
+ $Y2=0
cc_949 N_A_1252_451#_M1000_g N_VPWR_c_1648_n 0.0110999f $X=9.6 $Y=2.775 $X2=0
+ $Y2=0
cc_950 N_A_1252_451#_M1018_g N_VGND_c_1916_n 0.00146293f $X=8.25 $Y=0.835 $X2=0
+ $Y2=0
cc_951 N_A_1252_451#_c_1426_n N_VGND_c_1916_n 0.0108087f $X=8.685 $Y=1.41 $X2=0
+ $Y2=0
cc_952 N_A_1252_451#_M1013_g N_VGND_c_1917_n 0.00451113f $X=9.52 $Y=0.445 $X2=0
+ $Y2=0
cc_953 N_A_1252_451#_M1018_g N_VGND_c_1926_n 0.00400553f $X=8.25 $Y=0.835 $X2=0
+ $Y2=0
cc_954 N_A_1252_451#_M1013_g N_VGND_c_1926_n 0.00392529f $X=9.52 $Y=0.445 $X2=0
+ $Y2=0
cc_955 N_A_1252_451#_M1013_g N_VGND_c_1930_n 0.00951772f $X=9.52 $Y=0.445 $X2=0
+ $Y2=0
cc_956 N_A_1252_451#_M1018_g N_VGND_c_1931_n 0.00469432f $X=8.25 $Y=0.835 $X2=0
+ $Y2=0
cc_957 N_A_1252_451#_M1013_g N_VGND_c_1931_n 0.00678231f $X=9.52 $Y=0.445 $X2=0
+ $Y2=0
cc_958 N_A_1836_47#_c_1578_n N_VPWR_c_1653_n 0.023127f $X=9.385 $Y=2.61 $X2=0
+ $Y2=0
cc_959 N_A_1836_47#_M1029_g N_VPWR_c_1654_n 0.0241211f $X=10.11 $Y=2.465 $X2=0
+ $Y2=0
cc_960 N_A_1836_47#_M1033_g N_VPWR_c_1654_n 8.20832e-19 $X=10.54 $Y=2.465 $X2=0
+ $Y2=0
cc_961 N_A_1836_47#_c_1570_n N_VPWR_c_1654_n 0.0186313f $X=9.97 $Y=1.35 $X2=0
+ $Y2=0
cc_962 N_A_1836_47#_c_1572_n N_VPWR_c_1654_n 0.0717335f $X=9.387 $Y=2.515 $X2=0
+ $Y2=0
cc_963 N_A_1836_47#_c_1574_n N_VPWR_c_1654_n 0.00497129f $X=9.995 $Y=1.26 $X2=0
+ $Y2=0
cc_964 N_A_1836_47#_M1033_g N_VPWR_c_1656_n 0.00768196f $X=10.54 $Y=2.465 $X2=0
+ $Y2=0
cc_965 N_A_1836_47#_c_1578_n N_VPWR_c_1664_n 0.0212431f $X=9.385 $Y=2.61 $X2=0
+ $Y2=0
cc_966 N_A_1836_47#_M1029_g N_VPWR_c_1665_n 0.00486043f $X=10.11 $Y=2.465 $X2=0
+ $Y2=0
cc_967 N_A_1836_47#_M1033_g N_VPWR_c_1665_n 0.00585385f $X=10.54 $Y=2.465 $X2=0
+ $Y2=0
cc_968 N_A_1836_47#_M1000_s N_VPWR_c_1648_n 0.00215158f $X=9.26 $Y=2.455 $X2=0
+ $Y2=0
cc_969 N_A_1836_47#_M1029_g N_VPWR_c_1648_n 0.00824727f $X=10.11 $Y=2.465 $X2=0
+ $Y2=0
cc_970 N_A_1836_47#_M1033_g N_VPWR_c_1648_n 0.0114778f $X=10.54 $Y=2.465 $X2=0
+ $Y2=0
cc_971 N_A_1836_47#_c_1578_n N_VPWR_c_1648_n 0.0127122f $X=9.385 $Y=2.61 $X2=0
+ $Y2=0
cc_972 N_A_1836_47#_c_1564_n N_Q_c_1895_n 0.0159384f $X=10.465 $Y=1.26 $X2=0
+ $Y2=0
cc_973 N_A_1836_47#_c_1565_n N_Q_c_1895_n 0.00310445f $X=10.54 $Y=1.185 $X2=0
+ $Y2=0
cc_974 N_A_1836_47#_M1033_g N_Q_c_1895_n 0.0134794f $X=10.54 $Y=2.465 $X2=0
+ $Y2=0
cc_975 N_A_1836_47#_c_1570_n N_Q_c_1895_n 0.0262167f $X=9.97 $Y=1.35 $X2=0 $Y2=0
cc_976 N_A_1836_47#_c_1572_n N_Q_c_1895_n 0.00763602f $X=9.387 $Y=2.515 $X2=0
+ $Y2=0
cc_977 N_A_1836_47#_c_1574_n N_Q_c_1895_n 0.00633118f $X=9.995 $Y=1.26 $X2=0
+ $Y2=0
cc_978 N_A_1836_47#_c_1575_n N_Q_c_1895_n 0.00329488f $X=9.995 $Y=1.185 $X2=0
+ $Y2=0
cc_979 N_A_1836_47#_c_1569_n N_VGND_c_1917_n 0.0151926f $X=9.45 $Y=1.185 $X2=0
+ $Y2=0
cc_980 N_A_1836_47#_c_1570_n N_VGND_c_1917_n 0.0270048f $X=9.97 $Y=1.35 $X2=0
+ $Y2=0
cc_981 N_A_1836_47#_c_1571_n N_VGND_c_1917_n 0.0135994f $X=9.45 $Y=0.73 $X2=0
+ $Y2=0
cc_982 N_A_1836_47#_c_1574_n N_VGND_c_1917_n 0.00518432f $X=9.995 $Y=1.26 $X2=0
+ $Y2=0
cc_983 N_A_1836_47#_c_1575_n N_VGND_c_1917_n 0.00907365f $X=9.995 $Y=1.185 $X2=0
+ $Y2=0
cc_984 N_A_1836_47#_c_1565_n N_VGND_c_1919_n 0.00707803f $X=10.54 $Y=1.185 $X2=0
+ $Y2=0
cc_985 N_A_1836_47#_c_1568_n N_VGND_c_1926_n 0.0171244f $X=9.305 $Y=0.445 $X2=0
+ $Y2=0
cc_986 N_A_1836_47#_c_1571_n N_VGND_c_1926_n 0.00189247f $X=9.45 $Y=0.73 $X2=0
+ $Y2=0
cc_987 N_A_1836_47#_c_1565_n N_VGND_c_1927_n 0.00585385f $X=10.54 $Y=1.185 $X2=0
+ $Y2=0
cc_988 N_A_1836_47#_c_1575_n N_VGND_c_1927_n 0.00487821f $X=9.995 $Y=1.185 $X2=0
+ $Y2=0
cc_989 N_A_1836_47#_c_1565_n N_VGND_c_1930_n 6.87751e-19 $X=10.54 $Y=1.185 $X2=0
+ $Y2=0
cc_990 N_A_1836_47#_c_1575_n N_VGND_c_1930_n 0.0107919f $X=9.995 $Y=1.185 $X2=0
+ $Y2=0
cc_991 N_A_1836_47#_M1013_s N_VGND_c_1931_n 0.00233128f $X=9.18 $Y=0.235 $X2=0
+ $Y2=0
cc_992 N_A_1836_47#_c_1565_n N_VGND_c_1931_n 0.0114778f $X=10.54 $Y=1.185 $X2=0
+ $Y2=0
cc_993 N_A_1836_47#_c_1568_n N_VGND_c_1931_n 0.00989078f $X=9.305 $Y=0.445 $X2=0
+ $Y2=0
cc_994 N_A_1836_47#_c_1571_n N_VGND_c_1931_n 0.00343684f $X=9.45 $Y=0.73 $X2=0
+ $Y2=0
cc_995 N_A_1836_47#_c_1575_n N_VGND_c_1931_n 0.00824731f $X=9.995 $Y=1.185 $X2=0
+ $Y2=0
cc_996 N_VPWR_c_1648_n N_A_318_535#_M1001_s 0.00238695f $X=10.8 $Y=3.33 $X2=0
+ $Y2=0
cc_997 N_VPWR_c_1648_n N_A_318_535#_M1026_d 0.00254682f $X=10.8 $Y=3.33 $X2=0
+ $Y2=0
cc_998 N_VPWR_c_1662_n N_A_318_535#_c_1807_n 0.0152571f $X=1.98 $Y=3.33 $X2=0
+ $Y2=0
cc_999 N_VPWR_c_1648_n N_A_318_535#_c_1807_n 0.00988478f $X=10.8 $Y=3.33 $X2=0
+ $Y2=0
cc_1000 N_VPWR_c_1650_n N_A_318_535#_c_1808_n 0.0206626f $X=2.145 $Y=2.885 $X2=0
+ $Y2=0
cc_1001 N_VPWR_c_1657_n N_A_318_535#_c_1808_n 0.00229131f $X=3.755 $Y=3.33 $X2=0
+ $Y2=0
cc_1002 N_VPWR_c_1662_n N_A_318_535#_c_1808_n 0.00229131f $X=1.98 $Y=3.33 $X2=0
+ $Y2=0
cc_1003 N_VPWR_c_1648_n N_A_318_535#_c_1808_n 0.00901193f $X=10.8 $Y=3.33 $X2=0
+ $Y2=0
cc_1004 N_VPWR_c_1657_n N_A_318_535#_c_1810_n 0.0115999f $X=3.755 $Y=3.33 $X2=0
+ $Y2=0
cc_1005 N_VPWR_c_1648_n N_A_318_535#_c_1810_n 0.00835226f $X=10.8 $Y=3.33 $X2=0
+ $Y2=0
cc_1006 N_VPWR_c_1657_n N_A_318_535#_c_1811_n 0.00225293f $X=3.755 $Y=3.33 $X2=0
+ $Y2=0
cc_1007 N_VPWR_c_1648_n N_A_318_535#_c_1811_n 0.00408011f $X=10.8 $Y=3.33 $X2=0
+ $Y2=0
cc_1008 N_VPWR_c_1648_n A_667_535# 0.0016963f $X=10.8 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_1009 N_VPWR_c_1648_n A_1357_535# 0.00168881f $X=10.8 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_1010 N_VPWR_c_1648_n N_Q_M1029_d 0.0041489f $X=10.8 $Y=3.33 $X2=0 $Y2=0
cc_1011 N_VPWR_c_1654_n N_Q_c_1895_n 0.0481331f $X=9.895 $Y=1.98 $X2=0 $Y2=0
cc_1012 N_VPWR_c_1656_n N_Q_c_1895_n 0.0015231f $X=10.755 $Y=1.98 $X2=0 $Y2=0
cc_1013 N_VPWR_c_1665_n N_Q_c_1895_n 0.0136943f $X=10.625 $Y=3.33 $X2=0 $Y2=0
cc_1014 N_VPWR_c_1648_n N_Q_c_1895_n 0.00866972f $X=10.8 $Y=3.33 $X2=0 $Y2=0
cc_1015 N_Q_c_1895_n N_VGND_c_1919_n 0.0015231f $X=10.325 $Y=0.42 $X2=0 $Y2=0
cc_1016 N_Q_c_1895_n N_VGND_c_1927_n 0.0136943f $X=10.325 $Y=0.42 $X2=0 $Y2=0
cc_1017 N_Q_M1022_d N_VGND_c_1931_n 0.0041489f $X=10.185 $Y=0.235 $X2=0 $Y2=0
cc_1018 N_Q_c_1895_n N_VGND_c_1931_n 0.00866972f $X=10.325 $Y=0.42 $X2=0 $Y2=0
