* File: sky130_fd_sc_lp__or3_4.pxi.spice
* Created: Wed Sep  2 10:30:41 2020
* 
x_PM_SKY130_FD_SC_LP__OR3_4%C N_C_M1001_g N_C_M1000_g C C N_C_c_82_n
+ PM_SKY130_FD_SC_LP__OR3_4%C
x_PM_SKY130_FD_SC_LP__OR3_4%B N_B_M1003_g N_B_M1006_g B N_B_c_108_n N_B_c_109_n
+ PM_SKY130_FD_SC_LP__OR3_4%B
x_PM_SKY130_FD_SC_LP__OR3_4%A N_A_M1007_g N_A_M1013_g A N_A_c_141_n N_A_c_142_n
+ PM_SKY130_FD_SC_LP__OR3_4%A
x_PM_SKY130_FD_SC_LP__OR3_4%A_77_49# N_A_77_49#_M1001_s N_A_77_49#_M1006_d
+ N_A_77_49#_M1000_s N_A_77_49#_M1004_g N_A_77_49#_M1002_g N_A_77_49#_M1008_g
+ N_A_77_49#_M1005_g N_A_77_49#_M1009_g N_A_77_49#_M1010_g N_A_77_49#_M1012_g
+ N_A_77_49#_M1011_g N_A_77_49#_c_185_n N_A_77_49#_c_199_n N_A_77_49#_c_200_n
+ N_A_77_49#_c_186_n N_A_77_49#_c_187_n N_A_77_49#_c_212_n N_A_77_49#_c_230_n
+ N_A_77_49#_c_188_n N_A_77_49#_c_189_n N_A_77_49#_c_190_n N_A_77_49#_c_191_n
+ N_A_77_49#_c_192_n N_A_77_49#_c_193_n N_A_77_49#_c_194_n
+ PM_SKY130_FD_SC_LP__OR3_4%A_77_49#
x_PM_SKY130_FD_SC_LP__OR3_4%VPWR N_VPWR_M1007_d N_VPWR_M1005_s N_VPWR_M1011_s
+ N_VPWR_c_332_n N_VPWR_c_333_n N_VPWR_c_334_n N_VPWR_c_335_n N_VPWR_c_336_n
+ N_VPWR_c_337_n N_VPWR_c_338_n N_VPWR_c_339_n VPWR N_VPWR_c_340_n
+ N_VPWR_c_331_n N_VPWR_c_342_n PM_SKY130_FD_SC_LP__OR3_4%VPWR
x_PM_SKY130_FD_SC_LP__OR3_4%X N_X_M1004_d N_X_M1009_d N_X_M1002_d N_X_M1010_d
+ N_X_c_443_p N_X_c_429_n N_X_c_383_n N_X_c_384_n N_X_c_390_n N_X_c_391_n
+ N_X_c_440_p N_X_c_433_n N_X_c_392_n N_X_c_385_n N_X_c_386_n N_X_c_393_n X X X
+ X X PM_SKY130_FD_SC_LP__OR3_4%X
x_PM_SKY130_FD_SC_LP__OR3_4%VGND N_VGND_M1001_d N_VGND_M1013_d N_VGND_M1008_s
+ N_VGND_M1012_s N_VGND_c_450_n N_VGND_c_451_n N_VGND_c_452_n N_VGND_c_453_n
+ N_VGND_c_454_n N_VGND_c_455_n N_VGND_c_456_n N_VGND_c_457_n N_VGND_c_458_n
+ N_VGND_c_459_n N_VGND_c_460_n VGND N_VGND_c_461_n N_VGND_c_462_n
+ N_VGND_c_463_n PM_SKY130_FD_SC_LP__OR3_4%VGND
cc_1 VNB N_C_M1001_g 0.0295566f $X=-0.19 $Y=-0.245 $X2=0.725 $Y2=0.665
cc_2 VNB N_C_M1000_g 0.00158796f $X=-0.19 $Y=-0.245 $X2=0.725 $Y2=2.465
cc_3 VNB C 0.0268271f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_4 VNB N_C_c_82_n 0.0363925f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.46
cc_5 VNB N_B_M1006_g 0.0249911f $X=-0.19 $Y=-0.245 $X2=0.725 $Y2=2.465
cc_6 VNB N_B_c_108_n 0.0242554f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_B_c_109_n 0.00359456f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.46
cc_8 VNB N_A_M1013_g 0.0252226f $X=-0.19 $Y=-0.245 $X2=0.725 $Y2=2.465
cc_9 VNB N_A_c_141_n 0.0244148f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_c_142_n 0.00315322f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.46
cc_11 VNB N_A_77_49#_M1004_g 0.0239529f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_77_49#_M1008_g 0.0222554f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_77_49#_M1009_g 0.0222627f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_77_49#_M1012_g 0.0284259f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_77_49#_c_185_n 0.0285156f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_77_49#_c_186_n 0.00690176f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_77_49#_c_187_n 0.0097895f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_77_49#_c_188_n 0.00458312f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_77_49#_c_189_n 0.00227391f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_77_49#_c_190_n 3.45182e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_77_49#_c_191_n 0.0015776f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_77_49#_c_192_n 0.0805981f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_77_49#_c_193_n 0.00780685f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_77_49#_c_194_n 0.0010166f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_VPWR_c_331_n 0.183584f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_X_c_383_n 0.00310505f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_X_c_384_n 0.00266908f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_X_c_385_n 0.0102619f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_X_c_386_n 0.00180538f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB X 0.0368049f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB X 0.00815223f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB X 0.0202758f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_450_n 0.00537487f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.46
cc_34 VNB N_VGND_c_451_n 0.00266123f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_452_n 4.86514e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_453_n 0.0148369f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_454_n 0.00474568f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_455_n 0.0251627f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_456_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_457_n 0.0170188f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_458_n 0.00599098f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_459_n 0.0137079f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_460_n 0.00451663f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_461_n 0.0169569f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_462_n 0.248639f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_463_n 0.00452017f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VPB N_C_M1000_g 0.0249467f $X=-0.19 $Y=1.655 $X2=0.725 $Y2=2.465
cc_48 VPB C 0.0183042f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_49 VPB N_B_M1003_g 0.0192559f $X=-0.19 $Y=1.655 $X2=0.725 $Y2=0.665
cc_50 VPB N_B_c_108_n 0.00637381f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_51 VPB N_B_c_109_n 0.0023898f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.46
cc_52 VPB N_A_M1007_g 0.0210711f $X=-0.19 $Y=1.655 $X2=0.725 $Y2=0.665
cc_53 VPB N_A_c_141_n 0.00617736f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_54 VPB N_A_c_142_n 0.00234877f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.46
cc_55 VPB N_A_77_49#_M1002_g 0.0195509f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.295
cc_56 VPB N_A_77_49#_M1005_g 0.018006f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_57 VPB N_A_77_49#_M1010_g 0.0180133f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_58 VPB N_A_77_49#_M1011_g 0.0217749f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_59 VPB N_A_77_49#_c_199_n 0.00797287f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_60 VPB N_A_77_49#_c_200_n 0.0379885f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_61 VPB N_A_77_49#_c_190_n 0.00148424f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_62 VPB N_A_77_49#_c_192_n 0.0171987f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_63 VPB N_VPWR_c_332_n 0.00512086f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_64 VPB N_VPWR_c_333_n 3.177e-19 $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.295
cc_65 VPB N_VPWR_c_334_n 0.0129398f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_335_n 0.040815f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_67 VPB N_VPWR_c_336_n 0.0544595f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_337_n 0.00680245f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_69 VPB N_VPWR_c_338_n 0.0155777f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_70 VPB N_VPWR_c_339_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_71 VPB N_VPWR_c_340_n 0.0164632f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_72 VPB N_VPWR_c_331_n 0.0694175f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_73 VPB N_VPWR_c_342_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_74 VPB N_X_c_390_n 0.00310505f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_75 VPB N_X_c_391_n 0.00191858f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_76 VPB N_X_c_392_n 0.024814f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_77 VPB N_X_c_393_n 0.00147023f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_78 VPB X 0.00624245f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_79 N_C_M1000_g N_B_M1003_g 0.0589968f $X=0.725 $Y=2.465 $X2=0 $Y2=0
cc_80 N_C_M1001_g N_B_M1006_g 0.0196349f $X=0.725 $Y=0.665 $X2=0 $Y2=0
cc_81 C N_B_c_108_n 0.00231555f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_82 N_C_c_82_n N_B_c_108_n 0.0589968f $X=0.635 $Y=1.46 $X2=0 $Y2=0
cc_83 C N_B_c_109_n 0.0314179f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_84 N_C_c_82_n N_B_c_109_n 6.19219e-19 $X=0.635 $Y=1.46 $X2=0 $Y2=0
cc_85 N_C_M1000_g N_A_77_49#_c_199_n 7.54694e-19 $X=0.725 $Y=2.465 $X2=0 $Y2=0
cc_86 C N_A_77_49#_c_199_n 0.0261742f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_87 N_C_c_82_n N_A_77_49#_c_199_n 9.13663e-19 $X=0.635 $Y=1.46 $X2=0 $Y2=0
cc_88 N_C_M1000_g N_A_77_49#_c_200_n 0.0195724f $X=0.725 $Y=2.465 $X2=0 $Y2=0
cc_89 N_C_M1001_g N_A_77_49#_c_186_n 0.0152125f $X=0.725 $Y=0.665 $X2=0 $Y2=0
cc_90 C N_A_77_49#_c_186_n 0.0135541f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_91 N_C_c_82_n N_A_77_49#_c_186_n 2.37192e-19 $X=0.635 $Y=1.46 $X2=0 $Y2=0
cc_92 C N_A_77_49#_c_187_n 0.0219575f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_93 N_C_c_82_n N_A_77_49#_c_187_n 0.0042767f $X=0.635 $Y=1.46 $X2=0 $Y2=0
cc_94 N_C_M1000_g N_A_77_49#_c_212_n 0.0108953f $X=0.725 $Y=2.465 $X2=0 $Y2=0
cc_95 C N_A_77_49#_c_212_n 0.0113571f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_96 N_C_M1000_g N_VPWR_c_336_n 0.0054895f $X=0.725 $Y=2.465 $X2=0 $Y2=0
cc_97 N_C_M1000_g N_VPWR_c_331_n 0.0109514f $X=0.725 $Y=2.465 $X2=0 $Y2=0
cc_98 N_C_M1001_g N_VGND_c_450_n 0.00320431f $X=0.725 $Y=0.665 $X2=0 $Y2=0
cc_99 N_C_M1001_g N_VGND_c_455_n 0.00575161f $X=0.725 $Y=0.665 $X2=0 $Y2=0
cc_100 N_C_M1001_g N_VGND_c_462_n 0.0118402f $X=0.725 $Y=0.665 $X2=0 $Y2=0
cc_101 N_B_M1003_g N_A_M1007_g 0.051844f $X=1.085 $Y=2.465 $X2=0 $Y2=0
cc_102 N_B_M1006_g N_A_M1013_g 0.0238903f $X=1.235 $Y=0.665 $X2=0 $Y2=0
cc_103 N_B_c_108_n N_A_c_141_n 0.0214125f $X=1.175 $Y=1.51 $X2=0 $Y2=0
cc_104 N_B_c_109_n N_A_c_141_n 0.00129309f $X=1.175 $Y=1.51 $X2=0 $Y2=0
cc_105 N_B_c_108_n N_A_c_142_n 0.00102106f $X=1.175 $Y=1.51 $X2=0 $Y2=0
cc_106 N_B_c_109_n N_A_c_142_n 0.0333427f $X=1.175 $Y=1.51 $X2=0 $Y2=0
cc_107 N_B_M1003_g N_A_77_49#_c_200_n 0.0048871f $X=1.085 $Y=2.465 $X2=0 $Y2=0
cc_108 N_B_M1006_g N_A_77_49#_c_186_n 0.0134296f $X=1.235 $Y=0.665 $X2=0 $Y2=0
cc_109 N_B_c_108_n N_A_77_49#_c_186_n 0.00157771f $X=1.175 $Y=1.51 $X2=0 $Y2=0
cc_110 N_B_c_109_n N_A_77_49#_c_186_n 0.0202656f $X=1.175 $Y=1.51 $X2=0 $Y2=0
cc_111 N_B_M1003_g N_A_77_49#_c_212_n 0.0159785f $X=1.085 $Y=2.465 $X2=0 $Y2=0
cc_112 N_B_c_108_n N_A_77_49#_c_212_n 9.23487e-19 $X=1.175 $Y=1.51 $X2=0 $Y2=0
cc_113 N_B_c_109_n N_A_77_49#_c_212_n 0.0232322f $X=1.175 $Y=1.51 $X2=0 $Y2=0
cc_114 N_B_M1006_g N_A_77_49#_c_193_n 9.21681e-19 $X=1.235 $Y=0.665 $X2=0 $Y2=0
cc_115 N_B_c_108_n N_A_77_49#_c_193_n 2.35676e-19 $X=1.175 $Y=1.51 $X2=0 $Y2=0
cc_116 N_B_c_109_n N_A_77_49#_c_193_n 0.0036811f $X=1.175 $Y=1.51 $X2=0 $Y2=0
cc_117 N_B_M1003_g N_VPWR_c_336_n 0.00585385f $X=1.085 $Y=2.465 $X2=0 $Y2=0
cc_118 N_B_M1003_g N_VPWR_c_331_n 0.011101f $X=1.085 $Y=2.465 $X2=0 $Y2=0
cc_119 N_B_M1006_g N_VGND_c_450_n 0.00173997f $X=1.235 $Y=0.665 $X2=0 $Y2=0
cc_120 N_B_M1006_g N_VGND_c_457_n 0.00575161f $X=1.235 $Y=0.665 $X2=0 $Y2=0
cc_121 N_B_M1006_g N_VGND_c_462_n 0.0107942f $X=1.235 $Y=0.665 $X2=0 $Y2=0
cc_122 N_A_M1013_g N_A_77_49#_M1004_g 0.0155957f $X=1.665 $Y=0.665 $X2=0 $Y2=0
cc_123 N_A_M1007_g N_A_77_49#_M1002_g 0.0349521f $X=1.625 $Y=2.465 $X2=0 $Y2=0
cc_124 N_A_c_142_n N_A_77_49#_M1002_g 2.03002e-19 $X=1.715 $Y=1.51 $X2=0 $Y2=0
cc_125 N_A_M1007_g N_A_77_49#_c_212_n 0.0167565f $X=1.625 $Y=2.465 $X2=0 $Y2=0
cc_126 N_A_c_141_n N_A_77_49#_c_212_n 0.00299606f $X=1.715 $Y=1.51 $X2=0 $Y2=0
cc_127 N_A_c_142_n N_A_77_49#_c_212_n 0.0186451f $X=1.715 $Y=1.51 $X2=0 $Y2=0
cc_128 N_A_M1013_g N_A_77_49#_c_230_n 0.00943712f $X=1.665 $Y=0.665 $X2=0 $Y2=0
cc_129 N_A_M1013_g N_A_77_49#_c_188_n 0.0131755f $X=1.665 $Y=0.665 $X2=0 $Y2=0
cc_130 N_A_c_141_n N_A_77_49#_c_188_n 0.00311896f $X=1.715 $Y=1.51 $X2=0 $Y2=0
cc_131 N_A_c_142_n N_A_77_49#_c_188_n 0.0151419f $X=1.715 $Y=1.51 $X2=0 $Y2=0
cc_132 N_A_M1013_g N_A_77_49#_c_189_n 0.00357135f $X=1.665 $Y=0.665 $X2=0 $Y2=0
cc_133 N_A_c_141_n N_A_77_49#_c_189_n 5.26016e-19 $X=1.715 $Y=1.51 $X2=0 $Y2=0
cc_134 N_A_c_142_n N_A_77_49#_c_189_n 0.0059077f $X=1.715 $Y=1.51 $X2=0 $Y2=0
cc_135 N_A_M1007_g N_A_77_49#_c_190_n 0.00347303f $X=1.625 $Y=2.465 $X2=0 $Y2=0
cc_136 N_A_c_141_n N_A_77_49#_c_190_n 5.26016e-19 $X=1.715 $Y=1.51 $X2=0 $Y2=0
cc_137 N_A_c_142_n N_A_77_49#_c_190_n 0.0117847f $X=1.715 $Y=1.51 $X2=0 $Y2=0
cc_138 N_A_c_141_n N_A_77_49#_c_192_n 0.0168326f $X=1.715 $Y=1.51 $X2=0 $Y2=0
cc_139 N_A_c_142_n N_A_77_49#_c_192_n 2.91186e-19 $X=1.715 $Y=1.51 $X2=0 $Y2=0
cc_140 N_A_M1013_g N_A_77_49#_c_193_n 0.00106769f $X=1.665 $Y=0.665 $X2=0 $Y2=0
cc_141 N_A_c_141_n N_A_77_49#_c_193_n 3.10581e-19 $X=1.715 $Y=1.51 $X2=0 $Y2=0
cc_142 N_A_c_142_n N_A_77_49#_c_193_n 0.00575866f $X=1.715 $Y=1.51 $X2=0 $Y2=0
cc_143 N_A_c_141_n N_A_77_49#_c_194_n 0.00129183f $X=1.715 $Y=1.51 $X2=0 $Y2=0
cc_144 N_A_c_142_n N_A_77_49#_c_194_n 0.0141929f $X=1.715 $Y=1.51 $X2=0 $Y2=0
cc_145 N_A_M1007_g N_VPWR_c_332_n 0.00824772f $X=1.625 $Y=2.465 $X2=0 $Y2=0
cc_146 N_A_M1007_g N_VPWR_c_336_n 0.00585385f $X=1.625 $Y=2.465 $X2=0 $Y2=0
cc_147 N_A_M1007_g N_VPWR_c_331_n 0.011482f $X=1.625 $Y=2.465 $X2=0 $Y2=0
cc_148 N_A_M1013_g N_VGND_c_451_n 0.00176741f $X=1.665 $Y=0.665 $X2=0 $Y2=0
cc_149 N_A_M1013_g N_VGND_c_457_n 0.00569184f $X=1.665 $Y=0.665 $X2=0 $Y2=0
cc_150 N_A_M1013_g N_VGND_c_462_n 0.0107208f $X=1.665 $Y=0.665 $X2=0 $Y2=0
cc_151 N_A_77_49#_c_212_n A_160_367# 0.00737677f $X=1.98 $Y=2.01 $X2=-0.19
+ $Y2=-0.245
cc_152 N_A_77_49#_c_212_n A_232_367# 0.0174471f $X=1.98 $Y=2.01 $X2=-0.19
+ $Y2=-0.245
cc_153 N_A_77_49#_c_212_n N_VPWR_M1007_d 0.00909525f $X=1.98 $Y=2.01 $X2=-0.19
+ $Y2=-0.245
cc_154 N_A_77_49#_c_190_n N_VPWR_M1007_d 0.00106149f $X=2.065 $Y=1.92 $X2=-0.19
+ $Y2=-0.245
cc_155 N_A_77_49#_M1002_g N_VPWR_c_332_n 0.0070625f $X=2.2 $Y=2.465 $X2=0 $Y2=0
cc_156 N_A_77_49#_c_212_n N_VPWR_c_332_n 0.0260654f $X=1.98 $Y=2.01 $X2=0 $Y2=0
cc_157 N_A_77_49#_M1002_g N_VPWR_c_333_n 7.41729e-19 $X=2.2 $Y=2.465 $X2=0 $Y2=0
cc_158 N_A_77_49#_M1005_g N_VPWR_c_333_n 0.0141912f $X=2.63 $Y=2.465 $X2=0 $Y2=0
cc_159 N_A_77_49#_M1010_g N_VPWR_c_333_n 0.014077f $X=3.06 $Y=2.465 $X2=0 $Y2=0
cc_160 N_A_77_49#_M1011_g N_VPWR_c_333_n 7.21513e-19 $X=3.49 $Y=2.465 $X2=0
+ $Y2=0
cc_161 N_A_77_49#_M1010_g N_VPWR_c_334_n 0.00486043f $X=3.06 $Y=2.465 $X2=0
+ $Y2=0
cc_162 N_A_77_49#_M1011_g N_VPWR_c_334_n 0.00486043f $X=3.49 $Y=2.465 $X2=0
+ $Y2=0
cc_163 N_A_77_49#_M1010_g N_VPWR_c_335_n 7.21513e-19 $X=3.06 $Y=2.465 $X2=0
+ $Y2=0
cc_164 N_A_77_49#_M1011_g N_VPWR_c_335_n 0.0151817f $X=3.49 $Y=2.465 $X2=0 $Y2=0
cc_165 N_A_77_49#_c_200_n N_VPWR_c_336_n 0.0210467f $X=0.51 $Y=2.95 $X2=0 $Y2=0
cc_166 N_A_77_49#_M1002_g N_VPWR_c_338_n 0.00585385f $X=2.2 $Y=2.465 $X2=0 $Y2=0
cc_167 N_A_77_49#_M1005_g N_VPWR_c_338_n 0.00486043f $X=2.63 $Y=2.465 $X2=0
+ $Y2=0
cc_168 N_A_77_49#_M1000_s N_VPWR_c_331_n 0.00215158f $X=0.385 $Y=1.835 $X2=0
+ $Y2=0
cc_169 N_A_77_49#_M1002_g N_VPWR_c_331_n 0.0110314f $X=2.2 $Y=2.465 $X2=0 $Y2=0
cc_170 N_A_77_49#_M1005_g N_VPWR_c_331_n 0.00824727f $X=2.63 $Y=2.465 $X2=0
+ $Y2=0
cc_171 N_A_77_49#_M1010_g N_VPWR_c_331_n 0.00824727f $X=3.06 $Y=2.465 $X2=0
+ $Y2=0
cc_172 N_A_77_49#_M1011_g N_VPWR_c_331_n 0.00824727f $X=3.49 $Y=2.465 $X2=0
+ $Y2=0
cc_173 N_A_77_49#_c_200_n N_VPWR_c_331_n 0.0125689f $X=0.51 $Y=2.95 $X2=0 $Y2=0
cc_174 N_A_77_49#_M1008_g N_X_c_383_n 0.0138138f $X=2.63 $Y=0.665 $X2=0 $Y2=0
cc_175 N_A_77_49#_M1009_g N_X_c_383_n 0.01419f $X=3.06 $Y=0.665 $X2=0 $Y2=0
cc_176 N_A_77_49#_c_191_n N_X_c_383_n 0.0447065f $X=3.65 $Y=1.51 $X2=0 $Y2=0
cc_177 N_A_77_49#_c_192_n N_X_c_383_n 0.00244902f $X=3.65 $Y=1.51 $X2=0 $Y2=0
cc_178 N_A_77_49#_M1004_g N_X_c_384_n 0.00131418f $X=2.2 $Y=0.665 $X2=0 $Y2=0
cc_179 N_A_77_49#_c_188_n N_X_c_384_n 0.00750776f $X=1.98 $Y=1.08 $X2=0 $Y2=0
cc_180 N_A_77_49#_c_189_n N_X_c_384_n 0.00641961f $X=2.065 $Y=1.425 $X2=0 $Y2=0
cc_181 N_A_77_49#_c_191_n N_X_c_384_n 0.014687f $X=3.65 $Y=1.51 $X2=0 $Y2=0
cc_182 N_A_77_49#_c_192_n N_X_c_384_n 0.00255521f $X=3.65 $Y=1.51 $X2=0 $Y2=0
cc_183 N_A_77_49#_M1005_g N_X_c_390_n 0.0128776f $X=2.63 $Y=2.465 $X2=0 $Y2=0
cc_184 N_A_77_49#_M1010_g N_X_c_390_n 0.0129862f $X=3.06 $Y=2.465 $X2=0 $Y2=0
cc_185 N_A_77_49#_c_191_n N_X_c_390_n 0.0447065f $X=3.65 $Y=1.51 $X2=0 $Y2=0
cc_186 N_A_77_49#_c_192_n N_X_c_390_n 0.00244902f $X=3.65 $Y=1.51 $X2=0 $Y2=0
cc_187 N_A_77_49#_M1002_g N_X_c_391_n 4.90985e-19 $X=2.2 $Y=2.465 $X2=0 $Y2=0
cc_188 N_A_77_49#_c_190_n N_X_c_391_n 0.00765392f $X=2.065 $Y=1.92 $X2=0 $Y2=0
cc_189 N_A_77_49#_c_191_n N_X_c_391_n 0.014687f $X=3.65 $Y=1.51 $X2=0 $Y2=0
cc_190 N_A_77_49#_c_192_n N_X_c_391_n 0.00255521f $X=3.65 $Y=1.51 $X2=0 $Y2=0
cc_191 N_A_77_49#_M1011_g N_X_c_392_n 0.0149355f $X=3.49 $Y=2.465 $X2=0 $Y2=0
cc_192 N_A_77_49#_c_191_n N_X_c_392_n 0.0298871f $X=3.65 $Y=1.51 $X2=0 $Y2=0
cc_193 N_A_77_49#_c_192_n N_X_c_392_n 0.00612256f $X=3.65 $Y=1.51 $X2=0 $Y2=0
cc_194 N_A_77_49#_M1012_g N_X_c_385_n 0.0168733f $X=3.49 $Y=0.665 $X2=0 $Y2=0
cc_195 N_A_77_49#_c_191_n N_X_c_385_n 0.0274884f $X=3.65 $Y=1.51 $X2=0 $Y2=0
cc_196 N_A_77_49#_c_192_n N_X_c_385_n 0.00612256f $X=3.65 $Y=1.51 $X2=0 $Y2=0
cc_197 N_A_77_49#_c_191_n N_X_c_386_n 0.017393f $X=3.65 $Y=1.51 $X2=0 $Y2=0
cc_198 N_A_77_49#_c_192_n N_X_c_386_n 0.00255521f $X=3.65 $Y=1.51 $X2=0 $Y2=0
cc_199 N_A_77_49#_c_191_n N_X_c_393_n 0.014687f $X=3.65 $Y=1.51 $X2=0 $Y2=0
cc_200 N_A_77_49#_c_192_n N_X_c_393_n 0.00255521f $X=3.65 $Y=1.51 $X2=0 $Y2=0
cc_201 N_A_77_49#_M1012_g X 0.00330895f $X=3.49 $Y=0.665 $X2=0 $Y2=0
cc_202 N_A_77_49#_M1012_g X 0.00262005f $X=3.49 $Y=0.665 $X2=0 $Y2=0
cc_203 N_A_77_49#_M1011_g X 0.00262005f $X=3.49 $Y=2.465 $X2=0 $Y2=0
cc_204 N_A_77_49#_c_191_n X 0.0134813f $X=3.65 $Y=1.51 $X2=0 $Y2=0
cc_205 N_A_77_49#_c_192_n X 0.00793466f $X=3.65 $Y=1.51 $X2=0 $Y2=0
cc_206 N_A_77_49#_c_186_n N_VGND_M1001_d 0.00261503f $X=1.31 $Y=1.08 $X2=-0.19
+ $Y2=-0.245
cc_207 N_A_77_49#_c_188_n N_VGND_M1013_d 0.00303168f $X=1.98 $Y=1.08 $X2=0 $Y2=0
cc_208 N_A_77_49#_c_186_n N_VGND_c_450_n 0.0200142f $X=1.31 $Y=1.08 $X2=0 $Y2=0
cc_209 N_A_77_49#_M1004_g N_VGND_c_451_n 0.00869773f $X=2.2 $Y=0.665 $X2=0 $Y2=0
cc_210 N_A_77_49#_M1008_g N_VGND_c_451_n 5.89572e-19 $X=2.63 $Y=0.665 $X2=0
+ $Y2=0
cc_211 N_A_77_49#_c_188_n N_VGND_c_451_n 0.0230827f $X=1.98 $Y=1.08 $X2=0 $Y2=0
cc_212 N_A_77_49#_M1004_g N_VGND_c_452_n 6.23374e-19 $X=2.2 $Y=0.665 $X2=0 $Y2=0
cc_213 N_A_77_49#_M1008_g N_VGND_c_452_n 0.011284f $X=2.63 $Y=0.665 $X2=0 $Y2=0
cc_214 N_A_77_49#_M1009_g N_VGND_c_452_n 0.0113159f $X=3.06 $Y=0.665 $X2=0 $Y2=0
cc_215 N_A_77_49#_M1012_g N_VGND_c_452_n 6.29009e-19 $X=3.49 $Y=0.665 $X2=0
+ $Y2=0
cc_216 N_A_77_49#_M1009_g N_VGND_c_453_n 0.00477554f $X=3.06 $Y=0.665 $X2=0
+ $Y2=0
cc_217 N_A_77_49#_M1012_g N_VGND_c_453_n 0.00575161f $X=3.49 $Y=0.665 $X2=0
+ $Y2=0
cc_218 N_A_77_49#_M1012_g N_VGND_c_454_n 0.00332009f $X=3.49 $Y=0.665 $X2=0
+ $Y2=0
cc_219 N_A_77_49#_c_185_n N_VGND_c_455_n 0.0190529f $X=0.51 $Y=0.42 $X2=0 $Y2=0
cc_220 N_A_77_49#_c_230_n N_VGND_c_457_n 0.0159213f $X=1.45 $Y=0.42 $X2=0 $Y2=0
cc_221 N_A_77_49#_M1004_g N_VGND_c_459_n 0.00554242f $X=2.2 $Y=0.665 $X2=0 $Y2=0
cc_222 N_A_77_49#_M1008_g N_VGND_c_459_n 0.00477554f $X=2.63 $Y=0.665 $X2=0
+ $Y2=0
cc_223 N_A_77_49#_M1001_s N_VGND_c_462_n 0.00247088f $X=0.385 $Y=0.245 $X2=0
+ $Y2=0
cc_224 N_A_77_49#_M1006_d N_VGND_c_462_n 0.00223559f $X=1.31 $Y=0.245 $X2=0
+ $Y2=0
cc_225 N_A_77_49#_M1004_g N_VGND_c_462_n 0.00949547f $X=2.2 $Y=0.665 $X2=0 $Y2=0
cc_226 N_A_77_49#_M1008_g N_VGND_c_462_n 0.00825815f $X=2.63 $Y=0.665 $X2=0
+ $Y2=0
cc_227 N_A_77_49#_M1009_g N_VGND_c_462_n 0.00825815f $X=3.06 $Y=0.665 $X2=0
+ $Y2=0
cc_228 N_A_77_49#_M1012_g N_VGND_c_462_n 0.0118351f $X=3.49 $Y=0.665 $X2=0 $Y2=0
cc_229 N_A_77_49#_c_185_n N_VGND_c_462_n 0.0113912f $X=0.51 $Y=0.42 $X2=0 $Y2=0
cc_230 N_A_77_49#_c_230_n N_VGND_c_462_n 0.0109109f $X=1.45 $Y=0.42 $X2=0 $Y2=0
cc_231 A_160_367# N_VPWR_c_331_n 0.00899413f $X=0.8 $Y=1.835 $X2=0.51 $Y2=2.95
cc_232 A_232_367# N_VPWR_c_331_n 0.0167135f $X=1.16 $Y=1.835 $X2=0.51 $Y2=2.95
cc_233 N_VPWR_c_331_n N_X_M1002_d 0.00536646f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_234 N_VPWR_c_331_n N_X_M1010_d 0.00536646f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_235 N_VPWR_c_338_n N_X_c_429_n 0.0124525f $X=2.68 $Y=3.33 $X2=0 $Y2=0
cc_236 N_VPWR_c_331_n N_X_c_429_n 0.00730901f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_237 N_VPWR_M1005_s N_X_c_390_n 0.00176461f $X=2.705 $Y=1.835 $X2=0 $Y2=0
cc_238 N_VPWR_c_333_n N_X_c_390_n 0.0170777f $X=2.845 $Y=2.2 $X2=0 $Y2=0
cc_239 N_VPWR_c_334_n N_X_c_433_n 0.0124525f $X=3.54 $Y=3.33 $X2=0 $Y2=0
cc_240 N_VPWR_c_331_n N_X_c_433_n 0.00730901f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_241 N_VPWR_M1011_s N_X_c_392_n 0.0027239f $X=3.565 $Y=1.835 $X2=0 $Y2=0
cc_242 N_VPWR_c_335_n N_X_c_392_n 0.0220026f $X=3.705 $Y=2.2 $X2=0 $Y2=0
cc_243 N_X_c_383_n N_VGND_M1008_s 0.00176461f $X=3.18 $Y=1.16 $X2=0 $Y2=0
cc_244 N_X_c_385_n N_VGND_M1012_s 0.00283146f $X=3.98 $Y=1.16 $X2=0 $Y2=0
cc_245 N_X_c_383_n N_VGND_c_452_n 0.0170777f $X=3.18 $Y=1.16 $X2=0 $Y2=0
cc_246 N_X_c_440_p N_VGND_c_453_n 0.0136943f $X=3.275 $Y=0.42 $X2=0 $Y2=0
cc_247 N_X_c_385_n N_VGND_c_454_n 0.015214f $X=3.98 $Y=1.16 $X2=0 $Y2=0
cc_248 X N_VGND_c_454_n 0.0419418f $X=3.995 $Y=0.47 $X2=0 $Y2=0
cc_249 N_X_c_443_p N_VGND_c_459_n 0.0124525f $X=2.415 $Y=0.42 $X2=0 $Y2=0
cc_250 X N_VGND_c_461_n 0.00800499f $X=3.995 $Y=0.47 $X2=0 $Y2=0
cc_251 N_X_M1004_d N_VGND_c_462_n 0.00536646f $X=2.275 $Y=0.245 $X2=0 $Y2=0
cc_252 N_X_M1009_d N_VGND_c_462_n 0.0041489f $X=3.135 $Y=0.245 $X2=0 $Y2=0
cc_253 N_X_c_443_p N_VGND_c_462_n 0.00730901f $X=2.415 $Y=0.42 $X2=0 $Y2=0
cc_254 N_X_c_440_p N_VGND_c_462_n 0.00866972f $X=3.275 $Y=0.42 $X2=0 $Y2=0
cc_255 X N_VGND_c_462_n 0.00673845f $X=3.995 $Y=0.47 $X2=0 $Y2=0
