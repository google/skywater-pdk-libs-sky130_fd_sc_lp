* File: sky130_fd_sc_lp__o31ai_m.pex.spice
* Created: Wed Sep  2 10:25:43 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O31AI_M%A1 2 5 6 8 10 11 13 16 18 19 20 21 27
r38 27 28 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.385
+ $Y=1.34 $X2=0.385 $Y2=1.34
r39 20 21 13.5366 $w=3.13e-07 $l=3.7e-07 $layer=LI1_cond $X=0.312 $Y=2.035
+ $X2=0.312 $Y2=2.405
r40 19 20 13.5366 $w=3.13e-07 $l=3.7e-07 $layer=LI1_cond $X=0.312 $Y=1.665
+ $X2=0.312 $Y2=2.035
r41 19 28 11.8903 $w=3.13e-07 $l=3.25e-07 $layer=LI1_cond $X=0.312 $Y=1.665
+ $X2=0.312 $Y2=1.34
r42 18 28 1.64635 $w=3.13e-07 $l=4.5e-08 $layer=LI1_cond $X=0.312 $Y=1.295
+ $X2=0.312 $Y2=1.34
r43 14 16 112.809 $w=1.5e-07 $l=2.2e-07 $layer=POLY_cond $X=0.475 $Y=2.49
+ $X2=0.695 $Y2=2.49
r44 12 27 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.385 $Y=1.68
+ $X2=0.385 $Y2=1.34
r45 12 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.385 $Y=1.68
+ $X2=0.385 $Y2=1.845
r46 11 27 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=0.385 $Y=1.325
+ $X2=0.385 $Y2=1.34
r47 10 11 43.5886 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=0.425 $Y=1.175
+ $X2=0.425 $Y2=1.325
r48 6 16 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.695 $Y=2.565
+ $X2=0.695 $Y2=2.49
r49 6 8 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.695 $Y=2.565
+ $X2=0.695 $Y2=2.885
r50 5 10 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.555 $Y=0.855
+ $X2=0.555 $Y2=1.175
r51 2 14 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.475 $Y=2.415
+ $X2=0.475 $Y2=2.49
r52 2 13 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=0.475 $Y=2.415
+ $X2=0.475 $Y2=1.845
.ends

.subckt PM_SKY130_FD_SC_LP__O31AI_M%A2 3 7 11 12 13 14 15 20
r46 20 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.965
+ $Y=1.7 $X2=0.965 $Y2=1.7
r47 14 15 10.5285 $w=4.03e-07 $l=3.7e-07 $layer=LI1_cond $X=1.082 $Y=2.035
+ $X2=1.082 $Y2=2.405
r48 14 21 9.53255 $w=4.03e-07 $l=3.35e-07 $layer=LI1_cond $X=1.082 $Y=2.035
+ $X2=1.082 $Y2=1.7
r49 13 21 0.995938 $w=4.03e-07 $l=3.5e-08 $layer=LI1_cond $X=1.082 $Y=1.665
+ $X2=1.082 $Y2=1.7
r50 11 20 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.965 $Y=2.04
+ $X2=0.965 $Y2=1.7
r51 11 12 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.965 $Y=2.04
+ $X2=0.965 $Y2=2.205
r52 10 20 38.6168 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.965 $Y=1.535
+ $X2=0.965 $Y2=1.7
r53 7 12 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=1.055 $Y=2.885
+ $X2=1.055 $Y2=2.205
r54 3 10 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=0.985 $Y=0.855
+ $X2=0.985 $Y2=1.535
.ends

.subckt PM_SKY130_FD_SC_LP__O31AI_M%A3 3 7 11 14 15 16 20
r44 15 16 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=1.68 $Y=1.665
+ $X2=1.68 $Y2=2.035
r45 15 20 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.68 $Y=1.7
+ $X2=1.68 $Y2=1.7
r46 13 20 42.4591 $w=4.65e-07 $l=3.55e-07 $layer=POLY_cond $X=1.612 $Y=2.055
+ $X2=1.612 $Y2=1.7
r47 13 14 45.5629 $w=4.65e-07 $l=1.5e-07 $layer=POLY_cond $X=1.592 $Y=2.055
+ $X2=1.592 $Y2=2.205
r48 11 20 1.79404 $w=4.65e-07 $l=1.5e-08 $layer=POLY_cond $X=1.612 $Y=1.685
+ $X2=1.612 $Y2=1.7
r49 10 11 45.5629 $w=4.65e-07 $l=1.5e-07 $layer=POLY_cond $X=1.592 $Y=1.535
+ $X2=1.592 $Y2=1.685
r50 7 14 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=1.415 $Y=2.885
+ $X2=1.415 $Y2=2.205
r51 3 10 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=1.415 $Y=0.855
+ $X2=1.415 $Y2=1.535
.ends

.subckt PM_SKY130_FD_SC_LP__O31AI_M%B1 4 5 7 8 9 10 11 13 14 15 19
c43 10 0 1.13044e-19 $X=2.085 $Y=2.49
c44 4 0 9.98462e-20 $X=1.845 $Y=0.855
r45 19 22 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.935 $Y=0.37
+ $X2=1.935 $Y2=0.535
r46 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.935
+ $Y=0.37 $X2=1.935 $Y2=0.37
r47 15 20 7.30422 $w=3.53e-07 $l=2.25e-07 $layer=LI1_cond $X=2.16 $Y=0.462
+ $X2=1.935 $Y2=0.462
r48 14 20 8.27811 $w=3.53e-07 $l=2.55e-07 $layer=LI1_cond $X=1.68 $Y=0.462
+ $X2=1.935 $Y2=0.462
r49 12 13 558.915 $w=1.5e-07 $l=1.09e-06 $layer=POLY_cond $X=2.16 $Y=1.325
+ $X2=2.16 $Y2=2.415
r50 10 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.085 $Y=2.49
+ $X2=2.16 $Y2=2.415
r51 10 11 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.085 $Y=2.49
+ $X2=1.92 $Y2=2.49
r52 8 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.085 $Y=1.25
+ $X2=2.16 $Y2=1.325
r53 8 9 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.085 $Y=1.25
+ $X2=1.92 $Y2=1.25
r54 5 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.845 $Y=2.565
+ $X2=1.92 $Y2=2.49
r55 5 7 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.845 $Y=2.565
+ $X2=1.845 $Y2=2.885
r56 4 22 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.845 $Y=0.855
+ $X2=1.845 $Y2=0.535
r57 2 9 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.845 $Y=1.175
+ $X2=1.92 $Y2=1.25
r58 2 4 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.845 $Y=1.175
+ $X2=1.845 $Y2=0.855
.ends

.subckt PM_SKY130_FD_SC_LP__O31AI_M%VPWR 1 2 9 11 13 16 17 18 24 33
c34 24 0 1.13044e-19 $X=1.955 $Y=3.33
r35 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r36 30 33 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r37 29 30 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r38 26 29 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.72 $Y=3.33 $X2=1.68
+ $Y2=3.33
r39 26 27 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r40 24 32 3.62069 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=1.955 $Y=3.33
+ $X2=2.177 $Y2=3.33
r41 24 29 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=1.955 $Y=3.33
+ $X2=1.68 $Y2=3.33
r42 22 27 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r43 21 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r44 18 30 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r45 18 27 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r46 16 21 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=0.315 $Y=3.33
+ $X2=0.24 $Y2=3.33
r47 16 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.315 $Y=3.33
+ $X2=0.48 $Y2=3.33
r48 15 26 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=0.645 $Y=3.33
+ $X2=0.72 $Y2=3.33
r49 15 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.645 $Y=3.33
+ $X2=0.48 $Y2=3.33
r50 11 32 3.2945 $w=2.1e-07 $l=1.53734e-07 $layer=LI1_cond $X=2.06 $Y=3.245
+ $X2=2.177 $Y2=3.33
r51 11 13 15.5801 $w=2.08e-07 $l=2.95e-07 $layer=LI1_cond $X=2.06 $Y=3.245
+ $X2=2.06 $Y2=2.95
r52 7 17 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.48 $Y=3.245 $X2=0.48
+ $Y2=3.33
r53 7 9 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.48 $Y=3.245
+ $X2=0.48 $Y2=2.95
r54 2 13 600 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=1 $X=1.92
+ $Y=2.675 $X2=2.06 $Y2=2.95
r55 1 9 600 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_PDIFF $count=1 $X=0.355
+ $Y=2.675 $X2=0.48 $Y2=2.95
.ends

.subckt PM_SKY130_FD_SC_LP__O31AI_M%Y 1 2 7 11 13
r32 13 15 14.8852 $w=2.09e-07 $l=2.55e-07 $layer=LI1_cond $X=1.645 $Y=2.775
+ $X2=1.645 $Y2=2.52
r33 9 11 52.9076 $w=3.28e-07 $l=1.515e-06 $layer=LI1_cond $X=2.14 $Y=2.435
+ $X2=2.14 $Y2=0.92
r34 8 15 1.94907 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=1.765 $Y=2.52
+ $X2=1.645 $Y2=2.52
r35 7 9 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.975 $Y=2.52
+ $X2=2.14 $Y2=2.435
r36 7 8 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=1.975 $Y=2.52
+ $X2=1.765 $Y2=2.52
r37 2 13 600 $w=1.7e-07 $l=2.4e-07 $layer=licon1_PDIFF $count=1 $X=1.49 $Y=2.675
+ $X2=1.63 $Y2=2.855
r38 1 11 182 $w=1.7e-07 $l=3.68951e-07 $layer=licon1_NDIFF $count=1 $X=1.92
+ $Y=0.645 $X2=2.14 $Y2=0.92
.ends

.subckt PM_SKY130_FD_SC_LP__O31AI_M%VGND 1 2 7 9 13 15 17 24 25 31
r28 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r29 24 25 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r30 22 31 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.285 $Y=0 $X2=1.19
+ $Y2=0
r31 22 24 57.0856 $w=1.68e-07 $l=8.75e-07 $layer=LI1_cond $X=1.285 $Y=0 $X2=2.16
+ $Y2=0
r32 21 29 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r33 20 21 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r34 18 28 3.61992 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=0 $X2=0.222
+ $Y2=0
r35 18 20 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.445 $Y=0 $X2=0.72
+ $Y2=0
r36 17 31 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.095 $Y=0 $X2=1.19
+ $Y2=0
r37 17 20 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.095 $Y=0 $X2=0.72
+ $Y2=0
r38 15 25 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r39 15 21 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r40 15 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r41 11 31 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.19 $Y=0.085
+ $X2=1.19 $Y2=0
r42 11 13 39.9856 $w=1.88e-07 $l=6.85e-07 $layer=LI1_cond $X=1.19 $Y=0.085
+ $X2=1.19 $Y2=0.77
r43 7 28 3.29527 $w=2.1e-07 $l=1.54771e-07 $layer=LI1_cond $X=0.34 $Y=0.085
+ $X2=0.222 $Y2=0
r44 7 9 37.2338 $w=2.08e-07 $l=7.05e-07 $layer=LI1_cond $X=0.34 $Y=0.085
+ $X2=0.34 $Y2=0.79
r45 2 13 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=1.06
+ $Y=0.645 $X2=1.2 $Y2=0.77
r46 1 9 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.215
+ $Y=0.645 $X2=0.34 $Y2=0.79
.ends

.subckt PM_SKY130_FD_SC_LP__O31AI_M%A_126_129# 1 2 9 11 12 14
c24 11 0 9.98462e-20 $X=1.465 $Y=1.2
r25 14 16 9.7783 $w=3.28e-07 $l=2.8e-07 $layer=LI1_cond $X=1.63 $Y=0.92 $X2=1.63
+ $Y2=1.2
r26 11 16 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.465 $Y=1.2
+ $X2=1.63 $Y2=1.2
r27 11 12 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=1.465 $Y=1.2
+ $X2=0.875 $Y2=1.2
r28 7 12 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=0.77 $Y=1.115
+ $X2=0.875 $Y2=1.2
r29 7 9 9.24242 $w=2.08e-07 $l=1.75e-07 $layer=LI1_cond $X=0.77 $Y=1.115
+ $X2=0.77 $Y2=0.94
r30 2 14 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=1.49
+ $Y=0.645 $X2=1.63 $Y2=0.92
r31 1 9 182 $w=1.7e-07 $l=3.58225e-07 $layer=licon1_NDIFF $count=1 $X=0.63
+ $Y=0.645 $X2=0.77 $Y2=0.94
.ends

