* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__o41a_lp A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
X0 a_349_412# A4 a_457_412# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X1 VGND A2 a_31_57# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 a_457_412# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X3 VGND a_457_412# a_708_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 VPWR A1 a_137_412# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X5 a_137_412# A2 a_235_412# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X6 VPWR a_457_412# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X7 a_31_57# A1 VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 a_235_412# A3 a_349_412# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X9 a_31_57# A3 VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 a_708_47# a_457_412# X VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X11 VGND A4 a_31_57# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 a_31_57# B1 a_457_412# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
