* File: sky130_fd_sc_lp__iso0n_lp.spice
* Created: Wed Sep  2 09:57:41 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__iso0n_lp.pex.spice"
.subckt sky130_fd_sc_lp__iso0n_lp  VNB VPB A SLEEP_B VPWR X KAGND VGND
* 
* KAGND	KAGND
* X	X
* VPWR	VPWR
* SLEEP_B	SLEEP_B
* A	A
* VPB	VPB
* VNB	VNB
MM1007 A_221_93# N_A_M1007_g N_A_138_93#_M1007_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1113 PD=0.63 PS=1.37 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.9 A=0.063 P=1.14 MULT=1
MM1008 N_KAGND_M1008_d N_SLEEP_B_M1008_g A_221_93# VNB NSHORT L=0.15 W=0.42
+ AD=0.1785 AS=0.0441 PD=1.27 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6
+ SB=75001.6 A=0.063 P=1.14 MULT=1
MM1002 A_493_93# N_A_138_93#_M1002_g N_KAGND_M1008_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1785 PD=0.63 PS=1.27 NRD=14.28 NRS=1.428 M=1 R=2.8 SA=75001.6
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1004 N_X_M1004_d N_A_138_93#_M1004_g A_493_93# VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.0441 PD=1.37 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.9
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1009 A_149_489# N_A_M1009_g N_VPWR_M1009_s VPB PHIGHVT L=0.15 W=0.42 AD=0.0441
+ AS=0.1113 PD=0.63 PS=1.37 NRD=23.443 NRS=0 M=1 R=2.8 SA=75000.2 SB=75002.3
+ A=0.063 P=1.14 MULT=1
MM1005 N_A_138_93#_M1005_d N_A_M1005_g A_149_489# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=23.443 M=1 R=2.8 SA=75000.6
+ SB=75001.9 A=0.063 P=1.14 MULT=1
MM1000 A_307_489# N_SLEEP_B_M1000_g N_A_138_93#_M1005_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=23.443 NRS=0 M=1 R=2.8 SA=75001
+ SB=75001.5 A=0.063 P=1.14 MULT=1
MM1001 N_VPWR_M1001_d N_SLEEP_B_M1001_g A_307_489# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.09975 AS=0.0441 PD=0.84 PS=0.63 NRD=68.0044 NRS=23.443 M=1 R=2.8
+ SA=75001.3 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1003 A_493_367# N_A_138_93#_M1003_g N_VPWR_M1001_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1323 AS=0.29925 PD=1.47 PS=2.52 NRD=7.8012 NRS=0 M=1 R=8.4 SA=75000.8
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1006 N_X_M1006_d N_A_138_93#_M1006_g A_493_367# VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.1323 PD=3.05 PS=1.47 NRD=0 NRS=7.8012 M=1 R=8.4 SA=75001.1
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.96577 P=11.2
c_24 VNB 0 1.48936e-19 $X=0 $Y=0
*
.include "sky130_fd_sc_lp__iso0n_lp.pxi.spice"
*
.ends
*
*
