* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__or4b_m A B C D_N VGND VNB VPB VPWR X
X0 a_215_125# A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 a_38_125# D_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X2 a_215_125# a_38_125# a_338_397# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X3 VGND a_38_125# a_215_125# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 a_38_125# D_N VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 VGND B a_215_125# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 a_215_125# C VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 VGND a_215_125# X VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 VPWR a_215_125# X VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X9 a_338_397# C a_410_397# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X10 a_410_397# B a_482_397# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X11 a_482_397# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
.ends
