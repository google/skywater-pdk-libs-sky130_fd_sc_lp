* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__o22a_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
X0 X a_86_23# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X1 VPWR B1 a_608_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X2 a_86_23# A2 a_982_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X3 VPWR A1 a_982_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X4 VGND a_86_23# X VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X5 X a_86_23# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X6 a_86_23# B1 a_525_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X7 a_525_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X8 a_608_367# B2 a_86_23# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X9 a_982_367# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X10 VGND a_86_23# X VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X11 VGND A2 a_525_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X12 a_525_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X13 a_608_367# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X14 VGND A1 a_525_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X15 a_86_23# B2 a_608_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X16 VPWR a_86_23# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X17 X a_86_23# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X18 VPWR a_86_23# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X19 a_982_367# A2 a_86_23# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X20 a_525_47# B1 a_86_23# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X21 X a_86_23# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X22 a_86_23# B2 a_525_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X23 a_525_47# B2 a_86_23# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
.ends
