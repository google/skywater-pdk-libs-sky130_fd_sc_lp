* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
X0 a_80_237# B1 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X1 VGND A2 a_294_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X2 VGND C1 a_80_237# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X3 VPWR A1 a_217_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X4 X a_80_237# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X5 a_504_367# C1 a_80_237# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X6 a_217_367# B1 a_504_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X7 a_294_47# A1 a_80_237# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X8 X a_80_237# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X9 a_217_367# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
.ends
