* File: sky130_fd_sc_lp__xnor2_1.spice
* Created: Fri Aug 28 11:34:58 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__xnor2_1.pex.spice"
.subckt sky130_fd_sc_lp__xnor2_1  VNB VPB B A VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A	A
* B	B
* VPB	VPB
* VNB	VNB
MM1004 A_116_47# N_B_M1004_g N_A_33_47#_M1004_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1029 AS=0.2226 PD=1.085 PS=2.21 NRD=9.636 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1007 N_VGND_M1007_d N_A_M1007_g A_116_47# VNB NSHORT L=0.15 W=0.84 AD=0.2226
+ AS=0.1029 PD=2.21 PS=1.085 NRD=0 NRS=9.636 M=1 R=5.6 SA=75000.6 SB=75000.2
+ A=0.126 P=1.98 MULT=1
MM1009 N_VGND_M1009_d N_A_M1009_g N_A_302_47#_M1009_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1638 AS=0.2226 PD=1.23 PS=2.21 NRD=9.996 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75001.2 A=0.126 P=1.98 MULT=1
MM1000 N_A_302_47#_M1000_d N_B_M1000_g N_VGND_M1009_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1449 AS=0.1638 PD=1.185 PS=1.23 NRD=9.276 NRS=5.712 M=1 R=5.6 SA=75000.7
+ SB=75000.7 A=0.126 P=1.98 MULT=1
MM1003 N_Y_M1003_d N_A_33_47#_M1003_g N_A_302_47#_M1000_d VNB NSHORT L=0.15
+ W=0.84 AD=0.2226 AS=0.1449 PD=2.21 PS=1.185 NRD=0 NRS=0 M=1 R=5.6 SA=75001.2
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1002 N_A_33_47#_M1002_d N_B_M1002_g N_VPWR_M1002_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75002.6 A=0.189 P=2.82 MULT=1
MM1006 N_VPWR_M1006_d N_A_M1006_g N_A_33_47#_M1002_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.48195 AS=0.1764 PD=2.025 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75002.1 A=0.189 P=2.82 MULT=1
MM1008 A_385_367# N_A_M1008_g N_VPWR_M1006_d VPB PHIGHVT L=0.15 W=1.26 AD=0.2457
+ AS=0.48195 PD=1.65 PS=2.025 NRD=21.8867 NRS=0 M=1 R=8.4 SA=75001.5 SB=75001.2
+ A=0.189 P=2.82 MULT=1
MM1001 N_Y_M1001_d N_B_M1001_g A_385_367# VPB PHIGHVT L=0.15 W=1.26 AD=0.21735
+ AS=0.2457 PD=1.605 PS=1.65 NRD=10.1455 NRS=21.8867 M=1 R=8.4 SA=75002.1
+ SB=75000.7 A=0.189 P=2.82 MULT=1
MM1005 N_VPWR_M1005_d N_A_33_47#_M1005_g N_Y_M1001_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.21735 PD=3.05 PS=1.605 NRD=0 NRS=0 M=1 R=8.4 SA=75002.6
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9751 P=11.21
c_61 VPB 0 1.31259e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_lp__xnor2_1.pxi.spice"
*
.ends
*
*
