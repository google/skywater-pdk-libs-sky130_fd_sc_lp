* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__a32o_0 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
M1000 a_363_47# A2 a_275_47# VNB nshort w=420000u l=150000u
+  ad=1.302e+11p pd=1.46e+06u as=1.218e+11p ps=1.42e+06u
M1001 a_80_21# B1 a_269_429# VPB phighvt w=640000u l=150000u
+  ad=1.792e+11p pd=1.84e+06u as=6.016e+11p ps=5.72e+06u
M1002 VGND B2 a_563_47# VNB nshort w=420000u l=150000u
+  ad=4.011e+11p pd=3.59e+06u as=1.638e+11p ps=1.62e+06u
M1003 VPWR A2 a_269_429# VPB phighvt w=640000u l=150000u
+  ad=4.192e+11p pd=3.87e+06u as=0p ps=0u
M1004 a_275_47# A3 VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VGND a_80_21# X VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1006 a_269_429# A3 VPWR VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_80_21# A1 a_363_47# VNB nshort w=420000u l=150000u
+  ad=1.638e+11p pd=1.62e+06u as=0p ps=0u
M1008 a_269_429# B2 a_80_21# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR a_80_21# X VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.696e+11p ps=1.81e+06u
M1010 a_563_47# B1 a_80_21# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_269_429# A1 VPWR VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
