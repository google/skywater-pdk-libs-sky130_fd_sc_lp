* File: sky130_fd_sc_lp__a211o_0.pxi.spice
* Created: Fri Aug 28 09:47:18 2020
* 
x_PM_SKY130_FD_SC_LP__A211O_0%A_80_172# N_A_80_172#_M1002_d N_A_80_172#_M1000_d
+ N_A_80_172#_M1005_d N_A_80_172#_c_78_n N_A_80_172#_M1009_g N_A_80_172#_M1007_g
+ N_A_80_172#_c_81_n N_A_80_172#_c_82_n N_A_80_172#_c_83_n N_A_80_172#_c_84_n
+ N_A_80_172#_c_85_n N_A_80_172#_c_86_n N_A_80_172#_c_87_n N_A_80_172#_c_88_n
+ N_A_80_172#_c_89_n N_A_80_172#_c_90_n N_A_80_172#_c_93_n N_A_80_172#_c_91_n
+ PM_SKY130_FD_SC_LP__A211O_0%A_80_172#
x_PM_SKY130_FD_SC_LP__A211O_0%A2 N_A2_M1001_g N_A2_c_175_n N_A2_M1008_g
+ N_A2_c_172_n N_A2_c_178_n N_A2_c_179_n A2 A2 N_A2_c_174_n
+ PM_SKY130_FD_SC_LP__A211O_0%A2
x_PM_SKY130_FD_SC_LP__A211O_0%A1 N_A1_M1002_g N_A1_c_224_n N_A1_c_228_n
+ N_A1_M1006_g N_A1_c_230_n N_A1_c_231_n A1 A1 N_A1_c_226_n
+ PM_SKY130_FD_SC_LP__A211O_0%A1
x_PM_SKY130_FD_SC_LP__A211O_0%B1 N_B1_c_272_n N_B1_M1003_g N_B1_M1004_g
+ N_B1_c_273_n N_B1_c_274_n N_B1_c_275_n N_B1_c_280_n B1 B1 N_B1_c_277_n
+ PM_SKY130_FD_SC_LP__A211O_0%B1
x_PM_SKY130_FD_SC_LP__A211O_0%C1 N_C1_M1005_g N_C1_M1000_g C1 C1 C1 N_C1_c_320_n
+ PM_SKY130_FD_SC_LP__A211O_0%C1
x_PM_SKY130_FD_SC_LP__A211O_0%X N_X_M1007_s N_X_M1009_s X X X X X X X X
+ PM_SKY130_FD_SC_LP__A211O_0%X
x_PM_SKY130_FD_SC_LP__A211O_0%VPWR N_VPWR_M1009_d N_VPWR_M1008_d N_VPWR_c_361_n
+ N_VPWR_c_362_n VPWR N_VPWR_c_363_n N_VPWR_c_364_n N_VPWR_c_365_n
+ N_VPWR_c_360_n N_VPWR_c_367_n N_VPWR_c_368_n PM_SKY130_FD_SC_LP__A211O_0%VPWR
x_PM_SKY130_FD_SC_LP__A211O_0%A_224_482# N_A_224_482#_M1008_s
+ N_A_224_482#_M1006_d N_A_224_482#_c_401_n N_A_224_482#_c_402_n
+ N_A_224_482#_c_403_n N_A_224_482#_c_404_n
+ PM_SKY130_FD_SC_LP__A211O_0%A_224_482#
x_PM_SKY130_FD_SC_LP__A211O_0%VGND N_VGND_M1007_d N_VGND_M1003_d VGND
+ N_VGND_c_435_n N_VGND_c_436_n N_VGND_c_437_n N_VGND_c_438_n N_VGND_c_439_n
+ N_VGND_c_440_n PM_SKY130_FD_SC_LP__A211O_0%VGND
cc_1 VNB N_A_80_172#_c_78_n 0.0259237f $X=-0.19 $Y=-0.245 $X2=0.577 $Y2=1.353
cc_2 VNB N_A_80_172#_M1009_g 0.0076737f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.52
cc_3 VNB N_A_80_172#_M1007_g 0.0249177f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=0.51
cc_4 VNB N_A_80_172#_c_81_n 0.0197502f $X=-0.19 $Y=-0.245 $X2=0.577 $Y2=1.53
cc_5 VNB N_A_80_172#_c_82_n 0.0237457f $X=-0.19 $Y=-0.245 $X2=1.66 $Y2=0.945
cc_6 VNB N_A_80_172#_c_83_n 0.00133433f $X=-0.19 $Y=-0.245 $X2=1.825 $Y2=0.51
cc_7 VNB N_A_80_172#_c_84_n 0.0103222f $X=-0.19 $Y=-0.245 $X2=2.535 $Y2=0.945
cc_8 VNB N_A_80_172#_c_85_n 0.010396f $X=-0.19 $Y=-0.245 $X2=2.89 $Y2=0.945
cc_9 VNB N_A_80_172#_c_86_n 0.0217782f $X=-0.19 $Y=-0.245 $X2=3.025 $Y2=0.51
cc_10 VNB N_A_80_172#_c_87_n 0.00551996f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.025
cc_11 VNB N_A_80_172#_c_88_n 0.0199684f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.025
cc_12 VNB N_A_80_172#_c_89_n 0.00423472f $X=-0.19 $Y=-0.245 $X2=1.81 $Y2=0.945
cc_13 VNB N_A_80_172#_c_90_n 0.00168916f $X=-0.19 $Y=-0.245 $X2=2.62 $Y2=0.945
cc_14 VNB N_A_80_172#_c_91_n 0.0060222f $X=-0.19 $Y=-0.245 $X2=2.817 $Y2=2.39
cc_15 VNB N_A2_M1001_g 0.0377285f $X=-0.19 $Y=-0.245 $X2=2.795 $Y2=2.41
cc_16 VNB N_A2_c_172_n 0.0185318f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.52
cc_17 VNB A2 0.00479611f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A2_c_174_n 0.0155117f $X=-0.19 $Y=-0.245 $X2=0.755 $Y2=0.945
cc_19 VNB N_A1_M1002_g 0.0347158f $X=-0.19 $Y=-0.245 $X2=2.795 $Y2=2.41
cc_20 VNB N_A1_c_224_n 0.0165008f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB A1 0.00440518f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=0.51
cc_22 VNB N_A1_c_226_n 0.0175606f $X=-0.19 $Y=-0.245 $X2=1.66 $Y2=0.945
cc_23 VNB N_B1_c_272_n 0.0196f $X=-0.19 $Y=-0.245 $X2=1.685 $Y2=0.3
cc_24 VNB N_B1_c_273_n 0.0178057f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.53
cc_25 VNB N_B1_c_274_n 0.0142146f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_B1_c_275_n 0.0172247f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=0.86
cc_27 VNB B1 0.00443202f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=0.51
cc_28 VNB N_B1_c_277_n 0.0152463f $X=-0.19 $Y=-0.245 $X2=1.66 $Y2=0.945
cc_29 VNB N_C1_M1000_g 0.0513144f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB C1 0.0236409f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_C1_c_320_n 0.0499841f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=0.86
cc_32 VNB X 0.0130421f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB X 0.0495289f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VPWR_c_360_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_435_n 0.0176806f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_436_n 0.0266213f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.52
cc_37 VNB N_VGND_c_437_n 0.0201893f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_438_n 0.201261f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_439_n 0.0187734f $X=-0.19 $Y=-0.245 $X2=1.81 $Y2=0.51
cc_40 VNB N_VGND_c_440_n 0.0212819f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VPB N_A_80_172#_M1009_g 0.0479808f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.52
cc_42 VPB N_A_80_172#_c_93_n 0.0329665f $X=-0.19 $Y=1.655 $X2=2.935 $Y2=2.555
cc_43 VPB N_A_80_172#_c_91_n 0.005171f $X=-0.19 $Y=1.655 $X2=2.817 $Y2=2.39
cc_44 VPB N_A2_c_175_n 0.016337f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_45 VPB N_A2_M1008_g 0.0208376f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_46 VPB N_A2_c_172_n 0.00416442f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.52
cc_47 VPB N_A2_c_178_n 0.0167556f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.52
cc_48 VPB N_A2_c_179_n 0.0229577f $X=-0.19 $Y=1.655 $X2=0.48 $Y2=0.51
cc_49 VPB A2 0.00586982f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_50 VPB N_A1_c_224_n 0.00350805f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_51 VPB N_A1_c_228_n 0.0136953f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_52 VPB N_A1_M1006_g 0.0190001f $X=-0.19 $Y=1.655 $X2=0.577 $Y2=1.353
cc_53 VPB N_A1_c_230_n 0.0177576f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.52
cc_54 VPB N_A1_c_231_n 0.0146416f $X=-0.19 $Y=1.655 $X2=0.48 $Y2=0.86
cc_55 VPB A1 0.00350276f $X=-0.19 $Y=1.655 $X2=0.48 $Y2=0.51
cc_56 VPB N_B1_M1004_g 0.0386582f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_57 VPB N_B1_c_275_n 0.00364251f $X=-0.19 $Y=1.655 $X2=0.48 $Y2=0.86
cc_58 VPB N_B1_c_280_n 0.0153238f $X=-0.19 $Y=1.655 $X2=0.48 $Y2=0.51
cc_59 VPB B1 0.0042776f $X=-0.19 $Y=1.655 $X2=0.48 $Y2=0.51
cc_60 VPB N_C1_M1005_g 0.0435612f $X=-0.19 $Y=1.655 $X2=2.795 $Y2=2.41
cc_61 VPB C1 0.033732f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_62 VPB N_C1_c_320_n 0.0305085f $X=-0.19 $Y=1.655 $X2=0.48 $Y2=0.86
cc_63 VPB X 0.0283664f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_64 VPB X 0.00781704f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=1.53
cc_65 VPB X 0.0273039f $X=-0.19 $Y=1.655 $X2=2.89 $Y2=0.945
cc_66 VPB N_VPWR_c_361_n 0.0289083f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_67 VPB N_VPWR_c_362_n 0.00874354f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.52
cc_68 VPB N_VPWR_c_363_n 0.0176936f $X=-0.19 $Y=1.655 $X2=0.48 $Y2=0.51
cc_69 VPB N_VPWR_c_364_n 0.0192252f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_70 VPB N_VPWR_c_365_n 0.043613f $X=-0.19 $Y=1.655 $X2=2.62 $Y2=2.39
cc_71 VPB N_VPWR_c_360_n 0.0797527f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_72 VPB N_VPWR_c_367_n 0.00574453f $X=-0.19 $Y=1.655 $X2=2.705 $Y2=0.945
cc_73 VPB N_VPWR_c_368_n 0.00555219f $X=-0.19 $Y=1.655 $X2=3.025 $Y2=0.51
cc_74 VPB N_A_224_482#_c_401_n 0.0113905f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_75 VPB N_A_224_482#_c_402_n 0.016244f $X=-0.19 $Y=1.655 $X2=0.577 $Y2=1.353
cc_76 VPB N_A_224_482#_c_403_n 0.00452356f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=1.53
cc_77 VPB N_A_224_482#_c_404_n 0.00573488f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_78 N_A_80_172#_M1007_g N_A2_M1001_g 0.00572452f $X=0.48 $Y=0.51 $X2=0 $Y2=0
cc_79 N_A_80_172#_c_82_n N_A2_M1001_g 0.0120028f $X=1.66 $Y=0.945 $X2=0 $Y2=0
cc_80 N_A_80_172#_c_83_n N_A2_M1001_g 0.00182501f $X=1.825 $Y=0.51 $X2=0 $Y2=0
cc_81 N_A_80_172#_c_87_n N_A2_M1001_g 9.69962e-19 $X=0.59 $Y=1.025 $X2=0 $Y2=0
cc_82 N_A_80_172#_c_88_n N_A2_M1001_g 0.0099841f $X=0.59 $Y=1.025 $X2=0 $Y2=0
cc_83 N_A_80_172#_M1009_g N_A2_c_175_n 0.00663428f $X=0.475 $Y=2.52 $X2=0 $Y2=0
cc_84 N_A_80_172#_M1009_g N_A2_c_172_n 0.00860784f $X=0.475 $Y=2.52 $X2=0 $Y2=0
cc_85 N_A_80_172#_c_81_n N_A2_c_172_n 0.00830261f $X=0.577 $Y=1.53 $X2=0 $Y2=0
cc_86 N_A_80_172#_c_78_n A2 0.00127209f $X=0.577 $Y=1.353 $X2=0 $Y2=0
cc_87 N_A_80_172#_M1009_g A2 0.00135905f $X=0.475 $Y=2.52 $X2=0 $Y2=0
cc_88 N_A_80_172#_c_82_n A2 0.0281468f $X=1.66 $Y=0.945 $X2=0 $Y2=0
cc_89 N_A_80_172#_c_87_n A2 0.0184804f $X=0.59 $Y=1.025 $X2=0 $Y2=0
cc_90 N_A_80_172#_c_78_n N_A2_c_174_n 0.00830261f $X=0.577 $Y=1.353 $X2=0 $Y2=0
cc_91 N_A_80_172#_c_82_n N_A2_c_174_n 0.00121059f $X=1.66 $Y=0.945 $X2=0 $Y2=0
cc_92 N_A_80_172#_c_87_n N_A2_c_174_n 0.00117583f $X=0.59 $Y=1.025 $X2=0 $Y2=0
cc_93 N_A_80_172#_c_82_n N_A1_M1002_g 0.00819152f $X=1.66 $Y=0.945 $X2=0 $Y2=0
cc_94 N_A_80_172#_c_83_n N_A1_M1002_g 0.0102122f $X=1.825 $Y=0.51 $X2=0 $Y2=0
cc_95 N_A_80_172#_c_89_n N_A1_M1002_g 0.00293734f $X=1.81 $Y=0.945 $X2=0 $Y2=0
cc_96 N_A_80_172#_c_82_n A1 0.00983782f $X=1.66 $Y=0.945 $X2=0 $Y2=0
cc_97 N_A_80_172#_c_89_n A1 0.0161012f $X=1.81 $Y=0.945 $X2=0 $Y2=0
cc_98 N_A_80_172#_c_89_n N_A1_c_226_n 0.00396977f $X=1.81 $Y=0.945 $X2=0 $Y2=0
cc_99 N_A_80_172#_c_83_n N_B1_c_272_n 0.00400966f $X=1.825 $Y=0.51 $X2=-0.19
+ $Y2=-0.245
cc_100 N_A_80_172#_c_93_n N_B1_M1004_g 0.00130701f $X=2.935 $Y=2.555 $X2=0 $Y2=0
cc_101 N_A_80_172#_c_84_n N_B1_c_273_n 0.0135692f $X=2.535 $Y=0.945 $X2=0 $Y2=0
cc_102 N_A_80_172#_c_84_n N_B1_c_274_n 0.00430735f $X=2.535 $Y=0.945 $X2=0 $Y2=0
cc_103 N_A_80_172#_c_91_n N_B1_c_274_n 0.00336963f $X=2.817 $Y=2.39 $X2=0 $Y2=0
cc_104 N_A_80_172#_c_93_n N_B1_c_280_n 0.00574649f $X=2.935 $Y=2.555 $X2=0 $Y2=0
cc_105 N_A_80_172#_c_84_n B1 0.028991f $X=2.535 $Y=0.945 $X2=0 $Y2=0
cc_106 N_A_80_172#_c_91_n B1 0.0514096f $X=2.817 $Y=2.39 $X2=0 $Y2=0
cc_107 N_A_80_172#_c_84_n N_B1_c_277_n 0.00365181f $X=2.535 $Y=0.945 $X2=0 $Y2=0
cc_108 N_A_80_172#_c_91_n N_B1_c_277_n 0.00574649f $X=2.817 $Y=2.39 $X2=0 $Y2=0
cc_109 N_A_80_172#_c_93_n N_C1_M1005_g 0.017677f $X=2.935 $Y=2.555 $X2=0 $Y2=0
cc_110 N_A_80_172#_c_91_n N_C1_M1005_g 0.0148351f $X=2.817 $Y=2.39 $X2=0 $Y2=0
cc_111 N_A_80_172#_c_85_n N_C1_M1000_g 0.0186783f $X=2.89 $Y=0.945 $X2=0 $Y2=0
cc_112 N_A_80_172#_c_86_n N_C1_M1000_g 0.00640471f $X=3.025 $Y=0.51 $X2=0 $Y2=0
cc_113 N_A_80_172#_c_91_n N_C1_M1000_g 0.00469272f $X=2.817 $Y=2.39 $X2=0 $Y2=0
cc_114 N_A_80_172#_c_85_n C1 0.0291901f $X=2.89 $Y=0.945 $X2=0 $Y2=0
cc_115 N_A_80_172#_c_93_n C1 0.0189312f $X=2.935 $Y=2.555 $X2=0 $Y2=0
cc_116 N_A_80_172#_c_91_n C1 0.0734562f $X=2.817 $Y=2.39 $X2=0 $Y2=0
cc_117 N_A_80_172#_c_85_n N_C1_c_320_n 0.00310262f $X=2.89 $Y=0.945 $X2=0 $Y2=0
cc_118 N_A_80_172#_c_93_n N_C1_c_320_n 0.00361823f $X=2.935 $Y=2.555 $X2=0 $Y2=0
cc_119 N_A_80_172#_c_91_n N_C1_c_320_n 0.0172031f $X=2.817 $Y=2.39 $X2=0 $Y2=0
cc_120 N_A_80_172#_M1007_g X 0.00675353f $X=0.48 $Y=0.51 $X2=0 $Y2=0
cc_121 N_A_80_172#_c_87_n X 0.0516251f $X=0.59 $Y=1.025 $X2=0 $Y2=0
cc_122 N_A_80_172#_c_88_n X 0.0392073f $X=0.59 $Y=1.025 $X2=0 $Y2=0
cc_123 N_A_80_172#_M1009_g X 0.00268913f $X=0.475 $Y=2.52 $X2=0 $Y2=0
cc_124 N_A_80_172#_M1009_g N_VPWR_c_361_n 0.00403818f $X=0.475 $Y=2.52 $X2=0
+ $Y2=0
cc_125 N_A_80_172#_c_81_n N_VPWR_c_361_n 0.00120509f $X=0.577 $Y=1.53 $X2=0
+ $Y2=0
cc_126 N_A_80_172#_c_87_n N_VPWR_c_361_n 0.00633123f $X=0.59 $Y=1.025 $X2=0
+ $Y2=0
cc_127 N_A_80_172#_M1009_g N_VPWR_c_363_n 0.0049405f $X=0.475 $Y=2.52 $X2=0
+ $Y2=0
cc_128 N_A_80_172#_c_93_n N_VPWR_c_365_n 0.0310803f $X=2.935 $Y=2.555 $X2=0
+ $Y2=0
cc_129 N_A_80_172#_M1009_g N_VPWR_c_360_n 0.00508379f $X=0.475 $Y=2.52 $X2=0
+ $Y2=0
cc_130 N_A_80_172#_c_93_n N_VPWR_c_360_n 0.0212581f $X=2.935 $Y=2.555 $X2=0
+ $Y2=0
cc_131 N_A_80_172#_c_91_n N_A_224_482#_c_402_n 0.0106472f $X=2.817 $Y=2.39 $X2=0
+ $Y2=0
cc_132 N_A_80_172#_M1009_g N_A_224_482#_c_403_n 0.00251973f $X=0.475 $Y=2.52
+ $X2=0 $Y2=0
cc_133 N_A_80_172#_c_93_n N_A_224_482#_c_404_n 4.68793e-19 $X=2.935 $Y=2.555
+ $X2=0 $Y2=0
cc_134 N_A_80_172#_c_91_n N_A_224_482#_c_404_n 0.0152055f $X=2.817 $Y=2.39 $X2=0
+ $Y2=0
cc_135 N_A_80_172#_c_93_n A_487_482# 0.00267342f $X=2.935 $Y=2.555 $X2=-0.19
+ $Y2=-0.245
cc_136 N_A_80_172#_M1007_g N_VGND_c_435_n 0.00522039f $X=0.48 $Y=0.51 $X2=0
+ $Y2=0
cc_137 N_A_80_172#_c_83_n N_VGND_c_436_n 0.0108858f $X=1.825 $Y=0.51 $X2=0 $Y2=0
cc_138 N_A_80_172#_c_86_n N_VGND_c_437_n 0.0121922f $X=3.025 $Y=0.51 $X2=0 $Y2=0
cc_139 N_A_80_172#_M1007_g N_VGND_c_438_n 0.00944742f $X=0.48 $Y=0.51 $X2=0
+ $Y2=0
cc_140 N_A_80_172#_c_82_n N_VGND_c_438_n 0.0152774f $X=1.66 $Y=0.945 $X2=0 $Y2=0
cc_141 N_A_80_172#_c_83_n N_VGND_c_438_n 0.0109142f $X=1.825 $Y=0.51 $X2=0 $Y2=0
cc_142 N_A_80_172#_c_84_n N_VGND_c_438_n 0.00593056f $X=2.535 $Y=0.945 $X2=0
+ $Y2=0
cc_143 N_A_80_172#_c_85_n N_VGND_c_438_n 0.00476608f $X=2.89 $Y=0.945 $X2=0
+ $Y2=0
cc_144 N_A_80_172#_c_86_n N_VGND_c_438_n 0.0110418f $X=3.025 $Y=0.51 $X2=0 $Y2=0
cc_145 N_A_80_172#_c_87_n N_VGND_c_438_n 0.00240067f $X=0.59 $Y=1.025 $X2=0
+ $Y2=0
cc_146 N_A_80_172#_c_90_n N_VGND_c_438_n 6.26195e-19 $X=2.62 $Y=0.945 $X2=0
+ $Y2=0
cc_147 N_A_80_172#_M1007_g N_VGND_c_439_n 0.00435313f $X=0.48 $Y=0.51 $X2=0
+ $Y2=0
cc_148 N_A_80_172#_c_82_n N_VGND_c_439_n 0.0309723f $X=1.66 $Y=0.945 $X2=0 $Y2=0
cc_149 N_A_80_172#_c_83_n N_VGND_c_439_n 0.0115491f $X=1.825 $Y=0.51 $X2=0 $Y2=0
cc_150 N_A_80_172#_c_87_n N_VGND_c_439_n 0.0132598f $X=0.59 $Y=1.025 $X2=0 $Y2=0
cc_151 N_A_80_172#_c_88_n N_VGND_c_439_n 0.00134059f $X=0.59 $Y=1.025 $X2=0
+ $Y2=0
cc_152 N_A_80_172#_c_84_n N_VGND_c_440_n 0.0283672f $X=2.535 $Y=0.945 $X2=0
+ $Y2=0
cc_153 N_A_80_172#_c_90_n N_VGND_c_440_n 0.0131175f $X=2.62 $Y=0.945 $X2=0 $Y2=0
cc_154 N_A2_M1001_g N_A1_M1002_g 0.0270012f $X=1.25 $Y=0.51 $X2=0 $Y2=0
cc_155 A2 N_A1_M1002_g 0.00229092f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_156 N_A2_c_172_n N_A1_c_224_n 0.0270012f $X=1.16 $Y=1.715 $X2=0 $Y2=0
cc_157 N_A2_c_175_n N_A1_c_228_n 0.00773926f $X=1.25 $Y=2.13 $X2=0 $Y2=0
cc_158 N_A2_c_179_n N_A1_M1006_g 0.00995889f $X=1.46 $Y=2.205 $X2=0 $Y2=0
cc_159 N_A2_c_178_n N_A1_c_230_n 0.0270012f $X=1.16 $Y=1.88 $X2=0 $Y2=0
cc_160 N_A2_c_179_n N_A1_c_231_n 0.00909055f $X=1.46 $Y=2.205 $X2=0 $Y2=0
cc_161 N_A2_M1001_g A1 0.00215688f $X=1.25 $Y=0.51 $X2=0 $Y2=0
cc_162 N_A2_c_175_n A1 2.12641e-19 $X=1.25 $Y=2.13 $X2=0 $Y2=0
cc_163 A2 A1 0.0532499f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_164 N_A2_c_174_n N_A1_c_226_n 0.0270012f $X=1.16 $Y=1.375 $X2=0 $Y2=0
cc_165 A2 X 0.00953226f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_166 N_A2_M1008_g N_VPWR_c_361_n 0.00311854f $X=1.46 $Y=2.73 $X2=0 $Y2=0
cc_167 N_A2_c_179_n N_VPWR_c_361_n 3.60095e-19 $X=1.46 $Y=2.205 $X2=0 $Y2=0
cc_168 N_A2_M1008_g N_VPWR_c_362_n 0.00292665f $X=1.46 $Y=2.73 $X2=0 $Y2=0
cc_169 N_A2_M1008_g N_VPWR_c_364_n 0.00540763f $X=1.46 $Y=2.73 $X2=0 $Y2=0
cc_170 N_A2_M1008_g N_VPWR_c_360_n 0.0112907f $X=1.46 $Y=2.73 $X2=0 $Y2=0
cc_171 N_A2_M1008_g N_A_224_482#_c_401_n 0.00438514f $X=1.46 $Y=2.73 $X2=0 $Y2=0
cc_172 N_A2_c_179_n N_A_224_482#_c_401_n 0.0074367f $X=1.46 $Y=2.205 $X2=0 $Y2=0
cc_173 N_A2_c_179_n N_A_224_482#_c_402_n 0.011294f $X=1.46 $Y=2.205 $X2=0 $Y2=0
cc_174 N_A2_c_175_n N_A_224_482#_c_403_n 0.00511184f $X=1.25 $Y=2.13 $X2=0 $Y2=0
cc_175 N_A2_c_178_n N_A_224_482#_c_403_n 7.38424e-19 $X=1.16 $Y=1.88 $X2=0 $Y2=0
cc_176 N_A2_c_179_n N_A_224_482#_c_403_n 0.0039632f $X=1.46 $Y=2.205 $X2=0 $Y2=0
cc_177 A2 N_A_224_482#_c_403_n 0.0219404f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_178 N_A2_M1001_g N_VGND_c_436_n 0.00435032f $X=1.25 $Y=0.51 $X2=0 $Y2=0
cc_179 N_A2_M1001_g N_VGND_c_438_n 0.00423597f $X=1.25 $Y=0.51 $X2=0 $Y2=0
cc_180 N_A2_M1001_g N_VGND_c_439_n 0.0123515f $X=1.25 $Y=0.51 $X2=0 $Y2=0
cc_181 N_A1_M1002_g N_B1_c_272_n 0.0186455f $X=1.61 $Y=0.51 $X2=-0.19 $Y2=-0.245
cc_182 N_A1_c_230_n N_B1_M1004_g 0.00743089f $X=1.715 $Y=1.89 $X2=0 $Y2=0
cc_183 N_A1_c_231_n N_B1_M1004_g 0.0168223f $X=1.93 $Y=2.195 $X2=0 $Y2=0
cc_184 N_A1_M1002_g N_B1_c_274_n 0.00774433f $X=1.61 $Y=0.51 $X2=0 $Y2=0
cc_185 N_A1_c_224_n N_B1_c_275_n 0.0136898f $X=1.715 $Y=1.71 $X2=0 $Y2=0
cc_186 N_A1_c_230_n N_B1_c_280_n 0.0136898f $X=1.715 $Y=1.89 $X2=0 $Y2=0
cc_187 A1 B1 0.0538866f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_188 N_A1_c_226_n B1 0.00427463f $X=1.73 $Y=1.385 $X2=0 $Y2=0
cc_189 A1 N_B1_c_277_n 6.14e-19 $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_190 N_A1_c_226_n N_B1_c_277_n 0.0136898f $X=1.73 $Y=1.385 $X2=0 $Y2=0
cc_191 N_A1_M1006_g N_VPWR_c_362_n 0.00282761f $X=1.93 $Y=2.73 $X2=0 $Y2=0
cc_192 N_A1_c_231_n N_VPWR_c_362_n 0.00268539f $X=1.93 $Y=2.195 $X2=0 $Y2=0
cc_193 N_A1_M1006_g N_VPWR_c_365_n 0.00540763f $X=1.93 $Y=2.73 $X2=0 $Y2=0
cc_194 N_A1_M1006_g N_VPWR_c_360_n 0.0103595f $X=1.93 $Y=2.73 $X2=0 $Y2=0
cc_195 N_A1_c_228_n N_A_224_482#_c_402_n 0.00645249f $X=1.82 $Y=2.12 $X2=0 $Y2=0
cc_196 N_A1_c_230_n N_A_224_482#_c_402_n 0.00146114f $X=1.715 $Y=1.89 $X2=0
+ $Y2=0
cc_197 N_A1_c_231_n N_A_224_482#_c_402_n 0.0142751f $X=1.93 $Y=2.195 $X2=0 $Y2=0
cc_198 A1 N_A_224_482#_c_402_n 0.0239282f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_199 N_A1_c_231_n N_A_224_482#_c_404_n 0.00283028f $X=1.93 $Y=2.195 $X2=0
+ $Y2=0
cc_200 N_A1_M1002_g N_VGND_c_436_n 0.0049163f $X=1.61 $Y=0.51 $X2=0 $Y2=0
cc_201 N_A1_M1002_g N_VGND_c_438_n 0.00559291f $X=1.61 $Y=0.51 $X2=0 $Y2=0
cc_202 N_A1_M1002_g N_VGND_c_439_n 0.00205649f $X=1.61 $Y=0.51 $X2=0 $Y2=0
cc_203 N_B1_c_280_n N_C1_M1005_g 0.0594062f $X=2.27 $Y=1.88 $X2=0 $Y2=0
cc_204 N_B1_c_272_n N_C1_M1000_g 0.0051077f $X=2.04 $Y=0.83 $X2=0 $Y2=0
cc_205 N_B1_c_273_n N_C1_M1000_g 0.00727848f $X=2.18 $Y=0.905 $X2=0 $Y2=0
cc_206 B1 N_C1_c_320_n 5.99772e-19 $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_207 N_B1_c_277_n N_C1_c_320_n 0.0594062f $X=2.27 $Y=1.375 $X2=0 $Y2=0
cc_208 N_B1_M1004_g N_VPWR_c_365_n 0.00540763f $X=2.36 $Y=2.73 $X2=0 $Y2=0
cc_209 N_B1_M1004_g N_VPWR_c_360_n 0.0103881f $X=2.36 $Y=2.73 $X2=0 $Y2=0
cc_210 N_B1_M1004_g N_A_224_482#_c_402_n 0.00193812f $X=2.36 $Y=2.73 $X2=0 $Y2=0
cc_211 N_B1_c_280_n N_A_224_482#_c_402_n 0.00132014f $X=2.27 $Y=1.88 $X2=0 $Y2=0
cc_212 B1 N_A_224_482#_c_402_n 0.0230572f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_213 N_B1_M1004_g N_A_224_482#_c_404_n 0.0022302f $X=2.36 $Y=2.73 $X2=0 $Y2=0
cc_214 N_B1_c_272_n N_VGND_c_436_n 0.00522039f $X=2.04 $Y=0.83 $X2=0 $Y2=0
cc_215 N_B1_c_272_n N_VGND_c_438_n 0.00601774f $X=2.04 $Y=0.83 $X2=0 $Y2=0
cc_216 N_B1_c_273_n N_VGND_c_438_n 4.11751e-19 $X=2.18 $Y=0.905 $X2=0 $Y2=0
cc_217 N_B1_c_272_n N_VGND_c_440_n 0.00423713f $X=2.04 $Y=0.83 $X2=0 $Y2=0
cc_218 N_B1_c_273_n N_VGND_c_440_n 0.00333081f $X=2.18 $Y=0.905 $X2=0 $Y2=0
cc_219 N_C1_M1005_g N_VPWR_c_365_n 0.00331542f $X=2.72 $Y=2.73 $X2=0 $Y2=0
cc_220 N_C1_M1005_g N_VPWR_c_360_n 0.00558484f $X=2.72 $Y=2.73 $X2=0 $Y2=0
cc_221 N_C1_M1000_g N_VGND_c_437_n 0.00522039f $X=2.81 $Y=0.51 $X2=0 $Y2=0
cc_222 N_C1_M1000_g N_VGND_c_438_n 0.00657786f $X=2.81 $Y=0.51 $X2=0 $Y2=0
cc_223 N_C1_M1000_g N_VGND_c_440_n 0.00423713f $X=2.81 $Y=0.51 $X2=0 $Y2=0
cc_224 X N_VPWR_c_361_n 0.00924417f $X=0.155 $Y=2.32 $X2=0 $Y2=0
cc_225 X N_VPWR_c_363_n 0.0108785f $X=0.24 $Y=2.405 $X2=0 $Y2=0
cc_226 X N_VPWR_c_360_n 0.0103432f $X=0.24 $Y=2.405 $X2=0 $Y2=0
cc_227 X N_VGND_c_435_n 0.0121529f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_228 X N_VGND_c_438_n 0.0108082f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_229 N_VPWR_c_361_n N_A_224_482#_c_401_n 0.056642f $X=0.69 $Y=2.345 $X2=0
+ $Y2=0
cc_230 N_VPWR_c_362_n N_A_224_482#_c_401_n 0.00229059f $X=1.685 $Y=2.565 $X2=0
+ $Y2=0
cc_231 N_VPWR_c_364_n N_A_224_482#_c_401_n 0.0207086f $X=1.55 $Y=3.33 $X2=0
+ $Y2=0
cc_232 N_VPWR_c_360_n N_A_224_482#_c_401_n 0.0115583f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_233 N_VPWR_c_362_n N_A_224_482#_c_402_n 0.023969f $X=1.685 $Y=2.565 $X2=0
+ $Y2=0
cc_234 N_VPWR_c_361_n N_A_224_482#_c_403_n 0.00360703f $X=0.69 $Y=2.345 $X2=0
+ $Y2=0
cc_235 N_VPWR_c_362_n N_A_224_482#_c_404_n 0.00267444f $X=1.685 $Y=2.565 $X2=0
+ $Y2=0
cc_236 N_VPWR_c_365_n N_A_224_482#_c_404_n 0.0188536f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_237 N_VPWR_c_360_n N_A_224_482#_c_404_n 0.0102248f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
