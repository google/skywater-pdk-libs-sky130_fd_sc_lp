* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
M1000 a_58_65# A1 VGND VNB nshort w=840000u l=150000u
+  ad=1.2096e+12p pd=1.128e+07u as=1.0584e+12p ps=7.56e+06u
M1001 a_58_65# B1 Y VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=2.352e+11p ps=2.24e+06u
M1002 VPWR A1 a_44_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=7.056e+11p pd=6.16e+06u as=1.0206e+12p ps=9.18e+06u
M1003 VGND A2 a_58_65# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_299_367# A2 a_44_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=8.064e+11p pd=6.32e+06u as=0p ps=0u
M1005 a_299_367# A3 Y VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=1.2159e+12p ps=9.49e+06u
M1006 Y A3 a_299_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 Y B1 VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND A3 a_58_65# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_44_367# A1 VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND A1 a_58_65# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 Y B1 a_58_65# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VPWR B1 Y VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_58_65# A3 VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_58_65# A2 VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_44_367# A2 a_299_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
