* File: sky130_fd_sc_lp__nor2b_lp.spice
* Created: Wed Sep  2 10:08:34 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__nor2b_lp.pex.spice"
.subckt sky130_fd_sc_lp__nor2b_lp  VNB VPB A B_N VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B_N	B_N
* A	A
* VPB	VPB
* VNB	VNB
MM1000 A_195_57# N_A_M1000_g N_VGND_M1000_s VNB NSHORT L=0.15 W=0.42 AD=0.0441
+ AS=0.1197 PD=0.63 PS=1.41 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2 SB=75002.1
+ A=0.063 P=1.14 MULT=1
MM1001 N_Y_M1001_d N_A_M1001_g A_195_57# VNB NSHORT L=0.15 W=0.42 AD=0.0588
+ AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6 SB=75001.8
+ A=0.063 P=1.14 MULT=1
MM1005 A_353_57# N_A_303_300#_M1005_g N_Y_M1001_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75001
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1002 N_VGND_M1002_d N_A_303_300#_M1002_g A_353_57# VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.4
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1006 A_511_57# N_B_N_M1006_g N_VGND_M1002_d VNB NSHORT L=0.15 W=0.42 AD=0.0441
+ AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75001.8 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1007 N_A_303_300#_M1007_d N_B_N_M1007_g A_511_57# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75002.1
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1004 A_255_408# N_A_M1004_g N_VPWR_M1004_s VPB PHIGHVT L=0.25 W=1 AD=0.12
+ AS=0.285 PD=1.24 PS=2.57 NRD=12.7853 NRS=0 M=1 R=4 SA=125000 SB=125001 A=0.25
+ P=2.5 MULT=1
MM1008 N_Y_M1008_d N_A_303_300#_M1008_g A_255_408# VPB PHIGHVT L=0.25 W=1
+ AD=0.285 AS=0.12 PD=2.57 PS=1.24 NRD=0 NRS=12.7853 M=1 R=4 SA=125001 SB=125000
+ A=0.25 P=2.5 MULT=1
MM1003 N_A_303_300#_M1003_d N_B_N_M1003_g N_VPWR_M1003_s VPB PHIGHVT L=0.25 W=1
+ AD=0.285 AS=0.285 PD=2.57 PS=2.57 NRD=0 NRS=0 M=1 R=4 SA=125000 SB=125000
+ A=0.25 P=2.5 MULT=1
DX9_noxref VNB VPB NWDIODE A=6.9751 P=11.21
c_64 VPB 0 1.57071e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_lp__nor2b_lp.pxi.spice"
*
.ends
*
*
