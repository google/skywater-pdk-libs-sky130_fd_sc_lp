* File: sky130_fd_sc_lp__clkinv_0.pex.spice
* Created: Wed Sep  2 09:40:13 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__CLKINV_0%A 3 7 9 10 11 12 18
r21 18 21 88.6355 $w=4.55e-07 $l=5.05e-07 $layer=POLY_cond $X=0.332 $Y=1.12
+ $X2=0.332 $Y2=1.625
r22 18 20 47.0767 $w=4.55e-07 $l=1.65e-07 $layer=POLY_cond $X=0.332 $Y=1.12
+ $X2=0.332 $Y2=0.955
r23 18 19 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.27
+ $Y=1.12 $X2=0.27 $Y2=1.12
r24 11 12 13.5366 $w=3.13e-07 $l=3.7e-07 $layer=LI1_cond $X=0.242 $Y=1.665
+ $X2=0.242 $Y2=2.035
r25 10 11 13.5366 $w=3.13e-07 $l=3.7e-07 $layer=LI1_cond $X=0.242 $Y=1.295
+ $X2=0.242 $Y2=1.665
r26 10 19 6.40246 $w=3.13e-07 $l=1.75e-07 $layer=LI1_cond $X=0.242 $Y=1.295
+ $X2=0.242 $Y2=1.12
r27 9 19 7.13417 $w=3.13e-07 $l=1.95e-07 $layer=LI1_cond $X=0.242 $Y=0.925
+ $X2=0.242 $Y2=1.12
r28 7 21 515.33 $w=1.5e-07 $l=1.005e-06 $layer=POLY_cond $X=0.485 $Y=2.63
+ $X2=0.485 $Y2=1.625
r29 3 20 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.485 $Y=0.56
+ $X2=0.485 $Y2=0.955
.ends

.subckt PM_SKY130_FD_SC_LP__CLKINV_0%VPWR 1 4 6 8 12 13
r13 16 17 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r14 12 13 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r15 10 16 4.4377 $w=1.7e-07 $l=2e-07 $layer=LI1_cond $X=0.4 $Y=3.33 $X2=0.2
+ $Y2=3.33
r16 10 12 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=0.4 $Y=3.33 $X2=0.72
+ $Y2=3.33
r17 8 13 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=0.48 $Y=3.33
+ $X2=0.72 $Y2=3.33
r18 8 17 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=0.48 $Y=3.33
+ $X2=0.24 $Y2=3.33
r19 4 16 3.03982 $w=2.95e-07 $l=1.07912e-07 $layer=LI1_cond $X=0.252 $Y=3.245
+ $X2=0.2 $Y2=3.33
r20 4 6 30.4714 $w=2.93e-07 $l=7.8e-07 $layer=LI1_cond $X=0.252 $Y=3.245
+ $X2=0.252 $Y2=2.465
r21 1 6 300 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_PDIFF $count=2 $X=0.145
+ $Y=2.31 $X2=0.27 $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__CLKINV_0%Y 1 2 9 11 12 13 14 15 16 41
r13 24 41 0.264495 $w=3.03e-07 $l=7e-09 $layer=LI1_cond $X=0.722 $Y=0.932
+ $X2=0.722 $Y2=0.925
r14 15 16 13.9805 $w=3.03e-07 $l=3.7e-07 $layer=LI1_cond $X=0.722 $Y=2.405
+ $X2=0.722 $Y2=2.775
r15 14 15 13.9805 $w=3.03e-07 $l=3.7e-07 $layer=LI1_cond $X=0.722 $Y=2.035
+ $X2=0.722 $Y2=2.405
r16 13 14 13.9805 $w=3.03e-07 $l=3.7e-07 $layer=LI1_cond $X=0.722 $Y=1.665
+ $X2=0.722 $Y2=2.035
r17 12 13 13.9805 $w=3.03e-07 $l=3.7e-07 $layer=LI1_cond $X=0.722 $Y=1.295
+ $X2=0.722 $Y2=1.665
r18 11 41 1.47362 $w=3.03e-07 $l=3.9e-08 $layer=LI1_cond $X=0.722 $Y=0.886
+ $X2=0.722 $Y2=0.925
r19 11 39 4.18518 $w=3.03e-07 $l=1.06e-07 $layer=LI1_cond $X=0.722 $Y=0.886
+ $X2=0.722 $Y2=0.78
r20 11 12 12.2423 $w=3.03e-07 $l=3.24e-07 $layer=LI1_cond $X=0.722 $Y=0.971
+ $X2=0.722 $Y2=1.295
r21 11 24 1.47362 $w=3.03e-07 $l=3.9e-08 $layer=LI1_cond $X=0.722 $Y=0.971
+ $X2=0.722 $Y2=0.932
r22 9 39 9.39028 $w=2.68e-07 $l=2.2e-07 $layer=LI1_cond $X=0.74 $Y=0.56 $X2=0.74
+ $Y2=0.78
r23 2 15 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=0.56
+ $Y=2.31 $X2=0.7 $Y2=2.455
r24 1 9 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.56
+ $Y=0.35 $X2=0.7 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_LP__CLKINV_0%VGND 1 4 6 8 12 13
r13 16 17 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r14 12 13 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r15 10 16 4.75569 $w=1.7e-07 $l=2.18e-07 $layer=LI1_cond $X=0.435 $Y=0 $X2=0.217
+ $Y2=0
r16 10 12 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.435 $Y=0 $X2=0.72
+ $Y2=0
r17 8 13 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=0.48 $Y=0 $X2=0.72
+ $Y2=0
r18 8 17 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=0.48 $Y=0 $X2=0.24
+ $Y2=0
r19 4 16 3.01048 $w=3.3e-07 $l=1.08305e-07 $layer=LI1_cond $X=0.27 $Y=0.085
+ $X2=0.217 $Y2=0
r20 4 6 16.0644 $w=3.28e-07 $l=4.6e-07 $layer=LI1_cond $X=0.27 $Y=0.085 $X2=0.27
+ $Y2=0.545
r21 1 6 182 $w=1.7e-07 $l=2.498e-07 $layer=licon1_NDIFF $count=1 $X=0.145
+ $Y=0.35 $X2=0.27 $Y2=0.545
.ends

