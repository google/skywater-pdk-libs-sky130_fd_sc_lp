* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__sdfxtp_lp CLK D SCD SCE VGND VNB VPB VPWR Q
M1000 a_457_417# D a_351_417# VPB phighvt w=1e+06u l=250000u
+  ad=2.2e+11p pd=2.44e+06u as=5.65e+11p ps=5.13e+06u
M1001 VGND a_2148_185# a_1910_155# VNB nshort w=420000u l=150000u
+  ad=8.911e+11p pd=9.43e+06u as=2.289e+11p ps=2.77e+06u
M1002 a_2628_69# a_2148_185# Q VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=1.197e+11p ps=1.41e+06u
M1003 a_351_417# D a_351_125# VNB nshort w=420000u l=150000u
+  ad=2.688e+11p pd=2.96e+06u as=1.008e+11p ps=1.32e+06u
M1004 a_978_66# a_733_66# VGND VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1005 VPWR SCE a_27_409# VPB phighvt w=1e+06u l=250000u
+  ad=2.185e+12p pd=1.637e+07u as=2.85e+11p ps=2.57e+06u
M1006 VPWR a_2148_185# Q VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=2.85e+11p ps=2.57e+06u
M1007 a_1528_347# a_733_66# a_1263_155# VPB phighvt w=1e+06u l=250000u
+  ad=2.4e+11p pd=2.48e+06u as=2.8e+11p ps=2.56e+06u
M1008 a_1957_347# a_733_66# a_1910_155# VNB nshort w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=0p ps=0u
M1009 a_351_417# a_733_66# a_1263_155# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=2.31e+11p ps=1.94e+06u
M1010 a_1576_99# a_998_347# a_1957_347# VNB nshort w=420000u l=150000u
+  ad=3.697e+11p pd=4.11e+06u as=0p ps=0u
M1011 a_351_417# a_27_409# a_244_417# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=5.7e+11p ps=5.14e+06u
M1012 a_998_347# a_733_66# VPWR VPB phighvt w=1e+06u l=250000u
+  ad=2.85e+11p pd=2.57e+06u as=0p ps=0u
M1013 a_2148_185# a_1957_347# a_2359_69# VNB nshort w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=8.82e+10p ps=1.26e+06u
M1014 a_244_417# SCD VPWR VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VGND SCE a_159_125# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1016 a_1576_99# a_1263_155# a_1722_125# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1017 a_1957_347# a_733_66# a_1576_99# VPB phighvt w=1e+06u l=250000u
+  ad=4.603e+11p pd=3.02e+06u as=4.5e+11p ps=2.9e+06u
M1018 a_820_66# CLK a_733_66# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=1.197e+11p ps=1.41e+06u
M1019 VGND SCD a_531_125# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.302e+11p ps=1.46e+06u
M1020 VGND CLK a_820_66# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_1263_155# a_998_347# a_351_417# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VPWR a_1576_99# a_1528_347# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_1263_155# a_998_347# a_1160_155# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=2.73e+11p ps=2.98e+06u
M1024 a_2359_69# a_1957_347# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_351_125# a_27_409# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 VPWR a_2148_185# a_2095_361# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=2.65e+11p ps=2.53e+06u
M1027 a_998_347# a_733_66# a_978_66# VNB nshort w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=0p ps=0u
M1028 a_1722_125# a_1263_155# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 VPWR CLK a_733_66# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=2.85e+11p ps=2.57e+06u
M1030 VPWR SCE a_457_417# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_2148_185# a_1957_347# VPWR VPB phighvt w=1e+06u l=250000u
+  ad=2.85e+11p pd=2.57e+06u as=0p ps=0u
M1032 a_159_125# SCE a_27_409# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1033 a_2095_361# a_998_347# a_1957_347# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1034 a_531_125# SCE a_351_417# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1035 VGND a_2148_185# a_2628_69# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1036 a_1576_99# a_1263_155# VPWR VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1037 VGND a_1576_99# a_1160_155# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
