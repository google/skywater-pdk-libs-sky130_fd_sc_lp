* File: sky130_fd_sc_lp__and4b_2.pex.spice
* Created: Fri Aug 28 10:08:33 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__AND4B_2%A_N 5 8 10 11 12 13 17 19
r25 17 19 45.5639 $w=3.95e-07 $l=1.65e-07 $layer=POLY_cond $X=0.352 $Y=0.98
+ $X2=0.352 $Y2=0.815
r26 12 13 12.5413 $w=3.38e-07 $l=3.7e-07 $layer=LI1_cond $X=0.255 $Y=0.925
+ $X2=0.255 $Y2=1.295
r27 12 17 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.32
+ $Y=0.98 $X2=0.32 $Y2=0.98
r28 10 11 43.452 $w=3.95e-07 $l=1.5e-07 $layer=POLY_cond $X=0.417 $Y=1.335
+ $X2=0.417 $Y2=1.485
r29 8 11 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=0.605 $Y=2.085 $X2=0.605
+ $Y2=1.485
r30 5 19 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.475 $Y=0.495
+ $X2=0.475 $Y2=0.815
r31 1 17 4.50555 $w=3.95e-07 $l=3.2e-08 $layer=POLY_cond $X=0.352 $Y=1.012
+ $X2=0.352 $Y2=0.98
r32 1 10 45.4779 $w=3.95e-07 $l=3.23e-07 $layer=POLY_cond $X=0.352 $Y=1.012
+ $X2=0.352 $Y2=1.335
.ends

.subckt PM_SKY130_FD_SC_LP__AND4B_2%A_53_375# 1 2 11 13 15 16 17 18 19 22 24 25
+ 28
c49 28 0 7.49265e-20 $X=1.09 $Y=0.35
c50 17 0 1.4653e-20 $X=1 $Y=1.12
r51 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.09
+ $Y=0.35 $X2=1.09 $Y2=0.35
r52 26 36 2.75184 $w=3.4e-07 $l=1e-07 $layer=LI1_cond $X=0.795 $Y=0.425
+ $X2=0.695 $Y2=0.425
r53 26 28 9.99914 $w=3.38e-07 $l=2.95e-07 $layer=LI1_cond $X=0.795 $Y=0.425
+ $X2=1.09 $Y2=0.425
r54 24 36 4.67813 $w=2e-07 $l=1.7e-07 $layer=LI1_cond $X=0.695 $Y=0.595
+ $X2=0.695 $Y2=0.425
r55 24 25 61 $w=1.98e-07 $l=1.1e-06 $layer=LI1_cond $X=0.695 $Y=0.595 $X2=0.695
+ $Y2=1.695
r56 20 25 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.35 $Y=1.78
+ $X2=0.695 $Y2=1.78
r57 20 22 10.1415 $w=2.48e-07 $l=2.2e-07 $layer=LI1_cond $X=0.35 $Y=1.865
+ $X2=0.35 $Y2=2.085
r58 19 29 50.7098 $w=3.3e-07 $l=2.9e-07 $layer=POLY_cond $X=1.38 $Y=0.35
+ $X2=1.09 $Y2=0.35
r59 17 18 43.7534 $w=2.2e-07 $l=1.5e-07 $layer=POLY_cond $X=1 $Y=1.12 $X2=1
+ $Y2=1.27
r60 16 29 8.74306 $w=3.3e-07 $l=5e-08 $layer=POLY_cond $X=1.04 $Y=0.35 $X2=1.09
+ $Y2=0.35
r61 13 19 32.1775 $w=3.3e-07 $l=1.98997e-07 $layer=POLY_cond $X=1.455 $Y=0.515
+ $X2=1.38 $Y2=0.35
r62 13 15 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.455 $Y=0.515
+ $X2=1.455 $Y2=0.835
r63 11 18 417.904 $w=1.5e-07 $l=8.15e-07 $layer=POLY_cond $X=1.035 $Y=2.085
+ $X2=1.035 $Y2=1.27
r64 7 16 32.1775 $w=3.3e-07 $l=1.98997e-07 $layer=POLY_cond $X=0.965 $Y=0.515
+ $X2=1.04 $Y2=0.35
r65 7 17 310.223 $w=1.5e-07 $l=6.05e-07 $layer=POLY_cond $X=0.965 $Y=0.515
+ $X2=0.965 $Y2=1.12
r66 2 22 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=0.265
+ $Y=1.875 $X2=0.39 $Y2=2.085
r67 1 36 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.285 $X2=0.69 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__AND4B_2%B 3 7 9 10 18
c30 7 0 7.49265e-20 $X=1.815 $Y=0.835
r31 16 18 25.3549 $w=3.3e-07 $l=1.45e-07 $layer=POLY_cond $X=1.67 $Y=1.55
+ $X2=1.815 $Y2=1.55
r32 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.67
+ $Y=1.55 $X2=1.67 $Y2=1.55
r33 13 16 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=1.465 $Y=1.55
+ $X2=1.67 $Y2=1.55
r34 10 17 5.09734 $w=2.58e-07 $l=1.15e-07 $layer=LI1_cond $X=1.705 $Y=1.665
+ $X2=1.705 $Y2=1.55
r35 9 17 11.3028 $w=2.58e-07 $l=2.55e-07 $layer=LI1_cond $X=1.705 $Y=1.295
+ $X2=1.705 $Y2=1.55
r36 5 18 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.815 $Y=1.385
+ $X2=1.815 $Y2=1.55
r37 5 7 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=1.815 $Y=1.385
+ $X2=1.815 $Y2=0.835
r38 1 13 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.465 $Y=1.715
+ $X2=1.465 $Y2=1.55
r39 1 3 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=1.465 $Y=1.715
+ $X2=1.465 $Y2=2.085
.ends

.subckt PM_SKY130_FD_SC_LP__AND4B_2%C 3 7 9 10 14
c33 9 0 9.72756e-20 $X=2.16 $Y=1.295
c34 3 0 1.03285e-19 $X=2.175 $Y=0.835
r35 14 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.265 $Y=1.375
+ $X2=2.265 $Y2=1.54
r36 14 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.265 $Y=1.375
+ $X2=2.265 $Y2=1.21
r37 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.265
+ $Y=1.375 $X2=2.265 $Y2=1.375
r38 10 15 9.6872 $w=3.43e-07 $l=2.9e-07 $layer=LI1_cond $X=2.177 $Y=1.665
+ $X2=2.177 $Y2=1.375
r39 9 15 2.67233 $w=3.43e-07 $l=8e-08 $layer=LI1_cond $X=2.177 $Y=1.295
+ $X2=2.177 $Y2=1.375
r40 7 17 279.457 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=2.355 $Y=2.085
+ $X2=2.355 $Y2=1.54
r41 3 16 192.287 $w=1.5e-07 $l=3.75e-07 $layer=POLY_cond $X=2.175 $Y=0.835
+ $X2=2.175 $Y2=1.21
.ends

.subckt PM_SKY130_FD_SC_LP__AND4B_2%D 3 7 9 12 13
c34 13 0 2.00264e-19 $X=2.805 $Y=1.375
c35 12 0 6.06973e-20 $X=2.805 $Y=1.375
c36 3 0 9.72756e-20 $X=2.715 $Y=0.835
r37 12 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.805 $Y=1.375
+ $X2=2.805 $Y2=1.54
r38 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.805 $Y=1.375
+ $X2=2.805 $Y2=1.21
r39 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.805
+ $Y=1.375 $X2=2.805 $Y2=1.375
r40 9 13 5.20967 $w=3.63e-07 $l=1.65e-07 $layer=LI1_cond $X=2.64 $Y=1.357
+ $X2=2.805 $Y2=1.357
r41 7 15 279.457 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=2.83 $Y=2.085
+ $X2=2.83 $Y2=1.54
r42 3 14 192.287 $w=1.5e-07 $l=3.75e-07 $layer=POLY_cond $X=2.715 $Y=0.835
+ $X2=2.715 $Y2=1.21
.ends

.subckt PM_SKY130_FD_SC_LP__AND4B_2%A_222_375# 1 2 3 12 16 20 24 26 28 30 34 36
+ 37 39 41 47 55
c104 12 0 9.69794e-20 $X=3.29 $Y=0.655
r105 54 55 11.366 $w=3.3e-07 $l=6.5e-08 $layer=POLY_cond $X=3.72 $Y=1.375
+ $X2=3.785 $Y2=1.375
r106 53 54 63.8244 $w=3.3e-07 $l=3.65e-07 $layer=POLY_cond $X=3.355 $Y=1.375
+ $X2=3.72 $Y2=1.375
r107 48 53 1.74861 $w=3.3e-07 $l=1e-08 $layer=POLY_cond $X=3.345 $Y=1.375
+ $X2=3.355 $Y2=1.375
r108 48 50 9.61737 $w=3.3e-07 $l=5.5e-08 $layer=POLY_cond $X=3.345 $Y=1.375
+ $X2=3.29 $Y2=1.375
r109 47 48 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.345
+ $Y=1.375 $X2=3.345 $Y2=1.375
r110 44 47 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=3.155 $Y=1.375
+ $X2=3.345 $Y2=1.375
r111 40 44 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.155 $Y=1.54
+ $X2=3.155 $Y2=1.375
r112 40 41 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=3.155 $Y=1.54
+ $X2=3.155 $Y2=1.71
r113 39 44 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.155 $Y=1.21
+ $X2=3.155 $Y2=1.375
r114 38 39 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=3.155 $Y=1.005
+ $X2=3.155 $Y2=1.21
r115 36 41 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.07 $Y=1.795
+ $X2=3.155 $Y2=1.71
r116 36 37 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=3.07 $Y=1.795
+ $X2=2.71 $Y2=1.795
r117 32 37 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=2.615 $Y=1.88
+ $X2=2.71 $Y2=1.795
r118 32 34 11.9665 $w=1.88e-07 $l=2.05e-07 $layer=LI1_cond $X=2.615 $Y=1.88
+ $X2=2.615 $Y2=2.085
r119 31 43 3.66393 $w=2.1e-07 $l=1.65e-07 $layer=LI1_cond $X=1.405 $Y=0.9
+ $X2=1.24 $Y2=0.9
r120 30 38 6.91519 $w=2.1e-07 $l=1.41244e-07 $layer=LI1_cond $X=3.07 $Y=0.9
+ $X2=3.155 $Y2=1.005
r121 30 31 87.9351 $w=2.08e-07 $l=1.665e-06 $layer=LI1_cond $X=3.07 $Y=0.9
+ $X2=1.405 $Y2=0.9
r122 26 43 3.21982 $w=2.5e-07 $l=1.2339e-07 $layer=LI1_cond $X=1.28 $Y=1.005
+ $X2=1.24 $Y2=0.9
r123 26 28 49.7855 $w=2.48e-07 $l=1.08e-06 $layer=LI1_cond $X=1.28 $Y=1.005
+ $X2=1.28 $Y2=2.085
r124 22 55 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.785 $Y=1.54
+ $X2=3.785 $Y2=1.375
r125 22 24 474.309 $w=1.5e-07 $l=9.25e-07 $layer=POLY_cond $X=3.785 $Y=1.54
+ $X2=3.785 $Y2=2.465
r126 18 54 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.72 $Y=1.21
+ $X2=3.72 $Y2=1.375
r127 18 20 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=3.72 $Y=1.21
+ $X2=3.72 $Y2=0.655
r128 14 53 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.355 $Y=1.54
+ $X2=3.355 $Y2=1.375
r129 14 16 474.309 $w=1.5e-07 $l=9.25e-07 $layer=POLY_cond $X=3.355 $Y=1.54
+ $X2=3.355 $Y2=2.465
r130 10 50 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.29 $Y=1.21
+ $X2=3.29 $Y2=1.375
r131 10 12 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=3.29 $Y=1.21
+ $X2=3.29 $Y2=0.655
r132 3 34 600 $w=1.7e-07 $l=2.8801e-07 $layer=licon1_PDIFF $count=1 $X=2.43
+ $Y=1.875 $X2=2.615 $Y2=2.085
r133 2 28 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=1.11
+ $Y=1.875 $X2=1.25 $Y2=2.085
r134 1 43 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=1.115
+ $Y=0.625 $X2=1.24 $Y2=0.9
.ends

.subckt PM_SKY130_FD_SC_LP__AND4B_2%VPWR 1 2 3 4 17 21 25 29 30 32 35 37 42 47
+ 53 56 59 63
r44 62 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r45 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r46 53 54 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r47 51 63 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r48 51 60 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=3.12 $Y2=3.33
r49 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r50 48 59 10.2049 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=3.305 $Y=3.33
+ $X2=3.092 $Y2=3.33
r51 48 50 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=3.305 $Y=3.33
+ $X2=3.6 $Y2=3.33
r52 47 62 4.58008 $w=1.7e-07 $l=2.17e-07 $layer=LI1_cond $X=3.885 $Y=3.33
+ $X2=4.102 $Y2=3.33
r53 47 50 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=3.885 $Y=3.33
+ $X2=3.6 $Y2=3.33
r54 46 60 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r55 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r56 43 56 13.9655 $w=1.7e-07 $l=3.65e-07 $layer=LI1_cond $X=2.305 $Y=3.33
+ $X2=1.94 $Y2=3.33
r57 43 45 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=2.305 $Y=3.33
+ $X2=2.64 $Y2=3.33
r58 42 59 10.2049 $w=1.7e-07 $l=2.12e-07 $layer=LI1_cond $X=2.88 $Y=3.33
+ $X2=3.092 $Y2=3.33
r59 42 45 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=2.88 $Y=3.33
+ $X2=2.64 $Y2=3.33
r60 41 54 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r61 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r62 38 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.985 $Y=3.33
+ $X2=0.82 $Y2=3.33
r63 38 40 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=0.985 $Y=3.33
+ $X2=1.2 $Y2=3.33
r64 37 56 13.9655 $w=1.7e-07 $l=3.65e-07 $layer=LI1_cond $X=1.575 $Y=3.33
+ $X2=1.94 $Y2=3.33
r65 37 40 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.575 $Y=3.33
+ $X2=1.2 $Y2=3.33
r66 35 46 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r67 35 41 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.2 $Y2=3.33
r68 35 56 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r69 30 62 3.06042 $w=3.15e-07 $l=1.11018e-07 $layer=LI1_cond $X=4.042 $Y=3.245
+ $X2=4.102 $Y2=3.33
r70 30 32 28.3538 $w=3.13e-07 $l=7.75e-07 $layer=LI1_cond $X=4.042 $Y=3.245
+ $X2=4.042 $Y2=2.47
r71 29 34 9.01032 $w=3.15e-07 $l=2.27e-07 $layer=LI1_cond $X=4.042 $Y=2.207
+ $X2=4.042 $Y2=1.98
r72 29 32 9.62198 $w=3.13e-07 $l=2.63e-07 $layer=LI1_cond $X=4.042 $Y=2.207
+ $X2=4.042 $Y2=2.47
r73 25 28 11.2533 $w=4.23e-07 $l=4.15e-07 $layer=LI1_cond $X=3.092 $Y=2.135
+ $X2=3.092 $Y2=2.55
r74 23 59 1.63918 $w=4.25e-07 $l=8.5e-08 $layer=LI1_cond $X=3.092 $Y=3.245
+ $X2=3.092 $Y2=3.33
r75 23 28 18.8458 $w=4.23e-07 $l=6.95e-07 $layer=LI1_cond $X=3.092 $Y=3.245
+ $X2=3.092 $Y2=2.55
r76 19 56 2.94957 $w=7.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.94 $Y=3.245
+ $X2=1.94 $Y2=3.33
r77 19 21 19.0062 $w=7.28e-07 $l=1.16e-06 $layer=LI1_cond $X=1.94 $Y=3.245
+ $X2=1.94 $Y2=2.085
r78 15 53 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.82 $Y=3.245
+ $X2=0.82 $Y2=3.33
r79 15 17 38.4148 $w=3.28e-07 $l=1.1e-06 $layer=LI1_cond $X=0.82 $Y=3.245
+ $X2=0.82 $Y2=2.145
r80 4 34 600 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=3.86
+ $Y=1.835 $X2=4.035 $Y2=1.98
r81 4 32 300 $w=1.7e-07 $l=7.01516e-07 $layer=licon1_PDIFF $count=2 $X=3.86
+ $Y=1.835 $X2=4 $Y2=2.47
r82 3 28 300 $w=1.7e-07 $l=7.83741e-07 $layer=licon1_PDIFF $count=2 $X=2.905
+ $Y=1.875 $X2=3.14 $Y2=2.55
r83 3 25 600 $w=1.7e-07 $l=3.2249e-07 $layer=licon1_PDIFF $count=1 $X=2.905
+ $Y=1.875 $X2=3.045 $Y2=2.135
r84 2 21 300 $w=1.7e-07 $l=6.97137e-07 $layer=licon1_PDIFF $count=2 $X=1.54
+ $Y=1.875 $X2=2.14 $Y2=2.085
r85 1 17 600 $w=1.7e-07 $l=3.32716e-07 $layer=licon1_PDIFF $count=1 $X=0.68
+ $Y=1.875 $X2=0.82 $Y2=2.145
.ends

.subckt PM_SKY130_FD_SC_LP__AND4B_2%X 1 2 9 14 16 17 18 19 20
c28 16 0 9.96393e-20 $X=3.627 $Y=1.71
r29 20 32 6.91466 $w=2.23e-07 $l=1.35e-07 $layer=LI1_cond $X=3.587 $Y=2.775
+ $X2=3.587 $Y2=2.91
r30 19 20 18.9513 $w=2.23e-07 $l=3.7e-07 $layer=LI1_cond $X=3.587 $Y=2.405
+ $X2=3.587 $Y2=2.775
r31 18 19 19.9757 $w=2.23e-07 $l=3.9e-07 $layer=LI1_cond $X=3.587 $Y=2.015
+ $X2=3.587 $Y2=2.405
r32 17 18 6.91466 $w=2.23e-07 $l=1.35e-07 $layer=LI1_cond $X=3.587 $Y=1.88
+ $X2=3.587 $Y2=2.015
r33 16 17 9.2015 $w=2.23e-07 $l=1.7e-07 $layer=LI1_cond $X=3.627 $Y=1.71
+ $X2=3.627 $Y2=1.88
r34 14 16 41.2828 $w=1.78e-07 $l=6.7e-07 $layer=LI1_cond $X=3.69 $Y=1.04
+ $X2=3.69 $Y2=1.71
r35 13 14 9.21974 $w=2.48e-07 $l=1.8e-07 $layer=LI1_cond $X=3.595 $Y=0.86
+ $X2=3.595 $Y2=1.04
r36 9 13 20.283 $w=2.48e-07 $l=4.4e-07 $layer=LI1_cond $X=3.535 $Y=0.42
+ $X2=3.535 $Y2=0.86
r37 2 32 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=3.43
+ $Y=1.835 $X2=3.57 $Y2=2.91
r38 2 18 400 $w=1.7e-07 $l=2.4e-07 $layer=licon1_PDIFF $count=1 $X=3.43 $Y=1.835
+ $X2=3.57 $Y2=2.015
r39 1 9 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=3.365
+ $Y=0.235 $X2=3.505 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__AND4B_2%VGND 1 2 3 10 12 16 18 21 24 26 27 29 37 46
+ 50
c53 12 0 1.4653e-20 $X=0.26 $Y=0.495
r54 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r55 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r56 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r57 41 50 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r58 41 47 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=3.12
+ $Y2=0
r59 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r60 38 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.24 $Y=0 $X2=3.075
+ $Y2=0
r61 38 40 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=3.24 $Y=0 $X2=3.6
+ $Y2=0
r62 37 49 5.09459 $w=1.7e-07 $l=2.45e-07 $layer=LI1_cond $X=3.83 $Y=0 $X2=4.075
+ $Y2=0
r63 37 40 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=3.83 $Y=0 $X2=3.6
+ $Y2=0
r64 36 47 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r65 35 36 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r66 33 44 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r67 32 35 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=0.72 $Y=0 $X2=2.64
+ $Y2=0
r68 32 33 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r69 30 43 4.78091 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=0 $X2=0.212
+ $Y2=0
r70 30 32 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.425 $Y=0 $X2=0.72
+ $Y2=0
r71 29 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.91 $Y=0 $X2=3.075
+ $Y2=0
r72 29 35 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=2.91 $Y=0 $X2=2.64
+ $Y2=0
r73 27 36 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r74 27 33 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=2.16 $Y=0 $X2=0.72
+ $Y2=0
r75 24 26 10.833 $w=2.48e-07 $l=2.35e-07 $layer=LI1_cond $X=4.075 $Y=0.925
+ $X2=4.075 $Y2=0.69
r76 19 26 6.98016 $w=3.68e-07 $l=1.85e-07 $layer=LI1_cond $X=4.015 $Y=0.505
+ $X2=4.015 $Y2=0.69
r77 19 21 3.89339 $w=3.68e-07 $l=1.25e-07 $layer=LI1_cond $X=4.015 $Y=0.505
+ $X2=4.015 $Y2=0.38
r78 18 49 3.01517 $w=3.7e-07 $l=1.11018e-07 $layer=LI1_cond $X=4.015 $Y=0.085
+ $X2=4.075 $Y2=0
r79 18 21 9.1884 $w=3.68e-07 $l=2.95e-07 $layer=LI1_cond $X=4.015 $Y=0.085
+ $X2=4.015 $Y2=0.38
r80 14 46 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.075 $Y=0.085
+ $X2=3.075 $Y2=0
r81 14 16 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=3.075 $Y=0.085
+ $X2=3.075 $Y2=0.5
r82 10 43 2.98526 $w=3.3e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.212 $Y2=0
r83 10 12 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.26 $Y2=0.495
r84 3 24 182 $w=1.7e-07 $l=8.01062e-07 $layer=licon1_NDIFF $count=1 $X=3.795
+ $Y=0.235 $X2=4.035 $Y2=0.925
r85 3 21 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=3.795
+ $Y=0.235 $X2=3.935 $Y2=0.38
r86 2 16 182 $w=1.7e-07 $l=3.41833e-07 $layer=licon1_NDIFF $count=1 $X=2.79
+ $Y=0.625 $X2=3.075 $Y2=0.5
r87 1 12 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.285 $X2=0.26 $Y2=0.495
.ends

