* NGSPICE file created from sky130_fd_sc_lp__nor2_lp2.ext - technology: sky130A

.subckt sky130_fd_sc_lp__nor2_lp2 A B VGND VNB VPB VPWR Y
M1000 a_130_112# A VGND VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=2.394e+11p ps=2.82e+06u
M1001 VGND B a_294_112# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1002 Y A a_130_112# VNB nshort w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=0p ps=0u
M1003 a_294_112# B Y VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 Y B a_134_374# VPB phighvt w=1e+06u l=250000u
+  ad=2.65e+11p pd=2.53e+06u as=2.1e+11p ps=2.42e+06u
M1005 a_134_374# A VPWR VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=2.85e+11p ps=2.57e+06u
.ends

