* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__a41o_lp A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
M1000 a_428_47# A1 a_314_47# VNB nshort w=420000u l=150000u
+  ad=1.764e+11p pd=1.68e+06u as=1.764e+11p ps=1.68e+06u
M1001 VPWR A2 a_27_409# VPB phighvt w=1e+06u l=250000u
+  ad=8.65e+11p pd=7.73e+06u as=8.45e+11p ps=7.69e+06u
M1002 VPWR A4 a_27_409# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_428_47# B1 a_27_409# VPB phighvt w=1e+06u l=250000u
+  ad=2.85e+11p pd=2.57e+06u as=0p ps=0u
M1004 VGND B1 a_542_47# VNB nshort w=420000u l=150000u
+  ad=2.373e+11p pd=2.81e+06u as=8.82e+10p ps=1.26e+06u
M1005 a_206_47# A3 a_128_47# VNB nshort w=420000u l=150000u
+  ad=1.638e+11p pd=1.62e+06u as=1.008e+11p ps=1.32e+06u
M1006 a_27_409# A3 VPWR VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_314_47# A2 a_206_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_542_47# B1 a_428_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_700_47# a_428_47# VGND VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1010 a_128_47# A4 VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 X a_428_47# a_700_47# VNB nshort w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=0p ps=0u
M1012 a_27_409# A1 VPWR VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1013 X a_428_47# VPWR VPB phighvt w=1e+06u l=250000u
+  ad=2.85e+11p pd=2.57e+06u as=0p ps=0u
.ends
