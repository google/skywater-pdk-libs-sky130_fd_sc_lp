* File: sky130_fd_sc_lp__o21a_4.spice
* Created: Wed Sep  2 10:15:27 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__o21a_4.pex.spice"
.subckt sky130_fd_sc_lp__o21a_4  VNB VPB B1 A1 A2 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A2	A2
* A1	A1
* B1	B1
* VPB	VPB
* VNB	VNB
MM1001 N_X_M1001_d N_A_90_23#_M1001_g N_VGND_M1001_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75001.5 A=0.126 P=1.98 MULT=1
MM1003 N_X_M1001_d N_A_90_23#_M1003_g N_VGND_M1003_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1004 N_X_M1004_d N_A_90_23#_M1004_g N_VGND_M1003_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.1
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1010 N_X_M1004_d N_A_90_23#_M1010_g N_VGND_M1010_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75001.5
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1007 N_A_90_23#_M1007_d N_B1_M1007_g N_A_485_65#_M1007_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.3066 PD=1.12 PS=2.41 NRD=0 NRS=9.996 M=1 R=5.6
+ SA=75000.3 SB=75002.5 A=0.126 P=1.98 MULT=1
MM1013 N_A_90_23#_M1007_d N_B1_M1013_g N_A_485_65#_M1013_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1512 PD=1.12 PS=1.2 NRD=0 NRS=11.424 M=1 R=5.6
+ SA=75000.7 SB=75002.1 A=0.126 P=1.98 MULT=1
MM1016 N_A_485_65#_M1013_s N_A1_M1016_g N_VGND_M1016_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1512 AS=0.1512 PD=1.2 PS=1.2 NRD=0 NRS=9.996 M=1 R=5.6 SA=75001.2
+ SB=75001.6 A=0.126 P=1.98 MULT=1
MM1005 N_A_485_65#_M1005_d N_A2_M1005_g N_VGND_M1016_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1512 PD=1.12 PS=1.2 NRD=0 NRS=1.428 M=1 R=5.6 SA=75001.7
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1011 N_A_485_65#_M1005_d N_A2_M1011_g N_VGND_M1011_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002.2
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1019 N_A_485_65#_M1019_d N_A1_M1019_g N_VGND_M1011_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002.6
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1002 N_VPWR_M1002_d N_A_90_23#_M1002_g N_X_M1002_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75004.5 A=0.189 P=2.82 MULT=1
MM1009 N_VPWR_M1009_d N_A_90_23#_M1009_g N_X_M1002_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75004.1 A=0.189 P=2.82 MULT=1
MM1012 N_VPWR_M1009_d N_A_90_23#_M1012_g N_X_M1012_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75003.7 A=0.189 P=2.82 MULT=1
MM1018 N_VPWR_M1018_d N_A_90_23#_M1018_g N_X_M1012_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.5
+ SB=75003.2 A=0.189 P=2.82 MULT=1
MM1008 N_VPWR_M1018_d N_B1_M1008_g N_A_90_23#_M1008_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.9
+ SB=75002.8 A=0.189 P=2.82 MULT=1
MM1017 N_VPWR_M1017_d N_B1_M1017_g N_A_90_23#_M1008_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.4662 AS=0.1764 PD=2 PS=1.54 NRD=20.8426 NRS=0 M=1 R=8.4 SA=75002.3
+ SB=75002.4 A=0.189 P=2.82 MULT=1
MM1000 N_A_792_367#_M1000_d N_A1_M1000_g N_VPWR_M1017_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.4662 PD=1.54 PS=2 NRD=0 NRS=27.0875 M=1 R=8.4 SA=75003.2
+ SB=75001.5 A=0.189 P=2.82 MULT=1
MM1006 N_A_792_367#_M1000_d N_A2_M1006_g N_A_90_23#_M1006_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75003.7
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1014 N_A_792_367#_M1014_d N_A2_M1014_g N_A_90_23#_M1006_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75004.1
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1015 N_A_792_367#_M1014_d N_A1_M1015_g N_VPWR_M1015_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75004.5
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX20_noxref VNB VPB NWDIODE A=11.4511 P=16.01
c_55 VNB 0 5.42069e-20 $X=0 $Y=0
*
.include "sky130_fd_sc_lp__o21a_4.pxi.spice"
*
.ends
*
*
