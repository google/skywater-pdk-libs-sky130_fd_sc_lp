* File: sky130_fd_sc_lp__ha_m.spice
* Created: Fri Aug 28 10:36:53 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__ha_m.pex.spice"
.subckt sky130_fd_sc_lp__ha_m  VNB VPB B A SUM VPWR COUT VGND
* 
* VGND	VGND
* COUT	COUT
* VPWR	VPWR
* SUM	SUM
* A	A
* B	B
* VPB	VPB
* VNB	VNB
MM1001 N_VGND_M1001_d N_A_80_60#_M1001_g N_SUM_M1001_s VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.1113 PD=1.37 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1011 N_A_301_47#_M1011_d N_A_249_212#_M1011_g N_A_80_60#_M1011_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.2 A=0.063 P=1.14 MULT=1
MM1006 N_VGND_M1006_d N_B_M1006_g N_A_301_47#_M1011_d VNB NSHORT L=0.15 W=0.42
+ AD=0.09675 AS=0.0588 PD=0.89 PS=0.7 NRD=22.848 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.8 A=0.063 P=1.14 MULT=1
MM1007 N_A_301_47#_M1007_d N_A_M1007_g N_VGND_M1006_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.09675 PD=1.37 PS=0.89 NRD=0 NRS=22.848 M=1 R=2.8 SA=75001.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1005 A_720_125# N_B_M1005_g N_A_249_212#_M1005_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1512 PD=0.63 PS=1.56 NRD=14.28 NRS=27.132 M=1 R=2.8 SA=75000.3
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1000 N_VGND_M1000_d N_A_M1000_g A_720_125# VNB NSHORT L=0.15 W=0.42 AD=0.0588
+ AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1010 N_COUT_M1010_d N_A_249_212#_M1010_g N_VGND_M1000_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.1
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1002 N_VPWR_M1002_d N_A_80_60#_M1002_g N_SUM_M1002_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.09555 AS=0.1113 PD=0.875 PS=1.37 NRD=9.3772 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.2 A=0.063 P=1.14 MULT=1
MM1003 N_A_80_60#_M1003_d N_A_249_212#_M1003_g N_VPWR_M1002_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0588 AS=0.09555 PD=0.7 PS=0.875 NRD=0 NRS=72.693 M=1 R=2.8
+ SA=75000.8 SB=75001.6 A=0.063 P=1.14 MULT=1
MM1012 A_450_464# N_B_M1012_g N_A_80_60#_M1003_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0672 AS=0.0588 PD=0.74 PS=0.7 NRD=49.25 NRS=0 M=1 R=2.8 SA=75001.2
+ SB=75001.2 A=0.063 P=1.14 MULT=1
MM1009 N_VPWR_M1009_d N_A_M1009_g A_450_464# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.136825 AS=0.0672 PD=1.195 PS=0.74 NRD=44.5417 NRS=49.25 M=1 R=2.8
+ SA=75001.7 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1013 N_A_249_212#_M1013_d N_B_M1013_g N_VPWR_M1009_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0987 AS=0.136825 PD=0.89 PS=1.195 NRD=44.5417 NRS=126.986 M=1 R=2.8
+ SA=75000.8 SB=75001.2 A=0.063 P=1.14 MULT=1
MM1008 N_VPWR_M1008_d N_A_M1008_g N_A_249_212#_M1013_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0588 AS=0.0987 PD=0.7 PS=0.89 NRD=0 NRS=44.5417 M=1 R=2.8 SA=75001.5
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1004 N_COUT_M1004_d N_A_249_212#_M1004_g N_VPWR_M1008_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.9
+ SB=75000.2 A=0.063 P=1.14 MULT=1
DX14_noxref VNB VPB NWDIODE A=9.6607 P=14.09
c_95 VPB 0 1.9418e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_lp__ha_m.pxi.spice"
*
.ends
*
*
