* File: sky130_fd_sc_lp__nand4bb_lp.pxi.spice
* Created: Wed Sep  2 10:07:01 2020
* 
x_PM_SKY130_FD_SC_LP__NAND4BB_LP%A_N N_A_N_M1002_g N_A_N_M1008_g N_A_N_M1011_g
+ N_A_N_c_83_n N_A_N_c_84_n A_N N_A_N_c_85_n N_A_N_c_86_n
+ PM_SKY130_FD_SC_LP__NAND4BB_LP%A_N
x_PM_SKY130_FD_SC_LP__NAND4BB_LP%A_27_47# N_A_27_47#_M1002_s N_A_27_47#_M1008_s
+ N_A_27_47#_c_134_n N_A_27_47#_M1000_g N_A_27_47#_c_125_n N_A_27_47#_c_126_n
+ N_A_27_47#_c_127_n N_A_27_47#_M1003_g N_A_27_47#_c_128_n N_A_27_47#_c_129_n
+ N_A_27_47#_c_130_n N_A_27_47#_c_138_n N_A_27_47#_c_139_n N_A_27_47#_c_131_n
+ N_A_27_47#_c_132_n N_A_27_47#_c_133_n N_A_27_47#_c_140_n
+ PM_SKY130_FD_SC_LP__NAND4BB_LP%A_27_47#
x_PM_SKY130_FD_SC_LP__NAND4BB_LP%A_332_352# N_A_332_352#_M1001_d
+ N_A_332_352#_M1010_d N_A_332_352#_c_206_n N_A_332_352#_M1009_g
+ N_A_332_352#_M1005_g N_A_332_352#_c_208_n N_A_332_352#_c_209_n
+ N_A_332_352#_c_210_n N_A_332_352#_c_211_n N_A_332_352#_c_212_n
+ N_A_332_352#_c_213_n PM_SKY130_FD_SC_LP__NAND4BB_LP%A_332_352#
x_PM_SKY130_FD_SC_LP__NAND4BB_LP%C N_C_M1004_g N_C_M1006_g C N_C_c_281_n
+ N_C_c_284_n PM_SKY130_FD_SC_LP__NAND4BB_LP%C
x_PM_SKY130_FD_SC_LP__NAND4BB_LP%D N_D_c_322_n N_D_M1013_g N_D_M1012_g
+ N_D_c_323_n D N_D_c_324_n N_D_c_325_n N_D_c_326_n
+ PM_SKY130_FD_SC_LP__NAND4BB_LP%D
x_PM_SKY130_FD_SC_LP__NAND4BB_LP%B_N N_B_N_c_368_n N_B_N_M1007_g N_B_N_M1010_g
+ N_B_N_c_370_n N_B_N_M1001_g B_N B_N B_N N_B_N_c_372_n
+ PM_SKY130_FD_SC_LP__NAND4BB_LP%B_N
x_PM_SKY130_FD_SC_LP__NAND4BB_LP%VPWR N_VPWR_M1008_d N_VPWR_M1009_d
+ N_VPWR_M1012_d N_VPWR_c_409_n N_VPWR_c_410_n N_VPWR_c_411_n N_VPWR_c_412_n
+ N_VPWR_c_413_n N_VPWR_c_414_n N_VPWR_c_415_n VPWR N_VPWR_c_416_n
+ N_VPWR_c_417_n N_VPWR_c_408_n N_VPWR_c_419_n
+ PM_SKY130_FD_SC_LP__NAND4BB_LP%VPWR
x_PM_SKY130_FD_SC_LP__NAND4BB_LP%Y N_Y_M1003_s N_Y_M1000_d N_Y_M1004_d
+ N_Y_c_473_n N_Y_c_496_n N_Y_c_476_n N_Y_c_477_n N_Y_c_507_n N_Y_c_488_n
+ N_Y_c_474_n N_Y_c_509_n Y PM_SKY130_FD_SC_LP__NAND4BB_LP%Y
x_PM_SKY130_FD_SC_LP__NAND4BB_LP%VGND N_VGND_M1011_d N_VGND_M1013_d
+ N_VGND_c_540_n N_VGND_c_541_n VGND N_VGND_c_542_n N_VGND_c_543_n
+ N_VGND_c_544_n N_VGND_c_545_n N_VGND_c_546_n N_VGND_c_547_n
+ PM_SKY130_FD_SC_LP__NAND4BB_LP%VGND
cc_1 VNB N_A_N_M1002_g 0.0236161f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.445
cc_2 VNB N_A_N_M1011_g 0.0219604f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=0.445
cc_3 VNB N_A_N_c_83_n 0.0221011f $X=-0.19 $Y=-0.245 $X2=0.675 $Y2=0.985
cc_4 VNB N_A_N_c_84_n 0.0296113f $X=-0.19 $Y=-0.245 $X2=0.607 $Y2=1.338
cc_5 VNB N_A_N_c_85_n 0.0286479f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.02
cc_6 VNB N_A_N_c_86_n 0.00669918f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.02
cc_7 VNB N_A_27_47#_c_125_n 0.0352297f $X=-0.19 $Y=-0.245 $X2=0.607 $Y2=0.985
cc_8 VNB N_A_27_47#_c_126_n 0.0111957f $X=-0.19 $Y=-0.245 $X2=0.675 $Y2=0.835
cc_9 VNB N_A_27_47#_c_127_n 0.0170458f $X=-0.19 $Y=-0.245 $X2=0.675 $Y2=0.985
cc_10 VNB N_A_27_47#_c_128_n 0.0228304f $X=-0.19 $Y=-0.245 $X2=0.607 $Y2=1.02
cc_11 VNB N_A_27_47#_c_129_n 0.0199343f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.02
cc_12 VNB N_A_27_47#_c_130_n 0.0463979f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=1.02
cc_13 VNB N_A_27_47#_c_131_n 0.00370033f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_27_47#_c_132_n 0.0177285f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_27_47#_c_133_n 0.0209565f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_332_352#_c_206_n 0.0585696f $X=-0.19 $Y=-0.245 $X2=0.725 $Y2=2.595
cc_17 VNB N_A_332_352#_M1005_g 0.0347546f $X=-0.19 $Y=-0.245 $X2=0.607 $Y2=0.985
cc_18 VNB N_A_332_352#_c_208_n 0.0391906f $X=-0.19 $Y=-0.245 $X2=0.675 $Y2=0.985
cc_19 VNB N_A_332_352#_c_209_n 0.00971342f $X=-0.19 $Y=-0.245 $X2=0.607 $Y2=1.02
cc_20 VNB N_A_332_352#_c_210_n 0.0321883f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=1.02
cc_21 VNB N_A_332_352#_c_211_n 0.00727708f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=1.295
cc_22 VNB N_A_332_352#_c_212_n 0.010604f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_332_352#_c_213_n 0.01116f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_C_M1006_g 0.0582132f $X=-0.19 $Y=-0.245 $X2=0.725 $Y2=2.595
cc_25 VNB N_C_c_281_n 0.00796247f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_D_c_322_n 0.0145939f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.835
cc_27 VNB N_D_c_323_n 0.0145301f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_D_c_324_n 0.00777394f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_29 VNB N_D_c_325_n 4.80315e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_D_c_326_n 0.0388139f $X=-0.19 $Y=-0.245 $X2=0.607 $Y2=1.02
cc_31 VNB N_B_N_c_368_n 0.0159945f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.835
cc_32 VNB N_B_N_M1010_g 0.0435283f $X=-0.19 $Y=-0.245 $X2=0.725 $Y2=2.595
cc_33 VNB N_B_N_c_370_n 0.0185969f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB B_N 0.010963f $X=-0.19 $Y=-0.245 $X2=0.607 $Y2=0.985
cc_35 VNB N_B_N_c_372_n 0.0373839f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VPWR_c_408_n 0.183584f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_Y_c_473_n 0.00962766f $X=-0.19 $Y=-0.245 $X2=0.607 $Y2=0.985
cc_38 VNB N_Y_c_474_n 0.00503528f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_540_n 0.0152298f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=0.835
cc_40 VNB N_VGND_c_541_n 0.0028319f $X=-0.19 $Y=-0.245 $X2=0.607 $Y2=0.985
cc_41 VNB N_VGND_c_542_n 0.0268694f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_42 VNB N_VGND_c_543_n 0.0531396f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=1.02
cc_43 VNB N_VGND_c_544_n 0.0296796f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_545_n 0.235103f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_546_n 0.00513431f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_547_n 0.00510792f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VPB N_A_N_M1008_g 0.0500483f $X=-0.19 $Y=1.655 $X2=0.725 $Y2=2.595
cc_48 VPB N_A_27_47#_c_134_n 0.0120099f $X=-0.19 $Y=1.655 $X2=0.725 $Y2=2.595
cc_49 VPB N_A_27_47#_M1000_g 0.0281349f $X=-0.19 $Y=1.655 $X2=0.855 $Y2=0.835
cc_50 VPB N_A_27_47#_c_129_n 0.00535533f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=1.02
cc_51 VPB N_A_27_47#_c_130_n 0.00332766f $X=-0.19 $Y=1.655 $X2=0.65 $Y2=1.02
cc_52 VPB N_A_27_47#_c_138_n 0.0568014f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_53 VPB N_A_27_47#_c_139_n 0.0124129f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_54 VPB N_A_27_47#_c_140_n 0.0157504f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_55 VPB N_A_332_352#_c_206_n 0.0307515f $X=-0.19 $Y=1.655 $X2=0.725 $Y2=2.595
cc_56 VPB N_A_332_352#_M1009_g 0.0296551f $X=-0.19 $Y=1.655 $X2=0.855 $Y2=0.835
cc_57 VPB N_A_332_352#_c_209_n 0.0592826f $X=-0.19 $Y=1.655 $X2=0.607 $Y2=1.02
cc_58 VPB N_A_332_352#_c_211_n 0.00309745f $X=-0.19 $Y=1.655 $X2=0.65 $Y2=1.295
cc_59 VPB N_C_M1004_g 0.0264492f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=0.445
cc_60 VPB N_C_c_281_n 0.0235645f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_61 VPB N_C_c_284_n 0.00233215f $X=-0.19 $Y=1.655 $X2=0.607 $Y2=0.985
cc_62 VPB N_D_M1012_g 0.0241587f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_63 VPB N_D_c_324_n 0.0199423f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_64 VPB N_D_c_325_n 0.00424591f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_65 VPB N_B_N_M1010_g 0.0508518f $X=-0.19 $Y=1.655 $X2=0.725 $Y2=2.595
cc_66 VPB N_VPWR_c_409_n 0.00303789f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_67 VPB N_VPWR_c_410_n 0.00284591f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_411_n 0.00283153f $X=-0.19 $Y=1.655 $X2=0.65 $Y2=1.02
cc_69 VPB N_VPWR_c_412_n 0.022663f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_70 VPB N_VPWR_c_413_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_71 VPB N_VPWR_c_414_n 0.0289584f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_72 VPB N_VPWR_c_415_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_73 VPB N_VPWR_c_416_n 0.0180468f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_74 VPB N_VPWR_c_417_n 0.0220452f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_75 VPB N_VPWR_c_408_n 0.0481588f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_76 VPB N_VPWR_c_419_n 0.00511011f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_77 VPB N_Y_c_473_n 0.00190992f $X=-0.19 $Y=1.655 $X2=0.607 $Y2=0.985
cc_78 VPB N_Y_c_476_n 0.00451704f $X=-0.19 $Y=1.655 $X2=0.607 $Y2=1.338
cc_79 VPB N_Y_c_477_n 0.00176929f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_80 N_A_N_M1008_g N_A_27_47#_c_134_n 0.0104189f $X=0.725 $Y=2.595 $X2=0 $Y2=0
cc_81 N_A_N_M1008_g N_A_27_47#_M1000_g 0.0158144f $X=0.725 $Y=2.595 $X2=0 $Y2=0
cc_82 N_A_N_M1011_g N_A_27_47#_c_126_n 0.00524362f $X=0.855 $Y=0.445 $X2=0 $Y2=0
cc_83 N_A_N_c_86_n N_A_27_47#_c_126_n 6.72006e-19 $X=0.63 $Y=1.02 $X2=0 $Y2=0
cc_84 N_A_N_c_83_n N_A_27_47#_c_128_n 0.00524362f $X=0.675 $Y=0.985 $X2=0 $Y2=0
cc_85 N_A_N_c_85_n N_A_27_47#_c_128_n 0.00486487f $X=0.63 $Y=1.02 $X2=0 $Y2=0
cc_86 N_A_N_c_86_n N_A_27_47#_c_128_n 0.00454663f $X=0.63 $Y=1.02 $X2=0 $Y2=0
cc_87 N_A_N_c_84_n N_A_27_47#_c_129_n 0.0165389f $X=0.607 $Y=1.338 $X2=0 $Y2=0
cc_88 N_A_N_M1002_g N_A_27_47#_c_130_n 0.0210338f $X=0.495 $Y=0.445 $X2=0 $Y2=0
cc_89 N_A_N_c_84_n N_A_27_47#_c_130_n 0.00465147f $X=0.607 $Y=1.338 $X2=0 $Y2=0
cc_90 N_A_N_c_86_n N_A_27_47#_c_130_n 0.0485802f $X=0.63 $Y=1.02 $X2=0 $Y2=0
cc_91 N_A_N_M1008_g N_A_27_47#_c_138_n 0.0313747f $X=0.725 $Y=2.595 $X2=0 $Y2=0
cc_92 N_A_N_M1008_g N_A_27_47#_c_139_n 0.0181653f $X=0.725 $Y=2.595 $X2=0 $Y2=0
cc_93 N_A_N_c_86_n N_A_27_47#_c_139_n 0.0139211f $X=0.63 $Y=1.02 $X2=0 $Y2=0
cc_94 N_A_N_c_84_n N_A_27_47#_c_131_n 0.00135187f $X=0.607 $Y=1.338 $X2=0 $Y2=0
cc_95 N_A_N_c_85_n N_A_27_47#_c_131_n 3.60319e-19 $X=0.63 $Y=1.02 $X2=0 $Y2=0
cc_96 N_A_N_c_86_n N_A_27_47#_c_131_n 0.017691f $X=0.63 $Y=1.02 $X2=0 $Y2=0
cc_97 N_A_N_c_85_n N_A_27_47#_c_132_n 0.00612007f $X=0.63 $Y=1.02 $X2=0 $Y2=0
cc_98 N_A_N_c_86_n N_A_27_47#_c_132_n 0.0020313f $X=0.63 $Y=1.02 $X2=0 $Y2=0
cc_99 N_A_N_M1002_g N_A_27_47#_c_133_n 0.00850743f $X=0.495 $Y=0.445 $X2=0 $Y2=0
cc_100 N_A_N_M1011_g N_A_27_47#_c_133_n 0.00111595f $X=0.855 $Y=0.445 $X2=0
+ $Y2=0
cc_101 N_A_N_M1008_g N_A_27_47#_c_140_n 0.00459948f $X=0.725 $Y=2.595 $X2=0
+ $Y2=0
cc_102 N_A_N_c_84_n N_A_27_47#_c_140_n 0.00318244f $X=0.607 $Y=1.338 $X2=0 $Y2=0
cc_103 N_A_N_c_86_n N_A_27_47#_c_140_n 0.012405f $X=0.63 $Y=1.02 $X2=0 $Y2=0
cc_104 N_A_N_M1008_g N_VPWR_c_409_n 0.0239789f $X=0.725 $Y=2.595 $X2=0 $Y2=0
cc_105 N_A_N_M1008_g N_VPWR_c_412_n 0.00840199f $X=0.725 $Y=2.595 $X2=0 $Y2=0
cc_106 N_A_N_M1008_g N_VPWR_c_408_n 0.0146481f $X=0.725 $Y=2.595 $X2=0 $Y2=0
cc_107 N_A_N_M1011_g N_Y_c_473_n 0.00164942f $X=0.855 $Y=0.445 $X2=0 $Y2=0
cc_108 N_A_N_M1011_g N_Y_c_474_n 7.88281e-19 $X=0.855 $Y=0.445 $X2=0 $Y2=0
cc_109 N_A_N_M1002_g N_VGND_c_540_n 0.00239794f $X=0.495 $Y=0.445 $X2=0 $Y2=0
cc_110 N_A_N_M1011_g N_VGND_c_540_n 0.0150927f $X=0.855 $Y=0.445 $X2=0 $Y2=0
cc_111 N_A_N_M1002_g N_VGND_c_542_n 0.00549284f $X=0.495 $Y=0.445 $X2=0 $Y2=0
cc_112 N_A_N_M1011_g N_VGND_c_542_n 0.00486043f $X=0.855 $Y=0.445 $X2=0 $Y2=0
cc_113 N_A_N_M1002_g N_VGND_c_545_n 0.00784569f $X=0.495 $Y=0.445 $X2=0 $Y2=0
cc_114 N_A_N_M1011_g N_VGND_c_545_n 0.00655577f $X=0.855 $Y=0.445 $X2=0 $Y2=0
cc_115 N_A_N_c_83_n N_VGND_c_545_n 7.69802e-19 $X=0.675 $Y=0.985 $X2=0 $Y2=0
cc_116 N_A_N_c_86_n N_VGND_c_545_n 0.0122691f $X=0.63 $Y=1.02 $X2=0 $Y2=0
cc_117 N_A_27_47#_c_134_n N_A_332_352#_c_206_n 0.0073875f $X=1.255 $Y=1.895
+ $X2=0 $Y2=0
cc_118 N_A_27_47#_c_125_n N_A_332_352#_c_206_n 0.0130448f $X=1.77 $Y=0.805 $X2=0
+ $Y2=0
cc_119 N_A_27_47#_c_128_n N_A_332_352#_c_206_n 0.0219931f $X=1.255 $Y=1.225
+ $X2=0 $Y2=0
cc_120 N_A_27_47#_c_131_n N_A_332_352#_c_206_n 4.92733e-19 $X=1.255 $Y=1.39
+ $X2=0 $Y2=0
cc_121 N_A_27_47#_M1000_g N_A_332_352#_M1009_g 0.0253238f $X=1.255 $Y=2.595
+ $X2=0 $Y2=0
cc_122 N_A_27_47#_c_127_n N_A_332_352#_M1005_g 0.0496183f $X=1.845 $Y=0.73 $X2=0
+ $Y2=0
cc_123 N_A_27_47#_c_128_n N_A_332_352#_M1005_g 0.00187375f $X=1.255 $Y=1.225
+ $X2=0 $Y2=0
cc_124 N_A_27_47#_c_134_n N_VPWR_c_409_n 3.10915e-19 $X=1.255 $Y=1.895 $X2=0
+ $Y2=0
cc_125 N_A_27_47#_M1000_g N_VPWR_c_409_n 0.023424f $X=1.255 $Y=2.595 $X2=0 $Y2=0
cc_126 N_A_27_47#_c_138_n N_VPWR_c_409_n 0.067477f $X=0.46 $Y=2.24 $X2=0 $Y2=0
cc_127 N_A_27_47#_c_139_n N_VPWR_c_409_n 0.0265231f $X=1.09 $Y=1.81 $X2=0 $Y2=0
cc_128 N_A_27_47#_M1000_g N_VPWR_c_410_n 0.0010306f $X=1.255 $Y=2.595 $X2=0
+ $Y2=0
cc_129 N_A_27_47#_c_138_n N_VPWR_c_412_n 0.0318944f $X=0.46 $Y=2.24 $X2=0 $Y2=0
cc_130 N_A_27_47#_M1000_g N_VPWR_c_416_n 0.00840199f $X=1.255 $Y=2.595 $X2=0
+ $Y2=0
cc_131 N_A_27_47#_M1008_s N_VPWR_c_408_n 0.0023218f $X=0.315 $Y=2.095 $X2=0
+ $Y2=0
cc_132 N_A_27_47#_M1000_g N_VPWR_c_408_n 0.0136033f $X=1.255 $Y=2.595 $X2=0
+ $Y2=0
cc_133 N_A_27_47#_c_138_n N_VPWR_c_408_n 0.0194728f $X=0.46 $Y=2.24 $X2=0 $Y2=0
cc_134 N_A_27_47#_M1000_g N_Y_c_473_n 8.72896e-19 $X=1.255 $Y=2.595 $X2=0 $Y2=0
cc_135 N_A_27_47#_c_125_n N_Y_c_473_n 0.0151268f $X=1.77 $Y=0.805 $X2=0 $Y2=0
cc_136 N_A_27_47#_c_127_n N_Y_c_473_n 0.00222717f $X=1.845 $Y=0.73 $X2=0 $Y2=0
cc_137 N_A_27_47#_c_128_n N_Y_c_473_n 0.0113795f $X=1.255 $Y=1.225 $X2=0 $Y2=0
cc_138 N_A_27_47#_c_129_n N_Y_c_473_n 5.29e-19 $X=1.255 $Y=1.73 $X2=0 $Y2=0
cc_139 N_A_27_47#_c_139_n N_Y_c_473_n 0.0129673f $X=1.09 $Y=1.81 $X2=0 $Y2=0
cc_140 N_A_27_47#_c_131_n N_Y_c_473_n 0.0359225f $X=1.255 $Y=1.39 $X2=0 $Y2=0
cc_141 N_A_27_47#_M1000_g N_Y_c_477_n 0.00385494f $X=1.255 $Y=2.595 $X2=0 $Y2=0
cc_142 N_A_27_47#_M1000_g N_Y_c_488_n 0.0144755f $X=1.255 $Y=2.595 $X2=0 $Y2=0
cc_143 N_A_27_47#_c_139_n N_Y_c_488_n 0.0018973f $X=1.09 $Y=1.81 $X2=0 $Y2=0
cc_144 N_A_27_47#_c_125_n N_Y_c_474_n 0.00580169f $X=1.77 $Y=0.805 $X2=0 $Y2=0
cc_145 N_A_27_47#_c_127_n N_Y_c_474_n 0.00830278f $X=1.845 $Y=0.73 $X2=0 $Y2=0
cc_146 N_A_27_47#_c_127_n N_VGND_c_540_n 0.00336443f $X=1.845 $Y=0.73 $X2=0
+ $Y2=0
cc_147 N_A_27_47#_c_131_n N_VGND_c_540_n 0.00523728f $X=1.255 $Y=1.39 $X2=0
+ $Y2=0
cc_148 N_A_27_47#_c_132_n N_VGND_c_540_n 9.23947e-19 $X=1.255 $Y=1.39 $X2=0
+ $Y2=0
cc_149 N_A_27_47#_c_133_n N_VGND_c_540_n 0.0137175f $X=0.28 $Y=0.47 $X2=0 $Y2=0
cc_150 N_A_27_47#_c_133_n N_VGND_c_542_n 0.0195507f $X=0.28 $Y=0.47 $X2=0 $Y2=0
cc_151 N_A_27_47#_c_125_n N_VGND_c_543_n 3.99655e-19 $X=1.77 $Y=0.805 $X2=0
+ $Y2=0
cc_152 N_A_27_47#_c_126_n N_VGND_c_543_n 0.00392688f $X=1.42 $Y=0.805 $X2=0
+ $Y2=0
cc_153 N_A_27_47#_c_127_n N_VGND_c_543_n 0.00549284f $X=1.845 $Y=0.73 $X2=0
+ $Y2=0
cc_154 N_A_27_47#_M1002_s N_VGND_c_545_n 0.00232985f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_155 N_A_27_47#_c_126_n N_VGND_c_545_n 0.00509033f $X=1.42 $Y=0.805 $X2=0
+ $Y2=0
cc_156 N_A_27_47#_c_127_n N_VGND_c_545_n 0.0113234f $X=1.845 $Y=0.73 $X2=0 $Y2=0
cc_157 N_A_27_47#_c_133_n N_VGND_c_545_n 0.0124998f $X=0.28 $Y=0.47 $X2=0 $Y2=0
cc_158 N_A_332_352#_M1009_g N_C_M1004_g 0.0178841f $X=1.785 $Y=2.595 $X2=0 $Y2=0
cc_159 N_A_332_352#_M1005_g N_C_M1006_g 0.0851103f $X=2.205 $Y=0.445 $X2=0 $Y2=0
cc_160 N_A_332_352#_c_208_n N_C_M1006_g 0.0108447f $X=3.825 $Y=1.35 $X2=0 $Y2=0
cc_161 N_A_332_352#_c_211_n N_C_M1006_g 0.00235573f $X=2.115 $Y=1.255 $X2=0
+ $Y2=0
cc_162 N_A_332_352#_c_206_n N_C_c_281_n 0.0139099f $X=1.785 $Y=1.885 $X2=0 $Y2=0
cc_163 N_A_332_352#_c_208_n N_C_c_281_n 0.004479f $X=3.825 $Y=1.35 $X2=0 $Y2=0
cc_164 N_A_332_352#_c_211_n N_C_c_281_n 5.76377e-19 $X=2.115 $Y=1.255 $X2=0
+ $Y2=0
cc_165 N_A_332_352#_c_206_n N_C_c_284_n 0.0014981f $X=1.785 $Y=1.885 $X2=0 $Y2=0
cc_166 N_A_332_352#_M1009_g N_C_c_284_n 4.13831e-19 $X=1.785 $Y=2.595 $X2=0
+ $Y2=0
cc_167 N_A_332_352#_c_208_n N_C_c_284_n 0.0240581f $X=3.825 $Y=1.35 $X2=0 $Y2=0
cc_168 N_A_332_352#_c_211_n N_C_c_284_n 0.00918916f $X=2.115 $Y=1.255 $X2=0
+ $Y2=0
cc_169 N_A_332_352#_c_209_n N_D_M1012_g 0.00110956f $X=3.99 $Y=2.24 $X2=0 $Y2=0
cc_170 N_A_332_352#_c_208_n N_D_c_323_n 5.17254e-19 $X=3.825 $Y=1.35 $X2=0 $Y2=0
cc_171 N_A_332_352#_c_208_n N_D_c_324_n 0.00446396f $X=3.825 $Y=1.35 $X2=0 $Y2=0
cc_172 N_A_332_352#_c_209_n N_D_c_324_n 8.83015e-19 $X=3.99 $Y=2.24 $X2=0 $Y2=0
cc_173 N_A_332_352#_c_208_n N_D_c_325_n 0.0260416f $X=3.825 $Y=1.35 $X2=0 $Y2=0
cc_174 N_A_332_352#_c_209_n N_D_c_325_n 0.0188277f $X=3.99 $Y=2.24 $X2=0 $Y2=0
cc_175 N_A_332_352#_c_208_n N_D_c_326_n 0.0116388f $X=3.825 $Y=1.35 $X2=0 $Y2=0
cc_176 N_A_332_352#_c_209_n N_D_c_326_n 6.5549e-19 $X=3.99 $Y=2.24 $X2=0 $Y2=0
cc_177 N_A_332_352#_c_213_n N_B_N_c_368_n 8.11479e-19 $X=4.04 $Y=0.4 $X2=-0.19
+ $Y2=-0.245
cc_178 N_A_332_352#_c_208_n N_B_N_M1010_g 0.0224193f $X=3.825 $Y=1.35 $X2=0
+ $Y2=0
cc_179 N_A_332_352#_c_209_n N_B_N_M1010_g 0.0479717f $X=3.99 $Y=2.24 $X2=0 $Y2=0
cc_180 N_A_332_352#_c_210_n N_B_N_M1010_g 0.00427033f $X=4.12 $Y=1.265 $X2=0
+ $Y2=0
cc_181 N_A_332_352#_c_212_n N_B_N_M1010_g 0.00525478f $X=4.015 $Y=1.35 $X2=0
+ $Y2=0
cc_182 N_A_332_352#_c_210_n N_B_N_c_370_n 0.0137774f $X=4.12 $Y=1.265 $X2=0
+ $Y2=0
cc_183 N_A_332_352#_c_213_n N_B_N_c_370_n 0.00570002f $X=4.04 $Y=0.4 $X2=0 $Y2=0
cc_184 N_A_332_352#_M1005_g B_N 0.0020169f $X=2.205 $Y=0.445 $X2=0 $Y2=0
cc_185 N_A_332_352#_c_208_n B_N 0.0866224f $X=3.825 $Y=1.35 $X2=0 $Y2=0
cc_186 N_A_332_352#_c_210_n B_N 0.0159676f $X=4.12 $Y=1.265 $X2=0 $Y2=0
cc_187 N_A_332_352#_c_208_n N_B_N_c_372_n 0.00556062f $X=3.825 $Y=1.35 $X2=0
+ $Y2=0
cc_188 N_A_332_352#_c_212_n N_B_N_c_372_n 0.00207933f $X=4.015 $Y=1.35 $X2=0
+ $Y2=0
cc_189 N_A_332_352#_M1009_g N_VPWR_c_409_n 0.0018959f $X=1.785 $Y=2.595 $X2=0
+ $Y2=0
cc_190 N_A_332_352#_M1009_g N_VPWR_c_410_n 0.0127295f $X=1.785 $Y=2.595 $X2=0
+ $Y2=0
cc_191 N_A_332_352#_M1009_g N_VPWR_c_416_n 0.00840199f $X=1.785 $Y=2.595 $X2=0
+ $Y2=0
cc_192 N_A_332_352#_c_209_n N_VPWR_c_417_n 0.0231292f $X=3.99 $Y=2.24 $X2=0
+ $Y2=0
cc_193 N_A_332_352#_M1010_d N_VPWR_c_408_n 0.0023218f $X=3.85 $Y=2.095 $X2=0
+ $Y2=0
cc_194 N_A_332_352#_M1009_g N_VPWR_c_408_n 0.00749742f $X=1.785 $Y=2.595 $X2=0
+ $Y2=0
cc_195 N_A_332_352#_c_209_n N_VPWR_c_408_n 0.0144427f $X=3.99 $Y=2.24 $X2=0
+ $Y2=0
cc_196 N_A_332_352#_c_206_n N_Y_c_473_n 0.0251671f $X=1.785 $Y=1.885 $X2=0 $Y2=0
cc_197 N_A_332_352#_M1009_g N_Y_c_473_n 0.00282228f $X=1.785 $Y=2.595 $X2=0
+ $Y2=0
cc_198 N_A_332_352#_M1005_g N_Y_c_473_n 0.00478243f $X=2.205 $Y=0.445 $X2=0
+ $Y2=0
cc_199 N_A_332_352#_c_211_n N_Y_c_473_n 0.0457028f $X=2.115 $Y=1.255 $X2=0 $Y2=0
cc_200 N_A_332_352#_M1009_g N_Y_c_496_n 0.0157857f $X=1.785 $Y=2.595 $X2=0 $Y2=0
cc_201 N_A_332_352#_c_206_n N_Y_c_476_n 0.00406381f $X=1.785 $Y=1.885 $X2=0
+ $Y2=0
cc_202 N_A_332_352#_M1009_g N_Y_c_476_n 0.0130935f $X=1.785 $Y=2.595 $X2=0 $Y2=0
cc_203 N_A_332_352#_c_211_n N_Y_c_476_n 0.0265158f $X=2.115 $Y=1.255 $X2=0 $Y2=0
cc_204 N_A_332_352#_M1009_g N_Y_c_477_n 0.00407173f $X=1.785 $Y=2.595 $X2=0
+ $Y2=0
cc_205 N_A_332_352#_M1009_g N_Y_c_488_n 0.016659f $X=1.785 $Y=2.595 $X2=0 $Y2=0
cc_206 N_A_332_352#_M1005_g N_Y_c_474_n 0.00205641f $X=2.205 $Y=0.445 $X2=0
+ $Y2=0
cc_207 N_A_332_352#_M1009_g Y 0.00530319f $X=1.785 $Y=2.595 $X2=0 $Y2=0
cc_208 N_A_332_352#_M1005_g N_VGND_c_543_n 0.00585385f $X=2.205 $Y=0.445 $X2=0
+ $Y2=0
cc_209 N_A_332_352#_c_213_n N_VGND_c_544_n 0.0164114f $X=4.04 $Y=0.4 $X2=0 $Y2=0
cc_210 N_A_332_352#_M1001_d N_VGND_c_545_n 0.00234032f $X=3.9 $Y=0.235 $X2=0
+ $Y2=0
cc_211 N_A_332_352#_M1005_g N_VGND_c_545_n 0.0107317f $X=2.205 $Y=0.445 $X2=0
+ $Y2=0
cc_212 N_A_332_352#_c_213_n N_VGND_c_545_n 0.012174f $X=4.04 $Y=0.4 $X2=0 $Y2=0
cc_213 N_C_M1006_g N_D_c_322_n 0.0433949f $X=2.595 $Y=0.445 $X2=-0.19 $Y2=-0.245
cc_214 N_C_M1004_g N_D_M1012_g 0.0252409f $X=2.625 $Y=2.595 $X2=0 $Y2=0
cc_215 N_C_c_284_n N_D_M1012_g 7.25438e-19 $X=2.655 $Y=1.77 $X2=0 $Y2=0
cc_216 N_C_c_281_n N_D_c_324_n 0.0207936f $X=2.655 $Y=1.77 $X2=0 $Y2=0
cc_217 N_C_c_284_n N_D_c_324_n 3.82746e-19 $X=2.655 $Y=1.77 $X2=0 $Y2=0
cc_218 N_C_M1004_g N_D_c_325_n 5.28738e-19 $X=2.625 $Y=2.595 $X2=0 $Y2=0
cc_219 N_C_c_281_n N_D_c_325_n 0.00182931f $X=2.655 $Y=1.77 $X2=0 $Y2=0
cc_220 N_C_c_284_n N_D_c_325_n 0.0385571f $X=2.655 $Y=1.77 $X2=0 $Y2=0
cc_221 N_C_M1006_g N_D_c_326_n 0.0262255f $X=2.595 $Y=0.445 $X2=0 $Y2=0
cc_222 N_C_M1006_g B_N 0.0185416f $X=2.595 $Y=0.445 $X2=0 $Y2=0
cc_223 N_C_M1004_g N_VPWR_c_410_n 0.0067938f $X=2.625 $Y=2.595 $X2=0 $Y2=0
cc_224 N_C_M1004_g N_VPWR_c_411_n 0.00112815f $X=2.625 $Y=2.595 $X2=0 $Y2=0
cc_225 N_C_M1004_g N_VPWR_c_414_n 0.00939541f $X=2.625 $Y=2.595 $X2=0 $Y2=0
cc_226 N_C_M1004_g N_VPWR_c_408_n 0.0100563f $X=2.625 $Y=2.595 $X2=0 $Y2=0
cc_227 N_C_c_284_n N_Y_M1004_d 6.27237e-19 $X=2.655 $Y=1.77 $X2=0 $Y2=0
cc_228 N_C_M1004_g N_Y_c_476_n 8.20519e-19 $X=2.625 $Y=2.595 $X2=0 $Y2=0
cc_229 N_C_c_284_n N_Y_c_476_n 0.0121411f $X=2.655 $Y=1.77 $X2=0 $Y2=0
cc_230 N_C_M1004_g N_Y_c_507_n 0.0160838f $X=2.625 $Y=2.595 $X2=0 $Y2=0
cc_231 N_C_c_284_n N_Y_c_507_n 0.0161359f $X=2.655 $Y=1.77 $X2=0 $Y2=0
cc_232 N_C_M1004_g N_Y_c_509_n 0.0168898f $X=2.625 $Y=2.595 $X2=0 $Y2=0
cc_233 N_C_c_281_n N_Y_c_509_n 2.16536e-19 $X=2.655 $Y=1.77 $X2=0 $Y2=0
cc_234 N_C_c_284_n N_Y_c_509_n 0.00296201f $X=2.655 $Y=1.77 $X2=0 $Y2=0
cc_235 N_C_M1004_g Y 0.00444502f $X=2.625 $Y=2.595 $X2=0 $Y2=0
cc_236 N_C_M1006_g N_VGND_c_541_n 0.00282271f $X=2.595 $Y=0.445 $X2=0 $Y2=0
cc_237 N_C_M1006_g N_VGND_c_543_n 0.00585385f $X=2.595 $Y=0.445 $X2=0 $Y2=0
cc_238 N_C_M1006_g N_VGND_c_545_n 0.00633809f $X=2.595 $Y=0.445 $X2=0 $Y2=0
cc_239 N_D_c_322_n N_B_N_c_368_n 0.010977f $X=2.985 $Y=0.73 $X2=-0.19 $Y2=-0.245
cc_240 N_D_c_323_n N_B_N_c_368_n 0.0119223f $X=3.105 $Y=0.805 $X2=-0.19
+ $Y2=-0.245
cc_241 N_D_M1012_g N_B_N_M1010_g 0.021829f $X=3.155 $Y=2.595 $X2=0 $Y2=0
cc_242 N_D_c_324_n N_B_N_M1010_g 0.0176275f $X=3.195 $Y=1.77 $X2=0 $Y2=0
cc_243 N_D_c_325_n N_B_N_M1010_g 0.00326508f $X=3.195 $Y=1.77 $X2=0 $Y2=0
cc_244 N_D_c_326_n N_B_N_M1010_g 0.0160605f $X=3.195 $Y=1.605 $X2=0 $Y2=0
cc_245 N_D_c_323_n B_N 0.0113412f $X=3.105 $Y=0.805 $X2=0 $Y2=0
cc_246 N_D_c_326_n B_N 0.00974474f $X=3.195 $Y=1.605 $X2=0 $Y2=0
cc_247 N_D_c_326_n N_B_N_c_372_n 0.0119223f $X=3.195 $Y=1.605 $X2=0 $Y2=0
cc_248 N_D_c_325_n N_VPWR_M1012_d 9.87716e-19 $X=3.195 $Y=1.77 $X2=0 $Y2=0
cc_249 N_D_M1012_g N_VPWR_c_411_n 0.0189192f $X=3.155 $Y=2.595 $X2=0 $Y2=0
cc_250 N_D_c_324_n N_VPWR_c_411_n 2.65185e-19 $X=3.195 $Y=1.77 $X2=0 $Y2=0
cc_251 N_D_c_325_n N_VPWR_c_411_n 0.00373121f $X=3.195 $Y=1.77 $X2=0 $Y2=0
cc_252 N_D_M1012_g N_VPWR_c_414_n 0.00840199f $X=3.155 $Y=2.595 $X2=0 $Y2=0
cc_253 N_D_M1012_g N_VPWR_c_408_n 0.0136033f $X=3.155 $Y=2.595 $X2=0 $Y2=0
cc_254 N_D_M1012_g N_Y_c_509_n 0.0132063f $X=3.155 $Y=2.595 $X2=0 $Y2=0
cc_255 N_D_c_325_n N_Y_c_509_n 0.00194374f $X=3.195 $Y=1.77 $X2=0 $Y2=0
cc_256 N_D_c_322_n N_VGND_c_541_n 0.0113084f $X=2.985 $Y=0.73 $X2=0 $Y2=0
cc_257 N_D_c_323_n N_VGND_c_541_n 0.00319214f $X=3.105 $Y=0.805 $X2=0 $Y2=0
cc_258 N_D_c_322_n N_VGND_c_543_n 0.00486043f $X=2.985 $Y=0.73 $X2=0 $Y2=0
cc_259 N_D_c_322_n N_VGND_c_545_n 0.00438061f $X=2.985 $Y=0.73 $X2=0 $Y2=0
cc_260 N_B_N_M1010_g N_VPWR_c_411_n 0.00362166f $X=3.725 $Y=2.595 $X2=0 $Y2=0
cc_261 N_B_N_M1010_g N_VPWR_c_417_n 0.00939541f $X=3.725 $Y=2.595 $X2=0 $Y2=0
cc_262 N_B_N_M1010_g N_VPWR_c_408_n 0.0169788f $X=3.725 $Y=2.595 $X2=0 $Y2=0
cc_263 N_B_N_c_368_n N_VGND_c_541_n 0.00316183f $X=3.465 $Y=0.765 $X2=0 $Y2=0
cc_264 B_N N_VGND_c_541_n 0.0217614f $X=3.515 $Y=0.84 $X2=0 $Y2=0
cc_265 N_B_N_c_368_n N_VGND_c_544_n 0.00585385f $X=3.465 $Y=0.765 $X2=0 $Y2=0
cc_266 N_B_N_c_370_n N_VGND_c_544_n 0.00550269f $X=3.825 $Y=0.765 $X2=0 $Y2=0
cc_267 N_B_N_c_372_n N_VGND_c_544_n 5.95547e-19 $X=3.825 $Y=0.93 $X2=0 $Y2=0
cc_268 N_B_N_c_368_n N_VGND_c_545_n 0.00599793f $X=3.465 $Y=0.765 $X2=0 $Y2=0
cc_269 N_B_N_c_370_n N_VGND_c_545_n 0.0107628f $X=3.825 $Y=0.765 $X2=0 $Y2=0
cc_270 B_N N_VGND_c_545_n 0.0312296f $X=3.515 $Y=0.84 $X2=0 $Y2=0
cc_271 N_B_N_c_372_n N_VGND_c_545_n 8.01698e-19 $X=3.825 $Y=0.93 $X2=0 $Y2=0
cc_272 N_VPWR_c_408_n N_Y_M1000_d 0.00223819f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_273 N_VPWR_c_408_n N_Y_M1004_d 0.00223819f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_274 N_VPWR_M1009_d N_Y_c_496_n 0.0015061f $X=1.91 $Y=2.095 $X2=0 $Y2=0
cc_275 N_VPWR_c_410_n N_Y_c_496_n 0.00765546f $X=2.05 $Y=2.905 $X2=0 $Y2=0
cc_276 N_VPWR_c_408_n N_Y_c_496_n 0.00627166f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_277 N_VPWR_M1009_d N_Y_c_476_n 0.00105305f $X=1.91 $Y=2.095 $X2=0 $Y2=0
cc_278 N_VPWR_c_409_n N_Y_c_477_n 0.00140894f $X=0.99 $Y=2.24 $X2=0 $Y2=0
cc_279 N_VPWR_M1009_d N_Y_c_507_n 0.0102318f $X=1.91 $Y=2.095 $X2=0 $Y2=0
cc_280 N_VPWR_c_408_n N_Y_c_507_n 0.0144615f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_281 N_VPWR_c_409_n N_Y_c_488_n 0.0518318f $X=0.99 $Y=2.24 $X2=0 $Y2=0
cc_282 N_VPWR_c_410_n N_Y_c_488_n 0.0240501f $X=2.05 $Y=2.905 $X2=0 $Y2=0
cc_283 N_VPWR_c_416_n N_Y_c_488_n 0.0177952f $X=1.885 $Y=3.33 $X2=0 $Y2=0
cc_284 N_VPWR_c_408_n N_Y_c_488_n 0.0123247f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_285 N_VPWR_c_410_n N_Y_c_509_n 0.0120571f $X=2.05 $Y=2.905 $X2=0 $Y2=0
cc_286 N_VPWR_c_411_n N_Y_c_509_n 0.0491843f $X=3.42 $Y=2.495 $X2=0 $Y2=0
cc_287 N_VPWR_c_414_n N_Y_c_509_n 0.0177952f $X=3.255 $Y=3.33 $X2=0 $Y2=0
cc_288 N_VPWR_c_408_n N_Y_c_509_n 0.0123247f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_289 N_VPWR_M1009_d Y 0.0125321f $X=1.91 $Y=2.095 $X2=0 $Y2=0
cc_290 N_VPWR_c_410_n Y 0.0140272f $X=2.05 $Y=2.905 $X2=0 $Y2=0
cc_291 N_VPWR_c_408_n Y 0.0030818f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_292 N_Y_c_474_n N_VGND_c_540_n 0.0276416f $X=1.63 $Y=0.47 $X2=0 $Y2=0
cc_293 N_Y_c_474_n N_VGND_c_543_n 0.0194164f $X=1.63 $Y=0.47 $X2=0 $Y2=0
cc_294 N_Y_M1003_s N_VGND_c_545_n 0.00232985f $X=1.485 $Y=0.235 $X2=0 $Y2=0
cc_295 N_Y_c_474_n N_VGND_c_545_n 0.0125003f $X=1.63 $Y=0.47 $X2=0 $Y2=0
cc_296 A_114_47# N_VGND_c_545_n 0.00312559f $X=0.57 $Y=0.235 $X2=4.08 $Y2=0
cc_297 N_VGND_c_545_n A_384_47# 0.00899413f $X=4.08 $Y=0 $X2=-0.19 $Y2=-0.245
cc_298 N_VGND_c_545_n A_456_47# 0.010279f $X=4.08 $Y=0 $X2=-0.19 $Y2=-0.245
cc_299 N_VGND_c_545_n A_534_47# 0.00325212f $X=4.08 $Y=0 $X2=-0.19 $Y2=-0.245
cc_300 N_VGND_c_545_n A_708_47# 0.00372397f $X=4.08 $Y=0 $X2=-0.19 $Y2=-0.245
