* File: sky130_fd_sc_lp__o41a_0.spice
* Created: Fri Aug 28 11:19:00 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__o41a_0.pex.spice"
.subckt sky130_fd_sc_lp__o41a_0  VNB VPB B1 A4 A3 A2 A1 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* A1	A1
* A2	A2
* A3	A3
* A4	A4
* B1	B1
* VPB	VPB
* VNB	VNB
MM1003 N_VGND_M1003_d N_A_80_21#_M1003_g N_X_M1003_s VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.1113 PD=1.37 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1007 N_A_319_51#_M1007_d N_B1_M1007_g N_A_80_21#_M1007_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002 A=0.063 P=1.14 MULT=1
MM1009 N_VGND_M1009_d N_A4_M1009_g N_A_319_51#_M1007_d VNB NSHORT L=0.15 W=0.42
+ AD=0.063 AS=0.0588 PD=0.72 PS=0.7 NRD=4.284 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75001.5 A=0.063 P=1.14 MULT=1
MM1000 N_A_319_51#_M1000_d N_A3_M1000_g N_VGND_M1009_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.063 PD=0.7 PS=0.72 NRD=0 NRS=1.428 M=1 R=2.8 SA=75001.1
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1004 N_VGND_M1004_d N_A2_M1004_g N_A_319_51#_M1000_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0672 AS=0.0588 PD=0.74 PS=0.7 NRD=5.712 NRS=0 M=1 R=2.8 SA=75001.5
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1002 N_A_319_51#_M1002_d N_A1_M1002_g N_VGND_M1004_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.0672 PD=1.37 PS=0.74 NRD=0 NRS=5.712 M=1 R=2.8 SA=75002
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1010 N_VPWR_M1010_d N_A_80_21#_M1010_g N_X_M1010_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0896 AS=0.1696 PD=0.92 PS=1.81 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75002.8 A=0.096 P=1.58 MULT=1
MM1005 N_A_80_21#_M1005_d N_B1_M1005_g N_VPWR_M1010_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.256 AS=0.0896 PD=1.44 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.6
+ SB=75002.4 A=0.096 P=1.58 MULT=1
MM1006 A_423_483# N_A4_M1006_g N_A_80_21#_M1005_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.096 AS=0.256 PD=0.94 PS=1.44 NRD=29.2348 NRS=0 M=1 R=4.26667 SA=75001.6
+ SB=75001.4 A=0.096 P=1.58 MULT=1
MM1008 A_513_483# N_A3_M1008_g A_423_483# VPB PHIGHVT L=0.15 W=0.64 AD=0.096
+ AS=0.096 PD=0.94 PS=0.94 NRD=29.2348 NRS=29.2348 M=1 R=4.26667 SA=75002
+ SB=75001 A=0.096 P=1.58 MULT=1
MM1011 A_603_483# N_A2_M1011_g A_513_483# VPB PHIGHVT L=0.15 W=0.64 AD=0.0672
+ AS=0.096 PD=0.85 PS=0.94 NRD=15.3857 NRS=29.2348 M=1 R=4.26667 SA=75002.5
+ SB=75000.6 A=0.096 P=1.58 MULT=1
MM1001 N_VPWR_M1001_d N_A1_M1001_g A_603_483# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1696 AS=0.0672 PD=1.81 PS=0.85 NRD=0 NRS=15.3857 M=1 R=4.26667 SA=75002.8
+ SB=75000.2 A=0.096 P=1.58 MULT=1
DX12_noxref VNB VPB NWDIODE A=7.8703 P=12.17
*
.include "sky130_fd_sc_lp__o41a_0.pxi.spice"
*
.ends
*
*
