# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__dlxtn_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_lp__dlxtn_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.200000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.490000 1.200000 1.855000 1.490000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.588000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.370000 0.300000 6.635000 3.075000 ;
    END
  END Q
  PIN GATE_N
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 1.015000 0.275000 2.290000 0.640000 ;
    END
  END GATE_N
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 7.200000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 7.200000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.200000 0.085000 ;
      RECT 0.000000  3.245000 7.200000 3.415000 ;
      RECT 0.140000  0.695000 0.495000 1.025000 ;
      RECT 0.140000  1.025000 0.310000 1.660000 ;
      RECT 0.140000  1.660000 2.925000 1.855000 ;
      RECT 0.140000  1.855000 0.625000 3.055000 ;
      RECT 0.675000  0.085000 0.845000 0.810000 ;
      RECT 0.675000  0.810000 1.005000 1.025000 ;
      RECT 0.795000  2.415000 1.045000 3.245000 ;
      RECT 1.185000  0.810000 2.290000 0.995000 ;
      RECT 1.185000  0.995000 3.925000 1.030000 ;
      RECT 1.215000  2.395000 1.515000 2.905000 ;
      RECT 1.215000  2.905000 2.305000 3.075000 ;
      RECT 1.705000  2.035000 3.495000 2.205000 ;
      RECT 1.705000  2.205000 1.955000 2.735000 ;
      RECT 2.025000  1.030000 3.925000 1.165000 ;
      RECT 2.025000  1.165000 2.340000 1.490000 ;
      RECT 2.135000  2.375000 3.965000 2.545000 ;
      RECT 2.135000  2.545000 2.305000 2.905000 ;
      RECT 2.460000  0.275000 2.720000 0.645000 ;
      RECT 2.460000  0.645000 4.425000 0.815000 ;
      RECT 2.475000  2.715000 2.735000 3.245000 ;
      RECT 2.595000  1.345000 2.925000 1.660000 ;
      RECT 2.890000  0.085000 3.220000 0.475000 ;
      RECT 3.165000  1.535000 3.495000 2.035000 ;
      RECT 3.290000  2.715000 4.305000 3.065000 ;
      RECT 3.705000  1.165000 3.925000 1.915000 ;
      RECT 3.705000  1.915000 3.965000 2.375000 ;
      RECT 3.790000  0.255000 4.775000 0.475000 ;
      RECT 4.095000  0.815000 4.425000 1.100000 ;
      RECT 4.135000  1.270000 5.355000 1.450000 ;
      RECT 4.135000  1.450000 4.305000 2.715000 ;
      RECT 4.475000  2.495000 5.245000 3.245000 ;
      RECT 4.485000  1.620000 5.705000 1.790000 ;
      RECT 4.485000  1.790000 4.815000 2.245000 ;
      RECT 4.605000  0.475000 4.775000 1.260000 ;
      RECT 4.605000  1.260000 5.355000 1.270000 ;
      RECT 4.945000  0.085000 5.170000 1.090000 ;
      RECT 5.015000  1.960000 5.245000 2.495000 ;
      RECT 5.340000  0.255000 5.705000 1.090000 ;
      RECT 5.415000  1.790000 5.705000 2.960000 ;
      RECT 5.535000  1.090000 5.705000 1.270000 ;
      RECT 5.535000  1.270000 6.165000 1.600000 ;
      RECT 5.535000  1.600000 5.705000 1.620000 ;
      RECT 5.905000  0.085000 6.200000 1.100000 ;
      RECT 5.905000  1.815000 6.200000 3.245000 ;
      RECT 6.805000  0.085000 7.095000 1.180000 ;
      RECT 6.805000  1.815000 7.095000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
  END
END sky130_fd_sc_lp__dlxtn_2
END LIBRARY
