* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__nand3b_lp A_N B C VGND VNB VPB VPWR Y
X0 Y a_90_247# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X1 Y a_90_247# a_156_141# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 a_234_141# C VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 a_420_141# A_N a_90_247# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X5 a_156_141# B a_234_141# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 VGND A_N a_420_141# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X8 VPWR A_N a_90_247# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
.ends
