* File: sky130_fd_sc_lp__sdfrbp_lp.pex.spice
* Created: Wed Sep  2 10:34:20 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__SDFRBP_LP%SCE 3 7 11 15 17 19 21 24 28 30 33 34 35
+ 36 41
r72 41 42 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.64
+ $Y=1.48 $X2=0.64 $Y2=1.48
r73 35 36 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.64 $Y=1.665
+ $X2=0.64 $Y2=2.035
r74 35 42 6.46067 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=0.64 $Y=1.665
+ $X2=0.64 $Y2=1.48
r75 34 42 6.46067 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=0.64 $Y=1.295
+ $X2=0.64 $Y2=1.48
r76 31 41 38.3708 $w=4.95e-07 $l=3.55e-07 $layer=POLY_cond $X=0.722 $Y=1.835
+ $X2=0.722 $Y2=1.48
r77 30 31 7.86808 $w=5.1e-07 $l=7.5e-08 $layer=POLY_cond $X=0.73 $Y=1.91
+ $X2=0.73 $Y2=1.835
r78 28 41 1.6213 $w=4.95e-07 $l=1.5e-08 $layer=POLY_cond $X=0.722 $Y=1.465
+ $X2=0.722 $Y2=1.48
r79 22 33 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.635 $Y=1.985
+ $X2=1.635 $Y2=1.91
r80 22 24 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.635 $Y=1.985
+ $X2=1.635 $Y2=2.775
r81 19 33 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.635 $Y=1.835
+ $X2=1.635 $Y2=1.91
r82 19 21 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.635 $Y=1.835
+ $X2=1.635 $Y2=1.515
r83 18 30 31.9091 $w=1.5e-07 $l=2.55e-07 $layer=POLY_cond $X=0.985 $Y=1.91
+ $X2=0.73 $Y2=1.91
r84 17 33 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.56 $Y=1.91
+ $X2=1.635 $Y2=1.91
r85 17 18 294.84 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.56 $Y=1.91
+ $X2=0.985 $Y2=1.91
r86 5 30 37.3844 $w=5.1e-07 $l=7.5e-08 $layer=POLY_cond $X=0.73 $Y=1.985
+ $X2=0.73 $Y2=1.91
r87 5 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=0.91 $Y=1.985
+ $X2=0.91 $Y2=2.775
r88 5 7 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=0.55 $Y=1.985 $X2=0.55
+ $Y2=2.775
r89 1 28 24.455 $w=4.95e-07 $l=1.5e-07 $layer=POLY_cond $X=0.7 $Y=1.315 $X2=0.7
+ $Y2=1.465
r90 1 11 446.106 $w=1.5e-07 $l=8.7e-07 $layer=POLY_cond $X=0.895 $Y=1.315
+ $X2=0.895 $Y2=0.445
r91 1 3 446.106 $w=1.5e-07 $l=8.7e-07 $layer=POLY_cond $X=0.505 $Y=1.315
+ $X2=0.505 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRBP_LP%D 3 8 10 11 15 17 18 22
r49 18 22 10.2718 $w=2.28e-07 $l=2.05e-07 $layer=LI1_cond $X=3.12 $Y=0.555
+ $X2=3.12 $Y2=0.35
r50 15 21 18.3619 $w=3.15e-07 $l=1.2e-07 $layer=POLY_cond $X=1.945 $Y=0.4
+ $X2=2.065 $Y2=0.4
r51 14 17 8.61591 $w=2.68e-07 $l=1.65e-07 $layer=LI1_cond $X=1.945 $Y=0.4
+ $X2=2.11 $Y2=0.4
r52 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.945
+ $Y=0.4 $X2=1.945 $Y2=0.4
r53 11 22 2.50919 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=3.005 $Y=0.35
+ $X2=3.12 $Y2=0.35
r54 11 17 58.3904 $w=1.68e-07 $l=8.95e-07 $layer=LI1_cond $X=3.005 $Y=0.35
+ $X2=2.11 $Y2=0.35
r55 9 10 53.9552 $w=1.9e-07 $l=1.5e-07 $layer=POLY_cond $X=2.045 $Y=1.835
+ $X2=2.045 $Y2=1.985
r56 8 9 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.065 $Y=1.515
+ $X2=2.065 $Y2=1.835
r57 5 21 20.1192 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.065 $Y=0.565
+ $X2=2.065 $Y2=0.4
r58 5 8 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=2.065 $Y=0.565
+ $X2=2.065 $Y2=1.515
r59 3 10 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.025 $Y=2.775
+ $X2=2.025 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRBP_LP%A_29_47# 1 2 10 13 16 19 23 28 29 31 32 33
r71 32 37 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.515 $Y=0.75
+ $X2=2.515 $Y2=0.915
r72 31 33 10.9635 $w=2.68e-07 $l=2.2e-07 $layer=LI1_cond $X=2.515 $Y=0.75
+ $X2=2.295 $Y2=0.75
r73 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.515
+ $Y=0.75 $X2=2.515 $Y2=0.75
r74 27 28 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.455 $Y=0.8
+ $X2=0.29 $Y2=0.8
r75 27 33 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=0.455 $Y=0.8
+ $X2=2.295 $Y2=0.8
r76 23 29 9.23056 $w=3.73e-07 $l=1.87e-07 $layer=LI1_cond $X=0.312 $Y=2.622
+ $X2=0.312 $Y2=2.435
r77 23 25 4.16427 $w=3.75e-07 $l=1.28e-07 $layer=LI1_cond $X=0.312 $Y=2.622
+ $X2=0.312 $Y2=2.75
r78 21 28 3.70735 $w=2.5e-07 $l=1.18427e-07 $layer=LI1_cond $X=0.21 $Y=0.885
+ $X2=0.29 $Y2=0.8
r79 21 29 101.123 $w=1.68e-07 $l=1.55e-06 $layer=LI1_cond $X=0.21 $Y=0.885
+ $X2=0.21 $Y2=2.435
r80 17 28 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.29 $Y=0.715
+ $X2=0.29 $Y2=0.8
r81 17 19 8.55602 $w=3.28e-07 $l=2.45e-07 $layer=LI1_cond $X=0.29 $Y=0.715
+ $X2=0.29 $Y2=0.47
r82 15 16 58.3064 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=2.44 $Y=1.835
+ $X2=2.44 $Y2=1.985
r83 13 16 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.455 $Y=2.775
+ $X2=2.455 $Y2=1.985
r84 10 15 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.425 $Y=1.515
+ $X2=2.425 $Y2=1.835
r85 10 37 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=2.425 $Y=1.515
+ $X2=2.425 $Y2=0.915
r86 2 25 600 $w=1.7e-07 $l=3.60278e-07 $layer=licon1_PDIFF $count=1 $X=0.19
+ $Y=2.455 $X2=0.335 $Y2=2.75
r87 1 19 182 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_NDIFF $count=1 $X=0.145
+ $Y=0.235 $X2=0.29 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRBP_LP%SCD 3 5 7 8 10 11 14
c40 10 0 4.85838e-20 $X=2.85 $Y=1.91
r41 14 17 19.2347 $w=3.3e-07 $l=1.1e-07 $layer=POLY_cond $X=3.49 $Y=1.8 $X2=3.49
+ $Y2=1.91
r42 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.49
+ $Y=1.8 $X2=3.49 $Y2=1.8
r43 11 15 4.44514 $w=3.48e-07 $l=1.35e-07 $layer=LI1_cond $X=3.51 $Y=1.665
+ $X2=3.51 $Y2=1.8
r44 9 10 5.30422 $w=1.5e-07 $l=8e-08 $layer=POLY_cond $X=2.93 $Y=1.91 $X2=2.85
+ $Y2=1.91
r45 8 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.325 $Y=1.91
+ $X2=3.49 $Y2=1.91
r46 8 9 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=3.325 $Y=1.91
+ $X2=2.93 $Y2=1.91
r47 5 10 20.4101 $w=1.5e-07 $l=7.74597e-08 $layer=POLY_cond $X=2.855 $Y=1.835
+ $X2=2.85 $Y2=1.91
r48 5 7 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.855 $Y=1.835
+ $X2=2.855 $Y2=1.515
r49 1 10 20.4101 $w=1.5e-07 $l=7.74597e-08 $layer=POLY_cond $X=2.845 $Y=1.985
+ $X2=2.85 $Y2=1.91
r50 1 3 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.845 $Y=1.985
+ $X2=2.845 $Y2=2.775
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRBP_LP%A_876_93# 1 2 9 11 15 19 21 24 25 26 28 29
+ 30 32 33 34 37 40 43 47 50 54 56 57 62
c178 54 0 1.14697e-20 $X=4.545 $Y=0.63
c179 33 0 1.98701e-19 $X=9.765 $Y=0.73
c180 24 0 1.97601e-20 $X=6.655 $Y=0.715
r181 54 60 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.545 $Y=0.63
+ $X2=4.545 $Y2=0.795
r182 53 54 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.545
+ $Y=0.63 $X2=4.545 $Y2=0.63
r183 50 53 9.7783 $w=3.28e-07 $l=2.8e-07 $layer=LI1_cond $X=4.545 $Y=0.35
+ $X2=4.545 $Y2=0.63
r184 48 62 5.51908 $w=2.62e-07 $l=3e-08 $layer=POLY_cond $X=10.735 $Y=1.59
+ $X2=10.765 $Y2=1.59
r185 47 48 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.735
+ $Y=1.6 $X2=10.735 $Y2=1.6
r186 45 57 0.364692 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=10.095 $Y=1.6
+ $X2=9.93 $Y2=1.6
r187 45 47 22.3504 $w=3.28e-07 $l=6.4e-07 $layer=LI1_cond $X=10.095 $Y=1.6
+ $X2=10.735 $Y2=1.6
r188 41 57 6.46576 $w=2.5e-07 $l=2.0106e-07 $layer=LI1_cond $X=9.85 $Y=1.765
+ $X2=9.93 $Y2=1.6
r189 41 43 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=9.85 $Y=1.765
+ $X2=9.85 $Y2=1.98
r190 40 57 6.46576 $w=2.5e-07 $l=1.65e-07 $layer=LI1_cond $X=9.93 $Y=1.435
+ $X2=9.93 $Y2=1.6
r191 39 56 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.93 $Y=0.815
+ $X2=9.93 $Y2=0.73
r192 39 40 21.652 $w=3.28e-07 $l=6.2e-07 $layer=LI1_cond $X=9.93 $Y=0.815
+ $X2=9.93 $Y2=1.435
r193 35 56 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.93 $Y=0.645
+ $X2=9.93 $Y2=0.73
r194 35 37 7.50834 $w=3.28e-07 $l=2.15e-07 $layer=LI1_cond $X=9.93 $Y=0.645
+ $X2=9.93 $Y2=0.43
r195 33 56 3.80956 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.765 $Y=0.73
+ $X2=9.93 $Y2=0.73
r196 33 34 76.6578 $w=1.68e-07 $l=1.175e-06 $layer=LI1_cond $X=9.765 $Y=0.73
+ $X2=8.59 $Y2=0.73
r197 32 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.505 $Y=0.645
+ $X2=8.59 $Y2=0.73
r198 31 32 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=8.505 $Y=0.435
+ $X2=8.505 $Y2=0.645
r199 29 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.42 $Y=0.35
+ $X2=8.505 $Y2=0.435
r200 29 30 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=8.42 $Y=0.35
+ $X2=7.67 $Y2=0.35
r201 27 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.585 $Y=0.435
+ $X2=7.67 $Y2=0.35
r202 27 28 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=7.585 $Y=0.435
+ $X2=7.585 $Y2=0.715
r203 25 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.5 $Y=0.8
+ $X2=7.585 $Y2=0.715
r204 25 26 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=7.5 $Y=0.8 $X2=6.74
+ $Y2=0.8
r205 24 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.655 $Y=0.715
+ $X2=6.74 $Y2=0.8
r206 23 24 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=6.655 $Y=0.435
+ $X2=6.655 $Y2=0.715
r207 22 50 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.71 $Y=0.35
+ $X2=4.545 $Y2=0.35
r208 21 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.57 $Y=0.35
+ $X2=6.655 $Y2=0.435
r209 21 22 121.348 $w=1.68e-07 $l=1.86e-06 $layer=LI1_cond $X=6.57 $Y=0.35
+ $X2=4.71 $Y2=0.35
r210 17 62 57.9504 $w=2.62e-07 $l=3.92874e-07 $layer=POLY_cond $X=11.08 $Y=1.415
+ $X2=10.765 $Y2=1.59
r211 17 19 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=11.08 $Y=1.415
+ $X2=11.08 $Y2=0.915
r212 13 62 15.8058 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=10.765 $Y=1.765
+ $X2=10.765 $Y2=1.59
r213 13 15 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=10.765 $Y=1.765
+ $X2=10.765 $Y2=2.405
r214 9 11 697.362 $w=1.5e-07 $l=1.36e-06 $layer=POLY_cond $X=4.48 $Y=1.305
+ $X2=4.48 $Y2=2.665
r215 9 60 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=4.48 $Y=1.305
+ $X2=4.48 $Y2=0.795
r216 2 43 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=9.71
+ $Y=1.835 $X2=9.85 $Y2=1.98
r217 1 37 91 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_NDIFF $count=2 $X=9.79
+ $Y=0.235 $X2=9.93 $Y2=0.43
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRBP_LP%A_967_193# 1 2 9 13 15 16 19 23 27 31 33
+ 34 36 38 39 40 41 42 45 49 51 53 56 61 62 64 65 68 69 70 72 73 75 82 86 90 92
+ 96 100 101 103 107 109 125
c302 107 0 3.05635e-19 $X=14.85 $Y=1.405
c303 92 0 1.29593e-19 $X=12.855 $Y=0.35
c304 73 0 1.20402e-19 $X=8.59 $Y=1.51
c305 65 0 6.21055e-20 $X=7.64 $Y=1.97
c306 45 0 2.88191e-20 $X=11.31 $Y=2.355
c307 34 0 2.77482e-19 $X=9.79 $Y=1.42
c308 13 0 1.28847e-19 $X=5.025 $Y=2.665
r309 123 125 330.734 $w=1.5e-07 $l=6.45e-07 $layer=POLY_cond $X=14.76 $Y=0.595
+ $X2=14.76 $Y2=1.24
r310 119 120 47.738 $w=3.13e-07 $l=3.1e-07 $layer=POLY_cond $X=9.325 $Y=1.51
+ $X2=9.635 $Y2=1.51
r311 118 119 7.69968 $w=3.13e-07 $l=5e-08 $layer=POLY_cond $X=9.275 $Y=1.51
+ $X2=9.325 $Y2=1.51
r312 107 125 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=14.85 $Y=1.405
+ $X2=14.85 $Y2=1.24
r313 106 109 8.20679 $w=3.28e-07 $l=2.35e-07 $layer=LI1_cond $X=14.85 $Y=1.405
+ $X2=15.085 $Y2=1.405
r314 106 107 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=14.85
+ $Y=1.405 $X2=14.85 $Y2=1.405
r315 100 123 46.255 $w=3.35e-07 $l=1.65e-07 $layer=POLY_cond $X=14.667 $Y=0.43
+ $X2=14.667 $Y2=0.595
r316 99 103 10.877 $w=4.43e-07 $l=4.2e-07 $layer=LI1_cond $X=14.665 $Y=0.487
+ $X2=15.085 $Y2=0.487
r317 99 101 8.86124 $w=4.43e-07 $l=1.65e-07 $layer=LI1_cond $X=14.665 $Y=0.487
+ $X2=14.5 $Y2=0.487
r318 99 100 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=14.665
+ $Y=0.43 $X2=14.665 $Y2=0.43
r319 95 96 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=12.855
+ $Y=0.43 $X2=12.855 $Y2=0.43
r320 92 95 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=12.855 $Y=0.35
+ $X2=12.855 $Y2=0.43
r321 90 115 16.0872 $w=3.3e-07 $l=9.2e-08 $layer=POLY_cond $X=5.99 $Y=2.05
+ $X2=5.99 $Y2=2.142
r322 89 90 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.99
+ $Y=2.05 $X2=5.99 $Y2=2.05
r323 86 89 3.07318 $w=2.98e-07 $l=8e-08 $layer=LI1_cond $X=6.005 $Y=1.97
+ $X2=6.005 $Y2=2.05
r324 82 84 33.8748 $w=3.28e-07 $l=9.7e-07 $layer=LI1_cond $X=15.085 $Y=1.93
+ $X2=15.085 $Y2=2.9
r325 80 109 0.716491 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=15.085 $Y=1.57
+ $X2=15.085 $Y2=1.405
r326 80 82 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=15.085 $Y=1.57
+ $X2=15.085 $Y2=1.93
r327 79 92 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.02 $Y=0.35
+ $X2=12.855 $Y2=0.35
r328 79 101 96.5562 $w=1.68e-07 $l=1.48e-06 $layer=LI1_cond $X=13.02 $Y=0.35
+ $X2=14.5 $Y2=0.35
r329 76 118 26.9489 $w=3.13e-07 $l=1.75e-07 $layer=POLY_cond $X=9.1 $Y=1.51
+ $X2=9.275 $Y2=1.51
r330 75 76 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.1
+ $Y=1.51 $X2=9.1 $Y2=1.51
r331 73 75 17.8105 $w=3.28e-07 $l=5.1e-07 $layer=LI1_cond $X=8.59 $Y=1.51
+ $X2=9.1 $Y2=1.51
r332 71 73 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=8.505 $Y=1.675
+ $X2=8.59 $Y2=1.51
r333 71 72 79.5936 $w=1.68e-07 $l=1.22e-06 $layer=LI1_cond $X=8.505 $Y=1.675
+ $X2=8.505 $Y2=2.895
r334 69 72 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.42 $Y=2.98
+ $X2=8.505 $Y2=2.895
r335 69 70 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=8.42 $Y=2.98
+ $X2=7.81 $Y2=2.98
r336 68 70 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.725 $Y=2.895
+ $X2=7.81 $Y2=2.98
r337 67 68 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=7.725 $Y=2.055
+ $X2=7.725 $Y2=2.895
r338 66 86 4.061 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=6.155 $Y=1.97
+ $X2=6.005 $Y2=1.97
r339 65 67 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.64 $Y=1.97
+ $X2=7.725 $Y2=2.055
r340 65 66 96.8824 $w=1.68e-07 $l=1.485e-06 $layer=LI1_cond $X=7.64 $Y=1.97
+ $X2=6.155 $Y2=1.97
r341 63 96 30.6007 $w=3.3e-07 $l=1.75e-07 $layer=POLY_cond $X=12.855 $Y=0.255
+ $X2=12.855 $Y2=0.43
r342 63 64 5.03009 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=12.855 $Y=0.255
+ $X2=12.855 $Y2=0.18
r343 59 60 31.6743 $w=1.75e-07 $l=1.15e-07 $layer=POLY_cond $X=4.91 $Y=2.142
+ $X2=5.025 $Y2=2.142
r344 56 100 0.344503 $w=3.35e-07 $l=2e-09 $layer=POLY_cond $X=14.667 $Y=0.428
+ $X2=14.667 $Y2=0.43
r345 55 56 29.7995 $w=3.35e-07 $l=1.73e-07 $layer=POLY_cond $X=14.667 $Y=0.255
+ $X2=14.667 $Y2=0.428
r346 54 64 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=13.02 $Y=0.18
+ $X2=12.855 $Y2=0.18
r347 53 55 32.3722 $w=1.5e-07 $l=2.01032e-07 $layer=POLY_cond $X=14.5 $Y=0.18
+ $X2=14.667 $Y2=0.255
r348 53 54 758.894 $w=1.5e-07 $l=1.48e-06 $layer=POLY_cond $X=14.5 $Y=0.18
+ $X2=13.02 $Y2=0.18
r349 52 62 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=11.7 $Y=0.18
+ $X2=11.625 $Y2=0.18
r350 51 64 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=12.69 $Y=0.18
+ $X2=12.855 $Y2=0.18
r351 51 52 507.638 $w=1.5e-07 $l=9.9e-07 $layer=POLY_cond $X=12.69 $Y=0.18
+ $X2=11.7 $Y2=0.18
r352 47 62 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=11.625 $Y=0.255
+ $X2=11.625 $Y2=0.18
r353 47 49 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=11.625 $Y=0.255
+ $X2=11.625 $Y2=0.915
r354 43 45 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=11.31 $Y=2.985
+ $X2=11.31 $Y2=2.355
r355 41 43 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=11.235 $Y=3.06
+ $X2=11.31 $Y2=2.985
r356 41 42 464.053 $w=1.5e-07 $l=9.05e-07 $layer=POLY_cond $X=11.235 $Y=3.06
+ $X2=10.33 $Y2=3.06
r357 39 62 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=11.55 $Y=0.18
+ $X2=11.625 $Y2=0.18
r358 39 40 625.574 $w=1.5e-07 $l=1.22e-06 $layer=POLY_cond $X=11.55 $Y=0.18
+ $X2=10.33 $Y2=0.18
r359 38 42 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=10.255 $Y=2.985
+ $X2=10.33 $Y2=3.06
r360 37 61 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=10.255 $Y=1.495
+ $X2=10.255 $Y2=1.42
r361 37 38 764.021 $w=1.5e-07 $l=1.49e-06 $layer=POLY_cond $X=10.255 $Y=1.495
+ $X2=10.255 $Y2=2.985
r362 36 61 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=10.255 $Y=1.345
+ $X2=10.255 $Y2=1.42
r363 35 40 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=10.255 $Y=0.255
+ $X2=10.33 $Y2=0.18
r364 35 36 558.915 $w=1.5e-07 $l=1.09e-06 $layer=POLY_cond $X=10.255 $Y=0.255
+ $X2=10.255 $Y2=1.345
r365 33 61 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=10.18 $Y=1.42
+ $X2=10.255 $Y2=1.42
r366 33 34 199.979 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=10.18 $Y=1.42
+ $X2=9.79 $Y2=1.42
r367 29 34 24.674 $w=3.13e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.715 $Y=1.345
+ $X2=9.79 $Y2=1.42
r368 29 120 12.3195 $w=3.13e-07 $l=2.0106e-07 $layer=POLY_cond $X=9.715 $Y=1.345
+ $X2=9.635 $Y2=1.51
r369 29 31 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=9.715 $Y=1.345
+ $X2=9.715 $Y2=0.655
r370 25 120 19.9686 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.635 $Y=1.675
+ $X2=9.635 $Y2=1.51
r371 25 27 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=9.635 $Y=1.675
+ $X2=9.635 $Y2=2.465
r372 21 119 19.9686 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.325 $Y=1.345
+ $X2=9.325 $Y2=1.51
r373 21 23 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=9.325 $Y=1.345
+ $X2=9.325 $Y2=0.655
r374 17 118 19.9686 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.275 $Y=1.675
+ $X2=9.275 $Y2=1.51
r375 17 19 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=9.275 $Y=1.675
+ $X2=9.275 $Y2=2.465
r376 16 60 19.153 $w=1.95e-07 $l=7.5e-08 $layer=POLY_cond $X=5.1 $Y=2.142
+ $X2=5.025 $Y2=2.142
r377 15 115 15.146 $w=1.95e-07 $l=1.65e-07 $layer=POLY_cond $X=5.825 $Y=2.142
+ $X2=5.99 $Y2=2.142
r378 15 16 246.557 $w=1.95e-07 $l=7.25e-07 $layer=POLY_cond $X=5.825 $Y=2.142
+ $X2=5.1 $Y2=2.142
r379 11 60 6.48137 $w=1.5e-07 $l=9.8e-08 $layer=POLY_cond $X=5.025 $Y=2.24
+ $X2=5.025 $Y2=2.142
r380 11 13 217.926 $w=1.5e-07 $l=4.25e-07 $layer=POLY_cond $X=5.025 $Y=2.24
+ $X2=5.025 $Y2=2.665
r381 7 59 6.48137 $w=1.5e-07 $l=9.7e-08 $layer=POLY_cond $X=4.91 $Y=2.045
+ $X2=4.91 $Y2=2.142
r382 7 9 379.447 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=4.91 $Y=2.045
+ $X2=4.91 $Y2=1.305
r383 2 84 400 $w=1.7e-07 $l=1.18528e-06 $layer=licon1_PDIFF $count=1 $X=14.94
+ $Y=1.785 $X2=15.085 $Y2=2.9
r384 2 82 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=14.94
+ $Y=1.785 $X2=15.085 $Y2=1.93
r385 1 103 182 $w=1.7e-07 $l=3.14245e-07 $layer=licon1_NDIFF $count=1 $X=14.94
+ $Y=0.235 $X2=15.085 $Y2=0.485
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRBP_LP%A_1147_490# 1 2 3 4 13 15 16 17 20 22 23
+ 27 29 32 33 34 36 37 38 41 44 45 49 52 59 61 65
c194 59 0 2.88191e-20 $X=11.165 $Y=1.17
c195 32 0 9.44178e-20 $X=9.5 $Y=2.895
c196 29 0 1.85423e-19 $X=9.415 $Y=1.08
c197 27 0 1.14841e-19 $X=8.075 $Y=2.02
c198 23 0 6.21055e-20 $X=7.85 $Y=1.15
r199 61 63 16.8276 $w=2.61e-07 $l=3.6e-07 $layer=LI1_cond $X=11.165 $Y=2.08
+ $X2=11.525 $Y2=2.08
r200 55 56 3.99225 $w=3.88e-07 $l=8.5e-08 $layer=LI1_cond $X=8.045 $Y=1.15
+ $X2=8.045 $Y2=1.235
r201 54 55 2.06849 $w=3.88e-07 $l=7e-08 $layer=LI1_cond $X=8.045 $Y=1.08
+ $X2=8.045 $Y2=1.15
r202 52 54 6.64871 $w=3.88e-07 $l=2.25e-07 $layer=LI1_cond $X=8.045 $Y=0.855
+ $X2=8.045 $Y2=1.08
r203 49 66 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.35 $Y=1.29
+ $X2=6.35 $Y2=1.455
r204 49 65 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.35 $Y=1.29
+ $X2=6.35 $Y2=1.125
r205 48 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.35
+ $Y=1.29 $X2=6.35 $Y2=1.29
r206 45 48 4.88915 $w=3.28e-07 $l=1.4e-07 $layer=LI1_cond $X=6.35 $Y=1.15
+ $X2=6.35 $Y2=1.29
r207 44 61 3.24614 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.165 $Y=1.915
+ $X2=11.165 $Y2=2.08
r208 43 59 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.165 $Y=1.255
+ $X2=11.165 $Y2=1.17
r209 43 44 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=11.165 $Y=1.255
+ $X2=11.165 $Y2=1.915
r210 39 59 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=10.785 $Y=1.17
+ $X2=11.165 $Y2=1.17
r211 39 41 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=10.785 $Y=1.085
+ $X2=10.785 $Y2=0.74
r212 37 61 5.45457 $w=2.61e-07 $l=1.07121e-07 $layer=LI1_cond $X=11.08 $Y=2.03
+ $X2=11.165 $Y2=2.08
r213 37 38 51.8663 $w=1.68e-07 $l=7.95e-07 $layer=LI1_cond $X=11.08 $Y=2.03
+ $X2=10.285 $Y2=2.03
r214 35 38 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.2 $Y=2.115
+ $X2=10.285 $Y2=2.03
r215 35 36 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=10.2 $Y=2.115
+ $X2=10.2 $Y2=2.895
r216 33 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.115 $Y=2.98
+ $X2=10.2 $Y2=2.895
r217 33 34 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=10.115 $Y=2.98
+ $X2=9.585 $Y2=2.98
r218 32 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.5 $Y=2.895
+ $X2=9.585 $Y2=2.98
r219 31 32 112.866 $w=1.68e-07 $l=1.73e-06 $layer=LI1_cond $X=9.5 $Y=1.165
+ $X2=9.5 $Y2=2.895
r220 30 54 5.6248 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=8.24 $Y=1.08
+ $X2=8.045 $Y2=1.08
r221 29 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.415 $Y=1.08
+ $X2=9.5 $Y2=1.165
r222 29 30 76.6578 $w=1.68e-07 $l=1.175e-06 $layer=LI1_cond $X=9.415 $Y=1.08
+ $X2=8.24 $Y2=1.08
r223 27 56 36.1867 $w=2.48e-07 $l=7.85e-07 $layer=LI1_cond $X=8.115 $Y=2.02
+ $X2=8.115 $Y2=1.235
r224 24 45 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.515 $Y=1.15
+ $X2=6.35 $Y2=1.15
r225 23 55 5.6248 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=7.85 $Y=1.15
+ $X2=8.045 $Y2=1.15
r226 23 24 87.0963 $w=1.68e-07 $l=1.335e-06 $layer=LI1_cond $X=7.85 $Y=1.15
+ $X2=6.515 $Y2=1.15
r227 22 66 510.202 $w=1.5e-07 $l=9.95e-07 $layer=POLY_cond $X=6.44 $Y=2.45
+ $X2=6.44 $Y2=1.455
r228 20 65 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=6.44 $Y=0.805
+ $X2=6.44 $Y2=1.125
r229 16 22 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.365 $Y=2.525
+ $X2=6.44 $Y2=2.45
r230 16 17 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=6.365 $Y=2.525
+ $X2=5.885 $Y2=2.525
r231 13 17 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.81 $Y=2.6
+ $X2=5.885 $Y2=2.525
r232 13 15 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=5.81 $Y=2.6 $X2=5.81
+ $Y2=2.885
r233 4 63 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=11.385
+ $Y=1.935 $X2=11.525 $Y2=2.08
r234 3 27 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=7.93
+ $Y=1.875 $X2=8.075 $Y2=2.02
r235 2 41 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=10.64
+ $Y=0.595 $X2=10.785 $Y2=0.74
r236 1 52 182 $w=1.7e-07 $l=4.87134e-07 $layer=licon1_NDIFF $count=1 $X=7.87
+ $Y=0.435 $X2=8.015 $Y2=0.855
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRBP_LP%RESET_B 1 3 4 5 9 12 13 14 16 19 24 27 31
+ 34 37 41 45 48 49 50 53 55 56 57 58 63 64 66 69 70 74 75 82
c258 63 0 1.69588e-19 $X=14.16 $Y=2.405
c259 57 0 2.90512e-20 $X=14.015 $Y=2.405
c260 56 0 1.62564e-19 $X=4.225 $Y=2.405
c261 53 0 6.46456e-20 $X=13.52 $Y=1.7
c262 41 0 1.0756e-19 $X=13.88 $Y=2.8
c263 34 0 1.29974e-19 $X=13.52 $Y=2.1
c264 31 0 1.29593e-19 $X=13.335 $Y=0.915
c265 24 0 1.28843e-19 $X=6.83 $Y=0.805
r266 80 82 8.74306 $w=3.3e-07 $l=5e-08 $layer=POLY_cond $X=13.83 $Y=2.265
+ $X2=13.88 $Y2=2.265
r267 80 81 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=13.83
+ $Y=2.265 $X2=13.83 $Y2=2.265
r268 77 80 54.207 $w=3.3e-07 $l=3.1e-07 $layer=POLY_cond $X=13.52 $Y=2.265
+ $X2=13.83 $Y2=2.265
r269 74 76 36.2633 $w=3.19e-07 $l=2.4e-07 $layer=POLY_cond $X=6.92 $Y=2.35
+ $X2=7.16 $Y2=2.35
r270 74 75 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.92
+ $Y=2.35 $X2=6.92 $Y2=2.35
r271 72 74 13.5987 $w=3.19e-07 $l=9e-08 $layer=POLY_cond $X=6.83 $Y=2.35
+ $X2=6.92 $Y2=2.35
r272 71 72 4.53292 $w=3.19e-07 $l=3e-08 $layer=POLY_cond $X=6.8 $Y=2.35 $X2=6.83
+ $Y2=2.35
r273 70 87 21.4773 $w=3.28e-07 $l=6.15e-07 $layer=LI1_cond $X=4.03 $Y=1.79
+ $X2=4.03 $Y2=2.405
r274 69 70 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.03
+ $Y=1.79 $X2=4.03 $Y2=1.79
r275 66 87 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=2.405
+ $X2=4.08 $Y2=2.405
r276 64 81 9.05491 $w=4.18e-07 $l=3.3e-07 $layer=LI1_cond $X=14.16 $Y=2.31
+ $X2=13.83 $Y2=2.31
r277 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.16 $Y=2.405
+ $X2=14.16 $Y2=2.405
r278 60 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=2.405
+ $X2=6.96 $Y2=2.405
r279 58 60 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.105 $Y=2.405
+ $X2=6.96 $Y2=2.405
r280 57 63 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=14.015 $Y=2.405
+ $X2=14.16 $Y2=2.405
r281 57 58 8.55196 $w=1.4e-07 $l=6.91e-06 $layer=MET1_cond $X=14.015 $Y=2.405
+ $X2=7.105 $Y2=2.405
r282 56 66 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.225 $Y=2.405
+ $X2=4.08 $Y2=2.405
r283 55 60 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.815 $Y=2.405
+ $X2=6.96 $Y2=2.405
r284 55 56 3.20544 $w=1.4e-07 $l=2.59e-06 $layer=MET1_cond $X=6.815 $Y=2.405
+ $X2=4.225 $Y2=2.405
r285 51 53 94.8617 $w=1.5e-07 $l=1.85e-07 $layer=POLY_cond $X=13.335 $Y=1.7
+ $X2=13.52 $Y2=1.7
r286 49 69 70.8188 $w=3.3e-07 $l=4.05e-07 $layer=POLY_cond $X=4.03 $Y=2.195
+ $X2=4.03 $Y2=1.79
r287 49 50 13.5877 $w=2.4e-07 $l=7.5e-08 $layer=POLY_cond $X=4.03 $Y=2.195
+ $X2=4.03 $Y2=2.27
r288 48 69 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.03 $Y=1.625
+ $X2=4.03 $Y2=1.79
r289 43 45 51.2766 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=3.84 $Y=0.9 $X2=3.94
+ $Y2=0.9
r290 39 82 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=13.88 $Y=2.43
+ $X2=13.88 $Y2=2.265
r291 39 41 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=13.88 $Y=2.43
+ $X2=13.88 $Y2=2.8
r292 35 77 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=13.52 $Y=2.43
+ $X2=13.52 $Y2=2.265
r293 35 37 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=13.52 $Y=2.43
+ $X2=13.52 $Y2=2.8
r294 34 77 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=13.52 $Y=2.1
+ $X2=13.52 $Y2=2.265
r295 33 53 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=13.52 $Y=1.775
+ $X2=13.52 $Y2=1.7
r296 33 34 166.649 $w=1.5e-07 $l=3.25e-07 $layer=POLY_cond $X=13.52 $Y=1.775
+ $X2=13.52 $Y2=2.1
r297 29 51 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=13.335 $Y=1.625
+ $X2=13.335 $Y2=1.7
r298 29 31 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=13.335 $Y=1.625
+ $X2=13.335 $Y2=0.915
r299 25 76 20.418 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.16 $Y=2.515
+ $X2=7.16 $Y2=2.35
r300 25 27 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=7.16 $Y=2.515
+ $X2=7.16 $Y2=2.885
r301 22 72 20.418 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.83 $Y=2.185
+ $X2=6.83 $Y2=2.35
r302 22 24 707.617 $w=1.5e-07 $l=1.38e-06 $layer=POLY_cond $X=6.83 $Y=2.185
+ $X2=6.83 $Y2=0.805
r303 21 24 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=6.83 $Y=0.255
+ $X2=6.83 $Y2=0.805
r304 17 71 20.418 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.8 $Y=2.515
+ $X2=6.8 $Y2=2.35
r305 17 19 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=6.8 $Y=2.515
+ $X2=6.8 $Y2=2.885
r306 14 50 13.5877 $w=2.4e-07 $l=9.28709e-08 $layer=POLY_cond $X=3.99 $Y=2.345
+ $X2=4.03 $Y2=2.27
r307 14 16 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=3.99 $Y=2.345
+ $X2=3.99 $Y2=2.775
r308 12 21 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.755 $Y=0.18
+ $X2=6.83 $Y2=0.255
r309 12 13 1456.26 $w=1.5e-07 $l=2.84e-06 $layer=POLY_cond $X=6.755 $Y=0.18
+ $X2=3.915 $Y2=0.18
r310 10 45 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.94 $Y=0.975
+ $X2=3.94 $Y2=0.9
r311 10 48 333.298 $w=1.5e-07 $l=6.5e-07 $layer=POLY_cond $X=3.94 $Y=0.975
+ $X2=3.94 $Y2=1.625
r312 7 43 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.84 $Y=0.825
+ $X2=3.84 $Y2=0.9
r313 7 9 146.138 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.84 $Y=0.825
+ $X2=3.84 $Y2=0.54
r314 6 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.84 $Y=0.255
+ $X2=3.915 $Y2=0.18
r315 6 9 146.138 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.84 $Y=0.255
+ $X2=3.84 $Y2=0.54
r316 4 50 12.1617 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.865 $Y=2.27
+ $X2=4.03 $Y2=2.27
r317 4 5 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=3.865 $Y=2.27
+ $X2=3.675 $Y2=2.27
r318 1 5 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.6 $Y=2.345
+ $X2=3.675 $Y2=2.27
r319 1 3 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=3.6 $Y=2.345 $X2=3.6
+ $Y2=2.775
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRBP_LP%A_911_219# 1 2 3 10 14 18 20 24 28 30 31
+ 34 36 38 39 41 43 44 46 49 50 51 55 56 57 58 64 69
c186 69 0 2.90512e-20 $X=7.645 $Y=1.46
c187 31 0 2.7984e-19 $X=8.635 $Y=1.46
c188 24 0 3.6059e-20 $X=8.62 $Y=0.755
r189 65 69 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=7.645 $Y=1.55
+ $X2=7.645 $Y2=1.46
r190 64 67 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=7.645 $Y=1.55
+ $X2=7.645 $Y2=1.63
r191 64 65 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.645
+ $Y=1.55 $X2=7.645 $Y2=1.55
r192 58 61 4.37928 $w=2.48e-07 $l=9.5e-08 $layer=LI1_cond $X=7.335 $Y=2.785
+ $X2=7.335 $Y2=2.88
r193 53 55 8.48463 $w=2.98e-07 $l=1.65e-07 $layer=LI1_cond $X=4.695 $Y=1.385
+ $X2=4.86 $Y2=1.385
r194 50 58 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.21 $Y=2.785
+ $X2=7.335 $Y2=2.785
r195 50 51 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=7.21 $Y=2.785
+ $X2=6.54 $Y2=2.785
r196 49 51 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.455 $Y=2.7
+ $X2=6.54 $Y2=2.785
r197 48 49 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=6.455 $Y=2.555
+ $X2=6.455 $Y2=2.7
r198 47 57 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.675 $Y=2.47
+ $X2=5.59 $Y2=2.47
r199 46 48 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.37 $Y=2.47
+ $X2=6.455 $Y2=2.555
r200 46 47 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=6.37 $Y=2.47
+ $X2=5.675 $Y2=2.47
r201 45 56 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.675 $Y=1.63
+ $X2=5.59 $Y2=1.63
r202 44 67 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.48 $Y=1.63
+ $X2=7.645 $Y2=1.63
r203 44 45 117.759 $w=1.68e-07 $l=1.805e-06 $layer=LI1_cond $X=7.48 $Y=1.63
+ $X2=5.675 $Y2=1.63
r204 43 57 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.59 $Y=2.385
+ $X2=5.59 $Y2=2.47
r205 42 56 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.59 $Y=1.715
+ $X2=5.59 $Y2=1.63
r206 42 43 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.59 $Y=1.715
+ $X2=5.59 $Y2=2.385
r207 41 56 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.59 $Y=1.545
+ $X2=5.59 $Y2=1.63
r208 40 41 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=5.59 $Y=1.405
+ $X2=5.59 $Y2=1.545
r209 38 57 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.505 $Y=2.47
+ $X2=5.59 $Y2=2.47
r210 38 39 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=5.505 $Y=2.47
+ $X2=4.905 $Y2=2.47
r211 36 40 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.505 $Y=1.32
+ $X2=5.59 $Y2=1.405
r212 36 55 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=5.505 $Y=1.32
+ $X2=4.86 $Y2=1.32
r213 32 39 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=4.81 $Y=2.555
+ $X2=4.905 $Y2=2.47
r214 32 34 6.42105 $w=1.88e-07 $l=1.1e-07 $layer=LI1_cond $X=4.81 $Y=2.555
+ $X2=4.81 $Y2=2.665
r215 26 31 20.4101 $w=1.5e-07 $l=8.21584e-08 $layer=POLY_cond $X=8.65 $Y=1.535
+ $X2=8.635 $Y2=1.46
r216 26 28 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=8.65 $Y=1.535
+ $X2=8.65 $Y2=2.295
r217 22 31 20.4101 $w=1.5e-07 $l=8.21584e-08 $layer=POLY_cond $X=8.62 $Y=1.385
+ $X2=8.635 $Y2=1.46
r218 22 24 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=8.62 $Y=1.385
+ $X2=8.62 $Y2=0.755
r219 21 30 12.05 $w=1.5e-07 $l=1.05e-07 $layer=POLY_cond $X=8.365 $Y=1.46
+ $X2=8.26 $Y2=1.46
r220 20 31 5.30422 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=8.545 $Y=1.46
+ $X2=8.635 $Y2=1.46
r221 20 21 92.2979 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=8.545 $Y=1.46
+ $X2=8.365 $Y2=1.46
r222 16 30 12.05 $w=1.5e-07 $l=8.87412e-08 $layer=POLY_cond $X=8.29 $Y=1.535
+ $X2=8.26 $Y2=1.46
r223 16 18 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=8.29 $Y=1.535
+ $X2=8.29 $Y2=2.295
r224 12 30 12.05 $w=1.5e-07 $l=8.87412e-08 $layer=POLY_cond $X=8.23 $Y=1.385
+ $X2=8.26 $Y2=1.46
r225 12 14 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=8.23 $Y=1.385
+ $X2=8.23 $Y2=0.755
r226 11 69 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.81 $Y=1.46
+ $X2=7.645 $Y2=1.46
r227 10 30 12.05 $w=1.5e-07 $l=1.05e-07 $layer=POLY_cond $X=8.155 $Y=1.46
+ $X2=8.26 $Y2=1.46
r228 10 11 176.904 $w=1.5e-07 $l=3.45e-07 $layer=POLY_cond $X=8.155 $Y=1.46
+ $X2=7.81 $Y2=1.46
r229 3 61 600 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=1 $X=7.235
+ $Y=2.675 $X2=7.375 $Y2=2.88
r230 2 34 600 $w=1.7e-07 $l=3.44347e-07 $layer=licon1_PDIFF $count=1 $X=4.555
+ $Y=2.455 $X2=4.81 $Y2=2.665
r231 1 53 182 $w=1.7e-07 $l=3.27605e-07 $layer=licon1_NDIFF $count=1 $X=4.555
+ $Y=1.095 $X2=4.695 $Y2=1.36
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRBP_LP%A_2388_115# 1 2 7 9 14 18 21 23 24 25 29
+ 32 33 37 42 47 50
c110 47 0 2.42792e-20 $X=12.275 $Y=2.185
c111 21 0 1.69588e-19 $X=13.14 $Y=2.53
c112 18 0 8.97349e-20 $X=12.305 $Y=1.4
r113 42 44 4.84026 $w=2.48e-07 $l=1.05e-07 $layer=LI1_cond $X=14.015 $Y=0.87
+ $X2=14.015 $Y2=0.975
r114 37 39 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=12.775 $Y=0.975
+ $X2=12.775 $Y2=1.135
r115 33 48 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=12.275 $Y=2.35
+ $X2=12.275 $Y2=2.515
r116 33 47 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=12.275 $Y=2.35
+ $X2=12.275 $Y2=2.185
r117 32 35 7.54326 $w=2.73e-07 $l=1.8e-07 $layer=LI1_cond $X=12.277 $Y=2.35
+ $X2=12.277 $Y2=2.53
r118 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=12.275
+ $Y=2.35 $X2=12.275 $Y2=2.35
r119 27 29 6.46067 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=13.305 $Y=2.615
+ $X2=13.305 $Y2=2.8
r120 26 37 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=12.86 $Y=0.975
+ $X2=12.775 $Y2=0.975
r121 25 44 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=13.89 $Y=0.975
+ $X2=14.015 $Y2=0.975
r122 25 26 67.1979 $w=1.68e-07 $l=1.03e-06 $layer=LI1_cond $X=13.89 $Y=0.975
+ $X2=12.86 $Y2=0.975
r123 23 39 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=12.69 $Y=1.135
+ $X2=12.775 $Y2=1.135
r124 23 24 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=12.69 $Y=1.135
+ $X2=12.47 $Y2=1.135
r125 22 35 3.55113 $w=1.7e-07 $l=1.38e-07 $layer=LI1_cond $X=12.415 $Y=2.53
+ $X2=12.277 $Y2=2.53
r126 21 27 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=13.14 $Y=2.53
+ $X2=13.305 $Y2=2.615
r127 21 22 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=13.14 $Y=2.53
+ $X2=12.415 $Y2=2.53
r128 19 50 21.2647 $w=2.72e-07 $l=1.2e-07 $layer=POLY_cond $X=12.305 $Y=1.4
+ $X2=12.185 $Y2=1.4
r129 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=12.305
+ $Y=1.4 $X2=12.305 $Y2=1.4
r130 16 24 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=12.305 $Y=1.22
+ $X2=12.47 $Y2=1.135
r131 16 18 6.28605 $w=3.28e-07 $l=1.8e-07 $layer=LI1_cond $X=12.305 $Y=1.22
+ $X2=12.305 $Y2=1.4
r132 14 48 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=12.365 $Y=2.885
+ $X2=12.365 $Y2=2.515
r133 10 50 16.6763 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=12.185 $Y=1.565
+ $X2=12.185 $Y2=1.4
r134 10 47 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=12.185 $Y=1.565
+ $X2=12.185 $Y2=2.185
r135 7 50 30.125 $w=2.72e-07 $l=2.38642e-07 $layer=POLY_cond $X=12.015 $Y=1.235
+ $X2=12.185 $Y2=1.4
r136 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=12.015 $Y=1.235
+ $X2=12.015 $Y2=0.915
r137 2 29 600 $w=1.7e-07 $l=9.33836e-07 $layer=licon1_PDIFF $count=1 $X=13.05
+ $Y=1.985 $X2=13.305 $Y2=2.8
r138 1 42 182 $w=1.7e-07 $l=3.27261e-07 $layer=licon1_NDIFF $count=1 $X=13.8
+ $Y=0.705 $X2=14.055 $Y2=0.87
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRBP_LP%A_2168_439# 1 2 9 11 13 14 15 18 22 26 30
+ 34 36 40 44 46 50 54 56 57 58 62 65 67 68 73 74 76 78 79 80 86 87 91 92 95 97
+ 102 110
c244 79 0 1.97521e-19 $X=16.015 $Y=0.975
c245 76 0 2.42792e-20 $X=13.05 $Y=1.485
c246 74 0 8.97349e-20 $X=12.885 $Y=1.66
c247 68 0 1.9462e-19 $X=12.72 $Y=1.83
c248 9 0 1.41841e-19 $X=12.975 $Y=2.195
r249 109 110 30.474 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=16.45 $Y=1.42
+ $X2=16.525 $Y2=1.42
r250 96 109 47.2125 $w=3.3e-07 $l=2.7e-07 $layer=POLY_cond $X=16.18 $Y=1.42
+ $X2=16.45 $Y2=1.42
r251 96 106 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=16.18 $Y=1.42
+ $X2=16.09 $Y2=1.42
r252 95 97 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=16.18 $Y=1.42
+ $X2=16.18 $Y2=1.255
r253 95 96 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=16.18
+ $Y=1.42 $X2=16.18 $Y2=1.42
r254 90 105 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=14.22 $Y=1.405
+ $X2=14.22 $Y2=1.57
r255 90 102 16.6118 $w=3.3e-07 $l=9.5e-08 $layer=POLY_cond $X=14.22 $Y=1.405
+ $X2=14.22 $Y2=1.31
r256 89 92 6.46067 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=14.22 $Y=1.405
+ $X2=14.405 $Y2=1.405
r257 89 91 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=14.22 $Y=1.405
+ $X2=14.055 $Y2=1.405
r258 89 90 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=14.22
+ $Y=1.405 $X2=14.22 $Y2=1.405
r259 84 86 8.51388 $w=2.88e-07 $l=1.65e-07 $layer=LI1_cond $X=11.095 $Y=2.57
+ $X2=11.26 $Y2=2.57
r260 81 97 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=16.1 $Y=1.06
+ $X2=16.1 $Y2=1.255
r261 79 81 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=16.015 $Y=0.975
+ $X2=16.1 $Y2=1.06
r262 79 80 99.492 $w=1.68e-07 $l=1.525e-06 $layer=LI1_cond $X=16.015 $Y=0.975
+ $X2=14.49 $Y2=0.975
r263 78 92 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=14.405 $Y=1.24
+ $X2=14.405 $Y2=1.405
r264 77 80 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=14.405 $Y=1.06
+ $X2=14.49 $Y2=0.975
r265 77 78 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=14.405 $Y=1.06
+ $X2=14.405 $Y2=1.24
r266 76 91 65.5668 $w=1.68e-07 $l=1.005e-06 $layer=LI1_cond $X=13.05 $Y=1.485
+ $X2=14.055 $Y2=1.485
r267 74 101 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=12.885 $Y=1.66
+ $X2=12.885 $Y2=1.825
r268 73 74 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=12.885
+ $Y=1.66 $X2=12.885 $Y2=1.66
r269 71 73 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=12.885 $Y=1.745
+ $X2=12.885 $Y2=1.66
r270 70 76 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=12.885 $Y=1.57
+ $X2=13.05 $Y2=1.485
r271 70 73 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=12.885 $Y=1.57
+ $X2=12.885 $Y2=1.66
r272 69 87 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.96 $Y=1.83
+ $X2=11.875 $Y2=1.83
r273 68 71 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=12.72 $Y=1.83
+ $X2=12.885 $Y2=1.745
r274 68 69 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=12.72 $Y=1.83
+ $X2=11.96 $Y2=1.83
r275 66 87 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.875 $Y=1.915
+ $X2=11.875 $Y2=1.83
r276 66 67 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=11.875 $Y=1.915
+ $X2=11.875 $Y2=2.425
r277 65 87 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.875 $Y=1.745
+ $X2=11.875 $Y2=1.83
r278 64 65 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=11.875 $Y=0.905
+ $X2=11.875 $Y2=1.745
r279 62 67 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=11.79 $Y=2.51
+ $X2=11.875 $Y2=2.425
r280 62 86 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=11.79 $Y=2.51
+ $X2=11.26 $Y2=2.51
r281 58 64 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=11.79 $Y=0.74
+ $X2=11.875 $Y2=0.905
r282 58 60 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=11.79 $Y=0.74
+ $X2=11.295 $Y2=0.74
r283 52 57 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=17.8 $Y=1.405
+ $X2=17.8 $Y2=1.33
r284 52 54 384.574 $w=1.5e-07 $l=7.5e-07 $layer=POLY_cond $X=17.8 $Y=1.405
+ $X2=17.8 $Y2=2.155
r285 48 57 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=17.8 $Y=1.255
+ $X2=17.8 $Y2=1.33
r286 48 50 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=17.8 $Y=1.255
+ $X2=17.8 $Y2=0.895
r287 47 56 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=17.515 $Y=1.33
+ $X2=17.44 $Y2=1.33
r288 46 57 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=17.725 $Y=1.33
+ $X2=17.8 $Y2=1.33
r289 46 47 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=17.725 $Y=1.33
+ $X2=17.515 $Y2=1.33
r290 42 56 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=17.44 $Y=1.405
+ $X2=17.44 $Y2=1.33
r291 42 44 384.574 $w=1.5e-07 $l=7.5e-07 $layer=POLY_cond $X=17.44 $Y=1.405
+ $X2=17.44 $Y2=2.155
r292 38 56 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=17.44 $Y=1.255
+ $X2=17.44 $Y2=1.33
r293 38 40 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=17.44 $Y=1.255
+ $X2=17.44 $Y2=0.895
r294 36 56 24.1 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=17.365 $Y=1.33
+ $X2=17.44 $Y2=1.33
r295 36 110 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=17.365 $Y=1.33
+ $X2=16.525 $Y2=1.33
r296 32 109 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=16.45 $Y=1.585
+ $X2=16.45 $Y2=1.42
r297 32 34 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=16.45 $Y=1.585
+ $X2=16.45 $Y2=2.415
r298 28 109 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=16.45 $Y=1.255
+ $X2=16.45 $Y2=1.42
r299 28 30 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=16.45 $Y=1.255
+ $X2=16.45 $Y2=0.655
r300 24 106 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=16.09 $Y=1.585
+ $X2=16.09 $Y2=1.42
r301 24 26 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=16.09 $Y=1.585
+ $X2=16.09 $Y2=2.415
r302 20 106 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=16.09 $Y=1.255
+ $X2=16.09 $Y2=1.42
r303 20 22 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=16.09 $Y=1.255
+ $X2=16.09 $Y2=0.655
r304 18 105 630.702 $w=1.5e-07 $l=1.23e-06 $layer=POLY_cond $X=14.31 $Y=2.8
+ $X2=14.31 $Y2=1.57
r305 14 102 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=14.055 $Y=1.31
+ $X2=14.22 $Y2=1.31
r306 14 15 130.755 $w=1.5e-07 $l=2.55e-07 $layer=POLY_cond $X=14.055 $Y=1.31
+ $X2=13.8 $Y2=1.31
r307 11 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=13.725 $Y=1.235
+ $X2=13.8 $Y2=1.31
r308 11 13 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=13.725 $Y=1.235
+ $X2=13.725 $Y2=0.915
r309 9 101 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=12.975 $Y=2.195
+ $X2=12.975 $Y2=1.825
r310 2 84 600 $w=1.7e-07 $l=4.86056e-07 $layer=licon1_PDIFF $count=1 $X=10.84
+ $Y=2.195 $X2=11.095 $Y2=2.57
r311 1 60 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=11.155
+ $Y=0.595 $X2=11.295 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRBP_LP%CLK 3 7 11 15 17 23 24
c46 24 0 1.97521e-19 $X=15.66 $Y=1.46
c47 23 0 1.70221e-19 $X=15.595 $Y=1.46
r48 22 24 11.366 $w=3.3e-07 $l=6.5e-08 $layer=POLY_cond $X=15.595 $Y=1.46
+ $X2=15.66 $Y2=1.46
r49 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=15.595
+ $Y=1.46 $X2=15.595 $Y2=1.46
r50 19 22 51.5841 $w=3.3e-07 $l=2.95e-07 $layer=POLY_cond $X=15.3 $Y=1.46
+ $X2=15.595 $Y2=1.46
r51 17 23 7.15912 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=15.595 $Y=1.665
+ $X2=15.595 $Y2=1.46
r52 13 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=15.66 $Y=1.625
+ $X2=15.66 $Y2=1.46
r53 13 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=15.66 $Y=1.625
+ $X2=15.66 $Y2=2.415
r54 9 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=15.66 $Y=1.295
+ $X2=15.66 $Y2=1.46
r55 9 11 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=15.66 $Y=1.295
+ $X2=15.66 $Y2=0.655
r56 5 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=15.3 $Y=1.625
+ $X2=15.3 $Y2=1.46
r57 5 7 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=15.3 $Y=1.625 $X2=15.3
+ $Y2=2.415
r58 1 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=15.3 $Y=1.295
+ $X2=15.3 $Y2=1.46
r59 1 3 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=15.3 $Y=1.295 $X2=15.3
+ $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRBP_LP%A_3416_137# 1 2 9 13 17 21 25 29 33 36 40
r61 34 40 51.5841 $w=3.3e-07 $l=2.95e-07 $layer=POLY_cond $X=18.41 $Y=1.47
+ $X2=18.705 $Y2=1.47
r62 34 37 11.366 $w=3.3e-07 $l=6.5e-08 $layer=POLY_cond $X=18.41 $Y=1.47
+ $X2=18.345 $Y2=1.47
r63 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=18.41
+ $Y=1.47 $X2=18.41 $Y2=1.47
r64 31 36 1.34256 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=17.39 $Y=1.47
+ $X2=17.225 $Y2=1.47
r65 31 33 35.621 $w=3.28e-07 $l=1.02e-06 $layer=LI1_cond $X=17.39 $Y=1.47
+ $X2=18.41 $Y2=1.47
r66 27 36 5.16603 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=17.225 $Y=1.635
+ $X2=17.225 $Y2=1.47
r67 27 29 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=17.225 $Y=1.635
+ $X2=17.225 $Y2=1.98
r68 23 36 5.16603 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=17.225 $Y=1.305
+ $X2=17.225 $Y2=1.47
r69 23 25 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=17.225 $Y=1.305
+ $X2=17.225 $Y2=0.895
r70 19 40 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=18.705 $Y=1.635
+ $X2=18.705 $Y2=1.47
r71 19 21 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=18.705 $Y=1.635
+ $X2=18.705 $Y2=2.465
r72 15 40 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=18.705 $Y=1.305
+ $X2=18.705 $Y2=1.47
r73 15 17 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=18.705 $Y=1.305
+ $X2=18.705 $Y2=0.685
r74 11 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=18.345 $Y=1.635
+ $X2=18.345 $Y2=1.47
r75 11 13 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=18.345 $Y=1.635
+ $X2=18.345 $Y2=2.465
r76 7 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=18.345 $Y=1.305
+ $X2=18.345 $Y2=1.47
r77 7 9 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=18.345 $Y=1.305
+ $X2=18.345 $Y2=0.685
r78 2 29 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=17.08
+ $Y=1.835 $X2=17.225 $Y2=1.98
r79 1 25 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=17.08
+ $Y=0.685 $X2=17.225 $Y2=0.895
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRBP_LP%VPWR 1 2 3 4 5 6 7 8 27 31 35 39 45 49 53
+ 59 64 65 67 68 69 71 76 84 99 106 115 121 122 125 128 131 134 137 140
r215 140 141 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=18 $Y=3.33
+ $X2=18 $Y2=3.33
r216 137 138 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=14.16 $Y=3.33
+ $X2=14.16 $Y2=3.33
r217 134 135 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.72 $Y=3.33
+ $X2=12.72 $Y2=3.33
r218 131 132 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r219 128 129 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r220 125 126 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r221 122 141 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=18.96 $Y=3.33
+ $X2=18 $Y2=3.33
r222 121 122 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=18.96 $Y=3.33
+ $X2=18.96 $Y2=3.33
r223 119 140 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=18.295 $Y=3.33
+ $X2=18.13 $Y2=3.33
r224 119 121 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=18.295 $Y=3.33
+ $X2=18.96 $Y2=3.33
r225 118 141 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=16.08 $Y=3.33
+ $X2=18 $Y2=3.33
r226 117 118 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=16.08 $Y=3.33
+ $X2=16.08 $Y2=3.33
r227 115 140 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=17.965 $Y=3.33
+ $X2=18.13 $Y2=3.33
r228 115 117 122.979 $w=1.68e-07 $l=1.885e-06 $layer=LI1_cond $X=17.965 $Y=3.33
+ $X2=16.08 $Y2=3.33
r229 114 118 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=15.6 $Y=3.33
+ $X2=16.08 $Y2=3.33
r230 114 138 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=15.6 $Y=3.33
+ $X2=14.16 $Y2=3.33
r231 113 114 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=15.6 $Y=3.33
+ $X2=15.6 $Y2=3.33
r232 111 137 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=14.18 $Y=3.33
+ $X2=14.055 $Y2=3.33
r233 111 113 92.6417 $w=1.68e-07 $l=1.42e-06 $layer=LI1_cond $X=14.18 $Y=3.33
+ $X2=15.6 $Y2=3.33
r234 110 138 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.68 $Y=3.33
+ $X2=14.16 $Y2=3.33
r235 110 135 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=13.68 $Y=3.33
+ $X2=12.72 $Y2=3.33
r236 109 110 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=13.68 $Y=3.33
+ $X2=13.68 $Y2=3.33
r237 107 134 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.825 $Y=3.33
+ $X2=12.66 $Y2=3.33
r238 107 109 55.7807 $w=1.68e-07 $l=8.55e-07 $layer=LI1_cond $X=12.825 $Y=3.33
+ $X2=13.68 $Y2=3.33
r239 106 137 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=13.93 $Y=3.33
+ $X2=14.055 $Y2=3.33
r240 106 109 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=13.93 $Y=3.33
+ $X2=13.68 $Y2=3.33
r241 105 135 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.24 $Y=3.33
+ $X2=12.72 $Y2=3.33
r242 104 105 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=12.24
+ $Y=3.33 $X2=12.24 $Y2=3.33
r243 101 104 187.893 $w=1.68e-07 $l=2.88e-06 $layer=LI1_cond $X=9.36 $Y=3.33
+ $X2=12.24 $Y2=3.33
r244 101 102 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r245 99 134 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.495 $Y=3.33
+ $X2=12.66 $Y2=3.33
r246 99 104 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=12.495 $Y=3.33
+ $X2=12.24 $Y2=3.33
r247 98 102 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=9.36 $Y2=3.33
r248 97 98 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r249 95 98 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=8.88 $Y2=3.33
r250 95 132 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=6 $Y2=3.33
r251 94 97 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=6.48 $Y=3.33
+ $X2=8.88 $Y2=3.33
r252 94 95 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r253 92 131 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.19 $Y=3.33
+ $X2=6.025 $Y2=3.33
r254 92 94 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=6.19 $Y=3.33
+ $X2=6.48 $Y2=3.33
r255 91 132 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=6 $Y2=3.33
r256 90 91 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r257 88 91 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=5.52 $Y2=3.33
r258 88 129 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=3.12 $Y2=3.33
r259 87 90 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=3.6 $Y=3.33
+ $X2=5.52 $Y2=3.33
r260 87 88 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r261 85 128 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.225 $Y=3.33
+ $X2=3.06 $Y2=3.33
r262 85 87 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=3.225 $Y=3.33
+ $X2=3.6 $Y2=3.33
r263 84 131 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.86 $Y=3.33
+ $X2=6.025 $Y2=3.33
r264 84 90 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=5.86 $Y=3.33
+ $X2=5.52 $Y2=3.33
r265 83 129 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r266 82 83 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r267 80 83 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r268 80 126 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r269 79 82 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r270 79 80 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r271 77 125 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.29 $Y=3.33
+ $X2=1.125 $Y2=3.33
r272 77 79 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=1.29 $Y=3.33
+ $X2=1.68 $Y2=3.33
r273 76 128 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.895 $Y=3.33
+ $X2=3.06 $Y2=3.33
r274 76 82 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=2.895 $Y=3.33
+ $X2=2.64 $Y2=3.33
r275 74 126 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r276 73 74 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r277 71 125 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.96 $Y=3.33
+ $X2=1.125 $Y2=3.33
r278 71 73 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=0.96 $Y=3.33
+ $X2=0.72 $Y2=3.33
r279 69 105 0.73586 $w=4.9e-07 $l=2.64e-06 $layer=MET1_cond $X=9.6 $Y=3.33
+ $X2=12.24 $Y2=3.33
r280 69 102 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=9.6 $Y=3.33
+ $X2=9.36 $Y2=3.33
r281 67 113 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=15.71 $Y=3.33
+ $X2=15.6 $Y2=3.33
r282 67 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=15.71 $Y=3.33
+ $X2=15.875 $Y2=3.33
r283 66 117 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=16.04 $Y=3.33
+ $X2=16.08 $Y2=3.33
r284 66 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=16.04 $Y=3.33
+ $X2=15.875 $Y2=3.33
r285 64 97 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=8.895 $Y=3.33
+ $X2=8.88 $Y2=3.33
r286 64 65 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.895 $Y=3.33
+ $X2=9.06 $Y2=3.33
r287 63 101 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=9.225 $Y=3.33
+ $X2=9.36 $Y2=3.33
r288 63 65 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.225 $Y=3.33
+ $X2=9.06 $Y2=3.33
r289 59 62 16.9374 $w=3.28e-07 $l=4.85e-07 $layer=LI1_cond $X=18.13 $Y=1.98
+ $X2=18.13 $Y2=2.465
r290 57 140 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=18.13 $Y=3.245
+ $X2=18.13 $Y2=3.33
r291 57 62 27.2396 $w=3.28e-07 $l=7.8e-07 $layer=LI1_cond $X=18.13 $Y=3.245
+ $X2=18.13 $Y2=2.465
r292 53 56 27.0649 $w=3.28e-07 $l=7.75e-07 $layer=LI1_cond $X=15.875 $Y=2.125
+ $X2=15.875 $Y2=2.9
r293 51 68 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=15.875 $Y=3.245
+ $X2=15.875 $Y2=3.33
r294 51 56 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=15.875 $Y=3.245
+ $X2=15.875 $Y2=2.9
r295 47 137 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=14.055 $Y=3.245
+ $X2=14.055 $Y2=3.33
r296 47 49 17.5171 $w=2.48e-07 $l=3.8e-07 $layer=LI1_cond $X=14.055 $Y=3.245
+ $X2=14.055 $Y2=2.865
r297 43 134 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=12.66 $Y=3.245
+ $X2=12.66 $Y2=3.33
r298 43 45 11.5244 $w=3.28e-07 $l=3.3e-07 $layer=LI1_cond $X=12.66 $Y=3.245
+ $X2=12.66 $Y2=2.915
r299 39 42 32.4779 $w=3.28e-07 $l=9.3e-07 $layer=LI1_cond $X=9.06 $Y=2.02
+ $X2=9.06 $Y2=2.95
r300 37 65 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.06 $Y=3.245
+ $X2=9.06 $Y2=3.33
r301 37 42 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=9.06 $Y=3.245
+ $X2=9.06 $Y2=2.95
r302 33 131 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.025 $Y=3.245
+ $X2=6.025 $Y2=3.33
r303 33 35 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=6.025 $Y=3.245
+ $X2=6.025 $Y2=2.92
r304 29 128 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.06 $Y=3.245
+ $X2=3.06 $Y2=3.33
r305 29 31 15.3659 $w=3.28e-07 $l=4.4e-07 $layer=LI1_cond $X=3.06 $Y=3.245
+ $X2=3.06 $Y2=2.805
r306 25 125 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.125 $Y=3.245
+ $X2=1.125 $Y2=3.33
r307 25 27 15.3659 $w=3.28e-07 $l=4.4e-07 $layer=LI1_cond $X=1.125 $Y=3.245
+ $X2=1.125 $Y2=2.805
r308 8 62 300 $w=1.7e-07 $l=7.46693e-07 $layer=licon1_PDIFF $count=2 $X=17.875
+ $Y=1.835 $X2=18.13 $Y2=2.465
r309 8 59 600 $w=1.7e-07 $l=3.19374e-07 $layer=licon1_PDIFF $count=1 $X=17.875
+ $Y=1.835 $X2=18.13 $Y2=1.98
r310 7 56 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=15.735
+ $Y=1.785 $X2=15.875 $Y2=2.9
r311 7 53 400 $w=1.7e-07 $l=4.0398e-07 $layer=licon1_PDIFF $count=1 $X=15.735
+ $Y=1.785 $X2=15.875 $Y2=2.125
r312 6 49 600 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=1 $X=13.955
+ $Y=2.59 $X2=14.095 $Y2=2.865
r313 5 45 600 $w=1.7e-07 $l=3.32265e-07 $layer=licon1_PDIFF $count=1 $X=12.44
+ $Y=2.675 $X2=12.66 $Y2=2.915
r314 4 42 600 $w=1.7e-07 $l=1.23116e-06 $layer=licon1_PDIFF $count=1 $X=8.725
+ $Y=1.875 $X2=9.06 $Y2=2.95
r315 4 39 300 $w=1.7e-07 $l=4.00999e-07 $layer=licon1_PDIFF $count=2 $X=8.725
+ $Y=1.875 $X2=9.06 $Y2=2.02
r316 3 35 600 $w=1.7e-07 $l=3.07124e-07 $layer=licon1_PDIFF $count=1 $X=5.885
+ $Y=2.675 $X2=6.025 $Y2=2.92
r317 2 31 600 $w=1.7e-07 $l=4.14126e-07 $layer=licon1_PDIFF $count=1 $X=2.92
+ $Y=2.455 $X2=3.06 $Y2=2.805
r318 1 27 600 $w=1.7e-07 $l=4.14126e-07 $layer=licon1_PDIFF $count=1 $X=0.985
+ $Y=2.455 $X2=1.125 $Y2=2.805
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRBP_LP%A_342_261# 1 2 3 4 14 15 16 17 18 21 25 27
+ 30 31 32 36 37 38 41 43
c132 36 0 1.28847e-19 $X=4.46 $Y=2.7
c133 27 0 1.62564e-19 $X=3.405 $Y=2.23
r134 39 41 12.6769 $w=2.48e-07 $l=2.75e-07 $layer=LI1_cond $X=5.2 $Y=2.025
+ $X2=5.2 $Y2=1.75
r135 37 39 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=5.075 $Y=2.11
+ $X2=5.2 $Y2=2.025
r136 37 38 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=5.075 $Y=2.11
+ $X2=4.545 $Y2=2.11
r137 35 38 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.46 $Y=2.195
+ $X2=4.545 $Y2=2.11
r138 35 36 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=4.46 $Y=2.195
+ $X2=4.46 $Y2=2.7
r139 32 34 26.4014 $w=2.73e-07 $l=6.3e-07 $layer=LI1_cond $X=3.575 $Y=2.837
+ $X2=4.205 $Y2=2.837
r140 31 36 7.32204 $w=2.75e-07 $l=1.74396e-07 $layer=LI1_cond $X=4.375 $Y=2.837
+ $X2=4.46 $Y2=2.7
r141 31 34 7.12419 $w=2.73e-07 $l=1.7e-07 $layer=LI1_cond $X=4.375 $Y=2.837
+ $X2=4.205 $Y2=2.837
r142 30 32 7.32204 $w=2.75e-07 $l=1.74396e-07 $layer=LI1_cond $X=3.49 $Y=2.7
+ $X2=3.575 $Y2=2.837
r143 29 30 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=3.49 $Y=2.315
+ $X2=3.49 $Y2=2.7
r144 28 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.405 $Y=2.23
+ $X2=2.24 $Y2=2.23
r145 27 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.405 $Y=2.23
+ $X2=3.49 $Y2=2.315
r146 27 28 65.2406 $w=1.68e-07 $l=1e-06 $layer=LI1_cond $X=3.405 $Y=2.23
+ $X2=2.405 $Y2=2.23
r147 23 43 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.24 $Y=2.315
+ $X2=2.24 $Y2=2.23
r148 23 25 15.1913 $w=3.28e-07 $l=4.35e-07 $layer=LI1_cond $X=2.24 $Y=2.315
+ $X2=2.24 $Y2=2.75
r149 19 21 7.50834 $w=3.28e-07 $l=2.15e-07 $layer=LI1_cond $X=1.85 $Y=1.235
+ $X2=1.85 $Y2=1.45
r150 17 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.075 $Y=2.23
+ $X2=2.24 $Y2=2.23
r151 17 18 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=2.075 $Y=2.23
+ $X2=1.155 $Y2=2.23
r152 15 19 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.685 $Y=1.15
+ $X2=1.85 $Y2=1.235
r153 15 16 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=1.685 $Y=1.15
+ $X2=1.155 $Y2=1.15
r154 14 18 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.07 $Y=2.145
+ $X2=1.155 $Y2=2.23
r155 13 16 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.07 $Y=1.235
+ $X2=1.155 $Y2=1.15
r156 13 14 59.369 $w=1.68e-07 $l=9.1e-07 $layer=LI1_cond $X=1.07 $Y=1.235
+ $X2=1.07 $Y2=2.145
r157 4 34 600 $w=1.7e-07 $l=3.98905e-07 $layer=licon1_PDIFF $count=1 $X=4.065
+ $Y=2.455 $X2=4.205 $Y2=2.79
r158 3 25 600 $w=1.7e-07 $l=3.58225e-07 $layer=licon1_PDIFF $count=1 $X=2.1
+ $Y=2.455 $X2=2.24 $Y2=2.75
r159 2 41 182 $w=1.7e-07 $l=7.72043e-07 $layer=licon1_NDIFF $count=1 $X=4.985
+ $Y=1.095 $X2=5.24 $Y2=1.75
r160 1 21 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=1.71
+ $Y=1.305 $X2=1.85 $Y2=1.45
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRBP_LP%A_2081_439# 1 2 9 12 14 15
r30 14 15 8.61591 $w=2.68e-07 $l=1.65e-07 $layer=LI1_cond $X=12.15 $Y=2.93
+ $X2=11.985 $Y2=2.93
r31 12 15 82.8556 $w=1.68e-07 $l=1.27e-06 $layer=LI1_cond $X=10.715 $Y=2.98
+ $X2=11.985 $Y2=2.98
r32 7 12 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=10.59 $Y=2.895
+ $X2=10.715 $Y2=2.98
r33 7 9 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=10.59 $Y=2.895
+ $X2=10.59 $Y2=2.465
r34 2 14 600 $w=1.7e-07 $l=3.03974e-07 $layer=licon1_PDIFF $count=1 $X=12.005
+ $Y=2.675 $X2=12.15 $Y2=2.915
r35 1 9 600 $w=1.7e-07 $l=3.34739e-07 $layer=licon1_PDIFF $count=1 $X=10.405
+ $Y=2.195 $X2=10.55 $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRBP_LP%A_2523_397# 1 2 7 12 13 14 18 19
c49 18 0 1.0756e-19 $X=14.525 $Y=2.865
c50 14 0 1.41841e-19 $X=13.4 $Y=1.835
c51 13 0 1.35413e-19 $X=14.52 $Y=1.835
r52 18 19 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=14.525 $Y=2.865
+ $X2=14.525 $Y2=2.7
r53 15 19 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=14.605 $Y=1.92
+ $X2=14.605 $Y2=2.7
r54 13 15 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=14.52 $Y=1.835
+ $X2=14.605 $Y2=1.92
r55 13 14 73.0695 $w=1.68e-07 $l=1.12e-06 $layer=LI1_cond $X=14.52 $Y=1.835
+ $X2=13.4 $Y2=1.835
r56 11 14 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=13.315 $Y=1.92
+ $X2=13.4 $Y2=1.835
r57 11 12 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=13.315 $Y=1.92
+ $X2=13.315 $Y2=2.095
r58 7 12 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=13.23 $Y=2.18
+ $X2=13.315 $Y2=2.095
r59 7 9 30.6631 $w=1.68e-07 $l=4.7e-07 $layer=LI1_cond $X=13.23 $Y=2.18
+ $X2=12.76 $Y2=2.18
r60 2 18 600 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=1 $X=14.385
+ $Y=2.59 $X2=14.525 $Y2=2.865
r61 1 9 600 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_PDIFF $count=1 $X=12.615
+ $Y=1.985 $X2=12.76 $Y2=2.18
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRBP_LP%Q_N 1 2 9 11 15 16 17 23 29
r33 21 29 1.25721 $w=3.83e-07 $l=4.2e-08 $layer=LI1_cond $X=16.637 $Y=0.883
+ $X2=16.637 $Y2=0.925
r34 17 31 7.51133 $w=3.83e-07 $l=1.29e-07 $layer=LI1_cond $X=16.637 $Y=0.946
+ $X2=16.637 $Y2=1.075
r35 17 29 0.628605 $w=3.83e-07 $l=2.1e-08 $layer=LI1_cond $X=16.637 $Y=0.946
+ $X2=16.637 $Y2=0.925
r36 17 21 0.658539 $w=3.83e-07 $l=2.2e-08 $layer=LI1_cond $X=16.637 $Y=0.861
+ $X2=16.637 $Y2=0.883
r37 16 17 9.15968 $w=3.83e-07 $l=3.06e-07 $layer=LI1_cond $X=16.637 $Y=0.555
+ $X2=16.637 $Y2=0.861
r38 16 23 3.7417 $w=3.83e-07 $l=1.25e-07 $layer=LI1_cond $X=16.637 $Y=0.555
+ $X2=16.637 $Y2=0.43
r39 15 31 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=16.745 $Y=1.765
+ $X2=16.745 $Y2=1.075
r40 9 15 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=16.665 $Y=1.93
+ $X2=16.665 $Y2=1.765
r41 9 11 33.8748 $w=3.28e-07 $l=9.7e-07 $layer=LI1_cond $X=16.665 $Y=1.93
+ $X2=16.665 $Y2=2.9
r42 2 11 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=16.525
+ $Y=1.785 $X2=16.665 $Y2=2.9
r43 2 9 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=16.525
+ $Y=1.785 $X2=16.665 $Y2=1.93
r44 1 23 91 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_NDIFF $count=2 $X=16.525
+ $Y=0.235 $X2=16.665 $Y2=0.43
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRBP_LP%Q 1 2 7 8 9 10 11 12 13 22
r15 13 40 4.36531 $w=3.28e-07 $l=1.25e-07 $layer=LI1_cond $X=18.92 $Y=2.775
+ $X2=18.92 $Y2=2.9
r16 12 13 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=18.92 $Y=2.405
+ $X2=18.92 $Y2=2.775
r17 11 12 14.8421 $w=3.28e-07 $l=4.25e-07 $layer=LI1_cond $X=18.92 $Y=1.98
+ $X2=18.92 $Y2=2.405
r18 10 11 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=18.92 $Y=1.665
+ $X2=18.92 $Y2=1.98
r19 9 10 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=18.92 $Y=1.295
+ $X2=18.92 $Y2=1.665
r20 8 9 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=18.92 $Y=0.925
+ $X2=18.92 $Y2=1.295
r21 7 8 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=18.92 $Y=0.555
+ $X2=18.92 $Y2=0.925
r22 7 22 4.36531 $w=3.28e-07 $l=1.25e-07 $layer=LI1_cond $X=18.92 $Y=0.555
+ $X2=18.92 $Y2=0.43
r23 2 40 400 $w=1.7e-07 $l=1.13284e-06 $layer=licon1_PDIFF $count=1 $X=18.78
+ $Y=1.835 $X2=18.92 $Y2=2.9
r24 2 11 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=18.78
+ $Y=1.835 $X2=18.92 $Y2=1.98
r25 1 22 91 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=2 $X=18.78
+ $Y=0.265 $X2=18.92 $Y2=0.43
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRBP_LP%VGND 1 2 3 4 5 6 7 24 28 32 36 40 44 48 53
+ 54 56 57 58 60 65 74 78 90 96 97 100 103 106 109 112
c173 97 0 1.14697e-20 $X=18.96 $Y=0
r174 112 113 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=18 $Y=0 $X2=18
+ $Y2=0
r175 109 110 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=12.24 $Y=0
+ $X2=12.24 $Y2=0
r176 106 107 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.88 $Y=0
+ $X2=8.88 $Y2=0
r177 103 104 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=3.6 $Y=0
+ $X2=3.6 $Y2=0
r178 100 101 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.2 $Y=0
+ $X2=1.2 $Y2=0
r179 97 113 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=18.96 $Y=0 $X2=18
+ $Y2=0
r180 96 97 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=18.96 $Y=0
+ $X2=18.96 $Y2=0
r181 94 112 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=18.295 $Y=0
+ $X2=18.13 $Y2=0
r182 94 96 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=18.295 $Y=0
+ $X2=18.96 $Y2=0
r183 93 113 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=16.08 $Y=0
+ $X2=18 $Y2=0
r184 92 93 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=16.08 $Y=0
+ $X2=16.08 $Y2=0
r185 90 112 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=17.965 $Y=0
+ $X2=18.13 $Y2=0
r186 90 92 122.979 $w=1.68e-07 $l=1.885e-06 $layer=LI1_cond $X=17.965 $Y=0
+ $X2=16.08 $Y2=0
r187 89 93 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=15.6 $Y=0
+ $X2=16.08 $Y2=0
r188 88 89 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=15.6 $Y=0
+ $X2=15.6 $Y2=0
r189 86 89 0.802756 $w=4.9e-07 $l=2.88e-06 $layer=MET1_cond $X=12.72 $Y=0
+ $X2=15.6 $Y2=0
r190 86 110 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.72 $Y=0
+ $X2=12.24 $Y2=0
r191 85 88 187.893 $w=1.68e-07 $l=2.88e-06 $layer=LI1_cond $X=12.72 $Y=0
+ $X2=15.6 $Y2=0
r192 85 86 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=12.72 $Y=0
+ $X2=12.72 $Y2=0
r193 83 109 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.51 $Y=0
+ $X2=12.345 $Y2=0
r194 83 85 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=12.51 $Y=0
+ $X2=12.72 $Y2=0
r195 82 107 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=0
+ $X2=8.88 $Y2=0
r196 81 82 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=9.36 $Y=0
+ $X2=9.36 $Y2=0
r197 79 106 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.195 $Y=0
+ $X2=9.03 $Y2=0
r198 79 81 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=9.195 $Y=0
+ $X2=9.36 $Y2=0
r199 78 109 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.18 $Y=0
+ $X2=12.345 $Y2=0
r200 78 81 183.979 $w=1.68e-07 $l=2.82e-06 $layer=LI1_cond $X=12.18 $Y=0
+ $X2=9.36 $Y2=0
r201 77 107 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=7.44 $Y=0
+ $X2=8.88 $Y2=0
r202 76 77 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r203 74 106 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.865 $Y=0
+ $X2=9.03 $Y2=0
r204 74 76 92.9679 $w=1.68e-07 $l=1.425e-06 $layer=LI1_cond $X=8.865 $Y=0
+ $X2=7.44 $Y2=0
r205 73 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=7.44
+ $Y2=0
r206 73 104 0.936549 $w=4.9e-07 $l=3.36e-06 $layer=MET1_cond $X=6.96 $Y=0
+ $X2=3.6 $Y2=0
r207 72 73 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=6.96 $Y=0
+ $X2=6.96 $Y2=0
r208 70 103 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.65 $Y=0 $X2=3.565
+ $Y2=0
r209 70 72 215.947 $w=1.68e-07 $l=3.31e-06 $layer=LI1_cond $X=3.65 $Y=0 $X2=6.96
+ $Y2=0
r210 69 104 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r211 69 101 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=3.12 $Y=0
+ $X2=1.2 $Y2=0
r212 68 69 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=0
+ $X2=3.12 $Y2=0
r213 66 100 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.275 $Y=0
+ $X2=1.11 $Y2=0
r214 66 68 120.369 $w=1.68e-07 $l=1.845e-06 $layer=LI1_cond $X=1.275 $Y=0
+ $X2=3.12 $Y2=0
r215 65 103 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.48 $Y=0 $X2=3.565
+ $Y2=0
r216 65 68 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=3.48 $Y=0 $X2=3.12
+ $Y2=0
r217 63 101 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r218 62 63 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r219 60 100 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.945 $Y=0
+ $X2=1.11 $Y2=0
r220 60 62 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=0.945 $Y=0
+ $X2=0.72 $Y2=0
r221 58 110 0.73586 $w=4.9e-07 $l=2.64e-06 $layer=MET1_cond $X=9.6 $Y=0
+ $X2=12.24 $Y2=0
r222 58 82 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=9.6 $Y=0 $X2=9.36
+ $Y2=0
r223 56 88 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=15.71 $Y=0 $X2=15.6
+ $Y2=0
r224 56 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=15.71 $Y=0
+ $X2=15.875 $Y2=0
r225 55 92 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=16.04 $Y=0 $X2=16.08
+ $Y2=0
r226 55 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=16.04 $Y=0
+ $X2=15.875 $Y2=0
r227 53 72 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=6.995 $Y=0 $X2=6.96
+ $Y2=0
r228 53 54 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.995 $Y=0 $X2=7.12
+ $Y2=0
r229 52 76 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=7.245 $Y=0
+ $X2=7.44 $Y2=0
r230 52 54 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.245 $Y=0 $X2=7.12
+ $Y2=0
r231 48 50 19.2074 $w=3.28e-07 $l=5.5e-07 $layer=LI1_cond $X=18.13 $Y=0.41
+ $X2=18.13 $Y2=0.96
r232 46 112 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=18.13 $Y=0.085
+ $X2=18.13 $Y2=0
r233 46 48 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=18.13 $Y=0.085
+ $X2=18.13 $Y2=0.41
r234 42 57 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=15.875 $Y=0.085
+ $X2=15.875 $Y2=0
r235 42 44 13.0959 $w=3.28e-07 $l=3.75e-07 $layer=LI1_cond $X=15.875 $Y=0.085
+ $X2=15.875 $Y2=0.46
r236 38 109 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=12.345 $Y=0.085
+ $X2=12.345 $Y2=0
r237 38 40 21.652 $w=3.28e-07 $l=6.2e-07 $layer=LI1_cond $X=12.345 $Y=0.085
+ $X2=12.345 $Y2=0.705
r238 34 106 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.03 $Y=0.085
+ $X2=9.03 $Y2=0
r239 34 36 7.50834 $w=3.28e-07 $l=2.15e-07 $layer=LI1_cond $X=9.03 $Y=0.085
+ $X2=9.03 $Y2=0.3
r240 30 54 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.12 $Y=0.085
+ $X2=7.12 $Y2=0
r241 30 32 13.1378 $w=2.48e-07 $l=2.85e-07 $layer=LI1_cond $X=7.12 $Y=0.085
+ $X2=7.12 $Y2=0.37
r242 26 103 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.565 $Y=0.085
+ $X2=3.565 $Y2=0
r243 26 28 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=3.565 $Y=0.085
+ $X2=3.565 $Y2=0.38
r244 22 100 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.11 $Y=0.085
+ $X2=1.11 $Y2=0
r245 22 24 11.5244 $w=3.28e-07 $l=3.3e-07 $layer=LI1_cond $X=1.11 $Y=0.085
+ $X2=1.11 $Y2=0.415
r246 7 50 182 $w=1.7e-07 $l=3.81772e-07 $layer=licon1_NDIFF $count=1 $X=17.875
+ $Y=0.685 $X2=18.13 $Y2=0.96
r247 7 48 182 $w=1.7e-07 $l=3.81772e-07 $layer=licon1_NDIFF $count=1 $X=17.875
+ $Y=0.685 $X2=18.13 $Y2=0.41
r248 6 44 182 $w=1.7e-07 $l=2.86575e-07 $layer=licon1_NDIFF $count=1 $X=15.735
+ $Y=0.235 $X2=15.875 $Y2=0.46
r249 5 40 182 $w=1.7e-07 $l=2.55e-07 $layer=licon1_NDIFF $count=1 $X=12.09
+ $Y=0.705 $X2=12.345 $Y2=0.705
r250 4 36 182 $w=1.7e-07 $l=3.968e-07 $layer=licon1_NDIFF $count=1 $X=8.695
+ $Y=0.435 $X2=9.03 $Y2=0.3
r251 3 32 182 $w=1.7e-07 $l=3.49857e-07 $layer=licon1_NDIFF $count=1 $X=6.905
+ $Y=0.595 $X2=7.16 $Y2=0.37
r252 2 28 182 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=1 $X=3.44
+ $Y=0.215 $X2=3.565 $Y2=0.38
r253 1 24 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=0.97
+ $Y=0.235 $X2=1.11 $Y2=0.415
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRBP_LP%noxref_37 1 2 9 11 12 15
r34 13 15 9.91101 $w=2.48e-07 $l=2.15e-07 $layer=LI1_cond $X=3.03 $Y=1.795
+ $X2=3.03 $Y2=1.58
r35 11 13 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.905 $Y=1.88
+ $X2=3.03 $Y2=1.795
r36 11 12 91.3369 $w=1.68e-07 $l=1.4e-06 $layer=LI1_cond $X=2.905 $Y=1.88
+ $X2=1.505 $Y2=1.88
r37 7 12 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.42 $Y=1.795
+ $X2=1.505 $Y2=1.88
r38 7 9 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=1.42 $Y=1.795
+ $X2=1.42 $Y2=1.58
r39 2 15 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=2.93
+ $Y=1.305 $X2=3.07 $Y2=1.58
r40 1 9 182 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=1 $X=1.275
+ $Y=1.305 $X2=1.42 $Y2=1.58
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRBP_LP%noxref_39 1 2 9 11 12 14 15 16 18
c53 11 0 4.85838e-20 $X=3.415 $Y=1.15
r54 15 18 11.6281 $w=3.2e-07 $l=3.88555e-07 $layer=LI1_cond $X=3.83 $Y=0.81
+ $X2=4.02 $Y2=0.505
r55 15 16 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=3.83 $Y=0.81
+ $X2=3.585 $Y2=0.81
r56 13 16 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.5 $Y=0.895
+ $X2=3.585 $Y2=0.81
r57 13 14 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=3.5 $Y=0.895 $X2=3.5
+ $Y2=1.065
r58 11 14 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.415 $Y=1.15
+ $X2=3.5 $Y2=1.065
r59 11 12 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.415 $Y=1.15
+ $X2=2.725 $Y2=1.15
r60 7 12 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.6 $Y=1.235
+ $X2=2.725 $Y2=1.15
r61 7 9 9.91101 $w=2.48e-07 $l=2.15e-07 $layer=LI1_cond $X=2.6 $Y=1.235 $X2=2.6
+ $Y2=1.45
r62 2 18 182 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=1 $X=3.915
+ $Y=0.33 $X2=4.055 $Y2=0.505
r63 1 9 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=2.5
+ $Y=1.305 $X2=2.64 $Y2=1.45
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRBP_LP%A_824_219# 1 2 7 11 13 16
c30 11 0 1.28843e-19 $X=6.225 $Y=0.8
r31 16 18 6.53051 $w=2.98e-07 $l=1.7e-07 $layer=LI1_cond $X=5.62 $Y=0.8 $X2=5.62
+ $Y2=0.97
r32 13 15 17.036 $w=2.22e-07 $l=3.1e-07 $layer=LI1_cond $X=4.225 $Y=0.97
+ $X2=4.225 $Y2=1.28
r33 9 16 4.061 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=5.77 $Y=0.8 $X2=5.62
+ $Y2=0.8
r34 9 11 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=5.77 $Y=0.8
+ $X2=6.225 $Y2=0.8
r35 8 13 2.3025 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.35 $Y=0.97 $X2=4.225
+ $Y2=0.97
r36 7 18 4.061 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=5.47 $Y=0.97 $X2=5.62
+ $Y2=0.97
r37 7 8 73.0695 $w=1.68e-07 $l=1.12e-06 $layer=LI1_cond $X=5.47 $Y=0.97 $X2=4.35
+ $Y2=0.97
r38 2 11 182 $w=1.7e-07 $l=2.67862e-07 $layer=licon1_NDIFF $count=1 $X=6.08
+ $Y=0.595 $X2=6.225 $Y2=0.8
r39 1 15 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=4.12
+ $Y=1.095 $X2=4.265 $Y2=1.28
.ends

