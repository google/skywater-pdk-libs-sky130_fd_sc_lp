* NGSPICE file created from sky130_fd_sc_lp__o311ai_2.ext - technology: sky130A

.subckt sky130_fd_sc_lp__o311ai_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
M1000 a_35_47# B1 a_710_47# VNB nshort w=840000u l=150000u
+  ad=1.1844e+12p pd=1.122e+07u as=4.704e+11p ps=4.48e+06u
M1001 VPWR C1 Y VPB phighvt w=1.26e+06u l=150000u
+  ad=1.5372e+12p pd=1e+07u as=1.3734e+12p ps=1.226e+07u
M1002 a_35_47# A3 VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=9.912e+11p ps=7.4e+06u
M1003 a_290_367# A2 a_35_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=7.056e+11p pd=6.16e+06u as=1.0206e+12p ps=9.18e+06u
M1004 VPWR A1 a_35_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_290_367# A3 Y VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND A2 a_35_47# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 Y B1 VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_710_47# C1 Y VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=4.452e+11p ps=4.42e+06u
M1009 a_710_47# B1 a_35_47# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 Y C1 VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 Y C1 a_710_47# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_35_367# A1 VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VPWR B1 Y VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VGND A3 a_35_47# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_35_367# A2 a_290_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 Y A3 a_290_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_35_47# A2 VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VGND A1 a_35_47# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_35_47# A1 VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

