* File: sky130_fd_sc_lp__nand3b_2.pxi.spice
* Created: Wed Sep  2 10:04:52 2020
* 
x_PM_SKY130_FD_SC_LP__NAND3B_2%A_N N_A_N_M1009_g N_A_N_M1004_g A_N N_A_N_c_79_n
+ PM_SKY130_FD_SC_LP__NAND3B_2%A_N
x_PM_SKY130_FD_SC_LP__NAND3B_2%C N_C_M1005_g N_C_M1001_g N_C_M1007_g N_C_M1006_g
+ N_C_c_132_p N_C_c_165_p N_C_c_110_n N_C_c_111_n N_C_c_118_n C N_C_c_112_n
+ N_C_c_113_n PM_SKY130_FD_SC_LP__NAND3B_2%C
x_PM_SKY130_FD_SC_LP__NAND3B_2%B N_B_M1008_g N_B_M1012_g N_B_M1010_g N_B_M1013_g
+ N_B_c_207_n N_B_c_208_n N_B_c_215_n B B N_B_c_209_n N_B_c_210_n N_B_c_218_n
+ PM_SKY130_FD_SC_LP__NAND3B_2%B
x_PM_SKY130_FD_SC_LP__NAND3B_2%A_55_155# N_A_55_155#_M1009_s N_A_55_155#_M1004_s
+ N_A_55_155#_c_298_n N_A_55_155#_M1000_g N_A_55_155#_M1002_g
+ N_A_55_155#_M1011_g N_A_55_155#_c_301_n N_A_55_155#_M1003_g
+ N_A_55_155#_c_302_n N_A_55_155#_c_315_n N_A_55_155#_c_303_n
+ N_A_55_155#_c_304_n N_A_55_155#_c_345_n N_A_55_155#_c_305_n
+ N_A_55_155#_c_310_n N_A_55_155#_c_306_n PM_SKY130_FD_SC_LP__NAND3B_2%A_55_155#
x_PM_SKY130_FD_SC_LP__NAND3B_2%VPWR N_VPWR_M1004_d N_VPWR_M1012_s N_VPWR_M1011_s
+ N_VPWR_M1006_s N_VPWR_c_396_n N_VPWR_c_397_n N_VPWR_c_398_n N_VPWR_c_399_n
+ N_VPWR_c_400_n N_VPWR_c_401_n N_VPWR_c_402_n N_VPWR_c_403_n N_VPWR_c_404_n
+ N_VPWR_c_405_n N_VPWR_c_406_n N_VPWR_c_407_n VPWR N_VPWR_c_408_n
+ N_VPWR_c_395_n PM_SKY130_FD_SC_LP__NAND3B_2%VPWR
x_PM_SKY130_FD_SC_LP__NAND3B_2%Y N_Y_M1000_d N_Y_M1001_d N_Y_M1002_d N_Y_M1013_d
+ N_Y_c_476_n N_Y_c_467_n N_Y_c_480_n N_Y_c_481_n N_Y_c_483_n N_Y_c_501_n
+ N_Y_c_486_n N_Y_c_487_n Y Y Y Y N_Y_c_470_n Y PM_SKY130_FD_SC_LP__NAND3B_2%Y
x_PM_SKY130_FD_SC_LP__NAND3B_2%VGND N_VGND_M1009_d N_VGND_M1007_s N_VGND_c_556_n
+ N_VGND_c_557_n N_VGND_c_558_n N_VGND_c_559_n N_VGND_c_560_n N_VGND_c_561_n
+ VGND N_VGND_c_562_n N_VGND_c_563_n PM_SKY130_FD_SC_LP__NAND3B_2%VGND
x_PM_SKY130_FD_SC_LP__NAND3B_2%A_246_71# N_A_246_71#_M1005_d N_A_246_71#_M1010_d
+ N_A_246_71#_c_599_n N_A_246_71#_c_595_n N_A_246_71#_c_596_n
+ N_A_246_71#_c_612_n PM_SKY130_FD_SC_LP__NAND3B_2%A_246_71#
x_PM_SKY130_FD_SC_LP__NAND3B_2%A_332_71# N_A_332_71#_M1008_s N_A_332_71#_M1003_s
+ N_A_332_71#_c_625_n N_A_332_71#_c_622_n N_A_332_71#_c_630_n
+ PM_SKY130_FD_SC_LP__NAND3B_2%A_332_71#
cc_1 VNB N_A_N_M1009_g 0.0256745f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=0.985
cc_2 VNB A_N 0.00312827f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_3 VNB N_A_N_c_79_n 0.0258931f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.51
cc_4 VNB N_C_M1005_g 0.0217151f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=0.985
cc_5 VNB N_C_M1007_g 0.0222313f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.51
cc_6 VNB N_C_c_110_n 9.29659e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_C_c_111_n 0.0279932f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_C_c_112_n 0.0237517f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_C_c_113_n 0.00285359f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_B_M1008_g 0.019589f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=0.985
cc_11 VNB N_B_M1010_g 0.0192555f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.51
cc_12 VNB N_B_c_207_n 5.52202e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_B_c_208_n 0.0260562f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_B_c_209_n 0.0223664f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_B_c_210_n 0.0042783f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_55_155#_c_298_n 0.0180704f $X=-0.19 $Y=-0.245 $X2=0.615 $Y2=2.045
cc_17 VNB N_A_55_155#_M1002_g 0.00102808f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.51
cc_18 VNB N_A_55_155#_M1011_g 8.23994e-19 $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.547
cc_19 VNB N_A_55_155#_c_301_n 0.0180077f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.547
cc_20 VNB N_A_55_155#_c_302_n 0.0233776f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_55_155#_c_303_n 0.00149575f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_55_155#_c_304_n 0.00251167f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_55_155#_c_305_n 0.0207538f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_55_155#_c_306_n 0.0486854f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_VPWR_c_395_n 0.183584f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_Y_c_467_n 0.018807f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB Y 0.0258314f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_556_n 0.0218761f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_29 VNB N_VGND_c_557_n 0.0281161f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.51
cc_30 VNB N_VGND_c_558_n 0.0268053f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.547
cc_31 VNB N_VGND_c_559_n 0.00604418f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_560_n 0.0594397f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_561_n 0.00604418f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_562_n 0.0124854f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_563_n 0.264259f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_246_71#_c_595_n 0.0111775f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.51
cc_37 VNB N_A_246_71#_c_596_n 0.00245371f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=1.51
cc_38 VPB N_A_N_M1004_g 0.0294696f $X=-0.19 $Y=1.655 $X2=0.615 $Y2=2.045
cc_39 VPB A_N 0.00493805f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_40 VPB N_A_N_c_79_n 0.00631029f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=1.51
cc_41 VPB N_C_M1001_g 0.0213326f $X=-0.19 $Y=1.655 $X2=0.615 $Y2=2.045
cc_42 VPB N_C_M1006_g 0.0233956f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=1.675
cc_43 VPB N_C_c_110_n 0.00147968f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_44 VPB N_C_c_111_n 0.00846246f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_45 VPB N_C_c_118_n 8.2099e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_46 VPB N_C_c_112_n 0.00613587f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_47 VPB N_C_c_113_n 0.00463383f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_48 VPB N_B_M1012_g 0.0193613f $X=-0.19 $Y=1.655 $X2=0.615 $Y2=2.045
cc_49 VPB N_B_M1013_g 0.0188161f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=1.675
cc_50 VPB N_B_c_207_n 6.99739e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_51 VPB N_B_c_208_n 0.00623107f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_52 VPB N_B_c_215_n 6.3656e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_53 VPB N_B_c_209_n 0.00633055f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_54 VPB N_B_c_210_n 0.00217143f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_55 VPB N_B_c_218_n 0.0067513f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_56 VPB N_A_55_155#_M1002_g 0.0206828f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=1.51
cc_57 VPB N_A_55_155#_M1011_g 0.019666f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=1.547
cc_58 VPB N_A_55_155#_c_302_n 0.0135411f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_59 VPB N_A_55_155#_c_310_n 0.0205254f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_60 VPB N_VPWR_c_396_n 0.0343357f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=1.675
cc_61 VPB N_VPWR_c_397_n 0.00561774f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_62 VPB N_VPWR_c_398_n 0.0049444f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_63 VPB N_VPWR_c_399_n 0.017587f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_64 VPB N_VPWR_c_400_n 0.0255325f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_401_n 0.00545601f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_402_n 0.018723f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_67 VPB N_VPWR_c_403_n 0.00632057f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_404_n 0.0169969f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_69 VPB N_VPWR_c_405_n 0.0061216f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_70 VPB N_VPWR_c_406_n 0.0167176f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_71 VPB N_VPWR_c_407_n 0.00497102f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_72 VPB N_VPWR_c_408_n 0.0116219f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_73 VPB N_VPWR_c_395_n 0.0729343f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_74 VPB Y 0.0408781f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_75 VPB N_Y_c_470_n 0.0125371f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_76 N_A_N_M1009_g N_C_M1005_g 0.0179359f $X=0.615 $Y=0.985 $X2=0 $Y2=0
cc_77 N_A_N_M1004_g N_C_M1001_g 0.0120543f $X=0.615 $Y=2.045 $X2=0 $Y2=0
cc_78 A_N N_C_M1001_g 2.30766e-19 $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_79 N_A_N_M1004_g N_C_c_118_n 7.90859e-19 $X=0.615 $Y=2.045 $X2=0 $Y2=0
cc_80 A_N N_C_c_112_n 0.00232237f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_81 N_A_N_c_79_n N_C_c_112_n 0.0181789f $X=0.525 $Y=1.51 $X2=0 $Y2=0
cc_82 N_A_N_M1004_g N_C_c_113_n 2.07318e-19 $X=0.615 $Y=2.045 $X2=0 $Y2=0
cc_83 A_N N_C_c_113_n 0.0332136f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_84 N_A_N_c_79_n N_C_c_113_n 2.82114e-19 $X=0.525 $Y=1.51 $X2=0 $Y2=0
cc_85 N_A_N_M1009_g N_A_55_155#_c_302_n 0.00500856f $X=0.615 $Y=0.985 $X2=0
+ $Y2=0
cc_86 N_A_N_M1004_g N_A_55_155#_c_302_n 0.00439795f $X=0.615 $Y=2.045 $X2=0
+ $Y2=0
cc_87 A_N N_A_55_155#_c_302_n 0.0311998f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_88 N_A_N_c_79_n N_A_55_155#_c_302_n 0.00804858f $X=0.525 $Y=1.51 $X2=0 $Y2=0
cc_89 N_A_N_M1009_g N_A_55_155#_c_315_n 0.0112219f $X=0.615 $Y=0.985 $X2=0 $Y2=0
cc_90 N_A_N_M1009_g N_A_55_155#_c_305_n 0.00489447f $X=0.615 $Y=0.985 $X2=0
+ $Y2=0
cc_91 A_N N_A_55_155#_c_305_n 0.0263481f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_92 N_A_N_c_79_n N_A_55_155#_c_305_n 0.00521122f $X=0.525 $Y=1.51 $X2=0 $Y2=0
cc_93 N_A_N_M1004_g N_A_55_155#_c_310_n 0.00419903f $X=0.615 $Y=2.045 $X2=0
+ $Y2=0
cc_94 A_N N_A_55_155#_c_310_n 0.00864397f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_95 N_A_N_c_79_n N_A_55_155#_c_310_n 0.00310292f $X=0.525 $Y=1.51 $X2=0 $Y2=0
cc_96 N_A_N_M1004_g N_VPWR_c_396_n 0.00366166f $X=0.615 $Y=2.045 $X2=0 $Y2=0
cc_97 A_N N_VPWR_c_396_n 0.00777882f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_98 N_A_N_M1009_g N_VGND_c_556_n 0.00504443f $X=0.615 $Y=0.985 $X2=0 $Y2=0
cc_99 N_A_N_M1009_g N_VGND_c_558_n 0.00344367f $X=0.615 $Y=0.985 $X2=0 $Y2=0
cc_100 N_A_N_M1009_g N_VGND_c_563_n 0.00429888f $X=0.615 $Y=0.985 $X2=0 $Y2=0
cc_101 N_C_M1005_g N_B_M1008_g 0.0330976f $X=1.155 $Y=0.775 $X2=0 $Y2=0
cc_102 N_C_M1001_g N_B_M1012_g 0.0366395f $X=1.175 $Y=2.465 $X2=0 $Y2=0
cc_103 N_C_c_132_p N_B_M1012_g 0.01114f $X=3.54 $Y=2.16 $X2=0 $Y2=0
cc_104 N_C_c_118_n N_B_M1012_g 0.00398845f $X=1.275 $Y=2.075 $X2=0 $Y2=0
cc_105 N_C_c_113_n N_B_M1012_g 4.03537e-19 $X=1.275 $Y=1.547 $X2=0 $Y2=0
cc_106 N_C_M1007_g N_B_M1010_g 0.0287267f $X=3.615 $Y=0.775 $X2=0 $Y2=0
cc_107 N_C_M1006_g N_B_M1013_g 0.0368661f $X=3.615 $Y=2.465 $X2=0 $Y2=0
cc_108 N_C_c_132_p N_B_M1013_g 0.0110517f $X=3.54 $Y=2.16 $X2=0 $Y2=0
cc_109 N_C_c_110_n N_B_M1013_g 0.00133529f $X=3.705 $Y=1.51 $X2=0 $Y2=0
cc_110 N_C_c_112_n N_B_c_207_n 3.60495e-19 $X=1.085 $Y=1.51 $X2=0 $Y2=0
cc_111 N_C_c_113_n N_B_c_207_n 0.0298886f $X=1.275 $Y=1.547 $X2=0 $Y2=0
cc_112 N_C_c_132_p N_B_c_208_n 0.00143953f $X=3.54 $Y=2.16 $X2=0 $Y2=0
cc_113 N_C_c_112_n N_B_c_208_n 0.0204566f $X=1.085 $Y=1.51 $X2=0 $Y2=0
cc_114 N_C_c_113_n N_B_c_208_n 0.00215561f $X=1.275 $Y=1.547 $X2=0 $Y2=0
cc_115 N_C_c_132_p N_B_c_215_n 0.0111674f $X=3.54 $Y=2.16 $X2=0 $Y2=0
cc_116 N_C_c_118_n N_B_c_215_n 0.0122948f $X=1.275 $Y=2.075 $X2=0 $Y2=0
cc_117 N_C_c_113_n N_B_c_215_n 0.00118838f $X=1.275 $Y=1.547 $X2=0 $Y2=0
cc_118 N_C_c_132_p N_B_c_209_n 5.85248e-19 $X=3.54 $Y=2.16 $X2=0 $Y2=0
cc_119 N_C_c_110_n N_B_c_209_n 4.17019e-19 $X=3.705 $Y=1.51 $X2=0 $Y2=0
cc_120 N_C_c_111_n N_B_c_209_n 0.0207694f $X=3.705 $Y=1.51 $X2=0 $Y2=0
cc_121 N_C_M1006_g N_B_c_210_n 0.00149003f $X=3.615 $Y=2.465 $X2=0 $Y2=0
cc_122 N_C_c_110_n N_B_c_210_n 0.0377457f $X=3.705 $Y=1.51 $X2=0 $Y2=0
cc_123 N_C_c_111_n N_B_c_210_n 0.00114351f $X=3.705 $Y=1.51 $X2=0 $Y2=0
cc_124 N_C_c_132_p N_B_c_218_n 0.0929049f $X=3.54 $Y=2.16 $X2=0 $Y2=0
cc_125 N_C_c_132_p N_A_55_155#_M1002_g 0.01122f $X=3.54 $Y=2.16 $X2=0 $Y2=0
cc_126 N_C_c_132_p N_A_55_155#_M1011_g 0.0110982f $X=3.54 $Y=2.16 $X2=0 $Y2=0
cc_127 N_C_M1005_g N_A_55_155#_c_315_n 0.0148133f $X=1.155 $Y=0.775 $X2=0 $Y2=0
cc_128 N_C_c_112_n N_A_55_155#_c_315_n 0.0046739f $X=1.085 $Y=1.51 $X2=0 $Y2=0
cc_129 N_C_c_113_n N_A_55_155#_c_315_n 0.022973f $X=1.275 $Y=1.547 $X2=0 $Y2=0
cc_130 N_C_M1005_g N_A_55_155#_c_305_n 6.28513e-19 $X=1.155 $Y=0.775 $X2=0 $Y2=0
cc_131 N_C_c_132_p N_VPWR_M1012_s 0.00752485f $X=3.54 $Y=2.16 $X2=0 $Y2=0
cc_132 N_C_c_132_p N_VPWR_M1011_s 0.00666493f $X=3.54 $Y=2.16 $X2=0 $Y2=0
cc_133 N_C_c_132_p N_VPWR_M1006_s 0.00235182f $X=3.54 $Y=2.16 $X2=0 $Y2=0
cc_134 N_C_c_110_n N_VPWR_M1006_s 0.00257726f $X=3.705 $Y=1.51 $X2=0 $Y2=0
cc_135 N_C_M1001_g N_VPWR_c_396_n 0.0146561f $X=1.175 $Y=2.465 $X2=0 $Y2=0
cc_136 N_C_c_165_p N_VPWR_c_396_n 0.0138603f $X=1.36 $Y=2.16 $X2=0 $Y2=0
cc_137 N_C_c_118_n N_VPWR_c_396_n 0.0113004f $X=1.275 $Y=2.075 $X2=0 $Y2=0
cc_138 N_C_c_112_n N_VPWR_c_396_n 0.00340427f $X=1.085 $Y=1.51 $X2=0 $Y2=0
cc_139 N_C_c_113_n N_VPWR_c_396_n 0.00167209f $X=1.275 $Y=1.547 $X2=0 $Y2=0
cc_140 N_C_M1006_g N_VPWR_c_399_n 0.00327088f $X=3.615 $Y=2.465 $X2=0 $Y2=0
cc_141 N_C_M1001_g N_VPWR_c_402_n 0.0054895f $X=1.175 $Y=2.465 $X2=0 $Y2=0
cc_142 N_C_M1006_g N_VPWR_c_406_n 0.00428252f $X=3.615 $Y=2.465 $X2=0 $Y2=0
cc_143 N_C_M1001_g N_VPWR_c_395_n 0.0111864f $X=1.175 $Y=2.465 $X2=0 $Y2=0
cc_144 N_C_M1006_g N_VPWR_c_395_n 0.00696163f $X=3.615 $Y=2.465 $X2=0 $Y2=0
cc_145 N_C_c_132_p N_Y_M1001_d 0.00515101f $X=3.54 $Y=2.16 $X2=0 $Y2=0
cc_146 N_C_c_165_p N_Y_M1001_d 5.69898e-19 $X=1.36 $Y=2.16 $X2=0 $Y2=0
cc_147 N_C_c_118_n N_Y_M1001_d 0.00254467f $X=1.275 $Y=2.075 $X2=0 $Y2=0
cc_148 N_C_c_132_p N_Y_M1002_d 0.00339614f $X=3.54 $Y=2.16 $X2=0 $Y2=0
cc_149 N_C_c_132_p N_Y_M1013_d 0.00772134f $X=3.54 $Y=2.16 $X2=0 $Y2=0
cc_150 N_C_c_132_p N_Y_c_476_n 0.0405558f $X=3.54 $Y=2.16 $X2=0 $Y2=0
cc_151 N_C_M1007_g N_Y_c_467_n 0.0163373f $X=3.615 $Y=0.775 $X2=0 $Y2=0
cc_152 N_C_c_110_n N_Y_c_467_n 0.0170524f $X=3.705 $Y=1.51 $X2=0 $Y2=0
cc_153 N_C_c_111_n N_Y_c_467_n 0.0036164f $X=3.705 $Y=1.51 $X2=0 $Y2=0
cc_154 N_C_c_132_p N_Y_c_480_n 0.0383768f $X=3.54 $Y=2.16 $X2=0 $Y2=0
cc_155 N_C_M1006_g N_Y_c_481_n 0.0107018f $X=3.615 $Y=2.465 $X2=0 $Y2=0
cc_156 N_C_c_132_p N_Y_c_481_n 0.0129414f $X=3.54 $Y=2.16 $X2=0 $Y2=0
cc_157 N_C_M1001_g N_Y_c_483_n 0.00886145f $X=1.175 $Y=2.465 $X2=0 $Y2=0
cc_158 N_C_c_132_p N_Y_c_483_n 0.0109584f $X=3.54 $Y=2.16 $X2=0 $Y2=0
cc_159 N_C_c_165_p N_Y_c_483_n 0.00663472f $X=1.36 $Y=2.16 $X2=0 $Y2=0
cc_160 N_C_c_132_p N_Y_c_486_n 0.0171883f $X=3.54 $Y=2.16 $X2=0 $Y2=0
cc_161 N_C_M1006_g N_Y_c_487_n 0.0123522f $X=3.615 $Y=2.465 $X2=0 $Y2=0
cc_162 N_C_c_132_p N_Y_c_487_n 0.0173577f $X=3.54 $Y=2.16 $X2=0 $Y2=0
cc_163 N_C_M1007_g Y 0.00550655f $X=3.615 $Y=0.775 $X2=0 $Y2=0
cc_164 N_C_M1006_g Y 0.0087978f $X=3.615 $Y=2.465 $X2=0 $Y2=0
cc_165 N_C_c_132_p Y 0.0145426f $X=3.54 $Y=2.16 $X2=0 $Y2=0
cc_166 N_C_c_110_n Y 0.0570043f $X=3.705 $Y=1.51 $X2=0 $Y2=0
cc_167 N_C_c_111_n Y 0.00823336f $X=3.705 $Y=1.51 $X2=0 $Y2=0
cc_168 N_C_M1005_g N_VGND_c_556_n 0.0130612f $X=1.155 $Y=0.775 $X2=0 $Y2=0
cc_169 N_C_M1007_g N_VGND_c_557_n 0.0133941f $X=3.615 $Y=0.775 $X2=0 $Y2=0
cc_170 N_C_M1005_g N_VGND_c_560_n 0.00393414f $X=1.155 $Y=0.775 $X2=0 $Y2=0
cc_171 N_C_M1007_g N_VGND_c_560_n 0.00393414f $X=3.615 $Y=0.775 $X2=0 $Y2=0
cc_172 N_C_M1005_g N_VGND_c_563_n 0.00768358f $X=1.155 $Y=0.775 $X2=0 $Y2=0
cc_173 N_C_M1007_g N_VGND_c_563_n 0.00769799f $X=3.615 $Y=0.775 $X2=0 $Y2=0
cc_174 N_C_M1007_g N_A_246_71#_c_595_n 0.00121271f $X=3.615 $Y=0.775 $X2=0 $Y2=0
cc_175 N_C_M1005_g N_A_246_71#_c_596_n 0.00112235f $X=1.155 $Y=0.775 $X2=0 $Y2=0
cc_176 N_B_M1008_g N_A_55_155#_c_298_n 0.0299342f $X=1.585 $Y=0.775 $X2=0 $Y2=0
cc_177 N_B_M1012_g N_A_55_155#_M1002_g 0.0390416f $X=1.605 $Y=2.465 $X2=0 $Y2=0
cc_178 N_B_c_207_n N_A_55_155#_M1002_g 0.00122827f $X=1.625 $Y=1.51 $X2=0 $Y2=0
cc_179 N_B_c_208_n N_A_55_155#_M1002_g 0.00161716f $X=1.625 $Y=1.51 $X2=0 $Y2=0
cc_180 N_B_c_210_n N_A_55_155#_M1002_g 0.00250435f $X=3.165 $Y=1.51 $X2=0 $Y2=0
cc_181 N_B_c_218_n N_A_55_155#_M1002_g 0.011221f $X=2.52 $Y=1.625 $X2=0 $Y2=0
cc_182 N_B_M1013_g N_A_55_155#_M1011_g 0.0428741f $X=3.185 $Y=2.465 $X2=0 $Y2=0
cc_183 N_B_c_210_n N_A_55_155#_M1011_g 0.012396f $X=3.165 $Y=1.51 $X2=0 $Y2=0
cc_184 N_B_M1010_g N_A_55_155#_c_301_n 0.0346022f $X=3.145 $Y=0.775 $X2=0 $Y2=0
cc_185 N_B_M1008_g N_A_55_155#_c_315_n 0.0129959f $X=1.585 $Y=0.775 $X2=0 $Y2=0
cc_186 N_B_c_207_n N_A_55_155#_c_315_n 0.0121543f $X=1.625 $Y=1.51 $X2=0 $Y2=0
cc_187 N_B_c_208_n N_A_55_155#_c_315_n 0.00217672f $X=1.625 $Y=1.51 $X2=0 $Y2=0
cc_188 N_B_c_218_n N_A_55_155#_c_315_n 0.00528874f $X=2.52 $Y=1.625 $X2=0 $Y2=0
cc_189 N_B_M1008_g N_A_55_155#_c_303_n 0.00335936f $X=1.585 $Y=0.775 $X2=0 $Y2=0
cc_190 N_B_c_207_n N_A_55_155#_c_304_n 0.0172978f $X=1.625 $Y=1.51 $X2=0 $Y2=0
cc_191 N_B_c_208_n N_A_55_155#_c_304_n 0.00154753f $X=1.625 $Y=1.51 $X2=0 $Y2=0
cc_192 N_B_c_218_n N_A_55_155#_c_304_n 0.0139118f $X=2.52 $Y=1.625 $X2=0 $Y2=0
cc_193 N_B_c_210_n N_A_55_155#_c_345_n 0.0179211f $X=3.165 $Y=1.51 $X2=0 $Y2=0
cc_194 N_B_c_218_n N_A_55_155#_c_345_n 0.0205436f $X=2.52 $Y=1.625 $X2=0 $Y2=0
cc_195 N_B_c_207_n N_A_55_155#_c_306_n 6.50136e-19 $X=1.625 $Y=1.51 $X2=0 $Y2=0
cc_196 N_B_c_208_n N_A_55_155#_c_306_n 0.0167588f $X=1.625 $Y=1.51 $X2=0 $Y2=0
cc_197 N_B_c_209_n N_A_55_155#_c_306_n 0.0163218f $X=3.165 $Y=1.51 $X2=0 $Y2=0
cc_198 N_B_c_210_n N_A_55_155#_c_306_n 0.0212927f $X=3.165 $Y=1.51 $X2=0 $Y2=0
cc_199 N_B_c_218_n N_A_55_155#_c_306_n 0.00574937f $X=2.52 $Y=1.625 $X2=0 $Y2=0
cc_200 N_B_c_218_n N_VPWR_M1012_s 0.00373625f $X=2.52 $Y=1.625 $X2=0 $Y2=0
cc_201 N_B_c_210_n N_VPWR_M1011_s 0.00340752f $X=3.165 $Y=1.51 $X2=0 $Y2=0
cc_202 N_B_M1012_g N_VPWR_c_397_n 0.00522564f $X=1.605 $Y=2.465 $X2=0 $Y2=0
cc_203 N_B_M1013_g N_VPWR_c_398_n 0.00380557f $X=3.185 $Y=2.465 $X2=0 $Y2=0
cc_204 N_B_M1012_g N_VPWR_c_402_n 0.00428252f $X=1.605 $Y=2.465 $X2=0 $Y2=0
cc_205 N_B_M1013_g N_VPWR_c_406_n 0.00428252f $X=3.185 $Y=2.465 $X2=0 $Y2=0
cc_206 N_B_M1012_g N_VPWR_c_395_n 0.00636597f $X=1.605 $Y=2.465 $X2=0 $Y2=0
cc_207 N_B_M1013_g N_VPWR_c_395_n 0.00627835f $X=3.185 $Y=2.465 $X2=0 $Y2=0
cc_208 N_B_c_218_n N_Y_M1002_d 0.00176891f $X=2.52 $Y=1.625 $X2=0 $Y2=0
cc_209 N_B_c_210_n N_Y_M1013_d 8.06206e-19 $X=3.165 $Y=1.51 $X2=0 $Y2=0
cc_210 N_B_M1012_g N_Y_c_476_n 0.00959653f $X=1.605 $Y=2.465 $X2=0 $Y2=0
cc_211 N_B_M1010_g N_Y_c_467_n 0.0122651f $X=3.145 $Y=0.775 $X2=0 $Y2=0
cc_212 N_B_c_209_n N_Y_c_467_n 0.00394319f $X=3.165 $Y=1.51 $X2=0 $Y2=0
cc_213 N_B_M1013_g N_Y_c_480_n 0.00947478f $X=3.185 $Y=2.465 $X2=0 $Y2=0
cc_214 N_B_M1012_g N_Y_c_483_n 0.00849639f $X=1.605 $Y=2.465 $X2=0 $Y2=0
cc_215 N_B_c_210_n N_Y_c_501_n 0.0543481f $X=3.165 $Y=1.51 $X2=0 $Y2=0
cc_216 N_B_c_218_n N_Y_c_501_n 0.00542259f $X=2.52 $Y=1.625 $X2=0 $Y2=0
cc_217 N_B_M1012_g N_Y_c_486_n 8.29611e-19 $X=1.605 $Y=2.465 $X2=0 $Y2=0
cc_218 N_B_M1013_g N_Y_c_486_n 5.95738e-19 $X=3.185 $Y=2.465 $X2=0 $Y2=0
cc_219 N_B_M1013_g N_Y_c_487_n 0.00832365f $X=3.185 $Y=2.465 $X2=0 $Y2=0
cc_220 N_B_M1008_g N_VGND_c_556_n 4.68429e-19 $X=1.585 $Y=0.775 $X2=0 $Y2=0
cc_221 N_B_M1010_g N_VGND_c_557_n 4.23668e-19 $X=3.145 $Y=0.775 $X2=0 $Y2=0
cc_222 N_B_M1008_g N_VGND_c_560_n 0.00286088f $X=1.585 $Y=0.775 $X2=0 $Y2=0
cc_223 N_B_M1010_g N_VGND_c_560_n 0.00286113f $X=3.145 $Y=0.775 $X2=0 $Y2=0
cc_224 N_B_M1008_g N_VGND_c_563_n 0.00384131f $X=1.585 $Y=0.775 $X2=0 $Y2=0
cc_225 N_B_M1010_g N_VGND_c_563_n 0.00382792f $X=3.145 $Y=0.775 $X2=0 $Y2=0
cc_226 N_B_M1008_g N_A_246_71#_c_599_n 0.00644683f $X=1.585 $Y=0.775 $X2=0 $Y2=0
cc_227 N_B_M1008_g N_A_246_71#_c_595_n 0.00835001f $X=1.585 $Y=0.775 $X2=0 $Y2=0
cc_228 N_B_M1010_g N_A_246_71#_c_595_n 0.0106749f $X=3.145 $Y=0.775 $X2=0 $Y2=0
cc_229 N_B_M1008_g N_A_246_71#_c_596_n 0.00210524f $X=1.585 $Y=0.775 $X2=0 $Y2=0
cc_230 N_B_M1010_g N_A_332_71#_c_622_n 0.00309355f $X=3.145 $Y=0.775 $X2=0 $Y2=0
cc_231 N_A_55_155#_M1002_g N_VPWR_c_397_n 0.00522564f $X=2.195 $Y=2.465 $X2=0
+ $Y2=0
cc_232 N_A_55_155#_M1011_g N_VPWR_c_398_n 0.00516054f $X=2.625 $Y=2.465 $X2=0
+ $Y2=0
cc_233 N_A_55_155#_M1002_g N_VPWR_c_404_n 0.00428252f $X=2.195 $Y=2.465 $X2=0
+ $Y2=0
cc_234 N_A_55_155#_M1011_g N_VPWR_c_404_n 0.00428252f $X=2.625 $Y=2.465 $X2=0
+ $Y2=0
cc_235 N_A_55_155#_M1002_g N_VPWR_c_395_n 0.00634064f $X=2.195 $Y=2.465 $X2=0
+ $Y2=0
cc_236 N_A_55_155#_M1011_g N_VPWR_c_395_n 0.00625301f $X=2.625 $Y=2.465 $X2=0
+ $Y2=0
cc_237 N_A_55_155#_M1002_g N_Y_c_476_n 0.00959653f $X=2.195 $Y=2.465 $X2=0 $Y2=0
cc_238 N_A_55_155#_c_301_n N_Y_c_467_n 0.0113835f $X=2.715 $Y=1.305 $X2=0 $Y2=0
cc_239 N_A_55_155#_M1011_g N_Y_c_480_n 0.00947478f $X=2.625 $Y=2.465 $X2=0 $Y2=0
cc_240 N_A_55_155#_M1002_g N_Y_c_483_n 8.29611e-19 $X=2.195 $Y=2.465 $X2=0 $Y2=0
cc_241 N_A_55_155#_c_298_n N_Y_c_501_n 0.00373101f $X=2.095 $Y=1.305 $X2=0 $Y2=0
cc_242 N_A_55_155#_c_301_n N_Y_c_501_n 0.00199585f $X=2.715 $Y=1.305 $X2=0 $Y2=0
cc_243 N_A_55_155#_c_315_n N_Y_c_501_n 0.014126f $X=1.89 $Y=1.09 $X2=0 $Y2=0
cc_244 N_A_55_155#_c_345_n N_Y_c_501_n 0.00808512f $X=2.185 $Y=1.47 $X2=0 $Y2=0
cc_245 N_A_55_155#_c_306_n N_Y_c_501_n 0.00844527f $X=2.625 $Y=1.47 $X2=0 $Y2=0
cc_246 N_A_55_155#_M1002_g N_Y_c_486_n 0.00851302f $X=2.195 $Y=2.465 $X2=0 $Y2=0
cc_247 N_A_55_155#_M1011_g N_Y_c_486_n 0.00834028f $X=2.625 $Y=2.465 $X2=0 $Y2=0
cc_248 N_A_55_155#_M1011_g N_Y_c_487_n 5.95738e-19 $X=2.625 $Y=2.465 $X2=0 $Y2=0
cc_249 N_A_55_155#_c_315_n N_VGND_M1009_d 0.00943666f $X=1.89 $Y=1.09 $X2=-0.19
+ $Y2=-0.245
cc_250 N_A_55_155#_c_315_n N_VGND_c_556_n 0.0218816f $X=1.89 $Y=1.09 $X2=0 $Y2=0
cc_251 N_A_55_155#_c_305_n N_VGND_c_556_n 6.12601e-19 $X=0.565 $Y=1 $X2=0 $Y2=0
cc_252 N_A_55_155#_c_298_n N_VGND_c_560_n 0.00286113f $X=2.095 $Y=1.305 $X2=0
+ $Y2=0
cc_253 N_A_55_155#_c_301_n N_VGND_c_560_n 0.00286113f $X=2.715 $Y=1.305 $X2=0
+ $Y2=0
cc_254 N_A_55_155#_c_298_n N_VGND_c_563_n 0.00390141f $X=2.095 $Y=1.305 $X2=0
+ $Y2=0
cc_255 N_A_55_155#_c_301_n N_VGND_c_563_n 0.00387359f $X=2.715 $Y=1.305 $X2=0
+ $Y2=0
cc_256 N_A_55_155#_c_305_n N_VGND_c_563_n 0.0176415f $X=0.565 $Y=1 $X2=0 $Y2=0
cc_257 N_A_55_155#_c_315_n N_A_246_71#_M1005_d 0.00608032f $X=1.89 $Y=1.09
+ $X2=-0.19 $Y2=-0.245
cc_258 N_A_55_155#_c_298_n N_A_246_71#_c_599_n 6.12907e-19 $X=2.095 $Y=1.305
+ $X2=0 $Y2=0
cc_259 N_A_55_155#_c_315_n N_A_246_71#_c_599_n 0.0150947f $X=1.89 $Y=1.09 $X2=0
+ $Y2=0
cc_260 N_A_55_155#_c_298_n N_A_246_71#_c_595_n 0.0105551f $X=2.095 $Y=1.305
+ $X2=0 $Y2=0
cc_261 N_A_55_155#_c_301_n N_A_246_71#_c_595_n 0.0101273f $X=2.715 $Y=1.305
+ $X2=0 $Y2=0
cc_262 N_A_55_155#_c_315_n N_A_246_71#_c_595_n 0.00306745f $X=1.89 $Y=1.09 $X2=0
+ $Y2=0
cc_263 N_A_55_155#_c_315_n N_A_332_71#_M1008_s 0.0055015f $X=1.89 $Y=1.09
+ $X2=-0.19 $Y2=-0.245
cc_264 N_A_55_155#_c_303_n N_A_332_71#_M1008_s 2.30296e-19 $X=1.975 $Y=1.345
+ $X2=-0.19 $Y2=-0.245
cc_265 N_A_55_155#_c_298_n N_A_332_71#_c_625_n 0.00202075f $X=2.095 $Y=1.305
+ $X2=0 $Y2=0
cc_266 N_A_55_155#_c_301_n N_A_332_71#_c_625_n 3.02071e-19 $X=2.715 $Y=1.305
+ $X2=0 $Y2=0
cc_267 N_A_55_155#_c_315_n N_A_332_71#_c_625_n 0.0199658f $X=1.89 $Y=1.09 $X2=0
+ $Y2=0
cc_268 N_A_55_155#_c_298_n N_A_332_71#_c_622_n 3.06942e-19 $X=2.095 $Y=1.305
+ $X2=0 $Y2=0
cc_269 N_A_55_155#_c_301_n N_A_332_71#_c_622_n 0.00250667f $X=2.715 $Y=1.305
+ $X2=0 $Y2=0
cc_270 N_A_55_155#_c_298_n N_A_332_71#_c_630_n 0.0101929f $X=2.095 $Y=1.305
+ $X2=0 $Y2=0
cc_271 N_A_55_155#_c_301_n N_A_332_71#_c_630_n 0.00859579f $X=2.715 $Y=1.305
+ $X2=0 $Y2=0
cc_272 N_A_55_155#_c_315_n N_A_332_71#_c_630_n 0.00139466f $X=1.89 $Y=1.09 $X2=0
+ $Y2=0
cc_273 N_A_55_155#_c_345_n N_A_332_71#_c_630_n 0.00383839f $X=2.185 $Y=1.47
+ $X2=0 $Y2=0
cc_274 N_VPWR_c_395_n N_Y_M1001_d 0.00223559f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_275 N_VPWR_c_395_n N_Y_M1002_d 0.00223559f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_276 N_VPWR_c_395_n N_Y_M1013_d 0.00223559f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_277 N_VPWR_M1012_s N_Y_c_476_n 0.00760535f $X=1.68 $Y=1.835 $X2=0 $Y2=0
cc_278 N_VPWR_c_397_n N_Y_c_476_n 0.0256295f $X=1.9 $Y=2.92 $X2=0 $Y2=0
cc_279 N_VPWR_c_402_n N_Y_c_476_n 0.00199329f $X=1.735 $Y=3.33 $X2=0 $Y2=0
cc_280 N_VPWR_c_404_n N_Y_c_476_n 0.00199329f $X=2.745 $Y=3.33 $X2=0 $Y2=0
cc_281 N_VPWR_c_395_n N_Y_c_476_n 0.00939785f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_282 N_VPWR_M1011_s N_Y_c_480_n 0.00669496f $X=2.7 $Y=1.835 $X2=0 $Y2=0
cc_283 N_VPWR_c_398_n N_Y_c_480_n 0.023271f $X=2.905 $Y=2.92 $X2=0 $Y2=0
cc_284 N_VPWR_c_404_n N_Y_c_480_n 0.00191958f $X=2.745 $Y=3.33 $X2=0 $Y2=0
cc_285 N_VPWR_c_406_n N_Y_c_480_n 0.00191958f $X=3.735 $Y=3.33 $X2=0 $Y2=0
cc_286 N_VPWR_c_395_n N_Y_c_480_n 0.00883602f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_287 N_VPWR_M1006_s N_Y_c_481_n 0.00969392f $X=3.69 $Y=1.835 $X2=0 $Y2=0
cc_288 N_VPWR_c_399_n N_Y_c_481_n 0.0167255f $X=3.83 $Y=2.92 $X2=0 $Y2=0
cc_289 N_VPWR_c_406_n N_Y_c_481_n 0.00191958f $X=3.735 $Y=3.33 $X2=0 $Y2=0
cc_290 N_VPWR_c_395_n N_Y_c_481_n 0.00461984f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_291 N_VPWR_c_396_n N_Y_c_483_n 0.0445173f $X=0.875 $Y=2.085 $X2=0 $Y2=0
cc_292 N_VPWR_c_402_n N_Y_c_483_n 0.0188913f $X=1.735 $Y=3.33 $X2=0 $Y2=0
cc_293 N_VPWR_c_395_n N_Y_c_483_n 0.012376f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_294 N_VPWR_c_404_n N_Y_c_486_n 0.0188913f $X=2.745 $Y=3.33 $X2=0 $Y2=0
cc_295 N_VPWR_c_395_n N_Y_c_486_n 0.012376f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_296 N_VPWR_c_406_n N_Y_c_487_n 0.0188913f $X=3.735 $Y=3.33 $X2=0 $Y2=0
cc_297 N_VPWR_c_395_n N_Y_c_487_n 0.012376f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_298 N_VPWR_c_399_n N_Y_c_470_n 0.00302528f $X=3.83 $Y=2.92 $X2=0 $Y2=0
cc_299 N_VPWR_c_408_n N_Y_c_470_n 0.00391173f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_300 N_VPWR_c_395_n N_Y_c_470_n 0.00688996f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_301 N_Y_c_467_n N_VGND_M1007_s 0.00749256f $X=3.96 $Y=1.09 $X2=0 $Y2=0
cc_302 N_Y_c_467_n N_VGND_c_557_n 0.0222789f $X=3.96 $Y=1.09 $X2=0 $Y2=0
cc_303 N_Y_c_467_n N_A_246_71#_M1010_d 0.00847118f $X=3.96 $Y=1.09 $X2=0 $Y2=0
cc_304 N_Y_M1000_d N_A_246_71#_c_595_n 0.00421368f $X=2.17 $Y=0.355 $X2=0 $Y2=0
cc_305 N_Y_c_467_n N_A_246_71#_c_595_n 0.00307977f $X=3.96 $Y=1.09 $X2=0 $Y2=0
cc_306 N_Y_c_467_n N_A_246_71#_c_612_n 0.0165443f $X=3.96 $Y=1.09 $X2=0 $Y2=0
cc_307 N_Y_c_467_n N_A_332_71#_M1003_s 0.0035081f $X=3.96 $Y=1.09 $X2=0 $Y2=0
cc_308 N_Y_c_467_n N_A_332_71#_c_622_n 0.0157865f $X=3.96 $Y=1.09 $X2=0 $Y2=0
cc_309 N_Y_M1000_d N_A_332_71#_c_630_n 0.00826045f $X=2.17 $Y=0.355 $X2=0 $Y2=0
cc_310 N_Y_c_467_n N_A_332_71#_c_630_n 0.00711037f $X=3.96 $Y=1.09 $X2=0 $Y2=0
cc_311 N_Y_c_501_n N_A_332_71#_c_630_n 0.0246044f $X=2.57 $Y=1.055 $X2=0 $Y2=0
cc_312 N_VGND_c_557_n N_A_246_71#_c_595_n 0.0110244f $X=3.83 $Y=0.72 $X2=0 $Y2=0
cc_313 N_VGND_c_560_n N_A_246_71#_c_595_n 0.126007f $X=3.665 $Y=0 $X2=0 $Y2=0
cc_314 N_VGND_c_563_n N_A_246_71#_c_595_n 0.0713253f $X=4.08 $Y=0 $X2=0 $Y2=0
cc_315 N_VGND_c_556_n N_A_246_71#_c_596_n 0.0110244f $X=0.94 $Y=0.705 $X2=0
+ $Y2=0
cc_316 N_VGND_c_560_n N_A_246_71#_c_596_n 0.0183317f $X=3.665 $Y=0 $X2=0 $Y2=0
cc_317 N_VGND_c_563_n N_A_246_71#_c_596_n 0.00995233f $X=4.08 $Y=0 $X2=0 $Y2=0
cc_318 N_A_246_71#_c_595_n N_A_332_71#_M1008_s 0.0026214f $X=3.265 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_319 N_A_246_71#_c_595_n N_A_332_71#_M1003_s 0.00176891f $X=3.265 $Y=0.34
+ $X2=0 $Y2=0
cc_320 N_A_246_71#_c_595_n N_A_332_71#_c_625_n 0.0738724f $X=3.265 $Y=0.34 $X2=0
+ $Y2=0
