* File: sky130_fd_sc_lp__nand2_8.spice
* Created: Wed Sep  2 10:02:57 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__nand2_8.pex.spice"
.subckt sky130_fd_sc_lp__nand2_8  VNB VPB B A VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A	A
* B	B
* VPB	VPB
* VNB	VNB
MM1001 N_A_27_65#_M1001_d N_B_M1001_g N_VGND_M1001_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75006.9 A=0.126 P=1.98 MULT=1
MM1008 N_A_27_65#_M1008_d N_B_M1008_g N_VGND_M1001_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75006.5 A=0.126 P=1.98 MULT=1
MM1012 N_A_27_65#_M1008_d N_B_M1012_g N_VGND_M1012_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.1 SB=75006
+ A=0.126 P=1.98 MULT=1
MM1014 N_A_27_65#_M1014_d N_B_M1014_g N_VGND_M1012_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.5
+ SB=75005.6 A=0.126 P=1.98 MULT=1
MM1019 N_A_27_65#_M1014_d N_B_M1019_g N_VGND_M1019_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.9
+ SB=75005.2 A=0.126 P=1.98 MULT=1
MM1024 N_A_27_65#_M1024_d N_B_M1024_g N_VGND_M1019_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002.3
+ SB=75004.8 A=0.126 P=1.98 MULT=1
MM1029 N_A_27_65#_M1024_d N_B_M1029_g N_VGND_M1029_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002.8
+ SB=75004.3 A=0.126 P=1.98 MULT=1
MM1031 N_A_27_65#_M1031_d N_B_M1031_g N_VGND_M1029_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75003.2
+ SB=75003.9 A=0.126 P=1.98 MULT=1
MM1003 N_Y_M1003_d N_A_M1003_g N_A_27_65#_M1031_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75003.6
+ SB=75003.5 A=0.126 P=1.98 MULT=1
MM1006 N_Y_M1003_d N_A_M1006_g N_A_27_65#_M1006_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.147 PD=1.12 PS=1.19 NRD=0 NRS=9.996 M=1 R=5.6 SA=75004.1
+ SB=75003 A=0.126 P=1.98 MULT=1
MM1009 N_Y_M1009_d N_A_M1009_g N_A_27_65#_M1006_s VNB NSHORT L=0.15 W=0.84
+ AD=0.147 AS=0.147 PD=1.19 PS=1.19 NRD=9.996 NRS=0 M=1 R=5.6 SA=75004.6
+ SB=75002.5 A=0.126 P=1.98 MULT=1
MM1013 N_Y_M1009_d N_A_M1013_g N_A_27_65#_M1013_s VNB NSHORT L=0.15 W=0.84
+ AD=0.147 AS=0.147 PD=1.19 PS=1.19 NRD=0 NRS=9.996 M=1 R=5.6 SA=75005.1
+ SB=75002 A=0.126 P=1.98 MULT=1
MM1020 N_Y_M1020_d N_A_M1020_g N_A_27_65#_M1013_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1302 AS=0.147 PD=1.15 PS=1.19 NRD=4.284 NRS=0 M=1 R=5.6 SA=75005.6
+ SB=75001.5 A=0.126 P=1.98 MULT=1
MM1023 N_Y_M1020_d N_A_M1023_g N_A_27_65#_M1023_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1302 AS=0.1176 PD=1.15 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75006 SB=75001.1
+ A=0.126 P=1.98 MULT=1
MM1026 N_Y_M1026_d N_A_M1026_g N_A_27_65#_M1023_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75006.4
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1027 N_Y_M1026_d N_A_M1027_g N_A_27_65#_M1027_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2394 PD=1.12 PS=2.25 NRD=0 NRS=0 M=1 R=5.6 SA=75006.9
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1000 N_Y_M1000_d N_B_M1000_g N_VPWR_M1000_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75006.9 A=0.189 P=2.82 MULT=1
MM1004 N_Y_M1000_d N_B_M1004_g N_VPWR_M1004_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75006.4 A=0.189 P=2.82 MULT=1
MM1010 N_Y_M1010_d N_B_M1010_g N_VPWR_M1004_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1 SB=75006
+ A=0.189 P=2.82 MULT=1
MM1015 N_Y_M1010_d N_B_M1015_g N_VPWR_M1015_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.5
+ SB=75005.6 A=0.189 P=2.82 MULT=1
MM1021 N_Y_M1021_d N_B_M1021_g N_VPWR_M1015_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.9
+ SB=75005.2 A=0.189 P=2.82 MULT=1
MM1022 N_Y_M1021_d N_B_M1022_g N_VPWR_M1022_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.3
+ SB=75004.7 A=0.189 P=2.82 MULT=1
MM1028 N_Y_M1028_d N_B_M1028_g N_VPWR_M1022_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.8
+ SB=75004.3 A=0.189 P=2.82 MULT=1
MM1030 N_Y_M1028_d N_B_M1030_g N_VPWR_M1030_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75003.2
+ SB=75003.9 A=0.189 P=2.82 MULT=1
MM1002 N_VPWR_M1030_s N_A_M1002_g N_Y_M1002_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75003.6
+ SB=75003.4 A=0.189 P=2.82 MULT=1
MM1005 N_VPWR_M1005_d N_A_M1005_g N_Y_M1002_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.2205 AS=0.1764 PD=1.61 PS=1.54 NRD=5.4569 NRS=0 M=1 R=8.4 SA=75004.1
+ SB=75003 A=0.189 P=2.82 MULT=1
MM1007 N_VPWR_M1005_d N_A_M1007_g N_Y_M1007_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.2205 AS=0.2205 PD=1.61 PS=1.61 NRD=5.4569 NRS=5.4569 M=1 R=8.4 SA=75004.6
+ SB=75002.5 A=0.189 P=2.82 MULT=1
MM1011 N_VPWR_M1011_d N_A_M1011_g N_Y_M1007_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.2205 AS=0.2205 PD=1.61 PS=1.61 NRD=5.4569 NRS=5.4569 M=1 R=8.4 SA=75005.1
+ SB=75002 A=0.189 P=2.82 MULT=1
MM1016 N_VPWR_M1011_d N_A_M1016_g N_Y_M1016_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.2205 AS=0.1953 PD=1.61 PS=1.57 NRD=5.4569 NRS=4.6886 M=1 R=8.4 SA=75005.6
+ SB=75001.5 A=0.189 P=2.82 MULT=1
MM1017 N_VPWR_M1017_d N_A_M1017_g N_Y_M1016_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1953 PD=1.54 PS=1.57 NRD=0 NRS=0 M=1 R=8.4 SA=75006 SB=75001.1
+ A=0.189 P=2.82 MULT=1
MM1018 N_VPWR_M1017_d N_A_M1018_g N_Y_M1018_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75006.4
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1025 N_VPWR_M1025_d N_A_M1025_g N_Y_M1018_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75006.9
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX32_noxref VNB VPB NWDIODE A=15.0319 P=19.85
c_66 VNB 0 1.52615e-19 $X=0 $Y=0
*
.include "sky130_fd_sc_lp__nand2_8.pxi.spice"
*
.ends
*
*
