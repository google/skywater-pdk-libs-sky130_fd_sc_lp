* File: sky130_fd_sc_lp__a32o_lp.pex.spice
* Created: Wed Sep  2 09:27:55 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A32O_LP%B2 3 7 9 10 11 12 15 16
c32 3 0 4.58742e-20 $X=0.56 $Y=2.595
r33 15 16 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.52 $Y=1.4
+ $X2=0.52 $Y2=1.4
r34 12 16 4.99854 $w=6.68e-07 $l=2.8e-07 $layer=LI1_cond $X=0.24 $Y=1.57
+ $X2=0.52 $Y2=1.57
r35 10 15 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.52 $Y=1.74
+ $X2=0.52 $Y2=1.4
r36 10 11 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.52 $Y=1.74
+ $X2=0.52 $Y2=1.905
r37 9 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.52 $Y=1.235
+ $X2=0.52 $Y2=1.4
r38 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.61 $Y=0.915 $X2=0.61
+ $Y2=1.235
r39 3 11 171.433 $w=2.5e-07 $l=6.9e-07 $layer=POLY_cond $X=0.56 $Y=2.595
+ $X2=0.56 $Y2=1.905
.ends

.subckt PM_SKY130_FD_SC_LP__A32O_LP%B1 3 4 6 9 10 11 14
r45 14 15 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.09 $Y=1.4
+ $X2=1.09 $Y2=1.4
r46 11 15 1.96371 $w=6.68e-07 $l=1.1e-07 $layer=LI1_cond $X=1.2 $Y=1.57 $X2=1.09
+ $Y2=1.57
r47 10 14 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.09 $Y=1.74
+ $X2=1.09 $Y2=1.4
r48 9 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.09 $Y=1.235
+ $X2=1.09 $Y2=1.4
r49 4 10 30.6163 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.09 $Y=1.905
+ $X2=1.09 $Y2=1.74
r50 4 6 171.433 $w=2.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.09 $Y=1.905 $X2=1.09
+ $Y2=2.595
r51 3 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1 $Y=0.915 $X2=1
+ $Y2=1.235
.ends

.subckt PM_SKY130_FD_SC_LP__A32O_LP%A1 3 6 9 10 11 12 15 16
r44 15 16 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.66 $Y=1.4
+ $X2=1.66 $Y2=1.4
r45 12 16 9.25447 $w=3.28e-07 $l=2.65e-07 $layer=LI1_cond $X=1.66 $Y=1.665
+ $X2=1.66 $Y2=1.4
r46 10 15 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.66 $Y=1.74
+ $X2=1.66 $Y2=1.4
r47 10 11 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.66 $Y=1.74
+ $X2=1.66 $Y2=1.905
r48 9 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.66 $Y=1.235
+ $X2=1.66 $Y2=1.4
r49 6 11 171.433 $w=2.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.62 $Y=2.595
+ $X2=1.62 $Y2=1.905
r50 3 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.57 $Y=0.915 $X2=1.57
+ $Y2=1.235
.ends

.subckt PM_SKY130_FD_SC_LP__A32O_LP%A2 3 4 6 9 10 11 12 13 18
c45 9 0 1.03481e-19 $X=2.23 $Y=1.235
r46 18 19 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.23 $Y=1.4
+ $X2=2.23 $Y2=1.4
r47 13 19 8.72564 $w=3.48e-07 $l=2.65e-07 $layer=LI1_cond $X=2.22 $Y=1.665
+ $X2=2.22 $Y2=1.4
r48 12 19 3.45733 $w=3.48e-07 $l=1.05e-07 $layer=LI1_cond $X=2.22 $Y=1.295
+ $X2=2.22 $Y2=1.4
r49 11 12 12.183 $w=3.48e-07 $l=3.7e-07 $layer=LI1_cond $X=2.22 $Y=0.925
+ $X2=2.22 $Y2=1.295
r50 10 18 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.23 $Y=1.74
+ $X2=2.23 $Y2=1.4
r51 9 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.23 $Y=1.235
+ $X2=2.23 $Y2=1.4
r52 4 10 30.6163 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.23 $Y=1.905
+ $X2=2.23 $Y2=1.74
r53 4 6 171.433 $w=2.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.23 $Y=1.905 $X2=2.23
+ $Y2=2.595
r54 3 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.14 $Y=0.915 $X2=2.14
+ $Y2=1.235
.ends

.subckt PM_SKY130_FD_SC_LP__A32O_LP%A3 3 7 9 15
r39 13 15 57.7042 $w=3.3e-07 $l=3.3e-07 $layer=POLY_cond $X=2.76 $Y=1.715
+ $X2=3.09 $Y2=1.715
r40 11 13 8.74306 $w=3.3e-07 $l=5e-08 $layer=POLY_cond $X=2.71 $Y=1.715 $X2=2.76
+ $Y2=1.715
r41 9 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.09
+ $Y=1.715 $X2=3.09 $Y2=1.715
r42 5 13 9.34494 $w=2.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.76 $Y=1.88
+ $X2=2.76 $Y2=1.715
r43 5 7 177.644 $w=2.5e-07 $l=7.15e-07 $layer=POLY_cond $X=2.76 $Y=1.88 $X2=2.76
+ $Y2=2.595
r44 1 11 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.71 $Y=1.55
+ $X2=2.71 $Y2=1.715
r45 1 3 325.606 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=2.71 $Y=1.55 $X2=2.71
+ $Y2=0.915
.ends

.subckt PM_SKY130_FD_SC_LP__A32O_LP%A_137_419# 1 2 7 9 13 14 16 21 23 24 27 29
+ 30 32 34 35 39 42 46
c109 42 0 1.03481e-19 $X=2.66 $Y=1.285
r110 40 46 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=3.52 $Y=0.43
+ $X2=3.725 $Y2=0.43
r111 40 43 32.3493 $w=3.3e-07 $l=1.85e-07 $layer=POLY_cond $X=3.52 $Y=0.43
+ $X2=3.335 $Y2=0.43
r112 39 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.52
+ $Y=0.43 $X2=3.52 $Y2=0.43
r113 37 39 26.8903 $w=3.28e-07 $l=7.7e-07 $layer=LI1_cond $X=3.52 $Y=1.2
+ $X2=3.52 $Y2=0.43
r114 36 42 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.745 $Y=1.285
+ $X2=2.66 $Y2=1.285
r115 35 37 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.355 $Y=1.285
+ $X2=3.52 $Y2=1.2
r116 35 36 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=3.355 $Y=1.285
+ $X2=2.745 $Y2=1.285
r117 33 42 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.66 $Y=1.37
+ $X2=2.66 $Y2=1.285
r118 33 34 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=2.66 $Y=1.37
+ $X2=2.66 $Y2=2.085
r119 32 42 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.66 $Y=1.2 $X2=2.66
+ $Y2=1.285
r120 31 32 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=2.66 $Y=0.63
+ $X2=2.66 $Y2=1.2
r121 29 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.575 $Y=0.545
+ $X2=2.66 $Y2=0.63
r122 29 30 68.8289 $w=1.68e-07 $l=1.055e-06 $layer=LI1_cond $X=2.575 $Y=0.545
+ $X2=1.52 $Y2=0.545
r123 25 30 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.355 $Y=0.63
+ $X2=1.52 $Y2=0.545
r124 25 27 8.3814 $w=3.28e-07 $l=2.4e-07 $layer=LI1_cond $X=1.355 $Y=0.63
+ $X2=1.355 $Y2=0.87
r125 23 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.575 $Y=2.17
+ $X2=2.66 $Y2=2.085
r126 23 24 103.406 $w=1.68e-07 $l=1.585e-06 $layer=LI1_cond $X=2.575 $Y=2.17
+ $X2=0.99 $Y2=2.17
r127 19 24 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.825 $Y=2.255
+ $X2=0.99 $Y2=2.17
r128 19 21 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=0.825 $Y=2.255
+ $X2=0.825 $Y2=2.4
r129 14 18 40.9178 $w=2.5e-07 $l=1.25e-07 $layer=POLY_cond $X=3.775 $Y=1.475
+ $X2=3.775 $Y2=1.35
r130 14 16 278.268 $w=2.5e-07 $l=1.12e-06 $layer=POLY_cond $X=3.775 $Y=1.475
+ $X2=3.775 $Y2=2.595
r131 13 18 223.053 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.725 $Y=0.915
+ $X2=3.725 $Y2=1.35
r132 10 46 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.725 $Y=0.595
+ $X2=3.725 $Y2=0.43
r133 10 13 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=3.725 $Y=0.595
+ $X2=3.725 $Y2=0.915
r134 7 43 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.335 $Y=0.595
+ $X2=3.335 $Y2=0.43
r135 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=3.335 $Y=0.595
+ $X2=3.335 $Y2=0.915
r136 2 21 600 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_PDIFF $count=1 $X=0.685
+ $Y=2.095 $X2=0.825 $Y2=2.4
r137 1 27 182 $w=1.7e-07 $l=3.52987e-07 $layer=licon1_NDIFF $count=1 $X=1.075
+ $Y=0.705 $X2=1.355 $Y2=0.87
.ends

.subckt PM_SKY130_FD_SC_LP__A32O_LP%A_30_419# 1 2 3 12 14 15 19 20 21 24
c49 21 0 4.58742e-20 $X=1.52 $Y=2.52
r50 22 24 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=2.495 $Y=2.605
+ $X2=2.495 $Y2=2.75
r51 20 22 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.33 $Y=2.52
+ $X2=2.495 $Y2=2.605
r52 20 21 52.8449 $w=1.68e-07 $l=8.1e-07 $layer=LI1_cond $X=2.33 $Y=2.52
+ $X2=1.52 $Y2=2.52
r53 17 19 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=1.355 $Y=2.895
+ $X2=1.355 $Y2=2.75
r54 16 21 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.355 $Y=2.605
+ $X2=1.52 $Y2=2.52
r55 16 19 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=1.355 $Y=2.605
+ $X2=1.355 $Y2=2.75
r56 14 17 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.19 $Y=2.98
+ $X2=1.355 $Y2=2.895
r57 14 15 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=1.19 $Y=2.98
+ $X2=0.46 $Y2=2.98
r58 10 15 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.295 $Y=2.895
+ $X2=0.46 $Y2=2.98
r59 10 12 22.525 $w=3.28e-07 $l=6.45e-07 $layer=LI1_cond $X=0.295 $Y=2.895
+ $X2=0.295 $Y2=2.25
r60 3 24 600 $w=1.7e-07 $l=7.21613e-07 $layer=licon1_PDIFF $count=1 $X=2.355
+ $Y=2.095 $X2=2.495 $Y2=2.75
r61 2 19 600 $w=1.7e-07 $l=7.21613e-07 $layer=licon1_PDIFF $count=1 $X=1.215
+ $Y=2.095 $X2=1.355 $Y2=2.75
r62 1 12 300 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_PDIFF $count=2 $X=0.15
+ $Y=2.095 $X2=0.295 $Y2=2.25
.ends

.subckt PM_SKY130_FD_SC_LP__A32O_LP%VPWR 1 2 9 13 18 19 20 29 35 36 39
r52 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r53 36 40 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.12 $Y2=3.33
r54 35 36 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r55 33 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.255 $Y=3.33
+ $X2=3.09 $Y2=3.33
r56 33 35 53.8235 $w=1.68e-07 $l=8.25e-07 $layer=LI1_cond $X=3.255 $Y=3.33
+ $X2=4.08 $Y2=3.33
r57 32 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r58 31 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r59 29 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.925 $Y=3.33
+ $X2=3.09 $Y2=3.33
r60 29 31 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=2.925 $Y=3.33
+ $X2=2.64 $Y2=3.33
r61 27 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r62 24 28 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.68 $Y2=3.33
r63 23 27 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=0.24 $Y=3.33
+ $X2=1.68 $Y2=3.33
r64 23 24 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r65 20 32 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r66 20 28 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r67 18 27 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=1.72 $Y=3.33 $X2=1.68
+ $Y2=3.33
r68 18 19 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.72 $Y=3.33
+ $X2=1.885 $Y2=3.33
r69 17 31 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=2.05 $Y=3.33 $X2=2.64
+ $Y2=3.33
r70 17 19 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.05 $Y=3.33
+ $X2=1.885 $Y2=3.33
r71 13 16 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=3.09 $Y=2.24 $X2=3.09
+ $Y2=2.95
r72 11 39 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.09 $Y=3.245
+ $X2=3.09 $Y2=3.33
r73 11 16 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=3.09 $Y=3.245
+ $X2=3.09 $Y2=2.95
r74 7 19 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.885 $Y=3.245
+ $X2=1.885 $Y2=3.33
r75 7 9 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.885 $Y=3.245
+ $X2=1.885 $Y2=2.95
r76 2 16 400 $w=1.7e-07 $l=9.51998e-07 $layer=licon1_PDIFF $count=1 $X=2.885
+ $Y=2.095 $X2=3.09 $Y2=2.95
r77 2 13 400 $w=1.7e-07 $l=2.67862e-07 $layer=licon1_PDIFF $count=1 $X=2.885
+ $Y=2.095 $X2=3.09 $Y2=2.24
r78 1 9 600 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=1.745
+ $Y=2.095 $X2=1.885 $Y2=2.95
.ends

.subckt PM_SKY130_FD_SC_LP__A32O_LP%X 1 2 7 8 9 10 11 12 13
r15 12 13 12.5413 $w=3.38e-07 $l=3.7e-07 $layer=LI1_cond $X=4.035 $Y=2.405
+ $X2=4.035 $Y2=2.775
r16 12 34 5.59274 $w=3.38e-07 $l=1.65e-07 $layer=LI1_cond $X=4.035 $Y=2.405
+ $X2=4.035 $Y2=2.24
r17 11 34 6.94855 $w=3.38e-07 $l=2.05e-07 $layer=LI1_cond $X=4.035 $Y=2.035
+ $X2=4.035 $Y2=2.24
r18 10 11 12.5413 $w=3.38e-07 $l=3.7e-07 $layer=LI1_cond $X=4.035 $Y=1.665
+ $X2=4.035 $Y2=2.035
r19 9 10 12.5413 $w=3.38e-07 $l=3.7e-07 $layer=LI1_cond $X=4.035 $Y=1.295
+ $X2=4.035 $Y2=1.665
r20 8 9 12.8802 $w=3.38e-07 $l=3.8e-07 $layer=LI1_cond $X=4.035 $Y=0.915
+ $X2=4.035 $Y2=1.295
r21 7 8 12.2023 $w=3.38e-07 $l=3.6e-07 $layer=LI1_cond $X=4.035 $Y=0.555
+ $X2=4.035 $Y2=0.915
r22 2 34 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=3.9
+ $Y=2.095 $X2=4.04 $Y2=2.24
r23 1 8 182 $w=1.7e-07 $l=3.18119e-07 $layer=licon1_NDIFF $count=1 $X=3.8
+ $Y=0.705 $X2=4.03 $Y2=0.915
.ends

.subckt PM_SKY130_FD_SC_LP__A32O_LP%VGND 1 2 7 9 13 15 17 27 28 34
r37 34 35 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r38 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r39 28 35 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.12
+ $Y2=0
r40 27 28 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r41 25 34 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.175 $Y=0 $X2=3.05
+ $Y2=0
r42 25 27 59.0428 $w=1.68e-07 $l=9.05e-07 $layer=LI1_cond $X=3.175 $Y=0 $X2=4.08
+ $Y2=0
r43 24 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r44 23 24 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r45 21 32 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r46 20 23 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=0.72 $Y=0 $X2=2.64
+ $Y2=0
r47 20 21 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r48 18 31 4.53027 $w=1.7e-07 $l=2.8e-07 $layer=LI1_cond $X=0.56 $Y=0 $X2=0.28
+ $Y2=0
r49 18 20 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=0.56 $Y=0 $X2=0.72
+ $Y2=0
r50 17 34 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.925 $Y=0 $X2=3.05
+ $Y2=0
r51 17 23 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=2.925 $Y=0 $X2=2.64
+ $Y2=0
r52 15 24 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r53 15 21 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=2.16 $Y=0 $X2=0.72
+ $Y2=0
r54 11 34 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.05 $Y=0.085
+ $X2=3.05 $Y2=0
r55 11 13 35.2648 $w=2.48e-07 $l=7.65e-07 $layer=LI1_cond $X=3.05 $Y=0.085
+ $X2=3.05 $Y2=0.85
r56 7 31 3.23591 $w=3.3e-07 $l=1.51658e-07 $layer=LI1_cond $X=0.395 $Y=0.085
+ $X2=0.28 $Y2=0
r57 7 9 27.4142 $w=3.28e-07 $l=7.85e-07 $layer=LI1_cond $X=0.395 $Y=0.085
+ $X2=0.395 $Y2=0.87
r58 2 13 182 $w=1.7e-07 $l=2.88531e-07 $layer=licon1_NDIFF $count=1 $X=2.785
+ $Y=0.705 $X2=3.01 $Y2=0.85
r59 1 9 182 $w=1.7e-07 $l=2.26164e-07 $layer=licon1_NDIFF $count=1 $X=0.25
+ $Y=0.705 $X2=0.395 $Y2=0.87
.ends

