* NGSPICE file created from sky130_fd_sc_lp__nand3_lp.ext - technology: sky130A

.subckt sky130_fd_sc_lp__nand3_lp A B C VGND VNB VPB VPWR Y
M1000 Y C VPWR VPB phighvt w=1e+06u l=250000u
+  ad=5.65e+11p pd=5.13e+06u as=6.1e+11p ps=5.22e+06u
M1001 Y A a_233_47# VNB nshort w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=1.764e+11p ps=1.68e+06u
M1002 Y A VPWR VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1003 VPWR B Y VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_155_47# C VGND VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=1.197e+11p ps=1.41e+06u
M1005 a_233_47# B a_155_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

