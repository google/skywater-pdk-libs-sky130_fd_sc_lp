* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__einvp_1 A TE VGND VNB VPB VPWR Z
M1000 a_207_302# TE VPWR VPB phighvt w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=3.175e+11p ps=2.78e+06u
M1001 VGND TE a_128_47# VNB nshort w=840000u l=150000u
+  ad=4.347e+11p pd=3.22e+06u as=2.016e+11p ps=2.16e+06u
M1002 VPWR a_207_302# a_161_400# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=2.3e+11p ps=2.46e+06u
M1003 a_128_47# A Z VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=2.226e+11p ps=2.21e+06u
M1004 a_207_302# TE VGND VNB nshort w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=0p ps=0u
M1005 a_161_400# A Z VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=2.85e+11p ps=2.57e+06u
.ends
