* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__dlxtn_1 D GATE_N VGND VNB VPB VPWR Q
X0 VPWR a_842_413# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X1 a_656_47# a_228_129# a_656_481# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 VGND GATE_N a_228_129# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 VPWR GATE_N a_228_129# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X4 VPWR a_656_481# a_842_413# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X5 VGND a_656_481# a_842_413# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X6 VGND a_842_413# Q VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X7 a_342_481# a_228_129# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X8 a_342_481# a_228_129# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 a_656_481# a_342_481# a_836_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 a_764_481# a_842_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X11 a_836_47# a_842_413# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 a_59_129# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X13 a_656_481# a_228_129# a_764_481# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X14 VPWR a_59_129# a_584_481# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X15 a_584_481# a_342_481# a_656_481# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X16 VGND a_59_129# a_656_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X17 a_59_129# D VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
