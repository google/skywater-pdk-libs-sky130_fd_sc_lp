* File: sky130_fd_sc_lp__ebufn_8.pex.spice
* Created: Fri Aug 28 10:31:56 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__EBUFN_8%A_84_21# 1 2 9 13 17 21 25 29 33 37 41 45 49
+ 53 57 61 65 69 76 79 80 81 82 86 88 92 95 98 107 108 121
c276 97 0 1.11562e-19 $X=3.465 $Y=1.48
c277 82 0 1.46525e-19 $X=8.365 $Y=2.4
c278 81 0 5.76786e-20 $X=6.725 $Y=2.11
c279 69 0 1.61246e-19 $X=3.505 $Y=2.465
c280 13 0 1.6164e-19 $X=0.495 $Y=2.465
r281 118 119 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=2.645 $Y=1.48
+ $X2=3.075 $Y2=1.48
r282 117 118 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=2.215 $Y=1.48
+ $X2=2.645 $Y2=1.48
r283 116 117 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=1.785 $Y=1.48
+ $X2=2.215 $Y2=1.48
r284 115 116 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=1.355 $Y=1.48
+ $X2=1.785 $Y2=1.48
r285 111 113 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=0.495 $Y=1.48
+ $X2=0.925 $Y2=1.48
r286 109 110 4.5286 $w=6.58e-07 $l=8.5e-08 $layer=LI1_cond $X=8.695 $Y=2.4
+ $X2=8.695 $Y2=2.485
r287 107 109 7.61141 $w=6.58e-07 $l=4.2e-07 $layer=LI1_cond $X=8.695 $Y=1.98
+ $X2=8.695 $Y2=2.4
r288 107 108 10.5469 $w=6.58e-07 $l=1.65e-07 $layer=LI1_cond $X=8.695 $Y=1.98
+ $X2=8.695 $Y2=1.815
r289 98 100 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=7.58 $Y=2.11
+ $X2=7.58 $Y2=2.4
r290 96 121 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=3.3 $Y=1.48
+ $X2=3.505 $Y2=1.48
r291 96 119 39.3438 $w=3.3e-07 $l=2.25e-07 $layer=POLY_cond $X=3.3 $Y=1.48
+ $X2=3.075 $Y2=1.48
r292 95 97 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=3.3 $Y=1.48
+ $X2=3.465 $Y2=1.48
r293 95 96 41.5086 $w=1.7e-07 $l=5.95e-07 $layer=licon1_POLY $count=3 $X=3.3
+ $Y=1.48 $X2=3.3 $Y2=1.48
r294 92 110 14.8421 $w=3.28e-07 $l=4.25e-07 $layer=LI1_cond $X=8.86 $Y=2.91
+ $X2=8.86 $Y2=2.485
r295 86 102 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=8.86 $Y=0.925
+ $X2=8.45 $Y2=0.925
r296 86 88 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=8.86 $Y=0.84
+ $X2=8.86 $Y2=0.42
r297 84 102 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.45 $Y=1.01
+ $X2=8.45 $Y2=0.925
r298 84 108 52.5187 $w=1.68e-07 $l=8.05e-07 $layer=LI1_cond $X=8.45 $Y=1.01
+ $X2=8.45 $Y2=1.815
r299 83 100 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.665 $Y=2.4
+ $X2=7.58 $Y2=2.4
r300 82 109 8.93547 $w=1.7e-07 $l=3.3e-07 $layer=LI1_cond $X=8.365 $Y=2.4
+ $X2=8.695 $Y2=2.4
r301 82 83 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=8.365 $Y=2.4
+ $X2=7.665 $Y2=2.4
r302 80 98 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.495 $Y=2.11
+ $X2=7.58 $Y2=2.11
r303 80 81 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=7.495 $Y=2.11
+ $X2=6.725 $Y2=2.11
r304 79 81 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.64 $Y=2.025
+ $X2=6.725 $Y2=2.11
r305 78 79 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=6.64 $Y=1.645
+ $X2=6.64 $Y2=2.025
r306 76 78 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.555 $Y=1.56
+ $X2=6.64 $Y2=1.645
r307 76 97 201.594 $w=1.68e-07 $l=3.09e-06 $layer=LI1_cond $X=6.555 $Y=1.56
+ $X2=3.465 $Y2=1.56
r308 74 115 16.6118 $w=3.3e-07 $l=9.5e-08 $layer=POLY_cond $X=1.26 $Y=1.48
+ $X2=1.355 $Y2=1.48
r309 74 113 58.5785 $w=3.3e-07 $l=3.35e-07 $layer=POLY_cond $X=1.26 $Y=1.48
+ $X2=0.925 $Y2=1.48
r310 73 95 71.2419 $w=3.28e-07 $l=2.04e-06 $layer=LI1_cond $X=1.26 $Y=1.48
+ $X2=3.3 $Y2=1.48
r311 73 74 41.5086 $w=1.7e-07 $l=5.95e-07 $layer=licon1_POLY $count=3 $X=1.26
+ $Y=1.48 $X2=1.26 $Y2=1.48
r312 67 121 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.505 $Y=1.645
+ $X2=3.505 $Y2=1.48
r313 67 69 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=3.505 $Y=1.645
+ $X2=3.505 $Y2=2.465
r314 63 121 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.505 $Y=1.315
+ $X2=3.505 $Y2=1.48
r315 63 65 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.505 $Y=1.315
+ $X2=3.505 $Y2=0.655
r316 59 119 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.075 $Y=1.645
+ $X2=3.075 $Y2=1.48
r317 59 61 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=3.075 $Y=1.645
+ $X2=3.075 $Y2=2.465
r318 55 119 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.075 $Y=1.315
+ $X2=3.075 $Y2=1.48
r319 55 57 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.075 $Y=1.315
+ $X2=3.075 $Y2=0.655
r320 51 118 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.645 $Y=1.645
+ $X2=2.645 $Y2=1.48
r321 51 53 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=2.645 $Y=1.645
+ $X2=2.645 $Y2=2.465
r322 47 118 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.645 $Y=1.315
+ $X2=2.645 $Y2=1.48
r323 47 49 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.645 $Y=1.315
+ $X2=2.645 $Y2=0.655
r324 43 117 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.215 $Y=1.645
+ $X2=2.215 $Y2=1.48
r325 43 45 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=2.215 $Y=1.645
+ $X2=2.215 $Y2=2.465
r326 39 117 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.215 $Y=1.315
+ $X2=2.215 $Y2=1.48
r327 39 41 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.215 $Y=1.315
+ $X2=2.215 $Y2=0.655
r328 35 116 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.785 $Y=1.645
+ $X2=1.785 $Y2=1.48
r329 35 37 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=1.785 $Y=1.645
+ $X2=1.785 $Y2=2.465
r330 31 116 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.785 $Y=1.315
+ $X2=1.785 $Y2=1.48
r331 31 33 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.785 $Y=1.315
+ $X2=1.785 $Y2=0.655
r332 27 115 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.355 $Y=1.645
+ $X2=1.355 $Y2=1.48
r333 27 29 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=1.355 $Y=1.645
+ $X2=1.355 $Y2=2.465
r334 23 115 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.355 $Y=1.315
+ $X2=1.355 $Y2=1.48
r335 23 25 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.355 $Y=1.315
+ $X2=1.355 $Y2=0.655
r336 19 113 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.925 $Y=1.645
+ $X2=0.925 $Y2=1.48
r337 19 21 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=0.925 $Y=1.645
+ $X2=0.925 $Y2=2.465
r338 15 113 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.925 $Y=1.315
+ $X2=0.925 $Y2=1.48
r339 15 17 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.925 $Y=1.315
+ $X2=0.925 $Y2=0.655
r340 11 111 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=1.645
+ $X2=0.495 $Y2=1.48
r341 11 13 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=0.495 $Y=1.645
+ $X2=0.495 $Y2=2.465
r342 7 111 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=1.315
+ $X2=0.495 $Y2=1.48
r343 7 9 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.495 $Y=1.315
+ $X2=0.495 $Y2=0.655
r344 2 107 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=8.72
+ $Y=1.835 $X2=8.86 $Y2=1.98
r345 2 92 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=8.72
+ $Y=1.835 $X2=8.86 $Y2=2.91
r346 1 88 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=8.72
+ $Y=0.235 $X2=8.86 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__EBUFN_8%A_772_21# 1 2 7 9 10 11 12 14 15 17 19 20 22
+ 24 25 27 29 30 32 34 35 37 39 40 42 44 45 48 49 50 51 52 53 54 55 57 59 60 61
+ 63 64 68
c177 64 0 3.60707e-20 $X=7.58 $Y=0.42
c178 11 0 1.11562e-19 $X=4.01 $Y=1.26
c179 7 0 5.58653e-20 $X=3.935 $Y=1.185
r180 68 71 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=8 $Y=1.77 $X2=8
+ $Y2=1.98
r181 63 67 16.0268 $w=7.48e-07 $l=5.9e-07 $layer=LI1_cond $X=7.79 $Y=0.42
+ $X2=7.79 $Y2=1.01
r182 63 64 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.58
+ $Y=0.42 $X2=7.58 $Y2=0.42
r183 60 68 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.835 $Y=1.77 $X2=8
+ $Y2=1.77
r184 60 61 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=7.835 $Y=1.77
+ $X2=7.635 $Y2=1.77
r185 59 61 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=7.525 $Y=1.685
+ $X2=7.635 $Y2=1.77
r186 59 67 35.359 $w=2.18e-07 $l=6.75e-07 $layer=LI1_cond $X=7.525 $Y=1.685
+ $X2=7.525 $Y2=1.01
r187 56 64 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=7.58 $Y=0.76
+ $X2=7.58 $Y2=0.42
r188 56 57 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.58 $Y=0.76
+ $X2=7.58 $Y2=0.925
r189 48 57 133.319 $w=1.5e-07 $l=2.6e-07 $layer=POLY_cond $X=7.49 $Y=1.185
+ $X2=7.49 $Y2=0.925
r190 46 55 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.02 $Y=1.26
+ $X2=6.945 $Y2=1.26
r191 45 48 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.415 $Y=1.26
+ $X2=7.49 $Y2=1.185
r192 45 46 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=7.415 $Y=1.26
+ $X2=7.02 $Y2=1.26
r193 42 55 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.945 $Y=1.185
+ $X2=6.945 $Y2=1.26
r194 42 44 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=6.945 $Y=1.185
+ $X2=6.945 $Y2=0.655
r195 41 54 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.59 $Y=1.26
+ $X2=6.515 $Y2=1.26
r196 40 55 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.87 $Y=1.26
+ $X2=6.945 $Y2=1.26
r197 40 41 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=6.87 $Y=1.26
+ $X2=6.59 $Y2=1.26
r198 37 54 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.515 $Y=1.185
+ $X2=6.515 $Y2=1.26
r199 37 39 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=6.515 $Y=1.185
+ $X2=6.515 $Y2=0.655
r200 36 53 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.16 $Y=1.26
+ $X2=6.085 $Y2=1.26
r201 35 54 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.44 $Y=1.26
+ $X2=6.515 $Y2=1.26
r202 35 36 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=6.44 $Y=1.26
+ $X2=6.16 $Y2=1.26
r203 32 53 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.085 $Y=1.185
+ $X2=6.085 $Y2=1.26
r204 32 34 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=6.085 $Y=1.185
+ $X2=6.085 $Y2=0.655
r205 31 52 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.73 $Y=1.26
+ $X2=5.655 $Y2=1.26
r206 30 53 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.01 $Y=1.26
+ $X2=6.085 $Y2=1.26
r207 30 31 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=6.01 $Y=1.26
+ $X2=5.73 $Y2=1.26
r208 27 52 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.655 $Y=1.185
+ $X2=5.655 $Y2=1.26
r209 27 29 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=5.655 $Y=1.185
+ $X2=5.655 $Y2=0.655
r210 26 51 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.3 $Y=1.26
+ $X2=5.225 $Y2=1.26
r211 25 52 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.58 $Y=1.26
+ $X2=5.655 $Y2=1.26
r212 25 26 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=5.58 $Y=1.26
+ $X2=5.3 $Y2=1.26
r213 22 51 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.225 $Y=1.185
+ $X2=5.225 $Y2=1.26
r214 22 24 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=5.225 $Y=1.185
+ $X2=5.225 $Y2=0.655
r215 21 50 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.87 $Y=1.26
+ $X2=4.795 $Y2=1.26
r216 20 51 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.15 $Y=1.26
+ $X2=5.225 $Y2=1.26
r217 20 21 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=5.15 $Y=1.26
+ $X2=4.87 $Y2=1.26
r218 17 50 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.795 $Y=1.185
+ $X2=4.795 $Y2=1.26
r219 17 19 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=4.795 $Y=1.185
+ $X2=4.795 $Y2=0.655
r220 16 49 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.44 $Y=1.26
+ $X2=4.365 $Y2=1.26
r221 15 50 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.72 $Y=1.26
+ $X2=4.795 $Y2=1.26
r222 15 16 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=4.72 $Y=1.26
+ $X2=4.44 $Y2=1.26
r223 12 49 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.365 $Y=1.185
+ $X2=4.365 $Y2=1.26
r224 12 14 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=4.365 $Y=1.185
+ $X2=4.365 $Y2=0.655
r225 10 49 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.29 $Y=1.26
+ $X2=4.365 $Y2=1.26
r226 10 11 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=4.29 $Y=1.26
+ $X2=4.01 $Y2=1.26
r227 7 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.935 $Y=1.185
+ $X2=4.01 $Y2=1.26
r228 7 9 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=3.935 $Y=1.185
+ $X2=3.935 $Y2=0.655
r229 2 71 600 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=7.855
+ $Y=1.835 $X2=8 $Y2=1.98
r230 1 63 91 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=2 $X=7.855
+ $Y=0.235 $X2=8 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__EBUFN_8%TE_B 1 3 4 5 6 8 9 11 13 14 16 18 19 21 23
+ 24 26 28 29 31 33 34 36 38 39 43 46 47 48 49 50 51 52 53 54 57 58 59 61
c196 34 0 1.85809e-19 $X=6.87 $Y=1.65
c197 31 0 1.57686e-19 $X=6.515 $Y=1.725
c198 26 0 5.76786e-20 $X=6.085 $Y=1.725
c199 1 0 5.74299e-20 $X=3.935 $Y=1.725
r200 57 59 46.2775 $w=4.25e-07 $l=1.65e-07 $layer=POLY_cond $X=8.077 $Y=1.35
+ $X2=8.077 $Y2=1.185
r201 57 58 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.03
+ $Y=1.35 $X2=8.03 $Y2=1.35
r202 54 58 3.78414 $w=3.33e-07 $l=1.1e-07 $layer=LI1_cond $X=7.92 $Y=1.347
+ $X2=8.03 $Y2=1.347
r203 46 61 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=8.215 $Y=2.465
+ $X2=8.215 $Y2=1.725
r204 43 59 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=8.215 $Y=0.655
+ $X2=8.215 $Y2=1.185
r205 40 53 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.02 $Y=1.65
+ $X2=6.945 $Y2=1.65
r206 39 61 34.5001 $w=4.25e-07 $l=7.5e-08 $layer=POLY_cond $X=8.077 $Y=1.65
+ $X2=8.077 $Y2=1.725
r207 39 57 39.2579 $w=4.25e-07 $l=3e-07 $layer=POLY_cond $X=8.077 $Y=1.65
+ $X2=8.077 $Y2=1.35
r208 39 40 433.287 $w=1.5e-07 $l=8.45e-07 $layer=POLY_cond $X=7.865 $Y=1.65
+ $X2=7.02 $Y2=1.65
r209 36 53 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.945 $Y=1.725
+ $X2=6.945 $Y2=1.65
r210 36 38 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=6.945 $Y=1.725
+ $X2=6.945 $Y2=2.465
r211 35 52 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.59 $Y=1.65
+ $X2=6.515 $Y2=1.65
r212 34 53 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.87 $Y=1.65
+ $X2=6.945 $Y2=1.65
r213 34 35 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=6.87 $Y=1.65
+ $X2=6.59 $Y2=1.65
r214 31 52 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.515 $Y=1.725
+ $X2=6.515 $Y2=1.65
r215 31 33 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=6.515 $Y=1.725
+ $X2=6.515 $Y2=2.465
r216 30 51 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.16 $Y=1.65
+ $X2=6.085 $Y2=1.65
r217 29 52 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.44 $Y=1.65
+ $X2=6.515 $Y2=1.65
r218 29 30 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=6.44 $Y=1.65
+ $X2=6.16 $Y2=1.65
r219 26 51 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.085 $Y=1.725
+ $X2=6.085 $Y2=1.65
r220 26 28 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=6.085 $Y=1.725
+ $X2=6.085 $Y2=2.465
r221 25 50 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.73 $Y=1.65
+ $X2=5.655 $Y2=1.65
r222 24 51 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.01 $Y=1.65
+ $X2=6.085 $Y2=1.65
r223 24 25 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=6.01 $Y=1.65
+ $X2=5.73 $Y2=1.65
r224 21 50 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.655 $Y=1.725
+ $X2=5.655 $Y2=1.65
r225 21 23 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=5.655 $Y=1.725
+ $X2=5.655 $Y2=2.465
r226 20 49 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.3 $Y=1.65
+ $X2=5.225 $Y2=1.65
r227 19 50 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.58 $Y=1.65
+ $X2=5.655 $Y2=1.65
r228 19 20 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=5.58 $Y=1.65
+ $X2=5.3 $Y2=1.65
r229 16 49 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.225 $Y=1.725
+ $X2=5.225 $Y2=1.65
r230 16 18 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=5.225 $Y=1.725
+ $X2=5.225 $Y2=2.465
r231 15 48 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.87 $Y=1.65
+ $X2=4.795 $Y2=1.65
r232 14 49 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.15 $Y=1.65
+ $X2=5.225 $Y2=1.65
r233 14 15 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=5.15 $Y=1.65
+ $X2=4.87 $Y2=1.65
r234 11 48 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.795 $Y=1.725
+ $X2=4.795 $Y2=1.65
r235 11 13 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=4.795 $Y=1.725
+ $X2=4.795 $Y2=2.465
r236 10 47 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.44 $Y=1.65
+ $X2=4.365 $Y2=1.65
r237 9 48 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.72 $Y=1.65
+ $X2=4.795 $Y2=1.65
r238 9 10 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=4.72 $Y=1.65
+ $X2=4.44 $Y2=1.65
r239 6 47 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.365 $Y=1.725
+ $X2=4.365 $Y2=1.65
r240 6 8 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=4.365 $Y=1.725
+ $X2=4.365 $Y2=2.465
r241 4 47 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.29 $Y=1.65
+ $X2=4.365 $Y2=1.65
r242 4 5 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=4.29 $Y=1.65 $X2=4.01
+ $Y2=1.65
r243 1 5 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.935 $Y=1.725
+ $X2=4.01 $Y2=1.65
r244 1 3 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=3.935 $Y=1.725
+ $X2=3.935 $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__EBUFN_8%A 1 3 6 8 10 13 15 22
c39 6 0 1.46525e-19 $X=8.645 $Y=2.465
r40 20 22 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=8.87 $Y=1.35
+ $X2=9.075 $Y2=1.35
r41 17 20 39.3438 $w=3.3e-07 $l=2.25e-07 $layer=POLY_cond $X=8.645 $Y=1.35
+ $X2=8.87 $Y2=1.35
r42 15 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.87
+ $Y=1.35 $X2=8.87 $Y2=1.35
r43 11 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.075 $Y=1.515
+ $X2=9.075 $Y2=1.35
r44 11 13 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=9.075 $Y=1.515
+ $X2=9.075 $Y2=2.465
r45 8 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.075 $Y=1.185
+ $X2=9.075 $Y2=1.35
r46 8 10 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=9.075 $Y=1.185
+ $X2=9.075 $Y2=0.655
r47 4 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.645 $Y=1.515
+ $X2=8.645 $Y2=1.35
r48 4 6 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=8.645 $Y=1.515
+ $X2=8.645 $Y2=2.465
r49 1 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.645 $Y=1.185
+ $X2=8.645 $Y2=1.35
r50 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=8.645 $Y=1.185
+ $X2=8.645 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__EBUFN_8%A_27_367# 1 2 3 4 5 6 7 8 9 28 30 32 36 38
+ 42 44 48 50 52 53 54 58 60 64 66 68 69 72 74 80 81 82 88 90 93 95
c131 74 0 1.85809e-19 $X=6.995 $Y=2.45
c132 68 0 1.57686e-19 $X=6.26 $Y=1.985
c133 52 0 1.61246e-19 $X=3.72 $Y=1.985
r134 75 93 2.76166 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.385 $Y=2.45
+ $X2=6.26 $Y2=2.45
r135 74 95 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.995 $Y=2.45
+ $X2=7.16 $Y2=2.45
r136 74 75 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=6.995 $Y=2.45
+ $X2=6.385 $Y2=2.45
r137 70 93 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.26 $Y=2.535
+ $X2=6.26 $Y2=2.45
r138 70 72 17.2866 $w=2.48e-07 $l=3.75e-07 $layer=LI1_cond $X=6.26 $Y=2.535
+ $X2=6.26 $Y2=2.91
r139 69 93 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.26 $Y=2.365
+ $X2=6.26 $Y2=2.45
r140 68 92 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.26 $Y=1.985
+ $X2=6.26 $Y2=1.9
r141 68 69 17.5171 $w=2.48e-07 $l=3.8e-07 $layer=LI1_cond $X=6.26 $Y=1.985
+ $X2=6.26 $Y2=2.365
r142 67 90 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.605 $Y=1.9
+ $X2=5.44 $Y2=1.9
r143 66 92 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.135 $Y=1.9
+ $X2=6.26 $Y2=1.9
r144 66 67 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=6.135 $Y=1.9
+ $X2=5.605 $Y2=1.9
r145 62 90 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.44 $Y=1.985
+ $X2=5.44 $Y2=1.9
r146 62 64 32.3033 $w=3.28e-07 $l=9.25e-07 $layer=LI1_cond $X=5.44 $Y=1.985
+ $X2=5.44 $Y2=2.91
r147 61 88 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.745 $Y=1.9
+ $X2=4.58 $Y2=1.9
r148 60 90 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.275 $Y=1.9
+ $X2=5.44 $Y2=1.9
r149 60 61 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=5.275 $Y=1.9
+ $X2=4.745 $Y2=1.9
r150 56 88 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.58 $Y=1.985
+ $X2=4.58 $Y2=1.9
r151 56 58 32.3033 $w=3.28e-07 $l=9.25e-07 $layer=LI1_cond $X=4.58 $Y=1.985
+ $X2=4.58 $Y2=2.91
r152 55 84 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.805 $Y=1.9
+ $X2=3.72 $Y2=1.9
r153 54 88 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.415 $Y=1.9
+ $X2=4.58 $Y2=1.9
r154 54 55 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=4.415 $Y=1.9
+ $X2=3.805 $Y2=1.9
r155 53 86 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.72 $Y=2.905
+ $X2=3.72 $Y2=2.99
r156 52 84 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.72 $Y=1.985
+ $X2=3.72 $Y2=1.9
r157 52 53 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=3.72 $Y=1.985
+ $X2=3.72 $Y2=2.905
r158 51 82 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.945 $Y=2.99
+ $X2=2.86 $Y2=2.99
r159 50 86 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.635 $Y=2.99
+ $X2=3.72 $Y2=2.99
r160 50 51 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.635 $Y=2.99
+ $X2=2.945 $Y2=2.99
r161 46 82 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.86 $Y=2.905
+ $X2=2.86 $Y2=2.99
r162 46 48 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=2.86 $Y=2.905
+ $X2=2.86 $Y2=2.32
r163 45 81 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.085 $Y=2.99 $X2=2
+ $Y2=2.99
r164 44 82 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.775 $Y=2.99
+ $X2=2.86 $Y2=2.99
r165 44 45 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.775 $Y=2.99
+ $X2=2.085 $Y2=2.99
r166 40 81 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2 $Y=2.905 $X2=2
+ $Y2=2.99
r167 40 42 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=2 $Y=2.905 $X2=2
+ $Y2=2.32
r168 39 80 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.225 $Y=2.99
+ $X2=1.1 $Y2=2.99
r169 38 81 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.915 $Y=2.99 $X2=2
+ $Y2=2.99
r170 38 39 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.915 $Y=2.99
+ $X2=1.225 $Y2=2.99
r171 34 80 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.1 $Y=2.905
+ $X2=1.1 $Y2=2.99
r172 34 36 26.9672 $w=2.48e-07 $l=5.85e-07 $layer=LI1_cond $X=1.1 $Y=2.905
+ $X2=1.1 $Y2=2.32
r173 33 79 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.445 $Y=2.99
+ $X2=0.28 $Y2=2.99
r174 32 80 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.975 $Y=2.99
+ $X2=1.1 $Y2=2.99
r175 32 33 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=0.975 $Y=2.99
+ $X2=0.445 $Y2=2.99
r176 28 79 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.28 $Y=2.905
+ $X2=0.28 $Y2=2.99
r177 28 30 32.3033 $w=3.28e-07 $l=9.25e-07 $layer=LI1_cond $X=0.28 $Y=2.905
+ $X2=0.28 $Y2=1.98
r178 9 95 300 $w=1.7e-07 $l=7.61791e-07 $layer=licon1_PDIFF $count=2 $X=7.02
+ $Y=1.835 $X2=7.16 $Y2=2.53
r179 8 92 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=6.16
+ $Y=1.835 $X2=6.3 $Y2=1.98
r180 8 72 600 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=6.16
+ $Y=1.835 $X2=6.3 $Y2=2.91
r181 7 90 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=5.3
+ $Y=1.835 $X2=5.44 $Y2=1.98
r182 7 64 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=5.3
+ $Y=1.835 $X2=5.44 $Y2=2.91
r183 6 88 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=4.44
+ $Y=1.835 $X2=4.58 $Y2=1.98
r184 6 58 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=4.44
+ $Y=1.835 $X2=4.58 $Y2=2.91
r185 5 86 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=3.58
+ $Y=1.835 $X2=3.72 $Y2=2.91
r186 5 84 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=3.58
+ $Y=1.835 $X2=3.72 $Y2=1.98
r187 4 48 300 $w=1.7e-07 $l=5.50568e-07 $layer=licon1_PDIFF $count=2 $X=2.72
+ $Y=1.835 $X2=2.86 $Y2=2.32
r188 3 42 300 $w=1.7e-07 $l=5.50568e-07 $layer=licon1_PDIFF $count=2 $X=1.86
+ $Y=1.835 $X2=2 $Y2=2.32
r189 2 36 300 $w=1.7e-07 $l=5.50568e-07 $layer=licon1_PDIFF $count=2 $X=1
+ $Y=1.835 $X2=1.14 $Y2=2.32
r190 1 79 400 $w=1.7e-07 $l=1.14521e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.835 $X2=0.28 $Y2=2.91
r191 1 30 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.835 $X2=0.28 $Y2=1.98
.ends

.subckt PM_SKY130_FD_SC_LP__EBUFN_8%Z 1 2 3 4 5 6 7 8 27 29 30 33 35 39 43 45 49
+ 53 55 59 64 65 67 68 70 72 73 74 77
c136 72 0 5.74299e-20 $X=3.29 $Y=1.98
c137 64 0 2.92592e-19 $X=0.71 $Y=1.98
c138 53 0 5.58653e-20 $X=3.125 $Y=1.06
c139 30 0 1.81636e-19 $X=0.71 $Y=1.815
r140 74 81 9.4 $w=3.05e-07 $l=2.35e-07 $layer=LI1_cond $X=0.71 $Y=1.295 $X2=0.71
+ $Y2=1.06
r141 74 77 2.39218 $w=2.3e-07 $l=1.65e-07 $layer=LI1_cond $X=0.71 $Y=1.295
+ $X2=0.545 $Y2=1.295
r142 73 77 15.2824 $w=2.28e-07 $l=3.05e-07 $layer=LI1_cond $X=0.24 $Y=1.295
+ $X2=0.545 $Y2=1.295
r143 57 59 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=3.29 $Y=0.975
+ $X2=3.29 $Y2=0.805
r144 56 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.595 $Y=1.9
+ $X2=2.43 $Y2=1.9
r145 55 72 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.125 $Y=1.9
+ $X2=3.29 $Y2=1.9
r146 55 56 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=3.125 $Y=1.9
+ $X2=2.595 $Y2=1.9
r147 54 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.595 $Y=1.06
+ $X2=2.43 $Y2=1.06
r148 53 57 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.125 $Y=1.06
+ $X2=3.29 $Y2=0.975
r149 53 54 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=3.125 $Y=1.06
+ $X2=2.595 $Y2=1.06
r150 47 68 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.43 $Y=0.975
+ $X2=2.43 $Y2=1.06
r151 47 49 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=2.43 $Y=0.975
+ $X2=2.43 $Y2=0.805
r152 46 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.735 $Y=1.9
+ $X2=1.57 $Y2=1.9
r153 45 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.265 $Y=1.9
+ $X2=2.43 $Y2=1.9
r154 45 46 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=2.265 $Y=1.9
+ $X2=1.735 $Y2=1.9
r155 44 65 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.735 $Y=1.06
+ $X2=1.57 $Y2=1.06
r156 43 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.265 $Y=1.06
+ $X2=2.43 $Y2=1.06
r157 43 44 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=2.265 $Y=1.06
+ $X2=1.735 $Y2=1.06
r158 37 65 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.57 $Y=0.975
+ $X2=1.57 $Y2=1.06
r159 37 39 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=1.57 $Y=0.975
+ $X2=1.57 $Y2=0.805
r160 36 81 4.15824 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.875 $Y=1.06
+ $X2=0.71 $Y2=1.06
r161 35 65 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.405 $Y=1.06
+ $X2=1.57 $Y2=1.06
r162 35 36 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=1.405 $Y=1.06
+ $X2=0.875 $Y2=1.06
r163 34 64 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.795 $Y=1.9
+ $X2=0.71 $Y2=1.9
r164 33 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.405 $Y=1.9
+ $X2=1.57 $Y2=1.9
r165 33 34 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=1.405 $Y=1.9
+ $X2=0.795 $Y2=1.9
r166 30 64 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.71 $Y=1.815
+ $X2=0.71 $Y2=1.9
r167 29 74 6.97136 $w=3.05e-07 $l=1.15e-07 $layer=LI1_cond $X=0.71 $Y=1.41
+ $X2=0.71 $Y2=1.295
r168 29 30 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=0.71 $Y=1.41
+ $X2=0.71 $Y2=1.815
r169 25 81 3.23248 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.71 $Y=0.975
+ $X2=0.71 $Y2=1.06
r170 25 27 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=0.71 $Y=0.975
+ $X2=0.71 $Y2=0.805
r171 8 72 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=3.15
+ $Y=1.835 $X2=3.29 $Y2=1.98
r172 7 70 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=2.29
+ $Y=1.835 $X2=2.43 $Y2=1.98
r173 6 67 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=1.43
+ $Y=1.835 $X2=1.57 $Y2=1.98
r174 5 64 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=0.57
+ $Y=1.835 $X2=0.71 $Y2=1.98
r175 4 59 182 $w=1.7e-07 $l=6.3616e-07 $layer=licon1_NDIFF $count=1 $X=3.15
+ $Y=0.235 $X2=3.29 $Y2=0.805
r176 3 49 182 $w=1.7e-07 $l=6.3616e-07 $layer=licon1_NDIFF $count=1 $X=2.29
+ $Y=0.235 $X2=2.43 $Y2=0.805
r177 2 39 182 $w=1.7e-07 $l=6.3616e-07 $layer=licon1_NDIFF $count=1 $X=1.43
+ $Y=0.235 $X2=1.57 $Y2=0.805
r178 1 27 182 $w=1.7e-07 $l=6.3616e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.235 $X2=0.71 $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_LP__EBUFN_8%VPWR 1 2 3 4 5 6 21 25 29 33 37 39 41 46 47
+ 49 50 52 53 54 56 74 81 87 90 94
r134 93 94 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r135 90 91 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=3.33 $X2=8.4
+ $Y2=3.33
r136 87 88 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r137 85 94 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=9.36 $Y2=3.33
r138 85 91 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=8.4 $Y2=3.33
r139 84 85 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r140 82 90 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.515 $Y=3.33
+ $X2=8.39 $Y2=3.33
r141 82 84 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=8.515 $Y=3.33
+ $X2=8.88 $Y2=3.33
r142 81 93 3.97515 $w=1.7e-07 $l=1.97e-07 $layer=LI1_cond $X=9.205 $Y=3.33
+ $X2=9.402 $Y2=3.33
r143 81 84 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=9.205 $Y=3.33
+ $X2=8.88 $Y2=3.33
r144 80 91 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=8.4 $Y2=3.33
r145 79 80 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r146 77 80 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=7.92 $Y2=3.33
r147 76 79 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=6.96 $Y=3.33
+ $X2=7.92 $Y2=3.33
r148 76 77 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r149 74 90 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.265 $Y=3.33
+ $X2=8.39 $Y2=3.33
r150 74 79 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=8.265 $Y=3.33
+ $X2=7.92 $Y2=3.33
r151 73 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=6.96 $Y2=3.33
r152 72 73 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r153 70 73 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=6.48 $Y2=3.33
r154 69 70 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r155 67 88 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=4.08 $Y2=3.33
r156 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r157 64 87 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.235 $Y=3.33
+ $X2=4.11 $Y2=3.33
r158 64 66 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=4.235 $Y=3.33
+ $X2=4.56 $Y2=3.33
r159 63 88 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r160 62 63 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r161 59 63 0.936549 $w=4.9e-07 $l=3.36e-06 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=3.6 $Y2=3.33
r162 58 62 219.209 $w=1.68e-07 $l=3.36e-06 $layer=LI1_cond $X=0.24 $Y=3.33
+ $X2=3.6 $Y2=3.33
r163 58 59 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r164 56 87 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.985 $Y=3.33
+ $X2=4.11 $Y2=3.33
r165 56 62 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=3.985 $Y=3.33
+ $X2=3.6 $Y2=3.33
r166 54 70 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=4.8 $Y=3.33
+ $X2=5.52 $Y2=3.33
r167 54 67 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.8 $Y=3.33
+ $X2=4.56 $Y2=3.33
r168 52 72 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=6.565 $Y=3.33
+ $X2=6.48 $Y2=3.33
r169 52 53 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.565 $Y=3.33
+ $X2=6.69 $Y2=3.33
r170 51 76 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=6.815 $Y=3.33
+ $X2=6.96 $Y2=3.33
r171 51 53 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.815 $Y=3.33
+ $X2=6.69 $Y2=3.33
r172 49 69 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=5.785 $Y=3.33
+ $X2=5.52 $Y2=3.33
r173 49 50 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.785 $Y=3.33
+ $X2=5.87 $Y2=3.33
r174 48 72 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=5.955 $Y=3.33
+ $X2=6.48 $Y2=3.33
r175 48 50 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.955 $Y=3.33
+ $X2=5.87 $Y2=3.33
r176 46 66 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=4.925 $Y=3.33
+ $X2=4.56 $Y2=3.33
r177 46 47 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.925 $Y=3.33
+ $X2=5.01 $Y2=3.33
r178 45 69 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=5.095 $Y=3.33
+ $X2=5.52 $Y2=3.33
r179 45 47 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.095 $Y=3.33
+ $X2=5.01 $Y2=3.33
r180 41 44 44.7148 $w=2.48e-07 $l=9.7e-07 $layer=LI1_cond $X=9.33 $Y=1.98
+ $X2=9.33 $Y2=2.95
r181 39 93 3.16801 $w=2.5e-07 $l=1.15521e-07 $layer=LI1_cond $X=9.33 $Y=3.245
+ $X2=9.402 $Y2=3.33
r182 39 44 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=9.33 $Y=3.245
+ $X2=9.33 $Y2=2.95
r183 35 90 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=8.39 $Y=3.245
+ $X2=8.39 $Y2=3.33
r184 35 37 16.5952 $w=2.48e-07 $l=3.6e-07 $layer=LI1_cond $X=8.39 $Y=3.245
+ $X2=8.39 $Y2=2.885
r185 31 53 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.69 $Y=3.245
+ $X2=6.69 $Y2=3.33
r186 31 33 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=6.69 $Y=3.245
+ $X2=6.69 $Y2=2.91
r187 27 50 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.87 $Y=3.245
+ $X2=5.87 $Y2=3.33
r188 27 29 60.3476 $w=1.68e-07 $l=9.25e-07 $layer=LI1_cond $X=5.87 $Y=3.245
+ $X2=5.87 $Y2=2.32
r189 23 47 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.01 $Y=3.245
+ $X2=5.01 $Y2=3.33
r190 23 25 60.3476 $w=1.68e-07 $l=9.25e-07 $layer=LI1_cond $X=5.01 $Y=3.245
+ $X2=5.01 $Y2=2.32
r191 19 87 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.11 $Y=3.245
+ $X2=4.11 $Y2=3.33
r192 19 21 42.6404 $w=2.48e-07 $l=9.25e-07 $layer=LI1_cond $X=4.11 $Y=3.245
+ $X2=4.11 $Y2=2.32
r193 6 44 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=9.15
+ $Y=1.835 $X2=9.29 $Y2=2.95
r194 6 41 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=9.15
+ $Y=1.835 $X2=9.29 $Y2=1.98
r195 5 37 600 $w=1.7e-07 $l=1.11781e-06 $layer=licon1_PDIFF $count=1 $X=8.29
+ $Y=1.835 $X2=8.43 $Y2=2.885
r196 4 33 600 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=6.59
+ $Y=1.835 $X2=6.73 $Y2=2.91
r197 3 29 300 $w=1.7e-07 $l=5.50568e-07 $layer=licon1_PDIFF $count=2 $X=5.73
+ $Y=1.835 $X2=5.87 $Y2=2.32
r198 2 25 300 $w=1.7e-07 $l=5.50568e-07 $layer=licon1_PDIFF $count=2 $X=4.87
+ $Y=1.835 $X2=5.01 $Y2=2.32
r199 1 21 300 $w=1.7e-07 $l=5.50568e-07 $layer=licon1_PDIFF $count=2 $X=4.01
+ $Y=1.835 $X2=4.15 $Y2=2.32
.ends

.subckt PM_SKY130_FD_SC_LP__EBUFN_8%A_27_47# 1 2 3 4 5 6 7 8 9 30 34 36 40 42 46
+ 48 50 51 52 53 56 58 62 64 68 70 74 77 78 79 80 83 84 85
r152 72 74 32.9599 $w=2.48e-07 $l=7.15e-07 $layer=LI1_cond $X=7.12 $Y=1.135
+ $X2=7.12 $Y2=0.42
r153 71 85 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.465 $Y=1.22
+ $X2=6.3 $Y2=1.22
r154 70 72 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=6.995 $Y=1.22
+ $X2=7.12 $Y2=1.135
r155 70 71 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=6.995 $Y=1.22
+ $X2=6.465 $Y2=1.22
r156 66 85 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.3 $Y=1.135 $X2=6.3
+ $Y2=1.22
r157 66 68 24.9696 $w=3.28e-07 $l=7.15e-07 $layer=LI1_cond $X=6.3 $Y=1.135
+ $X2=6.3 $Y2=0.42
r158 65 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.605 $Y=1.22
+ $X2=5.44 $Y2=1.22
r159 64 85 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.135 $Y=1.22
+ $X2=6.3 $Y2=1.22
r160 64 65 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=6.135 $Y=1.22
+ $X2=5.605 $Y2=1.22
r161 60 84 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.44 $Y=1.135
+ $X2=5.44 $Y2=1.22
r162 60 62 26.3665 $w=3.28e-07 $l=7.55e-07 $layer=LI1_cond $X=5.44 $Y=1.135
+ $X2=5.44 $Y2=0.38
r163 59 83 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.745 $Y=1.22
+ $X2=4.58 $Y2=1.22
r164 58 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.275 $Y=1.22
+ $X2=5.44 $Y2=1.22
r165 58 59 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=5.275 $Y=1.22
+ $X2=4.745 $Y2=1.22
r166 54 83 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.58 $Y=1.135
+ $X2=4.58 $Y2=1.22
r167 54 56 24.9696 $w=3.28e-07 $l=7.15e-07 $layer=LI1_cond $X=4.58 $Y=1.135
+ $X2=4.58 $Y2=0.42
r168 52 83 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.415 $Y=1.22
+ $X2=4.58 $Y2=1.22
r169 52 53 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=4.415 $Y=1.22
+ $X2=3.805 $Y2=1.22
r170 51 53 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.72 $Y=1.135
+ $X2=3.805 $Y2=1.22
r171 50 82 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.72 $Y=0.425
+ $X2=3.72 $Y2=0.34
r172 50 51 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=3.72 $Y=0.425
+ $X2=3.72 $Y2=1.135
r173 49 80 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.945 $Y=0.34
+ $X2=2.86 $Y2=0.34
r174 48 82 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.635 $Y=0.34
+ $X2=3.72 $Y2=0.34
r175 48 49 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.635 $Y=0.34
+ $X2=2.945 $Y2=0.34
r176 44 80 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.86 $Y=0.425
+ $X2=2.86 $Y2=0.34
r177 44 46 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=2.86 $Y=0.425
+ $X2=2.86 $Y2=0.53
r178 43 79 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.085 $Y=0.34 $X2=2
+ $Y2=0.34
r179 42 80 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.775 $Y=0.34
+ $X2=2.86 $Y2=0.34
r180 42 43 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.775 $Y=0.34
+ $X2=2.085 $Y2=0.34
r181 38 79 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2 $Y=0.425 $X2=2
+ $Y2=0.34
r182 38 40 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=2 $Y=0.425 $X2=2
+ $Y2=0.53
r183 37 78 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.225 $Y=0.34
+ $X2=1.14 $Y2=0.34
r184 36 79 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.915 $Y=0.34 $X2=2
+ $Y2=0.34
r185 36 37 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.915 $Y=0.34
+ $X2=1.225 $Y2=0.34
r186 32 78 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.14 $Y=0.425
+ $X2=1.14 $Y2=0.34
r187 32 34 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=1.14 $Y=0.425
+ $X2=1.14 $Y2=0.53
r188 31 77 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.365 $Y=0.34
+ $X2=0.24 $Y2=0.34
r189 30 78 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.055 $Y=0.34
+ $X2=1.14 $Y2=0.34
r190 30 31 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.055 $Y=0.34
+ $X2=0.365 $Y2=0.34
r191 9 74 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=7.02
+ $Y=0.235 $X2=7.16 $Y2=0.42
r192 8 68 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=6.16
+ $Y=0.235 $X2=6.3 $Y2=0.42
r193 7 62 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.3
+ $Y=0.235 $X2=5.44 $Y2=0.38
r194 6 56 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=4.44
+ $Y=0.235 $X2=4.58 $Y2=0.42
r195 5 82 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=3.58
+ $Y=0.235 $X2=3.72 $Y2=0.42
r196 4 46 182 $w=1.7e-07 $l=3.58225e-07 $layer=licon1_NDIFF $count=1 $X=2.72
+ $Y=0.235 $X2=2.86 $Y2=0.53
r197 3 40 182 $w=1.7e-07 $l=3.58225e-07 $layer=licon1_NDIFF $count=1 $X=1.86
+ $Y=0.235 $X2=2 $Y2=0.53
r198 2 34 182 $w=1.7e-07 $l=3.58225e-07 $layer=licon1_NDIFF $count=1 $X=1
+ $Y=0.235 $X2=1.14 $Y2=0.53
r199 1 77 91 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.28 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__EBUFN_8%VGND 1 2 3 4 5 6 21 25 29 33 37 39 41 44 45
+ 47 48 50 51 52 54 72 76 82 85 89
c128 89 0 3.60707e-20 $X=9.36 $Y=0
r129 88 89 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=0 $X2=9.36
+ $Y2=0
r130 85 86 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r131 82 83 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r132 80 89 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=0 $X2=9.36
+ $Y2=0
r133 80 86 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=0 $X2=8.4
+ $Y2=0
r134 79 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=0 $X2=8.88
+ $Y2=0
r135 77 85 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.515 $Y=0 $X2=8.43
+ $Y2=0
r136 77 79 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=8.515 $Y=0
+ $X2=8.88 $Y2=0
r137 76 88 3.97515 $w=1.7e-07 $l=1.97e-07 $layer=LI1_cond $X=9.205 $Y=0
+ $X2=9.402 $Y2=0
r138 76 79 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=9.205 $Y=0
+ $X2=8.88 $Y2=0
r139 75 86 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=6.96 $Y=0 $X2=8.4
+ $Y2=0
r140 74 75 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r141 72 85 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.345 $Y=0 $X2=8.43
+ $Y2=0
r142 72 74 90.3583 $w=1.68e-07 $l=1.385e-06 $layer=LI1_cond $X=8.345 $Y=0
+ $X2=6.96 $Y2=0
r143 71 75 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6.96
+ $Y2=0
r144 70 71 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r145 68 71 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=6.48
+ $Y2=0
r146 67 68 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r147 65 83 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=4.08
+ $Y2=0
r148 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r149 62 82 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.235 $Y=0 $X2=4.11
+ $Y2=0
r150 62 64 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=4.235 $Y=0
+ $X2=4.56 $Y2=0
r151 61 83 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r152 60 61 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r153 57 61 0.936549 $w=4.9e-07 $l=3.36e-06 $layer=MET1_cond $X=0.24 $Y=0 $X2=3.6
+ $Y2=0
r154 56 60 219.209 $w=1.68e-07 $l=3.36e-06 $layer=LI1_cond $X=0.24 $Y=0 $X2=3.6
+ $Y2=0
r155 56 57 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=0.24 $Y=0
+ $X2=0.24 $Y2=0
r156 54 82 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.985 $Y=0 $X2=4.11
+ $Y2=0
r157 54 60 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=3.985 $Y=0 $X2=3.6
+ $Y2=0
r158 52 68 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=4.8 $Y=0 $X2=5.52
+ $Y2=0
r159 52 65 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.8 $Y=0 $X2=4.56
+ $Y2=0
r160 50 70 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=6.645 $Y=0
+ $X2=6.48 $Y2=0
r161 50 51 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.645 $Y=0 $X2=6.73
+ $Y2=0
r162 49 74 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=6.815 $Y=0
+ $X2=6.96 $Y2=0
r163 49 51 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.815 $Y=0 $X2=6.73
+ $Y2=0
r164 47 67 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=5.785 $Y=0
+ $X2=5.52 $Y2=0
r165 47 48 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.785 $Y=0 $X2=5.87
+ $Y2=0
r166 46 70 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=5.955 $Y=0
+ $X2=6.48 $Y2=0
r167 46 48 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.955 $Y=0 $X2=5.87
+ $Y2=0
r168 44 64 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=4.925 $Y=0
+ $X2=4.56 $Y2=0
r169 44 45 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.925 $Y=0 $X2=5.01
+ $Y2=0
r170 43 67 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=5.095 $Y=0
+ $X2=5.52 $Y2=0
r171 43 45 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.095 $Y=0 $X2=5.01
+ $Y2=0
r172 39 88 3.16801 $w=2.5e-07 $l=1.15521e-07 $layer=LI1_cond $X=9.33 $Y=0.085
+ $X2=9.402 $Y2=0
r173 39 41 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=9.33 $Y=0.085
+ $X2=9.33 $Y2=0.38
r174 35 85 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.43 $Y=0.085
+ $X2=8.43 $Y2=0
r175 35 37 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=8.43 $Y=0.085
+ $X2=8.43 $Y2=0.44
r176 31 51 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.73 $Y=0.085
+ $X2=6.73 $Y2=0
r177 31 33 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=6.73 $Y=0.085
+ $X2=6.73 $Y2=0.38
r178 27 48 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.87 $Y=0.085
+ $X2=5.87 $Y2=0
r179 27 29 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=5.87 $Y=0.085
+ $X2=5.87 $Y2=0.38
r180 23 45 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.01 $Y=0.085
+ $X2=5.01 $Y2=0
r181 23 25 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=5.01 $Y=0.085
+ $X2=5.01 $Y2=0.38
r182 19 82 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.11 $Y=0.085
+ $X2=4.11 $Y2=0
r183 19 21 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=4.11 $Y=0.085
+ $X2=4.11 $Y2=0.38
r184 6 41 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=9.15
+ $Y=0.235 $X2=9.29 $Y2=0.38
r185 5 37 182 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_NDIFF $count=1 $X=8.29
+ $Y=0.235 $X2=8.43 $Y2=0.44
r186 4 33 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.59
+ $Y=0.235 $X2=6.73 $Y2=0.38
r187 3 29 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.73
+ $Y=0.235 $X2=5.87 $Y2=0.38
r188 2 25 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.87
+ $Y=0.235 $X2=5.01 $Y2=0.38
r189 1 21 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.01
+ $Y=0.235 $X2=4.15 $Y2=0.38
.ends

