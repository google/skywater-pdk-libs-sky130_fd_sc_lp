* File: sky130_fd_sc_lp__or2_2.spice
* Created: Fri Aug 28 11:21:28 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__or2_2.pex.spice"
.subckt sky130_fd_sc_lp__or2_2  VNB VPB B A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* B	B
* VPB	VPB
* VNB	VNB
MM1004 N_A_48_390#_M1004_d N_B_M1004_g N_VGND_M1004_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75001.6
+ A=0.063 P=1.14 MULT=1
MM1003 N_VGND_M1003_d N_A_M1003_g N_A_48_390#_M1004_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0896 AS=0.0588 PD=0.81 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1002 N_VGND_M1003_d N_A_48_390#_M1002_g N_X_M1002_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1792 AS=0.1176 PD=1.62 PS=1.12 NRD=6.42 NRS=0 M=1 R=5.6 SA=75000.7
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1007 N_VGND_M1007_d N_A_48_390#_M1007_g N_X_M1002_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.1
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1000 A_131_390# N_B_M1000_g N_A_48_390#_M1000_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0441 AS=0.1113 PD=0.63 PS=1.37 NRD=23.443 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.5 A=0.063 P=1.14 MULT=1
MM1006 N_VPWR_M1006_d N_A_M1006_g A_131_390# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.095025 AS=0.0441 PD=0.8175 PS=0.63 NRD=0 NRS=23.443 M=1 R=2.8 SA=75000.6
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1001 N_VPWR_M1006_d N_A_48_390#_M1001_g N_X_M1001_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.285075 AS=0.1764 PD=2.4525 PS=1.54 NRD=4.9447 NRS=0 M=1 R=8.4 SA=75000.5
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1005 N_VPWR_M1005_d N_A_48_390#_M1005_g N_X_M1001_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.9
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX8_noxref VNB VPB NWDIODE A=5.1847 P=9.29
*
.include "sky130_fd_sc_lp__or2_2.pxi.spice"
*
.ends
*
*
