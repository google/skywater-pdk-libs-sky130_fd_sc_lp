* File: sky130_fd_sc_lp__o2111a_m.pex.spice
* Created: Fri Aug 28 11:00:30 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O2111A_M%A_80_21# 1 2 3 12 14 17 19 23 24 25 26 27
+ 28 31 35 37 41 43 45
c92 24 0 1.12474e-19 $X=0.63 $Y=0.93
r93 39 41 11.355 $w=2.08e-07 $l=2.15e-07 $layer=LI1_cond $X=2.53 $Y=2.605
+ $X2=2.53 $Y2=2.82
r94 38 43 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.51 $Y=2.52
+ $X2=1.405 $Y2=2.52
r95 37 39 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=2.425 $Y=2.52
+ $X2=2.53 $Y2=2.605
r96 37 38 59.6952 $w=1.68e-07 $l=9.15e-07 $layer=LI1_cond $X=2.425 $Y=2.52
+ $X2=1.51 $Y2=2.52
r97 33 43 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=1.405 $Y=2.605
+ $X2=1.405 $Y2=2.52
r98 33 35 11.355 $w=2.08e-07 $l=2.15e-07 $layer=LI1_cond $X=1.405 $Y=2.605
+ $X2=1.405 $Y2=2.82
r99 29 31 11.355 $w=2.08e-07 $l=2.15e-07 $layer=LI1_cond $X=1.215 $Y=0.725
+ $X2=1.215 $Y2=0.51
r100 27 43 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.3 $Y=2.52
+ $X2=1.405 $Y2=2.52
r101 27 28 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=1.3 $Y=2.52
+ $X2=0.715 $Y2=2.52
r102 25 29 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=1.11 $Y=0.81
+ $X2=1.215 $Y2=0.725
r103 25 26 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=1.11 $Y=0.81
+ $X2=0.715 $Y2=0.81
r104 24 45 45.5639 $w=3.95e-07 $l=1.65e-07 $layer=POLY_cond $X=0.597 $Y=0.93
+ $X2=0.597 $Y2=0.765
r105 23 24 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.63
+ $Y=0.93 $X2=0.63 $Y2=0.93
r106 21 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.63 $Y=2.435
+ $X2=0.715 $Y2=2.52
r107 21 23 98.1872 $w=1.68e-07 $l=1.505e-06 $layer=LI1_cond $X=0.63 $Y=2.435
+ $X2=0.63 $Y2=0.93
r108 20 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.63 $Y=0.895
+ $X2=0.715 $Y2=0.81
r109 20 23 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=0.63 $Y=0.895
+ $X2=0.63 $Y2=0.93
r110 17 19 743.511 $w=1.5e-07 $l=1.45e-06 $layer=POLY_cond $X=0.72 $Y=2.885
+ $X2=0.72 $Y2=1.435
r111 14 19 50.0695 $w=3.95e-07 $l=1.97e-07 $layer=POLY_cond $X=0.597 $Y=1.238
+ $X2=0.597 $Y2=1.435
r112 13 24 4.50555 $w=3.95e-07 $l=3.2e-08 $layer=POLY_cond $X=0.597 $Y=0.962
+ $X2=0.597 $Y2=0.93
r113 13 14 38.8604 $w=3.95e-07 $l=2.76e-07 $layer=POLY_cond $X=0.597 $Y=0.962
+ $X2=0.597 $Y2=1.238
r114 12 45 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.475 $Y=0.445
+ $X2=0.475 $Y2=0.765
r115 3 41 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.39
+ $Y=2.675 $X2=2.53 $Y2=2.82
r116 2 35 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.265
+ $Y=2.675 $X2=1.405 $Y2=2.82
r117 1 31 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=1.09
+ $Y=0.235 $X2=1.215 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_LP__O2111A_M%D1 3 7 8 9 11 13 14 15 16 17 18 23
c55 7 0 7.19238e-20 $X=1.59 $Y=0.84
r56 17 18 20.5182 $w=1.98e-07 $l=3.7e-07 $layer=LI1_cond $X=1.185 $Y=1.665
+ $X2=1.185 $Y2=2.035
r57 16 17 20.5182 $w=1.98e-07 $l=3.7e-07 $layer=LI1_cond $X=1.185 $Y=1.295
+ $X2=1.185 $Y2=1.665
r58 16 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.17
+ $Y=1.375 $X2=1.17 $Y2=1.375
r59 14 23 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.17 $Y=1.715
+ $X2=1.17 $Y2=1.375
r60 14 15 38.6168 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.17 $Y=1.715
+ $X2=1.17 $Y2=1.88
r61 13 23 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.17 $Y=1.21
+ $X2=1.17 $Y2=1.375
r62 9 11 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.665 $Y=0.765
+ $X2=1.665 $Y2=0.445
r63 7 9 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.59 $Y=0.84
+ $X2=1.665 $Y2=0.765
r64 7 8 130.755 $w=1.5e-07 $l=2.55e-07 $layer=POLY_cond $X=1.59 $Y=0.84
+ $X2=1.335 $Y2=0.84
r65 5 8 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.26 $Y=0.915
+ $X2=1.335 $Y2=0.84
r66 5 13 151.266 $w=1.5e-07 $l=2.95e-07 $layer=POLY_cond $X=1.26 $Y=0.915
+ $X2=1.26 $Y2=1.21
r67 3 15 515.33 $w=1.5e-07 $l=1.005e-06 $layer=POLY_cond $X=1.19 $Y=2.885
+ $X2=1.19 $Y2=1.88
.ends

.subckt PM_SKY130_FD_SC_LP__O2111A_M%C1 3 7 12 15 16 17 18 19 25
c48 25 0 1.4009e-19 $X=1.71 $Y=1.32
r49 18 19 20.5182 $w=1.98e-07 $l=3.7e-07 $layer=LI1_cond $X=1.695 $Y=1.665
+ $X2=1.695 $Y2=2.035
r50 17 18 20.5182 $w=1.98e-07 $l=3.7e-07 $layer=LI1_cond $X=1.695 $Y=1.295
+ $X2=1.695 $Y2=1.665
r51 17 25 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.71
+ $Y=1.32 $X2=1.71 $Y2=1.32
r52 16 17 20.5182 $w=1.98e-07 $l=3.7e-07 $layer=LI1_cond $X=1.695 $Y=0.925
+ $X2=1.695 $Y2=1.295
r53 14 25 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.71 $Y=1.66
+ $X2=1.71 $Y2=1.32
r54 14 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.71 $Y=1.66
+ $X2=1.71 $Y2=1.825
r55 10 25 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=1.71 $Y=1.305
+ $X2=1.71 $Y2=1.32
r56 10 12 161.521 $w=1.5e-07 $l=3.15e-07 $layer=POLY_cond $X=1.71 $Y=1.23
+ $X2=2.025 $Y2=1.23
r57 5 12 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.025 $Y=1.155
+ $X2=2.025 $Y2=1.23
r58 5 7 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=2.025 $Y=1.155
+ $X2=2.025 $Y2=0.445
r59 3 15 543.532 $w=1.5e-07 $l=1.06e-06 $layer=POLY_cond $X=1.62 $Y=2.885
+ $X2=1.62 $Y2=1.825
.ends

.subckt PM_SKY130_FD_SC_LP__O2111A_M%B1 2 5 9 11 12 13 14 15 21
c47 12 0 7.19238e-20 $X=2.16 $Y=0.925
r48 21 23 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=2.272 $Y=1.71
+ $X2=2.272 $Y2=1.545
r49 21 22 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.25
+ $Y=1.71 $X2=2.25 $Y2=1.71
r50 15 22 14.4055 $w=2.58e-07 $l=3.25e-07 $layer=LI1_cond $X=2.205 $Y=2.035
+ $X2=2.205 $Y2=1.71
r51 14 22 1.99461 $w=2.58e-07 $l=4.5e-08 $layer=LI1_cond $X=2.205 $Y=1.665
+ $X2=2.205 $Y2=1.71
r52 13 14 16.4002 $w=2.58e-07 $l=3.7e-07 $layer=LI1_cond $X=2.205 $Y=1.295
+ $X2=2.205 $Y2=1.665
r53 12 13 16.4002 $w=2.58e-07 $l=3.7e-07 $layer=LI1_cond $X=2.205 $Y=0.925
+ $X2=2.205 $Y2=1.295
r54 9 23 564.043 $w=1.5e-07 $l=1.1e-06 $layer=POLY_cond $X=2.385 $Y=0.445
+ $X2=2.385 $Y2=1.545
r55 5 11 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=2.315 $Y=2.885
+ $X2=2.315 $Y2=2.215
r56 2 11 40.5548 $w=3.75e-07 $l=1.87e-07 $layer=POLY_cond $X=2.272 $Y=2.028
+ $X2=2.272 $Y2=2.215
r57 1 21 3.26277 $w=3.75e-07 $l=2.2e-08 $layer=POLY_cond $X=2.272 $Y=1.732
+ $X2=2.272 $Y2=1.71
r58 1 2 43.8991 $w=3.75e-07 $l=2.96e-07 $layer=POLY_cond $X=2.272 $Y=1.732
+ $X2=2.272 $Y2=2.028
.ends

.subckt PM_SKY130_FD_SC_LP__O2111A_M%A2 3 7 11 12 13 14 15 20
r45 20 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.835
+ $Y=1.375 $X2=2.835 $Y2=1.375
r46 14 15 11.6823 $w=3.63e-07 $l=3.7e-07 $layer=LI1_cond $X=2.737 $Y=1.665
+ $X2=2.737 $Y2=2.035
r47 14 21 9.1564 $w=3.63e-07 $l=2.9e-07 $layer=LI1_cond $X=2.737 $Y=1.665
+ $X2=2.737 $Y2=1.375
r48 13 21 2.5259 $w=3.63e-07 $l=8e-08 $layer=LI1_cond $X=2.737 $Y=1.295
+ $X2=2.737 $Y2=1.375
r49 11 20 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.835 $Y=1.715
+ $X2=2.835 $Y2=1.375
r50 11 12 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.835 $Y=1.715
+ $X2=2.835 $Y2=1.88
r51 10 20 38.6168 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.835 $Y=1.21
+ $X2=2.835 $Y2=1.375
r52 7 10 392.266 $w=1.5e-07 $l=7.65e-07 $layer=POLY_cond $X=2.815 $Y=0.445
+ $X2=2.815 $Y2=1.21
r53 3 12 515.33 $w=1.5e-07 $l=1.005e-06 $layer=POLY_cond $X=2.745 $Y=2.885
+ $X2=2.745 $Y2=1.88
.ends

.subckt PM_SKY130_FD_SC_LP__O2111A_M%A1 3 7 14 18 21 22 23 24 25 31
c33 18 0 2.58839e-20 $X=3.365 $Y=0.895
r34 31 32 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.455
+ $Y=1.765 $X2=3.455 $Y2=1.765
r35 24 25 13.5366 $w=3.13e-07 $l=3.7e-07 $layer=LI1_cond $X=3.527 $Y=2.035
+ $X2=3.527 $Y2=2.405
r36 24 32 9.87808 $w=3.13e-07 $l=2.7e-07 $layer=LI1_cond $X=3.527 $Y=2.035
+ $X2=3.527 $Y2=1.765
r37 23 32 3.65855 $w=3.13e-07 $l=1e-07 $layer=LI1_cond $X=3.527 $Y=1.665
+ $X2=3.527 $Y2=1.765
r38 22 23 13.5366 $w=3.13e-07 $l=3.7e-07 $layer=LI1_cond $X=3.527 $Y=1.295
+ $X2=3.527 $Y2=1.665
r39 21 31 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.455 $Y=1.6
+ $X2=3.455 $Y2=1.765
r40 16 18 61.5319 $w=1.5e-07 $l=1.2e-07 $layer=POLY_cond $X=3.245 $Y=0.895
+ $X2=3.365 $Y2=0.895
r41 14 31 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=3.455 $Y=2.12
+ $X2=3.455 $Y2=1.765
r42 11 14 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=3.105 $Y=2.195
+ $X2=3.455 $Y2=2.195
r43 9 18 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.365 $Y=0.97
+ $X2=3.365 $Y2=0.895
r44 9 21 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=3.365 $Y=0.97
+ $X2=3.365 $Y2=1.6
r45 5 16 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.245 $Y=0.82
+ $X2=3.245 $Y2=0.895
r46 5 7 192.287 $w=1.5e-07 $l=3.75e-07 $layer=POLY_cond $X=3.245 $Y=0.82
+ $X2=3.245 $Y2=0.445
r47 1 11 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.105 $Y=2.27
+ $X2=3.105 $Y2=2.195
r48 1 3 315.351 $w=1.5e-07 $l=6.15e-07 $layer=POLY_cond $X=3.105 $Y=2.27
+ $X2=3.105 $Y2=2.885
.ends

.subckt PM_SKY130_FD_SC_LP__O2111A_M%X 1 2 9 11 12 13 14 15 16 17 26 28 44
r19 26 44 0.528139 $w=2.08e-07 $l=1e-08 $layer=LI1_cond $X=0.26 $Y=2.785
+ $X2=0.26 $Y2=2.775
r20 17 26 3.40825 $w=2.1e-07 $l=1.05e-07 $layer=LI1_cond $X=0.26 $Y=2.89
+ $X2=0.26 $Y2=2.785
r21 17 44 2.00693 $w=2.08e-07 $l=3.8e-08 $layer=LI1_cond $X=0.26 $Y=2.737
+ $X2=0.26 $Y2=2.775
r22 16 17 17.5342 $w=2.08e-07 $l=3.32e-07 $layer=LI1_cond $X=0.26 $Y=2.405
+ $X2=0.26 $Y2=2.737
r23 15 16 19.5411 $w=2.08e-07 $l=3.7e-07 $layer=LI1_cond $X=0.26 $Y=2.035
+ $X2=0.26 $Y2=2.405
r24 14 15 19.5411 $w=2.08e-07 $l=3.7e-07 $layer=LI1_cond $X=0.26 $Y=1.665
+ $X2=0.26 $Y2=2.035
r25 13 14 19.5411 $w=2.08e-07 $l=3.7e-07 $layer=LI1_cond $X=0.26 $Y=1.295
+ $X2=0.26 $Y2=1.665
r26 12 13 19.5411 $w=2.08e-07 $l=3.7e-07 $layer=LI1_cond $X=0.26 $Y=0.925
+ $X2=0.26 $Y2=1.295
r27 11 12 19.5411 $w=2.08e-07 $l=3.7e-07 $layer=LI1_cond $X=0.26 $Y=0.555
+ $X2=0.26 $Y2=0.925
r28 11 28 6.60173 $w=2.08e-07 $l=1.25e-07 $layer=LI1_cond $X=0.26 $Y=0.555
+ $X2=0.26 $Y2=0.43
r29 7 17 3.40825 $w=2.1e-07 $l=1.05e-07 $layer=LI1_cond $X=0.365 $Y=2.89
+ $X2=0.26 $Y2=2.89
r30 7 9 7.39394 $w=2.08e-07 $l=1.4e-07 $layer=LI1_cond $X=0.365 $Y=2.89
+ $X2=0.505 $Y2=2.89
r31 2 9 600 $w=1.7e-07 $l=2.7037e-07 $layer=licon1_PDIFF $count=1 $X=0.38
+ $Y=2.675 $X2=0.505 $Y2=2.89
r32 1 28 182 $w=1.7e-07 $l=2.498e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.43
.ends

.subckt PM_SKY130_FD_SC_LP__O2111A_M%VPWR 1 2 3 12 16 20 23 24 26 27 29 30 31 47
+ 48
r56 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r57 45 48 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r58 44 45 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r59 42 45 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r60 41 44 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.16 $Y=3.33 $X2=3.12
+ $Y2=3.33
r61 41 42 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r62 38 39 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r63 35 39 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r64 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r65 31 42 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=2.16 $Y2=3.33
r66 31 39 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=1.68 $Y2=3.33
r67 29 44 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=3.155 $Y=3.33
+ $X2=3.12 $Y2=3.33
r68 29 30 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.155 $Y=3.33
+ $X2=3.32 $Y2=3.33
r69 28 47 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=3.485 $Y=3.33
+ $X2=3.6 $Y2=3.33
r70 28 30 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.485 $Y=3.33
+ $X2=3.32 $Y2=3.33
r71 26 38 0.652406 $w=1.68e-07 $l=1e-08 $layer=LI1_cond $X=1.69 $Y=3.33 $X2=1.68
+ $Y2=3.33
r72 26 27 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.69 $Y=3.33
+ $X2=1.855 $Y2=3.33
r73 25 41 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=2.02 $Y=3.33
+ $X2=2.16 $Y2=3.33
r74 25 27 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.02 $Y=3.33
+ $X2=1.855 $Y2=3.33
r75 23 34 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=0.85 $Y=3.33
+ $X2=0.72 $Y2=3.33
r76 23 24 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=0.85 $Y=3.33
+ $X2=0.955 $Y2=3.33
r77 22 38 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=1.06 $Y=3.33
+ $X2=1.68 $Y2=3.33
r78 22 24 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.06 $Y=3.33
+ $X2=0.955 $Y2=3.33
r79 18 30 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.32 $Y=3.245
+ $X2=3.32 $Y2=3.33
r80 18 20 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=3.32 $Y=3.245
+ $X2=3.32 $Y2=2.95
r81 14 27 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.855 $Y=3.245
+ $X2=1.855 $Y2=3.33
r82 14 16 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.855 $Y=3.245
+ $X2=1.855 $Y2=2.95
r83 10 24 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=0.955 $Y=3.245
+ $X2=0.955 $Y2=3.33
r84 10 12 15.5801 $w=2.08e-07 $l=2.95e-07 $layer=LI1_cond $X=0.955 $Y=3.245
+ $X2=0.955 $Y2=2.95
r85 3 20 600 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=1 $X=3.18
+ $Y=2.675 $X2=3.32 $Y2=2.95
r86 2 16 600 $w=1.7e-07 $l=3.45868e-07 $layer=licon1_PDIFF $count=1 $X=1.695
+ $Y=2.675 $X2=1.855 $Y2=2.95
r87 1 12 600 $w=1.7e-07 $l=3.45868e-07 $layer=licon1_PDIFF $count=1 $X=0.795
+ $Y=2.675 $X2=0.955 $Y2=2.95
.ends

.subckt PM_SKY130_FD_SC_LP__O2111A_M%VGND 1 2 9 13 16 17 18 20 30 31 34
c53 31 0 2.58839e-20 $X=3.6 $Y=0
c54 20 0 1.12474e-19 $X=0.585 $Y=0
r55 34 35 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r56 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r57 28 31 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r58 27 28 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r59 25 34 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=0.795 $Y=0 $X2=0.69
+ $Y2=0
r60 25 27 120.369 $w=1.68e-07 $l=1.845e-06 $layer=LI1_cond $X=0.795 $Y=0
+ $X2=2.64 $Y2=0
r61 23 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r62 22 23 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r63 20 34 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=0.585 $Y=0 $X2=0.69
+ $Y2=0
r64 20 22 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.585 $Y=0 $X2=0.24
+ $Y2=0
r65 18 28 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=2.64
+ $Y2=0
r66 18 35 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=1.92 $Y=0 $X2=0.72
+ $Y2=0
r67 16 27 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=2.925 $Y=0 $X2=2.64
+ $Y2=0
r68 16 17 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=2.925 $Y=0 $X2=3.03
+ $Y2=0
r69 15 30 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=3.135 $Y=0 $X2=3.6
+ $Y2=0
r70 15 17 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=3.135 $Y=0 $X2=3.03
+ $Y2=0
r71 11 17 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=3.03 $Y=0.085
+ $X2=3.03 $Y2=0
r72 11 13 15.5801 $w=2.08e-07 $l=2.95e-07 $layer=LI1_cond $X=3.03 $Y=0.085
+ $X2=3.03 $Y2=0.38
r73 7 34 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=0.085
+ $X2=0.69 $Y2=0
r74 7 9 15.5801 $w=2.08e-07 $l=2.95e-07 $layer=LI1_cond $X=0.69 $Y=0.085
+ $X2=0.69 $Y2=0.38
r75 2 13 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=2.89
+ $Y=0.235 $X2=3.03 $Y2=0.38
r76 1 9 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.235 $X2=0.69 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_LP__O2111A_M%A_492_47# 1 2 9 11 12 15
r27 13 15 11.355 $w=2.08e-07 $l=2.15e-07 $layer=LI1_cond $X=3.46 $Y=0.725
+ $X2=3.46 $Y2=0.51
r28 11 13 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=3.355 $Y=0.81
+ $X2=3.46 $Y2=0.725
r29 11 12 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=3.355 $Y=0.81
+ $X2=2.705 $Y2=0.81
r30 7 12 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=2.61 $Y=0.725
+ $X2=2.705 $Y2=0.81
r31 7 9 12.5502 $w=1.88e-07 $l=2.15e-07 $layer=LI1_cond $X=2.61 $Y=0.725
+ $X2=2.61 $Y2=0.51
r32 2 15 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=3.32
+ $Y=0.235 $X2=3.46 $Y2=0.51
r33 1 9 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=2.46
+ $Y=0.235 $X2=2.6 $Y2=0.51
.ends

