* File: sky130_fd_sc_lp__nand3_lp.pex.spice
* Created: Wed Sep  2 10:04:31 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__NAND3_LP%C 3 7 11 12 13 14 18
r31 18 19 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.61
+ $Y=1.02 $X2=0.61 $Y2=1.02
r32 14 19 1.96371 $w=6.68e-07 $l=1.1e-07 $layer=LI1_cond $X=0.72 $Y=1.19
+ $X2=0.61 $Y2=1.19
r33 13 19 6.60521 $w=6.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.24 $Y=1.19
+ $X2=0.61 $Y2=1.19
r34 11 18 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.61 $Y=1.36
+ $X2=0.61 $Y2=1.02
r35 11 12 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.61 $Y=1.36
+ $X2=0.61 $Y2=1.525
r36 10 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.61 $Y=0.855
+ $X2=0.61 $Y2=1.02
r37 7 10 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=0.7 $Y=0.445 $X2=0.7
+ $Y2=0.855
r38 3 12 253.423 $w=2.5e-07 $l=1.02e-06 $layer=POLY_cond $X=0.65 $Y=2.545
+ $X2=0.65 $Y2=1.525
.ends

.subckt PM_SKY130_FD_SC_LP__NAND3_LP%B 3 4 6 9 10 11 12 13 18
c48 18 0 2.64121e-20 $X=1.18 $Y=0.93
r49 12 13 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.18 $Y=0.925
+ $X2=1.18 $Y2=1.295
r50 12 18 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.18
+ $Y=0.93 $X2=1.18 $Y2=0.93
r51 11 12 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.18 $Y=0.555
+ $X2=1.18 $Y2=0.925
r52 10 18 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.18 $Y=1.27
+ $X2=1.18 $Y2=0.93
r53 9 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.18 $Y=0.765
+ $X2=1.18 $Y2=0.93
r54 4 10 30.6163 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.18 $Y=1.435
+ $X2=1.18 $Y2=1.27
r55 4 6 275.784 $w=2.5e-07 $l=1.11e-06 $layer=POLY_cond $X=1.18 $Y=1.435
+ $X2=1.18 $Y2=2.545
r56 3 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.09 $Y=0.445 $X2=1.09
+ $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_LP__NAND3_LP%A 3 7 11 12 13 16 17
r37 16 17 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.75
+ $Y=1.02 $X2=1.75 $Y2=1.02
r38 13 17 9.05491 $w=3.48e-07 $l=2.75e-07 $layer=LI1_cond $X=1.74 $Y=1.295
+ $X2=1.74 $Y2=1.02
r39 11 16 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.75 $Y=1.36
+ $X2=1.75 $Y2=1.02
r40 11 12 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.75 $Y=1.36
+ $X2=1.75 $Y2=1.525
r41 10 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.75 $Y=0.855
+ $X2=1.75 $Y2=1.02
r42 7 12 253.423 $w=2.5e-07 $l=1.02e-06 $layer=POLY_cond $X=1.71 $Y=2.545
+ $X2=1.71 $Y2=1.525
r43 3 10 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=1.66 $Y=0.445
+ $X2=1.66 $Y2=0.855
.ends

.subckt PM_SKY130_FD_SC_LP__NAND3_LP%VPWR 1 2 7 9 15 20 21 22 29 30
r27 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r28 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r29 24 33 3.94169 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=3.33
+ $X2=0.212 $Y2=3.33
r30 24 26 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=0.425 $Y=3.33
+ $X2=1.2 $Y2=3.33
r31 22 30 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r32 22 34 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.24 $Y2=3.33
r33 22 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r34 20 26 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=1.28 $Y=3.33 $X2=1.2
+ $Y2=3.33
r35 20 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.28 $Y=3.33
+ $X2=1.445 $Y2=3.33
r36 19 29 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=1.61 $Y=3.33
+ $X2=2.16 $Y2=3.33
r37 19 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.61 $Y=3.33
+ $X2=1.445 $Y2=3.33
r38 15 18 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=1.445 $Y=2.22
+ $X2=1.445 $Y2=2.9
r39 13 21 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.445 $Y=3.245
+ $X2=1.445 $Y2=3.33
r40 13 18 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=1.445 $Y=3.245
+ $X2=1.445 $Y2=2.9
r41 9 12 32.7294 $w=2.48e-07 $l=7.1e-07 $layer=LI1_cond $X=0.3 $Y=2.19 $X2=0.3
+ $Y2=2.9
r42 7 33 3.20147 $w=2.5e-07 $l=1.23386e-07 $layer=LI1_cond $X=0.3 $Y=3.245
+ $X2=0.212 $Y2=3.33
r43 7 12 15.9037 $w=2.48e-07 $l=3.45e-07 $layer=LI1_cond $X=0.3 $Y=3.245 $X2=0.3
+ $Y2=2.9
r44 2 18 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=1.305
+ $Y=2.045 $X2=1.445 $Y2=2.9
r45 2 15 400 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_PDIFF $count=1 $X=1.305
+ $Y=2.045 $X2=1.445 $Y2=2.22
r46 1 12 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.195
+ $Y=2.045 $X2=0.34 $Y2=2.9
r47 1 9 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.195
+ $Y=2.045 $X2=0.34 $Y2=2.19
.ends

.subckt PM_SKY130_FD_SC_LP__NAND3_LP%Y 1 2 3 10 11 14 19 22 24 25 26 27
r46 27 40 3.14757 $w=4.73e-07 $l=1.25e-07 $layer=LI1_cond $X=0.842 $Y=2.775
+ $X2=0.842 $Y2=2.9
r47 26 27 9.31682 $w=4.73e-07 $l=3.7e-07 $layer=LI1_cond $X=0.842 $Y=2.405
+ $X2=0.842 $Y2=2.775
r48 26 34 5.41383 $w=4.73e-07 $l=2.15e-07 $layer=LI1_cond $X=0.842 $Y=2.405
+ $X2=0.842 $Y2=2.19
r49 25 34 3.90299 $w=4.73e-07 $l=1.55e-07 $layer=LI1_cond $X=0.842 $Y=2.035
+ $X2=0.842 $Y2=2.19
r50 20 25 4.0289 $w=4.73e-07 $l=1.6e-07 $layer=LI1_cond $X=0.842 $Y=1.875
+ $X2=0.842 $Y2=2.035
r51 19 24 3.03453 $w=3.12e-07 $l=1.80566e-07 $layer=LI1_cond $X=2.18 $Y=1.705
+ $X2=2.037 $Y2=1.79
r52 18 22 11.9263 $w=3.12e-07 $l=3.94398e-07 $layer=LI1_cond $X=2.18 $Y=0.675
+ $X2=1.875 $Y2=0.47
r53 18 19 67.1979 $w=1.68e-07 $l=1.03e-06 $layer=LI1_cond $X=2.18 $Y=0.675
+ $X2=2.18 $Y2=1.705
r54 14 16 18.6641 $w=4.53e-07 $l=7.1e-07 $layer=LI1_cond $X=2.037 $Y=2.19
+ $X2=2.037 $Y2=2.9
r55 12 24 3.03453 $w=3.12e-07 $l=8.5e-08 $layer=LI1_cond $X=2.037 $Y=1.875
+ $X2=2.037 $Y2=1.79
r56 12 14 8.28054 $w=4.53e-07 $l=3.15e-07 $layer=LI1_cond $X=2.037 $Y=1.875
+ $X2=2.037 $Y2=2.19
r57 11 20 9.01902 $w=1.7e-07 $l=2.77262e-07 $layer=LI1_cond $X=1.08 $Y=1.79
+ $X2=0.842 $Y2=1.875
r58 10 24 3.60271 $w=1.7e-07 $l=2.27e-07 $layer=LI1_cond $X=1.81 $Y=1.79
+ $X2=2.037 $Y2=1.79
r59 10 11 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=1.81 $Y=1.79
+ $X2=1.08 $Y2=1.79
r60 3 16 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=1.835
+ $Y=2.045 $X2=1.975 $Y2=2.9
r61 3 14 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.835
+ $Y=2.045 $X2=1.975 $Y2=2.19
r62 2 40 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=0.775
+ $Y=2.045 $X2=0.915 $Y2=2.9
r63 2 34 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.775
+ $Y=2.045 $X2=0.915 $Y2=2.19
r64 1 22 182 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=1 $X=1.735
+ $Y=0.235 $X2=1.875 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_LP__NAND3_LP%VGND 1 6 9 10 11 21 22
c26 22 0 2.64121e-20 $X=2.16 $Y=0
r27 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r28 18 21 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=0.72 $Y=0 $X2=2.16
+ $Y2=0
r29 18 19 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r30 15 19 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r31 14 15 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r32 11 22 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r33 11 19 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r34 9 14 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=0.32 $Y=0 $X2=0.24
+ $Y2=0
r35 9 10 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.32 $Y=0 $X2=0.485
+ $Y2=0
r36 8 18 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=0.65 $Y=0 $X2=0.72
+ $Y2=0
r37 8 10 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.65 $Y=0 $X2=0.485
+ $Y2=0
r38 4 10 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.485 $Y=0.085
+ $X2=0.485 $Y2=0
r39 4 6 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=0.485 $Y=0.085
+ $X2=0.485 $Y2=0.445
r40 1 6 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.34
+ $Y=0.235 $X2=0.485 $Y2=0.445
.ends

