* File: sky130_fd_sc_lp__o32ai_2.pxi.spice
* Created: Fri Aug 28 11:18:25 2020
* 
x_PM_SKY130_FD_SC_LP__O32AI_2%B2 N_B2_M1004_g N_B2_M1005_g N_B2_M1019_g
+ N_B2_M1015_g B2 B2 B2 N_B2_c_91_n PM_SKY130_FD_SC_LP__O32AI_2%B2
x_PM_SKY130_FD_SC_LP__O32AI_2%B1 N_B1_M1008_g N_B1_M1006_g N_B1_M1016_g
+ N_B1_M1012_g B1 N_B1_c_137_n N_B1_c_134_n PM_SKY130_FD_SC_LP__O32AI_2%B1
x_PM_SKY130_FD_SC_LP__O32AI_2%A3 N_A3_M1007_g N_A3_M1011_g N_A3_M1017_g
+ N_A3_M1018_g A3 A3 N_A3_c_184_n PM_SKY130_FD_SC_LP__O32AI_2%A3
x_PM_SKY130_FD_SC_LP__O32AI_2%A2 N_A2_M1003_g N_A2_c_241_n N_A2_M1002_g
+ N_A2_M1014_g N_A2_c_243_n N_A2_M1013_g A2 A2 A2 N_A2_c_245_n
+ PM_SKY130_FD_SC_LP__O32AI_2%A2
x_PM_SKY130_FD_SC_LP__O32AI_2%A1 N_A1_c_295_n N_A1_M1001_g N_A1_M1000_g
+ N_A1_c_297_n N_A1_M1010_g N_A1_M1009_g A1 A1 A1 N_A1_c_300_n
+ PM_SKY130_FD_SC_LP__O32AI_2%A1
x_PM_SKY130_FD_SC_LP__O32AI_2%A_39_367# N_A_39_367#_M1005_d N_A_39_367#_M1015_d
+ N_A_39_367#_M1016_d N_A_39_367#_c_334_n N_A_39_367#_c_335_n
+ N_A_39_367#_c_339_n N_A_39_367#_c_346_p N_A_39_367#_c_341_n
+ N_A_39_367#_c_336_n N_A_39_367#_c_337_n PM_SKY130_FD_SC_LP__O32AI_2%A_39_367#
x_PM_SKY130_FD_SC_LP__O32AI_2%Y N_Y_M1004_s N_Y_M1006_d N_Y_M1005_s N_Y_M1011_s
+ N_Y_c_371_n N_Y_c_364_n N_Y_c_365_n N_Y_c_370_n N_Y_c_393_n N_Y_c_366_n
+ N_Y_c_381_n N_Y_c_367_n Y Y Y Y N_Y_c_368_n Y PM_SKY130_FD_SC_LP__O32AI_2%Y
x_PM_SKY130_FD_SC_LP__O32AI_2%VPWR N_VPWR_M1008_s N_VPWR_M1000_d N_VPWR_M1009_d
+ N_VPWR_c_451_n N_VPWR_c_452_n N_VPWR_c_453_n N_VPWR_c_454_n VPWR
+ N_VPWR_c_455_n N_VPWR_c_456_n N_VPWR_c_457_n N_VPWR_c_458_n N_VPWR_c_459_n
+ N_VPWR_c_450_n PM_SKY130_FD_SC_LP__O32AI_2%VPWR
x_PM_SKY130_FD_SC_LP__O32AI_2%A_519_365# N_A_519_365#_M1011_d
+ N_A_519_365#_M1017_d N_A_519_365#_M1014_s N_A_519_365#_c_525_n
+ N_A_519_365#_c_530_n N_A_519_365#_c_526_n N_A_519_365#_c_527_n
+ N_A_519_365#_c_536_n N_A_519_365#_c_528_n N_A_519_365#_c_529_n
+ N_A_519_365#_c_560_n PM_SKY130_FD_SC_LP__O32AI_2%A_519_365#
x_PM_SKY130_FD_SC_LP__O32AI_2%A_778_365# N_A_778_365#_M1003_d
+ N_A_778_365#_M1000_s N_A_778_365#_c_570_n N_A_778_365#_c_567_n
+ N_A_778_365#_c_568_n N_A_778_365#_c_589_n
+ PM_SKY130_FD_SC_LP__O32AI_2%A_778_365#
x_PM_SKY130_FD_SC_LP__O32AI_2%A_39_65# N_A_39_65#_M1004_d N_A_39_65#_M1019_d
+ N_A_39_65#_M1012_s N_A_39_65#_M1018_d N_A_39_65#_M1013_s N_A_39_65#_M1010_s
+ N_A_39_65#_c_598_n N_A_39_65#_c_599_n N_A_39_65#_c_600_n N_A_39_65#_c_611_n
+ N_A_39_65#_c_601_n N_A_39_65#_c_617_n N_A_39_65#_c_618_n N_A_39_65#_c_621_n
+ N_A_39_65#_c_602_n N_A_39_65#_c_625_n N_A_39_65#_c_603_n N_A_39_65#_c_633_n
+ N_A_39_65#_c_604_n N_A_39_65#_c_605_n N_A_39_65#_c_606_n N_A_39_65#_c_623_n
+ N_A_39_65#_c_631_n PM_SKY130_FD_SC_LP__O32AI_2%A_39_65#
x_PM_SKY130_FD_SC_LP__O32AI_2%VGND N_VGND_M1007_s N_VGND_M1002_d N_VGND_M1001_d
+ N_VGND_c_687_n N_VGND_c_688_n VGND N_VGND_c_689_n N_VGND_c_690_n
+ N_VGND_c_691_n N_VGND_c_692_n N_VGND_c_693_n N_VGND_c_694_n N_VGND_c_695_n
+ N_VGND_c_696_n PM_SKY130_FD_SC_LP__O32AI_2%VGND
cc_1 VNB N_B2_M1004_g 0.0266153f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=0.745
cc_2 VNB N_B2_M1019_g 0.0202092f $X=-0.19 $Y=-0.245 $X2=0.965 $Y2=0.745
cc_3 VNB B2 0.0223688f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_4 VNB N_B2_c_91_n 0.036998f $X=-0.19 $Y=-0.245 $X2=0.965 $Y2=1.51
cc_5 VNB N_B1_M1006_g 0.0211501f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=2.465
cc_6 VNB N_B1_M1012_g 0.0211509f $X=-0.19 $Y=-0.245 $X2=0.965 $Y2=2.465
cc_7 VNB N_B1_c_134_n 0.0425442f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A3_M1007_g 0.0233101f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=0.745
cc_9 VNB N_A3_M1018_g 0.021653f $X=-0.19 $Y=-0.245 $X2=0.965 $Y2=2.465
cc_10 VNB A3 0.00334612f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_11 VNB N_A3_c_184_n 0.0624887f $X=-0.19 $Y=-0.245 $X2=0.965 $Y2=1.51
cc_12 VNB N_A2_M1003_g 0.00193877f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=0.745
cc_13 VNB N_A2_c_241_n 0.0164117f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=1.675
cc_14 VNB N_A2_M1014_g 0.0031385f $X=-0.19 $Y=-0.245 $X2=0.965 $Y2=0.745
cc_15 VNB N_A2_c_243_n 0.016814f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB A2 0.0143443f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_17 VNB N_A2_c_245_n 0.049318f $X=-0.19 $Y=-0.245 $X2=0.965 $Y2=1.51
cc_18 VNB N_A1_c_295_n 0.0163787f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=1.345
cc_19 VNB N_A1_M1000_g 0.00394324f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=2.465
cc_20 VNB N_A1_c_297_n 0.021262f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A1_M1009_g 0.00394324f $X=-0.19 $Y=-0.245 $X2=0.965 $Y2=1.675
cc_22 VNB A1 0.0514447f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_23 VNB N_A1_c_300_n 0.0789316f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_Y_c_364_n 0.00397373f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_25 VNB N_Y_c_365_n 0.00233022f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_Y_c_366_n 0.00682621f $X=-0.19 $Y=-0.245 $X2=0.625 $Y2=1.51
cc_27 VNB N_Y_c_367_n 0.00273928f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_Y_c_368_n 6.83794e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB Y 0.00168637f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VPWR_c_450_n 0.263193f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_39_65#_c_598_n 0.0315835f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_39_65#_c_599_n 0.0026914f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=1.51
cc_33 VNB N_A_39_65#_c_600_n 0.00928796f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_39_65#_c_601_n 0.00516631f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_39_65#_c_602_n 0.00177084f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_39_65#_c_603_n 0.00177527f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_39_65#_c_604_n 0.00742876f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_39_65#_c_605_n 0.0230663f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_39_65#_c_606_n 0.00221131f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_687_n 0.00392812f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_688_n 0.00231989f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_689_n 0.0139151f $X=-0.19 $Y=-0.245 $X2=0.625 $Y2=1.51
cc_43 VNB N_VGND_c_690_n 0.0155947f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.587
cc_44 VNB N_VGND_c_691_n 0.0337392f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_692_n 0.357705f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_693_n 0.0625057f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_694_n 0.023216f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_695_n 0.00581671f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_696_n 0.00549308f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VPB N_B2_M1005_g 0.0244533f $X=-0.19 $Y=1.655 $X2=0.535 $Y2=2.465
cc_51 VPB N_B2_M1015_g 0.0183424f $X=-0.19 $Y=1.655 $X2=0.965 $Y2=2.465
cc_52 VPB B2 0.0169798f $X=-0.19 $Y=1.655 $X2=1.115 $Y2=1.58
cc_53 VPB N_B2_c_91_n 0.00492723f $X=-0.19 $Y=1.655 $X2=0.965 $Y2=1.51
cc_54 VPB N_B1_M1008_g 0.0183955f $X=-0.19 $Y=1.655 $X2=0.535 $Y2=0.745
cc_55 VPB N_B1_M1016_g 0.0234657f $X=-0.19 $Y=1.655 $X2=0.965 $Y2=0.745
cc_56 VPB N_B1_c_137_n 0.00259635f $X=-0.19 $Y=1.655 $X2=0.535 $Y2=1.51
cc_57 VPB N_B1_c_134_n 0.0100899f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_58 VPB N_A3_M1011_g 0.0232781f $X=-0.19 $Y=1.655 $X2=0.535 $Y2=2.465
cc_59 VPB N_A3_M1017_g 0.0183784f $X=-0.19 $Y=1.655 $X2=0.965 $Y2=0.745
cc_60 VPB A3 0.00867f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_61 VPB N_A3_c_184_n 0.0220472f $X=-0.19 $Y=1.655 $X2=0.965 $Y2=1.51
cc_62 VPB N_A2_M1003_g 0.0195851f $X=-0.19 $Y=1.655 $X2=0.535 $Y2=0.745
cc_63 VPB N_A2_M1014_g 0.0250403f $X=-0.19 $Y=1.655 $X2=0.965 $Y2=0.745
cc_64 VPB N_A1_M1000_g 0.0239519f $X=-0.19 $Y=1.655 $X2=0.535 $Y2=2.465
cc_65 VPB N_A1_M1009_g 0.0272339f $X=-0.19 $Y=1.655 $X2=0.965 $Y2=1.675
cc_66 VPB N_A_39_367#_c_334_n 0.00746637f $X=-0.19 $Y=1.655 $X2=0.965 $Y2=0.745
cc_67 VPB N_A_39_367#_c_335_n 0.0374018f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_68 VPB N_A_39_367#_c_336_n 0.00261307f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_69 VPB N_A_39_367#_c_337_n 0.00747662f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_70 VPB N_Y_c_370_n 0.0188943f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_71 VPB N_VPWR_c_451_n 4.89148e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_72 VPB N_VPWR_c_452_n 0.0125161f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_73 VPB N_VPWR_c_453_n 0.0153455f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_74 VPB N_VPWR_c_454_n 0.0571176f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_75 VPB N_VPWR_c_455_n 0.0362774f $X=-0.19 $Y=1.655 $X2=0.965 $Y2=1.51
cc_76 VPB N_VPWR_c_456_n 0.0732202f $X=-0.19 $Y=1.655 $X2=1.2 $Y2=1.587
cc_77 VPB N_VPWR_c_457_n 0.0147711f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_78 VPB N_VPWR_c_458_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_79 VPB N_VPWR_c_459_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_80 VPB N_VPWR_c_450_n 0.0766113f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_81 VPB N_A_519_365#_c_525_n 0.0076747f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_82 VPB N_A_519_365#_c_526_n 0.00227906f $X=-0.19 $Y=1.655 $X2=0.965 $Y2=2.465
cc_83 VPB N_A_519_365#_c_527_n 0.00223364f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_84 VPB N_A_519_365#_c_528_n 0.001829f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_85 VPB N_A_519_365#_c_529_n 0.00801052f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_86 VPB N_A_778_365#_c_567_n 0.0200434f $X=-0.19 $Y=1.655 $X2=0.965 $Y2=1.675
cc_87 VPB N_A_778_365#_c_568_n 0.00233203f $X=-0.19 $Y=1.655 $X2=0.965 $Y2=2.465
cc_88 N_B2_M1015_g N_B1_M1008_g 0.0259112f $X=0.965 $Y=2.465 $X2=0 $Y2=0
cc_89 N_B2_M1019_g N_B1_M1006_g 0.0250346f $X=0.965 $Y=0.745 $X2=0 $Y2=0
cc_90 B2 N_B1_c_137_n 0.0273862f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_91 N_B2_c_91_n N_B1_c_137_n 2.20764e-19 $X=0.965 $Y=1.51 $X2=0 $Y2=0
cc_92 B2 N_B1_c_134_n 0.00325621f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_93 N_B2_c_91_n N_B1_c_134_n 0.0259112f $X=0.965 $Y=1.51 $X2=0 $Y2=0
cc_94 B2 N_A_39_367#_c_335_n 0.0219167f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_95 N_B2_M1005_g N_A_39_367#_c_339_n 0.0114565f $X=0.535 $Y=2.465 $X2=0 $Y2=0
cc_96 N_B2_M1015_g N_A_39_367#_c_339_n 0.0115031f $X=0.965 $Y=2.465 $X2=0 $Y2=0
cc_97 N_B2_M1004_g N_Y_c_371_n 0.0054303f $X=0.535 $Y=0.745 $X2=0 $Y2=0
cc_98 N_B2_M1019_g N_Y_c_371_n 0.00686014f $X=0.965 $Y=0.745 $X2=0 $Y2=0
cc_99 N_B2_M1019_g N_Y_c_364_n 0.00962413f $X=0.965 $Y=0.745 $X2=0 $Y2=0
cc_100 B2 N_Y_c_364_n 0.0278798f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_101 N_B2_M1004_g N_Y_c_365_n 0.00530981f $X=0.535 $Y=0.745 $X2=0 $Y2=0
cc_102 N_B2_M1019_g N_Y_c_365_n 0.00169298f $X=0.965 $Y=0.745 $X2=0 $Y2=0
cc_103 B2 N_Y_c_365_n 0.0263068f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_104 N_B2_c_91_n N_Y_c_365_n 0.00254667f $X=0.965 $Y=1.51 $X2=0 $Y2=0
cc_105 N_B2_M1015_g N_Y_c_370_n 0.0111034f $X=0.965 $Y=2.465 $X2=0 $Y2=0
cc_106 B2 N_Y_c_370_n 0.0255027f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_107 N_B2_M1005_g N_Y_c_381_n 0.0120634f $X=0.535 $Y=2.465 $X2=0 $Y2=0
cc_108 N_B2_M1015_g N_Y_c_381_n 0.0116361f $X=0.965 $Y=2.465 $X2=0 $Y2=0
cc_109 B2 N_Y_c_381_n 0.0230324f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_110 N_B2_c_91_n N_Y_c_381_n 6.52992e-19 $X=0.965 $Y=1.51 $X2=0 $Y2=0
cc_111 N_B2_M1015_g N_VPWR_c_451_n 0.00109252f $X=0.965 $Y=2.465 $X2=0 $Y2=0
cc_112 N_B2_M1005_g N_VPWR_c_455_n 0.00357877f $X=0.535 $Y=2.465 $X2=0 $Y2=0
cc_113 N_B2_M1015_g N_VPWR_c_455_n 0.00357877f $X=0.965 $Y=2.465 $X2=0 $Y2=0
cc_114 N_B2_M1005_g N_VPWR_c_450_n 0.00633582f $X=0.535 $Y=2.465 $X2=0 $Y2=0
cc_115 N_B2_M1015_g N_VPWR_c_450_n 0.00537654f $X=0.965 $Y=2.465 $X2=0 $Y2=0
cc_116 N_B2_M1004_g N_A_39_65#_c_598_n 0.00354524f $X=0.535 $Y=0.745 $X2=0 $Y2=0
cc_117 B2 N_A_39_65#_c_598_n 0.0179011f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_118 N_B2_M1004_g N_A_39_65#_c_599_n 0.0125492f $X=0.535 $Y=0.745 $X2=0 $Y2=0
cc_119 N_B2_M1019_g N_A_39_65#_c_599_n 0.0115989f $X=0.965 $Y=0.745 $X2=0 $Y2=0
cc_120 N_B2_M1004_g N_VGND_c_692_n 0.00472541f $X=0.535 $Y=0.745 $X2=0 $Y2=0
cc_121 N_B2_M1019_g N_VGND_c_692_n 0.00442601f $X=0.965 $Y=0.745 $X2=0 $Y2=0
cc_122 N_B2_M1004_g N_VGND_c_693_n 0.00302501f $X=0.535 $Y=0.745 $X2=0 $Y2=0
cc_123 N_B2_M1019_g N_VGND_c_693_n 0.00302501f $X=0.965 $Y=0.745 $X2=0 $Y2=0
cc_124 N_B1_M1012_g N_A3_M1007_g 0.0188067f $X=1.985 $Y=0.745 $X2=0 $Y2=0
cc_125 N_B1_M1016_g A3 0.00148355f $X=1.825 $Y=2.465 $X2=0 $Y2=0
cc_126 N_B1_c_137_n A3 0.0263254f $X=1.63 $Y=1.51 $X2=0 $Y2=0
cc_127 N_B1_c_134_n A3 0.011431f $X=1.825 $Y=1.512 $X2=0 $Y2=0
cc_128 N_B1_c_134_n N_A3_c_184_n 0.0188067f $X=1.825 $Y=1.512 $X2=0 $Y2=0
cc_129 N_B1_M1008_g N_A_39_367#_c_341_n 0.0127523f $X=1.395 $Y=2.465 $X2=0 $Y2=0
cc_130 N_B1_M1016_g N_A_39_367#_c_341_n 0.0128101f $X=1.825 $Y=2.465 $X2=0 $Y2=0
cc_131 N_B1_M1006_g N_Y_c_371_n 5.37284e-19 $X=1.475 $Y=0.745 $X2=0 $Y2=0
cc_132 N_B1_M1006_g N_Y_c_364_n 0.0141584f $X=1.475 $Y=0.745 $X2=0 $Y2=0
cc_133 N_B1_c_137_n N_Y_c_364_n 0.00968915f $X=1.63 $Y=1.51 $X2=0 $Y2=0
cc_134 N_B1_c_134_n N_Y_c_364_n 0.00273777f $X=1.825 $Y=1.512 $X2=0 $Y2=0
cc_135 N_B1_M1008_g N_Y_c_370_n 0.0123503f $X=1.395 $Y=2.465 $X2=0 $Y2=0
cc_136 N_B1_M1016_g N_Y_c_370_n 0.0135832f $X=1.825 $Y=2.465 $X2=0 $Y2=0
cc_137 N_B1_c_137_n N_Y_c_370_n 0.0236964f $X=1.63 $Y=1.51 $X2=0 $Y2=0
cc_138 N_B1_c_134_n N_Y_c_370_n 0.00343095f $X=1.825 $Y=1.512 $X2=0 $Y2=0
cc_139 N_B1_M1012_g N_Y_c_393_n 0.00685613f $X=1.985 $Y=0.745 $X2=0 $Y2=0
cc_140 N_B1_M1012_g N_Y_c_366_n 0.0103202f $X=1.985 $Y=0.745 $X2=0 $Y2=0
cc_141 N_B1_M1008_g N_Y_c_381_n 7.61713e-19 $X=1.395 $Y=2.465 $X2=0 $Y2=0
cc_142 N_B1_M1012_g N_Y_c_367_n 0.00215177f $X=1.985 $Y=0.745 $X2=0 $Y2=0
cc_143 N_B1_c_137_n N_Y_c_367_n 0.0180907f $X=1.63 $Y=1.51 $X2=0 $Y2=0
cc_144 N_B1_c_134_n N_Y_c_367_n 0.00526163f $X=1.825 $Y=1.512 $X2=0 $Y2=0
cc_145 N_B1_M1008_g N_VPWR_c_451_n 0.0119212f $X=1.395 $Y=2.465 $X2=0 $Y2=0
cc_146 N_B1_M1016_g N_VPWR_c_451_n 0.0124844f $X=1.825 $Y=2.465 $X2=0 $Y2=0
cc_147 N_B1_M1008_g N_VPWR_c_455_n 0.00486043f $X=1.395 $Y=2.465 $X2=0 $Y2=0
cc_148 N_B1_M1016_g N_VPWR_c_456_n 0.00486043f $X=1.825 $Y=2.465 $X2=0 $Y2=0
cc_149 N_B1_M1008_g N_VPWR_c_450_n 0.0082726f $X=1.395 $Y=2.465 $X2=0 $Y2=0
cc_150 N_B1_M1016_g N_VPWR_c_450_n 0.00954696f $X=1.825 $Y=2.465 $X2=0 $Y2=0
cc_151 N_B1_M1006_g N_A_39_65#_c_611_n 0.00686522f $X=1.475 $Y=0.745 $X2=0 $Y2=0
cc_152 N_B1_M1012_g N_A_39_65#_c_611_n 5.37284e-19 $X=1.985 $Y=0.745 $X2=0 $Y2=0
cc_153 N_B1_M1006_g N_A_39_65#_c_601_n 0.00872289f $X=1.475 $Y=0.745 $X2=0 $Y2=0
cc_154 N_B1_M1012_g N_A_39_65#_c_601_n 0.0120426f $X=1.985 $Y=0.745 $X2=0 $Y2=0
cc_155 N_B1_M1006_g N_A_39_65#_c_606_n 0.00152212f $X=1.475 $Y=0.745 $X2=0 $Y2=0
cc_156 N_B1_M1006_g N_VGND_c_692_n 0.00450051f $X=1.475 $Y=0.745 $X2=0 $Y2=0
cc_157 N_B1_M1012_g N_VGND_c_692_n 0.00450053f $X=1.985 $Y=0.745 $X2=0 $Y2=0
cc_158 N_B1_M1006_g N_VGND_c_693_n 0.00302473f $X=1.475 $Y=0.745 $X2=0 $Y2=0
cc_159 N_B1_M1012_g N_VGND_c_693_n 0.00302501f $X=1.985 $Y=0.745 $X2=0 $Y2=0
cc_160 N_A3_M1017_g N_A2_M1003_g 0.0183714f $X=3.385 $Y=2.455 $X2=0 $Y2=0
cc_161 N_A3_c_184_n N_A2_M1003_g 0.0134043f $X=3.455 $Y=1.5 $X2=0 $Y2=0
cc_162 N_A3_M1018_g N_A2_c_241_n 0.0138675f $X=3.455 $Y=0.745 $X2=0 $Y2=0
cc_163 N_A3_M1018_g A2 0.00296014f $X=3.455 $Y=0.745 $X2=0 $Y2=0
cc_164 N_A3_c_184_n A2 0.00520636f $X=3.455 $Y=1.5 $X2=0 $Y2=0
cc_165 N_A3_M1018_g N_A2_c_245_n 0.0134043f $X=3.455 $Y=0.745 $X2=0 $Y2=0
cc_166 N_A3_M1011_g N_Y_c_370_n 0.0148007f $X=2.955 $Y=2.455 $X2=0 $Y2=0
cc_167 A3 N_Y_c_370_n 0.0653048f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_168 N_A3_c_184_n N_Y_c_370_n 0.00230347f $X=3.455 $Y=1.5 $X2=0 $Y2=0
cc_169 N_A3_M1007_g N_Y_c_393_n 5.37284e-19 $X=2.495 $Y=0.745 $X2=0 $Y2=0
cc_170 N_A3_M1007_g N_Y_c_366_n 0.0129134f $X=2.495 $Y=0.745 $X2=0 $Y2=0
cc_171 A3 N_Y_c_366_n 0.0635312f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_172 N_A3_c_184_n N_Y_c_366_n 0.0100043f $X=3.455 $Y=1.5 $X2=0 $Y2=0
cc_173 N_A3_M1011_g Y 0.0132198f $X=2.955 $Y=2.455 $X2=0 $Y2=0
cc_174 N_A3_M1017_g Y 0.00856137f $X=3.385 $Y=2.455 $X2=0 $Y2=0
cc_175 N_A3_M1018_g N_Y_c_368_n 0.00467723f $X=3.455 $Y=0.745 $X2=0 $Y2=0
cc_176 N_A3_M1007_g Y 0.00249618f $X=2.495 $Y=0.745 $X2=0 $Y2=0
cc_177 N_A3_M1011_g Y 0.010152f $X=2.955 $Y=2.455 $X2=0 $Y2=0
cc_178 N_A3_M1017_g Y 0.00558299f $X=3.385 $Y=2.455 $X2=0 $Y2=0
cc_179 N_A3_M1018_g Y 0.00201636f $X=3.455 $Y=0.745 $X2=0 $Y2=0
cc_180 A3 Y 0.0269216f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_181 N_A3_c_184_n Y 0.0301779f $X=3.455 $Y=1.5 $X2=0 $Y2=0
cc_182 N_A3_M1011_g N_VPWR_c_456_n 0.00351226f $X=2.955 $Y=2.455 $X2=0 $Y2=0
cc_183 N_A3_M1017_g N_VPWR_c_456_n 0.00351226f $X=3.385 $Y=2.455 $X2=0 $Y2=0
cc_184 N_A3_M1011_g N_VPWR_c_450_n 0.00660267f $X=2.955 $Y=2.455 $X2=0 $Y2=0
cc_185 N_A3_M1017_g N_VPWR_c_450_n 0.00532831f $X=3.385 $Y=2.455 $X2=0 $Y2=0
cc_186 N_A3_M1011_g N_A_519_365#_c_530_n 0.0114688f $X=2.955 $Y=2.455 $X2=0
+ $Y2=0
cc_187 N_A3_M1017_g N_A_519_365#_c_530_n 0.0114688f $X=3.385 $Y=2.455 $X2=0
+ $Y2=0
cc_188 N_A3_M1017_g N_A_519_365#_c_527_n 7.13716e-19 $X=3.385 $Y=2.455 $X2=0
+ $Y2=0
cc_189 N_A3_c_184_n N_A_519_365#_c_527_n 7.16965e-19 $X=3.455 $Y=1.5 $X2=0 $Y2=0
cc_190 N_A3_M1017_g N_A_778_365#_c_568_n 3.39246e-19 $X=3.385 $Y=2.455 $X2=0
+ $Y2=0
cc_191 N_A3_M1007_g N_A_39_65#_c_601_n 0.00295806f $X=2.495 $Y=0.745 $X2=0 $Y2=0
cc_192 N_A3_M1007_g N_A_39_65#_c_617_n 0.00883436f $X=2.495 $Y=0.745 $X2=0 $Y2=0
cc_193 N_A3_M1007_g N_A_39_65#_c_618_n 0.0108024f $X=2.495 $Y=0.745 $X2=0 $Y2=0
cc_194 N_A3_M1018_g N_A_39_65#_c_618_n 0.0148893f $X=3.455 $Y=0.745 $X2=0 $Y2=0
cc_195 N_A3_c_184_n N_A_39_65#_c_618_n 0.00159091f $X=3.455 $Y=1.5 $X2=0 $Y2=0
cc_196 N_A3_M1007_g N_A_39_65#_c_621_n 7.31417e-19 $X=2.495 $Y=0.745 $X2=0 $Y2=0
cc_197 N_A3_M1018_g N_A_39_65#_c_602_n 3.36571e-19 $X=3.455 $Y=0.745 $X2=0 $Y2=0
cc_198 N_A3_M1018_g N_A_39_65#_c_623_n 0.00782491f $X=3.455 $Y=0.745 $X2=0 $Y2=0
cc_199 N_A3_M1018_g N_VGND_c_687_n 4.76318e-19 $X=3.455 $Y=0.745 $X2=0 $Y2=0
cc_200 N_A3_M1018_g N_VGND_c_689_n 0.00306556f $X=3.455 $Y=0.745 $X2=0 $Y2=0
cc_201 N_A3_M1007_g N_VGND_c_692_n 0.00551025f $X=2.495 $Y=0.745 $X2=0 $Y2=0
cc_202 N_A3_M1018_g N_VGND_c_692_n 0.00390569f $X=3.455 $Y=0.745 $X2=0 $Y2=0
cc_203 N_A3_M1007_g N_VGND_c_693_n 0.0035672f $X=2.495 $Y=0.745 $X2=0 $Y2=0
cc_204 N_A3_M1007_g N_VGND_c_694_n 0.00859154f $X=2.495 $Y=0.745 $X2=0 $Y2=0
cc_205 N_A3_M1018_g N_VGND_c_694_n 0.00839472f $X=3.455 $Y=0.745 $X2=0 $Y2=0
cc_206 N_A2_c_243_n N_A1_c_295_n 0.0142994f $X=4.355 $Y=1.275 $X2=-0.19
+ $Y2=-0.245
cc_207 A2 N_A1_c_295_n 0.00257327f $X=4.475 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_208 A2 A1 0.0278594f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_209 N_A2_c_245_n N_A1_c_300_n 0.0231325f $X=4.355 $Y=1.44 $X2=0 $Y2=0
cc_210 A2 N_Y_c_368_n 0.00303081f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_211 A2 Y 0.0225543f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_212 N_A2_c_245_n Y 0.00133436f $X=4.355 $Y=1.44 $X2=0 $Y2=0
cc_213 N_A2_M1014_g N_VPWR_c_452_n 0.00221807f $X=4.245 $Y=2.455 $X2=0 $Y2=0
cc_214 N_A2_M1003_g N_VPWR_c_456_n 0.00351226f $X=3.815 $Y=2.455 $X2=0 $Y2=0
cc_215 N_A2_M1014_g N_VPWR_c_456_n 0.00351226f $X=4.245 $Y=2.455 $X2=0 $Y2=0
cc_216 N_A2_M1003_g N_VPWR_c_450_n 0.00532831f $X=3.815 $Y=2.455 $X2=0 $Y2=0
cc_217 N_A2_M1014_g N_VPWR_c_450_n 0.00660267f $X=4.245 $Y=2.455 $X2=0 $Y2=0
cc_218 N_A2_M1003_g N_A_519_365#_c_527_n 7.13575e-19 $X=3.815 $Y=2.455 $X2=0
+ $Y2=0
cc_219 A2 N_A_519_365#_c_527_n 0.0113192f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_220 N_A2_M1003_g N_A_519_365#_c_536_n 0.0114688f $X=3.815 $Y=2.455 $X2=0
+ $Y2=0
cc_221 N_A2_M1014_g N_A_519_365#_c_536_n 0.0114688f $X=4.245 $Y=2.455 $X2=0
+ $Y2=0
cc_222 N_A2_M1003_g N_A_778_365#_c_570_n 0.00900833f $X=3.815 $Y=2.455 $X2=0
+ $Y2=0
cc_223 N_A2_M1014_g N_A_778_365#_c_570_n 0.0150032f $X=4.245 $Y=2.455 $X2=0
+ $Y2=0
cc_224 N_A2_M1014_g N_A_778_365#_c_567_n 0.0132413f $X=4.245 $Y=2.455 $X2=0
+ $Y2=0
cc_225 A2 N_A_778_365#_c_567_n 0.0323749f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_226 N_A2_c_245_n N_A_778_365#_c_567_n 0.00487589f $X=4.355 $Y=1.44 $X2=0
+ $Y2=0
cc_227 N_A2_M1003_g N_A_778_365#_c_568_n 0.00433988f $X=3.815 $Y=2.455 $X2=0
+ $Y2=0
cc_228 N_A2_M1014_g N_A_778_365#_c_568_n 0.00219014f $X=4.245 $Y=2.455 $X2=0
+ $Y2=0
cc_229 A2 N_A_778_365#_c_568_n 0.0263482f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_230 N_A2_c_245_n N_A_778_365#_c_568_n 0.00289569f $X=4.355 $Y=1.44 $X2=0
+ $Y2=0
cc_231 N_A2_c_241_n N_A_39_65#_c_602_n 4.47497e-19 $X=3.895 $Y=1.275 $X2=0 $Y2=0
cc_232 N_A2_c_241_n N_A_39_65#_c_625_n 0.0122731f $X=3.895 $Y=1.275 $X2=0 $Y2=0
cc_233 N_A2_c_243_n N_A_39_65#_c_625_n 0.0129225f $X=4.355 $Y=1.275 $X2=0 $Y2=0
cc_234 A2 N_A_39_65#_c_625_n 0.0445178f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_235 N_A2_c_245_n N_A_39_65#_c_625_n 7.61863e-19 $X=4.355 $Y=1.44 $X2=0 $Y2=0
cc_236 N_A2_c_243_n N_A_39_65#_c_603_n 4.46796e-19 $X=4.355 $Y=1.275 $X2=0 $Y2=0
cc_237 A2 N_A_39_65#_c_623_n 0.019785f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_238 A2 N_A_39_65#_c_631_n 0.0145642f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_239 N_A2_c_241_n N_VGND_c_687_n 0.00867825f $X=3.895 $Y=1.275 $X2=0 $Y2=0
cc_240 N_A2_c_243_n N_VGND_c_687_n 0.00205177f $X=4.355 $Y=1.275 $X2=0 $Y2=0
cc_241 N_A2_c_243_n N_VGND_c_688_n 4.84884e-19 $X=4.355 $Y=1.275 $X2=0 $Y2=0
cc_242 N_A2_c_241_n N_VGND_c_689_n 0.00414769f $X=3.895 $Y=1.275 $X2=0 $Y2=0
cc_243 N_A2_c_243_n N_VGND_c_690_n 0.00499542f $X=4.355 $Y=1.275 $X2=0 $Y2=0
cc_244 N_A2_c_241_n N_VGND_c_692_n 0.00789406f $X=3.895 $Y=1.275 $X2=0 $Y2=0
cc_245 N_A2_c_243_n N_VGND_c_692_n 0.00973406f $X=4.355 $Y=1.275 $X2=0 $Y2=0
cc_246 N_A2_c_241_n N_VGND_c_694_n 4.43819e-19 $X=3.895 $Y=1.275 $X2=0 $Y2=0
cc_247 N_A1_M1000_g N_VPWR_c_452_n 0.0166795f $X=5.195 $Y=2.465 $X2=0 $Y2=0
cc_248 N_A1_M1009_g N_VPWR_c_452_n 7.55536e-19 $X=5.625 $Y=2.465 $X2=0 $Y2=0
cc_249 N_A1_M1009_g N_VPWR_c_454_n 0.00768161f $X=5.625 $Y=2.465 $X2=0 $Y2=0
cc_250 A1 N_VPWR_c_454_n 0.0178016f $X=5.915 $Y=1.21 $X2=0 $Y2=0
cc_251 N_A1_M1000_g N_VPWR_c_457_n 0.00486043f $X=5.195 $Y=2.465 $X2=0 $Y2=0
cc_252 N_A1_M1009_g N_VPWR_c_457_n 0.00585385f $X=5.625 $Y=2.465 $X2=0 $Y2=0
cc_253 N_A1_M1000_g N_VPWR_c_450_n 0.00824727f $X=5.195 $Y=2.465 $X2=0 $Y2=0
cc_254 N_A1_M1009_g N_VPWR_c_450_n 0.0115632f $X=5.625 $Y=2.465 $X2=0 $Y2=0
cc_255 N_A1_M1000_g N_A_519_365#_c_529_n 0.00135858f $X=5.195 $Y=2.465 $X2=0
+ $Y2=0
cc_256 N_A1_M1000_g N_A_778_365#_c_567_n 0.0156548f $X=5.195 $Y=2.465 $X2=0
+ $Y2=0
cc_257 N_A1_M1009_g N_A_778_365#_c_567_n 0.0038539f $X=5.625 $Y=2.465 $X2=0
+ $Y2=0
cc_258 A1 N_A_778_365#_c_567_n 0.0533824f $X=5.915 $Y=1.21 $X2=0 $Y2=0
cc_259 N_A1_c_300_n N_A_778_365#_c_567_n 0.0144802f $X=5.625 $Y=1.44 $X2=0 $Y2=0
cc_260 N_A1_c_295_n N_A_39_65#_c_603_n 4.34728e-19 $X=4.785 $Y=1.275 $X2=0 $Y2=0
cc_261 N_A1_c_295_n N_A_39_65#_c_633_n 0.0134128f $X=4.785 $Y=1.275 $X2=0 $Y2=0
cc_262 N_A1_c_297_n N_A_39_65#_c_633_n 0.0120955f $X=5.215 $Y=1.275 $X2=0 $Y2=0
cc_263 A1 N_A_39_65#_c_633_n 0.0333046f $X=5.915 $Y=1.21 $X2=0 $Y2=0
cc_264 N_A1_c_300_n N_A_39_65#_c_633_n 5.92586e-19 $X=5.625 $Y=1.44 $X2=0 $Y2=0
cc_265 A1 N_A_39_65#_c_604_n 0.0219949f $X=5.915 $Y=1.21 $X2=0 $Y2=0
cc_266 N_A1_c_300_n N_A_39_65#_c_604_n 0.00169421f $X=5.625 $Y=1.44 $X2=0 $Y2=0
cc_267 N_A1_c_297_n N_A_39_65#_c_605_n 0.00186805f $X=5.215 $Y=1.275 $X2=0 $Y2=0
cc_268 N_A1_c_295_n N_VGND_c_688_n 0.00885412f $X=4.785 $Y=1.275 $X2=0 $Y2=0
cc_269 N_A1_c_297_n N_VGND_c_688_n 0.0112436f $X=5.215 $Y=1.275 $X2=0 $Y2=0
cc_270 N_A1_c_295_n N_VGND_c_690_n 0.00414769f $X=4.785 $Y=1.275 $X2=0 $Y2=0
cc_271 N_A1_c_297_n N_VGND_c_691_n 0.00414769f $X=5.215 $Y=1.275 $X2=0 $Y2=0
cc_272 N_A1_c_295_n N_VGND_c_692_n 0.0078848f $X=4.785 $Y=1.275 $X2=0 $Y2=0
cc_273 N_A1_c_297_n N_VGND_c_692_n 0.00837493f $X=5.215 $Y=1.275 $X2=0 $Y2=0
cc_274 N_A_39_367#_c_339_n N_Y_M1005_s 0.00332344f $X=1.085 $Y=2.99 $X2=0 $Y2=0
cc_275 N_A_39_367#_M1015_d N_Y_c_370_n 0.00353353f $X=1.04 $Y=1.835 $X2=0 $Y2=0
cc_276 N_A_39_367#_M1016_d N_Y_c_370_n 0.00526039f $X=1.9 $Y=1.835 $X2=0 $Y2=0
cc_277 N_A_39_367#_c_346_p N_Y_c_370_n 0.0135055f $X=1.18 $Y=2.45 $X2=0 $Y2=0
cc_278 N_A_39_367#_c_341_n N_Y_c_370_n 0.0325992f $X=1.945 $Y=2.355 $X2=0 $Y2=0
cc_279 N_A_39_367#_c_336_n N_Y_c_370_n 0.020301f $X=2.075 $Y=2.45 $X2=0 $Y2=0
cc_280 N_A_39_367#_c_339_n N_Y_c_381_n 0.0159805f $X=1.085 $Y=2.99 $X2=0 $Y2=0
cc_281 N_A_39_367#_c_341_n N_VPWR_M1008_s 0.00345035f $X=1.945 $Y=2.355
+ $X2=-0.19 $Y2=1.655
cc_282 N_A_39_367#_c_341_n N_VPWR_c_451_n 0.0172078f $X=1.945 $Y=2.355 $X2=0
+ $Y2=0
cc_283 N_A_39_367#_c_334_n N_VPWR_c_455_n 0.0179183f $X=0.285 $Y=2.905 $X2=0
+ $Y2=0
cc_284 N_A_39_367#_c_339_n N_VPWR_c_455_n 0.0486406f $X=1.085 $Y=2.99 $X2=0
+ $Y2=0
cc_285 N_A_39_367#_c_337_n N_VPWR_c_456_n 0.0178111f $X=2.04 $Y=2.91 $X2=0 $Y2=0
cc_286 N_A_39_367#_M1005_d N_VPWR_c_450_n 0.00215161f $X=0.195 $Y=1.835 $X2=0
+ $Y2=0
cc_287 N_A_39_367#_M1015_d N_VPWR_c_450_n 0.00376627f $X=1.04 $Y=1.835 $X2=0
+ $Y2=0
cc_288 N_A_39_367#_M1016_d N_VPWR_c_450_n 0.00371702f $X=1.9 $Y=1.835 $X2=0
+ $Y2=0
cc_289 N_A_39_367#_c_334_n N_VPWR_c_450_n 0.0101029f $X=0.285 $Y=2.905 $X2=0
+ $Y2=0
cc_290 N_A_39_367#_c_339_n N_VPWR_c_450_n 0.0310628f $X=1.085 $Y=2.99 $X2=0
+ $Y2=0
cc_291 N_A_39_367#_c_337_n N_VPWR_c_450_n 0.0100304f $X=2.04 $Y=2.91 $X2=0 $Y2=0
cc_292 N_A_39_367#_c_336_n N_A_519_365#_c_525_n 0.0100342f $X=2.075 $Y=2.45
+ $X2=0 $Y2=0
cc_293 N_A_39_367#_c_337_n N_A_519_365#_c_525_n 0.0221938f $X=2.04 $Y=2.91 $X2=0
+ $Y2=0
cc_294 N_A_39_367#_c_337_n N_A_519_365#_c_526_n 0.00895419f $X=2.04 $Y=2.91
+ $X2=0 $Y2=0
cc_295 N_Y_c_370_n N_VPWR_M1008_s 0.00332905f $X=3.005 $Y=2.005 $X2=-0.19
+ $Y2=-0.245
cc_296 N_Y_M1005_s N_VPWR_c_450_n 0.00225186f $X=0.61 $Y=1.835 $X2=0 $Y2=0
cc_297 N_Y_M1011_s N_VPWR_c_450_n 0.00225186f $X=3.03 $Y=1.825 $X2=0 $Y2=0
cc_298 N_Y_c_370_n N_A_519_365#_M1011_d 0.00536966f $X=3.005 $Y=2.005 $X2=-0.19
+ $Y2=-0.245
cc_299 N_Y_c_370_n N_A_519_365#_c_525_n 0.0218437f $X=3.005 $Y=2.005 $X2=0 $Y2=0
cc_300 N_Y_M1011_s N_A_519_365#_c_530_n 0.00332344f $X=3.03 $Y=1.825 $X2=0 $Y2=0
cc_301 Y N_A_519_365#_c_530_n 0.0159805f $X=3.035 $Y=1.95 $X2=0 $Y2=0
cc_302 Y N_A_519_365#_c_527_n 0.00424671f $X=3.12 $Y=1.295 $X2=0 $Y2=0
cc_303 Y N_A_778_365#_c_568_n 0.00344926f $X=3.12 $Y=1.295 $X2=0 $Y2=0
cc_304 N_Y_c_364_n N_A_39_65#_M1019_d 0.00261503f $X=1.605 $Y=1.16 $X2=0 $Y2=0
cc_305 N_Y_c_366_n N_A_39_65#_M1012_s 0.00261503f $X=3.005 $Y=1.16 $X2=0 $Y2=0
cc_306 N_Y_c_365_n N_A_39_65#_c_598_n 0.00539933f $X=0.915 $Y=1.16 $X2=0 $Y2=0
cc_307 N_Y_M1004_s N_A_39_65#_c_599_n 0.00176461f $X=0.61 $Y=0.325 $X2=0 $Y2=0
cc_308 N_Y_c_371_n N_A_39_65#_c_599_n 0.0159249f $X=0.75 $Y=0.68 $X2=0 $Y2=0
cc_309 N_Y_c_364_n N_A_39_65#_c_599_n 0.00275981f $X=1.605 $Y=1.16 $X2=0 $Y2=0
cc_310 N_Y_c_364_n N_A_39_65#_c_611_n 0.02172f $X=1.605 $Y=1.16 $X2=0 $Y2=0
cc_311 N_Y_M1006_d N_A_39_65#_c_601_n 0.00261503f $X=1.55 $Y=0.325 $X2=0 $Y2=0
cc_312 N_Y_c_364_n N_A_39_65#_c_601_n 0.00275981f $X=1.605 $Y=1.16 $X2=0 $Y2=0
cc_313 N_Y_c_393_n N_A_39_65#_c_601_n 0.0203258f $X=1.77 $Y=0.68 $X2=0 $Y2=0
cc_314 N_Y_c_366_n N_A_39_65#_c_601_n 0.00275981f $X=3.005 $Y=1.16 $X2=0 $Y2=0
cc_315 N_Y_c_366_n N_A_39_65#_c_618_n 0.0358577f $X=3.005 $Y=1.16 $X2=0 $Y2=0
cc_316 N_Y_c_368_n N_A_39_65#_c_618_n 0.025872f $X=3.17 $Y=1.245 $X2=0 $Y2=0
cc_317 N_Y_c_366_n N_A_39_65#_c_621_n 0.0217959f $X=3.005 $Y=1.16 $X2=0 $Y2=0
cc_318 N_Y_c_366_n N_VGND_M1007_s 0.00517008f $X=3.005 $Y=1.16 $X2=-0.19
+ $Y2=-0.245
cc_319 N_Y_c_368_n N_VGND_M1007_s 0.00487456f $X=3.17 $Y=1.245 $X2=-0.19
+ $Y2=-0.245
cc_320 N_VPWR_c_450_n N_A_519_365#_M1011_d 0.00228387f $X=6 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_321 N_VPWR_c_450_n N_A_519_365#_M1017_d 0.00223565f $X=6 $Y=3.33 $X2=0 $Y2=0
cc_322 N_VPWR_c_450_n N_A_519_365#_M1014_s 0.00212303f $X=6 $Y=3.33 $X2=0 $Y2=0
cc_323 N_VPWR_c_456_n N_A_519_365#_c_530_n 0.0364699f $X=4.815 $Y=3.33 $X2=0
+ $Y2=0
cc_324 N_VPWR_c_450_n N_A_519_365#_c_530_n 0.024052f $X=6 $Y=3.33 $X2=0 $Y2=0
cc_325 N_VPWR_c_456_n N_A_519_365#_c_526_n 0.0189697f $X=4.815 $Y=3.33 $X2=0
+ $Y2=0
cc_326 N_VPWR_c_450_n N_A_519_365#_c_526_n 0.0104864f $X=6 $Y=3.33 $X2=0 $Y2=0
cc_327 N_VPWR_c_456_n N_A_519_365#_c_536_n 0.0361172f $X=4.815 $Y=3.33 $X2=0
+ $Y2=0
cc_328 N_VPWR_c_450_n N_A_519_365#_c_536_n 0.023676f $X=6 $Y=3.33 $X2=0 $Y2=0
cc_329 N_VPWR_c_452_n N_A_519_365#_c_528_n 0.0139f $X=4.98 $Y=2.13 $X2=0 $Y2=0
cc_330 N_VPWR_c_456_n N_A_519_365#_c_528_n 0.0179183f $X=4.815 $Y=3.33 $X2=0
+ $Y2=0
cc_331 N_VPWR_c_450_n N_A_519_365#_c_528_n 0.0101082f $X=6 $Y=3.33 $X2=0 $Y2=0
cc_332 N_VPWR_c_452_n N_A_519_365#_c_529_n 0.0650111f $X=4.98 $Y=2.13 $X2=0
+ $Y2=0
cc_333 N_VPWR_c_456_n N_A_519_365#_c_560_n 0.0125234f $X=4.815 $Y=3.33 $X2=0
+ $Y2=0
cc_334 N_VPWR_c_450_n N_A_519_365#_c_560_n 0.0073762f $X=6 $Y=3.33 $X2=0 $Y2=0
cc_335 N_VPWR_c_450_n N_A_778_365#_M1003_d 0.00225186f $X=6 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_336 N_VPWR_c_450_n N_A_778_365#_M1000_s 0.0041489f $X=6 $Y=3.33 $X2=0 $Y2=0
cc_337 N_VPWR_M1000_d N_A_778_365#_c_567_n 0.00239457f $X=4.855 $Y=1.835 $X2=0
+ $Y2=0
cc_338 N_VPWR_c_452_n N_A_778_365#_c_567_n 0.0220025f $X=4.98 $Y=2.13 $X2=0
+ $Y2=0
cc_339 N_VPWR_c_454_n N_A_778_365#_c_567_n 0.00166618f $X=5.84 $Y=1.98 $X2=0
+ $Y2=0
cc_340 N_VPWR_c_457_n N_A_778_365#_c_589_n 0.0136943f $X=5.71 $Y=3.33 $X2=0
+ $Y2=0
cc_341 N_VPWR_c_450_n N_A_778_365#_c_589_n 0.00866972f $X=6 $Y=3.33 $X2=0 $Y2=0
cc_342 N_A_519_365#_c_536_n N_A_778_365#_M1003_d 0.00332344f $X=4.365 $Y=2.99
+ $X2=-0.19 $Y2=1.655
cc_343 N_A_519_365#_c_536_n N_A_778_365#_c_570_n 0.0159805f $X=4.365 $Y=2.99
+ $X2=0 $Y2=0
cc_344 N_A_519_365#_M1014_s N_A_778_365#_c_567_n 0.00244161f $X=4.32 $Y=1.825
+ $X2=0 $Y2=0
cc_345 N_A_519_365#_c_529_n N_A_778_365#_c_567_n 0.0202165f $X=4.46 $Y=2.21
+ $X2=0 $Y2=0
cc_346 N_A_519_365#_c_527_n N_A_778_365#_c_568_n 0.00287328f $X=3.6 $Y=1.98
+ $X2=0 $Y2=0
cc_347 N_A_778_365#_c_567_n N_A_39_65#_c_633_n 0.00327684f $X=5.315 $Y=1.79
+ $X2=0 $Y2=0
cc_348 N_A_778_365#_c_567_n N_A_39_65#_c_631_n 4.19026e-19 $X=5.315 $Y=1.79
+ $X2=0 $Y2=0
cc_349 N_A_39_65#_c_618_n N_VGND_M1007_s 0.0179394f $X=3.505 $Y=0.82 $X2=-0.19
+ $Y2=-0.245
cc_350 N_A_39_65#_c_625_n N_VGND_M1002_d 0.00390103f $X=4.465 $Y=0.955 $X2=0
+ $Y2=0
cc_351 N_A_39_65#_c_633_n N_VGND_M1001_d 0.003325f $X=5.335 $Y=0.955 $X2=0 $Y2=0
cc_352 N_A_39_65#_c_602_n N_VGND_c_687_n 0.0147932f $X=3.67 $Y=0.48 $X2=0 $Y2=0
cc_353 N_A_39_65#_c_625_n N_VGND_c_687_n 0.0177324f $X=4.465 $Y=0.955 $X2=0
+ $Y2=0
cc_354 N_A_39_65#_c_603_n N_VGND_c_687_n 6.67084e-19 $X=4.57 $Y=0.48 $X2=0 $Y2=0
cc_355 N_A_39_65#_c_603_n N_VGND_c_688_n 0.0147932f $X=4.57 $Y=0.48 $X2=0 $Y2=0
cc_356 N_A_39_65#_c_633_n N_VGND_c_688_n 0.0170777f $X=5.335 $Y=0.955 $X2=0
+ $Y2=0
cc_357 N_A_39_65#_c_605_n N_VGND_c_688_n 0.0148073f $X=5.43 $Y=0.48 $X2=0 $Y2=0
cc_358 N_A_39_65#_c_618_n N_VGND_c_689_n 0.0013004f $X=3.505 $Y=0.82 $X2=0 $Y2=0
cc_359 N_A_39_65#_c_602_n N_VGND_c_689_n 0.0102728f $X=3.67 $Y=0.48 $X2=0 $Y2=0
cc_360 N_A_39_65#_c_623_n N_VGND_c_689_n 6.68265e-19 $X=3.64 $Y=0.82 $X2=0 $Y2=0
cc_361 N_A_39_65#_c_603_n N_VGND_c_690_n 0.0102728f $X=4.57 $Y=0.48 $X2=0 $Y2=0
cc_362 N_A_39_65#_c_605_n N_VGND_c_691_n 0.0133857f $X=5.43 $Y=0.48 $X2=0 $Y2=0
cc_363 N_A_39_65#_c_599_n N_VGND_c_692_n 0.0241933f $X=1.095 $Y=0.34 $X2=0 $Y2=0
cc_364 N_A_39_65#_c_600_n N_VGND_c_692_n 0.0101082f $X=0.415 $Y=0.34 $X2=0 $Y2=0
cc_365 N_A_39_65#_c_601_n N_VGND_c_692_n 0.0373836f $X=2.115 $Y=0.34 $X2=0 $Y2=0
cc_366 N_A_39_65#_c_618_n N_VGND_c_692_n 0.00898798f $X=3.505 $Y=0.82 $X2=0
+ $Y2=0
cc_367 N_A_39_65#_c_602_n N_VGND_c_692_n 0.00746302f $X=3.67 $Y=0.48 $X2=0 $Y2=0
cc_368 N_A_39_65#_c_603_n N_VGND_c_692_n 0.00746302f $X=4.57 $Y=0.48 $X2=0 $Y2=0
cc_369 N_A_39_65#_c_605_n N_VGND_c_692_n 0.00972454f $X=5.43 $Y=0.48 $X2=0 $Y2=0
cc_370 N_A_39_65#_c_606_n N_VGND_c_692_n 0.0127001f $X=1.26 $Y=0.34 $X2=0 $Y2=0
cc_371 N_A_39_65#_c_623_n N_VGND_c_692_n 0.00175095f $X=3.64 $Y=0.82 $X2=0 $Y2=0
cc_372 N_A_39_65#_c_599_n N_VGND_c_693_n 0.0428729f $X=1.095 $Y=0.34 $X2=0 $Y2=0
cc_373 N_A_39_65#_c_600_n N_VGND_c_693_n 0.0186386f $X=0.415 $Y=0.34 $X2=0 $Y2=0
cc_374 N_A_39_65#_c_601_n N_VGND_c_693_n 0.0670812f $X=2.115 $Y=0.34 $X2=0 $Y2=0
cc_375 N_A_39_65#_c_618_n N_VGND_c_693_n 0.00196209f $X=3.505 $Y=0.82 $X2=0
+ $Y2=0
cc_376 N_A_39_65#_c_606_n N_VGND_c_693_n 0.023489f $X=1.26 $Y=0.34 $X2=0 $Y2=0
cc_377 N_A_39_65#_c_601_n N_VGND_c_694_n 0.0104256f $X=2.115 $Y=0.34 $X2=0 $Y2=0
cc_378 N_A_39_65#_c_618_n N_VGND_c_694_n 0.0560848f $X=3.505 $Y=0.82 $X2=0 $Y2=0
cc_379 N_A_39_65#_c_602_n N_VGND_c_694_n 0.0108374f $X=3.67 $Y=0.48 $X2=0 $Y2=0
