* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__sdfbbp_1 CLK D RESET_B SCD SCE SET_B VNB VPB Q Q_N
X0 a_290_119# a_332_93# VNB SUBS sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 VPB SET_B a_2064_453# w_n38_331# sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X2 VNB a_2064_453# Q_N SUBS sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X3 a_204_119# a_755_106# a_1216_457# SUBS sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 VPB SCE a_224_481# w_n38_331# sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X5 a_1302_457# a_1297_290# VPB w_n38_331# sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X6 a_1650_21# RESET_B VNB SUBS sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 VPB a_2892_137# Q w_n38_331# sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X8 a_204_119# D a_290_119# SUBS sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 a_27_481# SCD VPB w_n38_331# sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X10 a_2395_451# a_1650_21# VPB w_n38_331# sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X11 a_1318_47# a_1297_290# VNB SUBS sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 VNB SET_B a_2279_57# SUBS sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X13 a_204_119# a_893_101# a_1216_457# w_n38_331# sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X14 a_2279_57# a_1861_431# a_2064_453# SUBS sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X15 VNB SET_B a_1492_47# SUBS sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X16 VNB a_2892_137# Q SUBS sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X17 a_2064_453# a_1861_431# a_2395_451# w_n38_331# sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X18 a_893_101# a_755_106# VNB SUBS sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X19 a_1650_21# RESET_B VPB w_n38_331# sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X20 VPB SCE a_332_93# w_n38_331# sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X21 VPB SET_B a_1297_290# w_n38_331# sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X22 a_1963_515# a_2064_453# VPB w_n38_331# sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X23 VNB CLK a_755_106# SUBS sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X24 a_1880_57# a_893_101# a_1861_431# SUBS sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X25 a_1297_290# a_1650_21# a_1492_47# SUBS sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X26 VPB CLK a_755_106# w_n38_331# sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X27 a_1216_457# a_755_106# a_1302_457# w_n38_331# sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X28 a_1766_373# a_755_106# a_1861_431# w_n38_331# sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X29 VNB a_1297_290# a_1880_57# SUBS sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X30 a_1861_431# a_755_106# a_2066_101# SUBS sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X31 VNB SCD a_126_119# SUBS sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X32 a_1492_47# a_1216_457# a_1297_290# SUBS sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X33 a_2064_453# a_1650_21# a_2279_57# SUBS sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X34 a_893_101# a_755_106# VPB w_n38_331# sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X35 a_1297_290# a_1216_457# a_1584_373# w_n38_331# sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X36 VPB a_1297_290# a_1766_373# w_n38_331# sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X37 a_2892_137# a_2064_453# VNB SUBS sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X38 a_204_119# a_332_93# a_27_481# w_n38_331# sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X39 a_1584_373# a_1650_21# VPB w_n38_331# sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X40 a_224_481# D a_204_119# w_n38_331# sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X41 a_2892_137# a_2064_453# VPB w_n38_331# sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X42 a_2066_101# a_2064_453# VNB SUBS sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X43 a_1216_457# a_893_101# a_1318_47# SUBS sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X44 a_126_119# SCE a_204_119# SUBS sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X45 VNB SCE a_332_93# SUBS sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X46 a_1861_431# a_893_101# a_1963_515# w_n38_331# sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X47 VPB a_2064_453# Q_N w_n38_331# sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
.ends
