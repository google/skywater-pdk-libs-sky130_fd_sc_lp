* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__or4b_lp A B C D_N VGND VNB VPB VPWR X
X0 VPWR a_311_417# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X1 a_270_57# a_27_57# a_311_417# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 a_311_417# a_27_57# a_422_417# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X3 a_586_57# B a_311_417# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 a_311_417# A a_744_57# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 a_428_57# C VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 a_422_417# C a_520_417# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X7 a_744_57# A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 VGND a_311_417# a_902_57# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 a_112_57# D_N VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 a_27_57# D_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X11 a_27_57# D_N a_112_57# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 VGND a_27_57# a_270_57# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X13 a_520_417# B a_634_417# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X14 VGND B a_586_57# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X15 a_311_417# C a_428_57# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X16 a_634_417# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X17 a_902_57# a_311_417# X VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
