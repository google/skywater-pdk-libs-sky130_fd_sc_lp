# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_sc_lp__srsdfstp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_lp__srsdfstp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  18.72000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.085000 1.545000 1.430000 1.875000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.573300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 18.365000 0.255000 18.620000 3.075000 ;
    END
  END Q
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.205000 0.835000 1.875000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.725000 1.180000 3.235000 1.555000 ;
    END
  END SCE
  PIN SET_B
    ANTENNAGATEAREA  0.439000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 13.500000 1.580000 13.830000 1.840000 ;
    END
  END SET_B
  PIN SLEEP_B
    ANTENNAGATEAREA  0.598000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 15.935000 1.220000 16.260000 2.150000 ;
    END
  END SLEEP_B
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 14.965000 1.180000 15.235000 2.150000 ;
    END
  END CLK
  PIN KAPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.070000 2.675000 18.650000 2.945000 ;
    END
  END KAPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 18.720000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.000000 0.000000 18.720000 0.245000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.655000 18.910000 3.520000 ;
        RECT  2.245000 1.565000  4.025000 1.655000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 18.720000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 18.720000 0.085000 ;
      RECT  0.000000  3.245000 18.720000 3.415000 ;
      RECT  0.100000  0.085000  0.430000 1.035000 ;
      RECT  0.100000  2.045000  1.190000 2.215000 ;
      RECT  0.100000  2.215000  0.430000 3.065000 ;
      RECT  0.600000  2.385000  0.850000 3.245000 ;
      RECT  0.920000  0.575000  1.250000 0.865000 ;
      RECT  0.920000  0.865000  1.770000 1.035000 ;
      RECT  1.020000  2.215000  1.190000 2.905000 ;
      RECT  1.020000  2.905000  2.190000 3.075000 ;
      RECT  1.430000  2.225000  3.835000 2.395000 ;
      RECT  1.430000  2.395000  1.770000 2.735000 ;
      RECT  1.600000  1.035000  1.770000 2.225000 ;
      RECT  1.940000  0.085000  2.190000 1.035000 ;
      RECT  1.940000  1.305000  2.555000 1.725000 ;
      RECT  1.940000  1.725000  2.720000 2.055000 ;
      RECT  1.940000  2.565000  2.190000 2.905000 ;
      RECT  2.385000  0.675000  2.740000 1.010000 ;
      RECT  2.385000  1.010000  2.555000 1.305000 ;
      RECT  2.920000  0.085000  3.250000 1.010000 ;
      RECT  2.920000  2.565000  3.250000 3.245000 ;
      RECT  3.420000  0.255000  5.280000 0.425000 ;
      RECT  3.420000  0.425000  4.015000 0.585000 ;
      RECT  3.420000  0.585000  3.750000 1.725000 ;
      RECT  3.420000  1.725000  4.260000 2.055000 ;
      RECT  3.665000  2.395000  3.835000 2.655000 ;
      RECT  3.665000  2.655000  5.035000 2.825000 ;
      RECT  3.980000  0.755000  4.230000 1.385000 ;
      RECT  3.980000  1.385000  4.600000 1.555000 ;
      RECT  4.005000  2.055000  4.260000 2.395000 ;
      RECT  4.410000  0.675000  4.940000 1.135000 ;
      RECT  4.430000  1.555000  4.600000 2.655000 ;
      RECT  4.600000  2.825000  5.035000 3.075000 ;
      RECT  4.770000  1.135000  4.940000 1.905000 ;
      RECT  4.770000  1.905000  7.675000 2.075000 ;
      RECT  5.110000  0.425000  5.280000 1.545000 ;
      RECT  5.110000  1.545000  8.015000 1.640000 ;
      RECT  5.110000  1.640000  6.120000 1.715000 ;
      RECT  5.205000  2.075000  5.535000 3.075000 ;
      RECT  5.450000  0.675000  6.135000 0.845000 ;
      RECT  5.450000  0.845000  5.780000 1.375000 ;
      RECT  5.465000  0.085000  5.795000 0.505000 ;
      RECT  5.900000  2.245000  6.230000 2.265000 ;
      RECT  5.900000  2.265000  7.010000 2.485000 ;
      RECT  5.950000  1.470000  8.015000 1.545000 ;
      RECT  5.965000  0.255000  6.895000 0.425000 ;
      RECT  5.965000  0.425000  6.135000 0.675000 ;
      RECT  5.990000  1.015000  6.555000 1.300000 ;
      RECT  6.025000  2.655000  6.355000 3.245000 ;
      RECT  6.305000  0.595000  6.555000 1.015000 ;
      RECT  6.440000  1.810000  7.675000 1.905000 ;
      RECT  6.440000  2.075000  7.675000 2.095000 ;
      RECT  6.680000  2.485000  7.010000 2.695000 ;
      RECT  6.725000  0.425000  6.895000 1.130000 ;
      RECT  6.725000  1.130000  7.705000 1.300000 ;
      RECT  7.115000  0.085000  7.365000 0.960000 ;
      RECT  7.250000  2.265000  7.580000 3.245000 ;
      RECT  7.535000  0.255000 10.255000 0.425000 ;
      RECT  7.535000  0.425000  7.705000 1.130000 ;
      RECT  7.755000  2.905000  8.695000 3.075000 ;
      RECT  7.845000  1.640000  8.015000 2.905000 ;
      RECT  7.875000  0.595000  8.145000 1.095000 ;
      RECT  7.875000  1.095000  8.355000 1.265000 ;
      RECT  8.185000  1.265000  8.355000 2.565000 ;
      RECT  8.525000  0.595000  9.535000 0.765000 ;
      RECT  8.525000  0.765000  8.695000 1.410000 ;
      RECT  8.525000  1.410000  8.755000 1.740000 ;
      RECT  8.525000  1.740000  8.695000 2.905000 ;
      RECT  8.865000  0.935000  9.195000 1.225000 ;
      RECT  8.895000  2.235000  9.145000 2.745000 ;
      RECT  8.925000  1.225000  9.095000 2.235000 ;
      RECT  8.940000  2.745000 12.485000 3.075000 ;
      RECT  9.315000  1.885000  9.535000 2.135000 ;
      RECT  9.315000  2.135000  9.485000 2.405000 ;
      RECT  9.315000  2.405000 12.145000 2.575000 ;
      RECT  9.365000  0.765000  9.535000 1.885000 ;
      RECT 10.085000  0.425000 10.255000 1.545000 ;
      RECT 10.085000  1.545000 12.675000 1.715000 ;
      RECT 10.165000  1.715000 10.415000 2.145000 ;
      RECT 10.425000  0.605000 10.595000 1.205000 ;
      RECT 10.425000  1.205000 11.455000 1.375000 ;
      RECT 10.655000  1.885000 13.015000 2.055000 ;
      RECT 10.655000  2.055000 10.985000 2.215000 ;
      RECT 10.775000  0.085000 11.025000 1.035000 ;
      RECT 11.205000  0.605000 11.455000 1.205000 ;
      RECT 11.475000  2.055000 11.805000 2.235000 ;
      RECT 11.625000  1.125000 12.335000 1.375000 ;
      RECT 11.745000  0.085000 11.995000 0.955000 ;
      RECT 11.975000  2.225000 13.355000 2.395000 ;
      RECT 11.975000  2.395000 12.145000 2.405000 ;
      RECT 12.165000  0.255000 15.915000 0.425000 ;
      RECT 12.165000  0.425000 12.335000 1.125000 ;
      RECT 12.315000  2.565000 14.130000 2.735000 ;
      RECT 12.315000  2.735000 12.485000 2.745000 ;
      RECT 12.505000  0.595000 13.355000 0.765000 ;
      RECT 12.505000  0.765000 12.675000 1.545000 ;
      RECT 12.655000  2.905000 15.235000 3.075000 ;
      RECT 12.845000  0.935000 13.015000 1.240000 ;
      RECT 12.845000  1.240000 14.755000 1.410000 ;
      RECT 12.845000  1.410000 13.015000 1.885000 ;
      RECT 13.185000  0.765000 13.355000 0.900000 ;
      RECT 13.185000  0.900000 14.255000 1.070000 ;
      RECT 13.185000  2.010000 14.210000 2.180000 ;
      RECT 13.185000  2.180000 13.355000 2.225000 ;
      RECT 13.525000  0.425000 13.855000 0.730000 ;
      RECT 13.800000  2.350000 17.220000 2.490000 ;
      RECT 13.800000  2.490000 14.595000 2.520000 ;
      RECT 13.800000  2.520000 14.130000 2.565000 ;
      RECT 14.040000  1.580000 14.370000 1.910000 ;
      RECT 14.040000  1.910000 14.210000 2.010000 ;
      RECT 14.085000  0.595000 15.575000 0.845000 ;
      RECT 14.085000  0.845000 14.255000 0.900000 ;
      RECT 14.425000  1.040000 14.755000 1.240000 ;
      RECT 14.425000  2.320000 17.220000 2.350000 ;
      RECT 14.905000  2.660000 15.235000 2.905000 ;
      RECT 15.405000  0.845000 15.575000 1.900000 ;
      RECT 15.405000  1.900000 15.765000 2.150000 ;
      RECT 15.745000  0.425000 15.915000 0.880000 ;
      RECT 15.745000  0.880000 16.835000 1.050000 ;
      RECT 15.965000  2.660000 16.305000 2.940000 ;
      RECT 16.085000  0.085000 16.335000 0.710000 ;
      RECT 16.455000  1.050000 16.835000 2.150000 ;
      RECT 16.665000  0.630000 17.125000 0.800000 ;
      RECT 16.665000  0.800000 16.835000 0.880000 ;
      RECT 16.795000  0.420000 17.125000 0.630000 ;
      RECT 17.005000  1.495000 17.335000 1.825000 ;
      RECT 17.050000  1.825000 17.220000 2.320000 ;
      RECT 17.325000  0.295000 17.675000 0.675000 ;
      RECT 17.390000  1.995000 17.675000 2.675000 ;
      RECT 17.505000  0.675000 17.675000 1.185000 ;
      RECT 17.505000  1.185000 18.195000 1.515000 ;
      RECT 17.505000  1.515000 17.675000 1.995000 ;
      RECT 17.855000  1.815000 18.185000 3.245000 ;
      RECT 17.860000  0.085000 18.190000 1.015000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.245000 10.885000 3.415000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  3.245000 11.365000 3.415000 ;
      RECT 11.675000 -0.085000 11.845000 0.085000 ;
      RECT 11.675000  3.245000 11.845000 3.415000 ;
      RECT 12.155000 -0.085000 12.325000 0.085000 ;
      RECT 12.155000  3.245000 12.325000 3.415000 ;
      RECT 12.635000 -0.085000 12.805000 0.085000 ;
      RECT 12.635000  3.245000 12.805000 3.415000 ;
      RECT 13.115000 -0.085000 13.285000 0.085000 ;
      RECT 13.115000  3.245000 13.285000 3.415000 ;
      RECT 13.595000 -0.085000 13.765000 0.085000 ;
      RECT 13.595000  3.245000 13.765000 3.415000 ;
      RECT 14.075000 -0.085000 14.245000 0.085000 ;
      RECT 14.075000  3.245000 14.245000 3.415000 ;
      RECT 14.555000 -0.085000 14.725000 0.085000 ;
      RECT 14.555000  3.245000 14.725000 3.415000 ;
      RECT 15.035000 -0.085000 15.205000 0.085000 ;
      RECT 15.035000  2.735000 15.205000 2.905000 ;
      RECT 15.035000  3.245000 15.205000 3.415000 ;
      RECT 15.515000 -0.085000 15.685000 0.085000 ;
      RECT 15.515000  3.245000 15.685000 3.415000 ;
      RECT 15.995000 -0.085000 16.165000 0.085000 ;
      RECT 15.995000  2.735000 16.165000 2.905000 ;
      RECT 15.995000  3.245000 16.165000 3.415000 ;
      RECT 16.475000 -0.085000 16.645000 0.085000 ;
      RECT 16.475000  3.245000 16.645000 3.415000 ;
      RECT 16.955000 -0.085000 17.125000 0.085000 ;
      RECT 16.955000  3.245000 17.125000 3.415000 ;
      RECT 17.435000 -0.085000 17.605000 0.085000 ;
      RECT 17.435000  3.245000 17.605000 3.415000 ;
      RECT 17.915000 -0.085000 18.085000 0.085000 ;
      RECT 17.915000  3.245000 18.085000 3.415000 ;
      RECT 18.395000 -0.085000 18.565000 0.085000 ;
      RECT 18.395000  3.245000 18.565000 3.415000 ;
  END
END sky130_fd_sc_lp__srsdfstp_1
END LIBRARY
