* File: sky130_fd_sc_lp__a21o_m.pex.spice
* Created: Wed Sep  2 09:20:20 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A21O_M%A_80_153# 1 2 10 13 15 17 20 22 26 27 28 29
+ 30 31 34 38 41
r73 36 38 19.2771 $w=2.08e-07 $l=3.65e-07 $layer=LI1_cond $X=1.39 $Y=0.86
+ $X2=1.39 $Y2=0.495
r74 32 34 8.97835 $w=2.08e-07 $l=1.7e-07 $layer=LI1_cond $X=1.33 $Y=2.515
+ $X2=1.33 $Y2=2.685
r75 30 32 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=1.225 $Y=2.43
+ $X2=1.33 $Y2=2.515
r76 30 31 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=1.225 $Y=2.43
+ $X2=0.695 $Y2=2.43
r77 28 36 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=1.285 $Y=0.945
+ $X2=1.39 $Y2=0.86
r78 28 29 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=1.285 $Y=0.945
+ $X2=0.695 $Y2=0.945
r79 27 41 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=0.587 $Y=2.01
+ $X2=0.587 $Y2=1.845
r80 26 27 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.61
+ $Y=2.01 $X2=0.61 $Y2=2.01
r81 24 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.61 $Y=2.345
+ $X2=0.695 $Y2=2.43
r82 24 26 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=0.61 $Y=2.345
+ $X2=0.61 $Y2=2.01
r83 23 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.61 $Y=1.03
+ $X2=0.695 $Y2=0.945
r84 23 26 63.9358 $w=1.68e-07 $l=9.8e-07 $layer=LI1_cond $X=0.61 $Y=1.03
+ $X2=0.61 $Y2=2.01
r85 18 20 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=0.475 $Y=0.84
+ $X2=0.745 $Y2=0.84
r86 15 20 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.745 $Y=0.765
+ $X2=0.745 $Y2=0.84
r87 15 17 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.745 $Y=0.765
+ $X2=0.745 $Y2=0.445
r88 13 22 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=0.475 $Y=2.885
+ $X2=0.475 $Y2=2.515
r89 10 22 48.4185 $w=3.75e-07 $l=1.87e-07 $layer=POLY_cond $X=0.587 $Y=2.328
+ $X2=0.587 $Y2=2.515
r90 9 27 3.26277 $w=3.75e-07 $l=2.2e-08 $layer=POLY_cond $X=0.587 $Y=2.032
+ $X2=0.587 $Y2=2.01
r91 9 10 43.8991 $w=3.75e-07 $l=2.96e-07 $layer=POLY_cond $X=0.587 $Y=2.032
+ $X2=0.587 $Y2=2.328
r92 7 18 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.475 $Y=0.915
+ $X2=0.475 $Y2=0.84
r93 7 41 476.872 $w=1.5e-07 $l=9.3e-07 $layer=POLY_cond $X=0.475 $Y=0.915
+ $X2=0.475 $Y2=1.845
r94 2 34 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=1.205
+ $Y=2.54 $X2=1.33 $Y2=2.685
r95 1 38 182 $w=1.7e-07 $l=3.2249e-07 $layer=licon1_NDIFF $count=1 $X=1.25
+ $Y=0.235 $X2=1.39 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__A21O_M%B1 3 7 12 14 16 17 18 23
r47 17 18 22.5128 $w=2.13e-07 $l=4.2e-07 $layer=LI1_cond $X=1.177 $Y=1.615
+ $X2=1.177 $Y2=2.035
r48 17 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.155
+ $Y=1.615 $X2=1.155 $Y2=1.615
r49 16 17 17.1526 $w=2.13e-07 $l=3.2e-07 $layer=LI1_cond $X=1.177 $Y=1.295
+ $X2=1.177 $Y2=1.615
r50 12 23 78.6876 $w=3.3e-07 $l=4.5e-07 $layer=POLY_cond $X=1.155 $Y=2.065
+ $X2=1.155 $Y2=1.615
r51 12 14 199.979 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=1.155 $Y=2.14
+ $X2=1.545 $Y2=2.14
r52 10 23 38.6168 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.155 $Y=1.45
+ $X2=1.155 $Y2=1.615
r53 5 14 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.545 $Y=2.215
+ $X2=1.545 $Y2=2.14
r54 5 7 274.33 $w=1.5e-07 $l=5.35e-07 $layer=POLY_cond $X=1.545 $Y=2.215
+ $X2=1.545 $Y2=2.75
r55 3 10 515.33 $w=1.5e-07 $l=1.005e-06 $layer=POLY_cond $X=1.175 $Y=0.445
+ $X2=1.175 $Y2=1.45
.ends

.subckt PM_SKY130_FD_SC_LP__A21O_M%A1 3 7 9 10 11 12 18
c45 18 0 1.37919e-19 $X=1.885 $Y=1.32
r46 18 21 82.0993 $w=5.2e-07 $l=5.05e-07 $layer=POLY_cond $X=1.79 $Y=1.32
+ $X2=1.79 $Y2=1.825
r47 18 20 47.1166 $w=5.2e-07 $l=1.65e-07 $layer=POLY_cond $X=1.79 $Y=1.32
+ $X2=1.79 $Y2=1.155
r48 18 19 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.885
+ $Y=1.32 $X2=1.885 $Y2=1.32
r49 11 12 9.58211 $w=4.43e-07 $l=3.7e-07 $layer=LI1_cond $X=2.022 $Y=1.665
+ $X2=2.022 $Y2=2.035
r50 11 19 8.93467 $w=4.43e-07 $l=3.45e-07 $layer=LI1_cond $X=2.022 $Y=1.665
+ $X2=2.022 $Y2=1.32
r51 10 19 0.64744 $w=4.43e-07 $l=2.5e-08 $layer=LI1_cond $X=2.022 $Y=1.295
+ $X2=2.022 $Y2=1.32
r52 9 10 9.58211 $w=4.43e-07 $l=3.7e-07 $layer=LI1_cond $X=2.022 $Y=0.925
+ $X2=2.022 $Y2=1.295
r53 7 21 474.309 $w=1.5e-07 $l=9.25e-07 $layer=POLY_cond $X=1.975 $Y=2.75
+ $X2=1.975 $Y2=1.825
r54 3 20 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=1.605 $Y=0.445
+ $X2=1.605 $Y2=1.155
.ends

.subckt PM_SKY130_FD_SC_LP__A21O_M%A2 1 3 4 5 8 12 13 14 15 16 17 24
r34 16 17 20.5182 $w=1.98e-07 $l=3.7e-07 $layer=LI1_cond $X=2.625 $Y=1.665
+ $X2=2.625 $Y2=2.035
r35 15 16 20.5182 $w=1.98e-07 $l=3.7e-07 $layer=LI1_cond $X=2.625 $Y=1.295
+ $X2=2.625 $Y2=1.665
r36 14 15 20.5182 $w=1.98e-07 $l=3.7e-07 $layer=LI1_cond $X=2.625 $Y=0.925
+ $X2=2.625 $Y2=1.295
r37 14 24 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.61
+ $Y=0.93 $X2=2.61 $Y2=0.93
r38 13 14 20.5182 $w=1.98e-07 $l=3.7e-07 $layer=LI1_cond $X=2.625 $Y=0.555
+ $X2=2.625 $Y2=0.925
r39 11 24 35.3689 $w=4.45e-07 $l=2.83e-07 $layer=POLY_cond $X=2.552 $Y=1.213
+ $X2=2.552 $Y2=0.93
r40 11 12 53.9265 $w=4.45e-07 $l=2.22e-07 $layer=POLY_cond $X=2.552 $Y=1.213
+ $X2=2.552 $Y2=1.435
r41 10 24 1.87468 $w=4.45e-07 $l=1.5e-08 $layer=POLY_cond $X=2.552 $Y=0.915
+ $X2=2.552 $Y2=0.93
r42 8 12 674.287 $w=1.5e-07 $l=1.315e-06 $layer=POLY_cond $X=2.405 $Y=2.75
+ $X2=2.405 $Y2=1.435
r43 4 10 36.6125 $w=1.5e-07 $l=2.56776e-07 $layer=POLY_cond $X=2.33 $Y=0.84
+ $X2=2.552 $Y2=0.915
r44 4 5 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=2.33 $Y=0.84 $X2=2.04
+ $Y2=0.84
r45 1 5 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.965 $Y=0.765
+ $X2=2.04 $Y2=0.84
r46 1 3 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.965 $Y=0.765
+ $X2=1.965 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__A21O_M%X 1 2 7 8 9 10 11 12 13 41
r18 39 41 9.7783 $w=3.28e-07 $l=2.8e-07 $layer=LI1_cond $X=0.25 $Y=0.51 $X2=0.53
+ $Y2=0.51
r19 21 39 3.96751 $w=1.9e-07 $l=1.65e-07 $layer=LI1_cond $X=0.25 $Y=0.675
+ $X2=0.25 $Y2=0.51
r20 12 13 21.5981 $w=1.88e-07 $l=3.7e-07 $layer=LI1_cond $X=0.25 $Y=2.405
+ $X2=0.25 $Y2=2.775
r21 11 12 21.5981 $w=1.88e-07 $l=3.7e-07 $layer=LI1_cond $X=0.25 $Y=2.035
+ $X2=0.25 $Y2=2.405
r22 10 11 21.5981 $w=1.88e-07 $l=3.7e-07 $layer=LI1_cond $X=0.25 $Y=1.665
+ $X2=0.25 $Y2=2.035
r23 9 10 21.5981 $w=1.88e-07 $l=3.7e-07 $layer=LI1_cond $X=0.25 $Y=1.295
+ $X2=0.25 $Y2=1.665
r24 8 9 21.5981 $w=1.88e-07 $l=3.7e-07 $layer=LI1_cond $X=0.25 $Y=0.925 $X2=0.25
+ $Y2=1.295
r25 8 21 14.5933 $w=1.88e-07 $l=2.5e-07 $layer=LI1_cond $X=0.25 $Y=0.925
+ $X2=0.25 $Y2=0.675
r26 7 39 0.349225 $w=3.28e-07 $l=1e-08 $layer=LI1_cond $X=0.24 $Y=0.51 $X2=0.25
+ $Y2=0.51
r27 2 13 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.675 $X2=0.26 $Y2=2.82
r28 1 41 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=0.405
+ $Y=0.235 $X2=0.53 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_LP__A21O_M%VPWR 1 2 9 13 15 17 22 29 30 33 36
r38 36 37 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r39 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r40 30 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r41 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r42 27 36 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=2.295 $Y=3.33
+ $X2=2.19 $Y2=3.33
r43 27 29 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=2.295 $Y=3.33
+ $X2=2.64 $Y2=3.33
r44 26 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r45 25 26 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r46 23 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.855 $Y=3.33
+ $X2=0.69 $Y2=3.33
r47 23 25 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.855 $Y=3.33
+ $X2=1.2 $Y2=3.33
r48 22 36 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=2.085 $Y=3.33
+ $X2=2.19 $Y2=3.33
r49 22 25 57.738 $w=1.68e-07 $l=8.85e-07 $layer=LI1_cond $X=2.085 $Y=3.33
+ $X2=1.2 $Y2=3.33
r50 20 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r51 19 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r52 17 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.525 $Y=3.33
+ $X2=0.69 $Y2=3.33
r53 17 19 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.525 $Y=3.33
+ $X2=0.24 $Y2=3.33
r54 15 37 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=2.16 $Y2=3.33
r55 15 26 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=1.2 $Y2=3.33
r56 11 36 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=2.19 $Y=3.245
+ $X2=2.19 $Y2=3.33
r57 11 13 22.71 $w=2.08e-07 $l=4.3e-07 $layer=LI1_cond $X=2.19 $Y=3.245 $X2=2.19
+ $Y2=2.815
r58 7 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=3.245 $X2=0.69
+ $Y2=3.33
r59 7 9 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.69 $Y=3.245
+ $X2=0.69 $Y2=2.95
r60 2 13 600 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=1 $X=2.05
+ $Y=2.54 $X2=2.19 $Y2=2.815
r61 1 9 600 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=2.675 $X2=0.69 $Y2=2.95
.ends

.subckt PM_SKY130_FD_SC_LP__A21O_M%A_324_508# 1 2 9 11 12 15
c23 11 0 1.26348e-19 $X=2.515 $Y=2.385
r24 13 15 11.355 $w=2.08e-07 $l=2.15e-07 $layer=LI1_cond $X=2.62 $Y=2.47
+ $X2=2.62 $Y2=2.685
r25 11 13 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=2.515 $Y=2.385
+ $X2=2.62 $Y2=2.47
r26 11 12 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=2.515 $Y=2.385
+ $X2=1.865 $Y2=2.385
r27 7 12 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=1.76 $Y=2.47
+ $X2=1.865 $Y2=2.385
r28 7 9 11.355 $w=2.08e-07 $l=2.15e-07 $layer=LI1_cond $X=1.76 $Y=2.47 $X2=1.76
+ $Y2=2.685
r29 2 15 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.48
+ $Y=2.54 $X2=2.62 $Y2=2.685
r30 1 9 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.62
+ $Y=2.54 $X2=1.76 $Y2=2.685
.ends

.subckt PM_SKY130_FD_SC_LP__A21O_M%VGND 1 2 9 13 16 17 18 24 30 31 34
c40 13 0 1.15713e-20 $X=2.18 $Y=0.38
r41 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r42 31 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=2.16
+ $Y2=0
r43 30 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r44 28 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.345 $Y=0 $X2=2.18
+ $Y2=0
r45 28 30 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=2.345 $Y=0 $X2=2.64
+ $Y2=0
r46 27 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r47 26 27 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r48 24 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.015 $Y=0 $X2=2.18
+ $Y2=0
r49 24 26 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=2.015 $Y=0 $X2=1.68
+ $Y2=0
r50 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r51 18 27 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=1.68
+ $Y2=0
r52 18 22 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=0.72
+ $Y2=0
r53 16 21 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=0.855 $Y=0 $X2=0.72
+ $Y2=0
r54 16 17 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=0.855 $Y=0 $X2=0.96
+ $Y2=0
r55 15 26 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=1.065 $Y=0 $X2=1.68
+ $Y2=0
r56 15 17 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.065 $Y=0 $X2=0.96
+ $Y2=0
r57 11 34 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.18 $Y=0.085
+ $X2=2.18 $Y2=0
r58 11 13 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.18 $Y=0.085
+ $X2=2.18 $Y2=0.38
r59 7 17 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=0.96 $Y=0.085
+ $X2=0.96 $Y2=0
r60 7 9 15.5801 $w=2.08e-07 $l=2.95e-07 $layer=LI1_cond $X=0.96 $Y=0.085
+ $X2=0.96 $Y2=0.38
r61 2 13 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=2.04
+ $Y=0.235 $X2=2.18 $Y2=0.38
r62 1 9 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=0.82
+ $Y=0.235 $X2=0.96 $Y2=0.38
.ends

