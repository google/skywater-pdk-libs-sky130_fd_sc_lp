* File: sky130_fd_sc_lp__o311ai_0.pxi.spice
* Created: Fri Aug 28 11:14:19 2020
* 
x_PM_SKY130_FD_SC_LP__O311AI_0%A1 N_A1_c_78_n N_A1_c_79_n N_A1_M1005_g
+ N_A1_c_85_n N_A1_M1001_g N_A1_c_80_n N_A1_c_81_n N_A1_c_86_n A1 A1 A1
+ N_A1_c_83_n PM_SKY130_FD_SC_LP__O311AI_0%A1
x_PM_SKY130_FD_SC_LP__O311AI_0%A2 N_A2_M1002_g N_A2_M1000_g N_A2_c_118_n
+ N_A2_c_119_n N_A2_c_126_n N_A2_c_120_n N_A2_c_121_n A2 A2 N_A2_c_123_n
+ PM_SKY130_FD_SC_LP__O311AI_0%A2
x_PM_SKY130_FD_SC_LP__O311AI_0%A3 N_A3_c_165_n N_A3_M1004_g N_A3_M1006_g
+ N_A3_c_167_n A3 A3 N_A3_c_169_n PM_SKY130_FD_SC_LP__O311AI_0%A3
x_PM_SKY130_FD_SC_LP__O311AI_0%B1 N_B1_c_208_n N_B1_M1007_g N_B1_M1009_g
+ N_B1_c_209_n N_B1_c_210_n N_B1_c_205_n N_B1_c_212_n B1 B1 N_B1_c_207_n
+ PM_SKY130_FD_SC_LP__O311AI_0%B1
x_PM_SKY130_FD_SC_LP__O311AI_0%C1 N_C1_c_253_n N_C1_M1008_g N_C1_c_260_n
+ N_C1_M1003_g N_C1_c_254_n N_C1_c_255_n N_C1_c_261_n N_C1_c_262_n N_C1_c_256_n
+ N_C1_c_257_n C1 C1 C1 N_C1_c_259_n PM_SKY130_FD_SC_LP__O311AI_0%C1
x_PM_SKY130_FD_SC_LP__O311AI_0%VPWR N_VPWR_M1001_s N_VPWR_M1007_d N_VPWR_c_299_n
+ N_VPWR_c_300_n N_VPWR_c_301_n N_VPWR_c_302_n VPWR N_VPWR_c_303_n
+ N_VPWR_c_304_n N_VPWR_c_298_n N_VPWR_c_306_n PM_SKY130_FD_SC_LP__O311AI_0%VPWR
x_PM_SKY130_FD_SC_LP__O311AI_0%Y N_Y_M1008_d N_Y_M1004_d N_Y_M1003_d N_Y_c_333_n
+ N_Y_c_334_n N_Y_c_331_n Y Y Y Y N_Y_c_337_n Y PM_SKY130_FD_SC_LP__O311AI_0%Y
x_PM_SKY130_FD_SC_LP__O311AI_0%VGND N_VGND_M1005_s N_VGND_M1000_d N_VGND_c_383_n
+ N_VGND_c_384_n VGND N_VGND_c_385_n N_VGND_c_386_n N_VGND_c_387_n
+ N_VGND_c_388_n N_VGND_c_389_n N_VGND_c_390_n PM_SKY130_FD_SC_LP__O311AI_0%VGND
x_PM_SKY130_FD_SC_LP__O311AI_0%A_193_48# N_A_193_48#_M1005_d N_A_193_48#_M1006_d
+ N_A_193_48#_c_425_n N_A_193_48#_c_426_n N_A_193_48#_c_427_n
+ N_A_193_48#_c_428_n PM_SKY130_FD_SC_LP__O311AI_0%A_193_48#
cc_1 VNB N_A1_c_78_n 0.0117181f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=2.07
cc_2 VNB N_A1_c_79_n 0.0214152f $X=-0.19 $Y=-0.245 $X2=0.89 $Y2=0.77
cc_3 VNB N_A1_c_80_n 0.0377902f $X=-0.19 $Y=-0.245 $X2=0.89 $Y2=0.845
cc_4 VNB N_A1_c_81_n 0.0231487f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=1.44
cc_5 VNB A1 0.0158413f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.84
cc_6 VNB N_A1_c_83_n 0.0356623f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=0.935
cc_7 VNB N_A2_c_118_n 0.0140912f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A2_c_119_n 0.0203209f $X=-0.19 $Y=-0.245 $X2=0.89 $Y2=0.845
cc_9 VNB N_A2_c_120_n 0.0165601f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=1.275
cc_10 VNB N_A2_c_121_n 0.0114326f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=1.44
cc_11 VNB A2 0.00479768f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=2.145
cc_12 VNB N_A2_c_123_n 0.0157504f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_13 VNB N_A3_c_165_n 0.0210981f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=2.07
cc_14 VNB N_A3_M1006_g 0.0373446f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=0.845
cc_15 VNB N_A3_c_167_n 0.00151785f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB A3 0.00186576f $X=-0.19 $Y=-0.245 $X2=0.89 $Y2=0.845
cc_17 VNB N_A3_c_169_n 0.0215171f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_B1_M1009_g 0.0372183f $X=-0.19 $Y=-0.245 $X2=0.89 $Y2=2.22
cc_19 VNB N_B1_c_205_n 0.0233329f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=2.145
cc_20 VNB B1 0.0113711f $X=-0.19 $Y=-0.245 $X2=0.89 $Y2=2.145
cc_21 VNB N_B1_c_207_n 0.0168112f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_C1_c_253_n 0.0198811f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=1.44
cc_23 VNB N_C1_c_254_n 0.0397654f $X=-0.19 $Y=-0.245 $X2=0.89 $Y2=2.65
cc_24 VNB N_C1_c_255_n 0.0123824f $X=-0.19 $Y=-0.245 $X2=0.89 $Y2=2.65
cc_25 VNB N_C1_c_256_n 0.00981538f $X=-0.19 $Y=-0.245 $X2=0.89 $Y2=0.845
cc_26 VNB N_C1_c_257_n 0.0196204f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=1.44
cc_27 VNB C1 0.0300239f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=2.145
cc_28 VNB N_C1_c_259_n 0.0356283f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VPWR_c_298_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_Y_c_331_n 0.0134652f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB Y 0.0170327f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_32 VNB N_VGND_c_383_n 0.0170667f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=0.845
cc_33 VNB N_VGND_c_384_n 0.00486412f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_385_n 0.0183725f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_386_n 0.0154972f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_36 VNB N_VGND_c_387_n 0.0487307f $X=-0.19 $Y=-0.245 $X2=0.687 $Y2=0.925
cc_37 VNB N_VGND_c_388_n 0.207238f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_389_n 0.00514657f $X=-0.19 $Y=-0.245 $X2=0.687 $Y2=1.295
cc_39 VNB N_VGND_c_390_n 0.00545686f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_193_48#_c_425_n 0.00111702f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=0.845
cc_41 VNB N_A_193_48#_c_426_n 0.0174597f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_193_48#_c_427_n 0.00224477f $X=-0.19 $Y=-0.245 $X2=0.89 $Y2=0.845
cc_43 VNB N_A_193_48#_c_428_n 0.00101617f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=1.44
cc_44 VPB N_A1_c_78_n 0.030038f $X=-0.19 $Y=1.655 $X2=0.71 $Y2=2.07
cc_45 VPB N_A1_c_85_n 0.0211787f $X=-0.19 $Y=1.655 $X2=0.89 $Y2=2.22
cc_46 VPB N_A1_c_86_n 0.0281753f $X=-0.19 $Y=1.655 $X2=0.89 $Y2=2.145
cc_47 VPB A1 0.00971323f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=0.84
cc_48 VPB N_A2_M1002_g 0.0370252f $X=-0.19 $Y=1.655 $X2=0.89 $Y2=0.45
cc_49 VPB N_A2_c_119_n 5.55892e-19 $X=-0.19 $Y=1.655 $X2=0.89 $Y2=0.845
cc_50 VPB N_A2_c_126_n 0.0157504f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_51 VPB A2 0.00915027f $X=-0.19 $Y=1.655 $X2=0.71 $Y2=2.145
cc_52 VPB N_A3_M1004_g 0.0394374f $X=-0.19 $Y=1.655 $X2=0.89 $Y2=0.45
cc_53 VPB N_A3_c_167_n 0.0199887f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_54 VPB N_B1_c_208_n 0.0184915f $X=-0.19 $Y=1.655 $X2=0.71 $Y2=1.44
cc_55 VPB N_B1_c_209_n 0.0158403f $X=-0.19 $Y=1.655 $X2=0.62 $Y2=0.845
cc_56 VPB N_B1_c_210_n 0.0177367f $X=-0.19 $Y=1.655 $X2=0.89 $Y2=0.845
cc_57 VPB N_B1_c_205_n 6.38287e-19 $X=-0.19 $Y=1.655 $X2=0.71 $Y2=2.145
cc_58 VPB N_B1_c_212_n 0.0165812f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_59 VPB B1 0.00158781f $X=-0.19 $Y=1.655 $X2=0.89 $Y2=2.145
cc_60 VPB N_C1_c_260_n 0.021842f $X=-0.19 $Y=1.655 $X2=0.89 $Y2=0.45
cc_61 VPB N_C1_c_261_n 0.0268813f $X=-0.19 $Y=1.655 $X2=0.62 $Y2=0.845
cc_62 VPB N_C1_c_262_n 0.00902828f $X=-0.19 $Y=1.655 $X2=0.62 $Y2=0.92
cc_63 VPB N_C1_c_256_n 0.0297168f $X=-0.19 $Y=1.655 $X2=0.89 $Y2=0.845
cc_64 VPB C1 0.00647366f $X=-0.19 $Y=1.655 $X2=0.71 $Y2=2.145
cc_65 VPB N_VPWR_c_299_n 0.0386796f $X=-0.19 $Y=1.655 $X2=0.62 $Y2=0.845
cc_66 VPB N_VPWR_c_300_n 0.0121481f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_67 VPB N_VPWR_c_301_n 0.0405616f $X=-0.19 $Y=1.655 $X2=0.71 $Y2=2.145
cc_68 VPB N_VPWR_c_302_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_69 VPB N_VPWR_c_303_n 0.0183725f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=0.84
cc_70 VPB N_VPWR_c_304_n 0.0238586f $X=-0.19 $Y=1.655 $X2=0.687 $Y2=1.295
cc_71 VPB N_VPWR_c_298_n 0.0872647f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_72 VPB N_VPWR_c_306_n 0.0060562f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_73 VPB N_Y_c_333_n 0.00598453f $X=-0.19 $Y=1.655 $X2=0.89 $Y2=0.845
cc_74 VPB N_Y_c_334_n 0.00875598f $X=-0.19 $Y=1.655 $X2=0.62 $Y2=1.275
cc_75 VPB Y 0.0179719f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_76 VPB Y 0.0474588f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_77 VPB N_Y_c_337_n 0.0108869f $X=-0.19 $Y=1.655 $X2=0.687 $Y2=1.665
cc_78 N_A1_c_78_n N_A2_M1002_g 0.008947f $X=0.71 $Y=2.07 $X2=0 $Y2=0
cc_79 N_A1_c_86_n N_A2_M1002_g 0.065003f $X=0.89 $Y=2.145 $X2=0 $Y2=0
cc_80 A1 N_A2_c_118_n 0.00356342f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_81 N_A1_c_83_n N_A2_c_118_n 0.00652152f $X=0.62 $Y=0.935 $X2=0 $Y2=0
cc_82 N_A1_c_81_n N_A2_c_119_n 0.0138553f $X=0.62 $Y=1.44 $X2=0 $Y2=0
cc_83 N_A1_c_78_n N_A2_c_126_n 0.0138553f $X=0.71 $Y=2.07 $X2=0 $Y2=0
cc_84 N_A1_c_79_n N_A2_c_120_n 0.0121583f $X=0.89 $Y=0.77 $X2=0 $Y2=0
cc_85 N_A1_c_80_n N_A2_c_121_n 0.00953079f $X=0.89 $Y=0.845 $X2=0 $Y2=0
cc_86 A1 A2 0.052788f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_87 N_A1_c_83_n A2 7.3276e-19 $X=0.62 $Y=0.935 $X2=0 $Y2=0
cc_88 A1 N_A2_c_123_n 0.00385203f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_89 N_A1_c_83_n N_A2_c_123_n 0.0138553f $X=0.62 $Y=0.935 $X2=0 $Y2=0
cc_90 N_A1_c_85_n N_VPWR_c_299_n 0.0172898f $X=0.89 $Y=2.22 $X2=0 $Y2=0
cc_91 N_A1_c_86_n N_VPWR_c_299_n 0.00604348f $X=0.89 $Y=2.145 $X2=0 $Y2=0
cc_92 A1 N_VPWR_c_299_n 0.012827f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_93 N_A1_c_85_n N_VPWR_c_301_n 0.00389963f $X=0.89 $Y=2.22 $X2=0 $Y2=0
cc_94 N_A1_c_85_n N_VPWR_c_298_n 0.00762892f $X=0.89 $Y=2.22 $X2=0 $Y2=0
cc_95 N_A1_c_79_n N_VGND_c_383_n 0.00918295f $X=0.89 $Y=0.77 $X2=0 $Y2=0
cc_96 N_A1_c_80_n N_VGND_c_383_n 0.00320107f $X=0.89 $Y=0.845 $X2=0 $Y2=0
cc_97 A1 N_VGND_c_383_n 0.0230368f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_98 N_A1_c_80_n N_VGND_c_385_n 0.00106709f $X=0.89 $Y=0.845 $X2=0 $Y2=0
cc_99 N_A1_c_79_n N_VGND_c_386_n 0.0048178f $X=0.89 $Y=0.77 $X2=0 $Y2=0
cc_100 N_A1_c_79_n N_VGND_c_388_n 0.00835603f $X=0.89 $Y=0.77 $X2=0 $Y2=0
cc_101 N_A1_c_80_n N_VGND_c_388_n 0.00147479f $X=0.89 $Y=0.845 $X2=0 $Y2=0
cc_102 A1 N_VGND_c_388_n 0.00111334f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_103 N_A1_c_79_n N_A_193_48#_c_425_n 0.0030097f $X=0.89 $Y=0.77 $X2=0 $Y2=0
cc_104 A1 N_A_193_48#_c_425_n 0.00111458f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_105 N_A1_c_80_n N_A_193_48#_c_427_n 0.00112636f $X=0.89 $Y=0.845 $X2=0 $Y2=0
cc_106 A1 N_A_193_48#_c_427_n 0.0174786f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_107 N_A1_c_83_n N_A_193_48#_c_427_n 2.63243e-19 $X=0.62 $Y=0.935 $X2=0 $Y2=0
cc_108 N_A2_c_119_n N_A3_c_165_n 0.0300975f $X=1.16 $Y=1.665 $X2=0 $Y2=0
cc_109 N_A2_M1002_g N_A3_M1004_g 0.0300975f $X=1.25 $Y=2.65 $X2=0 $Y2=0
cc_110 N_A2_c_118_n N_A3_M1006_g 0.0079383f $X=1.16 $Y=1.16 $X2=0 $Y2=0
cc_111 N_A2_c_120_n N_A3_M1006_g 0.0150019f $X=1.285 $Y=0.77 $X2=0 $Y2=0
cc_112 N_A2_c_126_n N_A3_c_167_n 0.0300975f $X=1.16 $Y=1.83 $X2=0 $Y2=0
cc_113 A2 A3 0.0471f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_114 N_A2_c_123_n A3 7.30456e-19 $X=1.16 $Y=1.325 $X2=0 $Y2=0
cc_115 A2 N_A3_c_169_n 0.0047586f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_116 N_A2_c_123_n N_A3_c_169_n 0.0300975f $X=1.16 $Y=1.325 $X2=0 $Y2=0
cc_117 N_A2_M1002_g N_VPWR_c_299_n 0.00396356f $X=1.25 $Y=2.65 $X2=0 $Y2=0
cc_118 N_A2_M1002_g N_VPWR_c_301_n 0.00469667f $X=1.25 $Y=2.65 $X2=0 $Y2=0
cc_119 N_A2_M1002_g N_VPWR_c_298_n 0.00923821f $X=1.25 $Y=2.65 $X2=0 $Y2=0
cc_120 N_A2_c_120_n N_VGND_c_383_n 5.18826e-19 $X=1.285 $Y=0.77 $X2=0 $Y2=0
cc_121 N_A2_c_120_n N_VGND_c_384_n 0.00167407f $X=1.285 $Y=0.77 $X2=0 $Y2=0
cc_122 N_A2_c_120_n N_VGND_c_386_n 0.00559736f $X=1.285 $Y=0.77 $X2=0 $Y2=0
cc_123 N_A2_c_120_n N_VGND_c_388_n 0.00625648f $X=1.285 $Y=0.77 $X2=0 $Y2=0
cc_124 N_A2_c_120_n N_A_193_48#_c_425_n 0.00728821f $X=1.285 $Y=0.77 $X2=0 $Y2=0
cc_125 N_A2_c_121_n N_A_193_48#_c_425_n 0.00200465f $X=1.285 $Y=0.92 $X2=0 $Y2=0
cc_126 N_A2_c_118_n N_A_193_48#_c_426_n 0.00234813f $X=1.16 $Y=1.16 $X2=0 $Y2=0
cc_127 N_A2_c_121_n N_A_193_48#_c_426_n 0.00765737f $X=1.285 $Y=0.92 $X2=0 $Y2=0
cc_128 A2 N_A_193_48#_c_426_n 0.00745249f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_129 N_A2_c_118_n N_A_193_48#_c_427_n 0.00246371f $X=1.16 $Y=1.16 $X2=0 $Y2=0
cc_130 N_A2_c_121_n N_A_193_48#_c_427_n 0.00189237f $X=1.285 $Y=0.92 $X2=0 $Y2=0
cc_131 A2 N_A_193_48#_c_427_n 0.0218543f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_132 N_A2_c_123_n N_A_193_48#_c_427_n 0.00128156f $X=1.16 $Y=1.325 $X2=0 $Y2=0
cc_133 N_A3_M1006_g N_B1_M1009_g 0.0306579f $X=1.81 $Y=0.45 $X2=0 $Y2=0
cc_134 N_A3_M1004_g N_B1_c_209_n 0.00585083f $X=1.61 $Y=2.65 $X2=0 $Y2=0
cc_135 N_A3_M1004_g N_B1_c_210_n 0.012834f $X=1.61 $Y=2.65 $X2=0 $Y2=0
cc_136 N_A3_c_165_n N_B1_c_205_n 0.0119992f $X=1.73 $Y=1.635 $X2=0 $Y2=0
cc_137 N_A3_c_167_n N_B1_c_212_n 0.0119992f $X=1.73 $Y=1.83 $X2=0 $Y2=0
cc_138 A3 B1 0.0503154f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_139 N_A3_c_169_n B1 0.00444885f $X=1.7 $Y=1.325 $X2=0 $Y2=0
cc_140 A3 N_B1_c_207_n 5.60537e-19 $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_141 N_A3_c_169_n N_B1_c_207_n 0.0119992f $X=1.7 $Y=1.325 $X2=0 $Y2=0
cc_142 N_A3_M1004_g N_VPWR_c_301_n 0.00469667f $X=1.61 $Y=2.65 $X2=0 $Y2=0
cc_143 N_A3_M1004_g N_VPWR_c_298_n 0.00927506f $X=1.61 $Y=2.65 $X2=0 $Y2=0
cc_144 N_A3_M1004_g N_Y_c_333_n 0.00634268f $X=1.61 $Y=2.65 $X2=0 $Y2=0
cc_145 N_A3_M1004_g N_Y_c_334_n 0.00597017f $X=1.61 $Y=2.65 $X2=0 $Y2=0
cc_146 N_A3_c_167_n N_Y_c_334_n 0.00768116f $X=1.73 $Y=1.83 $X2=0 $Y2=0
cc_147 A3 N_Y_c_334_n 0.0140807f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_148 N_A3_M1006_g N_VGND_c_384_n 0.00319125f $X=1.81 $Y=0.45 $X2=0 $Y2=0
cc_149 N_A3_M1006_g N_VGND_c_387_n 0.0058025f $X=1.81 $Y=0.45 $X2=0 $Y2=0
cc_150 N_A3_M1006_g N_VGND_c_388_n 0.00632127f $X=1.81 $Y=0.45 $X2=0 $Y2=0
cc_151 N_A3_M1006_g N_A_193_48#_c_425_n 5.25359e-19 $X=1.81 $Y=0.45 $X2=0 $Y2=0
cc_152 N_A3_M1006_g N_A_193_48#_c_426_n 0.0142033f $X=1.81 $Y=0.45 $X2=0 $Y2=0
cc_153 A3 N_A_193_48#_c_426_n 0.0258824f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_154 N_A3_c_169_n N_A_193_48#_c_426_n 0.00331883f $X=1.7 $Y=1.325 $X2=0 $Y2=0
cc_155 N_A3_M1006_g N_A_193_48#_c_428_n 0.00197359f $X=1.81 $Y=0.45 $X2=0 $Y2=0
cc_156 N_B1_M1009_g N_C1_c_253_n 0.0419948f $X=2.24 $Y=0.45 $X2=-0.19 $Y2=-0.245
cc_157 N_B1_c_208_n N_C1_c_260_n 0.006119f $X=2.1 $Y=2.22 $X2=0 $Y2=0
cc_158 N_B1_c_210_n N_C1_c_262_n 0.00857218f $X=2.24 $Y=2.145 $X2=0 $Y2=0
cc_159 N_B1_c_209_n N_C1_c_256_n 0.00175337f $X=2.24 $Y=2.07 $X2=0 $Y2=0
cc_160 N_B1_c_212_n N_C1_c_256_n 0.00458825f $X=2.33 $Y=1.83 $X2=0 $Y2=0
cc_161 N_B1_c_205_n N_C1_c_257_n 0.00458825f $X=2.33 $Y=1.665 $X2=0 $Y2=0
cc_162 N_B1_M1009_g N_C1_c_259_n 0.00179346f $X=2.24 $Y=0.45 $X2=0 $Y2=0
cc_163 N_B1_c_207_n N_C1_c_259_n 0.00458825f $X=2.33 $Y=1.325 $X2=0 $Y2=0
cc_164 N_B1_c_208_n N_VPWR_c_300_n 0.0036132f $X=2.1 $Y=2.22 $X2=0 $Y2=0
cc_165 N_B1_c_210_n N_VPWR_c_300_n 0.00329f $X=2.24 $Y=2.145 $X2=0 $Y2=0
cc_166 N_B1_c_208_n N_VPWR_c_301_n 0.00459311f $X=2.1 $Y=2.22 $X2=0 $Y2=0
cc_167 N_B1_c_208_n N_VPWR_c_298_n 0.00894505f $X=2.1 $Y=2.22 $X2=0 $Y2=0
cc_168 N_B1_c_208_n N_Y_c_333_n 0.00949421f $X=2.1 $Y=2.22 $X2=0 $Y2=0
cc_169 N_B1_c_210_n N_Y_c_333_n 0.00333139f $X=2.24 $Y=2.145 $X2=0 $Y2=0
cc_170 N_B1_c_210_n N_Y_c_334_n 8.16348e-19 $X=2.24 $Y=2.145 $X2=0 $Y2=0
cc_171 N_B1_M1009_g N_Y_c_331_n 9.51964e-19 $X=2.24 $Y=0.45 $X2=0 $Y2=0
cc_172 N_B1_M1009_g Y 0.00554701f $X=2.24 $Y=0.45 $X2=0 $Y2=0
cc_173 N_B1_c_209_n Y 0.00226014f $X=2.24 $Y=2.07 $X2=0 $Y2=0
cc_174 B1 Y 0.0477306f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_175 N_B1_c_207_n Y 0.0061041f $X=2.33 $Y=1.325 $X2=0 $Y2=0
cc_176 N_B1_c_210_n Y 3.20171e-19 $X=2.24 $Y=2.145 $X2=0 $Y2=0
cc_177 N_B1_c_209_n N_Y_c_337_n 0.00834538f $X=2.24 $Y=2.07 $X2=0 $Y2=0
cc_178 N_B1_c_210_n N_Y_c_337_n 0.0121977f $X=2.24 $Y=2.145 $X2=0 $Y2=0
cc_179 N_B1_c_212_n N_Y_c_337_n 0.00496807f $X=2.33 $Y=1.83 $X2=0 $Y2=0
cc_180 B1 N_Y_c_337_n 0.0363483f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_181 N_B1_M1009_g N_VGND_c_387_n 0.00545083f $X=2.24 $Y=0.45 $X2=0 $Y2=0
cc_182 N_B1_M1009_g N_VGND_c_388_n 0.00998575f $X=2.24 $Y=0.45 $X2=0 $Y2=0
cc_183 N_B1_M1009_g N_A_193_48#_c_426_n 0.0062501f $X=2.24 $Y=0.45 $X2=0 $Y2=0
cc_184 B1 N_A_193_48#_c_426_n 0.0141436f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_185 N_B1_M1009_g N_A_193_48#_c_428_n 0.00974667f $X=2.24 $Y=0.45 $X2=0 $Y2=0
cc_186 N_C1_c_260_n N_VPWR_c_300_n 0.00346101f $X=2.63 $Y=2.22 $X2=0 $Y2=0
cc_187 N_C1_c_260_n N_VPWR_c_304_n 0.00469667f $X=2.63 $Y=2.22 $X2=0 $Y2=0
cc_188 N_C1_c_260_n N_VPWR_c_298_n 0.00937668f $X=2.63 $Y=2.22 $X2=0 $Y2=0
cc_189 N_C1_c_262_n N_Y_c_333_n 7.16877e-19 $X=2.705 $Y=2.145 $X2=0 $Y2=0
cc_190 N_C1_c_253_n N_Y_c_331_n 0.00620624f $X=2.63 $Y=0.77 $X2=0 $Y2=0
cc_191 N_C1_c_254_n N_Y_c_331_n 0.00791789f $X=2.925 $Y=0.845 $X2=0 $Y2=0
cc_192 N_C1_c_253_n Y 0.00501086f $X=2.63 $Y=0.77 $X2=0 $Y2=0
cc_193 N_C1_c_254_n Y 0.0111024f $X=2.925 $Y=0.845 $X2=0 $Y2=0
cc_194 N_C1_c_255_n Y 0.00359231f $X=2.705 $Y=0.845 $X2=0 $Y2=0
cc_195 N_C1_c_261_n Y 0.00724596f $X=2.925 $Y=2.145 $X2=0 $Y2=0
cc_196 N_C1_c_262_n Y 0.00327044f $X=2.705 $Y=2.145 $X2=0 $Y2=0
cc_197 N_C1_c_256_n Y 0.00965477f $X=3 $Y=2.07 $X2=0 $Y2=0
cc_198 N_C1_c_257_n Y 7.78193e-19 $X=3.09 $Y=1.51 $X2=0 $Y2=0
cc_199 C1 Y 0.0936527f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_200 N_C1_c_259_n Y 0.0115959f $X=3.09 $Y=1.005 $X2=0 $Y2=0
cc_201 N_C1_c_260_n Y 0.00399546f $X=2.63 $Y=2.22 $X2=0 $Y2=0
cc_202 N_C1_c_261_n Y 0.0160298f $X=2.925 $Y=2.145 $X2=0 $Y2=0
cc_203 N_C1_c_262_n N_Y_c_337_n 0.00765066f $X=2.705 $Y=2.145 $X2=0 $Y2=0
cc_204 N_C1_c_253_n N_VGND_c_387_n 0.00521691f $X=2.63 $Y=0.77 $X2=0 $Y2=0
cc_205 N_C1_c_254_n N_VGND_c_387_n 0.0049319f $X=2.925 $Y=0.845 $X2=0 $Y2=0
cc_206 N_C1_c_253_n N_VGND_c_388_n 0.0105015f $X=2.63 $Y=0.77 $X2=0 $Y2=0
cc_207 N_C1_c_254_n N_VGND_c_388_n 0.00652821f $X=2.925 $Y=0.845 $X2=0 $Y2=0
cc_208 C1 N_VGND_c_388_n 0.00951602f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_209 N_C1_c_255_n N_A_193_48#_c_426_n 4.92446e-19 $X=2.705 $Y=0.845 $X2=0
+ $Y2=0
cc_210 N_C1_c_253_n N_A_193_48#_c_428_n 0.00141921f $X=2.63 $Y=0.77 $X2=0 $Y2=0
cc_211 N_VPWR_c_300_n N_Y_c_333_n 0.0255136f $X=2.37 $Y=2.485 $X2=0 $Y2=0
cc_212 N_VPWR_c_301_n N_Y_c_333_n 0.0146088f $X=2.205 $Y=3.33 $X2=0 $Y2=0
cc_213 N_VPWR_c_298_n N_Y_c_333_n 0.0120707f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_214 N_VPWR_c_300_n Y 0.0313483f $X=2.37 $Y=2.485 $X2=0 $Y2=0
cc_215 N_VPWR_c_304_n Y 0.0264029f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_216 N_VPWR_c_298_n Y 0.0211034f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_217 N_VPWR_c_300_n N_Y_c_337_n 0.0242776f $X=2.37 $Y=2.485 $X2=0 $Y2=0
cc_218 N_Y_c_331_n N_VGND_c_387_n 0.0176903f $X=2.845 $Y=0.45 $X2=0 $Y2=0
cc_219 N_Y_M1008_d N_VGND_c_388_n 0.00215838f $X=2.705 $Y=0.24 $X2=0 $Y2=0
cc_220 N_Y_c_331_n N_VGND_c_388_n 0.0127506f $X=2.845 $Y=0.45 $X2=0 $Y2=0
cc_221 Y N_A_193_48#_c_426_n 0.00701666f $X=2.555 $Y=1.95 $X2=0 $Y2=0
cc_222 N_Y_c_331_n N_A_193_48#_c_428_n 0.010672f $X=2.845 $Y=0.45 $X2=0 $Y2=0
cc_223 Y N_A_193_48#_c_428_n 0.00520122f $X=2.555 $Y=1.95 $X2=0 $Y2=0
cc_224 N_VGND_c_388_n N_A_193_48#_M1005_d 0.00386283f $X=3.12 $Y=0 $X2=-0.19
+ $Y2=-0.245
cc_225 N_VGND_c_388_n N_A_193_48#_M1006_d 0.00225666f $X=3.12 $Y=0 $X2=0 $Y2=0
cc_226 N_VGND_c_386_n N_A_193_48#_c_425_n 0.0126287f $X=1.43 $Y=0 $X2=0 $Y2=0
cc_227 N_VGND_c_388_n N_A_193_48#_c_425_n 0.00943397f $X=3.12 $Y=0 $X2=0 $Y2=0
cc_228 N_VGND_c_384_n N_A_193_48#_c_426_n 0.0205333f $X=1.57 $Y=0.45 $X2=0 $Y2=0
cc_229 N_VGND_c_388_n N_A_193_48#_c_426_n 0.0114202f $X=3.12 $Y=0 $X2=0 $Y2=0
cc_230 N_VGND_c_387_n N_A_193_48#_c_428_n 0.0145575f $X=3.12 $Y=0 $X2=0 $Y2=0
cc_231 N_VGND_c_388_n N_A_193_48#_c_428_n 0.0114964f $X=3.12 $Y=0 $X2=0 $Y2=0
cc_232 N_VGND_c_388_n A_463_48# 0.010279f $X=3.12 $Y=0 $X2=-0.19 $Y2=-0.245
