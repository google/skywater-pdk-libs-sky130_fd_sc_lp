* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__or4b_1 A B C D_N VGND VNB VPB VPWR X
X0 a_483_367# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X1 a_220_367# a_64_131# a_303_367# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X2 VGND a_64_131# a_220_367# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 a_220_367# C VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 VGND B a_220_367# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 a_303_367# C a_397_367# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X6 VPWR a_220_367# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X7 VGND a_220_367# X VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X8 a_220_367# A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 a_64_131# D_N VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 a_64_131# D_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X11 a_397_367# B a_483_367# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
.ends
