* File: sky130_fd_sc_lp__sdfrtp_2.pex.spice
* Created: Fri Aug 28 11:28:28 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__SDFRTP_2%A_35_74# 1 2 7 9 12 16 22 27 28 30 31 32 38
r69 31 34 6.16778 $w=8.98e-07 $l=4.55e-07 $layer=LI1_cond $X=0.585 $Y=2.03
+ $X2=0.585 $Y2=2.485
r70 31 32 7.94142 $w=8.98e-07 $l=1e-07 $layer=LI1_cond $X=0.585 $Y=2.03
+ $X2=0.585 $Y2=1.93
r71 28 42 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.395 $Y=2.015
+ $X2=2.395 $Y2=2.18
r72 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.395
+ $Y=2.015 $X2=2.395 $Y2=2.015
r73 25 31 9.90988 $w=2e-07 $l=4.5e-07 $layer=LI1_cond $X=1.035 $Y=2.03 $X2=0.585
+ $Y2=2.03
r74 25 27 75.4182 $w=1.98e-07 $l=1.36e-06 $layer=LI1_cond $X=1.035 $Y=2.03
+ $X2=2.395 $Y2=2.03
r75 23 38 20.9834 $w=3.3e-07 $l=1.2e-07 $layer=POLY_cond $X=1.345 $Y=0.945
+ $X2=1.465 $Y2=0.945
r76 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.345
+ $Y=0.945 $X2=1.345 $Y2=0.945
r77 20 30 2.98021 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=0.405 $Y=0.945
+ $X2=0.27 $Y2=0.945
r78 20 22 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=0.405 $Y=0.945
+ $X2=1.345 $Y2=0.945
r79 18 30 3.52026 $w=2.65e-07 $l=8.5e-08 $layer=LI1_cond $X=0.27 $Y=1.03
+ $X2=0.27 $Y2=0.945
r80 18 32 38.4148 $w=2.68e-07 $l=9e-07 $layer=LI1_cond $X=0.27 $Y=1.03 $X2=0.27
+ $Y2=1.93
r81 14 30 3.52026 $w=2.65e-07 $l=8.74643e-08 $layer=LI1_cond $X=0.265 $Y=0.86
+ $X2=0.27 $Y2=0.945
r82 14 16 12.4109 $w=2.58e-07 $l=2.8e-07 $layer=LI1_cond $X=0.265 $Y=0.86
+ $X2=0.265 $Y2=0.58
r83 12 42 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.375 $Y=2.66
+ $X2=2.375 $Y2=2.18
r84 7 38 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.465 $Y=0.78
+ $X2=1.465 $Y2=0.945
r85 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.465 $Y=0.78
+ $X2=1.465 $Y2=0.46
r86 2 34 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.815
+ $Y=2.34 $X2=0.94 $Y2=2.485
r87 1 16 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.175
+ $Y=0.37 $X2=0.3 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRTP_2%SCE 3 6 7 8 11 13 17 21 23 24 25 26 27 28
+ 35 39
c67 39 0 1.61331e-19 $X=2.395 $Y=1.295
r68 39 41 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.395 $Y=1.295
+ $X2=2.395 $Y2=1.13
r69 39 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.395
+ $Y=1.295 $X2=2.395 $Y2=1.295
r70 35 37 47.6426 $w=4.75e-07 $l=1.65e-07 $layer=POLY_cond $X=0.677 $Y=1.295
+ $X2=0.677 $Y2=1.13
r71 28 40 15.096 $w=1.78e-07 $l=2.45e-07 $layer=LI1_cond $X=2.64 $Y=1.29
+ $X2=2.395 $Y2=1.29
r72 27 40 14.4798 $w=1.78e-07 $l=2.35e-07 $layer=LI1_cond $X=2.16 $Y=1.29
+ $X2=2.395 $Y2=1.29
r73 26 27 29.5758 $w=1.78e-07 $l=4.8e-07 $layer=LI1_cond $X=1.68 $Y=1.29
+ $X2=2.16 $Y2=1.29
r74 25 26 29.5758 $w=1.78e-07 $l=4.8e-07 $layer=LI1_cond $X=1.2 $Y=1.29 $X2=1.68
+ $Y2=1.29
r75 24 25 29.5758 $w=1.78e-07 $l=4.8e-07 $layer=LI1_cond $X=0.72 $Y=1.29 $X2=1.2
+ $Y2=1.29
r76 24 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.75
+ $Y=1.295 $X2=0.75 $Y2=1.295
r77 21 41 264.074 $w=1.5e-07 $l=5.15e-07 $layer=POLY_cond $X=2.485 $Y=0.615
+ $X2=2.485 $Y2=1.13
r78 15 17 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=1.585 $Y=2.21
+ $X2=1.585 $Y2=2.66
r79 14 23 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.23 $Y=2.135
+ $X2=1.155 $Y2=2.135
r80 13 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.51 $Y=2.135
+ $X2=1.585 $Y2=2.21
r81 13 14 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=1.51 $Y=2.135
+ $X2=1.23 $Y2=2.135
r82 9 23 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.155 $Y=2.21
+ $X2=1.155 $Y2=2.135
r83 9 11 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=1.155 $Y=2.21
+ $X2=1.155 $Y2=2.66
r84 7 23 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.08 $Y=2.135
+ $X2=1.155 $Y2=2.135
r85 7 8 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.08 $Y=2.135
+ $X2=0.915 $Y2=2.135
r86 6 8 37.7275 $w=1.5e-07 $l=2.72936e-07 $layer=POLY_cond $X=0.677 $Y=2.06
+ $X2=0.915 $Y2=2.135
r87 5 35 8.43012 $w=4.75e-07 $l=7.2e-08 $layer=POLY_cond $X=0.677 $Y=1.367
+ $X2=0.677 $Y2=1.295
r88 5 6 81.1399 $w=4.75e-07 $l=6.93e-07 $layer=POLY_cond $X=0.677 $Y=1.367
+ $X2=0.677 $Y2=2.06
r89 3 37 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=0.515 $Y=0.58
+ $X2=0.515 $Y2=1.13
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRTP_2%D 3 5 7 9 10 11 12 13
r36 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.825
+ $Y=1.655 $X2=1.825 $Y2=1.655
r37 12 13 25.3506 $w=2.08e-07 $l=4.8e-07 $layer=LI1_cond $X=2.16 $Y=1.655
+ $X2=2.64 $Y2=1.655
r38 12 21 17.6926 $w=2.08e-07 $l=3.35e-07 $layer=LI1_cond $X=2.16 $Y=1.655
+ $X2=1.825 $Y2=1.655
r39 11 21 7.65801 $w=2.08e-07 $l=1.45e-07 $layer=LI1_cond $X=1.68 $Y=1.655
+ $X2=1.825 $Y2=1.655
r40 10 11 25.3506 $w=2.08e-07 $l=4.8e-07 $layer=LI1_cond $X=1.2 $Y=1.655
+ $X2=1.68 $Y2=1.655
r41 9 10 25.3506 $w=2.08e-07 $l=4.8e-07 $layer=LI1_cond $X=0.72 $Y=1.655 $X2=1.2
+ $Y2=1.655
r42 5 20 38.7084 $w=3.43e-07 $l=2.11069e-07 $layer=POLY_cond $X=1.945 $Y=1.82
+ $X2=1.84 $Y2=1.655
r43 5 7 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=1.945 $Y=1.82
+ $X2=1.945 $Y2=2.66
r44 1 20 38.7084 $w=3.43e-07 $l=1.72337e-07 $layer=POLY_cond $X=1.825 $Y=1.49
+ $X2=1.84 $Y2=1.655
r45 1 3 528.149 $w=1.5e-07 $l=1.03e-06 $layer=POLY_cond $X=1.825 $Y=1.49
+ $X2=1.825 $Y2=0.46
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRTP_2%SCD 1 3 7 12 13 14 15 20
c46 3 0 1.91378e-19 $X=2.845 $Y=0.615
r47 20 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.99
+ $Y=1.49 $X2=2.99 $Y2=1.49
r48 14 15 11.2212 $w=3.78e-07 $l=3.7e-07 $layer=LI1_cond $X=3.095 $Y=1.665
+ $X2=3.095 $Y2=2.035
r49 14 21 5.3073 $w=3.78e-07 $l=1.75e-07 $layer=LI1_cond $X=3.095 $Y=1.665
+ $X2=3.095 $Y2=1.49
r50 13 21 5.91385 $w=3.78e-07 $l=1.95e-07 $layer=LI1_cond $X=3.095 $Y=1.295
+ $X2=3.095 $Y2=1.49
r51 11 20 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=2.99 $Y=1.845
+ $X2=2.99 $Y2=1.49
r52 11 12 43.5886 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=2.962 $Y=1.845
+ $X2=2.962 $Y2=1.995
r53 9 20 27.1035 $w=3.3e-07 $l=1.55e-07 $layer=POLY_cond $X=2.99 $Y=1.335
+ $X2=2.99 $Y2=1.49
r54 7 12 340.989 $w=1.5e-07 $l=6.65e-07 $layer=POLY_cond $X=2.845 $Y=2.66
+ $X2=2.845 $Y2=1.995
r55 1 9 33.318 $w=2.17e-07 $l=2.10357e-07 $layer=POLY_cond $X=2.845 $Y=1.185
+ $X2=2.99 $Y2=1.335
r56 1 3 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=2.845 $Y=1.185
+ $X2=2.845 $Y2=0.615
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRTP_2%A_756_265# 1 2 9 13 14 16 17 18 21 24 26 27
+ 29 31 35 36 38 39 40 41 42 43 46 55 59 63 64 65 67
c202 43 0 2.29156e-19 $X=7.585 $Y=1.295
c203 39 0 1.50829e-19 $X=4.225 $Y=1.295
c204 36 0 3.488e-20 $X=7.91 $Y=2.26
c205 35 0 7.03183e-20 $X=7.91 $Y=2.26
c206 31 0 1.46831e-19 $X=7.725 $Y=1.26
c207 9 0 1.50059e-19 $X=3.965 $Y=2.525
r208 70 71 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.44
+ $Y=1.26 $X2=7.44 $Y2=1.26
r209 67 70 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=7.44 $Y=1.17 $X2=7.44
+ $Y2=1.26
r210 63 65 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.9 $Y=1.29
+ $X2=4.9 $Y2=1.125
r211 63 64 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.9
+ $Y=1.29 $X2=4.9 $Y2=1.29
r212 59 60 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.945
+ $Y=1.49 $X2=3.945 $Y2=1.49
r213 56 87 5.81596 $w=4.51e-07 $l=2.15e-07 $layer=LI1_cond $X=10.455 $Y=1.295
+ $X2=10.455 $Y2=1.08
r214 55 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.32 $Y=1.295
+ $X2=10.32 $Y2=1.295
r215 52 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=1.295
+ $X2=7.44 $Y2=1.295
r216 49 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=1.295
+ $X2=5.04 $Y2=1.295
r217 46 60 6.15689 $w=3.63e-07 $l=1.95e-07 $layer=LI1_cond $X=4.032 $Y=1.295
+ $X2=4.032 $Y2=1.49
r218 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=1.295
+ $X2=4.08 $Y2=1.295
r219 43 52 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.585 $Y=1.295
+ $X2=7.44 $Y2=1.295
r220 42 55 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=10.175 $Y=1.295
+ $X2=10.32 $Y2=1.295
r221 42 43 3.20544 $w=1.4e-07 $l=2.59e-06 $layer=MET1_cond $X=10.175 $Y=1.295
+ $X2=7.585 $Y2=1.295
r222 41 49 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.185 $Y=1.295
+ $X2=5.04 $Y2=1.295
r223 40 52 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.295 $Y=1.295
+ $X2=7.44 $Y2=1.295
r224 40 41 2.61138 $w=1.4e-07 $l=2.11e-06 $layer=MET1_cond $X=7.295 $Y=1.295
+ $X2=5.185 $Y2=1.295
r225 39 45 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.225 $Y=1.295
+ $X2=4.08 $Y2=1.295
r226 38 49 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.895 $Y=1.295
+ $X2=5.04 $Y2=1.295
r227 38 39 0.829206 $w=1.4e-07 $l=6.7e-07 $layer=MET1_cond $X=4.895 $Y=1.295
+ $X2=4.225 $Y2=1.295
r228 36 73 24.4806 $w=3.3e-07 $l=1.4e-07 $layer=POLY_cond $X=7.91 $Y=2.26
+ $X2=7.77 $Y2=2.26
r229 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.91
+ $Y=2.26 $X2=7.91 $Y2=2.26
r230 32 35 4.43247 $w=2.58e-07 $l=1e-07 $layer=LI1_cond $X=7.81 $Y=2.225
+ $X2=7.91 $Y2=2.225
r231 31 71 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=7.725 $Y=1.26
+ $X2=7.44 $Y2=1.26
r232 27 56 5.68638 $w=4.51e-07 $l=1.52971e-07 $layer=LI1_cond $X=10.505 $Y=1.425
+ $X2=10.455 $Y2=1.295
r233 27 29 24.6002 $w=2.58e-07 $l=5.55e-07 $layer=LI1_cond $X=10.505 $Y=1.425
+ $X2=10.505 $Y2=1.98
r234 26 32 3.22376 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=7.81 $Y=2.095
+ $X2=7.81 $Y2=2.225
r235 25 31 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=7.81 $Y=1.425
+ $X2=7.725 $Y2=1.26
r236 25 26 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=7.81 $Y=1.425
+ $X2=7.81 $Y2=2.095
r237 23 59 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=3.945 $Y=1.83
+ $X2=3.945 $Y2=1.49
r238 23 24 38.6168 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.945 $Y=1.83
+ $X2=3.945 $Y2=1.995
r239 19 73 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.77 $Y=2.425
+ $X2=7.77 $Y2=2.26
r240 19 21 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=7.77 $Y=2.425
+ $X2=7.77 $Y2=2.88
r241 17 67 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.275 $Y=1.17
+ $X2=7.44 $Y2=1.17
r242 17 18 125.628 $w=1.5e-07 $l=2.45e-07 $layer=POLY_cond $X=7.275 $Y=1.17
+ $X2=7.03 $Y2=1.17
r243 14 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.955 $Y=1.095
+ $X2=7.03 $Y2=1.17
r244 14 16 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=6.955 $Y=1.095
+ $X2=6.955 $Y2=0.665
r245 13 65 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=4.88 $Y=0.805
+ $X2=4.88 $Y2=1.125
r246 9 24 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=3.965 $Y=2.525
+ $X2=3.965 $Y2=1.995
r247 2 29 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=10.415
+ $Y=1.835 $X2=10.54 $Y2=1.98
r248 1 87 182 $w=1.7e-07 $l=7.84156e-07 $layer=licon1_NDIFF $count=1 $X=10.39
+ $Y=0.365 $X2=10.535 $Y2=1.08
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRTP_2%A_936_333# 1 2 9 11 15 18 20 21 25 28 29 35
+ 39 44
c99 29 0 1.20546e-19 $X=4.867 $Y=1.685
r100 36 39 11.0909 $w=1.88e-07 $l=1.9e-07 $layer=LI1_cond $X=6.745 $Y=2.04
+ $X2=6.935 $Y2=2.04
r101 33 44 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.845 $Y=1.83
+ $X2=5.01 $Y2=1.83
r102 33 41 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=4.845 $Y=1.83
+ $X2=4.755 $Y2=1.83
r103 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.845
+ $Y=1.83 $X2=4.845 $Y2=1.83
r104 29 32 5.86331 $w=2.83e-07 $l=1.45e-07 $layer=LI1_cond $X=4.867 $Y=1.685
+ $X2=4.867 $Y2=1.83
r105 28 36 1.04402 $w=1.8e-07 $l=9.5e-08 $layer=LI1_cond $X=6.745 $Y=1.945
+ $X2=6.745 $Y2=2.04
r106 27 35 4.81226 $w=1.85e-07 $l=8.74643e-08 $layer=LI1_cond $X=6.745 $Y=1.77
+ $X2=6.74 $Y2=1.685
r107 27 28 10.7828 $w=1.78e-07 $l=1.75e-07 $layer=LI1_cond $X=6.745 $Y=1.77
+ $X2=6.745 $Y2=1.945
r108 23 35 4.81226 $w=1.85e-07 $l=8.5e-08 $layer=LI1_cond $X=6.74 $Y=1.6
+ $X2=6.74 $Y2=1.685
r109 23 25 64.7943 $w=1.88e-07 $l=1.11e-06 $layer=LI1_cond $X=6.74 $Y=1.6
+ $X2=6.74 $Y2=0.49
r110 22 29 3.76007 $w=1.7e-07 $l=1.43e-07 $layer=LI1_cond $X=5.01 $Y=1.685
+ $X2=4.867 $Y2=1.685
r111 21 35 1.64875 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=6.645 $Y=1.685
+ $X2=6.74 $Y2=1.685
r112 21 22 106.668 $w=1.68e-07 $l=1.635e-06 $layer=LI1_cond $X=6.645 $Y=1.685
+ $X2=5.01 $Y2=1.685
r113 19 20 58.3064 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=5.365 $Y=1.275
+ $X2=5.365 $Y2=1.425
r114 18 20 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=5.38 $Y=1.695
+ $X2=5.38 $Y2=1.425
r115 15 19 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=5.35 $Y=0.805 $X2=5.35
+ $Y2=1.275
r116 11 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.305 $Y=1.77
+ $X2=5.38 $Y2=1.695
r117 11 44 151.266 $w=1.5e-07 $l=2.95e-07 $layer=POLY_cond $X=5.305 $Y=1.77
+ $X2=5.01 $Y2=1.77
r118 7 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.755 $Y=1.995
+ $X2=4.755 $Y2=1.83
r119 7 9 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=4.755 $Y=1.995
+ $X2=4.755 $Y2=2.525
r120 2 39 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=6.795
+ $Y=1.895 $X2=6.935 $Y2=2.04
r121 1 25 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.6
+ $Y=0.345 $X2=6.74 $Y2=0.49
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRTP_2%RESET_B 4 5 6 9 11 12 14 15 17 19 20 21 27
+ 30 32 33 36 43 45 46 47 48 51 56 57 61 64 66 70
c203 56 0 9.68445e-20 $X=9.24 $Y=2.345
c204 30 0 2.88588e-20 $X=8.97 $Y=0.805
c205 4 0 1.06522e-19 $X=3.29 $Y=0.615
r206 64 67 14.8159 $w=3.7e-07 $l=9.5e-08 $layer=POLY_cond $X=5.94 $Y=2.035
+ $X2=5.94 $Y2=2.13
r207 64 66 46.7569 $w=3.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.94 $Y=2.035
+ $X2=5.94 $Y2=1.87
r208 61 64 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.96
+ $Y=2.035 $X2=5.96 $Y2=2.035
r209 57 71 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=9.24 $Y=2.345
+ $X2=9.24 $Y2=2.51
r210 57 70 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=9.24 $Y=2.345
+ $X2=9.24 $Y2=2.18
r211 56 59 9.25447 $w=3.28e-07 $l=2.65e-07 $layer=LI1_cond $X=9.24 $Y=2.345
+ $X2=9.24 $Y2=2.61
r212 56 57 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.24
+ $Y=2.345 $X2=9.24 $Y2=2.345
r213 51 53 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=6.84 $Y=2.39
+ $X2=6.84 $Y2=2.61
r214 50 61 9.42908 $w=3.28e-07 $l=2.7e-07 $layer=LI1_cond $X=5.96 $Y=2.305
+ $X2=5.96 $Y2=2.035
r215 49 53 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.925 $Y=2.61
+ $X2=6.84 $Y2=2.61
r216 48 59 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.075 $Y=2.61
+ $X2=9.24 $Y2=2.61
r217 48 49 140.267 $w=1.68e-07 $l=2.15e-06 $layer=LI1_cond $X=9.075 $Y=2.61
+ $X2=6.925 $Y2=2.61
r218 47 50 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.125 $Y=2.39
+ $X2=5.96 $Y2=2.305
r219 46 51 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.755 $Y=2.39
+ $X2=6.84 $Y2=2.39
r220 46 47 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=6.755 $Y=2.39
+ $X2=6.125 $Y2=2.39
r221 45 66 320.479 $w=1.5e-07 $l=6.25e-07 $layer=POLY_cond $X=5.83 $Y=1.245
+ $X2=5.83 $Y2=1.87
r222 44 45 58.3064 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=5.845 $Y=1.095
+ $X2=5.845 $Y2=1.245
r223 40 42 76.9149 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=3.29 $Y=1.01
+ $X2=3.44 $Y2=1.01
r224 38 70 264.074 $w=1.5e-07 $l=5.15e-07 $layer=POLY_cond $X=9.33 $Y=1.665
+ $X2=9.33 $Y2=2.18
r225 36 71 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=9.26 $Y=2.88
+ $X2=9.26 $Y2=2.51
r226 32 38 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.255 $Y=1.59
+ $X2=9.33 $Y2=1.665
r227 32 33 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=9.255 $Y=1.59
+ $X2=9.045 $Y2=1.59
r228 28 33 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.97 $Y=1.515
+ $X2=9.045 $Y2=1.59
r229 28 30 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=8.97 $Y=1.515
+ $X2=8.97 $Y2=0.805
r230 27 44 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=5.86 $Y=0.775
+ $X2=5.86 $Y2=1.095
r231 24 27 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=5.86 $Y=0.255
+ $X2=5.86 $Y2=0.775
r232 20 67 23.9667 $w=1.5e-07 $l=1.85e-07 $layer=POLY_cond $X=5.755 $Y=2.13
+ $X2=5.94 $Y2=2.13
r233 20 21 197.415 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=5.755 $Y=2.13
+ $X2=5.37 $Y2=2.13
r234 17 21 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.295 $Y=2.205
+ $X2=5.37 $Y2=2.13
r235 17 19 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=5.295 $Y=2.205
+ $X2=5.295 $Y2=2.525
r236 16 43 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.92 $Y=0.18
+ $X2=3.845 $Y2=0.18
r237 15 24 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.785 $Y=0.18
+ $X2=5.86 $Y2=0.255
r238 15 16 956.309 $w=1.5e-07 $l=1.865e-06 $layer=POLY_cond $X=5.785 $Y=0.18
+ $X2=3.92 $Y2=0.18
r239 13 43 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.845 $Y=0.255
+ $X2=3.845 $Y2=0.18
r240 13 14 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=3.845 $Y=0.255
+ $X2=3.845 $Y2=0.935
r241 12 42 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.515 $Y=1.01
+ $X2=3.44 $Y2=1.01
r242 11 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.77 $Y=1.01
+ $X2=3.845 $Y2=0.935
r243 11 12 130.755 $w=1.5e-07 $l=2.55e-07 $layer=POLY_cond $X=3.77 $Y=1.01
+ $X2=3.515 $Y2=1.01
r244 7 42 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.44 $Y=1.085
+ $X2=3.44 $Y2=1.01
r245 7 9 794.787 $w=1.5e-07 $l=1.55e-06 $layer=POLY_cond $X=3.44 $Y=1.085
+ $X2=3.44 $Y2=2.635
r246 5 43 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.77 $Y=0.18
+ $X2=3.845 $Y2=0.18
r247 5 6 207.67 $w=1.5e-07 $l=4.05e-07 $layer=POLY_cond $X=3.77 $Y=0.18
+ $X2=3.365 $Y2=0.18
r248 2 40 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.29 $Y=0.935
+ $X2=3.29 $Y2=1.01
r249 2 4 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=3.29 $Y=0.935
+ $X2=3.29 $Y2=0.615
r250 1 6 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.29 $Y=0.255
+ $X2=3.365 $Y2=0.18
r251 1 4 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=3.29 $Y=0.255
+ $X2=3.29 $Y2=0.615
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRTP_2%A_808_463# 1 2 3 10 12 15 19 22 23 25 29 33
+ 36 41 43
c119 41 0 1.20546e-19 $X=4.8 $Y=0.817
c120 15 0 9.3538e-21 $X=6.72 $Y=2.315
r121 40 41 6.28949 $w=3.53e-07 $l=1.35e-07 $layer=LI1_cond $X=4.665 $Y=0.817
+ $X2=4.8 $Y2=0.817
r122 37 40 6.33032 $w=3.53e-07 $l=1.95e-07 $layer=LI1_cond $X=4.47 $Y=0.817
+ $X2=4.665 $Y2=0.817
r123 34 43 31.9846 $w=3.24e-07 $l=2.15e-07 $layer=POLY_cond $X=6.31 $Y=1.365
+ $X2=6.525 $Y2=1.365
r124 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.31
+ $Y=1.26 $X2=6.31 $Y2=1.26
r125 31 33 9.25447 $w=3.28e-07 $l=2.65e-07 $layer=LI1_cond $X=6.31 $Y=0.995
+ $X2=6.31 $Y2=1.26
r126 27 29 7.89637 $w=2.68e-07 $l=1.85e-07 $layer=LI1_cond $X=5.49 $Y=2.345
+ $X2=5.49 $Y2=2.53
r127 25 31 7.26367 $w=2.1e-07 $l=2.11069e-07 $layer=LI1_cond $X=6.145 $Y=0.89
+ $X2=6.31 $Y2=0.995
r128 25 41 71.0346 $w=2.08e-07 $l=1.345e-06 $layer=LI1_cond $X=6.145 $Y=0.89
+ $X2=4.8 $Y2=0.89
r129 24 36 2.76166 $w=1.7e-07 $l=2.5e-07 $layer=LI1_cond $X=4.555 $Y=2.26
+ $X2=4.305 $Y2=2.26
r130 23 27 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=5.355 $Y=2.26
+ $X2=5.49 $Y2=2.345
r131 23 24 52.1925 $w=1.68e-07 $l=8e-07 $layer=LI1_cond $X=5.355 $Y=2.26
+ $X2=4.555 $Y2=2.26
r132 22 36 3.70735 $w=2.5e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.47 $Y=2.175
+ $X2=4.305 $Y2=2.26
r133 21 37 5.0588 $w=1.7e-07 $l=1.78e-07 $layer=LI1_cond $X=4.47 $Y=0.995
+ $X2=4.47 $Y2=0.817
r134 21 22 76.984 $w=1.68e-07 $l=1.18e-06 $layer=LI1_cond $X=4.47 $Y=0.995
+ $X2=4.47 $Y2=2.175
r135 17 36 3.70735 $w=2.5e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.22 $Y=2.345
+ $X2=4.305 $Y2=2.26
r136 17 19 6.46067 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=4.22 $Y=2.345
+ $X2=4.22 $Y2=2.53
r137 13 43 29.0093 $w=3.24e-07 $l=3.5433e-07 $layer=POLY_cond $X=6.72 $Y=1.635
+ $X2=6.525 $Y2=1.365
r138 13 15 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=6.72 $Y=1.635
+ $X2=6.72 $Y2=2.315
r139 10 43 20.7868 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=6.525 $Y=1.095
+ $X2=6.525 $Y2=1.365
r140 10 12 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=6.525 $Y=1.095
+ $X2=6.525 $Y2=0.665
r141 3 29 600 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_PDIFF $count=1 $X=5.37
+ $Y=2.315 $X2=5.51 $Y2=2.53
r142 2 19 600 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_PDIFF $count=1 $X=4.04
+ $Y=2.315 $X2=4.18 $Y2=2.53
r143 1 40 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=4.525
+ $Y=0.595 $X2=4.665 $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRTP_2%A_864_255# 1 2 10 13 15 16 20 21 22 25 29
+ 33 36 38 39 40 42 43 44 45 46 48 51 56 57 61
c198 56 0 3.25675e-20 $X=10.89 $Y=1.51
c199 51 0 1.2669e-20 $X=8.16 $Y=1.72
c200 45 0 1.04785e-19 $X=11.132 $Y=1.672
c201 40 0 1.90875e-19 $X=8.325 $Y=1.645
c202 39 0 1.47127e-19 $X=9.935 $Y=1.645
c203 38 0 1.77274e-19 $X=7.89 $Y=1.72
c204 21 0 5.76493e-20 $X=7.815 $Y=1.71
r205 58 61 7.40856 $w=2.78e-07 $l=1.8e-07 $layer=LI1_cond $X=11.375 $Y=2.8
+ $X2=11.555 $Y2=2.8
r206 56 67 45.2517 $w=3.8e-07 $l=1.65e-07 $layer=POLY_cond $X=10.865 $Y=1.51
+ $X2=10.865 $Y2=1.675
r207 56 66 45.2517 $w=3.8e-07 $l=1.65e-07 $layer=POLY_cond $X=10.865 $Y=1.51
+ $X2=10.865 $Y2=1.345
r208 55 56 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.89
+ $Y=1.51 $X2=10.89 $Y2=1.51
r209 53 55 10.513 $w=4.99e-07 $l=6.90293e-07 $layer=LI1_cond $X=11.555 $Y=1.08
+ $X2=11.047 $Y2=1.51
r210 50 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.16
+ $Y=1.72 $X2=8.16 $Y2=1.72
r211 48 58 3.65648 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=11.375 $Y=2.66
+ $X2=11.375 $Y2=2.8
r212 47 57 2.35019 $w=4.12e-07 $l=2.82319e-07 $layer=LI1_cond $X=11.375 $Y=2.495
+ $X2=11.132 $Y2=2.41
r213 47 48 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=11.375 $Y=2.495
+ $X2=11.375 $Y2=2.66
r214 46 57 2.35019 $w=4.12e-07 $l=8.5e-08 $layer=LI1_cond $X=11.132 $Y=2.325
+ $X2=11.132 $Y2=2.41
r215 45 55 3.73927 $w=6.55e-07 $l=2.00035e-07 $layer=LI1_cond $X=11.132 $Y=1.672
+ $X2=11.047 $Y2=1.51
r216 45 46 11.9243 $w=6.53e-07 $l=6.53e-07 $layer=LI1_cond $X=11.132 $Y=1.672
+ $X2=11.132 $Y2=2.325
r217 43 57 4.66114 $w=1.7e-07 $l=3.27e-07 $layer=LI1_cond $X=10.805 $Y=2.41
+ $X2=11.132 $Y2=2.41
r218 43 44 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=10.805 $Y=2.41
+ $X2=10.105 $Y2=2.41
r219 42 44 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.02 $Y=2.325
+ $X2=10.105 $Y2=2.41
r220 41 42 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=10.02 $Y=1.73
+ $X2=10.02 $Y2=2.325
r221 40 50 8.95713 $w=3.28e-07 $l=1.98997e-07 $layer=LI1_cond $X=8.325 $Y=1.645
+ $X2=8.16 $Y2=1.72
r222 39 41 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.935 $Y=1.645
+ $X2=10.02 $Y2=1.73
r223 39 40 105.037 $w=1.68e-07 $l=1.61e-06 $layer=LI1_cond $X=9.935 $Y=1.645
+ $X2=8.325 $Y2=1.645
r224 37 51 34.0979 $w=3.3e-07 $l=1.95e-07 $layer=POLY_cond $X=7.965 $Y=1.72
+ $X2=8.16 $Y2=1.72
r225 37 38 13.5877 $w=2.4e-07 $l=7.5e-08 $layer=POLY_cond $X=7.965 $Y=1.72
+ $X2=7.89 $Y2=1.72
r226 35 36 48.5235 $w=2.05e-07 $l=1.5e-07 $layer=POLY_cond $X=4.422 $Y=1.275
+ $X2=4.422 $Y2=1.425
r227 33 67 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=10.755 $Y=2.465
+ $X2=10.755 $Y2=1.675
r228 29 66 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=10.75 $Y=0.785
+ $X2=10.75 $Y2=1.345
r229 23 38 12.1617 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.89 $Y=1.555
+ $X2=7.89 $Y2=1.72
r230 23 25 399.957 $w=1.5e-07 $l=7.8e-07 $layer=POLY_cond $X=7.89 $Y=1.555
+ $X2=7.89 $Y2=0.775
r231 21 38 13.5877 $w=2.4e-07 $l=7.98436e-08 $layer=POLY_cond $X=7.815 $Y=1.71
+ $X2=7.89 $Y2=1.72
r232 21 22 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=7.815 $Y=1.71
+ $X2=7.225 $Y2=1.71
r233 18 20 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=7.15 $Y=3.075
+ $X2=7.15 $Y2=2.315
r234 17 22 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.15 $Y=1.785
+ $X2=7.225 $Y2=1.71
r235 17 20 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=7.15 $Y=1.785
+ $X2=7.15 $Y2=2.315
r236 15 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.075 $Y=3.15
+ $X2=7.15 $Y2=3.075
r237 15 16 1335.76 $w=1.5e-07 $l=2.605e-06 $layer=POLY_cond $X=7.075 $Y=3.15
+ $X2=4.47 $Y2=3.15
r238 13 35 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=4.45 $Y=0.805 $X2=4.45
+ $Y2=1.275
r239 10 36 564.043 $w=1.5e-07 $l=1.1e-06 $layer=POLY_cond $X=4.395 $Y=2.525
+ $X2=4.395 $Y2=1.425
r240 8 16 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.395 $Y=3.075
+ $X2=4.47 $Y2=3.15
r241 8 10 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=4.395 $Y=3.075
+ $X2=4.395 $Y2=2.525
r242 2 61 600 $w=1.7e-07 $l=9.97547e-07 $layer=licon1_PDIFF $count=1 $X=11.415
+ $Y=1.835 $X2=11.555 $Y2=2.765
r243 1 53 182 $w=1.7e-07 $l=7.81873e-07 $layer=licon1_NDIFF $count=1 $X=11.415
+ $Y=0.365 $X2=11.555 $Y2=1.08
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRTP_2%A_1406_69# 1 2 7 9 10 11 14 18 22 24 27 28
+ 29 30 34 36 39 40 41 46 47 48 50 60 62
c197 41 0 1.33016e-19 $X=8.235 $Y=1.29
c198 39 0 9.61405e-20 $X=8.15 $Y=1.205
c199 36 0 9.3538e-21 $X=7.405 $Y=2.19
c200 34 0 1.77274e-19 $X=7.412 $Y=1.775
c201 11 0 1.47127e-19 $X=9.405 $Y=1.2
r202 59 60 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=12.375
+ $Y=1.08 $X2=12.375 $Y2=1.08
r203 50 59 12.3906 $w=3.84e-07 $l=5.01548e-07 $layer=LI1_cond $X=11.985 $Y=0.995
+ $X2=12.375 $Y2=1.25
r204 49 50 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=11.985 $Y=0.815
+ $X2=11.985 $Y2=0.995
r205 47 49 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=11.9 $Y=0.73
+ $X2=11.985 $Y2=0.815
r206 47 48 123.957 $w=1.68e-07 $l=1.9e-06 $layer=LI1_cond $X=11.9 $Y=0.73 $X2=10
+ $Y2=0.73
r207 45 48 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.915 $Y=0.815
+ $X2=10 $Y2=0.73
r208 45 46 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=9.915 $Y=0.815
+ $X2=9.915 $Y2=1.205
r209 44 65 53.2059 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=9.78 $Y=1.29
+ $X2=9.78 $Y2=1.495
r210 44 62 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=9.78 $Y=1.29 $X2=9.78
+ $Y2=1.2
r211 43 44 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.78
+ $Y=1.29 $X2=9.78 $Y2=1.29
r212 41 43 100.797 $w=1.68e-07 $l=1.545e-06 $layer=LI1_cond $X=8.235 $Y=1.29
+ $X2=9.78 $Y2=1.29
r213 40 46 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.83 $Y=1.29
+ $X2=9.915 $Y2=1.205
r214 40 43 3.26203 $w=1.68e-07 $l=5e-08 $layer=LI1_cond $X=9.83 $Y=1.29 $X2=9.78
+ $Y2=1.29
r215 39 41 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.15 $Y=1.205
+ $X2=8.235 $Y2=1.29
r216 38 39 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=8.15 $Y=0.925
+ $X2=8.15 $Y2=1.205
r217 34 53 21.0075 $w=1.68e-07 $l=3.22e-07 $layer=LI1_cond $X=7.412 $Y=1.69
+ $X2=7.09 $Y2=1.69
r218 34 36 16.7812 $w=2.83e-07 $l=4.15e-07 $layer=LI1_cond $X=7.412 $Y=1.775
+ $X2=7.412 $Y2=2.19
r219 31 52 2.21775 $w=6e-07 $l=8.5e-08 $layer=LI1_cond $X=7.175 $Y=0.625
+ $X2=7.09 $Y2=0.625
r220 31 33 9.96732 $w=5.98e-07 $l=5e-07 $layer=LI1_cond $X=7.175 $Y=0.625
+ $X2=7.675 $Y2=0.625
r221 30 38 10.0451 $w=6e-07 $l=3.39853e-07 $layer=LI1_cond $X=8.065 $Y=0.625
+ $X2=8.15 $Y2=0.925
r222 30 33 7.77451 $w=5.98e-07 $l=3.9e-07 $layer=LI1_cond $X=8.065 $Y=0.625
+ $X2=7.675 $Y2=0.625
r223 29 53 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.09 $Y=1.605
+ $X2=7.09 $Y2=1.69
r224 28 52 7.82736 $w=1.7e-07 $l=3e-07 $layer=LI1_cond $X=7.09 $Y=0.925 $X2=7.09
+ $Y2=0.625
r225 28 29 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=7.09 $Y=0.925
+ $X2=7.09 $Y2=1.605
r226 26 60 52.0941 $w=3.6e-07 $l=3.25e-07 $layer=POLY_cond $X=12.39 $Y=1.405
+ $X2=12.39 $Y2=1.08
r227 26 27 48.987 $w=3.6e-07 $l=1.8e-07 $layer=POLY_cond $X=12.39 $Y=1.405
+ $X2=12.39 $Y2=1.585
r228 24 60 7.21303 $w=3.6e-07 $l=4.5e-08 $layer=POLY_cond $X=12.39 $Y=1.035
+ $X2=12.39 $Y2=1.08
r229 24 25 48.987 $w=3.6e-07 $l=1.8e-07 $layer=POLY_cond $X=12.39 $Y=1.035
+ $X2=12.39 $Y2=0.855
r230 22 27 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=12.495 $Y=2.155
+ $X2=12.495 $Y2=1.585
r231 18 25 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=12.495 $Y=0.445
+ $X2=12.495 $Y2=0.855
r232 14 65 710.181 $w=1.5e-07 $l=1.385e-06 $layer=POLY_cond $X=9.69 $Y=2.88
+ $X2=9.69 $Y2=1.495
r233 10 62 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.615 $Y=1.2
+ $X2=9.78 $Y2=1.2
r234 10 11 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=9.615 $Y=1.2
+ $X2=9.405 $Y2=1.2
r235 7 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.33 $Y=1.125
+ $X2=9.405 $Y2=1.2
r236 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=9.33 $Y=1.125
+ $X2=9.33 $Y2=0.805
r237 2 36 600 $w=1.7e-07 $l=3.74333e-07 $layer=licon1_PDIFF $count=1 $X=7.225
+ $Y=1.895 $X2=7.405 $Y2=2.19
r238 1 52 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=7.03
+ $Y=0.345 $X2=7.17 $Y2=0.49
r239 1 33 182 $w=1.7e-07 $l=8.26862e-07 $layer=licon1_NDIFF $count=1 $X=7.03
+ $Y=0.345 $X2=7.675 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRTP_2%A_1635_21# 1 2 10 13 15 16 17 18 20 21 23
+ 29 32 33 35 38 45 47
c117 45 0 9.68445e-20 $X=8.61 $Y=2.11
c118 33 0 2.88588e-20 $X=9.66 $Y=0.365
c119 18 0 3.02826e-19 $X=8.325 $Y=1.17
r120 42 45 17.2143 $w=2.52e-07 $l=9e-08 $layer=POLY_cond $X=8.7 $Y=2.11 $X2=8.61
+ $Y2=2.11
r121 41 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.7
+ $Y=2.11 $X2=8.7 $Y2=2.11
r122 38 41 4.01609 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=8.7 $Y=1.995
+ $X2=8.7 $Y2=2.11
r123 36 47 29.7264 $w=3.3e-07 $l=1.7e-07 $layer=POLY_cond $X=9.945 $Y=0.35
+ $X2=9.945 $Y2=0.18
r124 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.945
+ $Y=0.35 $X2=9.945 $Y2=0.35
r125 33 35 14.9294 $w=2.18e-07 $l=2.85e-07 $layer=LI1_cond $X=9.66 $Y=0.365
+ $X2=9.945 $Y2=0.365
r126 31 32 51.2139 $w=1.68e-07 $l=7.85e-07 $layer=LI1_cond $X=9.67 $Y=2.08
+ $X2=9.67 $Y2=2.865
r127 27 33 6.94494 $w=2.2e-07 $l=1.87083e-07 $layer=LI1_cond $X=9.52 $Y=0.475
+ $X2=9.66 $Y2=0.365
r128 27 29 13.5824 $w=2.78e-07 $l=3.3e-07 $layer=LI1_cond $X=9.52 $Y=0.475
+ $X2=9.52 $Y2=0.805
r129 23 32 6.91519 $w=2.1e-07 $l=1.41244e-07 $layer=LI1_cond $X=9.585 $Y=2.97
+ $X2=9.67 $Y2=2.865
r130 23 25 5.80952 $w=2.08e-07 $l=1.1e-07 $layer=LI1_cond $X=9.585 $Y=2.97
+ $X2=9.475 $Y2=2.97
r131 22 38 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.865 $Y=1.995
+ $X2=8.7 $Y2=1.995
r132 21 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.585 $Y=1.995
+ $X2=9.67 $Y2=2.08
r133 21 22 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=9.585 $Y=1.995
+ $X2=8.865 $Y2=1.995
r134 20 45 14.904 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.61 $Y=1.945
+ $X2=8.61 $Y2=2.11
r135 19 20 358.936 $w=1.5e-07 $l=7e-07 $layer=POLY_cond $X=8.61 $Y=1.245
+ $X2=8.61 $Y2=1.945
r136 17 19 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.535 $Y=1.17
+ $X2=8.61 $Y2=1.245
r137 17 18 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=8.535 $Y=1.17
+ $X2=8.325 $Y2=1.17
r138 15 47 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.78 $Y=0.18
+ $X2=9.945 $Y2=0.18
r139 15 16 746.074 $w=1.5e-07 $l=1.455e-06 $layer=POLY_cond $X=9.78 $Y=0.18
+ $X2=8.325 $Y2=0.18
r140 11 45 47.8175 $w=2.52e-07 $l=3.22102e-07 $layer=POLY_cond $X=8.36 $Y=2.275
+ $X2=8.61 $Y2=2.11
r141 11 13 310.223 $w=1.5e-07 $l=6.05e-07 $layer=POLY_cond $X=8.36 $Y=2.275
+ $X2=8.36 $Y2=2.88
r142 8 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.25 $Y=1.095
+ $X2=8.325 $Y2=1.17
r143 8 10 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=8.25 $Y=1.095
+ $X2=8.25 $Y2=0.775
r144 7 16 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.25 $Y=0.255
+ $X2=8.325 $Y2=0.18
r145 7 10 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=8.25 $Y=0.255
+ $X2=8.25 $Y2=0.775
r146 2 25 600 $w=1.7e-07 $l=3.53129e-07 $layer=licon1_PDIFF $count=1 $X=9.335
+ $Y=2.67 $X2=9.475 $Y2=2.96
r147 1 29 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=9.405
+ $Y=0.595 $X2=9.545 $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRTP_2%CLK 3 7 9 11 12 13 14 18 22
c46 22 0 3.25675e-20 $X=11.805 $Y=1.51
r47 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.805
+ $Y=1.51 $X2=11.805 $Y2=1.51
r48 18 21 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=11.805 $Y=1.42
+ $X2=11.805 $Y2=1.51
r49 13 14 11.3708 $w=3.73e-07 $l=3.7e-07 $layer=LI1_cond $X=11.817 $Y=2.035
+ $X2=11.817 $Y2=2.405
r50 12 13 11.3708 $w=3.73e-07 $l=3.7e-07 $layer=LI1_cond $X=11.817 $Y=1.665
+ $X2=11.817 $Y2=2.035
r51 12 22 4.76343 $w=3.73e-07 $l=1.55e-07 $layer=LI1_cond $X=11.817 $Y=1.665
+ $X2=11.817 $Y2=1.51
r52 10 11 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=11.415 $Y=1.42
+ $X2=11.34 $Y2=1.42
r53 9 18 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=11.64 $Y=1.42
+ $X2=11.805 $Y2=1.42
r54 9 10 115.372 $w=1.5e-07 $l=2.25e-07 $layer=POLY_cond $X=11.64 $Y=1.42
+ $X2=11.415 $Y2=1.42
r55 5 11 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=11.34 $Y=1.495
+ $X2=11.34 $Y2=1.42
r56 5 7 497.383 $w=1.5e-07 $l=9.7e-07 $layer=POLY_cond $X=11.34 $Y=1.495
+ $X2=11.34 $Y2=2.465
r57 1 11 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=11.34 $Y=1.345
+ $X2=11.34 $Y2=1.42
r58 1 3 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=11.34 $Y=1.345
+ $X2=11.34 $Y2=0.785
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRTP_2%A_2431_47# 1 2 9 13 17 21 25 28 29 30 31 32
+ 34 36 40 46
r88 45 46 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=13.005 $Y=1.41
+ $X2=13.435 $Y2=1.41
r89 41 45 10.4917 $w=3.3e-07 $l=6e-08 $layer=POLY_cond $X=12.945 $Y=1.41
+ $X2=13.005 $Y2=1.41
r90 40 42 17.2874 $w=2.47e-07 $l=3.5e-07 $layer=LI1_cond $X=12.875 $Y=1.41
+ $X2=12.875 $Y2=1.76
r91 40 41 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=12.945
+ $Y=1.41 $X2=12.945 $Y2=1.41
r92 34 40 8.27038 $w=2.47e-07 $l=1.85257e-07 $layer=LI1_cond $X=12.832 $Y=1.245
+ $X2=12.875 $Y2=1.41
r93 33 34 22.0245 $w=2.23e-07 $l=4.3e-07 $layer=LI1_cond $X=12.832 $Y=0.815
+ $X2=12.832 $Y2=1.245
r94 31 33 6.9898 $w=1.7e-07 $l=1.4854e-07 $layer=LI1_cond $X=12.72 $Y=0.73
+ $X2=12.832 $Y2=0.815
r95 31 32 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=12.72 $Y=0.73
+ $X2=12.445 $Y2=0.73
r96 29 42 2.92482 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=12.72 $Y=1.76
+ $X2=12.875 $Y2=1.76
r97 29 30 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=12.72 $Y=1.76
+ $X2=12.375 $Y2=1.76
r98 28 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=12.36 $Y=0.645
+ $X2=12.445 $Y2=0.73
r99 27 36 1.386 $w=1.7e-07 $l=1.28938e-07 $layer=LI1_cond $X=12.36 $Y=0.465
+ $X2=12.28 $Y2=0.37
r100 27 28 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=12.36 $Y=0.465
+ $X2=12.36 $Y2=0.645
r101 23 30 6.87494 $w=1.7e-07 $l=1.36015e-07 $layer=LI1_cond $X=12.275 $Y=1.845
+ $X2=12.375 $Y2=1.76
r102 23 25 7.48636 $w=1.98e-07 $l=1.35e-07 $layer=LI1_cond $X=12.275 $Y=1.845
+ $X2=12.275 $Y2=1.98
r103 19 46 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=13.435 $Y=1.575
+ $X2=13.435 $Y2=1.41
r104 19 21 456.362 $w=1.5e-07 $l=8.9e-07 $layer=POLY_cond $X=13.435 $Y=1.575
+ $X2=13.435 $Y2=2.465
r105 15 46 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=13.435 $Y=1.245
+ $X2=13.435 $Y2=1.41
r106 15 17 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=13.435 $Y=1.245
+ $X2=13.435 $Y2=0.655
r107 11 45 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=13.005 $Y=1.575
+ $X2=13.005 $Y2=1.41
r108 11 13 456.362 $w=1.5e-07 $l=8.9e-07 $layer=POLY_cond $X=13.005 $Y=1.575
+ $X2=13.005 $Y2=2.465
r109 7 45 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=13.005 $Y=1.245
+ $X2=13.005 $Y2=1.41
r110 7 9 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=13.005 $Y=1.245
+ $X2=13.005 $Y2=0.655
r111 2 25 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=12.155
+ $Y=1.835 $X2=12.28 $Y2=1.98
r112 1 36 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=12.155
+ $Y=0.235 $X2=12.28 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRTP_2%VPWR 1 2 3 4 5 6 7 8 9 30 34 38 42 46 50 54
+ 58 60 65 66 68 69 71 72 73 82 89 97 117 124 130 133 136 141 144 146 150
r161 149 150 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.68 $Y=3.33
+ $X2=13.68 $Y2=3.33
r162 146 147 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.72 $Y=3.33
+ $X2=12.72 $Y2=3.33
r163 143 144 9.83198 $w=5.48e-07 $l=1.65e-07 $layer=LI1_cond $X=8.975 $Y=3.14
+ $X2=9.14 $Y2=3.14
r164 139 143 2.06595 $w=5.48e-07 $l=9.5e-08 $layer=LI1_cond $X=8.88 $Y=3.14
+ $X2=8.975 $Y2=3.14
r165 139 141 16.4648 $w=5.48e-07 $l=4.7e-07 $layer=LI1_cond $X=8.88 $Y=3.14
+ $X2=8.41 $Y2=3.14
r166 139 140 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r167 136 137 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r168 133 134 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r169 130 131 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r170 128 150 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.2 $Y=3.33
+ $X2=13.68 $Y2=3.33
r171 128 147 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.2 $Y=3.33
+ $X2=12.72 $Y2=3.33
r172 127 128 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.2 $Y=3.33
+ $X2=13.2 $Y2=3.33
r173 125 146 9.81116 $w=1.7e-07 $l=2e-07 $layer=LI1_cond $X=12.945 $Y=3.33
+ $X2=12.745 $Y2=3.33
r174 125 127 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=12.945 $Y=3.33
+ $X2=13.2 $Y2=3.33
r175 124 149 4.20444 $w=1.7e-07 $l=1.87e-07 $layer=LI1_cond $X=13.545 $Y=3.33
+ $X2=13.732 $Y2=3.33
r176 124 127 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=13.545 $Y=3.33
+ $X2=13.2 $Y2=3.33
r177 123 147 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.24 $Y=3.33
+ $X2=12.72 $Y2=3.33
r178 122 123 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=12.24 $Y=3.33
+ $X2=12.24 $Y2=3.33
r179 120 123 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=11.28 $Y=3.33
+ $X2=12.24 $Y2=3.33
r180 119 122 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=11.28 $Y=3.33
+ $X2=12.24 $Y2=3.33
r181 119 120 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=11.28 $Y=3.33
+ $X2=11.28 $Y2=3.33
r182 117 146 9.81116 $w=1.7e-07 $l=2e-07 $layer=LI1_cond $X=12.545 $Y=3.33
+ $X2=12.745 $Y2=3.33
r183 117 122 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=12.545 $Y=3.33
+ $X2=12.24 $Y2=3.33
r184 116 120 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.8 $Y=3.33
+ $X2=11.28 $Y2=3.33
r185 115 116 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.8 $Y=3.33
+ $X2=10.8 $Y2=3.33
r186 113 116 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=9.84 $Y=3.33
+ $X2=10.8 $Y2=3.33
r187 113 140 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=9.84 $Y=3.33
+ $X2=8.88 $Y2=3.33
r188 112 144 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=9.84 $Y=3.33
+ $X2=9.14 $Y2=3.33
r189 112 113 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r190 109 140 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=8.88 $Y2=3.33
r191 108 141 0.652406 $w=1.68e-07 $l=1e-08 $layer=LI1_cond $X=8.4 $Y=3.33
+ $X2=8.41 $Y2=3.33
r192 108 109 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r193 105 108 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=6.96 $Y=3.33
+ $X2=8.4 $Y2=3.33
r194 103 136 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.575 $Y=3.33
+ $X2=6.41 $Y2=3.33
r195 103 105 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=6.575 $Y=3.33
+ $X2=6.96 $Y2=3.33
r196 101 137 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33
+ $X2=6.48 $Y2=3.33
r197 101 134 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=3.33
+ $X2=5.04 $Y2=3.33
r198 100 101 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r199 98 133 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.185 $Y=3.33
+ $X2=5.02 $Y2=3.33
r200 98 100 53.1711 $w=1.68e-07 $l=8.15e-07 $layer=LI1_cond $X=5.185 $Y=3.33
+ $X2=6 $Y2=3.33
r201 97 136 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.245 $Y=3.33
+ $X2=6.41 $Y2=3.33
r202 97 100 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=6.245 $Y=3.33
+ $X2=6 $Y2=3.33
r203 96 134 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.04 $Y2=3.33
r204 95 96 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r205 93 96 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.56 $Y2=3.33
r206 93 131 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=3.12 $Y2=3.33
r207 92 95 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=3.6 $Y=3.33 $X2=4.56
+ $Y2=3.33
r208 92 93 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r209 90 130 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.3 $Y=3.33
+ $X2=3.135 $Y2=3.33
r210 90 92 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=3.3 $Y=3.33 $X2=3.6
+ $Y2=3.33
r211 89 133 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.855 $Y=3.33
+ $X2=5.02 $Y2=3.33
r212 89 95 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=4.855 $Y=3.33
+ $X2=4.56 $Y2=3.33
r213 88 131 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r214 87 88 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r215 85 88 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r216 84 87 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r217 84 85 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r218 82 130 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.97 $Y=3.33
+ $X2=3.135 $Y2=3.33
r219 82 87 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=2.97 $Y=3.33
+ $X2=2.64 $Y2=3.33
r220 81 85 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r221 80 81 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r222 77 81 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.2 $Y2=3.33
r223 76 80 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.24 $Y=3.33 $X2=1.2
+ $Y2=3.33
r224 76 77 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r225 73 109 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=8.4 $Y2=3.33
r226 73 137 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=6.48 $Y2=3.33
r227 73 105 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r228 71 115 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=10.805 $Y=3.33
+ $X2=10.8 $Y2=3.33
r229 71 72 8.33247 $w=1.7e-07 $l=1.57e-07 $layer=LI1_cond $X=10.805 $Y=3.33
+ $X2=10.962 $Y2=3.33
r230 70 119 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=11.12 $Y=3.33
+ $X2=11.28 $Y2=3.33
r231 70 72 8.33247 $w=1.7e-07 $l=1.58e-07 $layer=LI1_cond $X=11.12 $Y=3.33
+ $X2=10.962 $Y2=3.33
r232 68 112 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=9.925 $Y=3.33
+ $X2=9.84 $Y2=3.33
r233 68 69 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.925 $Y=3.33
+ $X2=10.05 $Y2=3.33
r234 67 115 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=10.175 $Y=3.33
+ $X2=10.8 $Y2=3.33
r235 67 69 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.175 $Y=3.33
+ $X2=10.05 $Y2=3.33
r236 65 80 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=1.205 $Y=3.33
+ $X2=1.2 $Y2=3.33
r237 65 66 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=1.205 $Y=3.33
+ $X2=1.34 $Y2=3.33
r238 64 84 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=1.475 $Y=3.33
+ $X2=1.68 $Y2=3.33
r239 64 66 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=1.475 $Y=3.33
+ $X2=1.34 $Y2=3.33
r240 60 63 41.4026 $w=2.68e-07 $l=9.7e-07 $layer=LI1_cond $X=13.68 $Y=1.98
+ $X2=13.68 $Y2=2.95
r241 58 149 3.08026 $w=2.7e-07 $l=1.07912e-07 $layer=LI1_cond $X=13.68 $Y=3.245
+ $X2=13.732 $Y2=3.33
r242 58 63 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=13.68 $Y=3.245
+ $X2=13.68 $Y2=2.95
r243 54 57 12.2447 $w=3.98e-07 $l=4.25e-07 $layer=LI1_cond $X=12.745 $Y=2.1
+ $X2=12.745 $Y2=2.525
r244 52 146 1.46811 $w=4e-07 $l=8.5e-08 $layer=LI1_cond $X=12.745 $Y=3.245
+ $X2=12.745 $Y2=3.33
r245 52 57 20.744 $w=3.98e-07 $l=7.2e-07 $layer=LI1_cond $X=12.745 $Y=3.245
+ $X2=12.745 $Y2=2.525
r246 48 72 0.751525 $w=3.15e-07 $l=8.5e-08 $layer=LI1_cond $X=10.962 $Y=3.245
+ $X2=10.962 $Y2=3.33
r247 48 50 15.183 $w=3.13e-07 $l=4.15e-07 $layer=LI1_cond $X=10.962 $Y=3.245
+ $X2=10.962 $Y2=2.83
r248 44 69 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=10.05 $Y=3.245
+ $X2=10.05 $Y2=3.33
r249 44 46 17.2866 $w=2.48e-07 $l=3.75e-07 $layer=LI1_cond $X=10.05 $Y=3.245
+ $X2=10.05 $Y2=2.87
r250 40 136 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.41 $Y=3.245
+ $X2=6.41 $Y2=3.33
r251 40 42 17.6359 $w=3.28e-07 $l=5.05e-07 $layer=LI1_cond $X=6.41 $Y=3.245
+ $X2=6.41 $Y2=2.74
r252 36 133 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.02 $Y=3.245
+ $X2=5.02 $Y2=3.33
r253 36 38 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=5.02 $Y=3.245
+ $X2=5.02 $Y2=2.61
r254 32 130 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.135 $Y=3.245
+ $X2=3.135 $Y2=3.33
r255 32 34 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=3.135 $Y=3.245
+ $X2=3.135 $Y2=2.765
r256 28 66 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.34 $Y=3.245
+ $X2=1.34 $Y2=3.33
r257 28 30 32.4391 $w=2.68e-07 $l=7.6e-07 $layer=LI1_cond $X=1.34 $Y=3.245
+ $X2=1.34 $Y2=2.485
r258 9 63 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=13.51
+ $Y=1.835 $X2=13.65 $Y2=2.95
r259 9 60 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=13.51
+ $Y=1.835 $X2=13.65 $Y2=1.98
r260 8 57 300 $w=1.7e-07 $l=7.92401e-07 $layer=licon1_PDIFF $count=2 $X=12.57
+ $Y=1.835 $X2=12.79 $Y2=2.525
r261 8 54 600 $w=1.7e-07 $l=3.27605e-07 $layer=licon1_PDIFF $count=1 $X=12.57
+ $Y=1.835 $X2=12.71 $Y2=2.1
r262 7 50 600 $w=1.7e-07 $l=1.08356e-06 $layer=licon1_PDIFF $count=1 $X=10.83
+ $Y=1.835 $X2=11.015 $Y2=2.83
r263 6 46 600 $w=1.7e-07 $l=3.30189e-07 $layer=licon1_PDIFF $count=1 $X=9.765
+ $Y=2.67 $X2=10.01 $Y2=2.87
r264 5 143 300 $w=1.7e-07 $l=6.71491e-07 $layer=licon1_PDIFF $count=2 $X=8.435
+ $Y=2.67 $X2=8.975 $Y2=2.965
r265 4 42 600 $w=1.7e-07 $l=9.05345e-07 $layer=licon1_PDIFF $count=1 $X=6.285
+ $Y=1.895 $X2=6.41 $Y2=2.74
r266 3 38 600 $w=1.7e-07 $l=3.78253e-07 $layer=licon1_PDIFF $count=1 $X=4.83
+ $Y=2.315 $X2=5.02 $Y2=2.61
r267 2 34 600 $w=1.7e-07 $l=5.21536e-07 $layer=licon1_PDIFF $count=1 $X=2.92
+ $Y=2.34 $X2=3.135 $Y2=2.765
r268 1 30 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=1.23
+ $Y=2.34 $X2=1.37 $Y2=2.485
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRTP_2%A_380_50# 1 2 3 4 15 17 20 23 26 31 32 34
+ 36
c99 34 0 1.50059e-19 $X=3.75 $Y=2.465
c100 23 0 1.50829e-19 $X=3.955 $Y=0.92
r101 36 38 5.09734 $w=2.58e-07 $l=1.15e-07 $layer=LI1_cond $X=4.085 $Y=0.805
+ $X2=4.085 $Y2=0.92
r102 26 28 7.68295 $w=3.28e-07 $l=2.2e-07 $layer=LI1_cond $X=2.155 $Y=0.7
+ $X2=2.155 $Y2=0.92
r103 24 32 6.47928 $w=1.7e-07 $l=1.13e-07 $layer=LI1_cond $X=3.68 $Y=0.92
+ $X2=3.567 $Y2=0.92
r104 23 38 3.22376 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.955 $Y=0.92
+ $X2=4.085 $Y2=0.92
r105 23 24 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=3.955 $Y=0.92
+ $X2=3.68 $Y2=0.92
r106 20 34 3.14896 $w=3e-07 $l=1.39155e-07 $layer=LI1_cond $X=3.567 $Y=2.3
+ $X2=3.67 $Y2=2.385
r107 19 32 0.355529 $w=2.25e-07 $l=8.5e-08 $layer=LI1_cond $X=3.567 $Y=1.005
+ $X2=3.567 $Y2=0.92
r108 19 20 66.3295 $w=2.23e-07 $l=1.295e-06 $layer=LI1_cond $X=3.567 $Y=1.005
+ $X2=3.567 $Y2=2.3
r109 18 31 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.325 $Y=2.385
+ $X2=2.16 $Y2=2.385
r110 17 34 3.44808 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=3.455 $Y=2.385
+ $X2=3.67 $Y2=2.385
r111 17 18 73.7219 $w=1.68e-07 $l=1.13e-06 $layer=LI1_cond $X=3.455 $Y=2.385
+ $X2=2.325 $Y2=2.385
r112 16 28 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.32 $Y=0.92
+ $X2=2.155 $Y2=0.92
r113 15 32 6.47928 $w=1.7e-07 $l=1.12e-07 $layer=LI1_cond $X=3.455 $Y=0.92
+ $X2=3.567 $Y2=0.92
r114 15 16 74.0481 $w=1.68e-07 $l=1.135e-06 $layer=LI1_cond $X=3.455 $Y=0.92
+ $X2=2.32 $Y2=0.92
r115 4 34 300 $w=1.7e-07 $l=3.00791e-07 $layer=licon1_PDIFF $count=2 $X=3.515
+ $Y=2.315 $X2=3.75 $Y2=2.465
r116 3 31 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=2.02
+ $Y=2.34 $X2=2.16 $Y2=2.465
r117 2 36 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=3.995
+ $Y=0.595 $X2=4.13 $Y2=0.805
r118 1 26 182 $w=1.7e-07 $l=5.6325e-07 $layer=licon1_NDIFF $count=1 $X=1.9
+ $Y=0.25 $X2=2.155 $Y2=0.7
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRTP_2%Q 1 2 9 13 14 15 16 17 18
r26 18 30 5.98384 $w=2.58e-07 $l=1.35e-07 $layer=LI1_cond $X=13.245 $Y=2.775
+ $X2=13.245 $Y2=2.91
r27 17 18 16.4002 $w=2.58e-07 $l=3.7e-07 $layer=LI1_cond $X=13.245 $Y=2.405
+ $X2=13.245 $Y2=2.775
r28 16 17 19.7245 $w=2.58e-07 $l=4.45e-07 $layer=LI1_cond $X=13.245 $Y=1.96
+ $X2=13.245 $Y2=2.405
r29 14 16 3.32435 $w=2.58e-07 $l=7.5e-08 $layer=LI1_cond $X=13.245 $Y=1.885
+ $X2=13.245 $Y2=1.96
r30 14 15 6.99888 $w=2.58e-07 $l=1.3e-07 $layer=LI1_cond $X=13.245 $Y=1.885
+ $X2=13.245 $Y2=1.755
r31 13 15 43.7299 $w=1.73e-07 $l=6.9e-07 $layer=LI1_cond $X=13.287 $Y=1.065
+ $X2=13.287 $Y2=1.755
r32 7 13 6.99888 $w=2.58e-07 $l=1.3e-07 $layer=LI1_cond $X=13.245 $Y=0.935
+ $X2=13.245 $Y2=1.065
r33 7 9 22.8272 $w=2.58e-07 $l=5.15e-07 $layer=LI1_cond $X=13.245 $Y=0.935
+ $X2=13.245 $Y2=0.42
r34 2 30 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=13.08
+ $Y=1.835 $X2=13.22 $Y2=2.91
r35 2 16 400 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=13.08
+ $Y=1.835 $X2=13.22 $Y2=1.96
r36 1 9 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=13.08
+ $Y=0.235 $X2=13.22 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRTP_2%VGND 1 2 3 4 5 6 7 24 28 32 36 40 44 46 48
+ 51 52 54 55 57 58 59 61 66 93 100 106 109 112 116
c143 116 0 3.56444e-20 $X=13.68 $Y=0
c144 28 0 1.55733e-19 $X=3.57 $Y=0.55
r145 115 116 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.68 $Y=0
+ $X2=13.68 $Y2=0
r146 112 113 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.72 $Y=0
+ $X2=12.72 $Y2=0
r147 109 110 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r148 106 107 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0
+ $X2=0.72 $Y2=0
r149 104 116 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.2 $Y=0
+ $X2=13.68 $Y2=0
r150 104 113 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.2 $Y=0
+ $X2=12.72 $Y2=0
r151 103 104 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.2 $Y=0
+ $X2=13.2 $Y2=0
r152 101 112 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.945 $Y=0
+ $X2=12.78 $Y2=0
r153 101 103 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=12.945 $Y=0
+ $X2=13.2 $Y2=0
r154 100 115 4.20444 $w=1.7e-07 $l=1.87e-07 $layer=LI1_cond $X=13.545 $Y=0
+ $X2=13.732 $Y2=0
r155 100 103 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=13.545 $Y=0
+ $X2=13.2 $Y2=0
r156 99 113 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.24 $Y=0
+ $X2=12.72 $Y2=0
r157 98 99 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=12.24 $Y=0
+ $X2=12.24 $Y2=0
r158 96 99 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=11.28 $Y=0
+ $X2=12.24 $Y2=0
r159 95 98 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=11.28 $Y=0 $X2=12.24
+ $Y2=0
r160 95 96 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=11.28 $Y=0
+ $X2=11.28 $Y2=0
r161 93 112 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.615 $Y=0
+ $X2=12.78 $Y2=0
r162 93 98 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=12.615 $Y=0
+ $X2=12.24 $Y2=0
r163 92 96 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.8 $Y=0
+ $X2=11.28 $Y2=0
r164 91 92 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=10.8 $Y=0
+ $X2=10.8 $Y2=0
r165 89 92 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=8.88 $Y=0
+ $X2=10.8 $Y2=0
r166 88 91 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=8.88 $Y=0 $X2=10.8
+ $Y2=0
r167 88 89 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=8.88 $Y=0
+ $X2=8.88 $Y2=0
r168 86 89 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=0 $X2=8.88
+ $Y2=0
r169 85 86 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r170 82 85 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=6.48 $Y=0 $X2=8.4
+ $Y2=0
r171 82 83 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.48 $Y=0
+ $X2=6.48 $Y2=0
r172 80 83 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.48
+ $Y2=0
r173 79 80 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6 $Y=0 $X2=6
+ $Y2=0
r174 77 80 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=4.08 $Y=0 $X2=6
+ $Y2=0
r175 77 110 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.6
+ $Y2=0
r176 76 79 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=4.08 $Y=0 $X2=6
+ $Y2=0
r177 76 77 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.08 $Y=0
+ $X2=4.08 $Y2=0
r178 74 109 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.735 $Y=0
+ $X2=3.57 $Y2=0
r179 74 76 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=3.735 $Y=0 $X2=4.08
+ $Y2=0
r180 73 110 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r181 72 73 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=0
+ $X2=3.12 $Y2=0
r182 70 73 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=1.2 $Y=0 $X2=3.12
+ $Y2=0
r183 70 107 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r184 69 72 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=3.12
+ $Y2=0
r185 69 70 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r186 67 106 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.895 $Y=0
+ $X2=0.73 $Y2=0
r187 67 69 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.895 $Y=0 $X2=1.2
+ $Y2=0
r188 66 109 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.405 $Y=0
+ $X2=3.57 $Y2=0
r189 66 72 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=3.405 $Y=0
+ $X2=3.12 $Y2=0
r190 64 107 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0
+ $X2=0.72 $Y2=0
r191 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r192 61 106 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.565 $Y=0
+ $X2=0.73 $Y2=0
r193 61 63 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.565 $Y=0
+ $X2=0.24 $Y2=0
r194 59 86 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=6.96 $Y=0 $X2=8.4
+ $Y2=0
r195 59 83 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=6.48
+ $Y2=0
r196 57 91 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=10.88 $Y=0 $X2=10.8
+ $Y2=0
r197 57 58 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.88 $Y=0
+ $X2=11.045 $Y2=0
r198 56 95 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=11.21 $Y=0 $X2=11.28
+ $Y2=0
r199 56 58 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.21 $Y=0
+ $X2=11.045 $Y2=0
r200 54 85 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=8.47 $Y=0 $X2=8.4
+ $Y2=0
r201 54 55 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.47 $Y=0 $X2=8.635
+ $Y2=0
r202 53 88 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=8.8 $Y=0 $X2=8.88
+ $Y2=0
r203 53 55 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.8 $Y=0 $X2=8.635
+ $Y2=0
r204 51 79 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=6.145 $Y=0 $X2=6
+ $Y2=0
r205 51 52 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.145 $Y=0 $X2=6.31
+ $Y2=0
r206 50 82 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=6.475 $Y=0 $X2=6.48
+ $Y2=0
r207 50 52 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.475 $Y=0 $X2=6.31
+ $Y2=0
r208 46 115 3.08026 $w=2.7e-07 $l=1.07912e-07 $layer=LI1_cond $X=13.68 $Y=0.085
+ $X2=13.732 $Y2=0
r209 46 48 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=13.68 $Y=0.085
+ $X2=13.68 $Y2=0.38
r210 42 112 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=12.78 $Y=0.085
+ $X2=12.78 $Y2=0
r211 42 44 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=12.78 $Y=0.085
+ $X2=12.78 $Y2=0.36
r212 38 58 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=11.045 $Y=0.085
+ $X2=11.045 $Y2=0
r213 38 40 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=11.045 $Y=0.085
+ $X2=11.045 $Y2=0.38
r214 34 55 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.635 $Y=0.085
+ $X2=8.635 $Y2=0
r215 34 36 24.6204 $w=3.28e-07 $l=7.05e-07 $layer=LI1_cond $X=8.635 $Y=0.085
+ $X2=8.635 $Y2=0.79
r216 30 52 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.31 $Y=0.085
+ $X2=6.31 $Y2=0
r217 30 32 14.8421 $w=3.28e-07 $l=4.25e-07 $layer=LI1_cond $X=6.31 $Y=0.085
+ $X2=6.31 $Y2=0.51
r218 26 109 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.57 $Y=0.085
+ $X2=3.57 $Y2=0
r219 26 28 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=3.57 $Y=0.085
+ $X2=3.57 $Y2=0.55
r220 22 106 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=0.085
+ $X2=0.73 $Y2=0
r221 22 24 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=0.73 $Y=0.085
+ $X2=0.73 $Y2=0.565
r222 7 48 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=13.51
+ $Y=0.235 $X2=13.65 $Y2=0.38
r223 6 44 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=12.57
+ $Y=0.235 $X2=12.78 $Y2=0.36
r224 5 40 182 $w=1.7e-07 $l=2.27376e-07 $layer=licon1_NDIFF $count=1 $X=10.825
+ $Y=0.365 $X2=11.045 $Y2=0.38
r225 4 36 182 $w=1.7e-07 $l=4.07247e-07 $layer=licon1_NDIFF $count=1 $X=8.325
+ $Y=0.565 $X2=8.635 $Y2=0.79
r226 3 32 182 $w=1.7e-07 $l=4.01559e-07 $layer=licon1_NDIFF $count=1 $X=5.935
+ $Y=0.565 $X2=6.31 $Y2=0.51
r227 2 28 182 $w=1.7e-07 $l=2.67862e-07 $layer=licon1_NDIFF $count=1 $X=3.365
+ $Y=0.405 $X2=3.57 $Y2=0.55
r228 1 24 182 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_NDIFF $count=1 $X=0.59
+ $Y=0.37 $X2=0.73 $Y2=0.565
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRTP_2%noxref_24 1 2 7 9 14
c32 7 0 2.67853e-19 $X=2.895 $Y=0.35
r33 14 17 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=3.06 $Y=0.35 $X2=3.06
+ $Y2=0.55
r34 9 12 3.84148 $w=3.28e-07 $l=1.1e-07 $layer=LI1_cond $X=1.25 $Y=0.35 $X2=1.25
+ $Y2=0.46
r35 8 9 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.415 $Y=0.35 $X2=1.25
+ $Y2=0.35
r36 7 14 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.895 $Y=0.35
+ $X2=3.06 $Y2=0.35
r37 7 8 96.5562 $w=1.68e-07 $l=1.48e-06 $layer=LI1_cond $X=2.895 $Y=0.35
+ $X2=1.415 $Y2=0.35
r38 2 17 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=2.92
+ $Y=0.405 $X2=3.06 $Y2=0.55
r39 1 12 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=1.125
+ $Y=0.25 $X2=1.25 $Y2=0.46
.ends

