# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_sc_lp__and4bb_m
  CLASS CORE ;
  FOREIGN sky130_fd_sc_lp__and4bb_m ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.320000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.475000 0.805000 0.805000 1.475000 ;
    END
  END A_N
  PIN B_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.045000 0.805000 1.285000 1.475000 ;
    END
  END B_N
  PIN C
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.075000 1.210000 2.975000 1.405000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.005000 1.950000 3.335000 2.120000 ;
    END
  END D
  PIN X
    ANTENNADIFFAREA  0.222600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.730000 2.655000 4.165000 2.985000 ;
        RECT 3.975000 0.470000 4.165000 2.655000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.320000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.000000 0.000000 4.320000 0.245000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.655000 4.510000 3.520000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.320000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.320000 0.085000 ;
      RECT 0.000000  3.245000 4.320000 3.415000 ;
      RECT 0.125000  0.295000 0.500000 0.625000 ;
      RECT 0.125000  0.625000 0.295000 1.655000 ;
      RECT 0.125000  1.655000 1.785000 1.825000 ;
      RECT 0.125000  1.825000 0.500000 2.295000 ;
      RECT 0.720000  0.085000 0.930000 0.585000 ;
      RECT 0.720000  2.095000 0.930000 3.245000 ;
      RECT 1.150000  0.265000 2.615000 0.435000 ;
      RECT 1.150000  0.435000 1.360000 0.595000 ;
      RECT 1.150000  2.005000 2.435000 2.175000 ;
      RECT 1.150000  2.175000 1.360000 2.335000 ;
      RECT 1.540000  2.785000 1.750000 3.245000 ;
      RECT 1.615000  1.155000 1.785000 1.655000 ;
      RECT 1.680000  0.645000 3.325000 0.975000 ;
      RECT 1.970000  2.435000 3.040000 2.605000 ;
      RECT 1.970000  2.605000 2.180000 2.985000 ;
      RECT 2.105000  1.615000 2.435000 2.005000 ;
      RECT 2.400000  2.785000 2.610000 3.245000 ;
      RECT 2.655000  1.585000 3.795000 1.755000 ;
      RECT 2.655000  1.755000 2.825000 2.435000 ;
      RECT 2.830000  2.605000 3.040000 2.985000 ;
      RECT 3.155000  0.975000 3.325000 1.585000 ;
      RECT 3.220000  2.845000 3.550000 3.245000 ;
      RECT 3.505000  0.085000 3.715000 0.935000 ;
      RECT 3.625000  1.755000 3.795000 2.255000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
  END
END sky130_fd_sc_lp__and4bb_m
END LIBRARY
