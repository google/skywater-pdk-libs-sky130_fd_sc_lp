* File: sky130_fd_sc_lp__or2b_2.pxi.spice
* Created: Fri Aug 28 11:22:21 2020
* 
x_PM_SKY130_FD_SC_LP__OR2B_2%B_N N_B_N_M1001_g N_B_N_M1005_g N_B_N_c_57_n
+ N_B_N_c_58_n B_N N_B_N_c_59_n N_B_N_c_60_n PM_SKY130_FD_SC_LP__OR2B_2%B_N
x_PM_SKY130_FD_SC_LP__OR2B_2%A_191_254# N_A_191_254#_M1004_d
+ N_A_191_254#_M1007_d N_A_191_254#_M1002_g N_A_191_254#_c_83_n
+ N_A_191_254#_M1000_g N_A_191_254#_M1008_g N_A_191_254#_c_85_n
+ N_A_191_254#_M1003_g N_A_191_254#_c_86_n N_A_191_254#_c_87_n
+ N_A_191_254#_c_88_n N_A_191_254#_c_106_p N_A_191_254#_c_136_p
+ N_A_191_254#_c_93_n N_A_191_254#_c_89_n PM_SKY130_FD_SC_LP__OR2B_2%A_191_254#
x_PM_SKY130_FD_SC_LP__OR2B_2%A N_A_M1004_g N_A_M1006_g A A N_A_c_165_n
+ PM_SKY130_FD_SC_LP__OR2B_2%A
x_PM_SKY130_FD_SC_LP__OR2B_2%A_27_49# N_A_27_49#_M1001_s N_A_27_49#_M1005_s
+ N_A_27_49#_c_200_n N_A_27_49#_M1009_g N_A_27_49#_M1007_g N_A_27_49#_c_202_n
+ N_A_27_49#_c_203_n N_A_27_49#_c_204_n N_A_27_49#_c_205_n N_A_27_49#_c_234_n
+ N_A_27_49#_c_206_n N_A_27_49#_c_211_n N_A_27_49#_c_260_p N_A_27_49#_c_207_n
+ N_A_27_49#_c_208_n PM_SKY130_FD_SC_LP__OR2B_2%A_27_49#
x_PM_SKY130_FD_SC_LP__OR2B_2%VPWR N_VPWR_M1005_d N_VPWR_M1008_d N_VPWR_c_284_n
+ N_VPWR_c_285_n VPWR N_VPWR_c_286_n N_VPWR_c_287_n N_VPWR_c_283_n
+ N_VPWR_c_289_n N_VPWR_c_290_n PM_SKY130_FD_SC_LP__OR2B_2%VPWR
x_PM_SKY130_FD_SC_LP__OR2B_2%X N_X_M1000_d N_X_M1002_s N_X_c_311_n X X X X X
+ PM_SKY130_FD_SC_LP__OR2B_2%X
x_PM_SKY130_FD_SC_LP__OR2B_2%VGND N_VGND_M1001_d N_VGND_M1003_s N_VGND_M1009_d
+ N_VGND_c_329_n N_VGND_c_330_n VGND N_VGND_c_331_n N_VGND_c_332_n
+ N_VGND_c_333_n N_VGND_c_334_n N_VGND_c_335_n N_VGND_c_336_n
+ PM_SKY130_FD_SC_LP__OR2B_2%VGND
cc_1 VNB N_B_N_M1001_g 0.0314471f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.455
cc_2 VNB N_B_N_M1005_g 0.00914145f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=2.045
cc_3 VNB N_B_N_c_57_n 0.0309647f $X=-0.19 $Y=-0.245 $X2=0.417 $Y2=1.395
cc_4 VNB N_B_N_c_58_n 0.0237317f $X=-0.19 $Y=-0.245 $X2=0.417 $Y2=1.545
cc_5 VNB N_B_N_c_59_n 0.0192047f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.04
cc_6 VNB N_B_N_c_60_n 0.030631f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.04
cc_7 VNB N_A_191_254#_M1002_g 0.00646903f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.04
cc_8 VNB N_A_191_254#_c_83_n 0.0172093f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.395
cc_9 VNB N_A_191_254#_M1008_g 0.00713075f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.04
cc_10 VNB N_A_191_254#_c_85_n 0.0196644f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.04
cc_11 VNB N_A_191_254#_c_86_n 0.00156678f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_191_254#_c_87_n 0.0027935f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_191_254#_c_88_n 0.010005f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_191_254#_c_89_n 0.0674824f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_M1004_g 0.0261156f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.455
cc_16 VNB A 0.0122514f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=0.875
cc_17 VNB N_A_c_165_n 0.0244758f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_18 VNB N_A_27_49#_c_200_n 0.0195433f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=2.045
cc_19 VNB N_A_27_49#_M1007_g 0.0070637f $X=-0.19 $Y=-0.245 $X2=0.417 $Y2=1.395
cc_20 VNB N_A_27_49#_c_202_n 0.0112022f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_27_49#_c_203_n 0.003401f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.04
cc_22 VNB N_A_27_49#_c_204_n 0.013487f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.21
cc_23 VNB N_A_27_49#_c_205_n 0.0116788f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_27_49#_c_206_n 0.0183396f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_27_49#_c_207_n 0.0532278f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_27_49#_c_208_n 0.0904527f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_VPWR_c_283_n 0.163682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB X 6.5803e-19 $X=-0.19 $Y=-0.245 $X2=0.417 $Y2=1.395
cc_29 VNB N_VGND_c_329_n 0.0181447f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=0.875
cc_30 VNB N_VGND_c_330_n 0.0476757f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_31 VNB N_VGND_c_331_n 0.0286702f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.04
cc_32 VNB N_VGND_c_332_n 0.0291746f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_333_n 0.0174178f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_334_n 0.240078f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_335_n 0.0155415f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_336_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VPB N_B_N_M1005_g 0.0313917f $X=-0.19 $Y=1.655 $X2=0.54 $Y2=2.045
cc_38 VPB N_A_191_254#_M1002_g 0.0223201f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.04
cc_39 VPB N_A_191_254#_M1008_g 0.0237899f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.04
cc_40 VPB N_A_191_254#_c_86_n 0.00384419f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_41 VPB N_A_191_254#_c_93_n 0.0244957f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_42 VPB N_A_M1006_g 0.0254752f $X=-0.19 $Y=1.655 $X2=0.54 $Y2=2.045
cc_43 VPB A 0.0094008f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=0.875
cc_44 VPB N_A_c_165_n 0.0064595f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_45 VPB N_A_27_49#_M1007_g 0.0300978f $X=-0.19 $Y=1.655 $X2=0.417 $Y2=1.395
cc_46 VPB N_A_27_49#_c_204_n 9.86942e-19 $X=-0.19 $Y=1.655 $X2=0.24 $Y2=1.21
cc_47 VPB N_A_27_49#_c_211_n 0.0248004f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_48 VPB N_VPWR_c_284_n 0.0308435f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.395
cc_49 VPB N_VPWR_c_285_n 0.0331033f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.04
cc_50 VPB N_VPWR_c_286_n 0.017949f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_51 VPB N_VPWR_c_287_n 0.0657873f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_52 VPB N_VPWR_c_283_n 0.147377f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_53 VPB N_VPWR_c_289_n 0.02824f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_54 VPB N_VPWR_c_290_n 0.00497181f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_55 N_B_N_M1005_g N_A_191_254#_M1002_g 0.0119185f $X=0.54 $Y=2.045 $X2=0 $Y2=0
cc_56 N_B_N_M1001_g N_A_191_254#_c_83_n 0.0128996f $X=0.475 $Y=0.455 $X2=0 $Y2=0
cc_57 N_B_N_c_57_n N_A_191_254#_c_89_n 0.00305605f $X=0.417 $Y=1.395 $X2=0 $Y2=0
cc_58 N_B_N_c_58_n N_A_191_254#_c_89_n 0.0119185f $X=0.417 $Y=1.545 $X2=0 $Y2=0
cc_59 N_B_N_c_59_n N_A_191_254#_c_89_n 0.0128996f $X=0.385 $Y=1.04 $X2=0 $Y2=0
cc_60 N_B_N_M1001_g N_A_27_49#_c_203_n 0.0120676f $X=0.475 $Y=0.455 $X2=0 $Y2=0
cc_61 N_B_N_c_60_n N_A_27_49#_c_203_n 0.00361551f $X=0.385 $Y=1.04 $X2=0 $Y2=0
cc_62 N_B_N_M1001_g N_A_27_49#_c_204_n 0.0092083f $X=0.475 $Y=0.455 $X2=0 $Y2=0
cc_63 N_B_N_c_58_n N_A_27_49#_c_204_n 0.00571753f $X=0.417 $Y=1.545 $X2=0 $Y2=0
cc_64 N_B_N_c_60_n N_A_27_49#_c_204_n 0.0488038f $X=0.385 $Y=1.04 $X2=0 $Y2=0
cc_65 N_B_N_M1001_g N_A_27_49#_c_206_n 0.00628757f $X=0.475 $Y=0.455 $X2=0 $Y2=0
cc_66 N_B_N_c_59_n N_A_27_49#_c_206_n 0.00473499f $X=0.385 $Y=1.04 $X2=0 $Y2=0
cc_67 N_B_N_c_60_n N_A_27_49#_c_206_n 0.0268247f $X=0.385 $Y=1.04 $X2=0 $Y2=0
cc_68 N_B_N_M1005_g N_A_27_49#_c_211_n 0.024323f $X=0.54 $Y=2.045 $X2=0 $Y2=0
cc_69 N_B_N_c_58_n N_A_27_49#_c_211_n 0.00654169f $X=0.417 $Y=1.545 $X2=0 $Y2=0
cc_70 N_B_N_c_60_n N_A_27_49#_c_211_n 0.0270559f $X=0.385 $Y=1.04 $X2=0 $Y2=0
cc_71 N_B_N_M1005_g N_VPWR_c_284_n 0.00570632f $X=0.54 $Y=2.045 $X2=0 $Y2=0
cc_72 N_B_N_M1005_g X 7.39028e-19 $X=0.54 $Y=2.045 $X2=0 $Y2=0
cc_73 N_B_N_M1001_g N_VGND_c_331_n 0.00780554f $X=0.475 $Y=0.455 $X2=0 $Y2=0
cc_74 N_B_N_M1001_g N_VGND_c_334_n 0.00674166f $X=0.475 $Y=0.455 $X2=0 $Y2=0
cc_75 N_A_191_254#_c_85_n N_A_M1004_g 0.0137786f $X=1.495 $Y=1.195 $X2=0 $Y2=0
cc_76 N_A_191_254#_c_86_n N_A_M1004_g 9.17641e-19 $X=1.665 $Y=1.36 $X2=0 $Y2=0
cc_77 N_A_191_254#_c_87_n N_A_M1004_g 0.0021183f $X=1.83 $Y=0.995 $X2=0 $Y2=0
cc_78 N_A_191_254#_c_88_n N_A_M1004_g 0.0132149f $X=2.355 $Y=0.96 $X2=0 $Y2=0
cc_79 N_A_191_254#_c_89_n N_A_M1004_g 0.019202f $X=1.495 $Y=1.36 $X2=0 $Y2=0
cc_80 N_A_191_254#_M1008_g N_A_M1006_g 0.00760725f $X=1.46 $Y=2.465 $X2=0 $Y2=0
cc_81 N_A_191_254#_c_86_n N_A_M1006_g 0.00350347f $X=1.665 $Y=1.36 $X2=0 $Y2=0
cc_82 N_A_191_254#_c_106_p N_A_M1006_g 0.0153676f $X=2.73 $Y=2.015 $X2=0 $Y2=0
cc_83 N_A_191_254#_c_93_n N_A_M1006_g 8.79113e-19 $X=2.895 $Y=2.015 $X2=0 $Y2=0
cc_84 N_A_191_254#_c_86_n A 0.0293164f $X=1.665 $Y=1.36 $X2=0 $Y2=0
cc_85 N_A_191_254#_c_88_n A 0.0274247f $X=2.355 $Y=0.96 $X2=0 $Y2=0
cc_86 N_A_191_254#_c_106_p A 0.0490945f $X=2.73 $Y=2.015 $X2=0 $Y2=0
cc_87 N_A_191_254#_c_93_n A 0.00262073f $X=2.895 $Y=2.015 $X2=0 $Y2=0
cc_88 N_A_191_254#_c_89_n A 7.77521e-19 $X=1.495 $Y=1.36 $X2=0 $Y2=0
cc_89 N_A_191_254#_M1008_g N_A_c_165_n 0.00227616f $X=1.46 $Y=2.465 $X2=0 $Y2=0
cc_90 N_A_191_254#_c_86_n N_A_c_165_n 6.30719e-19 $X=1.665 $Y=1.36 $X2=0 $Y2=0
cc_91 N_A_191_254#_c_88_n N_A_c_165_n 0.00465154f $X=2.355 $Y=0.96 $X2=0 $Y2=0
cc_92 N_A_191_254#_c_106_p N_A_c_165_n 8.99471e-19 $X=2.73 $Y=2.015 $X2=0 $Y2=0
cc_93 N_A_191_254#_c_88_n N_A_27_49#_c_200_n 0.00229625f $X=2.355 $Y=0.96 $X2=0
+ $Y2=0
cc_94 N_A_191_254#_c_106_p N_A_27_49#_M1007_g 0.01071f $X=2.73 $Y=2.015 $X2=0
+ $Y2=0
cc_95 N_A_191_254#_c_93_n N_A_27_49#_M1007_g 0.0049628f $X=2.895 $Y=2.015 $X2=0
+ $Y2=0
cc_96 N_A_191_254#_c_83_n N_A_27_49#_c_204_n 0.00723473f $X=1.065 $Y=1.195 $X2=0
+ $Y2=0
cc_97 N_A_191_254#_c_89_n N_A_27_49#_c_204_n 0.0040092f $X=1.495 $Y=1.36 $X2=0
+ $Y2=0
cc_98 N_A_191_254#_M1004_d N_A_27_49#_c_205_n 0.00366138f $X=2.215 $Y=0.665
+ $X2=0 $Y2=0
cc_99 N_A_191_254#_c_83_n N_A_27_49#_c_205_n 0.0148329f $X=1.065 $Y=1.195 $X2=0
+ $Y2=0
cc_100 N_A_191_254#_c_85_n N_A_27_49#_c_205_n 0.0161627f $X=1.495 $Y=1.195 $X2=0
+ $Y2=0
cc_101 N_A_191_254#_c_87_n N_A_27_49#_c_205_n 0.0161097f $X=1.83 $Y=0.995 $X2=0
+ $Y2=0
cc_102 N_A_191_254#_c_88_n N_A_27_49#_c_205_n 0.0423932f $X=2.355 $Y=0.96 $X2=0
+ $Y2=0
cc_103 N_A_191_254#_c_89_n N_A_27_49#_c_205_n 0.00115549f $X=1.495 $Y=1.36 $X2=0
+ $Y2=0
cc_104 N_A_191_254#_c_88_n N_A_27_49#_c_234_n 0.0164623f $X=2.355 $Y=0.96 $X2=0
+ $Y2=0
cc_105 N_A_191_254#_c_83_n N_A_27_49#_c_206_n 8.54725e-19 $X=1.065 $Y=1.195
+ $X2=0 $Y2=0
cc_106 N_A_191_254#_M1002_g N_A_27_49#_c_211_n 0.00201891f $X=1.03 $Y=2.465
+ $X2=0 $Y2=0
cc_107 N_A_191_254#_c_88_n N_A_27_49#_c_207_n 0.00435067f $X=2.355 $Y=0.96 $X2=0
+ $Y2=0
cc_108 N_A_191_254#_c_93_n N_A_27_49#_c_207_n 0.00472759f $X=2.895 $Y=2.015
+ $X2=0 $Y2=0
cc_109 N_A_191_254#_c_93_n N_A_27_49#_c_208_n 0.00550552f $X=2.895 $Y=2.015
+ $X2=0 $Y2=0
cc_110 N_A_191_254#_c_86_n N_VPWR_M1008_d 0.00263887f $X=1.665 $Y=1.36 $X2=0
+ $Y2=0
cc_111 N_A_191_254#_c_106_p N_VPWR_M1008_d 0.0237807f $X=2.73 $Y=2.015 $X2=0
+ $Y2=0
cc_112 N_A_191_254#_c_136_p N_VPWR_M1008_d 0.00486217f $X=1.83 $Y=2.015 $X2=0
+ $Y2=0
cc_113 N_A_191_254#_M1002_g N_VPWR_c_284_n 0.00325151f $X=1.03 $Y=2.465 $X2=0
+ $Y2=0
cc_114 N_A_191_254#_M1008_g N_VPWR_c_285_n 0.00569178f $X=1.46 $Y=2.465 $X2=0
+ $Y2=0
cc_115 N_A_191_254#_c_106_p N_VPWR_c_285_n 7.11687e-19 $X=2.73 $Y=2.015 $X2=0
+ $Y2=0
cc_116 N_A_191_254#_c_136_p N_VPWR_c_285_n 0.0214665f $X=1.83 $Y=2.015 $X2=0
+ $Y2=0
cc_117 N_A_191_254#_M1002_g N_VPWR_c_286_n 0.0054895f $X=1.03 $Y=2.465 $X2=0
+ $Y2=0
cc_118 N_A_191_254#_M1008_g N_VPWR_c_286_n 0.0054895f $X=1.46 $Y=2.465 $X2=0
+ $Y2=0
cc_119 N_A_191_254#_M1002_g N_VPWR_c_283_n 0.0110654f $X=1.03 $Y=2.465 $X2=0
+ $Y2=0
cc_120 N_A_191_254#_M1008_g N_VPWR_c_283_n 0.0110654f $X=1.46 $Y=2.465 $X2=0
+ $Y2=0
cc_121 N_A_191_254#_c_83_n N_X_c_311_n 0.00351196f $X=1.065 $Y=1.195 $X2=0 $Y2=0
cc_122 N_A_191_254#_c_85_n N_X_c_311_n 0.00319821f $X=1.495 $Y=1.195 $X2=0 $Y2=0
cc_123 N_A_191_254#_M1002_g X 0.024262f $X=1.03 $Y=2.465 $X2=0 $Y2=0
cc_124 N_A_191_254#_c_83_n X 0.00327589f $X=1.065 $Y=1.195 $X2=0 $Y2=0
cc_125 N_A_191_254#_M1008_g X 0.0279715f $X=1.46 $Y=2.465 $X2=0 $Y2=0
cc_126 N_A_191_254#_c_85_n X 9.36079e-19 $X=1.495 $Y=1.195 $X2=0 $Y2=0
cc_127 N_A_191_254#_c_86_n X 0.0454529f $X=1.665 $Y=1.36 $X2=0 $Y2=0
cc_128 N_A_191_254#_c_87_n X 0.0147029f $X=1.83 $Y=0.995 $X2=0 $Y2=0
cc_129 N_A_191_254#_c_89_n X 0.0225585f $X=1.495 $Y=1.36 $X2=0 $Y2=0
cc_130 N_A_191_254#_c_106_p A_479_367# 0.00468592f $X=2.73 $Y=2.015 $X2=-0.19
+ $Y2=-0.245
cc_131 N_A_191_254#_c_87_n N_VGND_M1003_s 0.00384935f $X=1.83 $Y=0.995 $X2=0
+ $Y2=0
cc_132 N_A_191_254#_c_88_n N_VGND_M1003_s 0.00235634f $X=2.355 $Y=0.96 $X2=0
+ $Y2=0
cc_133 N_A_191_254#_c_83_n N_VGND_c_329_n 0.00400062f $X=1.065 $Y=1.195 $X2=0
+ $Y2=0
cc_134 N_A_191_254#_c_85_n N_VGND_c_329_n 0.00400062f $X=1.495 $Y=1.195 $X2=0
+ $Y2=0
cc_135 N_A_191_254#_c_83_n N_VGND_c_331_n 0.00373415f $X=1.065 $Y=1.195 $X2=0
+ $Y2=0
cc_136 N_A_191_254#_c_83_n N_VGND_c_334_n 0.00590457f $X=1.065 $Y=1.195 $X2=0
+ $Y2=0
cc_137 N_A_191_254#_c_85_n N_VGND_c_334_n 0.00684172f $X=1.495 $Y=1.195 $X2=0
+ $Y2=0
cc_138 N_A_191_254#_c_85_n N_VGND_c_335_n 0.00659856f $X=1.495 $Y=1.195 $X2=0
+ $Y2=0
cc_139 N_A_M1004_g N_A_27_49#_c_200_n 0.0204625f $X=2.14 $Y=0.875 $X2=0 $Y2=0
cc_140 N_A_M1006_g N_A_27_49#_M1007_g 0.0338974f $X=2.32 $Y=2.045 $X2=0 $Y2=0
cc_141 A N_A_27_49#_M1007_g 0.0108016f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_142 A N_A_27_49#_c_202_n 0.00753481f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_143 N_A_c_165_n N_A_27_49#_c_202_n 0.0338974f $X=2.23 $Y=1.51 $X2=0 $Y2=0
cc_144 N_A_M1004_g N_A_27_49#_c_205_n 0.0115624f $X=2.14 $Y=0.875 $X2=0 $Y2=0
cc_145 N_A_M1004_g N_A_27_49#_c_234_n 5.92513e-19 $X=2.14 $Y=0.875 $X2=0 $Y2=0
cc_146 N_A_M1004_g N_A_27_49#_c_207_n 6.24844e-19 $X=2.14 $Y=0.875 $X2=0 $Y2=0
cc_147 A N_A_27_49#_c_207_n 0.015995f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_148 N_A_c_165_n N_A_27_49#_c_207_n 3.02661e-19 $X=2.23 $Y=1.51 $X2=0 $Y2=0
cc_149 A N_A_27_49#_c_208_n 0.00239908f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_150 N_A_M1006_g N_VPWR_c_285_n 0.00226799f $X=2.32 $Y=2.045 $X2=0 $Y2=0
cc_151 N_A_M1004_g N_VGND_c_332_n 6.65218e-19 $X=2.14 $Y=0.875 $X2=0 $Y2=0
cc_152 N_A_27_49#_c_211_n N_VPWR_M1005_d 0.00269442f $X=0.325 $Y=2.045 $X2=-0.19
+ $Y2=-0.245
cc_153 N_A_27_49#_c_211_n N_VPWR_c_284_n 0.022641f $X=0.325 $Y=2.045 $X2=0 $Y2=0
cc_154 N_A_27_49#_c_205_n N_X_M1000_d 0.00415657f $X=2.69 $Y=0.61 $X2=-0.19
+ $Y2=-0.245
cc_155 N_A_27_49#_c_204_n N_X_c_311_n 0.0461456f $X=0.735 $Y=1.715 $X2=0 $Y2=0
cc_156 N_A_27_49#_c_205_n N_X_c_311_n 0.0190902f $X=2.69 $Y=0.61 $X2=0 $Y2=0
cc_157 N_A_27_49#_c_211_n X 0.0148947f $X=0.325 $Y=2.045 $X2=0 $Y2=0
cc_158 N_A_27_49#_c_203_n N_VGND_M1001_d 4.18348e-19 $X=0.65 $Y=0.61 $X2=-0.19
+ $Y2=-0.245
cc_159 N_A_27_49#_c_204_n N_VGND_M1001_d 0.00678716f $X=0.735 $Y=1.715 $X2=-0.19
+ $Y2=-0.245
cc_160 N_A_27_49#_c_205_n N_VGND_M1001_d 0.00538902f $X=2.69 $Y=0.61 $X2=-0.19
+ $Y2=-0.245
cc_161 N_A_27_49#_c_260_p N_VGND_M1001_d 0.00251533f $X=0.735 $Y=0.61 $X2=-0.19
+ $Y2=-0.245
cc_162 N_A_27_49#_c_205_n N_VGND_M1003_s 0.00813814f $X=2.69 $Y=0.61 $X2=0 $Y2=0
cc_163 N_A_27_49#_c_205_n N_VGND_M1009_d 3.32804e-19 $X=2.69 $Y=0.61 $X2=0 $Y2=0
cc_164 N_A_27_49#_c_234_n N_VGND_M1009_d 0.00867541f $X=2.775 $Y=1.075 $X2=0
+ $Y2=0
cc_165 N_A_27_49#_c_207_n N_VGND_M1009_d 0.0100983f $X=3.03 $Y=1.36 $X2=0 $Y2=0
cc_166 N_A_27_49#_c_205_n N_VGND_c_329_n 0.0131559f $X=2.69 $Y=0.61 $X2=0 $Y2=0
cc_167 N_A_27_49#_c_200_n N_VGND_c_330_n 0.00214003f $X=2.68 $Y=1.195 $X2=0
+ $Y2=0
cc_168 N_A_27_49#_c_205_n N_VGND_c_330_n 0.0149385f $X=2.69 $Y=0.61 $X2=0 $Y2=0
cc_169 N_A_27_49#_c_234_n N_VGND_c_330_n 0.0160122f $X=2.775 $Y=1.075 $X2=0
+ $Y2=0
cc_170 N_A_27_49#_c_207_n N_VGND_c_330_n 0.0288267f $X=3.03 $Y=1.36 $X2=0 $Y2=0
cc_171 N_A_27_49#_c_208_n N_VGND_c_330_n 0.00192991f $X=3.47 $Y=1.36 $X2=0 $Y2=0
cc_172 N_A_27_49#_c_203_n N_VGND_c_331_n 0.00643851f $X=0.65 $Y=0.61 $X2=0 $Y2=0
cc_173 N_A_27_49#_c_205_n N_VGND_c_331_n 0.00825314f $X=2.69 $Y=0.61 $X2=0 $Y2=0
cc_174 N_A_27_49#_c_206_n N_VGND_c_331_n 0.0163719f $X=0.26 $Y=0.455 $X2=0 $Y2=0
cc_175 N_A_27_49#_c_260_p N_VGND_c_331_n 0.013757f $X=0.735 $Y=0.61 $X2=0 $Y2=0
cc_176 N_A_27_49#_c_200_n N_VGND_c_332_n 6.80511e-19 $X=2.68 $Y=1.195 $X2=0
+ $Y2=0
cc_177 N_A_27_49#_c_205_n N_VGND_c_332_n 0.021679f $X=2.69 $Y=0.61 $X2=0 $Y2=0
cc_178 N_A_27_49#_M1001_s N_VGND_c_334_n 0.00214692f $X=0.135 $Y=0.245 $X2=0
+ $Y2=0
cc_179 N_A_27_49#_c_203_n N_VGND_c_334_n 0.00496331f $X=0.65 $Y=0.61 $X2=0 $Y2=0
cc_180 N_A_27_49#_c_205_n N_VGND_c_334_n 0.0509261f $X=2.69 $Y=0.61 $X2=0 $Y2=0
cc_181 N_A_27_49#_c_206_n N_VGND_c_334_n 0.0120621f $X=0.26 $Y=0.455 $X2=0 $Y2=0
cc_182 N_A_27_49#_c_260_p N_VGND_c_334_n 0.00107416f $X=0.735 $Y=0.61 $X2=0
+ $Y2=0
cc_183 N_A_27_49#_c_205_n N_VGND_c_335_n 0.0240258f $X=2.69 $Y=0.61 $X2=0 $Y2=0
cc_184 N_VPWR_c_283_n N_X_M1002_s 0.00223559f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_185 N_VPWR_c_286_n X 0.0189236f $X=1.58 $Y=3.33 $X2=0 $Y2=0
cc_186 N_VPWR_c_283_n X 0.0123859f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_187 N_X_M1000_d N_VGND_c_334_n 0.00283464f $X=1.14 $Y=0.245 $X2=0 $Y2=0
