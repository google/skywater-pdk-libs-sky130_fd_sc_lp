* File: sky130_fd_sc_lp__a2bb2o_1.pxi.spice
* Created: Fri Aug 28 09:55:45 2020
* 
x_PM_SKY130_FD_SC_LP__A2BB2O_1%A_91_269# N_A_91_269#_M1008_d N_A_91_269#_M1010_s
+ N_A_91_269#_M1011_g N_A_91_269#_M1009_g N_A_91_269#_c_92_n N_A_91_269#_c_99_n
+ N_A_91_269#_c_165_p N_A_91_269#_c_100_n N_A_91_269#_c_101_n
+ N_A_91_269#_c_102_n N_A_91_269#_c_93_n N_A_91_269#_c_94_n N_A_91_269#_c_95_n
+ N_A_91_269#_c_96_n PM_SKY130_FD_SC_LP__A2BB2O_1%A_91_269#
x_PM_SKY130_FD_SC_LP__A2BB2O_1%A1_N N_A1_N_c_187_n N_A1_N_M1005_g N_A1_N_M1000_g
+ N_A1_N_c_189_n A1_N A1_N A1_N A1_N A1_N N_A1_N_c_191_n
+ PM_SKY130_FD_SC_LP__A2BB2O_1%A1_N
x_PM_SKY130_FD_SC_LP__A2BB2O_1%A2_N N_A2_N_M1007_g N_A2_N_M1006_g N_A2_N_c_237_n
+ N_A2_N_c_238_n A2_N N_A2_N_c_239_n N_A2_N_c_240_n
+ PM_SKY130_FD_SC_LP__A2BB2O_1%A2_N
x_PM_SKY130_FD_SC_LP__A2BB2O_1%A_271_47# N_A_271_47#_M1005_d N_A_271_47#_M1007_d
+ N_A_271_47#_M1008_g N_A_271_47#_M1010_g N_A_271_47#_c_285_n
+ N_A_271_47#_c_286_n N_A_271_47#_c_295_n N_A_271_47#_c_296_n
+ N_A_271_47#_c_318_n N_A_271_47#_c_287_n N_A_271_47#_c_288_n
+ N_A_271_47#_c_289_n N_A_271_47#_c_290_n N_A_271_47#_c_291_n
+ N_A_271_47#_c_298_n N_A_271_47#_c_292_n PM_SKY130_FD_SC_LP__A2BB2O_1%A_271_47#
x_PM_SKY130_FD_SC_LP__A2BB2O_1%B2 N_B2_M1002_g N_B2_M1004_g B2 B2 B2 B2 B2
+ N_B2_c_376_n PM_SKY130_FD_SC_LP__A2BB2O_1%B2
x_PM_SKY130_FD_SC_LP__A2BB2O_1%B1 N_B1_M1003_g N_B1_M1001_g N_B1_c_424_n
+ N_B1_c_425_n N_B1_c_426_n N_B1_c_432_n N_B1_c_427_n B1 B1 B1 B1 N_B1_c_429_n
+ PM_SKY130_FD_SC_LP__A2BB2O_1%B1
x_PM_SKY130_FD_SC_LP__A2BB2O_1%X N_X_M1011_s N_X_M1009_s N_X_c_466_n N_X_c_467_n
+ N_X_c_463_n X X N_X_c_464_n X PM_SKY130_FD_SC_LP__A2BB2O_1%X
x_PM_SKY130_FD_SC_LP__A2BB2O_1%VPWR N_VPWR_M1009_d N_VPWR_M1004_d N_VPWR_c_489_n
+ N_VPWR_c_490_n N_VPWR_c_491_n N_VPWR_c_492_n VPWR N_VPWR_c_493_n
+ N_VPWR_c_494_n N_VPWR_c_488_n N_VPWR_c_496_n PM_SKY130_FD_SC_LP__A2BB2O_1%VPWR
x_PM_SKY130_FD_SC_LP__A2BB2O_1%A_505_529# N_A_505_529#_M1010_d
+ N_A_505_529#_M1001_d N_A_505_529#_c_528_n N_A_505_529#_c_529_n
+ N_A_505_529#_c_530_n N_A_505_529#_c_531_n
+ PM_SKY130_FD_SC_LP__A2BB2O_1%A_505_529#
x_PM_SKY130_FD_SC_LP__A2BB2O_1%VGND N_VGND_M1011_d N_VGND_M1006_d N_VGND_M1003_d
+ N_VGND_c_553_n N_VGND_c_554_n N_VGND_c_555_n N_VGND_c_556_n VGND
+ N_VGND_c_557_n N_VGND_c_558_n N_VGND_c_559_n N_VGND_c_560_n N_VGND_c_561_n
+ PM_SKY130_FD_SC_LP__A2BB2O_1%VGND
cc_1 VNB N_A_91_269#_M1011_g 0.0319838f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=0.655
cc_2 VNB N_A_91_269#_c_92_n 4.56378e-19 $X=-0.19 $Y=-0.245 $X2=0.84 $Y2=2.325
cc_3 VNB N_A_91_269#_c_93_n 0.00618206f $X=-0.19 $Y=-0.245 $X2=2.65 $Y2=2.055
cc_4 VNB N_A_91_269#_c_94_n 0.0285788f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=1.51
cc_5 VNB N_A_91_269#_c_95_n 0.0064741f $X=-0.19 $Y=-0.245 $X2=0.84 $Y2=1.495
cc_6 VNB N_A_91_269#_c_96_n 0.00416839f $X=-0.19 $Y=-0.245 $X2=2.565 $Y2=0.445
cc_7 VNB N_A1_N_c_187_n 0.0239769f $X=-0.19 $Y=-0.245 $X2=2.11 $Y2=2.645
cc_8 VNB N_A1_N_M1005_g 0.0320536f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A1_N_c_189_n 0.0108881f $X=-0.19 $Y=-0.245 $X2=0.685 $Y2=1.675
cc_10 VNB A1_N 0.00243711f $X=-0.19 $Y=-0.245 $X2=0.685 $Y2=2.465
cc_11 VNB N_A1_N_c_191_n 0.0211876f $X=-0.19 $Y=-0.245 $X2=2.565 $Y2=2.14
cc_12 VNB N_A2_N_M1007_g 0.00271115f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A2_N_M1006_g 0.0267857f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.345
cc_14 VNB N_A2_N_c_237_n 0.0189612f $X=-0.19 $Y=-0.245 $X2=0.685 $Y2=1.675
cc_15 VNB N_A2_N_c_238_n 0.0158791f $X=-0.19 $Y=-0.245 $X2=0.685 $Y2=2.465
cc_16 VNB N_A2_N_c_239_n 0.0152407f $X=-0.19 $Y=-0.245 $X2=0.84 $Y2=2.325
cc_17 VNB N_A2_N_c_240_n 0.0125896f $X=-0.19 $Y=-0.245 $X2=2.07 $Y2=2.41
cc_18 VNB N_A_271_47#_M1008_g 0.0299539f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=0.655
cc_19 VNB N_A_271_47#_c_285_n 0.0212765f $X=-0.19 $Y=-0.245 $X2=2.217 $Y2=2.495
cc_20 VNB N_A_271_47#_c_286_n 0.0094814f $X=-0.19 $Y=-0.245 $X2=2.217 $Y2=2.855
cc_21 VNB N_A_271_47#_c_287_n 0.0114293f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=1.495
cc_22 VNB N_A_271_47#_c_288_n 0.00305302f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=1.51
cc_23 VNB N_A_271_47#_c_289_n 9.00408e-19 $X=-0.19 $Y=-0.245 $X2=0.84 $Y2=1.495
cc_24 VNB N_A_271_47#_c_290_n 0.00381439f $X=-0.19 $Y=-0.245 $X2=2.217 $Y2=2.41
cc_25 VNB N_A_271_47#_c_291_n 0.0162183f $X=-0.19 $Y=-0.245 $X2=2.592 $Y2=0.445
cc_26 VNB N_A_271_47#_c_292_n 0.00169713f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=1.51
cc_27 VNB N_B2_M1002_g 0.0390906f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB B2 0.00749442f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=0.655
cc_29 VNB N_B2_c_376_n 0.0398886f $X=-0.19 $Y=-0.245 $X2=2.217 $Y2=2.855
cc_30 VNB N_B1_M1003_g 0.0268545f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_B1_c_424_n 0.0341557f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=0.655
cc_32 VNB N_B1_c_425_n 0.00804628f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_B1_c_426_n 0.00809048f $X=-0.19 $Y=-0.245 $X2=0.685 $Y2=2.465
cc_34 VNB N_B1_c_427_n 0.0175475f $X=-0.19 $Y=-0.245 $X2=2.217 $Y2=2.495
cc_35 VNB B1 0.0399056f $X=-0.19 $Y=-0.245 $X2=2.217 $Y2=2.855
cc_36 VNB N_B1_c_429_n 0.0288598f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=1.51
cc_37 VNB N_X_c_463_n 0.0270545f $X=-0.19 $Y=-0.245 $X2=0.84 $Y2=1.645
cc_38 VNB N_X_c_464_n 0.0288337f $X=-0.19 $Y=-0.245 $X2=2.565 $Y2=2.14
cc_39 VNB X 0.016273f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=1.51
cc_40 VNB N_VPWR_c_488_n 0.163682f $X=-0.19 $Y=-0.245 $X2=2.217 $Y2=2.41
cc_41 VNB N_VGND_c_553_n 0.010977f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_554_n 0.00560269f $X=-0.19 $Y=-0.245 $X2=2.217 $Y2=2.855
cc_43 VNB N_VGND_c_555_n 0.0132703f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_556_n 0.0194804f $X=-0.19 $Y=-0.245 $X2=2.365 $Y2=2.14
cc_45 VNB N_VGND_c_557_n 0.0259513f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=1.51
cc_46 VNB N_VGND_c_558_n 0.0315563f $X=-0.19 $Y=-0.245 $X2=2.217 $Y2=2.14
cc_47 VNB N_VGND_c_559_n 0.0248799f $X=-0.19 $Y=-0.245 $X2=0.62 $Y2=1.51
cc_48 VNB N_VGND_c_560_n 0.00631622f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_561_n 0.210148f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VPB N_A_91_269#_M1009_g 0.0255881f $X=-0.19 $Y=1.655 $X2=0.685 $Y2=2.465
cc_51 VPB N_A_91_269#_c_92_n 0.00115408f $X=-0.19 $Y=1.655 $X2=0.84 $Y2=2.325
cc_52 VPB N_A_91_269#_c_99_n 0.032617f $X=-0.19 $Y=1.655 $X2=2.07 $Y2=2.41
cc_53 VPB N_A_91_269#_c_100_n 0.00755783f $X=-0.19 $Y=1.655 $X2=2.217 $Y2=2.495
cc_54 VPB N_A_91_269#_c_101_n 0.0225831f $X=-0.19 $Y=1.655 $X2=2.235 $Y2=2.855
cc_55 VPB N_A_91_269#_c_102_n 0.00676831f $X=-0.19 $Y=1.655 $X2=2.565 $Y2=2.14
cc_56 VPB N_A_91_269#_c_93_n 0.00384004f $X=-0.19 $Y=1.655 $X2=2.65 $Y2=2.055
cc_57 VPB N_A_91_269#_c_94_n 0.0073607f $X=-0.19 $Y=1.655 $X2=0.62 $Y2=1.51
cc_58 VPB N_A1_N_M1000_g 0.0193984f $X=-0.19 $Y=1.655 $X2=0.59 $Y2=0.655
cc_59 VPB N_A1_N_c_189_n 0.00774305f $X=-0.19 $Y=1.655 $X2=0.685 $Y2=1.675
cc_60 VPB A1_N 0.00107592f $X=-0.19 $Y=1.655 $X2=0.685 $Y2=2.465
cc_61 VPB N_A2_N_M1007_g 0.0224105f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_62 VPB N_A_271_47#_M1010_g 0.0342057f $X=-0.19 $Y=1.655 $X2=0.84 $Y2=1.645
cc_63 VPB N_A_271_47#_c_286_n 0.00653818f $X=-0.19 $Y=1.655 $X2=2.217 $Y2=2.855
cc_64 VPB N_A_271_47#_c_295_n 0.0269016f $X=-0.19 $Y=1.655 $X2=2.235 $Y2=2.855
cc_65 VPB N_A_271_47#_c_296_n 0.0126856f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_66 VPB N_A_271_47#_c_290_n 5.88549e-19 $X=-0.19 $Y=1.655 $X2=2.217 $Y2=2.41
cc_67 VPB N_A_271_47#_c_298_n 0.0131511f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_68 VPB N_B2_M1004_g 0.0486415f $X=-0.19 $Y=1.655 $X2=0.59 $Y2=1.345
cc_69 VPB B2 0.00624493f $X=-0.19 $Y=1.655 $X2=0.59 $Y2=0.655
cc_70 VPB N_B2_c_376_n 0.0268047f $X=-0.19 $Y=1.655 $X2=2.217 $Y2=2.855
cc_71 VPB N_B1_M1001_g 0.0387273f $X=-0.19 $Y=1.655 $X2=0.59 $Y2=1.345
cc_72 VPB N_B1_c_426_n 0.0270476f $X=-0.19 $Y=1.655 $X2=0.685 $Y2=2.465
cc_73 VPB N_B1_c_432_n 0.0261846f $X=-0.19 $Y=1.655 $X2=0.84 $Y2=1.645
cc_74 VPB B1 0.0287903f $X=-0.19 $Y=1.655 $X2=2.217 $Y2=2.855
cc_75 VPB N_X_c_466_n 0.050776f $X=-0.19 $Y=1.655 $X2=0.685 $Y2=1.675
cc_76 VPB N_X_c_467_n 0.0187259f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_77 VPB N_X_c_463_n 0.00781712f $X=-0.19 $Y=1.655 $X2=0.84 $Y2=1.645
cc_78 VPB N_VPWR_c_489_n 0.0196139f $X=-0.19 $Y=1.655 $X2=0.59 $Y2=0.655
cc_79 VPB N_VPWR_c_490_n 0.00126149f $X=-0.19 $Y=1.655 $X2=0.685 $Y2=2.465
cc_80 VPB N_VPWR_c_491_n 0.0201769f $X=-0.19 $Y=1.655 $X2=0.84 $Y2=2.325
cc_81 VPB N_VPWR_c_492_n 0.00510842f $X=-0.19 $Y=1.655 $X2=2.07 $Y2=2.41
cc_82 VPB N_VPWR_c_493_n 0.0540757f $X=-0.19 $Y=1.655 $X2=2.365 $Y2=2.14
cc_83 VPB N_VPWR_c_494_n 0.0175582f $X=-0.19 $Y=1.655 $X2=2.217 $Y2=2.14
cc_84 VPB N_VPWR_c_488_n 0.0708572f $X=-0.19 $Y=1.655 $X2=2.217 $Y2=2.41
cc_85 VPB N_VPWR_c_496_n 0.00473485f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_86 VPB N_A_505_529#_c_528_n 0.00137967f $X=-0.19 $Y=1.655 $X2=0.59 $Y2=0.655
cc_87 VPB N_A_505_529#_c_529_n 0.0169498f $X=-0.19 $Y=1.655 $X2=0.685 $Y2=1.675
cc_88 VPB N_A_505_529#_c_530_n 0.00365501f $X=-0.19 $Y=1.655 $X2=0.685 $Y2=2.465
cc_89 VPB N_A_505_529#_c_531_n 0.0183176f $X=-0.19 $Y=1.655 $X2=0.84 $Y2=1.645
cc_90 N_A_91_269#_c_94_n N_A1_N_c_187_n 0.0172692f $X=0.62 $Y=1.51 $X2=0 $Y2=0
cc_91 N_A_91_269#_c_95_n N_A1_N_c_187_n 0.00220457f $X=0.84 $Y=1.495 $X2=0 $Y2=0
cc_92 N_A_91_269#_M1011_g N_A1_N_M1005_g 0.0102239f $X=0.59 $Y=0.655 $X2=0 $Y2=0
cc_93 N_A_91_269#_M1009_g N_A1_N_M1000_g 0.016263f $X=0.685 $Y=2.465 $X2=0 $Y2=0
cc_94 N_A_91_269#_c_92_n N_A1_N_M1000_g 0.0046648f $X=0.84 $Y=2.325 $X2=0 $Y2=0
cc_95 N_A_91_269#_c_99_n N_A1_N_M1000_g 0.00878163f $X=2.07 $Y=2.41 $X2=0 $Y2=0
cc_96 N_A_91_269#_c_92_n N_A1_N_c_189_n 2.01257e-19 $X=0.84 $Y=2.325 $X2=0 $Y2=0
cc_97 N_A_91_269#_c_99_n N_A1_N_c_189_n 0.00266904f $X=2.07 $Y=2.41 $X2=0 $Y2=0
cc_98 N_A_91_269#_M1011_g A1_N 0.00130008f $X=0.59 $Y=0.655 $X2=0 $Y2=0
cc_99 N_A_91_269#_M1009_g A1_N 0.00120295f $X=0.685 $Y=2.465 $X2=0 $Y2=0
cc_100 N_A_91_269#_c_92_n A1_N 0.0362041f $X=0.84 $Y=2.325 $X2=0 $Y2=0
cc_101 N_A_91_269#_c_99_n A1_N 0.0124076f $X=2.07 $Y=2.41 $X2=0 $Y2=0
cc_102 N_A_91_269#_c_94_n A1_N 2.86961e-19 $X=0.62 $Y=1.51 $X2=0 $Y2=0
cc_103 N_A_91_269#_c_95_n A1_N 0.0224445f $X=0.84 $Y=1.495 $X2=0 $Y2=0
cc_104 N_A_91_269#_M1011_g N_A1_N_c_191_n 0.0108447f $X=0.59 $Y=0.655 $X2=0
+ $Y2=0
cc_105 N_A_91_269#_c_99_n N_A2_N_M1007_g 0.011688f $X=2.07 $Y=2.41 $X2=0 $Y2=0
cc_106 N_A_91_269#_c_100_n N_A2_N_M1007_g 0.00353586f $X=2.217 $Y=2.495 $X2=0
+ $Y2=0
cc_107 N_A_91_269#_c_93_n N_A_271_47#_M1008_g 0.00238649f $X=2.65 $Y=2.055 $X2=0
+ $Y2=0
cc_108 N_A_91_269#_c_96_n N_A_271_47#_M1008_g 3.95974e-19 $X=2.565 $Y=0.445
+ $X2=0 $Y2=0
cc_109 N_A_91_269#_c_100_n N_A_271_47#_M1010_g 0.00624846f $X=2.217 $Y=2.495
+ $X2=0 $Y2=0
cc_110 N_A_91_269#_c_101_n N_A_271_47#_M1010_g 0.00383455f $X=2.235 $Y=2.855
+ $X2=0 $Y2=0
cc_111 N_A_91_269#_c_100_n N_A_271_47#_c_286_n 8.89446e-19 $X=2.217 $Y=2.495
+ $X2=0 $Y2=0
cc_112 N_A_91_269#_c_100_n N_A_271_47#_c_295_n 0.00218262f $X=2.217 $Y=2.495
+ $X2=0 $Y2=0
cc_113 N_A_91_269#_c_102_n N_A_271_47#_c_295_n 0.00549761f $X=2.565 $Y=2.14
+ $X2=0 $Y2=0
cc_114 N_A_91_269#_c_100_n N_A_271_47#_c_296_n 0.00485183f $X=2.217 $Y=2.495
+ $X2=0 $Y2=0
cc_115 N_A_91_269#_c_102_n N_A_271_47#_c_296_n 0.00991677f $X=2.565 $Y=2.14
+ $X2=0 $Y2=0
cc_116 N_A_91_269#_c_93_n N_A_271_47#_c_287_n 0.00863569f $X=2.65 $Y=2.055 $X2=0
+ $Y2=0
cc_117 N_A_91_269#_c_96_n N_A_271_47#_c_287_n 8.2986e-19 $X=2.565 $Y=0.445 $X2=0
+ $Y2=0
cc_118 N_A_91_269#_c_93_n N_A_271_47#_c_289_n 0.0495206f $X=2.65 $Y=2.055 $X2=0
+ $Y2=0
cc_119 N_A_91_269#_c_93_n N_A_271_47#_c_291_n 0.00773397f $X=2.65 $Y=2.055 $X2=0
+ $Y2=0
cc_120 N_A_91_269#_c_96_n N_A_271_47#_c_291_n 5.34646e-19 $X=2.565 $Y=0.445
+ $X2=0 $Y2=0
cc_121 N_A_91_269#_c_99_n N_A_271_47#_c_298_n 0.0182359f $X=2.07 $Y=2.41 $X2=0
+ $Y2=0
cc_122 N_A_91_269#_c_100_n N_A_271_47#_c_298_n 0.0288702f $X=2.217 $Y=2.495
+ $X2=0 $Y2=0
cc_123 N_A_91_269#_c_102_n N_A_271_47#_c_298_n 0.00138211f $X=2.565 $Y=2.14
+ $X2=0 $Y2=0
cc_124 N_A_91_269#_c_93_n N_A_271_47#_c_298_n 0.0184633f $X=2.65 $Y=2.055 $X2=0
+ $Y2=0
cc_125 N_A_91_269#_c_93_n N_A_271_47#_c_292_n 0.00823056f $X=2.65 $Y=2.055 $X2=0
+ $Y2=0
cc_126 N_A_91_269#_c_93_n N_B2_M1002_g 0.00975187f $X=2.65 $Y=2.055 $X2=0 $Y2=0
cc_127 N_A_91_269#_c_96_n N_B2_M1002_g 0.00479906f $X=2.565 $Y=0.445 $X2=0 $Y2=0
cc_128 N_A_91_269#_c_100_n N_B2_M1004_g 2.99919e-19 $X=2.217 $Y=2.495 $X2=0
+ $Y2=0
cc_129 N_A_91_269#_c_102_n N_B2_M1004_g 0.00139315f $X=2.565 $Y=2.14 $X2=0 $Y2=0
cc_130 N_A_91_269#_c_93_n N_B2_M1004_g 0.00118103f $X=2.65 $Y=2.055 $X2=0 $Y2=0
cc_131 N_A_91_269#_c_102_n B2 0.0134326f $X=2.565 $Y=2.14 $X2=0 $Y2=0
cc_132 N_A_91_269#_c_96_n B2 0.124961f $X=2.565 $Y=0.445 $X2=0 $Y2=0
cc_133 N_A_91_269#_c_93_n N_B2_c_376_n 0.0157628f $X=2.65 $Y=2.055 $X2=0 $Y2=0
cc_134 N_A_91_269#_c_96_n N_B1_M1003_g 2.78053e-19 $X=2.565 $Y=0.445 $X2=0 $Y2=0
cc_135 N_A_91_269#_c_93_n N_B1_c_425_n 2.78053e-19 $X=2.65 $Y=2.055 $X2=0 $Y2=0
cc_136 N_A_91_269#_M1009_g N_X_c_467_n 0.00336744f $X=0.685 $Y=2.465 $X2=0 $Y2=0
cc_137 N_A_91_269#_c_92_n N_X_c_467_n 0.016548f $X=0.84 $Y=2.325 $X2=0 $Y2=0
cc_138 N_A_91_269#_c_94_n N_X_c_467_n 0.00283243f $X=0.62 $Y=1.51 $X2=0 $Y2=0
cc_139 N_A_91_269#_c_95_n N_X_c_467_n 0.00913238f $X=0.84 $Y=1.495 $X2=0 $Y2=0
cc_140 N_A_91_269#_M1011_g N_X_c_463_n 0.00644694f $X=0.59 $Y=0.655 $X2=0 $Y2=0
cc_141 N_A_91_269#_M1009_g N_X_c_463_n 0.0016442f $X=0.685 $Y=2.465 $X2=0 $Y2=0
cc_142 N_A_91_269#_c_92_n N_X_c_463_n 0.00401392f $X=0.84 $Y=2.325 $X2=0 $Y2=0
cc_143 N_A_91_269#_c_94_n N_X_c_463_n 0.00291743f $X=0.62 $Y=1.51 $X2=0 $Y2=0
cc_144 N_A_91_269#_c_95_n N_X_c_463_n 0.0232272f $X=0.84 $Y=1.495 $X2=0 $Y2=0
cc_145 N_A_91_269#_M1011_g X 0.00288913f $X=0.59 $Y=0.655 $X2=0 $Y2=0
cc_146 N_A_91_269#_c_94_n X 0.0010927f $X=0.62 $Y=1.51 $X2=0 $Y2=0
cc_147 N_A_91_269#_c_95_n X 0.00307952f $X=0.84 $Y=1.495 $X2=0 $Y2=0
cc_148 N_A_91_269#_c_92_n N_VPWR_M1009_d 0.00498935f $X=0.84 $Y=2.325 $X2=-0.19
+ $Y2=-0.245
cc_149 N_A_91_269#_c_99_n N_VPWR_M1009_d 0.00560553f $X=2.07 $Y=2.41 $X2=-0.19
+ $Y2=-0.245
cc_150 N_A_91_269#_c_165_p N_VPWR_M1009_d 0.00116756f $X=0.925 $Y=2.41 $X2=-0.19
+ $Y2=-0.245
cc_151 N_A_91_269#_M1009_g N_VPWR_c_489_n 0.0140949f $X=0.685 $Y=2.465 $X2=0
+ $Y2=0
cc_152 N_A_91_269#_c_99_n N_VPWR_c_489_n 0.01114f $X=2.07 $Y=2.41 $X2=0 $Y2=0
cc_153 N_A_91_269#_c_165_p N_VPWR_c_489_n 0.0097857f $X=0.925 $Y=2.41 $X2=0
+ $Y2=0
cc_154 N_A_91_269#_M1009_g N_VPWR_c_491_n 0.00486043f $X=0.685 $Y=2.465 $X2=0
+ $Y2=0
cc_155 N_A_91_269#_c_101_n N_VPWR_c_493_n 0.0140996f $X=2.235 $Y=2.855 $X2=0
+ $Y2=0
cc_156 N_A_91_269#_M1009_g N_VPWR_c_488_n 0.0093271f $X=0.685 $Y=2.465 $X2=0
+ $Y2=0
cc_157 N_A_91_269#_c_99_n N_VPWR_c_488_n 0.0353481f $X=2.07 $Y=2.41 $X2=0 $Y2=0
cc_158 N_A_91_269#_c_165_p N_VPWR_c_488_n 6.1821e-19 $X=0.925 $Y=2.41 $X2=0
+ $Y2=0
cc_159 N_A_91_269#_c_101_n N_VPWR_c_488_n 0.0110771f $X=2.235 $Y=2.855 $X2=0
+ $Y2=0
cc_160 N_A_91_269#_c_101_n N_A_505_529#_c_528_n 0.00629364f $X=2.235 $Y=2.855
+ $X2=0 $Y2=0
cc_161 N_A_91_269#_c_100_n N_A_505_529#_c_530_n 0.00936298f $X=2.217 $Y=2.495
+ $X2=0 $Y2=0
cc_162 N_A_91_269#_c_101_n N_A_505_529#_c_530_n 0.00609749f $X=2.235 $Y=2.855
+ $X2=0 $Y2=0
cc_163 N_A_91_269#_c_102_n N_A_505_529#_c_530_n 0.0182603f $X=2.565 $Y=2.14
+ $X2=0 $Y2=0
cc_164 N_A_91_269#_M1011_g N_VGND_c_553_n 0.00493472f $X=0.59 $Y=0.655 $X2=0
+ $Y2=0
cc_165 N_A_91_269#_c_94_n N_VGND_c_553_n 0.00273476f $X=0.62 $Y=1.51 $X2=0 $Y2=0
cc_166 N_A_91_269#_c_95_n N_VGND_c_553_n 0.0162398f $X=0.84 $Y=1.495 $X2=0 $Y2=0
cc_167 N_A_91_269#_c_96_n N_VGND_c_558_n 0.0142541f $X=2.565 $Y=0.445 $X2=0
+ $Y2=0
cc_168 N_A_91_269#_M1011_g N_VGND_c_559_n 0.00585385f $X=0.59 $Y=0.655 $X2=0
+ $Y2=0
cc_169 N_A_91_269#_M1008_d N_VGND_c_561_n 0.00316506f $X=2.425 $Y=0.235 $X2=0
+ $Y2=0
cc_170 N_A_91_269#_M1011_g N_VGND_c_561_n 0.0120756f $X=0.59 $Y=0.655 $X2=0
+ $Y2=0
cc_171 N_A_91_269#_c_96_n N_VGND_c_561_n 0.0106583f $X=2.565 $Y=0.445 $X2=0
+ $Y2=0
cc_172 N_A1_N_M1000_g N_A2_N_M1007_g 0.0361689f $X=1.28 $Y=2.045 $X2=0 $Y2=0
cc_173 N_A1_N_M1005_g N_A2_N_M1006_g 0.0158124f $X=1.28 $Y=0.445 $X2=0 $Y2=0
cc_174 A1_N N_A2_N_M1006_g 7.82713e-19 $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_175 N_A1_N_c_187_n N_A2_N_c_237_n 0.0129593f $X=1.197 $Y=1.503 $X2=0 $Y2=0
cc_176 N_A1_N_c_189_n N_A2_N_c_238_n 0.0129593f $X=1.197 $Y=1.675 $X2=0 $Y2=0
cc_177 A1_N N_A2_N_c_238_n 0.00253242f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_178 N_A1_N_M1005_g N_A2_N_c_239_n 0.00387383f $X=1.28 $Y=0.445 $X2=0 $Y2=0
cc_179 A1_N N_A2_N_c_239_n 9.38761e-19 $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_180 N_A1_N_c_191_n N_A2_N_c_239_n 0.0129593f $X=1.205 $Y=1.17 $X2=0 $Y2=0
cc_181 A1_N N_A2_N_c_240_n 0.0398604f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_182 N_A1_N_c_191_n N_A2_N_c_240_n 0.00358175f $X=1.205 $Y=1.17 $X2=0 $Y2=0
cc_183 N_A1_N_M1005_g N_A_271_47#_c_318_n 0.00155924f $X=1.28 $Y=0.445 $X2=0
+ $Y2=0
cc_184 A1_N N_A_271_47#_c_318_n 0.0214943f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_185 N_A1_N_M1005_g N_A_271_47#_c_288_n 0.00133491f $X=1.28 $Y=0.445 $X2=0
+ $Y2=0
cc_186 A1_N N_A_271_47#_c_288_n 0.013815f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_187 A1_N N_A_271_47#_c_298_n 0.00929965f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_188 A1_N N_VPWR_M1009_d 0.00340567f $X=1.115 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_189 A1_N N_VGND_M1011_d 0.00317155f $X=1.115 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_190 N_A1_N_M1005_g N_VGND_c_553_n 0.00591665f $X=1.28 $Y=0.445 $X2=0 $Y2=0
cc_191 A1_N N_VGND_c_553_n 0.055724f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_192 N_A1_N_c_191_n N_VGND_c_553_n 7.86781e-19 $X=1.205 $Y=1.17 $X2=0 $Y2=0
cc_193 N_A1_N_M1005_g N_VGND_c_557_n 0.00463859f $X=1.28 $Y=0.445 $X2=0 $Y2=0
cc_194 A1_N N_VGND_c_557_n 0.00631844f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_195 N_A1_N_M1005_g N_VGND_c_561_n 0.00846256f $X=1.28 $Y=0.445 $X2=0 $Y2=0
cc_196 A1_N N_VGND_c_561_n 0.00642626f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_197 N_A2_N_M1006_g N_A_271_47#_M1008_g 0.0191985f $X=1.765 $Y=0.445 $X2=0
+ $Y2=0
cc_198 N_A2_N_c_239_n N_A_271_47#_M1008_g 0.00219611f $X=1.76 $Y=1.1 $X2=0 $Y2=0
cc_199 N_A2_N_M1007_g N_A_271_47#_M1010_g 0.00104312f $X=1.67 $Y=2.045 $X2=0
+ $Y2=0
cc_200 N_A2_N_c_237_n N_A_271_47#_c_285_n 0.012865f $X=1.76 $Y=1.44 $X2=0 $Y2=0
cc_201 N_A2_N_M1007_g N_A_271_47#_c_286_n 0.00187502f $X=1.67 $Y=2.045 $X2=0
+ $Y2=0
cc_202 N_A2_N_c_238_n N_A_271_47#_c_286_n 0.012865f $X=1.76 $Y=1.605 $X2=0 $Y2=0
cc_203 N_A2_N_M1007_g N_A_271_47#_c_295_n 0.00627003f $X=1.67 $Y=2.045 $X2=0
+ $Y2=0
cc_204 N_A2_N_M1006_g N_A_271_47#_c_318_n 0.00609829f $X=1.765 $Y=0.445 $X2=0
+ $Y2=0
cc_205 N_A2_N_M1006_g N_A_271_47#_c_287_n 0.00936626f $X=1.765 $Y=0.445 $X2=0
+ $Y2=0
cc_206 N_A2_N_c_239_n N_A_271_47#_c_287_n 0.00240694f $X=1.76 $Y=1.1 $X2=0 $Y2=0
cc_207 N_A2_N_c_240_n N_A_271_47#_c_287_n 0.0151307f $X=1.76 $Y=1.1 $X2=0 $Y2=0
cc_208 N_A2_N_M1006_g N_A_271_47#_c_288_n 0.00250553f $X=1.765 $Y=0.445 $X2=0
+ $Y2=0
cc_209 N_A2_N_c_239_n N_A_271_47#_c_288_n 0.00281149f $X=1.76 $Y=1.1 $X2=0 $Y2=0
cc_210 N_A2_N_c_240_n N_A_271_47#_c_288_n 0.0209431f $X=1.76 $Y=1.1 $X2=0 $Y2=0
cc_211 N_A2_N_c_239_n N_A_271_47#_c_289_n 8.2468e-19 $X=1.76 $Y=1.1 $X2=0 $Y2=0
cc_212 N_A2_N_c_240_n N_A_271_47#_c_289_n 0.0381725f $X=1.76 $Y=1.1 $X2=0 $Y2=0
cc_213 N_A2_N_M1007_g N_A_271_47#_c_290_n 0.00190348f $X=1.67 $Y=2.045 $X2=0
+ $Y2=0
cc_214 N_A2_N_c_237_n N_A_271_47#_c_290_n 8.2468e-19 $X=1.76 $Y=1.44 $X2=0 $Y2=0
cc_215 N_A2_N_c_238_n N_A_271_47#_c_290_n 0.00178597f $X=1.76 $Y=1.605 $X2=0
+ $Y2=0
cc_216 N_A2_N_c_239_n N_A_271_47#_c_291_n 0.012865f $X=1.76 $Y=1.1 $X2=0 $Y2=0
cc_217 N_A2_N_c_240_n N_A_271_47#_c_291_n 6.05912e-19 $X=1.76 $Y=1.1 $X2=0 $Y2=0
cc_218 N_A2_N_M1007_g N_A_271_47#_c_298_n 0.00226798f $X=1.67 $Y=2.045 $X2=0
+ $Y2=0
cc_219 N_A2_N_c_238_n N_A_271_47#_c_298_n 0.00422898f $X=1.76 $Y=1.605 $X2=0
+ $Y2=0
cc_220 N_A2_N_c_240_n N_A_271_47#_c_298_n 0.0116597f $X=1.76 $Y=1.1 $X2=0 $Y2=0
cc_221 N_A2_N_M1006_g N_A_271_47#_c_292_n 0.00194466f $X=1.765 $Y=0.445 $X2=0
+ $Y2=0
cc_222 N_A2_N_c_239_n N_A_271_47#_c_292_n 0.00175078f $X=1.76 $Y=1.1 $X2=0 $Y2=0
cc_223 N_A2_N_M1006_g N_VGND_c_554_n 0.0047565f $X=1.765 $Y=0.445 $X2=0 $Y2=0
cc_224 N_A2_N_M1006_g N_VGND_c_557_n 0.00419847f $X=1.765 $Y=0.445 $X2=0 $Y2=0
cc_225 N_A2_N_M1006_g N_VGND_c_561_n 0.00638767f $X=1.765 $Y=0.445 $X2=0 $Y2=0
cc_226 N_A_271_47#_M1008_g N_B2_M1002_g 0.0219787f $X=2.35 $Y=0.445 $X2=0 $Y2=0
cc_227 N_A_271_47#_c_289_n N_B2_M1002_g 3.04926e-19 $X=2.247 $Y=1.142 $X2=0
+ $Y2=0
cc_228 N_A_271_47#_c_291_n N_B2_M1002_g 0.0229881f $X=2.3 $Y=1.17 $X2=0 $Y2=0
cc_229 N_A_271_47#_c_295_n N_B2_M1004_g 0.00667567f $X=2.42 $Y=2.14 $X2=0 $Y2=0
cc_230 N_A_271_47#_c_296_n N_B2_M1004_g 0.0285069f $X=2.42 $Y=2.29 $X2=0 $Y2=0
cc_231 N_A_271_47#_c_295_n B2 2.83745e-19 $X=2.42 $Y=2.14 $X2=0 $Y2=0
cc_232 N_A_271_47#_c_286_n N_B2_c_376_n 0.0229881f $X=2.3 $Y=1.675 $X2=0 $Y2=0
cc_233 N_A_271_47#_c_290_n N_B2_c_376_n 3.04926e-19 $X=2.3 $Y=1.17 $X2=0 $Y2=0
cc_234 N_A_271_47#_M1010_g N_VPWR_c_490_n 0.00118108f $X=2.45 $Y=2.855 $X2=0
+ $Y2=0
cc_235 N_A_271_47#_M1010_g N_VPWR_c_493_n 0.00555245f $X=2.45 $Y=2.855 $X2=0
+ $Y2=0
cc_236 N_A_271_47#_M1010_g N_VPWR_c_488_n 0.0117713f $X=2.45 $Y=2.855 $X2=0
+ $Y2=0
cc_237 N_A_271_47#_M1010_g N_A_505_529#_c_528_n 6.94016e-19 $X=2.45 $Y=2.855
+ $X2=0 $Y2=0
cc_238 N_A_271_47#_M1010_g N_A_505_529#_c_530_n 0.00150843f $X=2.45 $Y=2.855
+ $X2=0 $Y2=0
cc_239 N_A_271_47#_c_318_n N_VGND_c_553_n 0.00297469f $X=1.55 $Y=0.445 $X2=0
+ $Y2=0
cc_240 N_A_271_47#_M1008_g N_VGND_c_554_n 0.00470957f $X=2.35 $Y=0.445 $X2=0
+ $Y2=0
cc_241 N_A_271_47#_c_287_n N_VGND_c_554_n 0.0262111f $X=2.11 $Y=0.75 $X2=0 $Y2=0
cc_242 N_A_271_47#_c_291_n N_VGND_c_554_n 3.1304e-19 $X=2.3 $Y=1.17 $X2=0 $Y2=0
cc_243 N_A_271_47#_c_318_n N_VGND_c_557_n 0.0130869f $X=1.55 $Y=0.445 $X2=0
+ $Y2=0
cc_244 N_A_271_47#_c_287_n N_VGND_c_557_n 0.00274686f $X=2.11 $Y=0.75 $X2=0
+ $Y2=0
cc_245 N_A_271_47#_M1008_g N_VGND_c_558_n 0.00580182f $X=2.35 $Y=0.445 $X2=0
+ $Y2=0
cc_246 N_A_271_47#_c_287_n N_VGND_c_558_n 0.00112271f $X=2.11 $Y=0.75 $X2=0
+ $Y2=0
cc_247 N_A_271_47#_M1005_d N_VGND_c_561_n 0.00656323f $X=1.355 $Y=0.235 $X2=0
+ $Y2=0
cc_248 N_A_271_47#_M1008_g N_VGND_c_561_n 0.0111056f $X=2.35 $Y=0.445 $X2=0
+ $Y2=0
cc_249 N_A_271_47#_c_318_n N_VGND_c_561_n 0.0093482f $X=1.55 $Y=0.445 $X2=0
+ $Y2=0
cc_250 N_A_271_47#_c_287_n N_VGND_c_561_n 0.00746008f $X=2.11 $Y=0.75 $X2=0
+ $Y2=0
cc_251 N_B2_M1002_g N_B1_M1003_g 0.0450939f $X=2.78 $Y=0.445 $X2=0 $Y2=0
cc_252 B2 N_B1_M1003_g 0.0223278f $X=3.035 $Y=0.47 $X2=0 $Y2=0
cc_253 B2 N_B1_c_425_n 0.00681618f $X=3.035 $Y=0.47 $X2=0 $Y2=0
cc_254 N_B2_c_376_n N_B1_c_425_n 0.00387985f $X=3 $Y=1.395 $X2=0 $Y2=0
cc_255 N_B2_M1004_g N_B1_c_426_n 0.00480583f $X=2.88 $Y=2.855 $X2=0 $Y2=0
cc_256 N_B2_M1004_g N_B1_c_432_n 0.0317096f $X=2.88 $Y=2.855 $X2=0 $Y2=0
cc_257 B2 N_B1_c_432_n 0.00101149f $X=3.035 $Y=0.47 $X2=0 $Y2=0
cc_258 N_B2_M1004_g B1 5.53266e-19 $X=2.88 $Y=2.855 $X2=0 $Y2=0
cc_259 B2 B1 0.113764f $X=3.035 $Y=0.47 $X2=0 $Y2=0
cc_260 N_B2_c_376_n B1 0.00204885f $X=3 $Y=1.395 $X2=0 $Y2=0
cc_261 N_B2_M1002_g N_B1_c_429_n 0.00340754f $X=2.78 $Y=0.445 $X2=0 $Y2=0
cc_262 B2 N_B1_c_429_n 0.00387347f $X=3.035 $Y=0.47 $X2=0 $Y2=0
cc_263 N_B2_c_376_n N_B1_c_429_n 0.0367742f $X=3 $Y=1.395 $X2=0 $Y2=0
cc_264 N_B2_M1004_g N_VPWR_c_490_n 0.00891614f $X=2.88 $Y=2.855 $X2=0 $Y2=0
cc_265 N_B2_M1004_g N_VPWR_c_493_n 0.00461019f $X=2.88 $Y=2.855 $X2=0 $Y2=0
cc_266 N_B2_M1004_g N_VPWR_c_488_n 0.00433009f $X=2.88 $Y=2.855 $X2=0 $Y2=0
cc_267 N_B2_M1004_g N_A_505_529#_c_528_n 0.00115618f $X=2.88 $Y=2.855 $X2=0
+ $Y2=0
cc_268 N_B2_M1004_g N_A_505_529#_c_529_n 0.0145015f $X=2.88 $Y=2.855 $X2=0 $Y2=0
cc_269 B2 N_A_505_529#_c_529_n 0.024846f $X=3.035 $Y=0.47 $X2=0 $Y2=0
cc_270 N_B2_c_376_n N_A_505_529#_c_529_n 0.0020414f $X=3 $Y=1.395 $X2=0 $Y2=0
cc_271 N_B2_c_376_n N_A_505_529#_c_530_n 9.77949e-19 $X=3 $Y=1.395 $X2=0 $Y2=0
cc_272 B2 N_VGND_c_556_n 0.0250463f $X=3.035 $Y=0.47 $X2=0 $Y2=0
cc_273 N_B2_M1002_g N_VGND_c_558_n 0.00542362f $X=2.78 $Y=0.445 $X2=0 $Y2=0
cc_274 B2 N_VGND_c_558_n 0.0161138f $X=3.035 $Y=0.47 $X2=0 $Y2=0
cc_275 N_B2_M1002_g N_VGND_c_561_n 0.00985329f $X=2.78 $Y=0.445 $X2=0 $Y2=0
cc_276 B2 N_VGND_c_561_n 0.0108915f $X=3.035 $Y=0.47 $X2=0 $Y2=0
cc_277 B2 A_571_47# 0.00443436f $X=3.035 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_278 N_B1_M1001_g N_VPWR_c_490_n 0.0107019f $X=3.31 $Y=2.855 $X2=0 $Y2=0
cc_279 N_B1_M1001_g N_VPWR_c_494_n 0.00461019f $X=3.31 $Y=2.855 $X2=0 $Y2=0
cc_280 N_B1_M1001_g N_VPWR_c_488_n 0.00513842f $X=3.31 $Y=2.855 $X2=0 $Y2=0
cc_281 N_B1_M1001_g N_A_505_529#_c_529_n 0.0167746f $X=3.31 $Y=2.855 $X2=0 $Y2=0
cc_282 N_B1_c_432_n N_A_505_529#_c_529_n 0.00461385f $X=3.48 $Y=2.185 $X2=0
+ $Y2=0
cc_283 B1 N_A_505_529#_c_529_n 0.027119f $X=3.515 $Y=0.84 $X2=0 $Y2=0
cc_284 N_B1_M1001_g N_A_505_529#_c_531_n 0.00261315f $X=3.31 $Y=2.855 $X2=0
+ $Y2=0
cc_285 N_B1_M1003_g N_VGND_c_556_n 0.0120429f $X=3.17 $Y=0.445 $X2=0 $Y2=0
cc_286 N_B1_c_424_n N_VGND_c_556_n 0.00201481f $X=3.405 $Y=0.915 $X2=0 $Y2=0
cc_287 B1 N_VGND_c_556_n 0.0176563f $X=3.515 $Y=0.84 $X2=0 $Y2=0
cc_288 N_B1_M1003_g N_VGND_c_558_n 0.00408844f $X=3.17 $Y=0.445 $X2=0 $Y2=0
cc_289 N_B1_M1003_g N_VGND_c_561_n 0.00764877f $X=3.17 $Y=0.445 $X2=0 $Y2=0
cc_290 N_B1_c_424_n N_VGND_c_561_n 0.00286559f $X=3.405 $Y=0.915 $X2=0 $Y2=0
cc_291 B1 N_VGND_c_561_n 0.00463609f $X=3.515 $Y=0.84 $X2=0 $Y2=0
cc_292 N_X_c_466_n N_VPWR_c_491_n 0.0321484f $X=0.47 $Y=2.91 $X2=0 $Y2=0
cc_293 N_X_M1009_s N_VPWR_c_488_n 0.00371702f $X=0.345 $Y=1.835 $X2=0 $Y2=0
cc_294 N_X_c_466_n N_VPWR_c_488_n 0.017806f $X=0.47 $Y=2.91 $X2=0 $Y2=0
cc_295 X N_VGND_c_553_n 0.00157626f $X=0.24 $Y=0.925 $X2=0 $Y2=0
cc_296 N_X_c_464_n N_VGND_c_559_n 0.02658f $X=0.375 $Y=0.42 $X2=0 $Y2=0
cc_297 N_X_M1011_s N_VGND_c_561_n 0.00249946f $X=0.25 $Y=0.235 $X2=0 $Y2=0
cc_298 N_X_c_464_n N_VGND_c_561_n 0.0154733f $X=0.375 $Y=0.42 $X2=0 $Y2=0
cc_299 N_VPWR_c_493_n N_A_505_529#_c_528_n 0.0100873f $X=2.93 $Y=3.33 $X2=0
+ $Y2=0
cc_300 N_VPWR_c_488_n N_A_505_529#_c_528_n 0.00840669f $X=3.6 $Y=3.33 $X2=0
+ $Y2=0
cc_301 N_VPWR_c_490_n N_A_505_529#_c_529_n 0.0208172f $X=3.095 $Y=2.855 $X2=0
+ $Y2=0
cc_302 N_VPWR_c_488_n N_A_505_529#_c_529_n 0.0119053f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_303 N_VPWR_c_494_n N_A_505_529#_c_531_n 0.0130724f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_304 N_VPWR_c_488_n N_A_505_529#_c_531_n 0.00972613f $X=3.6 $Y=3.33 $X2=0
+ $Y2=0
cc_305 N_VGND_c_561_n A_571_47# 0.00405832f $X=3.6 $Y=0 $X2=-0.19 $Y2=-0.245
