# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__o41ai_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_lp__o41ai_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.240000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.320000 1.335000 6.115000 1.750000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.930000 1.335000 5.150000 1.750000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.385000 1.335000 3.760000 1.750000 ;
    END
  END A3
  PIN A4
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.455000 1.335000 3.215000 1.750000 ;
    END
  END A4
  PIN B1
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.155000 1.015000 1.065000 1.525000 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  0.940800 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.615000 1.705000 2.285000 1.875000 ;
        RECT 0.615000 1.875000 0.835000 3.075000 ;
        RECT 1.235000 0.595000 1.485000 1.335000 ;
        RECT 1.235000 1.335000 2.285000 1.705000 ;
        RECT 1.955000 1.875000 2.285000 2.715000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 6.240000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 6.240000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.240000 0.085000 ;
      RECT 0.000000  3.245000 6.240000 3.415000 ;
      RECT 0.145000  1.815000 0.445000 3.245000 ;
      RECT 0.735000  0.255000 1.925000 0.425000 ;
      RECT 0.735000  0.425000 1.065000 0.845000 ;
      RECT 1.005000  2.045000 1.335000 3.245000 ;
      RECT 1.525000  2.045000 1.785000 2.895000 ;
      RECT 1.525000  2.895000 2.840000 3.075000 ;
      RECT 1.655000  0.425000 1.925000 0.995000 ;
      RECT 1.655000  0.995000 5.610000 1.165000 ;
      RECT 2.100000  0.085000 2.430000 0.825000 ;
      RECT 2.510000  1.920000 3.810000 2.090000 ;
      RECT 2.510000  2.090000 2.840000 2.895000 ;
      RECT 2.620000  0.255000 2.900000 0.995000 ;
      RECT 3.050000  2.260000 3.380000 2.905000 ;
      RECT 3.050000  2.905000 4.760000 3.075000 ;
      RECT 3.070000  0.085000 3.400000 0.825000 ;
      RECT 3.550000  2.090000 3.810000 2.735000 ;
      RECT 3.570000  0.255000 3.800000 0.995000 ;
      RECT 3.970000  0.085000 4.300000 0.825000 ;
      RECT 4.000000  1.920000 6.050000 2.090000 ;
      RECT 4.000000  2.090000 4.260000 2.735000 ;
      RECT 4.430000  2.260000 4.760000 2.905000 ;
      RECT 4.470000  0.255000 4.660000 0.995000 ;
      RECT 4.830000  0.085000 5.160000 0.825000 ;
      RECT 4.930000  2.090000 5.120000 3.075000 ;
      RECT 5.290000  2.260000 5.620000 3.245000 ;
      RECT 5.340000  0.255000 5.610000 0.995000 ;
      RECT 5.790000  2.090000 6.050000 3.075000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
  END
END sky130_fd_sc_lp__o41ai_2
END LIBRARY
