* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__or3b_m A B C_N VGND VNB VPB VPWR X
M1000 a_112_55# C_N VGND VNB nshort w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=3.465e+11p ps=4.17e+06u
M1001 X a_212_418# VGND VNB nshort w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1002 a_212_418# B VGND VNB nshort w=420000u l=150000u
+  ad=2.289e+11p pd=2.77e+06u as=0p ps=0u
M1003 a_371_418# B a_299_418# VPB phighvt w=420000u l=150000u
+  ad=1.638e+11p pd=1.62e+06u as=8.82e+10p ps=1.26e+06u
M1004 a_299_418# a_112_55# a_212_418# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.16025e+11p ps=1.41e+06u
M1005 a_112_55# C_N VPWR VPB phighvt w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=2.478e+11p ps=2.86e+06u
M1006 X a_212_418# VPWR VPB phighvt w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=0p ps=0u
M1007 VGND A a_212_418# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND a_112_55# a_212_418# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR A a_371_418# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
