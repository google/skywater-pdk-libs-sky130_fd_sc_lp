* File: sky130_fd_sc_lp__sregsbp_1.pex.spice
* Created: Fri Aug 28 11:33:43 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__SREGSBP_1%SCE 3 7 9 13 17 19 23 24 26 27 37 41 47 49
c83 24 0 2.8797e-19 $X=2.295 $Y=1.45
c84 13 0 1.19902e-19 $X=1.245 $Y=2.865
r85 41 47 1.74613 $w=3.28e-07 $l=5e-08 $layer=LI1_cond $X=1.15 $Y=1.64 $X2=1.2
+ $Y2=1.64
r86 36 37 30.474 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=0.735 $Y=1.64
+ $X2=0.81 $Y2=1.64
r87 34 36 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=0.645 $Y=1.64
+ $X2=0.735 $Y2=1.64
r88 31 34 26.2292 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=0.495 $Y=1.64
+ $X2=0.645 $Y2=1.64
r89 27 49 6.12237 $w=3.28e-07 $l=9.8e-08 $layer=LI1_cond $X=1.217 $Y=1.64
+ $X2=1.315 $Y2=1.64
r90 27 47 0.593683 $w=3.28e-07 $l=1.7e-08 $layer=LI1_cond $X=1.217 $Y=1.64
+ $X2=1.2 $Y2=1.64
r91 27 41 0.628605 $w=3.28e-07 $l=1.8e-08 $layer=LI1_cond $X=1.132 $Y=1.64
+ $X2=1.15 $Y2=1.64
r92 26 27 17.0073 $w=3.28e-07 $l=4.87e-07 $layer=LI1_cond $X=0.645 $Y=1.64
+ $X2=1.132 $Y2=1.64
r93 26 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.645
+ $Y=1.64 $X2=0.645 $Y2=1.64
r94 24 39 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.295 $Y=1.45
+ $X2=2.295 $Y2=1.285
r95 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.295
+ $Y=1.45 $X2=2.295 $Y2=1.45
r96 21 23 6.66256 $w=3.18e-07 $l=1.85e-07 $layer=LI1_cond $X=2.29 $Y=1.635
+ $X2=2.29 $Y2=1.45
r97 19 21 7.68211 $w=1.7e-07 $l=1.9799e-07 $layer=LI1_cond $X=2.13 $Y=1.72
+ $X2=2.29 $Y2=1.635
r98 19 49 53.1711 $w=1.68e-07 $l=8.15e-07 $layer=LI1_cond $X=2.13 $Y=1.72
+ $X2=1.315 $Y2=1.72
r99 17 39 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=2.355 $Y=0.445
+ $X2=2.355 $Y2=1.285
r100 11 13 543.532 $w=1.5e-07 $l=1.06e-06 $layer=POLY_cond $X=1.245 $Y=1.805
+ $X2=1.245 $Y2=2.865
r101 9 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.17 $Y=1.73
+ $X2=1.245 $Y2=1.805
r102 9 37 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=1.17 $Y=1.73
+ $X2=0.81 $Y2=1.73
r103 5 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.735 $Y=1.805
+ $X2=0.735 $Y2=1.64
r104 5 7 543.532 $w=1.5e-07 $l=1.06e-06 $layer=POLY_cond $X=0.735 $Y=1.805
+ $X2=0.735 $Y2=2.865
r105 1 31 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=1.475
+ $X2=0.495 $Y2=1.64
r106 1 3 510.202 $w=1.5e-07 $l=9.95e-07 $layer=POLY_cond $X=0.495 $Y=1.475
+ $X2=0.495 $Y2=0.48
.ends

.subckt PM_SKY130_FD_SC_LP__SREGSBP_1%A_75_531# 1 2 7 9 11 14 17 19 22 23 27 33
+ 36 40 42
c75 42 0 1.14682e-19 $X=0.975 $Y=0.84
c76 40 0 1.19902e-19 $X=0.52 $Y=2.85
c77 23 0 3.55192e-19 $X=2.115 $Y=2.15
c78 22 0 1.42481e-19 $X=2.115 $Y=2.15
r79 37 40 8.1743 $w=4.28e-07 $l=3.05e-07 $layer=LI1_cond $X=0.215 $Y=2.85
+ $X2=0.52 $Y2=2.85
r80 34 42 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=0.975 $Y=1.055
+ $X2=0.975 $Y2=0.84
r81 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.975
+ $Y=1.055 $X2=0.975 $Y2=1.055
r82 31 33 9.25447 $w=3.28e-07 $l=2.65e-07 $layer=LI1_cond $X=0.71 $Y=1.055
+ $X2=0.975 $Y2=1.055
r83 29 31 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=0.215 $Y=1.055
+ $X2=0.71 $Y2=1.055
r84 25 31 0.716491 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=0.71 $Y=0.89
+ $X2=0.71 $Y2=1.055
r85 25 27 14.1436 $w=3.28e-07 $l=4.05e-07 $layer=LI1_cond $X=0.71 $Y=0.89
+ $X2=0.71 $Y2=0.485
r86 23 48 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.115 $Y=2.15
+ $X2=2.115 $Y2=2.315
r87 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.115
+ $Y=2.15 $X2=2.115 $Y2=2.15
r88 20 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.3 $Y=2.15 $X2=0.215
+ $Y2=2.15
r89 20 22 63.3844 $w=3.28e-07 $l=1.815e-06 $layer=LI1_cond $X=0.3 $Y=2.15
+ $X2=2.115 $Y2=2.15
r90 19 37 6.22023 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=0.215 $Y=2.635
+ $X2=0.215 $Y2=2.85
r91 18 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.215 $Y=2.315
+ $X2=0.215 $Y2=2.15
r92 18 19 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=0.215 $Y=2.315
+ $X2=0.215 $Y2=2.635
r93 17 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.215 $Y=1.985
+ $X2=0.215 $Y2=2.15
r94 16 29 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.215 $Y=1.22
+ $X2=0.215 $Y2=1.055
r95 16 17 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=0.215 $Y=1.22
+ $X2=0.215 $Y2=1.985
r96 14 48 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=2.065 $Y=2.865
+ $X2=2.065 $Y2=2.315
r97 9 11 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.485 $Y=0.765
+ $X2=1.485 $Y2=0.445
r98 8 42 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.14 $Y=0.84
+ $X2=0.975 $Y2=0.84
r99 7 9 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.41 $Y=0.84
+ $X2=1.485 $Y2=0.765
r100 7 8 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=1.41 $Y=0.84 $X2=1.14
+ $Y2=0.84
r101 2 40 600 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_PDIFF $count=1 $X=0.375
+ $Y=2.655 $X2=0.52 $Y2=2.85
r102 1 27 182 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.27 $X2=0.71 $Y2=0.485
.ends

.subckt PM_SKY130_FD_SC_LP__SREGSBP_1%D 1 3 7 9
c37 9 0 1.14682e-19 $X=1.68 $Y=1.295
c38 3 0 1.45489e-19 $X=1.635 $Y=2.865
r39 9 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.725
+ $Y=1.29 $X2=1.725 $Y2=1.29
r40 5 12 75.7623 $w=2.98e-07 $l=4.51027e-07 $layer=POLY_cond $X=1.875 $Y=0.895
+ $X2=1.755 $Y2=1.29
r41 5 7 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=1.875 $Y=0.895
+ $X2=1.875 $Y2=0.445
r42 1 12 63.6315 $w=2.98e-07 $l=3.75233e-07 $layer=POLY_cond $X=1.635 $Y=1.61
+ $X2=1.755 $Y2=1.29
r43 1 3 643.521 $w=1.5e-07 $l=1.255e-06 $layer=POLY_cond $X=1.635 $Y=1.61
+ $X2=1.635 $Y2=2.865
.ends

.subckt PM_SKY130_FD_SC_LP__SREGSBP_1%SCD 1 3 7 9 10
c49 7 0 1.94003e-19 $X=2.745 $Y=0.445
c50 1 0 2.24855e-20 $X=2.595 $Y=2.005
r51 9 10 13.3251 $w=3.18e-07 $l=3.7e-07 $layer=LI1_cond $X=3.14 $Y=1.295
+ $X2=3.14 $Y2=1.665
r52 9 14 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.135
+ $Y=1.35 $X2=3.135 $Y2=1.35
r53 5 14 43.7503 $w=5.69e-07 $l=2.33345e-07 $layer=POLY_cond $X=2.745 $Y=1.185
+ $X2=2.91 $Y2=1.35
r54 5 7 379.447 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=2.745 $Y=1.185
+ $X2=2.745 $Y2=0.445
r55 1 14 85.2582 $w=5.69e-07 $l=7.97088e-07 $layer=POLY_cond $X=2.595 $Y=2.005
+ $X2=2.91 $Y2=1.35
r56 1 3 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=2.595 $Y=2.005
+ $X2=2.595 $Y2=2.865
.ends

.subckt PM_SKY130_FD_SC_LP__SREGSBP_1%A_342_531# 1 2 3 4 15 17 19 20 21 23 26 28
+ 29 31 32 33 35 38 39 43 45 46 48 49 50 51 57 64 71
c202 71 0 1.41824e-19 $X=5.955 $Y=0.737
c203 51 0 1.96333e-19 $X=2.305 $Y=0.555
c204 50 0 1.92092e-20 $X=5.375 $Y=0.555
c205 49 0 1.60209e-19 $X=2.715 $Y=2.415
c206 48 0 7.16051e-20 $X=5.955 $Y=2.085
c207 45 0 6.03758e-20 $X=5.87 $Y=2.17
c208 35 0 1.94983e-19 $X=2.715 $Y=2.165
r209 70 71 4.72401 $w=5.93e-07 $l=2.35e-07 $layer=LI1_cond $X=5.72 $Y=0.737
+ $X2=5.955 $Y2=0.737
r210 64 66 9.85908 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=2.14 $Y=0.47
+ $X2=2.14 $Y2=0.675
r211 58 70 4.02043 $w=5.93e-07 $l=2e-07 $layer=LI1_cond $X=5.52 $Y=0.737
+ $X2=5.72 $Y2=0.737
r212 57 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0.555
+ $X2=5.52 $Y2=0.555
r213 53 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0.555
+ $X2=2.16 $Y2=0.555
r214 51 53 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.305 $Y=0.555
+ $X2=2.16 $Y2=0.555
r215 50 57 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.375 $Y=0.555
+ $X2=5.52 $Y2=0.555
r216 50 51 3.7995 $w=1.4e-07 $l=3.07e-06 $layer=MET1_cond $X=5.375 $Y=0.555
+ $X2=2.305 $Y2=0.555
r217 47 71 8.26286 $w=1.7e-07 $l=2.98e-07 $layer=LI1_cond $X=5.955 $Y=1.035
+ $X2=5.955 $Y2=0.737
r218 47 48 68.5027 $w=1.68e-07 $l=1.05e-06 $layer=LI1_cond $X=5.955 $Y=1.035
+ $X2=5.955 $Y2=2.085
r219 45 48 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.87 $Y=2.17
+ $X2=5.955 $Y2=2.085
r220 45 46 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=5.87 $Y=2.17
+ $X2=5.49 $Y2=2.17
r221 41 46 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=5.365 $Y=2.255
+ $X2=5.49 $Y2=2.17
r222 41 43 12.4464 $w=2.48e-07 $l=2.7e-07 $layer=LI1_cond $X=5.365 $Y=2.255
+ $X2=5.365 $Y2=2.525
r223 39 60 17.7787 $w=2.44e-07 $l=9e-08 $layer=POLY_cond $X=3.195 $Y=2.33
+ $X2=3.105 $Y2=2.33
r224 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.195
+ $Y=2.33 $X2=3.195 $Y2=2.33
r225 36 49 3.70735 $w=2.5e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.8 $Y=2.33
+ $X2=2.715 $Y2=2.415
r226 36 38 13.7944 $w=3.28e-07 $l=3.95e-07 $layer=LI1_cond $X=2.8 $Y=2.33
+ $X2=3.195 $Y2=2.33
r227 35 49 2.76166 $w=1.7e-07 $l=2.5e-07 $layer=LI1_cond $X=2.715 $Y=2.165
+ $X2=2.715 $Y2=2.415
r228 34 35 74.3743 $w=1.68e-07 $l=1.14e-06 $layer=LI1_cond $X=2.715 $Y=1.025
+ $X2=2.715 $Y2=2.165
r229 32 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.63 $Y=0.94
+ $X2=2.715 $Y2=1.025
r230 32 33 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=2.63 $Y=0.94
+ $X2=2.305 $Y2=0.94
r231 31 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.22 $Y=0.855
+ $X2=2.305 $Y2=0.94
r232 31 66 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=2.22 $Y=0.855
+ $X2=2.22 $Y2=0.675
r233 28 49 3.70735 $w=2.5e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.63 $Y=2.58
+ $X2=2.715 $Y2=2.415
r234 28 29 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=2.63 $Y=2.58
+ $X2=2.015 $Y2=2.58
r235 24 29 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.85 $Y=2.665
+ $X2=2.015 $Y2=2.58
r236 24 26 6.46067 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=1.85 $Y=2.665
+ $X2=1.85 $Y2=2.85
r237 23 39 77.041 $w=2.44e-07 $l=4.65242e-07 $layer=POLY_cond $X=3.585 $Y=2.165
+ $X2=3.195 $Y2=2.33
r238 22 23 640.957 $w=1.5e-07 $l=1.25e-06 $layer=POLY_cond $X=3.585 $Y=0.915
+ $X2=3.585 $Y2=2.165
r239 20 22 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.51 $Y=0.84
+ $X2=3.585 $Y2=0.915
r240 20 21 133.319 $w=1.5e-07 $l=2.6e-07 $layer=POLY_cond $X=3.51 $Y=0.84
+ $X2=3.25 $Y2=0.84
r241 17 21 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.175 $Y=0.765
+ $X2=3.25 $Y2=0.84
r242 17 19 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=3.175 $Y=0.765
+ $X2=3.175 $Y2=0.445
r243 13 60 14.1583 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.105 $Y=2.495
+ $X2=3.105 $Y2=2.33
r244 13 15 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=3.105 $Y=2.495
+ $X2=3.105 $Y2=2.865
r245 4 43 600 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=1 $X=5.26
+ $Y=2.315 $X2=5.405 $Y2=2.525
r246 3 26 600 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_PDIFF $count=1 $X=1.71
+ $Y=2.655 $X2=1.85 $Y2=2.85
r247 2 70 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=5.575
+ $Y=0.595 $X2=5.72 $Y2=0.805
r248 1 64 182 $w=1.7e-07 $l=3.1603e-07 $layer=licon1_NDIFF $count=1 $X=1.95
+ $Y=0.235 $X2=2.14 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_LP__SREGSBP_1%CLK 1 3 5 7 8
c44 5 0 1.72328e-20 $X=4.205 $Y=1.185
c45 1 0 1.92092e-20 $X=4.165 $Y=1.515
r46 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.035
+ $Y=1.35 $X2=4.035 $Y2=1.35
r47 5 11 39.3587 $w=3.88e-07 $l=2.20624e-07 $layer=POLY_cond $X=4.205 $Y=1.185
+ $X2=4.075 $Y2=1.35
r48 5 7 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=4.205 $Y=1.185
+ $X2=4.205 $Y2=0.655
r49 1 11 39.3587 $w=3.88e-07 $l=2.05122e-07 $layer=POLY_cond $X=4.165 $Y=1.515
+ $X2=4.075 $Y2=1.35
r50 1 3 461.489 $w=1.5e-07 $l=9e-07 $layer=POLY_cond $X=4.165 $Y=1.515 $X2=4.165
+ $Y2=2.415
.ends

.subckt PM_SKY130_FD_SC_LP__SREGSBP_1%A_934_357# 1 2 9 11 15 19 20 24 29 35 38
+ 40 41 42 43 46 49 50 52 59 61
c178 59 0 1.95779e-19 $X=9.53 $Y=1.54
c179 41 0 1.72328e-20 $X=5.022 $Y=1.045
c180 11 0 2.06024e-19 $X=6.22 $Y=1.65
r181 59 62 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=9.53 $Y=1.54 $X2=9.53
+ $Y2=1.63
r182 59 61 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=9.53 $Y=1.54
+ $X2=9.53 $Y2=1.375
r183 55 57 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.555 $Y=1.74
+ $X2=5.555 $Y2=1.905
r184 52 55 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=5.555 $Y=1.65
+ $X2=5.555 $Y2=1.74
r185 50 59 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.53
+ $Y=1.54 $X2=9.53 $Y2=1.54
r186 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=1.665
+ $X2=9.36 $Y2=1.665
r187 46 55 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.555
+ $Y=1.74 $X2=5.555 $Y2=1.74
r188 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=1.665
+ $X2=5.52 $Y2=1.665
r189 43 45 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.665 $Y=1.665
+ $X2=5.52 $Y2=1.665
r190 42 49 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=9.215 $Y=1.665
+ $X2=9.36 $Y2=1.665
r191 42 43 4.39356 $w=1.4e-07 $l=3.55e-06 $layer=MET1_cond $X=9.215 $Y=1.665
+ $X2=5.665 $Y2=1.665
r192 39 46 10.3882 $w=3.53e-07 $l=3.2e-07 $layer=LI1_cond $X=5.2 $Y=1.727
+ $X2=5.52 $Y2=1.727
r193 39 40 0.0561152 $w=3.55e-07 $l=4.78983e-07 $layer=LI1_cond $X=5.2 $Y=1.727
+ $X2=4.725 $Y2=1.735
r194 38 40 7.11569 $w=2.37e-07 $l=4.7355e-07 $layer=LI1_cond $X=5.115 $Y=1.55
+ $X2=4.725 $Y2=1.735
r195 38 41 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=5.115 $Y=1.55
+ $X2=5.115 $Y2=1.045
r196 33 41 8.88861 $w=3.53e-07 $l=1.77e-07 $layer=LI1_cond $X=5.022 $Y=0.868
+ $X2=5.022 $Y2=1.045
r197 33 35 14.2189 $w=3.53e-07 $l=4.38e-07 $layer=LI1_cond $X=5.022 $Y=0.868
+ $X2=5.022 $Y2=0.43
r198 29 31 36.6515 $w=3.03e-07 $l=9.7e-07 $layer=LI1_cond $X=4.877 $Y=1.93
+ $X2=4.877 $Y2=2.9
r199 27 40 7.11569 $w=2.37e-07 $l=2.33966e-07 $layer=LI1_cond $X=4.877 $Y=1.905
+ $X2=4.725 $Y2=1.735
r200 27 29 0.944625 $w=3.03e-07 $l=2.5e-08 $layer=LI1_cond $X=4.877 $Y=1.905
+ $X2=4.877 $Y2=1.93
r201 22 24 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=10.135 $Y=1.705
+ $X2=10.135 $Y2=2.465
r202 21 62 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.695 $Y=1.63
+ $X2=9.53 $Y2=1.63
r203 20 22 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=10.06 $Y=1.63
+ $X2=10.135 $Y2=1.705
r204 20 21 187.16 $w=1.5e-07 $l=3.65e-07 $layer=POLY_cond $X=10.06 $Y=1.63
+ $X2=9.695 $Y2=1.63
r205 19 61 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=9.44 $Y=0.945
+ $X2=9.44 $Y2=1.375
r206 13 26 11.9802 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=6.52 $Y=1.395
+ $X2=6.52 $Y2=1.545
r207 13 15 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=6.52 $Y=1.395
+ $X2=6.52 $Y2=0.805
r208 12 52 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.72 $Y=1.65
+ $X2=5.555 $Y2=1.65
r209 11 26 70.2291 $w=2.22e-07 $l=3.48569e-07 $layer=POLY_cond $X=6.22 $Y=1.65
+ $X2=6.52 $Y2=1.545
r210 11 12 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=6.22 $Y=1.65 $X2=5.72
+ $Y2=1.65
r211 9 57 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=5.62 $Y=2.525
+ $X2=5.62 $Y2=1.905
r212 2 31 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=4.67
+ $Y=1.785 $X2=4.81 $Y2=2.9
r213 2 29 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=4.67
+ $Y=1.785 $X2=4.81 $Y2=1.93
r214 1 35 91 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_NDIFF $count=2 $X=4.87
+ $Y=0.235 $X2=5.01 $Y2=0.43
.ends

.subckt PM_SKY130_FD_SC_LP__SREGSBP_1%A_1273_393# 1 2 3 12 16 18 20 23 26 27 28
+ 29 32 34 39 44 46 50 52 53 57 62
c142 46 0 2.41575e-19 $X=7.215 $Y=2.05
c143 12 0 6.03758e-20 $X=6.44 $Y=2.525
r144 62 63 4.56151 $w=3.17e-07 $l=3e-08 $layer=POLY_cond $X=9.05 $Y=1.54
+ $X2=9.08 $Y2=1.54
r145 53 55 6.68417 $w=2.48e-07 $l=1.45e-07 $layer=LI1_cond $X=8.345 $Y=2.415
+ $X2=8.345 $Y2=2.56
r146 48 50 5.88393 $w=6.18e-07 $l=3.05e-07 $layer=LI1_cond $X=8.035 $Y=0.885
+ $X2=8.34 $Y2=0.885
r147 44 60 24.6477 $w=2.64e-07 $l=1.35e-07 $layer=POLY_cond $X=6.745 $Y=1.95
+ $X2=6.88 $Y2=1.95
r148 43 46 21.1587 $w=2.71e-07 $l=4.7e-07 $layer=LI1_cond $X=6.745 $Y=1.95
+ $X2=7.215 $Y2=1.95
r149 43 44 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.745
+ $Y=1.95 $X2=6.745 $Y2=1.95
r150 40 62 22.8076 $w=3.17e-07 $l=1.5e-07 $layer=POLY_cond $X=8.9 $Y=1.54
+ $X2=9.05 $Y2=1.54
r151 39 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.9
+ $Y=1.54 $X2=8.9 $Y2=1.54
r152 37 57 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.425 $Y=1.54
+ $X2=8.34 $Y2=1.54
r153 37 39 16.5882 $w=3.28e-07 $l=4.75e-07 $layer=LI1_cond $X=8.425 $Y=1.54
+ $X2=8.9 $Y2=1.54
r154 35 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.34 $Y=1.705
+ $X2=8.34 $Y2=1.54
r155 35 52 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=8.34 $Y=1.705
+ $X2=8.34 $Y2=1.885
r156 34 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.34 $Y=1.375
+ $X2=8.34 $Y2=1.54
r157 33 50 8.52869 $w=1.7e-07 $l=3.1e-07 $layer=LI1_cond $X=8.34 $Y=1.195
+ $X2=8.34 $Y2=0.885
r158 33 34 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=8.34 $Y=1.195
+ $X2=8.34 $Y2=1.375
r159 30 53 3.91831 $w=2.48e-07 $l=8.5e-08 $layer=LI1_cond $X=8.345 $Y=2.33
+ $X2=8.345 $Y2=2.415
r160 30 32 12.9074 $w=2.48e-07 $l=2.8e-07 $layer=LI1_cond $X=8.345 $Y=2.33
+ $X2=8.345 $Y2=2.05
r161 29 52 6.39536 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=8.345 $Y=2.01
+ $X2=8.345 $Y2=1.885
r162 29 32 1.84391 $w=2.48e-07 $l=4e-08 $layer=LI1_cond $X=8.345 $Y=2.01
+ $X2=8.345 $Y2=2.05
r163 27 53 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.22 $Y=2.415
+ $X2=8.345 $Y2=2.415
r164 27 28 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=8.22 $Y=2.415
+ $X2=7.38 $Y2=2.415
r165 26 28 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=7.215 $Y=2.33
+ $X2=7.38 $Y2=2.415
r166 26 46 7.50834 $w=3.28e-07 $l=2.15e-07 $layer=LI1_cond $X=7.215 $Y=2.33
+ $X2=7.215 $Y2=2.115
r167 21 63 20.269 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.08 $Y=1.705
+ $X2=9.08 $Y2=1.54
r168 21 23 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=9.08 $Y=1.705
+ $X2=9.08 $Y2=2.285
r169 18 62 20.269 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.05 $Y=1.375
+ $X2=9.05 $Y2=1.54
r170 18 20 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=9.05 $Y=1.375
+ $X2=9.05 $Y2=0.945
r171 14 60 15.9823 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.88 $Y=1.785
+ $X2=6.88 $Y2=1.95
r172 14 16 502.511 $w=1.5e-07 $l=9.8e-07 $layer=POLY_cond $X=6.88 $Y=1.785
+ $X2=6.88 $Y2=0.805
r173 10 44 55.6856 $w=2.64e-07 $l=3.78616e-07 $layer=POLY_cond $X=6.44 $Y=2.115
+ $X2=6.745 $Y2=1.95
r174 10 12 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=6.44 $Y=2.115
+ $X2=6.44 $Y2=2.525
r175 3 55 600 $w=1.7e-07 $l=7.61791e-07 $layer=licon1_PDIFF $count=1 $X=8.165
+ $Y=1.865 $X2=8.305 $Y2=2.56
r176 3 32 600 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_PDIFF $count=1 $X=8.165
+ $Y=1.865 $X2=8.305 $Y2=2.05
r177 2 46 300 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_PDIFF $count=2 $X=7.07
+ $Y=1.865 $X2=7.215 $Y2=2.05
r178 1 48 182 $w=1.7e-07 $l=3.53129e-07 $layer=licon1_NDIFF $count=1 $X=7.895
+ $Y=0.595 $X2=8.035 $Y2=0.885
.ends

.subckt PM_SKY130_FD_SC_LP__SREGSBP_1%A_1139_463# 1 2 9 13 15 21 24 25 27 28 32
r89 32 36 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.34 $Y=1.54
+ $X2=7.34 $Y2=1.705
r90 32 35 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.34 $Y=1.54
+ $X2=7.34 $Y2=1.375
r91 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.34
+ $Y=1.54 $X2=7.34 $Y2=1.54
r92 28 31 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=7.34 $Y=1.46 $X2=7.34
+ $Y2=1.54
r93 26 27 2.11342 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.47 $Y=1.46
+ $X2=6.345 $Y2=1.46
r94 25 28 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.175 $Y=1.46
+ $X2=7.34 $Y2=1.46
r95 25 26 45.9947 $w=1.68e-07 $l=7.05e-07 $layer=LI1_cond $X=7.175 $Y=1.46
+ $X2=6.47 $Y2=1.46
r96 23 27 4.3182 $w=2.1e-07 $l=1.03078e-07 $layer=LI1_cond $X=6.305 $Y=1.545
+ $X2=6.345 $Y2=1.46
r97 23 24 58.0642 $w=1.68e-07 $l=8.9e-07 $layer=LI1_cond $X=6.305 $Y=1.545
+ $X2=6.305 $Y2=2.435
r98 19 27 4.3182 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=6.345 $Y=1.375
+ $X2=6.345 $Y2=1.46
r99 19 21 26.2757 $w=2.48e-07 $l=5.7e-07 $layer=LI1_cond $X=6.345 $Y=1.375
+ $X2=6.345 $Y2=0.805
r100 15 24 7.68211 $w=3.2e-07 $l=1.9799e-07 $layer=LI1_cond $X=6.22 $Y=2.595
+ $X2=6.305 $Y2=2.435
r101 15 17 13.8653 $w=3.18e-07 $l=3.85e-07 $layer=LI1_cond $X=6.22 $Y=2.595
+ $X2=5.835 $Y2=2.595
r102 13 36 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=7.43 $Y=2.285
+ $X2=7.43 $Y2=1.705
r103 9 35 235.872 $w=1.5e-07 $l=4.6e-07 $layer=POLY_cond $X=7.43 $Y=0.915
+ $X2=7.43 $Y2=1.375
r104 2 17 600 $w=1.7e-07 $l=3.01993e-07 $layer=licon1_PDIFF $count=1 $X=5.695
+ $Y=2.315 $X2=5.835 $Y2=2.555
r105 1 21 182 $w=1.7e-07 $l=3.85973e-07 $layer=licon1_NDIFF $count=1 $X=6.01
+ $Y=0.595 $X2=6.305 $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_LP__SREGSBP_1%ASYNC 3 7 9 11 16 20 24 25 29 33 34 37 39
+ 44 47 55
c134 55 0 7.80799e-20 $X=11.395 $Y=1.977
c135 47 0 1.61879e-19 $X=11.697 $Y=1.765
c136 25 0 1.44748e-19 $X=11.67 $Y=1.93
c137 7 0 1.77375e-19 $X=8.09 $Y=2.285
r138 52 55 4.16805 $w=3.43e-07 $l=1.15e-07 $layer=LI1_cond $X=11.28 $Y=1.977
+ $X2=11.395 $Y2=1.977
r139 39 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.28 $Y=2.035
+ $X2=11.28 $Y2=2.035
r140 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=2.035
+ $X2=7.92 $Y2=2.035
r141 34 36 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.065 $Y=2.035
+ $X2=7.92 $Y2=2.035
r142 33 39 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=11.135 $Y=2.035
+ $X2=11.28 $Y2=2.035
r143 33 34 3.7995 $w=1.4e-07 $l=3.07e-06 $layer=MET1_cond $X=11.135 $Y=2.035
+ $X2=8.065 $Y2=2.035
r144 32 37 13.114 $w=2.88e-07 $l=3.3e-07 $layer=LI1_cond $X=7.89 $Y=1.705
+ $X2=7.89 $Y2=2.035
r145 30 44 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=7.91 $Y=1.54
+ $X2=8.09 $Y2=1.54
r146 30 41 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=7.91 $Y=1.54 $X2=7.82
+ $Y2=1.54
r147 29 32 5.96091 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=7.91 $Y=1.54
+ $X2=7.91 $Y2=1.705
r148 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.91
+ $Y=1.54 $X2=7.91 $Y2=1.54
r149 25 48 45.3519 $w=3.85e-07 $l=1.65e-07 $layer=POLY_cond $X=11.697 $Y=1.93
+ $X2=11.697 $Y2=2.095
r150 25 47 45.3519 $w=3.85e-07 $l=1.65e-07 $layer=POLY_cond $X=11.697 $Y=1.93
+ $X2=11.697 $Y2=1.765
r151 24 55 10.9283 $w=2.88e-07 $l=2.75e-07 $layer=LI1_cond $X=11.67 $Y=1.95
+ $X2=11.395 $Y2=1.95
r152 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.67
+ $Y=1.93 $X2=11.67 $Y2=1.93
r153 18 20 94.8617 $w=1.5e-07 $l=1.85e-07 $layer=POLY_cond $X=11.395 $Y=1.06
+ $X2=11.58 $Y2=1.06
r154 16 48 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=11.58 $Y=2.675
+ $X2=11.58 $Y2=2.095
r155 12 20 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=11.58 $Y=1.135
+ $X2=11.58 $Y2=1.06
r156 12 47 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=11.58 $Y=1.135
+ $X2=11.58 $Y2=1.765
r157 9 18 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=11.395 $Y=0.985
+ $X2=11.395 $Y2=1.06
r158 9 11 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=11.395 $Y=0.985
+ $X2=11.395 $Y2=0.555
r159 5 44 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.09 $Y=1.705
+ $X2=8.09 $Y2=1.54
r160 5 7 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=8.09 $Y=1.705
+ $X2=8.09 $Y2=2.285
r161 1 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.82 $Y=1.375
+ $X2=7.82 $Y2=1.54
r162 1 3 235.872 $w=1.5e-07 $l=4.6e-07 $layer=POLY_cond $X=7.82 $Y=1.375
+ $X2=7.82 $Y2=0.915
.ends

.subckt PM_SKY130_FD_SC_LP__SREGSBP_1%A_761_357# 1 2 9 11 13 15 16 18 19 23 26
+ 28 29 30 34 38 40 43 49 51 52 53 54 56 58 62 70
c182 15 0 7.16051e-20 $X=5.105 $Y=3.075
r183 69 70 32.7208 $w=3.7e-07 $l=7.5e-08 $layer=POLY_cond $X=5.105 $Y=1.37
+ $X2=5.18 $Y2=1.37
r184 68 69 48.3468 $w=3.7e-07 $l=3.1e-07 $layer=POLY_cond $X=4.795 $Y=1.37
+ $X2=5.105 $Y2=1.37
r185 63 68 17.1553 $w=3.7e-07 $l=1.1e-07 $layer=POLY_cond $X=4.685 $Y=1.37
+ $X2=4.795 $Y2=1.37
r186 63 65 14.0362 $w=3.7e-07 $l=9e-08 $layer=POLY_cond $X=4.685 $Y=1.37
+ $X2=4.595 $Y2=1.37
r187 62 63 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.685
+ $Y=1.39 $X2=4.685 $Y2=1.39
r188 59 62 7.85757 $w=3.28e-07 $l=2.25e-07 $layer=LI1_cond $X=4.46 $Y=1.39
+ $X2=4.685 $Y2=1.39
r189 57 59 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.46 $Y=1.555
+ $X2=4.46 $Y2=1.39
r190 57 58 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=4.46 $Y=1.555
+ $X2=4.46 $Y2=1.695
r191 56 59 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.46 $Y=1.225
+ $X2=4.46 $Y2=1.39
r192 55 56 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=4.46 $Y=1 $X2=4.46
+ $Y2=1.225
r193 53 55 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.375 $Y=0.915
+ $X2=4.46 $Y2=1
r194 53 54 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=4.375 $Y=0.915
+ $X2=4.155 $Y2=0.915
r195 51 58 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.375 $Y=1.78
+ $X2=4.46 $Y2=1.695
r196 51 52 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=4.375 $Y=1.78
+ $X2=4.035 $Y2=1.78
r197 47 54 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=4.03 $Y=0.83
+ $X2=4.155 $Y2=0.915
r198 47 49 18.4391 $w=2.48e-07 $l=4e-07 $layer=LI1_cond $X=4.03 $Y=0.83 $X2=4.03
+ $Y2=0.43
r199 43 45 63.2834 $w=1.68e-07 $l=9.7e-07 $layer=LI1_cond $X=3.95 $Y=1.93
+ $X2=3.95 $Y2=2.9
r200 41 52 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.95 $Y=1.865
+ $X2=4.035 $Y2=1.78
r201 41 43 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=3.95 $Y=1.865
+ $X2=3.95 $Y2=1.93
r202 36 38 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=10.1 $Y=0.255
+ $X2=10.1 $Y2=0.665
r203 32 34 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=9.59 $Y=3.075
+ $X2=9.59 $Y2=2.465
r204 31 40 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.125 $Y=3.15
+ $X2=6.05 $Y2=3.15
r205 30 32 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.515 $Y=3.15
+ $X2=9.59 $Y2=3.075
r206 30 31 1738.28 $w=1.5e-07 $l=3.39e-06 $layer=POLY_cond $X=9.515 $Y=3.15
+ $X2=6.125 $Y2=3.15
r207 28 36 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=10.025 $Y=0.18
+ $X2=10.1 $Y2=0.255
r208 28 29 2058.76 $w=1.5e-07 $l=4.015e-06 $layer=POLY_cond $X=10.025 $Y=0.18
+ $X2=6.01 $Y2=0.18
r209 24 40 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.05 $Y=3.075
+ $X2=6.05 $Y2=3.15
r210 24 26 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=6.05 $Y=3.075
+ $X2=6.05 $Y2=2.525
r211 21 23 194.851 $w=1.5e-07 $l=3.8e-07 $layer=POLY_cond $X=5.935 $Y=1.185
+ $X2=5.935 $Y2=0.805
r212 20 29 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.935 $Y=0.255
+ $X2=6.01 $Y2=0.18
r213 20 23 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=5.935 $Y=0.255
+ $X2=5.935 $Y2=0.805
r214 18 40 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.975 $Y=3.15
+ $X2=6.05 $Y2=3.15
r215 18 19 407.649 $w=1.5e-07 $l=7.95e-07 $layer=POLY_cond $X=5.975 $Y=3.15
+ $X2=5.18 $Y2=3.15
r216 16 21 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.86 $Y=1.26
+ $X2=5.935 $Y2=1.185
r217 16 70 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=5.86 $Y=1.26
+ $X2=5.18 $Y2=1.26
r218 15 19 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.105 $Y=3.075
+ $X2=5.18 $Y2=3.15
r219 14 69 23.9667 $w=1.5e-07 $l=1.85e-07 $layer=POLY_cond $X=5.105 $Y=1.555
+ $X2=5.105 $Y2=1.37
r220 14 15 779.404 $w=1.5e-07 $l=1.52e-06 $layer=POLY_cond $X=5.105 $Y=1.555
+ $X2=5.105 $Y2=3.075
r221 11 68 23.9667 $w=1.5e-07 $l=1.85e-07 $layer=POLY_cond $X=4.795 $Y=1.185
+ $X2=4.795 $Y2=1.37
r222 11 13 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=4.795 $Y=1.185
+ $X2=4.795 $Y2=0.655
r223 7 65 23.9667 $w=1.5e-07 $l=1.85e-07 $layer=POLY_cond $X=4.595 $Y=1.555
+ $X2=4.595 $Y2=1.37
r224 7 9 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=4.595 $Y=1.555
+ $X2=4.595 $Y2=2.415
r225 2 45 400 $w=1.7e-07 $l=1.18528e-06 $layer=licon1_PDIFF $count=1 $X=3.805
+ $Y=1.785 $X2=3.95 $Y2=2.9
r226 2 43 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=3.805
+ $Y=1.785 $X2=3.95 $Y2=1.93
r227 1 49 91 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_NDIFF $count=2 $X=3.845
+ $Y=0.235 $X2=3.99 $Y2=0.43
.ends

.subckt PM_SKY130_FD_SC_LP__SREGSBP_1%A_2083_65# 1 2 9 14 18 22 24 28 32 34 35
+ 36 40 41 42 43 44 49 51 54 55 56 59 60 61 68 70
c167 61 0 1.44748e-19 $X=12.265 $Y=1.54
c168 28 0 1.66705e-19 $X=13.345 $Y=2.465
c169 14 0 7.80799e-20 $X=10.525 $Y=2.465
r170 70 71 32.1566 $w=3.6e-07 $l=7.5e-08 $layer=POLY_cond $X=12.28 $Y=1.53
+ $X2=12.28 $Y2=1.455
r171 65 73 46.5827 $w=3.6e-07 $l=1.65e-07 $layer=POLY_cond $X=12.28 $Y=1.62
+ $X2=12.28 $Y2=1.785
r172 65 70 14.4261 $w=3.6e-07 $l=9e-08 $layer=POLY_cond $X=12.28 $Y=1.62
+ $X2=12.28 $Y2=1.53
r173 64 65 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=12.265
+ $Y=1.62 $X2=12.265 $Y2=1.62
r174 61 64 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=12.265 $Y=1.54
+ $X2=12.265 $Y2=1.62
r175 55 69 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=10.585 $Y=1.93
+ $X2=10.585 $Y2=2.095
r176 55 68 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=10.585 $Y=1.93
+ $X2=10.585 $Y2=1.765
r177 54 57 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=10.585 $Y=1.93
+ $X2=10.585 $Y2=2.095
r178 54 56 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=10.585 $Y=1.93
+ $X2=10.585 $Y2=1.765
r179 54 55 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.585
+ $Y=1.93 $X2=10.585 $Y2=1.93
r180 52 60 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.775 $Y=1.54
+ $X2=11.61 $Y2=1.54
r181 51 61 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.1 $Y=1.54
+ $X2=12.265 $Y2=1.54
r182 51 52 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=12.1 $Y=1.54
+ $X2=11.775 $Y2=1.54
r183 47 60 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=11.61 $Y=1.455
+ $X2=11.61 $Y2=1.54
r184 47 49 30.5572 $w=3.28e-07 $l=8.75e-07 $layer=LI1_cond $X=11.61 $Y=1.455
+ $X2=11.61 $Y2=0.58
r185 43 59 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.2 $Y=2.415
+ $X2=11.365 $Y2=2.415
r186 43 44 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=11.2 $Y=2.415
+ $X2=10.75 $Y2=2.415
r187 41 60 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.445 $Y=1.54
+ $X2=11.61 $Y2=1.54
r188 41 42 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=11.445 $Y=1.54
+ $X2=10.75 $Y2=1.54
r189 40 44 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.665 $Y=2.33
+ $X2=10.75 $Y2=2.415
r190 40 57 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=10.665 $Y=2.33
+ $X2=10.665 $Y2=2.095
r191 37 42 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.665 $Y=1.625
+ $X2=10.75 $Y2=1.54
r192 37 56 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=10.665 $Y=1.625
+ $X2=10.665 $Y2=1.765
r193 35 68 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=10.495 $Y=1.135
+ $X2=10.495 $Y2=1.765
r194 34 35 71.7618 $w=1.55e-07 $l=1.5e-07 $layer=POLY_cond $X=10.492 $Y=0.985
+ $X2=10.492 $Y2=1.135
r195 30 36 20.4101 $w=1.5e-07 $l=8.21584e-08 $layer=POLY_cond $X=13.375 $Y=1.455
+ $X2=13.36 $Y2=1.53
r196 30 32 384.574 $w=1.5e-07 $l=7.5e-07 $layer=POLY_cond $X=13.375 $Y=1.455
+ $X2=13.375 $Y2=0.705
r197 26 36 20.4101 $w=1.5e-07 $l=8.21584e-08 $layer=POLY_cond $X=13.345 $Y=1.605
+ $X2=13.36 $Y2=1.53
r198 26 28 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=13.345 $Y=1.605
+ $X2=13.345 $Y2=2.465
r199 25 70 23.3057 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=12.46 $Y=1.53
+ $X2=12.28 $Y2=1.53
r200 24 36 5.30422 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=13.27 $Y=1.53
+ $X2=13.36 $Y2=1.53
r201 24 25 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=13.27 $Y=1.53
+ $X2=12.46 $Y2=1.53
r202 22 71 492.255 $w=1.5e-07 $l=9.6e-07 $layer=POLY_cond $X=12.385 $Y=0.495
+ $X2=12.385 $Y2=1.455
r203 18 73 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=12.205 $Y=2.575
+ $X2=12.205 $Y2=1.785
r204 14 69 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=10.525 $Y=2.465
+ $X2=10.525 $Y2=2.095
r205 9 34 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=10.49 $Y=0.665
+ $X2=10.49 $Y2=0.985
r206 2 59 300 $w=1.7e-07 $l=3.01993e-07 $layer=licon1_PDIFF $count=2 $X=11.225
+ $Y=2.255 $X2=11.365 $Y2=2.495
r207 1 49 182 $w=1.7e-07 $l=4.09054e-07 $layer=licon1_NDIFF $count=1 $X=11.47
+ $Y=0.235 $X2=11.61 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_LP__SREGSBP_1%A_1903_125# 1 2 9 12 15 17 18 21 30 32 33
+ 36 37 38
c92 36 0 1.61879e-19 $X=10.945 $Y=1.15
c93 32 0 1.95779e-19 $X=9.805 $Y=2.19
c94 30 0 4.80826e-20 $X=9.77 $Y=1.03
r95 36 38 7.45374 $w=2.88e-07 $l=1.65e-07 $layer=LI1_cond $X=10.945 $Y=1.13
+ $X2=10.78 $Y2=1.13
r96 36 37 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.945
+ $Y=1.15 $X2=10.945 $Y2=1.15
r97 32 33 8.6688 $w=4.03e-07 $l=1.65e-07 $layer=LI1_cond $X=9.842 $Y=2.19
+ $X2=9.842 $Y2=2.025
r98 28 30 2.71504 $w=2.1e-07 $l=2.2e-07 $layer=LI1_cond $X=10.045 $Y=1.09
+ $X2=9.825 $Y2=1.09
r99 28 38 38.8182 $w=2.08e-07 $l=7.35e-07 $layer=LI1_cond $X=10.045 $Y=1.09
+ $X2=10.78 $Y2=1.09
r100 25 30 3.74844 $w=3.05e-07 $l=1.8e-07 $layer=LI1_cond $X=9.96 $Y=1.195
+ $X2=9.825 $Y2=1.09
r101 25 33 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=9.96 $Y=1.195
+ $X2=9.96 $Y2=2.025
r102 19 30 3.74844 $w=3.05e-07 $l=1.05e-07 $layer=LI1_cond $X=9.825 $Y=0.985
+ $X2=9.825 $Y2=1.09
r103 19 21 10.0839 $w=4.38e-07 $l=3.85e-07 $layer=LI1_cond $X=9.825 $Y=0.985
+ $X2=9.825 $Y2=0.6
r104 17 37 39.3438 $w=3.3e-07 $l=2.25e-07 $layer=POLY_cond $X=10.945 $Y=1.375
+ $X2=10.945 $Y2=1.15
r105 17 18 43.5886 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=11.002 $Y=1.375
+ $X2=11.002 $Y2=1.525
r106 15 37 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=10.945 $Y=0.985
+ $X2=10.945 $Y2=1.15
r107 12 18 589.681 $w=1.5e-07 $l=1.15e-06 $layer=POLY_cond $X=11.15 $Y=2.675
+ $X2=11.15 $Y2=1.525
r108 9 15 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=11.035 $Y=0.555
+ $X2=11.035 $Y2=0.985
r109 2 32 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=9.665
+ $Y=2.045 $X2=9.805 $Y2=2.19
r110 1 30 182 $w=1.7e-07 $l=5.17011e-07 $layer=licon1_NDIFF $count=1 $X=9.515
+ $Y=0.625 $X2=9.77 $Y2=1.03
r111 1 21 182 $w=1.7e-07 $l=2.67208e-07 $layer=licon1_NDIFF $count=1 $X=9.515
+ $Y=0.625 $X2=9.77 $Y2=0.6
.ends

.subckt PM_SKY130_FD_SC_LP__SREGSBP_1%A_2456_451# 1 2 9 13 18 19 22 24 27 29 35
+ 36
r98 36 40 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=13.825 $Y=1.49
+ $X2=13.825 $Y2=1.655
r99 36 39 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=13.825 $Y=1.49
+ $X2=13.825 $Y2=1.325
r100 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=13.825
+ $Y=1.49 $X2=13.825 $Y2=1.49
r101 32 35 6.46067 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=13.64 $Y=1.49
+ $X2=13.825 $Y2=1.49
r102 29 31 10.6507 $w=3.43e-07 $l=2.3e-07 $layer=LI1_cond $X=12.607 $Y=0.495
+ $X2=12.607 $Y2=0.725
r103 26 27 5.14764 $w=2.58e-07 $l=8.5e-08 $layer=LI1_cond $X=12.695 $Y=2.365
+ $X2=12.78 $Y2=2.365
r104 24 26 12.1893 $w=2.58e-07 $l=2.75e-07 $layer=LI1_cond $X=12.42 $Y=2.365
+ $X2=12.695 $Y2=2.365
r105 21 32 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.64 $Y=1.655
+ $X2=13.64 $Y2=1.49
r106 21 22 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=13.64 $Y=1.655
+ $X2=13.64 $Y2=2.325
r107 19 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=13.555 $Y=2.41
+ $X2=13.64 $Y2=2.325
r108 19 27 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=13.555 $Y=2.41
+ $X2=12.78 $Y2=2.41
r109 18 26 3.22376 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=12.695 $Y=2.235
+ $X2=12.695 $Y2=2.365
r110 18 31 98.5134 $w=1.68e-07 $l=1.51e-06 $layer=LI1_cond $X=12.695 $Y=2.235
+ $X2=12.695 $Y2=0.725
r111 13 39 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=13.885 $Y=0.705
+ $X2=13.885 $Y2=1.325
r112 9 40 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=13.855 $Y=2.465
+ $X2=13.855 $Y2=1.655
r113 2 24 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=12.28
+ $Y=2.255 $X2=12.42 $Y2=2.4
r114 1 29 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=12.46
+ $Y=0.285 $X2=12.6 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__SREGSBP_1%VPWR 1 2 3 4 5 6 7 8 9 30 34 38 44 48 52
+ 56 58 62 68 71 72 74 75 77 78 80 81 83 84 86 87 88 115 119 135 136 139 142 145
r187 145 146 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.76 $Y=3.33
+ $X2=11.76 $Y2=3.33
r188 143 146 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=10.8 $Y=3.33
+ $X2=11.76 $Y2=3.33
r189 142 143 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=3.33
+ $X2=10.8 $Y2=3.33
r190 139 140 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r191 135 136 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=14.16 $Y=3.33
+ $X2=14.16 $Y2=3.33
r192 133 136 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=13.2 $Y=3.33
+ $X2=14.16 $Y2=3.33
r193 132 133 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=13.2 $Y=3.33
+ $X2=13.2 $Y2=3.33
r194 130 133 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=12.24 $Y=3.33
+ $X2=13.2 $Y2=3.33
r195 130 146 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.24 $Y=3.33
+ $X2=11.76 $Y2=3.33
r196 129 132 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=12.24 $Y=3.33
+ $X2=13.2 $Y2=3.33
r197 129 130 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=12.24 $Y=3.33
+ $X2=12.24 $Y2=3.33
r198 127 145 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.04 $Y=3.33
+ $X2=11.875 $Y2=3.33
r199 127 129 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=12.04 $Y=3.33
+ $X2=12.24 $Y2=3.33
r200 126 143 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=3.33
+ $X2=10.8 $Y2=3.33
r201 125 126 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=10.32 $Y=3.33
+ $X2=10.32 $Y2=3.33
r202 123 126 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=10.32 $Y2=3.33
r203 123 140 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=8.88 $Y2=3.33
r204 122 125 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=9.36 $Y=3.33
+ $X2=10.32 $Y2=3.33
r205 122 123 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r206 120 139 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.03 $Y=3.33
+ $X2=8.865 $Y2=3.33
r207 120 122 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=9.03 $Y=3.33
+ $X2=9.36 $Y2=3.33
r208 119 142 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.69 $Y=3.33
+ $X2=10.855 $Y2=3.33
r209 119 125 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=10.69 $Y=3.33
+ $X2=10.32 $Y2=3.33
r210 118 140 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=8.88 $Y2=3.33
r211 117 118 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r212 115 139 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.7 $Y=3.33
+ $X2=8.865 $Y2=3.33
r213 115 117 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=8.7 $Y=3.33 $X2=8.4
+ $Y2=3.33
r214 114 118 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=8.4 $Y2=3.33
r215 113 114 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r216 110 111 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r217 108 111 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=6.48 $Y2=3.33
r218 107 110 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=4.56 $Y=3.33
+ $X2=6.48 $Y2=3.33
r219 107 108 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r220 105 108 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r221 104 105 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r222 102 105 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=4.08 $Y2=3.33
r223 101 104 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=3.12 $Y=3.33
+ $X2=4.08 $Y2=3.33
r224 101 102 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r225 99 102 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r226 98 99 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r227 96 99 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r228 95 98 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r229 95 96 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r230 92 96 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r231 91 92 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r232 88 114 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=7.2 $Y=3.33
+ $X2=7.44 $Y2=3.33
r233 88 111 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=7.2 $Y=3.33
+ $X2=6.48 $Y2=3.33
r234 86 132 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=13.395 $Y=3.33
+ $X2=13.2 $Y2=3.33
r235 86 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.395 $Y=3.33
+ $X2=13.56 $Y2=3.33
r236 85 135 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=13.725 $Y=3.33
+ $X2=14.16 $Y2=3.33
r237 85 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.725 $Y=3.33
+ $X2=13.56 $Y2=3.33
r238 83 113 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=7.595 $Y=3.33
+ $X2=7.44 $Y2=3.33
r239 83 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.595 $Y=3.33
+ $X2=7.76 $Y2=3.33
r240 82 117 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=7.925 $Y=3.33
+ $X2=8.4 $Y2=3.33
r241 82 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.925 $Y=3.33
+ $X2=7.76 $Y2=3.33
r242 80 110 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=6.57 $Y=3.33
+ $X2=6.48 $Y2=3.33
r243 80 81 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.57 $Y=3.33
+ $X2=6.695 $Y2=3.33
r244 79 113 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=6.82 $Y=3.33
+ $X2=7.44 $Y2=3.33
r245 79 81 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.82 $Y=3.33
+ $X2=6.695 $Y2=3.33
r246 77 104 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=4.215 $Y=3.33
+ $X2=4.08 $Y2=3.33
r247 77 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.215 $Y=3.33
+ $X2=4.38 $Y2=3.33
r248 76 107 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=4.545 $Y=3.33
+ $X2=4.56 $Y2=3.33
r249 76 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.545 $Y=3.33
+ $X2=4.38 $Y2=3.33
r250 74 98 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=2.645 $Y=3.33
+ $X2=2.64 $Y2=3.33
r251 74 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.645 $Y=3.33
+ $X2=2.81 $Y2=3.33
r252 73 101 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=2.975 $Y=3.33
+ $X2=3.12 $Y2=3.33
r253 73 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.975 $Y=3.33
+ $X2=2.81 $Y2=3.33
r254 71 91 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=0.865 $Y=3.33
+ $X2=0.72 $Y2=3.33
r255 71 72 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.865 $Y=3.33
+ $X2=1.03 $Y2=3.33
r256 70 95 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=1.195 $Y=3.33
+ $X2=1.2 $Y2=3.33
r257 70 72 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.195 $Y=3.33
+ $X2=1.03 $Y2=3.33
r258 66 87 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=13.56 $Y=3.245
+ $X2=13.56 $Y2=3.33
r259 66 68 12.2229 $w=3.28e-07 $l=3.5e-07 $layer=LI1_cond $X=13.56 $Y=3.245
+ $X2=13.56 $Y2=2.895
r260 62 65 17.8105 $w=3.28e-07 $l=5.1e-07 $layer=LI1_cond $X=11.875 $Y=2.44
+ $X2=11.875 $Y2=2.95
r261 60 145 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=11.875 $Y=3.245
+ $X2=11.875 $Y2=3.33
r262 60 65 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=11.875 $Y=3.245
+ $X2=11.875 $Y2=2.95
r263 59 142 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.02 $Y=3.33
+ $X2=10.855 $Y2=3.33
r264 58 145 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.71 $Y=3.33
+ $X2=11.875 $Y2=3.33
r265 58 59 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=11.71 $Y=3.33
+ $X2=11.02 $Y2=3.33
r266 54 142 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.855 $Y=3.245
+ $X2=10.855 $Y2=3.33
r267 54 56 12.2229 $w=3.28e-07 $l=3.5e-07 $layer=LI1_cond $X=10.855 $Y=3.245
+ $X2=10.855 $Y2=2.895
r268 50 139 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.865 $Y=3.245
+ $X2=8.865 $Y2=3.33
r269 50 52 41.7324 $w=3.28e-07 $l=1.195e-06 $layer=LI1_cond $X=8.865 $Y=3.245
+ $X2=8.865 $Y2=2.05
r270 46 84 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.76 $Y=3.245
+ $X2=7.76 $Y2=3.33
r271 46 48 13.969 $w=3.28e-07 $l=4e-07 $layer=LI1_cond $X=7.76 $Y=3.245 $X2=7.76
+ $Y2=2.845
r272 42 81 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.695 $Y=3.245
+ $X2=6.695 $Y2=3.33
r273 42 44 33.1904 $w=2.48e-07 $l=7.2e-07 $layer=LI1_cond $X=6.695 $Y=3.245
+ $X2=6.695 $Y2=2.525
r274 38 41 24.0965 $w=3.28e-07 $l=6.9e-07 $layer=LI1_cond $X=4.38 $Y=2.21
+ $X2=4.38 $Y2=2.9
r275 36 78 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.38 $Y=3.245
+ $X2=4.38 $Y2=3.33
r276 36 41 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=4.38 $Y=3.245
+ $X2=4.38 $Y2=2.9
r277 32 75 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.81 $Y=3.245
+ $X2=2.81 $Y2=3.33
r278 32 34 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=2.81 $Y=3.245
+ $X2=2.81 $Y2=2.93
r279 28 72 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.03 $Y=3.245
+ $X2=1.03 $Y2=3.33
r280 28 30 13.2706 $w=3.28e-07 $l=3.8e-07 $layer=LI1_cond $X=1.03 $Y=3.245
+ $X2=1.03 $Y2=2.865
r281 9 68 600 $w=1.7e-07 $l=1.12783e-06 $layer=licon1_PDIFF $count=1 $X=13.42
+ $Y=1.835 $X2=13.56 $Y2=2.895
r282 8 65 600 $w=1.7e-07 $l=7.97449e-07 $layer=licon1_PDIFF $count=1 $X=11.655
+ $Y=2.255 $X2=11.875 $Y2=2.95
r283 8 62 600 $w=1.7e-07 $l=2.98496e-07 $layer=licon1_PDIFF $count=1 $X=11.655
+ $Y=2.255 $X2=11.875 $Y2=2.44
r284 7 56 600 $w=1.7e-07 $l=7.56836e-07 $layer=licon1_PDIFF $count=1 $X=10.6
+ $Y=2.255 $X2=10.855 $Y2=2.895
r285 6 52 300 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_PDIFF $count=2 $X=8.72
+ $Y=1.865 $X2=8.865 $Y2=2.05
r286 5 48 600 $w=1.7e-07 $l=1.10014e-06 $layer=licon1_PDIFF $count=1 $X=7.505
+ $Y=1.865 $X2=7.76 $Y2=2.845
r287 4 44 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=6.515
+ $Y=2.315 $X2=6.655 $Y2=2.525
r288 3 41 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=4.24
+ $Y=1.785 $X2=4.38 $Y2=2.9
r289 3 38 400 $w=1.7e-07 $l=4.90026e-07 $layer=licon1_PDIFF $count=1 $X=4.24
+ $Y=1.785 $X2=4.38 $Y2=2.21
r290 2 34 600 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=1 $X=2.67
+ $Y=2.655 $X2=2.81 $Y2=2.93
r291 1 30 600 $w=1.7e-07 $l=3.07571e-07 $layer=licon1_PDIFF $count=1 $X=0.81
+ $Y=2.655 $X2=1.03 $Y2=2.865
.ends

.subckt PM_SKY130_FD_SC_LP__SREGSBP_1%A_636_531# 1 2 8 10 15
c39 15 0 2.16488e-19 $X=3.6 $Y=0.47
r40 13 15 5.90276 $w=4.08e-07 $l=2.1e-07 $layer=LI1_cond $X=3.39 $Y=0.47 $X2=3.6
+ $Y2=0.47
r41 8 10 11.1634 $w=3.06e-07 $l=3.64692e-07 $layer=LI1_cond $X=3.6 $Y=2.675
+ $X2=3.32 $Y2=2.87
r42 7 15 5.92876 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=3.6 $Y=0.675 $X2=3.6
+ $Y2=0.47
r43 7 8 130.481 $w=1.68e-07 $l=2e-06 $layer=LI1_cond $X=3.6 $Y=0.675 $X2=3.6
+ $Y2=2.675
r44 2 10 600 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_PDIFF $count=1 $X=3.18
+ $Y=2.655 $X2=3.32 $Y2=2.87
r45 1 13 182 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=1 $X=3.25
+ $Y=0.235 $X2=3.39 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_LP__SREGSBP_1%Q_N 1 2 9 11 14 17
r37 12 21 21.9284 $w=3.58e-07 $l=6.85e-07 $layer=LI1_cond $X=13.145 $Y=1.295
+ $X2=13.145 $Y2=1.98
r38 12 17 27.6906 $w=3.58e-07 $l=8.65e-07 $layer=LI1_cond $X=13.145 $Y=1.295
+ $X2=13.145 $Y2=0.43
r39 11 12 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.2 $Y=1.295
+ $X2=13.2 $Y2=1.295
r40 9 14 0.414603 $w=1.4e-07 $l=3.35e-07 $layer=MET1_cond $X=13.345 $Y=1.295
+ $X2=13.68 $Y2=1.295
r41 9 11 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=13.345 $Y=1.295
+ $X2=13.2 $Y2=1.295
r42 2 21 600 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=12.985
+ $Y=1.835 $X2=13.13 $Y2=1.98
r43 1 17 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=13.015
+ $Y=0.285 $X2=13.16 $Y2=0.43
.ends

.subckt PM_SKY130_FD_SC_LP__SREGSBP_1%Q 1 2 9 13 17 20 22 25 28 29
c44 28 0 1.66705e-19 $X=14.07 $Y=2
r45 28 29 8.6688 $w=4.03e-07 $l=1.65e-07 $layer=LI1_cond $X=14.107 $Y=2
+ $X2=14.107 $Y2=1.835
r46 22 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.16 $Y=2.035
+ $X2=14.16 $Y2=2.035
r47 20 25 0.414603 $w=1.4e-07 $l=3.35e-07 $layer=MET1_cond $X=14.015 $Y=2.035
+ $X2=13.68 $Y2=2.035
r48 20 22 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=14.015 $Y=2.035
+ $X2=14.16 $Y2=2.035
r49 17 29 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=14.225 $Y=1.145
+ $X2=14.225 $Y2=1.835
r50 11 17 9.23056 $w=3.73e-07 $l=1.87e-07 $layer=LI1_cond $X=14.122 $Y=0.958
+ $X2=14.122 $Y2=1.145
r51 11 13 16.2264 $w=3.73e-07 $l=5.28e-07 $layer=LI1_cond $X=14.122 $Y=0.958
+ $X2=14.122 $Y2=0.43
r52 7 28 1.05285 $w=4.03e-07 $l=3.7e-08 $layer=LI1_cond $X=14.107 $Y=2.037
+ $X2=14.107 $Y2=2
r53 7 9 24.557 $w=4.03e-07 $l=8.63e-07 $layer=LI1_cond $X=14.107 $Y=2.037
+ $X2=14.107 $Y2=2.9
r54 2 28 400 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_PDIFF $count=1 $X=13.93
+ $Y=1.835 $X2=14.07 $Y2=2
r55 2 9 400 $w=1.7e-07 $l=1.13284e-06 $layer=licon1_PDIFF $count=1 $X=13.93
+ $Y=1.835 $X2=14.07 $Y2=2.9
r56 1 13 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=13.96
+ $Y=0.285 $X2=14.1 $Y2=0.43
.ends

.subckt PM_SKY130_FD_SC_LP__SREGSBP_1%VGND 1 2 3 4 5 6 7 8 9 28 30 34 38 42 46
+ 50 54 58 62 65 66 68 69 71 72 73 75 87 101 108 113 123 124 130 133 136 139 142
c177 65 0 1.96333e-19 $X=2.795 $Y=0
r178 142 143 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=12.24 $Y=0
+ $X2=12.24 $Y2=0
r179 139 140 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=0
+ $X2=10.8 $Y2=0
r180 136 137 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.88 $Y=0
+ $X2=8.88 $Y2=0
r181 133 134 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=0
+ $X2=4.56 $Y2=0
r182 130 131 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r183 127 128 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0
+ $X2=0.24 $Y2=0
r184 123 124 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=14.16 $Y=0
+ $X2=14.16 $Y2=0
r185 121 124 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=13.2 $Y=0
+ $X2=14.16 $Y2=0
r186 121 143 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=13.2 $Y=0
+ $X2=12.24 $Y2=0
r187 120 121 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=13.2 $Y=0
+ $X2=13.2 $Y2=0
r188 118 142 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=12.255 $Y=0
+ $X2=12.13 $Y2=0
r189 118 120 61.6524 $w=1.68e-07 $l=9.45e-07 $layer=LI1_cond $X=12.255 $Y=0
+ $X2=13.2 $Y2=0
r190 117 143 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.76 $Y=0
+ $X2=12.24 $Y2=0
r191 117 140 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=11.76 $Y=0
+ $X2=10.8 $Y2=0
r192 116 117 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.76 $Y=0
+ $X2=11.76 $Y2=0
r193 114 139 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.985 $Y=0
+ $X2=10.82 $Y2=0
r194 114 116 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=10.985 $Y=0
+ $X2=11.76 $Y2=0
r195 113 142 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=12.005 $Y=0
+ $X2=12.13 $Y2=0
r196 113 116 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=12.005 $Y=0
+ $X2=11.76 $Y2=0
r197 112 140 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=0
+ $X2=10.8 $Y2=0
r198 112 137 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=10.32 $Y=0
+ $X2=8.88 $Y2=0
r199 111 112 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.32 $Y=0
+ $X2=10.32 $Y2=0
r200 109 136 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.885 $Y=0
+ $X2=8.76 $Y2=0
r201 109 111 93.6203 $w=1.68e-07 $l=1.435e-06 $layer=LI1_cond $X=8.885 $Y=0
+ $X2=10.32 $Y2=0
r202 108 139 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.655 $Y=0
+ $X2=10.82 $Y2=0
r203 108 111 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=10.655 $Y=0
+ $X2=10.32 $Y2=0
r204 107 137 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=0
+ $X2=8.88 $Y2=0
r205 106 107 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r206 104 107 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.44 $Y=0
+ $X2=8.4 $Y2=0
r207 103 106 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=7.44 $Y=0 $X2=8.4
+ $Y2=0
r208 103 104 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=7.44 $Y=0
+ $X2=7.44 $Y2=0
r209 101 136 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.635 $Y=0
+ $X2=8.76 $Y2=0
r210 101 106 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=8.635 $Y=0
+ $X2=8.4 $Y2=0
r211 99 100 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.96 $Y=0
+ $X2=6.96 $Y2=0
r212 97 100 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=5.04 $Y=0
+ $X2=6.96 $Y2=0
r213 97 134 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0
+ $X2=4.56 $Y2=0
r214 96 99 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=5.04 $Y=0 $X2=6.96
+ $Y2=0
r215 96 97 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.04 $Y=0
+ $X2=5.04 $Y2=0
r216 94 133 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.665 $Y=0 $X2=4.5
+ $Y2=0
r217 94 96 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=4.665 $Y=0
+ $X2=5.04 $Y2=0
r218 93 134 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0
+ $X2=4.56 $Y2=0
r219 92 93 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r220 90 93 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=4.08
+ $Y2=0
r221 89 92 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=3.12 $Y=0 $X2=4.08
+ $Y2=0
r222 89 90 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r223 87 133 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.335 $Y=0 $X2=4.5
+ $Y2=0
r224 87 92 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=4.335 $Y=0
+ $X2=4.08 $Y2=0
r225 86 90 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r226 85 86 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r227 83 86 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r228 83 131 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r229 82 85 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r230 82 83 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r231 80 130 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.435 $Y=0
+ $X2=1.27 $Y2=0
r232 80 82 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=1.435 $Y=0 $X2=1.68
+ $Y2=0
r233 79 131 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r234 79 128 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0
+ $X2=0.24 $Y2=0
r235 78 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r236 76 127 4.00981 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=0.365 $Y=0
+ $X2=0.182 $Y2=0
r237 76 78 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=0.365 $Y=0
+ $X2=0.72 $Y2=0
r238 75 130 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.105 $Y=0
+ $X2=1.27 $Y2=0
r239 75 78 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=1.105 $Y=0
+ $X2=0.72 $Y2=0
r240 73 104 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=7.2 $Y=0
+ $X2=7.44 $Y2=0
r241 73 100 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=7.2 $Y=0
+ $X2=6.96 $Y2=0
r242 71 120 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=13.505 $Y=0
+ $X2=13.2 $Y2=0
r243 71 72 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=13.505 $Y=0
+ $X2=13.63 $Y2=0
r244 70 123 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=13.755 $Y=0
+ $X2=14.16 $Y2=0
r245 70 72 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=13.755 $Y=0
+ $X2=13.63 $Y2=0
r246 68 99 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=7.05 $Y=0 $X2=6.96
+ $Y2=0
r247 68 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.05 $Y=0 $X2=7.215
+ $Y2=0
r248 67 103 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=7.38 $Y=0 $X2=7.44
+ $Y2=0
r249 67 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.38 $Y=0 $X2=7.215
+ $Y2=0
r250 65 85 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=2.795 $Y=0
+ $X2=2.64 $Y2=0
r251 65 66 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.795 $Y=0 $X2=2.92
+ $Y2=0
r252 64 89 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=3.045 $Y=0 $X2=3.12
+ $Y2=0
r253 64 66 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.045 $Y=0 $X2=2.92
+ $Y2=0
r254 60 72 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=13.63 $Y=0.085
+ $X2=13.63 $Y2=0
r255 60 62 15.9037 $w=2.48e-07 $l=3.45e-07 $layer=LI1_cond $X=13.63 $Y=0.085
+ $X2=13.63 $Y2=0.43
r256 56 142 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=12.13 $Y=0.085
+ $X2=12.13 $Y2=0
r257 56 58 18.9001 $w=2.48e-07 $l=4.1e-07 $layer=LI1_cond $X=12.13 $Y=0.085
+ $X2=12.13 $Y2=0.495
r258 52 139 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.82 $Y=0.085
+ $X2=10.82 $Y2=0
r259 52 54 14.8421 $w=3.28e-07 $l=4.25e-07 $layer=LI1_cond $X=10.82 $Y=0.085
+ $X2=10.82 $Y2=0.51
r260 48 136 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=8.76 $Y=0.085
+ $X2=8.76 $Y2=0
r261 48 50 37.5696 $w=2.48e-07 $l=8.15e-07 $layer=LI1_cond $X=8.76 $Y=0.085
+ $X2=8.76 $Y2=0.9
r262 44 69 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.215 $Y=0.085
+ $X2=7.215 $Y2=0
r263 44 46 27.938 $w=3.28e-07 $l=8e-07 $layer=LI1_cond $X=7.215 $Y=0.085
+ $X2=7.215 $Y2=0.885
r264 40 133 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.5 $Y=0.085
+ $X2=4.5 $Y2=0
r265 40 42 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=4.5 $Y=0.085
+ $X2=4.5 $Y2=0.43
r266 36 66 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.92 $Y=0.085
+ $X2=2.92 $Y2=0
r267 36 38 16.5952 $w=2.48e-07 $l=3.6e-07 $layer=LI1_cond $X=2.92 $Y=0.085
+ $X2=2.92 $Y2=0.445
r268 32 130 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.27 $Y=0.085
+ $X2=1.27 $Y2=0
r269 32 34 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=1.27 $Y=0.085
+ $X2=1.27 $Y2=0.445
r270 28 127 3.13335 $w=2.5e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.24 $Y=0.085
+ $X2=0.182 $Y2=0
r271 28 30 18.2086 $w=2.48e-07 $l=3.95e-07 $layer=LI1_cond $X=0.24 $Y=0.085
+ $X2=0.24 $Y2=0.48
r272 9 62 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=13.45
+ $Y=0.285 $X2=13.59 $Y2=0.43
r273 8 58 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=12.025
+ $Y=0.285 $X2=12.17 $Y2=0.495
r274 7 54 182 $w=1.7e-07 $l=2.81158e-07 $layer=licon1_NDIFF $count=1 $X=10.565
+ $Y=0.455 $X2=10.82 $Y2=0.51
r275 6 50 182 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=1 $X=8.575
+ $Y=0.625 $X2=8.72 $Y2=0.9
r276 5 46 182 $w=1.7e-07 $l=3.99375e-07 $layer=licon1_NDIFF $count=1 $X=6.955
+ $Y=0.595 $X2=7.215 $Y2=0.885
r277 4 42 182 $w=1.7e-07 $l=3.02159e-07 $layer=licon1_NDIFF $count=1 $X=4.28
+ $Y=0.235 $X2=4.5 $Y2=0.43
r278 3 38 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.82
+ $Y=0.235 $X2=2.96 $Y2=0.445
r279 2 34 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=1.125
+ $Y=0.235 $X2=1.27 $Y2=0.445
r280 1 30 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.27 $X2=0.28 $Y2=0.48
.ends

