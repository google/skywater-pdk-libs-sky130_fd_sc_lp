* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__a221oi_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
M1000 a_1334_47# A1 Y VNB nshort w=840000u l=150000u
+  ad=9.408e+11p pd=8.96e+06u as=1.4112e+12p ps=1.344e+07u
M1001 a_546_47# B2 VGND VNB nshort w=840000u l=150000u
+  ad=1.2936e+12p pd=9.8e+06u as=1.6884e+12p ps=1.578e+07u
M1002 VGND B2 a_546_47# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_533_367# B1 a_85_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=3.2886e+12p pd=2.79e+07u as=2.4318e+12p ps=2.15e+07u
M1004 a_533_367# B2 a_85_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_533_367# A2 VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=1.449e+12p ps=1.238e+07u
M1006 a_546_47# B1 Y VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND C1 Y VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_85_367# B2 a_533_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_533_367# A1 VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR A1 a_533_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_533_367# B1 a_85_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 Y B1 a_546_47# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VGND A2 a_1334_47# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VPWR A2 a_533_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VGND A2 a_1334_47# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 Y C1 a_85_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=7.056e+11p pd=6.16e+06u as=0p ps=0u
M1017 Y A1 a_1334_47# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_1334_47# A2 VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VPWR A2 a_533_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 Y A1 a_1334_47# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_546_47# B2 VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 Y C1 a_85_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_85_367# B2 a_533_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_533_367# A1 VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 Y C1 VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 Y B1 a_546_47# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_546_47# B1 Y VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 Y C1 VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 a_1334_47# A2 VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 a_85_367# B1 a_533_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_85_367# C1 Y VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 a_533_367# B2 a_85_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 a_533_367# A2 VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1034 VGND B2 a_546_47# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1035 a_85_367# B1 a_533_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1036 VGND C1 Y VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1037 a_85_367# C1 Y VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1038 VPWR A1 a_533_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1039 a_1334_47# A1 Y VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
