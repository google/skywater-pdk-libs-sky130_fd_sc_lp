* NGSPICE file created from sky130_fd_sc_lp__dlxtn_1.ext - technology: sky130A

.subckt sky130_fd_sc_lp__dlxtn_1 D GATE_N VGND VNB VPB VPWR Q
M1000 VPWR a_228_129# a_342_481# VPB phighvt w=640000u l=150000u
+  ad=1.5034e+12p pd=1.167e+07u as=1.696e+11p ps=1.81e+06u
M1001 VPWR D a_59_129# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.696e+11p ps=1.81e+06u
M1002 a_764_481# a_228_129# a_656_481# VPB phighvt w=420000u l=150000u
+  ad=1.638e+11p pd=1.62e+06u as=2.221e+11p ps=2.06e+06u
M1003 a_656_47# a_59_129# VGND VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=7.266e+11p ps=7.44e+06u
M1004 a_228_129# GATE_N VGND VNB nshort w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1005 a_228_129# GATE_N VPWR VPB phighvt w=640000u l=150000u
+  ad=1.696e+11p pd=1.81e+06u as=0p ps=0u
M1006 Q a_842_413# VGND VNB nshort w=840000u l=150000u
+  ad=2.226e+11p pd=2.21e+06u as=0p ps=0u
M1007 VPWR a_842_413# a_764_481# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_836_47# a_342_481# a_656_481# VNB nshort w=420000u l=150000u
+  ad=1.638e+11p pd=1.62e+06u as=1.638e+11p ps=1.62e+06u
M1009 VGND D a_59_129# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1010 a_842_413# a_656_481# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=3.339e+11p pd=3.05e+06u as=0p ps=0u
M1011 VGND a_228_129# a_342_481# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1012 a_584_481# a_59_129# VPWR VPB phighvt w=640000u l=150000u
+  ad=1.344e+11p pd=1.7e+06u as=0p ps=0u
M1013 a_656_481# a_342_481# a_584_481# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VGND a_842_413# a_836_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 Q a_842_413# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=3.339e+11p pd=3.05e+06u as=0p ps=0u
M1016 a_656_481# a_228_129# a_656_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_842_413# a_656_481# VGND VNB nshort w=840000u l=150000u
+  ad=2.226e+11p pd=2.21e+06u as=0p ps=0u
.ends

