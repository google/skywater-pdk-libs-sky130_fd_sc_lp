# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_sc_lp__srdlrtp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_lp__srdlrtp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  12.00000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 1.080000 0.435000 1.410000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.598500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.555000 0.255000 11.915000 1.135000 ;
        RECT 11.555000 1.815000 11.915000 3.075000 ;
        RECT 11.745000 1.135000 11.915000 1.815000 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  0.472000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1.055000 1.920000 1.345000 1.965000 ;
        RECT 1.055000 1.965000 9.505000 2.105000 ;
        RECT 1.055000 2.105000 1.345000 2.150000 ;
        RECT 9.215000 1.920000 9.505000 1.965000 ;
        RECT 9.215000 2.105000 9.505000 2.150000 ;
    END
  END RESET_B
  PIN SLEEP_B
    ANTENNAGATEAREA  0.598000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.885000 1.140000 6.595000 1.470000 ;
    END
  END SLEEP_B
  PIN GATE
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 5.045000 1.090000 5.635000 1.420000 ;
    END
  END GATE
  PIN KAPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.070000 2.675000 11.930000 2.945000 ;
    END
  END KAPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 12.000000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.000000 0.000000 12.000000 0.245000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.655000 12.190000 3.520000 ;
        RECT  5.055000 1.400000  7.200000 1.655000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 12.000000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 12.000000 0.085000 ;
      RECT  0.000000  3.245000 12.000000 3.415000 ;
      RECT  0.115000  0.465000  0.445000 0.740000 ;
      RECT  0.115000  0.740000  0.775000 0.910000 ;
      RECT  0.115000  2.765000  0.445000 3.245000 ;
      RECT  0.605000  0.910000  0.775000 1.580000 ;
      RECT  0.605000  1.580000  1.470000 1.750000 ;
      RECT  0.605000  1.750000  0.775000 2.425000 ;
      RECT  0.605000  2.425000  0.945000 2.595000 ;
      RECT  0.615000  2.595000  0.945000 3.075000 ;
      RECT  0.945000  0.085000  1.195000 0.845000 ;
      RECT  0.945000  1.920000  1.315000 2.255000 ;
      RECT  1.140000  1.015000  1.470000 1.580000 ;
      RECT  1.160000  2.425000  1.490000 3.245000 ;
      RECT  1.375000  0.465000  1.830000 0.845000 ;
      RECT  1.660000  0.845000  1.830000 2.415000 ;
      RECT  1.660000  2.415000  1.990000 3.075000 ;
      RECT  2.000000  0.255000  3.010000 0.425000 ;
      RECT  2.000000  0.425000  2.170000 1.095000 ;
      RECT  2.000000  1.095000  2.330000 1.425000 ;
      RECT  2.360000  0.595000  2.670000 0.865000 ;
      RECT  2.360000  0.865000  3.730000 0.925000 ;
      RECT  2.450000  2.415000  2.780000 3.075000 ;
      RECT  2.500000  0.925000  3.730000 1.035000 ;
      RECT  2.500000  1.035000  2.780000 2.415000 ;
      RECT  2.840000  0.425000  3.010000 0.525000 ;
      RECT  2.840000  0.525000  4.535000 0.695000 ;
      RECT  2.960000  1.205000  3.390000 1.445000 ;
      RECT  2.960000  1.445000  3.130000 2.635000 ;
      RECT  2.960000  2.635000  4.770000 2.805000 ;
      RECT  3.300000  1.615000  3.730000 1.785000 ;
      RECT  3.300000  1.785000  3.470000 2.295000 ;
      RECT  3.300000  2.295000  4.430000 2.465000 ;
      RECT  3.560000  1.035000  3.730000 1.615000 ;
      RECT  3.640000  1.955000  4.070000 2.125000 ;
      RECT  3.660000  0.085000  3.990000 0.355000 ;
      RECT  3.900000  0.695000  4.535000 0.925000 ;
      RECT  3.900000  0.925000  4.070000 1.955000 ;
      RECT  4.205000  0.255000  5.975000 0.425000 ;
      RECT  4.205000  0.425000  4.535000 0.525000 ;
      RECT  4.260000  1.980000  7.760000 2.150000 ;
      RECT  4.260000  2.150000  4.430000 2.295000 ;
      RECT  4.300000  2.975000  4.630000 3.245000 ;
      RECT  4.375000  1.105000  4.875000 1.640000 ;
      RECT  4.375000  1.640000  5.735000 1.810000 ;
      RECT  4.600000  2.320000  6.735000 2.490000 ;
      RECT  4.600000  2.490000  4.770000 2.635000 ;
      RECT  4.705000  0.595000  5.220000 0.920000 ;
      RECT  4.705000  0.920000  4.875000 1.105000 ;
      RECT  4.940000  2.660000  5.635000 2.990000 ;
      RECT  5.805000  0.425000  5.975000 0.800000 ;
      RECT  5.805000  0.800000  7.000000 0.970000 ;
      RECT  5.885000  2.660000  6.395000 2.990000 ;
      RECT  6.150000  0.085000  6.480000 0.630000 ;
      RECT  6.565000  2.490000  6.735000 2.905000 ;
      RECT  6.565000  2.905000  8.100000 3.075000 ;
      RECT  6.710000  1.640000  7.040000 1.810000 ;
      RECT  6.830000  0.255000  7.920000 0.425000 ;
      RECT  6.830000  0.425000  7.000000 0.800000 ;
      RECT  6.870000  1.140000  7.420000 1.310000 ;
      RECT  6.870000  1.310000  7.040000 1.640000 ;
      RECT  7.170000  0.595000  7.420000 0.875000 ;
      RECT  7.170000  0.875000  8.715000 1.135000 ;
      RECT  7.170000  1.135000  7.420000 1.140000 ;
      RECT  7.270000  2.150000  7.760000 2.735000 ;
      RECT  7.590000  0.425000  7.920000 0.585000 ;
      RECT  7.590000  1.305000  9.765000 1.365000 ;
      RECT  7.590000  1.365000  9.055000 1.475000 ;
      RECT  7.590000  1.475000  7.760000 1.980000 ;
      RECT  7.930000  1.645000  8.365000 1.935000 ;
      RECT  7.930000  1.935000  8.100000 2.320000 ;
      RECT  7.930000  2.320000 10.295000 2.490000 ;
      RECT  7.930000  2.490000  8.100000 2.905000 ;
      RECT  8.180000  0.255000  8.430000 0.535000 ;
      RECT  8.180000  0.535000  9.455000 0.705000 ;
      RECT  8.270000  2.660000  8.600000 3.075000 ;
      RECT  8.610000  0.085000  8.940000 0.365000 ;
      RECT  8.885000  1.035000  9.765000 1.305000 ;
      RECT  9.125000  0.255000  9.455000 0.535000 ;
      RECT  9.225000  1.550000  9.955000 2.150000 ;
      RECT  9.375000  2.490000  9.705000 3.075000 ;
      RECT  9.920000  0.255000 10.295000 0.675000 ;
      RECT 10.020000  2.660000 10.435000 3.075000 ;
      RECT 10.125000  0.675000 10.295000 2.320000 ;
      RECT 10.580000  0.255000 10.910000 1.315000 ;
      RECT 10.580000  1.315000 11.575000 1.645000 ;
      RECT 10.580000  1.645000 10.910000 2.490000 ;
      RECT 11.125000  0.085000 11.375000 0.965000 ;
      RECT 11.125000  1.815000 11.375000 3.245000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  1.950000  1.285000 2.120000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  2.735000  5.605000 2.905000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  2.735000  6.085000 2.905000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  2.735000  8.485000 2.905000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  1.950000  9.445000 2.120000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  2.735000 10.405000 2.905000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.245000 10.885000 3.415000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  3.245000 11.365000 3.415000 ;
      RECT 11.675000 -0.085000 11.845000 0.085000 ;
      RECT 11.675000  3.245000 11.845000 3.415000 ;
  END
END sky130_fd_sc_lp__srdlrtp_1
END LIBRARY
