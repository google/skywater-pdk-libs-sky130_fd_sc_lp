* File: sky130_fd_sc_lp__a21oi_lp.pex.spice
* Created: Fri Aug 28 09:51:58 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A21OI_LP%A2 2 5 7 11 13 14 15 18 19
r38 18 20 46.6684 $w=4.4e-07 $l=1.65e-07 $layer=POLY_cond $X=0.44 $Y=1.02
+ $X2=0.44 $Y2=0.855
r39 18 19 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.385
+ $Y=1.02 $X2=0.385 $Y2=1.02
r40 15 19 2.58853 $w=6.68e-07 $l=1.45e-07 $layer=LI1_cond $X=0.24 $Y=1.19
+ $X2=0.385 $Y2=1.19
r41 13 14 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=0.515 $Y=1.525
+ $X2=0.515 $Y2=1.765
r42 11 20 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=0.585 $Y=0.445
+ $X2=0.585 $Y2=0.855
r43 5 14 40.9178 $w=2.5e-07 $l=1.25e-07 $layer=POLY_cond $X=0.565 $Y=1.89
+ $X2=0.565 $Y2=1.765
r44 5 7 162.737 $w=2.5e-07 $l=6.55e-07 $layer=POLY_cond $X=0.565 $Y=1.89
+ $X2=0.565 $Y2=2.545
r45 2 13 45.2162 $w=4.4e-07 $l=2.2e-07 $layer=POLY_cond $X=0.44 $Y=1.305
+ $X2=0.44 $Y2=1.525
r46 1 18 6.95192 $w=4.4e-07 $l=5.5e-08 $layer=POLY_cond $X=0.44 $Y=1.075
+ $X2=0.44 $Y2=1.02
r47 1 2 29.0717 $w=4.4e-07 $l=2.3e-07 $layer=POLY_cond $X=0.44 $Y=1.075 $X2=0.44
+ $Y2=1.305
.ends

.subckt PM_SKY130_FD_SC_LP__A21OI_LP%A1 3 7 11 12 13 16
r41 16 17 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.065
+ $Y=1.24 $X2=1.065 $Y2=1.24
r42 13 17 2.41001 $w=6.68e-07 $l=1.35e-07 $layer=LI1_cond $X=1.2 $Y=1.41
+ $X2=1.065 $Y2=1.41
r43 11 16 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.065 $Y=1.58
+ $X2=1.065 $Y2=1.24
r44 11 12 31.6748 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.065 $Y=1.58
+ $X2=1.065 $Y2=1.745
r45 10 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.065 $Y=1.075
+ $X2=1.065 $Y2=1.24
r46 7 12 198.763 $w=2.5e-07 $l=8e-07 $layer=POLY_cond $X=1.095 $Y=2.545
+ $X2=1.095 $Y2=1.745
r47 3 10 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=0.975 $Y=0.445
+ $X2=0.975 $Y2=1.075
.ends

.subckt PM_SKY130_FD_SC_LP__A21OI_LP%B1 3 7 11 13 16
r40 16 18 66.9034 $w=5.1e-07 $l=5.05e-07 $layer=POLY_cond $X=1.725 $Y=1.24
+ $X2=1.725 $Y2=1.745
r41 13 16 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.66
+ $Y=1.24 $X2=1.66 $Y2=1.24
r42 9 16 32.933 $w=2.55e-07 $l=2.49199e-07 $layer=POLY_cond $X=1.905 $Y=1.075
+ $X2=1.725 $Y2=1.24
r43 9 11 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=1.905 $Y=1.075
+ $X2=1.905 $Y2=0.445
r44 7 18 198.763 $w=2.5e-07 $l=8e-07 $layer=POLY_cond $X=1.625 $Y=2.545
+ $X2=1.625 $Y2=1.745
r45 1 16 32.933 $w=2.55e-07 $l=2.49199e-07 $layer=POLY_cond $X=1.545 $Y=1.075
+ $X2=1.725 $Y2=1.24
r46 1 3 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=1.545 $Y=1.075
+ $X2=1.545 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__A21OI_LP%A_31_409# 1 2 9 13 14 17
r32 17 19 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=1.36 $Y=2.19 $X2=1.36
+ $Y2=2.9
r33 15 17 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=1.36 $Y=2.095
+ $X2=1.36 $Y2=2.19
r34 13 15 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.195 $Y=2.01
+ $X2=1.36 $Y2=2.095
r35 13 14 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=1.195 $Y=2.01
+ $X2=0.465 $Y2=2.01
r36 9 11 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=0.3 $Y=2.19 $X2=0.3
+ $Y2=2.9
r37 7 14 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.3 $Y=2.095
+ $X2=0.465 $Y2=2.01
r38 7 9 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=0.3 $Y=2.095 $X2=0.3
+ $Y2=2.19
r39 2 19 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=1.22
+ $Y=2.045 $X2=1.36 $Y2=2.9
r40 2 17 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.22
+ $Y=2.045 $X2=1.36 $Y2=2.19
r41 1 11 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.155
+ $Y=2.045 $X2=0.3 $Y2=2.9
r42 1 9 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.155
+ $Y=2.045 $X2=0.3 $Y2=2.19
.ends

.subckt PM_SKY130_FD_SC_LP__A21OI_LP%VPWR 1 8 10 17 18 21
r24 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r25 17 18 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r26 14 17 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=3.33 $X2=2.16
+ $Y2=3.33
r27 12 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.995 $Y=3.33
+ $X2=0.83 $Y2=3.33
r28 12 14 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=0.995 $Y=3.33
+ $X2=1.2 $Y2=3.33
r29 10 18 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r30 10 22 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r31 10 14 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r32 6 21 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.83 $Y=3.245 $X2=0.83
+ $Y2=3.33
r33 6 8 28.1126 $w=3.28e-07 $l=8.05e-07 $layer=LI1_cond $X=0.83 $Y=3.245
+ $X2=0.83 $Y2=2.44
r34 1 8 300 $w=1.7e-07 $l=4.59701e-07 $layer=licon1_PDIFF $count=2 $X=0.69
+ $Y=2.045 $X2=0.83 $Y2=2.44
.ends

.subckt PM_SKY130_FD_SC_LP__A21OI_LP%Y 1 2 9 11 12 13 14 15 16 17 27 30 49
r43 49 50 5.31909 $w=5.48e-07 $l=1e-08 $layer=LI1_cond $X=2 $Y=2.035 $X2=2
+ $Y2=2.025
r44 37 53 2.39216 $w=5.48e-07 $l=1.1e-07 $layer=LI1_cond $X=2 $Y=2.3 $X2=2
+ $Y2=2.19
r45 27 30 1.66364 $w=1.98e-07 $l=3e-08 $layer=LI1_cond $X=2.175 $Y=0.895
+ $X2=2.175 $Y2=0.925
r46 17 43 2.71836 $w=5.48e-07 $l=1.25e-07 $layer=LI1_cond $X=2 $Y=2.775 $X2=2
+ $Y2=2.9
r47 16 17 8.04635 $w=5.48e-07 $l=3.7e-07 $layer=LI1_cond $X=2 $Y=2.405 $X2=2
+ $Y2=2.775
r48 16 37 2.28342 $w=5.48e-07 $l=1.05e-07 $layer=LI1_cond $X=2 $Y=2.405 $X2=2
+ $Y2=2.3
r49 15 53 2.56613 $w=5.48e-07 $l=1.18e-07 $layer=LI1_cond $X=2 $Y=2.072 $X2=2
+ $Y2=2.19
r50 15 49 0.804635 $w=5.48e-07 $l=3.7e-08 $layer=LI1_cond $X=2 $Y=2.072 $X2=2
+ $Y2=2.035
r51 15 50 2.10727 $w=1.98e-07 $l=3.8e-08 $layer=LI1_cond $X=2.175 $Y=1.987
+ $X2=2.175 $Y2=2.025
r52 14 15 17.8564 $w=1.98e-07 $l=3.22e-07 $layer=LI1_cond $X=2.175 $Y=1.665
+ $X2=2.175 $Y2=1.987
r53 13 14 20.5182 $w=1.98e-07 $l=3.7e-07 $layer=LI1_cond $X=2.175 $Y=1.295
+ $X2=2.175 $Y2=1.665
r54 12 27 3.15876 $w=2e-07 $l=8.5e-08 $layer=LI1_cond $X=2.175 $Y=0.81 $X2=2.175
+ $Y2=0.895
r55 12 13 19.0209 $w=1.98e-07 $l=3.43e-07 $layer=LI1_cond $X=2.175 $Y=0.952
+ $X2=2.175 $Y2=1.295
r56 12 30 1.49727 $w=1.98e-07 $l=2.7e-08 $layer=LI1_cond $X=2.175 $Y=0.952
+ $X2=2.175 $Y2=0.925
r57 11 12 30.423 $w=2.23e-07 $l=5.8e-07 $layer=LI1_cond $X=1.495 $Y=0.81
+ $X2=2.075 $Y2=0.81
r58 7 11 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.33 $Y=0.725
+ $X2=1.495 $Y2=0.81
r59 7 9 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=1.33 $Y=0.725
+ $X2=1.33 $Y2=0.47
r60 2 53 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.75
+ $Y=2.045 $X2=1.89 $Y2=2.19
r61 2 43 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=1.75
+ $Y=2.045 $X2=1.89 $Y2=2.9
r62 1 9 182 $w=1.7e-07 $l=3.79737e-07 $layer=licon1_NDIFF $count=1 $X=1.05
+ $Y=0.235 $X2=1.33 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_LP__A21OI_LP%VGND 1 2 7 9 11 13 15 17 30
r33 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r34 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r35 24 30 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r36 23 24 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r37 21 27 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r38 20 23 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r39 20 21 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r40 18 26 4.56433 $w=1.7e-07 $l=2.68e-07 $layer=LI1_cond $X=0.535 $Y=0 $X2=0.267
+ $Y2=0
r41 18 20 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=0.535 $Y=0 $X2=0.72
+ $Y2=0
r42 17 29 4.73651 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=1.955 $Y=0 $X2=2.177
+ $Y2=0
r43 17 23 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=1.955 $Y=0 $X2=1.68
+ $Y2=0
r44 15 24 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r45 15 21 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r46 11 29 3.02966 $w=3.3e-07 $l=1.09864e-07 $layer=LI1_cond $X=2.12 $Y=0.085
+ $X2=2.177 $Y2=0
r47 11 13 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.12 $Y=0.085
+ $X2=2.12 $Y2=0.38
r48 7 26 3.20184 $w=3.3e-07 $l=1.39155e-07 $layer=LI1_cond $X=0.37 $Y=0.085
+ $X2=0.267 $Y2=0
r49 7 9 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=0.37 $Y=0.085 $X2=0.37
+ $Y2=0.445
r50 2 13 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=1.98
+ $Y=0.235 $X2=2.12 $Y2=0.38
r51 1 9 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.225
+ $Y=0.235 $X2=0.37 $Y2=0.445
.ends

