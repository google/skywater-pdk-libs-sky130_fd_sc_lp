* NGSPICE file created from sky130_fd_sc_lp__einvn_lp.ext - technology: sky130A

.subckt sky130_fd_sc_lp__einvn_lp A TE_B VGND VNB VPB VPWR Z
M1000 a_284_148# a_28_148# VGND VNB nshort w=420000u l=150000u
+  ad=1.365e+11p pd=1.49e+06u as=1.407e+11p ps=1.51e+06u
M1001 VGND TE_B a_115_148# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1002 a_252_414# TE_B VPWR VPB phighvt w=1e+06u l=250000u
+  ad=2.4e+11p pd=2.48e+06u as=2.8e+11p ps=2.56e+06u
M1003 a_115_148# TE_B a_28_148# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1004 VPWR TE_B a_28_148# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=2.85e+11p ps=2.57e+06u
M1005 Z A a_284_148# VNB nshort w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=0p ps=0u
M1006 Z A a_252_414# VPB phighvt w=1e+06u l=250000u
+  ad=2.85e+11p pd=2.57e+06u as=0p ps=0u
.ends

