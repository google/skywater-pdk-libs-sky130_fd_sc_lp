* File: sky130_fd_sc_lp__and4bb_lp.pex.spice
* Created: Fri Aug 28 10:09:35 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__AND4BB_LP%A_N 1 3 6 8 10 11 16
r38 16 18 65.7961 $w=5.35e-07 $l=5.05e-07 $layer=POLY_cond $X=0.687 $Y=0.95
+ $X2=0.687 $Y2=1.455
r39 16 17 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.79
+ $Y=0.95 $X2=0.79 $Y2=0.95
r40 11 17 7.31929 $w=6.68e-07 $l=4.1e-07 $layer=LI1_cond $X=1.2 $Y=1.12 $X2=0.79
+ $Y2=1.12
r41 8 16 31.8222 $w=2.67e-07 $l=2.36525e-07 $layer=POLY_cond $X=0.855 $Y=0.785
+ $X2=0.687 $Y2=0.95
r42 8 10 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.855 $Y=0.785
+ $X2=0.855 $Y2=0.465
r43 6 18 260.876 $w=2.5e-07 $l=1.05e-06 $layer=POLY_cond $X=0.545 $Y=2.505
+ $X2=0.545 $Y2=1.455
r44 1 16 31.8222 $w=2.67e-07 $l=2.61809e-07 $layer=POLY_cond $X=0.495 $Y=0.785
+ $X2=0.687 $Y2=0.95
r45 1 3 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.495 $Y=0.785
+ $X2=0.495 $Y2=0.465
.ends

.subckt PM_SKY130_FD_SC_LP__AND4BB_LP%B_N 3 5 6 9 13 15 19
c49 19 0 1.86394e-19 $X=1.725 $Y=1.29
c50 15 0 4.45047e-20 $X=1.68 $Y=1.295
c51 13 0 1.52904e-19 $X=1.865 $Y=2.545
r52 19 21 23.4306 $w=2.88e-07 $l=1.4e-07 $layer=POLY_cond $X=1.725 $Y=1.29
+ $X2=1.865 $Y2=1.29
r53 17 19 8.36806 $w=2.88e-07 $l=5e-08 $layer=POLY_cond $X=1.675 $Y=1.29
+ $X2=1.725 $Y2=1.29
r54 15 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.725
+ $Y=1.29 $X2=1.725 $Y2=1.29
r55 11 21 6.18571 $w=2.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.865 $Y=1.455
+ $X2=1.865 $Y2=1.29
r56 11 13 270.814 $w=2.5e-07 $l=1.09e-06 $layer=POLY_cond $X=1.865 $Y=1.455
+ $X2=1.865 $Y2=2.545
r57 7 17 18.0107 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.675 $Y=1.125
+ $X2=1.675 $Y2=1.29
r58 7 9 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.675 $Y=1.125
+ $X2=1.675 $Y2=0.465
r59 5 17 30.2662 $w=2.88e-07 $l=1.53542e-07 $layer=POLY_cond $X=1.56 $Y=1.2
+ $X2=1.675 $Y2=1.29
r60 5 6 102.553 $w=1.5e-07 $l=2e-07 $layer=POLY_cond $X=1.56 $Y=1.2 $X2=1.36
+ $Y2=1.2
r61 1 6 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.285 $Y=1.125
+ $X2=1.36 $Y2=1.2
r62 1 3 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.285 $Y=1.125
+ $X2=1.285 $Y2=0.465
.ends

.subckt PM_SKY130_FD_SC_LP__AND4BB_LP%A_27_51# 1 2 7 9 15 18 19 22 26 30 34 38
+ 39 41
c79 34 0 1.07824e-19 $X=2.23 $Y=1.72
c80 18 0 2.30899e-19 $X=2.395 $Y=1.135
c81 7 0 1.08877e-19 $X=2.395 $Y=1.805
r82 38 39 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.395
+ $Y=1.3 $X2=2.395 $Y2=1.3
r83 36 38 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=2.395 $Y=1.635
+ $X2=2.395 $Y2=1.3
r84 35 41 3.80956 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.445 $Y=1.72
+ $X2=0.28 $Y2=1.72
r85 34 36 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.23 $Y=1.72
+ $X2=2.395 $Y2=1.635
r86 34 35 116.455 $w=1.68e-07 $l=1.785e-06 $layer=LI1_cond $X=2.23 $Y=1.72
+ $X2=0.445 $Y2=1.72
r87 30 32 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=0.28 $Y=2.15 $X2=0.28
+ $Y2=2.86
r88 28 41 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.28 $Y=1.805
+ $X2=0.28 $Y2=1.72
r89 28 30 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=0.28 $Y=1.805
+ $X2=0.28 $Y2=2.15
r90 24 41 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.28 $Y=1.635
+ $X2=0.28 $Y2=1.72
r91 24 26 40.3355 $w=3.28e-07 $l=1.155e-06 $layer=LI1_cond $X=0.28 $Y=1.635
+ $X2=0.28 $Y2=0.48
r92 20 22 92.2979 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=2.485 $Y=0.9
+ $X2=2.665 $Y2=0.9
r93 19 39 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.395 $Y=1.64
+ $X2=2.395 $Y2=1.3
r94 18 39 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.395 $Y=1.135
+ $X2=2.395 $Y2=1.3
r95 13 22 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.665 $Y=0.825
+ $X2=2.665 $Y2=0.9
r96 13 15 194.851 $w=1.5e-07 $l=3.8e-07 $layer=POLY_cond $X=2.665 $Y=0.825
+ $X2=2.665 $Y2=0.445
r97 11 20 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.485 $Y=0.975
+ $X2=2.485 $Y2=0.9
r98 11 18 82.0426 $w=1.5e-07 $l=1.6e-07 $layer=POLY_cond $X=2.485 $Y=0.975
+ $X2=2.485 $Y2=1.135
r99 7 19 30.6163 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.395 $Y=1.805
+ $X2=2.395 $Y2=1.64
r100 7 9 183.856 $w=2.5e-07 $l=7.4e-07 $layer=POLY_cond $X=2.395 $Y=1.805
+ $X2=2.395 $Y2=2.545
r101 2 32 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.005 $X2=0.28 $Y2=2.86
r102 2 30 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.005 $X2=0.28 $Y2=2.15
r103 1 26 182 $w=1.7e-07 $l=2.88531e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.255 $X2=0.28 $Y2=0.48
.ends

.subckt PM_SKY130_FD_SC_LP__AND4BB_LP%A_291_409# 1 2 9 13 17 18 21 27 29 30 31
+ 32 36 38 39 40
c100 38 0 1.66554e-19 $X=2.965 $Y=1.38
c101 36 0 1.08877e-19 $X=2.965 $Y=1.72
c102 18 0 1.97298e-19 $X=2.965 $Y=1.885
r103 38 40 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=2.965 $Y=1.38
+ $X2=2.965 $Y2=1.215
r104 38 39 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.965
+ $Y=1.38 $X2=2.965 $Y2=1.38
r105 36 41 14.0725 $w=3.3e-07 $l=3.5e-07 $layer=LI1_cond $X=2.965 $Y=1.72
+ $X2=2.965 $Y2=2.07
r106 36 38 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=2.965 $Y=1.72
+ $X2=2.965 $Y2=1.38
r107 33 40 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=2.885 $Y=0.945
+ $X2=2.885 $Y2=1.215
r108 31 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.8 $Y=0.86
+ $X2=2.885 $Y2=0.945
r109 31 32 48.6043 $w=1.68e-07 $l=7.45e-07 $layer=LI1_cond $X=2.8 $Y=0.86
+ $X2=2.055 $Y2=0.86
r110 29 41 2.50919 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.8 $Y=2.07
+ $X2=2.965 $Y2=2.07
r111 29 30 67.5241 $w=1.68e-07 $l=1.035e-06 $layer=LI1_cond $X=2.8 $Y=2.07
+ $X2=1.765 $Y2=2.07
r112 25 32 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.89 $Y=0.775
+ $X2=2.055 $Y2=0.86
r113 25 27 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.89 $Y=0.775
+ $X2=1.89 $Y2=0.48
r114 21 23 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=1.6 $Y=2.19 $X2=1.6
+ $Y2=2.9
r115 19 30 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.6 $Y=2.155
+ $X2=1.765 $Y2=2.07
r116 19 21 1.22229 $w=3.28e-07 $l=3.5e-08 $layer=LI1_cond $X=1.6 $Y=2.155
+ $X2=1.6 $Y2=2.19
r117 17 39 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.965 $Y=1.72
+ $X2=2.965 $Y2=1.38
r118 17 18 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.965 $Y=1.72
+ $X2=2.965 $Y2=1.885
r119 16 39 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.965 $Y=1.215
+ $X2=2.965 $Y2=1.38
r120 13 16 394.83 $w=1.5e-07 $l=7.7e-07 $layer=POLY_cond $X=3.055 $Y=0.445
+ $X2=3.055 $Y2=1.215
r121 9 18 163.979 $w=2.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.925 $Y=2.545
+ $X2=2.925 $Y2=1.885
r122 2 23 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=1.455
+ $Y=2.045 $X2=1.6 $Y2=2.9
r123 2 21 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=1.455
+ $Y=2.045 $X2=1.6 $Y2=2.19
r124 1 27 182 $w=1.7e-07 $l=2.86575e-07 $layer=licon1_NDIFF $count=1 $X=1.75
+ $Y=0.255 $X2=1.89 $Y2=0.48
.ends

.subckt PM_SKY130_FD_SC_LP__AND4BB_LP%C 3 5 7 11 12 13 17
c54 12 0 8.94739e-20 $X=3.6 $Y=1.295
r55 12 13 12.6936 $w=3.43e-07 $l=3.8e-07 $layer=LI1_cond $X=3.542 $Y=1.285
+ $X2=3.542 $Y2=1.665
r56 12 17 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.535
+ $Y=1.285 $X2=3.535 $Y2=1.285
r57 11 17 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=3.535 $Y=1.625
+ $X2=3.535 $Y2=1.285
r58 10 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.535 $Y=1.12
+ $X2=3.535 $Y2=1.285
r59 5 11 30.6163 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.535 $Y=1.79
+ $X2=3.535 $Y2=1.625
r60 5 7 187.582 $w=2.5e-07 $l=7.55e-07 $layer=POLY_cond $X=3.535 $Y=1.79
+ $X2=3.535 $Y2=2.545
r61 3 10 346.117 $w=1.5e-07 $l=6.75e-07 $layer=POLY_cond $X=3.445 $Y=0.445
+ $X2=3.445 $Y2=1.12
.ends

.subckt PM_SKY130_FD_SC_LP__AND4BB_LP%D 1 3 8 12 15 16 17 18 19 23
c56 23 0 9.23532e-20 $X=4.105 $Y=1.285
c57 18 0 1.86771e-19 $X=4.08 $Y=1.295
c58 8 0 1.02627e-19 $X=4.065 $Y=2.545
r59 18 19 13.2706 $w=3.28e-07 $l=3.8e-07 $layer=LI1_cond $X=4.105 $Y=1.285
+ $X2=4.105 $Y2=1.665
r60 18 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.105
+ $Y=1.285 $X2=4.105 $Y2=1.285
r61 16 23 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=4.105 $Y=1.625
+ $X2=4.105 $Y2=1.285
r62 16 17 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.105 $Y=1.625
+ $X2=4.105 $Y2=1.79
r63 15 23 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.105 $Y=1.12
+ $X2=4.105 $Y2=1.285
r64 10 12 92.2979 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=3.835 $Y=0.805
+ $X2=4.015 $Y2=0.805
r65 8 17 187.582 $w=2.5e-07 $l=7.55e-07 $layer=POLY_cond $X=4.065 $Y=2.545
+ $X2=4.065 $Y2=1.79
r66 4 12 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.015 $Y=0.88
+ $X2=4.015 $Y2=0.805
r67 4 15 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=4.015 $Y=0.88
+ $X2=4.015 $Y2=1.12
r68 1 10 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.835 $Y=0.73
+ $X2=3.835 $Y2=0.805
r69 1 3 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.835 $Y=0.73 $X2=3.835
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__AND4BB_LP%A_461_47# 1 2 3 10 12 15 17 19 24 27 28 34
+ 37 38 39 43 46 48 49 50 51 53 55 56 60 61
c137 55 0 1.52904e-19 $X=2.66 $Y=2.5
c138 50 0 9.23532e-20 $X=4.645 $Y=1.135
c139 27 0 1.0197e-19 $X=4.675 $Y=1.61
c140 15 0 1.86771e-19 $X=4.7 $Y=2.545
r141 59 60 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.675
+ $Y=1.105 $X2=4.675 $Y2=1.105
r142 53 61 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=4.535 $Y=1.97
+ $X2=4.535 $Y2=1.61
r143 51 61 9.49412 $w=3.88e-07 $l=1.95e-07 $layer=LI1_cond $X=4.645 $Y=1.415
+ $X2=4.645 $Y2=1.61
r144 50 59 1.81342 $w=3.9e-07 $l=3e-08 $layer=LI1_cond $X=4.645 $Y=1.135
+ $X2=4.645 $Y2=1.105
r145 50 51 8.27395 $w=3.88e-07 $l=2.8e-07 $layer=LI1_cond $X=4.645 $Y=1.135
+ $X2=4.645 $Y2=1.415
r146 48 53 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.45 $Y=2.055
+ $X2=4.535 $Y2=1.97
r147 48 49 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=4.45 $Y=2.055
+ $X2=3.965 $Y2=2.055
r148 44 56 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.8 $Y=2.505 $X2=3.8
+ $Y2=2.42
r149 44 46 13.7944 $w=3.28e-07 $l=3.95e-07 $layer=LI1_cond $X=3.8 $Y=2.505
+ $X2=3.8 $Y2=2.9
r150 41 56 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.8 $Y=2.335 $X2=3.8
+ $Y2=2.42
r151 41 43 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=3.8 $Y=2.335
+ $X2=3.8 $Y2=2.19
r152 40 49 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.8 $Y=2.14
+ $X2=3.965 $Y2=2.055
r153 40 43 1.74613 $w=3.28e-07 $l=5e-08 $layer=LI1_cond $X=3.8 $Y=2.14 $X2=3.8
+ $Y2=2.19
r154 38 59 10.6272 $w=2.87e-07 $l=3.33542e-07 $layer=LI1_cond $X=4.45 $Y=0.855
+ $X2=4.645 $Y2=1.105
r155 38 39 63.2834 $w=1.68e-07 $l=9.7e-07 $layer=LI1_cond $X=4.45 $Y=0.855
+ $X2=3.48 $Y2=0.855
r156 37 39 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.395 $Y=0.77
+ $X2=3.48 $Y2=0.855
r157 36 37 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=3.395 $Y=0.595
+ $X2=3.395 $Y2=0.77
r158 35 55 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.825 $Y=2.42
+ $X2=2.66 $Y2=2.42
r159 34 56 3.80956 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.635 $Y=2.42
+ $X2=3.8 $Y2=2.42
r160 34 35 52.8449 $w=1.68e-07 $l=8.1e-07 $layer=LI1_cond $X=3.635 $Y=2.42
+ $X2=2.825 $Y2=2.42
r161 28 36 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.31 $Y=0.43
+ $X2=3.395 $Y2=0.595
r162 28 30 30.0334 $w=3.28e-07 $l=8.6e-07 $layer=LI1_cond $X=3.31 $Y=0.43
+ $X2=2.45 $Y2=0.43
r163 26 60 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=4.675 $Y=1.445
+ $X2=4.675 $Y2=1.105
r164 26 27 31.4182 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.675 $Y=1.445
+ $X2=4.675 $Y2=1.61
r165 23 60 39.3438 $w=3.3e-07 $l=2.25e-07 $layer=POLY_cond $X=4.675 $Y=0.88
+ $X2=4.675 $Y2=1.105
r166 23 24 46.1489 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=4.675 $Y=0.805
+ $X2=4.765 $Y2=0.805
r167 20 23 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=4.405 $Y=0.805
+ $X2=4.675 $Y2=0.805
r168 17 24 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.765 $Y=0.73
+ $X2=4.765 $Y2=0.805
r169 17 19 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=4.765 $Y=0.73
+ $X2=4.765 $Y2=0.445
r170 15 27 232.304 $w=2.5e-07 $l=9.35e-07 $layer=POLY_cond $X=4.7 $Y=2.545
+ $X2=4.7 $Y2=1.61
r171 10 20 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.405 $Y=0.73
+ $X2=4.405 $Y2=0.805
r172 10 12 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=4.405 $Y=0.73
+ $X2=4.405 $Y2=0.445
r173 3 46 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=3.66
+ $Y=2.045 $X2=3.8 $Y2=2.9
r174 3 43 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=3.66
+ $Y=2.045 $X2=3.8 $Y2=2.19
r175 2 55 300 $w=1.7e-07 $l=5.20312e-07 $layer=licon1_PDIFF $count=2 $X=2.52
+ $Y=2.045 $X2=2.66 $Y2=2.5
r176 1 30 182 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_NDIFF $count=1 $X=2.305
+ $Y=0.235 $X2=2.45 $Y2=0.43
.ends

.subckt PM_SKY130_FD_SC_LP__AND4BB_LP%VPWR 1 2 3 4 17 23 27 31 34 35 36 38 43 53
+ 54 57 60 63
r67 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r68 60 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r69 57 58 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r70 53 54 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r71 51 54 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=5.04 $Y2=3.33
r72 51 64 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.12 $Y2=3.33
r73 50 51 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r74 48 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.355 $Y=3.33
+ $X2=3.19 $Y2=3.33
r75 48 50 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=3.355 $Y=3.33
+ $X2=4.08 $Y2=3.33
r76 44 60 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.295 $Y=3.33
+ $X2=2.13 $Y2=3.33
r77 44 46 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=2.295 $Y=3.33
+ $X2=2.64 $Y2=3.33
r78 43 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.025 $Y=3.33
+ $X2=3.19 $Y2=3.33
r79 43 46 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=3.025 $Y=3.33
+ $X2=2.64 $Y2=3.33
r80 42 61 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r81 42 58 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.72 $Y2=3.33
r82 41 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r83 39 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.975 $Y=3.33
+ $X2=0.81 $Y2=3.33
r84 39 41 45.9947 $w=1.68e-07 $l=7.05e-07 $layer=LI1_cond $X=0.975 $Y=3.33
+ $X2=1.68 $Y2=3.33
r85 38 60 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.965 $Y=3.33
+ $X2=2.13 $Y2=3.33
r86 38 41 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.965 $Y=3.33
+ $X2=1.68 $Y2=3.33
r87 36 64 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r88 36 61 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r89 36 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r90 34 50 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=4.165 $Y=3.33
+ $X2=4.08 $Y2=3.33
r91 34 35 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.165 $Y=3.33
+ $X2=4.33 $Y2=3.33
r92 33 53 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=4.495 $Y=3.33
+ $X2=5.04 $Y2=3.33
r93 33 35 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.495 $Y=3.33
+ $X2=4.33 $Y2=3.33
r94 29 35 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.33 $Y=3.245
+ $X2=4.33 $Y2=3.33
r95 29 31 26.5411 $w=3.28e-07 $l=7.6e-07 $layer=LI1_cond $X=4.33 $Y=3.245
+ $X2=4.33 $Y2=2.485
r96 25 63 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.19 $Y=3.245
+ $X2=3.19 $Y2=3.33
r97 25 27 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=3.19 $Y=3.245
+ $X2=3.19 $Y2=2.875
r98 21 60 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.13 $Y=3.245
+ $X2=2.13 $Y2=3.33
r99 21 23 26.0173 $w=3.28e-07 $l=7.45e-07 $layer=LI1_cond $X=2.13 $Y=3.245
+ $X2=2.13 $Y2=2.5
r100 17 20 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=0.81 $Y=2.15
+ $X2=0.81 $Y2=2.86
r101 15 57 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.81 $Y=3.245
+ $X2=0.81 $Y2=3.33
r102 15 20 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=0.81 $Y=3.245
+ $X2=0.81 $Y2=2.86
r103 4 31 300 $w=1.7e-07 $l=5.05173e-07 $layer=licon1_PDIFF $count=2 $X=4.19
+ $Y=2.045 $X2=4.33 $Y2=2.485
r104 3 27 600 $w=1.7e-07 $l=8.97274e-07 $layer=licon1_PDIFF $count=1 $X=3.05
+ $Y=2.045 $X2=3.19 $Y2=2.875
r105 2 23 300 $w=1.7e-07 $l=5.20312e-07 $layer=licon1_PDIFF $count=2 $X=1.99
+ $Y=2.045 $X2=2.13 $Y2=2.5
r106 1 20 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=0.67
+ $Y=2.005 $X2=0.81 $Y2=2.86
r107 1 17 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.67
+ $Y=2.005 $X2=0.81 $Y2=2.15
.ends

.subckt PM_SKY130_FD_SC_LP__AND4BB_LP%X 1 2 12 14 15 16 32 34
c25 14 0 2.04597e-19 $X=4.955 $Y=1.95
r26 21 34 2.36399 $w=3.88e-07 $l=8e-08 $layer=LI1_cond $X=4.995 $Y=2.115
+ $X2=4.995 $Y2=2.035
r27 16 29 3.69373 $w=3.88e-07 $l=1.25e-07 $layer=LI1_cond $X=4.995 $Y=2.775
+ $X2=4.995 $Y2=2.9
r28 15 16 10.9334 $w=3.88e-07 $l=3.7e-07 $layer=LI1_cond $X=4.995 $Y=2.405
+ $X2=4.995 $Y2=2.775
r29 14 34 0.0886495 $w=3.88e-07 $l=3e-09 $layer=LI1_cond $X=4.995 $Y=2.032
+ $X2=4.995 $Y2=2.035
r30 14 32 7.04148 $w=3.88e-07 $l=1.12e-07 $layer=LI1_cond $X=4.995 $Y=2.032
+ $X2=4.995 $Y2=1.92
r31 14 15 8.51035 $w=3.88e-07 $l=2.88e-07 $layer=LI1_cond $X=4.995 $Y=2.117
+ $X2=4.995 $Y2=2.405
r32 14 21 0.0590996 $w=3.88e-07 $l=2e-09 $layer=LI1_cond $X=4.995 $Y=2.117
+ $X2=4.995 $Y2=2.115
r33 10 12 3.51355 $w=4.08e-07 $l=1.25e-07 $layer=LI1_cond $X=4.98 $Y=0.47
+ $X2=5.105 $Y2=0.47
r34 7 12 5.92876 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=5.105 $Y=0.675
+ $X2=5.105 $Y2=0.47
r35 7 32 81.2246 $w=1.68e-07 $l=1.245e-06 $layer=LI1_cond $X=5.105 $Y=0.675
+ $X2=5.105 $Y2=1.92
r36 2 29 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=4.825
+ $Y=2.045 $X2=4.965 $Y2=2.9
r37 2 14 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=4.825
+ $Y=2.045 $X2=4.965 $Y2=2.19
r38 1 10 182 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=1 $X=4.84
+ $Y=0.235 $X2=4.98 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_LP__AND4BB_LP%VGND 1 2 9 13 15 17 22 29 30 33 36
r63 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r64 33 34 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r65 30 37 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=4.08
+ $Y2=0
r66 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r67 27 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.215 $Y=0 $X2=4.05
+ $Y2=0
r68 27 29 53.8235 $w=1.68e-07 $l=8.25e-07 $layer=LI1_cond $X=4.215 $Y=0 $X2=5.04
+ $Y2=0
r69 26 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r70 25 26 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r71 23 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.235 $Y=0 $X2=1.07
+ $Y2=0
r72 23 25 154.294 $w=1.68e-07 $l=2.365e-06 $layer=LI1_cond $X=1.235 $Y=0 $X2=3.6
+ $Y2=0
r73 22 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.885 $Y=0 $X2=4.05
+ $Y2=0
r74 22 25 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=3.885 $Y=0 $X2=3.6
+ $Y2=0
r75 20 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r76 19 20 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r77 17 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.905 $Y=0 $X2=1.07
+ $Y2=0
r78 17 19 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=0.905 $Y=0 $X2=0.72
+ $Y2=0
r79 15 26 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r80 15 34 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=2.64 $Y=0 $X2=1.2
+ $Y2=0
r81 11 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.05 $Y=0.085
+ $X2=4.05 $Y2=0
r82 11 13 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=4.05 $Y=0.085
+ $X2=4.05 $Y2=0.4
r83 7 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.07 $Y=0.085 $X2=1.07
+ $Y2=0
r84 7 9 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=1.07 $Y=0.085 $X2=1.07
+ $Y2=0.42
r85 2 13 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=3.91
+ $Y=0.235 $X2=4.05 $Y2=0.4
r86 1 9 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=0.93
+ $Y=0.255 $X2=1.07 $Y2=0.42
.ends

