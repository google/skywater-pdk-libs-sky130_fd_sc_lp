* File: sky130_fd_sc_lp__o211ai_4.pxi.spice
* Created: Fri Aug 28 11:03:09 2020
* 
x_PM_SKY130_FD_SC_LP__O211AI_4%A1 N_A1_M1010_g N_A1_M1004_g N_A1_M1020_g
+ N_A1_M1005_g N_A1_M1027_g N_A1_M1013_g N_A1_M1031_g N_A1_M1028_g N_A1_c_122_n
+ N_A1_c_123_n N_A1_c_145_p N_A1_c_159_p N_A1_c_124_n N_A1_c_125_n A1 A1 A1 A1
+ A1 A1 N_A1_c_126_n N_A1_c_127_n N_A1_c_136_p PM_SKY130_FD_SC_LP__O211AI_4%A1
x_PM_SKY130_FD_SC_LP__O211AI_4%A2 N_A2_M1006_g N_A2_c_243_n N_A2_M1011_g
+ N_A2_M1008_g N_A2_c_244_n N_A2_M1018_g N_A2_M1017_g N_A2_c_245_n N_A2_M1021_g
+ N_A2_M1023_g N_A2_c_246_n N_A2_M1025_g A2 A2 A2 N_A2_c_242_n
+ PM_SKY130_FD_SC_LP__O211AI_4%A2
x_PM_SKY130_FD_SC_LP__O211AI_4%B1 N_B1_M1001_g N_B1_M1000_g N_B1_M1002_g
+ N_B1_M1007_g N_B1_M1014_g N_B1_M1026_g N_B1_M1030_g N_B1_M1015_g N_B1_c_321_n
+ N_B1_c_330_n N_B1_c_346_p N_B1_c_384_p N_B1_c_331_n N_B1_c_322_n B1 B1 B1
+ N_B1_c_324_n PM_SKY130_FD_SC_LP__O211AI_4%B1
x_PM_SKY130_FD_SC_LP__O211AI_4%C1 N_C1_M1009_g N_C1_M1003_g N_C1_M1012_g
+ N_C1_M1016_g N_C1_M1019_g N_C1_M1022_g N_C1_M1029_g N_C1_M1024_g C1 C1 C1 C1
+ N_C1_c_447_n PM_SKY130_FD_SC_LP__O211AI_4%C1
x_PM_SKY130_FD_SC_LP__O211AI_4%VPWR N_VPWR_M1004_s N_VPWR_M1005_s N_VPWR_M1031_s
+ N_VPWR_M1007_s N_VPWR_M1009_s N_VPWR_M1019_s N_VPWR_M1030_s N_VPWR_c_521_n
+ N_VPWR_c_522_n N_VPWR_c_523_n N_VPWR_c_524_n N_VPWR_c_525_n N_VPWR_c_526_n
+ N_VPWR_c_527_n N_VPWR_c_528_n N_VPWR_c_529_n N_VPWR_c_530_n N_VPWR_c_531_n
+ N_VPWR_c_532_n N_VPWR_c_533_n N_VPWR_c_534_n VPWR N_VPWR_c_535_n
+ N_VPWR_c_536_n N_VPWR_c_537_n N_VPWR_c_520_n N_VPWR_c_539_n N_VPWR_c_540_n
+ N_VPWR_c_541_n PM_SKY130_FD_SC_LP__O211AI_4%VPWR
x_PM_SKY130_FD_SC_LP__O211AI_4%A_140_367# N_A_140_367#_M1004_d
+ N_A_140_367#_M1013_d N_A_140_367#_M1018_d N_A_140_367#_M1025_d
+ N_A_140_367#_c_645_n N_A_140_367#_c_655_n N_A_140_367#_c_660_n
+ N_A_140_367#_c_673_n N_A_140_367#_c_675_n N_A_140_367#_c_683_p
+ N_A_140_367#_c_661_n PM_SKY130_FD_SC_LP__O211AI_4%A_140_367#
x_PM_SKY130_FD_SC_LP__O211AI_4%Y N_Y_M1003_s N_Y_M1022_s N_Y_M1011_s N_Y_M1021_s
+ N_Y_M1000_d N_Y_M1026_d N_Y_M1012_d N_Y_M1029_d N_Y_c_694_n N_Y_c_709_n
+ N_Y_c_711_n N_Y_c_716_n N_Y_c_686_n N_Y_c_759_n N_Y_c_687_n N_Y_c_761_n
+ N_Y_c_688_n N_Y_c_698_n N_Y_c_763_n N_Y_c_726_n N_Y_c_689_n N_Y_c_729_n
+ N_Y_c_730_n N_Y_c_691_n Y Y Y Y PM_SKY130_FD_SC_LP__O211AI_4%Y
x_PM_SKY130_FD_SC_LP__O211AI_4%A_57_47# N_A_57_47#_M1010_s N_A_57_47#_M1020_s
+ N_A_57_47#_M1006_s N_A_57_47#_M1017_s N_A_57_47#_M1028_s N_A_57_47#_M1002_s
+ N_A_57_47#_M1015_s N_A_57_47#_c_878_p N_A_57_47#_c_790_n N_A_57_47#_c_791_n
+ N_A_57_47#_c_867_p N_A_57_47#_c_792_n N_A_57_47#_c_868_p N_A_57_47#_c_793_n
+ N_A_57_47#_c_866_p N_A_57_47#_c_794_n N_A_57_47#_c_869_p N_A_57_47#_c_795_n
+ N_A_57_47#_c_835_n N_A_57_47#_c_836_n N_A_57_47#_c_837_n N_A_57_47#_c_796_n
+ N_A_57_47#_c_797_n N_A_57_47#_c_798_n N_A_57_47#_c_799_n N_A_57_47#_c_800_n
+ PM_SKY130_FD_SC_LP__O211AI_4%A_57_47#
x_PM_SKY130_FD_SC_LP__O211AI_4%VGND N_VGND_M1010_d N_VGND_M1027_d N_VGND_M1008_d
+ N_VGND_M1023_d N_VGND_c_895_n N_VGND_c_896_n N_VGND_c_897_n N_VGND_c_898_n
+ N_VGND_c_899_n N_VGND_c_900_n VGND N_VGND_c_901_n N_VGND_c_902_n
+ N_VGND_c_903_n N_VGND_c_904_n N_VGND_c_905_n N_VGND_c_906_n N_VGND_c_907_n
+ PM_SKY130_FD_SC_LP__O211AI_4%VGND
x_PM_SKY130_FD_SC_LP__O211AI_4%A_836_47# N_A_836_47#_M1001_d N_A_836_47#_M1014_d
+ N_A_836_47#_M1016_d N_A_836_47#_M1024_d N_A_836_47#_c_991_n
+ N_A_836_47#_c_995_n PM_SKY130_FD_SC_LP__O211AI_4%A_836_47#
cc_1 VNB N_A1_M1010_g 0.0284365f $X=-0.19 $Y=-0.245 $X2=0.625 $Y2=0.655
cc_2 VNB N_A1_M1004_g 0.0021209f $X=-0.19 $Y=-0.245 $X2=0.625 $Y2=2.465
cc_3 VNB N_A1_M1020_g 0.0207302f $X=-0.19 $Y=-0.245 $X2=1.055 $Y2=0.655
cc_4 VNB N_A1_M1005_g 0.00123474f $X=-0.19 $Y=-0.245 $X2=1.055 $Y2=2.465
cc_5 VNB N_A1_M1027_g 0.0209507f $X=-0.19 $Y=-0.245 $X2=1.485 $Y2=0.655
cc_6 VNB N_A1_M1013_g 0.00125594f $X=-0.19 $Y=-0.245 $X2=1.485 $Y2=2.465
cc_7 VNB N_A1_M1028_g 0.0245991f $X=-0.19 $Y=-0.245 $X2=3.645 $Y2=0.655
cc_8 VNB N_A1_c_122_n 0.0192323f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.487
cc_9 VNB N_A1_c_123_n 0.00256364f $X=-0.19 $Y=-0.245 $X2=1.337 $Y2=1.63
cc_10 VNB N_A1_c_124_n 0.00120154f $X=-0.19 $Y=-0.245 $X2=3.655 $Y2=1.51
cc_11 VNB N_A1_c_125_n 0.0260373f $X=-0.19 $Y=-0.245 $X2=3.655 $Y2=1.51
cc_12 VNB N_A1_c_126_n 0.042941f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=1.46
cc_13 VNB N_A1_c_127_n 0.0505289f $X=-0.19 $Y=-0.245 $X2=1.485 $Y2=1.46
cc_14 VNB N_A2_M1006_g 0.0235785f $X=-0.19 $Y=-0.245 $X2=0.625 $Y2=0.655
cc_15 VNB N_A2_M1008_g 0.023273f $X=-0.19 $Y=-0.245 $X2=1.055 $Y2=0.655
cc_16 VNB N_A2_M1017_g 0.023273f $X=-0.19 $Y=-0.245 $X2=1.485 $Y2=1.295
cc_17 VNB N_A2_M1023_g 0.0237353f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB A2 0.0019354f $X=-0.19 $Y=-0.245 $X2=3.645 $Y2=0.655
cc_19 VNB N_A2_c_242_n 0.0645734f $X=-0.19 $Y=-0.245 $X2=3.655 $Y2=1.51
cc_20 VNB N_B1_M1001_g 0.0242801f $X=-0.19 $Y=-0.245 $X2=0.625 $Y2=0.655
cc_21 VNB N_B1_M1002_g 0.0234721f $X=-0.19 $Y=-0.245 $X2=1.055 $Y2=0.655
cc_22 VNB N_B1_M1014_g 0.0287886f $X=-0.19 $Y=-0.245 $X2=1.485 $Y2=0.655
cc_23 VNB N_B1_M1015_g 0.0257974f $X=-0.19 $Y=-0.245 $X2=3.645 $Y2=0.655
cc_24 VNB N_B1_c_321_n 0.00383433f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.487
cc_25 VNB N_B1_c_322_n 0.0301585f $X=-0.19 $Y=-0.245 $X2=0.715 $Y2=1.46
cc_26 VNB B1 0.00261207f $X=-0.19 $Y=-0.245 $X2=3.64 $Y2=1.51
cc_27 VNB N_B1_c_324_n 0.0453212f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_C1_M1003_g 0.0210171f $X=-0.19 $Y=-0.245 $X2=0.625 $Y2=2.465
cc_29 VNB N_C1_M1016_g 0.0198617f $X=-0.19 $Y=-0.245 $X2=1.055 $Y2=2.465
cc_30 VNB N_C1_M1022_g 0.0198617f $X=-0.19 $Y=-0.245 $X2=1.485 $Y2=2.465
cc_31 VNB N_C1_M1024_g 0.020008f $X=-0.19 $Y=-0.245 $X2=3.645 $Y2=0.655
cc_32 VNB N_C1_c_447_n 0.0922966f $X=-0.19 $Y=-0.245 $X2=3.515 $Y2=1.95
cc_33 VNB N_VPWR_c_520_n 0.342803f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_Y_c_686_n 0.00687867f $X=-0.19 $Y=-0.245 $X2=1.337 $Y2=1.63
cc_35 VNB N_Y_c_687_n 0.0196201f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.95
cc_36 VNB N_Y_c_688_n 0.0191582f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_Y_c_689_n 0.00101109f $X=-0.19 $Y=-0.245 $X2=1.055 $Y2=1.46
cc_38 VNB N_A_57_47#_c_790_n 0.00290783f $X=-0.19 $Y=-0.245 $X2=3.635 $Y2=2.465
cc_39 VNB N_A_57_47#_c_791_n 0.00549523f $X=-0.19 $Y=-0.245 $X2=3.635 $Y2=2.465
cc_40 VNB N_A_57_47#_c_792_n 0.0105569f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_57_47#_c_793_n 0.00352066f $X=-0.19 $Y=-0.245 $X2=0.715 $Y2=1.487
cc_42 VNB N_A_57_47#_c_794_n 0.00725601f $X=-0.19 $Y=-0.245 $X2=3.64 $Y2=1.51
cc_43 VNB N_A_57_47#_c_795_n 0.00494069f $X=-0.19 $Y=-0.245 $X2=1.395 $Y2=1.46
cc_44 VNB N_A_57_47#_c_796_n 0.00144427f $X=-0.19 $Y=-0.245 $X2=3.515 $Y2=1.95
cc_45 VNB N_A_57_47#_c_797_n 0.0016721f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_57_47#_c_798_n 0.0016721f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_57_47#_c_799_n 0.00623654f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_57_47#_c_800_n 0.0208484f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=1.46
cc_49 VNB N_VGND_c_895_n 3.99129e-19 $X=-0.19 $Y=-0.245 $X2=1.485 $Y2=1.295
cc_50 VNB N_VGND_c_896_n 3.0911e-19 $X=-0.19 $Y=-0.245 $X2=1.485 $Y2=1.625
cc_51 VNB N_VGND_c_897_n 3.0911e-19 $X=-0.19 $Y=-0.245 $X2=3.635 $Y2=1.675
cc_52 VNB N_VGND_c_898_n 3.99129e-19 $X=-0.19 $Y=-0.245 $X2=3.645 $Y2=1.345
cc_53 VNB N_VGND_c_899_n 0.0129398f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_900_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.487
cc_55 VNB N_VGND_c_901_n 0.0129398f $X=-0.19 $Y=-0.245 $X2=0.375 $Y2=1.46
cc_56 VNB N_VGND_c_902_n 0.0129398f $X=-0.19 $Y=-0.245 $X2=1.337 $Y2=1.63
cc_57 VNB N_VGND_c_903_n 0.110093f $X=-0.19 $Y=-0.245 $X2=2.555 $Y2=1.95
cc_58 VNB N_VGND_c_904_n 0.405913f $X=-0.19 $Y=-0.245 $X2=3.035 $Y2=1.95
cc_59 VNB N_VGND_c_905_n 0.0251082f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_906_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_907_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0.375 $Y2=1.46
cc_62 VNB N_A_836_47#_c_991_n 0.00754019f $X=-0.19 $Y=-0.245 $X2=1.485 $Y2=1.625
cc_63 VPB N_A1_M1004_g 0.0272589f $X=-0.19 $Y=1.655 $X2=0.625 $Y2=2.465
cc_64 VPB N_A1_M1005_g 0.0188433f $X=-0.19 $Y=1.655 $X2=1.055 $Y2=2.465
cc_65 VPB N_A1_M1013_g 0.0191608f $X=-0.19 $Y=1.655 $X2=1.485 $Y2=2.465
cc_66 VPB N_A1_M1031_g 0.0177081f $X=-0.19 $Y=1.655 $X2=3.635 $Y2=2.465
cc_67 VPB N_A1_c_124_n 0.0027229f $X=-0.19 $Y=1.655 $X2=3.655 $Y2=1.51
cc_68 VPB N_A1_c_125_n 0.00663035f $X=-0.19 $Y=1.655 $X2=3.655 $Y2=1.51
cc_69 VPB N_A2_c_243_n 0.0163296f $X=-0.19 $Y=1.655 $X2=0.625 $Y2=1.625
cc_70 VPB N_A2_c_244_n 0.0160131f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_71 VPB N_A2_c_245_n 0.016012f $X=-0.19 $Y=1.655 $X2=1.485 $Y2=0.655
cc_72 VPB N_A2_c_246_n 0.0161953f $X=-0.19 $Y=1.655 $X2=3.635 $Y2=2.465
cc_73 VPB A2 0.00892978f $X=-0.19 $Y=1.655 $X2=3.645 $Y2=0.655
cc_74 VPB N_A2_c_242_n 0.0215314f $X=-0.19 $Y=1.655 $X2=3.655 $Y2=1.51
cc_75 VPB N_B1_M1000_g 0.0184222f $X=-0.19 $Y=1.655 $X2=0.625 $Y2=2.465
cc_76 VPB N_B1_M1007_g 0.0178289f $X=-0.19 $Y=1.655 $X2=1.055 $Y2=2.465
cc_77 VPB N_B1_M1026_g 0.0175527f $X=-0.19 $Y=1.655 $X2=1.485 $Y2=2.465
cc_78 VPB N_B1_M1030_g 0.0225752f $X=-0.19 $Y=1.655 $X2=3.635 $Y2=2.465
cc_79 VPB N_B1_c_321_n 7.11043e-19 $X=-0.19 $Y=1.655 $X2=1.115 $Y2=1.487
cc_80 VPB N_B1_c_330_n 7.2292e-19 $X=-0.19 $Y=1.655 $X2=0.375 $Y2=1.487
cc_81 VPB N_B1_c_331_n 0.00148678f $X=-0.19 $Y=1.655 $X2=0.715 $Y2=1.46
cc_82 VPB N_B1_c_322_n 0.00777567f $X=-0.19 $Y=1.655 $X2=0.715 $Y2=1.46
cc_83 VPB B1 0.00904201f $X=-0.19 $Y=1.655 $X2=3.64 $Y2=1.51
cc_84 VPB N_B1_c_324_n 0.00833062f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_85 VPB N_C1_M1009_g 0.0186861f $X=-0.19 $Y=1.655 $X2=0.625 $Y2=0.655
cc_86 VPB N_C1_M1012_g 0.0180356f $X=-0.19 $Y=1.655 $X2=1.055 $Y2=0.655
cc_87 VPB N_C1_M1019_g 0.0206874f $X=-0.19 $Y=1.655 $X2=1.485 $Y2=0.655
cc_88 VPB N_C1_M1029_g 0.0213329f $X=-0.19 $Y=1.655 $X2=3.635 $Y2=2.465
cc_89 VPB C1 0.0109678f $X=-0.19 $Y=1.655 $X2=0.375 $Y2=1.46
cc_90 VPB N_C1_c_447_n 0.0228423f $X=-0.19 $Y=1.655 $X2=3.515 $Y2=1.95
cc_91 VPB N_VPWR_c_521_n 0.0155683f $X=-0.19 $Y=1.655 $X2=1.485 $Y2=2.465
cc_92 VPB N_VPWR_c_522_n 0.0554469f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_93 VPB N_VPWR_c_523_n 4.06069e-19 $X=-0.19 $Y=1.655 $X2=3.645 $Y2=0.655
cc_94 VPB N_VPWR_c_524_n 4.02668e-19 $X=-0.19 $Y=1.655 $X2=0.375 $Y2=1.487
cc_95 VPB N_VPWR_c_525_n 3.18751e-19 $X=-0.19 $Y=1.655 $X2=0.715 $Y2=1.487
cc_96 VPB N_VPWR_c_526_n 0.0147711f $X=-0.19 $Y=1.655 $X2=0.715 $Y2=1.46
cc_97 VPB N_VPWR_c_527_n 0.00387954f $X=-0.19 $Y=1.655 $X2=3.64 $Y2=1.51
cc_98 VPB N_VPWR_c_528_n 0.0191368f $X=-0.19 $Y=1.655 $X2=1.337 $Y2=1.487
cc_99 VPB N_VPWR_c_529_n 0.0515153f $X=-0.19 $Y=1.655 $X2=1.115 $Y2=1.95
cc_100 VPB N_VPWR_c_530_n 0.00436868f $X=-0.19 $Y=1.655 $X2=1.595 $Y2=1.95
cc_101 VPB N_VPWR_c_531_n 0.0133881f $X=-0.19 $Y=1.655 $X2=2.075 $Y2=1.95
cc_102 VPB N_VPWR_c_532_n 0.00436868f $X=-0.19 $Y=1.655 $X2=2.555 $Y2=1.95
cc_103 VPB N_VPWR_c_533_n 0.0129657f $X=-0.19 $Y=1.655 $X2=3.515 $Y2=1.95
cc_104 VPB N_VPWR_c_534_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_105 VPB N_VPWR_c_535_n 0.0149772f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_106 VPB N_VPWR_c_536_n 0.0150084f $X=-0.19 $Y=1.655 $X2=3.5 $Y2=2.022
cc_107 VPB N_VPWR_c_537_n 0.0124854f $X=-0.19 $Y=1.655 $X2=1.337 $Y2=2.022
cc_108 VPB N_VPWR_c_520_n 0.0534729f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_109 VPB N_VPWR_c_539_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_110 VPB N_VPWR_c_540_n 0.0047828f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_111 VPB N_VPWR_c_541_n 0.0122104f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_112 VPB N_A_140_367#_c_645_n 0.00216024f $X=-0.19 $Y=1.655 $X2=1.055
+ $Y2=2.465
cc_113 VPB N_Y_c_688_n 0.0300903f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_114 VPB N_Y_c_691_n 0.0202062f $X=-0.19 $Y=1.655 $X2=3.655 $Y2=1.345
cc_115 N_A1_M1027_g N_A2_M1006_g 0.0259842f $X=1.485 $Y=0.655 $X2=0 $Y2=0
cc_116 N_A1_M1013_g N_A2_c_243_n 0.0259842f $X=1.485 $Y=2.465 $X2=0 $Y2=0
cc_117 N_A1_c_136_p N_A2_c_243_n 0.0165846f $X=3.5 $Y=2.022 $X2=0 $Y2=0
cc_118 N_A1_c_136_p N_A2_c_244_n 0.0114985f $X=3.5 $Y=2.022 $X2=0 $Y2=0
cc_119 N_A1_c_136_p N_A2_c_245_n 0.0114985f $X=3.5 $Y=2.022 $X2=0 $Y2=0
cc_120 N_A1_M1028_g N_A2_M1023_g 0.0250747f $X=3.645 $Y=0.655 $X2=0 $Y2=0
cc_121 N_A1_c_124_n N_A2_c_246_n 0.0037593f $X=3.655 $Y=1.51 $X2=0 $Y2=0
cc_122 N_A1_c_136_p N_A2_c_246_n 0.011445f $X=3.5 $Y=2.022 $X2=0 $Y2=0
cc_123 N_A1_M1013_g A2 3.88715e-19 $X=1.485 $Y=2.465 $X2=0 $Y2=0
cc_124 N_A1_M1031_g A2 2.57243e-19 $X=3.635 $Y=2.465 $X2=0 $Y2=0
cc_125 N_A1_c_123_n A2 0.0110419f $X=1.337 $Y=1.63 $X2=0 $Y2=0
cc_126 N_A1_c_145_p A2 0.00618362f $X=1.337 $Y=1.925 $X2=0 $Y2=0
cc_127 N_A1_c_124_n A2 0.0272336f $X=3.655 $Y=1.51 $X2=0 $Y2=0
cc_128 N_A1_c_125_n A2 0.00155774f $X=3.655 $Y=1.51 $X2=0 $Y2=0
cc_129 N_A1_c_127_n A2 2.50929e-19 $X=1.485 $Y=1.46 $X2=0 $Y2=0
cc_130 N_A1_c_136_p A2 0.0954675f $X=3.5 $Y=2.022 $X2=0 $Y2=0
cc_131 N_A1_M1031_g N_A2_c_242_n 0.0538749f $X=3.635 $Y=2.465 $X2=0 $Y2=0
cc_132 N_A1_c_123_n N_A2_c_242_n 0.0015237f $X=1.337 $Y=1.63 $X2=0 $Y2=0
cc_133 N_A1_c_145_p N_A2_c_242_n 0.00160411f $X=1.337 $Y=1.925 $X2=0 $Y2=0
cc_134 N_A1_c_124_n N_A2_c_242_n 0.00110395f $X=3.655 $Y=1.51 $X2=0 $Y2=0
cc_135 N_A1_c_125_n N_A2_c_242_n 0.021402f $X=3.655 $Y=1.51 $X2=0 $Y2=0
cc_136 N_A1_c_127_n N_A2_c_242_n 0.0259842f $X=1.485 $Y=1.46 $X2=0 $Y2=0
cc_137 N_A1_c_136_p N_A2_c_242_n 0.00197832f $X=3.5 $Y=2.022 $X2=0 $Y2=0
cc_138 N_A1_M1028_g N_B1_M1001_g 0.0212431f $X=3.645 $Y=0.655 $X2=0 $Y2=0
cc_139 N_A1_M1031_g N_B1_M1000_g 0.0433281f $X=3.635 $Y=2.465 $X2=0 $Y2=0
cc_140 N_A1_c_159_p N_B1_M1000_g 0.00189179f $X=3.64 $Y=1.925 $X2=0 $Y2=0
cc_141 N_A1_c_124_n N_B1_M1000_g 0.00372471f $X=3.655 $Y=1.51 $X2=0 $Y2=0
cc_142 N_A1_M1031_g B1 2.93401e-19 $X=3.635 $Y=2.465 $X2=0 $Y2=0
cc_143 N_A1_c_124_n B1 0.0347784f $X=3.655 $Y=1.51 $X2=0 $Y2=0
cc_144 N_A1_c_125_n B1 0.00218633f $X=3.655 $Y=1.51 $X2=0 $Y2=0
cc_145 N_A1_c_124_n N_B1_c_324_n 3.2456e-19 $X=3.655 $Y=1.51 $X2=0 $Y2=0
cc_146 N_A1_c_125_n N_B1_c_324_n 0.0206161f $X=3.655 $Y=1.51 $X2=0 $Y2=0
cc_147 N_A1_c_145_p N_VPWR_M1005_s 0.00184152f $X=1.337 $Y=1.925 $X2=0 $Y2=0
cc_148 N_A1_c_159_p N_VPWR_M1031_s 0.00275169f $X=3.64 $Y=1.925 $X2=0 $Y2=0
cc_149 N_A1_c_124_n N_VPWR_M1031_s 0.00116461f $X=3.655 $Y=1.51 $X2=0 $Y2=0
cc_150 N_A1_M1004_g N_VPWR_c_522_n 0.0076281f $X=0.625 $Y=2.465 $X2=0 $Y2=0
cc_151 N_A1_c_122_n N_VPWR_c_522_n 0.0237411f $X=1.115 $Y=1.487 $X2=0 $Y2=0
cc_152 N_A1_c_126_n N_VPWR_c_522_n 0.00222894f $X=0.55 $Y=1.46 $X2=0 $Y2=0
cc_153 N_A1_M1004_g N_VPWR_c_523_n 5.81037e-19 $X=0.625 $Y=2.465 $X2=0 $Y2=0
cc_154 N_A1_M1005_g N_VPWR_c_523_n 0.00942207f $X=1.055 $Y=2.465 $X2=0 $Y2=0
cc_155 N_A1_M1013_g N_VPWR_c_523_n 0.0104125f $X=1.485 $Y=2.465 $X2=0 $Y2=0
cc_156 N_A1_M1031_g N_VPWR_c_524_n 0.00942951f $X=3.635 $Y=2.465 $X2=0 $Y2=0
cc_157 N_A1_M1013_g N_VPWR_c_529_n 0.00486043f $X=1.485 $Y=2.465 $X2=0 $Y2=0
cc_158 N_A1_M1031_g N_VPWR_c_529_n 0.00564095f $X=3.635 $Y=2.465 $X2=0 $Y2=0
cc_159 N_A1_M1004_g N_VPWR_c_535_n 0.00585385f $X=0.625 $Y=2.465 $X2=0 $Y2=0
cc_160 N_A1_M1005_g N_VPWR_c_535_n 0.00486043f $X=1.055 $Y=2.465 $X2=0 $Y2=0
cc_161 N_A1_M1004_g N_VPWR_c_520_n 0.0115829f $X=0.625 $Y=2.465 $X2=0 $Y2=0
cc_162 N_A1_M1005_g N_VPWR_c_520_n 0.00447879f $X=1.055 $Y=2.465 $X2=0 $Y2=0
cc_163 N_A1_M1013_g N_VPWR_c_520_n 0.00450413f $X=1.485 $Y=2.465 $X2=0 $Y2=0
cc_164 N_A1_M1031_g N_VPWR_c_520_n 0.00524073f $X=3.635 $Y=2.465 $X2=0 $Y2=0
cc_165 N_A1_c_136_p N_A_140_367#_M1013_d 0.00821203f $X=3.5 $Y=2.022 $X2=0 $Y2=0
cc_166 N_A1_c_136_p N_A_140_367#_M1018_d 0.00334999f $X=3.5 $Y=2.022 $X2=0 $Y2=0
cc_167 N_A1_c_124_n N_A_140_367#_M1025_d 0.00113684f $X=3.655 $Y=1.51 $X2=0
+ $Y2=0
cc_168 N_A1_c_136_p N_A_140_367#_M1025_d 0.00778195f $X=3.5 $Y=2.022 $X2=0 $Y2=0
cc_169 N_A1_M1004_g N_A_140_367#_c_645_n 4.83072e-19 $X=0.625 $Y=2.465 $X2=0
+ $Y2=0
cc_170 N_A1_M1005_g N_A_140_367#_c_645_n 4.40781e-19 $X=1.055 $Y=2.465 $X2=0
+ $Y2=0
cc_171 N_A1_c_122_n N_A_140_367#_c_645_n 0.0179731f $X=1.115 $Y=1.487 $X2=0
+ $Y2=0
cc_172 N_A1_c_145_p N_A_140_367#_c_645_n 0.0046037f $X=1.337 $Y=1.925 $X2=0
+ $Y2=0
cc_173 N_A1_c_127_n N_A_140_367#_c_645_n 7.73936e-19 $X=1.485 $Y=1.46 $X2=0
+ $Y2=0
cc_174 N_A1_M1005_g N_A_140_367#_c_655_n 0.0133285f $X=1.055 $Y=2.465 $X2=0
+ $Y2=0
cc_175 N_A1_M1013_g N_A_140_367#_c_655_n 0.0112861f $X=1.485 $Y=2.465 $X2=0
+ $Y2=0
cc_176 N_A1_c_122_n N_A_140_367#_c_655_n 0.0039872f $X=1.115 $Y=1.487 $X2=0
+ $Y2=0
cc_177 N_A1_c_145_p N_A_140_367#_c_655_n 0.0265866f $X=1.337 $Y=1.925 $X2=0
+ $Y2=0
cc_178 N_A1_c_127_n N_A_140_367#_c_655_n 2.70813e-19 $X=1.485 $Y=1.46 $X2=0
+ $Y2=0
cc_179 N_A1_c_136_p N_A_140_367#_c_660_n 0.0136314f $X=3.5 $Y=2.022 $X2=0 $Y2=0
cc_180 N_A1_c_136_p N_Y_M1011_s 0.00334566f $X=3.5 $Y=2.022 $X2=0 $Y2=0
cc_181 N_A1_c_136_p N_Y_M1021_s 0.00334999f $X=3.5 $Y=2.022 $X2=0 $Y2=0
cc_182 N_A1_M1031_g N_Y_c_694_n 0.0140867f $X=3.635 $Y=2.465 $X2=0 $Y2=0
cc_183 N_A1_c_159_p N_Y_c_694_n 0.0127022f $X=3.64 $Y=1.925 $X2=0 $Y2=0
cc_184 N_A1_c_125_n N_Y_c_694_n 0.00115422f $X=3.655 $Y=1.51 $X2=0 $Y2=0
cc_185 N_A1_c_136_p N_Y_c_694_n 0.0683359f $X=3.5 $Y=2.022 $X2=0 $Y2=0
cc_186 N_A1_c_136_p N_Y_c_698_n 0.0129035f $X=3.5 $Y=2.022 $X2=0 $Y2=0
cc_187 N_A1_M1010_g N_A_57_47#_c_790_n 0.0144681f $X=0.625 $Y=0.655 $X2=0 $Y2=0
cc_188 N_A1_M1020_g N_A_57_47#_c_790_n 0.0137055f $X=1.055 $Y=0.655 $X2=0 $Y2=0
cc_189 N_A1_c_122_n N_A_57_47#_c_790_n 0.0443533f $X=1.115 $Y=1.487 $X2=0 $Y2=0
cc_190 N_A1_c_123_n N_A_57_47#_c_790_n 0.0047208f $X=1.337 $Y=1.63 $X2=0 $Y2=0
cc_191 N_A1_c_126_n N_A_57_47#_c_790_n 0.00104779f $X=0.55 $Y=1.46 $X2=0 $Y2=0
cc_192 N_A1_c_127_n N_A_57_47#_c_790_n 0.00238134f $X=1.485 $Y=1.46 $X2=0 $Y2=0
cc_193 N_A1_c_122_n N_A_57_47#_c_791_n 0.016698f $X=1.115 $Y=1.487 $X2=0 $Y2=0
cc_194 N_A1_c_126_n N_A_57_47#_c_791_n 0.00494971f $X=0.55 $Y=1.46 $X2=0 $Y2=0
cc_195 N_A1_M1027_g N_A_57_47#_c_792_n 0.0137195f $X=1.485 $Y=0.655 $X2=0 $Y2=0
cc_196 N_A1_c_123_n N_A_57_47#_c_792_n 0.0150451f $X=1.337 $Y=1.63 $X2=0 $Y2=0
cc_197 N_A1_M1028_g N_A_57_47#_c_794_n 0.0141429f $X=3.645 $Y=0.655 $X2=0 $Y2=0
cc_198 N_A1_c_124_n N_A_57_47#_c_794_n 0.0197789f $X=3.655 $Y=1.51 $X2=0 $Y2=0
cc_199 N_A1_c_125_n N_A_57_47#_c_794_n 0.00114877f $X=3.655 $Y=1.51 $X2=0 $Y2=0
cc_200 N_A1_c_123_n N_A_57_47#_c_796_n 0.0169405f $X=1.337 $Y=1.63 $X2=0 $Y2=0
cc_201 N_A1_c_127_n N_A_57_47#_c_796_n 0.00247302f $X=1.485 $Y=1.46 $X2=0 $Y2=0
cc_202 N_A1_c_124_n N_A_57_47#_c_799_n 0.00213971f $X=3.655 $Y=1.51 $X2=0 $Y2=0
cc_203 N_A1_c_125_n N_A_57_47#_c_799_n 0.00201205f $X=3.655 $Y=1.51 $X2=0 $Y2=0
cc_204 N_A1_M1010_g N_VGND_c_895_n 0.0118316f $X=0.625 $Y=0.655 $X2=0 $Y2=0
cc_205 N_A1_M1020_g N_VGND_c_895_n 0.010076f $X=1.055 $Y=0.655 $X2=0 $Y2=0
cc_206 N_A1_M1027_g N_VGND_c_895_n 6.11179e-19 $X=1.485 $Y=0.655 $X2=0 $Y2=0
cc_207 N_A1_M1020_g N_VGND_c_896_n 6.05521e-19 $X=1.055 $Y=0.655 $X2=0 $Y2=0
cc_208 N_A1_M1027_g N_VGND_c_896_n 0.00985804f $X=1.485 $Y=0.655 $X2=0 $Y2=0
cc_209 N_A1_M1028_g N_VGND_c_898_n 0.0104772f $X=3.645 $Y=0.655 $X2=0 $Y2=0
cc_210 N_A1_M1020_g N_VGND_c_901_n 0.00486043f $X=1.055 $Y=0.655 $X2=0 $Y2=0
cc_211 N_A1_M1027_g N_VGND_c_901_n 0.00486043f $X=1.485 $Y=0.655 $X2=0 $Y2=0
cc_212 N_A1_M1028_g N_VGND_c_903_n 0.00525069f $X=3.645 $Y=0.655 $X2=0 $Y2=0
cc_213 N_A1_M1010_g N_VGND_c_904_n 0.00929414f $X=0.625 $Y=0.655 $X2=0 $Y2=0
cc_214 N_A1_M1020_g N_VGND_c_904_n 0.00824727f $X=1.055 $Y=0.655 $X2=0 $Y2=0
cc_215 N_A1_M1027_g N_VGND_c_904_n 0.00824727f $X=1.485 $Y=0.655 $X2=0 $Y2=0
cc_216 N_A1_M1028_g N_VGND_c_904_n 0.00896134f $X=3.645 $Y=0.655 $X2=0 $Y2=0
cc_217 N_A1_M1010_g N_VGND_c_905_n 0.00486043f $X=0.625 $Y=0.655 $X2=0 $Y2=0
cc_218 N_A2_c_243_n N_VPWR_c_523_n 0.00109252f $X=1.915 $Y=1.725 $X2=0 $Y2=0
cc_219 N_A2_c_246_n N_VPWR_c_524_n 0.0011792f $X=3.205 $Y=1.725 $X2=0 $Y2=0
cc_220 N_A2_c_243_n N_VPWR_c_529_n 0.00357877f $X=1.915 $Y=1.725 $X2=0 $Y2=0
cc_221 N_A2_c_244_n N_VPWR_c_529_n 0.00357877f $X=2.345 $Y=1.725 $X2=0 $Y2=0
cc_222 N_A2_c_245_n N_VPWR_c_529_n 0.00357877f $X=2.775 $Y=1.725 $X2=0 $Y2=0
cc_223 N_A2_c_246_n N_VPWR_c_529_n 0.00357877f $X=3.205 $Y=1.725 $X2=0 $Y2=0
cc_224 N_A2_c_243_n N_VPWR_c_520_n 0.00537654f $X=1.915 $Y=1.725 $X2=0 $Y2=0
cc_225 N_A2_c_244_n N_VPWR_c_520_n 0.0053512f $X=2.345 $Y=1.725 $X2=0 $Y2=0
cc_226 N_A2_c_245_n N_VPWR_c_520_n 0.0053512f $X=2.775 $Y=1.725 $X2=0 $Y2=0
cc_227 N_A2_c_246_n N_VPWR_c_520_n 0.00544922f $X=3.205 $Y=1.725 $X2=0 $Y2=0
cc_228 N_A2_c_243_n N_A_140_367#_c_661_n 0.0150519f $X=1.915 $Y=1.725 $X2=0
+ $Y2=0
cc_229 N_A2_c_244_n N_A_140_367#_c_661_n 0.0108707f $X=2.345 $Y=1.725 $X2=0
+ $Y2=0
cc_230 N_A2_c_245_n N_A_140_367#_c_661_n 0.0108707f $X=2.775 $Y=1.725 $X2=0
+ $Y2=0
cc_231 N_A2_c_246_n N_A_140_367#_c_661_n 0.011277f $X=3.205 $Y=1.725 $X2=0 $Y2=0
cc_232 N_A2_c_244_n N_Y_c_694_n 0.0105121f $X=2.345 $Y=1.725 $X2=0 $Y2=0
cc_233 N_A2_c_245_n N_Y_c_694_n 0.0104517f $X=2.775 $Y=1.725 $X2=0 $Y2=0
cc_234 N_A2_c_246_n N_Y_c_694_n 0.0104517f $X=3.205 $Y=1.725 $X2=0 $Y2=0
cc_235 N_A2_M1006_g N_A_57_47#_c_792_n 0.0146113f $X=1.915 $Y=0.655 $X2=0 $Y2=0
cc_236 A2 N_A_57_47#_c_792_n 0.00962057f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_237 N_A2_M1008_g N_A_57_47#_c_793_n 0.0142261f $X=2.345 $Y=0.655 $X2=0 $Y2=0
cc_238 N_A2_M1017_g N_A_57_47#_c_793_n 0.0142261f $X=2.775 $Y=0.655 $X2=0 $Y2=0
cc_239 A2 N_A_57_47#_c_793_n 0.0366479f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_240 N_A2_c_242_n N_A_57_47#_c_793_n 0.00240471f $X=3.205 $Y=1.535 $X2=0 $Y2=0
cc_241 N_A2_M1023_g N_A_57_47#_c_794_n 0.0142387f $X=3.205 $Y=0.655 $X2=0 $Y2=0
cc_242 A2 N_A_57_47#_c_794_n 0.0134492f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_243 A2 N_A_57_47#_c_797_n 0.0120054f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_244 N_A2_c_242_n N_A_57_47#_c_797_n 0.00252486f $X=3.205 $Y=1.535 $X2=0 $Y2=0
cc_245 A2 N_A_57_47#_c_798_n 0.0120054f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_246 N_A2_c_242_n N_A_57_47#_c_798_n 0.00252486f $X=3.205 $Y=1.535 $X2=0 $Y2=0
cc_247 N_A2_M1006_g N_VGND_c_896_n 0.00985804f $X=1.915 $Y=0.655 $X2=0 $Y2=0
cc_248 N_A2_M1008_g N_VGND_c_896_n 6.05521e-19 $X=2.345 $Y=0.655 $X2=0 $Y2=0
cc_249 N_A2_M1006_g N_VGND_c_897_n 6.11179e-19 $X=1.915 $Y=0.655 $X2=0 $Y2=0
cc_250 N_A2_M1008_g N_VGND_c_897_n 0.010076f $X=2.345 $Y=0.655 $X2=0 $Y2=0
cc_251 N_A2_M1017_g N_VGND_c_897_n 0.010076f $X=2.775 $Y=0.655 $X2=0 $Y2=0
cc_252 N_A2_M1023_g N_VGND_c_897_n 6.11179e-19 $X=3.205 $Y=0.655 $X2=0 $Y2=0
cc_253 N_A2_M1017_g N_VGND_c_898_n 6.11179e-19 $X=2.775 $Y=0.655 $X2=0 $Y2=0
cc_254 N_A2_M1023_g N_VGND_c_898_n 0.0100851f $X=3.205 $Y=0.655 $X2=0 $Y2=0
cc_255 N_A2_M1017_g N_VGND_c_899_n 0.00486043f $X=2.775 $Y=0.655 $X2=0 $Y2=0
cc_256 N_A2_M1023_g N_VGND_c_899_n 0.00486043f $X=3.205 $Y=0.655 $X2=0 $Y2=0
cc_257 N_A2_M1006_g N_VGND_c_902_n 0.00486043f $X=1.915 $Y=0.655 $X2=0 $Y2=0
cc_258 N_A2_M1008_g N_VGND_c_902_n 0.00486043f $X=2.345 $Y=0.655 $X2=0 $Y2=0
cc_259 N_A2_M1006_g N_VGND_c_904_n 0.00824727f $X=1.915 $Y=0.655 $X2=0 $Y2=0
cc_260 N_A2_M1008_g N_VGND_c_904_n 0.00824727f $X=2.345 $Y=0.655 $X2=0 $Y2=0
cc_261 N_A2_M1017_g N_VGND_c_904_n 0.00824727f $X=2.775 $Y=0.655 $X2=0 $Y2=0
cc_262 N_A2_M1023_g N_VGND_c_904_n 0.00824727f $X=3.205 $Y=0.655 $X2=0 $Y2=0
cc_263 N_B1_M1026_g N_C1_M1009_g 0.024313f $X=4.965 $Y=2.465 $X2=0 $Y2=0
cc_264 N_B1_c_330_n N_C1_M1009_g 0.00337642f $X=5.04 $Y=1.93 $X2=0 $Y2=0
cc_265 N_B1_c_346_p N_C1_M1009_g 0.0114498f $X=7.39 $Y=2.015 $X2=0 $Y2=0
cc_266 N_B1_M1014_g N_C1_M1003_g 0.0260155f $X=4.965 $Y=0.655 $X2=0 $Y2=0
cc_267 N_B1_c_346_p N_C1_M1012_g 0.0104926f $X=7.39 $Y=2.015 $X2=0 $Y2=0
cc_268 N_B1_c_346_p N_C1_M1019_g 0.0118664f $X=7.39 $Y=2.015 $X2=0 $Y2=0
cc_269 N_B1_M1030_g N_C1_M1029_g 0.0205623f $X=7.455 $Y=2.465 $X2=0 $Y2=0
cc_270 N_B1_c_346_p N_C1_M1029_g 0.0126613f $X=7.39 $Y=2.015 $X2=0 $Y2=0
cc_271 N_B1_M1015_g N_C1_M1024_g 0.0301291f $X=7.665 $Y=0.765 $X2=0 $Y2=0
cc_272 N_B1_c_321_n C1 0.0236004f $X=5.04 $Y=1.76 $X2=0 $Y2=0
cc_273 N_B1_c_346_p C1 0.116139f $X=7.39 $Y=2.015 $X2=0 $Y2=0
cc_274 N_B1_c_331_n C1 0.0149888f $X=7.555 $Y=1.51 $X2=0 $Y2=0
cc_275 N_B1_c_322_n C1 0.00113056f $X=7.555 $Y=1.51 $X2=0 $Y2=0
cc_276 N_B1_c_324_n C1 3.46547e-19 $X=4.965 $Y=1.51 $X2=0 $Y2=0
cc_277 N_B1_c_321_n N_C1_c_447_n 0.00497369f $X=5.04 $Y=1.76 $X2=0 $Y2=0
cc_278 N_B1_c_346_p N_C1_c_447_n 0.00357502f $X=7.39 $Y=2.015 $X2=0 $Y2=0
cc_279 N_B1_c_331_n N_C1_c_447_n 0.00247078f $X=7.555 $Y=1.51 $X2=0 $Y2=0
cc_280 N_B1_c_322_n N_C1_c_447_n 0.0314662f $X=7.555 $Y=1.51 $X2=0 $Y2=0
cc_281 N_B1_c_324_n N_C1_c_447_n 0.024313f $X=4.965 $Y=1.51 $X2=0 $Y2=0
cc_282 N_B1_c_346_p N_VPWR_M1009_s 0.00333608f $X=7.39 $Y=2.015 $X2=0 $Y2=0
cc_283 N_B1_c_346_p N_VPWR_M1019_s 0.012314f $X=7.39 $Y=2.015 $X2=0 $Y2=0
cc_284 N_B1_c_346_p N_VPWR_M1030_s 0.00344399f $X=7.39 $Y=2.015 $X2=0 $Y2=0
cc_285 N_B1_c_331_n N_VPWR_M1030_s 0.0010592f $X=7.555 $Y=1.51 $X2=0 $Y2=0
cc_286 N_B1_M1000_g N_VPWR_c_524_n 0.00822115f $X=4.105 $Y=2.465 $X2=0 $Y2=0
cc_287 N_B1_M1007_g N_VPWR_c_524_n 5.41941e-19 $X=4.535 $Y=2.465 $X2=0 $Y2=0
cc_288 N_B1_M1000_g N_VPWR_c_525_n 5.89638e-19 $X=4.105 $Y=2.465 $X2=0 $Y2=0
cc_289 N_B1_M1007_g N_VPWR_c_525_n 0.0109392f $X=4.535 $Y=2.465 $X2=0 $Y2=0
cc_290 N_B1_M1026_g N_VPWR_c_525_n 0.0109734f $X=4.965 $Y=2.465 $X2=0 $Y2=0
cc_291 N_B1_M1026_g N_VPWR_c_526_n 0.00486043f $X=4.965 $Y=2.465 $X2=0 $Y2=0
cc_292 N_B1_M1030_g N_VPWR_c_528_n 0.010963f $X=7.455 $Y=2.465 $X2=0 $Y2=0
cc_293 N_B1_M1000_g N_VPWR_c_531_n 0.00564095f $X=4.105 $Y=2.465 $X2=0 $Y2=0
cc_294 N_B1_M1007_g N_VPWR_c_531_n 0.00486043f $X=4.535 $Y=2.465 $X2=0 $Y2=0
cc_295 N_B1_M1030_g N_VPWR_c_533_n 0.00486043f $X=7.455 $Y=2.465 $X2=0 $Y2=0
cc_296 N_B1_M1000_g N_VPWR_c_520_n 0.00513564f $X=4.105 $Y=2.465 $X2=0 $Y2=0
cc_297 N_B1_M1007_g N_VPWR_c_520_n 0.00824727f $X=4.535 $Y=2.465 $X2=0 $Y2=0
cc_298 N_B1_M1026_g N_VPWR_c_520_n 0.0082726f $X=4.965 $Y=2.465 $X2=0 $Y2=0
cc_299 N_B1_M1030_g N_VPWR_c_520_n 0.00453535f $X=7.455 $Y=2.465 $X2=0 $Y2=0
cc_300 N_B1_M1030_g N_VPWR_c_541_n 5.78042e-19 $X=7.455 $Y=2.465 $X2=0 $Y2=0
cc_301 N_B1_c_330_n N_Y_M1026_d 0.00110935f $X=5.04 $Y=1.93 $X2=0 $Y2=0
cc_302 N_B1_c_346_p N_Y_M1026_d 0.00668365f $X=7.39 $Y=2.015 $X2=0 $Y2=0
cc_303 N_B1_c_384_p N_Y_M1026_d 2.98789e-19 $X=5.125 $Y=2.015 $X2=0 $Y2=0
cc_304 N_B1_c_346_p N_Y_M1012_d 0.00333177f $X=7.39 $Y=2.015 $X2=0 $Y2=0
cc_305 N_B1_c_346_p N_Y_M1029_d 0.00528167f $X=7.39 $Y=2.015 $X2=0 $Y2=0
cc_306 N_B1_M1000_g N_Y_c_694_n 0.0135363f $X=4.105 $Y=2.465 $X2=0 $Y2=0
cc_307 B1 N_Y_c_694_n 0.00681482f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_308 B1 N_Y_c_709_n 0.0164531f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_309 N_B1_c_324_n N_Y_c_709_n 6.37898e-19 $X=4.965 $Y=1.51 $X2=0 $Y2=0
cc_310 N_B1_M1007_g N_Y_c_711_n 0.0141904f $X=4.535 $Y=2.465 $X2=0 $Y2=0
cc_311 N_B1_M1026_g N_Y_c_711_n 0.0129881f $X=4.965 $Y=2.465 $X2=0 $Y2=0
cc_312 N_B1_c_384_p N_Y_c_711_n 0.00644085f $X=5.125 $Y=2.015 $X2=0 $Y2=0
cc_313 B1 N_Y_c_711_n 0.0153666f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_314 N_B1_c_324_n N_Y_c_711_n 4.70485e-19 $X=4.965 $Y=1.51 $X2=0 $Y2=0
cc_315 N_B1_c_346_p N_Y_c_716_n 0.0323235f $X=7.39 $Y=2.015 $X2=0 $Y2=0
cc_316 N_B1_M1014_g N_Y_c_686_n 0.00124217f $X=4.965 $Y=0.655 $X2=0 $Y2=0
cc_317 N_B1_M1015_g N_Y_c_687_n 0.0142815f $X=7.665 $Y=0.765 $X2=0 $Y2=0
cc_318 N_B1_c_346_p N_Y_c_687_n 0.00742542f $X=7.39 $Y=2.015 $X2=0 $Y2=0
cc_319 N_B1_c_331_n N_Y_c_687_n 0.0258173f $X=7.555 $Y=1.51 $X2=0 $Y2=0
cc_320 N_B1_c_322_n N_Y_c_687_n 0.00582955f $X=7.555 $Y=1.51 $X2=0 $Y2=0
cc_321 N_B1_M1030_g N_Y_c_688_n 0.00672688f $X=7.455 $Y=2.465 $X2=0 $Y2=0
cc_322 N_B1_M1015_g N_Y_c_688_n 0.0120828f $X=7.665 $Y=0.765 $X2=0 $Y2=0
cc_323 N_B1_c_346_p N_Y_c_688_n 0.0141128f $X=7.39 $Y=2.015 $X2=0 $Y2=0
cc_324 N_B1_c_331_n N_Y_c_688_n 0.0389862f $X=7.555 $Y=1.51 $X2=0 $Y2=0
cc_325 N_B1_c_346_p N_Y_c_726_n 0.011191f $X=7.39 $Y=2.015 $X2=0 $Y2=0
cc_326 N_B1_c_384_p N_Y_c_726_n 0.00247945f $X=5.125 $Y=2.015 $X2=0 $Y2=0
cc_327 N_B1_M1015_g N_Y_c_689_n 4.88604e-19 $X=7.665 $Y=0.765 $X2=0 $Y2=0
cc_328 N_B1_c_346_p N_Y_c_729_n 0.0584476f $X=7.39 $Y=2.015 $X2=0 $Y2=0
cc_329 N_B1_c_346_p N_Y_c_730_n 0.0135055f $X=7.39 $Y=2.015 $X2=0 $Y2=0
cc_330 N_B1_M1030_g N_Y_c_691_n 0.0140565f $X=7.455 $Y=2.465 $X2=0 $Y2=0
cc_331 N_B1_c_346_p N_Y_c_691_n 0.0224952f $X=7.39 $Y=2.015 $X2=0 $Y2=0
cc_332 N_B1_c_322_n N_Y_c_691_n 0.00107403f $X=7.555 $Y=1.51 $X2=0 $Y2=0
cc_333 N_B1_c_346_p Y 0.0135055f $X=7.39 $Y=2.015 $X2=0 $Y2=0
cc_334 N_B1_M1001_g N_A_57_47#_c_795_n 0.013828f $X=4.105 $Y=0.655 $X2=0 $Y2=0
cc_335 N_B1_M1002_g N_A_57_47#_c_795_n 0.0123883f $X=4.535 $Y=0.655 $X2=0 $Y2=0
cc_336 N_B1_M1014_g N_A_57_47#_c_795_n 0.00676029f $X=4.965 $Y=0.655 $X2=0 $Y2=0
cc_337 B1 N_A_57_47#_c_795_n 0.0722485f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_338 N_B1_c_324_n N_A_57_47#_c_795_n 0.00455638f $X=4.965 $Y=1.51 $X2=0 $Y2=0
cc_339 N_B1_M1014_g N_A_57_47#_c_835_n 7.24563e-19 $X=4.965 $Y=0.655 $X2=0 $Y2=0
cc_340 N_B1_M1014_g N_A_57_47#_c_836_n 0.00427771f $X=4.965 $Y=0.655 $X2=0 $Y2=0
cc_341 N_B1_M1014_g N_A_57_47#_c_837_n 0.00985252f $X=4.965 $Y=0.655 $X2=0 $Y2=0
cc_342 N_B1_M1015_g N_A_57_47#_c_837_n 0.010167f $X=7.665 $Y=0.765 $X2=0 $Y2=0
cc_343 N_B1_c_321_n N_A_57_47#_c_837_n 0.00463886f $X=5.04 $Y=1.76 $X2=0 $Y2=0
cc_344 B1 N_A_57_47#_c_837_n 0.00108207f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_345 B1 N_A_57_47#_c_799_n 0.00314774f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_346 N_B1_M1015_g N_A_57_47#_c_800_n 0.00825439f $X=7.665 $Y=0.765 $X2=0 $Y2=0
cc_347 N_B1_M1001_g N_VGND_c_898_n 0.00117355f $X=4.105 $Y=0.655 $X2=0 $Y2=0
cc_348 N_B1_M1001_g N_VGND_c_903_n 0.0054778f $X=4.105 $Y=0.655 $X2=0 $Y2=0
cc_349 N_B1_M1002_g N_VGND_c_903_n 0.0035993f $X=4.535 $Y=0.655 $X2=0 $Y2=0
cc_350 N_B1_M1014_g N_VGND_c_903_n 0.00359964f $X=4.965 $Y=0.655 $X2=0 $Y2=0
cc_351 N_B1_M1015_g N_VGND_c_903_n 0.00336885f $X=7.665 $Y=0.765 $X2=0 $Y2=0
cc_352 N_B1_M1001_g N_VGND_c_904_n 0.00997231f $X=4.105 $Y=0.655 $X2=0 $Y2=0
cc_353 N_B1_M1002_g N_VGND_c_904_n 0.00535284f $X=4.535 $Y=0.655 $X2=0 $Y2=0
cc_354 N_B1_M1014_g N_VGND_c_904_n 0.00663456f $X=4.965 $Y=0.655 $X2=0 $Y2=0
cc_355 N_B1_M1015_g N_VGND_c_904_n 0.0047742f $X=7.665 $Y=0.765 $X2=0 $Y2=0
cc_356 N_B1_M1002_g N_A_836_47#_c_991_n 0.00878231f $X=4.535 $Y=0.655 $X2=0
+ $Y2=0
cc_357 N_B1_M1014_g N_A_836_47#_c_991_n 0.0116629f $X=4.965 $Y=0.655 $X2=0 $Y2=0
cc_358 N_B1_M1015_g N_A_836_47#_c_991_n 0.0033042f $X=7.665 $Y=0.765 $X2=0 $Y2=0
cc_359 N_B1_M1001_g N_A_836_47#_c_995_n 0.00622367f $X=4.105 $Y=0.655 $X2=0
+ $Y2=0
cc_360 N_B1_M1002_g N_A_836_47#_c_995_n 0.00605622f $X=4.535 $Y=0.655 $X2=0
+ $Y2=0
cc_361 N_B1_M1014_g N_A_836_47#_c_995_n 7.61432e-19 $X=4.965 $Y=0.655 $X2=0
+ $Y2=0
cc_362 N_C1_M1009_g N_VPWR_c_525_n 5.95693e-19 $X=5.395 $Y=2.465 $X2=0 $Y2=0
cc_363 N_C1_M1009_g N_VPWR_c_526_n 0.00585385f $X=5.395 $Y=2.465 $X2=0 $Y2=0
cc_364 N_C1_M1009_g N_VPWR_c_527_n 0.00215341f $X=5.395 $Y=2.465 $X2=0 $Y2=0
cc_365 N_C1_M1012_g N_VPWR_c_527_n 0.00211296f $X=5.825 $Y=2.465 $X2=0 $Y2=0
cc_366 N_C1_M1029_g N_VPWR_c_528_n 5.63085e-19 $X=7.025 $Y=2.465 $X2=0 $Y2=0
cc_367 N_C1_M1029_g N_VPWR_c_533_n 0.00487821f $X=7.025 $Y=2.465 $X2=0 $Y2=0
cc_368 N_C1_M1012_g N_VPWR_c_536_n 0.00585385f $X=5.825 $Y=2.465 $X2=0 $Y2=0
cc_369 N_C1_M1019_g N_VPWR_c_536_n 0.00487821f $X=6.255 $Y=2.465 $X2=0 $Y2=0
cc_370 N_C1_M1009_g N_VPWR_c_520_n 0.0106551f $X=5.395 $Y=2.465 $X2=0 $Y2=0
cc_371 N_C1_M1012_g N_VPWR_c_520_n 0.0106571f $X=5.825 $Y=2.465 $X2=0 $Y2=0
cc_372 N_C1_M1019_g N_VPWR_c_520_n 0.00451006f $X=6.255 $Y=2.465 $X2=0 $Y2=0
cc_373 N_C1_M1029_g N_VPWR_c_520_n 0.0045354f $X=7.025 $Y=2.465 $X2=0 $Y2=0
cc_374 N_C1_M1012_g N_VPWR_c_541_n 5.97452e-19 $X=5.825 $Y=2.465 $X2=0 $Y2=0
cc_375 N_C1_M1019_g N_VPWR_c_541_n 0.0114568f $X=6.255 $Y=2.465 $X2=0 $Y2=0
cc_376 N_C1_M1029_g N_VPWR_c_541_n 0.0113537f $X=7.025 $Y=2.465 $X2=0 $Y2=0
cc_377 N_C1_M1009_g N_Y_c_716_n 0.0129934f $X=5.395 $Y=2.465 $X2=0 $Y2=0
cc_378 N_C1_M1012_g N_Y_c_716_n 0.0129934f $X=5.825 $Y=2.465 $X2=0 $Y2=0
cc_379 N_C1_M1003_g N_Y_c_686_n 0.00828011f $X=5.625 $Y=0.765 $X2=0 $Y2=0
cc_380 N_C1_M1016_g N_Y_c_686_n 0.0138625f $X=6.055 $Y=0.765 $X2=0 $Y2=0
cc_381 N_C1_M1022_g N_Y_c_686_n 0.0138625f $X=6.645 $Y=0.765 $X2=0 $Y2=0
cc_382 C1 N_Y_c_686_n 0.105825f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_383 N_C1_c_447_n N_Y_c_686_n 0.0129945f $X=7.025 $Y=1.51 $X2=0 $Y2=0
cc_384 N_C1_M1024_g N_Y_c_687_n 0.0101933f $X=7.075 $Y=0.765 $X2=0 $Y2=0
cc_385 N_C1_M1024_g N_Y_c_689_n 0.00434837f $X=7.075 $Y=0.765 $X2=0 $Y2=0
cc_386 N_C1_M1019_g N_Y_c_729_n 0.0134403f $X=6.255 $Y=2.465 $X2=0 $Y2=0
cc_387 N_C1_M1029_g N_Y_c_729_n 0.0134403f $X=7.025 $Y=2.465 $X2=0 $Y2=0
cc_388 N_C1_M1003_g N_A_57_47#_c_795_n 7.76353e-19 $X=5.625 $Y=0.765 $X2=0 $Y2=0
cc_389 N_C1_M1003_g N_A_57_47#_c_836_n 8.66905e-19 $X=5.625 $Y=0.765 $X2=0 $Y2=0
cc_390 N_C1_M1003_g N_A_57_47#_c_837_n 0.0132324f $X=5.625 $Y=0.765 $X2=0 $Y2=0
cc_391 N_C1_M1016_g N_A_57_47#_c_837_n 0.0112681f $X=6.055 $Y=0.765 $X2=0 $Y2=0
cc_392 N_C1_M1022_g N_A_57_47#_c_837_n 0.0112681f $X=6.645 $Y=0.765 $X2=0 $Y2=0
cc_393 N_C1_M1024_g N_A_57_47#_c_837_n 0.011723f $X=7.075 $Y=0.765 $X2=0 $Y2=0
cc_394 C1 N_A_57_47#_c_837_n 0.00735546f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_395 N_C1_c_447_n N_A_57_47#_c_837_n 0.00463668f $X=7.025 $Y=1.51 $X2=0 $Y2=0
cc_396 N_C1_M1024_g N_A_57_47#_c_800_n 0.00141389f $X=7.075 $Y=0.765 $X2=0 $Y2=0
cc_397 N_C1_M1003_g N_VGND_c_903_n 0.00293025f $X=5.625 $Y=0.765 $X2=0 $Y2=0
cc_398 N_C1_M1016_g N_VGND_c_903_n 0.00293025f $X=6.055 $Y=0.765 $X2=0 $Y2=0
cc_399 N_C1_M1022_g N_VGND_c_903_n 0.00293025f $X=6.645 $Y=0.765 $X2=0 $Y2=0
cc_400 N_C1_M1024_g N_VGND_c_903_n 0.00293025f $X=7.075 $Y=0.765 $X2=0 $Y2=0
cc_401 N_C1_M1003_g N_VGND_c_904_n 0.00409921f $X=5.625 $Y=0.765 $X2=0 $Y2=0
cc_402 N_C1_M1016_g N_VGND_c_904_n 0.00407106f $X=6.055 $Y=0.765 $X2=0 $Y2=0
cc_403 N_C1_M1022_g N_VGND_c_904_n 0.00407106f $X=6.645 $Y=0.765 $X2=0 $Y2=0
cc_404 N_C1_M1024_g N_VGND_c_904_n 0.00407167f $X=7.075 $Y=0.765 $X2=0 $Y2=0
cc_405 N_C1_M1003_g N_A_836_47#_c_991_n 0.0112452f $X=5.625 $Y=0.765 $X2=0 $Y2=0
cc_406 N_C1_M1016_g N_A_836_47#_c_991_n 0.0110477f $X=6.055 $Y=0.765 $X2=0 $Y2=0
cc_407 N_C1_M1022_g N_A_836_47#_c_991_n 0.0110477f $X=6.645 $Y=0.765 $X2=0 $Y2=0
cc_408 N_C1_M1024_g N_A_836_47#_c_991_n 0.0106892f $X=7.075 $Y=0.765 $X2=0 $Y2=0
cc_409 N_VPWR_c_520_n N_A_140_367#_M1004_d 0.00273541f $X=7.92 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_410 N_VPWR_c_520_n N_A_140_367#_M1013_d 0.00250769f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_411 N_VPWR_c_520_n N_A_140_367#_M1018_d 0.00223577f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_412 N_VPWR_c_520_n N_A_140_367#_M1025_d 0.00247351f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_413 N_VPWR_c_522_n N_A_140_367#_c_645_n 0.00151856f $X=0.41 $Y=1.98 $X2=0
+ $Y2=0
cc_414 N_VPWR_M1005_s N_A_140_367#_c_655_n 0.00345715f $X=1.13 $Y=1.835 $X2=0
+ $Y2=0
cc_415 N_VPWR_c_523_n N_A_140_367#_c_655_n 0.0169953f $X=1.27 $Y=2.815 $X2=0
+ $Y2=0
cc_416 N_VPWR_c_520_n N_A_140_367#_c_655_n 0.0119319f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_417 N_VPWR_c_529_n N_A_140_367#_c_673_n 0.0128782f $X=3.705 $Y=3.33 $X2=0
+ $Y2=0
cc_418 N_VPWR_c_520_n N_A_140_367#_c_673_n 0.00777554f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_419 N_VPWR_c_535_n N_A_140_367#_c_675_n 0.0135169f $X=1.105 $Y=3.33 $X2=0
+ $Y2=0
cc_420 N_VPWR_c_520_n N_A_140_367#_c_675_n 0.00847005f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_421 N_VPWR_c_529_n N_A_140_367#_c_661_n 0.0976286f $X=3.705 $Y=3.33 $X2=0
+ $Y2=0
cc_422 N_VPWR_c_520_n N_A_140_367#_c_661_n 0.0624058f $X=7.92 $Y=3.33 $X2=0
+ $Y2=0
cc_423 N_VPWR_c_520_n N_Y_M1011_s 0.00224381f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_424 N_VPWR_c_520_n N_Y_M1021_s 0.00225186f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_425 N_VPWR_c_520_n N_Y_M1000_d 0.00394499f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_426 N_VPWR_c_520_n N_Y_M1026_d 0.0041489f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_427 N_VPWR_c_520_n N_Y_M1012_d 0.00250952f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_428 N_VPWR_c_520_n N_Y_M1029_d 0.00278345f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_429 N_VPWR_M1031_s N_Y_c_694_n 0.00854213f $X=3.71 $Y=1.835 $X2=0 $Y2=0
cc_430 N_VPWR_c_524_n N_Y_c_694_n 0.0171653f $X=3.87 $Y=2.805 $X2=0 $Y2=0
cc_431 N_VPWR_c_520_n N_Y_c_694_n 0.0144204f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_432 N_VPWR_M1007_s N_Y_c_711_n 0.00456103f $X=4.61 $Y=1.835 $X2=0 $Y2=0
cc_433 N_VPWR_c_525_n N_Y_c_711_n 0.0170777f $X=4.75 $Y=2.745 $X2=0 $Y2=0
cc_434 N_VPWR_M1009_s N_Y_c_716_n 0.00344105f $X=5.47 $Y=1.835 $X2=0 $Y2=0
cc_435 N_VPWR_c_527_n N_Y_c_716_n 0.0135055f $X=5.61 $Y=2.775 $X2=0 $Y2=0
cc_436 N_VPWR_c_536_n N_Y_c_759_n 0.0140491f $X=6.305 $Y=3.33 $X2=0 $Y2=0
cc_437 N_VPWR_c_520_n N_Y_c_759_n 0.0090585f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_438 N_VPWR_c_533_n N_Y_c_761_n 0.0124525f $X=7.505 $Y=3.33 $X2=0 $Y2=0
cc_439 N_VPWR_c_520_n N_Y_c_761_n 0.00730901f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_440 N_VPWR_c_531_n N_Y_c_763_n 0.0131621f $X=4.585 $Y=3.33 $X2=0 $Y2=0
cc_441 N_VPWR_c_520_n N_Y_c_763_n 0.00808656f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_442 N_VPWR_c_526_n N_Y_c_726_n 0.0136943f $X=5.48 $Y=3.33 $X2=0 $Y2=0
cc_443 N_VPWR_c_520_n N_Y_c_726_n 0.00866972f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_444 N_VPWR_M1019_s N_Y_c_729_n 0.0137412f $X=6.33 $Y=1.835 $X2=0 $Y2=0
cc_445 N_VPWR_c_520_n N_Y_c_729_n 0.0125576f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_446 N_VPWR_c_541_n N_Y_c_729_n 0.0446491f $X=6.81 $Y=2.805 $X2=0 $Y2=0
cc_447 N_VPWR_M1030_s N_Y_c_691_n 0.00712074f $X=7.53 $Y=1.835 $X2=0 $Y2=0
cc_448 N_VPWR_c_528_n N_Y_c_691_n 0.0219591f $X=7.67 $Y=2.825 $X2=0 $Y2=0
cc_449 N_VPWR_c_520_n N_Y_c_691_n 0.0154106f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_450 N_A_140_367#_c_661_n N_Y_M1011_s 0.00341273f $X=3.315 $Y=2.877 $X2=0
+ $Y2=0
cc_451 N_A_140_367#_c_661_n N_Y_M1021_s 0.00391015f $X=3.315 $Y=2.877 $X2=0
+ $Y2=0
cc_452 N_A_140_367#_M1018_d N_Y_c_694_n 0.00394558f $X=2.42 $Y=1.835 $X2=0 $Y2=0
cc_453 N_A_140_367#_M1025_d N_Y_c_694_n 0.00347683f $X=3.28 $Y=1.835 $X2=0 $Y2=0
cc_454 N_A_140_367#_c_683_p N_Y_c_694_n 0.0126145f $X=3.42 $Y=2.845 $X2=0 $Y2=0
cc_455 N_A_140_367#_c_661_n N_Y_c_694_n 0.0335956f $X=3.315 $Y=2.877 $X2=0 $Y2=0
cc_456 N_A_140_367#_c_661_n N_Y_c_698_n 0.0120339f $X=3.315 $Y=2.877 $X2=0 $Y2=0
cc_457 N_Y_c_687_n N_A_57_47#_M1015_s 0.00311294f $X=7.89 $Y=1.165 $X2=0 $Y2=0
cc_458 N_Y_M1003_s N_A_57_47#_c_837_n 0.00336136f $X=5.7 $Y=0.345 $X2=0 $Y2=0
cc_459 N_Y_M1022_s N_A_57_47#_c_837_n 0.00336136f $X=6.72 $Y=0.345 $X2=0 $Y2=0
cc_460 N_Y_c_686_n N_A_57_47#_c_837_n 0.074332f $X=6.88 $Y=1.11 $X2=0 $Y2=0
cc_461 N_Y_c_687_n N_A_57_47#_c_837_n 0.0278733f $X=7.89 $Y=1.165 $X2=0 $Y2=0
cc_462 N_Y_c_687_n N_A_57_47#_c_800_n 0.0228956f $X=7.89 $Y=1.165 $X2=0 $Y2=0
cc_463 N_Y_c_686_n N_A_836_47#_M1016_d 0.00450125f $X=6.88 $Y=1.11 $X2=0 $Y2=0
cc_464 N_Y_c_687_n N_A_836_47#_M1024_d 0.00484944f $X=7.89 $Y=1.165 $X2=0 $Y2=0
cc_465 N_Y_M1003_s N_A_836_47#_c_991_n 0.001775f $X=5.7 $Y=0.345 $X2=0 $Y2=0
cc_466 N_Y_M1022_s N_A_836_47#_c_991_n 0.001775f $X=6.72 $Y=0.345 $X2=0 $Y2=0
cc_467 N_A_57_47#_c_790_n N_VGND_M1010_d 0.00176773f $X=1.175 $Y=1.085 $X2=-0.19
+ $Y2=-0.245
cc_468 N_A_57_47#_c_792_n N_VGND_M1027_d 0.00185322f $X=2.035 $Y=1.085 $X2=0
+ $Y2=0
cc_469 N_A_57_47#_c_793_n N_VGND_M1008_d 0.00176773f $X=2.895 $Y=1.085 $X2=0
+ $Y2=0
cc_470 N_A_57_47#_c_794_n N_VGND_M1023_d 0.00187422f $X=3.755 $Y=1.085 $X2=0
+ $Y2=0
cc_471 N_A_57_47#_c_790_n N_VGND_c_895_n 0.0171443f $X=1.175 $Y=1.085 $X2=0
+ $Y2=0
cc_472 N_A_57_47#_c_792_n N_VGND_c_896_n 0.0157565f $X=2.035 $Y=1.085 $X2=0
+ $Y2=0
cc_473 N_A_57_47#_c_793_n N_VGND_c_897_n 0.0171443f $X=2.895 $Y=1.085 $X2=0
+ $Y2=0
cc_474 N_A_57_47#_c_794_n N_VGND_c_898_n 0.0171962f $X=3.755 $Y=1.085 $X2=0
+ $Y2=0
cc_475 N_A_57_47#_c_866_p N_VGND_c_899_n 0.0124525f $X=2.99 $Y=0.42 $X2=0 $Y2=0
cc_476 N_A_57_47#_c_867_p N_VGND_c_901_n 0.0124525f $X=1.27 $Y=0.42 $X2=0 $Y2=0
cc_477 N_A_57_47#_c_868_p N_VGND_c_902_n 0.0124525f $X=2.13 $Y=0.42 $X2=0 $Y2=0
cc_478 N_A_57_47#_c_869_p N_VGND_c_903_n 0.0149167f $X=3.87 $Y=0.42 $X2=0 $Y2=0
cc_479 N_A_57_47#_c_837_n N_VGND_c_903_n 0.00264215f $X=7.715 $Y=0.71 $X2=0
+ $Y2=0
cc_480 N_A_57_47#_c_800_n N_VGND_c_903_n 0.0121119f $X=7.88 $Y=0.47 $X2=0 $Y2=0
cc_481 N_A_57_47#_M1010_s N_VGND_c_904_n 0.00444756f $X=0.285 $Y=0.235 $X2=0
+ $Y2=0
cc_482 N_A_57_47#_M1020_s N_VGND_c_904_n 0.00536646f $X=1.13 $Y=0.235 $X2=0
+ $Y2=0
cc_483 N_A_57_47#_M1006_s N_VGND_c_904_n 0.00536646f $X=1.99 $Y=0.235 $X2=0
+ $Y2=0
cc_484 N_A_57_47#_M1017_s N_VGND_c_904_n 0.00536646f $X=2.85 $Y=0.235 $X2=0
+ $Y2=0
cc_485 N_A_57_47#_M1028_s N_VGND_c_904_n 0.00525984f $X=3.72 $Y=0.235 $X2=0
+ $Y2=0
cc_486 N_A_57_47#_M1002_s N_VGND_c_904_n 0.00225465f $X=4.61 $Y=0.235 $X2=0
+ $Y2=0
cc_487 N_A_57_47#_c_878_p N_VGND_c_904_n 0.00769778f $X=0.41 $Y=0.42 $X2=0 $Y2=0
cc_488 N_A_57_47#_c_867_p N_VGND_c_904_n 0.00730901f $X=1.27 $Y=0.42 $X2=0 $Y2=0
cc_489 N_A_57_47#_c_868_p N_VGND_c_904_n 0.00730901f $X=2.13 $Y=0.42 $X2=0 $Y2=0
cc_490 N_A_57_47#_c_866_p N_VGND_c_904_n 0.00730901f $X=2.99 $Y=0.42 $X2=0 $Y2=0
cc_491 N_A_57_47#_c_869_p N_VGND_c_904_n 0.00886411f $X=3.87 $Y=0.42 $X2=0 $Y2=0
cc_492 N_A_57_47#_c_837_n N_VGND_c_904_n 0.00951814f $X=7.715 $Y=0.71 $X2=0
+ $Y2=0
cc_493 N_A_57_47#_c_800_n N_VGND_c_904_n 0.0117806f $X=7.88 $Y=0.47 $X2=0 $Y2=0
cc_494 N_A_57_47#_c_878_p N_VGND_c_905_n 0.0135387f $X=0.41 $Y=0.42 $X2=0 $Y2=0
cc_495 N_A_57_47#_c_795_n N_A_836_47#_M1001_d 0.00176773f $X=4.655 $Y=1.085
+ $X2=-0.19 $Y2=-0.245
cc_496 N_A_57_47#_c_837_n N_A_836_47#_M1014_d 0.0163535f $X=7.715 $Y=0.71 $X2=0
+ $Y2=0
cc_497 N_A_57_47#_c_837_n N_A_836_47#_M1016_d 0.00727881f $X=7.715 $Y=0.71 $X2=0
+ $Y2=0
cc_498 N_A_57_47#_c_837_n N_A_836_47#_M1024_d 0.00820897f $X=7.715 $Y=0.71 $X2=0
+ $Y2=0
cc_499 N_A_57_47#_M1002_s N_A_836_47#_c_991_n 0.00336963f $X=4.61 $Y=0.235 $X2=0
+ $Y2=0
cc_500 N_A_57_47#_c_795_n N_A_836_47#_c_991_n 0.00331416f $X=4.655 $Y=1.085
+ $X2=0 $Y2=0
cc_501 N_A_57_47#_c_835_n N_A_836_47#_c_991_n 0.0143514f $X=4.785 $Y=0.795 $X2=0
+ $Y2=0
cc_502 N_A_57_47#_c_837_n N_A_836_47#_c_991_n 0.142608f $X=7.715 $Y=0.71 $X2=0
+ $Y2=0
cc_503 N_A_57_47#_c_795_n N_A_836_47#_c_995_n 0.0168764f $X=4.655 $Y=1.085 $X2=0
+ $Y2=0
cc_504 N_VGND_c_904_n N_A_836_47#_M1001_d 0.00223819f $X=7.92 $Y=0 $X2=-0.19
+ $Y2=-0.245
cc_505 N_VGND_c_904_n N_A_836_47#_M1014_d 0.00327137f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_506 N_VGND_c_904_n N_A_836_47#_M1016_d 0.00236207f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_507 N_VGND_c_904_n N_A_836_47#_M1024_d 0.00236207f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_508 N_VGND_c_903_n N_A_836_47#_c_991_n 0.177893f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_509 N_VGND_c_904_n N_A_836_47#_c_991_n 0.110256f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_510 N_VGND_c_903_n N_A_836_47#_c_995_n 0.0177289f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_511 N_VGND_c_904_n N_A_836_47#_c_995_n 0.0123275f $X=7.92 $Y=0 $X2=0 $Y2=0
