# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__dfrbp_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_lp__dfrbp_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  12.00000 BY  3.330000 ;
  SYMMETRY R90 ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.060000 1.210000 2.640000 2.155000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.588000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.185000 0.335000 11.410000 3.075000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.588000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.195000 0.820000 9.455000 2.920000 ;
        RECT 9.265000 0.255000 9.455000 0.820000 ;
    END
  END Q_N
  PIN RESET_B
    ANTENNAGATEAREA  0.378000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1.535000 1.920000 1.825000 1.965000 ;
        RECT 1.535000 1.965000 8.065000 2.105000 ;
        RECT 1.535000 2.105000 1.825000 2.150000 ;
        RECT 4.415000 1.920000 4.705000 1.965000 ;
        RECT 4.415000 2.105000 4.705000 2.150000 ;
        RECT 7.775000 1.920000 8.065000 1.965000 ;
        RECT 7.775000 2.105000 8.065000 2.150000 ;
    END
  END RESET_B
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.525000 1.495000 0.905000 2.165000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 12.000000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 12.000000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 12.000000 0.085000 ;
      RECT  0.000000  3.245000 12.000000 3.415000 ;
      RECT  0.120000  0.425000  0.400000 0.925000 ;
      RECT  0.120000  0.925000  1.055000 1.255000 ;
      RECT  0.120000  1.255000  0.355000 2.335000 ;
      RECT  0.120000  2.335000  0.380000 3.020000 ;
      RECT  0.550000  2.335000  0.880000 3.245000 ;
      RECT  0.570000  0.085000  0.830000 0.755000 ;
      RECT  1.000000  0.395000  1.405000 0.755000 ;
      RECT  1.050000  2.335000  1.380000 3.020000 ;
      RECT  1.110000  2.305000  1.380000 2.335000 ;
      RECT  1.210000  1.935000  1.415000 2.155000 ;
      RECT  1.210000  2.155000  1.380000 2.305000 ;
      RECT  1.235000  0.755000  1.405000 0.870000 ;
      RECT  1.235000  0.870000  2.315000 1.040000 ;
      RECT  1.235000  1.040000  1.415000 1.935000 ;
      RECT  1.550000  2.325000  3.365000 2.495000 ;
      RECT  1.550000  2.495000  1.750000 2.735000 ;
      RECT  1.575000  0.085000  1.905000 0.700000 ;
      RECT  1.585000  1.450000  1.890000 2.155000 ;
      RECT  1.990000  2.665000  2.340000 3.245000 ;
      RECT  2.075000  0.630000  4.775000 0.720000 ;
      RECT  2.075000  0.720000  6.470000 0.800000 ;
      RECT  2.075000  0.800000  2.315000 0.870000 ;
      RECT  2.560000  2.495000  3.365000 2.735000 ;
      RECT  2.810000  0.980000  3.035000 2.115000 ;
      RECT  2.810000  2.115000  3.170000 2.300000 ;
      RECT  2.810000  2.300000  3.365000 2.325000 ;
      RECT  3.205000  0.800000  3.375000 1.615000 ;
      RECT  3.205000  1.615000  3.625000 1.945000 ;
      RECT  3.535000  2.370000  5.115000 2.470000 ;
      RECT  3.535000  2.470000  3.985000 2.735000 ;
      RECT  3.545000  0.970000  4.235000 1.060000 ;
      RECT  3.545000  1.060000  5.620000 1.260000 ;
      RECT  3.545000  1.260000  3.965000 1.300000 ;
      RECT  3.795000  1.300000  3.965000 2.300000 ;
      RECT  3.795000  2.300000  5.115000 2.370000 ;
      RECT  4.135000  1.440000  5.260000 1.610000 ;
      RECT  4.135000  1.610000  4.305000 2.030000 ;
      RECT  4.360000  2.650000  4.690000 3.245000 ;
      RECT  4.475000  1.950000  4.920000 2.120000 ;
      RECT  4.495000  1.790000  4.920000 1.950000 ;
      RECT  4.560000  0.800000  6.470000 0.890000 ;
      RECT  4.870000  2.470000  5.115000 2.735000 ;
      RECT  5.090000  1.610000  5.260000 1.900000 ;
      RECT  5.090000  1.900000  6.165000 2.070000 ;
      RECT  5.245000  0.085000  5.575000 0.550000 ;
      RECT  5.370000  2.240000  5.700000 3.245000 ;
      RECT  5.430000  1.260000  5.620000 1.720000 ;
      RECT  5.790000  1.060000  6.120000 1.320000 ;
      RECT  5.950000  1.320000  6.120000 1.900000 ;
      RECT  5.950000  2.070000  6.165000 2.910000 ;
      RECT  6.290000  0.890000  6.470000 1.720000 ;
      RECT  6.520000  2.040000  6.840000 2.915000 ;
      RECT  6.640000  0.630000  6.840000 1.240000 ;
      RECT  6.640000  1.240000  8.565000 1.430000 ;
      RECT  6.640000  1.430000  6.840000 2.040000 ;
      RECT  7.220000  1.600000  9.025000 1.770000 ;
      RECT  7.220000  1.770000  8.490000 1.780000 ;
      RECT  7.220000  1.780000  7.550000 2.270000 ;
      RECT  7.345000  2.525000  8.025000 3.245000 ;
      RECT  7.455000  0.085000  7.785000 1.015000 ;
      RECT  7.760000  1.950000  8.050000 2.280000 ;
      RECT  8.220000  1.780000  8.490000 2.855000 ;
      RECT  8.245000  0.820000  9.025000 1.070000 ;
      RECT  8.685000  1.940000  9.015000 3.245000 ;
      RECT  8.745000  1.070000  9.025000 1.600000 ;
      RECT  8.765000  0.085000  9.095000 0.650000 ;
      RECT  9.625000  0.085000  9.955000 1.110000 ;
      RECT  9.625000  1.620000  9.875000 3.245000 ;
      RECT 10.125000  0.385000 10.490000 1.295000 ;
      RECT 10.125000  1.295000 11.015000 1.625000 ;
      RECT 10.125000  1.625000 10.430000 2.485000 ;
      RECT 10.600000  1.815000 10.955000 3.245000 ;
      RECT 10.660000  0.085000 11.015000 1.125000 ;
      RECT 11.580000  0.085000 11.875000 1.205000 ;
      RECT 11.580000  1.815000 11.875000 3.245000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  1.950000  1.765000 2.120000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  1.950000  8.005000 2.120000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.245000 10.885000 3.415000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  3.245000 11.365000 3.415000 ;
      RECT 11.675000 -0.085000 11.845000 0.085000 ;
      RECT 11.675000  3.245000 11.845000 3.415000 ;
  END
END sky130_fd_sc_lp__dfrbp_2
END LIBRARY
