* File: sky130_fd_sc_lp__sdfrtp_2.spice
* Created: Wed Sep  2 10:34:43 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__sdfrtp_2.pex.spice"
.subckt sky130_fd_sc_lp__sdfrtp_2  VNB VPB SCE D SCD RESET_B CLK VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* CLK	CLK
* RESET_B	RESET_B
* SCD	SCD
* D	D
* SCE	SCE
* VPB	VPB
* VNB	VNB
MM1023 N_VGND_M1023_d N_SCE_M1023_g N_A_35_74#_M1023_s VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.1113 PD=1.37 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1003 noxref_25 N_A_35_74#_M1003_g N_noxref_24_M1003_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1113 PD=0.63 PS=1.37 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.6 A=0.063 P=1.14 MULT=1
MM1033 N_A_380_50#_M1033_d N_D_M1033_g noxref_25 VNB NSHORT L=0.15 W=0.42
+ AD=0.129575 AS=0.0441 PD=1.085 PS=0.63 NRD=34.284 NRS=14.28 M=1 R=2.8
+ SA=75000.6 SB=75001.2 A=0.063 P=1.14 MULT=1
MM1039 noxref_26 N_SCE_M1039_g N_A_380_50#_M1033_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.129575 PD=0.63 PS=1.085 NRD=14.28 NRS=32.856 M=1 R=2.8
+ SA=75000.9 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1000 N_noxref_24_M1000_d N_SCD_M1000_g noxref_26 VNB NSHORT L=0.15 W=0.42
+ AD=0.06195 AS=0.0441 PD=0.715 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.2
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1019 N_VGND_M1019_d N_RESET_B_M1019_g N_noxref_24_M1000_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1386 AS=0.06195 PD=1.5 PS=0.715 NRD=18.564 NRS=4.284 M=1 R=2.8
+ SA=75001.7 SB=75000.3 A=0.063 P=1.14 MULT=1
MM1031 N_A_808_463#_M1031_d N_A_864_255#_M1031_g N_A_380_50#_M1031_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.0588 AS=0.1596 PD=0.7 PS=1.6 NRD=0 NRS=30 M=1 R=2.8
+ SA=75000.3 SB=75004.8 A=0.063 P=1.14 MULT=1
MM1036 A_991_119# N_A_756_265#_M1036_g N_A_808_463#_M1031_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0672 AS=0.0588 PD=0.74 PS=0.7 NRD=30 NRS=0 M=1 R=2.8 SA=75000.7
+ SB=75004.4 A=0.063 P=1.14 MULT=1
MM1005 A_1085_119# N_A_936_333#_M1005_g A_991_119# VNB NSHORT L=0.15 W=0.42
+ AD=0.0777 AS=0.0672 PD=0.81 PS=0.74 NRD=37.14 NRS=30 M=1 R=2.8 SA=75001.2
+ SB=75003.9 A=0.063 P=1.14 MULT=1
MM1037 N_VGND_M1037_d N_RESET_B_M1037_g A_1085_119# VNB NSHORT L=0.15 W=0.42
+ AD=0.108804 AS=0.0777 PD=0.915283 PS=0.81 NRD=68.568 NRS=37.14 M=1 R=2.8
+ SA=75001.6 SB=75003.6 A=0.063 P=1.14 MULT=1
MM1030 N_A_936_333#_M1030_d N_A_808_463#_M1030_g N_VGND_M1037_d VNB NSHORT
+ L=0.15 W=0.64 AD=0.0896 AS=0.165796 PD=0.92 PS=1.39472 NRD=0 NRS=0 M=1
+ R=4.26667 SA=75001.6 SB=75002.1 A=0.096 P=1.58 MULT=1
MM1015 N_A_1406_69#_M1015_d N_A_756_265#_M1015_g N_A_936_333#_M1030_d VNB NSHORT
+ L=0.15 W=0.64 AD=0.234264 AS=0.0896 PD=1.72075 PS=0.92 NRD=0 NRS=0 M=1
+ R=4.26667 SA=75002 SB=75001.7 A=0.096 P=1.58 MULT=1
MM1027 A_1593_113# N_A_864_255#_M1027_g N_A_1406_69#_M1015_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.153736 PD=0.63 PS=1.12925 NRD=14.28 NRS=145.704 M=1
+ R=2.8 SA=75003.6 SB=75001.6 A=0.063 P=1.14 MULT=1
MM1017 N_VGND_M1017_d N_A_1635_21#_M1017_g A_1593_113# VNB NSHORT L=0.15 W=0.42
+ AD=0.12345 AS=0.0441 PD=1.02 PS=0.63 NRD=48.564 NRS=14.28 M=1 R=2.8 SA=75004
+ SB=75001.2 A=0.063 P=1.14 MULT=1
MM1034 A_1809_119# N_RESET_B_M1034_g N_VGND_M1017_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.12345 PD=0.63 PS=1.02 NRD=14.28 NRS=34.284 M=1 R=2.8 SA=75004.5
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1040 N_A_1635_21#_M1040_d N_A_1406_69#_M1040_g A_1809_119# VNB NSHORT L=0.15
+ W=0.42 AD=0.1113 AS=0.0441 PD=1.37 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8
+ SA=75004.9 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1006 N_VGND_M1006_d N_A_864_255#_M1006_g N_A_756_265#_M1006_s VNB NSHORT
+ L=0.15 W=0.84 AD=0.20075 AS=0.2394 PD=1.39 PS=2.25 NRD=12.132 NRS=0 M=1 R=5.6
+ SA=75000.2 SB=75000.8 A=0.126 P=1.98 MULT=1
MM1008 N_A_864_255#_M1008_d N_CLK_M1008_g N_VGND_M1006_d VNB NSHORT L=0.15
+ W=0.84 AD=0.2394 AS=0.20075 PD=2.25 PS=1.39 NRD=0 NRS=12.132 M=1 R=5.6
+ SA=75000.8 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1011 N_VGND_M1011_d N_A_1406_69#_M1011_g N_A_2431_47#_M1011_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.0854 AS=0.1113 PD=0.8 PS=1.37 NRD=19.992 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1024 N_Q_M1024_d N_A_2431_47#_M1024_g N_VGND_M1011_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1708 PD=1.12 PS=1.6 NRD=0 NRS=1.428 M=1 R=5.6 SA=75000.4
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1041 N_Q_M1024_d N_A_2431_47#_M1041_g N_VGND_M1041_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.9
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1022 N_VPWR_M1022_d N_SCE_M1022_g N_A_35_74#_M1022_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0896 AS=0.1696 PD=0.92 PS=1.81 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75003.6 A=0.096 P=1.58 MULT=1
MM1007 A_332_468# N_SCE_M1007_g N_VPWR_M1022_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0672 AS=0.0896 PD=0.85 PS=0.92 NRD=15.3857 NRS=0 M=1 R=4.26667 SA=75000.6
+ SB=75003.2 A=0.096 P=1.58 MULT=1
MM1032 N_A_380_50#_M1032_d N_D_M1032_g A_332_468# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0896 AS=0.0672 PD=0.92 PS=0.85 NRD=0 NRS=15.3857 M=1 R=4.26667 SA=75001
+ SB=75002.8 A=0.096 P=1.58 MULT=1
MM1018 A_490_468# N_A_35_74#_M1018_g N_A_380_50#_M1032_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1024 AS=0.0896 PD=0.96 PS=0.92 NRD=32.308 NRS=0 M=1 R=4.26667
+ SA=75001.4 SB=75002.4 A=0.096 P=1.58 MULT=1
MM1012 N_VPWR_M1012_d N_SCD_M1012_g A_490_468# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.143275 AS=0.1024 PD=1.11 PS=0.96 NRD=23.0687 NRS=32.308 M=1 R=4.26667
+ SA=75001.9 SB=75001.9 A=0.096 P=1.58 MULT=1
MM1026 N_A_380_50#_M1026_d N_RESET_B_M1026_g N_VPWR_M1012_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.130294 AS=0.143275 PD=1.22566 PS=1.11 NRD=14.6174 NRS=27.6982 M=1
+ R=4.26667 SA=75002.4 SB=75001.4 A=0.096 P=1.58 MULT=1
MM1016 N_A_808_463#_M1016_d N_A_756_265#_M1016_g N_A_380_50#_M1026_d VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.0588 AS=0.0855057 PD=0.7 PS=0.80434 NRD=0 NRS=23.443 M=1
+ R=2.8 SA=75002.9 SB=75001.5 A=0.063 P=1.14 MULT=1
MM1001 A_894_463# N_A_864_255#_M1001_g N_A_808_463#_M1016_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=23.443 NRS=0 M=1 R=2.8
+ SA=75003.3 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1004 N_VPWR_M1004_d N_A_936_333#_M1004_g A_894_463# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0819 AS=0.0441 PD=0.81 PS=0.63 NRD=23.443 NRS=23.443 M=1 R=2.8 SA=75003.7
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1013 N_A_808_463#_M1013_d N_RESET_B_M1013_g N_VPWR_M1004_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1113 AS=0.0819 PD=1.37 PS=0.81 NRD=0 NRS=28.1316 M=1 R=2.8
+ SA=75004.2 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1025 N_A_936_333#_M1025_d N_A_808_463#_M1025_g N_VPWR_M1025_s VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.1176 AS=0.3399 PD=1.12 PS=2.7 NRD=0 NRS=23.443 M=1 R=5.6
+ SA=75000.3 SB=75000.9 A=0.126 P=1.98 MULT=1
MM1009 N_A_1406_69#_M1009_d N_A_864_255#_M1009_g N_A_936_333#_M1025_d VPB
+ PHIGHVT L=0.15 W=0.84 AD=0.291567 AS=0.1176 PD=2.22 PS=1.12 NRD=9.3772 NRS=0
+ M=1 R=5.6 SA=75000.7 SB=75000.5 A=0.126 P=1.98 MULT=1
MM1021 A_1569_534# N_A_756_265#_M1021_g N_A_1406_69#_M1009_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0924 AS=0.145783 PD=0.86 PS=1.11 NRD=77.3816 NRS=136.994 M=1 R=2.8
+ SA=75000.4 SB=75002.2 A=0.063 P=1.14 MULT=1
MM1035 N_VPWR_M1035_d N_A_1635_21#_M1035_g A_1569_534# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.1575 AS=0.0924 PD=1.17 PS=0.86 NRD=0 NRS=77.3816 M=1 R=2.8 SA=75001
+ SB=75001.6 A=0.063 P=1.14 MULT=1
MM1014 N_A_1635_21#_M1014_d N_RESET_B_M1014_g N_VPWR_M1035_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0588 AS=0.1575 PD=0.7 PS=1.17 NRD=0 NRS=32.8202 M=1 R=2.8
+ SA=75001.9 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1038 N_VPWR_M1038_d N_A_1406_69#_M1038_g N_A_1635_21#_M1014_d VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.1596 AS=0.0588 PD=1.6 PS=0.7 NRD=49.25 NRS=0 M=1 R=2.8
+ SA=75002.4 SB=75000.3 A=0.063 P=1.14 MULT=1
MM1002 N_VPWR_M1002_d N_A_864_255#_M1002_g N_A_756_265#_M1002_s VPB PHIGHVT
+ L=0.15 W=1.26 AD=0.27405 AS=0.3339 PD=1.695 PS=3.05 NRD=7.0329 NRS=0 M=1 R=8.4
+ SA=75000.2 SB=75000.8 A=0.189 P=2.82 MULT=1
MM1020 N_A_864_255#_M1020_d N_CLK_M1020_g N_VPWR_M1002_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.27405 PD=3.05 PS=1.695 NRD=0 NRS=17.1981 M=1 R=8.4
+ SA=75000.8 SB=75000.2 A=0.189 P=2.82 MULT=1
MM1028 N_VPWR_M1028_d N_A_1406_69#_M1028_g N_A_2431_47#_M1028_s VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.132952 AS=0.1696 PD=1.09137 PS=1.81 NRD=43.0839 NRS=0 M=1
+ R=4.26667 SA=75000.2 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1010 N_VPWR_M1028_d N_A_2431_47#_M1010_g N_Q_M1010_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.261748 AS=0.1764 PD=2.14863 PS=1.54 NRD=4.1567 NRS=0 M=1 R=8.4 SA=75000.4
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1029 N_VPWR_M1029_d N_A_2431_47#_M1029_g N_Q_M1010_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.9
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX42_noxref VNB VPB NWDIODE A=26.6695 P=32.33
c_282 VPB 0 1.04785e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_lp__sdfrtp_2.pxi.spice"
*
.ends
*
*
