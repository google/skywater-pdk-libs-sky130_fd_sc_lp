* File: sky130_fd_sc_lp__a211oi_0.pex.spice
* Created: Wed Sep  2 09:17:57 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A211OI_0%A2 2 3 4 7 11 15 18 20 21 22 27
c39 15 0 1.46445e-19 $X=0.27 $Y=1.51
r40 21 22 12.5413 $w=3.38e-07 $l=3.7e-07 $layer=LI1_cond $X=0.255 $Y=1.295
+ $X2=0.255 $Y2=1.665
r41 20 21 12.5413 $w=3.38e-07 $l=3.7e-07 $layer=LI1_cond $X=0.255 $Y=0.925
+ $X2=0.255 $Y2=1.295
r42 20 27 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.27
+ $Y=1.005 $X2=0.27 $Y2=1.005
r43 16 18 135.883 $w=1.5e-07 $l=2.65e-07 $layer=POLY_cond $X=0.36 $Y=2.19
+ $X2=0.625 $Y2=2.19
r44 14 27 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.27 $Y=1.345
+ $X2=0.27 $Y2=1.005
r45 14 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.27 $Y=1.345
+ $X2=0.27 $Y2=1.51
r46 13 27 6.99445 $w=3.3e-07 $l=4e-08 $layer=POLY_cond $X=0.27 $Y=0.965 $X2=0.27
+ $Y2=1.005
r47 9 11 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=0.665 $Y=0.815
+ $X2=0.665 $Y2=0.445
r48 5 18 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.625 $Y=2.265
+ $X2=0.625 $Y2=2.19
r49 5 7 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=0.625 $Y=2.265 $X2=0.625
+ $Y2=2.735
r50 4 13 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=0.435 $Y=0.89
+ $X2=0.27 $Y2=0.965
r51 3 9 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.59 $Y=0.89
+ $X2=0.665 $Y2=0.815
r52 3 4 79.4787 $w=1.5e-07 $l=1.55e-07 $layer=POLY_cond $X=0.59 $Y=0.89
+ $X2=0.435 $Y2=0.89
r53 2 16 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.36 $Y=2.115
+ $X2=0.36 $Y2=2.19
r54 2 15 310.223 $w=1.5e-07 $l=6.05e-07 $layer=POLY_cond $X=0.36 $Y=2.115
+ $X2=0.36 $Y2=1.51
.ends

.subckt PM_SKY130_FD_SC_LP__A211OI_0%A1 3 7 9 10 11 16
c40 7 0 1.12335e-19 $X=1.055 $Y=2.735
r41 16 19 88.6355 $w=4.55e-07 $l=5.05e-07 $layer=POLY_cond $X=0.902 $Y=1.37
+ $X2=0.902 $Y2=1.875
r42 16 18 47.0767 $w=4.55e-07 $l=1.65e-07 $layer=POLY_cond $X=0.902 $Y=1.37
+ $X2=0.902 $Y2=1.205
r43 16 17 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.84
+ $Y=1.37 $X2=0.84 $Y2=1.37
r44 11 17 8.83041 $w=3.83e-07 $l=2.95e-07 $layer=LI1_cond $X=0.787 $Y=1.665
+ $X2=0.787 $Y2=1.37
r45 10 17 2.24502 $w=3.83e-07 $l=7.5e-08 $layer=LI1_cond $X=0.787 $Y=1.295
+ $X2=0.787 $Y2=1.37
r46 9 10 11.0754 $w=3.83e-07 $l=3.7e-07 $layer=LI1_cond $X=0.787 $Y=0.925
+ $X2=0.787 $Y2=1.295
r47 7 19 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=1.055 $Y=2.735
+ $X2=1.055 $Y2=1.875
r48 3 18 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=1.055 $Y=0.445
+ $X2=1.055 $Y2=1.205
.ends

.subckt PM_SKY130_FD_SC_LP__A211OI_0%B1 3 6 9 11 12 13 17
c38 12 0 1.05268e-19 $X=1.68 $Y=1.295
r39 17 19 46.536 $w=4.35e-07 $l=1.65e-07 $layer=POLY_cond $X=1.627 $Y=1.32
+ $X2=1.627 $Y2=1.155
r40 12 13 12.3595 $w=3.43e-07 $l=3.7e-07 $layer=LI1_cond $X=1.642 $Y=1.295
+ $X2=1.642 $Y2=1.665
r41 12 17 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.68
+ $Y=1.32 $X2=1.68 $Y2=1.32
r42 9 11 466.617 $w=1.5e-07 $l=9.1e-07 $layer=POLY_cond $X=1.485 $Y=2.735
+ $X2=1.485 $Y2=1.825
r43 6 11 53.1843 $w=4.35e-07 $l=2.17e-07 $layer=POLY_cond $X=1.627 $Y=1.608
+ $X2=1.627 $Y2=1.825
r44 5 17 6.64828 $w=4.35e-07 $l=5.2e-08 $layer=POLY_cond $X=1.627 $Y=1.372
+ $X2=1.627 $Y2=1.32
r45 5 6 30.1729 $w=4.35e-07 $l=2.36e-07 $layer=POLY_cond $X=1.627 $Y=1.372
+ $X2=1.627 $Y2=1.608
r46 3 19 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=1.485 $Y=0.445
+ $X2=1.485 $Y2=1.155
.ends

.subckt PM_SKY130_FD_SC_LP__A211OI_0%C1 3 5 7 8 9 10 11 15 17 18 19 20 21 22 23
+ 24 31
c46 9 0 1.05268e-19 $X=1.95 $Y=2.14
r47 31 32 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.495
+ $Y=1.375 $X2=2.495 $Y2=1.375
r48 23 24 10.4001 $w=4.08e-07 $l=3.7e-07 $layer=LI1_cond $X=2.59 $Y=2.405
+ $X2=2.59 $Y2=2.775
r49 22 23 10.4001 $w=4.08e-07 $l=3.7e-07 $layer=LI1_cond $X=2.59 $Y=2.035
+ $X2=2.59 $Y2=2.405
r50 21 22 10.4001 $w=4.08e-07 $l=3.7e-07 $layer=LI1_cond $X=2.59 $Y=1.665
+ $X2=2.59 $Y2=2.035
r51 21 32 8.15143 $w=4.08e-07 $l=2.9e-07 $layer=LI1_cond $X=2.59 $Y=1.665
+ $X2=2.59 $Y2=1.375
r52 20 32 2.24867 $w=4.08e-07 $l=8e-08 $layer=LI1_cond $X=2.59 $Y=1.295 $X2=2.59
+ $Y2=1.375
r53 18 31 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.495 $Y=1.715
+ $X2=2.495 $Y2=1.375
r54 18 19 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.495 $Y=1.715
+ $X2=2.495 $Y2=1.88
r55 17 31 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.495 $Y=1.21
+ $X2=2.495 $Y2=1.375
r56 15 19 94.8617 $w=1.5e-07 $l=1.85e-07 $layer=POLY_cond $X=2.405 $Y=2.065
+ $X2=2.405 $Y2=1.88
r57 12 17 151.266 $w=1.5e-07 $l=2.95e-07 $layer=POLY_cond $X=2.405 $Y=0.915
+ $X2=2.405 $Y2=1.21
r58 10 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.33 $Y=0.84
+ $X2=2.405 $Y2=0.915
r59 10 11 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=2.33 $Y=0.84 $X2=1.99
+ $Y2=0.84
r60 8 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.33 $Y=2.14
+ $X2=2.405 $Y2=2.065
r61 8 9 194.851 $w=1.5e-07 $l=3.8e-07 $layer=POLY_cond $X=2.33 $Y=2.14 $X2=1.95
+ $Y2=2.14
r62 5 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.915 $Y=0.765
+ $X2=1.99 $Y2=0.84
r63 5 7 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.915 $Y=0.765
+ $X2=1.915 $Y2=0.445
r64 1 9 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.875 $Y=2.215
+ $X2=1.95 $Y2=2.14
r65 1 3 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=1.875 $Y=2.215
+ $X2=1.875 $Y2=2.735
.ends

.subckt PM_SKY130_FD_SC_LP__A211OI_0%A_57_483# 1 2 9 11 12 15
c28 12 0 1.46445e-19 $X=0.54 $Y=2.135
c29 9 0 1.12335e-19 $X=0.41 $Y=2.56
r30 13 15 13.0871 $w=2.93e-07 $l=3.35e-07 $layer=LI1_cond $X=1.287 $Y=2.225
+ $X2=1.287 $Y2=2.56
r31 11 13 7.34943 $w=1.8e-07 $l=1.86652e-07 $layer=LI1_cond $X=1.14 $Y=2.135
+ $X2=1.287 $Y2=2.225
r32 11 12 36.9697 $w=1.78e-07 $l=6e-07 $layer=LI1_cond $X=1.14 $Y=2.135 $X2=0.54
+ $Y2=2.135
r33 7 12 7.34943 $w=1.8e-07 $l=1.87681e-07 $layer=LI1_cond $X=0.392 $Y=2.225
+ $X2=0.54 $Y2=2.135
r34 7 9 13.0871 $w=2.93e-07 $l=3.35e-07 $layer=LI1_cond $X=0.392 $Y=2.225
+ $X2=0.392 $Y2=2.56
r35 2 15 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=1.13
+ $Y=2.415 $X2=1.27 $Y2=2.56
r36 1 9 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.285
+ $Y=2.415 $X2=0.41 $Y2=2.56
.ends

.subckt PM_SKY130_FD_SC_LP__A211OI_0%VPWR 1 8 10 17 18 21
r26 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r27 17 18 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r28 15 22 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r29 14 17 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r30 14 15 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r31 12 21 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.97 $Y=3.33 $X2=0.84
+ $Y2=3.33
r32 12 14 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=0.97 $Y=3.33 $X2=1.2
+ $Y2=3.33
r33 10 18 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=2.64 $Y2=3.33
r34 10 15 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=1.2 $Y2=3.33
r35 6 21 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=0.84 $Y=3.245
+ $X2=0.84 $Y2=3.33
r36 6 8 30.3624 $w=2.58e-07 $l=6.85e-07 $layer=LI1_cond $X=0.84 $Y=3.245
+ $X2=0.84 $Y2=2.56
r37 1 8 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=0.7
+ $Y=2.415 $X2=0.84 $Y2=2.56
.ends

.subckt PM_SKY130_FD_SC_LP__A211OI_0%Y 1 2 3 12 14 15 16 18 22 23 25
r48 25 36 2.76533 $w=7.5e-07 $l=1.7e-07 $layer=LI1_cond $X=2.64 $Y=0.66 $X2=2.47
+ $Y2=0.66
r49 23 36 5.04267 $w=7.5e-07 $l=3.1e-07 $layer=LI1_cond $X=2.16 $Y=0.66 $X2=2.47
+ $Y2=0.66
r50 23 31 0.976 $w=7.5e-07 $l=6e-08 $layer=LI1_cond $X=2.16 $Y=0.66 $X2=2.1
+ $Y2=0.66
r51 20 31 7.80943 $w=2.3e-07 $l=3.8e-07 $layer=LI1_cond $X=2.1 $Y=1.04 $X2=2.1
+ $Y2=0.66
r52 20 22 67.8939 $w=2.28e-07 $l=1.355e-06 $layer=LI1_cond $X=2.1 $Y=1.04
+ $X2=2.1 $Y2=2.395
r53 16 22 6.28811 $w=2.88e-07 $l=1.45e-07 $layer=LI1_cond $X=2.07 $Y=2.54
+ $X2=2.07 $Y2=2.395
r54 16 18 0.794788 $w=2.88e-07 $l=2e-08 $layer=LI1_cond $X=2.07 $Y=2.54 $X2=2.07
+ $Y2=2.56
r55 14 31 9.13929 $w=7.5e-07 $l=2.73521e-07 $layer=LI1_cond $X=1.985 $Y=0.882
+ $X2=2.1 $Y2=0.66
r56 14 15 31.6497 $w=2.03e-07 $l=5.85e-07 $layer=LI1_cond $X=1.985 $Y=0.882
+ $X2=1.4 $Y2=0.882
r57 10 15 6.90357 $w=2.05e-07 $l=1.68449e-07 $layer=LI1_cond $X=1.275 $Y=0.78
+ $X2=1.4 $Y2=0.882
r58 10 12 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=1.275 $Y=0.78
+ $X2=1.275 $Y2=0.445
r59 3 18 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=1.95
+ $Y=2.415 $X2=2.09 $Y2=2.56
r60 2 36 91 $w=1.7e-07 $l=5.755e-07 $layer=licon1_NDIFF $count=2 $X=1.99
+ $Y=0.235 $X2=2.47 $Y2=0.445
r61 1 12 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.13
+ $Y=0.235 $X2=1.27 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__A211OI_0%VGND 1 2 9 13 16 17 18 23 29 30 33
r36 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r37 30 34 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=1.68
+ $Y2=0
r38 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r39 27 33 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.83 $Y=0 $X2=1.7
+ $Y2=0
r40 27 29 52.8449 $w=1.68e-07 $l=8.1e-07 $layer=LI1_cond $X=1.83 $Y=0 $X2=2.64
+ $Y2=0
r41 25 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r42 23 33 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.57 $Y=0 $X2=1.7
+ $Y2=0
r43 23 25 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=1.57 $Y=0 $X2=1.2
+ $Y2=0
r44 22 26 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r45 21 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r46 18 34 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=1.68
+ $Y2=0
r47 18 26 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=1.2
+ $Y2=0
r48 16 21 3.22941 $w=1.7e-07 $l=4.5e-08 $layer=LI1_cond $X=0.285 $Y=0 $X2=0.24
+ $Y2=0
r49 16 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.285 $Y=0 $X2=0.45
+ $Y2=0
r50 15 25 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=0.615 $Y=0 $X2=1.2
+ $Y2=0
r51 15 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.615 $Y=0 $X2=0.45
+ $Y2=0
r52 11 33 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=1.7 $Y=0.085 $X2=1.7
+ $Y2=0
r53 11 13 15.9569 $w=2.58e-07 $l=3.6e-07 $layer=LI1_cond $X=1.7 $Y=0.085 $X2=1.7
+ $Y2=0.445
r54 7 17 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.45 $Y=0.085 $X2=0.45
+ $Y2=0
r55 7 9 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=0.45 $Y=0.085 $X2=0.45
+ $Y2=0.445
r56 2 13 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.56
+ $Y=0.235 $X2=1.7 $Y2=0.445
r57 1 9 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.325
+ $Y=0.235 $X2=0.45 $Y2=0.445
.ends

