* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__maj3_lp A B C VGND VNB VPB VPWR X
X0 a_548_419# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X1 a_530_68# C VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 VPWR A a_350_419# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X3 a_350_419# C a_29_419# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X4 a_29_419# B a_154_125# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 a_29_419# B a_530_68# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 VGND a_29_419# a_708_68# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 VPWR a_29_419# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X8 VGND A a_350_125# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 a_154_125# A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 a_350_125# C a_29_419# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X11 a_29_419# B a_548_419# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X12 a_708_68# a_29_419# X VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X13 a_29_419# B a_152_419# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X14 a_152_419# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
.ends
