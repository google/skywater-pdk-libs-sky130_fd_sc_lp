* File: sky130_fd_sc_lp__o311ai_m.pxi.spice
* Created: Fri Aug 28 11:15:08 2020
* 
x_PM_SKY130_FD_SC_LP__O311AI_M%A1 N_A1_M1008_g N_A1_M1005_g N_A1_c_68_n
+ N_A1_c_69_n A1 A1 A1 N_A1_c_71_n N_A1_c_72_n PM_SKY130_FD_SC_LP__O311AI_M%A1
x_PM_SKY130_FD_SC_LP__O311AI_M%A2 N_A2_M1001_g N_A2_M1009_g N_A2_c_105_n
+ N_A2_c_107_n A2 PM_SKY130_FD_SC_LP__O311AI_M%A2
x_PM_SKY130_FD_SC_LP__O311AI_M%A3 N_A3_M1002_g N_A3_M1004_g N_A3_c_146_n
+ N_A3_c_150_n N_A3_c_147_n A3 A3 N_A3_c_152_n PM_SKY130_FD_SC_LP__O311AI_M%A3
x_PM_SKY130_FD_SC_LP__O311AI_M%B1 N_B1_M1000_g N_B1_M1006_g B1 B1 B1
+ N_B1_c_192_n PM_SKY130_FD_SC_LP__O311AI_M%B1
x_PM_SKY130_FD_SC_LP__O311AI_M%C1 N_C1_M1007_g N_C1_M1003_g N_C1_c_234_n
+ N_C1_c_235_n N_C1_c_236_n C1 C1 C1 N_C1_c_237_n N_C1_c_238_n N_C1_c_239_n
+ PM_SKY130_FD_SC_LP__O311AI_M%C1
x_PM_SKY130_FD_SC_LP__O311AI_M%VPWR N_VPWR_M1005_s N_VPWR_M1000_d N_VPWR_c_273_n
+ N_VPWR_c_274_n N_VPWR_c_275_n VPWR N_VPWR_c_276_n N_VPWR_c_277_n
+ N_VPWR_c_272_n N_VPWR_c_279_n PM_SKY130_FD_SC_LP__O311AI_M%VPWR
x_PM_SKY130_FD_SC_LP__O311AI_M%Y N_Y_M1007_d N_Y_M1002_d N_Y_M1003_d N_Y_c_319_n
+ N_Y_c_320_n N_Y_c_314_n N_Y_c_365_n N_Y_c_315_n N_Y_c_321_n N_Y_c_316_n
+ N_Y_c_322_n Y Y Y Y PM_SKY130_FD_SC_LP__O311AI_M%Y
x_PM_SKY130_FD_SC_LP__O311AI_M%VGND N_VGND_M1008_s N_VGND_M1009_d N_VGND_c_391_n
+ N_VGND_c_392_n N_VGND_c_393_n VGND N_VGND_c_394_n N_VGND_c_395_n
+ N_VGND_c_396_n N_VGND_c_397_n PM_SKY130_FD_SC_LP__O311AI_M%VGND
x_PM_SKY130_FD_SC_LP__O311AI_M%A_136_82# N_A_136_82#_M1008_d N_A_136_82#_M1004_d
+ N_A_136_82#_c_442_n N_A_136_82#_c_428_n N_A_136_82#_c_429_n
+ N_A_136_82#_c_435_n PM_SKY130_FD_SC_LP__O311AI_M%A_136_82#
cc_1 VNB N_A1_M1005_g 0.0021123f $X=-0.19 $Y=-0.245 $X2=0.665 $Y2=2.225
cc_2 VNB N_A1_c_68_n 0.0260905f $X=-0.19 $Y=-0.245 $X2=0.472 $Y2=1.46
cc_3 VNB N_A1_c_69_n 0.0306304f $X=-0.19 $Y=-0.245 $X2=0.472 $Y2=1.61
cc_4 VNB A1 0.0344779f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_5 VNB N_A1_c_71_n 0.0326182f $X=-0.19 $Y=-0.245 $X2=0.37 $Y2=1.105
cc_6 VNB N_A1_c_72_n 0.0186228f $X=-0.19 $Y=-0.245 $X2=0.442 $Y2=0.94
cc_7 VNB N_A2_M1001_g 0.00694488f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=0.62
cc_8 VNB N_A2_M1009_g 0.0350467f $X=-0.19 $Y=-0.245 $X2=0.665 $Y2=2.225
cc_9 VNB N_A2_c_105_n 0.00850351f $X=-0.19 $Y=-0.245 $X2=0.472 $Y2=1.46
cc_10 VNB N_A3_M1004_g 0.0233532f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A3_c_146_n 0.0186433f $X=-0.19 $Y=-0.245 $X2=0.472 $Y2=1.61
cc_12 VNB N_A3_c_147_n 0.0101198f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_13 VNB N_B1_M1006_g 0.0455879f $X=-0.19 $Y=-0.245 $X2=0.665 $Y2=2.225
cc_14 VNB B1 0.00725959f $X=-0.19 $Y=-0.245 $X2=0.472 $Y2=1.61
cc_15 VNB N_B1_c_192_n 0.014586f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_C1_M1003_g 0.00160246f $X=-0.19 $Y=-0.245 $X2=0.665 $Y2=1.61
cc_17 VNB N_C1_c_234_n 0.0210382f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_C1_c_235_n 0.0373737f $X=-0.19 $Y=-0.245 $X2=0.472 $Y2=1.46
cc_19 VNB N_C1_c_236_n 0.0364663f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_20 VNB N_C1_c_237_n 0.0345008f $X=-0.19 $Y=-0.245 $X2=0.37 $Y2=1.105
cc_21 VNB N_C1_c_238_n 0.001256f $X=-0.19 $Y=-0.245 $X2=0.442 $Y2=0.94
cc_22 VNB N_C1_c_239_n 0.00762655f $X=-0.19 $Y=-0.245 $X2=0.305 $Y2=0.925
cc_23 VNB N_VPWR_c_272_n 0.123877f $X=-0.19 $Y=-0.245 $X2=0.305 $Y2=1.665
cc_24 VNB N_Y_c_314_n 0.0048476f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_Y_c_315_n 0.00904332f $X=-0.19 $Y=-0.245 $X2=0.37 $Y2=1.105
cc_26 VNB N_Y_c_316_n 0.0280035f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB Y 0.00293469f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB Y 0.00242664f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_391_n 0.0157256f $X=-0.19 $Y=-0.245 $X2=0.665 $Y2=2.225
cc_30 VNB N_VGND_c_392_n 0.021474f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_393_n 0.00527219f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_32 VNB N_VGND_c_394_n 0.0158627f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_395_n 0.0447624f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_396_n 0.204624f $X=-0.19 $Y=-0.245 $X2=0.305 $Y2=1.665
cc_35 VNB N_VGND_c_397_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_136_82#_c_428_n 0.01146f $X=-0.19 $Y=-0.245 $X2=0.472 $Y2=1.61
cc_37 VNB N_A_136_82#_c_429_n 0.00309077f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_38 VPB N_A1_M1005_g 0.03349f $X=-0.19 $Y=1.655 $X2=0.665 $Y2=2.225
cc_39 VPB A1 0.0109847f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_40 VPB N_A2_M1001_g 0.0353057f $X=-0.19 $Y=1.655 $X2=0.605 $Y2=0.62
cc_41 VPB N_A2_c_107_n 0.0553099f $X=-0.19 $Y=1.655 $X2=0.472 $Y2=1.61
cc_42 VPB A2 0.00414759f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_43 VPB N_A3_M1002_g 0.0237083f $X=-0.19 $Y=1.655 $X2=0.605 $Y2=0.62
cc_44 VPB N_A3_c_146_n 0.00398183f $X=-0.19 $Y=1.655 $X2=0.472 $Y2=1.61
cc_45 VPB N_A3_c_150_n 0.0103581f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_46 VPB A3 0.0127622f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_47 VPB N_A3_c_152_n 0.0439967f $X=-0.19 $Y=1.655 $X2=0.305 $Y2=0.925
cc_48 VPB N_B1_M1000_g 0.0227744f $X=-0.19 $Y=1.655 $X2=0.605 $Y2=0.94
cc_49 VPB B1 0.00878744f $X=-0.19 $Y=1.655 $X2=0.472 $Y2=1.61
cc_50 VPB N_B1_c_192_n 0.0157365f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_51 VPB N_C1_M1003_g 0.0427388f $X=-0.19 $Y=1.655 $X2=0.665 $Y2=1.61
cc_52 VPB N_C1_c_238_n 0.00586282f $X=-0.19 $Y=1.655 $X2=0.442 $Y2=0.94
cc_53 VPB N_VPWR_c_273_n 0.0133258f $X=-0.19 $Y=1.655 $X2=0.665 $Y2=2.225
cc_54 VPB N_VPWR_c_274_n 0.0378285f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_55 VPB N_VPWR_c_275_n 0.0397098f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_56 VPB N_VPWR_c_276_n 0.0399599f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_57 VPB N_VPWR_c_277_n 0.0213956f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_58 VPB N_VPWR_c_272_n 0.0806306f $X=-0.19 $Y=1.655 $X2=0.305 $Y2=1.665
cc_59 VPB N_VPWR_c_279_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_60 VPB N_Y_c_319_n 0.00502652f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_61 VPB N_Y_c_320_n 0.00302846f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_62 VPB N_Y_c_321_n 0.00511866f $X=-0.19 $Y=1.655 $X2=0.305 $Y2=0.925
cc_63 VPB N_Y_c_322_n 0.00478481f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_64 VPB Y 0.00319533f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_65 VPB Y 4.15375e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_66 N_A1_M1005_g N_A2_M1001_g 0.0330734f $X=0.665 $Y=2.225 $X2=0 $Y2=0
cc_67 A1 N_A2_M1009_g 9.56215e-19 $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_68 N_A1_c_72_n N_A2_M1009_g 0.0330932f $X=0.442 $Y=0.94 $X2=0 $Y2=0
cc_69 N_A1_c_68_n N_A2_c_105_n 0.00412334f $X=0.472 $Y=1.46 $X2=0 $Y2=0
cc_70 N_A1_c_69_n N_A2_c_105_n 0.0330734f $X=0.472 $Y=1.61 $X2=0 $Y2=0
cc_71 N_A1_M1005_g N_A2_c_107_n 0.00889917f $X=0.665 $Y=2.225 $X2=0 $Y2=0
cc_72 N_A1_M1005_g A2 0.00149944f $X=0.665 $Y=2.225 $X2=0 $Y2=0
cc_73 N_A1_M1005_g N_VPWR_c_274_n 0.00982163f $X=0.665 $Y=2.225 $X2=0 $Y2=0
cc_74 N_A1_c_69_n N_VPWR_c_274_n 0.00103848f $X=0.472 $Y=1.61 $X2=0 $Y2=0
cc_75 A1 N_VPWR_c_274_n 0.00978823f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_76 N_A1_M1005_g N_VPWR_c_276_n 2.99266e-19 $X=0.665 $Y=2.225 $X2=0 $Y2=0
cc_77 N_A1_M1005_g N_VPWR_c_272_n 4.05263e-19 $X=0.665 $Y=2.225 $X2=0 $Y2=0
cc_78 N_A1_c_68_n Y 0.0076092f $X=0.472 $Y=1.46 $X2=0 $Y2=0
cc_79 A1 Y 0.01287f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_80 N_A1_M1005_g Y 0.0254625f $X=0.665 $Y=2.225 $X2=0 $Y2=0
cc_81 N_A1_c_68_n Y 0.00193154f $X=0.472 $Y=1.46 $X2=0 $Y2=0
cc_82 N_A1_c_69_n Y 0.00523259f $X=0.472 $Y=1.61 $X2=0 $Y2=0
cc_83 A1 Y 0.0254845f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_84 N_A1_M1005_g Y 0.00516388f $X=0.665 $Y=2.225 $X2=0 $Y2=0
cc_85 A1 N_VGND_c_392_n 0.0195848f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_86 N_A1_c_71_n N_VGND_c_392_n 0.00340418f $X=0.37 $Y=1.105 $X2=0 $Y2=0
cc_87 N_A1_c_72_n N_VGND_c_392_n 0.00995023f $X=0.442 $Y=0.94 $X2=0 $Y2=0
cc_88 N_A1_c_72_n N_VGND_c_393_n 6.8348e-19 $X=0.442 $Y=0.94 $X2=0 $Y2=0
cc_89 N_A1_c_72_n N_VGND_c_394_n 0.00455951f $X=0.442 $Y=0.94 $X2=0 $Y2=0
cc_90 A1 N_VGND_c_396_n 0.00361332f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_91 N_A1_c_72_n N_VGND_c_396_n 0.00447788f $X=0.442 $Y=0.94 $X2=0 $Y2=0
cc_92 A1 N_A_136_82#_c_429_n 0.0102309f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_93 N_A1_c_72_n N_A_136_82#_c_429_n 0.00183015f $X=0.442 $Y=0.94 $X2=0 $Y2=0
cc_94 N_A2_c_107_n N_A3_M1002_g 0.0425291f $X=0.95 $Y=2.94 $X2=0 $Y2=0
cc_95 N_A2_M1009_g N_A3_M1004_g 0.0223441f $X=1.035 $Y=0.62 $X2=0 $Y2=0
cc_96 N_A2_M1001_g N_A3_c_146_n 0.0115393f $X=1.025 $Y=2.225 $X2=0 $Y2=0
cc_97 N_A2_c_105_n N_A3_c_146_n 0.011329f $X=1.03 $Y=1.515 $X2=0 $Y2=0
cc_98 N_A2_M1001_g N_A3_c_150_n 0.0425291f $X=1.025 $Y=2.225 $X2=0 $Y2=0
cc_99 N_A2_M1009_g N_A3_c_147_n 0.011329f $X=1.035 $Y=0.62 $X2=0 $Y2=0
cc_100 N_A2_M1001_g A3 0.00289649f $X=1.025 $Y=2.225 $X2=0 $Y2=0
cc_101 A2 A3 0.0271391f $X=0.635 $Y=2.69 $X2=0 $Y2=0
cc_102 N_A2_M1001_g B1 0.00190431f $X=1.025 $Y=2.225 $X2=0 $Y2=0
cc_103 N_A2_M1001_g N_VPWR_c_274_n 0.00319843f $X=1.025 $Y=2.225 $X2=0 $Y2=0
cc_104 N_A2_c_107_n N_VPWR_c_274_n 0.00901957f $X=0.95 $Y=2.94 $X2=0 $Y2=0
cc_105 A2 N_VPWR_c_274_n 0.0246768f $X=0.635 $Y=2.69 $X2=0 $Y2=0
cc_106 N_A2_c_107_n N_VPWR_c_276_n 0.011133f $X=0.95 $Y=2.94 $X2=0 $Y2=0
cc_107 A2 N_VPWR_c_276_n 0.015991f $X=0.635 $Y=2.69 $X2=0 $Y2=0
cc_108 N_A2_c_107_n N_VPWR_c_272_n 0.0129615f $X=0.95 $Y=2.94 $X2=0 $Y2=0
cc_109 A2 N_VPWR_c_272_n 0.0106361f $X=0.635 $Y=2.69 $X2=0 $Y2=0
cc_110 N_A2_M1001_g N_Y_c_321_n 0.0154897f $X=1.025 $Y=2.225 $X2=0 $Y2=0
cc_111 N_A2_c_107_n N_Y_c_321_n 0.00122708f $X=0.95 $Y=2.94 $X2=0 $Y2=0
cc_112 A2 N_Y_c_321_n 0.00880675f $X=0.635 $Y=2.69 $X2=0 $Y2=0
cc_113 N_A2_M1009_g N_Y_c_316_n 0.00773845f $X=1.035 $Y=0.62 $X2=0 $Y2=0
cc_114 N_A2_c_105_n N_Y_c_316_n 0.00770324f $X=1.03 $Y=1.515 $X2=0 $Y2=0
cc_115 N_A2_c_105_n Y 0.016982f $X=1.03 $Y=1.515 $X2=0 $Y2=0
cc_116 N_A2_c_107_n Y 5.08257e-19 $X=0.95 $Y=2.94 $X2=0 $Y2=0
cc_117 A2 Y 0.0124104f $X=0.635 $Y=2.69 $X2=0 $Y2=0
cc_118 N_A2_M1009_g N_VGND_c_392_n 6.8348e-19 $X=1.035 $Y=0.62 $X2=0 $Y2=0
cc_119 N_A2_M1009_g N_VGND_c_393_n 0.00800037f $X=1.035 $Y=0.62 $X2=0 $Y2=0
cc_120 N_A2_M1009_g N_VGND_c_394_n 0.00455951f $X=1.035 $Y=0.62 $X2=0 $Y2=0
cc_121 N_A2_M1009_g N_VGND_c_396_n 0.00447788f $X=1.035 $Y=0.62 $X2=0 $Y2=0
cc_122 N_A2_M1009_g N_A_136_82#_c_428_n 0.011321f $X=1.035 $Y=0.62 $X2=0 $Y2=0
cc_123 N_A3_M1002_g N_B1_M1000_g 0.0135092f $X=1.385 $Y=2.225 $X2=0 $Y2=0
cc_124 N_A3_c_150_n N_B1_M1000_g 0.0118733f $X=1.405 $Y=1.905 $X2=0 $Y2=0
cc_125 A3 N_B1_M1000_g 8.39511e-19 $X=1.595 $Y=2.69 $X2=0 $Y2=0
cc_126 N_A3_M1004_g N_B1_M1006_g 0.0284211f $X=1.465 $Y=0.62 $X2=0 $Y2=0
cc_127 N_A3_c_146_n N_B1_M1006_g 0.00991391f $X=1.405 $Y=1.755 $X2=0 $Y2=0
cc_128 N_A3_c_146_n B1 0.011382f $X=1.405 $Y=1.755 $X2=0 $Y2=0
cc_129 N_A3_c_150_n B1 0.001503f $X=1.405 $Y=1.905 $X2=0 $Y2=0
cc_130 N_A3_c_147_n B1 2.03629e-19 $X=1.445 $Y=1.26 $X2=0 $Y2=0
cc_131 N_A3_c_146_n N_B1_c_192_n 0.0118733f $X=1.405 $Y=1.755 $X2=0 $Y2=0
cc_132 N_A3_M1002_g N_VPWR_c_275_n 0.00382443f $X=1.385 $Y=2.225 $X2=0 $Y2=0
cc_133 A3 N_VPWR_c_275_n 0.0281844f $X=1.595 $Y=2.69 $X2=0 $Y2=0
cc_134 N_A3_c_152_n N_VPWR_c_275_n 0.00416045f $X=1.505 $Y=2.94 $X2=0 $Y2=0
cc_135 A3 N_VPWR_c_276_n 0.0323672f $X=1.595 $Y=2.69 $X2=0 $Y2=0
cc_136 N_A3_c_152_n N_VPWR_c_276_n 0.00671525f $X=1.505 $Y=2.94 $X2=0 $Y2=0
cc_137 A3 N_VPWR_c_272_n 0.0224213f $X=1.595 $Y=2.69 $X2=0 $Y2=0
cc_138 N_A3_c_152_n N_VPWR_c_272_n 0.0087784f $X=1.505 $Y=2.94 $X2=0 $Y2=0
cc_139 A3 N_Y_c_319_n 0.00133974f $X=1.595 $Y=2.69 $X2=0 $Y2=0
cc_140 N_A3_M1002_g N_Y_c_320_n 0.00272888f $X=1.385 $Y=2.225 $X2=0 $Y2=0
cc_141 N_A3_M1002_g N_Y_c_321_n 0.0112485f $X=1.385 $Y=2.225 $X2=0 $Y2=0
cc_142 A3 N_Y_c_321_n 0.0404028f $X=1.595 $Y=2.69 $X2=0 $Y2=0
cc_143 N_A3_c_152_n N_Y_c_321_n 0.00127779f $X=1.505 $Y=2.94 $X2=0 $Y2=0
cc_144 N_A3_c_146_n N_Y_c_316_n 0.00663758f $X=1.405 $Y=1.755 $X2=0 $Y2=0
cc_145 N_A3_c_147_n N_Y_c_316_n 0.00519752f $X=1.445 $Y=1.26 $X2=0 $Y2=0
cc_146 N_A3_M1004_g N_VGND_c_393_n 0.00819747f $X=1.465 $Y=0.62 $X2=0 $Y2=0
cc_147 N_A3_M1004_g N_VGND_c_395_n 0.00455951f $X=1.465 $Y=0.62 $X2=0 $Y2=0
cc_148 N_A3_M1004_g N_VGND_c_396_n 0.00447788f $X=1.465 $Y=0.62 $X2=0 $Y2=0
cc_149 N_A3_M1004_g N_A_136_82#_c_428_n 0.0113853f $X=1.465 $Y=0.62 $X2=0 $Y2=0
cc_150 N_A3_c_147_n N_A_136_82#_c_428_n 0.00116041f $X=1.445 $Y=1.26 $X2=0 $Y2=0
cc_151 N_A3_M1004_g N_A_136_82#_c_435_n 2.03427e-19 $X=1.465 $Y=0.62 $X2=0 $Y2=0
cc_152 N_B1_M1000_g N_C1_M1003_g 0.0168637f $X=1.815 $Y=2.225 $X2=0 $Y2=0
cc_153 N_B1_M1006_g N_C1_c_234_n 0.050007f $X=1.895 $Y=0.62 $X2=0 $Y2=0
cc_154 B1 N_C1_c_235_n 2.45628e-19 $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_155 B1 N_C1_c_236_n 0.00162172f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_156 N_B1_c_192_n N_C1_c_236_n 0.0169435f $X=1.905 $Y=1.665 $X2=0 $Y2=0
cc_157 N_B1_M1006_g N_C1_c_237_n 0.0132467f $X=1.895 $Y=0.62 $X2=0 $Y2=0
cc_158 N_B1_M1006_g N_C1_c_238_n 6.37539e-19 $X=1.895 $Y=0.62 $X2=0 $Y2=0
cc_159 B1 N_C1_c_238_n 0.0099345f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_160 N_B1_c_192_n N_C1_c_238_n 4.15568e-19 $X=1.905 $Y=1.665 $X2=0 $Y2=0
cc_161 N_B1_M1000_g N_VPWR_c_275_n 0.00371759f $X=1.815 $Y=2.225 $X2=0 $Y2=0
cc_162 N_B1_M1000_g N_VPWR_c_276_n 0.00249672f $X=1.815 $Y=2.225 $X2=0 $Y2=0
cc_163 N_B1_M1000_g N_VPWR_c_272_n 0.00334041f $X=1.815 $Y=2.225 $X2=0 $Y2=0
cc_164 N_B1_M1000_g N_Y_c_319_n 0.0137659f $X=1.815 $Y=2.225 $X2=0 $Y2=0
cc_165 B1 N_Y_c_319_n 0.0371961f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_166 N_B1_c_192_n N_Y_c_319_n 0.00474835f $X=1.905 $Y=1.665 $X2=0 $Y2=0
cc_167 B1 N_Y_c_320_n 0.0167423f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_168 N_B1_M1006_g N_Y_c_314_n 0.0055697f $X=1.895 $Y=0.62 $X2=0 $Y2=0
cc_169 N_B1_M1000_g N_Y_c_321_n 8.90842e-19 $X=1.815 $Y=2.225 $X2=0 $Y2=0
cc_170 B1 N_Y_c_321_n 0.00890597f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_171 N_B1_M1006_g N_Y_c_316_n 0.0157496f $X=1.895 $Y=0.62 $X2=0 $Y2=0
cc_172 B1 N_Y_c_316_n 0.0734543f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_173 N_B1_c_192_n N_Y_c_316_n 0.00468341f $X=1.905 $Y=1.665 $X2=0 $Y2=0
cc_174 B1 Y 0.00931443f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_175 N_B1_M1006_g N_VGND_c_393_n 0.00114726f $X=1.895 $Y=0.62 $X2=0 $Y2=0
cc_176 N_B1_M1006_g N_VGND_c_395_n 0.00548708f $X=1.895 $Y=0.62 $X2=0 $Y2=0
cc_177 N_B1_M1006_g N_VGND_c_396_n 0.00533081f $X=1.895 $Y=0.62 $X2=0 $Y2=0
cc_178 N_B1_M1006_g N_A_136_82#_c_428_n 0.00217059f $X=1.895 $Y=0.62 $X2=0 $Y2=0
cc_179 N_C1_M1003_g N_VPWR_c_275_n 0.00471632f $X=2.405 $Y=2.225 $X2=0 $Y2=0
cc_180 N_C1_M1003_g N_VPWR_c_277_n 0.00297774f $X=2.405 $Y=2.225 $X2=0 $Y2=0
cc_181 N_C1_M1003_g N_VPWR_c_272_n 0.00400849f $X=2.405 $Y=2.225 $X2=0 $Y2=0
cc_182 N_C1_M1003_g N_Y_c_319_n 0.0188509f $X=2.405 $Y=2.225 $X2=0 $Y2=0
cc_183 N_C1_c_236_n N_Y_c_319_n 0.00124575f $X=2.552 $Y=1.625 $X2=0 $Y2=0
cc_184 N_C1_c_234_n N_Y_c_314_n 0.00735955f $X=2.477 $Y=0.955 $X2=0 $Y2=0
cc_185 N_C1_c_235_n N_Y_c_314_n 0.00788312f $X=2.477 $Y=1.105 $X2=0 $Y2=0
cc_186 N_C1_c_237_n N_Y_c_314_n 0.00253972f $X=2.61 $Y=1.12 $X2=0 $Y2=0
cc_187 N_C1_c_238_n N_Y_c_314_n 0.0100312f $X=2.61 $Y=1.12 $X2=0 $Y2=0
cc_188 N_C1_c_239_n N_Y_c_314_n 0.0140882f $X=2.625 $Y=1.055 $X2=0 $Y2=0
cc_189 N_C1_c_234_n N_Y_c_365_n 0.00523899f $X=2.477 $Y=0.955 $X2=0 $Y2=0
cc_190 N_C1_c_235_n N_Y_c_315_n 0.00660087f $X=2.477 $Y=1.105 $X2=0 $Y2=0
cc_191 N_C1_c_239_n N_Y_c_315_n 0.00788189f $X=2.625 $Y=1.055 $X2=0 $Y2=0
cc_192 N_C1_c_237_n N_Y_c_316_n 0.00559196f $X=2.61 $Y=1.12 $X2=0 $Y2=0
cc_193 N_C1_c_238_n N_Y_c_316_n 0.0125062f $X=2.61 $Y=1.12 $X2=0 $Y2=0
cc_194 N_C1_M1003_g N_Y_c_322_n 9.28094e-19 $X=2.405 $Y=2.225 $X2=0 $Y2=0
cc_195 N_C1_c_236_n N_Y_c_322_n 0.00146803f $X=2.552 $Y=1.625 $X2=0 $Y2=0
cc_196 N_C1_c_238_n N_Y_c_322_n 0.0171108f $X=2.61 $Y=1.12 $X2=0 $Y2=0
cc_197 N_C1_c_234_n N_VGND_c_395_n 0.00400834f $X=2.477 $Y=0.955 $X2=0 $Y2=0
cc_198 N_C1_c_234_n N_VGND_c_396_n 0.00533081f $X=2.477 $Y=0.955 $X2=0 $Y2=0
cc_199 N_C1_c_239_n N_VGND_c_396_n 0.00370453f $X=2.625 $Y=1.055 $X2=0 $Y2=0
cc_200 N_VPWR_M1000_d N_Y_c_319_n 0.00392154f $X=1.89 $Y=2.015 $X2=0 $Y2=0
cc_201 N_VPWR_c_275_n N_Y_c_319_n 0.0254128f $X=2.11 $Y=2.365 $X2=0 $Y2=0
cc_202 N_VPWR_c_275_n N_Y_c_321_n 0.0037449f $X=2.11 $Y=2.365 $X2=0 $Y2=0
cc_203 N_VPWR_c_272_n N_Y_c_321_n 0.00588281f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_204 N_VPWR_c_274_n Y 0.0117101f $X=0.34 $Y=2.29 $X2=0 $Y2=0
cc_205 N_VPWR_c_274_n Y 0.0115071f $X=0.34 $Y=2.29 $X2=0 $Y2=0
cc_206 A_148_403# N_Y_c_321_n 0.00331953f $X=0.74 $Y=2.015 $X2=1.495 $Y2=2.405
cc_207 A_148_403# Y 0.00347104f $X=0.74 $Y=2.015 $X2=0.635 $Y2=1.58
cc_208 A_220_403# N_Y_c_321_n 0.00185966f $X=1.1 $Y=2.015 $X2=1.495 $Y2=2.405
cc_209 N_Y_c_365_n N_VGND_c_395_n 0.00468431f $X=2.345 $Y=0.555 $X2=0 $Y2=0
cc_210 N_Y_c_315_n N_VGND_c_395_n 0.00773979f $X=2.47 $Y=0.555 $X2=0 $Y2=0
cc_211 N_Y_c_365_n N_VGND_c_396_n 0.00572537f $X=2.345 $Y=0.555 $X2=0 $Y2=0
cc_212 N_Y_c_315_n N_VGND_c_396_n 0.00960518f $X=2.47 $Y=0.555 $X2=0 $Y2=0
cc_213 N_Y_c_314_n N_A_136_82#_c_428_n 0.0080348f $X=2.26 $Y=1.21 $X2=0 $Y2=0
cc_214 N_Y_c_316_n N_A_136_82#_c_428_n 0.0577648f $X=2.175 $Y=1.295 $X2=0 $Y2=0
cc_215 N_Y_c_316_n N_A_136_82#_c_429_n 0.00729871f $X=2.175 $Y=1.295 $X2=0 $Y2=0
cc_216 Y N_A_136_82#_c_429_n 0.00570533f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_217 N_Y_c_314_n N_A_136_82#_c_435_n 3.61971e-19 $X=2.26 $Y=1.21 $X2=0 $Y2=0
cc_218 N_VGND_c_394_n N_A_136_82#_c_442_n 0.00412673f $X=1.085 $Y=0 $X2=0 $Y2=0
cc_219 N_VGND_c_396_n N_A_136_82#_c_442_n 0.00545208f $X=2.64 $Y=0 $X2=0 $Y2=0
cc_220 N_VGND_c_393_n N_A_136_82#_c_428_n 0.0200383f $X=1.25 $Y=0.555 $X2=0
+ $Y2=0
cc_221 N_VGND_c_396_n N_A_136_82#_c_428_n 0.0126889f $X=2.64 $Y=0 $X2=0 $Y2=0
cc_222 N_VGND_c_395_n N_A_136_82#_c_435_n 0.00439471f $X=2.64 $Y=0 $X2=0 $Y2=0
cc_223 N_VGND_c_396_n N_A_136_82#_c_435_n 0.00610964f $X=2.64 $Y=0 $X2=0 $Y2=0
