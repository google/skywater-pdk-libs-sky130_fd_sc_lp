* File: sky130_fd_sc_lp__sdlclkp_4.spice
* Created: Wed Sep  2 10:37:18 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__sdlclkp_4.pex.spice"
.subckt sky130_fd_sc_lp__sdlclkp_4  VNB VPB SCE GATE CLK VPWR GCLK VGND
* 
* VGND	VGND
* GCLK	GCLK
* VPWR	VPWR
* CLK	CLK
* GATE	GATE
* SCE	SCE
* VPB	VPB
* VNB	VNB
MM1014 N_A_134_70#_M1014_d N_SCE_M1014_g N_VGND_M1014_s VNB NSHORT L=0.15 W=0.42
+ AD=0.06615 AS=0.1155 PD=0.735 PS=1.39 NRD=0 NRS=2.856 M=1 R=2.8 SA=75000.2
+ SB=75001.2 A=0.063 P=1.14 MULT=1
MM1012 N_VGND_M1012_d N_GATE_M1012_g N_A_134_70#_M1014_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0819 AS=0.06615 PD=0.81 PS=0.735 NRD=17.136 NRS=9.996 M=1 R=2.8
+ SA=75000.7 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1027 N_A_335_70#_M1027_d N_A_252_361#_M1027_g N_VGND_M1012_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1113 AS=0.0819 PD=1.37 PS=0.81 NRD=0 NRS=14.28 M=1 R=2.8
+ SA=75001.2 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1011 N_A_634_133#_M1011_d N_A_252_361#_M1011_g N_A_134_70#_M1011_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.6 A=0.063 P=1.14 MULT=1
MM1016 A_720_133# N_A_335_70#_M1016_g N_A_634_133#_M1011_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75001.2 A=0.063 P=1.14 MULT=1
MM1009 N_VGND_M1009_d N_A_762_107#_M1009_g A_720_133# VNB NSHORT L=0.15 W=0.42
+ AD=0.128233 AS=0.0441 PD=0.95 PS=0.63 NRD=71.508 NRS=14.28 M=1 R=2.8 SA=75001
+ SB=75000.8 A=0.063 P=1.14 MULT=1
MM1004 N_A_762_107#_M1004_d N_A_634_133#_M1004_g N_VGND_M1009_d VNB NSHORT
+ L=0.15 W=0.84 AD=0.2394 AS=0.256467 PD=2.25 PS=1.9 NRD=0 NRS=12.132 M=1 R=5.6
+ SA=75000.9 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1017 N_VGND_M1017_d N_CLK_M1017_g N_A_252_361#_M1017_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0896 AS=0.1113 PD=0.81 PS=1.37 NRD=27.132 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1002 A_1216_47# N_CLK_M1002_g N_VGND_M1017_d VNB NSHORT L=0.15 W=0.84
+ AD=0.0882 AS=0.1792 PD=1.05 PS=1.62 NRD=7.14 NRS=0 M=1 R=5.6 SA=75000.5
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1003 N_A_1275_367#_M1003_d N_A_762_107#_M1003_g A_1216_47# VNB NSHORT L=0.15
+ W=0.84 AD=0.2226 AS=0.0882 PD=2.21 PS=1.05 NRD=0 NRS=7.14 M=1 R=5.6 SA=75000.8
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1006 N_GCLK_M1006_d N_A_1275_367#_M1006_g N_VGND_M1006_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75001.5 A=0.126 P=1.98 MULT=1
MM1010 N_GCLK_M1006_d N_A_1275_367#_M1010_g N_VGND_M1010_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1021 N_GCLK_M1021_d N_A_1275_367#_M1021_g N_VGND_M1010_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.1
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1024 N_GCLK_M1021_d N_A_1275_367#_M1024_g N_VGND_M1024_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75001.5
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1022 A_110_468# N_SCE_M1022_g N_VPWR_M1022_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0672 AS=0.1696 PD=0.85 PS=1.81 NRD=15.3857 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75000.6 A=0.096 P=1.58 MULT=1
MM1019 N_A_134_70#_M1019_d N_GATE_M1019_g A_110_468# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1696 AS=0.0672 PD=1.81 PS=0.85 NRD=0 NRS=15.3857 M=1 R=4.26667 SA=75000.6
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1015 N_A_335_70#_M1015_d N_A_252_361#_M1015_g N_VPWR_M1015_s VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.2112 AS=0.3008 PD=1.94 PS=2.22 NRD=19.9955 NRS=63.0991 M=1
+ R=4.26667 SA=75000.4 SB=75000.3 A=0.096 P=1.58 MULT=1
MM1020 N_A_634_133#_M1020_d N_A_335_70#_M1020_g N_A_134_70#_M1020_s VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.8 A=0.063 P=1.14 MULT=1
MM1025 A_720_463# N_A_252_361#_M1025_g N_A_634_133#_M1020_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=23.443 NRS=0 M=1 R=2.8
+ SA=75000.6 SB=75001.3 A=0.063 P=1.14 MULT=1
MM1000 N_VPWR_M1000_d N_A_762_107#_M1000_g A_720_463# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.125475 AS=0.0441 PD=0.9425 PS=0.63 NRD=114.319 NRS=23.443 M=1 R=2.8
+ SA=75001 SB=75001 A=0.063 P=1.14 MULT=1
MM1005 N_A_762_107#_M1005_d N_A_634_133#_M1005_g N_VPWR_M1000_d VPB PHIGHVT
+ L=0.15 W=1.26 AD=0.3339 AS=0.376425 PD=3.05 PS=2.8275 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.7 SB=75000.2 A=0.189 P=2.82 MULT=1
MM1026 N_VPWR_M1026_d N_CLK_M1026_g N_A_252_361#_M1026_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.136185 AS=0.1696 PD=1.10147 PS=1.81 NRD=48.5605 NRS=0 M=1
+ R=4.26667 SA=75000.2 SB=75003 A=0.096 P=1.58 MULT=1
MM1018 N_A_1275_367#_M1018_d N_CLK_M1018_g N_VPWR_M1026_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.268115 PD=1.54 PS=2.16853 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.5 SB=75002.4 A=0.189 P=2.82 MULT=1
MM1007 N_VPWR_M1007_d N_A_762_107#_M1007_g N_A_1275_367#_M1018_d VPB PHIGHVT
+ L=0.15 W=1.26 AD=0.24255 AS=0.1764 PD=1.645 PS=1.54 NRD=16.4101 NRS=0 M=1
+ R=8.4 SA=75000.9 SB=75002 A=0.189 P=2.82 MULT=1
MM1001 N_GCLK_M1001_d N_A_1275_367#_M1001_g N_VPWR_M1007_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.24255 PD=1.54 PS=1.645 NRD=0 NRS=0 M=1 R=8.4 SA=75001.4
+ SB=75001.5 A=0.189 P=2.82 MULT=1
MM1008 N_GCLK_M1001_d N_A_1275_367#_M1008_g N_VPWR_M1008_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.9
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1013 N_GCLK_M1013_d N_A_1275_367#_M1013_g N_VPWR_M1008_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.3
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1023 N_GCLK_M1013_d N_A_1275_367#_M1023_g N_VPWR_M1023_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75002.7
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX28_noxref VNB VPB NWDIODE A=17.8659 P=23.01
*
.include "sky130_fd_sc_lp__sdlclkp_4.pxi.spice"
*
.ends
*
*
