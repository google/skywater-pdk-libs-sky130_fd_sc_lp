* File: sky130_fd_sc_lp__sdlclkp_2.spice
* Created: Wed Sep  2 10:37:10 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__sdlclkp_2.pex.spice"
.subckt sky130_fd_sc_lp__sdlclkp_2  VNB VPB SCE GATE CLK VPWR GCLK VGND
* 
* VGND	VGND
* GCLK	GCLK
* VPWR	VPWR
* CLK	CLK
* GATE	GATE
* SCE	SCE
* VPB	VPB
* VNB	VNB
MM1005 N_A_110_70#_M1005_d N_SCE_M1005_g N_VGND_M1005_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75001.1
+ A=0.063 P=1.14 MULT=1
MM1010 N_VGND_M1010_d N_GATE_M1010_g N_A_110_70#_M1005_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1020 N_A_282_70#_M1020_d N_A_250_443#_M1020_g N_VGND_M1010_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.1
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1014 N_A_614_133#_M1014_d N_A_250_443#_M1014_g N_A_110_70#_M1014_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.0588 AS=0.1533 PD=0.7 PS=1.57 NRD=0 NRS=22.848 M=1 R=2.8
+ SA=75000.3 SB=75001.6 A=0.063 P=1.14 MULT=1
MM1015 A_700_133# N_A_282_70#_M1015_g N_A_614_133#_M1014_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.7
+ SB=75001.2 A=0.063 P=1.14 MULT=1
MM1013 N_VGND_M1013_d N_A_742_107#_M1013_g A_700_133# VNB NSHORT L=0.15 W=0.42
+ AD=0.123333 AS=0.0441 PD=0.926667 PS=0.63 NRD=68.184 NRS=14.28 M=1 R=2.8
+ SA=75001.1 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1016 N_A_742_107#_M1016_d N_A_614_133#_M1016_g N_VGND_M1013_d VNB NSHORT
+ L=0.15 W=0.84 AD=0.2394 AS=0.246667 PD=2.25 PS=1.85333 NRD=0 NRS=12.132 M=1
+ R=5.6 SA=75001 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1023 N_VGND_M1023_d N_CLK_M1023_g N_A_250_443#_M1023_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1006 A_1174_74# N_CLK_M1006_g N_VGND_M1023_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1008 N_A_1235_429#_M1008_d N_A_742_107#_M1008_g A_1174_74# VNB NSHORT L=0.15
+ W=0.42 AD=0.1113 AS=0.0441 PD=1.37 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1001 N_VGND_M1001_d N_A_1235_429#_M1001_g N_GCLK_M1001_s VNB NSHORT L=0.15
+ W=0.84 AD=0.231 AS=0.1176 PD=2.23 PS=1.12 NRD=1.428 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1012 N_VGND_M1012_d N_A_1235_429#_M1012_g N_GCLK_M1001_s VNB NSHORT L=0.15
+ W=0.84 AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1021 A_110_468# N_SCE_M1021_g N_VPWR_M1021_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0672 AS=0.1696 PD=0.85 PS=1.81 NRD=15.3857 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75000.6 A=0.096 P=1.58 MULT=1
MM1017 N_A_110_70#_M1017_d N_GATE_M1017_g A_110_468# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1696 AS=0.0672 PD=1.81 PS=0.85 NRD=0 NRS=15.3857 M=1 R=4.26667 SA=75000.6
+ SB=75000.2 A=0.096 P=1.58 MULT=1
MM1007 N_A_282_70#_M1007_d N_A_250_443#_M1007_g N_VPWR_M1007_s VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.3136 AS=0.2113 PD=2.26 PS=2.14 NRD=60.0062 NRS=41.5473 M=1
+ R=4.26667 SA=75000.3 SB=75000.4 A=0.096 P=1.58 MULT=1
MM1002 N_A_614_133#_M1002_d N_A_282_70#_M1002_g N_A_110_70#_M1002_s VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.5 A=0.063 P=1.14 MULT=1
MM1018 A_746_457# N_A_250_443#_M1018_g N_A_614_133#_M1002_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=23.443 NRS=0 M=1 R=2.8
+ SA=75000.6 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1011 N_VPWR_M1011_d N_A_742_107#_M1011_g A_746_457# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.095025 AS=0.0441 PD=0.8175 PS=0.63 NRD=0 NRS=23.443 M=1 R=2.8 SA=75001
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1019 N_A_742_107#_M1019_d N_A_614_133#_M1019_g N_VPWR_M1011_d VPB PHIGHVT
+ L=0.15 W=1.26 AD=0.3339 AS=0.285075 PD=3.05 PS=2.4525 NRD=0 NRS=4.9447 M=1
+ R=8.4 SA=75000.6 SB=75000.2 A=0.189 P=2.82 MULT=1
MM1003 N_VPWR_M1003_d N_CLK_M1003_g N_A_250_443#_M1003_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.18575 AS=0.1824 PD=1.39 PS=1.85 NRD=72.3975 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75002.3 A=0.096 P=1.58 MULT=1
MM1022 N_A_1235_429#_M1022_d N_CLK_M1022_g N_VPWR_M1003_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.0896 AS=0.18575 PD=0.92 PS=1.39 NRD=0 NRS=72.3975 M=1 R=4.26667
+ SA=75000.8 SB=75001.8 A=0.096 P=1.58 MULT=1
MM1000 N_VPWR_M1000_d N_A_742_107#_M1000_g N_A_1235_429#_M1022_d VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.179166 AS=0.0896 PD=1.22274 PS=0.92 NRD=0 NRS=0 M=1
+ R=4.26667 SA=75001.2 SB=75001.3 A=0.096 P=1.58 MULT=1
MM1004 N_VPWR_M1000_d N_A_1235_429#_M1004_g N_GCLK_M1004_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.352734 AS=0.1764 PD=2.40726 PS=1.54 NRD=21.4927 NRS=0 M=1 R=8.4
+ SA=75001.1 SB=75000.6 A=0.189 P=2.82 MULT=1
MM1009 N_VPWR_M1009_d N_A_1235_429#_M1009_g N_GCLK_M1004_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.5
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX24_noxref VNB VPB NWDIODE A=15.9375 P=20.83
*
.include "sky130_fd_sc_lp__sdlclkp_2.pxi.spice"
*
.ends
*
*
