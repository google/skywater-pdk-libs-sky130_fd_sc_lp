* File: sky130_fd_sc_lp__o31a_1.pxi.spice
* Created: Fri Aug 28 11:15:23 2020
* 
x_PM_SKY130_FD_SC_LP__O31A_1%A_86_23# N_A_86_23#_M1008_d N_A_86_23#_M1001_d
+ N_A_86_23#_M1005_g N_A_86_23#_M1003_g N_A_86_23#_c_57_n N_A_86_23#_c_58_n
+ N_A_86_23#_c_69_p N_A_86_23#_c_102_p N_A_86_23#_c_109_p N_A_86_23#_c_65_n
+ N_A_86_23#_c_59_n N_A_86_23#_c_60_n N_A_86_23#_c_84_p N_A_86_23#_c_61_n
+ N_A_86_23#_c_62_n PM_SKY130_FD_SC_LP__O31A_1%A_86_23#
x_PM_SKY130_FD_SC_LP__O31A_1%A1 N_A1_M1002_g N_A1_M1007_g A1 A1 N_A1_c_127_n
+ N_A1_c_128_n PM_SKY130_FD_SC_LP__O31A_1%A1
x_PM_SKY130_FD_SC_LP__O31A_1%A2 N_A2_M1000_g N_A2_M1009_g A2 N_A2_c_162_n
+ N_A2_c_163_n PM_SKY130_FD_SC_LP__O31A_1%A2
x_PM_SKY130_FD_SC_LP__O31A_1%A3 N_A3_M1001_g N_A3_M1004_g A3 N_A3_c_200_n
+ N_A3_c_201_n PM_SKY130_FD_SC_LP__O31A_1%A3
x_PM_SKY130_FD_SC_LP__O31A_1%B1 N_B1_M1008_g N_B1_M1006_g B1 N_B1_c_236_n
+ N_B1_c_237_n PM_SKY130_FD_SC_LP__O31A_1%B1
x_PM_SKY130_FD_SC_LP__O31A_1%X N_X_M1005_s N_X_M1003_s X X X X X X X N_X_c_267_n
+ PM_SKY130_FD_SC_LP__O31A_1%X
x_PM_SKY130_FD_SC_LP__O31A_1%VPWR N_VPWR_M1003_d N_VPWR_M1006_d N_VPWR_c_278_n
+ N_VPWR_c_279_n N_VPWR_c_280_n VPWR N_VPWR_c_281_n N_VPWR_c_282_n
+ N_VPWR_c_283_n N_VPWR_c_277_n PM_SKY130_FD_SC_LP__O31A_1%VPWR
x_PM_SKY130_FD_SC_LP__O31A_1%VGND N_VGND_M1005_d N_VGND_M1000_d N_VGND_c_319_n
+ N_VGND_c_320_n VGND N_VGND_c_321_n N_VGND_c_322_n N_VGND_c_323_n
+ N_VGND_c_324_n N_VGND_c_325_n N_VGND_c_326_n PM_SKY130_FD_SC_LP__O31A_1%VGND
x_PM_SKY130_FD_SC_LP__O31A_1%A_275_49# N_A_275_49#_M1002_d N_A_275_49#_M1004_d
+ N_A_275_49#_c_366_n N_A_275_49#_c_362_n N_A_275_49#_c_363_n
+ N_A_275_49#_c_375_n PM_SKY130_FD_SC_LP__O31A_1%A_275_49#
cc_1 VNB N_A_86_23#_M1003_g 0.00770473f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.465
cc_2 VNB N_A_86_23#_c_57_n 0.00308053f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.36
cc_3 VNB N_A_86_23#_c_58_n 0.0395191f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.36
cc_4 VNB N_A_86_23#_c_59_n 0.0300449f $X=-0.19 $Y=-0.245 $X2=2.955 $Y2=0.42
cc_5 VNB N_A_86_23#_c_60_n 0.0266612f $X=-0.19 $Y=-0.245 $X2=3.185 $Y2=1.93
cc_6 VNB N_A_86_23#_c_61_n 0.0162378f $X=-0.19 $Y=-0.245 $X2=3.05 $Y2=1.105
cc_7 VNB N_A_86_23#_c_62_n 0.0217126f $X=-0.19 $Y=-0.245 $X2=0.617 $Y2=1.195
cc_8 VNB N_A1_M1007_g 0.00628176f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB A1 0.00271182f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=0.665
cc_10 VNB N_A1_c_127_n 0.0345992f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A1_c_128_n 0.0199915f $X=-0.19 $Y=-0.245 $X2=0.68 $Y2=1.36
cc_12 VNB N_A2_M1000_g 0.0258094f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A2_c_162_n 0.02377f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.465
cc_14 VNB N_A2_c_163_n 0.00365498f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A3_M1004_g 0.0254494f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.195
cc_16 VNB N_A3_c_200_n 0.0239519f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.465
cc_17 VNB N_A3_c_201_n 0.00396526f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_B1_M1008_g 0.0285741f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_B1_c_236_n 0.0260747f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.465
cc_20 VNB N_B1_c_237_n 0.0031748f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_X_c_267_n 0.0644279f $X=-0.19 $Y=-0.245 $X2=2.455 $Y2=2.485
cc_22 VNB N_VPWR_c_277_n 0.143779f $X=-0.19 $Y=-0.245 $X2=2.455 $Y2=2.015
cc_23 VNB N_VGND_c_319_n 0.00231017f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=0.665
cc_24 VNB N_VGND_c_320_n 0.00527679f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_321_n 0.0160201f $X=-0.19 $Y=-0.245 $X2=0.64 $Y2=1.36
cc_26 VNB N_VGND_c_322_n 0.0162765f $X=-0.19 $Y=-0.245 $X2=2.455 $Y2=2.485
cc_27 VNB N_VGND_c_323_n 0.032059f $X=-0.19 $Y=-0.245 $X2=2.955 $Y2=0.42
cc_28 VNB N_VGND_c_324_n 0.189321f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_325_n 0.0110935f $X=-0.19 $Y=-0.245 $X2=2.455 $Y2=2.015
cc_30 VNB N_VGND_c_326_n 0.00634081f $X=-0.19 $Y=-0.245 $X2=0.617 $Y2=1.36
cc_31 VNB N_A_275_49#_c_362_n 0.0125542f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.465
cc_32 VNB N_A_275_49#_c_363_n 0.00432564f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.465
cc_33 VPB N_A_86_23#_M1003_g 0.0251635f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=2.465
cc_34 VPB N_A_86_23#_c_57_n 0.00197515f $X=-0.19 $Y=1.655 $X2=0.64 $Y2=1.36
cc_35 VPB N_A_86_23#_c_65_n 0.0152801f $X=-0.19 $Y=1.655 $X2=3.095 $Y2=2.015
cc_36 VPB N_A_86_23#_c_60_n 0.0136606f $X=-0.19 $Y=1.655 $X2=3.185 $Y2=1.93
cc_37 VPB N_A1_M1007_g 0.0229955f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_38 VPB A1 0.0025755f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=0.665
cc_39 VPB N_A2_M1009_g 0.0193303f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=1.195
cc_40 VPB N_A2_c_162_n 0.00613609f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=2.465
cc_41 VPB N_A2_c_163_n 0.00240649f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_42 VPB N_A3_M1001_g 0.0196534f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_43 VPB N_A3_c_200_n 0.00615025f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=2.465
cc_44 VPB N_A3_c_201_n 0.00321714f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_45 VPB N_B1_M1006_g 0.0229308f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=1.195
cc_46 VPB N_B1_c_236_n 0.00630358f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=2.465
cc_47 VPB N_B1_c_237_n 0.00350186f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_48 VPB N_X_c_267_n 0.0594775f $X=-0.19 $Y=1.655 $X2=2.455 $Y2=2.485
cc_49 VPB N_VPWR_c_278_n 0.0020627f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=0.665
cc_50 VPB N_VPWR_c_279_n 0.014965f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=2.465
cc_51 VPB N_VPWR_c_280_n 0.034895f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_52 VPB N_VPWR_c_281_n 0.0159542f $X=-0.19 $Y=1.655 $X2=0.64 $Y2=1.36
cc_53 VPB N_VPWR_c_282_n 0.0437629f $X=-0.19 $Y=1.655 $X2=2.455 $Y2=2.485
cc_54 VPB N_VPWR_c_283_n 0.0109159f $X=-0.19 $Y=1.655 $X2=3.05 $Y2=0.42
cc_55 VPB N_VPWR_c_277_n 0.050049f $X=-0.19 $Y=1.655 $X2=2.455 $Y2=2.015
cc_56 N_A_86_23#_M1003_g N_A1_M1007_g 0.0118392f $X=0.505 $Y=2.465 $X2=0 $Y2=0
cc_57 N_A_86_23#_c_57_n N_A1_M1007_g 0.00391153f $X=0.64 $Y=1.36 $X2=0 $Y2=0
cc_58 N_A_86_23#_c_69_p N_A1_M1007_g 0.0186005f $X=2.29 $Y=2.015 $X2=0 $Y2=0
cc_59 N_A_86_23#_M1003_g A1 5.92362e-19 $X=0.505 $Y=2.465 $X2=0 $Y2=0
cc_60 N_A_86_23#_c_57_n A1 0.0325977f $X=0.64 $Y=1.36 $X2=0 $Y2=0
cc_61 N_A_86_23#_c_58_n A1 0.00116942f $X=0.64 $Y=1.36 $X2=0 $Y2=0
cc_62 N_A_86_23#_c_69_p A1 0.0173766f $X=2.29 $Y=2.015 $X2=0 $Y2=0
cc_63 N_A_86_23#_M1003_g N_A1_c_127_n 3.11697e-19 $X=0.505 $Y=2.465 $X2=0 $Y2=0
cc_64 N_A_86_23#_c_57_n N_A1_c_127_n 0.00127241f $X=0.64 $Y=1.36 $X2=0 $Y2=0
cc_65 N_A_86_23#_c_58_n N_A1_c_127_n 0.0173859f $X=0.64 $Y=1.36 $X2=0 $Y2=0
cc_66 N_A_86_23#_c_69_p N_A1_c_127_n 7.2381e-19 $X=2.29 $Y=2.015 $X2=0 $Y2=0
cc_67 N_A_86_23#_c_58_n N_A1_c_128_n 4.65474e-19 $X=0.64 $Y=1.36 $X2=0 $Y2=0
cc_68 N_A_86_23#_c_62_n N_A1_c_128_n 0.00594269f $X=0.617 $Y=1.195 $X2=0 $Y2=0
cc_69 N_A_86_23#_c_69_p N_A2_M1009_g 0.0151461f $X=2.29 $Y=2.015 $X2=0 $Y2=0
cc_70 N_A_86_23#_c_69_p N_A2_c_162_n 0.00229911f $X=2.29 $Y=2.015 $X2=0 $Y2=0
cc_71 N_A_86_23#_c_69_p N_A2_c_163_n 0.0234981f $X=2.29 $Y=2.015 $X2=0 $Y2=0
cc_72 N_A_86_23#_c_69_p N_A3_M1001_g 0.0129992f $X=2.29 $Y=2.015 $X2=0 $Y2=0
cc_73 N_A_86_23#_c_84_p N_A3_c_200_n 0.00374626f $X=2.455 $Y=2.015 $X2=0 $Y2=0
cc_74 N_A_86_23#_c_69_p N_A3_c_201_n 0.0190005f $X=2.29 $Y=2.015 $X2=0 $Y2=0
cc_75 N_A_86_23#_c_84_p N_A3_c_201_n 0.00554706f $X=2.455 $Y=2.015 $X2=0 $Y2=0
cc_76 N_A_86_23#_c_60_n N_B1_M1008_g 0.00653474f $X=3.185 $Y=1.93 $X2=0 $Y2=0
cc_77 N_A_86_23#_c_61_n N_B1_M1008_g 0.00309198f $X=3.05 $Y=1.105 $X2=0 $Y2=0
cc_78 N_A_86_23#_c_65_n N_B1_M1006_g 0.0165738f $X=3.095 $Y=2.015 $X2=0 $Y2=0
cc_79 N_A_86_23#_c_60_n N_B1_M1006_g 0.00567484f $X=3.185 $Y=1.93 $X2=0 $Y2=0
cc_80 N_A_86_23#_c_65_n N_B1_c_236_n 0.00291568f $X=3.095 $Y=2.015 $X2=0 $Y2=0
cc_81 N_A_86_23#_c_60_n N_B1_c_236_n 0.00805981f $X=3.185 $Y=1.93 $X2=0 $Y2=0
cc_82 N_A_86_23#_c_61_n N_B1_c_236_n 0.00510637f $X=3.05 $Y=1.105 $X2=0 $Y2=0
cc_83 N_A_86_23#_c_65_n N_B1_c_237_n 0.0195184f $X=3.095 $Y=2.015 $X2=0 $Y2=0
cc_84 N_A_86_23#_c_60_n N_B1_c_237_n 0.0319519f $X=3.185 $Y=1.93 $X2=0 $Y2=0
cc_85 N_A_86_23#_c_84_p N_B1_c_237_n 0.00519213f $X=2.455 $Y=2.015 $X2=0 $Y2=0
cc_86 N_A_86_23#_c_61_n N_B1_c_237_n 0.00655466f $X=3.05 $Y=1.105 $X2=0 $Y2=0
cc_87 N_A_86_23#_c_57_n N_X_c_267_n 0.0525633f $X=0.64 $Y=1.36 $X2=0 $Y2=0
cc_88 N_A_86_23#_c_62_n N_X_c_267_n 0.0259311f $X=0.617 $Y=1.195 $X2=0 $Y2=0
cc_89 N_A_86_23#_c_57_n N_VPWR_M1003_d 0.00164112f $X=0.64 $Y=1.36 $X2=-0.19
+ $Y2=-0.245
cc_90 N_A_86_23#_c_69_p N_VPWR_M1003_d 0.0160602f $X=2.29 $Y=2.015 $X2=-0.19
+ $Y2=-0.245
cc_91 N_A_86_23#_c_102_p N_VPWR_M1003_d 0.00227149f $X=0.805 $Y=2.015 $X2=-0.19
+ $Y2=-0.245
cc_92 N_A_86_23#_c_65_n N_VPWR_M1006_d 0.00756851f $X=3.095 $Y=2.015 $X2=0 $Y2=0
cc_93 N_A_86_23#_M1003_g N_VPWR_c_278_n 0.0195205f $X=0.505 $Y=2.465 $X2=0 $Y2=0
cc_94 N_A_86_23#_c_69_p N_VPWR_c_278_n 0.0312828f $X=2.29 $Y=2.015 $X2=0 $Y2=0
cc_95 N_A_86_23#_c_102_p N_VPWR_c_278_n 0.0170914f $X=0.805 $Y=2.015 $X2=0 $Y2=0
cc_96 N_A_86_23#_c_65_n N_VPWR_c_280_n 0.0221397f $X=3.095 $Y=2.015 $X2=0 $Y2=0
cc_97 N_A_86_23#_M1003_g N_VPWR_c_281_n 0.00486043f $X=0.505 $Y=2.465 $X2=0
+ $Y2=0
cc_98 N_A_86_23#_c_109_p N_VPWR_c_282_n 0.0212513f $X=2.455 $Y=2.485 $X2=0 $Y2=0
cc_99 N_A_86_23#_M1001_d N_VPWR_c_277_n 0.00526034f $X=2.275 $Y=1.835 $X2=0
+ $Y2=0
cc_100 N_A_86_23#_M1003_g N_VPWR_c_277_n 0.00920706f $X=0.505 $Y=2.465 $X2=0
+ $Y2=0
cc_101 N_A_86_23#_c_109_p N_VPWR_c_277_n 0.0127519f $X=2.455 $Y=2.485 $X2=0
+ $Y2=0
cc_102 N_A_86_23#_c_69_p A_275_367# 0.0113748f $X=2.29 $Y=2.015 $X2=-0.19
+ $Y2=-0.245
cc_103 N_A_86_23#_c_69_p A_367_367# 0.0111311f $X=2.29 $Y=2.015 $X2=-0.19
+ $Y2=-0.245
cc_104 N_A_86_23#_c_57_n N_VGND_c_319_n 0.0189984f $X=0.64 $Y=1.36 $X2=0 $Y2=0
cc_105 N_A_86_23#_c_58_n N_VGND_c_319_n 0.00160017f $X=0.64 $Y=1.36 $X2=0 $Y2=0
cc_106 N_A_86_23#_c_62_n N_VGND_c_319_n 0.0180351f $X=0.617 $Y=1.195 $X2=0 $Y2=0
cc_107 N_A_86_23#_c_62_n N_VGND_c_321_n 0.00477554f $X=0.617 $Y=1.195 $X2=0
+ $Y2=0
cc_108 N_A_86_23#_c_59_n N_VGND_c_323_n 0.0301644f $X=2.955 $Y=0.42 $X2=0 $Y2=0
cc_109 N_A_86_23#_M1008_d N_VGND_c_324_n 0.00247088f $X=2.815 $Y=0.245 $X2=0
+ $Y2=0
cc_110 N_A_86_23#_c_59_n N_VGND_c_324_n 0.0174172f $X=2.955 $Y=0.42 $X2=0 $Y2=0
cc_111 N_A_86_23#_c_62_n N_VGND_c_324_n 0.00921794f $X=0.617 $Y=1.195 $X2=0
+ $Y2=0
cc_112 N_A_86_23#_c_60_n N_A_275_49#_c_362_n 0.00303221f $X=3.185 $Y=1.93 $X2=0
+ $Y2=0
cc_113 N_A_86_23#_c_61_n N_A_275_49#_c_362_n 0.00171763f $X=3.05 $Y=1.105 $X2=0
+ $Y2=0
cc_114 A1 N_A2_M1000_g 6.9501e-19 $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_115 N_A1_c_128_n N_A2_M1000_g 0.0214229f $X=1.205 $Y=1.21 $X2=0 $Y2=0
cc_116 N_A1_M1007_g N_A2_M1009_g 0.0652339f $X=1.3 $Y=2.465 $X2=0 $Y2=0
cc_117 A1 N_A2_c_162_n 3.1061e-19 $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_118 N_A1_c_127_n N_A2_c_162_n 0.0200527f $X=1.2 $Y=1.375 $X2=0 $Y2=0
cc_119 A1 N_A2_c_163_n 0.0266906f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_120 N_A1_c_127_n N_A2_c_163_n 0.00291121f $X=1.2 $Y=1.375 $X2=0 $Y2=0
cc_121 N_A1_M1007_g N_VPWR_c_278_n 0.0269504f $X=1.3 $Y=2.465 $X2=0 $Y2=0
cc_122 N_A1_M1007_g N_VPWR_c_282_n 0.00486043f $X=1.3 $Y=2.465 $X2=0 $Y2=0
cc_123 N_A1_M1007_g N_VPWR_c_277_n 0.00845871f $X=1.3 $Y=2.465 $X2=0 $Y2=0
cc_124 A1 N_VGND_c_319_n 0.0146319f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_125 N_A1_c_127_n N_VGND_c_319_n 0.00129819f $X=1.2 $Y=1.375 $X2=0 $Y2=0
cc_126 N_A1_c_128_n N_VGND_c_319_n 0.0170765f $X=1.205 $Y=1.21 $X2=0 $Y2=0
cc_127 N_A1_c_128_n N_VGND_c_322_n 0.00477554f $X=1.205 $Y=1.21 $X2=0 $Y2=0
cc_128 N_A1_c_128_n N_VGND_c_324_n 0.00834285f $X=1.205 $Y=1.21 $X2=0 $Y2=0
cc_129 N_A1_c_128_n N_A_275_49#_c_366_n 0.00310763f $X=1.205 $Y=1.21 $X2=0 $Y2=0
cc_130 N_A1_c_128_n N_A_275_49#_c_363_n 0.00447809f $X=1.205 $Y=1.21 $X2=0 $Y2=0
cc_131 N_A2_M1009_g N_A3_M1001_g 0.0694856f $X=1.76 $Y=2.465 $X2=0 $Y2=0
cc_132 N_A2_M1000_g N_A3_M1004_g 0.0313619f $X=1.755 $Y=0.665 $X2=0 $Y2=0
cc_133 N_A2_c_162_n N_A3_c_200_n 0.0204266f $X=1.75 $Y=1.51 $X2=0 $Y2=0
cc_134 N_A2_c_163_n N_A3_c_200_n 3.76435e-19 $X=1.75 $Y=1.51 $X2=0 $Y2=0
cc_135 N_A2_M1009_g N_A3_c_201_n 5.12465e-19 $X=1.76 $Y=2.465 $X2=0 $Y2=0
cc_136 N_A2_c_162_n N_A3_c_201_n 0.00221329f $X=1.75 $Y=1.51 $X2=0 $Y2=0
cc_137 N_A2_c_163_n N_A3_c_201_n 0.0331397f $X=1.75 $Y=1.51 $X2=0 $Y2=0
cc_138 N_A2_M1009_g N_VPWR_c_278_n 0.00498086f $X=1.76 $Y=2.465 $X2=0 $Y2=0
cc_139 N_A2_M1009_g N_VPWR_c_282_n 0.00585385f $X=1.76 $Y=2.465 $X2=0 $Y2=0
cc_140 N_A2_M1009_g N_VPWR_c_277_n 0.0111377f $X=1.76 $Y=2.465 $X2=0 $Y2=0
cc_141 N_A2_M1000_g N_VGND_c_319_n 7.67654e-19 $X=1.755 $Y=0.665 $X2=0 $Y2=0
cc_142 N_A2_M1000_g N_VGND_c_320_n 0.00521996f $X=1.755 $Y=0.665 $X2=0 $Y2=0
cc_143 N_A2_M1000_g N_VGND_c_322_n 0.0054677f $X=1.755 $Y=0.665 $X2=0 $Y2=0
cc_144 N_A2_M1000_g N_VGND_c_324_n 0.0103781f $X=1.755 $Y=0.665 $X2=0 $Y2=0
cc_145 N_A2_M1000_g N_A_275_49#_c_366_n 0.0105566f $X=1.755 $Y=0.665 $X2=0 $Y2=0
cc_146 N_A2_M1000_g N_A_275_49#_c_362_n 0.0120988f $X=1.755 $Y=0.665 $X2=0 $Y2=0
cc_147 N_A2_c_162_n N_A_275_49#_c_362_n 0.00304681f $X=1.75 $Y=1.51 $X2=0 $Y2=0
cc_148 N_A2_c_163_n N_A_275_49#_c_362_n 0.00977984f $X=1.75 $Y=1.51 $X2=0 $Y2=0
cc_149 N_A2_M1000_g N_A_275_49#_c_363_n 0.00146026f $X=1.755 $Y=0.665 $X2=0
+ $Y2=0
cc_150 N_A2_c_162_n N_A_275_49#_c_363_n 7.519e-19 $X=1.75 $Y=1.51 $X2=0 $Y2=0
cc_151 N_A2_c_163_n N_A_275_49#_c_363_n 0.0173993f $X=1.75 $Y=1.51 $X2=0 $Y2=0
cc_152 N_A2_M1000_g N_A_275_49#_c_375_n 6.4041e-19 $X=1.755 $Y=0.665 $X2=0 $Y2=0
cc_153 N_A3_M1004_g N_B1_M1008_g 0.0239076f $X=2.31 $Y=0.665 $X2=0 $Y2=0
cc_154 N_A3_M1001_g N_B1_M1006_g 0.0263515f $X=2.2 $Y=2.465 $X2=0 $Y2=0
cc_155 N_A3_c_201_n N_B1_M1006_g 2.53873e-19 $X=2.29 $Y=1.51 $X2=0 $Y2=0
cc_156 N_A3_c_200_n N_B1_c_236_n 0.0204543f $X=2.29 $Y=1.51 $X2=0 $Y2=0
cc_157 N_A3_c_201_n N_B1_c_236_n 2.93393e-19 $X=2.29 $Y=1.51 $X2=0 $Y2=0
cc_158 N_A3_M1001_g N_B1_c_237_n 2.60445e-19 $X=2.2 $Y=2.465 $X2=0 $Y2=0
cc_159 N_A3_c_200_n N_B1_c_237_n 0.00221553f $X=2.29 $Y=1.51 $X2=0 $Y2=0
cc_160 N_A3_c_201_n N_B1_c_237_n 0.0323586f $X=2.29 $Y=1.51 $X2=0 $Y2=0
cc_161 N_A3_M1001_g N_VPWR_c_280_n 0.00110954f $X=2.2 $Y=2.465 $X2=0 $Y2=0
cc_162 N_A3_M1001_g N_VPWR_c_282_n 0.00585385f $X=2.2 $Y=2.465 $X2=0 $Y2=0
cc_163 N_A3_M1001_g N_VPWR_c_277_n 0.0111937f $X=2.2 $Y=2.465 $X2=0 $Y2=0
cc_164 N_A3_M1004_g N_VGND_c_320_n 0.00666369f $X=2.31 $Y=0.665 $X2=0 $Y2=0
cc_165 N_A3_M1004_g N_VGND_c_323_n 0.00554241f $X=2.31 $Y=0.665 $X2=0 $Y2=0
cc_166 N_A3_M1004_g N_VGND_c_324_n 0.0104903f $X=2.31 $Y=0.665 $X2=0 $Y2=0
cc_167 N_A3_M1004_g N_A_275_49#_c_366_n 6.47401e-19 $X=2.31 $Y=0.665 $X2=0 $Y2=0
cc_168 N_A3_M1004_g N_A_275_49#_c_362_n 0.0141182f $X=2.31 $Y=0.665 $X2=0 $Y2=0
cc_169 N_A3_c_200_n N_A_275_49#_c_362_n 0.00387598f $X=2.29 $Y=1.51 $X2=0 $Y2=0
cc_170 N_A3_c_201_n N_A_275_49#_c_362_n 0.0279468f $X=2.29 $Y=1.51 $X2=0 $Y2=0
cc_171 N_A3_M1004_g N_A_275_49#_c_375_n 0.0102914f $X=2.31 $Y=0.665 $X2=0 $Y2=0
cc_172 N_B1_M1006_g N_VPWR_c_280_n 0.0184095f $X=2.74 $Y=2.465 $X2=0 $Y2=0
cc_173 N_B1_M1006_g N_VPWR_c_282_n 0.00486043f $X=2.74 $Y=2.465 $X2=0 $Y2=0
cc_174 N_B1_M1006_g N_VPWR_c_277_n 0.00864313f $X=2.74 $Y=2.465 $X2=0 $Y2=0
cc_175 N_B1_M1008_g N_VGND_c_323_n 0.00575161f $X=2.74 $Y=0.665 $X2=0 $Y2=0
cc_176 N_B1_M1008_g N_VGND_c_324_n 0.0118478f $X=2.74 $Y=0.665 $X2=0 $Y2=0
cc_177 N_B1_M1008_g N_A_275_49#_c_362_n 0.00117868f $X=2.74 $Y=0.665 $X2=0 $Y2=0
cc_178 N_B1_c_237_n N_A_275_49#_c_362_n 0.00899355f $X=2.83 $Y=1.51 $X2=0 $Y2=0
cc_179 N_X_c_267_n N_VPWR_c_281_n 0.0206786f $X=0.29 $Y=0.42 $X2=0 $Y2=0
cc_180 N_X_M1003_s N_VPWR_c_277_n 0.00371702f $X=0.165 $Y=1.835 $X2=0 $Y2=0
cc_181 N_X_c_267_n N_VPWR_c_277_n 0.0115856f $X=0.29 $Y=0.42 $X2=0 $Y2=0
cc_182 N_X_c_267_n N_VGND_c_321_n 0.0206786f $X=0.29 $Y=0.42 $X2=0 $Y2=0
cc_183 N_X_M1005_s N_VGND_c_324_n 0.00368844f $X=0.165 $Y=0.245 $X2=0 $Y2=0
cc_184 N_X_c_267_n N_VGND_c_324_n 0.0115856f $X=0.29 $Y=0.42 $X2=0 $Y2=0
cc_185 N_VPWR_c_277_n A_275_367# 0.0132771f $X=3.12 $Y=3.33 $X2=-0.19 $Y2=-0.245
cc_186 N_VPWR_c_277_n A_367_367# 0.0124205f $X=3.12 $Y=3.33 $X2=-0.19 $Y2=-0.245
cc_187 N_VGND_c_324_n N_A_275_49#_M1002_d 0.00521963f $X=3.12 $Y=0 $X2=-0.19
+ $Y2=-0.245
cc_188 N_VGND_c_324_n N_A_275_49#_M1004_d 0.00258346f $X=3.12 $Y=0 $X2=0 $Y2=0
cc_189 N_VGND_c_319_n N_A_275_49#_c_366_n 0.0521562f $X=1.085 $Y=0.39 $X2=0
+ $Y2=0
cc_190 N_VGND_c_322_n N_A_275_49#_c_366_n 0.0150272f $X=1.87 $Y=0 $X2=0 $Y2=0
cc_191 N_VGND_c_324_n N_A_275_49#_c_366_n 0.00928716f $X=3.12 $Y=0 $X2=0 $Y2=0
cc_192 N_VGND_M1000_d N_A_275_49#_c_362_n 0.00329016f $X=1.83 $Y=0.245 $X2=0
+ $Y2=0
cc_193 N_VGND_c_320_n N_A_275_49#_c_362_n 0.0236753f $X=2.035 $Y=0.37 $X2=0
+ $Y2=0
cc_194 N_VGND_c_319_n N_A_275_49#_c_363_n 0.00150747f $X=1.085 $Y=0.39 $X2=0
+ $Y2=0
cc_195 N_VGND_c_323_n N_A_275_49#_c_375_n 0.0162482f $X=3.12 $Y=0 $X2=0 $Y2=0
cc_196 N_VGND_c_324_n N_A_275_49#_c_375_n 0.0108651f $X=3.12 $Y=0 $X2=0 $Y2=0
