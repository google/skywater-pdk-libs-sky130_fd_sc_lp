* File: sky130_fd_sc_lp__or3b_1.pex.spice
* Created: Fri Aug 28 11:23:55 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__OR3B_1%C_N 2 5 8 10 11 12 13 14 15 22 24
r25 22 24 45.5639 $w=3.95e-07 $l=1.65e-07 $layer=POLY_cond $X=0.352 $Y=1.045
+ $X2=0.352 $Y2=0.88
r26 22 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.32
+ $Y=1.045 $X2=0.32 $Y2=1.045
r27 14 15 13.3251 $w=3.18e-07 $l=3.7e-07 $layer=LI1_cond $X=0.245 $Y=2.035
+ $X2=0.245 $Y2=2.405
r28 13 14 13.3251 $w=3.18e-07 $l=3.7e-07 $layer=LI1_cond $X=0.245 $Y=1.665
+ $X2=0.245 $Y2=2.035
r29 12 13 13.3251 $w=3.18e-07 $l=3.7e-07 $layer=LI1_cond $X=0.245 $Y=1.295
+ $X2=0.245 $Y2=1.665
r30 12 23 9.00346 $w=3.18e-07 $l=2.5e-07 $layer=LI1_cond $X=0.245 $Y=1.295
+ $X2=0.245 $Y2=1.045
r31 11 23 4.32166 $w=3.18e-07 $l=1.2e-07 $layer=LI1_cond $X=0.245 $Y=0.925
+ $X2=0.245 $Y2=1.045
r32 8 10 625.574 $w=1.5e-07 $l=1.22e-06 $layer=POLY_cond $X=0.475 $Y=2.77
+ $X2=0.475 $Y2=1.55
r33 5 24 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.475 $Y=0.56
+ $X2=0.475 $Y2=0.88
r34 2 10 50.0695 $w=3.95e-07 $l=1.97e-07 $layer=POLY_cond $X=0.352 $Y=1.353
+ $X2=0.352 $Y2=1.55
r35 1 22 4.50555 $w=3.95e-07 $l=3.2e-08 $layer=POLY_cond $X=0.352 $Y=1.077
+ $X2=0.352 $Y2=1.045
r36 1 2 38.8604 $w=3.95e-07 $l=2.76e-07 $layer=POLY_cond $X=0.352 $Y=1.077
+ $X2=0.352 $Y2=1.353
.ends

.subckt PM_SKY130_FD_SC_LP__OR3B_1%A_110_70# 1 2 9 13 17 21 24 25
r44 25 30 75.2115 $w=7.25e-07 $l=5.05e-07 $layer=POLY_cond $X=1.152 $Y=1.165
+ $X2=1.152 $Y2=1.67
r45 25 29 51.0986 $w=7.25e-07 $l=1.65e-07 $layer=POLY_cond $X=1.152 $Y=1.165
+ $X2=1.152 $Y2=1
r46 24 27 15.4537 $w=4.53e-07 $l=5.05e-07 $layer=LI1_cond $X=0.822 $Y=1.165
+ $X2=0.822 $Y2=1.67
r47 24 26 6.51597 $w=4.53e-07 $l=1.65e-07 $layer=LI1_cond $X=0.822 $Y=1.165
+ $X2=0.822 $Y2=1
r48 24 25 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.955
+ $Y=1.165 $X2=0.955 $Y2=1.165
r49 21 27 48.7572 $w=2.58e-07 $l=1.1e-06 $layer=LI1_cond $X=0.725 $Y=2.77
+ $X2=0.725 $Y2=1.67
r50 17 26 19.5029 $w=2.58e-07 $l=4.4e-07 $layer=LI1_cond $X=0.725 $Y=0.56
+ $X2=0.725 $Y2=1
r51 13 30 192.287 $w=1.5e-07 $l=3.75e-07 $layer=POLY_cond $X=1.44 $Y=2.045
+ $X2=1.44 $Y2=1.67
r52 9 29 215.362 $w=1.5e-07 $l=4.2e-07 $layer=POLY_cond $X=1.44 $Y=0.58 $X2=1.44
+ $Y2=1
r53 2 21 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=2.56 $X2=0.69 $Y2=2.77
r54 1 17 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.35 $X2=0.69 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_LP__OR3B_1%B 3 7 9 10 11 12 13 14 15 21
c45 9 0 4.27728e-20 $X=1.89 $Y=0.9
r46 21 22 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.89
+ $Y=1.065 $X2=1.89 $Y2=1.065
r47 14 15 10.2748 $w=4.13e-07 $l=3.7e-07 $layer=LI1_cond $X=1.767 $Y=1.665
+ $X2=1.767 $Y2=2.035
r48 13 14 10.2748 $w=4.13e-07 $l=3.7e-07 $layer=LI1_cond $X=1.767 $Y=1.295
+ $X2=1.767 $Y2=1.665
r49 13 22 6.38703 $w=4.13e-07 $l=2.3e-07 $layer=LI1_cond $X=1.767 $Y=1.295
+ $X2=1.767 $Y2=1.065
r50 12 22 3.88776 $w=4.13e-07 $l=1.4e-07 $layer=LI1_cond $X=1.767 $Y=0.925
+ $X2=1.767 $Y2=1.065
r51 10 21 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.89 $Y=1.405
+ $X2=1.89 $Y2=1.065
r52 10 11 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.89 $Y=1.405
+ $X2=1.89 $Y2=1.57
r53 9 21 38.6168 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.89 $Y=0.9 $X2=1.89
+ $Y2=1.065
r54 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.91 $Y=0.58 $X2=1.91
+ $Y2=0.9
r55 3 11 243.564 $w=1.5e-07 $l=4.75e-07 $layer=POLY_cond $X=1.8 $Y=2.045 $X2=1.8
+ $Y2=1.57
.ends

.subckt PM_SKY130_FD_SC_LP__OR3B_1%A 3 6 7 8 15
r31 12 15 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=2.16 $Y=2.855
+ $X2=2.34 $Y2=2.855
r32 8 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.16
+ $Y=2.855 $X2=2.16 $Y2=2.855
r33 7 8 14.5572 $w=3.78e-07 $l=4.8e-07 $layer=LI1_cond $X=1.68 $Y=2.83 $X2=2.16
+ $Y2=2.83
r34 3 6 751.202 $w=1.5e-07 $l=1.465e-06 $layer=POLY_cond $X=2.34 $Y=0.58
+ $X2=2.34 $Y2=2.045
r35 1 15 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.34 $Y=2.69
+ $X2=2.34 $Y2=2.855
r36 1 6 330.734 $w=1.5e-07 $l=6.45e-07 $layer=POLY_cond $X=2.34 $Y=2.69 $X2=2.34
+ $Y2=2.045
.ends

.subckt PM_SKY130_FD_SC_LP__OR3B_1%A_220_74# 1 2 3 12 15 18 20 23 24 26 28 31 32
+ 35 38 42 44 46
c88 38 0 4.27728e-20 $X=1.225 $Y=1.88
c89 28 0 1.33431e-19 $X=2.24 $Y=2.3
c90 15 0 6.36774e-20 $X=2.865 $Y=2.465
r91 40 42 4.73325 $w=2.78e-07 $l=1.15e-07 $layer=LI1_cond $X=2.125 $Y=0.53
+ $X2=2.24 $Y2=0.53
r92 37 38 73.7219 $w=1.68e-07 $l=1.13e-06 $layer=LI1_cond $X=1.305 $Y=0.75
+ $X2=1.305 $Y2=1.88
r93 35 37 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=1.225 $Y=0.585
+ $X2=1.225 $Y2=0.75
r94 32 47 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.82 $Y=1.485
+ $X2=2.82 $Y2=1.65
r95 32 46 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.82 $Y=1.485
+ $X2=2.82 $Y2=1.32
r96 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.82
+ $Y=1.485 $X2=2.82 $Y2=1.485
r97 29 44 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.325 $Y=1.485
+ $X2=2.24 $Y2=1.485
r98 29 31 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=2.325 $Y=1.485
+ $X2=2.82 $Y2=1.485
r99 27 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.24 $Y=1.65
+ $X2=2.24 $Y2=1.485
r100 27 28 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=2.24 $Y=1.65
+ $X2=2.24 $Y2=2.3
r101 26 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.24 $Y=1.32
+ $X2=2.24 $Y2=1.485
r102 25 42 3.65648 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=2.24 $Y=0.67
+ $X2=2.24 $Y2=0.53
r103 25 26 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=2.24 $Y=0.67
+ $X2=2.24 $Y2=1.32
r104 23 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.155 $Y=2.385
+ $X2=2.24 $Y2=2.3
r105 23 24 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=2.155 $Y=2.385
+ $X2=1.39 $Y2=2.385
r106 20 38 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=1.225 $Y=2.045
+ $X2=1.225 $Y2=1.88
r107 18 24 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.225 $Y=2.3
+ $X2=1.39 $Y2=2.385
r108 18 20 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=1.225 $Y=2.3
+ $X2=1.225 $Y2=2.045
r109 15 47 417.904 $w=1.5e-07 $l=8.15e-07 $layer=POLY_cond $X=2.865 $Y=2.465
+ $X2=2.865 $Y2=1.65
r110 12 46 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.865 $Y=0.79
+ $X2=2.865 $Y2=1.32
r111 3 20 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=1.1
+ $Y=1.835 $X2=1.225 $Y2=2.045
r112 2 40 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=1.985
+ $Y=0.37 $X2=2.125 $Y2=0.555
r113 1 35 182 $w=1.7e-07 $l=2.7037e-07 $layer=licon1_NDIFF $count=1 $X=1.1
+ $Y=0.37 $X2=1.225 $Y2=0.585
.ends

.subckt PM_SKY130_FD_SC_LP__OR3B_1%VPWR 1 2 7 9 13 17 19 29 30 36
r34 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r35 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r36 30 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.64 $Y2=3.33
r37 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r38 27 36 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.755 $Y=3.33
+ $X2=2.625 $Y2=3.33
r39 27 29 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=2.755 $Y=3.33
+ $X2=3.12 $Y2=3.33
r40 26 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r41 25 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r42 23 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r43 22 25 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=0.72 $Y=3.33
+ $X2=2.16 $Y2=3.33
r44 22 23 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r45 20 33 4.78091 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=3.33
+ $X2=0.212 $Y2=3.33
r46 20 22 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.425 $Y=3.33
+ $X2=0.72 $Y2=3.33
r47 19 36 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.495 $Y=3.33
+ $X2=2.625 $Y2=3.33
r48 19 25 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=2.495 $Y=3.33
+ $X2=2.16 $Y2=3.33
r49 17 26 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r50 17 23 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.72 $Y2=3.33
r51 13 16 21.7191 $w=2.58e-07 $l=4.9e-07 $layer=LI1_cond $X=2.625 $Y=1.985
+ $X2=2.625 $Y2=2.475
r52 11 36 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=2.625 $Y=3.245
+ $X2=2.625 $Y2=3.33
r53 11 16 34.13 $w=2.58e-07 $l=7.7e-07 $layer=LI1_cond $X=2.625 $Y=3.245
+ $X2=2.625 $Y2=2.475
r54 7 33 2.98526 $w=3.3e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.26 $Y=3.245
+ $X2=0.212 $Y2=3.33
r55 7 9 16.5882 $w=3.28e-07 $l=4.75e-07 $layer=LI1_cond $X=0.26 $Y=3.245
+ $X2=0.26 $Y2=2.77
r56 2 16 300 $w=1.7e-07 $l=7.48331e-07 $layer=licon1_PDIFF $count=2 $X=2.415
+ $Y=1.835 $X2=2.65 $Y2=2.475
r57 2 13 600 $w=1.7e-07 $l=2.54165e-07 $layer=licon1_PDIFF $count=1 $X=2.415
+ $Y=1.835 $X2=2.605 $Y2=1.985
r58 1 9 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.56 $X2=0.26 $Y2=2.77
.ends

.subckt PM_SKY130_FD_SC_LP__OR3B_1%X 1 2 10 11 12 13 14 15 31 41
c20 13 0 1.33431e-19 $X=3.035 $Y=1.95
r21 28 31 1.02897 $w=2.78e-07 $l=2.5e-08 $layer=LI1_cond $X=3.115 $Y=1.955
+ $X2=3.115 $Y2=1.98
r22 15 38 5.55642 $w=2.78e-07 $l=1.35e-07 $layer=LI1_cond $X=3.115 $Y=2.775
+ $X2=3.115 $Y2=2.91
r23 14 15 15.2287 $w=2.78e-07 $l=3.7e-07 $layer=LI1_cond $X=3.115 $Y=2.405
+ $X2=3.115 $Y2=2.775
r24 13 28 0.123476 $w=2.78e-07 $l=3e-09 $layer=LI1_cond $X=3.115 $Y=1.952
+ $X2=3.115 $Y2=1.955
r25 13 41 7.40445 $w=2.78e-07 $l=1.37e-07 $layer=LI1_cond $X=3.115 $Y=1.952
+ $X2=3.115 $Y2=1.815
r26 13 14 15.1464 $w=2.78e-07 $l=3.68e-07 $layer=LI1_cond $X=3.115 $Y=2.037
+ $X2=3.115 $Y2=2.405
r27 13 31 2.34604 $w=2.78e-07 $l=5.7e-08 $layer=LI1_cond $X=3.115 $Y=2.037
+ $X2=3.115 $Y2=1.98
r28 11 12 16.8751 $w=2.78e-07 $l=4.1e-07 $layer=LI1_cond $X=3.115 $Y=0.515
+ $X2=3.115 $Y2=0.925
r29 10 41 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=3.17 $Y=1.16
+ $X2=3.17 $Y2=1.815
r30 9 12 3.91007 $w=2.78e-07 $l=9.5e-08 $layer=LI1_cond $X=3.115 $Y=1.02
+ $X2=3.115 $Y2=0.925
r31 9 10 7.52792 $w=2.78e-07 $l=1.4e-07 $layer=LI1_cond $X=3.115 $Y=1.02
+ $X2=3.115 $Y2=1.16
r32 2 38 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=2.94
+ $Y=1.835 $X2=3.08 $Y2=2.91
r33 2 31 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.94
+ $Y=1.835 $X2=3.08 $Y2=1.98
r34 1 11 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.94
+ $Y=0.37 $X2=3.08 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LP__OR3B_1%VGND 1 2 3 10 12 16 20 24 26 31 38 39 45 48
r44 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r45 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r46 39 49 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.64
+ $Y2=0
r47 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r48 36 48 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.755 $Y=0 $X2=2.625
+ $Y2=0
r49 36 38 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=2.755 $Y=0 $X2=3.12
+ $Y2=0
r50 35 49 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r51 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r52 32 45 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=1.79 $Y=0 $X2=1.675
+ $Y2=0
r53 32 34 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=1.79 $Y=0 $X2=2.16
+ $Y2=0
r54 31 48 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.495 $Y=0 $X2=2.625
+ $Y2=0
r55 31 34 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=2.495 $Y=0 $X2=2.16
+ $Y2=0
r56 30 43 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.24
+ $Y2=0
r57 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r58 27 42 4.78091 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=0 $X2=0.212
+ $Y2=0
r59 27 29 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=0.425 $Y=0 $X2=1.2
+ $Y2=0
r60 26 45 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=1.56 $Y=0 $X2=1.675
+ $Y2=0
r61 26 29 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=1.56 $Y=0 $X2=1.2
+ $Y2=0
r62 24 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r63 24 30 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r64 24 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r65 20 22 20.8326 $w=2.58e-07 $l=4.7e-07 $layer=LI1_cond $X=2.625 $Y=0.515
+ $X2=2.625 $Y2=0.985
r66 18 48 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=2.625 $Y=0.085
+ $X2=2.625 $Y2=0
r67 18 20 19.0596 $w=2.58e-07 $l=4.3e-07 $layer=LI1_cond $X=2.625 $Y=0.085
+ $X2=2.625 $Y2=0.515
r68 14 45 0.280307 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.675 $Y=0.085
+ $X2=1.675 $Y2=0
r69 14 16 21.0446 $w=2.28e-07 $l=4.2e-07 $layer=LI1_cond $X=1.675 $Y=0.085
+ $X2=1.675 $Y2=0.505
r70 10 42 2.98526 $w=3.3e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.212 $Y2=0
r71 10 12 16.5882 $w=3.28e-07 $l=4.75e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.26 $Y2=0.56
r72 3 22 182 $w=1.7e-07 $l=7.23015e-07 $layer=licon1_NDIFF $count=1 $X=2.415
+ $Y=0.37 $X2=2.65 $Y2=0.985
r73 3 20 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=2.415
+ $Y=0.37 $X2=2.6 $Y2=0.515
r74 2 16 182 $w=1.7e-07 $l=2.17256e-07 $layer=licon1_NDIFF $count=1 $X=1.515
+ $Y=0.37 $X2=1.675 $Y2=0.505
r75 1 12 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.35 $X2=0.26 $Y2=0.56
.ends

