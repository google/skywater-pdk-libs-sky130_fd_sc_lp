* File: sky130_fd_sc_lp__srsdfstp_1.spice
* Created: Fri Aug 28 11:34:09 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__srsdfstp_1.pex.spice"
.subckt sky130_fd_sc_lp__srsdfstp_1  VNB VPB SCD D SCE SET_B CLK SLEEP_B VPWR
+ KAPWR Q VGND
* 
* VGND	VGND
* Q	Q
* KAPWR	KAPWR
* VPWR	VPWR
* SLEEP_B	SLEEP_B
* CLK	CLK
* SET_B	SET_B
* SCE	SCE
* D	D
* SCD	SCD
* VPB	VPB
* VNB	VNB
MM1001 A_111_119# N_SCD_M1001_g N_VGND_M1001_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.1134 PD=0.66 PS=1.38 NRD=18.564 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.5 A=0.063 P=1.14 MULT=1
MM1013 N_A_189_119#_M1013_d N_SCE_M1013_g A_111_119# VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0504 PD=0.7 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75000.6
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1016 A_275_119# N_D_M1016_g N_A_189_119#_M1013_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0672 AS=0.0588 PD=0.74 PS=0.7 NRD=30 NRS=0 M=1 R=2.8 SA=75001 SB=75000.7
+ A=0.063 P=1.14 MULT=1
MM1023 N_VGND_M1023_d N_A_339_93#_M1023_g A_275_119# VNB NSHORT L=0.15 W=0.42
+ AD=0.1365 AS=0.0672 PD=1.49 PS=0.74 NRD=11.424 NRS=30 M=1 R=2.8 SA=75001.5
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1029 N_VGND_M1029_d N_SCE_M1029_g N_A_339_93#_M1029_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0735 AS=0.1197 PD=0.77 PS=1.41 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1028 N_A_689_139#_M1028_d N_A_659_113#_M1028_g N_VGND_M1029_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.1197 AS=0.0735 PD=1.41 PS=0.77 NRD=0 NRS=19.992 M=1 R=2.8
+ SA=75000.7 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1047 N_A_887_139#_M1047_d N_A_659_113#_M1047_g N_A_189_119#_M1047_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.113475 AS=0.1197 PD=1.145 PS=1.41 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.3 A=0.063 P=1.14 MULT=1
MM1031 A_996_73# N_A_689_139#_M1031_g N_A_887_139#_M1047_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0847 AS=0.113475 PD=0.91 PS=1.145 NRD=41.904 NRS=61.476 M=1 R=2.8
+ SA=75000.3 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1002 N_VGND_M1002_d N_A_1068_21#_M1002_g A_996_73# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0847 PD=1.41 PS=0.91 NRD=0 NRS=41.904 M=1 R=2.8 SA=75000.5
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1038 A_1336_97# N_A_887_139#_M1038_g N_A_1068_21#_M1038_s VNB NSHORT L=0.15
+ W=0.42 AD=0.05145 AS=0.1197 PD=0.665 PS=1.41 NRD=19.284 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75003.4 A=0.063 P=1.14 MULT=1
MM1003 N_VGND_M1003_d N_SET_B_M1003_g A_1336_97# VNB NSHORT L=0.15 W=0.42
+ AD=0.131547 AS=0.05145 PD=0.998491 PS=0.665 NRD=18.564 NRS=19.284 M=1 R=2.8
+ SA=75000.6 SB=75003 A=0.063 P=1.14 MULT=1
MM1040 N_A_1541_125#_M1040_d N_A_887_139#_M1040_g N_VGND_M1003_d VNB NSHORT
+ L=0.15 W=0.64 AD=0.136 AS=0.200453 PD=1.065 PS=1.52151 NRD=27.18 NRS=26.244
+ M=1 R=4.26667 SA=75000.7 SB=75003 A=0.096 P=1.58 MULT=1
MM1025 A_1656_125# N_A_689_139#_M1025_g N_A_1541_125#_M1040_d VNB NSHORT L=0.15
+ W=0.64 AD=0.0672 AS=0.136 PD=0.85 PS=1.065 NRD=9.372 NRS=0 M=1 R=4.26667
+ SA=75001.3 SB=75002.4 A=0.096 P=1.58 MULT=1
MM1017 N_A_1728_125#_M1017_d N_A_689_139#_M1017_g A_1656_125# VNB NSHORT L=0.15
+ W=0.64 AD=0.322355 AS=0.0672 PD=1.81132 PS=0.85 NRD=46.872 NRS=9.372 M=1
+ R=4.26667 SA=75001.7 SB=75002.1 A=0.096 P=1.58 MULT=1
MM1050 A_1930_125# N_A_659_113#_M1050_g N_A_1728_125#_M1017_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.211545 PD=0.63 PS=1.18868 NRD=14.28 NRS=128.184 M=1
+ R=2.8 SA=75002.9 SB=75001.8 A=0.063 P=1.14 MULT=1
MM1046 A_2002_125# N_A_1972_99#_M1046_g A_1930_125# VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0441 PD=0.63 PS=0.63 NRD=14.28 NRS=14.28 M=1 R=2.8 SA=75003.2
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1006 N_A_2074_125#_M1006_d N_A_1972_99#_M1006_g A_2002_125# VNB NSHORT L=0.15
+ W=0.42 AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75003.6
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1008 N_VGND_M1008_d N_SET_B_M1008_g N_A_2074_125#_M1006_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75004
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1044 N_A_2074_125#_M1044_d N_A_2216_99#_M1044_g N_VGND_M1008_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.1155 AS=0.0588 PD=1.39 PS=0.7 NRD=0 NRS=0 M=1 R=2.8
+ SA=75004.5 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1051 A_2463_119# N_A_1728_125#_M1051_g N_VGND_M1051_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1638 PD=0.63 PS=1.62 NRD=14.28 NRS=32.856 M=1 R=2.8 SA=75000.3
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1041 N_A_1972_99#_M1041_d N_A_1728_125#_M1041_g A_2463_119# VNB NSHORT L=0.15
+ W=0.42 AD=0.2282 AS=0.0441 PD=2.08 PS=0.63 NRD=139.512 NRS=14.28 M=1 R=2.8
+ SA=75000.7 SB=75000.3 A=0.063 P=1.14 MULT=1
MM1015 A_3056_72# N_CLK_M1015_g N_A_659_113#_M1015_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.18105 PD=0.66 PS=1.73 NRD=18.564 NRS=32.856 M=1 R=2.8
+ SA=75000.3 SB=75001.7 A=0.063 P=1.14 MULT=1
MM1014 A_3134_72# N_SLEEP_B_M1014_g A_3056_72# VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0504 PD=0.63 PS=0.66 NRD=14.28 NRS=18.564 M=1 R=2.8 SA=75000.7
+ SB=75001.3 A=0.063 P=1.14 MULT=1
MM1049 N_VGND_M1049_d N_SLEEP_B_M1049_g A_3134_72# VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.1
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1020 A_3292_72# N_SLEEP_B_M1020_g N_VGND_M1049_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75001.5
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1022 N_A_2216_99#_M1022_d N_SLEEP_B_M1022_g A_3292_72# VNB NSHORT L=0.15
+ W=0.42 AD=0.1134 AS=0.0441 PD=1.38 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8
+ SA=75001.9 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1007 N_VGND_M1007_d N_A_1728_125#_M1007_g N_A_3466_403#_M1007_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.0924 AS=0.1134 PD=0.816667 PS=1.38 NRD=30 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1033 N_Q_M1033_d N_A_3466_403#_M1033_g N_VGND_M1007_d VNB NSHORT L=0.15 W=0.84
+ AD=0.2268 AS=0.1848 PD=2.22 PS=1.63333 NRD=0 NRS=0 M=1 R=5.6 SA=75000.5
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1000 N_VPWR_M1000_d N_SCD_M1000_g N_A_27_481#_M1000_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1152 AS=0.1728 PD=1 PS=1.82 NRD=21.5321 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75001.5 A=0.096 P=1.58 MULT=1
MM1042 A_213_481# N_SCE_M1042_g N_VPWR_M1000_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0768 AS=0.1152 PD=0.88 PS=1 NRD=19.9955 NRS=3.0732 M=1 R=4.26667
+ SA=75000.7 SB=75001 A=0.096 P=1.58 MULT=1
MM1012 N_A_189_119#_M1012_d N_D_M1012_g A_213_481# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0896 AS=0.0768 PD=0.92 PS=0.88 NRD=0 NRS=19.9955 M=1 R=4.26667 SA=75001.1
+ SB=75000.6 A=0.096 P=1.58 MULT=1
MM1048 N_A_27_481#_M1048_d N_A_339_93#_M1048_g N_A_189_119#_M1012_d VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.1728 AS=0.0896 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75001.5 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1036 N_VPWR_M1036_d N_SCE_M1036_g N_A_339_93#_M1036_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.2428 AS=0.1728 PD=1.66 PS=1.82 NRD=99.8396 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75000.9 A=0.096 P=1.58 MULT=1
MM1010 N_A_689_139#_M1010_d N_A_659_113#_M1010_g N_VPWR_M1036_d VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.1728 AS=0.2428 PD=1.82 PS=1.66 NRD=0 NRS=99.8396 M=1
+ R=4.26667 SA=75000.9 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1005 N_A_887_139#_M1005_d N_A_689_139#_M1005_g N_A_189_119#_M1005_s VPB
+ PHIGHVT L=0.15 W=0.42 AD=0.0588 AS=0.1491 PD=0.7 PS=1.55 NRD=0 NRS=32.8202 M=1
+ R=2.8 SA=75000.3 SB=75001.6 A=0.063 P=1.14 MULT=1
MM1034 A_1132_535# N_A_659_113#_M1034_g N_A_887_139#_M1005_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0504 AS=0.0588 PD=0.66 PS=0.7 NRD=30.4759 NRS=0 M=1 R=2.8
+ SA=75000.7 SB=75001.2 A=0.063 P=1.14 MULT=1
MM1035 N_VPWR_M1035_d N_A_1068_21#_M1035_g A_1132_535# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0819 AS=0.0504 PD=0.81 PS=0.66 NRD=0 NRS=30.4759 M=1 R=2.8 SA=75001.1
+ SB=75000.8 A=0.063 P=1.14 MULT=1
MM1009 N_A_1068_21#_M1009_d N_A_887_139#_M1009_g N_VPWR_M1035_d VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.12705 AS=0.0819 PD=1.235 PS=0.81 NRD=116.072 NRS=51.5943
+ M=1 R=2.8 SA=75001.6 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1027 N_VPWR_M1027_d N_SET_B_M1027_g N_A_1068_21#_M1009_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0987 AS=0.12705 PD=0.84 PS=1.235 NRD=65.6601 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75002 A=0.063 P=1.14 MULT=1
MM1032 N_A_1541_125#_M1032_d N_A_887_139#_M1032_g N_VPWR_M1027_d VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.2961 AS=0.1974 PD=1.545 PS=1.68 NRD=99.6623 NRS=0 M=1 R=5.6
+ SA=75000.5 SB=75001.4 A=0.126 P=1.98 MULT=1
MM1030 A_1712_451# N_A_659_113#_M1030_g N_A_1541_125#_M1032_d VPB PHIGHVT L=0.15
+ W=0.84 AD=0.0882 AS=0.2961 PD=1.05 PS=1.545 NRD=11.7215 NRS=0 M=1 R=5.6
+ SA=75001.3 SB=75000.6 A=0.126 P=1.98 MULT=1
MM1037 N_A_1728_125#_M1037_d N_A_659_113#_M1037_g A_1712_451# VPB PHIGHVT L=0.15
+ W=0.84 AD=0.2394 AS=0.0882 PD=2.25 PS=1.05 NRD=0 NRS=11.7215 M=1 R=5.6
+ SA=75001.7 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1018 N_KAPWR_M1018_d N_A_1728_125#_M1018_g N_A_1972_99#_M1018_s VPB PHIGHVT
+ L=0.25 W=1 AD=0.235112 AS=0.855 PD=1.57 PS=3.71 NRD=16.7253 NRS=112.27 M=1 R=4
+ SA=125001 SB=125003 A=0.25 P=2.5 MULT=1
MM1024 A_2658_414# N_A_2216_99#_M1024_g N_KAPWR_M1018_d VPB PHIGHVT L=0.25 W=1
+ AD=0.12 AS=0.235112 PD=1.24 PS=1.57 NRD=12.7853 NRS=16.7253 M=1 R=4 SA=125001
+ SB=125003 A=0.25 P=2.5 MULT=1
MM1043 N_A_1728_125#_M1043_d N_SET_B_M1043_g A_2658_414# VPB PHIGHVT L=0.25 W=1
+ AD=0.14 AS=0.12 PD=1.28 PS=1.24 NRD=0 NRS=12.7853 M=1 R=4 SA=125002 SB=125002
+ A=0.25 P=2.5 MULT=1
MM1021 A_2862_414# N_A_689_139#_M1021_g N_A_1728_125#_M1043_d VPB PHIGHVT L=0.25
+ W=1 AD=0.135 AS=0.14 PD=1.27 PS=1.28 NRD=15.7403 NRS=0 M=1 R=4 SA=125002
+ SB=125002 A=0.25 P=2.5 MULT=1
MM1011 N_KAPWR_M1011_d N_A_1972_99#_M1011_g A_2862_414# VPB PHIGHVT L=0.25 W=1
+ AD=0.292317 AS=0.135 PD=1.9878 PS=1.27 NRD=19.7 NRS=15.7403 M=1 R=4 SA=125003
+ SB=125001 A=0.25 P=2.5 MULT=1
MM1039 N_A_659_113#_M1039_d N_CLK_M1039_g N_KAPWR_M1011_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.0896 AS=0.187083 PD=0.92 PS=1.2722 NRD=0 NRS=73.0476 M=1 R=4.26667
+ SA=75002.9 SB=75001.3 A=0.096 P=1.58 MULT=1
MM1026 N_KAPWR_M1026_d N_SLEEP_B_M1026_g N_A_659_113#_M1039_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.136741 AS=0.0896 PD=1.08488 PS=0.92 NRD=48.8363 NRS=0 M=1
+ R=4.26667 SA=75003.4 SB=75000.8 A=0.096 P=1.58 MULT=1
MM1045 N_A_2216_99#_M1045_d N_SLEEP_B_M1045_g N_KAPWR_M1026_d VPB PHIGHVT L=0.25
+ W=1 AD=0.285 AS=0.213659 PD=2.57 PS=1.69512 NRD=0 NRS=0 M=1 R=4 SA=125003
+ SB=125000 A=0.25 P=2.5 MULT=1
MM1019 N_VPWR_M1019_d N_A_1728_125#_M1019_g N_A_3466_403#_M1019_s VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.144674 AS=0.1824 PD=1.11495 PS=1.85 NRD=36.1495 NRS=0 M=1
+ R=4.26667 SA=75000.2 SB=75000.7 A=0.096 P=1.58 MULT=1
MM1004 N_Q_M1004_d N_A_3466_403#_M1004_g N_VPWR_M1019_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3465 AS=0.284826 PD=3.07 PS=2.19505 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.5 SB=75000.2 A=0.189 P=2.82 MULT=1
DX52_noxref VNB VPB NWDIODE A=35.7817 P=42.11
c_3020 A_1656_125# 0 5.02674e-20 $X=8.28 $Y=0.625
*
.include "sky130_fd_sc_lp__srsdfstp_1.pxi.spice"
*
.ends
*
*
