* File: sky130_fd_sc_lp__sregrbp_1.pxi.spice
* Created: Wed Sep  2 10:38:50 2020
* 
x_PM_SKY130_FD_SC_LP__SREGRBP_1%SCE N_SCE_M1022_g N_SCE_M1041_g N_SCE_c_296_n
+ N_SCE_M1000_g N_SCE_M1024_g N_SCE_c_298_n N_SCE_c_299_n N_SCE_c_300_n SCE SCE
+ N_SCE_c_301_n N_SCE_c_302_n SCE N_SCE_c_303_n
+ PM_SKY130_FD_SC_LP__SREGRBP_1%SCE
x_PM_SKY130_FD_SC_LP__SREGRBP_1%A_75_531# N_A_75_531#_M1022_d
+ N_A_75_531#_M1041_s N_A_75_531#_c_375_n N_A_75_531#_c_376_n
+ N_A_75_531#_M1012_g N_A_75_531#_M1030_g N_A_75_531#_c_377_n
+ N_A_75_531#_c_383_n N_A_75_531#_c_384_n N_A_75_531#_c_385_n
+ N_A_75_531#_c_378_n N_A_75_531#_c_379_n N_A_75_531#_c_386_n
+ N_A_75_531#_c_387_n N_A_75_531#_c_380_n
+ PM_SKY130_FD_SC_LP__SREGRBP_1%A_75_531#
x_PM_SKY130_FD_SC_LP__SREGRBP_1%D N_D_c_450_n N_D_M1020_g N_D_M1013_g D
+ PM_SKY130_FD_SC_LP__SREGRBP_1%D
x_PM_SKY130_FD_SC_LP__SREGRBP_1%SCD N_SCD_c_487_n N_SCD_M1028_g N_SCD_M1025_g
+ SCD SCD PM_SKY130_FD_SC_LP__SREGRBP_1%SCD
x_PM_SKY130_FD_SC_LP__SREGRBP_1%A_342_531# N_A_342_531#_M1013_d
+ N_A_342_531#_M1020_d N_A_342_531#_M1031_g N_A_342_531#_c_533_n
+ N_A_342_531#_M1036_g N_A_342_531#_c_534_n N_A_342_531#_c_535_n
+ N_A_342_531#_c_536_n N_A_342_531#_c_550_n N_A_342_531#_c_544_n
+ N_A_342_531#_c_545_n N_A_342_531#_c_537_n N_A_342_531#_c_538_n
+ N_A_342_531#_c_539_n N_A_342_531#_c_540_n N_A_342_531#_c_547_n
+ N_A_342_531#_c_548_n N_A_342_531#_c_541_n N_A_342_531#_c_549_n
+ PM_SKY130_FD_SC_LP__SREGRBP_1%A_342_531#
x_PM_SKY130_FD_SC_LP__SREGRBP_1%CLK N_CLK_c_645_n N_CLK_M1005_g N_CLK_c_647_n
+ N_CLK_M1039_g CLK PM_SKY130_FD_SC_LP__SREGRBP_1%CLK
x_PM_SKY130_FD_SC_LP__SREGRBP_1%A_934_357# N_A_934_357#_M1043_d
+ N_A_934_357#_M1029_d N_A_934_357#_M1009_g N_A_934_357#_c_689_n
+ N_A_934_357#_M1037_g N_A_934_357#_M1027_g N_A_934_357#_c_691_n
+ N_A_934_357#_M1007_g N_A_934_357#_c_708_n N_A_934_357#_c_692_n
+ N_A_934_357#_c_693_n N_A_934_357#_c_694_n N_A_934_357#_c_695_n
+ N_A_934_357#_c_696_n N_A_934_357#_c_697_n N_A_934_357#_c_698_n
+ N_A_934_357#_c_699_n N_A_934_357#_c_700_n N_A_934_357#_c_701_n
+ N_A_934_357#_c_702_n N_A_934_357#_c_703_n
+ PM_SKY130_FD_SC_LP__SREGRBP_1%A_934_357#
x_PM_SKY130_FD_SC_LP__SREGRBP_1%A_1273_393# N_A_1273_393#_M1010_d
+ N_A_1273_393#_M1019_s N_A_1273_393#_M1034_d N_A_1273_393#_M1033_g
+ N_A_1273_393#_M1001_g N_A_1273_393#_c_868_n N_A_1273_393#_M1002_g
+ N_A_1273_393#_M1018_g N_A_1273_393#_c_877_n N_A_1273_393#_c_894_n
+ N_A_1273_393#_c_878_n N_A_1273_393#_c_879_n N_A_1273_393#_c_880_n
+ N_A_1273_393#_c_869_n N_A_1273_393#_c_870_n N_A_1273_393#_c_882_n
+ N_A_1273_393#_c_883_n N_A_1273_393#_c_871_n N_A_1273_393#_c_884_n
+ N_A_1273_393#_c_885_n N_A_1273_393#_c_872_n N_A_1273_393#_c_873_n
+ PM_SKY130_FD_SC_LP__SREGRBP_1%A_1273_393#
x_PM_SKY130_FD_SC_LP__SREGRBP_1%A_1139_463# N_A_1139_463#_M1032_d
+ N_A_1139_463#_M1009_d N_A_1139_463#_M1038_g N_A_1139_463#_M1019_g
+ N_A_1139_463#_c_1017_n N_A_1139_463#_c_1010_n N_A_1139_463#_c_1011_n
+ N_A_1139_463#_c_1012_n N_A_1139_463#_c_1013_n N_A_1139_463#_c_1014_n
+ N_A_1139_463#_c_1015_n PM_SKY130_FD_SC_LP__SREGRBP_1%A_1139_463#
x_PM_SKY130_FD_SC_LP__SREGRBP_1%ASYNC N_ASYNC_M1010_g N_ASYNC_M1034_g
+ N_ASYNC_c_1099_n N_ASYNC_M1003_g N_ASYNC_M1035_g N_ASYNC_c_1100_n
+ N_ASYNC_c_1106_n N_ASYNC_c_1107_n N_ASYNC_c_1101_n N_ASYNC_c_1108_n
+ N_ASYNC_c_1121_n N_ASYNC_c_1109_n ASYNC N_ASYNC_c_1102_n N_ASYNC_c_1103_n
+ N_ASYNC_c_1113_n PM_SKY130_FD_SC_LP__SREGRBP_1%ASYNC
x_PM_SKY130_FD_SC_LP__SREGRBP_1%A_761_357# N_A_761_357#_M1039_s
+ N_A_761_357#_M1005_s N_A_761_357#_M1029_g N_A_761_357#_c_1233_n
+ N_A_761_357#_M1043_g N_A_761_357#_c_1234_n N_A_761_357#_c_1235_n
+ N_A_761_357#_c_1246_n N_A_761_357#_c_1247_n N_A_761_357#_M1032_g
+ N_A_761_357#_M1017_g N_A_761_357#_c_1237_n N_A_761_357#_c_1238_n
+ N_A_761_357#_c_1249_n N_A_761_357#_M1042_g N_A_761_357#_M1021_g
+ N_A_761_357#_c_1251_n N_A_761_357#_c_1252_n N_A_761_357#_c_1257_n
+ N_A_761_357#_c_1253_n N_A_761_357#_c_1254_n N_A_761_357#_c_1270_n
+ N_A_761_357#_c_1260_n N_A_761_357#_c_1240_n N_A_761_357#_c_1241_n
+ N_A_761_357#_c_1242_n N_A_761_357#_c_1243_n
+ PM_SKY130_FD_SC_LP__SREGRBP_1%A_761_357#
x_PM_SKY130_FD_SC_LP__SREGRBP_1%A_2083_65# N_A_2083_65#_M1003_d
+ N_A_2083_65#_M1015_d N_A_2083_65#_M1006_g N_A_2083_65#_M1008_g
+ N_A_2083_65#_M1023_g N_A_2083_65#_M1026_g N_A_2083_65#_c_1416_n
+ N_A_2083_65#_M1011_g N_A_2083_65#_M1004_g N_A_2083_65#_c_1419_n
+ N_A_2083_65#_c_1420_n N_A_2083_65#_c_1421_n N_A_2083_65#_c_1434_n
+ N_A_2083_65#_c_1422_n N_A_2083_65#_c_1423_n N_A_2083_65#_c_1458_n
+ N_A_2083_65#_c_1443_n N_A_2083_65#_c_1424_n N_A_2083_65#_c_1425_n
+ N_A_2083_65#_c_1435_n N_A_2083_65#_c_1436_n N_A_2083_65#_c_1426_n
+ N_A_2083_65#_c_1472_n N_A_2083_65#_c_1427_n N_A_2083_65#_c_1428_n
+ N_A_2083_65#_c_1429_n N_A_2083_65#_c_1430_n
+ PM_SKY130_FD_SC_LP__SREGRBP_1%A_2083_65#
x_PM_SKY130_FD_SC_LP__SREGRBP_1%A_1903_125# N_A_1903_125#_M1027_d
+ N_A_1903_125#_M1042_d N_A_1903_125#_M1040_g N_A_1903_125#_M1015_g
+ N_A_1903_125#_c_1585_n N_A_1903_125#_c_1586_n N_A_1903_125#_c_1587_n
+ N_A_1903_125#_c_1588_n N_A_1903_125#_c_1597_n N_A_1903_125#_c_1594_n
+ N_A_1903_125#_c_1589_n N_A_1903_125#_c_1590_n N_A_1903_125#_c_1591_n
+ N_A_1903_125#_c_1592_n PM_SKY130_FD_SC_LP__SREGRBP_1%A_1903_125#
x_PM_SKY130_FD_SC_LP__SREGRBP_1%A_2456_451# N_A_2456_451#_M1026_d
+ N_A_2456_451#_M1023_d N_A_2456_451#_M1014_g N_A_2456_451#_M1016_g
+ N_A_2456_451#_c_1677_n N_A_2456_451#_c_1684_n N_A_2456_451#_c_1678_n
+ N_A_2456_451#_c_1686_n N_A_2456_451#_c_1687_n N_A_2456_451#_c_1679_n
+ N_A_2456_451#_c_1680_n N_A_2456_451#_c_1681_n
+ PM_SKY130_FD_SC_LP__SREGRBP_1%A_2456_451#
x_PM_SKY130_FD_SC_LP__SREGRBP_1%VPWR N_VPWR_M1041_d N_VPWR_M1028_d
+ N_VPWR_M1005_d N_VPWR_M1033_d N_VPWR_M1019_d N_VPWR_M1018_s N_VPWR_M1008_d
+ N_VPWR_M1035_d N_VPWR_M1011_d N_VPWR_c_1776_n N_VPWR_c_1777_n N_VPWR_c_1778_n
+ N_VPWR_c_1779_n N_VPWR_c_1780_n N_VPWR_c_1781_n N_VPWR_c_1782_n
+ N_VPWR_c_1783_n N_VPWR_c_1784_n N_VPWR_c_1785_n N_VPWR_c_1786_n
+ N_VPWR_c_1787_n N_VPWR_c_1788_n N_VPWR_c_1789_n N_VPWR_c_1790_n
+ N_VPWR_c_1791_n N_VPWR_c_1792_n N_VPWR_c_1793_n N_VPWR_c_1794_n
+ N_VPWR_c_1795_n N_VPWR_c_1796_n N_VPWR_c_1797_n VPWR N_VPWR_c_1798_n
+ N_VPWR_c_1799_n N_VPWR_c_1800_n N_VPWR_c_1775_n N_VPWR_c_1802_n
+ N_VPWR_c_1803_n N_VPWR_c_1804_n PM_SKY130_FD_SC_LP__SREGRBP_1%VPWR
x_PM_SKY130_FD_SC_LP__SREGRBP_1%A_636_531# N_A_636_531#_M1036_d
+ N_A_636_531#_M1032_s N_A_636_531#_M1031_d N_A_636_531#_M1009_s
+ N_A_636_531#_c_1963_n N_A_636_531#_c_1971_n N_A_636_531#_c_1972_n
+ N_A_636_531#_c_1973_n N_A_636_531#_c_1964_n N_A_636_531#_c_1975_n
+ N_A_636_531#_c_1965_n N_A_636_531#_c_1966_n N_A_636_531#_c_1967_n
+ N_A_636_531#_c_1968_n N_A_636_531#_c_1969_n
+ PM_SKY130_FD_SC_LP__SREGRBP_1%A_636_531#
x_PM_SKY130_FD_SC_LP__SREGRBP_1%Q N_Q_M1004_s N_Q_M1011_s N_Q_c_2095_n
+ N_Q_c_2086_n N_Q_c_2101_n Q N_Q_c_2084_n PM_SKY130_FD_SC_LP__SREGRBP_1%Q
x_PM_SKY130_FD_SC_LP__SREGRBP_1%Q_N N_Q_N_M1016_d N_Q_N_M1014_d N_Q_N_c_2128_n
+ N_Q_N_c_2123_n N_Q_N_c_2124_n N_Q_N_c_2125_n N_Q_N_c_2143_n N_Q_N_c_2126_n Q_N
+ N_Q_N_c_2130_n N_Q_N_c_2127_n PM_SKY130_FD_SC_LP__SREGRBP_1%Q_N
x_PM_SKY130_FD_SC_LP__SREGRBP_1%VGND N_VGND_M1022_s N_VGND_M1012_s
+ N_VGND_M1025_d N_VGND_M1039_d N_VGND_M1001_d N_VGND_M1002_s N_VGND_M1006_d
+ N_VGND_M1026_s N_VGND_M1004_d N_VGND_c_2168_n N_VGND_c_2169_n N_VGND_c_2170_n
+ N_VGND_c_2171_n N_VGND_c_2172_n N_VGND_c_2173_n N_VGND_c_2174_n
+ N_VGND_c_2175_n N_VGND_c_2176_n N_VGND_c_2177_n N_VGND_c_2178_n
+ N_VGND_c_2179_n N_VGND_c_2180_n N_VGND_c_2181_n N_VGND_c_2182_n
+ N_VGND_c_2183_n VGND N_VGND_c_2184_n N_VGND_c_2185_n N_VGND_c_2186_n
+ N_VGND_c_2187_n N_VGND_c_2188_n N_VGND_c_2189_n N_VGND_c_2190_n
+ N_VGND_c_2191_n N_VGND_c_2192_n N_VGND_c_2193_n N_VGND_c_2194_n
+ N_VGND_c_2195_n PM_SKY130_FD_SC_LP__SREGRBP_1%VGND
cc_1 VNB N_SCE_M1022_g 0.0710623f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.48
cc_2 VNB N_SCE_c_296_n 0.0110437f $X=-0.19 $Y=-0.245 $X2=1.17 $Y2=1.73
cc_3 VNB N_SCE_M1024_g 0.0420922f $X=-0.19 $Y=-0.245 $X2=2.355 $Y2=0.445
cc_4 VNB N_SCE_c_298_n 0.0164454f $X=-0.19 $Y=-0.245 $X2=2.13 $Y2=1.72
cc_5 VNB N_SCE_c_299_n 0.00216011f $X=-0.19 $Y=-0.245 $X2=2.295 $Y2=1.45
cc_6 VNB N_SCE_c_300_n 0.0354022f $X=-0.19 $Y=-0.245 $X2=2.295 $Y2=1.45
cc_7 VNB N_SCE_c_301_n 0.0233261f $X=-0.19 $Y=-0.245 $X2=0.81 $Y2=1.64
cc_8 VNB N_SCE_c_302_n 0.0025232f $X=-0.19 $Y=-0.245 $X2=1.15 $Y2=1.64
cc_9 VNB N_SCE_c_303_n 0.00433576f $X=-0.19 $Y=-0.245 $X2=1.315 $Y2=1.64
cc_10 VNB N_A_75_531#_c_375_n 0.0329769f $X=-0.19 $Y=-0.245 $X2=0.735 $Y2=2.865
cc_11 VNB N_A_75_531#_c_376_n 0.0190473f $X=-0.19 $Y=-0.245 $X2=1.17 $Y2=1.73
cc_12 VNB N_A_75_531#_c_377_n 0.0211908f $X=-0.19 $Y=-0.245 $X2=2.355 $Y2=0.445
cc_13 VNB N_A_75_531#_c_378_n 0.00769483f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_14 VNB N_A_75_531#_c_379_n 0.0308856f $X=-0.19 $Y=-0.245 $X2=0.645 $Y2=1.64
cc_15 VNB N_A_75_531#_c_380_n 0.0466874f $X=-0.19 $Y=-0.245 $X2=0.645 $Y2=1.64
cc_16 VNB N_D_c_450_n 0.0754631f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.475
cc_17 VNB N_D_M1020_g 0.00288266f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.48
cc_18 VNB N_D_M1013_g 0.0237457f $X=-0.19 $Y=-0.245 $X2=0.735 $Y2=2.865
cc_19 VNB D 0.00966136f $X=-0.19 $Y=-0.245 $X2=1.17 $Y2=1.73
cc_20 VNB N_SCD_c_487_n 0.0563146f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.475
cc_21 VNB N_SCD_M1025_g 0.0391519f $X=-0.19 $Y=-0.245 $X2=0.735 $Y2=2.865
cc_22 VNB SCD 0.00552779f $X=-0.19 $Y=-0.245 $X2=1.17 $Y2=1.73
cc_23 VNB N_A_342_531#_c_533_n 0.0196904f $X=-0.19 $Y=-0.245 $X2=1.245 $Y2=1.805
cc_24 VNB N_A_342_531#_c_534_n 0.0299508f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_342_531#_c_535_n 0.00828572f $X=-0.19 $Y=-0.245 $X2=2.355
+ $Y2=1.285
cc_26 VNB N_A_342_531#_c_536_n 0.0351055f $X=-0.19 $Y=-0.245 $X2=2.355 $Y2=0.445
cc_27 VNB N_A_342_531#_c_537_n 0.00172632f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_342_531#_c_538_n 0.0103581f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_29 VNB N_A_342_531#_c_539_n 0.00301951f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_30 VNB N_A_342_531#_c_540_n 0.00493076f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_342_531#_c_541_n 0.00634756f $X=-0.19 $Y=-0.245 $X2=0.735 $Y2=1.64
cc_32 VNB N_CLK_c_645_n 0.0400996f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.475
cc_33 VNB N_CLK_M1005_g 0.00522655f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.48
cc_34 VNB N_CLK_c_647_n 0.0210779f $X=-0.19 $Y=-0.245 $X2=0.735 $Y2=1.805
cc_35 VNB CLK 0.00470615f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_934_357#_c_689_n 0.0452783f $X=-0.19 $Y=-0.245 $X2=1.245 $Y2=1.805
cc_37 VNB N_A_934_357#_M1037_g 0.029448f $X=-0.19 $Y=-0.245 $X2=2.355 $Y2=1.285
cc_38 VNB N_A_934_357#_c_691_n 0.0211034f $X=-0.19 $Y=-0.245 $X2=1.315 $Y2=1.72
cc_39 VNB N_A_934_357#_c_692_n 0.00690511f $X=-0.19 $Y=-0.245 $X2=0.645 $Y2=1.64
cc_40 VNB N_A_934_357#_c_693_n 0.00637357f $X=-0.19 $Y=-0.245 $X2=2.295 $Y2=1.45
cc_41 VNB N_A_934_357#_c_694_n 4.91165e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_934_357#_c_695_n 0.00172668f $X=-0.19 $Y=-0.245 $X2=1.15 $Y2=1.64
cc_43 VNB N_A_934_357#_c_696_n 0.0156744f $X=-0.19 $Y=-0.245 $X2=0.645 $Y2=1.64
cc_44 VNB N_A_934_357#_c_697_n 0.0032936f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_934_357#_c_698_n 0.00478873f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=1.64
cc_46 VNB N_A_934_357#_c_699_n 0.00144069f $X=-0.19 $Y=-0.245 $X2=1.315 $Y2=1.64
cc_47 VNB N_A_934_357#_c_700_n 0.00771921f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_934_357#_c_701_n 0.00763098f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_934_357#_c_702_n 0.0247947f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_934_357#_c_703_n 0.0168702f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_1273_393#_M1001_g 0.0414798f $X=-0.19 $Y=-0.245 $X2=2.355
+ $Y2=0.445
cc_52 VNB N_A_1273_393#_c_868_n 0.0167358f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_1273_393#_c_869_n 0.00600968f $X=-0.19 $Y=-0.245 $X2=0.645
+ $Y2=1.64
cc_54 VNB N_A_1273_393#_c_870_n 0.0100937f $X=-0.19 $Y=-0.245 $X2=2.295
+ $Y2=1.285
cc_55 VNB N_A_1273_393#_c_871_n 0.0166226f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_1273_393#_c_872_n 0.00331131f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_1273_393#_c_873_n 0.0323801f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_1139_463#_M1038_g 0.0169117f $X=-0.19 $Y=-0.245 $X2=1.17 $Y2=1.73
cc_59 VNB N_A_1139_463#_c_1010_n 0.00466651f $X=-0.19 $Y=-0.245 $X2=2.29
+ $Y2=1.635
cc_60 VNB N_A_1139_463#_c_1011_n 0.00134958f $X=-0.19 $Y=-0.245 $X2=2.295
+ $Y2=1.45
cc_61 VNB N_A_1139_463#_c_1012_n 0.0147685f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_A_1139_463#_c_1013_n 0.00196047f $X=-0.19 $Y=-0.245 $X2=1.115
+ $Y2=1.58
cc_63 VNB N_A_1139_463#_c_1014_n 0.00168955f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_A_1139_463#_c_1015_n 0.0229051f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_ASYNC_M1010_g 0.020844f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.48
cc_66 VNB N_ASYNC_c_1099_n 0.0195829f $X=-0.19 $Y=-0.245 $X2=1.17 $Y2=1.73
cc_67 VNB N_ASYNC_c_1100_n 0.021871f $X=-0.19 $Y=-0.245 $X2=1.315 $Y2=1.72
cc_68 VNB N_ASYNC_c_1101_n 0.0017094f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_ASYNC_c_1102_n 0.0321502f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_ASYNC_c_1103_n 0.0276015f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=1.665
cc_71 VNB N_A_761_357#_M1029_g 0.00243562f $X=-0.19 $Y=-0.245 $X2=1.17 $Y2=1.73
cc_72 VNB N_A_761_357#_c_1233_n 0.0207501f $X=-0.19 $Y=-0.245 $X2=1.245
+ $Y2=1.805
cc_73 VNB N_A_761_357#_c_1234_n 0.00317772f $X=-0.19 $Y=-0.245 $X2=2.355
+ $Y2=1.285
cc_74 VNB N_A_761_357#_c_1235_n 0.0468598f $X=-0.19 $Y=-0.245 $X2=2.355
+ $Y2=0.445
cc_75 VNB N_A_761_357#_M1032_g 0.0384531f $X=-0.19 $Y=-0.245 $X2=2.295 $Y2=1.45
cc_76 VNB N_A_761_357#_c_1237_n 0.326967f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_A_761_357#_c_1238_n 0.012806f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_A_761_357#_M1021_g 0.0263479f $X=-0.19 $Y=-0.245 $X2=2.295 $Y2=1.45
cc_79 VNB N_A_761_357#_c_1240_n 0.00260863f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_A_761_357#_c_1241_n 8.80678e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_A_761_357#_c_1242_n 0.00298293f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_A_761_357#_c_1243_n 0.0519986f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_A_2083_65#_M1026_g 0.0662089f $X=-0.19 $Y=-0.245 $X2=2.29 $Y2=1.45
cc_84 VNB N_A_2083_65#_c_1416_n 0.0637166f $X=-0.19 $Y=-0.245 $X2=2.295 $Y2=1.45
cc_85 VNB N_A_2083_65#_M1011_g 0.00301752f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_A_2083_65#_M1004_g 0.0351674f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_A_2083_65#_c_1419_n 0.0175793f $X=-0.19 $Y=-0.245 $X2=0.645 $Y2=1.64
cc_88 VNB N_A_2083_65#_c_1420_n 0.00834971f $X=-0.19 $Y=-0.245 $X2=0.645
+ $Y2=1.64
cc_89 VNB N_A_2083_65#_c_1421_n 0.00661055f $X=-0.19 $Y=-0.245 $X2=0.735
+ $Y2=1.64
cc_90 VNB N_A_2083_65#_c_1422_n 0.0110145f $X=-0.19 $Y=-0.245 $X2=1.15 $Y2=1.64
cc_91 VNB N_A_2083_65#_c_1423_n 0.00348886f $X=-0.19 $Y=-0.245 $X2=0.645
+ $Y2=1.64
cc_92 VNB N_A_2083_65#_c_1424_n 0.0179606f $X=-0.19 $Y=-0.245 $X2=1.315 $Y2=1.64
cc_93 VNB N_A_2083_65#_c_1425_n 0.0171095f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_94 VNB N_A_2083_65#_c_1426_n 5.68065e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_95 VNB N_A_2083_65#_c_1427_n 0.00131482f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_96 VNB N_A_2083_65#_c_1428_n 0.0077949f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_97 VNB N_A_2083_65#_c_1429_n 0.0301054f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_98 VNB N_A_2083_65#_c_1430_n 0.0187633f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_99 VNB N_A_1903_125#_M1015_g 0.00673344f $X=-0.19 $Y=-0.245 $X2=1.245
+ $Y2=2.865
cc_100 VNB N_A_1903_125#_c_1585_n 0.0181538f $X=-0.19 $Y=-0.245 $X2=2.355
+ $Y2=1.285
cc_101 VNB N_A_1903_125#_c_1586_n 0.0152279f $X=-0.19 $Y=-0.245 $X2=2.355
+ $Y2=0.445
cc_102 VNB N_A_1903_125#_c_1587_n 0.0264141f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_103 VNB N_A_1903_125#_c_1588_n 0.00690059f $X=-0.19 $Y=-0.245 $X2=2.29
+ $Y2=1.635
cc_104 VNB N_A_1903_125#_c_1589_n 0.00743296f $X=-0.19 $Y=-0.245 $X2=0.645
+ $Y2=1.64
cc_105 VNB N_A_1903_125#_c_1590_n 0.00323287f $X=-0.19 $Y=-0.245 $X2=0.735
+ $Y2=1.64
cc_106 VNB N_A_1903_125#_c_1591_n 0.013823f $X=-0.19 $Y=-0.245 $X2=0.81 $Y2=1.64
cc_107 VNB N_A_1903_125#_c_1592_n 0.023883f $X=-0.19 $Y=-0.245 $X2=2.295
+ $Y2=1.45
cc_108 VNB N_A_2456_451#_M1016_g 0.0279996f $X=-0.19 $Y=-0.245 $X2=1.245
+ $Y2=2.865
cc_109 VNB N_A_2456_451#_c_1677_n 0.0158726f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_110 VNB N_A_2456_451#_c_1678_n 2.75776e-19 $X=-0.19 $Y=-0.245 $X2=2.29
+ $Y2=1.45
cc_111 VNB N_A_2456_451#_c_1679_n 0.0123747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_112 VNB N_A_2456_451#_c_1680_n 0.00268035f $X=-0.19 $Y=-0.245 $X2=0.645
+ $Y2=1.64
cc_113 VNB N_A_2456_451#_c_1681_n 0.0293591f $X=-0.19 $Y=-0.245 $X2=0.735
+ $Y2=1.64
cc_114 VNB N_VPWR_c_1775_n 0.601534f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_115 VNB N_A_636_531#_c_1963_n 0.00911435f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_116 VNB N_A_636_531#_c_1964_n 0.00701325f $X=-0.19 $Y=-0.245 $X2=2.29
+ $Y2=1.45
cc_117 VNB N_A_636_531#_c_1965_n 0.00764552f $X=-0.19 $Y=-0.245 $X2=0.635
+ $Y2=1.58
cc_118 VNB N_A_636_531#_c_1966_n 0.001907f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.58
cc_119 VNB N_A_636_531#_c_1967_n 0.00974815f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_120 VNB N_A_636_531#_c_1968_n 0.00245596f $X=-0.19 $Y=-0.245 $X2=0.645
+ $Y2=1.64
cc_121 VNB N_A_636_531#_c_1969_n 0.0183354f $X=-0.19 $Y=-0.245 $X2=1.132
+ $Y2=1.64
cc_122 VNB N_Q_c_2084_n 0.0142306f $X=-0.19 $Y=-0.245 $X2=2.355 $Y2=0.445
cc_123 VNB N_Q_N_c_2123_n 0.0304981f $X=-0.19 $Y=-0.245 $X2=1.245 $Y2=2.865
cc_124 VNB N_Q_N_c_2124_n 0.00952577f $X=-0.19 $Y=-0.245 $X2=2.355 $Y2=0.445
cc_125 VNB N_Q_N_c_2125_n 0.0018979f $X=-0.19 $Y=-0.245 $X2=2.13 $Y2=1.72
cc_126 VNB N_Q_N_c_2126_n 0.00530503f $X=-0.19 $Y=-0.245 $X2=2.295 $Y2=1.45
cc_127 VNB N_Q_N_c_2127_n 0.0237016f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_128 VNB N_VGND_c_2168_n 0.010678f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_129 VNB N_VGND_c_2169_n 0.026105f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_130 VNB N_VGND_c_2170_n 0.0101458f $X=-0.19 $Y=-0.245 $X2=0.645 $Y2=1.64
cc_131 VNB N_VGND_c_2171_n 0.00566391f $X=-0.19 $Y=-0.245 $X2=2.295 $Y2=1.45
cc_132 VNB N_VGND_c_2172_n 0.00561774f $X=-0.19 $Y=-0.245 $X2=0.645 $Y2=1.64
cc_133 VNB N_VGND_c_2173_n 0.0201098f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=1.64
cc_134 VNB N_VGND_c_2174_n 0.0241786f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_135 VNB N_VGND_c_2175_n 0.00550687f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_136 VNB N_VGND_c_2176_n 0.0209096f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_137 VNB N_VGND_c_2177_n 0.0102417f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_138 VNB N_VGND_c_2178_n 0.0380947f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_139 VNB N_VGND_c_2179_n 0.00359553f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_140 VNB N_VGND_c_2180_n 0.066136f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_141 VNB N_VGND_c_2181_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_142 VNB N_VGND_c_2182_n 0.0332467f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_143 VNB N_VGND_c_2183_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_144 VNB N_VGND_c_2184_n 0.0204586f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_145 VNB N_VGND_c_2185_n 0.034187f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_146 VNB N_VGND_c_2186_n 0.0350017f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_147 VNB N_VGND_c_2187_n 0.0523189f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_148 VNB N_VGND_c_2188_n 0.028322f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_149 VNB N_VGND_c_2189_n 0.0192273f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_150 VNB N_VGND_c_2190_n 0.712208f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_151 VNB N_VGND_c_2191_n 0.00513431f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_152 VNB N_VGND_c_2192_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_153 VNB N_VGND_c_2193_n 0.00332923f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_154 VNB N_VGND_c_2194_n 0.00513431f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_155 VNB N_VGND_c_2195_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_156 VPB N_SCE_M1041_g 0.0660819f $X=-0.19 $Y=1.655 $X2=0.735 $Y2=2.865
cc_157 VPB N_SCE_c_296_n 0.0248918f $X=-0.19 $Y=1.655 $X2=1.17 $Y2=1.73
cc_158 VPB N_SCE_M1000_g 0.0531565f $X=-0.19 $Y=1.655 $X2=1.245 $Y2=2.865
cc_159 VPB N_SCE_c_298_n 0.0146609f $X=-0.19 $Y=1.655 $X2=2.13 $Y2=1.72
cc_160 VPB N_SCE_c_301_n 0.0161725f $X=-0.19 $Y=1.655 $X2=0.81 $Y2=1.64
cc_161 VPB N_A_75_531#_M1030_g 0.0290178f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_162 VPB N_A_75_531#_c_377_n 0.0162548f $X=-0.19 $Y=1.655 $X2=2.355 $Y2=0.445
cc_163 VPB N_A_75_531#_c_383_n 0.0169846f $X=-0.19 $Y=1.655 $X2=2.13 $Y2=1.72
cc_164 VPB N_A_75_531#_c_384_n 0.0381863f $X=-0.19 $Y=1.655 $X2=2.29 $Y2=1.45
cc_165 VPB N_A_75_531#_c_385_n 0.0315753f $X=-0.19 $Y=1.655 $X2=2.295 $Y2=1.45
cc_166 VPB N_A_75_531#_c_386_n 0.015515f $X=-0.19 $Y=1.655 $X2=0.735 $Y2=1.64
cc_167 VPB N_A_75_531#_c_387_n 0.0266481f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_168 VPB N_D_M1020_g 0.0635012f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=0.48
cc_169 VPB N_SCD_c_487_n 0.0602671f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=1.475
cc_170 VPB N_SCD_M1028_g 0.0464325f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=0.48
cc_171 VPB SCD 0.00276926f $X=-0.19 $Y=1.655 $X2=1.17 $Y2=1.73
cc_172 VPB N_A_342_531#_M1031_g 0.0238846f $X=-0.19 $Y=1.655 $X2=1.17 $Y2=1.73
cc_173 VPB N_A_342_531#_c_536_n 0.0298391f $X=-0.19 $Y=1.655 $X2=2.355 $Y2=0.445
cc_174 VPB N_A_342_531#_c_544_n 0.00922203f $X=-0.19 $Y=1.655 $X2=2.29 $Y2=1.45
cc_175 VPB N_A_342_531#_c_545_n 0.00254143f $X=-0.19 $Y=1.655 $X2=2.295 $Y2=1.45
cc_176 VPB N_A_342_531#_c_540_n 0.00858203f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_177 VPB N_A_342_531#_c_547_n 0.00551021f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_178 VPB N_A_342_531#_c_548_n 0.0569269f $X=-0.19 $Y=1.655 $X2=0.645 $Y2=1.64
cc_179 VPB N_A_342_531#_c_549_n 0.00190264f $X=-0.19 $Y=1.655 $X2=2.295
+ $Y2=1.285
cc_180 VPB N_CLK_M1005_g 0.0226807f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=0.48
cc_181 VPB N_A_934_357#_M1009_g 0.0336635f $X=-0.19 $Y=1.655 $X2=1.17 $Y2=1.73
cc_182 VPB N_A_934_357#_c_689_n 0.024417f $X=-0.19 $Y=1.655 $X2=1.245 $Y2=1.805
cc_183 VPB N_A_934_357#_c_691_n 0.0133115f $X=-0.19 $Y=1.655 $X2=1.315 $Y2=1.72
cc_184 VPB N_A_934_357#_M1007_g 0.0405869f $X=-0.19 $Y=1.655 $X2=2.295 $Y2=1.45
cc_185 VPB N_A_934_357#_c_708_n 0.0140892f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_186 VPB N_A_934_357#_c_694_n 0.00823874f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_187 VPB N_A_934_357#_c_696_n 0.0202058f $X=-0.19 $Y=1.655 $X2=0.645 $Y2=1.64
cc_188 VPB N_A_934_357#_c_698_n 0.00288672f $X=-0.19 $Y=1.655 $X2=1.2 $Y2=1.64
cc_189 VPB N_A_934_357#_c_699_n 0.00303615f $X=-0.19 $Y=1.655 $X2=1.315 $Y2=1.64
cc_190 VPB N_A_934_357#_c_700_n 0.00594476f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_191 VPB N_A_934_357#_c_701_n 0.0200642f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_192 VPB N_A_934_357#_c_702_n 0.00891327f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_193 VPB N_A_1273_393#_M1033_g 0.021428f $X=-0.19 $Y=1.655 $X2=1.245 $Y2=2.865
cc_194 VPB N_A_1273_393#_M1001_g 0.00728893f $X=-0.19 $Y=1.655 $X2=2.355
+ $Y2=0.445
cc_195 VPB N_A_1273_393#_M1018_g 0.0245022f $X=-0.19 $Y=1.655 $X2=2.295 $Y2=1.45
cc_196 VPB N_A_1273_393#_c_877_n 0.00252725f $X=-0.19 $Y=1.655 $X2=0.635
+ $Y2=1.58
cc_197 VPB N_A_1273_393#_c_878_n 0.00621672f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_198 VPB N_A_1273_393#_c_879_n 0.0010399f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_199 VPB N_A_1273_393#_c_880_n 0.00245813f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_200 VPB N_A_1273_393#_c_870_n 0.00348441f $X=-0.19 $Y=1.655 $X2=2.295
+ $Y2=1.285
cc_201 VPB N_A_1273_393#_c_882_n 0.0564459f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_202 VPB N_A_1273_393#_c_883_n 0.0152468f $X=-0.19 $Y=1.655 $X2=1.2 $Y2=1.64
cc_203 VPB N_A_1273_393#_c_884_n 0.00409487f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_204 VPB N_A_1273_393#_c_885_n 0.00590959f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_205 VPB N_A_1273_393#_c_872_n 4.94381e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_206 VPB N_A_1273_393#_c_873_n 0.0129879f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_207 VPB N_A_1139_463#_M1019_g 0.0219666f $X=-0.19 $Y=1.655 $X2=1.245
+ $Y2=2.865
cc_208 VPB N_A_1139_463#_c_1017_n 0.00487107f $X=-0.19 $Y=1.655 $X2=2.355
+ $Y2=1.285
cc_209 VPB N_A_1139_463#_c_1011_n 0.00701418f $X=-0.19 $Y=1.655 $X2=2.295
+ $Y2=1.45
cc_210 VPB N_A_1139_463#_c_1014_n 6.39154e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_211 VPB N_A_1139_463#_c_1015_n 0.00804f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_212 VPB N_ASYNC_M1034_g 0.0212978f $X=-0.19 $Y=1.655 $X2=0.735 $Y2=2.865
cc_213 VPB N_ASYNC_M1035_g 0.0229992f $X=-0.19 $Y=1.655 $X2=2.355 $Y2=0.445
cc_214 VPB N_ASYNC_c_1106_n 0.00181908f $X=-0.19 $Y=1.655 $X2=2.295 $Y2=1.45
cc_215 VPB N_ASYNC_c_1107_n 0.0368598f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_216 VPB N_ASYNC_c_1108_n 0.0352224f $X=-0.19 $Y=1.655 $X2=0.645 $Y2=1.64
cc_217 VPB N_ASYNC_c_1109_n 0.00177791f $X=-0.19 $Y=1.655 $X2=0.81 $Y2=1.64
cc_218 VPB ASYNC 0.00229403f $X=-0.19 $Y=1.655 $X2=2.295 $Y2=1.285
cc_219 VPB N_ASYNC_c_1102_n 0.0116521f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_220 VPB N_ASYNC_c_1103_n 0.00651044f $X=-0.19 $Y=1.655 $X2=1.2 $Y2=1.665
cc_221 VPB N_ASYNC_c_1113_n 0.00280008f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_222 VPB N_A_761_357#_M1029_g 0.0199261f $X=-0.19 $Y=1.655 $X2=1.17 $Y2=1.73
cc_223 VPB N_A_761_357#_c_1234_n 0.0806358f $X=-0.19 $Y=1.655 $X2=2.355
+ $Y2=1.285
cc_224 VPB N_A_761_357#_c_1246_n 0.0546513f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_225 VPB N_A_761_357#_c_1247_n 0.0108815f $X=-0.19 $Y=1.655 $X2=2.13 $Y2=1.72
cc_226 VPB N_A_761_357#_M1017_g 0.0353294f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_227 VPB N_A_761_357#_c_1249_n 0.273687f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_228 VPB N_A_761_357#_M1042_g 0.0263823f $X=-0.19 $Y=1.655 $X2=0.645 $Y2=1.64
cc_229 VPB N_A_761_357#_c_1251_n 0.00749069f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_230 VPB N_A_761_357#_c_1252_n 0.00168903f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_231 VPB N_A_761_357#_c_1253_n 0.00401098f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_232 VPB N_A_761_357#_c_1254_n 0.00199332f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_233 VPB N_A_761_357#_c_1241_n 8.35774e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_234 VPB N_A_2083_65#_M1008_g 0.0206956f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_235 VPB N_A_2083_65#_M1023_g 0.0437306f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_236 VPB N_A_2083_65#_M1011_g 0.0253738f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_237 VPB N_A_2083_65#_c_1434_n 0.00154814f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_238 VPB N_A_2083_65#_c_1435_n 5.30273e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_239 VPB N_A_2083_65#_c_1436_n 0.0327416f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_240 VPB N_A_2083_65#_c_1426_n 0.00213514f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_241 VPB N_A_2083_65#_c_1428_n 0.00315917f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_242 VPB N_A_2083_65#_c_1429_n 0.0062895f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_243 VPB N_A_2083_65#_c_1430_n 0.0173179f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_244 VPB N_A_1903_125#_M1015_g 0.0454468f $X=-0.19 $Y=1.655 $X2=1.245
+ $Y2=2.865
cc_245 VPB N_A_1903_125#_c_1594_n 0.0163062f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_246 VPB N_A_1903_125#_c_1589_n 0.0091936f $X=-0.19 $Y=1.655 $X2=0.645
+ $Y2=1.64
cc_247 VPB N_A_2456_451#_M1014_g 0.0250215f $X=-0.19 $Y=1.655 $X2=1.17 $Y2=1.73
cc_248 VPB N_A_2456_451#_c_1677_n 0.0133331f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_249 VPB N_A_2456_451#_c_1684_n 0.0113012f $X=-0.19 $Y=1.655 $X2=2.13 $Y2=1.72
cc_250 VPB N_A_2456_451#_c_1678_n 0.00232453f $X=-0.19 $Y=1.655 $X2=2.29
+ $Y2=1.45
cc_251 VPB N_A_2456_451#_c_1686_n 0.0101388f $X=-0.19 $Y=1.655 $X2=2.295
+ $Y2=1.45
cc_252 VPB N_A_2456_451#_c_1687_n 0.0115895f $X=-0.19 $Y=1.655 $X2=1.115
+ $Y2=1.58
cc_253 VPB N_A_2456_451#_c_1681_n 0.00562432f $X=-0.19 $Y=1.655 $X2=0.735
+ $Y2=1.64
cc_254 VPB N_VPWR_c_1776_n 0.00727356f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_255 VPB N_VPWR_c_1777_n 0.00341245f $X=-0.19 $Y=1.655 $X2=0.645 $Y2=1.64
cc_256 VPB N_VPWR_c_1778_n 0.00177638f $X=-0.19 $Y=1.655 $X2=2.295 $Y2=1.45
cc_257 VPB N_VPWR_c_1779_n 0.0215003f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_258 VPB N_VPWR_c_1780_n 0.0211064f $X=-0.19 $Y=1.655 $X2=1.217 $Y2=1.64
cc_259 VPB N_VPWR_c_1781_n 0.022087f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_260 VPB N_VPWR_c_1782_n 0.0178711f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_261 VPB N_VPWR_c_1783_n 0.0188675f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_262 VPB N_VPWR_c_1784_n 0.00935938f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_263 VPB N_VPWR_c_1785_n 0.002833f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_264 VPB N_VPWR_c_1786_n 0.0245555f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_265 VPB N_VPWR_c_1787_n 0.00526006f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_266 VPB N_VPWR_c_1788_n 0.0385678f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_267 VPB N_VPWR_c_1789_n 0.00525412f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_268 VPB N_VPWR_c_1790_n 0.0328786f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_269 VPB N_VPWR_c_1791_n 0.00497896f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_270 VPB N_VPWR_c_1792_n 0.0549467f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_271 VPB N_VPWR_c_1793_n 0.00330333f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_272 VPB N_VPWR_c_1794_n 0.0209455f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_273 VPB N_VPWR_c_1795_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_274 VPB N_VPWR_c_1796_n 0.039753f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_275 VPB N_VPWR_c_1797_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_276 VPB N_VPWR_c_1798_n 0.021333f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_277 VPB N_VPWR_c_1799_n 0.0495026f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_278 VPB N_VPWR_c_1800_n 0.0199052f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_279 VPB N_VPWR_c_1775_n 0.127546f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_280 VPB N_VPWR_c_1802_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_281 VPB N_VPWR_c_1803_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_282 VPB N_VPWR_c_1804_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_283 VPB N_A_636_531#_c_1963_n 0.0120047f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_284 VPB N_A_636_531#_c_1971_n 0.00665077f $X=-0.19 $Y=1.655 $X2=2.355
+ $Y2=0.445
cc_285 VPB N_A_636_531#_c_1972_n 0.00620592f $X=-0.19 $Y=1.655 $X2=2.13 $Y2=1.72
cc_286 VPB N_A_636_531#_c_1973_n 0.00380503f $X=-0.19 $Y=1.655 $X2=1.315
+ $Y2=1.72
cc_287 VPB N_A_636_531#_c_1964_n 0.00597269f $X=-0.19 $Y=1.655 $X2=2.29 $Y2=1.45
cc_288 VPB N_A_636_531#_c_1975_n 0.00784607f $X=-0.19 $Y=1.655 $X2=2.295
+ $Y2=1.45
cc_289 VPB N_Q_c_2084_n 0.00450473f $X=-0.19 $Y=1.655 $X2=2.355 $Y2=0.445
cc_290 VPB N_Q_N_c_2128_n 0.0435135f $X=-0.19 $Y=1.655 $X2=1.17 $Y2=1.73
cc_291 VPB N_Q_N_c_2125_n 0.00156922f $X=-0.19 $Y=1.655 $X2=2.13 $Y2=1.72
cc_292 VPB N_Q_N_c_2130_n 0.0108816f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_293 VPB N_Q_N_c_2127_n 0.00848377f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_294 N_SCE_c_302_n N_A_75_531#_c_375_n 0.00429869f $X=1.15 $Y=1.64 $X2=0 $Y2=0
cc_295 N_SCE_M1022_g N_A_75_531#_c_377_n 0.0178906f $X=0.495 $Y=0.48 $X2=0 $Y2=0
cc_296 N_SCE_M1041_g N_A_75_531#_c_377_n 0.00500796f $X=0.735 $Y=2.865 $X2=0
+ $Y2=0
cc_297 N_SCE_c_302_n N_A_75_531#_c_377_n 0.0250949f $X=1.15 $Y=1.64 $X2=0 $Y2=0
cc_298 N_SCE_M1041_g N_A_75_531#_c_383_n 0.00893862f $X=0.735 $Y=2.865 $X2=0
+ $Y2=0
cc_299 N_SCE_M1041_g N_A_75_531#_c_384_n 0.0254817f $X=0.735 $Y=2.865 $X2=0
+ $Y2=0
cc_300 N_SCE_c_296_n N_A_75_531#_c_384_n 0.00348417f $X=1.17 $Y=1.73 $X2=0 $Y2=0
cc_301 N_SCE_M1000_g N_A_75_531#_c_384_n 0.0214255f $X=1.245 $Y=2.865 $X2=0
+ $Y2=0
cc_302 N_SCE_c_298_n N_A_75_531#_c_384_n 0.0118533f $X=2.13 $Y=1.72 $X2=0 $Y2=0
cc_303 N_SCE_c_301_n N_A_75_531#_c_384_n 0.00706118f $X=0.81 $Y=1.64 $X2=0 $Y2=0
cc_304 N_SCE_c_302_n N_A_75_531#_c_384_n 0.121998f $X=1.15 $Y=1.64 $X2=0 $Y2=0
cc_305 N_SCE_c_298_n N_A_75_531#_c_385_n 0.00575476f $X=2.13 $Y=1.72 $X2=0 $Y2=0
cc_306 N_SCE_c_300_n N_A_75_531#_c_385_n 0.00441123f $X=2.295 $Y=1.45 $X2=0
+ $Y2=0
cc_307 N_SCE_M1022_g N_A_75_531#_c_378_n 0.0163639f $X=0.495 $Y=0.48 $X2=0 $Y2=0
cc_308 N_SCE_M1022_g N_A_75_531#_c_379_n 0.0249258f $X=0.495 $Y=0.48 $X2=0 $Y2=0
cc_309 N_SCE_c_296_n N_A_75_531#_c_379_n 3.2663e-19 $X=1.17 $Y=1.73 $X2=0 $Y2=0
cc_310 N_SCE_c_301_n N_A_75_531#_c_379_n 0.00572422f $X=0.81 $Y=1.64 $X2=0 $Y2=0
cc_311 N_SCE_c_302_n N_A_75_531#_c_379_n 0.0382378f $X=1.15 $Y=1.64 $X2=0 $Y2=0
cc_312 N_SCE_M1041_g N_A_75_531#_c_387_n 0.00601092f $X=0.735 $Y=2.865 $X2=0
+ $Y2=0
cc_313 N_SCE_M1022_g N_A_75_531#_c_380_n 0.0249774f $X=0.495 $Y=0.48 $X2=0 $Y2=0
cc_314 N_SCE_c_296_n N_A_75_531#_c_380_n 0.0078743f $X=1.17 $Y=1.73 $X2=0 $Y2=0
cc_315 N_SCE_c_302_n N_A_75_531#_c_380_n 0.00281168f $X=1.15 $Y=1.64 $X2=0 $Y2=0
cc_316 N_SCE_M1024_g N_D_c_450_n 0.00920164f $X=2.355 $Y=0.445 $X2=-0.19
+ $Y2=-0.245
cc_317 N_SCE_c_298_n N_D_c_450_n 0.00777507f $X=2.13 $Y=1.72 $X2=-0.19
+ $Y2=-0.245
cc_318 N_SCE_c_299_n N_D_c_450_n 0.00173431f $X=2.295 $Y=1.45 $X2=-0.19
+ $Y2=-0.245
cc_319 N_SCE_c_300_n N_D_c_450_n 0.0210326f $X=2.295 $Y=1.45 $X2=-0.19
+ $Y2=-0.245
cc_320 N_SCE_c_303_n N_D_c_450_n 0.0064771f $X=1.315 $Y=1.64 $X2=-0.19
+ $Y2=-0.245
cc_321 N_SCE_c_296_n N_D_M1020_g 0.0838128f $X=1.17 $Y=1.73 $X2=0 $Y2=0
cc_322 N_SCE_c_298_n N_D_M1020_g 0.0126236f $X=2.13 $Y=1.72 $X2=0 $Y2=0
cc_323 N_SCE_c_299_n N_D_M1020_g 5.7739e-19 $X=2.295 $Y=1.45 $X2=0 $Y2=0
cc_324 N_SCE_M1024_g N_D_M1013_g 0.01995f $X=2.355 $Y=0.445 $X2=0 $Y2=0
cc_325 N_SCE_M1024_g D 8.8592e-19 $X=2.355 $Y=0.445 $X2=0 $Y2=0
cc_326 N_SCE_c_298_n D 0.0231875f $X=2.13 $Y=1.72 $X2=0 $Y2=0
cc_327 N_SCE_c_299_n D 0.00964191f $X=2.295 $Y=1.45 $X2=0 $Y2=0
cc_328 N_SCE_c_300_n D 5.63661e-19 $X=2.295 $Y=1.45 $X2=0 $Y2=0
cc_329 N_SCE_c_298_n N_SCD_c_487_n 0.00119376f $X=2.13 $Y=1.72 $X2=-0.19
+ $Y2=-0.245
cc_330 N_SCE_c_299_n N_SCD_c_487_n 5.00583e-19 $X=2.295 $Y=1.45 $X2=-0.19
+ $Y2=-0.245
cc_331 N_SCE_c_300_n N_SCD_c_487_n 0.0207009f $X=2.295 $Y=1.45 $X2=-0.19
+ $Y2=-0.245
cc_332 N_SCE_M1024_g N_SCD_M1025_g 0.0611447f $X=2.355 $Y=0.445 $X2=0 $Y2=0
cc_333 N_SCE_M1000_g N_A_342_531#_c_550_n 0.00113139f $X=1.245 $Y=2.865 $X2=0
+ $Y2=0
cc_334 N_SCE_M1000_g N_A_342_531#_c_545_n 7.71857e-19 $X=1.245 $Y=2.865 $X2=0
+ $Y2=0
cc_335 N_SCE_M1024_g N_A_342_531#_c_537_n 0.00445341f $X=2.355 $Y=0.445 $X2=0
+ $Y2=0
cc_336 N_SCE_M1024_g N_A_342_531#_c_538_n 0.00881891f $X=2.355 $Y=0.445 $X2=0
+ $Y2=0
cc_337 N_SCE_c_299_n N_A_342_531#_c_538_n 0.00767558f $X=2.295 $Y=1.45 $X2=0
+ $Y2=0
cc_338 N_SCE_c_300_n N_A_342_531#_c_538_n 4.9771e-19 $X=2.295 $Y=1.45 $X2=0
+ $Y2=0
cc_339 N_SCE_M1024_g N_A_342_531#_c_539_n 0.00228437f $X=2.355 $Y=0.445 $X2=0
+ $Y2=0
cc_340 N_SCE_c_299_n N_A_342_531#_c_539_n 0.0106895f $X=2.295 $Y=1.45 $X2=0
+ $Y2=0
cc_341 N_SCE_c_300_n N_A_342_531#_c_539_n 0.00108988f $X=2.295 $Y=1.45 $X2=0
+ $Y2=0
cc_342 N_SCE_M1024_g N_A_342_531#_c_540_n 0.00505798f $X=2.355 $Y=0.445 $X2=0
+ $Y2=0
cc_343 N_SCE_c_298_n N_A_342_531#_c_540_n 0.0137852f $X=2.13 $Y=1.72 $X2=0 $Y2=0
cc_344 N_SCE_c_299_n N_A_342_531#_c_540_n 0.0251795f $X=2.295 $Y=1.45 $X2=0
+ $Y2=0
cc_345 N_SCE_c_300_n N_A_342_531#_c_540_n 0.00177932f $X=2.295 $Y=1.45 $X2=0
+ $Y2=0
cc_346 N_SCE_M1024_g N_A_342_531#_c_541_n 0.00735269f $X=2.355 $Y=0.445 $X2=0
+ $Y2=0
cc_347 N_SCE_M1041_g N_VPWR_c_1776_n 0.00536123f $X=0.735 $Y=2.865 $X2=0 $Y2=0
cc_348 N_SCE_M1000_g N_VPWR_c_1776_n 0.0131472f $X=1.245 $Y=2.865 $X2=0 $Y2=0
cc_349 N_SCE_M1041_g N_VPWR_c_1786_n 0.0052871f $X=0.735 $Y=2.865 $X2=0 $Y2=0
cc_350 N_SCE_M1000_g N_VPWR_c_1788_n 0.00469214f $X=1.245 $Y=2.865 $X2=0 $Y2=0
cc_351 N_SCE_M1041_g N_VPWR_c_1775_n 0.0109112f $X=0.735 $Y=2.865 $X2=0 $Y2=0
cc_352 N_SCE_M1000_g N_VPWR_c_1775_n 0.00818361f $X=1.245 $Y=2.865 $X2=0 $Y2=0
cc_353 N_SCE_M1022_g N_VGND_c_2169_n 0.00551061f $X=0.495 $Y=0.48 $X2=0 $Y2=0
cc_354 N_SCE_M1022_g N_VGND_c_2170_n 0.00283338f $X=0.495 $Y=0.48 $X2=0 $Y2=0
cc_355 N_SCE_M1024_g N_VGND_c_2171_n 0.00237638f $X=2.355 $Y=0.445 $X2=0 $Y2=0
cc_356 N_SCE_M1024_g N_VGND_c_2178_n 0.00549284f $X=2.355 $Y=0.445 $X2=0 $Y2=0
cc_357 N_SCE_M1022_g N_VGND_c_2184_n 0.00516215f $X=0.495 $Y=0.48 $X2=0 $Y2=0
cc_358 N_SCE_M1022_g N_VGND_c_2190_n 0.0114031f $X=0.495 $Y=0.48 $X2=0 $Y2=0
cc_359 N_SCE_M1024_g N_VGND_c_2190_n 0.00644159f $X=2.355 $Y=0.445 $X2=0 $Y2=0
cc_360 N_A_75_531#_c_375_n N_D_c_450_n 0.00140609f $X=1.41 $Y=0.84 $X2=-0.19
+ $Y2=-0.245
cc_361 N_A_75_531#_c_379_n N_D_c_450_n 0.00120837f $X=0.975 $Y=1.055 $X2=-0.19
+ $Y2=-0.245
cc_362 N_A_75_531#_c_380_n N_D_c_450_n 0.00530356f $X=0.975 $Y=0.84 $X2=-0.19
+ $Y2=-0.245
cc_363 N_A_75_531#_M1030_g N_D_M1020_g 0.0242768f $X=2.065 $Y=2.865 $X2=0 $Y2=0
cc_364 N_A_75_531#_c_384_n N_D_M1020_g 0.0198182f $X=2.115 $Y=2.15 $X2=0 $Y2=0
cc_365 N_A_75_531#_c_385_n N_D_M1020_g 0.0180926f $X=2.115 $Y=2.15 $X2=0 $Y2=0
cc_366 N_A_75_531#_c_376_n N_D_M1013_g 0.0425173f $X=1.485 $Y=0.765 $X2=0 $Y2=0
cc_367 N_A_75_531#_c_379_n D 0.00357528f $X=0.975 $Y=1.055 $X2=0 $Y2=0
cc_368 N_A_75_531#_c_384_n N_SCD_c_487_n 0.00112915f $X=2.115 $Y=2.15 $X2=-0.19
+ $Y2=-0.245
cc_369 N_A_75_531#_c_385_n N_SCD_c_487_n 0.0167057f $X=2.115 $Y=2.15 $X2=-0.19
+ $Y2=-0.245
cc_370 N_A_75_531#_M1030_g N_SCD_M1028_g 0.0282049f $X=2.065 $Y=2.865 $X2=0
+ $Y2=0
cc_371 N_A_75_531#_M1030_g N_A_342_531#_c_550_n 0.00827807f $X=2.065 $Y=2.865
+ $X2=0 $Y2=0
cc_372 N_A_75_531#_M1030_g N_A_342_531#_c_544_n 0.00911372f $X=2.065 $Y=2.865
+ $X2=0 $Y2=0
cc_373 N_A_75_531#_c_384_n N_A_342_531#_c_544_n 0.0185727f $X=2.115 $Y=2.15
+ $X2=0 $Y2=0
cc_374 N_A_75_531#_c_385_n N_A_342_531#_c_544_n 0.00311872f $X=2.115 $Y=2.15
+ $X2=0 $Y2=0
cc_375 N_A_75_531#_M1030_g N_A_342_531#_c_545_n 0.00260994f $X=2.065 $Y=2.865
+ $X2=0 $Y2=0
cc_376 N_A_75_531#_c_384_n N_A_342_531#_c_545_n 0.0270504f $X=2.115 $Y=2.15
+ $X2=0 $Y2=0
cc_377 N_A_75_531#_c_385_n N_A_342_531#_c_545_n 9.20695e-19 $X=2.115 $Y=2.15
+ $X2=0 $Y2=0
cc_378 N_A_75_531#_c_384_n N_A_342_531#_c_540_n 0.00758316f $X=2.115 $Y=2.15
+ $X2=0 $Y2=0
cc_379 N_A_75_531#_M1030_g N_A_342_531#_c_549_n 8.51233e-19 $X=2.065 $Y=2.865
+ $X2=0 $Y2=0
cc_380 N_A_75_531#_c_384_n N_A_342_531#_c_549_n 0.00705202f $X=2.115 $Y=2.15
+ $X2=0 $Y2=0
cc_381 N_A_75_531#_c_384_n N_VPWR_c_1776_n 0.0184717f $X=2.115 $Y=2.15 $X2=0
+ $Y2=0
cc_382 N_A_75_531#_c_387_n N_VPWR_c_1776_n 0.0174148f $X=0.52 $Y=2.85 $X2=0
+ $Y2=0
cc_383 N_A_75_531#_M1030_g N_VPWR_c_1777_n 0.00158451f $X=2.065 $Y=2.865 $X2=0
+ $Y2=0
cc_384 N_A_75_531#_c_387_n N_VPWR_c_1786_n 0.0337539f $X=0.52 $Y=2.85 $X2=0
+ $Y2=0
cc_385 N_A_75_531#_M1030_g N_VPWR_c_1788_n 0.00403185f $X=2.065 $Y=2.865 $X2=0
+ $Y2=0
cc_386 N_A_75_531#_M1030_g N_VPWR_c_1775_n 0.00600782f $X=2.065 $Y=2.865 $X2=0
+ $Y2=0
cc_387 N_A_75_531#_c_387_n N_VPWR_c_1775_n 0.021083f $X=0.52 $Y=2.85 $X2=0 $Y2=0
cc_388 N_A_75_531#_c_378_n N_VGND_c_2169_n 0.0168306f $X=0.71 $Y=0.485 $X2=0
+ $Y2=0
cc_389 N_A_75_531#_c_379_n N_VGND_c_2169_n 0.0198777f $X=0.975 $Y=1.055 $X2=0
+ $Y2=0
cc_390 N_A_75_531#_c_376_n N_VGND_c_2170_n 0.0156898f $X=1.485 $Y=0.765 $X2=0
+ $Y2=0
cc_391 N_A_75_531#_c_378_n N_VGND_c_2170_n 0.0276416f $X=0.71 $Y=0.485 $X2=0
+ $Y2=0
cc_392 N_A_75_531#_c_379_n N_VGND_c_2170_n 0.00240426f $X=0.975 $Y=1.055 $X2=0
+ $Y2=0
cc_393 N_A_75_531#_c_380_n N_VGND_c_2170_n 0.0130308f $X=0.975 $Y=0.84 $X2=0
+ $Y2=0
cc_394 N_A_75_531#_c_376_n N_VGND_c_2178_n 0.00486043f $X=1.485 $Y=0.765 $X2=0
+ $Y2=0
cc_395 N_A_75_531#_c_378_n N_VGND_c_2184_n 0.0218928f $X=0.71 $Y=0.485 $X2=0
+ $Y2=0
cc_396 N_A_75_531#_c_380_n N_VGND_c_2184_n 0.00439215f $X=0.975 $Y=0.84 $X2=0
+ $Y2=0
cc_397 N_A_75_531#_c_376_n N_VGND_c_2190_n 0.00827383f $X=1.485 $Y=0.765 $X2=0
+ $Y2=0
cc_398 N_A_75_531#_c_378_n N_VGND_c_2190_n 0.0125518f $X=0.71 $Y=0.485 $X2=0
+ $Y2=0
cc_399 N_A_75_531#_c_380_n N_VGND_c_2190_n 0.00576584f $X=0.975 $Y=0.84 $X2=0
+ $Y2=0
cc_400 N_D_M1020_g N_A_342_531#_c_550_n 0.00705574f $X=1.635 $Y=2.865 $X2=0
+ $Y2=0
cc_401 N_D_M1020_g N_A_342_531#_c_545_n 0.00540615f $X=1.635 $Y=2.865 $X2=0
+ $Y2=0
cc_402 N_D_M1013_g N_A_342_531#_c_537_n 0.00371231f $X=1.875 $Y=0.445 $X2=0
+ $Y2=0
cc_403 N_D_M1013_g N_A_342_531#_c_539_n 0.00463014f $X=1.875 $Y=0.445 $X2=0
+ $Y2=0
cc_404 N_D_M1013_g N_A_342_531#_c_541_n 3.31023e-19 $X=1.875 $Y=0.445 $X2=0
+ $Y2=0
cc_405 N_D_M1020_g N_VPWR_c_1776_n 0.0022911f $X=1.635 $Y=2.865 $X2=0 $Y2=0
cc_406 N_D_M1020_g N_VPWR_c_1788_n 0.00530134f $X=1.635 $Y=2.865 $X2=0 $Y2=0
cc_407 N_D_M1020_g N_VPWR_c_1775_n 0.0098253f $X=1.635 $Y=2.865 $X2=0 $Y2=0
cc_408 N_D_M1013_g N_VGND_c_2170_n 0.00242534f $X=1.875 $Y=0.445 $X2=0 $Y2=0
cc_409 N_D_M1013_g N_VGND_c_2178_n 0.00585385f $X=1.875 $Y=0.445 $X2=0 $Y2=0
cc_410 N_D_M1013_g N_VGND_c_2190_n 0.0110519f $X=1.875 $Y=0.445 $X2=0 $Y2=0
cc_411 N_SCD_M1025_g N_A_342_531#_c_533_n 0.0201484f $X=2.745 $Y=0.445 $X2=0
+ $Y2=0
cc_412 N_SCD_c_487_n N_A_342_531#_c_535_n 0.00954206f $X=2.595 $Y=2.005 $X2=0
+ $Y2=0
cc_413 SCD N_A_342_531#_c_535_n 0.00388693f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_414 N_SCD_c_487_n N_A_342_531#_c_536_n 0.0434038f $X=2.595 $Y=2.005 $X2=0
+ $Y2=0
cc_415 N_SCD_M1025_g N_A_342_531#_c_536_n 0.00310134f $X=2.745 $Y=0.445 $X2=0
+ $Y2=0
cc_416 SCD N_A_342_531#_c_536_n 0.00207658f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_417 N_SCD_M1028_g N_A_342_531#_c_550_n 0.00151887f $X=2.595 $Y=2.865 $X2=0
+ $Y2=0
cc_418 N_SCD_M1028_g N_A_342_531#_c_544_n 0.0114306f $X=2.595 $Y=2.865 $X2=0
+ $Y2=0
cc_419 N_SCD_M1025_g N_A_342_531#_c_538_n 0.0130785f $X=2.745 $Y=0.445 $X2=0
+ $Y2=0
cc_420 N_SCD_c_487_n N_A_342_531#_c_540_n 0.0393467f $X=2.595 $Y=2.005 $X2=0
+ $Y2=0
cc_421 N_SCD_M1028_g N_A_342_531#_c_540_n 0.00504997f $X=2.595 $Y=2.865 $X2=0
+ $Y2=0
cc_422 N_SCD_M1025_g N_A_342_531#_c_540_n 0.0080848f $X=2.745 $Y=0.445 $X2=0
+ $Y2=0
cc_423 SCD N_A_342_531#_c_540_n 0.0459184f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_424 N_SCD_c_487_n N_A_342_531#_c_547_n 0.00763969f $X=2.595 $Y=2.005 $X2=0
+ $Y2=0
cc_425 SCD N_A_342_531#_c_547_n 0.0158615f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_426 N_SCD_c_487_n N_A_342_531#_c_548_n 0.0108856f $X=2.595 $Y=2.005 $X2=0
+ $Y2=0
cc_427 N_SCD_M1028_g N_A_342_531#_c_548_n 0.0276531f $X=2.595 $Y=2.865 $X2=0
+ $Y2=0
cc_428 SCD N_A_342_531#_c_548_n 0.00117466f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_429 N_SCD_M1025_g N_A_342_531#_c_541_n 0.00205573f $X=2.745 $Y=0.445 $X2=0
+ $Y2=0
cc_430 N_SCD_M1028_g N_A_342_531#_c_549_n 0.0137814f $X=2.595 $Y=2.865 $X2=0
+ $Y2=0
cc_431 N_SCD_M1028_g N_VPWR_c_1777_n 0.00964326f $X=2.595 $Y=2.865 $X2=0 $Y2=0
cc_432 N_SCD_M1028_g N_VPWR_c_1788_n 0.00343267f $X=2.595 $Y=2.865 $X2=0 $Y2=0
cc_433 N_SCD_M1028_g N_VPWR_c_1775_n 0.00437946f $X=2.595 $Y=2.865 $X2=0 $Y2=0
cc_434 N_SCD_c_487_n N_A_636_531#_c_1963_n 0.00339915f $X=2.595 $Y=2.005 $X2=0
+ $Y2=0
cc_435 N_SCD_M1025_g N_A_636_531#_c_1963_n 0.00230768f $X=2.745 $Y=0.445 $X2=0
+ $Y2=0
cc_436 SCD N_A_636_531#_c_1963_n 0.0398719f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_437 N_SCD_M1028_g N_A_636_531#_c_1975_n 5.35812e-19 $X=2.595 $Y=2.865 $X2=0
+ $Y2=0
cc_438 SCD N_A_636_531#_c_1967_n 0.00299441f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_439 N_SCD_c_487_n N_VGND_c_2171_n 0.00582527f $X=2.595 $Y=2.005 $X2=0 $Y2=0
cc_440 N_SCD_M1025_g N_VGND_c_2171_n 0.0134276f $X=2.745 $Y=0.445 $X2=0 $Y2=0
cc_441 SCD N_VGND_c_2171_n 0.00276073f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_442 N_SCD_M1025_g N_VGND_c_2178_n 0.00486043f $X=2.745 $Y=0.445 $X2=0 $Y2=0
cc_443 N_SCD_M1025_g N_VGND_c_2190_n 0.00456736f $X=2.745 $Y=0.445 $X2=0 $Y2=0
cc_444 N_A_342_531#_c_536_n N_CLK_c_645_n 0.0208368f $X=3.585 $Y=2.165 $X2=-0.19
+ $Y2=-0.245
cc_445 N_A_342_531#_c_536_n N_CLK_M1005_g 0.0138961f $X=3.585 $Y=2.165 $X2=0
+ $Y2=0
cc_446 N_A_342_531#_c_534_n N_CLK_c_647_n 0.00605793f $X=3.51 $Y=0.84 $X2=0
+ $Y2=0
cc_447 N_A_342_531#_c_536_n CLK 4.18192e-19 $X=3.585 $Y=2.165 $X2=0 $Y2=0
cc_448 N_A_342_531#_c_536_n N_A_761_357#_c_1252_n 0.00151414f $X=3.585 $Y=2.165
+ $X2=0 $Y2=0
cc_449 N_A_342_531#_c_533_n N_A_761_357#_c_1257_n 5.68634e-19 $X=3.175 $Y=0.765
+ $X2=0 $Y2=0
cc_450 N_A_342_531#_c_534_n N_A_761_357#_c_1257_n 2.40674e-19 $X=3.51 $Y=0.84
+ $X2=0 $Y2=0
cc_451 N_A_342_531#_c_536_n N_A_761_357#_c_1254_n 7.14402e-19 $X=3.585 $Y=2.165
+ $X2=0 $Y2=0
cc_452 N_A_342_531#_c_534_n N_A_761_357#_c_1260_n 7.41751e-19 $X=3.51 $Y=0.84
+ $X2=0 $Y2=0
cc_453 N_A_342_531#_c_549_n N_VPWR_M1028_d 9.42151e-19 $X=2.715 $Y=2.415 $X2=0
+ $Y2=0
cc_454 N_A_342_531#_c_550_n N_VPWR_c_1776_n 0.0126564f $X=1.85 $Y=2.85 $X2=0
+ $Y2=0
cc_455 N_A_342_531#_c_545_n N_VPWR_c_1776_n 0.00100797f $X=2.015 $Y=2.58 $X2=0
+ $Y2=0
cc_456 N_A_342_531#_M1031_g N_VPWR_c_1777_n 0.00417866f $X=3.105 $Y=2.865 $X2=0
+ $Y2=0
cc_457 N_A_342_531#_c_550_n N_VPWR_c_1777_n 0.00555787f $X=1.85 $Y=2.85 $X2=0
+ $Y2=0
cc_458 N_A_342_531#_c_547_n N_VPWR_c_1777_n 0.00780288f $X=3.195 $Y=2.33 $X2=0
+ $Y2=0
cc_459 N_A_342_531#_c_549_n N_VPWR_c_1777_n 0.00766691f $X=2.715 $Y=2.415 $X2=0
+ $Y2=0
cc_460 N_A_342_531#_c_550_n N_VPWR_c_1788_n 0.0176777f $X=1.85 $Y=2.85 $X2=0
+ $Y2=0
cc_461 N_A_342_531#_c_544_n N_VPWR_c_1788_n 0.00895434f $X=2.63 $Y=2.58 $X2=0
+ $Y2=0
cc_462 N_A_342_531#_c_549_n N_VPWR_c_1788_n 2.34538e-19 $X=2.715 $Y=2.415 $X2=0
+ $Y2=0
cc_463 N_A_342_531#_M1031_g N_VPWR_c_1790_n 0.00528677f $X=3.105 $Y=2.865 $X2=0
+ $Y2=0
cc_464 N_A_342_531#_M1031_g N_VPWR_c_1775_n 0.00738776f $X=3.105 $Y=2.865 $X2=0
+ $Y2=0
cc_465 N_A_342_531#_c_550_n N_VPWR_c_1775_n 0.0124101f $X=1.85 $Y=2.85 $X2=0
+ $Y2=0
cc_466 N_A_342_531#_c_544_n N_VPWR_c_1775_n 0.0159829f $X=2.63 $Y=2.58 $X2=0
+ $Y2=0
cc_467 N_A_342_531#_c_547_n N_VPWR_c_1775_n 0.00684847f $X=3.195 $Y=2.33 $X2=0
+ $Y2=0
cc_468 N_A_342_531#_c_549_n N_VPWR_c_1775_n 0.00115251f $X=2.715 $Y=2.415 $X2=0
+ $Y2=0
cc_469 N_A_342_531#_c_544_n A_428_531# 0.00479126f $X=2.63 $Y=2.58 $X2=-0.19
+ $Y2=-0.245
cc_470 N_A_342_531#_M1031_g N_A_636_531#_c_1963_n 0.00512655f $X=3.105 $Y=2.865
+ $X2=0 $Y2=0
cc_471 N_A_342_531#_c_533_n N_A_636_531#_c_1963_n 0.00276776f $X=3.175 $Y=0.765
+ $X2=0 $Y2=0
cc_472 N_A_342_531#_c_534_n N_A_636_531#_c_1963_n 0.00850882f $X=3.51 $Y=0.84
+ $X2=0 $Y2=0
cc_473 N_A_342_531#_c_536_n N_A_636_531#_c_1963_n 0.0418976f $X=3.585 $Y=2.165
+ $X2=0 $Y2=0
cc_474 N_A_342_531#_c_547_n N_A_636_531#_c_1963_n 0.0246071f $X=3.195 $Y=2.33
+ $X2=0 $Y2=0
cc_475 N_A_342_531#_c_548_n N_A_636_531#_c_1963_n 0.0125575f $X=3.195 $Y=2.33
+ $X2=0 $Y2=0
cc_476 N_A_342_531#_M1031_g N_A_636_531#_c_1975_n 0.00635632f $X=3.105 $Y=2.865
+ $X2=0 $Y2=0
cc_477 N_A_342_531#_c_547_n N_A_636_531#_c_1975_n 0.010867f $X=3.195 $Y=2.33
+ $X2=0 $Y2=0
cc_478 N_A_342_531#_c_548_n N_A_636_531#_c_1975_n 0.00914168f $X=3.195 $Y=2.33
+ $X2=0 $Y2=0
cc_479 N_A_342_531#_c_533_n N_A_636_531#_c_1967_n 0.00541367f $X=3.175 $Y=0.765
+ $X2=0 $Y2=0
cc_480 N_A_342_531#_c_534_n N_A_636_531#_c_1967_n 0.0113113f $X=3.51 $Y=0.84
+ $X2=0 $Y2=0
cc_481 N_A_342_531#_c_541_n N_VGND_c_2170_n 0.0063109f $X=2.14 $Y=0.47 $X2=0
+ $Y2=0
cc_482 N_A_342_531#_c_533_n N_VGND_c_2171_n 0.00311162f $X=3.175 $Y=0.765 $X2=0
+ $Y2=0
cc_483 N_A_342_531#_c_541_n N_VGND_c_2171_n 0.0127186f $X=2.14 $Y=0.47 $X2=0
+ $Y2=0
cc_484 N_A_342_531#_c_541_n N_VGND_c_2178_n 0.0184519f $X=2.14 $Y=0.47 $X2=0
+ $Y2=0
cc_485 N_A_342_531#_c_533_n N_VGND_c_2185_n 0.00547815f $X=3.175 $Y=0.765 $X2=0
+ $Y2=0
cc_486 N_A_342_531#_M1013_d N_VGND_c_2190_n 0.00356108f $X=1.95 $Y=0.235 $X2=0
+ $Y2=0
cc_487 N_A_342_531#_c_533_n N_VGND_c_2190_n 0.0113613f $X=3.175 $Y=0.765 $X2=0
+ $Y2=0
cc_488 N_A_342_531#_c_538_n N_VGND_c_2190_n 0.0156578f $X=2.63 $Y=0.94 $X2=0
+ $Y2=0
cc_489 N_A_342_531#_c_541_n N_VGND_c_2190_n 0.0124996f $X=2.14 $Y=0.47 $X2=0
+ $Y2=0
cc_490 N_CLK_c_647_n N_A_934_357#_c_692_n 0.00105968f $X=4.205 $Y=1.185 $X2=0
+ $Y2=0
cc_491 N_CLK_M1005_g N_A_761_357#_M1029_g 0.0174217f $X=4.165 $Y=2.415 $X2=0
+ $Y2=0
cc_492 N_CLK_c_647_n N_A_761_357#_c_1233_n 0.0242116f $X=4.205 $Y=1.185 $X2=0
+ $Y2=0
cc_493 N_CLK_M1005_g N_A_761_357#_c_1252_n 0.00283499f $X=4.165 $Y=2.415 $X2=0
+ $Y2=0
cc_494 N_CLK_c_647_n N_A_761_357#_c_1257_n 0.00766071f $X=4.205 $Y=1.185 $X2=0
+ $Y2=0
cc_495 N_CLK_c_645_n N_A_761_357#_c_1253_n 0.00173739f $X=4.165 $Y=1.515 $X2=0
+ $Y2=0
cc_496 N_CLK_M1005_g N_A_761_357#_c_1253_n 0.0147518f $X=4.165 $Y=2.415 $X2=0
+ $Y2=0
cc_497 CLK N_A_761_357#_c_1253_n 0.011084f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_498 N_CLK_c_645_n N_A_761_357#_c_1254_n 0.00128836f $X=4.165 $Y=1.515 $X2=0
+ $Y2=0
cc_499 CLK N_A_761_357#_c_1254_n 0.0133227f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_500 N_CLK_c_647_n N_A_761_357#_c_1270_n 0.0103353f $X=4.205 $Y=1.185 $X2=0
+ $Y2=0
cc_501 CLK N_A_761_357#_c_1270_n 0.00255004f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_502 N_CLK_c_645_n N_A_761_357#_c_1260_n 0.00156296f $X=4.165 $Y=1.515 $X2=0
+ $Y2=0
cc_503 N_CLK_c_647_n N_A_761_357#_c_1260_n 7.41524e-19 $X=4.205 $Y=1.185 $X2=0
+ $Y2=0
cc_504 CLK N_A_761_357#_c_1260_n 0.01757f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_505 N_CLK_c_647_n N_A_761_357#_c_1240_n 0.00470977f $X=4.205 $Y=1.185 $X2=0
+ $Y2=0
cc_506 CLK N_A_761_357#_c_1240_n 0.00319955f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_507 N_CLK_M1005_g N_A_761_357#_c_1241_n 0.00300433f $X=4.165 $Y=2.415 $X2=0
+ $Y2=0
cc_508 N_CLK_c_645_n N_A_761_357#_c_1242_n 0.00321979f $X=4.165 $Y=1.515 $X2=0
+ $Y2=0
cc_509 CLK N_A_761_357#_c_1242_n 0.0226395f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_510 N_CLK_c_645_n N_A_761_357#_c_1243_n 0.0254154f $X=4.165 $Y=1.515 $X2=0
+ $Y2=0
cc_511 CLK N_A_761_357#_c_1243_n 2.92218e-19 $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_512 N_CLK_M1005_g N_VPWR_c_1778_n 0.0161534f $X=4.165 $Y=2.415 $X2=0 $Y2=0
cc_513 N_CLK_M1005_g N_VPWR_c_1790_n 0.00445056f $X=4.165 $Y=2.415 $X2=0 $Y2=0
cc_514 N_CLK_M1005_g N_VPWR_c_1775_n 0.00899805f $X=4.165 $Y=2.415 $X2=0 $Y2=0
cc_515 N_CLK_c_645_n N_A_636_531#_c_1963_n 0.00178325f $X=4.165 $Y=1.515 $X2=0
+ $Y2=0
cc_516 N_CLK_M1005_g N_A_636_531#_c_1963_n 0.00331335f $X=4.165 $Y=2.415 $X2=0
+ $Y2=0
cc_517 N_CLK_c_647_n N_A_636_531#_c_1963_n 0.00282475f $X=4.205 $Y=1.185 $X2=0
+ $Y2=0
cc_518 CLK N_A_636_531#_c_1963_n 0.0236179f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_519 N_CLK_c_647_n N_A_636_531#_c_1965_n 0.00338803f $X=4.205 $Y=1.185 $X2=0
+ $Y2=0
cc_520 CLK N_A_636_531#_c_1965_n 0.00219352f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_521 N_CLK_c_647_n N_A_636_531#_c_1967_n 6.54556e-19 $X=4.205 $Y=1.185 $X2=0
+ $Y2=0
cc_522 N_CLK_c_647_n N_VGND_c_2172_n 0.0057576f $X=4.205 $Y=1.185 $X2=0 $Y2=0
cc_523 N_CLK_c_647_n N_VGND_c_2185_n 0.00549284f $X=4.205 $Y=1.185 $X2=0 $Y2=0
cc_524 N_CLK_c_647_n N_VGND_c_2190_n 0.00682088f $X=4.205 $Y=1.185 $X2=0 $Y2=0
cc_525 N_A_934_357#_c_689_n N_A_1273_393#_M1001_g 0.00473157f $X=6.22 $Y=1.65
+ $X2=0 $Y2=0
cc_526 N_A_934_357#_M1037_g N_A_1273_393#_M1001_g 0.0646955f $X=6.52 $Y=0.805
+ $X2=0 $Y2=0
cc_527 N_A_934_357#_c_696_n N_A_1273_393#_M1001_g 0.00541313f $X=9.215 $Y=1.665
+ $X2=0 $Y2=0
cc_528 N_A_934_357#_c_703_n N_A_1273_393#_c_868_n 0.0277336f $X=9.53 $Y=1.375
+ $X2=0 $Y2=0
cc_529 N_A_934_357#_c_696_n N_A_1273_393#_M1018_g 0.00233565f $X=9.215 $Y=1.665
+ $X2=0 $Y2=0
cc_530 N_A_934_357#_c_699_n N_A_1273_393#_M1018_g 0.00114441f $X=9.36 $Y=1.665
+ $X2=0 $Y2=0
cc_531 N_A_934_357#_c_696_n N_A_1273_393#_c_894_n 0.00938854f $X=9.215 $Y=1.665
+ $X2=0 $Y2=0
cc_532 N_A_934_357#_c_696_n N_A_1273_393#_c_879_n 0.00150641f $X=9.215 $Y=1.665
+ $X2=0 $Y2=0
cc_533 N_A_934_357#_c_696_n N_A_1273_393#_c_870_n 0.0364201f $X=9.215 $Y=1.665
+ $X2=0 $Y2=0
cc_534 N_A_934_357#_c_699_n N_A_1273_393#_c_870_n 0.00134414f $X=9.36 $Y=1.665
+ $X2=0 $Y2=0
cc_535 N_A_934_357#_c_700_n N_A_1273_393#_c_870_n 0.0245638f $X=9.36 $Y=1.665
+ $X2=0 $Y2=0
cc_536 N_A_934_357#_c_702_n N_A_1273_393#_c_870_n 3.53194e-19 $X=9.53 $Y=1.54
+ $X2=0 $Y2=0
cc_537 N_A_934_357#_M1009_g N_A_1273_393#_c_882_n 0.00226576f $X=5.62 $Y=2.525
+ $X2=0 $Y2=0
cc_538 N_A_934_357#_c_689_n N_A_1273_393#_c_882_n 0.0072092f $X=6.22 $Y=1.65
+ $X2=0 $Y2=0
cc_539 N_A_934_357#_c_696_n N_A_1273_393#_c_882_n 0.00267908f $X=9.215 $Y=1.665
+ $X2=0 $Y2=0
cc_540 N_A_934_357#_c_696_n N_A_1273_393#_c_883_n 0.0226264f $X=9.215 $Y=1.665
+ $X2=0 $Y2=0
cc_541 N_A_934_357#_c_696_n N_A_1273_393#_c_871_n 0.0088021f $X=9.215 $Y=1.665
+ $X2=0 $Y2=0
cc_542 N_A_934_357#_c_696_n N_A_1273_393#_c_884_n 0.00475473f $X=9.215 $Y=1.665
+ $X2=0 $Y2=0
cc_543 N_A_934_357#_c_696_n N_A_1273_393#_c_872_n 0.00594361f $X=9.215 $Y=1.665
+ $X2=0 $Y2=0
cc_544 N_A_934_357#_c_696_n N_A_1273_393#_c_873_n 0.00633316f $X=9.215 $Y=1.665
+ $X2=0 $Y2=0
cc_545 N_A_934_357#_c_699_n N_A_1273_393#_c_873_n 7.49209e-19 $X=9.36 $Y=1.665
+ $X2=0 $Y2=0
cc_546 N_A_934_357#_c_700_n N_A_1273_393#_c_873_n 0.00472342f $X=9.36 $Y=1.665
+ $X2=0 $Y2=0
cc_547 N_A_934_357#_c_702_n N_A_1273_393#_c_873_n 0.0377904f $X=9.53 $Y=1.54
+ $X2=0 $Y2=0
cc_548 N_A_934_357#_c_696_n N_A_1139_463#_M1019_g 0.00258175f $X=9.215 $Y=1.665
+ $X2=0 $Y2=0
cc_549 N_A_934_357#_M1009_g N_A_1139_463#_c_1017_n 0.00417666f $X=5.62 $Y=2.525
+ $X2=0 $Y2=0
cc_550 N_A_934_357#_M1037_g N_A_1139_463#_c_1010_n 0.0196453f $X=6.52 $Y=0.805
+ $X2=0 $Y2=0
cc_551 N_A_934_357#_M1009_g N_A_1139_463#_c_1011_n 4.35326e-19 $X=5.62 $Y=2.525
+ $X2=0 $Y2=0
cc_552 N_A_934_357#_c_689_n N_A_1139_463#_c_1011_n 0.00876203f $X=6.22 $Y=1.65
+ $X2=0 $Y2=0
cc_553 N_A_934_357#_c_696_n N_A_1139_463#_c_1011_n 0.025556f $X=9.215 $Y=1.665
+ $X2=0 $Y2=0
cc_554 N_A_934_357#_c_689_n N_A_1139_463#_c_1012_n 0.00368728f $X=6.22 $Y=1.65
+ $X2=0 $Y2=0
cc_555 N_A_934_357#_M1037_g N_A_1139_463#_c_1012_n 0.00585587f $X=6.52 $Y=0.805
+ $X2=0 $Y2=0
cc_556 N_A_934_357#_c_696_n N_A_1139_463#_c_1012_n 0.0230002f $X=9.215 $Y=1.665
+ $X2=0 $Y2=0
cc_557 N_A_934_357#_c_689_n N_A_1139_463#_c_1013_n 0.00950994f $X=6.22 $Y=1.65
+ $X2=0 $Y2=0
cc_558 N_A_934_357#_M1037_g N_A_1139_463#_c_1013_n 4.02994e-19 $X=6.52 $Y=0.805
+ $X2=0 $Y2=0
cc_559 N_A_934_357#_c_696_n N_A_1139_463#_c_1013_n 0.00444405f $X=9.215 $Y=1.665
+ $X2=0 $Y2=0
cc_560 N_A_934_357#_c_696_n N_A_1139_463#_c_1014_n 0.0189445f $X=9.215 $Y=1.665
+ $X2=0 $Y2=0
cc_561 N_A_934_357#_c_696_n N_A_1139_463#_c_1015_n 0.00268026f $X=9.215 $Y=1.665
+ $X2=0 $Y2=0
cc_562 N_A_934_357#_c_696_n N_ASYNC_M1034_g 0.00157252f $X=9.215 $Y=1.665 $X2=0
+ $Y2=0
cc_563 N_A_934_357#_c_696_n N_ASYNC_c_1101_n 0.0156503f $X=9.215 $Y=1.665 $X2=0
+ $Y2=0
cc_564 N_A_934_357#_c_691_n N_ASYNC_c_1108_n 0.00393745f $X=10.06 $Y=1.63 $X2=0
+ $Y2=0
cc_565 N_A_934_357#_M1007_g N_ASYNC_c_1108_n 0.0139725f $X=10.135 $Y=2.465 $X2=0
+ $Y2=0
cc_566 N_A_934_357#_c_696_n N_ASYNC_c_1108_n 0.0854784f $X=9.215 $Y=1.665 $X2=0
+ $Y2=0
cc_567 N_A_934_357#_c_699_n N_ASYNC_c_1108_n 0.0257814f $X=9.36 $Y=1.665 $X2=0
+ $Y2=0
cc_568 N_A_934_357#_c_700_n N_ASYNC_c_1108_n 0.00943217f $X=9.36 $Y=1.665 $X2=0
+ $Y2=0
cc_569 N_A_934_357#_c_696_n N_ASYNC_c_1121_n 0.0231704f $X=9.215 $Y=1.665 $X2=0
+ $Y2=0
cc_570 N_A_934_357#_c_696_n N_ASYNC_c_1109_n 0.00665253f $X=9.215 $Y=1.665 $X2=0
+ $Y2=0
cc_571 N_A_934_357#_c_696_n N_ASYNC_c_1102_n 0.00273582f $X=9.215 $Y=1.665 $X2=0
+ $Y2=0
cc_572 N_A_934_357#_c_708_n N_A_761_357#_M1029_g 0.00116223f $X=4.81 $Y=1.93
+ $X2=0 $Y2=0
cc_573 N_A_934_357#_c_694_n N_A_761_357#_M1029_g 0.00113087f $X=4.725 $Y=1.735
+ $X2=0 $Y2=0
cc_574 N_A_934_357#_c_692_n N_A_761_357#_c_1233_n 0.00925585f $X=5.01 $Y=0.43
+ $X2=0 $Y2=0
cc_575 N_A_934_357#_c_693_n N_A_761_357#_c_1233_n 0.00264333f $X=5.115 $Y=1.55
+ $X2=0 $Y2=0
cc_576 N_A_934_357#_c_695_n N_A_761_357#_c_1233_n 0.00348785f $X=5.022 $Y=1.045
+ $X2=0 $Y2=0
cc_577 N_A_934_357#_M1009_g N_A_761_357#_c_1234_n 0.0213561f $X=5.62 $Y=2.525
+ $X2=0 $Y2=0
cc_578 N_A_934_357#_c_708_n N_A_761_357#_c_1234_n 0.0215836f $X=4.81 $Y=1.93
+ $X2=0 $Y2=0
cc_579 N_A_934_357#_c_694_n N_A_761_357#_c_1234_n 0.0191445f $X=4.725 $Y=1.735
+ $X2=0 $Y2=0
cc_580 N_A_934_357#_c_701_n N_A_761_357#_c_1234_n 0.0213699f $X=5.555 $Y=1.65
+ $X2=0 $Y2=0
cc_581 N_A_934_357#_c_693_n N_A_761_357#_c_1235_n 0.00543494f $X=5.115 $Y=1.55
+ $X2=0 $Y2=0
cc_582 N_A_934_357#_c_696_n N_A_761_357#_c_1235_n 9.99416e-19 $X=9.215 $Y=1.665
+ $X2=0 $Y2=0
cc_583 N_A_934_357#_c_697_n N_A_761_357#_c_1235_n 0.00408074f $X=5.665 $Y=1.665
+ $X2=0 $Y2=0
cc_584 N_A_934_357#_c_698_n N_A_761_357#_c_1235_n 0.0089927f $X=5.52 $Y=1.665
+ $X2=0 $Y2=0
cc_585 N_A_934_357#_c_701_n N_A_761_357#_c_1235_n 0.0332091f $X=5.555 $Y=1.65
+ $X2=0 $Y2=0
cc_586 N_A_934_357#_M1009_g N_A_761_357#_c_1246_n 0.0102957f $X=5.62 $Y=2.525
+ $X2=0 $Y2=0
cc_587 N_A_934_357#_M1037_g N_A_761_357#_M1032_g 0.0162801f $X=6.52 $Y=0.805
+ $X2=0 $Y2=0
cc_588 N_A_934_357#_c_692_n N_A_761_357#_M1032_g 0.00501062f $X=5.01 $Y=0.43
+ $X2=0 $Y2=0
cc_589 N_A_934_357#_c_695_n N_A_761_357#_M1032_g 0.00201544f $X=5.022 $Y=1.045
+ $X2=0 $Y2=0
cc_590 N_A_934_357#_M1009_g N_A_761_357#_M1017_g 0.0140822f $X=5.62 $Y=2.525
+ $X2=0 $Y2=0
cc_591 N_A_934_357#_c_689_n N_A_761_357#_M1017_g 0.00404223f $X=6.22 $Y=1.65
+ $X2=0 $Y2=0
cc_592 N_A_934_357#_c_696_n N_A_761_357#_M1017_g 0.00107473f $X=9.215 $Y=1.665
+ $X2=0 $Y2=0
cc_593 N_A_934_357#_M1037_g N_A_761_357#_c_1237_n 0.0103003f $X=6.52 $Y=0.805
+ $X2=0 $Y2=0
cc_594 N_A_934_357#_c_703_n N_A_761_357#_c_1237_n 0.00907339f $X=9.53 $Y=1.375
+ $X2=0 $Y2=0
cc_595 N_A_934_357#_M1007_g N_A_761_357#_M1042_g 0.0143828f $X=10.135 $Y=2.465
+ $X2=0 $Y2=0
cc_596 N_A_934_357#_c_700_n N_A_761_357#_M1042_g 0.00345817f $X=9.36 $Y=1.665
+ $X2=0 $Y2=0
cc_597 N_A_934_357#_c_702_n N_A_761_357#_M1042_g 0.00989034f $X=9.53 $Y=1.54
+ $X2=0 $Y2=0
cc_598 N_A_934_357#_c_691_n N_A_761_357#_M1021_g 0.00257732f $X=10.06 $Y=1.63
+ $X2=0 $Y2=0
cc_599 N_A_934_357#_c_703_n N_A_761_357#_M1021_g 0.00831166f $X=9.53 $Y=1.375
+ $X2=0 $Y2=0
cc_600 N_A_934_357#_c_694_n N_A_761_357#_c_1253_n 0.00888568f $X=4.725 $Y=1.735
+ $X2=0 $Y2=0
cc_601 N_A_934_357#_c_692_n N_A_761_357#_c_1270_n 0.00905117f $X=5.01 $Y=0.43
+ $X2=0 $Y2=0
cc_602 N_A_934_357#_c_693_n N_A_761_357#_c_1240_n 0.00612248f $X=5.115 $Y=1.55
+ $X2=0 $Y2=0
cc_603 N_A_934_357#_c_695_n N_A_761_357#_c_1240_n 0.00213618f $X=5.022 $Y=1.045
+ $X2=0 $Y2=0
cc_604 N_A_934_357#_c_694_n N_A_761_357#_c_1241_n 0.00447149f $X=4.725 $Y=1.735
+ $X2=0 $Y2=0
cc_605 N_A_934_357#_c_693_n N_A_761_357#_c_1242_n 0.0228436f $X=5.115 $Y=1.55
+ $X2=0 $Y2=0
cc_606 N_A_934_357#_c_694_n N_A_761_357#_c_1242_n 0.0100983f $X=4.725 $Y=1.735
+ $X2=0 $Y2=0
cc_607 N_A_934_357#_c_693_n N_A_761_357#_c_1243_n 0.0161313f $X=5.115 $Y=1.55
+ $X2=0 $Y2=0
cc_608 N_A_934_357#_c_694_n N_A_761_357#_c_1243_n 0.00681598f $X=4.725 $Y=1.735
+ $X2=0 $Y2=0
cc_609 N_A_934_357#_c_695_n N_A_761_357#_c_1243_n 0.00349887f $X=5.022 $Y=1.045
+ $X2=0 $Y2=0
cc_610 N_A_934_357#_M1007_g N_A_2083_65#_M1008_g 0.0362531f $X=10.135 $Y=2.465
+ $X2=0 $Y2=0
cc_611 N_A_934_357#_M1007_g N_A_2083_65#_c_1434_n 6.90596e-19 $X=10.135 $Y=2.465
+ $X2=0 $Y2=0
cc_612 N_A_934_357#_M1007_g N_A_2083_65#_c_1443_n 5.01056e-19 $X=10.135 $Y=2.465
+ $X2=0 $Y2=0
cc_613 N_A_934_357#_M1007_g N_A_2083_65#_c_1435_n 0.00122016f $X=10.135 $Y=2.465
+ $X2=0 $Y2=0
cc_614 N_A_934_357#_M1007_g N_A_2083_65#_c_1436_n 0.0170651f $X=10.135 $Y=2.465
+ $X2=0 $Y2=0
cc_615 N_A_934_357#_c_691_n N_A_2083_65#_c_1429_n 0.0170651f $X=10.06 $Y=1.63
+ $X2=0 $Y2=0
cc_616 N_A_934_357#_c_703_n N_A_1903_125#_c_1588_n 0.0146966f $X=9.53 $Y=1.375
+ $X2=0 $Y2=0
cc_617 N_A_934_357#_c_691_n N_A_1903_125#_c_1597_n 0.00603263f $X=10.06 $Y=1.63
+ $X2=0 $Y2=0
cc_618 N_A_934_357#_c_700_n N_A_1903_125#_c_1597_n 0.00717041f $X=9.36 $Y=1.665
+ $X2=0 $Y2=0
cc_619 N_A_934_357#_c_702_n N_A_1903_125#_c_1597_n 0.00208313f $X=9.53 $Y=1.54
+ $X2=0 $Y2=0
cc_620 N_A_934_357#_c_703_n N_A_1903_125#_c_1597_n 0.00917886f $X=9.53 $Y=1.375
+ $X2=0 $Y2=0
cc_621 N_A_934_357#_c_691_n N_A_1903_125#_c_1594_n 0.00483908f $X=10.06 $Y=1.63
+ $X2=0 $Y2=0
cc_622 N_A_934_357#_M1007_g N_A_1903_125#_c_1594_n 0.0126603f $X=10.135 $Y=2.465
+ $X2=0 $Y2=0
cc_623 N_A_934_357#_c_700_n N_A_1903_125#_c_1594_n 0.00255235f $X=9.36 $Y=1.665
+ $X2=0 $Y2=0
cc_624 N_A_934_357#_c_691_n N_A_1903_125#_c_1589_n 0.0147182f $X=10.06 $Y=1.63
+ $X2=0 $Y2=0
cc_625 N_A_934_357#_M1007_g N_A_1903_125#_c_1589_n 0.00923562f $X=10.135
+ $Y=2.465 $X2=0 $Y2=0
cc_626 N_A_934_357#_c_699_n N_A_1903_125#_c_1589_n 0.00102978f $X=9.36 $Y=1.665
+ $X2=0 $Y2=0
cc_627 N_A_934_357#_c_700_n N_A_1903_125#_c_1589_n 0.0286472f $X=9.36 $Y=1.665
+ $X2=0 $Y2=0
cc_628 N_A_934_357#_c_702_n N_A_1903_125#_c_1589_n 0.00124625f $X=9.53 $Y=1.54
+ $X2=0 $Y2=0
cc_629 N_A_934_357#_c_703_n N_A_1903_125#_c_1589_n 0.00362326f $X=9.53 $Y=1.375
+ $X2=0 $Y2=0
cc_630 N_A_934_357#_c_691_n N_A_1903_125#_c_1592_n 0.00388433f $X=10.06 $Y=1.63
+ $X2=0 $Y2=0
cc_631 N_A_934_357#_c_708_n N_VPWR_c_1778_n 0.0373084f $X=4.81 $Y=1.93 $X2=0
+ $Y2=0
cc_632 N_A_934_357#_c_696_n N_VPWR_c_1779_n 8.1649e-19 $X=9.215 $Y=1.665 $X2=0
+ $Y2=0
cc_633 N_A_934_357#_c_696_n N_VPWR_c_1781_n 0.00259861f $X=9.215 $Y=1.665 $X2=0
+ $Y2=0
cc_634 N_A_934_357#_c_708_n N_VPWR_c_1792_n 0.0204296f $X=4.81 $Y=1.93 $X2=0
+ $Y2=0
cc_635 N_A_934_357#_M1007_g N_VPWR_c_1799_n 0.00399858f $X=10.135 $Y=2.465 $X2=0
+ $Y2=0
cc_636 N_A_934_357#_M1009_g N_VPWR_c_1775_n 9.39239e-19 $X=5.62 $Y=2.525 $X2=0
+ $Y2=0
cc_637 N_A_934_357#_M1007_g N_VPWR_c_1775_n 0.0046122f $X=10.135 $Y=2.465 $X2=0
+ $Y2=0
cc_638 N_A_934_357#_c_708_n N_VPWR_c_1775_n 0.011724f $X=4.81 $Y=1.93 $X2=0
+ $Y2=0
cc_639 N_A_934_357#_M1009_g N_A_636_531#_c_1971_n 0.00190702f $X=5.62 $Y=2.525
+ $X2=0 $Y2=0
cc_640 N_A_934_357#_c_708_n N_A_636_531#_c_1971_n 0.0348782f $X=4.81 $Y=1.93
+ $X2=0 $Y2=0
cc_641 N_A_934_357#_M1009_g N_A_636_531#_c_1972_n 0.0147177f $X=5.62 $Y=2.525
+ $X2=0 $Y2=0
cc_642 N_A_934_357#_c_689_n N_A_636_531#_c_1972_n 0.00354579f $X=6.22 $Y=1.65
+ $X2=0 $Y2=0
cc_643 N_A_934_357#_c_696_n N_A_636_531#_c_1972_n 0.00682551f $X=9.215 $Y=1.665
+ $X2=0 $Y2=0
cc_644 N_A_934_357#_c_697_n N_A_636_531#_c_1972_n 9.24148e-19 $X=5.665 $Y=1.665
+ $X2=0 $Y2=0
cc_645 N_A_934_357#_c_698_n N_A_636_531#_c_1972_n 0.0129062f $X=5.52 $Y=1.665
+ $X2=0 $Y2=0
cc_646 N_A_934_357#_c_701_n N_A_636_531#_c_1972_n 0.00215202f $X=5.555 $Y=1.65
+ $X2=0 $Y2=0
cc_647 N_A_934_357#_c_708_n N_A_636_531#_c_1973_n 0.0128704f $X=4.81 $Y=1.93
+ $X2=0 $Y2=0
cc_648 N_A_934_357#_c_697_n N_A_636_531#_c_1973_n 7.27918e-19 $X=5.665 $Y=1.665
+ $X2=0 $Y2=0
cc_649 N_A_934_357#_c_698_n N_A_636_531#_c_1973_n 0.020133f $X=5.52 $Y=1.665
+ $X2=0 $Y2=0
cc_650 N_A_934_357#_c_701_n N_A_636_531#_c_1973_n 0.00231301f $X=5.555 $Y=1.65
+ $X2=0 $Y2=0
cc_651 N_A_934_357#_M1009_g N_A_636_531#_c_1964_n 0.00490161f $X=5.62 $Y=2.525
+ $X2=0 $Y2=0
cc_652 N_A_934_357#_c_689_n N_A_636_531#_c_1964_n 0.0121281f $X=6.22 $Y=1.65
+ $X2=0 $Y2=0
cc_653 N_A_934_357#_M1037_g N_A_636_531#_c_1964_n 9.10352e-19 $X=6.52 $Y=0.805
+ $X2=0 $Y2=0
cc_654 N_A_934_357#_c_695_n N_A_636_531#_c_1964_n 0.013198f $X=5.022 $Y=1.045
+ $X2=0 $Y2=0
cc_655 N_A_934_357#_c_696_n N_A_636_531#_c_1964_n 0.015671f $X=9.215 $Y=1.665
+ $X2=0 $Y2=0
cc_656 N_A_934_357#_c_697_n N_A_636_531#_c_1964_n 6.13261e-19 $X=5.665 $Y=1.665
+ $X2=0 $Y2=0
cc_657 N_A_934_357#_c_698_n N_A_636_531#_c_1964_n 0.0243745f $X=5.52 $Y=1.665
+ $X2=0 $Y2=0
cc_658 N_A_934_357#_c_701_n N_A_636_531#_c_1964_n 0.00410885f $X=5.555 $Y=1.65
+ $X2=0 $Y2=0
cc_659 N_A_934_357#_c_692_n N_A_636_531#_c_1965_n 0.0256632f $X=5.01 $Y=0.43
+ $X2=0 $Y2=0
cc_660 N_A_934_357#_c_692_n N_A_636_531#_c_1968_n 0.00267978f $X=5.01 $Y=0.43
+ $X2=0 $Y2=0
cc_661 N_A_934_357#_M1037_g N_A_636_531#_c_1969_n 0.00248996f $X=6.52 $Y=0.805
+ $X2=0 $Y2=0
cc_662 N_A_934_357#_c_692_n N_A_636_531#_c_1969_n 0.0419128f $X=5.01 $Y=0.43
+ $X2=0 $Y2=0
cc_663 N_A_934_357#_c_696_n N_A_636_531#_c_1969_n 0.00635375f $X=9.215 $Y=1.665
+ $X2=0 $Y2=0
cc_664 N_A_934_357#_c_697_n N_A_636_531#_c_1969_n 0.00604343f $X=5.665 $Y=1.665
+ $X2=0 $Y2=0
cc_665 N_A_934_357#_c_698_n N_A_636_531#_c_1969_n 0.00689343f $X=5.52 $Y=1.665
+ $X2=0 $Y2=0
cc_666 N_A_934_357#_c_701_n N_A_636_531#_c_1969_n 0.00167557f $X=5.555 $Y=1.65
+ $X2=0 $Y2=0
cc_667 N_A_934_357#_c_692_n N_VGND_c_2172_n 0.0155501f $X=5.01 $Y=0.43 $X2=0
+ $Y2=0
cc_668 N_A_934_357#_c_696_n N_VGND_c_2173_n 0.00107779f $X=9.215 $Y=1.665 $X2=0
+ $Y2=0
cc_669 N_A_934_357#_c_696_n N_VGND_c_2174_n 0.00133308f $X=9.215 $Y=1.665 $X2=0
+ $Y2=0
cc_670 N_A_934_357#_c_692_n N_VGND_c_2180_n 0.0214436f $X=5.01 $Y=0.43 $X2=0
+ $Y2=0
cc_671 N_A_934_357#_M1043_d N_VGND_c_2190_n 0.00140449f $X=4.87 $Y=0.235 $X2=0
+ $Y2=0
cc_672 N_A_934_357#_M1037_g N_VGND_c_2190_n 9.39239e-19 $X=6.52 $Y=0.805 $X2=0
+ $Y2=0
cc_673 N_A_934_357#_c_692_n N_VGND_c_2190_n 0.00419796f $X=5.01 $Y=0.43 $X2=0
+ $Y2=0
cc_674 N_A_934_357#_c_703_n N_VGND_c_2190_n 9.49986e-19 $X=9.53 $Y=1.375 $X2=0
+ $Y2=0
cc_675 N_A_1273_393#_M1001_g N_A_1139_463#_M1038_g 0.0188657f $X=6.88 $Y=0.805
+ $X2=0 $Y2=0
cc_676 N_A_1273_393#_c_871_n N_A_1139_463#_M1038_g 0.00174543f $X=8.34 $Y=0.885
+ $X2=0 $Y2=0
cc_677 N_A_1273_393#_M1001_g N_A_1139_463#_M1019_g 0.00915307f $X=6.88 $Y=0.805
+ $X2=0 $Y2=0
cc_678 N_A_1273_393#_c_877_n N_A_1139_463#_M1019_g 0.00609153f $X=7.215 $Y=2.33
+ $X2=0 $Y2=0
cc_679 N_A_1273_393#_c_894_n N_A_1139_463#_M1019_g 0.00952625f $X=8.22 $Y=2.415
+ $X2=0 $Y2=0
cc_680 N_A_1273_393#_c_878_n N_A_1139_463#_M1019_g 0.00625608f $X=7.38 $Y=2.415
+ $X2=0 $Y2=0
cc_681 N_A_1273_393#_c_883_n N_A_1139_463#_M1019_g 0.00422398f $X=7.215 $Y=2.05
+ $X2=0 $Y2=0
cc_682 N_A_1273_393#_M1033_g N_A_1139_463#_c_1017_n 0.00709057f $X=6.44 $Y=2.525
+ $X2=0 $Y2=0
cc_683 N_A_1273_393#_M1001_g N_A_1139_463#_c_1010_n 0.00270661f $X=6.88 $Y=0.805
+ $X2=0 $Y2=0
cc_684 N_A_1273_393#_M1033_g N_A_1139_463#_c_1011_n 0.00801673f $X=6.44 $Y=2.525
+ $X2=0 $Y2=0
cc_685 N_A_1273_393#_M1001_g N_A_1139_463#_c_1011_n 0.00372318f $X=6.88 $Y=0.805
+ $X2=0 $Y2=0
cc_686 N_A_1273_393#_c_877_n N_A_1139_463#_c_1011_n 0.00484066f $X=7.215 $Y=2.33
+ $X2=0 $Y2=0
cc_687 N_A_1273_393#_c_882_n N_A_1139_463#_c_1011_n 0.00614067f $X=6.745 $Y=1.95
+ $X2=0 $Y2=0
cc_688 N_A_1273_393#_c_883_n N_A_1139_463#_c_1011_n 0.0232652f $X=7.215 $Y=2.05
+ $X2=0 $Y2=0
cc_689 N_A_1273_393#_M1001_g N_A_1139_463#_c_1012_n 0.0145201f $X=6.88 $Y=0.805
+ $X2=0 $Y2=0
cc_690 N_A_1273_393#_c_882_n N_A_1139_463#_c_1012_n 0.0020797f $X=6.745 $Y=1.95
+ $X2=0 $Y2=0
cc_691 N_A_1273_393#_c_883_n N_A_1139_463#_c_1012_n 0.0192669f $X=7.215 $Y=2.05
+ $X2=0 $Y2=0
cc_692 N_A_1273_393#_c_882_n N_A_1139_463#_c_1013_n 5.54033e-19 $X=6.745 $Y=1.95
+ $X2=0 $Y2=0
cc_693 N_A_1273_393#_M1001_g N_A_1139_463#_c_1014_n 0.00162701f $X=6.88 $Y=0.805
+ $X2=0 $Y2=0
cc_694 N_A_1273_393#_c_894_n N_A_1139_463#_c_1014_n 0.00140716f $X=8.22 $Y=2.415
+ $X2=0 $Y2=0
cc_695 N_A_1273_393#_c_883_n N_A_1139_463#_c_1014_n 0.0112419f $X=7.215 $Y=2.05
+ $X2=0 $Y2=0
cc_696 N_A_1273_393#_M1001_g N_A_1139_463#_c_1015_n 0.0207485f $X=6.88 $Y=0.805
+ $X2=0 $Y2=0
cc_697 N_A_1273_393#_c_883_n N_A_1139_463#_c_1015_n 0.00122759f $X=7.215 $Y=2.05
+ $X2=0 $Y2=0
cc_698 N_A_1273_393#_c_869_n N_ASYNC_M1010_g 0.00500796f $X=8.34 $Y=1.375 $X2=0
+ $Y2=0
cc_699 N_A_1273_393#_c_871_n N_ASYNC_M1010_g 0.0161876f $X=8.34 $Y=0.885 $X2=0
+ $Y2=0
cc_700 N_A_1273_393#_c_877_n N_ASYNC_M1034_g 8.06571e-19 $X=7.215 $Y=2.33 $X2=0
+ $Y2=0
cc_701 N_A_1273_393#_c_894_n N_ASYNC_M1034_g 0.0100574f $X=8.22 $Y=2.415 $X2=0
+ $Y2=0
cc_702 N_A_1273_393#_c_878_n N_ASYNC_M1034_g 7.91781e-19 $X=7.38 $Y=2.415 $X2=0
+ $Y2=0
cc_703 N_A_1273_393#_c_879_n N_ASYNC_M1034_g 0.00183335f $X=8.345 $Y=2.01 $X2=0
+ $Y2=0
cc_704 N_A_1273_393#_c_884_n N_ASYNC_M1034_g 0.00341054f $X=8.345 $Y=1.885 $X2=0
+ $Y2=0
cc_705 N_A_1273_393#_c_885_n N_ASYNC_M1034_g 4.77545e-19 $X=8.345 $Y=2.415 $X2=0
+ $Y2=0
cc_706 N_A_1273_393#_c_894_n N_ASYNC_c_1101_n 3.60586e-19 $X=8.22 $Y=2.415 $X2=0
+ $Y2=0
cc_707 N_A_1273_393#_c_871_n N_ASYNC_c_1101_n 0.0135129f $X=8.34 $Y=0.885 $X2=0
+ $Y2=0
cc_708 N_A_1273_393#_c_872_n N_ASYNC_c_1101_n 0.0250074f $X=8.34 $Y=1.54 $X2=0
+ $Y2=0
cc_709 N_A_1273_393#_c_873_n N_ASYNC_c_1101_n 2.25027e-19 $X=9.05 $Y=1.54 $X2=0
+ $Y2=0
cc_710 N_A_1273_393#_M1034_d N_ASYNC_c_1108_n 9.51227e-19 $X=8.165 $Y=1.865
+ $X2=0 $Y2=0
cc_711 N_A_1273_393#_M1018_g N_ASYNC_c_1108_n 0.0076249f $X=9.08 $Y=2.285 $X2=0
+ $Y2=0
cc_712 N_A_1273_393#_c_894_n N_ASYNC_c_1108_n 0.00572645f $X=8.22 $Y=2.415 $X2=0
+ $Y2=0
cc_713 N_A_1273_393#_c_879_n N_ASYNC_c_1108_n 0.00594611f $X=8.345 $Y=2.01 $X2=0
+ $Y2=0
cc_714 N_A_1273_393#_c_880_n N_ASYNC_c_1108_n 0.0181179f $X=8.305 $Y=2.05 $X2=0
+ $Y2=0
cc_715 N_A_1273_393#_c_870_n N_ASYNC_c_1108_n 0.00272101f $X=8.9 $Y=1.54 $X2=0
+ $Y2=0
cc_716 N_A_1273_393#_c_877_n N_ASYNC_c_1121_n 2.15063e-19 $X=7.215 $Y=2.33 $X2=0
+ $Y2=0
cc_717 N_A_1273_393#_c_894_n N_ASYNC_c_1121_n 0.00283116f $X=8.22 $Y=2.415 $X2=0
+ $Y2=0
cc_718 N_A_1273_393#_c_879_n N_ASYNC_c_1121_n 0.00115685f $X=8.345 $Y=2.01 $X2=0
+ $Y2=0
cc_719 N_A_1273_393#_c_880_n N_ASYNC_c_1121_n 0.00115685f $X=8.305 $Y=2.05 $X2=0
+ $Y2=0
cc_720 N_A_1273_393#_c_883_n N_ASYNC_c_1121_n 0.00132026f $X=7.215 $Y=2.05 $X2=0
+ $Y2=0
cc_721 N_A_1273_393#_c_877_n N_ASYNC_c_1109_n 0.00123834f $X=7.215 $Y=2.33 $X2=0
+ $Y2=0
cc_722 N_A_1273_393#_c_894_n N_ASYNC_c_1109_n 0.0155118f $X=8.22 $Y=2.415 $X2=0
+ $Y2=0
cc_723 N_A_1273_393#_c_879_n N_ASYNC_c_1109_n 0.0103082f $X=8.345 $Y=2.01 $X2=0
+ $Y2=0
cc_724 N_A_1273_393#_c_883_n N_ASYNC_c_1109_n 0.008879f $X=7.215 $Y=2.05 $X2=0
+ $Y2=0
cc_725 N_A_1273_393#_c_884_n N_ASYNC_c_1109_n 0.0106461f $X=8.345 $Y=1.885 $X2=0
+ $Y2=0
cc_726 N_A_1273_393#_c_894_n N_ASYNC_c_1102_n 7.08417e-19 $X=8.22 $Y=2.415 $X2=0
+ $Y2=0
cc_727 N_A_1273_393#_c_871_n N_ASYNC_c_1102_n 0.0054841f $X=8.34 $Y=0.885 $X2=0
+ $Y2=0
cc_728 N_A_1273_393#_c_872_n N_ASYNC_c_1102_n 0.00385396f $X=8.34 $Y=1.54 $X2=0
+ $Y2=0
cc_729 N_A_1273_393#_c_873_n N_ASYNC_c_1102_n 0.00520091f $X=9.05 $Y=1.54 $X2=0
+ $Y2=0
cc_730 N_A_1273_393#_M1033_g N_A_761_357#_M1017_g 0.0357064f $X=6.44 $Y=2.525
+ $X2=0 $Y2=0
cc_731 N_A_1273_393#_M1001_g N_A_761_357#_c_1237_n 0.0104164f $X=6.88 $Y=0.805
+ $X2=0 $Y2=0
cc_732 N_A_1273_393#_c_868_n N_A_761_357#_c_1237_n 0.00907339f $X=9.05 $Y=1.375
+ $X2=0 $Y2=0
cc_733 N_A_1273_393#_c_871_n N_A_761_357#_c_1237_n 0.0107219f $X=8.34 $Y=0.885
+ $X2=0 $Y2=0
cc_734 N_A_1273_393#_M1033_g N_A_761_357#_c_1249_n 0.0102955f $X=6.44 $Y=2.525
+ $X2=0 $Y2=0
cc_735 N_A_1273_393#_M1018_g N_A_761_357#_c_1249_n 0.00894529f $X=9.08 $Y=2.285
+ $X2=0 $Y2=0
cc_736 N_A_1273_393#_c_894_n N_A_761_357#_c_1249_n 0.0047676f $X=8.22 $Y=2.415
+ $X2=0 $Y2=0
cc_737 N_A_1273_393#_c_878_n N_A_761_357#_c_1249_n 0.00612696f $X=7.38 $Y=2.415
+ $X2=0 $Y2=0
cc_738 N_A_1273_393#_c_885_n N_A_761_357#_c_1249_n 0.00492264f $X=8.345 $Y=2.415
+ $X2=0 $Y2=0
cc_739 N_A_1273_393#_M1018_g N_A_761_357#_M1042_g 0.0290071f $X=9.08 $Y=2.285
+ $X2=0 $Y2=0
cc_740 N_A_1273_393#_M1018_g N_A_1903_125#_c_1594_n 0.00250624f $X=9.08 $Y=2.285
+ $X2=0 $Y2=0
cc_741 N_A_1273_393#_c_894_n N_VPWR_M1019_d 0.0108204f $X=8.22 $Y=2.415 $X2=0
+ $Y2=0
cc_742 N_A_1273_393#_M1033_g N_VPWR_c_1779_n 0.00593231f $X=6.44 $Y=2.525 $X2=0
+ $Y2=0
cc_743 N_A_1273_393#_c_877_n N_VPWR_c_1779_n 0.00227737f $X=7.215 $Y=2.33 $X2=0
+ $Y2=0
cc_744 N_A_1273_393#_c_878_n N_VPWR_c_1779_n 0.0268338f $X=7.38 $Y=2.415 $X2=0
+ $Y2=0
cc_745 N_A_1273_393#_c_882_n N_VPWR_c_1779_n 0.00224227f $X=6.745 $Y=1.95 $X2=0
+ $Y2=0
cc_746 N_A_1273_393#_c_883_n N_VPWR_c_1779_n 0.0187004f $X=7.215 $Y=2.05 $X2=0
+ $Y2=0
cc_747 N_A_1273_393#_c_894_n N_VPWR_c_1780_n 0.0244147f $X=8.22 $Y=2.415 $X2=0
+ $Y2=0
cc_748 N_A_1273_393#_c_878_n N_VPWR_c_1780_n 0.00295942f $X=7.38 $Y=2.415 $X2=0
+ $Y2=0
cc_749 N_A_1273_393#_c_885_n N_VPWR_c_1780_n 0.00175107f $X=8.345 $Y=2.415 $X2=0
+ $Y2=0
cc_750 N_A_1273_393#_M1018_g N_VPWR_c_1781_n 0.0242972f $X=9.08 $Y=2.285 $X2=0
+ $Y2=0
cc_751 N_A_1273_393#_c_879_n N_VPWR_c_1781_n 0.0536278f $X=8.345 $Y=2.01 $X2=0
+ $Y2=0
cc_752 N_A_1273_393#_c_870_n N_VPWR_c_1781_n 0.0193293f $X=8.9 $Y=1.54 $X2=0
+ $Y2=0
cc_753 N_A_1273_393#_c_873_n N_VPWR_c_1781_n 0.00465478f $X=9.05 $Y=1.54 $X2=0
+ $Y2=0
cc_754 N_A_1273_393#_c_878_n N_VPWR_c_1794_n 0.00704253f $X=7.38 $Y=2.415 $X2=0
+ $Y2=0
cc_755 N_A_1273_393#_c_885_n N_VPWR_c_1798_n 0.00534275f $X=8.345 $Y=2.415 $X2=0
+ $Y2=0
cc_756 N_A_1273_393#_M1033_g N_VPWR_c_1775_n 9.39239e-19 $X=6.44 $Y=2.525 $X2=0
+ $Y2=0
cc_757 N_A_1273_393#_M1018_g N_VPWR_c_1775_n 7.97988e-19 $X=9.08 $Y=2.285 $X2=0
+ $Y2=0
cc_758 N_A_1273_393#_c_894_n N_VPWR_c_1775_n 0.0160107f $X=8.22 $Y=2.415 $X2=0
+ $Y2=0
cc_759 N_A_1273_393#_c_878_n N_VPWR_c_1775_n 0.00889837f $X=7.38 $Y=2.415 $X2=0
+ $Y2=0
cc_760 N_A_1273_393#_c_885_n N_VPWR_c_1775_n 0.00671416f $X=8.345 $Y=2.415 $X2=0
+ $Y2=0
cc_761 N_A_1273_393#_c_882_n N_A_636_531#_c_1972_n 3.56662e-19 $X=6.745 $Y=1.95
+ $X2=0 $Y2=0
cc_762 N_A_1273_393#_c_882_n N_A_636_531#_c_1964_n 3.43685e-19 $X=6.745 $Y=1.95
+ $X2=0 $Y2=0
cc_763 N_A_1273_393#_M1001_g N_VGND_c_2173_n 0.0115588f $X=6.88 $Y=0.805 $X2=0
+ $Y2=0
cc_764 N_A_1273_393#_c_871_n N_VGND_c_2173_n 0.0204307f $X=8.34 $Y=0.885 $X2=0
+ $Y2=0
cc_765 N_A_1273_393#_c_868_n N_VGND_c_2174_n 0.0273746f $X=9.05 $Y=1.375 $X2=0
+ $Y2=0
cc_766 N_A_1273_393#_c_870_n N_VGND_c_2174_n 0.0188002f $X=8.9 $Y=1.54 $X2=0
+ $Y2=0
cc_767 N_A_1273_393#_c_871_n N_VGND_c_2174_n 0.0445769f $X=8.34 $Y=0.885 $X2=0
+ $Y2=0
cc_768 N_A_1273_393#_c_873_n N_VGND_c_2174_n 0.00345394f $X=9.05 $Y=1.54 $X2=0
+ $Y2=0
cc_769 N_A_1273_393#_c_871_n N_VGND_c_2186_n 0.0125992f $X=8.34 $Y=0.885 $X2=0
+ $Y2=0
cc_770 N_A_1273_393#_M1001_g N_VGND_c_2190_n 9.39239e-19 $X=6.88 $Y=0.805 $X2=0
+ $Y2=0
cc_771 N_A_1273_393#_c_868_n N_VGND_c_2190_n 9.49986e-19 $X=9.05 $Y=1.375 $X2=0
+ $Y2=0
cc_772 N_A_1273_393#_c_871_n N_VGND_c_2190_n 0.0152817f $X=8.34 $Y=0.885 $X2=0
+ $Y2=0
cc_773 N_A_1139_463#_M1038_g N_ASYNC_M1010_g 0.0323631f $X=7.43 $Y=0.915 $X2=0
+ $Y2=0
cc_774 N_A_1139_463#_M1019_g N_ASYNC_M1034_g 0.0218515f $X=7.43 $Y=2.285 $X2=0
+ $Y2=0
cc_775 N_A_1139_463#_c_1014_n N_ASYNC_c_1101_n 0.0174154f $X=7.34 $Y=1.46 $X2=0
+ $Y2=0
cc_776 N_A_1139_463#_c_1015_n N_ASYNC_c_1101_n 0.00119627f $X=7.34 $Y=1.54 $X2=0
+ $Y2=0
cc_777 N_A_1139_463#_M1019_g N_ASYNC_c_1109_n 0.00638448f $X=7.43 $Y=2.285 $X2=0
+ $Y2=0
cc_778 N_A_1139_463#_c_1014_n N_ASYNC_c_1102_n 0.0012411f $X=7.34 $Y=1.46 $X2=0
+ $Y2=0
cc_779 N_A_1139_463#_c_1015_n N_ASYNC_c_1102_n 0.0323631f $X=7.34 $Y=1.54 $X2=0
+ $Y2=0
cc_780 N_A_1139_463#_c_1017_n N_A_761_357#_c_1246_n 0.0037375f $X=6.22 $Y=2.595
+ $X2=0 $Y2=0
cc_781 N_A_1139_463#_c_1010_n N_A_761_357#_M1032_g 0.00269029f $X=6.305 $Y=0.805
+ $X2=0 $Y2=0
cc_782 N_A_1139_463#_c_1017_n N_A_761_357#_M1017_g 0.0156027f $X=6.22 $Y=2.595
+ $X2=0 $Y2=0
cc_783 N_A_1139_463#_c_1011_n N_A_761_357#_M1017_g 0.00439957f $X=6.305 $Y=2.435
+ $X2=0 $Y2=0
cc_784 N_A_1139_463#_M1038_g N_A_761_357#_c_1237_n 0.0103107f $X=7.43 $Y=0.915
+ $X2=0 $Y2=0
cc_785 N_A_1139_463#_c_1010_n N_A_761_357#_c_1237_n 0.00461852f $X=6.305
+ $Y=0.805 $X2=0 $Y2=0
cc_786 N_A_1139_463#_M1019_g N_A_761_357#_c_1249_n 0.00856127f $X=7.43 $Y=2.285
+ $X2=0 $Y2=0
cc_787 N_A_1139_463#_c_1017_n N_A_761_357#_c_1249_n 0.00310727f $X=6.22 $Y=2.595
+ $X2=0 $Y2=0
cc_788 N_A_1139_463#_M1019_g N_VPWR_c_1779_n 0.00359689f $X=7.43 $Y=2.285 $X2=0
+ $Y2=0
cc_789 N_A_1139_463#_c_1017_n N_VPWR_c_1779_n 0.0137149f $X=6.22 $Y=2.595 $X2=0
+ $Y2=0
cc_790 N_A_1139_463#_c_1011_n N_VPWR_c_1779_n 0.00522766f $X=6.305 $Y=2.435
+ $X2=0 $Y2=0
cc_791 N_A_1139_463#_M1019_g N_VPWR_c_1780_n 0.00359875f $X=7.43 $Y=2.285 $X2=0
+ $Y2=0
cc_792 N_A_1139_463#_c_1017_n N_VPWR_c_1792_n 0.0154231f $X=6.22 $Y=2.595 $X2=0
+ $Y2=0
cc_793 N_A_1139_463#_M1019_g N_VPWR_c_1775_n 9.49986e-19 $X=7.43 $Y=2.285 $X2=0
+ $Y2=0
cc_794 N_A_1139_463#_c_1017_n N_VPWR_c_1775_n 0.019134f $X=6.22 $Y=2.595 $X2=0
+ $Y2=0
cc_795 N_A_1139_463#_c_1017_n N_A_636_531#_c_1971_n 0.013596f $X=6.22 $Y=2.595
+ $X2=0 $Y2=0
cc_796 N_A_1139_463#_c_1017_n N_A_636_531#_c_1972_n 0.0239287f $X=6.22 $Y=2.595
+ $X2=0 $Y2=0
cc_797 N_A_1139_463#_c_1011_n N_A_636_531#_c_1972_n 0.0134653f $X=6.305 $Y=2.435
+ $X2=0 $Y2=0
cc_798 N_A_1139_463#_c_1010_n N_A_636_531#_c_1964_n 0.0252895f $X=6.305 $Y=0.805
+ $X2=0 $Y2=0
cc_799 N_A_1139_463#_c_1011_n N_A_636_531#_c_1964_n 0.0369722f $X=6.305 $Y=2.435
+ $X2=0 $Y2=0
cc_800 N_A_1139_463#_c_1013_n N_A_636_531#_c_1964_n 0.0130993f $X=6.345 $Y=1.46
+ $X2=0 $Y2=0
cc_801 N_A_1139_463#_c_1010_n N_A_636_531#_c_1968_n 3.44058e-19 $X=6.305
+ $Y=0.805 $X2=0 $Y2=0
cc_802 N_A_1139_463#_c_1010_n N_A_636_531#_c_1969_n 0.0184563f $X=6.305 $Y=0.805
+ $X2=0 $Y2=0
cc_803 N_A_1139_463#_c_1017_n A_1225_463# 0.00152387f $X=6.22 $Y=2.595 $X2=-0.19
+ $Y2=-0.245
cc_804 N_A_1139_463#_c_1011_n A_1225_463# 0.00132484f $X=6.305 $Y=2.435
+ $X2=-0.19 $Y2=-0.245
cc_805 N_A_1139_463#_M1038_g N_VGND_c_2173_n 0.0172156f $X=7.43 $Y=0.915 $X2=0
+ $Y2=0
cc_806 N_A_1139_463#_c_1010_n N_VGND_c_2173_n 0.0182894f $X=6.305 $Y=0.805 $X2=0
+ $Y2=0
cc_807 N_A_1139_463#_c_1012_n N_VGND_c_2173_n 0.009263f $X=7.175 $Y=1.46 $X2=0
+ $Y2=0
cc_808 N_A_1139_463#_c_1014_n N_VGND_c_2173_n 0.0128905f $X=7.34 $Y=1.46 $X2=0
+ $Y2=0
cc_809 N_A_1139_463#_c_1015_n N_VGND_c_2173_n 0.00122759f $X=7.34 $Y=1.54 $X2=0
+ $Y2=0
cc_810 N_A_1139_463#_c_1010_n N_VGND_c_2180_n 0.00565285f $X=6.305 $Y=0.805
+ $X2=0 $Y2=0
cc_811 N_A_1139_463#_M1038_g N_VGND_c_2190_n 7.88961e-19 $X=7.43 $Y=0.915 $X2=0
+ $Y2=0
cc_812 N_A_1139_463#_c_1010_n N_VGND_c_2190_n 0.00685297f $X=6.305 $Y=0.805
+ $X2=0 $Y2=0
cc_813 N_ASYNC_M1010_g N_A_761_357#_c_1237_n 0.0102957f $X=7.82 $Y=0.915 $X2=0
+ $Y2=0
cc_814 N_ASYNC_M1034_g N_A_761_357#_c_1249_n 0.00861299f $X=8.09 $Y=2.285 $X2=0
+ $Y2=0
cc_815 N_ASYNC_c_1108_n N_A_761_357#_M1042_g 0.00809106f $X=11.135 $Y=2.035
+ $X2=0 $Y2=0
cc_816 N_ASYNC_c_1108_n N_A_2083_65#_M1008_g 0.00543237f $X=11.135 $Y=2.035
+ $X2=0 $Y2=0
cc_817 N_ASYNC_M1035_g N_A_2083_65#_M1023_g 0.0172056f $X=11.58 $Y=2.675 $X2=0
+ $Y2=0
cc_818 N_ASYNC_c_1106_n N_A_2083_65#_M1023_g 0.00163399f $X=11.67 $Y=1.93 $X2=0
+ $Y2=0
cc_819 N_ASYNC_c_1107_n N_A_2083_65#_M1023_g 0.017824f $X=11.67 $Y=1.93 $X2=0
+ $Y2=0
cc_820 N_ASYNC_c_1100_n N_A_2083_65#_M1026_g 0.00560936f $X=11.58 $Y=1.06 $X2=0
+ $Y2=0
cc_821 N_ASYNC_c_1108_n N_A_2083_65#_c_1434_n 0.00691819f $X=11.135 $Y=2.035
+ $X2=0 $Y2=0
cc_822 ASYNC N_A_2083_65#_c_1434_n 9.82613e-19 $X=11.195 $Y=1.95 $X2=0 $Y2=0
cc_823 N_ASYNC_c_1100_n N_A_2083_65#_c_1422_n 0.00440649f $X=11.58 $Y=1.06 $X2=0
+ $Y2=0
cc_824 N_ASYNC_c_1108_n N_A_2083_65#_c_1422_n 0.0143321f $X=11.135 $Y=2.035
+ $X2=0 $Y2=0
cc_825 ASYNC N_A_2083_65#_c_1422_n 0.00249744f $X=11.195 $Y=1.95 $X2=0 $Y2=0
cc_826 N_ASYNC_c_1113_n N_A_2083_65#_c_1422_n 0.0193697f $X=11.395 $Y=1.977
+ $X2=0 $Y2=0
cc_827 N_ASYNC_c_1108_n N_A_2083_65#_c_1458_n 0.0160689f $X=11.135 $Y=2.035
+ $X2=0 $Y2=0
cc_828 ASYNC N_A_2083_65#_c_1458_n 0.00199287f $X=11.195 $Y=1.95 $X2=0 $Y2=0
cc_829 N_ASYNC_c_1113_n N_A_2083_65#_c_1458_n 0.00194862f $X=11.395 $Y=1.977
+ $X2=0 $Y2=0
cc_830 N_ASYNC_c_1099_n N_A_2083_65#_c_1424_n 0.0185806f $X=11.395 $Y=0.985
+ $X2=0 $Y2=0
cc_831 N_ASYNC_c_1100_n N_A_2083_65#_c_1424_n 0.0125016f $X=11.58 $Y=1.06 $X2=0
+ $Y2=0
cc_832 N_ASYNC_c_1103_n N_A_2083_65#_c_1424_n 0.0106767f $X=11.697 $Y=1.765
+ $X2=0 $Y2=0
cc_833 N_ASYNC_c_1106_n N_A_2083_65#_c_1425_n 0.00424076f $X=11.67 $Y=1.93 $X2=0
+ $Y2=0
cc_834 N_ASYNC_c_1107_n N_A_2083_65#_c_1425_n 0.00295162f $X=11.67 $Y=1.93 $X2=0
+ $Y2=0
cc_835 N_ASYNC_c_1108_n N_A_2083_65#_c_1435_n 0.0271963f $X=11.135 $Y=2.035
+ $X2=0 $Y2=0
cc_836 ASYNC N_A_2083_65#_c_1435_n 9.55543e-19 $X=11.195 $Y=1.95 $X2=0 $Y2=0
cc_837 N_ASYNC_c_1113_n N_A_2083_65#_c_1435_n 0.0094469f $X=11.395 $Y=1.977
+ $X2=0 $Y2=0
cc_838 N_ASYNC_c_1108_n N_A_2083_65#_c_1436_n 0.00180829f $X=11.135 $Y=2.035
+ $X2=0 $Y2=0
cc_839 ASYNC N_A_2083_65#_c_1436_n 2.41601e-19 $X=11.195 $Y=1.95 $X2=0 $Y2=0
cc_840 N_ASYNC_c_1113_n N_A_2083_65#_c_1436_n 0.00103358f $X=11.395 $Y=1.977
+ $X2=0 $Y2=0
cc_841 N_ASYNC_M1035_g N_A_2083_65#_c_1472_n 0.00861087f $X=11.58 $Y=2.675 $X2=0
+ $Y2=0
cc_842 N_ASYNC_c_1106_n N_A_2083_65#_c_1472_n 0.00642584f $X=11.67 $Y=1.93 $X2=0
+ $Y2=0
cc_843 ASYNC N_A_2083_65#_c_1472_n 0.00628386f $X=11.195 $Y=1.95 $X2=0 $Y2=0
cc_844 N_ASYNC_c_1113_n N_A_2083_65#_c_1472_n 0.0112416f $X=11.395 $Y=1.977
+ $X2=0 $Y2=0
cc_845 N_ASYNC_c_1106_n N_A_2083_65#_c_1427_n 0.0259869f $X=11.67 $Y=1.93 $X2=0
+ $Y2=0
cc_846 N_ASYNC_c_1107_n N_A_2083_65#_c_1427_n 0.00291956f $X=11.67 $Y=1.93 $X2=0
+ $Y2=0
cc_847 N_ASYNC_c_1103_n N_A_2083_65#_c_1427_n 0.00937882f $X=11.697 $Y=1.765
+ $X2=0 $Y2=0
cc_848 N_ASYNC_c_1103_n N_A_2083_65#_c_1428_n 8.86512e-19 $X=11.697 $Y=1.765
+ $X2=0 $Y2=0
cc_849 N_ASYNC_c_1107_n N_A_2083_65#_c_1430_n 0.00137668f $X=11.67 $Y=1.93 $X2=0
+ $Y2=0
cc_850 N_ASYNC_c_1103_n N_A_2083_65#_c_1430_n 0.00819877f $X=11.697 $Y=1.765
+ $X2=0 $Y2=0
cc_851 N_ASYNC_c_1107_n N_A_1903_125#_M1015_g 0.025269f $X=11.67 $Y=1.93 $X2=0
+ $Y2=0
cc_852 N_ASYNC_c_1108_n N_A_1903_125#_M1015_g 0.00222784f $X=11.135 $Y=2.035
+ $X2=0 $Y2=0
cc_853 ASYNC N_A_1903_125#_M1015_g 0.002102f $X=11.195 $Y=1.95 $X2=0 $Y2=0
cc_854 N_ASYNC_c_1113_n N_A_1903_125#_M1015_g 0.010307f $X=11.395 $Y=1.977 $X2=0
+ $Y2=0
cc_855 N_ASYNC_c_1099_n N_A_1903_125#_c_1585_n 0.0309549f $X=11.395 $Y=0.985
+ $X2=0 $Y2=0
cc_856 N_ASYNC_c_1103_n N_A_1903_125#_c_1587_n 0.025269f $X=11.697 $Y=1.765
+ $X2=0 $Y2=0
cc_857 N_ASYNC_c_1108_n N_A_1903_125#_c_1594_n 0.0319254f $X=11.135 $Y=2.035
+ $X2=0 $Y2=0
cc_858 N_ASYNC_c_1108_n N_A_1903_125#_c_1589_n 0.00702355f $X=11.135 $Y=2.035
+ $X2=0 $Y2=0
cc_859 N_ASYNC_c_1100_n N_A_1903_125#_c_1590_n 5.67729e-19 $X=11.58 $Y=1.06
+ $X2=0 $Y2=0
cc_860 N_ASYNC_c_1100_n N_A_1903_125#_c_1591_n 0.0309549f $X=11.58 $Y=1.06 $X2=0
+ $Y2=0
cc_861 N_ASYNC_c_1103_n N_A_1903_125#_c_1591_n 0.00668295f $X=11.697 $Y=1.765
+ $X2=0 $Y2=0
cc_862 N_ASYNC_M1035_g N_A_2456_451#_c_1687_n 2.19003e-19 $X=11.58 $Y=2.675
+ $X2=0 $Y2=0
cc_863 N_ASYNC_c_1121_n N_VPWR_M1019_d 0.00153076f $X=8.065 $Y=2.035 $X2=0 $Y2=0
cc_864 N_ASYNC_c_1109_n N_VPWR_M1019_d 0.00599344f $X=7.92 $Y=2.035 $X2=0 $Y2=0
cc_865 N_ASYNC_M1034_g N_VPWR_c_1780_n 0.00365382f $X=8.09 $Y=2.285 $X2=0 $Y2=0
cc_866 N_ASYNC_M1034_g N_VPWR_c_1781_n 0.00317893f $X=8.09 $Y=2.285 $X2=0 $Y2=0
cc_867 N_ASYNC_c_1108_n N_VPWR_c_1781_n 0.0308426f $X=11.135 $Y=2.035 $X2=0
+ $Y2=0
cc_868 N_ASYNC_c_1108_n N_VPWR_c_1782_n 7.89152e-19 $X=11.135 $Y=2.035 $X2=0
+ $Y2=0
cc_869 N_ASYNC_M1035_g N_VPWR_c_1783_n 0.00549284f $X=11.58 $Y=2.675 $X2=0 $Y2=0
cc_870 N_ASYNC_M1035_g N_VPWR_c_1784_n 0.0108315f $X=11.58 $Y=2.675 $X2=0 $Y2=0
cc_871 N_ASYNC_c_1106_n N_VPWR_c_1784_n 0.0096659f $X=11.67 $Y=1.93 $X2=0 $Y2=0
cc_872 N_ASYNC_c_1107_n N_VPWR_c_1784_n 0.0044969f $X=11.67 $Y=1.93 $X2=0 $Y2=0
cc_873 N_ASYNC_M1034_g N_VPWR_c_1775_n 9.49986e-19 $X=8.09 $Y=2.285 $X2=0 $Y2=0
cc_874 N_ASYNC_M1035_g N_VPWR_c_1775_n 0.0113256f $X=11.58 $Y=2.675 $X2=0 $Y2=0
cc_875 N_ASYNC_c_1108_n A_1831_373# 0.015295f $X=11.135 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_876 N_ASYNC_M1010_g N_VGND_c_2173_n 0.00230357f $X=7.82 $Y=0.915 $X2=0 $Y2=0
cc_877 N_ASYNC_c_1099_n N_VGND_c_2175_n 0.00275178f $X=11.395 $Y=0.985 $X2=0
+ $Y2=0
cc_878 N_ASYNC_c_1099_n N_VGND_c_2176_n 0.00354497f $X=11.395 $Y=0.985 $X2=0
+ $Y2=0
cc_879 N_ASYNC_c_1099_n N_VGND_c_2188_n 0.00549284f $X=11.395 $Y=0.985 $X2=0
+ $Y2=0
cc_880 N_ASYNC_M1010_g N_VGND_c_2190_n 9.39239e-19 $X=7.82 $Y=0.915 $X2=0 $Y2=0
cc_881 N_ASYNC_c_1099_n N_VGND_c_2190_n 0.0113234f $X=11.395 $Y=0.985 $X2=0
+ $Y2=0
cc_882 N_A_761_357#_M1021_g N_A_2083_65#_c_1419_n 0.0350573f $X=10.1 $Y=0.665
+ $X2=0 $Y2=0
cc_883 N_A_761_357#_c_1237_n N_A_1903_125#_c_1588_n 0.00739039f $X=10.025
+ $Y=0.18 $X2=0 $Y2=0
cc_884 N_A_761_357#_M1021_g N_A_1903_125#_c_1588_n 0.0195267f $X=10.1 $Y=0.665
+ $X2=0 $Y2=0
cc_885 N_A_761_357#_M1021_g N_A_1903_125#_c_1597_n 7.43301e-19 $X=10.1 $Y=0.665
+ $X2=0 $Y2=0
cc_886 N_A_761_357#_M1042_g N_A_1903_125#_c_1594_n 0.0198042f $X=9.59 $Y=2.465
+ $X2=0 $Y2=0
cc_887 N_A_761_357#_M1042_g N_A_1903_125#_c_1589_n 0.00119912f $X=9.59 $Y=2.465
+ $X2=0 $Y2=0
cc_888 N_A_761_357#_M1021_g N_A_1903_125#_c_1592_n 0.00796874f $X=10.1 $Y=0.665
+ $X2=0 $Y2=0
cc_889 N_A_761_357#_c_1253_n N_VPWR_M1005_d 0.00180133f $X=4.375 $Y=1.78 $X2=0
+ $Y2=0
cc_890 N_A_761_357#_M1029_g N_VPWR_c_1778_n 0.0153164f $X=4.595 $Y=2.415 $X2=0
+ $Y2=0
cc_891 N_A_761_357#_c_1234_n N_VPWR_c_1778_n 0.0010106f $X=5.105 $Y=3.075 $X2=0
+ $Y2=0
cc_892 N_A_761_357#_c_1247_n N_VPWR_c_1778_n 8.93566e-19 $X=5.18 $Y=3.15 $X2=0
+ $Y2=0
cc_893 N_A_761_357#_c_1252_n N_VPWR_c_1778_n 0.0372447f $X=3.95 $Y=1.93 $X2=0
+ $Y2=0
cc_894 N_A_761_357#_c_1253_n N_VPWR_c_1778_n 0.0167279f $X=4.375 $Y=1.78 $X2=0
+ $Y2=0
cc_895 N_A_761_357#_M1017_g N_VPWR_c_1779_n 0.00581491f $X=6.05 $Y=2.525 $X2=0
+ $Y2=0
cc_896 N_A_761_357#_c_1249_n N_VPWR_c_1779_n 0.0216291f $X=9.515 $Y=3.15 $X2=0
+ $Y2=0
cc_897 N_A_761_357#_c_1249_n N_VPWR_c_1780_n 0.0252872f $X=9.515 $Y=3.15 $X2=0
+ $Y2=0
cc_898 N_A_761_357#_c_1249_n N_VPWR_c_1781_n 0.0257368f $X=9.515 $Y=3.15 $X2=0
+ $Y2=0
cc_899 N_A_761_357#_M1042_g N_VPWR_c_1781_n 0.00883595f $X=9.59 $Y=2.465 $X2=0
+ $Y2=0
cc_900 N_A_761_357#_c_1252_n N_VPWR_c_1790_n 0.0113273f $X=3.95 $Y=1.93 $X2=0
+ $Y2=0
cc_901 N_A_761_357#_M1029_g N_VPWR_c_1792_n 0.00445056f $X=4.595 $Y=2.415 $X2=0
+ $Y2=0
cc_902 N_A_761_357#_c_1247_n N_VPWR_c_1792_n 0.0454664f $X=5.18 $Y=3.15 $X2=0
+ $Y2=0
cc_903 N_A_761_357#_c_1249_n N_VPWR_c_1794_n 0.0236924f $X=9.515 $Y=3.15 $X2=0
+ $Y2=0
cc_904 N_A_761_357#_c_1249_n N_VPWR_c_1798_n 0.024594f $X=9.515 $Y=3.15 $X2=0
+ $Y2=0
cc_905 N_A_761_357#_c_1249_n N_VPWR_c_1799_n 0.0229586f $X=9.515 $Y=3.15 $X2=0
+ $Y2=0
cc_906 N_A_761_357#_M1029_g N_VPWR_c_1775_n 0.0082324f $X=4.595 $Y=2.415 $X2=0
+ $Y2=0
cc_907 N_A_761_357#_c_1246_n N_VPWR_c_1775_n 0.0253712f $X=5.975 $Y=3.15 $X2=0
+ $Y2=0
cc_908 N_A_761_357#_c_1247_n N_VPWR_c_1775_n 0.0107868f $X=5.18 $Y=3.15 $X2=0
+ $Y2=0
cc_909 N_A_761_357#_c_1249_n N_VPWR_c_1775_n 0.103074f $X=9.515 $Y=3.15 $X2=0
+ $Y2=0
cc_910 N_A_761_357#_c_1251_n N_VPWR_c_1775_n 0.00416972f $X=6.05 $Y=3.15 $X2=0
+ $Y2=0
cc_911 N_A_761_357#_c_1252_n N_VPWR_c_1775_n 0.00650045f $X=3.95 $Y=1.93 $X2=0
+ $Y2=0
cc_912 N_A_761_357#_c_1252_n N_A_636_531#_c_1963_n 0.0574121f $X=3.95 $Y=1.93
+ $X2=0 $Y2=0
cc_913 N_A_761_357#_c_1257_n N_A_636_531#_c_1963_n 0.00976949f $X=3.99 $Y=0.43
+ $X2=0 $Y2=0
cc_914 N_A_761_357#_c_1254_n N_A_636_531#_c_1963_n 0.0136422f $X=4.035 $Y=1.78
+ $X2=0 $Y2=0
cc_915 N_A_761_357#_c_1260_n N_A_636_531#_c_1963_n 0.0116035f $X=4.155 $Y=0.915
+ $X2=0 $Y2=0
cc_916 N_A_761_357#_c_1234_n N_A_636_531#_c_1971_n 0.00443646f $X=5.105 $Y=3.075
+ $X2=0 $Y2=0
cc_917 N_A_761_357#_c_1246_n N_A_636_531#_c_1971_n 0.00442759f $X=5.975 $Y=3.15
+ $X2=0 $Y2=0
cc_918 N_A_761_357#_M1017_g N_A_636_531#_c_1972_n 0.00381988f $X=6.05 $Y=2.525
+ $X2=0 $Y2=0
cc_919 N_A_761_357#_c_1234_n N_A_636_531#_c_1973_n 0.00168005f $X=5.105 $Y=3.075
+ $X2=0 $Y2=0
cc_920 N_A_761_357#_c_1235_n N_A_636_531#_c_1964_n 0.00879203f $X=5.86 $Y=1.26
+ $X2=0 $Y2=0
cc_921 N_A_761_357#_M1032_g N_A_636_531#_c_1964_n 0.00597368f $X=5.935 $Y=0.805
+ $X2=0 $Y2=0
cc_922 N_A_761_357#_c_1243_n N_A_636_531#_c_1964_n 6.66351e-19 $X=5.18 $Y=1.37
+ $X2=0 $Y2=0
cc_923 N_A_761_357#_c_1252_n N_A_636_531#_c_1975_n 0.0230052f $X=3.95 $Y=1.93
+ $X2=0 $Y2=0
cc_924 N_A_761_357#_M1039_s N_A_636_531#_c_1965_n 0.00177172f $X=3.845 $Y=0.235
+ $X2=0 $Y2=0
cc_925 N_A_761_357#_c_1233_n N_A_636_531#_c_1965_n 0.00408701f $X=4.795 $Y=1.185
+ $X2=0 $Y2=0
cc_926 N_A_761_357#_c_1257_n N_A_636_531#_c_1965_n 0.0147405f $X=3.99 $Y=0.43
+ $X2=0 $Y2=0
cc_927 N_A_761_357#_c_1270_n N_A_636_531#_c_1965_n 0.00854757f $X=4.375 $Y=0.915
+ $X2=0 $Y2=0
cc_928 N_A_761_357#_c_1242_n N_A_636_531#_c_1965_n 0.00549366f $X=4.685 $Y=1.39
+ $X2=0 $Y2=0
cc_929 N_A_761_357#_c_1243_n N_A_636_531#_c_1965_n 0.00419774f $X=5.18 $Y=1.37
+ $X2=0 $Y2=0
cc_930 N_A_761_357#_c_1257_n N_A_636_531#_c_1966_n 0.00265521f $X=3.99 $Y=0.43
+ $X2=0 $Y2=0
cc_931 N_A_761_357#_c_1257_n N_A_636_531#_c_1967_n 0.0280113f $X=3.99 $Y=0.43
+ $X2=0 $Y2=0
cc_932 N_A_761_357#_c_1235_n N_A_636_531#_c_1968_n 5.61748e-19 $X=5.86 $Y=1.26
+ $X2=0 $Y2=0
cc_933 N_A_761_357#_c_1233_n N_A_636_531#_c_1969_n 0.00100798f $X=4.795 $Y=1.185
+ $X2=0 $Y2=0
cc_934 N_A_761_357#_c_1235_n N_A_636_531#_c_1969_n 0.0104783f $X=5.86 $Y=1.26
+ $X2=0 $Y2=0
cc_935 N_A_761_357#_M1032_g N_A_636_531#_c_1969_n 0.0201556f $X=5.935 $Y=0.805
+ $X2=0 $Y2=0
cc_936 N_A_761_357#_c_1270_n N_VGND_M1039_d 0.00616544f $X=4.375 $Y=0.915 $X2=0
+ $Y2=0
cc_937 N_A_761_357#_c_1240_n N_VGND_M1039_d 0.00169703f $X=4.46 $Y=1.225 $X2=0
+ $Y2=0
cc_938 N_A_761_357#_c_1233_n N_VGND_c_2172_n 0.0057576f $X=4.795 $Y=1.185 $X2=0
+ $Y2=0
cc_939 N_A_761_357#_c_1257_n N_VGND_c_2172_n 0.0150732f $X=3.99 $Y=0.43 $X2=0
+ $Y2=0
cc_940 N_A_761_357#_c_1270_n N_VGND_c_2172_n 0.0155101f $X=4.375 $Y=0.915 $X2=0
+ $Y2=0
cc_941 N_A_761_357#_c_1242_n N_VGND_c_2172_n 0.00311983f $X=4.685 $Y=1.39 $X2=0
+ $Y2=0
cc_942 N_A_761_357#_c_1243_n N_VGND_c_2172_n 0.0026277f $X=5.18 $Y=1.37 $X2=0
+ $Y2=0
cc_943 N_A_761_357#_c_1237_n N_VGND_c_2173_n 0.025796f $X=10.025 $Y=0.18 $X2=0
+ $Y2=0
cc_944 N_A_761_357#_c_1237_n N_VGND_c_2174_n 0.0216291f $X=10.025 $Y=0.18 $X2=0
+ $Y2=0
cc_945 N_A_761_357#_c_1237_n N_VGND_c_2175_n 0.00549693f $X=10.025 $Y=0.18 $X2=0
+ $Y2=0
cc_946 N_A_761_357#_c_1233_n N_VGND_c_2180_n 0.00549284f $X=4.795 $Y=1.185 $X2=0
+ $Y2=0
cc_947 N_A_761_357#_c_1238_n N_VGND_c_2180_n 0.0377554f $X=6.01 $Y=0.18 $X2=0
+ $Y2=0
cc_948 N_A_761_357#_c_1257_n N_VGND_c_2185_n 0.014447f $X=3.99 $Y=0.43 $X2=0
+ $Y2=0
cc_949 N_A_761_357#_c_1237_n N_VGND_c_2186_n 0.0379965f $X=10.025 $Y=0.18 $X2=0
+ $Y2=0
cc_950 N_A_761_357#_c_1237_n N_VGND_c_2187_n 0.0407578f $X=10.025 $Y=0.18 $X2=0
+ $Y2=0
cc_951 N_A_761_357#_M1039_s N_VGND_c_2190_n 0.00170858f $X=3.845 $Y=0.235 $X2=0
+ $Y2=0
cc_952 N_A_761_357#_c_1233_n N_VGND_c_2190_n 0.00710682f $X=4.795 $Y=1.185 $X2=0
+ $Y2=0
cc_953 N_A_761_357#_c_1237_n N_VGND_c_2190_n 0.143367f $X=10.025 $Y=0.18 $X2=0
+ $Y2=0
cc_954 N_A_761_357#_c_1238_n N_VGND_c_2190_n 0.00622941f $X=6.01 $Y=0.18 $X2=0
+ $Y2=0
cc_955 N_A_761_357#_c_1257_n N_VGND_c_2190_n 0.00293246f $X=3.99 $Y=0.43 $X2=0
+ $Y2=0
cc_956 N_A_2083_65#_M1008_g N_A_1903_125#_M1015_g 0.014947f $X=10.525 $Y=2.465
+ $X2=0 $Y2=0
cc_957 N_A_2083_65#_c_1434_n N_A_1903_125#_M1015_g 0.00375014f $X=10.665 $Y=2.33
+ $X2=0 $Y2=0
cc_958 N_A_2083_65#_c_1422_n N_A_1903_125#_M1015_g 0.0066805f $X=11.445 $Y=1.54
+ $X2=0 $Y2=0
cc_959 N_A_2083_65#_c_1458_n N_A_1903_125#_M1015_g 0.00971003f $X=11.2 $Y=2.415
+ $X2=0 $Y2=0
cc_960 N_A_2083_65#_c_1435_n N_A_1903_125#_M1015_g 0.00132561f $X=10.585 $Y=1.93
+ $X2=0 $Y2=0
cc_961 N_A_2083_65#_c_1436_n N_A_1903_125#_M1015_g 0.0127829f $X=10.585 $Y=1.93
+ $X2=0 $Y2=0
cc_962 N_A_2083_65#_c_1426_n N_A_1903_125#_M1015_g 0.00261342f $X=10.585
+ $Y=1.765 $X2=0 $Y2=0
cc_963 N_A_2083_65#_c_1472_n N_A_1903_125#_M1015_g 0.0090699f $X=11.365 $Y=2.495
+ $X2=0 $Y2=0
cc_964 N_A_2083_65#_c_1429_n N_A_1903_125#_M1015_g 0.00376465f $X=10.585
+ $Y=1.765 $X2=0 $Y2=0
cc_965 N_A_2083_65#_c_1419_n N_A_1903_125#_c_1585_n 0.0131311f $X=10.492
+ $Y=0.985 $X2=0 $Y2=0
cc_966 N_A_2083_65#_c_1424_n N_A_1903_125#_c_1585_n 0.00237297f $X=11.61 $Y=0.58
+ $X2=0 $Y2=0
cc_967 N_A_2083_65#_c_1424_n N_A_1903_125#_c_1586_n 0.00210955f $X=11.61 $Y=0.58
+ $X2=0 $Y2=0
cc_968 N_A_2083_65#_c_1429_n N_A_1903_125#_c_1586_n 0.0175527f $X=10.585
+ $Y=1.765 $X2=0 $Y2=0
cc_969 N_A_2083_65#_c_1422_n N_A_1903_125#_c_1587_n 0.0179312f $X=11.445 $Y=1.54
+ $X2=0 $Y2=0
cc_970 N_A_2083_65#_c_1424_n N_A_1903_125#_c_1587_n 0.00182301f $X=11.61 $Y=0.58
+ $X2=0 $Y2=0
cc_971 N_A_2083_65#_c_1419_n N_A_1903_125#_c_1588_n 0.001968f $X=10.492 $Y=0.985
+ $X2=0 $Y2=0
cc_972 N_A_2083_65#_c_1434_n N_A_1903_125#_c_1594_n 0.00679569f $X=10.665
+ $Y=2.33 $X2=0 $Y2=0
cc_973 N_A_2083_65#_c_1443_n N_A_1903_125#_c_1594_n 0.00507581f $X=10.75
+ $Y=2.415 $X2=0 $Y2=0
cc_974 N_A_2083_65#_c_1423_n N_A_1903_125#_c_1589_n 0.0061555f $X=10.75 $Y=1.54
+ $X2=0 $Y2=0
cc_975 N_A_2083_65#_c_1435_n N_A_1903_125#_c_1589_n 0.012051f $X=10.585 $Y=1.93
+ $X2=0 $Y2=0
cc_976 N_A_2083_65#_c_1426_n N_A_1903_125#_c_1589_n 0.00438521f $X=10.585
+ $Y=1.765 $X2=0 $Y2=0
cc_977 N_A_2083_65#_c_1429_n N_A_1903_125#_c_1589_n 0.00958141f $X=10.585
+ $Y=1.765 $X2=0 $Y2=0
cc_978 N_A_2083_65#_c_1422_n N_A_1903_125#_c_1590_n 0.0222786f $X=11.445 $Y=1.54
+ $X2=0 $Y2=0
cc_979 N_A_2083_65#_c_1424_n N_A_1903_125#_c_1590_n 0.0136811f $X=11.61 $Y=0.58
+ $X2=0 $Y2=0
cc_980 N_A_2083_65#_c_1429_n N_A_1903_125#_c_1590_n 5.27994e-19 $X=10.585
+ $Y=1.765 $X2=0 $Y2=0
cc_981 N_A_2083_65#_c_1420_n N_A_1903_125#_c_1591_n 0.0175527f $X=10.492
+ $Y=1.135 $X2=0 $Y2=0
cc_982 N_A_2083_65#_c_1424_n N_A_1903_125#_c_1591_n 7.37985e-19 $X=11.61 $Y=0.58
+ $X2=0 $Y2=0
cc_983 N_A_2083_65#_c_1420_n N_A_1903_125#_c_1592_n 0.0136762f $X=10.492
+ $Y=1.135 $X2=0 $Y2=0
cc_984 N_A_2083_65#_c_1422_n N_A_1903_125#_c_1592_n 0.00165131f $X=11.445
+ $Y=1.54 $X2=0 $Y2=0
cc_985 N_A_2083_65#_c_1423_n N_A_1903_125#_c_1592_n 0.0108227f $X=10.75 $Y=1.54
+ $X2=0 $Y2=0
cc_986 N_A_2083_65#_c_1435_n N_A_1903_125#_c_1592_n 0.00430615f $X=10.585
+ $Y=1.93 $X2=0 $Y2=0
cc_987 N_A_2083_65#_c_1436_n N_A_1903_125#_c_1592_n 6.72609e-19 $X=10.585
+ $Y=1.93 $X2=0 $Y2=0
cc_988 N_A_2083_65#_c_1429_n N_A_1903_125#_c_1592_n 0.00672982f $X=10.585
+ $Y=1.765 $X2=0 $Y2=0
cc_989 N_A_2083_65#_M1011_g N_A_2456_451#_M1014_g 0.0385825f $X=13.345 $Y=2.465
+ $X2=0 $Y2=0
cc_990 N_A_2083_65#_M1004_g N_A_2456_451#_M1016_g 0.0231625f $X=13.375 $Y=0.705
+ $X2=0 $Y2=0
cc_991 N_A_2083_65#_M1023_g N_A_2456_451#_c_1677_n 0.0129774f $X=12.205 $Y=2.575
+ $X2=0 $Y2=0
cc_992 N_A_2083_65#_M1026_g N_A_2456_451#_c_1677_n 0.0255047f $X=12.385 $Y=0.495
+ $X2=0 $Y2=0
cc_993 N_A_2083_65#_c_1416_n N_A_2456_451#_c_1677_n 0.0145698f $X=13.27 $Y=1.53
+ $X2=0 $Y2=0
cc_994 N_A_2083_65#_M1011_g N_A_2456_451#_c_1677_n 0.00309097f $X=13.345
+ $Y=2.465 $X2=0 $Y2=0
cc_995 N_A_2083_65#_c_1428_n N_A_2456_451#_c_1677_n 0.0231893f $X=12.265 $Y=1.54
+ $X2=0 $Y2=0
cc_996 N_A_2083_65#_c_1430_n N_A_2456_451#_c_1677_n 0.00422829f $X=12.28 $Y=1.53
+ $X2=0 $Y2=0
cc_997 N_A_2083_65#_M1011_g N_A_2456_451#_c_1684_n 0.0141394f $X=13.345 $Y=2.465
+ $X2=0 $Y2=0
cc_998 N_A_2083_65#_M1011_g N_A_2456_451#_c_1678_n 0.00753132f $X=13.345
+ $Y=2.465 $X2=0 $Y2=0
cc_999 N_A_2083_65#_M1023_g N_A_2456_451#_c_1686_n 0.00554972f $X=12.205
+ $Y=2.575 $X2=0 $Y2=0
cc_1000 N_A_2083_65#_M1011_g N_A_2456_451#_c_1686_n 0.00917211f $X=13.345
+ $Y=2.465 $X2=0 $Y2=0
cc_1001 N_A_2083_65#_M1023_g N_A_2456_451#_c_1687_n 0.00453109f $X=12.205
+ $Y=2.575 $X2=0 $Y2=0
cc_1002 N_A_2083_65#_c_1416_n N_A_2456_451#_c_1687_n 0.00408648f $X=13.27
+ $Y=1.53 $X2=0 $Y2=0
cc_1003 N_A_2083_65#_M1011_g N_A_2456_451#_c_1687_n 0.00250775f $X=13.345
+ $Y=2.465 $X2=0 $Y2=0
cc_1004 N_A_2083_65#_c_1428_n N_A_2456_451#_c_1687_n 0.00644293f $X=12.265
+ $Y=1.54 $X2=0 $Y2=0
cc_1005 N_A_2083_65#_c_1430_n N_A_2456_451#_c_1687_n 0.00188047f $X=12.28
+ $Y=1.53 $X2=0 $Y2=0
cc_1006 N_A_2083_65#_M1026_g N_A_2456_451#_c_1679_n 0.00783423f $X=12.385
+ $Y=0.495 $X2=0 $Y2=0
cc_1007 N_A_2083_65#_M1004_g N_A_2456_451#_c_1679_n 0.00272797f $X=13.375
+ $Y=0.705 $X2=0 $Y2=0
cc_1008 N_A_2083_65#_M1011_g N_A_2456_451#_c_1680_n 3.35186e-19 $X=13.345
+ $Y=2.465 $X2=0 $Y2=0
cc_1009 N_A_2083_65#_M1004_g N_A_2456_451#_c_1680_n 0.00212764f $X=13.375
+ $Y=0.705 $X2=0 $Y2=0
cc_1010 N_A_2083_65#_M1011_g N_A_2456_451#_c_1681_n 0.00246846f $X=13.345
+ $Y=2.465 $X2=0 $Y2=0
cc_1011 N_A_2083_65#_M1004_g N_A_2456_451#_c_1681_n 0.0174608f $X=13.375
+ $Y=0.705 $X2=0 $Y2=0
cc_1012 N_A_2083_65#_c_1434_n N_VPWR_M1008_d 9.73102e-19 $X=10.665 $Y=2.33 $X2=0
+ $Y2=0
cc_1013 N_A_2083_65#_c_1458_n N_VPWR_M1008_d 0.00759485f $X=11.2 $Y=2.415 $X2=0
+ $Y2=0
cc_1014 N_A_2083_65#_c_1443_n N_VPWR_M1008_d 0.0014484f $X=10.75 $Y=2.415 $X2=0
+ $Y2=0
cc_1015 N_A_2083_65#_M1008_g N_VPWR_c_1782_n 0.00352209f $X=10.525 $Y=2.465
+ $X2=0 $Y2=0
cc_1016 N_A_2083_65#_c_1458_n N_VPWR_c_1782_n 0.0195804f $X=11.2 $Y=2.415 $X2=0
+ $Y2=0
cc_1017 N_A_2083_65#_c_1443_n N_VPWR_c_1782_n 0.00478003f $X=10.75 $Y=2.415
+ $X2=0 $Y2=0
cc_1018 N_A_2083_65#_c_1436_n N_VPWR_c_1782_n 2.02124e-19 $X=10.585 $Y=1.93
+ $X2=0 $Y2=0
cc_1019 N_A_2083_65#_c_1472_n N_VPWR_c_1783_n 0.0177952f $X=11.365 $Y=2.495
+ $X2=0 $Y2=0
cc_1020 N_A_2083_65#_M1023_g N_VPWR_c_1784_n 0.00942857f $X=12.205 $Y=2.575
+ $X2=0 $Y2=0
cc_1021 N_A_2083_65#_c_1425_n N_VPWR_c_1784_n 0.00632748f $X=12.1 $Y=1.54 $X2=0
+ $Y2=0
cc_1022 N_A_2083_65#_M1011_g N_VPWR_c_1785_n 0.0235342f $X=13.345 $Y=2.465 $X2=0
+ $Y2=0
cc_1023 N_A_2083_65#_M1023_g N_VPWR_c_1796_n 0.00507528f $X=12.205 $Y=2.575
+ $X2=0 $Y2=0
cc_1024 N_A_2083_65#_M1011_g N_VPWR_c_1796_n 0.00486043f $X=13.345 $Y=2.465
+ $X2=0 $Y2=0
cc_1025 N_A_2083_65#_M1008_g N_VPWR_c_1799_n 0.00399858f $X=10.525 $Y=2.465
+ $X2=0 $Y2=0
cc_1026 N_A_2083_65#_M1015_d N_VPWR_c_1775_n 0.00223819f $X=11.225 $Y=2.255
+ $X2=0 $Y2=0
cc_1027 N_A_2083_65#_M1008_g N_VPWR_c_1775_n 0.0046122f $X=10.525 $Y=2.465 $X2=0
+ $Y2=0
cc_1028 N_A_2083_65#_M1023_g N_VPWR_c_1775_n 0.00525227f $X=12.205 $Y=2.575
+ $X2=0 $Y2=0
cc_1029 N_A_2083_65#_M1011_g N_VPWR_c_1775_n 0.00600853f $X=13.345 $Y=2.465
+ $X2=0 $Y2=0
cc_1030 N_A_2083_65#_c_1458_n N_VPWR_c_1775_n 0.00625607f $X=11.2 $Y=2.415 $X2=0
+ $Y2=0
cc_1031 N_A_2083_65#_c_1443_n N_VPWR_c_1775_n 0.00455894f $X=10.75 $Y=2.415
+ $X2=0 $Y2=0
cc_1032 N_A_2083_65#_c_1472_n N_VPWR_c_1775_n 0.0123247f $X=11.365 $Y=2.495
+ $X2=0 $Y2=0
cc_1033 N_A_2083_65#_M1004_g N_Q_c_2086_n 0.00310294f $X=13.375 $Y=0.705 $X2=0
+ $Y2=0
cc_1034 N_A_2083_65#_M1011_g Q 0.00498682f $X=13.345 $Y=2.465 $X2=0 $Y2=0
cc_1035 N_A_2083_65#_c_1421_n Q 7.47331e-19 $X=13.36 $Y=1.53 $X2=0 $Y2=0
cc_1036 N_A_2083_65#_M1026_g N_Q_c_2084_n 8.61087e-19 $X=12.385 $Y=0.495 $X2=0
+ $Y2=0
cc_1037 N_A_2083_65#_c_1416_n N_Q_c_2084_n 0.0192979f $X=13.27 $Y=1.53 $X2=0
+ $Y2=0
cc_1038 N_A_2083_65#_M1011_g N_Q_c_2084_n 0.012209f $X=13.345 $Y=2.465 $X2=0
+ $Y2=0
cc_1039 N_A_2083_65#_M1004_g N_Q_c_2084_n 0.0248646f $X=13.375 $Y=0.705 $X2=0
+ $Y2=0
cc_1040 N_A_2083_65#_c_1421_n N_Q_c_2084_n 0.00213235f $X=13.36 $Y=1.53 $X2=0
+ $Y2=0
cc_1041 N_A_2083_65#_M1011_g N_Q_N_c_2128_n 0.00107114f $X=13.345 $Y=2.465 $X2=0
+ $Y2=0
cc_1042 N_A_2083_65#_M1004_g N_Q_N_c_2126_n 5.88656e-19 $X=13.375 $Y=0.705 $X2=0
+ $Y2=0
cc_1043 N_A_2083_65#_c_1419_n N_VGND_c_2175_n 0.00827139f $X=10.492 $Y=0.985
+ $X2=0 $Y2=0
cc_1044 N_A_2083_65#_c_1424_n N_VGND_c_2175_n 0.018067f $X=11.61 $Y=0.58 $X2=0
+ $Y2=0
cc_1045 N_A_2083_65#_M1026_g N_VGND_c_2176_n 0.00533583f $X=12.385 $Y=0.495
+ $X2=0 $Y2=0
cc_1046 N_A_2083_65#_c_1424_n N_VGND_c_2176_n 0.0303742f $X=11.61 $Y=0.58 $X2=0
+ $Y2=0
cc_1047 N_A_2083_65#_M1004_g N_VGND_c_2177_n 0.00368477f $X=13.375 $Y=0.705
+ $X2=0 $Y2=0
cc_1048 N_A_2083_65#_M1026_g N_VGND_c_2182_n 0.00502664f $X=12.385 $Y=0.495
+ $X2=0 $Y2=0
cc_1049 N_A_2083_65#_M1004_g N_VGND_c_2182_n 0.00502664f $X=13.375 $Y=0.705
+ $X2=0 $Y2=0
cc_1050 N_A_2083_65#_c_1419_n N_VGND_c_2187_n 0.00517164f $X=10.492 $Y=0.985
+ $X2=0 $Y2=0
cc_1051 N_A_2083_65#_c_1424_n N_VGND_c_2188_n 0.0197885f $X=11.61 $Y=0.58 $X2=0
+ $Y2=0
cc_1052 N_A_2083_65#_M1003_d N_VGND_c_2190_n 0.00232985f $X=11.47 $Y=0.235 $X2=0
+ $Y2=0
cc_1053 N_A_2083_65#_M1026_g N_VGND_c_2190_n 0.011218f $X=12.385 $Y=0.495 $X2=0
+ $Y2=0
cc_1054 N_A_2083_65#_M1004_g N_VGND_c_2190_n 0.0104609f $X=13.375 $Y=0.705 $X2=0
+ $Y2=0
cc_1055 N_A_2083_65#_c_1419_n N_VGND_c_2190_n 0.00519032f $X=10.492 $Y=0.985
+ $X2=0 $Y2=0
cc_1056 N_A_2083_65#_c_1424_n N_VGND_c_2190_n 0.0125808f $X=11.61 $Y=0.58 $X2=0
+ $Y2=0
cc_1057 N_A_1903_125#_c_1594_n N_VPWR_c_1781_n 0.0219664f $X=9.805 $Y=2.19 $X2=0
+ $Y2=0
cc_1058 N_A_1903_125#_M1015_g N_VPWR_c_1782_n 0.0109329f $X=11.15 $Y=2.675 $X2=0
+ $Y2=0
cc_1059 N_A_1903_125#_M1015_g N_VPWR_c_1783_n 0.00549284f $X=11.15 $Y=2.675
+ $X2=0 $Y2=0
cc_1060 N_A_1903_125#_c_1594_n N_VPWR_c_1799_n 0.0111657f $X=9.805 $Y=2.19 $X2=0
+ $Y2=0
cc_1061 N_A_1903_125#_M1015_g N_VPWR_c_1775_n 0.0075526f $X=11.15 $Y=2.675 $X2=0
+ $Y2=0
cc_1062 N_A_1903_125#_c_1594_n N_VPWR_c_1775_n 0.0114323f $X=9.805 $Y=2.19 $X2=0
+ $Y2=0
cc_1063 N_A_1903_125#_c_1585_n N_VGND_c_2175_n 0.0182963f $X=10.945 $Y=0.985
+ $X2=0 $Y2=0
cc_1064 N_A_1903_125#_c_1588_n N_VGND_c_2175_n 0.0107144f $X=9.77 $Y=0.6 $X2=0
+ $Y2=0
cc_1065 N_A_1903_125#_c_1591_n N_VGND_c_2175_n 0.00442171f $X=10.945 $Y=1.15
+ $X2=0 $Y2=0
cc_1066 N_A_1903_125#_c_1592_n N_VGND_c_2175_n 0.0233988f $X=10.78 $Y=1.13 $X2=0
+ $Y2=0
cc_1067 N_A_1903_125#_c_1588_n N_VGND_c_2187_n 0.0144759f $X=9.77 $Y=0.6 $X2=0
+ $Y2=0
cc_1068 N_A_1903_125#_c_1585_n N_VGND_c_2188_n 0.00486043f $X=10.945 $Y=0.985
+ $X2=0 $Y2=0
cc_1069 N_A_1903_125#_c_1585_n N_VGND_c_2190_n 0.00818711f $X=10.945 $Y=0.985
+ $X2=0 $Y2=0
cc_1070 N_A_1903_125#_c_1588_n N_VGND_c_2190_n 0.0135253f $X=9.77 $Y=0.6 $X2=0
+ $Y2=0
cc_1071 N_A_2456_451#_c_1684_n N_VPWR_M1011_d 0.00489995f $X=13.555 $Y=2.41
+ $X2=0 $Y2=0
cc_1072 N_A_2456_451#_c_1678_n N_VPWR_M1011_d 0.00850272f $X=13.64 $Y=2.325
+ $X2=0 $Y2=0
cc_1073 N_A_2456_451#_c_1686_n N_VPWR_c_1784_n 0.0272489f $X=12.42 $Y=2.4 $X2=0
+ $Y2=0
cc_1074 N_A_2456_451#_c_1687_n N_VPWR_c_1784_n 0.0149774f $X=12.78 $Y=2.365
+ $X2=0 $Y2=0
cc_1075 N_A_2456_451#_M1014_g N_VPWR_c_1785_n 0.00521498f $X=13.855 $Y=2.465
+ $X2=0 $Y2=0
cc_1076 N_A_2456_451#_c_1684_n N_VPWR_c_1785_n 0.0209079f $X=13.555 $Y=2.41
+ $X2=0 $Y2=0
cc_1077 N_A_2456_451#_c_1686_n N_VPWR_c_1796_n 0.0111416f $X=12.42 $Y=2.4 $X2=0
+ $Y2=0
cc_1078 N_A_2456_451#_M1014_g N_VPWR_c_1800_n 0.00549284f $X=13.855 $Y=2.465
+ $X2=0 $Y2=0
cc_1079 N_A_2456_451#_M1014_g N_VPWR_c_1775_n 0.011115f $X=13.855 $Y=2.465 $X2=0
+ $Y2=0
cc_1080 N_A_2456_451#_c_1684_n N_VPWR_c_1775_n 0.00114993f $X=13.555 $Y=2.41
+ $X2=0 $Y2=0
cc_1081 N_A_2456_451#_c_1686_n N_VPWR_c_1775_n 0.0114016f $X=12.42 $Y=2.4 $X2=0
+ $Y2=0
cc_1082 N_A_2456_451#_c_1687_n N_VPWR_c_1775_n 0.0275472f $X=12.78 $Y=2.365
+ $X2=0 $Y2=0
cc_1083 N_A_2456_451#_c_1684_n N_Q_M1011_s 0.00795069f $X=13.555 $Y=2.41 $X2=0
+ $Y2=0
cc_1084 N_A_2456_451#_c_1677_n N_Q_c_2095_n 0.00354781f $X=12.695 $Y=2.235 $X2=0
+ $Y2=0
cc_1085 N_A_2456_451#_c_1678_n N_Q_c_2095_n 0.00203796f $X=13.64 $Y=2.325 $X2=0
+ $Y2=0
cc_1086 N_A_2456_451#_c_1680_n N_Q_c_2095_n 0.00174554f $X=13.825 $Y=1.49 $X2=0
+ $Y2=0
cc_1087 N_A_2456_451#_M1016_g N_Q_c_2086_n 3.01349e-19 $X=13.885 $Y=0.705 $X2=0
+ $Y2=0
cc_1088 N_A_2456_451#_c_1677_n N_Q_c_2086_n 0.00137447f $X=12.695 $Y=2.235 $X2=0
+ $Y2=0
cc_1089 N_A_2456_451#_c_1680_n N_Q_c_2086_n 0.00143394f $X=13.825 $Y=1.49 $X2=0
+ $Y2=0
cc_1090 N_A_2456_451#_c_1684_n N_Q_c_2101_n 0.00125447f $X=13.555 $Y=2.41 $X2=0
+ $Y2=0
cc_1091 N_A_2456_451#_M1014_g Q 9.97718e-19 $X=13.855 $Y=2.465 $X2=0 $Y2=0
cc_1092 N_A_2456_451#_c_1684_n Q 0.00925086f $X=13.555 $Y=2.41 $X2=0 $Y2=0
cc_1093 N_A_2456_451#_c_1678_n Q 0.0103002f $X=13.64 $Y=2.325 $X2=0 $Y2=0
cc_1094 N_A_2456_451#_c_1680_n Q 0.0020906f $X=13.825 $Y=1.49 $X2=0 $Y2=0
cc_1095 N_A_2456_451#_c_1681_n Q 8.91972e-19 $X=13.825 $Y=1.49 $X2=0 $Y2=0
cc_1096 N_A_2456_451#_M1016_g N_Q_c_2084_n 0.00142519f $X=13.885 $Y=0.705 $X2=0
+ $Y2=0
cc_1097 N_A_2456_451#_c_1684_n N_Q_c_2084_n 0.022339f $X=13.555 $Y=2.41 $X2=0
+ $Y2=0
cc_1098 N_A_2456_451#_c_1678_n N_Q_c_2084_n 0.0254743f $X=13.64 $Y=2.325 $X2=0
+ $Y2=0
cc_1099 N_A_2456_451#_c_1679_n N_Q_c_2084_n 0.137253f $X=12.6 $Y=0.495 $X2=0
+ $Y2=0
cc_1100 N_A_2456_451#_c_1680_n N_Q_c_2084_n 0.0178517f $X=13.825 $Y=1.49 $X2=0
+ $Y2=0
cc_1101 N_A_2456_451#_c_1681_n N_Q_c_2084_n 3.3588e-19 $X=13.825 $Y=1.49 $X2=0
+ $Y2=0
cc_1102 N_A_2456_451#_M1014_g N_Q_N_c_2128_n 0.0151652f $X=13.855 $Y=2.465 $X2=0
+ $Y2=0
cc_1103 N_A_2456_451#_M1016_g N_Q_N_c_2123_n 0.0111798f $X=13.885 $Y=0.705 $X2=0
+ $Y2=0
cc_1104 N_A_2456_451#_M1016_g N_Q_N_c_2124_n 0.0026953f $X=13.885 $Y=0.705 $X2=0
+ $Y2=0
cc_1105 N_A_2456_451#_c_1680_n N_Q_N_c_2124_n 0.00147869f $X=13.825 $Y=1.49
+ $X2=0 $Y2=0
cc_1106 N_A_2456_451#_c_1681_n N_Q_N_c_2124_n 0.00115575f $X=13.825 $Y=1.49
+ $X2=0 $Y2=0
cc_1107 N_A_2456_451#_M1014_g N_Q_N_c_2125_n 0.00381435f $X=13.855 $Y=2.465
+ $X2=0 $Y2=0
cc_1108 N_A_2456_451#_c_1678_n N_Q_N_c_2125_n 0.00529764f $X=13.64 $Y=2.325
+ $X2=0 $Y2=0
cc_1109 N_A_2456_451#_c_1680_n N_Q_N_c_2125_n 0.00767639f $X=13.825 $Y=1.49
+ $X2=0 $Y2=0
cc_1110 N_A_2456_451#_c_1681_n N_Q_N_c_2125_n 0.00728458f $X=13.825 $Y=1.49
+ $X2=0 $Y2=0
cc_1111 N_A_2456_451#_c_1678_n N_Q_N_c_2143_n 6.44547e-19 $X=13.64 $Y=2.325
+ $X2=0 $Y2=0
cc_1112 N_A_2456_451#_M1016_g N_Q_N_c_2126_n 0.00692296f $X=13.885 $Y=0.705
+ $X2=0 $Y2=0
cc_1113 N_A_2456_451#_c_1678_n N_Q_N_c_2126_n 4.44926e-19 $X=13.64 $Y=2.325
+ $X2=0 $Y2=0
cc_1114 N_A_2456_451#_c_1680_n N_Q_N_c_2126_n 0.0171136f $X=13.825 $Y=1.49 $X2=0
+ $Y2=0
cc_1115 N_A_2456_451#_c_1681_n N_Q_N_c_2126_n 0.0025683f $X=13.825 $Y=1.49 $X2=0
+ $Y2=0
cc_1116 N_A_2456_451#_M1014_g N_Q_N_c_2130_n 0.0024291f $X=13.855 $Y=2.465 $X2=0
+ $Y2=0
cc_1117 N_A_2456_451#_c_1678_n N_Q_N_c_2130_n 0.0192938f $X=13.64 $Y=2.325 $X2=0
+ $Y2=0
cc_1118 N_A_2456_451#_c_1680_n N_Q_N_c_2130_n 0.00278627f $X=13.825 $Y=1.49
+ $X2=0 $Y2=0
cc_1119 N_A_2456_451#_c_1681_n N_Q_N_c_2130_n 0.00139072f $X=13.825 $Y=1.49
+ $X2=0 $Y2=0
cc_1120 N_A_2456_451#_M1014_g N_Q_N_c_2127_n 0.00253526f $X=13.855 $Y=2.465
+ $X2=0 $Y2=0
cc_1121 N_A_2456_451#_M1016_g N_Q_N_c_2127_n 0.00366557f $X=13.885 $Y=0.705
+ $X2=0 $Y2=0
cc_1122 N_A_2456_451#_c_1678_n N_Q_N_c_2127_n 0.00339775f $X=13.64 $Y=2.325
+ $X2=0 $Y2=0
cc_1123 N_A_2456_451#_c_1680_n N_Q_N_c_2127_n 0.0205721f $X=13.825 $Y=1.49 $X2=0
+ $Y2=0
cc_1124 N_A_2456_451#_c_1681_n N_Q_N_c_2127_n 0.00726364f $X=13.825 $Y=1.49
+ $X2=0 $Y2=0
cc_1125 N_A_2456_451#_c_1679_n N_VGND_c_2176_n 0.0180555f $X=12.6 $Y=0.495 $X2=0
+ $Y2=0
cc_1126 N_A_2456_451#_M1016_g N_VGND_c_2177_n 0.00724214f $X=13.885 $Y=0.705
+ $X2=0 $Y2=0
cc_1127 N_A_2456_451#_c_1680_n N_VGND_c_2177_n 0.0139708f $X=13.825 $Y=1.49
+ $X2=0 $Y2=0
cc_1128 N_A_2456_451#_c_1681_n N_VGND_c_2177_n 0.00166772f $X=13.825 $Y=1.49
+ $X2=0 $Y2=0
cc_1129 N_A_2456_451#_c_1679_n N_VGND_c_2182_n 0.0227108f $X=12.6 $Y=0.495 $X2=0
+ $Y2=0
cc_1130 N_A_2456_451#_M1016_g N_VGND_c_2189_n 0.00502664f $X=13.885 $Y=0.705
+ $X2=0 $Y2=0
cc_1131 N_A_2456_451#_M1016_g N_VGND_c_2190_n 0.0102315f $X=13.885 $Y=0.705
+ $X2=0 $Y2=0
cc_1132 N_A_2456_451#_c_1679_n N_VGND_c_2190_n 0.0130919f $X=12.6 $Y=0.495 $X2=0
+ $Y2=0
cc_1133 N_VPWR_c_1792_n N_A_636_531#_c_1971_n 0.00570423f $X=6.57 $Y=3.33 $X2=0
+ $Y2=0
cc_1134 N_VPWR_c_1775_n N_A_636_531#_c_1971_n 0.0068754f $X=14.16 $Y=3.33 $X2=0
+ $Y2=0
cc_1135 N_VPWR_c_1790_n N_A_636_531#_c_1975_n 0.0248505f $X=4.215 $Y=3.33 $X2=0
+ $Y2=0
cc_1136 N_VPWR_c_1775_n N_A_636_531#_c_1975_n 0.0191634f $X=14.16 $Y=3.33 $X2=0
+ $Y2=0
cc_1137 N_VPWR_c_1775_n N_Q_M1011_s 0.00419625f $X=14.16 $Y=3.33 $X2=0 $Y2=0
cc_1138 N_VPWR_M1011_d Q 0.00838058f $X=13.42 $Y=1.835 $X2=0 $Y2=0
cc_1139 N_VPWR_c_1785_n Q 0.00100968f $X=13.56 $Y=2.895 $X2=0 $Y2=0
cc_1140 N_VPWR_c_1775_n N_Q_N_M1014_d 0.0023218f $X=14.16 $Y=3.33 $X2=0 $Y2=0
cc_1141 N_VPWR_c_1800_n N_Q_N_c_2128_n 0.0248149f $X=14.16 $Y=3.33 $X2=0 $Y2=0
cc_1142 N_VPWR_c_1775_n N_Q_N_c_2128_n 0.01541f $X=14.16 $Y=3.33 $X2=0 $Y2=0
cc_1143 N_A_636_531#_c_1965_n N_VGND_M1039_d 0.00183001f $X=5.375 $Y=0.555 $X2=0
+ $Y2=0
cc_1144 N_A_636_531#_c_1966_n N_VGND_c_2171_n 0.00105387f $X=3.745 $Y=0.555
+ $X2=0 $Y2=0
cc_1145 N_A_636_531#_c_1967_n N_VGND_c_2171_n 0.0162475f $X=3.6 $Y=0.555 $X2=0
+ $Y2=0
cc_1146 N_A_636_531#_c_1965_n N_VGND_c_2172_n 0.018244f $X=5.375 $Y=0.555 $X2=0
+ $Y2=0
cc_1147 N_A_636_531#_c_1965_n N_VGND_c_2180_n 0.00203161f $X=5.375 $Y=0.555
+ $X2=0 $Y2=0
cc_1148 N_A_636_531#_c_1968_n N_VGND_c_2180_n 9.72113e-19 $X=5.52 $Y=0.555 $X2=0
+ $Y2=0
cc_1149 N_A_636_531#_c_1969_n N_VGND_c_2180_n 0.0206756f $X=5.955 $Y=0.737 $X2=0
+ $Y2=0
cc_1150 N_A_636_531#_c_1965_n N_VGND_c_2185_n 0.00188203f $X=5.375 $Y=0.555
+ $X2=0 $Y2=0
cc_1151 N_A_636_531#_c_1966_n N_VGND_c_2185_n 3.39548e-19 $X=3.745 $Y=0.555
+ $X2=0 $Y2=0
cc_1152 N_A_636_531#_c_1967_n N_VGND_c_2185_n 0.0294816f $X=3.6 $Y=0.555 $X2=0
+ $Y2=0
cc_1153 N_A_636_531#_M1036_d N_VGND_c_2190_n 0.00204599f $X=3.25 $Y=0.235 $X2=0
+ $Y2=0
cc_1154 N_A_636_531#_c_1965_n N_VGND_c_2190_n 0.127104f $X=5.375 $Y=0.555 $X2=0
+ $Y2=0
cc_1155 N_A_636_531#_c_1966_n N_VGND_c_2190_n 0.0257798f $X=3.745 $Y=0.555 $X2=0
+ $Y2=0
cc_1156 N_A_636_531#_c_1967_n N_VGND_c_2190_n 0.011368f $X=3.6 $Y=0.555 $X2=0
+ $Y2=0
cc_1157 N_A_636_531#_c_1968_n N_VGND_c_2190_n 0.0272763f $X=5.52 $Y=0.555 $X2=0
+ $Y2=0
cc_1158 N_A_636_531#_c_1969_n N_VGND_c_2190_n 0.013362f $X=5.955 $Y=0.737 $X2=0
+ $Y2=0
cc_1159 Q N_Q_N_c_2143_n 0.0111805f $X=13.595 $Y=1.965 $X2=0 $Y2=0
cc_1160 N_Q_c_2086_n N_Q_N_c_2126_n 0.0116635f $X=13.2 $Y=1.295 $X2=0 $Y2=0
cc_1161 N_Q_c_2084_n N_Q_N_c_2126_n 0.00173764f $X=13.16 $Y=0.43 $X2=0 $Y2=0
cc_1162 Q N_Q_N_c_2130_n 0.00125449f $X=13.595 $Y=1.965 $X2=0 $Y2=0
cc_1163 N_Q_c_2084_n N_VGND_c_2177_n 0.0334192f $X=13.16 $Y=0.43 $X2=0 $Y2=0
cc_1164 N_Q_c_2084_n N_VGND_c_2182_n 0.0240548f $X=13.16 $Y=0.43 $X2=0 $Y2=0
cc_1165 N_Q_c_2084_n N_VGND_c_2190_n 0.0137416f $X=13.16 $Y=0.43 $X2=0 $Y2=0
cc_1166 N_Q_N_c_2123_n N_VGND_c_2177_n 0.0335829f $X=14.1 $Y=0.43 $X2=0 $Y2=0
cc_1167 N_Q_N_c_2126_n N_VGND_c_2177_n 0.00465703f $X=14.09 $Y=1.295 $X2=0 $Y2=0
cc_1168 N_Q_N_c_2123_n N_VGND_c_2189_n 0.0250662f $X=14.1 $Y=0.43 $X2=0 $Y2=0
cc_1169 N_Q_N_c_2123_n N_VGND_c_2190_n 0.014322f $X=14.1 $Y=0.43 $X2=0 $Y2=0
cc_1170 N_VGND_c_2190_n A_312_47# 0.010279f $X=14.16 $Y=0 $X2=-0.19 $Y2=-0.245
cc_1171 N_VGND_c_2190_n A_486_47# 0.00357508f $X=14.16 $Y=0 $X2=-0.19 $Y2=-0.245
cc_1172 N_VGND_c_2190_n A_2222_47# 0.00899413f $X=14.16 $Y=0 $X2=-0.19
+ $Y2=-0.245
