* NGSPICE file created from sky130_fd_sc_lp__and2b_2.ext - technology: sky130A

.subckt sky130_fd_sc_lp__and2b_2 A_N B VGND VNB VPB VPWR X
M1000 VPWR a_186_239# X VPB phighvt w=1.26e+06u l=150000u
+  ad=9.429e+11p pd=8.25e+06u as=3.528e+11p ps=3.08e+06u
M1001 X a_186_239# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1002 VGND a_186_239# X VNB nshort w=840000u l=150000u
+  ad=7.4e+11p pd=5.56e+06u as=2.352e+11p ps=2.24e+06u
M1003 a_186_239# B VPWR VPB phighvt w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=0p ps=0u
M1004 VGND A_N a_28_367# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1005 a_186_239# a_28_367# a_455_133# VNB nshort w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=8.82e+10p ps=1.26e+06u
M1006 VPWR A_N a_28_367# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1007 VPWR a_28_367# a_186_239# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 X a_186_239# VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_455_133# B VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

