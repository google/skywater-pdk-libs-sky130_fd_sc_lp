* File: sky130_fd_sc_lp__a2bb2oi_m.pxi.spice
* Created: Fri Aug 28 09:57:08 2020
* 
x_PM_SKY130_FD_SC_LP__A2BB2OI_M%A1_N N_A1_N_c_76_n N_A1_N_c_84_n N_A1_N_c_85_n
+ N_A1_N_c_77_n N_A1_N_c_78_n N_A1_N_M1007_g N_A1_N_c_79_n N_A1_N_M1005_g
+ N_A1_N_c_80_n A1_N A1_N A1_N A1_N A1_N A1_N N_A1_N_c_82_n
+ PM_SKY130_FD_SC_LP__A2BB2OI_M%A1_N
x_PM_SKY130_FD_SC_LP__A2BB2OI_M%A2_N N_A2_N_M1002_g N_A2_N_c_122_n
+ N_A2_N_c_123_n N_A2_N_M1000_g N_A2_N_c_125_n A2_N A2_N A2_N A2_N A2_N A2_N
+ N_A2_N_c_127_n PM_SKY130_FD_SC_LP__A2BB2OI_M%A2_N
x_PM_SKY130_FD_SC_LP__A2BB2OI_M%A_202_47# N_A_202_47#_M1005_d
+ N_A_202_47#_M1002_d N_A_202_47#_c_178_n N_A_202_47#_c_179_n
+ N_A_202_47#_c_180_n N_A_202_47#_c_173_n N_A_202_47#_c_174_n
+ N_A_202_47#_M1001_g N_A_202_47#_c_182_n N_A_202_47#_M1006_g
+ N_A_202_47#_c_183_n N_A_202_47#_c_176_n N_A_202_47#_c_177_n
+ N_A_202_47#_c_185_n N_A_202_47#_c_186_n
+ PM_SKY130_FD_SC_LP__A2BB2OI_M%A_202_47#
x_PM_SKY130_FD_SC_LP__A2BB2OI_M%B2 N_B2_M1008_g N_B2_M1003_g N_B2_c_239_n
+ N_B2_c_240_n N_B2_c_241_n B2 B2 N_B2_c_243_n PM_SKY130_FD_SC_LP__A2BB2OI_M%B2
x_PM_SKY130_FD_SC_LP__A2BB2OI_M%B1 N_B1_M1004_g N_B1_M1009_g N_B1_c_283_n
+ N_B1_c_284_n N_B1_c_285_n B1 B1 N_B1_c_287_n PM_SKY130_FD_SC_LP__A2BB2OI_M%B1
x_PM_SKY130_FD_SC_LP__A2BB2OI_M%VPWR N_VPWR_M1007_s N_VPWR_M1003_d
+ N_VPWR_c_314_n N_VPWR_c_315_n N_VPWR_c_316_n VPWR N_VPWR_c_317_n
+ N_VPWR_c_318_n N_VPWR_c_313_n N_VPWR_c_320_n
+ PM_SKY130_FD_SC_LP__A2BB2OI_M%VPWR
x_PM_SKY130_FD_SC_LP__A2BB2OI_M%Y N_Y_M1001_d N_Y_M1006_s N_Y_c_346_n
+ N_Y_c_347_n N_Y_c_359_n Y PM_SKY130_FD_SC_LP__A2BB2OI_M%Y
x_PM_SKY130_FD_SC_LP__A2BB2OI_M%A_403_387# N_A_403_387#_M1006_d
+ N_A_403_387#_M1009_d N_A_403_387#_c_389_n N_A_403_387#_c_385_n
+ N_A_403_387#_c_386_n N_A_403_387#_c_387_n
+ PM_SKY130_FD_SC_LP__A2BB2OI_M%A_403_387#
x_PM_SKY130_FD_SC_LP__A2BB2OI_M%VGND N_VGND_M1005_s N_VGND_M1000_d
+ N_VGND_M1004_d N_VGND_c_402_n N_VGND_c_403_n N_VGND_c_404_n N_VGND_c_405_n
+ N_VGND_c_406_n N_VGND_c_407_n VGND N_VGND_c_408_n N_VGND_c_409_n
+ N_VGND_c_410_n N_VGND_c_411_n PM_SKY130_FD_SC_LP__A2BB2OI_M%VGND
cc_1 VNB N_A1_N_c_76_n 0.017584f $X=-0.19 $Y=-0.245 $X2=0.18 $Y2=2.065
cc_2 VNB N_A1_N_c_77_n 0.0376441f $X=-0.19 $Y=-0.245 $X2=0.86 $Y2=0.84
cc_3 VNB N_A1_N_c_78_n 0.0240808f $X=-0.19 $Y=-0.245 $X2=0.435 $Y2=0.84
cc_4 VNB N_A1_N_c_79_n 0.0193697f $X=-0.19 $Y=-0.245 $X2=0.935 $Y2=0.765
cc_5 VNB N_A1_N_c_80_n 0.0215434f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.435
cc_6 VNB A1_N 0.0187093f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.47
cc_7 VNB N_A1_N_c_82_n 0.0381518f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=0.93
cc_8 VNB N_A2_N_c_122_n 0.033781f $X=-0.19 $Y=-0.245 $X2=0.86 $Y2=0.84
cc_9 VNB N_A2_N_c_123_n 0.0130616f $X=-0.19 $Y=-0.245 $X2=0.435 $Y2=0.84
cc_10 VNB N_A2_N_M1000_g 0.0390038f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=2.795
cc_11 VNB N_A2_N_c_125_n 0.0014849f $X=-0.19 $Y=-0.245 $X2=0.935 $Y2=0.445
cc_12 VNB A2_N 0.00720045f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=0.915
cc_13 VNB N_A2_N_c_127_n 0.0270736f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_202_47#_c_173_n 0.00627889f $X=-0.19 $Y=-0.245 $X2=0.935 $Y2=0.765
cc_15 VNB N_A_202_47#_c_174_n 0.00822778f $X=-0.19 $Y=-0.245 $X2=0.935 $Y2=0.445
cc_16 VNB N_A_202_47#_M1001_g 0.048511f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.27
cc_17 VNB N_A_202_47#_c_176_n 0.0171699f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_202_47#_c_177_n 4.40119e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_B2_M1003_g 0.0126593f $X=-0.19 $Y=-0.245 $X2=0.435 $Y2=0.84
cc_20 VNB N_B2_c_239_n 0.0170155f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=2.795
cc_21 VNB N_B2_c_240_n 0.0229352f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_B2_c_241_n 0.0158934f $X=-0.19 $Y=-0.245 $X2=0.935 $Y2=0.765
cc_23 VNB B2 0.0150123f $X=-0.19 $Y=-0.245 $X2=0.935 $Y2=0.445
cc_24 VNB N_B2_c_243_n 0.015247f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.47
cc_25 VNB N_B1_M1009_g 0.0179962f $X=-0.19 $Y=-0.245 $X2=0.435 $Y2=0.84
cc_26 VNB N_B1_c_283_n 0.0218131f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=2.795
cc_27 VNB N_B1_c_284_n 0.0273299f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_B1_c_285_n 0.0237174f $X=-0.19 $Y=-0.245 $X2=0.935 $Y2=0.445
cc_29 VNB B1 0.0342382f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=0.915
cc_30 VNB N_B1_c_287_n 0.0323097f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_31 VNB N_VPWR_c_313_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_Y_c_346_n 0.00508628f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=2.795
cc_33 VNB N_Y_c_347_n 0.0104704f $X=-0.19 $Y=-0.245 $X2=0.935 $Y2=0.445
cc_34 VNB Y 0.00112415f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_35 VNB N_VGND_c_402_n 0.0123699f $X=-0.19 $Y=-0.245 $X2=0.935 $Y2=0.445
cc_36 VNB N_VGND_c_403_n 0.00425268f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.435
cc_37 VNB N_VGND_c_404_n 0.0149546f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_38 VNB N_VGND_c_405_n 0.0125783f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_39 VNB N_VGND_c_406_n 0.0165299f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_407_n 0.00362723f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_408_n 0.0179462f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_409_n 0.0316561f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_410_n 0.00522083f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_411_n 0.197744f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VPB N_A1_N_c_76_n 0.0340869f $X=-0.19 $Y=1.655 $X2=0.18 $Y2=2.065
cc_46 VPB N_A1_N_c_84_n 0.031698f $X=-0.19 $Y=1.655 $X2=0.51 $Y2=2.14
cc_47 VPB N_A1_N_c_85_n 0.0154685f $X=-0.19 $Y=1.655 $X2=0.255 $Y2=2.14
cc_48 VPB N_A1_N_M1007_g 0.0325543f $X=-0.19 $Y=1.655 $X2=0.585 $Y2=2.795
cc_49 VPB A1_N 0.0176913f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.47
cc_50 VPB N_A2_N_M1002_g 0.0528973f $X=-0.19 $Y=1.655 $X2=0.51 $Y2=2.14
cc_51 VPB N_A2_N_c_125_n 0.0197612f $X=-0.19 $Y=1.655 $X2=0.935 $Y2=0.445
cc_52 VPB A2_N 0.0032884f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=0.915
cc_53 VPB N_A_202_47#_c_178_n 0.0493779f $X=-0.19 $Y=1.655 $X2=0.585 $Y2=2.795
cc_54 VPB N_A_202_47#_c_179_n 0.0138067f $X=-0.19 $Y=1.655 $X2=0.585 $Y2=2.795
cc_55 VPB N_A_202_47#_c_180_n 0.0119609f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_56 VPB N_A_202_47#_c_174_n 0.00125732f $X=-0.19 $Y=1.655 $X2=0.935 $Y2=0.445
cc_57 VPB N_A_202_47#_c_182_n 0.0195634f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.47
cc_58 VPB N_A_202_47#_c_183_n 0.0117753f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.95
cc_59 VPB N_A_202_47#_c_176_n 0.0193395f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_60 VPB N_A_202_47#_c_185_n 0.00595771f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_61 VPB N_A_202_47#_c_186_n 0.0498016f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_62 VPB N_B2_M1003_g 0.0255919f $X=-0.19 $Y=1.655 $X2=0.435 $Y2=0.84
cc_63 VPB N_B1_M1009_g 0.0345609f $X=-0.19 $Y=1.655 $X2=0.435 $Y2=0.84
cc_64 VPB N_VPWR_c_314_n 0.0125089f $X=-0.19 $Y=1.655 $X2=0.585 $Y2=2.215
cc_65 VPB N_VPWR_c_315_n 0.0209705f $X=-0.19 $Y=1.655 $X2=0.585 $Y2=2.795
cc_66 VPB N_VPWR_c_316_n 0.0487408f $X=-0.19 $Y=1.655 $X2=0.935 $Y2=0.445
cc_67 VPB N_VPWR_c_317_n 0.055591f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.47
cc_68 VPB N_VPWR_c_318_n 0.0215547f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_69 VPB N_VPWR_c_313_n 0.0967232f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_70 VPB N_VPWR_c_320_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_71 VPB Y 0.00416556f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_72 VPB N_A_403_387#_c_385_n 0.0194358f $X=-0.19 $Y=1.655 $X2=0.935 $Y2=0.765
cc_73 VPB N_A_403_387#_c_386_n 0.00535629f $X=-0.19 $Y=1.655 $X2=0.935 $Y2=0.445
cc_74 VPB N_A_403_387#_c_387_n 4.08405e-19 $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.27
cc_75 N_A1_N_c_76_n N_A2_N_M1002_g 0.00307633f $X=0.18 $Y=2.065 $X2=0 $Y2=0
cc_76 N_A1_N_c_84_n N_A2_N_M1002_g 0.0679956f $X=0.51 $Y=2.14 $X2=0 $Y2=0
cc_77 A1_N N_A2_N_M1002_g 7.15449e-19 $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_78 N_A1_N_c_77_n N_A2_N_c_123_n 0.0222683f $X=0.86 $Y=0.84 $X2=0 $Y2=0
cc_79 A1_N N_A2_N_c_123_n 3.0834e-19 $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_80 N_A1_N_c_82_n N_A2_N_c_123_n 0.00878425f $X=0.27 $Y=0.93 $X2=0 $Y2=0
cc_81 N_A1_N_c_79_n N_A2_N_M1000_g 0.0190745f $X=0.935 $Y=0.765 $X2=0 $Y2=0
cc_82 N_A1_N_c_84_n N_A2_N_c_125_n 8.31396e-19 $X=0.51 $Y=2.14 $X2=0 $Y2=0
cc_83 N_A1_N_c_76_n A2_N 0.00210492f $X=0.18 $Y=2.065 $X2=0 $Y2=0
cc_84 N_A1_N_c_84_n A2_N 0.00483066f $X=0.51 $Y=2.14 $X2=0 $Y2=0
cc_85 N_A1_N_c_77_n A2_N 0.00999259f $X=0.86 $Y=0.84 $X2=0 $Y2=0
cc_86 N_A1_N_M1007_g A2_N 0.0222401f $X=0.585 $Y=2.795 $X2=0 $Y2=0
cc_87 A1_N A2_N 0.0867533f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_88 N_A1_N_c_82_n A2_N 0.00735645f $X=0.27 $Y=0.93 $X2=0 $Y2=0
cc_89 N_A1_N_c_76_n N_A2_N_c_127_n 0.0112261f $X=0.18 $Y=2.065 $X2=0 $Y2=0
cc_90 N_A1_N_c_80_n N_A2_N_c_127_n 0.00878425f $X=0.27 $Y=1.435 $X2=0 $Y2=0
cc_91 A1_N N_A2_N_c_127_n 0.00143519f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_92 N_A1_N_c_79_n N_A_202_47#_c_176_n 0.00510427f $X=0.935 $Y=0.765 $X2=0
+ $Y2=0
cc_93 N_A1_N_c_84_n N_VPWR_c_315_n 0.0027446f $X=0.51 $Y=2.14 $X2=0 $Y2=0
cc_94 N_A1_N_c_85_n N_VPWR_c_315_n 0.00184964f $X=0.255 $Y=2.14 $X2=0 $Y2=0
cc_95 N_A1_N_M1007_g N_VPWR_c_315_n 0.00962334f $X=0.585 $Y=2.795 $X2=0 $Y2=0
cc_96 A1_N N_VPWR_c_315_n 0.0122248f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_97 N_A1_N_M1007_g N_VPWR_c_317_n 0.00473177f $X=0.585 $Y=2.795 $X2=0 $Y2=0
cc_98 N_A1_N_M1007_g N_VPWR_c_313_n 0.00928834f $X=0.585 $Y=2.795 $X2=0 $Y2=0
cc_99 A1_N N_VPWR_c_313_n 9.09196e-19 $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_100 N_A1_N_c_77_n N_VGND_c_402_n 0.00765496f $X=0.86 $Y=0.84 $X2=0 $Y2=0
cc_101 N_A1_N_c_79_n N_VGND_c_402_n 0.00729952f $X=0.935 $Y=0.765 $X2=0 $Y2=0
cc_102 A1_N N_VGND_c_402_n 0.00115588f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_103 N_A1_N_c_79_n N_VGND_c_406_n 0.00564095f $X=0.935 $Y=0.765 $X2=0 $Y2=0
cc_104 N_A1_N_c_78_n N_VGND_c_408_n 0.00467355f $X=0.435 $Y=0.84 $X2=0 $Y2=0
cc_105 A1_N N_VGND_c_408_n 0.0059365f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_106 N_A1_N_c_78_n N_VGND_c_411_n 0.0056437f $X=0.435 $Y=0.84 $X2=0 $Y2=0
cc_107 N_A1_N_c_79_n N_VGND_c_411_n 0.00872803f $X=0.935 $Y=0.765 $X2=0 $Y2=0
cc_108 A1_N N_VGND_c_411_n 0.00676397f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_109 N_A2_N_M1002_g N_A_202_47#_c_178_n 0.015976f $X=0.945 $Y=2.795 $X2=0
+ $Y2=0
cc_110 N_A2_N_c_122_n N_A_202_47#_c_180_n 0.00325335f $X=1.29 $Y=1.23 $X2=0
+ $Y2=0
cc_111 N_A2_N_c_125_n N_A_202_47#_c_180_n 0.015976f $X=0.832 $Y=1.825 $X2=0
+ $Y2=0
cc_112 N_A2_N_c_127_n N_A_202_47#_c_173_n 0.00111538f $X=0.81 $Y=1.32 $X2=0
+ $Y2=0
cc_113 N_A2_N_c_125_n N_A_202_47#_c_174_n 0.00111538f $X=0.832 $Y=1.825 $X2=0
+ $Y2=0
cc_114 N_A2_N_M1000_g N_A_202_47#_M1001_g 0.0321953f $X=1.365 $Y=0.445 $X2=0
+ $Y2=0
cc_115 N_A2_N_c_122_n N_A_202_47#_c_176_n 0.016408f $X=1.29 $Y=1.23 $X2=0 $Y2=0
cc_116 A2_N N_A_202_47#_c_176_n 0.128489f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_117 N_A2_N_c_127_n N_A_202_47#_c_176_n 0.0148012f $X=0.81 $Y=1.32 $X2=0 $Y2=0
cc_118 N_A2_N_c_122_n N_A_202_47#_c_177_n 7.66338e-19 $X=1.29 $Y=1.23 $X2=0
+ $Y2=0
cc_119 N_A2_N_M1000_g N_A_202_47#_c_177_n 0.0101892f $X=1.365 $Y=0.445 $X2=0
+ $Y2=0
cc_120 N_A2_N_M1002_g N_A_202_47#_c_185_n 3.00499e-19 $X=0.945 $Y=2.795 $X2=0
+ $Y2=0
cc_121 A2_N N_A_202_47#_c_186_n 3.718e-19 $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_122 N_A2_N_M1002_g N_VPWR_c_317_n 0.00473177f $X=0.945 $Y=2.795 $X2=0 $Y2=0
cc_123 A2_N N_VPWR_c_317_n 0.0058573f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_124 N_A2_N_M1002_g N_VPWR_c_313_n 0.00949399f $X=0.945 $Y=2.795 $X2=0 $Y2=0
cc_125 A2_N N_VPWR_c_313_n 0.00857257f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_126 A2_N A_132_517# 0.00139886f $X=0.635 $Y=0.84 $X2=-0.19 $Y2=-0.245
cc_127 N_A2_N_M1000_g N_Y_c_346_n 0.00250196f $X=1.365 $Y=0.445 $X2=0 $Y2=0
cc_128 N_A2_N_M1000_g N_VGND_c_402_n 6.9394e-19 $X=1.365 $Y=0.445 $X2=0 $Y2=0
cc_129 A2_N N_VGND_c_402_n 0.0083714f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_130 N_A2_N_M1000_g N_VGND_c_403_n 0.0015556f $X=1.365 $Y=0.445 $X2=0 $Y2=0
cc_131 N_A2_N_M1000_g N_VGND_c_406_n 0.00585385f $X=1.365 $Y=0.445 $X2=0 $Y2=0
cc_132 N_A2_N_M1000_g N_VGND_c_411_n 0.0108335f $X=1.365 $Y=0.445 $X2=0 $Y2=0
cc_133 A2_N N_VGND_c_411_n 0.00203126f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_134 N_A_202_47#_c_173_n N_B2_M1003_g 0.00689858f $X=1.815 $Y=1.525 $X2=0
+ $Y2=0
cc_135 N_A_202_47#_c_183_n N_B2_M1003_g 0.0211889f $X=1.87 $Y=1.75 $X2=0 $Y2=0
cc_136 N_A_202_47#_M1001_g N_B2_c_239_n 0.0133574f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_137 N_A_202_47#_M1001_g B2 6.00516e-19 $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_138 N_A_202_47#_M1001_g N_B2_c_243_n 0.0412537f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_139 N_A_202_47#_c_185_n N_VPWR_c_315_n 6.28954e-19 $X=1.61 $Y=2.86 $X2=0
+ $Y2=0
cc_140 N_A_202_47#_c_182_n N_VPWR_c_316_n 0.00114726f $X=1.94 $Y=1.825 $X2=0
+ $Y2=0
cc_141 N_A_202_47#_c_186_n N_VPWR_c_316_n 0.00834975f $X=1.61 $Y=2.86 $X2=0
+ $Y2=0
cc_142 N_A_202_47#_c_185_n N_VPWR_c_317_n 0.0308858f $X=1.61 $Y=2.86 $X2=0 $Y2=0
cc_143 N_A_202_47#_c_186_n N_VPWR_c_317_n 0.00983957f $X=1.61 $Y=2.86 $X2=0
+ $Y2=0
cc_144 N_A_202_47#_c_182_n N_VPWR_c_313_n 0.0038268f $X=1.94 $Y=1.825 $X2=0
+ $Y2=0
cc_145 N_A_202_47#_c_185_n N_VPWR_c_313_n 0.0227624f $X=1.61 $Y=2.86 $X2=0 $Y2=0
cc_146 N_A_202_47#_c_186_n N_VPWR_c_313_n 0.0130133f $X=1.61 $Y=2.86 $X2=0 $Y2=0
cc_147 N_A_202_47#_M1001_g N_Y_c_346_n 0.0215024f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_148 N_A_202_47#_c_177_n N_Y_c_346_n 0.0216132f $X=1.15 $Y=0.495 $X2=0 $Y2=0
cc_149 N_A_202_47#_c_179_n N_Y_c_347_n 8.47438e-19 $X=1.725 $Y=1.75 $X2=0 $Y2=0
cc_150 N_A_202_47#_c_173_n N_Y_c_347_n 0.00396515f $X=1.815 $Y=1.525 $X2=0 $Y2=0
cc_151 N_A_202_47#_c_174_n N_Y_c_347_n 0.00557223f $X=1.815 $Y=1.675 $X2=0 $Y2=0
cc_152 N_A_202_47#_M1001_g N_Y_c_347_n 0.00522793f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_153 N_A_202_47#_c_183_n N_Y_c_347_n 0.00492656f $X=1.87 $Y=1.75 $X2=0 $Y2=0
cc_154 N_A_202_47#_c_176_n N_Y_c_347_n 0.00866886f $X=1.17 $Y=2.695 $X2=0 $Y2=0
cc_155 N_A_202_47#_M1001_g N_Y_c_359_n 0.00397125f $X=1.83 $Y=0.445 $X2=0 $Y2=0
cc_156 N_A_202_47#_c_178_n Y 0.00332229f $X=1.45 $Y=2.695 $X2=0 $Y2=0
cc_157 N_A_202_47#_c_179_n Y 0.00835565f $X=1.725 $Y=1.75 $X2=0 $Y2=0
cc_158 N_A_202_47#_c_174_n Y 0.0042305f $X=1.815 $Y=1.675 $X2=0 $Y2=0
cc_159 N_A_202_47#_c_182_n Y 0.00227501f $X=1.94 $Y=1.825 $X2=0 $Y2=0
cc_160 N_A_202_47#_c_183_n Y 0.00461176f $X=1.87 $Y=1.75 $X2=0 $Y2=0
cc_161 N_A_202_47#_c_176_n Y 0.032276f $X=1.17 $Y=2.695 $X2=0 $Y2=0
cc_162 N_A_202_47#_c_185_n Y 0.00385411f $X=1.61 $Y=2.86 $X2=0 $Y2=0
cc_163 N_A_202_47#_c_186_n Y 0.00454239f $X=1.61 $Y=2.86 $X2=0 $Y2=0
cc_164 N_A_202_47#_c_183_n N_A_403_387#_c_386_n 0.00172956f $X=1.87 $Y=1.75
+ $X2=0 $Y2=0
cc_165 N_A_202_47#_M1001_g N_VGND_c_403_n 0.00571639f $X=1.83 $Y=0.445 $X2=0
+ $Y2=0
cc_166 N_A_202_47#_c_177_n N_VGND_c_406_n 0.0091159f $X=1.15 $Y=0.495 $X2=0
+ $Y2=0
cc_167 N_A_202_47#_M1001_g N_VGND_c_409_n 0.00503909f $X=1.83 $Y=0.445 $X2=0
+ $Y2=0
cc_168 N_A_202_47#_M1005_d N_VGND_c_411_n 0.00445618f $X=1.01 $Y=0.235 $X2=0
+ $Y2=0
cc_169 N_A_202_47#_M1001_g N_VGND_c_411_n 0.00878501f $X=1.83 $Y=0.445 $X2=0
+ $Y2=0
cc_170 N_A_202_47#_c_177_n N_VGND_c_411_n 0.008123f $X=1.15 $Y=0.495 $X2=0 $Y2=0
cc_171 N_B2_M1003_g N_B1_M1009_g 0.0199797f $X=2.37 $Y=2.145 $X2=0 $Y2=0
cc_172 N_B2_c_239_n N_B1_c_283_n 0.0264348f $X=2.28 $Y=0.765 $X2=0 $Y2=0
cc_173 B2 N_B1_c_284_n 0.00788111f $X=2.555 $Y=0.84 $X2=0 $Y2=0
cc_174 N_B2_c_243_n N_B1_c_284_n 0.0097538f $X=2.28 $Y=0.93 $X2=0 $Y2=0
cc_175 N_B2_c_241_n N_B1_c_285_n 0.0199797f $X=2.28 $Y=1.435 $X2=0 $Y2=0
cc_176 B2 N_B1_c_285_n 0.00154284f $X=2.555 $Y=0.84 $X2=0 $Y2=0
cc_177 B2 B1 0.0516964f $X=2.555 $Y=0.84 $X2=0 $Y2=0
cc_178 N_B2_c_243_n B1 4.53546e-19 $X=2.28 $Y=0.93 $X2=0 $Y2=0
cc_179 B2 N_B1_c_287_n 0.00355507f $X=2.555 $Y=0.84 $X2=0 $Y2=0
cc_180 N_B2_c_243_n N_B1_c_287_n 0.011053f $X=2.28 $Y=0.93 $X2=0 $Y2=0
cc_181 N_B2_M1003_g N_VPWR_c_316_n 0.00829547f $X=2.37 $Y=2.145 $X2=0 $Y2=0
cc_182 N_B2_M1003_g N_VPWR_c_313_n 0.00321451f $X=2.37 $Y=2.145 $X2=0 $Y2=0
cc_183 N_B2_c_239_n N_Y_c_346_n 0.00348516f $X=2.28 $Y=0.765 $X2=0 $Y2=0
cc_184 B2 N_Y_c_346_n 0.0477136f $X=2.555 $Y=0.84 $X2=0 $Y2=0
cc_185 N_B2_c_243_n N_Y_c_346_n 0.00396771f $X=2.28 $Y=0.93 $X2=0 $Y2=0
cc_186 N_B2_M1003_g N_Y_c_347_n 0.00314573f $X=2.37 $Y=2.145 $X2=0 $Y2=0
cc_187 B2 N_Y_c_347_n 0.00233005f $X=2.555 $Y=0.84 $X2=0 $Y2=0
cc_188 N_B2_c_239_n N_Y_c_359_n 0.00487762f $X=2.28 $Y=0.765 $X2=0 $Y2=0
cc_189 B2 N_Y_c_359_n 9.89683e-19 $X=2.555 $Y=0.84 $X2=0 $Y2=0
cc_190 N_B2_c_243_n N_Y_c_359_n 0.00188037f $X=2.28 $Y=0.93 $X2=0 $Y2=0
cc_191 N_B2_M1003_g Y 9.06541e-19 $X=2.37 $Y=2.145 $X2=0 $Y2=0
cc_192 N_B2_M1003_g N_A_403_387#_c_389_n 2.03427e-19 $X=2.37 $Y=2.145 $X2=0
+ $Y2=0
cc_193 N_B2_M1003_g N_A_403_387#_c_385_n 0.0144668f $X=2.37 $Y=2.145 $X2=0 $Y2=0
cc_194 N_B2_c_241_n N_A_403_387#_c_385_n 3.32529e-19 $X=2.28 $Y=1.435 $X2=0
+ $Y2=0
cc_195 B2 N_A_403_387#_c_385_n 0.0247246f $X=2.555 $Y=0.84 $X2=0 $Y2=0
cc_196 N_B2_c_241_n N_A_403_387#_c_386_n 0.00348027f $X=2.28 $Y=1.435 $X2=0
+ $Y2=0
cc_197 B2 N_A_403_387#_c_386_n 0.00237654f $X=2.555 $Y=0.84 $X2=0 $Y2=0
cc_198 N_B2_c_239_n N_VGND_c_405_n 0.0019812f $X=2.28 $Y=0.765 $X2=0 $Y2=0
cc_199 N_B2_c_239_n N_VGND_c_409_n 0.00551436f $X=2.28 $Y=0.765 $X2=0 $Y2=0
cc_200 N_B2_c_243_n N_VGND_c_409_n 7.94643e-19 $X=2.28 $Y=0.93 $X2=0 $Y2=0
cc_201 N_B2_c_239_n N_VGND_c_411_n 0.00635977f $X=2.28 $Y=0.765 $X2=0 $Y2=0
cc_202 B2 N_VGND_c_411_n 0.0197031f $X=2.555 $Y=0.84 $X2=0 $Y2=0
cc_203 N_B1_M1009_g N_VPWR_c_316_n 0.0143932f $X=2.8 $Y=2.145 $X2=0 $Y2=0
cc_204 N_B1_M1009_g N_VPWR_c_313_n 0.00321451f $X=2.8 $Y=2.145 $X2=0 $Y2=0
cc_205 N_B1_c_283_n N_Y_c_359_n 8.04745e-19 $X=2.905 $Y=0.765 $X2=0 $Y2=0
cc_206 N_B1_M1009_g N_A_403_387#_c_385_n 0.0196354f $X=2.8 $Y=2.145 $X2=0 $Y2=0
cc_207 N_B1_c_285_n N_A_403_387#_c_385_n 0.0025444f $X=2.94 $Y=1.435 $X2=0 $Y2=0
cc_208 B1 N_A_403_387#_c_385_n 0.0114252f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_209 N_B1_M1009_g N_A_403_387#_c_387_n 3.52891e-19 $X=2.8 $Y=2.145 $X2=0 $Y2=0
cc_210 B1 N_VGND_c_404_n 0.00138566f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_211 N_B1_c_283_n N_VGND_c_405_n 0.0116066f $X=2.905 $Y=0.765 $X2=0 $Y2=0
cc_212 N_B1_c_284_n N_VGND_c_405_n 0.00451659f $X=2.905 $Y=0.915 $X2=0 $Y2=0
cc_213 B1 N_VGND_c_405_n 0.0108758f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_214 N_B1_c_283_n N_VGND_c_409_n 0.00486043f $X=2.905 $Y=0.765 $X2=0 $Y2=0
cc_215 N_B1_c_283_n N_VGND_c_411_n 0.00635011f $X=2.905 $Y=0.765 $X2=0 $Y2=0
cc_216 B1 N_VGND_c_411_n 0.00352163f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_217 N_VPWR_c_316_n N_A_403_387#_c_385_n 0.0207154f $X=2.585 $Y=2.21 $X2=0
+ $Y2=0
cc_218 Y N_A_403_387#_c_389_n 5.52253e-19 $X=1.595 $Y=1.95 $X2=0 $Y2=0
cc_219 Y N_A_403_387#_c_386_n 0.0119514f $X=1.595 $Y=1.95 $X2=0 $Y2=0
cc_220 N_Y_c_359_n N_VGND_c_403_n 0.0121894f $X=2.045 $Y=0.48 $X2=0 $Y2=0
cc_221 N_Y_c_359_n N_VGND_c_405_n 0.00304905f $X=2.045 $Y=0.48 $X2=0 $Y2=0
cc_222 N_Y_c_359_n N_VGND_c_409_n 0.0113299f $X=2.045 $Y=0.48 $X2=0 $Y2=0
cc_223 N_Y_M1001_d N_VGND_c_411_n 0.00239483f $X=1.905 $Y=0.235 $X2=0 $Y2=0
cc_224 N_Y_c_359_n N_VGND_c_411_n 0.0123334f $X=2.045 $Y=0.48 $X2=0 $Y2=0
cc_225 N_VGND_c_411_n A_467_47# 0.00433137f $X=3.12 $Y=0 $X2=-0.19 $Y2=-0.245
