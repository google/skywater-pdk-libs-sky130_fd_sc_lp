* File: sky130_fd_sc_lp__and3_m.pxi.spice
* Created: Wed Sep  2 09:31:59 2020
* 
x_PM_SKY130_FD_SC_LP__AND3_M%A N_A_M1004_g N_A_M1006_g A A N_A_c_57_n
+ PM_SKY130_FD_SC_LP__AND3_M%A
x_PM_SKY130_FD_SC_LP__AND3_M%B N_B_M1002_g N_B_M1000_g N_B_c_79_n N_B_c_80_n
+ N_B_c_81_n B B B N_B_c_83_n PM_SKY130_FD_SC_LP__AND3_M%B
x_PM_SKY130_FD_SC_LP__AND3_M%C N_C_M1005_g N_C_M1003_g N_C_c_120_n N_C_c_125_n C
+ C C N_C_c_122_n PM_SKY130_FD_SC_LP__AND3_M%C
x_PM_SKY130_FD_SC_LP__AND3_M%A_51_47# N_A_51_47#_M1004_s N_A_51_47#_M1006_s
+ N_A_51_47#_M1000_d N_A_51_47#_c_170_n N_A_51_47#_M1001_g N_A_51_47#_c_165_n
+ N_A_51_47#_M1007_g N_A_51_47#_c_166_n N_A_51_47#_c_173_n N_A_51_47#_c_167_n
+ N_A_51_47#_c_168_n N_A_51_47#_c_169_n N_A_51_47#_c_175_n N_A_51_47#_c_176_n
+ N_A_51_47#_c_177_n N_A_51_47#_c_178_n N_A_51_47#_c_179_n N_A_51_47#_c_180_n
+ PM_SKY130_FD_SC_LP__AND3_M%A_51_47#
x_PM_SKY130_FD_SC_LP__AND3_M%VPWR N_VPWR_M1006_d N_VPWR_M1005_d N_VPWR_c_254_n
+ N_VPWR_c_255_n N_VPWR_c_256_n N_VPWR_c_257_n N_VPWR_c_258_n N_VPWR_c_259_n
+ VPWR N_VPWR_c_260_n N_VPWR_c_253_n N_VPWR_c_262_n
+ PM_SKY130_FD_SC_LP__AND3_M%VPWR
x_PM_SKY130_FD_SC_LP__AND3_M%X N_X_M1007_d N_X_M1001_d X X X X X X X
+ PM_SKY130_FD_SC_LP__AND3_M%X
x_PM_SKY130_FD_SC_LP__AND3_M%VGND N_VGND_M1003_d N_VGND_c_316_n VGND
+ N_VGND_c_317_n N_VGND_c_318_n N_VGND_c_319_n N_VGND_c_320_n
+ PM_SKY130_FD_SC_LP__AND3_M%VGND
cc_1 VNB N_A_M1004_g 0.0261778f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=0.445
cc_2 VNB N_A_M1006_g 0.0109967f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=2.165
cc_3 VNB A 0.0327846f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_4 VNB N_A_c_57_n 0.0800314f $X=-0.19 $Y=-0.245 $X2=0.345 $Y2=1.005
cc_5 VNB N_B_M1000_g 0.0121256f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=2.165
cc_6 VNB N_B_c_79_n 0.0162506f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_7 VNB N_B_c_80_n 0.0208673f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_8 VNB N_B_c_81_n 0.0152974f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB B 0.00780412f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_B_c_83_n 0.0153242f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_C_M1003_g 0.0368799f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=2.165
cc_12 VNB N_C_c_120_n 0.00924947f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB C 0.00808111f $X=-0.19 $Y=-0.245 $X2=0.425 $Y2=1.005
cc_14 VNB N_C_c_122_n 0.0313688f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_51_47#_c_165_n 0.0202769f $X=-0.19 $Y=-0.245 $X2=0.425 $Y2=0.84
cc_16 VNB N_A_51_47#_c_166_n 0.048317f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_51_47#_c_167_n 0.0235426f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_51_47#_c_168_n 0.00191853f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_51_47#_c_169_n 0.00671778f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_VPWR_c_253_n 0.103974f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB X 0.0360215f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=2.165
cc_22 VNB N_VGND_c_316_n 0.00494119f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=2.165
cc_23 VNB N_VGND_c_317_n 0.0471271f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_24 VNB N_VGND_c_318_n 0.0187831f $X=-0.19 $Y=-0.245 $X2=0.425 $Y2=1.51
cc_25 VNB N_VGND_c_319_n 0.15343f $X=-0.19 $Y=-0.245 $X2=0.292 $Y2=0.925
cc_26 VNB N_VGND_c_320_n 0.00401177f $X=-0.19 $Y=-0.245 $X2=0.292 $Y2=1.005
cc_27 VPB N_A_M1006_g 0.0358236f $X=-0.19 $Y=1.655 $X2=0.595 $Y2=2.165
cc_28 VPB N_B_M1000_g 0.0275526f $X=-0.19 $Y=1.655 $X2=0.595 $Y2=2.165
cc_29 VPB N_C_M1005_g 0.0166659f $X=-0.19 $Y=1.655 $X2=0.595 $Y2=0.445
cc_30 VPB N_C_c_120_n 0.00103988f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_31 VPB N_C_c_125_n 0.0126304f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_32 VPB C 0.00298794f $X=-0.19 $Y=1.655 $X2=0.425 $Y2=1.005
cc_33 VPB N_A_51_47#_c_170_n 0.0355226f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_34 VPB N_A_51_47#_M1001_g 0.028381f $X=-0.19 $Y=1.655 $X2=0.345 $Y2=1.005
cc_35 VPB N_A_51_47#_c_166_n 0.00265628f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_36 VPB N_A_51_47#_c_173_n 0.0278128f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_37 VPB N_A_51_47#_c_169_n 5.66269e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_38 VPB N_A_51_47#_c_175_n 0.00803715f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_39 VPB N_A_51_47#_c_176_n 0.0271166f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_40 VPB N_A_51_47#_c_177_n 0.00701902f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_41 VPB N_A_51_47#_c_178_n 0.00264527f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_42 VPB N_A_51_47#_c_179_n 0.00764809f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_43 VPB N_A_51_47#_c_180_n 0.0426505f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_44 VPB N_VPWR_c_254_n 0.0375579f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_45 VPB N_VPWR_c_255_n 0.020512f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_46 VPB N_VPWR_c_256_n 0.0168972f $X=-0.19 $Y=1.655 $X2=0.345 $Y2=1.005
cc_47 VPB N_VPWR_c_257_n 0.0252142f $X=-0.19 $Y=1.655 $X2=0.345 $Y2=1.005
cc_48 VPB N_VPWR_c_258_n 0.00362871f $X=-0.19 $Y=1.655 $X2=0.425 $Y2=0.84
cc_49 VPB N_VPWR_c_259_n 0.00112291f $X=-0.19 $Y=1.655 $X2=0.292 $Y2=0.925
cc_50 VPB N_VPWR_c_260_n 0.0192288f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_51 VPB N_VPWR_c_253_n 0.0867763f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_52 VPB N_VPWR_c_262_n 0.00324402f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_53 VPB X 0.0545807f $X=-0.19 $Y=1.655 $X2=0.595 $Y2=2.165
cc_54 N_A_c_57_n N_B_M1000_g 0.0296884f $X=0.345 $Y=1.005 $X2=0 $Y2=0
cc_55 N_A_M1004_g N_B_c_79_n 0.0410696f $X=0.595 $Y=0.445 $X2=0 $Y2=0
cc_56 N_A_c_57_n N_B_c_80_n 0.0410696f $X=0.345 $Y=1.005 $X2=0 $Y2=0
cc_57 N_A_M1004_g B 8.64076e-19 $X=0.595 $Y=0.445 $X2=0 $Y2=0
cc_58 N_A_M1004_g N_A_51_47#_c_168_n 0.0121006f $X=0.595 $Y=0.445 $X2=0 $Y2=0
cc_59 A N_A_51_47#_c_168_n 0.0120027f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_60 N_A_c_57_n N_A_51_47#_c_168_n 0.00507518f $X=0.345 $Y=1.005 $X2=0 $Y2=0
cc_61 N_A_M1004_g N_A_51_47#_c_169_n 0.00851049f $X=0.595 $Y=0.445 $X2=0 $Y2=0
cc_62 N_A_M1006_g N_A_51_47#_c_169_n 0.0100625f $X=0.595 $Y=2.165 $X2=0 $Y2=0
cc_63 A N_A_51_47#_c_169_n 0.0450414f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_64 N_A_c_57_n N_A_51_47#_c_169_n 0.0163785f $X=0.345 $Y=1.005 $X2=0 $Y2=0
cc_65 N_A_M1006_g N_A_51_47#_c_176_n 0.024908f $X=0.595 $Y=2.165 $X2=0 $Y2=0
cc_66 A N_A_51_47#_c_176_n 0.0161191f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_67 N_A_c_57_n N_A_51_47#_c_176_n 0.00560486f $X=0.345 $Y=1.005 $X2=0 $Y2=0
cc_68 N_A_M1006_g N_VPWR_c_254_n 0.00314874f $X=0.595 $Y=2.165 $X2=0 $Y2=0
cc_69 N_A_M1006_g N_VPWR_c_253_n 0.00387136f $X=0.595 $Y=2.165 $X2=0 $Y2=0
cc_70 N_A_M1004_g N_VGND_c_317_n 0.00372993f $X=0.595 $Y=0.445 $X2=0 $Y2=0
cc_71 N_A_M1004_g N_VGND_c_319_n 0.00639832f $X=0.595 $Y=0.445 $X2=0 $Y2=0
cc_72 A N_VGND_c_319_n 0.00455527f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_73 N_B_c_79_n N_C_M1003_g 0.0190955f $X=1.045 $Y=0.765 $X2=0 $Y2=0
cc_74 B N_C_M1003_g 0.0119503f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_75 N_B_c_83_n N_C_M1003_g 0.0201419f $X=1.045 $Y=0.93 $X2=0 $Y2=0
cc_76 N_B_M1000_g N_C_c_125_n 0.0183424f $X=1.025 $Y=2.165 $X2=0 $Y2=0
cc_77 N_B_M1000_g C 0.00147107f $X=1.025 $Y=2.165 $X2=0 $Y2=0
cc_78 B C 0.0388108f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_79 N_B_c_83_n C 5.77029e-19 $X=1.045 $Y=0.93 $X2=0 $Y2=0
cc_80 N_B_M1000_g N_C_c_122_n 0.0086346f $X=1.025 $Y=2.165 $X2=0 $Y2=0
cc_81 N_B_c_80_n N_C_c_122_n 0.0201419f $X=1.045 $Y=1.27 $X2=0 $Y2=0
cc_82 N_B_c_79_n N_A_51_47#_c_168_n 0.00500134f $X=1.045 $Y=0.765 $X2=0 $Y2=0
cc_83 B N_A_51_47#_c_168_n 0.0146519f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_84 N_B_M1000_g N_A_51_47#_c_169_n 0.00576954f $X=1.025 $Y=2.165 $X2=0 $Y2=0
cc_85 N_B_c_79_n N_A_51_47#_c_169_n 0.00473923f $X=1.045 $Y=0.765 $X2=0 $Y2=0
cc_86 B N_A_51_47#_c_169_n 0.0555762f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_87 N_B_M1000_g N_A_51_47#_c_175_n 0.015149f $X=1.025 $Y=2.165 $X2=0 $Y2=0
cc_88 N_B_c_81_n N_A_51_47#_c_175_n 0.00279988f $X=1.045 $Y=1.435 $X2=0 $Y2=0
cc_89 B N_A_51_47#_c_175_n 0.0089875f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_90 N_B_M1000_g N_A_51_47#_c_176_n 5.20386e-19 $X=1.025 $Y=2.165 $X2=0 $Y2=0
cc_91 N_B_M1000_g N_A_51_47#_c_177_n 8.9241e-19 $X=1.025 $Y=2.165 $X2=0 $Y2=0
cc_92 N_B_c_81_n N_A_51_47#_c_177_n 5.53883e-19 $X=1.045 $Y=1.435 $X2=0 $Y2=0
cc_93 B N_A_51_47#_c_177_n 0.00948297f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_94 N_B_M1000_g N_A_51_47#_c_179_n 0.00141726f $X=1.025 $Y=2.165 $X2=0 $Y2=0
cc_95 N_B_M1000_g N_VPWR_c_254_n 0.00105495f $X=1.025 $Y=2.165 $X2=0 $Y2=0
cc_96 N_B_M1000_g N_VPWR_c_253_n 0.00387136f $X=1.025 $Y=2.165 $X2=0 $Y2=0
cc_97 B A_206_47# 0.00551255f $X=1.115 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_98 N_B_c_79_n N_VGND_c_317_n 0.00499463f $X=1.045 $Y=0.765 $X2=0 $Y2=0
cc_99 B N_VGND_c_317_n 0.00847263f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_100 N_B_c_83_n N_VGND_c_317_n 4.84097e-19 $X=1.045 $Y=0.93 $X2=0 $Y2=0
cc_101 N_B_c_79_n N_VGND_c_319_n 0.00865283f $X=1.045 $Y=0.765 $X2=0 $Y2=0
cc_102 B N_VGND_c_319_n 0.0106876f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_103 N_C_M1003_g N_A_51_47#_c_165_n 0.0209764f $X=1.495 $Y=0.445 $X2=0 $Y2=0
cc_104 N_C_M1003_g N_A_51_47#_c_166_n 0.00550988f $X=1.495 $Y=0.445 $X2=0 $Y2=0
cc_105 N_C_c_120_n N_A_51_47#_c_166_n 0.00480605f $X=1.475 $Y=1.675 $X2=0 $Y2=0
cc_106 C N_A_51_47#_c_166_n 0.00502703f $X=1.595 $Y=0.84 $X2=0 $Y2=0
cc_107 N_C_c_122_n N_A_51_47#_c_166_n 0.0166105f $X=1.585 $Y=1.32 $X2=0 $Y2=0
cc_108 N_C_M1005_g N_A_51_47#_c_173_n 0.0139977f $X=1.455 $Y=2.165 $X2=0 $Y2=0
cc_109 N_C_c_125_n N_A_51_47#_c_173_n 0.00693566f $X=1.475 $Y=1.825 $X2=0 $Y2=0
cc_110 C N_A_51_47#_c_173_n 4.73927e-19 $X=1.595 $Y=0.84 $X2=0 $Y2=0
cc_111 C N_A_51_47#_c_167_n 6.30053e-19 $X=1.595 $Y=0.84 $X2=0 $Y2=0
cc_112 N_C_M1005_g N_A_51_47#_c_177_n 2.67283e-19 $X=1.455 $Y=2.165 $X2=0 $Y2=0
cc_113 N_C_c_125_n N_A_51_47#_c_177_n 0.00564503f $X=1.475 $Y=1.825 $X2=0 $Y2=0
cc_114 C N_A_51_47#_c_177_n 0.00262304f $X=1.595 $Y=0.84 $X2=0 $Y2=0
cc_115 N_C_M1005_g N_A_51_47#_c_178_n 5.45931e-19 $X=1.455 $Y=2.165 $X2=0 $Y2=0
cc_116 N_C_M1005_g N_A_51_47#_c_179_n 0.00154996f $X=1.455 $Y=2.165 $X2=0 $Y2=0
cc_117 N_C_M1005_g N_A_51_47#_c_180_n 0.00954305f $X=1.455 $Y=2.165 $X2=0 $Y2=0
cc_118 N_C_M1005_g N_VPWR_c_256_n 8.55012e-19 $X=1.455 $Y=2.165 $X2=0 $Y2=0
cc_119 C N_VPWR_c_259_n 0.0105759f $X=1.595 $Y=0.84 $X2=0 $Y2=0
cc_120 N_C_c_122_n N_VPWR_c_259_n 7.52351e-19 $X=1.585 $Y=1.32 $X2=0 $Y2=0
cc_121 N_C_M1003_g X 0.00167598f $X=1.495 $Y=0.445 $X2=0 $Y2=0
cc_122 N_C_c_120_n X 2.43546e-19 $X=1.475 $Y=1.675 $X2=0 $Y2=0
cc_123 N_C_c_125_n X 3.40634e-19 $X=1.475 $Y=1.825 $X2=0 $Y2=0
cc_124 C X 0.0552958f $X=1.595 $Y=0.84 $X2=0 $Y2=0
cc_125 N_C_c_122_n X 4.09003e-19 $X=1.585 $Y=1.32 $X2=0 $Y2=0
cc_126 N_C_M1003_g N_VGND_c_316_n 0.00288714f $X=1.495 $Y=0.445 $X2=0 $Y2=0
cc_127 C N_VGND_c_316_n 0.00821138f $X=1.595 $Y=0.84 $X2=0 $Y2=0
cc_128 N_C_c_122_n N_VGND_c_316_n 5.47722e-19 $X=1.585 $Y=1.32 $X2=0 $Y2=0
cc_129 N_C_M1003_g N_VGND_c_317_n 0.00585385f $X=1.495 $Y=0.445 $X2=0 $Y2=0
cc_130 N_C_M1003_g N_VGND_c_319_n 0.0089947f $X=1.495 $Y=0.445 $X2=0 $Y2=0
cc_131 C N_VGND_c_319_n 0.00430742f $X=1.595 $Y=0.84 $X2=0 $Y2=0
cc_132 N_A_51_47#_c_175_n N_VPWR_c_254_n 0.00968807f $X=1.135 $Y=1.8 $X2=0 $Y2=0
cc_133 N_A_51_47#_c_176_n N_VPWR_c_254_n 0.00467243f $X=0.78 $Y=1.8 $X2=0 $Y2=0
cc_134 N_A_51_47#_c_178_n N_VPWR_c_254_n 0.0105383f $X=1.24 $Y=2.825 $X2=0 $Y2=0
cc_135 N_A_51_47#_c_179_n N_VPWR_c_254_n 0.0286013f $X=1.24 $Y=2.1 $X2=0 $Y2=0
cc_136 N_A_51_47#_c_180_n N_VPWR_c_254_n 0.00612344f $X=1.3 $Y=2.82 $X2=0 $Y2=0
cc_137 N_A_51_47#_c_170_n N_VPWR_c_255_n 0.00427618f $X=1.81 $Y=2.82 $X2=0 $Y2=0
cc_138 N_A_51_47#_c_178_n N_VPWR_c_255_n 0.013307f $X=1.24 $Y=2.825 $X2=0 $Y2=0
cc_139 N_A_51_47#_c_180_n N_VPWR_c_255_n 0.00748434f $X=1.3 $Y=2.82 $X2=0 $Y2=0
cc_140 N_A_51_47#_c_170_n N_VPWR_c_256_n 0.014786f $X=1.81 $Y=2.82 $X2=0 $Y2=0
cc_141 N_A_51_47#_M1001_g N_VPWR_c_256_n 0.00841415f $X=1.885 $Y=2.165 $X2=0
+ $Y2=0
cc_142 N_A_51_47#_c_178_n N_VPWR_c_256_n 0.0118902f $X=1.24 $Y=2.825 $X2=0 $Y2=0
cc_143 N_A_51_47#_c_179_n N_VPWR_c_256_n 0.0215252f $X=1.24 $Y=2.1 $X2=0 $Y2=0
cc_144 N_A_51_47#_c_180_n N_VPWR_c_256_n 0.00369946f $X=1.3 $Y=2.82 $X2=0 $Y2=0
cc_145 N_A_51_47#_c_170_n N_VPWR_c_259_n 0.00242431f $X=1.81 $Y=2.82 $X2=0 $Y2=0
cc_146 N_A_51_47#_M1001_g N_VPWR_c_259_n 0.00332502f $X=1.885 $Y=2.165 $X2=0
+ $Y2=0
cc_147 N_A_51_47#_c_179_n N_VPWR_c_259_n 0.00124848f $X=1.24 $Y=2.1 $X2=0 $Y2=0
cc_148 N_A_51_47#_c_170_n N_VPWR_c_260_n 0.00432443f $X=1.81 $Y=2.82 $X2=0 $Y2=0
cc_149 N_A_51_47#_c_170_n N_VPWR_c_253_n 0.009398f $X=1.81 $Y=2.82 $X2=0 $Y2=0
cc_150 N_A_51_47#_c_178_n N_VPWR_c_253_n 0.0115437f $X=1.24 $Y=2.825 $X2=0 $Y2=0
cc_151 N_A_51_47#_c_180_n N_VPWR_c_253_n 0.0105534f $X=1.3 $Y=2.82 $X2=0 $Y2=0
cc_152 N_A_51_47#_M1001_g X 0.0179259f $X=1.885 $Y=2.165 $X2=0 $Y2=0
cc_153 N_A_51_47#_c_165_n X 0.00743422f $X=1.925 $Y=0.765 $X2=0 $Y2=0
cc_154 N_A_51_47#_c_166_n X 0.0278837f $X=2.065 $Y=1.695 $X2=0 $Y2=0
cc_155 N_A_51_47#_c_173_n X 0.0102393f $X=2.065 $Y=1.77 $X2=0 $Y2=0
cc_156 N_A_51_47#_c_167_n X 0.0094603f $X=2.065 $Y=0.84 $X2=0 $Y2=0
cc_157 N_A_51_47#_c_177_n X 5.76623e-19 $X=1.24 $Y=2.04 $X2=0 $Y2=0
cc_158 N_A_51_47#_c_168_n A_134_47# 0.0039738f $X=0.61 $Y=0.495 $X2=-0.19
+ $Y2=-0.245
cc_159 N_A_51_47#_c_165_n N_VGND_c_316_n 0.00288714f $X=1.925 $Y=0.765 $X2=0
+ $Y2=0
cc_160 N_A_51_47#_c_168_n N_VGND_c_317_n 0.0203008f $X=0.61 $Y=0.495 $X2=0 $Y2=0
cc_161 N_A_51_47#_c_165_n N_VGND_c_318_n 0.00579795f $X=1.925 $Y=0.765 $X2=0
+ $Y2=0
cc_162 N_A_51_47#_c_167_n N_VGND_c_318_n 3.33196e-19 $X=2.065 $Y=0.84 $X2=0
+ $Y2=0
cc_163 N_A_51_47#_M1004_s N_VGND_c_319_n 0.00234684f $X=0.255 $Y=0.235 $X2=0
+ $Y2=0
cc_164 N_A_51_47#_c_165_n N_VGND_c_319_n 0.0115436f $X=1.925 $Y=0.765 $X2=0
+ $Y2=0
cc_165 N_A_51_47#_c_168_n N_VGND_c_319_n 0.0178558f $X=0.61 $Y=0.495 $X2=0 $Y2=0
cc_166 N_VPWR_c_259_n X 0.0448667f $X=1.67 $Y=2.23 $X2=0 $Y2=0
cc_167 N_VPWR_c_260_n X 0.00743562f $X=2.16 $Y=3.33 $X2=0 $Y2=0
cc_168 N_VPWR_c_253_n X 0.00847205f $X=2.16 $Y=3.33 $X2=0 $Y2=0
cc_169 X N_VGND_c_318_n 0.0097709f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_170 N_X_M1007_d N_VGND_c_319_n 0.00296381f $X=2 $Y=0.235 $X2=0 $Y2=0
cc_171 X N_VGND_c_319_n 0.00915554f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_172 A_134_47# N_VGND_c_319_n 0.00519157f $X=0.67 $Y=0.235 $X2=1.925 $Y2=0.445
cc_173 A_206_47# N_VGND_c_319_n 0.00823499f $X=1.03 $Y=0.235 $X2=1.045 $Y2=0.93
