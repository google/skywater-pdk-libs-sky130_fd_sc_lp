* File: sky130_fd_sc_lp__a311o_4.spice
* Created: Wed Sep  2 09:25:14 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__a311o_4.pex.spice"
.subckt sky130_fd_sc_lp__a311o_4  VNB VPB C1 B1 A3 A2 A1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A1	A1
* A2	A2
* A3	A3
* B1	B1
* C1	C1
* VPB	VPB
* VNB	VNB
MM1002 N_A_111_47#_M1002_d N_C1_M1002_g N_VGND_M1002_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75004.5 A=0.126 P=1.98 MULT=1
MM1010 N_A_111_47#_M1002_d N_C1_M1010_g N_VGND_M1010_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1344 PD=1.12 PS=1.16 NRD=0 NRS=2.136 M=1 R=5.6 SA=75000.6
+ SB=75004.1 A=0.126 P=1.98 MULT=1
MM1000 N_A_111_47#_M1000_d N_B1_M1000_g N_VGND_M1010_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1344 PD=1.12 PS=1.16 NRD=0 NRS=3.564 M=1 R=5.6 SA=75001.1
+ SB=75003.6 A=0.126 P=1.98 MULT=1
MM1020 N_A_111_47#_M1000_d N_B1_M1020_g N_VGND_M1020_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1218 PD=1.12 PS=1.13 NRD=0 NRS=0 M=1 R=5.6 SA=75001.5
+ SB=75003.2 A=0.126 P=1.98 MULT=1
MM1011 N_X_M1011_d N_A_111_47#_M1011_g N_VGND_M1020_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1218 PD=1.12 PS=1.13 NRD=0 NRS=1.428 M=1 R=5.6 SA=75002
+ SB=75002.8 A=0.126 P=1.98 MULT=1
MM1012 N_X_M1011_d N_A_111_47#_M1012_g N_VGND_M1012_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002.4
+ SB=75002.3 A=0.126 P=1.98 MULT=1
MM1014 N_X_M1014_d N_A_111_47#_M1014_g N_VGND_M1012_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002.8
+ SB=75001.9 A=0.126 P=1.98 MULT=1
MM1021 N_X_M1014_d N_A_111_47#_M1021_g N_VGND_M1021_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2604 PD=1.12 PS=1.46 NRD=0 NRS=0 M=1 R=5.6 SA=75003.2
+ SB=75001.5 A=0.126 P=1.98 MULT=1
MM1005 N_A_877_47#_M1005_d N_A3_M1005_g N_VGND_M1021_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2604 PD=1.12 PS=1.46 NRD=0 NRS=0 M=1 R=5.6 SA=75004 SB=75000.7
+ A=0.126 P=1.98 MULT=1
MM1016 N_A_877_47#_M1005_d N_A3_M1016_g N_VGND_M1016_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2814 PD=1.12 PS=2.35 NRD=0 NRS=0 M=1 R=5.6 SA=75004.4
+ SB=75000.3 A=0.126 P=1.98 MULT=1
MM1006 N_A_1098_69#_M1006_d N_A2_M1006_g N_A_877_47#_M1006_s VNB NSHORT L=0.15
+ W=0.84 AD=0.2226 AS=0.1491 PD=2.21 PS=1.195 NRD=0 NRS=4.992 M=1 R=5.6
+ SA=75000.2 SB=75001.6 A=0.126 P=1.98 MULT=1
MM1018 N_A_1098_69#_M1018_d N_A2_M1018_g N_A_877_47#_M1006_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1491 PD=1.12 PS=1.195 NRD=0 NRS=5.712 M=1 R=5.6
+ SA=75000.7 SB=75001.1 A=0.126 P=1.98 MULT=1
MM1004 N_A_1098_69#_M1018_d N_A1_M1004_g N_A_111_47#_M1004_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.1
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1022 N_A_1098_69#_M1022_d N_A1_M1022_g N_A_111_47#_M1004_s VNB NSHORT L=0.15
+ W=0.84 AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.6
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1013 N_A_28_367#_M1013_d N_C1_M1013_g N_A_111_47#_M1013_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75001.5 A=0.189 P=2.82 MULT=1
MM1026 N_A_28_367#_M1026_d N_C1_M1026_g N_A_111_47#_M1013_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1024 N_A_28_367#_M1026_d N_B1_M1024_g N_A_283_367#_M1024_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.2016 PD=1.54 PS=1.58 NRD=0 NRS=3.1126 M=1 R=8.4
+ SA=75001.1 SB=75000.7 A=0.189 P=2.82 MULT=1
MM1027 N_A_28_367#_M1027_d N_B1_M1027_g N_A_283_367#_M1024_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.2016 PD=3.05 PS=1.58 NRD=0 NRS=3.1126 M=1 R=8.4
+ SA=75001.5 SB=75000.2 A=0.189 P=2.82 MULT=1
MM1001 N_VPWR_M1001_d N_A_111_47#_M1001_g N_X_M1001_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.4686 AS=0.1764 PD=3.36 PS=1.54 NRD=15.6221 NRS=0 M=1 R=8.4 SA=75000.3
+ SB=75004.3 A=0.189 P=2.82 MULT=1
MM1003 N_VPWR_M1003_d N_A_111_47#_M1003_g N_X_M1001_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.262 AS=0.1764 PD=1.74 PS=1.54 NRD=10.1455 NRS=0 M=1 R=8.4 SA=75000.7
+ SB=75003.9 A=0.189 P=2.82 MULT=1
MM1009 N_VPWR_M1003_d N_A_111_47#_M1009_g N_X_M1009_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.262 AS=0.3036 PD=1.74 PS=1.79 NRD=10.1455 NRS=14.8341 M=1 R=8.4
+ SA=75001.3 SB=75003.3 A=0.189 P=2.82 MULT=1
MM1015 N_VPWR_M1015_d N_A_111_47#_M1015_g N_X_M1009_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.3036 PD=1.54 PS=1.79 NRD=0 NRS=15.6221 M=1 R=8.4 SA=75001.8
+ SB=75002.8 A=0.189 P=2.82 MULT=1
MM1007 N_VPWR_M1015_d N_A3_M1007_g N_A_283_367#_M1007_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.2
+ SB=75002.4 A=0.189 P=2.82 MULT=1
MM1023 N_VPWR_M1023_d N_A3_M1023_g N_A_283_367#_M1007_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.7
+ SB=75002 A=0.189 P=2.82 MULT=1
MM1017 N_VPWR_M1023_d N_A2_M1017_g N_A_283_367#_M1017_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75003.1
+ SB=75001.6 A=0.189 P=2.82 MULT=1
MM1025 N_VPWR_M1025_d N_A2_M1025_g N_A_283_367#_M1017_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.22365 AS=0.1764 PD=1.615 PS=1.54 NRD=5.4569 NRS=0 M=1 R=8.4
+ SA=75003.5 SB=75001.1 A=0.189 P=2.82 MULT=1
MM1008 N_VPWR_M1025_d N_A1_M1008_g N_A_283_367#_M1008_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.22365 AS=0.1764 PD=1.615 PS=1.54 NRD=6.2449 NRS=0 M=1 R=8.4
+ SA=75004 SB=75000.6 A=0.189 P=2.82 MULT=1
MM1019 N_VPWR_M1019_d N_A1_M1019_g N_A_283_367#_M1008_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75004.5
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX28_noxref VNB VPB NWDIODE A=15.1645 P=19.97
*
.include "sky130_fd_sc_lp__a311o_4.pxi.spice"
*
.ends
*
*
