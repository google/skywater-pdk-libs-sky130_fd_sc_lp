* File: sky130_fd_sc_lp__o41ai_m.pex.spice
* Created: Fri Aug 28 11:20:53 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O41AI_M%B1 2 5 9 10 11 12 13 18 20
r39 18 20 45.5639 $w=3.95e-07 $l=1.65e-07 $layer=POLY_cond $X=0.677 $Y=0.93
+ $X2=0.677 $Y2=0.765
r40 12 13 22.798 $w=1.78e-07 $l=3.7e-07 $layer=LI1_cond $X=0.715 $Y=0.925
+ $X2=0.715 $Y2=1.295
r41 12 18 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.71
+ $Y=0.93 $X2=0.71 $Y2=0.93
r42 11 12 22.798 $w=1.78e-07 $l=3.7e-07 $layer=LI1_cond $X=0.715 $Y=0.555
+ $X2=0.715 $Y2=0.925
r43 9 20 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.8 $Y=0.445 $X2=0.8
+ $Y2=0.765
r44 5 10 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=0.555 $Y=2.065
+ $X2=0.555 $Y2=1.435
r45 2 10 50.0695 $w=3.95e-07 $l=1.97e-07 $layer=POLY_cond $X=0.677 $Y=1.238
+ $X2=0.677 $Y2=1.435
r46 1 18 4.50555 $w=3.95e-07 $l=3.2e-08 $layer=POLY_cond $X=0.677 $Y=0.962
+ $X2=0.677 $Y2=0.93
r47 1 2 38.8604 $w=3.95e-07 $l=2.76e-07 $layer=POLY_cond $X=0.677 $Y=0.962
+ $X2=0.677 $Y2=1.238
.ends

.subckt PM_SKY130_FD_SC_LP__O41AI_M%A4 3 7 11 12 13 14 15 20 21
r42 20 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.25
+ $Y=1.19 $X2=1.25 $Y2=1.19
r43 14 15 19.382 $w=2.18e-07 $l=3.7e-07 $layer=LI1_cond $X=1.225 $Y=1.665
+ $X2=1.225 $Y2=2.035
r44 13 14 19.382 $w=2.18e-07 $l=3.7e-07 $layer=LI1_cond $X=1.225 $Y=1.295
+ $X2=1.225 $Y2=1.665
r45 13 21 5.5003 $w=2.18e-07 $l=1.05e-07 $layer=LI1_cond $X=1.225 $Y=1.295
+ $X2=1.225 $Y2=1.19
r46 11 20 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.25 $Y=1.53
+ $X2=1.25 $Y2=1.19
r47 11 12 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.25 $Y=1.53
+ $X2=1.25 $Y2=1.695
r48 10 20 39.6269 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.25 $Y=1.025
+ $X2=1.25 $Y2=1.19
r49 7 10 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=1.285 $Y=0.445
+ $X2=1.285 $Y2=1.025
r50 3 12 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=1.16 $Y=2.065
+ $X2=1.16 $Y2=1.695
.ends

.subckt PM_SKY130_FD_SC_LP__O41AI_M%A3 3 7 11 12 13 14 15 20 21
c37 3 0 1.9275e-19 $X=1.7 $Y=2.065
r38 20 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.79
+ $Y=1.19 $X2=1.79 $Y2=1.19
r39 14 15 15.2287 $w=2.78e-07 $l=3.7e-07 $layer=LI1_cond $X=1.735 $Y=1.665
+ $X2=1.735 $Y2=2.035
r40 13 14 15.2287 $w=2.78e-07 $l=3.7e-07 $layer=LI1_cond $X=1.735 $Y=1.295
+ $X2=1.735 $Y2=1.665
r41 13 21 4.32166 $w=2.78e-07 $l=1.05e-07 $layer=LI1_cond $X=1.735 $Y=1.295
+ $X2=1.735 $Y2=1.19
r42 11 20 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.79 $Y=1.53
+ $X2=1.79 $Y2=1.19
r43 11 12 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.79 $Y=1.53
+ $X2=1.79 $Y2=1.695
r44 10 20 38.6168 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.79 $Y=1.025
+ $X2=1.79 $Y2=1.19
r45 7 10 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=1.81 $Y=0.445
+ $X2=1.81 $Y2=1.025
r46 3 12 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=1.7 $Y=2.065 $X2=1.7
+ $Y2=1.695
.ends

.subckt PM_SKY130_FD_SC_LP__O41AI_M%A2 3 6 9 11 13 15 17 30
r37 30 31 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.15 $Y=2.6
+ $X2=2.15 $Y2=2.6
r38 15 17 8.14351 $w=7.03e-07 $l=4.8e-07 $layer=LI1_cond $X=2.16 $Y=2.672
+ $X2=2.64 $Y2=2.672
r39 15 31 0.169657 $w=7.03e-07 $l=1e-08 $layer=LI1_cond $X=2.16 $Y=2.672
+ $X2=2.15 $Y2=2.672
r40 13 31 7.97386 $w=7.03e-07 $l=4.7e-07 $layer=LI1_cond $X=1.68 $Y=2.672
+ $X2=2.15 $Y2=2.672
r41 11 13 8.14351 $w=7.03e-07 $l=4.8e-07 $layer=LI1_cond $X=1.2 $Y=2.672
+ $X2=1.68 $Y2=2.672
r42 9 11 8.14351 $w=7.03e-07 $l=4.8e-07 $layer=LI1_cond $X=0.72 $Y=2.672 $X2=1.2
+ $Y2=2.672
r43 8 30 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.15 $Y=2.435
+ $X2=2.15 $Y2=2.6
r44 6 8 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=2.24 $Y=2.065 $X2=2.24
+ $Y2=2.435
r45 3 6 830.681 $w=1.5e-07 $l=1.62e-06 $layer=POLY_cond $X=2.24 $Y=0.445
+ $X2=2.24 $Y2=2.065
.ends

.subckt PM_SKY130_FD_SC_LP__O41AI_M%A1 3 7 10 11 12 14 16 25
c28 16 0 1.9275e-19 $X=3.12 $Y=1.665
r29 25 26 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.69
+ $Y=1.14 $X2=2.69 $Y2=1.14
r30 16 26 7.4002 $w=6.93e-07 $l=4.3e-07 $layer=LI1_cond $X=3.12 $Y=1.402
+ $X2=2.69 $Y2=1.402
r31 14 26 0.860488 $w=6.93e-07 $l=5e-08 $layer=LI1_cond $X=2.64 $Y=1.402
+ $X2=2.69 $Y2=1.402
r32 12 14 8.26068 $w=6.93e-07 $l=4.8e-07 $layer=LI1_cond $X=2.16 $Y=1.402
+ $X2=2.64 $Y2=1.402
r33 10 25 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.69 $Y=1.48
+ $X2=2.69 $Y2=1.14
r34 10 11 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.69 $Y=1.48
+ $X2=2.69 $Y2=1.645
r35 5 25 37.5318 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.69 $Y=0.975
+ $X2=2.69 $Y2=1.14
r36 5 7 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.69 $Y=0.975 $X2=2.69
+ $Y2=0.445
r37 3 11 215.362 $w=1.5e-07 $l=4.2e-07 $layer=POLY_cond $X=2.6 $Y=2.065 $X2=2.6
+ $Y2=1.645
.ends

.subckt PM_SKY130_FD_SC_LP__O41AI_M%VPWR 1 2 7 9 12 16 18 19 20 21 32
r26 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r27 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r28 29 32 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r29 28 29 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r30 26 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r31 25 28 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=0.72 $Y=3.33
+ $X2=2.64 $Y2=3.33
r32 25 26 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r33 23 34 3.5042 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=3.33
+ $X2=0.212 $Y2=3.33
r34 23 25 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.425 $Y=3.33
+ $X2=0.72 $Y2=3.33
r35 21 29 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r36 21 26 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.72 $Y2=3.33
r37 19 28 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=2.905 $Y=3.33
+ $X2=2.64 $Y2=3.33
r38 19 20 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.905 $Y=3.33
+ $X2=2.99 $Y2=3.33
r39 18 31 3.22941 $w=1.7e-07 $l=4.5e-08 $layer=LI1_cond $X=3.075 $Y=3.33
+ $X2=3.12 $Y2=3.33
r40 18 20 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.075 $Y=3.33
+ $X2=2.99 $Y2=3.33
r41 14 16 9.24242 $w=2.08e-07 $l=1.75e-07 $layer=LI1_cond $X=2.815 $Y=2.035
+ $X2=2.99 $Y2=2.035
r42 12 20 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.99 $Y=3.245
+ $X2=2.99 $Y2=3.33
r43 11 16 1.9771 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=2.99 $Y=2.14 $X2=2.99
+ $Y2=2.035
r44 11 12 72.0909 $w=1.68e-07 $l=1.105e-06 $layer=LI1_cond $X=2.99 $Y=2.14
+ $X2=2.99 $Y2=3.245
r45 7 34 3.33969 $w=1.9e-07 $l=1.54771e-07 $layer=LI1_cond $X=0.33 $Y=3.245
+ $X2=0.212 $Y2=3.33
r46 7 9 65.0861 $w=1.88e-07 $l=1.115e-06 $layer=LI1_cond $X=0.33 $Y=3.245
+ $X2=0.33 $Y2=2.13
r47 2 14 600 $w=1.7e-07 $l=2.4e-07 $layer=licon1_PDIFF $count=1 $X=2.675
+ $Y=1.855 $X2=2.815 $Y2=2.035
r48 1 9 600 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_PDIFF $count=1 $X=0.215
+ $Y=1.855 $X2=0.34 $Y2=2.13
.ends

.subckt PM_SKY130_FD_SC_LP__O41AI_M%Y 1 2 7 8 13 14 15 16 25 38
r27 16 25 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.24 $Y=1.7 $X2=0.24
+ $Y2=1.615
r28 16 25 1.17433 $w=1.68e-07 $l=1.8e-08 $layer=LI1_cond $X=0.24 $Y=1.597
+ $X2=0.24 $Y2=1.615
r29 15 16 19.7027 $w=1.68e-07 $l=3.02e-07 $layer=LI1_cond $X=0.24 $Y=1.295
+ $X2=0.24 $Y2=1.597
r30 14 15 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.24 $Y=0.925
+ $X2=0.24 $Y2=1.295
r31 13 38 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=0.24 $Y=0.43 $X2=0.36
+ $Y2=0.43
r32 13 24 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.24 $Y=0.43
+ $X2=0.24 $Y2=0.595
r33 13 14 20.0941 $w=1.68e-07 $l=3.08e-07 $layer=LI1_cond $X=0.24 $Y=0.617
+ $X2=0.24 $Y2=0.925
r34 13 24 1.43529 $w=1.68e-07 $l=2.2e-08 $layer=LI1_cond $X=0.24 $Y=0.617
+ $X2=0.24 $Y2=0.595
r35 8 16 11.8777 $w=3.03e-07 $l=2.8e-07 $layer=LI1_cond $X=0.605 $Y=1.7
+ $X2=0.325 $Y2=1.7
r36 7 11 10.4768 $w=3.28e-07 $l=3e-07 $layer=LI1_cond $X=0.77 $Y=1.7 $X2=0.77
+ $Y2=2
r37 7 8 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.77 $Y=1.7 $X2=0.605
+ $Y2=1.7
r38 2 11 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.63
+ $Y=1.855 $X2=0.77 $Y2=2
r39 1 38 182 $w=1.7e-07 $l=2.498e-07 $layer=licon1_NDIFF $count=1 $X=0.235
+ $Y=0.235 $X2=0.36 $Y2=0.43
.ends

.subckt PM_SKY130_FD_SC_LP__O41AI_M%A_175_47# 1 2 3 12 14 15 18 20 24 26
c45 18 0 1.48511e-19 $X=2.025 $Y=0.51
c46 12 0 1.4103e-19 $X=1.07 $Y=0.51
r47 22 24 9.04785 $w=1.88e-07 $l=1.55e-07 $layer=LI1_cond $X=2.915 $Y=0.665
+ $X2=2.915 $Y2=0.51
r48 21 26 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=2.13 $Y=0.75
+ $X2=2.025 $Y2=0.75
r49 20 22 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=2.82 $Y=0.75
+ $X2=2.915 $Y2=0.665
r50 20 21 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.82 $Y=0.75 $X2=2.13
+ $Y2=0.75
r51 16 26 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=2.025 $Y=0.665
+ $X2=2.025 $Y2=0.75
r52 16 18 8.18615 $w=2.08e-07 $l=1.55e-07 $layer=LI1_cond $X=2.025 $Y=0.665
+ $X2=2.025 $Y2=0.51
r53 14 26 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.92 $Y=0.75
+ $X2=2.025 $Y2=0.75
r54 14 15 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=1.92 $Y=0.75
+ $X2=1.155 $Y2=0.75
r55 10 15 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.07 $Y=0.665
+ $X2=1.155 $Y2=0.75
r56 10 12 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=1.07 $Y=0.665
+ $X2=1.07 $Y2=0.51
r57 3 24 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=2.765
+ $Y=0.235 $X2=2.905 $Y2=0.51
r58 2 18 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=1.885
+ $Y=0.235 $X2=2.025 $Y2=0.51
r59 1 12 182 $w=1.7e-07 $l=3.59514e-07 $layer=licon1_NDIFF $count=1 $X=0.875
+ $Y=0.235 $X2=1.07 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_LP__O41AI_M%VGND 1 2 9 13 16 17 19 20 21 34 35
r48 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r49 32 35 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r50 31 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r51 28 29 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r52 25 29 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r53 24 28 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r54 24 25 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r55 21 32 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r56 21 29 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r57 19 31 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=2.31 $Y=0 $X2=2.16
+ $Y2=0
r58 19 20 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.31 $Y=0 $X2=2.475
+ $Y2=0
r59 18 34 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r60 18 20 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.64 $Y=0 $X2=2.475
+ $Y2=0
r61 16 28 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=1.335 $Y=0 $X2=1.2
+ $Y2=0
r62 16 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.335 $Y=0 $X2=1.5
+ $Y2=0
r63 15 31 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=1.665 $Y=0 $X2=2.16
+ $Y2=0
r64 15 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.665 $Y=0 $X2=1.5
+ $Y2=0
r65 11 20 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.475 $Y=0.085
+ $X2=2.475 $Y2=0
r66 11 13 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.475 $Y=0.085
+ $X2=2.475 $Y2=0.38
r67 7 17 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.5 $Y=0.085 $X2=1.5
+ $Y2=0
r68 7 9 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.5 $Y=0.085 $X2=1.5
+ $Y2=0.38
r69 2 13 182 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_NDIFF $count=1 $X=2.315
+ $Y=0.235 $X2=2.475 $Y2=0.38
r70 1 9 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=1.36
+ $Y=0.235 $X2=1.5 $Y2=0.38
.ends

