* File: sky130_fd_sc_lp__a21oi_m.pex.spice
* Created: Wed Sep  2 09:20:57 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A21OI_M%A2 2 5 9 13 15 18 20 21 22 23 29
r39 22 23 20.0177 $w=2.03e-07 $l=3.7e-07 $layer=LI1_cond $X=0.257 $Y=1.665
+ $X2=0.257 $Y2=2.035
r40 21 22 20.0177 $w=2.03e-07 $l=3.7e-07 $layer=LI1_cond $X=0.257 $Y=1.295
+ $X2=0.257 $Y2=1.665
r41 20 21 20.0177 $w=2.03e-07 $l=3.7e-07 $layer=LI1_cond $X=0.257 $Y=0.925
+ $X2=0.257 $Y2=1.295
r42 20 29 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.275
+ $Y=1.005 $X2=0.275 $Y2=1.005
r43 16 18 71.7872 $w=1.5e-07 $l=1.4e-07 $layer=POLY_cond $X=0.335 $Y=2.215
+ $X2=0.475 $Y2=2.215
r44 14 29 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.275 $Y=1.345
+ $X2=0.275 $Y2=1.005
r45 14 15 41.8716 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.275 $Y=1.345
+ $X2=0.275 $Y2=1.51
r46 13 29 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=0.275 $Y=0.99
+ $X2=0.275 $Y2=1.005
r47 12 13 43.5886 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=0.35 $Y=0.84
+ $X2=0.35 $Y2=0.99
r48 9 12 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.515 $Y=0.445
+ $X2=0.515 $Y2=0.84
r49 3 18 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.475 $Y=2.29
+ $X2=0.475 $Y2=2.215
r50 3 5 225.617 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=0.475 $Y=2.29
+ $X2=0.475 $Y2=2.73
r51 2 16 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.335 $Y=2.14
+ $X2=0.335 $Y2=2.215
r52 2 15 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=0.335 $Y=2.14
+ $X2=0.335 $Y2=1.51
.ends

.subckt PM_SKY130_FD_SC_LP__A21OI_M%A1 3 7 11 12 13 14 15 16 22
r47 22 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.815
+ $Y=1.395 $X2=0.815 $Y2=1.395
r48 15 16 16.0907 $w=2.63e-07 $l=3.7e-07 $layer=LI1_cond $X=0.767 $Y=1.665
+ $X2=0.767 $Y2=2.035
r49 15 23 11.7419 $w=2.63e-07 $l=2.7e-07 $layer=LI1_cond $X=0.767 $Y=1.665
+ $X2=0.767 $Y2=1.395
r50 14 23 4.34884 $w=2.63e-07 $l=1e-07 $layer=LI1_cond $X=0.767 $Y=1.295
+ $X2=0.767 $Y2=1.395
r51 13 14 16.0907 $w=2.63e-07 $l=3.7e-07 $layer=LI1_cond $X=0.767 $Y=0.925
+ $X2=0.767 $Y2=1.295
r52 11 22 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.815 $Y=1.735
+ $X2=0.815 $Y2=1.395
r53 11 12 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.815 $Y=1.735
+ $X2=0.815 $Y2=1.9
r54 10 22 41.8716 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.815 $Y=1.23
+ $X2=0.815 $Y2=1.395
r55 7 12 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=0.905 $Y=2.73
+ $X2=0.905 $Y2=1.9
r56 3 10 402.521 $w=1.5e-07 $l=7.85e-07 $layer=POLY_cond $X=0.875 $Y=0.445
+ $X2=0.875 $Y2=1.23
.ends

.subckt PM_SKY130_FD_SC_LP__A21OI_M%B1 3 7 11 12 13 14 18 19
c38 12 0 3.09864e-20 $X=1.385 $Y=1.75
r39 18 19 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.385
+ $Y=1.245 $X2=1.385 $Y2=1.245
r40 13 14 12.0114 $w=3.53e-07 $l=3.7e-07 $layer=LI1_cond $X=1.292 $Y=1.295
+ $X2=1.292 $Y2=1.665
r41 13 19 1.62316 $w=3.53e-07 $l=5e-08 $layer=LI1_cond $X=1.292 $Y=1.295
+ $X2=1.292 $Y2=1.245
r42 11 18 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.385 $Y=1.585
+ $X2=1.385 $Y2=1.245
r43 11 12 40.8701 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.385 $Y=1.585
+ $X2=1.385 $Y2=1.75
r44 10 18 37.7798 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.385 $Y=1.08
+ $X2=1.385 $Y2=1.245
r45 7 10 325.606 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=1.38 $Y=0.445
+ $X2=1.38 $Y2=1.08
r46 3 12 502.511 $w=1.5e-07 $l=9.8e-07 $layer=POLY_cond $X=1.335 $Y=2.73
+ $X2=1.335 $Y2=1.75
.ends

.subckt PM_SKY130_FD_SC_LP__A21OI_M%A_27_504# 1 2 9 11 12 15
c24 11 0 3.09864e-20 $X=1.015 $Y=2.385
r25 13 15 9.24242 $w=2.08e-07 $l=1.75e-07 $layer=LI1_cond $X=1.12 $Y=2.47
+ $X2=1.12 $Y2=2.645
r26 11 13 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=1.015 $Y=2.385
+ $X2=1.12 $Y2=2.47
r27 11 12 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=1.015 $Y=2.385
+ $X2=0.365 $Y2=2.385
r28 7 12 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=0.26 $Y=2.47
+ $X2=0.365 $Y2=2.385
r29 7 9 10.2987 $w=2.08e-07 $l=1.95e-07 $layer=LI1_cond $X=0.26 $Y=2.47 $X2=0.26
+ $Y2=2.665
r30 2 15 600 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=0.98
+ $Y=2.52 $X2=1.12 $Y2=2.645
r31 1 9 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.52 $X2=0.26 $Y2=2.665
.ends

.subckt PM_SKY130_FD_SC_LP__A21OI_M%VPWR 1 6 8 10 17 18 21
r22 21 22 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r23 17 18 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r24 15 21 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=0.795 $Y=3.33
+ $X2=0.69 $Y2=3.33
r25 15 17 57.738 $w=1.68e-07 $l=8.85e-07 $layer=LI1_cond $X=0.795 $Y=3.33
+ $X2=1.68 $Y2=3.33
r26 13 22 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r27 12 13 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r28 10 21 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=0.585 $Y=3.33
+ $X2=0.69 $Y2=3.33
r29 10 12 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.585 $Y=3.33
+ $X2=0.24 $Y2=3.33
r30 8 18 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=0.96 $Y=3.33
+ $X2=1.68 $Y2=3.33
r31 8 22 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=0.96 $Y=3.33
+ $X2=0.72 $Y2=3.33
r32 4 21 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=3.245
+ $X2=0.69 $Y2=3.33
r33 4 6 22.71 $w=2.08e-07 $l=4.3e-07 $layer=LI1_cond $X=0.69 $Y=3.245 $X2=0.69
+ $Y2=2.815
r34 1 6 600 $w=1.7e-07 $l=3.58225e-07 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=2.52 $X2=0.69 $Y2=2.815
.ends

.subckt PM_SKY130_FD_SC_LP__A21OI_M%Y 1 2 9 11 12 14 15 22
c28 9 0 1.71582e-19 $X=1.165 $Y=0.51
r29 15 22 1.92074 $w=3.28e-07 $l=5.5e-08 $layer=LI1_cond $X=1.68 $Y=2.695
+ $X2=1.735 $Y2=2.695
r30 15 18 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=1.68 $Y=2.695
+ $X2=1.55 $Y2=2.695
r31 14 22 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.735 $Y=2.53
+ $X2=1.735 $Y2=2.695
r32 13 14 110.583 $w=1.68e-07 $l=1.695e-06 $layer=LI1_cond $X=1.735 $Y=0.835
+ $X2=1.735 $Y2=2.53
r33 11 13 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.65 $Y=0.75
+ $X2=1.735 $Y2=0.835
r34 11 12 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=1.65 $Y=0.75 $X2=1.25
+ $Y2=0.75
r35 7 12 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.165 $Y=0.665
+ $X2=1.25 $Y2=0.75
r36 7 9 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=1.165 $Y=0.665
+ $X2=1.165 $Y2=0.51
r37 2 18 600 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_PDIFF $count=1 $X=1.41
+ $Y=2.52 $X2=1.55 $Y2=2.695
r38 1 9 182 $w=1.7e-07 $l=3.67083e-07 $layer=licon1_NDIFF $count=1 $X=0.95
+ $Y=0.235 $X2=1.165 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_LP__A21OI_M%VGND 1 2 7 9 11 13 15 17 27
r28 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r29 23 24 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r30 21 27 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r31 20 21 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r32 18 23 3.63675 $w=1.7e-07 $l=2.03e-07 $layer=LI1_cond $X=0.405 $Y=0 $X2=0.202
+ $Y2=0
r33 18 20 51.8663 $w=1.68e-07 $l=7.95e-07 $layer=LI1_cond $X=0.405 $Y=0 $X2=1.2
+ $Y2=0
r34 17 26 4.64076 $w=1.7e-07 $l=2.45e-07 $layer=LI1_cond $X=1.43 $Y=0 $X2=1.675
+ $Y2=0
r35 17 20 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=1.43 $Y=0 $X2=1.2
+ $Y2=0
r36 15 21 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=0.96 $Y=0 $X2=1.2
+ $Y2=0
r37 15 24 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=0.96 $Y=0 $X2=0.24
+ $Y2=0
r38 11 26 3.12541 $w=3.3e-07 $l=1.18427e-07 $layer=LI1_cond $X=1.595 $Y=0.085
+ $X2=1.675 $Y2=0
r39 11 13 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.595 $Y=0.085
+ $X2=1.595 $Y2=0.38
r40 7 23 3.27845 $w=2.1e-07 $l=1.33918e-07 $layer=LI1_cond $X=0.3 $Y=0.085
+ $X2=0.202 $Y2=0
r41 7 9 15.5801 $w=2.08e-07 $l=2.95e-07 $layer=LI1_cond $X=0.3 $Y=0.085 $X2=0.3
+ $Y2=0.38
r42 2 13 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=1.455
+ $Y=0.235 $X2=1.595 $Y2=0.38
r43 1 9 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.175
+ $Y=0.235 $X2=0.3 $Y2=0.38
.ends

