* File: sky130_fd_sc_lp__clkbuflp_4.pxi.spice
* Created: Wed Sep  2 09:39:07 2020
* 
x_PM_SKY130_FD_SC_LP__CLKBUFLP_4%A N_A_M1006_g N_A_M1005_g N_A_M1000_g
+ N_A_M1010_g A A N_A_c_65_n PM_SKY130_FD_SC_LP__CLKBUFLP_4%A
x_PM_SKY130_FD_SC_LP__CLKBUFLP_4%A_130_417# N_A_130_417#_M1000_d
+ N_A_130_417#_M1005_s N_A_130_417#_M1001_g N_A_130_417#_M1002_g
+ N_A_130_417#_M1008_g N_A_130_417#_M1003_g N_A_130_417#_M1007_g
+ N_A_130_417#_M1009_g N_A_130_417#_M1004_g N_A_130_417#_M1011_g
+ N_A_130_417#_c_126_n N_A_130_417#_c_114_n N_A_130_417#_c_115_n
+ N_A_130_417#_c_123_n N_A_130_417#_c_116_n N_A_130_417#_c_117_n
+ N_A_130_417#_c_118_n PM_SKY130_FD_SC_LP__CLKBUFLP_4%A_130_417#
x_PM_SKY130_FD_SC_LP__CLKBUFLP_4%VPWR N_VPWR_M1005_d N_VPWR_M1010_d
+ N_VPWR_M1008_d N_VPWR_M1011_d N_VPWR_c_222_n N_VPWR_c_223_n N_VPWR_c_224_n
+ N_VPWR_c_225_n N_VPWR_c_226_n N_VPWR_c_227_n N_VPWR_c_228_n N_VPWR_c_229_n
+ N_VPWR_c_230_n N_VPWR_c_231_n VPWR N_VPWR_c_232_n N_VPWR_c_221_n
+ PM_SKY130_FD_SC_LP__CLKBUFLP_4%VPWR
x_PM_SKY130_FD_SC_LP__CLKBUFLP_4%X N_X_M1003_s N_X_M1001_s N_X_M1009_s
+ N_X_c_285_n N_X_c_280_n N_X_c_281_n X X X X X X N_X_c_305_n N_X_c_283_n
+ N_X_c_279_n PM_SKY130_FD_SC_LP__CLKBUFLP_4%X
x_PM_SKY130_FD_SC_LP__CLKBUFLP_4%VGND N_VGND_M1006_s N_VGND_M1002_d
+ N_VGND_M1004_d N_VGND_c_341_n N_VGND_c_342_n N_VGND_c_343_n N_VGND_c_344_n
+ VGND N_VGND_c_345_n N_VGND_c_346_n N_VGND_c_347_n N_VGND_c_348_n
+ N_VGND_c_349_n N_VGND_c_350_n PM_SKY130_FD_SC_LP__CLKBUFLP_4%VGND
cc_1 VNB N_A_M1006_g 0.0371616f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.555
cc_2 VNB N_A_M1005_g 0.00644544f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=2.585
cc_3 VNB N_A_M1000_g 0.0337887f $X=-0.19 $Y=-0.245 $X2=0.835 $Y2=0.555
cc_4 VNB N_A_M1010_g 0.00527519f $X=-0.19 $Y=-0.245 $X2=1.055 $Y2=2.585
cc_5 VNB A 0.0321953f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_6 VNB N_A_c_65_n 0.0532012f $X=-0.19 $Y=-0.245 $X2=1.055 $Y2=1.4
cc_7 VNB N_A_130_417#_M1001_g 0.00690599f $X=-0.19 $Y=-0.245 $X2=0.835 $Y2=1.235
cc_8 VNB N_A_130_417#_M1002_g 0.0363957f $X=-0.19 $Y=-0.245 $X2=1.055 $Y2=1.565
cc_9 VNB N_A_130_417#_M1008_g 0.00666918f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_10 VNB N_A_130_417#_M1003_g 0.0301622f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.4
cc_11 VNB N_A_130_417#_M1007_g 0.0266424f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=1.4
cc_12 VNB N_A_130_417#_M1009_g 0.00578869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_130_417#_M1004_g 0.0436494f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.665
cc_14 VNB N_A_130_417#_M1011_g 0.00745847f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_130_417#_c_114_n 0.0129998f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_130_417#_c_115_n 0.0108178f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_130_417#_c_116_n 8.06543e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_130_417#_c_117_n 0.00203637f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_130_417#_c_118_n 0.111445f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_VPWR_c_221_n 0.163682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB X 0.00865464f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=1.4
cc_22 VNB X 0.0451127f $X=-0.19 $Y=-0.245 $X2=0.42 $Y2=1.295
cc_23 VNB N_X_c_279_n 0.00685644f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_VGND_c_341_n 0.0107456f $X=-0.19 $Y=-0.245 $X2=0.835 $Y2=0.555
cc_25 VNB N_VGND_c_342_n 0.02995f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_343_n 0.00724798f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_344_n 0.0193592f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_345_n 0.0267208f $X=-0.19 $Y=-0.245 $X2=0.565 $Y2=1.4
cc_29 VNB N_VGND_c_346_n 0.0328783f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_347_n 0.0188498f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_348_n 0.234131f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_349_n 0.00513431f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_350_n 0.00513431f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VPB N_A_M1005_g 0.0549057f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=2.585
cc_35 VPB N_A_M1010_g 0.0414578f $X=-0.19 $Y=1.655 $X2=1.055 $Y2=2.585
cc_36 VPB A 0.0081482f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_37 VPB N_A_130_417#_M1001_g 0.0412785f $X=-0.19 $Y=1.655 $X2=0.835 $Y2=1.235
cc_38 VPB N_A_130_417#_M1008_g 0.039811f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_39 VPB N_A_130_417#_M1009_g 0.0394204f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_40 VPB N_A_130_417#_M1011_g 0.0534647f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_41 VPB N_A_130_417#_c_123_n 0.00533931f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_42 VPB N_A_130_417#_c_116_n 0.00398282f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_43 VPB N_VPWR_c_222_n 0.0107197f $X=-0.19 $Y=1.655 $X2=1.055 $Y2=1.565
cc_44 VPB N_VPWR_c_223_n 0.0439499f $X=-0.19 $Y=1.655 $X2=1.055 $Y2=2.585
cc_45 VPB N_VPWR_c_224_n 0.00622359f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=1.4
cc_46 VPB N_VPWR_c_225_n 0.00195694f $X=-0.19 $Y=1.655 $X2=0.835 $Y2=1.4
cc_47 VPB N_VPWR_c_226_n 0.0148055f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_48 VPB N_VPWR_c_227_n 0.0446022f $X=-0.19 $Y=1.655 $X2=0.24 $Y2=1.665
cc_49 VPB N_VPWR_c_228_n 0.0201143f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_50 VPB N_VPWR_c_229_n 0.00375865f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_51 VPB N_VPWR_c_230_n 0.0178633f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_52 VPB N_VPWR_c_231_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_53 VPB N_VPWR_c_232_n 0.0178633f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_54 VPB N_VPWR_c_221_n 0.050578f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_55 VPB N_X_c_280_n 0.00230158f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_56 VPB N_X_c_281_n 7.23973e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_57 VPB X 0.0157477f $X=-0.19 $Y=1.655 $X2=0.42 $Y2=1.295
cc_58 VPB N_X_c_283_n 0.00444666f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_59 VPB N_X_c_279_n 0.00302133f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_60 N_A_M1010_g N_A_130_417#_M1001_g 0.022949f $X=1.055 $Y=2.585 $X2=0 $Y2=0
cc_61 N_A_M1005_g N_A_130_417#_c_126_n 0.0142364f $X=0.525 $Y=2.585 $X2=0 $Y2=0
cc_62 N_A_M1010_g N_A_130_417#_c_126_n 0.0165535f $X=1.055 $Y=2.585 $X2=0 $Y2=0
cc_63 N_A_M1006_g N_A_130_417#_c_114_n 0.0029976f $X=0.475 $Y=0.555 $X2=0 $Y2=0
cc_64 N_A_M1000_g N_A_130_417#_c_114_n 0.0219672f $X=0.835 $Y=0.555 $X2=0 $Y2=0
cc_65 A N_A_130_417#_c_114_n 0.00581356f $X=0.155 $Y=1.58 $X2=0 $Y2=0
cc_66 N_A_M1005_g N_A_130_417#_c_123_n 0.00466227f $X=0.525 $Y=2.585 $X2=0 $Y2=0
cc_67 N_A_M1010_g N_A_130_417#_c_123_n 0.00442588f $X=1.055 $Y=2.585 $X2=0 $Y2=0
cc_68 A N_A_130_417#_c_123_n 0.00330371f $X=0.155 $Y=1.58 $X2=0 $Y2=0
cc_69 N_A_c_65_n N_A_130_417#_c_123_n 0.00342304f $X=1.055 $Y=1.4 $X2=0 $Y2=0
cc_70 N_A_M1005_g N_A_130_417#_c_116_n 0.00727613f $X=0.525 $Y=2.585 $X2=0 $Y2=0
cc_71 N_A_M1010_g N_A_130_417#_c_116_n 0.0161008f $X=1.055 $Y=2.585 $X2=0 $Y2=0
cc_72 A N_A_130_417#_c_116_n 0.00960507f $X=0.155 $Y=1.58 $X2=0 $Y2=0
cc_73 N_A_c_65_n N_A_130_417#_c_116_n 0.00128669f $X=1.055 $Y=1.4 $X2=0 $Y2=0
cc_74 N_A_M1000_g N_A_130_417#_c_117_n 8.29209e-19 $X=0.835 $Y=0.555 $X2=0 $Y2=0
cc_75 A N_A_130_417#_c_117_n 0.0277261f $X=0.155 $Y=1.58 $X2=0 $Y2=0
cc_76 N_A_c_65_n N_A_130_417#_c_117_n 0.0295332f $X=1.055 $Y=1.4 $X2=0 $Y2=0
cc_77 N_A_M1000_g N_A_130_417#_c_118_n 4.88583e-19 $X=0.835 $Y=0.555 $X2=0 $Y2=0
cc_78 N_A_c_65_n N_A_130_417#_c_118_n 0.022949f $X=1.055 $Y=1.4 $X2=0 $Y2=0
cc_79 N_A_M1005_g N_VPWR_c_223_n 0.0243876f $X=0.525 $Y=2.585 $X2=0 $Y2=0
cc_80 N_A_M1010_g N_VPWR_c_223_n 0.00118407f $X=1.055 $Y=2.585 $X2=0 $Y2=0
cc_81 A N_VPWR_c_223_n 0.0188297f $X=0.155 $Y=1.58 $X2=0 $Y2=0
cc_82 N_A_M1010_g N_VPWR_c_224_n 0.00321157f $X=1.055 $Y=2.585 $X2=0 $Y2=0
cc_83 N_A_M1005_g N_VPWR_c_228_n 0.00839865f $X=0.525 $Y=2.585 $X2=0 $Y2=0
cc_84 N_A_M1010_g N_VPWR_c_228_n 0.00787395f $X=1.055 $Y=2.585 $X2=0 $Y2=0
cc_85 N_A_M1005_g N_VPWR_c_221_n 0.0136348f $X=0.525 $Y=2.585 $X2=0 $Y2=0
cc_86 N_A_M1010_g N_VPWR_c_221_n 0.012393f $X=1.055 $Y=2.585 $X2=0 $Y2=0
cc_87 N_A_M1010_g N_X_c_285_n 7.78968e-19 $X=1.055 $Y=2.585 $X2=0 $Y2=0
cc_88 N_A_M1010_g N_X_c_280_n 4.65654e-19 $X=1.055 $Y=2.585 $X2=0 $Y2=0
cc_89 N_A_M1006_g N_VGND_c_342_n 0.0171478f $X=0.475 $Y=0.555 $X2=0 $Y2=0
cc_90 N_A_M1000_g N_VGND_c_342_n 0.00296662f $X=0.835 $Y=0.555 $X2=0 $Y2=0
cc_91 A N_VGND_c_342_n 0.0215578f $X=0.155 $Y=1.58 $X2=0 $Y2=0
cc_92 N_A_M1000_g N_VGND_c_343_n 0.00230008f $X=0.835 $Y=0.555 $X2=0 $Y2=0
cc_93 N_A_M1006_g N_VGND_c_345_n 0.00486043f $X=0.475 $Y=0.555 $X2=0 $Y2=0
cc_94 N_A_M1000_g N_VGND_c_345_n 0.0054895f $X=0.835 $Y=0.555 $X2=0 $Y2=0
cc_95 N_A_M1006_g N_VGND_c_348_n 0.00814425f $X=0.475 $Y=0.555 $X2=0 $Y2=0
cc_96 N_A_M1000_g N_VGND_c_348_n 0.0111095f $X=0.835 $Y=0.555 $X2=0 $Y2=0
cc_97 N_A_130_417#_c_123_n N_VPWR_c_223_n 0.0674082f $X=0.79 $Y=2.23 $X2=0 $Y2=0
cc_98 N_A_130_417#_M1001_g N_VPWR_c_224_n 0.0227327f $X=1.585 $Y=2.585 $X2=0
+ $Y2=0
cc_99 N_A_130_417#_M1008_g N_VPWR_c_224_n 0.00117568f $X=2.115 $Y=2.585 $X2=0
+ $Y2=0
cc_100 N_A_130_417#_c_115_n N_VPWR_c_224_n 0.00996389f $X=1.965 $Y=1.37 $X2=0
+ $Y2=0
cc_101 N_A_130_417#_c_123_n N_VPWR_c_224_n 0.0401872f $X=0.79 $Y=2.23 $X2=0
+ $Y2=0
cc_102 N_A_130_417#_M1001_g N_VPWR_c_225_n 9.25377e-19 $X=1.585 $Y=2.585 $X2=0
+ $Y2=0
cc_103 N_A_130_417#_M1008_g N_VPWR_c_225_n 0.0224727f $X=2.115 $Y=2.585 $X2=0
+ $Y2=0
cc_104 N_A_130_417#_M1009_g N_VPWR_c_225_n 0.0224727f $X=2.645 $Y=2.585 $X2=0
+ $Y2=0
cc_105 N_A_130_417#_M1011_g N_VPWR_c_225_n 9.25377e-19 $X=3.175 $Y=2.585 $X2=0
+ $Y2=0
cc_106 N_A_130_417#_c_118_n N_VPWR_c_225_n 3.00486e-19 $X=3.175 $Y=1.375 $X2=0
+ $Y2=0
cc_107 N_A_130_417#_M1009_g N_VPWR_c_227_n 9.25377e-19 $X=2.645 $Y=2.585 $X2=0
+ $Y2=0
cc_108 N_A_130_417#_M1011_g N_VPWR_c_227_n 0.0236961f $X=3.175 $Y=2.585 $X2=0
+ $Y2=0
cc_109 N_A_130_417#_c_126_n N_VPWR_c_228_n 0.0257409f $X=0.79 $Y=2.91 $X2=0
+ $Y2=0
cc_110 N_A_130_417#_M1001_g N_VPWR_c_230_n 0.00839865f $X=1.585 $Y=2.585 $X2=0
+ $Y2=0
cc_111 N_A_130_417#_M1008_g N_VPWR_c_230_n 0.00839865f $X=2.115 $Y=2.585 $X2=0
+ $Y2=0
cc_112 N_A_130_417#_M1009_g N_VPWR_c_232_n 0.00839865f $X=2.645 $Y=2.585 $X2=0
+ $Y2=0
cc_113 N_A_130_417#_M1011_g N_VPWR_c_232_n 0.00839865f $X=3.175 $Y=2.585 $X2=0
+ $Y2=0
cc_114 N_A_130_417#_M1005_s N_VPWR_c_221_n 0.00223559f $X=0.65 $Y=2.085 $X2=0
+ $Y2=0
cc_115 N_A_130_417#_M1001_g N_VPWR_c_221_n 0.0136348f $X=1.585 $Y=2.585 $X2=0
+ $Y2=0
cc_116 N_A_130_417#_M1008_g N_VPWR_c_221_n 0.0136348f $X=2.115 $Y=2.585 $X2=0
+ $Y2=0
cc_117 N_A_130_417#_M1009_g N_VPWR_c_221_n 0.0136348f $X=2.645 $Y=2.585 $X2=0
+ $Y2=0
cc_118 N_A_130_417#_M1011_g N_VPWR_c_221_n 0.0136348f $X=3.175 $Y=2.585 $X2=0
+ $Y2=0
cc_119 N_A_130_417#_c_126_n N_VPWR_c_221_n 0.0158161f $X=0.79 $Y=2.91 $X2=0
+ $Y2=0
cc_120 N_A_130_417#_M1001_g N_X_c_285_n 0.0236657f $X=1.585 $Y=2.585 $X2=0 $Y2=0
cc_121 N_A_130_417#_M1008_g N_X_c_285_n 0.0235159f $X=2.115 $Y=2.585 $X2=0 $Y2=0
cc_122 N_A_130_417#_M1009_g N_X_c_285_n 8.9921e-19 $X=2.645 $Y=2.585 $X2=0 $Y2=0
cc_123 N_A_130_417#_c_116_n N_X_c_285_n 0.00454232f $X=0.84 $Y=2.065 $X2=0 $Y2=0
cc_124 N_A_130_417#_M1001_g N_X_c_280_n 0.00606303f $X=1.585 $Y=2.585 $X2=0
+ $Y2=0
cc_125 N_A_130_417#_M1008_g N_X_c_280_n 0.00279308f $X=2.115 $Y=2.585 $X2=0
+ $Y2=0
cc_126 N_A_130_417#_c_115_n N_X_c_280_n 0.027608f $X=1.965 $Y=1.37 $X2=0 $Y2=0
cc_127 N_A_130_417#_c_116_n N_X_c_280_n 0.00434411f $X=0.84 $Y=2.065 $X2=0 $Y2=0
cc_128 N_A_130_417#_c_118_n N_X_c_280_n 0.00275645f $X=3.175 $Y=1.375 $X2=0
+ $Y2=0
cc_129 N_A_130_417#_M1008_g N_X_c_281_n 9.0147e-19 $X=2.115 $Y=2.585 $X2=0 $Y2=0
cc_130 N_A_130_417#_M1009_g N_X_c_281_n 0.0236239f $X=2.645 $Y=2.585 $X2=0 $Y2=0
cc_131 N_A_130_417#_M1011_g N_X_c_281_n 0.0294748f $X=3.175 $Y=2.585 $X2=0 $Y2=0
cc_132 N_A_130_417#_c_118_n N_X_c_281_n 3.1299e-19 $X=3.175 $Y=1.375 $X2=0 $Y2=0
cc_133 N_A_130_417#_M1003_g X 0.0131321f $X=2.145 $Y=0.51 $X2=0 $Y2=0
cc_134 N_A_130_417#_M1007_g X 0.0138274f $X=2.575 $Y=0.51 $X2=0 $Y2=0
cc_135 N_A_130_417#_c_118_n X 9.15772e-19 $X=3.175 $Y=1.375 $X2=0 $Y2=0
cc_136 N_A_130_417#_M1011_g X 0.0211949f $X=3.175 $Y=2.585 $X2=0 $Y2=0
cc_137 N_A_130_417#_c_118_n X 0.0179061f $X=3.175 $Y=1.375 $X2=0 $Y2=0
cc_138 N_A_130_417#_M1002_g N_X_c_305_n 8.94287e-19 $X=1.785 $Y=0.51 $X2=0 $Y2=0
cc_139 N_A_130_417#_M1003_g N_X_c_305_n 0.00662055f $X=2.145 $Y=0.51 $X2=0 $Y2=0
cc_140 N_A_130_417#_M1007_g N_X_c_305_n 0.00801674f $X=2.575 $Y=0.51 $X2=0 $Y2=0
cc_141 N_A_130_417#_M1004_g N_X_c_305_n 0.0160006f $X=2.935 $Y=0.51 $X2=0 $Y2=0
cc_142 N_A_130_417#_c_118_n N_X_c_305_n 0.00128119f $X=3.175 $Y=1.375 $X2=0
+ $Y2=0
cc_143 N_A_130_417#_M1008_g N_X_c_283_n 0.0211879f $X=2.115 $Y=2.585 $X2=0 $Y2=0
cc_144 N_A_130_417#_c_115_n N_X_c_283_n 0.00817855f $X=1.965 $Y=1.37 $X2=0 $Y2=0
cc_145 N_A_130_417#_c_118_n N_X_c_283_n 9.35333e-19 $X=3.175 $Y=1.375 $X2=0
+ $Y2=0
cc_146 N_A_130_417#_M1008_g N_X_c_279_n 0.00477565f $X=2.115 $Y=2.585 $X2=0
+ $Y2=0
cc_147 N_A_130_417#_M1003_g N_X_c_279_n 9.72672e-19 $X=2.145 $Y=0.51 $X2=0 $Y2=0
cc_148 N_A_130_417#_M1007_g N_X_c_279_n 0.00148077f $X=2.575 $Y=0.51 $X2=0 $Y2=0
cc_149 N_A_130_417#_M1009_g N_X_c_279_n 0.0258871f $X=2.645 $Y=2.585 $X2=0 $Y2=0
cc_150 N_A_130_417#_M1004_g N_X_c_279_n 0.00876684f $X=2.935 $Y=0.51 $X2=0 $Y2=0
cc_151 N_A_130_417#_M1011_g N_X_c_279_n 0.00860892f $X=3.175 $Y=2.585 $X2=0
+ $Y2=0
cc_152 N_A_130_417#_c_115_n N_X_c_279_n 0.0221393f $X=1.965 $Y=1.37 $X2=0 $Y2=0
cc_153 N_A_130_417#_c_118_n N_X_c_279_n 0.0349052f $X=3.175 $Y=1.375 $X2=0 $Y2=0
cc_154 N_A_130_417#_c_114_n N_VGND_c_342_n 0.0213307f $X=1.05 $Y=0.39 $X2=0
+ $Y2=0
cc_155 N_A_130_417#_M1002_g N_VGND_c_343_n 0.0145684f $X=1.785 $Y=0.51 $X2=0
+ $Y2=0
cc_156 N_A_130_417#_M1003_g N_VGND_c_343_n 0.00248113f $X=2.145 $Y=0.51 $X2=0
+ $Y2=0
cc_157 N_A_130_417#_c_114_n N_VGND_c_343_n 0.032743f $X=1.05 $Y=0.39 $X2=0 $Y2=0
cc_158 N_A_130_417#_c_115_n N_VGND_c_343_n 0.0099824f $X=1.965 $Y=1.37 $X2=0
+ $Y2=0
cc_159 N_A_130_417#_c_118_n N_VGND_c_343_n 0.00491971f $X=3.175 $Y=1.375 $X2=0
+ $Y2=0
cc_160 N_A_130_417#_M1007_g N_VGND_c_344_n 0.0018613f $X=2.575 $Y=0.51 $X2=0
+ $Y2=0
cc_161 N_A_130_417#_M1004_g N_VGND_c_344_n 0.0128807f $X=2.935 $Y=0.51 $X2=0
+ $Y2=0
cc_162 N_A_130_417#_c_118_n N_VGND_c_344_n 0.00158209f $X=3.175 $Y=1.375 $X2=0
+ $Y2=0
cc_163 N_A_130_417#_c_114_n N_VGND_c_345_n 0.022122f $X=1.05 $Y=0.39 $X2=0 $Y2=0
cc_164 N_A_130_417#_M1002_g N_VGND_c_346_n 0.00486043f $X=1.785 $Y=0.51 $X2=0
+ $Y2=0
cc_165 N_A_130_417#_M1003_g N_VGND_c_346_n 0.00551226f $X=2.145 $Y=0.51 $X2=0
+ $Y2=0
cc_166 N_A_130_417#_M1007_g N_VGND_c_346_n 0.00371894f $X=2.575 $Y=0.51 $X2=0
+ $Y2=0
cc_167 N_A_130_417#_M1004_g N_VGND_c_346_n 0.00486043f $X=2.935 $Y=0.51 $X2=0
+ $Y2=0
cc_168 N_A_130_417#_M1000_d N_VGND_c_348_n 0.00215158f $X=0.91 $Y=0.235 $X2=0
+ $Y2=0
cc_169 N_A_130_417#_M1002_g N_VGND_c_348_n 0.00814425f $X=1.785 $Y=0.51 $X2=0
+ $Y2=0
cc_170 N_A_130_417#_M1003_g N_VGND_c_348_n 0.00988581f $X=2.145 $Y=0.51 $X2=0
+ $Y2=0
cc_171 N_A_130_417#_M1007_g N_VGND_c_348_n 0.00524368f $X=2.575 $Y=0.51 $X2=0
+ $Y2=0
cc_172 N_A_130_417#_M1004_g N_VGND_c_348_n 0.00814425f $X=2.935 $Y=0.51 $X2=0
+ $Y2=0
cc_173 N_A_130_417#_c_114_n N_VGND_c_348_n 0.0131521f $X=1.05 $Y=0.39 $X2=0
+ $Y2=0
cc_174 N_VPWR_c_221_n N_X_M1001_s 0.00223559f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_175 N_VPWR_c_221_n N_X_M1009_s 0.00223559f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_176 N_VPWR_c_224_n N_X_c_285_n 0.065356f $X=1.32 $Y=2.23 $X2=0 $Y2=0
cc_177 N_VPWR_c_225_n N_X_c_285_n 0.0652318f $X=2.38 $Y=2.23 $X2=0 $Y2=0
cc_178 N_VPWR_c_230_n N_X_c_285_n 0.0189236f $X=2.215 $Y=3.33 $X2=0 $Y2=0
cc_179 N_VPWR_c_221_n N_X_c_285_n 0.0123859f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_180 N_VPWR_c_225_n N_X_c_281_n 0.0652318f $X=2.38 $Y=2.23 $X2=0 $Y2=0
cc_181 N_VPWR_c_227_n N_X_c_281_n 0.0652318f $X=3.44 $Y=2.23 $X2=0 $Y2=0
cc_182 N_VPWR_c_232_n N_X_c_281_n 0.0189236f $X=3.275 $Y=3.33 $X2=0 $Y2=0
cc_183 N_VPWR_c_221_n N_X_c_281_n 0.0123859f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_184 N_VPWR_c_227_n X 0.0182353f $X=3.44 $Y=2.23 $X2=0 $Y2=0
cc_185 N_VPWR_c_225_n N_X_c_283_n 0.0199276f $X=2.38 $Y=2.23 $X2=0 $Y2=0
cc_186 N_X_c_305_n N_VGND_c_343_n 0.011538f $X=2.36 $Y=0.49 $X2=0 $Y2=0
cc_187 N_X_c_305_n N_VGND_c_344_n 0.0227658f $X=2.36 $Y=0.49 $X2=0 $Y2=0
cc_188 N_X_c_279_n N_VGND_c_344_n 0.0122118f $X=3.075 $Y=1.522 $X2=0 $Y2=0
cc_189 N_X_c_305_n N_VGND_c_346_n 0.0233911f $X=2.36 $Y=0.49 $X2=0 $Y2=0
cc_190 N_X_M1003_s N_VGND_c_348_n 0.00230594f $X=2.22 $Y=0.235 $X2=0 $Y2=0
cc_191 N_X_c_305_n N_VGND_c_348_n 0.0206818f $X=2.36 $Y=0.49 $X2=0 $Y2=0
cc_192 X A_530_47# 0.00159552f $X=2.555 $Y=0.84 $X2=-0.19 $Y2=-0.245
cc_193 N_X_c_305_n A_530_47# 0.00379922f $X=2.36 $Y=0.49 $X2=-0.19 $Y2=-0.245
cc_194 N_VGND_c_348_n A_110_47# 0.00899413f $X=3.6 $Y=0 $X2=-0.19 $Y2=-0.245
cc_195 N_VGND_c_348_n A_372_47# 0.00899413f $X=3.6 $Y=0 $X2=-0.19 $Y2=-0.245
cc_196 N_VGND_c_348_n A_530_47# 0.00470451f $X=3.6 $Y=0 $X2=-0.19 $Y2=-0.245
