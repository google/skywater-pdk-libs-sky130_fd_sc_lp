* File: sky130_fd_sc_lp__nor2b_m.spice
* Created: Fri Aug 28 10:54:59 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__nor2b_m.pex.spice"
.subckt sky130_fd_sc_lp__nor2b_m  VNB VPB B_N A VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A	A
* B_N	B_N
* VPB	VPB
* VNB	VNB
MM1003 N_VGND_M1003_d N_B_N_M1003_g N_A_47_70#_M1003_s VNB NSHORT L=0.15 W=0.42
+ AD=0.1176 AS=0.1113 PD=0.98 PS=1.37 NRD=79.992 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.3 A=0.063 P=1.14 MULT=1
MM1005 N_Y_M1005_d N_A_M1005_g N_VGND_M1003_d VNB NSHORT L=0.15 W=0.42 AD=0.0588
+ AS=0.1176 PD=0.7 PS=0.98 NRD=0 NRS=0 M=1 R=2.8 SA=75000.9 SB=75000.6 A=0.063
+ P=1.14 MULT=1
MM1002 N_VGND_M1002_d N_A_47_70#_M1002_g N_Y_M1005_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0588 PD=1.41 PS=0.7 NRD=5.712 NRS=0 M=1 R=2.8 SA=75001.3
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1004 N_VPWR_M1004_d N_B_N_M1004_g N_A_47_70#_M1004_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.09135 AS=0.1197 PD=0.855 PS=1.41 NRD=28.1316 NRS=9.3772 M=1 R=2.8
+ SA=75000.2 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1001 A_328_492# N_A_M1001_g N_VPWR_M1004_d VPB PHIGHVT L=0.15 W=0.42 AD=0.0441
+ AS=0.09135 PD=0.63 PS=0.855 NRD=23.443 NRS=44.5417 M=1 R=2.8 SA=75000.8
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1000 N_Y_M1000_d N_A_47_70#_M1000_g A_328_492# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.1113 AS=0.0441 PD=1.37 PS=0.63 NRD=0 NRS=23.443 M=1 R=2.8 SA=75001.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
DX6_noxref VNB VPB NWDIODE A=5.1847 P=9.29
*
.include "sky130_fd_sc_lp__nor2b_m.pxi.spice"
*
.ends
*
*
