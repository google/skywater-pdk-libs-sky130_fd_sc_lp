* File: sky130_fd_sc_lp__o221ai_1.pxi.spice
* Created: Wed Sep  2 10:19:04 2020
* 
x_PM_SKY130_FD_SC_LP__O221AI_1%C1 N_C1_M1002_g N_C1_M1000_g C1 N_C1_c_61_n
+ N_C1_c_62_n PM_SKY130_FD_SC_LP__O221AI_1%C1
x_PM_SKY130_FD_SC_LP__O221AI_1%B1 N_B1_M1008_g N_B1_M1007_g B1 N_B1_c_90_n
+ N_B1_c_91_n PM_SKY130_FD_SC_LP__O221AI_1%B1
x_PM_SKY130_FD_SC_LP__O221AI_1%B2 N_B2_M1009_g N_B2_M1001_g B2 N_B2_c_127_n
+ N_B2_c_128_n PM_SKY130_FD_SC_LP__O221AI_1%B2
x_PM_SKY130_FD_SC_LP__O221AI_1%A2 N_A2_M1006_g N_A2_M1004_g A2 A2 A2 A2
+ N_A2_c_166_n PM_SKY130_FD_SC_LP__O221AI_1%A2
x_PM_SKY130_FD_SC_LP__O221AI_1%A1 N_A1_M1003_g N_A1_M1005_g A1 N_A1_c_207_n
+ N_A1_c_208_n PM_SKY130_FD_SC_LP__O221AI_1%A1
x_PM_SKY130_FD_SC_LP__O221AI_1%Y N_Y_M1002_s N_Y_M1000_s N_Y_M1009_d N_Y_c_233_n
+ N_Y_c_229_n N_Y_c_249_n N_Y_c_260_n N_Y_c_262_n Y Y Y Y Y N_Y_c_231_n
+ N_Y_c_232_n Y N_Y_c_235_n PM_SKY130_FD_SC_LP__O221AI_1%Y
x_PM_SKY130_FD_SC_LP__O221AI_1%VPWR N_VPWR_M1000_d N_VPWR_M1005_d N_VPWR_c_289_n
+ N_VPWR_c_290_n N_VPWR_c_291_n VPWR N_VPWR_c_292_n N_VPWR_c_293_n
+ N_VPWR_c_294_n N_VPWR_c_288_n PM_SKY130_FD_SC_LP__O221AI_1%VPWR
x_PM_SKY130_FD_SC_LP__O221AI_1%A_114_47# N_A_114_47#_M1002_d N_A_114_47#_M1008_d
+ N_A_114_47#_c_334_n N_A_114_47#_c_335_n N_A_114_47#_c_348_p
+ PM_SKY130_FD_SC_LP__O221AI_1%A_114_47#
x_PM_SKY130_FD_SC_LP__O221AI_1%A_221_49# N_A_221_49#_M1008_s N_A_221_49#_M1001_d
+ N_A_221_49#_M1003_d N_A_221_49#_c_357_n N_A_221_49#_c_358_n
+ N_A_221_49#_c_359_n N_A_221_49#_c_370_n N_A_221_49#_c_360_n
+ N_A_221_49#_c_361_n N_A_221_49#_c_362_n PM_SKY130_FD_SC_LP__O221AI_1%A_221_49#
x_PM_SKY130_FD_SC_LP__O221AI_1%VGND N_VGND_M1006_d N_VGND_c_402_n VGND
+ N_VGND_c_403_n N_VGND_c_404_n N_VGND_c_405_n N_VGND_c_406_n
+ PM_SKY130_FD_SC_LP__O221AI_1%VGND
cc_1 VNB N_C1_M1002_g 0.0332231f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.655
cc_2 VNB N_C1_M1000_g 0.00154808f $X=-0.19 $Y=-0.245 $X2=0.675 $Y2=2.465
cc_3 VNB N_C1_c_61_n 0.00129844f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.46
cc_4 VNB N_C1_c_62_n 0.0683907f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.46
cc_5 VNB N_B1_M1008_g 0.0307002f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.655
cc_6 VNB N_B1_c_90_n 0.00529209f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.46
cc_7 VNB N_B1_c_91_n 0.0330459f $X=-0.19 $Y=-0.245 $X2=0.675 $Y2=1.625
cc_8 VNB N_B2_M1001_g 0.025264f $X=-0.19 $Y=-0.245 $X2=0.675 $Y2=2.465
cc_9 VNB N_B2_c_127_n 0.0217697f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.46
cc_10 VNB N_B2_c_128_n 0.00559372f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.46
cc_11 VNB N_A2_M1006_g 0.0243346f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.655
cc_12 VNB A2 0.0051285f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_13 VNB N_A2_c_166_n 0.0217149f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A1_M1003_g 0.0286513f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.655
cc_15 VNB N_A1_M1005_g 0.00176104f $X=-0.19 $Y=-0.245 $X2=0.675 $Y2=2.465
cc_16 VNB N_A1_c_207_n 0.045552f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.46
cc_17 VNB N_A1_c_208_n 0.012339f $X=-0.19 $Y=-0.245 $X2=0.675 $Y2=1.625
cc_18 VNB N_Y_c_229_n 0.00324534f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.46
cc_19 VNB Y 0.00711519f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_Y_c_231_n 0.00934659f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_Y_c_232_n 0.0284746f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_VPWR_c_288_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_114_47#_c_334_n 0.00976939f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_24 VNB N_A_114_47#_c_335_n 0.00513623f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.46
cc_25 VNB N_A_221_49#_c_357_n 0.00488388f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.46
cc_26 VNB N_A_221_49#_c_358_n 0.00373846f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.46
cc_27 VNB N_A_221_49#_c_359_n 0.00382096f $X=-0.19 $Y=-0.245 $X2=0.675 $Y2=1.625
cc_28 VNB N_A_221_49#_c_360_n 0.0138813f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_221_49#_c_361_n 0.0286004f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_221_49#_c_362_n 0.00889046f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_402_n 0.00319327f $X=-0.19 $Y=-0.245 $X2=0.675 $Y2=2.465
cc_32 VNB N_VGND_c_403_n 0.0635447f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_404_n 0.0156658f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_405_n 0.191922f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_406_n 0.00526561f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VPB N_C1_M1000_g 0.026905f $X=-0.19 $Y=1.655 $X2=0.675 $Y2=2.465
cc_37 VPB N_C1_c_61_n 0.0124971f $X=-0.19 $Y=1.655 $X2=0.29 $Y2=1.46
cc_38 VPB N_B1_M1007_g 0.0203979f $X=-0.19 $Y=1.655 $X2=0.675 $Y2=2.465
cc_39 VPB N_B1_c_90_n 0.00374106f $X=-0.19 $Y=1.655 $X2=0.29 $Y2=1.46
cc_40 VPB N_B1_c_91_n 0.0097125f $X=-0.19 $Y=1.655 $X2=0.675 $Y2=1.625
cc_41 VPB N_B2_M1009_g 0.0199048f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=0.655
cc_42 VPB N_B2_c_127_n 0.00623577f $X=-0.19 $Y=1.655 $X2=0.29 $Y2=1.46
cc_43 VPB N_B2_c_128_n 0.0052204f $X=-0.19 $Y=1.655 $X2=0.29 $Y2=1.46
cc_44 VPB N_A2_M1004_g 0.0201232f $X=-0.19 $Y=1.655 $X2=0.675 $Y2=2.465
cc_45 VPB A2 0.00225429f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_46 VPB N_A2_c_166_n 0.00948199f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_47 VPB N_A1_M1005_g 0.0245897f $X=-0.19 $Y=1.655 $X2=0.675 $Y2=2.465
cc_48 VPB N_A1_c_208_n 0.00679678f $X=-0.19 $Y=1.655 $X2=0.675 $Y2=1.625
cc_49 VPB N_Y_c_233_n 0.036317f $X=-0.19 $Y=1.655 $X2=0.29 $Y2=1.46
cc_50 VPB Y 0.00160851f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_51 VPB N_Y_c_235_n 0.00829097f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_52 VPB N_VPWR_c_289_n 0.00192478f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_53 VPB N_VPWR_c_290_n 0.0103398f $X=-0.19 $Y=1.655 $X2=0.29 $Y2=1.46
cc_54 VPB N_VPWR_c_291_n 0.0484246f $X=-0.19 $Y=1.655 $X2=0.29 $Y2=1.46
cc_55 VPB N_VPWR_c_292_n 0.0217403f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_56 VPB N_VPWR_c_293_n 0.0419248f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_57 VPB N_VPWR_c_294_n 0.0104351f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_58 VPB N_VPWR_c_288_n 0.0526623f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_59 N_C1_M1000_g N_B1_M1007_g 0.0114548f $X=0.675 $Y=2.465 $X2=0 $Y2=0
cc_60 N_C1_c_62_n N_B1_c_90_n 8.5988e-19 $X=0.495 $Y=1.46 $X2=0 $Y2=0
cc_61 N_C1_c_62_n N_B1_c_91_n 0.00942882f $X=0.495 $Y=1.46 $X2=0 $Y2=0
cc_62 N_C1_M1002_g N_Y_c_229_n 0.0188868f $X=0.495 $Y=0.655 $X2=0 $Y2=0
cc_63 N_C1_c_61_n N_Y_c_229_n 0.00590726f $X=0.29 $Y=1.46 $X2=0 $Y2=0
cc_64 N_C1_c_62_n N_Y_c_229_n 0.00284905f $X=0.495 $Y=1.46 $X2=0 $Y2=0
cc_65 N_C1_M1002_g Y 0.00873796f $X=0.495 $Y=0.655 $X2=0 $Y2=0
cc_66 N_C1_M1000_g Y 0.0149252f $X=0.675 $Y=2.465 $X2=0 $Y2=0
cc_67 N_C1_c_61_n Y 0.0316153f $X=0.29 $Y=1.46 $X2=0 $Y2=0
cc_68 N_C1_c_62_n Y 0.00783647f $X=0.495 $Y=1.46 $X2=0 $Y2=0
cc_69 N_C1_c_61_n N_Y_c_231_n 0.021435f $X=0.29 $Y=1.46 $X2=0 $Y2=0
cc_70 N_C1_c_62_n N_Y_c_231_n 0.00620474f $X=0.495 $Y=1.46 $X2=0 $Y2=0
cc_71 N_C1_M1000_g N_Y_c_235_n 0.0135644f $X=0.675 $Y=2.465 $X2=0 $Y2=0
cc_72 N_C1_c_61_n N_Y_c_235_n 0.0128386f $X=0.29 $Y=1.46 $X2=0 $Y2=0
cc_73 N_C1_c_62_n N_Y_c_235_n 0.00504195f $X=0.495 $Y=1.46 $X2=0 $Y2=0
cc_74 N_C1_M1000_g N_VPWR_c_289_n 0.0183024f $X=0.675 $Y=2.465 $X2=0 $Y2=0
cc_75 N_C1_M1000_g N_VPWR_c_292_n 0.00486043f $X=0.675 $Y=2.465 $X2=0 $Y2=0
cc_76 N_C1_M1000_g N_VPWR_c_288_n 0.00932201f $X=0.675 $Y=2.465 $X2=0 $Y2=0
cc_77 N_C1_M1002_g N_A_114_47#_c_335_n 0.00670331f $X=0.495 $Y=0.655 $X2=0 $Y2=0
cc_78 N_C1_c_62_n N_A_114_47#_c_335_n 3.73041e-19 $X=0.495 $Y=1.46 $X2=0 $Y2=0
cc_79 N_C1_M1002_g N_A_221_49#_c_357_n 0.00322073f $X=0.495 $Y=0.655 $X2=0 $Y2=0
cc_80 N_C1_M1002_g N_A_221_49#_c_359_n 9.95316e-19 $X=0.495 $Y=0.655 $X2=0 $Y2=0
cc_81 N_C1_M1002_g N_VGND_c_403_n 0.00547432f $X=0.495 $Y=0.655 $X2=0 $Y2=0
cc_82 N_C1_M1002_g N_VGND_c_405_n 0.0121265f $X=0.495 $Y=0.655 $X2=0 $Y2=0
cc_83 N_B1_M1007_g N_B2_M1009_g 0.0577034f $X=1.445 $Y=2.465 $X2=0 $Y2=0
cc_84 N_B1_M1008_g N_B2_M1001_g 0.0185175f $X=1.445 $Y=0.665 $X2=0 $Y2=0
cc_85 N_B1_c_90_n N_B2_c_127_n 3.06477e-19 $X=1.25 $Y=1.51 $X2=0 $Y2=0
cc_86 N_B1_c_91_n N_B2_c_127_n 0.0577034f $X=1.445 $Y=1.51 $X2=0 $Y2=0
cc_87 N_B1_c_90_n N_B2_c_128_n 0.0351587f $X=1.25 $Y=1.51 $X2=0 $Y2=0
cc_88 N_B1_c_91_n N_B2_c_128_n 0.00342916f $X=1.445 $Y=1.51 $X2=0 $Y2=0
cc_89 N_B1_M1008_g N_Y_c_229_n 7.09747e-19 $X=1.445 $Y=0.665 $X2=0 $Y2=0
cc_90 N_B1_M1007_g N_Y_c_249_n 0.0194762f $X=1.445 $Y=2.465 $X2=0 $Y2=0
cc_91 N_B1_c_90_n N_Y_c_249_n 0.0233653f $X=1.25 $Y=1.51 $X2=0 $Y2=0
cc_92 N_B1_c_91_n N_Y_c_249_n 0.00143225f $X=1.445 $Y=1.51 $X2=0 $Y2=0
cc_93 N_B1_M1008_g Y 0.00437288f $X=1.445 $Y=0.665 $X2=0 $Y2=0
cc_94 N_B1_M1007_g Y 0.00284616f $X=1.445 $Y=2.465 $X2=0 $Y2=0
cc_95 N_B1_c_90_n Y 0.0354896f $X=1.25 $Y=1.51 $X2=0 $Y2=0
cc_96 N_B1_c_91_n Y 0.00113614f $X=1.445 $Y=1.51 $X2=0 $Y2=0
cc_97 N_B1_M1007_g N_Y_c_235_n 3.87416e-19 $X=1.445 $Y=2.465 $X2=0 $Y2=0
cc_98 N_B1_M1007_g N_VPWR_c_289_n 0.0237928f $X=1.445 $Y=2.465 $X2=0 $Y2=0
cc_99 N_B1_M1007_g N_VPWR_c_293_n 0.00486043f $X=1.445 $Y=2.465 $X2=0 $Y2=0
cc_100 N_B1_M1007_g N_VPWR_c_288_n 0.00818711f $X=1.445 $Y=2.465 $X2=0 $Y2=0
cc_101 N_B1_M1008_g N_A_114_47#_c_334_n 0.0114689f $X=1.445 $Y=0.665 $X2=0 $Y2=0
cc_102 N_B1_M1008_g N_A_114_47#_c_335_n 0.00248909f $X=1.445 $Y=0.665 $X2=0
+ $Y2=0
cc_103 N_B1_M1008_g N_A_221_49#_c_357_n 0.00637118f $X=1.445 $Y=0.665 $X2=0
+ $Y2=0
cc_104 N_B1_M1008_g N_A_221_49#_c_358_n 0.0148984f $X=1.445 $Y=0.665 $X2=0 $Y2=0
cc_105 N_B1_M1008_g N_A_221_49#_c_359_n 0.004061f $X=1.445 $Y=0.665 $X2=0 $Y2=0
cc_106 N_B1_c_90_n N_A_221_49#_c_359_n 0.0264163f $X=1.25 $Y=1.51 $X2=0 $Y2=0
cc_107 N_B1_c_91_n N_A_221_49#_c_359_n 0.00221413f $X=1.445 $Y=1.51 $X2=0 $Y2=0
cc_108 N_B1_M1008_g N_A_221_49#_c_370_n 4.18786e-19 $X=1.445 $Y=0.665 $X2=0
+ $Y2=0
cc_109 N_B1_M1008_g N_VGND_c_403_n 0.00351226f $X=1.445 $Y=0.665 $X2=0 $Y2=0
cc_110 N_B1_M1008_g N_VGND_c_405_n 0.00687017f $X=1.445 $Y=0.665 $X2=0 $Y2=0
cc_111 N_B2_M1001_g N_A2_M1006_g 0.0243706f $X=1.985 $Y=0.665 $X2=0 $Y2=0
cc_112 N_B2_M1009_g N_A2_M1004_g 0.0219509f $X=1.805 $Y=2.465 $X2=0 $Y2=0
cc_113 N_B2_c_128_n N_A2_M1004_g 8.33509e-19 $X=1.895 $Y=1.51 $X2=0 $Y2=0
cc_114 N_B2_M1009_g A2 0.00120158f $X=1.805 $Y=2.465 $X2=0 $Y2=0
cc_115 N_B2_c_127_n A2 4.13162e-19 $X=1.895 $Y=1.51 $X2=0 $Y2=0
cc_116 N_B2_c_128_n A2 0.0262482f $X=1.895 $Y=1.51 $X2=0 $Y2=0
cc_117 N_B2_c_127_n N_A2_c_166_n 0.0214266f $X=1.895 $Y=1.51 $X2=0 $Y2=0
cc_118 N_B2_c_128_n N_A2_c_166_n 4.12637e-19 $X=1.895 $Y=1.51 $X2=0 $Y2=0
cc_119 N_B2_M1009_g N_Y_c_249_n 0.0155045f $X=1.805 $Y=2.465 $X2=0 $Y2=0
cc_120 N_B2_c_127_n N_Y_c_249_n 4.86217e-19 $X=1.895 $Y=1.51 $X2=0 $Y2=0
cc_121 N_B2_c_128_n N_Y_c_249_n 0.0284779f $X=1.895 $Y=1.51 $X2=0 $Y2=0
cc_122 N_B2_c_127_n N_Y_c_260_n 4.26566e-19 $X=1.895 $Y=1.51 $X2=0 $Y2=0
cc_123 N_B2_c_128_n N_Y_c_260_n 0.00605827f $X=1.895 $Y=1.51 $X2=0 $Y2=0
cc_124 N_B2_M1009_g N_Y_c_262_n 0.0168149f $X=1.805 $Y=2.465 $X2=0 $Y2=0
cc_125 N_B2_M1009_g N_VPWR_c_289_n 0.00357776f $X=1.805 $Y=2.465 $X2=0 $Y2=0
cc_126 N_B2_M1009_g N_VPWR_c_293_n 0.00585385f $X=1.805 $Y=2.465 $X2=0 $Y2=0
cc_127 N_B2_M1009_g N_VPWR_c_288_n 0.0114297f $X=1.805 $Y=2.465 $X2=0 $Y2=0
cc_128 N_B2_M1001_g N_A_221_49#_c_357_n 3.82796e-19 $X=1.985 $Y=0.665 $X2=0
+ $Y2=0
cc_129 N_B2_M1001_g N_A_221_49#_c_358_n 0.013103f $X=1.985 $Y=0.665 $X2=0 $Y2=0
cc_130 N_B2_c_127_n N_A_221_49#_c_358_n 0.00463193f $X=1.895 $Y=1.51 $X2=0 $Y2=0
cc_131 N_B2_c_128_n N_A_221_49#_c_358_n 0.0391321f $X=1.895 $Y=1.51 $X2=0 $Y2=0
cc_132 N_B2_M1001_g N_A_221_49#_c_370_n 0.00994111f $X=1.985 $Y=0.665 $X2=0
+ $Y2=0
cc_133 N_B2_M1001_g N_A_221_49#_c_362_n 0.00134433f $X=1.985 $Y=0.665 $X2=0
+ $Y2=0
cc_134 N_B2_c_128_n N_A_221_49#_c_362_n 8.13827e-19 $X=1.895 $Y=1.51 $X2=0 $Y2=0
cc_135 N_B2_M1001_g N_VGND_c_403_n 0.00561712f $X=1.985 $Y=0.665 $X2=0 $Y2=0
cc_136 N_B2_M1001_g N_VGND_c_405_n 0.010775f $X=1.985 $Y=0.665 $X2=0 $Y2=0
cc_137 N_A2_M1006_g N_A1_M1003_g 0.023077f $X=2.415 $Y=0.665 $X2=0 $Y2=0
cc_138 N_A2_M1004_g N_A1_M1005_g 0.0561821f $X=2.525 $Y=2.465 $X2=0 $Y2=0
cc_139 A2 N_A1_M1005_g 0.0112765f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_140 A2 N_A1_c_207_n 0.00235445f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_141 N_A2_c_166_n N_A1_c_207_n 0.0561821f $X=2.435 $Y=1.51 $X2=0 $Y2=0
cc_142 A2 N_A1_c_208_n 0.0328353f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_143 N_A2_c_166_n N_A1_c_208_n 2.71878e-19 $X=2.435 $Y=1.51 $X2=0 $Y2=0
cc_144 N_A2_M1004_g N_Y_c_260_n 0.001682f $X=2.525 $Y=2.465 $X2=0 $Y2=0
cc_145 A2 N_Y_c_260_n 0.0166061f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_146 N_A2_c_166_n N_Y_c_260_n 0.00109807f $X=2.435 $Y=1.51 $X2=0 $Y2=0
cc_147 N_A2_M1004_g N_Y_c_262_n 0.0095686f $X=2.525 $Y=2.465 $X2=0 $Y2=0
cc_148 A2 N_Y_c_262_n 0.0637588f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_149 N_A2_M1004_g N_VPWR_c_291_n 0.00242923f $X=2.525 $Y=2.465 $X2=0 $Y2=0
cc_150 A2 N_VPWR_c_291_n 0.0696263f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_151 N_A2_M1004_g N_VPWR_c_293_n 0.0043655f $X=2.525 $Y=2.465 $X2=0 $Y2=0
cc_152 A2 N_VPWR_c_293_n 0.00849121f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_153 N_A2_M1004_g N_VPWR_c_288_n 0.00744729f $X=2.525 $Y=2.465 $X2=0 $Y2=0
cc_154 A2 N_VPWR_c_288_n 0.00833565f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_155 A2 A_520_367# 0.0110648f $X=2.555 $Y=1.58 $X2=-0.19 $Y2=-0.245
cc_156 N_A2_M1006_g N_A_221_49#_c_360_n 0.0142207f $X=2.415 $Y=0.665 $X2=0 $Y2=0
cc_157 A2 N_A_221_49#_c_360_n 0.0307724f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_158 N_A2_c_166_n N_A_221_49#_c_360_n 0.00323377f $X=2.435 $Y=1.51 $X2=0 $Y2=0
cc_159 A2 N_A_221_49#_c_362_n 0.00463833f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_160 N_A2_c_166_n N_A_221_49#_c_362_n 0.00128126f $X=2.435 $Y=1.51 $X2=0 $Y2=0
cc_161 N_A2_M1006_g N_VGND_c_402_n 0.00317214f $X=2.415 $Y=0.665 $X2=0 $Y2=0
cc_162 N_A2_M1006_g N_VGND_c_403_n 0.00575161f $X=2.415 $Y=0.665 $X2=0 $Y2=0
cc_163 N_A2_M1006_g N_VGND_c_405_n 0.0106661f $X=2.415 $Y=0.665 $X2=0 $Y2=0
cc_164 N_A1_M1005_g N_VPWR_c_291_n 0.0230926f $X=2.885 $Y=2.465 $X2=0 $Y2=0
cc_165 N_A1_c_207_n N_VPWR_c_291_n 0.00146498f $X=3.07 $Y=1.46 $X2=0 $Y2=0
cc_166 N_A1_c_208_n N_VPWR_c_291_n 0.0262905f $X=3.07 $Y=1.46 $X2=0 $Y2=0
cc_167 N_A1_M1005_g N_VPWR_c_293_n 0.00486043f $X=2.885 $Y=2.465 $X2=0 $Y2=0
cc_168 N_A1_M1005_g N_VPWR_c_288_n 0.00818711f $X=2.885 $Y=2.465 $X2=0 $Y2=0
cc_169 N_A1_M1003_g N_A_221_49#_c_360_n 0.0174735f $X=2.885 $Y=0.665 $X2=0 $Y2=0
cc_170 N_A1_c_207_n N_A_221_49#_c_360_n 0.00676472f $X=3.07 $Y=1.46 $X2=0 $Y2=0
cc_171 N_A1_c_208_n N_A_221_49#_c_360_n 0.0299192f $X=3.07 $Y=1.46 $X2=0 $Y2=0
cc_172 N_A1_M1003_g N_VGND_c_402_n 0.0108377f $X=2.885 $Y=0.665 $X2=0 $Y2=0
cc_173 N_A1_M1003_g N_VGND_c_404_n 0.00515898f $X=2.885 $Y=0.665 $X2=0 $Y2=0
cc_174 N_A1_M1003_g N_VGND_c_405_n 0.00980941f $X=2.885 $Y=0.665 $X2=0 $Y2=0
cc_175 N_Y_c_249_n N_VPWR_M1000_d 0.0157325f $X=1.99 $Y=2.035 $X2=-0.19
+ $Y2=-0.245
cc_176 Y N_VPWR_M1000_d 0.00174802f $X=0.635 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_177 N_Y_c_235_n N_VPWR_M1000_d 0.00138445f $X=0.885 $Y=2.025 $X2=-0.19
+ $Y2=-0.245
cc_178 N_Y_c_262_n N_VPWR_c_289_n 0.0238926f $X=2.155 $Y=2.48 $X2=0 $Y2=0
cc_179 N_Y_c_235_n N_VPWR_c_289_n 0.044728f $X=0.885 $Y=2.025 $X2=0 $Y2=0
cc_180 N_Y_c_262_n N_VPWR_c_291_n 0.00323087f $X=2.155 $Y=2.48 $X2=0 $Y2=0
cc_181 N_Y_c_233_n N_VPWR_c_292_n 0.0178111f $X=0.46 $Y=2.48 $X2=0 $Y2=0
cc_182 N_Y_c_262_n N_VPWR_c_293_n 0.0230625f $X=2.155 $Y=2.48 $X2=0 $Y2=0
cc_183 N_Y_M1000_s N_VPWR_c_288_n 0.00371702f $X=0.335 $Y=1.835 $X2=0 $Y2=0
cc_184 N_Y_M1009_d N_VPWR_c_288_n 0.0130729f $X=1.88 $Y=1.835 $X2=0 $Y2=0
cc_185 N_Y_c_233_n N_VPWR_c_288_n 0.0100304f $X=0.46 $Y=2.48 $X2=0 $Y2=0
cc_186 N_Y_c_262_n N_VPWR_c_288_n 0.0127519f $X=2.155 $Y=2.48 $X2=0 $Y2=0
cc_187 N_Y_c_249_n A_304_367# 0.00469833f $X=1.99 $Y=2.035 $X2=-0.19 $Y2=-0.245
cc_188 N_Y_c_229_n N_A_114_47#_M1002_d 0.00263111f $X=0.625 $Y=1.09 $X2=-0.19
+ $Y2=-0.245
cc_189 N_Y_c_229_n N_A_114_47#_c_334_n 3.43077e-19 $X=0.625 $Y=1.09 $X2=0 $Y2=0
cc_190 N_Y_c_229_n N_A_114_47#_c_335_n 0.023909f $X=0.625 $Y=1.09 $X2=0 $Y2=0
cc_191 N_Y_c_229_n N_A_221_49#_c_359_n 0.0152916f $X=0.625 $Y=1.09 $X2=0 $Y2=0
cc_192 N_Y_c_232_n N_VGND_c_403_n 0.0178111f $X=0.28 $Y=0.42 $X2=0 $Y2=0
cc_193 N_Y_M1002_s N_VGND_c_405_n 0.00371702f $X=0.155 $Y=0.235 $X2=0 $Y2=0
cc_194 N_Y_c_232_n N_VGND_c_405_n 0.0100304f $X=0.28 $Y=0.42 $X2=0 $Y2=0
cc_195 N_VPWR_c_288_n A_304_367# 0.00899413f $X=3.12 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_196 N_VPWR_c_288_n A_520_367# 0.00439517f $X=3.12 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_197 N_A_114_47#_c_334_n N_A_221_49#_M1008_s 0.00495471f $X=1.55 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_198 N_A_114_47#_c_334_n N_A_221_49#_c_357_n 0.0192796f $X=1.55 $Y=0.34 $X2=0
+ $Y2=0
cc_199 N_A_114_47#_c_335_n N_A_221_49#_c_357_n 0.0184158f $X=0.71 $Y=0.38 $X2=0
+ $Y2=0
cc_200 N_A_114_47#_M1008_d N_A_221_49#_c_358_n 0.00315828f $X=1.52 $Y=0.245
+ $X2=0 $Y2=0
cc_201 N_A_114_47#_c_334_n N_A_221_49#_c_358_n 0.00349462f $X=1.55 $Y=0.34 $X2=0
+ $Y2=0
cc_202 N_A_114_47#_c_348_p N_A_221_49#_c_358_n 0.0212613f $X=1.715 $Y=0.37 $X2=0
+ $Y2=0
cc_203 N_A_114_47#_c_334_n N_VGND_c_403_n 0.0402398f $X=1.55 $Y=0.34 $X2=0 $Y2=0
cc_204 N_A_114_47#_c_335_n N_VGND_c_403_n 0.0209663f $X=0.71 $Y=0.38 $X2=0 $Y2=0
cc_205 N_A_114_47#_c_348_p N_VGND_c_403_n 0.0210494f $X=1.715 $Y=0.37 $X2=0
+ $Y2=0
cc_206 N_A_114_47#_M1002_d N_VGND_c_405_n 0.00215158f $X=0.57 $Y=0.235 $X2=0
+ $Y2=0
cc_207 N_A_114_47#_M1008_d N_VGND_c_405_n 0.00412903f $X=1.52 $Y=0.245 $X2=0
+ $Y2=0
cc_208 N_A_114_47#_c_334_n N_VGND_c_405_n 0.0246172f $X=1.55 $Y=0.34 $X2=0 $Y2=0
cc_209 N_A_114_47#_c_335_n N_VGND_c_405_n 0.0125896f $X=0.71 $Y=0.38 $X2=0 $Y2=0
cc_210 N_A_114_47#_c_348_p N_VGND_c_405_n 0.0127654f $X=1.715 $Y=0.37 $X2=0
+ $Y2=0
cc_211 N_A_221_49#_c_360_n N_VGND_M1006_d 0.00218982f $X=2.995 $Y=1.09 $X2=-0.19
+ $Y2=-0.245
cc_212 N_A_221_49#_c_360_n N_VGND_c_402_n 0.0177842f $X=2.995 $Y=1.09 $X2=0
+ $Y2=0
cc_213 N_A_221_49#_c_370_n N_VGND_c_403_n 0.0157299f $X=2.2 $Y=0.42 $X2=0 $Y2=0
cc_214 N_A_221_49#_c_361_n N_VGND_c_404_n 0.0181659f $X=3.1 $Y=0.42 $X2=0 $Y2=0
cc_215 N_A_221_49#_M1008_s N_VGND_c_405_n 0.00213122f $X=1.105 $Y=0.245 $X2=0
+ $Y2=0
cc_216 N_A_221_49#_M1001_d N_VGND_c_405_n 0.0027574f $X=2.06 $Y=0.245 $X2=0
+ $Y2=0
cc_217 N_A_221_49#_M1003_d N_VGND_c_405_n 0.00334057f $X=2.96 $Y=0.245 $X2=0
+ $Y2=0
cc_218 N_A_221_49#_c_370_n N_VGND_c_405_n 0.0104992f $X=2.2 $Y=0.42 $X2=0 $Y2=0
cc_219 N_A_221_49#_c_361_n N_VGND_c_405_n 0.0104192f $X=3.1 $Y=0.42 $X2=0 $Y2=0
