* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__a2bb2o_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
X0 a_742_367# A2_N a_436_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X1 VGND A1_N a_436_21# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X2 VGND a_200_47# X VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X3 VGND B1 a_114_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X4 X a_200_47# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X5 VPWR a_200_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X6 a_436_21# A1_N VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X7 a_436_21# A2_N a_742_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X8 VGND a_200_47# X VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X9 a_114_47# B2 a_200_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X10 VGND a_436_21# a_200_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X11 X a_200_47# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X12 a_200_47# a_436_21# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X13 X a_200_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X14 VPWR A1_N a_742_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X15 a_742_367# A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X16 a_27_367# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X17 a_27_367# a_436_21# a_200_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X18 VPWR B1 a_27_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X19 VPWR B2 a_27_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X20 a_27_367# B2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X21 a_200_47# B2 a_114_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X22 VPWR a_200_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X23 X a_200_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X24 a_114_47# B1 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X25 a_436_21# A2_N VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X26 a_200_47# a_436_21# a_27_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X27 VGND A2_N a_436_21# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
.ends
