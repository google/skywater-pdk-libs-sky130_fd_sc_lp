* File: sky130_fd_sc_lp__o21ai_2.spice
* Created: Fri Aug 28 11:04:48 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__o21ai_2.pex.spice"
.subckt sky130_fd_sc_lp__o21ai_2  VNB VPB A1 A2 B1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B1	B1
* A2	A2
* A1	A1
* VPB	VPB
* VNB	VNB
MM1005 N_VGND_M1005_d N_A1_M1005_g N_A_30_47#_M1005_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75002.5 A=0.126 P=1.98 MULT=1
MM1001 N_VGND_M1005_d N_A2_M1001_g N_A_30_47#_M1001_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75002.1 A=0.126 P=1.98 MULT=1
MM1009 N_VGND_M1009_d N_A2_M1009_g N_A_30_47#_M1001_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1995 AS=0.1176 PD=1.315 PS=1.12 NRD=19.284 NRS=0 M=1 R=5.6 SA=75001.1
+ SB=75001.7 A=0.126 P=1.98 MULT=1
MM1010 N_VGND_M1009_d N_A1_M1010_g N_A_30_47#_M1010_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1995 AS=0.1176 PD=1.315 PS=1.12 NRD=8.568 NRS=0 M=1 R=5.6 SA=75001.7
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1004 N_Y_M1004_d N_B1_M1004_g N_A_30_47#_M1010_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002.1
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1008 N_Y_M1004_d N_B1_M1008_g N_A_30_47#_M1008_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75002.5
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1003 N_VPWR_M1003_d N_A1_M1003_g N_A_113_367#_M1003_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75002.5 A=0.189 P=2.82 MULT=1
MM1002 N_Y_M1002_d N_A2_M1002_g N_A_113_367#_M1003_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75002.1 A=0.189 P=2.82 MULT=1
MM1011 N_Y_M1002_d N_A2_M1011_g N_A_113_367#_M1011_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.27405 PD=1.54 PS=1.695 NRD=0 NRS=11.7215 M=1 R=8.4 SA=75001.1
+ SB=75001.7 A=0.189 P=2.82 MULT=1
MM1007 N_VPWR_M1007_d N_A1_M1007_g N_A_113_367#_M1011_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.2016 AS=0.27405 PD=1.58 PS=1.695 NRD=2.3443 NRS=12.4898 M=1 R=8.4
+ SA=75001.6 SB=75001.1 A=0.189 P=2.82 MULT=1
MM1000 N_Y_M1000_d N_B1_M1000_g N_VPWR_M1007_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.2016 PD=1.54 PS=1.58 NRD=0 NRS=3.9006 M=1 R=8.4 SA=75002.1
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1006 N_Y_M1000_d N_B1_M1006_g N_VPWR_M1006_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75002.5
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX12_noxref VNB VPB NWDIODE A=6.9751 P=11.21
*
.include "sky130_fd_sc_lp__o21ai_2.pxi.spice"
*
.ends
*
*
