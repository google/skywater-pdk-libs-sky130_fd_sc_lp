* File: sky130_fd_sc_lp__dlrtp_2.pex.spice
* Created: Wed Sep  2 09:47:24 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__DLRTP_2%D 3 5 8 10 11 12 13 14 15 23 25 42
c44 12 0 6.23206e-20 $X=0.635 $Y=0.84
r45 23 25 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=0.652 $Y=0.965
+ $X2=0.652 $Y2=0.8
r46 14 15 14.2135 $w=2.98e-07 $l=3.7e-07 $layer=LI1_cond $X=0.73 $Y=1.665
+ $X2=0.73 $Y2=2.035
r47 13 14 14.2135 $w=2.98e-07 $l=3.7e-07 $layer=LI1_cond $X=0.73 $Y=1.295
+ $X2=0.73 $Y2=1.665
r48 12 42 1.53659 $w=2.98e-07 $l=4e-08 $layer=LI1_cond $X=0.73 $Y=0.965 $X2=0.73
+ $Y2=0.925
r49 12 42 0.88354 $w=2.98e-07 $l=2.3e-08 $layer=LI1_cond $X=0.73 $Y=0.902
+ $X2=0.73 $Y2=0.925
r50 12 40 4.08822 $w=2.98e-07 $l=8.7e-08 $layer=LI1_cond $X=0.73 $Y=0.902
+ $X2=0.73 $Y2=0.815
r51 12 13 12.6769 $w=2.98e-07 $l=3.3e-07 $layer=LI1_cond $X=0.73 $Y=0.965
+ $X2=0.73 $Y2=1.295
r52 12 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.675
+ $Y=0.965 $X2=0.675 $Y2=0.965
r53 11 40 13.3171 $w=2.23e-07 $l=2.6e-07 $layer=LI1_cond $X=0.692 $Y=0.555
+ $X2=0.692 $Y2=0.815
r54 8 10 628.138 $w=1.5e-07 $l=1.225e-06 $layer=POLY_cond $X=0.54 $Y=2.695
+ $X2=0.54 $Y2=1.47
r55 5 10 48.4185 $w=3.75e-07 $l=1.87e-07 $layer=POLY_cond $X=0.652 $Y=1.283
+ $X2=0.652 $Y2=1.47
r56 4 23 3.26277 $w=3.75e-07 $l=2.2e-08 $layer=POLY_cond $X=0.652 $Y=0.987
+ $X2=0.652 $Y2=0.965
r57 4 5 43.8991 $w=3.75e-07 $l=2.96e-07 $layer=POLY_cond $X=0.652 $Y=0.987
+ $X2=0.652 $Y2=1.283
r58 3 25 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.54 $Y=0.48 $X2=0.54
+ $Y2=0.8
.ends

.subckt PM_SKY130_FD_SC_LP__DLRTP_2%GATE 3 7 11 12 13 14 15 16 22
c54 7 0 6.23206e-20 $X=1.295 $Y=0.48
r55 15 16 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=1.175 $Y=1.665
+ $X2=1.175 $Y2=2.035
r56 14 15 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=1.175 $Y=1.295
+ $X2=1.175 $Y2=1.665
r57 13 14 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=1.175 $Y=0.925
+ $X2=1.175 $Y2=1.295
r58 13 22 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.215
+ $Y=1.005 $X2=1.215 $Y2=1.005
r59 11 22 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.215 $Y=1.345
+ $X2=1.215 $Y2=1.005
r60 11 12 39.6269 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.215 $Y=1.345
+ $X2=1.215 $Y2=1.51
r61 10 22 44.4756 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.215 $Y=0.84
+ $X2=1.215 $Y2=1.005
r62 7 10 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=1.295 $Y=0.48
+ $X2=1.295 $Y2=0.84
r63 3 12 607.628 $w=1.5e-07 $l=1.185e-06 $layer=POLY_cond $X=1.18 $Y=2.695
+ $X2=1.18 $Y2=1.51
.ends

.subckt PM_SKY130_FD_SC_LP__DLRTP_2%A_251_475# 1 2 9 13 15 17 20 22 23 26 30 33
+ 36 37 40 43 44 46 50 53 56 60 61 65 71
c154 46 0 1.63114e-19 $X=3.675 $Y=1.125
c155 43 0 1.934e-19 $X=3.59 $Y=0.79
c156 26 0 9.36306e-20 $X=3.695 $Y=0.445
c157 9 0 4.84857e-20 $X=2.18 $Y=2.14
r158 60 61 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.785
+ $Y=1.29 $X2=3.785 $Y2=1.29
r159 57 60 4.87572 $w=2.58e-07 $l=1.1e-07 $layer=LI1_cond $X=3.675 $Y=1.255
+ $X2=3.785 $Y2=1.255
r160 55 56 79.9198 $w=1.68e-07 $l=1.225e-06 $layer=LI1_cond $X=1.565 $Y=0.66
+ $X2=1.565 $Y2=1.885
r161 53 55 9.16686 $w=2.23e-07 $l=1.65e-07 $layer=LI1_cond $X=1.537 $Y=0.495
+ $X2=1.537 $Y2=0.66
r162 48 50 4.86587 $w=3.58e-07 $l=1.52e-07 $layer=LI1_cond $X=1.445 $Y=2.535
+ $X2=1.597 $Y2=2.535
r163 46 57 3.22376 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.675 $Y=1.125
+ $X2=3.675 $Y2=1.255
r164 45 46 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=3.675 $Y=0.875
+ $X2=3.675 $Y2=1.125
r165 43 45 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.59 $Y=0.79
+ $X2=3.675 $Y2=0.875
r166 43 44 70.4599 $w=1.68e-07 $l=1.08e-06 $layer=LI1_cond $X=3.59 $Y=0.79
+ $X2=2.51 $Y2=0.79
r167 41 71 1.5971 $w=6.7e-07 $l=2e-08 $layer=POLY_cond $X=2.345 $Y=1.1 $X2=2.365
+ $Y2=1.1
r168 41 68 49.9095 $w=6.7e-07 $l=6.25e-07 $layer=POLY_cond $X=2.345 $Y=1.1
+ $X2=1.72 $Y2=1.1
r169 40 41 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.345
+ $Y=0.93 $X2=2.345 $Y2=0.93
r170 38 44 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.345 $Y=0.875
+ $X2=2.51 $Y2=0.79
r171 38 40 1.92074 $w=3.28e-07 $l=5.5e-08 $layer=LI1_cond $X=2.345 $Y=0.875
+ $X2=2.345 $Y2=0.93
r172 37 66 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=1.63 $Y=2.05 $X2=1.63
+ $Y2=2.14
r173 37 65 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.63 $Y=2.05
+ $X2=1.63 $Y2=1.885
r174 36 37 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.63
+ $Y=2.05 $X2=1.63 $Y2=2.05
r175 34 50 3.25024 $w=2.35e-07 $l=1.8e-07 $layer=LI1_cond $X=1.597 $Y=2.355
+ $X2=1.597 $Y2=2.535
r176 34 36 14.9572 $w=2.33e-07 $l=3.05e-07 $layer=LI1_cond $X=1.597 $Y=2.355
+ $X2=1.597 $Y2=2.05
r177 33 56 6.63891 $w=2.33e-07 $l=1.17e-07 $layer=LI1_cond $X=1.597 $Y=2.002
+ $X2=1.597 $Y2=1.885
r178 33 36 2.35393 $w=2.33e-07 $l=4.8e-08 $layer=LI1_cond $X=1.597 $Y=2.002
+ $X2=1.597 $Y2=2.05
r179 30 61 39.3438 $w=3.3e-07 $l=2.25e-07 $layer=POLY_cond $X=3.785 $Y=1.515
+ $X2=3.785 $Y2=1.29
r180 29 61 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.785 $Y=1.125
+ $X2=3.785 $Y2=1.29
r181 26 29 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=3.695 $Y=0.445
+ $X2=3.695 $Y2=1.125
r182 22 30 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=3.62 $Y=1.59
+ $X2=3.785 $Y2=1.515
r183 22 23 105.117 $w=1.5e-07 $l=2.05e-07 $layer=POLY_cond $X=3.62 $Y=1.59
+ $X2=3.415 $Y2=1.59
r184 18 23 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.34 $Y=1.665
+ $X2=3.415 $Y2=1.59
r185 18 20 538.404 $w=1.5e-07 $l=1.05e-06 $layer=POLY_cond $X=3.34 $Y=1.665
+ $X2=3.34 $Y2=2.715
r186 15 71 38.9565 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=2.365 $Y=0.765
+ $X2=2.365 $Y2=1.1
r187 15 17 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.365 $Y=0.765
+ $X2=2.365 $Y2=0.445
r188 11 13 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=2.255 $Y=2.215
+ $X2=2.255 $Y2=2.715
r189 10 66 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.795 $Y=2.14
+ $X2=1.63 $Y2=2.14
r190 9 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.18 $Y=2.14
+ $X2=2.255 $Y2=2.215
r191 9 10 197.415 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=2.18 $Y=2.14
+ $X2=1.795 $Y2=2.14
r192 7 68 38.9565 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=1.72 $Y=1.435
+ $X2=1.72 $Y2=1.1
r193 7 65 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=1.72 $Y=1.435
+ $X2=1.72 $Y2=1.885
r194 2 48 600 $w=1.7e-07 $l=2.63344e-07 $layer=licon1_PDIFF $count=1 $X=1.255
+ $Y=2.375 $X2=1.445 $Y2=2.55
r195 1 53 182 $w=1.7e-07 $l=2.94321e-07 $layer=licon1_NDIFF $count=1 $X=1.37
+ $Y=0.27 $X2=1.53 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__DLRTP_2%A_40_54# 1 2 9 13 17 21 24 25 26 28 30 34 38
c90 9 0 1.17851e-19 $X=2.795 $Y=0.445
r91 35 38 16.3698 $w=2.65e-07 $l=9e-08 $layer=POLY_cond $X=2.705 $Y=2.06
+ $X2=2.795 $Y2=2.06
r92 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.705
+ $Y=2.06 $X2=2.705 $Y2=2.06
r93 31 34 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=2.39 $Y=2.06
+ $X2=2.705 $Y2=2.06
r94 27 31 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.39 $Y=2.225
+ $X2=2.39 $Y2=2.06
r95 27 28 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=2.39 $Y=2.225
+ $X2=2.39 $Y2=2.885
r96 25 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.305 $Y=2.97
+ $X2=2.39 $Y2=2.885
r97 25 26 72.7433 $w=1.68e-07 $l=1.115e-06 $layer=LI1_cond $X=2.305 $Y=2.97
+ $X2=1.19 $Y2=2.97
r98 24 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.105 $Y=2.885
+ $X2=1.19 $Y2=2.97
r99 23 24 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=1.105 $Y=2.525
+ $X2=1.105 $Y2=2.885
r100 22 30 2.90867 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=0.43 $Y=2.44
+ $X2=0.295 $Y2=2.44
r101 21 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.02 $Y=2.44
+ $X2=1.105 $Y2=2.525
r102 21 22 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=1.02 $Y=2.44
+ $X2=0.43 $Y2=2.44
r103 15 30 3.58051 $w=2.6e-07 $l=8.9861e-08 $layer=LI1_cond $X=0.285 $Y=2.355
+ $X2=0.295 $Y2=2.44
r104 15 17 86.4332 $w=2.48e-07 $l=1.875e-06 $layer=LI1_cond $X=0.285 $Y=2.355
+ $X2=0.285 $Y2=0.48
r105 11 38 33.6491 $w=2.65e-07 $l=2.5446e-07 $layer=POLY_cond $X=2.98 $Y=2.225
+ $X2=2.795 $Y2=2.06
r106 11 13 251.255 $w=1.5e-07 $l=4.9e-07 $layer=POLY_cond $X=2.98 $Y=2.225
+ $X2=2.98 $Y2=2.715
r107 7 38 16.0701 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.795 $Y=1.895
+ $X2=2.795 $Y2=2.06
r108 7 9 743.511 $w=1.5e-07 $l=1.45e-06 $layer=POLY_cond $X=2.795 $Y=1.895
+ $X2=2.795 $Y2=0.445
r109 2 30 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.2
+ $Y=2.375 $X2=0.325 $Y2=2.52
r110 1 17 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.2
+ $Y=0.27 $X2=0.325 $Y2=0.48
.ends

.subckt PM_SKY130_FD_SC_LP__DLRTP_2%A_383_479# 1 2 9 13 16 19 21 24 26 27 28 30
+ 34 36 40 41 43 46 48
c135 41 0 1.80031e-19 $X=3.245 $Y=1.14
c136 40 0 9.36306e-20 $X=3.245 $Y=1.14
c137 26 0 4.84857e-20 $X=3.09 $Y=2.825
r138 46 55 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.79 $Y=2.07
+ $X2=3.79 $Y2=2.235
r139 45 48 6.80989 $w=3.28e-07 $l=1.95e-07 $layer=LI1_cond $X=3.79 $Y=2.07
+ $X2=3.985 $Y2=2.07
r140 45 46 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.79
+ $Y=2.07 $X2=3.79 $Y2=2.07
r141 41 51 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.245 $Y=1.14
+ $X2=3.245 $Y2=0.975
r142 40 41 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.245
+ $Y=1.14 $X2=3.245 $Y2=1.14
r143 37 40 6.87033 $w=2.58e-07 $l=1.55e-07 $layer=LI1_cond $X=3.09 $Y=1.175
+ $X2=3.245 $Y2=1.175
r144 31 34 8.84912 $w=2.78e-07 $l=2.15e-07 $layer=LI1_cond $X=1.915 $Y=0.395
+ $X2=2.13 $Y2=0.395
r145 29 48 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.985 $Y=2.235
+ $X2=3.985 $Y2=2.07
r146 29 30 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=3.985 $Y=2.235
+ $X2=3.985 $Y2=2.825
r147 27 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.9 $Y=2.91
+ $X2=3.985 $Y2=2.825
r148 27 28 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=3.9 $Y=2.91
+ $X2=3.175 $Y2=2.91
r149 26 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.09 $Y=2.825
+ $X2=3.175 $Y2=2.91
r150 25 43 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.09 $Y=1.705
+ $X2=3.09 $Y2=1.62
r151 25 26 73.0695 $w=1.68e-07 $l=1.12e-06 $layer=LI1_cond $X=3.09 $Y=1.705
+ $X2=3.09 $Y2=2.825
r152 24 43 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.09 $Y=1.535
+ $X2=3.09 $Y2=1.62
r153 23 37 3.22376 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.09 $Y=1.305
+ $X2=3.09 $Y2=1.175
r154 23 24 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=3.09 $Y=1.305
+ $X2=3.09 $Y2=1.535
r155 22 36 2.28545 $w=1.7e-07 $l=1.58e-07 $layer=LI1_cond $X=2.135 $Y=1.62
+ $X2=1.977 $Y2=1.62
r156 21 43 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.005 $Y=1.62
+ $X2=3.09 $Y2=1.62
r157 21 22 56.7594 $w=1.68e-07 $l=8.7e-07 $layer=LI1_cond $X=3.005 $Y=1.62
+ $X2=2.135 $Y2=1.62
r158 17 36 4.14756 $w=2.2e-07 $l=1.0015e-07 $layer=LI1_cond $X=2.01 $Y=1.705
+ $X2=1.977 $Y2=1.62
r159 17 19 38.9526 $w=2.48e-07 $l=8.45e-07 $layer=LI1_cond $X=2.01 $Y=1.705
+ $X2=2.01 $Y2=2.55
r160 16 36 4.14756 $w=2.2e-07 $l=1.11781e-07 $layer=LI1_cond $X=1.915 $Y=1.535
+ $X2=1.977 $Y2=1.62
r161 15 31 3.00742 $w=1.9e-07 $l=1.4e-07 $layer=LI1_cond $X=1.915 $Y=0.535
+ $X2=1.915 $Y2=0.395
r162 15 16 58.3732 $w=1.88e-07 $l=1e-06 $layer=LI1_cond $X=1.915 $Y=0.535
+ $X2=1.915 $Y2=1.535
r163 13 55 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=3.85 $Y=2.605
+ $X2=3.85 $Y2=2.235
r164 9 51 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=3.155 $Y=0.445
+ $X2=3.155 $Y2=0.975
r165 2 19 600 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_PDIFF $count=1 $X=1.915
+ $Y=2.395 $X2=2.04 $Y2=2.55
r166 1 34 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=2.005
+ $Y=0.235 $X2=2.13 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__DLRTP_2%A_796_21# 1 2 7 9 14 18 22 24 28 32 36 39 41
+ 44 48 51 54 58 61 66 68 74
c138 66 0 1.89225e-19 $X=5.355 $Y=2.445
c139 58 0 8.43473e-20 $X=6.13 $Y=1.51
c140 51 0 1.22782e-19 $X=5.04 $Y=1.905
c141 36 0 1.63114e-19 $X=4.24 $Y=0.84
c142 7 0 1.934e-19 $X=4.055 $Y=0.765
r143 73 74 30.474 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=6.265 $Y=1.51
+ $X2=6.34 $Y2=1.51
r144 64 66 9.11355 $w=5.02e-07 $l=3.75e-07 $layer=LI1_cond $X=5.212 $Y=2.07
+ $X2=5.212 $Y2=2.445
r145 63 64 1.45817 $w=5.02e-07 $l=6e-08 $layer=LI1_cond $X=5.212 $Y=2.01
+ $X2=5.212 $Y2=2.07
r146 59 73 23.6063 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=6.13 $Y=1.51
+ $X2=6.265 $Y2=1.51
r147 59 70 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=6.13 $Y=1.51 $X2=6.04
+ $Y2=1.51
r148 58 59 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.13
+ $Y=1.51 $X2=6.13 $Y2=1.51
r149 56 58 19.1306 $w=2.48e-07 $l=4.15e-07 $layer=LI1_cond $X=6.09 $Y=1.925
+ $X2=6.09 $Y2=1.51
r150 55 63 7.18174 $w=1.7e-07 $l=2.58e-07 $layer=LI1_cond $X=5.47 $Y=2.01
+ $X2=5.212 $Y2=2.01
r151 54 56 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=5.965 $Y=2.01
+ $X2=6.09 $Y2=1.925
r152 54 55 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=5.965 $Y=2.01
+ $X2=5.47 $Y2=2.01
r153 51 63 8.26182 $w=5.02e-07 $l=2.18275e-07 $layer=LI1_cond $X=5.04 $Y=1.905
+ $X2=5.212 $Y2=2.01
r154 51 61 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=5.04 $Y=1.905
+ $X2=5.04 $Y2=1.165
r155 46 61 8.16989 $w=3.13e-07 $l=1.57e-07 $layer=LI1_cond $X=4.967 $Y=1.008
+ $X2=4.967 $Y2=1.165
r156 46 48 18.2196 $w=3.13e-07 $l=4.98e-07 $layer=LI1_cond $X=4.967 $Y=1.008
+ $X2=4.967 $Y2=0.51
r157 44 69 46.255 $w=3.35e-07 $l=1.65e-07 $layer=POLY_cond $X=4.332 $Y=2.07
+ $X2=4.332 $Y2=2.235
r158 44 68 46.255 $w=3.35e-07 $l=1.65e-07 $layer=POLY_cond $X=4.332 $Y=2.07
+ $X2=4.332 $Y2=1.905
r159 43 44 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.335
+ $Y=2.07 $X2=4.335 $Y2=2.07
r160 41 64 3.19241 $w=3.3e-07 $l=2.57e-07 $layer=LI1_cond $X=4.955 $Y=2.07
+ $X2=5.212 $Y2=2.07
r161 41 43 21.652 $w=3.28e-07 $l=6.2e-07 $layer=LI1_cond $X=4.955 $Y=2.07
+ $X2=4.335 $Y2=2.07
r162 38 39 56.4043 $w=1.5e-07 $l=1.1e-07 $layer=POLY_cond $X=6.585 $Y=1.42
+ $X2=6.695 $Y2=1.42
r163 34 36 94.8617 $w=1.5e-07 $l=1.85e-07 $layer=POLY_cond $X=4.055 $Y=0.84
+ $X2=4.24 $Y2=0.84
r164 30 39 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.695 $Y=1.495
+ $X2=6.695 $Y2=1.42
r165 30 32 497.383 $w=1.5e-07 $l=9.7e-07 $layer=POLY_cond $X=6.695 $Y=1.495
+ $X2=6.695 $Y2=2.465
r166 26 38 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.585 $Y=1.345
+ $X2=6.585 $Y2=1.42
r167 26 28 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=6.585 $Y=1.345
+ $X2=6.585 $Y2=0.785
r168 24 38 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.51 $Y=1.42
+ $X2=6.585 $Y2=1.42
r169 24 74 87.1702 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=6.51 $Y=1.42
+ $X2=6.34 $Y2=1.42
r170 20 73 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.265 $Y=1.675
+ $X2=6.265 $Y2=1.51
r171 20 22 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=6.265 $Y=1.675
+ $X2=6.265 $Y2=2.465
r172 16 70 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.04 $Y=1.345
+ $X2=6.04 $Y2=1.51
r173 16 18 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=6.04 $Y=1.345
+ $X2=6.04 $Y2=0.785
r174 14 69 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=4.24 $Y=2.605
+ $X2=4.24 $Y2=2.235
r175 10 36 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.24 $Y=0.915
+ $X2=4.24 $Y2=0.84
r176 10 68 507.638 $w=1.5e-07 $l=9.9e-07 $layer=POLY_cond $X=4.24 $Y=0.915
+ $X2=4.24 $Y2=1.905
r177 7 34 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.055 $Y=0.765
+ $X2=4.055 $Y2=0.84
r178 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=4.055 $Y=0.765
+ $X2=4.055 $Y2=0.445
r179 2 66 300 $w=1.7e-07 $l=6.76387e-07 $layer=licon1_PDIFF $count=2 $X=5.215
+ $Y=1.835 $X2=5.355 $Y2=2.445
r180 2 63 600 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_PDIFF $count=1 $X=5.215
+ $Y=1.835 $X2=5.355 $Y2=2.01
r181 1 48 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=4.8
+ $Y=0.365 $X2=4.925 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_LP__DLRTP_2%A_646_47# 1 2 8 9 10 11 13 15 18 20 25 26 27
+ 29 30 31 37 40 41 42
c118 27 0 2.97881e-19 $X=3.525 $Y=1.64
r119 41 46 18.3619 $w=3.15e-07 $l=1.2e-07 $layer=POLY_cond $X=4.69 $Y=1.5
+ $X2=4.69 $Y2=1.62
r120 40 42 8.47458 $w=3.03e-07 $l=1.65e-07 $layer=LI1_cond $X=4.622 $Y=1.5
+ $X2=4.622 $Y2=1.335
r121 40 41 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.69
+ $Y=1.5 $X2=4.69 $Y2=1.5
r122 34 37 5.30124 $w=2.48e-07 $l=1.15e-07 $layer=LI1_cond $X=3.44 $Y=2.53
+ $X2=3.555 $Y2=2.53
r123 32 42 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=4.555 $Y=0.895
+ $X2=4.555 $Y2=1.335
r124 30 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.47 $Y=0.81
+ $X2=4.555 $Y2=0.895
r125 30 31 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=4.47 $Y=0.81
+ $X2=4.11 $Y2=0.81
r126 29 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.025 $Y=0.725
+ $X2=4.11 $Y2=0.81
r127 28 29 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=4.025 $Y=0.535
+ $X2=4.025 $Y2=0.725
r128 26 40 5.2899 $w=3.03e-07 $l=1.4e-07 $layer=LI1_cond $X=4.622 $Y=1.64
+ $X2=4.622 $Y2=1.5
r129 26 27 61.6524 $w=1.68e-07 $l=9.45e-07 $layer=LI1_cond $X=4.47 $Y=1.64
+ $X2=3.525 $Y2=1.64
r130 25 34 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.44 $Y=2.405
+ $X2=3.44 $Y2=2.53
r131 24 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.44 $Y=1.725
+ $X2=3.525 $Y2=1.64
r132 24 25 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=3.44 $Y=1.725
+ $X2=3.44 $Y2=2.405
r133 20 28 7.36005 $w=2.8e-07 $l=1.77482e-07 $layer=LI1_cond $X=3.94 $Y=0.395
+ $X2=4.025 $Y2=0.535
r134 20 22 18.933 $w=2.78e-07 $l=4.6e-07 $layer=LI1_cond $X=3.94 $Y=0.395
+ $X2=3.48 $Y2=0.395
r135 16 18 394.83 $w=1.5e-07 $l=7.7e-07 $layer=POLY_cond $X=5.14 $Y=1.695
+ $X2=5.14 $Y2=2.465
r136 13 15 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=5.14 $Y=0.255
+ $X2=5.14 $Y2=0.785
r137 12 46 20.1192 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.855 $Y=1.62
+ $X2=4.69 $Y2=1.62
r138 11 16 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.065 $Y=1.62
+ $X2=5.14 $Y2=1.695
r139 11 12 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=5.065 $Y=1.62
+ $X2=4.855 $Y2=1.62
r140 9 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.065 $Y=0.18
+ $X2=5.14 $Y2=0.255
r141 9 10 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=5.065 $Y=0.18
+ $X2=4.725 $Y2=0.18
r142 8 41 38.5363 $w=3.15e-07 $l=1.83916e-07 $layer=POLY_cond $X=4.65 $Y=1.335
+ $X2=4.69 $Y2=1.5
r143 7 10 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.65 $Y=0.255
+ $X2=4.725 $Y2=0.18
r144 7 8 553.787 $w=1.5e-07 $l=1.08e-06 $layer=POLY_cond $X=4.65 $Y=0.255
+ $X2=4.65 $Y2=1.335
r145 2 37 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=3.415
+ $Y=2.395 $X2=3.555 $Y2=2.54
r146 1 22 182 $w=1.7e-07 $l=3.29773e-07 $layer=licon1_NDIFF $count=1 $X=3.23
+ $Y=0.235 $X2=3.48 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__DLRTP_2%RESET_B 3 6 8 9 13 15
c39 15 0 1.22782e-19 $X=5.59 $Y=1.315
c40 13 0 1.89225e-19 $X=5.59 $Y=1.48
r41 13 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.59 $Y=1.48
+ $X2=5.59 $Y2=1.645
r42 13 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.59 $Y=1.48
+ $X2=5.59 $Y2=1.315
r43 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.59
+ $Y=1.48 $X2=5.59 $Y2=1.48
r44 9 14 6.66256 $w=3.18e-07 $l=1.85e-07 $layer=LI1_cond $X=5.515 $Y=1.665
+ $X2=5.515 $Y2=1.48
r45 8 14 6.66256 $w=3.18e-07 $l=1.85e-07 $layer=LI1_cond $X=5.515 $Y=1.295
+ $X2=5.515 $Y2=1.48
r46 6 16 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=5.57 $Y=2.465
+ $X2=5.57 $Y2=1.645
r47 3 15 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=5.5 $Y=0.785 $X2=5.5
+ $Y2=1.315
.ends

.subckt PM_SKY130_FD_SC_LP__DLRTP_2%VPWR 1 2 3 4 5 18 22 26 28 30 35 36 38 39 40
+ 42 54 65 70 77 81
r94 80 81 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r95 77 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r96 75 77 9.21893 $w=7.08e-07 $l=5.35e-07 $layer=LI1_cond $X=4.67 $Y=2.795
+ $X2=4.67 $Y2=3.33
r97 73 75 3.27401 $w=7.08e-07 $l=1.9e-07 $layer=LI1_cond $X=4.67 $Y=2.605
+ $X2=4.67 $Y2=2.795
r98 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r99 68 81 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=6.96 $Y2=3.33
r100 67 68 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r101 65 80 4.80598 $w=1.7e-07 $l=2.32e-07 $layer=LI1_cond $X=6.735 $Y=3.33
+ $X2=6.967 $Y2=3.33
r102 65 67 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=6.735 $Y=3.33
+ $X2=6.48 $Y2=3.33
r103 64 68 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=6.48 $Y2=3.33
r104 64 78 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=4.56 $Y2=3.33
r105 63 64 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r106 61 77 9.39643 $w=1.7e-07 $l=3.8e-07 $layer=LI1_cond $X=5.05 $Y=3.33
+ $X2=4.67 $Y2=3.33
r107 61 63 30.6631 $w=1.68e-07 $l=4.7e-07 $layer=LI1_cond $X=5.05 $Y=3.33
+ $X2=5.52 $Y2=3.33
r108 60 78 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r109 59 60 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r110 56 59 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=3.12 $Y=3.33
+ $X2=4.08 $Y2=3.33
r111 56 57 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r112 54 77 9.39643 $w=1.7e-07 $l=3.8e-07 $layer=LI1_cond $X=4.29 $Y=3.33
+ $X2=4.67 $Y2=3.33
r113 54 59 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=4.29 $Y=3.33
+ $X2=4.08 $Y2=3.33
r114 53 57 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r115 52 53 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r116 50 53 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r117 50 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r118 49 52 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r119 49 50 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r120 47 70 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.85 $Y=3.33
+ $X2=0.725 $Y2=3.33
r121 47 49 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=0.85 $Y=3.33
+ $X2=1.2 $Y2=3.33
r122 45 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r123 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r124 42 70 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.6 $Y=3.33
+ $X2=0.725 $Y2=3.33
r125 42 44 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=0.6 $Y=3.33
+ $X2=0.24 $Y2=3.33
r126 40 60 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r127 40 57 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=3.12 $Y2=3.33
r128 38 63 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=5.75 $Y=3.33
+ $X2=5.52 $Y2=3.33
r129 38 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.75 $Y=3.33
+ $X2=5.915 $Y2=3.33
r130 37 67 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=6.08 $Y=3.33 $X2=6.48
+ $Y2=3.33
r131 37 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.08 $Y=3.33
+ $X2=5.915 $Y2=3.33
r132 35 52 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=2.645 $Y=3.33
+ $X2=2.64 $Y2=3.33
r133 35 36 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.645 $Y=3.33
+ $X2=2.74 $Y2=3.33
r134 34 56 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=2.835 $Y=3.33
+ $X2=3.12 $Y2=3.33
r135 34 36 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.835 $Y=3.33
+ $X2=2.74 $Y2=3.33
r136 30 33 32.8785 $w=3.38e-07 $l=9.7e-07 $layer=LI1_cond $X=6.905 $Y=1.98
+ $X2=6.905 $Y2=2.95
r137 28 80 3.04517 $w=3.4e-07 $l=1.11781e-07 $layer=LI1_cond $X=6.905 $Y=3.245
+ $X2=6.967 $Y2=3.33
r138 28 33 9.99914 $w=3.38e-07 $l=2.95e-07 $layer=LI1_cond $X=6.905 $Y=3.245
+ $X2=6.905 $Y2=2.95
r139 24 39 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.915 $Y=3.245
+ $X2=5.915 $Y2=3.33
r140 24 26 30.208 $w=3.28e-07 $l=8.65e-07 $layer=LI1_cond $X=5.915 $Y=3.245
+ $X2=5.915 $Y2=2.38
r141 20 36 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=2.74 $Y=3.245
+ $X2=2.74 $Y2=3.33
r142 20 22 39.4019 $w=1.88e-07 $l=6.75e-07 $layer=LI1_cond $X=2.74 $Y=3.245
+ $X2=2.74 $Y2=2.57
r143 16 70 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.725 $Y=3.245
+ $X2=0.725 $Y2=3.33
r144 16 18 17.2866 $w=2.48e-07 $l=3.75e-07 $layer=LI1_cond $X=0.725 $Y=3.245
+ $X2=0.725 $Y2=2.87
r145 5 33 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=6.77
+ $Y=1.835 $X2=6.91 $Y2=2.95
r146 5 30 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=6.77
+ $Y=1.835 $X2=6.91 $Y2=1.98
r147 4 26 300 $w=1.7e-07 $l=6.66465e-07 $layer=licon1_PDIFF $count=2 $X=5.645
+ $Y=1.835 $X2=5.915 $Y2=2.38
r148 3 75 600 $w=1.7e-07 $l=7.8492e-07 $layer=licon1_PDIFF $count=1 $X=4.315
+ $Y=2.395 $X2=4.925 $Y2=2.795
r149 3 73 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=4.315
+ $Y=2.395 $X2=4.455 $Y2=2.605
r150 2 22 300 $w=1.7e-07 $l=4.89745e-07 $layer=licon1_PDIFF $count=2 $X=2.33
+ $Y=2.395 $X2=2.74 $Y2=2.57
r151 1 18 600 $w=1.7e-07 $l=5.60647e-07 $layer=licon1_PDIFF $count=1 $X=0.615
+ $Y=2.375 $X2=0.755 $Y2=2.87
.ends

.subckt PM_SKY130_FD_SC_LP__DLRTP_2%Q 1 2 7 8 9 10 11 12 13 24 30
r23 22 30 1.36586 $w=4.03e-07 $l=4.8e-08 $layer=LI1_cond $X=6.362 $Y=0.973
+ $X2=6.362 $Y2=0.925
r24 13 44 8.31818 $w=1.78e-07 $l=1.35e-07 $layer=LI1_cond $X=6.475 $Y=2.775
+ $X2=6.475 $Y2=2.91
r25 12 13 22.798 $w=1.78e-07 $l=3.7e-07 $layer=LI1_cond $X=6.475 $Y=2.405
+ $X2=6.475 $Y2=2.775
r26 11 12 26.1869 $w=1.78e-07 $l=4.25e-07 $layer=LI1_cond $X=6.475 $Y=1.98
+ $X2=6.475 $Y2=2.405
r27 10 11 19.4091 $w=1.78e-07 $l=3.15e-07 $layer=LI1_cond $X=6.475 $Y=1.665
+ $X2=6.475 $Y2=1.98
r28 9 10 22.798 $w=1.78e-07 $l=3.7e-07 $layer=LI1_cond $X=6.475 $Y=1.295
+ $X2=6.475 $Y2=1.665
r29 9 47 7.39394 $w=1.78e-07 $l=1.2e-07 $layer=LI1_cond $X=6.475 $Y=1.295
+ $X2=6.475 $Y2=1.175
r30 8 47 8.84441 $w=4.03e-07 $l=1.84e-07 $layer=LI1_cond $X=6.362 $Y=0.991
+ $X2=6.362 $Y2=1.175
r31 8 22 0.512197 $w=4.03e-07 $l=1.8e-08 $layer=LI1_cond $X=6.362 $Y=0.991
+ $X2=6.362 $Y2=0.973
r32 8 30 0.540652 $w=4.03e-07 $l=1.9e-08 $layer=LI1_cond $X=6.362 $Y=0.906
+ $X2=6.362 $Y2=0.925
r33 7 8 9.98784 $w=4.03e-07 $l=3.51e-07 $layer=LI1_cond $X=6.362 $Y=0.555
+ $X2=6.362 $Y2=0.906
r34 7 24 1.28049 $w=4.03e-07 $l=4.5e-08 $layer=LI1_cond $X=6.362 $Y=0.555
+ $X2=6.362 $Y2=0.51
r35 2 44 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=6.34
+ $Y=1.835 $X2=6.48 $Y2=2.91
r36 2 11 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=6.34
+ $Y=1.835 $X2=6.48 $Y2=1.98
r37 1 24 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=6.115
+ $Y=0.365 $X2=6.325 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_LP__DLRTP_2%VGND 1 2 3 4 5 18 22 26 30 32 34 37 38 40 41
+ 43 44 45 51 71 76 80
r103 79 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r104 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r105 74 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6.96
+ $Y2=0
r106 73 74 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r107 71 79 3.90852 $w=1.7e-07 $l=2.32e-07 $layer=LI1_cond $X=6.735 $Y=0
+ $X2=6.967 $Y2=0
r108 71 73 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=6.735 $Y=0
+ $X2=6.48 $Y2=0
r109 70 74 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=6.48
+ $Y2=0
r110 69 70 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r111 67 70 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.52
+ $Y2=0
r112 66 69 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=4.56 $Y=0 $X2=5.52
+ $Y2=0
r113 66 67 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r114 64 67 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=4.56
+ $Y2=0
r115 63 64 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r116 61 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.64
+ $Y2=0
r117 60 63 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=3.12 $Y=0 $X2=4.08
+ $Y2=0
r118 60 61 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r119 58 76 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=2.745 $Y=0 $X2=2.605
+ $Y2=0
r120 58 60 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=2.745 $Y=0
+ $X2=3.12 $Y2=0
r121 57 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r122 56 57 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r123 54 57 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r124 53 56 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r125 53 54 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r126 51 76 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=2.465 $Y=0 $X2=2.605
+ $Y2=0
r127 51 56 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.465 $Y=0
+ $X2=2.16 $Y2=0
r128 49 54 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r129 48 49 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r130 45 64 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r131 45 61 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=3.12
+ $Y2=0
r132 43 69 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=5.605 $Y=0 $X2=5.52
+ $Y2=0
r133 43 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.605 $Y=0 $X2=5.77
+ $Y2=0
r134 42 73 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=5.935 $Y=0
+ $X2=6.48 $Y2=0
r135 42 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.935 $Y=0 $X2=5.77
+ $Y2=0
r136 40 63 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=4.28 $Y=0 $X2=4.08
+ $Y2=0
r137 40 41 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=4.28 $Y=0 $X2=4.38
+ $Y2=0
r138 39 66 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=4.48 $Y=0 $X2=4.56
+ $Y2=0
r139 39 41 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=4.48 $Y=0 $X2=4.38
+ $Y2=0
r140 37 48 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.975 $Y=0
+ $X2=0.72 $Y2=0
r141 37 38 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=0.975 $Y=0 $X2=1.075
+ $Y2=0
r142 36 53 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=1.175 $Y=0 $X2=1.2
+ $Y2=0
r143 36 38 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=1.175 $Y=0 $X2=1.075
+ $Y2=0
r144 32 79 3.23464 $w=2.5e-07 $l=1.43332e-07 $layer=LI1_cond $X=6.86 $Y=0.085
+ $X2=6.967 $Y2=0
r145 32 34 19.5915 $w=2.48e-07 $l=4.25e-07 $layer=LI1_cond $X=6.86 $Y=0.085
+ $X2=6.86 $Y2=0.51
r146 28 44 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.77 $Y=0.085
+ $X2=5.77 $Y2=0
r147 28 30 14.8421 $w=3.28e-07 $l=4.25e-07 $layer=LI1_cond $X=5.77 $Y=0.085
+ $X2=5.77 $Y2=0.51
r148 24 41 0.764409 $w=2e-07 $l=8.5e-08 $layer=LI1_cond $X=4.38 $Y=0.085
+ $X2=4.38 $Y2=0
r149 24 26 16.9136 $w=1.98e-07 $l=3.05e-07 $layer=LI1_cond $X=4.38 $Y=0.085
+ $X2=4.38 $Y2=0.39
r150 20 76 0.375625 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.605 $Y=0.085
+ $X2=2.605 $Y2=0
r151 20 22 11.7302 $w=2.78e-07 $l=2.85e-07 $layer=LI1_cond $X=2.605 $Y=0.085
+ $X2=2.605 $Y2=0.37
r152 16 38 0.764409 $w=2e-07 $l=8.5e-08 $layer=LI1_cond $X=1.075 $Y=0.085
+ $X2=1.075 $Y2=0
r153 16 18 21.9045 $w=1.98e-07 $l=3.95e-07 $layer=LI1_cond $X=1.075 $Y=0.085
+ $X2=1.075 $Y2=0.48
r154 5 34 91 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_NDIFF $count=2 $X=6.66
+ $Y=0.365 $X2=6.82 $Y2=0.51
r155 4 30 91 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_NDIFF $count=2 $X=5.575
+ $Y=0.365 $X2=5.77 $Y2=0.51
r156 3 26 182 $w=1.7e-07 $l=3.02738e-07 $layer=licon1_NDIFF $count=1 $X=4.13
+ $Y=0.235 $X2=4.365 $Y2=0.39
r157 2 22 182 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_NDIFF $count=1 $X=2.44
+ $Y=0.235 $X2=2.58 $Y2=0.37
r158 1 18 182 $w=1.7e-07 $l=5.50068e-07 $layer=licon1_NDIFF $count=1 $X=0.615
+ $Y=0.27 $X2=1.07 $Y2=0.48
.ends

