* File: sky130_fd_sc_lp__or4b_2.spice
* Created: Wed Sep  2 10:32:34 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__or4b_2.pex.spice"
.subckt sky130_fd_sc_lp__or4b_2  VNB VPB D_N A B C VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* C	C
* B	B
* A	A
* D_N	D_N
* VPB	VPB
* VNB	VNB
MM1012 N_VGND_M1012_d N_D_N_M1012_g N_A_31_131#_M1012_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0896 AS=0.1113 PD=0.81 PS=1.37 NRD=28.56 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1002 N_X_M1002_d N_A_189_21#_M1002_g N_VGND_M1012_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1792 PD=1.12 PS=1.62 NRD=0 NRS=0 M=1 R=5.6 SA=75000.5
+ SB=75001.6 A=0.126 P=1.98 MULT=1
MM1007 N_X_M1002_d N_A_189_21#_M1007_g N_VGND_M1007_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1792 PD=1.12 PS=1.62 NRD=0 NRS=6.78 M=1 R=5.6 SA=75000.9
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1010 N_A_189_21#_M1010_d N_A_M1010_g N_VGND_M1007_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0896 PD=0.7 PS=0.81 NRD=0 NRS=0 M=1 R=2.8 SA=75001.1 SB=75001.6
+ A=0.063 P=1.14 MULT=1
MM1005 N_VGND_M1005_d N_B_M1005_g N_A_189_21#_M1010_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0798 AS=0.0588 PD=0.8 PS=0.7 NRD=8.568 NRS=0 M=1 R=2.8 SA=75001.6
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1001 N_A_189_21#_M1001_d N_C_M1001_g N_VGND_M1005_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0798 PD=0.7 PS=0.8 NRD=0 NRS=19.992 M=1 R=2.8 SA=75002.1
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1011 N_VGND_M1011_d N_A_31_131#_M1011_g N_A_189_21#_M1001_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75002.5
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1008 N_VPWR_M1008_d N_D_N_M1008_g N_A_31_131#_M1008_s VPB PHIGHVT L=0.15
+ W=0.42 AD=0.095025 AS=0.1113 PD=0.8175 PS=1.37 NRD=80.3169 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75002.6 A=0.063 P=1.14 MULT=1
MM1000 N_X_M1000_d N_A_189_21#_M1000_g N_VPWR_M1008_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.285075 PD=1.54 PS=2.4525 NRD=0 NRS=0 M=1 R=8.4 SA=75000.4
+ SB=75001.3 A=0.189 P=2.82 MULT=1
MM1009 N_X_M1000_d N_A_189_21#_M1009_g N_VPWR_M1009_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.326025 PD=1.54 PS=2.6475 NRD=0 NRS=0 M=1 R=8.4 SA=75000.8
+ SB=75000.8 A=0.189 P=2.82 MULT=1
MM1003 A_436_385# N_A_M1003_g N_VPWR_M1009_s VPB PHIGHVT L=0.15 W=0.42 AD=0.0441
+ AS=0.108675 PD=0.63 PS=0.8825 NRD=23.443 NRS=95.5647 M=1 R=2.8 SA=75001.7
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1013 A_508_385# N_B_M1013_g A_436_385# VPB PHIGHVT L=0.15 W=0.42 AD=0.0819
+ AS=0.0441 PD=0.81 PS=0.63 NRD=65.6601 NRS=23.443 M=1 R=2.8 SA=75002 SB=75001.1
+ A=0.063 P=1.14 MULT=1
MM1004 A_616_385# N_C_M1004_g A_508_385# VPB PHIGHVT L=0.15 W=0.42 AD=0.0441
+ AS=0.0819 PD=0.63 PS=0.81 NRD=23.443 NRS=65.6601 M=1 R=2.8 SA=75002.6
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1006 N_A_189_21#_M1006_d N_A_31_131#_M1006_g A_616_385# VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1113 AS=0.0441 PD=1.37 PS=0.63 NRD=0 NRS=23.443 M=1 R=2.8
+ SA=75002.9 SB=75000.2 A=0.063 P=1.14 MULT=1
DX14_noxref VNB VPB NWDIODE A=7.8703 P=12.17
c_79 VPB 0 6.20762e-20 $X=0 $Y=3.085
*
.include "sky130_fd_sc_lp__or4b_2.pxi.spice"
*
.ends
*
*
