# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__ebufn_lp
  CLASS CORE ;
  FOREIGN sky130_fd_sc_lp__ebufn_lp ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.320000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.490000 1.245000 0.835000 2.150000 ;
    END
  END A
  PIN TE_B
    ANTENNAGATEAREA  0.507000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.440000 1.175000 3.770000 1.780000 ;
    END
  END TE_B
  PIN Z
    ANTENNADIFFAREA  0.598500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.905000 0.595000 2.405000 1.005000 ;
        RECT 1.905000 1.005000 2.575000 1.175000 ;
        RECT 2.120000 2.025000 2.755000 2.890000 ;
        RECT 2.120000 2.890000 2.450000 3.075000 ;
        RECT 2.405000 1.175000 2.755000 2.025000 ;
    END
  END Z
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.320000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.320000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.320000 0.085000 ;
      RECT 0.000000  3.245000 4.320000 3.415000 ;
      RECT 0.125000  0.635000 0.485000 1.075000 ;
      RECT 0.125000  1.075000 0.295000 2.395000 ;
      RECT 0.125000  2.395000 1.175000 2.565000 ;
      RECT 0.125000  2.565000 0.455000 3.075000 ;
      RECT 1.005000  1.685000 2.235000 1.855000 ;
      RECT 1.005000  1.855000 1.175000 2.395000 ;
      RECT 1.065000  0.085000 1.395000 1.015000 ;
      RECT 1.210000  1.185000 1.735000 1.515000 ;
      RECT 1.345000  2.395000 1.675000 3.245000 ;
      RECT 1.565000  0.255000 2.915000 0.425000 ;
      RECT 1.565000  0.425000 1.735000 1.185000 ;
      RECT 1.905000  1.345000 2.235000 1.685000 ;
      RECT 2.745000  0.425000 2.915000 0.835000 ;
      RECT 2.745000  0.835000 4.205000 1.005000 ;
      RECT 2.940000  1.815000 3.270000 3.245000 ;
      RECT 3.085000  0.085000 3.415000 0.665000 ;
      RECT 3.875000  0.255000 4.205000 0.835000 ;
      RECT 3.875000  1.985000 4.205000 2.665000 ;
      RECT 4.035000  1.005000 4.205000 1.985000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
  END
END sky130_fd_sc_lp__ebufn_lp
END LIBRARY
