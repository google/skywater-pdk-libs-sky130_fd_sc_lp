* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__o32ai_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
X0 a_778_365# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X1 Y B2 a_39_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X2 VGND A1 a_39_65# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X3 a_39_367# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X4 VGND A2 a_39_65# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X5 a_519_365# A3 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X6 a_39_65# A1 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X7 a_39_367# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X8 a_39_65# B1 Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X9 a_519_365# A2 a_778_365# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X10 Y B1 a_39_65# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X11 VGND A3 a_39_65# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X12 Y A3 a_519_365# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X13 Y B2 a_39_65# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X14 a_39_65# A3 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X15 VPWR B1 a_39_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X16 a_778_365# A2 a_519_365# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X17 VPWR A1 a_778_365# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X18 a_39_65# B2 Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X19 a_39_65# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
.ends
