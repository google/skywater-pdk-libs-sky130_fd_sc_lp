* File: sky130_fd_sc_lp__o221a_m.pex.spice
* Created: Wed Sep  2 10:18:45 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O221A_M%C1 2 6 7 9 12 16 18 19 23
c43 6 0 7.46275e-20 $X=0.475 $Y=1.105
r44 23 26 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.455 $Y=0.555
+ $X2=0.455 $Y2=0.72
r45 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.455
+ $Y=0.555 $X2=0.455 $Y2=0.555
r46 19 24 9.25447 $w=3.28e-07 $l=2.65e-07 $layer=LI1_cond $X=0.72 $Y=0.555
+ $X2=0.455 $Y2=0.555
r47 18 24 7.50834 $w=3.28e-07 $l=2.15e-07 $layer=LI1_cond $X=0.24 $Y=0.555
+ $X2=0.455 $Y2=0.555
r48 14 16 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=0.28 $Y=2.49
+ $X2=0.52 $Y2=2.49
r49 10 12 99.9894 $w=1.5e-07 $l=1.95e-07 $layer=POLY_cond $X=0.28 $Y=1.53
+ $X2=0.475 $Y2=1.53
r50 7 16 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.52 $Y=2.565
+ $X2=0.52 $Y2=2.49
r51 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.52 $Y=2.565 $X2=0.52
+ $Y2=2.885
r52 6 26 197.415 $w=1.5e-07 $l=3.85e-07 $layer=POLY_cond $X=0.475 $Y=1.105
+ $X2=0.475 $Y2=0.72
r53 4 12 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.475 $Y=1.455
+ $X2=0.475 $Y2=1.53
r54 4 6 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=0.475 $Y=1.455
+ $X2=0.475 $Y2=1.105
r55 2 14 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.28 $Y=2.415
+ $X2=0.28 $Y2=2.49
r56 1 10 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.28 $Y=1.605
+ $X2=0.28 $Y2=1.53
r57 1 2 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=0.28 $Y=1.605 $X2=0.28
+ $Y2=2.415
.ends

.subckt PM_SKY130_FD_SC_LP__O221A_M%B1 4 7 10 12 13 16 18 21 23
c59 21 0 1.90606e-19 $X=0.76 $Y=2.01
c60 16 0 1.6235e-20 $X=1.115 $Y=2.46
r61 21 24 46.5827 $w=3.6e-07 $l=1.65e-07 $layer=POLY_cond $X=0.775 $Y=2.01
+ $X2=0.775 $Y2=2.175
r62 21 23 46.5827 $w=3.6e-07 $l=1.65e-07 $layer=POLY_cond $X=0.775 $Y=2.01
+ $X2=0.775 $Y2=1.845
r63 18 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.76
+ $Y=2.01 $X2=0.76 $Y2=2.01
r64 14 16 120.5 $w=1.5e-07 $l=2.35e-07 $layer=POLY_cond $X=0.88 $Y=2.46
+ $X2=1.115 $Y2=2.46
r65 13 23 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=0.85 $Y=1.575
+ $X2=0.85 $Y2=1.845
r66 12 13 48.5235 $w=2.05e-07 $l=1.5e-07 $layer=POLY_cond $X=0.877 $Y=1.425
+ $X2=0.877 $Y2=1.575
r67 8 16 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.115 $Y=2.535
+ $X2=1.115 $Y2=2.46
r68 8 10 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=1.115 $Y=2.535
+ $X2=1.115 $Y2=2.885
r69 7 12 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.905 $Y=1.105
+ $X2=0.905 $Y2=1.425
r70 4 14 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.88 $Y=2.385
+ $X2=0.88 $Y2=2.46
r71 4 24 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=0.88 $Y=2.385
+ $X2=0.88 $Y2=2.175
.ends

.subckt PM_SKY130_FD_SC_LP__O221A_M%B2 5 9 10 11 12 15 16 17
c44 16 0 1.3013e-19 $X=1.33 $Y=1.98
c45 5 0 1.39673e-19 $X=1.475 $Y=2.885
r46 15 18 45.3519 $w=3.85e-07 $l=1.65e-07 $layer=POLY_cond $X=1.357 $Y=1.98
+ $X2=1.357 $Y2=2.145
r47 15 17 45.3519 $w=3.85e-07 $l=1.65e-07 $layer=POLY_cond $X=1.357 $Y=1.98
+ $X2=1.357 $Y2=1.815
r48 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.33
+ $Y=1.98 $X2=1.33 $Y2=1.98
r49 12 16 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=1.2 $Y=1.98 $X2=1.33
+ $Y2=1.98
r50 11 17 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=1.475 $Y=1.605
+ $X2=1.475 $Y2=1.815
r51 10 11 49.7366 $w=2e-07 $l=1.5e-07 $layer=POLY_cond $X=1.5 $Y=1.455 $X2=1.5
+ $Y2=1.605
r52 9 10 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.525 $Y=1.135
+ $X2=1.525 $Y2=1.455
r53 5 18 379.447 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=1.475 $Y=2.885
+ $X2=1.475 $Y2=2.145
.ends

.subckt PM_SKY130_FD_SC_LP__O221A_M%A2 3 9 11 12 13 14 15 16 17 21 22
c50 15 0 7.74767e-20 $X=2.02 $Y=0.915
c51 13 0 1.52574e-20 $X=1.925 $Y=2.515
c52 11 0 1.3013e-19 $X=1.925 $Y=1.845
r53 21 22 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.925
+ $Y=2.01 $X2=1.925 $Y2=2.01
r54 16 17 10.2748 $w=4.13e-07 $l=3.7e-07 $layer=LI1_cond $X=1.802 $Y=2.035
+ $X2=1.802 $Y2=2.405
r55 16 22 0.694243 $w=4.13e-07 $l=2.5e-08 $layer=LI1_cond $X=1.802 $Y=2.035
+ $X2=1.802 $Y2=2.01
r56 14 15 69.5192 $w=1.6e-07 $l=1.5e-07 $layer=POLY_cond $X=2.02 $Y=0.765
+ $X2=2.02 $Y2=0.915
r57 12 21 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.925 $Y=2.35
+ $X2=1.925 $Y2=2.01
r58 12 13 38.6168 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.925 $Y=2.35
+ $X2=1.925 $Y2=2.515
r59 11 21 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.925 $Y=1.845
+ $X2=1.925 $Y2=2.01
r60 11 15 476.872 $w=1.5e-07 $l=9.3e-07 $layer=POLY_cond $X=2.015 $Y=1.845
+ $X2=2.015 $Y2=0.915
r61 9 14 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.025 $Y=0.445
+ $X2=2.025 $Y2=0.765
r62 3 13 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=1.905 $Y=2.885
+ $X2=1.905 $Y2=2.515
.ends

.subckt PM_SKY130_FD_SC_LP__O221A_M%A1 3 7 11 12 13 14 18 19
c51 7 0 1.19165e-19 $X=2.455 $Y=0.445
r52 18 19 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.465
+ $Y=1.255 $X2=2.465 $Y2=1.255
r53 13 14 9.31682 $w=4.73e-07 $l=3.7e-07 $layer=LI1_cond $X=2.537 $Y=1.295
+ $X2=2.537 $Y2=1.665
r54 13 19 1.00722 $w=4.73e-07 $l=4e-08 $layer=LI1_cond $X=2.537 $Y=1.295
+ $X2=2.537 $Y2=1.255
r55 11 18 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.465 $Y=1.595
+ $X2=2.465 $Y2=1.255
r56 11 12 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.465 $Y=1.595
+ $X2=2.465 $Y2=1.76
r57 10 18 38.0424 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.465 $Y=1.09
+ $X2=2.465 $Y2=1.255
r58 7 10 330.734 $w=1.5e-07 $l=6.45e-07 $layer=POLY_cond $X=2.455 $Y=0.445
+ $X2=2.455 $Y2=1.09
r59 3 12 576.862 $w=1.5e-07 $l=1.125e-06 $layer=POLY_cond $X=2.375 $Y=2.885
+ $X2=2.375 $Y2=1.76
.ends

.subckt PM_SKY130_FD_SC_LP__O221A_M%A_27_179# 1 2 3 12 16 19 20 23 25 27 32 33
+ 35 36 38 43 48
c106 43 0 1.52574e-20 $X=1.33 $Y=2.58
c107 38 0 1.6235e-20 $X=0.305 $Y=2.58
c108 25 0 1.39673e-19 $X=1.245 $Y=2.58
r109 38 41 8.3814 $w=3.28e-07 $l=2.4e-07 $layer=LI1_cond $X=0.305 $Y=2.58
+ $X2=0.305 $Y2=2.82
r110 38 39 4.14275 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=0.305 $Y=2.58
+ $X2=0.305 $Y2=2.495
r111 36 48 46.5827 $w=3.6e-07 $l=1.65e-07 $layer=POLY_cond $X=2.84 $Y=2.135
+ $X2=2.84 $Y2=1.97
r112 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.825
+ $Y=2.135 $X2=2.825 $Y2=2.135
r113 33 35 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=2.36 $Y=2.135
+ $X2=2.825 $Y2=2.135
r114 31 33 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.275 $Y=2.3
+ $X2=2.36 $Y2=2.135
r115 31 32 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=2.275 $Y=2.3
+ $X2=2.275 $Y2=2.695
r116 28 43 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=1.33 $Y=2.86
+ $X2=1.33 $Y2=2.58
r117 28 30 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=1.415 $Y=2.86
+ $X2=1.69 $Y2=2.86
r118 27 32 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.19 $Y=2.86
+ $X2=2.275 $Y2=2.695
r119 27 30 17.4613 $w=3.28e-07 $l=5e-07 $layer=LI1_cond $X=2.19 $Y=2.86 $X2=1.69
+ $Y2=2.86
r120 26 38 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.47 $Y=2.58
+ $X2=0.305 $Y2=2.58
r121 25 43 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.245 $Y=2.58
+ $X2=1.33 $Y2=2.58
r122 25 26 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=1.245 $Y=2.58
+ $X2=0.47 $Y2=2.58
r123 23 39 67.8661 $w=2.23e-07 $l=1.325e-06 $layer=LI1_cond $X=0.252 $Y=1.17
+ $X2=0.252 $Y2=2.495
r124 20 48 558.915 $w=1.5e-07 $l=1.09e-06 $layer=POLY_cond $X=2.945 $Y=0.88
+ $X2=2.945 $Y2=1.97
r125 19 20 47.3682 $w=2.1e-07 $l=1.5e-07 $layer=POLY_cond $X=2.915 $Y=0.73
+ $X2=2.915 $Y2=0.88
r126 16 19 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.885 $Y=0.445
+ $X2=2.885 $Y2=0.73
r127 10 36 46.5827 $w=3.6e-07 $l=1.65e-07 $layer=POLY_cond $X=2.84 $Y=2.3
+ $X2=2.84 $Y2=2.135
r128 10 12 299.968 $w=1.5e-07 $l=5.85e-07 $layer=POLY_cond $X=2.84 $Y=2.3
+ $X2=2.84 $Y2=2.885
r129 3 30 600 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_PDIFF $count=1 $X=1.55
+ $Y=2.675 $X2=1.69 $Y2=2.86
r130 2 41 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.18
+ $Y=2.675 $X2=0.305 $Y2=2.82
r131 1 23 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.895 $X2=0.26 $Y2=1.17
.ends

.subckt PM_SKY130_FD_SC_LP__O221A_M%VPWR 1 2 11 15 17 19 29 30 33 36
r46 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r47 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r48 30 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.64 $Y2=3.33
r49 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r50 27 36 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.73 $Y=3.33
+ $X2=2.635 $Y2=3.33
r51 27 29 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=2.73 $Y=3.33
+ $X2=3.12 $Y2=3.33
r52 26 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r53 25 26 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r54 23 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r55 22 25 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=3.33 $X2=2.16
+ $Y2=3.33
r56 22 23 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r57 20 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.98 $Y=3.33
+ $X2=0.815 $Y2=3.33
r58 20 22 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=0.98 $Y=3.33 $X2=1.2
+ $Y2=3.33
r59 19 36 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.54 $Y=3.33
+ $X2=2.635 $Y2=3.33
r60 19 25 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=2.54 $Y=3.33
+ $X2=2.16 $Y2=3.33
r61 17 26 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r62 17 23 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r63 13 36 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=2.635 $Y=3.245
+ $X2=2.635 $Y2=3.33
r64 13 15 17.2201 $w=1.88e-07 $l=2.95e-07 $layer=LI1_cond $X=2.635 $Y=3.245
+ $X2=2.635 $Y2=2.95
r65 9 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.815 $Y=3.245
+ $X2=0.815 $Y2=3.33
r66 9 11 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.815 $Y=3.245
+ $X2=0.815 $Y2=2.95
r67 2 15 600 $w=1.7e-07 $l=3.51781e-07 $layer=licon1_PDIFF $count=1 $X=2.45
+ $Y=2.675 $X2=2.625 $Y2=2.95
r68 1 11 600 $w=1.7e-07 $l=3.68951e-07 $layer=licon1_PDIFF $count=1 $X=0.595
+ $Y=2.675 $X2=0.815 $Y2=2.95
.ends

.subckt PM_SKY130_FD_SC_LP__O221A_M%X 1 2 10 11 13 14 15 16 36
r28 23 36 2.04396 $w=2.63e-07 $l=4.7e-08 $layer=LI1_cond $X=3.127 $Y=1.618
+ $X2=3.127 $Y2=1.665
r29 16 36 0.82628 $w=2.63e-07 $l=1.9e-08 $layer=LI1_cond $X=3.127 $Y=1.684
+ $X2=3.127 $Y2=1.665
r30 16 23 0.82628 $w=2.63e-07 $l=1.9e-08 $layer=LI1_cond $X=3.127 $Y=1.599
+ $X2=3.127 $Y2=1.618
r31 15 16 13.2205 $w=2.63e-07 $l=3.04e-07 $layer=LI1_cond $X=3.127 $Y=1.295
+ $X2=3.127 $Y2=1.599
r32 14 15 16.0907 $w=2.63e-07 $l=3.7e-07 $layer=LI1_cond $X=3.127 $Y=0.925
+ $X2=3.127 $Y2=1.295
r33 13 14 18.0477 $w=2.63e-07 $l=4.15e-07 $layer=LI1_cond $X=3.127 $Y=0.51
+ $X2=3.127 $Y2=0.925
r34 11 16 37.8325 $w=2.83e-07 $l=9.05e-07 $layer=LI1_cond $X=3.175 $Y=2.655
+ $X2=3.175 $Y2=1.75
r35 10 11 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.175 $Y=2.82
+ $X2=3.175 $Y2=2.655
r36 8 10 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=3.055 $Y=2.82
+ $X2=3.175 $Y2=2.82
r37 2 8 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.915
+ $Y=2.675 $X2=3.055 $Y2=2.82
r38 1 13 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=2.96
+ $Y=0.235 $X2=3.1 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_LP__O221A_M%A_110_179# 1 2 9 11 12 15
c29 11 0 1.90606e-19 $X=1.635 $Y=1.41
c30 9 0 1.99117e-19 $X=0.69 $Y=1.17
r31 13 15 6.60173 $w=2.08e-07 $l=1.25e-07 $layer=LI1_cond $X=1.74 $Y=1.325
+ $X2=1.74 $Y2=1.2
r32 11 13 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=1.635 $Y=1.41
+ $X2=1.74 $Y2=1.325
r33 11 12 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=1.635 $Y=1.41
+ $X2=0.795 $Y2=1.41
r34 7 12 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=0.69 $Y=1.325
+ $X2=0.795 $Y2=1.41
r35 7 9 8.18615 $w=2.08e-07 $l=1.55e-07 $layer=LI1_cond $X=0.69 $Y=1.325
+ $X2=0.69 $Y2=1.17
r36 2 15 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=1.6
+ $Y=0.925 $X2=1.74 $Y2=1.2
r37 1 9 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.895 $X2=0.69 $Y2=1.17
.ends

.subckt PM_SKY130_FD_SC_LP__O221A_M%A_196_179# 1 2 7 11 13
c31 13 0 7.74767e-20 $X=1.215 $Y=0.75
c32 11 0 2.89257e-19 $X=2.24 $Y=0.51
r33 13 16 10.1275 $w=3.28e-07 $l=2.9e-07 $layer=LI1_cond $X=1.215 $Y=0.75
+ $X2=1.215 $Y2=1.04
r34 9 11 8.18615 $w=2.08e-07 $l=1.55e-07 $layer=LI1_cond $X=2.24 $Y=0.665
+ $X2=2.24 $Y2=0.51
r35 8 13 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.38 $Y=0.75
+ $X2=1.215 $Y2=0.75
r36 7 9 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=2.135 $Y=0.75
+ $X2=2.24 $Y2=0.665
r37 7 8 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=2.135 $Y=0.75
+ $X2=1.38 $Y2=0.75
r38 2 11 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=2.1
+ $Y=0.235 $X2=2.24 $Y2=0.51
r39 1 16 182 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_NDIFF $count=1 $X=0.98
+ $Y=0.895 $X2=1.215 $Y2=1.04
.ends

.subckt PM_SKY130_FD_SC_LP__O221A_M%VGND 1 2 9 11 15 17 19 26 27 30 33
r40 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r41 27 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.64
+ $Y2=0
r42 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r43 24 33 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=2.775 $Y=0 $X2=2.67
+ $Y2=0
r44 24 26 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=2.775 $Y=0 $X2=3.12
+ $Y2=0
r45 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r46 19 30 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.625 $Y=0 $X2=1.79
+ $Y2=0
r47 19 21 90.3583 $w=1.68e-07 $l=1.385e-06 $layer=LI1_cond $X=1.625 $Y=0
+ $X2=0.24 $Y2=0
r48 17 34 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r49 17 22 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.68 $Y=0 $X2=0.24
+ $Y2=0
r50 17 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r51 13 33 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=2.67 $Y=0.085
+ $X2=2.67 $Y2=0
r52 13 15 15.5801 $w=2.08e-07 $l=2.95e-07 $layer=LI1_cond $X=2.67 $Y=0.085
+ $X2=2.67 $Y2=0.38
r53 12 30 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.955 $Y=0 $X2=1.79
+ $Y2=0
r54 11 33 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=2.565 $Y=0 $X2=2.67
+ $Y2=0
r55 11 12 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=2.565 $Y=0 $X2=1.955
+ $Y2=0
r56 7 30 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.79 $Y=0.085 $X2=1.79
+ $Y2=0
r57 7 9 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.79 $Y=0.085
+ $X2=1.79 $Y2=0.38
r58 2 15 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=2.53
+ $Y=0.235 $X2=2.67 $Y2=0.38
r59 1 9 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=1.665
+ $Y=0.235 $X2=1.79 $Y2=0.38
.ends

