* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__busdriver_20 A TE_B VGND VNB VPB VPWR Z
X0 VPWR a_286_367# a_630_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X1 a_630_367# a_286_367# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X2 a_1909_21# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X3 Z a_1909_21# a_584_47# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X4 a_584_47# a_114_47# VGND VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X5 VPWR a_286_367# a_630_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X6 a_630_367# a_286_367# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X7 VGND TE_B a_114_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X8 a_584_47# a_114_47# VGND VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X9 VGND a_114_47# a_584_47# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X10 Z a_1909_21# a_584_47# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X11 a_584_47# a_1909_21# Z VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X12 VGND A a_1909_21# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X13 a_630_367# a_286_367# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X14 a_630_367# a_1909_21# Z VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X15 VGND a_114_47# a_584_47# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X16 VGND a_114_47# a_584_47# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X17 a_584_47# a_114_47# VGND VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X18 a_286_367# a_114_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X19 VPWR a_286_367# a_630_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X20 Z a_1909_21# a_630_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X21 a_630_367# a_1909_21# Z VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X22 Z a_1909_21# a_630_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X23 VGND a_114_47# a_584_47# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X24 a_584_47# a_1909_21# Z VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X25 Z a_1909_21# a_630_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X26 a_1909_21# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X27 VPWR a_286_367# a_630_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X28 VPWR a_286_367# a_630_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X29 a_630_367# a_1909_21# Z VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X30 VPWR A a_1909_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X31 Z a_1909_21# a_584_47# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X32 a_630_367# a_286_367# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X33 a_584_47# a_1909_21# Z VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X34 a_630_367# a_286_367# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X35 a_630_367# a_286_367# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X36 VGND a_114_47# a_584_47# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X37 VPWR a_286_367# a_630_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X38 VPWR a_286_367# a_630_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X39 Z a_1909_21# a_584_47# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X40 a_630_367# a_286_367# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X41 a_630_367# a_1909_21# Z VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X42 a_286_367# a_114_47# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X43 a_584_47# a_1909_21# Z VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X44 VGND A a_1909_21# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X45 VPWR a_286_367# a_630_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X46 a_630_367# a_1909_21# Z VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X47 Z a_1909_21# a_630_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X48 Z a_1909_21# a_630_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X49 a_114_47# TE_B VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X50 a_584_47# a_114_47# VGND VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X51 Z a_1909_21# a_584_47# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X52 a_1909_21# A VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X53 VPWR a_286_367# a_630_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X54 Z a_1909_21# a_630_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X55 VGND a_114_47# a_584_47# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X56 a_584_47# a_114_47# VGND VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X57 a_1909_21# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X58 VGND a_114_47# a_584_47# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X59 a_584_47# a_1909_21# Z VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X60 a_1909_21# A VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X61 VPWR A a_1909_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X62 VGND a_114_47# a_286_367# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X63 VPWR TE_B a_114_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X64 a_630_367# a_286_367# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X65 a_630_367# a_286_367# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X66 VPWR a_286_367# a_630_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X67 Z a_1909_21# a_630_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X68 Z a_1909_21# a_630_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X69 a_114_47# TE_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X70 VPWR a_114_47# a_286_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X71 Z a_1909_21# a_630_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X72 a_630_367# a_1909_21# Z VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X73 a_630_367# a_1909_21# Z VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X74 a_584_47# a_1909_21# Z VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X75 a_630_367# a_1909_21# Z VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X76 VPWR A a_1909_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X77 Z a_1909_21# a_584_47# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X78 a_584_47# a_1909_21# Z VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X79 a_584_47# a_114_47# VGND VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X80 a_584_47# a_114_47# VGND VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X81 VPWR a_114_47# a_286_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X82 a_630_367# a_286_367# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X83 a_630_367# a_1909_21# Z VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X84 a_286_367# a_114_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X85 Z a_1909_21# a_630_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X86 a_630_367# a_1909_21# Z VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X87 VPWR A a_1909_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X88 a_1909_21# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X89 Z a_1909_21# a_584_47# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
.ends
