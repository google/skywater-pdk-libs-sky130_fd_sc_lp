* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__xnor3_1 A B C VGND VNB VPB VPWR X
M1000 a_354_109# a_754_367# a_871_373# VNB nshort w=640000u l=150000u
+  ad=4.032e+11p pd=3.82e+06u as=5.701e+11p ps=4.79e+06u
M1001 a_355_451# a_754_367# a_1090_373# VNB nshort w=420000u l=150000u
+  ad=4.846e+11p pd=4.15e+06u as=4.173e+11p ps=4.01e+06u
M1002 a_754_367# B VGND VNB nshort w=840000u l=150000u
+  ad=2.394e+11p pd=2.25e+06u as=1.10875e+12p ps=7.97e+06u
M1003 VGND A a_871_373# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_1090_373# B a_354_109# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_1090_373# a_871_373# VPWR VPB phighvt w=1e+06u l=150000u
+  ad=4.642e+11p pd=4.41e+06u as=1.26e+12p ps=9.44e+06u
M1006 a_244_137# C VGND VNB nshort w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=0p ps=0u
M1007 a_871_373# B a_355_451# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_354_109# a_754_367# a_1090_373# VPB phighvt w=640000u l=150000u
+  ad=6.356e+11p pd=4.99e+06u as=0p ps=0u
M1009 a_355_451# a_244_137# a_81_259# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=2.24e+11p ps=1.98e+06u
M1010 a_81_259# C a_354_109# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_81_259# C a_355_451# VPB phighvt w=840000u l=150000u
+  ad=3.612e+11p pd=2.89e+06u as=5.408e+11p ps=4.7e+06u
M1012 a_355_451# a_754_367# a_871_373# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=9.1105e+11p ps=6.07e+06u
M1013 a_871_373# B a_354_109# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_244_137# C VPWR VPB phighvt w=640000u l=150000u
+  ad=1.728e+11p pd=1.82e+06u as=0p ps=0u
M1015 a_1090_373# a_871_373# VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_354_109# a_244_137# a_81_259# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_1090_373# B a_355_451# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VPWR A a_871_373# VPB phighvt w=1e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VGND a_81_259# X VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=2.352e+11p ps=2.24e+06u
M1020 VPWR a_81_259# X VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=3.402e+11p ps=3.06e+06u
M1021 a_754_367# B VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=3.591e+11p pd=3.09e+06u as=0p ps=0u
.ends
