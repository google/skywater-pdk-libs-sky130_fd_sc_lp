* File: sky130_fd_sc_lp__and4b_2.pxi.spice
* Created: Wed Sep  2 09:33:34 2020
* 
x_PM_SKY130_FD_SC_LP__AND4B_2%A_N N_A_N_M1008_g N_A_N_M1012_g N_A_N_c_82_n
+ N_A_N_c_83_n A_N A_N N_A_N_c_85_n N_A_N_c_86_n PM_SKY130_FD_SC_LP__AND4B_2%A_N
x_PM_SKY130_FD_SC_LP__AND4B_2%A_53_375# N_A_53_375#_M1008_d N_A_53_375#_M1012_s
+ N_A_53_375#_M1002_g N_A_53_375#_c_107_n N_A_53_375#_M1001_g
+ N_A_53_375#_c_108_n N_A_53_375#_c_109_n N_A_53_375#_c_110_n
+ N_A_53_375#_c_111_n N_A_53_375#_c_116_n N_A_53_375#_c_112_n
+ N_A_53_375#_c_113_n N_A_53_375#_c_114_n PM_SKY130_FD_SC_LP__AND4B_2%A_53_375#
x_PM_SKY130_FD_SC_LP__AND4B_2%B N_B_M1009_g N_B_M1010_g B B N_B_c_157_n
+ PM_SKY130_FD_SC_LP__AND4B_2%B
x_PM_SKY130_FD_SC_LP__AND4B_2%C N_C_M1011_g N_C_M1005_g C C N_C_c_188_n
+ PM_SKY130_FD_SC_LP__AND4B_2%C
x_PM_SKY130_FD_SC_LP__AND4B_2%D N_D_M1013_g N_D_M1003_g D N_D_c_220_n
+ N_D_c_221_n PM_SKY130_FD_SC_LP__AND4B_2%D
x_PM_SKY130_FD_SC_LP__AND4B_2%A_222_375# N_A_222_375#_M1001_s
+ N_A_222_375#_M1002_d N_A_222_375#_M1005_d N_A_222_375#_M1004_g
+ N_A_222_375#_M1000_g N_A_222_375#_M1007_g N_A_222_375#_M1006_g
+ N_A_222_375#_c_256_n N_A_222_375#_c_257_n N_A_222_375#_c_278_n
+ N_A_222_375#_c_290_n N_A_222_375#_c_265_n N_A_222_375#_c_266_n
+ N_A_222_375#_c_258_n N_A_222_375#_c_259_n N_A_222_375#_c_260_n
+ N_A_222_375#_c_261_n PM_SKY130_FD_SC_LP__AND4B_2%A_222_375#
x_PM_SKY130_FD_SC_LP__AND4B_2%VPWR N_VPWR_M1012_d N_VPWR_M1009_d N_VPWR_M1003_d
+ N_VPWR_M1006_d N_VPWR_c_357_n N_VPWR_c_358_n N_VPWR_c_359_n N_VPWR_c_360_n
+ N_VPWR_c_361_n N_VPWR_c_362_n VPWR N_VPWR_c_363_n N_VPWR_c_364_n
+ N_VPWR_c_365_n N_VPWR_c_366_n N_VPWR_c_367_n N_VPWR_c_368_n N_VPWR_c_356_n
+ PM_SKY130_FD_SC_LP__AND4B_2%VPWR
x_PM_SKY130_FD_SC_LP__AND4B_2%X N_X_M1004_s N_X_M1000_s N_X_c_402_n N_X_c_403_n
+ N_X_c_400_n N_X_c_401_n X X X PM_SKY130_FD_SC_LP__AND4B_2%X
x_PM_SKY130_FD_SC_LP__AND4B_2%VGND N_VGND_M1008_s N_VGND_M1013_d N_VGND_M1007_d
+ N_VGND_c_428_n N_VGND_c_429_n N_VGND_c_430_n N_VGND_c_431_n N_VGND_c_432_n
+ N_VGND_c_433_n N_VGND_c_434_n VGND N_VGND_c_435_n N_VGND_c_436_n
+ N_VGND_c_437_n N_VGND_c_438_n PM_SKY130_FD_SC_LP__AND4B_2%VGND
cc_1 VNB N_A_N_M1012_g 0.0129058f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=2.085
cc_2 VNB N_A_N_c_82_n 0.0296608f $X=-0.19 $Y=-0.245 $X2=0.417 $Y2=1.335
cc_3 VNB N_A_N_c_83_n 0.0300707f $X=-0.19 $Y=-0.245 $X2=0.417 $Y2=1.485
cc_4 VNB A_N 0.0356094f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_5 VNB N_A_N_c_85_n 0.0251095f $X=-0.19 $Y=-0.245 $X2=0.32 $Y2=0.98
cc_6 VNB N_A_N_c_86_n 0.0226592f $X=-0.19 $Y=-0.245 $X2=0.352 $Y2=0.815
cc_7 VNB N_A_53_375#_M1002_g 0.02193f $X=-0.19 $Y=-0.245 $X2=0.417 $Y2=1.485
cc_8 VNB N_A_53_375#_c_107_n 0.0142692f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_9 VNB N_A_53_375#_c_108_n 0.0156001f $X=-0.19 $Y=-0.245 $X2=0.352 $Y2=0.98
cc_10 VNB N_A_53_375#_c_109_n 0.0332628f $X=-0.19 $Y=-0.245 $X2=0.32 $Y2=0.98
cc_11 VNB N_A_53_375#_c_110_n 0.0162387f $X=-0.19 $Y=-0.245 $X2=0.32 $Y2=0.98
cc_12 VNB N_A_53_375#_c_111_n 0.0541903f $X=-0.19 $Y=-0.245 $X2=0.352 $Y2=0.815
cc_13 VNB N_A_53_375#_c_112_n 0.00173877f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_53_375#_c_113_n 0.0142689f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_53_375#_c_114_n 0.00654796f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_B_M1010_g 0.0289646f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=2.085
cc_17 VNB B 0.00288003f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_B_c_157_n 0.0314547f $X=-0.19 $Y=-0.245 $X2=0.32 $Y2=0.98
cc_19 VNB N_C_M1011_g 0.0205068f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.815
cc_20 VNB N_C_M1005_g 0.00615862f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=2.085
cc_21 VNB C 0.00500475f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_C_c_188_n 0.0304695f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_D_M1013_g 0.0227114f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.815
cc_24 VNB N_D_M1003_g 0.00669635f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=2.085
cc_25 VNB N_D_c_220_n 0.029769f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_26 VNB N_D_c_221_n 0.00554982f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_27 VNB N_A_222_375#_M1004_g 0.019328f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_28 VNB N_A_222_375#_M1000_g 0.00628238f $X=-0.19 $Y=-0.245 $X2=0.352 $Y2=0.98
cc_29 VNB N_A_222_375#_M1007_g 0.0230058f $X=-0.19 $Y=-0.245 $X2=0.255 $Y2=0.925
cc_30 VNB N_A_222_375#_M1006_g 0.00869743f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_222_375#_c_256_n 0.00264988f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_222_375#_c_257_n 0.00723086f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_222_375#_c_258_n 0.00158873f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_222_375#_c_259_n 0.00226986f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_222_375#_c_260_n 0.00259297f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_222_375#_c_261_n 0.0574066f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VPWR_c_356_n 0.183584f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_X_c_400_n 0.00186216f $X=-0.19 $Y=-0.245 $X2=0.352 $Y2=0.98
cc_39 VNB N_VGND_c_428_n 0.0107448f $X=-0.19 $Y=-0.245 $X2=0.417 $Y2=1.335
cc_40 VNB N_VGND_c_429_n 0.0196254f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_41 VNB N_VGND_c_430_n 0.0140752f $X=-0.19 $Y=-0.245 $X2=0.352 $Y2=0.98
cc_42 VNB N_VGND_c_431_n 0.0131423f $X=-0.19 $Y=-0.245 $X2=0.32 $Y2=0.98
cc_43 VNB N_VGND_c_432_n 0.0154922f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_433_n 0.0255047f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_434_n 0.0072588f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_435_n 0.0718813f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_436_n 0.0152106f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_437_n 0.00510987f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_438_n 0.250483f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VPB N_A_N_M1012_g 0.0310067f $X=-0.19 $Y=1.655 $X2=0.605 $Y2=2.085
cc_51 VPB N_A_53_375#_M1002_g 0.0256887f $X=-0.19 $Y=1.655 $X2=0.417 $Y2=1.485
cc_52 VPB N_A_53_375#_c_116_n 0.0165579f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_53 VPB N_A_53_375#_c_113_n 0.0157935f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_54 VPB N_B_M1009_g 0.0268444f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.815
cc_55 VPB B 0.00285762f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_56 VPB N_B_c_157_n 0.016072f $X=-0.19 $Y=1.655 $X2=0.32 $Y2=0.98
cc_57 VPB N_C_M1005_g 0.0320469f $X=-0.19 $Y=1.655 $X2=0.605 $Y2=2.085
cc_58 VPB C 0.00326249f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_59 VPB N_D_M1003_g 0.0256484f $X=-0.19 $Y=1.655 $X2=0.605 $Y2=2.085
cc_60 VPB N_A_222_375#_M1000_g 0.0223652f $X=-0.19 $Y=1.655 $X2=0.352 $Y2=0.98
cc_61 VPB N_A_222_375#_M1006_g 0.0264962f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_62 VPB N_A_222_375#_c_257_n 0.00209297f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_63 VPB N_A_222_375#_c_265_n 0.00576678f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_64 VPB N_A_222_375#_c_266_n 0.00340963f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_65 VPB N_A_222_375#_c_259_n 9.97414e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_357_n 0.0450259f $X=-0.19 $Y=1.655 $X2=0.32 $Y2=0.98
cc_67 VPB N_VPWR_c_358_n 0.0452979f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_359_n 0.0142562f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_69 VPB N_VPWR_c_360_n 0.0253235f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_70 VPB N_VPWR_c_361_n 0.0120619f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_71 VPB N_VPWR_c_362_n 0.0388188f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_72 VPB N_VPWR_c_363_n 0.0187113f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_73 VPB N_VPWR_c_364_n 0.018234f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_74 VPB N_VPWR_c_365_n 0.0152484f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_75 VPB N_VPWR_c_366_n 0.0293083f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_76 VPB N_VPWR_c_367_n 0.0140155f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_77 VPB N_VPWR_c_368_n 0.00693572f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_78 VPB N_VPWR_c_356_n 0.115938f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_79 VPB N_X_c_401_n 0.00240734f $X=-0.19 $Y=1.655 $X2=0.32 $Y2=0.98
cc_80 N_A_N_c_82_n N_A_53_375#_M1002_g 0.00138629f $X=0.417 $Y=1.335 $X2=0 $Y2=0
cc_81 N_A_N_c_83_n N_A_53_375#_M1002_g 0.0309327f $X=0.417 $Y=1.485 $X2=0 $Y2=0
cc_82 N_A_N_c_86_n N_A_53_375#_c_108_n 0.00902153f $X=0.352 $Y=0.815 $X2=0 $Y2=0
cc_83 N_A_N_c_85_n N_A_53_375#_c_109_n 0.00902153f $X=0.32 $Y=0.98 $X2=0 $Y2=0
cc_84 N_A_N_c_82_n N_A_53_375#_c_110_n 0.00902153f $X=0.417 $Y=1.335 $X2=0 $Y2=0
cc_85 N_A_N_M1012_g N_A_53_375#_c_116_n 6.72223e-19 $X=0.605 $Y=2.085 $X2=0
+ $Y2=0
cc_86 N_A_N_c_86_n N_A_53_375#_c_112_n 3.41499e-19 $X=0.352 $Y=0.815 $X2=0 $Y2=0
cc_87 N_A_N_M1012_g N_A_53_375#_c_113_n 0.0267521f $X=0.605 $Y=2.085 $X2=0 $Y2=0
cc_88 N_A_N_c_83_n N_A_53_375#_c_113_n 0.0118795f $X=0.417 $Y=1.485 $X2=0 $Y2=0
cc_89 A_N N_A_53_375#_c_113_n 0.0639814f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_90 N_A_N_c_86_n N_A_53_375#_c_113_n 0.00776673f $X=0.352 $Y=0.815 $X2=0 $Y2=0
cc_91 N_A_N_M1012_g N_VPWR_c_357_n 0.0123844f $X=0.605 $Y=2.085 $X2=0 $Y2=0
cc_92 A_N N_VGND_c_429_n 0.0255463f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_93 N_A_N_c_85_n N_VGND_c_429_n 0.00174534f $X=0.32 $Y=0.98 $X2=0 $Y2=0
cc_94 N_A_N_c_86_n N_VGND_c_429_n 0.00980982f $X=0.352 $Y=0.815 $X2=0 $Y2=0
cc_95 N_A_N_c_86_n N_VGND_c_435_n 0.00445056f $X=0.352 $Y=0.815 $X2=0 $Y2=0
cc_96 A_N N_VGND_c_438_n 0.00154298f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_97 N_A_N_c_86_n N_VGND_c_438_n 0.00847361f $X=0.352 $Y=0.815 $X2=0 $Y2=0
cc_98 N_A_53_375#_c_110_n N_B_M1010_g 0.0023063f $X=1 $Y=1.27 $X2=0 $Y2=0
cc_99 N_A_53_375#_c_111_n N_B_M1010_g 0.0435326f $X=1.38 $Y=0.35 $X2=0 $Y2=0
cc_100 N_A_53_375#_M1002_g N_B_c_157_n 0.0261935f $X=1.035 $Y=2.085 $X2=0 $Y2=0
cc_101 N_A_53_375#_c_107_n N_B_c_157_n 0.0107831f $X=1.455 $Y=0.515 $X2=0 $Y2=0
cc_102 N_A_53_375#_c_107_n N_A_222_375#_c_256_n 0.00109708f $X=1.455 $Y=0.515
+ $X2=0 $Y2=0
cc_103 N_A_53_375#_c_109_n N_A_222_375#_c_256_n 0.00241716f $X=1 $Y=1.12 $X2=0
+ $Y2=0
cc_104 N_A_53_375#_c_110_n N_A_222_375#_c_256_n 0.00157744f $X=1 $Y=1.27 $X2=0
+ $Y2=0
cc_105 N_A_53_375#_c_111_n N_A_222_375#_c_256_n 0.00216885f $X=1.38 $Y=0.35
+ $X2=0 $Y2=0
cc_106 N_A_53_375#_c_113_n N_A_222_375#_c_256_n 0.0126329f $X=0.695 $Y=1.695
+ $X2=0 $Y2=0
cc_107 N_A_53_375#_c_114_n N_A_222_375#_c_256_n 0.0128503f $X=1.09 $Y=0.35 $X2=0
+ $Y2=0
cc_108 N_A_53_375#_c_107_n N_A_222_375#_c_257_n 0.00448534f $X=1.455 $Y=0.515
+ $X2=0 $Y2=0
cc_109 N_A_53_375#_c_109_n N_A_222_375#_c_257_n 0.00109923f $X=1 $Y=1.12 $X2=0
+ $Y2=0
cc_110 N_A_53_375#_c_110_n N_A_222_375#_c_257_n 0.00894471f $X=1 $Y=1.27 $X2=0
+ $Y2=0
cc_111 N_A_53_375#_c_113_n N_A_222_375#_c_257_n 0.0405425f $X=0.695 $Y=1.695
+ $X2=0 $Y2=0
cc_112 N_A_53_375#_c_107_n N_A_222_375#_c_278_n 0.00899459f $X=1.455 $Y=0.515
+ $X2=0 $Y2=0
cc_113 N_A_53_375#_M1002_g N_VPWR_c_357_n 0.00870678f $X=1.035 $Y=2.085 $X2=0
+ $Y2=0
cc_114 N_A_53_375#_c_113_n N_VPWR_c_357_n 0.00869932f $X=0.695 $Y=1.695 $X2=0
+ $Y2=0
cc_115 N_A_53_375#_c_108_n N_VGND_c_429_n 7.37936e-19 $X=1.04 $Y=0.35 $X2=0
+ $Y2=0
cc_116 N_A_53_375#_c_112_n N_VGND_c_429_n 0.0141643f $X=0.695 $Y=0.595 $X2=0
+ $Y2=0
cc_117 N_A_53_375#_c_108_n N_VGND_c_435_n 0.0165132f $X=1.04 $Y=0.35 $X2=0 $Y2=0
cc_118 N_A_53_375#_c_112_n N_VGND_c_435_n 0.0143373f $X=0.695 $Y=0.595 $X2=0
+ $Y2=0
cc_119 N_A_53_375#_c_114_n N_VGND_c_435_n 0.0298901f $X=1.09 $Y=0.35 $X2=0 $Y2=0
cc_120 N_A_53_375#_c_108_n N_VGND_c_438_n 0.00424196f $X=1.04 $Y=0.35 $X2=0
+ $Y2=0
cc_121 N_A_53_375#_c_111_n N_VGND_c_438_n 0.0149418f $X=1.38 $Y=0.35 $X2=0 $Y2=0
cc_122 N_A_53_375#_c_112_n N_VGND_c_438_n 0.00777554f $X=0.695 $Y=0.595 $X2=0
+ $Y2=0
cc_123 N_A_53_375#_c_114_n N_VGND_c_438_n 0.0158597f $X=1.09 $Y=0.35 $X2=0 $Y2=0
cc_124 N_B_M1010_g N_C_M1011_g 0.0332006f $X=1.815 $Y=0.835 $X2=0 $Y2=0
cc_125 B N_C_M1005_g 2.81182e-19 $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_126 N_B_c_157_n N_C_M1005_g 0.00477613f $X=1.815 $Y=1.55 $X2=0 $Y2=0
cc_127 N_B_M1010_g C 0.0040857f $X=1.815 $Y=0.835 $X2=0 $Y2=0
cc_128 B C 0.0422608f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_129 B N_C_c_188_n 3.13252e-19 $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_130 N_B_c_157_n N_C_c_188_n 0.0332006f $X=1.815 $Y=1.55 $X2=0 $Y2=0
cc_131 N_B_M1009_g N_A_222_375#_c_257_n 0.0128493f $X=1.465 $Y=2.085 $X2=0 $Y2=0
cc_132 N_B_M1010_g N_A_222_375#_c_257_n 0.00171105f $X=1.815 $Y=0.835 $X2=0
+ $Y2=0
cc_133 B N_A_222_375#_c_257_n 0.0404451f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_134 N_B_c_157_n N_A_222_375#_c_257_n 0.00815137f $X=1.815 $Y=1.55 $X2=0 $Y2=0
cc_135 N_B_M1010_g N_A_222_375#_c_278_n 0.0138514f $X=1.815 $Y=0.835 $X2=0 $Y2=0
cc_136 B N_A_222_375#_c_278_n 0.0157529f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_137 N_B_c_157_n N_A_222_375#_c_278_n 0.0013115f $X=1.815 $Y=1.55 $X2=0 $Y2=0
cc_138 N_B_M1009_g N_VPWR_c_357_n 4.63085e-19 $X=1.465 $Y=2.085 $X2=0 $Y2=0
cc_139 N_B_M1009_g N_VPWR_c_358_n 0.00433917f $X=1.465 $Y=2.085 $X2=0 $Y2=0
cc_140 B N_VPWR_c_358_n 0.0223591f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_141 N_B_c_157_n N_VPWR_c_358_n 0.00439771f $X=1.815 $Y=1.55 $X2=0 $Y2=0
cc_142 N_B_M1010_g N_VGND_c_435_n 0.00415323f $X=1.815 $Y=0.835 $X2=0 $Y2=0
cc_143 N_B_M1010_g N_VGND_c_438_n 0.00469432f $X=1.815 $Y=0.835 $X2=0 $Y2=0
cc_144 N_C_M1011_g N_D_M1013_g 0.0241861f $X=2.175 $Y=0.835 $X2=0 $Y2=0
cc_145 N_C_M1005_g N_D_M1003_g 0.0166827f $X=2.355 $Y=2.085 $X2=0 $Y2=0
cc_146 C N_D_M1003_g 9.10382e-19 $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_147 C N_D_c_220_n 2.86533e-19 $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_148 N_C_c_188_n N_D_c_220_n 0.0204371f $X=2.265 $Y=1.375 $X2=0 $Y2=0
cc_149 C N_D_c_221_n 0.029364f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_150 N_C_c_188_n N_D_c_221_n 0.00220692f $X=2.265 $Y=1.375 $X2=0 $Y2=0
cc_151 C N_A_222_375#_c_257_n 0.00117965f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_152 N_C_M1011_g N_A_222_375#_c_278_n 0.0132157f $X=2.175 $Y=0.835 $X2=0 $Y2=0
cc_153 C N_A_222_375#_c_278_n 0.0231899f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_154 N_C_c_188_n N_A_222_375#_c_278_n 0.00381993f $X=2.265 $Y=1.375 $X2=0
+ $Y2=0
cc_155 N_C_M1005_g N_A_222_375#_c_290_n 0.00188396f $X=2.355 $Y=2.085 $X2=0
+ $Y2=0
cc_156 N_C_M1005_g N_A_222_375#_c_266_n 0.00433484f $X=2.355 $Y=2.085 $X2=0
+ $Y2=0
cc_157 C N_A_222_375#_c_266_n 0.00339935f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_158 N_C_M1005_g N_VPWR_c_358_n 0.0113297f $X=2.355 $Y=2.085 $X2=0 $Y2=0
cc_159 C N_VPWR_c_358_n 0.0242631f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_160 N_C_c_188_n N_VPWR_c_358_n 7.56645e-19 $X=2.265 $Y=1.375 $X2=0 $Y2=0
cc_161 N_C_M1005_g N_VPWR_c_359_n 5.11579e-19 $X=2.355 $Y=2.085 $X2=0 $Y2=0
cc_162 N_C_M1011_g N_VGND_c_435_n 0.00415323f $X=2.175 $Y=0.835 $X2=0 $Y2=0
cc_163 N_C_M1011_g N_VGND_c_438_n 0.00469432f $X=2.175 $Y=0.835 $X2=0 $Y2=0
cc_164 N_D_M1013_g N_A_222_375#_M1004_g 0.0152164f $X=2.715 $Y=0.835 $X2=0 $Y2=0
cc_165 N_D_M1003_g N_A_222_375#_M1000_g 0.0184408f $X=2.83 $Y=2.085 $X2=0 $Y2=0
cc_166 N_D_M1013_g N_A_222_375#_c_278_n 0.0146712f $X=2.715 $Y=0.835 $X2=0 $Y2=0
cc_167 N_D_c_220_n N_A_222_375#_c_278_n 0.0035369f $X=2.805 $Y=1.375 $X2=0 $Y2=0
cc_168 N_D_c_221_n N_A_222_375#_c_278_n 0.0242411f $X=2.805 $Y=1.375 $X2=0 $Y2=0
cc_169 N_D_M1003_g N_A_222_375#_c_265_n 0.0143844f $X=2.83 $Y=2.085 $X2=0 $Y2=0
cc_170 N_D_c_220_n N_A_222_375#_c_265_n 0.00362584f $X=2.805 $Y=1.375 $X2=0
+ $Y2=0
cc_171 N_D_c_221_n N_A_222_375#_c_265_n 0.0130901f $X=2.805 $Y=1.375 $X2=0 $Y2=0
cc_172 N_D_c_220_n N_A_222_375#_c_266_n 0.00189343f $X=2.805 $Y=1.375 $X2=0
+ $Y2=0
cc_173 N_D_c_221_n N_A_222_375#_c_266_n 0.0163381f $X=2.805 $Y=1.375 $X2=0 $Y2=0
cc_174 N_D_M1013_g N_A_222_375#_c_258_n 0.00338389f $X=2.715 $Y=0.835 $X2=0
+ $Y2=0
cc_175 N_D_c_221_n N_A_222_375#_c_258_n 0.00262394f $X=2.805 $Y=1.375 $X2=0
+ $Y2=0
cc_176 N_D_M1003_g N_A_222_375#_c_259_n 0.00368269f $X=2.83 $Y=2.085 $X2=0 $Y2=0
cc_177 N_D_c_220_n N_A_222_375#_c_260_n 0.00219699f $X=2.805 $Y=1.375 $X2=0
+ $Y2=0
cc_178 N_D_c_221_n N_A_222_375#_c_260_n 0.0254789f $X=2.805 $Y=1.375 $X2=0 $Y2=0
cc_179 N_D_c_220_n N_A_222_375#_c_261_n 0.0205522f $X=2.805 $Y=1.375 $X2=0 $Y2=0
cc_180 N_D_c_221_n N_A_222_375#_c_261_n 2.89895e-19 $X=2.805 $Y=1.375 $X2=0
+ $Y2=0
cc_181 N_D_M1003_g N_VPWR_c_358_n 5.61107e-19 $X=2.83 $Y=2.085 $X2=0 $Y2=0
cc_182 N_D_M1003_g N_VPWR_c_359_n 0.00809429f $X=2.83 $Y=2.085 $X2=0 $Y2=0
cc_183 N_D_M1013_g N_VGND_c_430_n 0.00345938f $X=2.715 $Y=0.835 $X2=0 $Y2=0
cc_184 N_D_M1013_g N_VGND_c_435_n 0.00415323f $X=2.715 $Y=0.835 $X2=0 $Y2=0
cc_185 N_D_M1013_g N_VGND_c_438_n 0.00469432f $X=2.715 $Y=0.835 $X2=0 $Y2=0
cc_186 N_A_222_375#_c_265_n N_VPWR_M1003_d 0.00305996f $X=3.07 $Y=1.795 $X2=0
+ $Y2=0
cc_187 N_A_222_375#_c_290_n N_VPWR_c_358_n 0.0217079f $X=2.615 $Y=2.085 $X2=0
+ $Y2=0
cc_188 N_A_222_375#_M1000_g N_VPWR_c_359_n 0.021032f $X=3.355 $Y=2.465 $X2=0
+ $Y2=0
cc_189 N_A_222_375#_M1006_g N_VPWR_c_359_n 7.64614e-19 $X=3.785 $Y=2.465 $X2=0
+ $Y2=0
cc_190 N_A_222_375#_c_265_n N_VPWR_c_359_n 0.0236616f $X=3.07 $Y=1.795 $X2=0
+ $Y2=0
cc_191 N_A_222_375#_c_260_n N_VPWR_c_359_n 0.00142686f $X=3.345 $Y=1.375 $X2=0
+ $Y2=0
cc_192 N_A_222_375#_c_261_n N_VPWR_c_359_n 2.00935e-19 $X=3.785 $Y=1.375 $X2=0
+ $Y2=0
cc_193 N_A_222_375#_M1006_g N_VPWR_c_360_n 0.00123232f $X=3.785 $Y=2.465 $X2=0
+ $Y2=0
cc_194 N_A_222_375#_M1006_g N_VPWR_c_362_n 0.00644397f $X=3.785 $Y=2.465 $X2=0
+ $Y2=0
cc_195 N_A_222_375#_M1000_g N_VPWR_c_365_n 0.00486043f $X=3.355 $Y=2.465 $X2=0
+ $Y2=0
cc_196 N_A_222_375#_M1006_g N_VPWR_c_365_n 0.00585385f $X=3.785 $Y=2.465 $X2=0
+ $Y2=0
cc_197 N_A_222_375#_M1000_g N_VPWR_c_356_n 0.00824727f $X=3.355 $Y=2.465 $X2=0
+ $Y2=0
cc_198 N_A_222_375#_M1006_g N_VPWR_c_356_n 0.011548f $X=3.785 $Y=2.465 $X2=0
+ $Y2=0
cc_199 N_A_222_375#_M1007_g N_X_c_402_n 0.00717014f $X=3.72 $Y=0.655 $X2=0 $Y2=0
cc_200 N_A_222_375#_M1007_g N_X_c_403_n 0.00661708f $X=3.72 $Y=0.655 $X2=0 $Y2=0
cc_201 N_A_222_375#_c_260_n N_X_c_403_n 0.00107537f $X=3.345 $Y=1.375 $X2=0
+ $Y2=0
cc_202 N_A_222_375#_c_261_n N_X_c_403_n 0.00357268f $X=3.785 $Y=1.375 $X2=0
+ $Y2=0
cc_203 N_A_222_375#_M1004_g N_X_c_400_n 8.12475e-19 $X=3.29 $Y=0.655 $X2=0 $Y2=0
cc_204 N_A_222_375#_M1000_g N_X_c_400_n 9.1981e-19 $X=3.355 $Y=2.465 $X2=0 $Y2=0
cc_205 N_A_222_375#_M1007_g N_X_c_400_n 0.00748758f $X=3.72 $Y=0.655 $X2=0 $Y2=0
cc_206 N_A_222_375#_M1006_g N_X_c_400_n 0.00909433f $X=3.785 $Y=2.465 $X2=0
+ $Y2=0
cc_207 N_A_222_375#_c_258_n N_X_c_400_n 0.00491548f $X=3.155 $Y=1.21 $X2=0 $Y2=0
cc_208 N_A_222_375#_c_259_n N_X_c_400_n 0.00538246f $X=3.155 $Y=1.71 $X2=0 $Y2=0
cc_209 N_A_222_375#_c_260_n N_X_c_400_n 0.0238097f $X=3.345 $Y=1.375 $X2=0 $Y2=0
cc_210 N_A_222_375#_c_261_n N_X_c_400_n 0.0228345f $X=3.785 $Y=1.375 $X2=0 $Y2=0
cc_211 N_A_222_375#_M1000_g N_X_c_401_n 0.00156857f $X=3.355 $Y=2.465 $X2=0
+ $Y2=0
cc_212 N_A_222_375#_M1006_g N_X_c_401_n 0.0104693f $X=3.785 $Y=2.465 $X2=0 $Y2=0
cc_213 N_A_222_375#_c_265_n N_X_c_401_n 0.00871733f $X=3.07 $Y=1.795 $X2=0 $Y2=0
cc_214 N_A_222_375#_c_261_n N_X_c_401_n 0.00259069f $X=3.785 $Y=1.375 $X2=0
+ $Y2=0
cc_215 N_A_222_375#_c_278_n N_VGND_M1013_d 0.00982834f $X=3.07 $Y=0.9 $X2=0
+ $Y2=0
cc_216 N_A_222_375#_c_258_n N_VGND_M1013_d 8.71942e-19 $X=3.155 $Y=1.21 $X2=0
+ $Y2=0
cc_217 N_A_222_375#_M1004_g N_VGND_c_430_n 0.0106944f $X=3.29 $Y=0.655 $X2=0
+ $Y2=0
cc_218 N_A_222_375#_M1007_g N_VGND_c_430_n 5.83321e-19 $X=3.72 $Y=0.655 $X2=0
+ $Y2=0
cc_219 N_A_222_375#_c_278_n N_VGND_c_430_n 0.0221262f $X=3.07 $Y=0.9 $X2=0 $Y2=0
cc_220 N_A_222_375#_M1007_g N_VGND_c_432_n 0.00553513f $X=3.72 $Y=0.655 $X2=0
+ $Y2=0
cc_221 N_A_222_375#_M1007_g N_VGND_c_433_n 0.00821263f $X=3.72 $Y=0.655 $X2=0
+ $Y2=0
cc_222 N_A_222_375#_c_261_n N_VGND_c_434_n 6.20567e-19 $X=3.785 $Y=1.375 $X2=0
+ $Y2=0
cc_223 N_A_222_375#_M1004_g N_VGND_c_436_n 0.00486043f $X=3.29 $Y=0.655 $X2=0
+ $Y2=0
cc_224 N_A_222_375#_M1007_g N_VGND_c_436_n 0.00564131f $X=3.72 $Y=0.655 $X2=0
+ $Y2=0
cc_225 N_A_222_375#_M1004_g N_VGND_c_438_n 0.00824727f $X=3.29 $Y=0.655 $X2=0
+ $Y2=0
cc_226 N_A_222_375#_M1007_g N_VGND_c_438_n 0.00760335f $X=3.72 $Y=0.655 $X2=0
+ $Y2=0
cc_227 N_A_222_375#_c_256_n N_VGND_c_438_n 0.00580461f $X=1.28 $Y=1.005 $X2=0
+ $Y2=0
cc_228 N_A_222_375#_c_278_n N_VGND_c_438_n 0.0538467f $X=3.07 $Y=0.9 $X2=0 $Y2=0
cc_229 N_A_222_375#_c_278_n A_306_125# 0.00284626f $X=3.07 $Y=0.9 $X2=-0.19
+ $Y2=-0.245
cc_230 N_A_222_375#_c_278_n A_378_125# 0.0046088f $X=3.07 $Y=0.9 $X2=-0.19
+ $Y2=-0.245
cc_231 N_A_222_375#_c_278_n A_450_125# 0.0113618f $X=3.07 $Y=0.9 $X2=-0.19
+ $Y2=-0.245
cc_232 N_VPWR_c_356_n N_X_M1000_s 0.0041489f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_233 N_VPWR_c_360_n N_X_c_401_n 0.00496438f $X=4.042 $Y=2.207 $X2=0 $Y2=0
cc_234 N_VPWR_c_365_n X 0.0136943f $X=3.885 $Y=3.33 $X2=0 $Y2=0
cc_235 N_VPWR_c_356_n X 0.00866972f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_236 N_X_c_402_n N_VGND_c_433_n 0.00835387f $X=3.505 $Y=0.42 $X2=0 $Y2=0
cc_237 N_X_c_403_n N_VGND_c_433_n 0.0181686f $X=3.595 $Y=1.04 $X2=0 $Y2=0
cc_238 N_X_c_402_n N_VGND_c_436_n 0.0150063f $X=3.505 $Y=0.42 $X2=0 $Y2=0
cc_239 N_X_M1004_s N_VGND_c_438_n 0.00380103f $X=3.365 $Y=0.235 $X2=0 $Y2=0
cc_240 N_X_c_402_n N_VGND_c_438_n 0.00950443f $X=3.505 $Y=0.42 $X2=0 $Y2=0
cc_241 N_X_c_403_n N_VGND_c_438_n 0.00369804f $X=3.595 $Y=1.04 $X2=0 $Y2=0
