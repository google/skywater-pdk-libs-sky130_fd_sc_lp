* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__dlxtp_lp2 D GATE VGND VNB VPB VPWR Q
X0 VPWR GATE a_240_409# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X1 VPWR a_778_47# a_928_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X2 a_452_419# a_240_409# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X3 a_972_419# a_928_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X4 VPWR a_27_57# a_766_419# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X5 a_778_47# a_452_419# a_972_419# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X6 VGND a_928_21# a_1477_83# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 a_1207_47# a_778_47# a_928_21# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 a_766_419# a_240_409# a_778_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X9 a_27_57# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X10 a_880_47# a_928_21# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X11 a_272_57# GATE a_240_409# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 a_778_47# a_240_409# a_880_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X13 a_452_419# a_240_409# a_542_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X14 a_700_47# a_452_419# a_778_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X15 VGND a_778_47# a_1207_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X16 a_542_47# a_240_409# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X17 a_114_57# D VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X18 a_27_57# D a_114_57# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X19 VGND GATE a_272_57# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X20 VGND a_27_57# a_700_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X21 VPWR a_928_21# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X22 a_1477_83# a_928_21# Q VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
