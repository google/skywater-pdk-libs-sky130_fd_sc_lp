* NGSPICE file created from sky130_fd_sc_lp__xor3_lp.ext - technology: sky130A

.subckt sky130_fd_sc_lp__xor3_lp A B C VGND VNB VPB VPWR X
M1000 a_430_113# a_57_113# VGND VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=6.825e+11p ps=5.77e+06u
M1001 VGND C a_1860_141# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1002 a_144_113# A a_57_113# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=3.22525e+11p ps=3.56e+06u
M1003 a_388_419# a_57_113# VPWR VPB phighvt w=1e+06u l=250000u
+  ad=5.65e+11p pd=5.13e+06u as=1.785e+12p ps=9.57e+06u
M1004 X a_1459_406# a_2046_141# VNB nshort w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=1.008e+11p ps=1.32e+06u
M1005 a_1459_406# C a_494_419# VNB nshort w=420000u l=150000u
+  ad=1.302e+11p pd=1.46e+06u as=3.954e+11p ps=3.6e+06u
M1006 a_57_113# B a_494_419# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_388_419# a_580_21# a_855_66# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=5.75e+11p ps=5.15e+06u
M1008 a_1860_141# C a_1393_300# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.659e+11p ps=1.63e+06u
M1009 a_494_419# a_580_21# a_388_419# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=2.709e+11p ps=2.97e+06u
M1010 VGND B a_1245_89# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1011 a_2046_141# a_1459_406# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_855_66# C a_1459_406# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=2.8e+11p ps=2.56e+06u
M1013 a_388_419# a_57_113# a_430_113# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VPWR B a_580_21# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=3.75e+11p ps=2.75e+06u
M1015 a_1245_89# B a_580_21# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1016 a_388_419# B a_855_66# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=4.1495e+11p ps=3.82e+06u
M1017 a_494_419# B a_388_419# VPB phighvt w=1e+06u l=250000u
+  ad=1.1e+12p pd=6.2e+06u as=0p ps=0u
M1018 a_855_66# a_580_21# a_57_113# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_57_113# a_580_21# a_494_419# VPB phighvt w=1e+06u l=250000u
+  ad=9.05e+11p pd=5.81e+06u as=0p ps=0u
M1020 a_855_66# B a_57_113# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1021 X a_1459_406# VPWR VPB phighvt w=1e+06u l=250000u
+  ad=2.85e+11p pd=2.57e+06u as=0p ps=0u
M1022 a_855_66# a_1393_300# a_1459_406# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 VPWR A a_57_113# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_1459_406# a_1393_300# a_494_419# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1025 VGND A a_144_113# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 VPWR C a_1393_300# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=2.85e+11p ps=2.57e+06u
.ends

