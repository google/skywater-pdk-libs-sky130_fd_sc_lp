* File: sky130_fd_sc_lp__a22o_1.pxi.spice
* Created: Wed Sep  2 09:22:27 2020
* 
x_PM_SKY130_FD_SC_LP__A22O_1%A_80_246# N_A_80_246#_M1004_d N_A_80_246#_M1002_d
+ N_A_80_246#_M1009_g N_A_80_246#_c_57_n N_A_80_246#_M1006_g N_A_80_246#_c_58_n
+ N_A_80_246#_c_59_n N_A_80_246#_c_67_p N_A_80_246#_c_112_p N_A_80_246#_c_60_n
+ N_A_80_246#_c_64_n N_A_80_246#_c_70_p N_A_80_246#_c_82_p N_A_80_246#_c_61_n
+ PM_SKY130_FD_SC_LP__A22O_1%A_80_246#
x_PM_SKY130_FD_SC_LP__A22O_1%B2 N_B2_c_123_n N_B2_M1003_g N_B2_M1002_g B2
+ N_B2_c_126_n PM_SKY130_FD_SC_LP__A22O_1%B2
x_PM_SKY130_FD_SC_LP__A22O_1%B1 N_B1_M1004_g N_B1_M1005_g B1 N_B1_c_157_n
+ N_B1_c_158_n N_B1_c_159_n PM_SKY130_FD_SC_LP__A22O_1%B1
x_PM_SKY130_FD_SC_LP__A22O_1%A1 N_A1_M1007_g N_A1_M1008_g A1 A1 A1 N_A1_c_195_n
+ N_A1_c_196_n PM_SKY130_FD_SC_LP__A22O_1%A1
x_PM_SKY130_FD_SC_LP__A22O_1%A2 N_A2_M1001_g N_A2_M1000_g A2 N_A2_c_232_n
+ N_A2_c_233_n PM_SKY130_FD_SC_LP__A22O_1%A2
x_PM_SKY130_FD_SC_LP__A22O_1%X N_X_M1006_s N_X_M1009_s X X X X X X X N_X_c_257_n
+ X PM_SKY130_FD_SC_LP__A22O_1%X
x_PM_SKY130_FD_SC_LP__A22O_1%VPWR N_VPWR_M1009_d N_VPWR_M1008_d N_VPWR_c_273_n
+ N_VPWR_c_274_n VPWR N_VPWR_c_275_n N_VPWR_c_276_n N_VPWR_c_277_n
+ N_VPWR_c_272_n N_VPWR_c_279_n N_VPWR_c_280_n PM_SKY130_FD_SC_LP__A22O_1%VPWR
x_PM_SKY130_FD_SC_LP__A22O_1%A_217_367# N_A_217_367#_M1002_s
+ N_A_217_367#_M1005_d N_A_217_367#_M1000_d N_A_217_367#_c_317_n
+ N_A_217_367#_c_318_n N_A_217_367#_c_323_n N_A_217_367#_c_332_n
+ N_A_217_367#_c_333_n N_A_217_367#_c_319_n N_A_217_367#_c_320_n
+ N_A_217_367#_c_321_n PM_SKY130_FD_SC_LP__A22O_1%A_217_367#
x_PM_SKY130_FD_SC_LP__A22O_1%VGND N_VGND_M1006_d N_VGND_M1001_d N_VGND_c_359_n
+ N_VGND_c_360_n VGND N_VGND_c_361_n N_VGND_c_362_n N_VGND_c_363_n
+ N_VGND_c_364_n PM_SKY130_FD_SC_LP__A22O_1%VGND
cc_1 VNB N_A_80_246#_M1009_g 0.00548882f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.465
cc_2 VNB N_A_80_246#_c_57_n 0.0209106f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=1.23
cc_3 VNB N_A_80_246#_c_58_n 0.00309511f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=1.395
cc_4 VNB N_A_80_246#_c_59_n 0.0504129f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=1.395
cc_5 VNB N_A_80_246#_c_60_n 0.00736132f $X=-0.19 $Y=-0.245 $X2=1.475 $Y2=1.735
cc_6 VNB N_A_80_246#_c_61_n 0.00313833f $X=-0.19 $Y=-0.245 $X2=2.06 $Y2=0.42
cc_7 VNB N_B2_c_123_n 0.0186912f $X=-0.19 $Y=-0.245 $X2=1.86 $Y2=0.28
cc_8 VNB N_B2_M1002_g 0.0058622f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB B2 0.00508982f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.465
cc_10 VNB N_B2_c_126_n 0.0374157f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=0.7
cc_11 VNB N_B1_M1005_g 0.00521331f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_B1_c_157_n 0.0298407f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=1.23
cc_13 VNB N_B1_c_158_n 0.00756677f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=0.7
cc_14 VNB N_B1_c_159_n 0.017352f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=0.7
cc_15 VNB N_A1_M1008_g 0.00553928f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB A1 0.00170212f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.465
cc_17 VNB A1 0.00705046f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A1_c_195_n 0.0306857f $X=-0.19 $Y=-0.245 $X2=0.725 $Y2=1.395
cc_19 VNB N_A1_c_196_n 0.018719f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=1.395
cc_20 VNB N_A2_M1000_g 0.00809292f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB A2 0.0191086f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.465
cc_22 VNB N_A2_c_232_n 0.0389946f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=1.23
cc_23 VNB N_A2_c_233_n 0.0221737f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=0.7
cc_24 VNB X 0.00916912f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.465
cc_25 VNB X 0.0271351f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.465
cc_26 VNB N_X_c_257_n 0.0326457f $X=-0.19 $Y=-0.245 $X2=1.64 $Y2=1.98
cc_27 VNB N_VPWR_c_272_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_359_n 0.0113448f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.56
cc_29 VNB N_VGND_c_360_n 0.0348513f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.465
cc_30 VNB N_VGND_c_361_n 0.0174909f $X=-0.19 $Y=-0.245 $X2=0.555 $Y2=0.7
cc_31 VNB N_VGND_c_362_n 0.0433138f $X=-0.19 $Y=-0.245 $X2=0.71 $Y2=1.395
cc_32 VNB N_VGND_c_363_n 0.0165489f $X=-0.19 $Y=-0.245 $X2=2.06 $Y2=0.42
cc_33 VNB N_VGND_c_364_n 0.213661f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VPB N_A_80_246#_M1009_g 0.0268543f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.465
cc_35 VPB N_A_80_246#_c_60_n 0.0119937f $X=-0.19 $Y=1.655 $X2=1.475 $Y2=1.735
cc_36 VPB N_A_80_246#_c_64_n 0.0040507f $X=-0.19 $Y=1.655 $X2=0.845 $Y2=1.735
cc_37 VPB N_B2_M1002_g 0.0242982f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_38 VPB N_B1_M1005_g 0.0199009f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_39 VPB N_A1_M1008_g 0.02073f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_40 VPB N_A2_M1000_g 0.0267712f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_41 VPB X 0.056696f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.465
cc_42 VPB N_VPWR_c_273_n 0.0154975f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.465
cc_43 VPB N_VPWR_c_274_n 0.00557848f $X=-0.19 $Y=1.655 $X2=0.725 $Y2=1.65
cc_44 VPB N_VPWR_c_275_n 0.0182379f $X=-0.19 $Y=1.655 $X2=1.475 $Y2=1.735
cc_45 VPB N_VPWR_c_276_n 0.0381285f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_46 VPB N_VPWR_c_277_n 0.0180487f $X=-0.19 $Y=1.655 $X2=0.71 $Y2=1.395
cc_47 VPB N_VPWR_c_272_n 0.0537482f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_48 VPB N_VPWR_c_279_n 0.00516749f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_49 VPB N_VPWR_c_280_n 0.0065069f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_50 VPB N_A_217_367#_c_317_n 0.001829f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_51 VPB N_A_217_367#_c_318_n 0.00849997f $X=-0.19 $Y=1.655 $X2=0.555 $Y2=0.7
cc_52 VPB N_A_217_367#_c_319_n 0.0141496f $X=-0.19 $Y=1.655 $X2=0.845 $Y2=0.955
cc_53 VPB N_A_217_367#_c_320_n 0.00994699f $X=-0.19 $Y=1.655 $X2=1.475 $Y2=1.735
cc_54 VPB N_A_217_367#_c_321_n 0.0453969f $X=-0.19 $Y=1.655 $X2=1.64 $Y2=1.98
cc_55 N_A_80_246#_c_57_n N_B2_c_123_n 0.00818263f $X=0.555 $Y=1.23 $X2=-0.19
+ $Y2=-0.245
cc_56 N_A_80_246#_c_58_n N_B2_c_123_n 0.00305753f $X=0.71 $Y=1.395 $X2=-0.19
+ $Y2=-0.245
cc_57 N_A_80_246#_c_67_p N_B2_c_123_n 0.0162269f $X=1.895 $Y=0.955 $X2=-0.19
+ $Y2=-0.245
cc_58 N_A_80_246#_c_58_n N_B2_M1002_g 0.00223473f $X=0.71 $Y=1.395 $X2=0 $Y2=0
cc_59 N_A_80_246#_c_60_n N_B2_M1002_g 0.0168142f $X=1.475 $Y=1.735 $X2=0 $Y2=0
cc_60 N_A_80_246#_c_70_p N_B2_M1002_g 0.0192365f $X=1.64 $Y=1.98 $X2=0 $Y2=0
cc_61 N_A_80_246#_c_58_n B2 0.0212949f $X=0.71 $Y=1.395 $X2=0 $Y2=0
cc_62 N_A_80_246#_c_59_n B2 0.0015973f $X=0.71 $Y=1.395 $X2=0 $Y2=0
cc_63 N_A_80_246#_c_67_p B2 0.0279942f $X=1.895 $Y=0.955 $X2=0 $Y2=0
cc_64 N_A_80_246#_c_60_n B2 0.029644f $X=1.475 $Y=1.735 $X2=0 $Y2=0
cc_65 N_A_80_246#_c_58_n N_B2_c_126_n 8.03e-19 $X=0.71 $Y=1.395 $X2=0 $Y2=0
cc_66 N_A_80_246#_c_59_n N_B2_c_126_n 0.0216899f $X=0.71 $Y=1.395 $X2=0 $Y2=0
cc_67 N_A_80_246#_c_67_p N_B2_c_126_n 0.00144428f $X=1.895 $Y=0.955 $X2=0 $Y2=0
cc_68 N_A_80_246#_c_60_n N_B2_c_126_n 0.00665676f $X=1.475 $Y=1.735 $X2=0 $Y2=0
cc_69 N_A_80_246#_c_60_n N_B1_M1005_g 0.00446989f $X=1.475 $Y=1.735 $X2=0 $Y2=0
cc_70 N_A_80_246#_c_70_p N_B1_M1005_g 0.0116513f $X=1.64 $Y=1.98 $X2=0 $Y2=0
cc_71 N_A_80_246#_c_60_n N_B1_c_157_n 0.00269808f $X=1.475 $Y=1.735 $X2=0 $Y2=0
cc_72 N_A_80_246#_c_82_p N_B1_c_157_n 0.00101827f $X=2.06 $Y=0.87 $X2=0 $Y2=0
cc_73 N_A_80_246#_c_67_p N_B1_c_158_n 0.0194733f $X=1.895 $Y=0.955 $X2=0 $Y2=0
cc_74 N_A_80_246#_c_60_n N_B1_c_158_n 0.0187812f $X=1.475 $Y=1.735 $X2=0 $Y2=0
cc_75 N_A_80_246#_c_82_p N_B1_c_158_n 0.0114012f $X=2.06 $Y=0.87 $X2=0 $Y2=0
cc_76 N_A_80_246#_c_67_p N_B1_c_159_n 0.015067f $X=1.895 $Y=0.955 $X2=0 $Y2=0
cc_77 N_A_80_246#_c_61_n N_B1_c_159_n 0.00380582f $X=2.06 $Y=0.42 $X2=0 $Y2=0
cc_78 N_A_80_246#_c_60_n N_A1_M1008_g 4.31297e-19 $X=1.475 $Y=1.735 $X2=0 $Y2=0
cc_79 N_A_80_246#_c_70_p N_A1_M1008_g 3.04372e-19 $X=1.64 $Y=1.98 $X2=0 $Y2=0
cc_80 N_A_80_246#_c_61_n N_A1_c_196_n 0.00157944f $X=2.06 $Y=0.42 $X2=0 $Y2=0
cc_81 N_A_80_246#_c_58_n X 0.00433183f $X=0.71 $Y=1.395 $X2=0 $Y2=0
cc_82 N_A_80_246#_c_59_n X 0.00179468f $X=0.71 $Y=1.395 $X2=0 $Y2=0
cc_83 N_A_80_246#_c_57_n X 0.00192838f $X=0.555 $Y=1.23 $X2=0 $Y2=0
cc_84 N_A_80_246#_c_58_n X 0.0302765f $X=0.71 $Y=1.395 $X2=0 $Y2=0
cc_85 N_A_80_246#_c_59_n X 0.0189298f $X=0.71 $Y=1.395 $X2=0 $Y2=0
cc_86 N_A_80_246#_c_64_n X 0.0116228f $X=0.845 $Y=1.735 $X2=0 $Y2=0
cc_87 N_A_80_246#_c_57_n N_X_c_257_n 0.00411342f $X=0.555 $Y=1.23 $X2=0 $Y2=0
cc_88 N_A_80_246#_M1009_g N_VPWR_c_273_n 0.00507622f $X=0.475 $Y=2.465 $X2=0
+ $Y2=0
cc_89 N_A_80_246#_c_59_n N_VPWR_c_273_n 0.00109093f $X=0.71 $Y=1.395 $X2=0 $Y2=0
cc_90 N_A_80_246#_c_60_n N_VPWR_c_273_n 7.2232e-19 $X=1.475 $Y=1.735 $X2=0 $Y2=0
cc_91 N_A_80_246#_c_64_n N_VPWR_c_273_n 0.0220259f $X=0.845 $Y=1.735 $X2=0 $Y2=0
cc_92 N_A_80_246#_M1009_g N_VPWR_c_275_n 0.00585385f $X=0.475 $Y=2.465 $X2=0
+ $Y2=0
cc_93 N_A_80_246#_M1002_d N_VPWR_c_272_n 0.0024127f $X=1.5 $Y=1.835 $X2=0 $Y2=0
cc_94 N_A_80_246#_M1009_g N_VPWR_c_272_n 0.012823f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_95 N_A_80_246#_c_60_n N_A_217_367#_c_318_n 0.0209093f $X=1.475 $Y=1.735 $X2=0
+ $Y2=0
cc_96 N_A_80_246#_M1002_d N_A_217_367#_c_323_n 0.00372385f $X=1.5 $Y=1.835 $X2=0
+ $Y2=0
cc_97 N_A_80_246#_c_70_p N_A_217_367#_c_323_n 0.0160777f $X=1.64 $Y=1.98 $X2=0
+ $Y2=0
cc_98 N_A_80_246#_c_60_n N_A_217_367#_c_320_n 0.00802266f $X=1.475 $Y=1.735
+ $X2=0 $Y2=0
cc_99 N_A_80_246#_c_70_p N_A_217_367#_c_320_n 0.00363101f $X=1.64 $Y=1.98 $X2=0
+ $Y2=0
cc_100 N_A_80_246#_c_58_n N_VGND_M1006_d 0.00125798f $X=0.71 $Y=1.395 $X2=-0.19
+ $Y2=-0.245
cc_101 N_A_80_246#_c_67_p N_VGND_M1006_d 0.0124545f $X=1.895 $Y=0.955 $X2=-0.19
+ $Y2=-0.245
cc_102 N_A_80_246#_c_112_p N_VGND_M1006_d 0.0020778f $X=0.845 $Y=0.955 $X2=-0.19
+ $Y2=-0.245
cc_103 N_A_80_246#_c_57_n N_VGND_c_361_n 0.00450636f $X=0.555 $Y=1.23 $X2=0
+ $Y2=0
cc_104 N_A_80_246#_c_61_n N_VGND_c_362_n 0.0235133f $X=2.06 $Y=0.42 $X2=0 $Y2=0
cc_105 N_A_80_246#_c_57_n N_VGND_c_363_n 0.0127851f $X=0.555 $Y=1.23 $X2=0 $Y2=0
cc_106 N_A_80_246#_c_59_n N_VGND_c_363_n 7.72205e-19 $X=0.71 $Y=1.395 $X2=0
+ $Y2=0
cc_107 N_A_80_246#_c_67_p N_VGND_c_363_n 0.0357575f $X=1.895 $Y=0.955 $X2=0
+ $Y2=0
cc_108 N_A_80_246#_c_112_p N_VGND_c_363_n 0.0162349f $X=0.845 $Y=0.955 $X2=0
+ $Y2=0
cc_109 N_A_80_246#_c_61_n N_VGND_c_363_n 0.00754689f $X=2.06 $Y=0.42 $X2=0 $Y2=0
cc_110 N_A_80_246#_c_57_n N_VGND_c_364_n 0.00885506f $X=0.555 $Y=1.23 $X2=0
+ $Y2=0
cc_111 N_A_80_246#_c_61_n N_VGND_c_364_n 0.0127519f $X=2.06 $Y=0.42 $X2=0 $Y2=0
cc_112 N_A_80_246#_c_67_p A_294_56# 0.0066275f $X=1.895 $Y=0.955 $X2=-0.19
+ $Y2=-0.245
cc_113 N_B2_M1002_g N_B1_M1005_g 0.039741f $X=1.425 $Y=2.465 $X2=0 $Y2=0
cc_114 N_B2_c_126_n N_B1_c_157_n 0.0439053f $X=1.395 $Y=1.395 $X2=0 $Y2=0
cc_115 N_B2_c_123_n N_B1_c_158_n 0.00139426f $X=1.395 $Y=1.23 $X2=0 $Y2=0
cc_116 B2 N_B1_c_158_n 0.0221298f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_117 N_B2_c_126_n N_B1_c_158_n 4.91622e-19 $X=1.395 $Y=1.395 $X2=0 $Y2=0
cc_118 N_B2_c_123_n N_B1_c_159_n 0.03344f $X=1.395 $Y=1.23 $X2=0 $Y2=0
cc_119 B2 N_B1_c_159_n 2.40881e-19 $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_120 N_B2_M1002_g N_VPWR_c_273_n 0.0022664f $X=1.425 $Y=2.465 $X2=0 $Y2=0
cc_121 N_B2_M1002_g N_VPWR_c_276_n 0.00357877f $X=1.425 $Y=2.465 $X2=0 $Y2=0
cc_122 N_B2_M1002_g N_VPWR_c_272_n 0.00672955f $X=1.425 $Y=2.465 $X2=0 $Y2=0
cc_123 N_B2_M1002_g N_A_217_367#_c_323_n 0.011572f $X=1.425 $Y=2.465 $X2=0 $Y2=0
cc_124 N_B2_c_123_n N_VGND_c_362_n 0.00450636f $X=1.395 $Y=1.23 $X2=0 $Y2=0
cc_125 N_B2_c_123_n N_VGND_c_363_n 0.0155803f $X=1.395 $Y=1.23 $X2=0 $Y2=0
cc_126 N_B2_c_123_n N_VGND_c_364_n 0.00806919f $X=1.395 $Y=1.23 $X2=0 $Y2=0
cc_127 N_B1_M1005_g N_A1_M1008_g 0.0229977f $X=1.875 $Y=2.465 $X2=0 $Y2=0
cc_128 N_B1_c_157_n A1 7.56264e-19 $X=1.875 $Y=1.395 $X2=0 $Y2=0
cc_129 N_B1_c_158_n A1 0.0137631f $X=1.875 $Y=1.395 $X2=0 $Y2=0
cc_130 N_B1_c_157_n N_A1_c_195_n 0.021213f $X=1.875 $Y=1.395 $X2=0 $Y2=0
cc_131 N_B1_c_158_n N_A1_c_195_n 9.20483e-19 $X=1.875 $Y=1.395 $X2=0 $Y2=0
cc_132 N_B1_c_159_n N_A1_c_196_n 0.0190524f $X=1.875 $Y=1.23 $X2=0 $Y2=0
cc_133 N_B1_M1005_g N_VPWR_c_276_n 0.00357877f $X=1.875 $Y=2.465 $X2=0 $Y2=0
cc_134 N_B1_M1005_g N_VPWR_c_272_n 0.00546654f $X=1.875 $Y=2.465 $X2=0 $Y2=0
cc_135 N_B1_M1005_g N_A_217_367#_c_323_n 0.012129f $X=1.875 $Y=2.465 $X2=0 $Y2=0
cc_136 N_B1_M1005_g N_A_217_367#_c_320_n 9.26765e-19 $X=1.875 $Y=2.465 $X2=0
+ $Y2=0
cc_137 N_B1_c_157_n N_A_217_367#_c_320_n 0.00159811f $X=1.875 $Y=1.395 $X2=0
+ $Y2=0
cc_138 N_B1_c_158_n N_A_217_367#_c_320_n 0.00405564f $X=1.875 $Y=1.395 $X2=0
+ $Y2=0
cc_139 N_B1_c_159_n N_VGND_c_362_n 0.00540763f $X=1.875 $Y=1.23 $X2=0 $Y2=0
cc_140 N_B1_c_159_n N_VGND_c_363_n 0.00215724f $X=1.875 $Y=1.23 $X2=0 $Y2=0
cc_141 N_B1_c_159_n N_VGND_c_364_n 0.0106239f $X=1.875 $Y=1.23 $X2=0 $Y2=0
cc_142 N_A1_M1008_g N_A2_M1000_g 0.0300385f $X=2.325 $Y=2.465 $X2=0 $Y2=0
cc_143 A1 A2 0.0283208f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_144 N_A1_c_195_n A2 2.5763e-19 $X=2.415 $Y=1.395 $X2=0 $Y2=0
cc_145 A1 N_A2_c_232_n 0.00457637f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_146 N_A1_c_195_n N_A2_c_232_n 0.0205208f $X=2.415 $Y=1.395 $X2=0 $Y2=0
cc_147 A1 N_A2_c_233_n 0.00457637f $X=2.555 $Y=0.47 $X2=0 $Y2=0
cc_148 N_A1_c_196_n N_A2_c_233_n 0.0253341f $X=2.415 $Y=1.23 $X2=0 $Y2=0
cc_149 N_A1_M1008_g N_VPWR_c_274_n 0.00935148f $X=2.325 $Y=2.465 $X2=0 $Y2=0
cc_150 N_A1_M1008_g N_VPWR_c_276_n 0.00577794f $X=2.325 $Y=2.465 $X2=0 $Y2=0
cc_151 N_A1_M1008_g N_VPWR_c_272_n 0.0108473f $X=2.325 $Y=2.465 $X2=0 $Y2=0
cc_152 N_A1_M1008_g N_A_217_367#_c_332_n 0.00152007f $X=2.325 $Y=2.465 $X2=0
+ $Y2=0
cc_153 N_A1_M1008_g N_A_217_367#_c_333_n 0.0120559f $X=2.325 $Y=2.465 $X2=0
+ $Y2=0
cc_154 N_A1_M1008_g N_A_217_367#_c_319_n 0.0154326f $X=2.325 $Y=2.465 $X2=0
+ $Y2=0
cc_155 A1 N_A_217_367#_c_319_n 0.032166f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_156 N_A1_c_195_n N_A_217_367#_c_319_n 0.00126891f $X=2.415 $Y=1.395 $X2=0
+ $Y2=0
cc_157 N_A1_M1008_g N_A_217_367#_c_320_n 0.00142064f $X=2.325 $Y=2.465 $X2=0
+ $Y2=0
cc_158 N_A1_M1008_g N_A_217_367#_c_321_n 9.65196e-19 $X=2.325 $Y=2.465 $X2=0
+ $Y2=0
cc_159 N_A1_c_196_n N_VGND_c_360_n 0.00147184f $X=2.415 $Y=1.23 $X2=0 $Y2=0
cc_160 A1 N_VGND_c_362_n 0.0102499f $X=2.555 $Y=0.47 $X2=0 $Y2=0
cc_161 N_A1_c_196_n N_VGND_c_362_n 0.00540763f $X=2.415 $Y=1.23 $X2=0 $Y2=0
cc_162 A1 N_VGND_c_364_n 0.0101568f $X=2.555 $Y=0.47 $X2=0 $Y2=0
cc_163 N_A1_c_196_n N_VGND_c_364_n 0.0108745f $X=2.415 $Y=1.23 $X2=0 $Y2=0
cc_164 A1 A_480_56# 0.0134139f $X=2.555 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_165 N_A2_M1000_g N_VPWR_c_274_n 0.00334987f $X=2.865 $Y=2.465 $X2=0 $Y2=0
cc_166 N_A2_M1000_g N_VPWR_c_277_n 0.00579312f $X=2.865 $Y=2.465 $X2=0 $Y2=0
cc_167 N_A2_M1000_g N_VPWR_c_272_n 0.0116435f $X=2.865 $Y=2.465 $X2=0 $Y2=0
cc_168 N_A2_M1000_g N_A_217_367#_c_333_n 6.74841e-19 $X=2.865 $Y=2.465 $X2=0
+ $Y2=0
cc_169 N_A2_M1000_g N_A_217_367#_c_319_n 0.0189046f $X=2.865 $Y=2.465 $X2=0
+ $Y2=0
cc_170 A2 N_A_217_367#_c_319_n 0.0287197f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_171 N_A2_c_232_n N_A_217_367#_c_319_n 0.00500857f $X=2.99 $Y=1.395 $X2=0
+ $Y2=0
cc_172 N_A2_M1000_g N_A_217_367#_c_321_n 0.0150759f $X=2.865 $Y=2.465 $X2=0
+ $Y2=0
cc_173 A2 N_VGND_c_360_n 0.02586f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_174 N_A2_c_232_n N_VGND_c_360_n 0.00144567f $X=2.99 $Y=1.395 $X2=0 $Y2=0
cc_175 N_A2_c_233_n N_VGND_c_360_n 0.0180503f $X=2.972 $Y=1.23 $X2=0 $Y2=0
cc_176 N_A2_c_233_n N_VGND_c_362_n 0.00448994f $X=2.972 $Y=1.23 $X2=0 $Y2=0
cc_177 N_A2_c_233_n N_VGND_c_364_n 0.00831975f $X=2.972 $Y=1.23 $X2=0 $Y2=0
cc_178 X N_VPWR_c_275_n 0.0181659f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_179 N_X_M1009_s N_VPWR_c_272_n 0.00336915f $X=0.135 $Y=1.835 $X2=0 $Y2=0
cc_180 X N_VPWR_c_272_n 0.0104192f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_181 N_X_c_257_n N_VGND_c_361_n 0.0242301f $X=0.34 $Y=0.425 $X2=0 $Y2=0
cc_182 N_X_c_257_n N_VGND_c_363_n 0.0196597f $X=0.34 $Y=0.425 $X2=0 $Y2=0
cc_183 N_X_c_257_n N_VGND_c_364_n 0.0131407f $X=0.34 $Y=0.425 $X2=0 $Y2=0
cc_184 N_VPWR_c_272_n N_A_217_367#_M1002_s 0.00215161f $X=3.12 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_185 N_VPWR_c_272_n N_A_217_367#_M1005_d 0.00239644f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_186 N_VPWR_c_272_n N_A_217_367#_M1000_d 0.00215158f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_187 N_VPWR_c_273_n N_A_217_367#_c_317_n 0.0137034f $X=0.69 $Y=2.155 $X2=0
+ $Y2=0
cc_188 N_VPWR_c_276_n N_A_217_367#_c_317_n 0.0179183f $X=2.425 $Y=3.33 $X2=0
+ $Y2=0
cc_189 N_VPWR_c_272_n N_A_217_367#_c_317_n 0.0101082f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_190 N_VPWR_c_273_n N_A_217_367#_c_318_n 0.0681172f $X=0.69 $Y=2.155 $X2=0
+ $Y2=0
cc_191 N_VPWR_c_276_n N_A_217_367#_c_323_n 0.0366794f $X=2.425 $Y=3.33 $X2=0
+ $Y2=0
cc_192 N_VPWR_c_272_n N_A_217_367#_c_323_n 0.023676f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_193 N_VPWR_c_276_n N_A_217_367#_c_332_n 0.0165441f $X=2.425 $Y=3.33 $X2=0
+ $Y2=0
cc_194 N_VPWR_c_272_n N_A_217_367#_c_332_n 0.0107897f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_195 N_VPWR_M1008_d N_A_217_367#_c_319_n 0.00304021f $X=2.4 $Y=1.835 $X2=0
+ $Y2=0
cc_196 N_VPWR_c_274_n N_A_217_367#_c_319_n 0.022455f $X=2.6 $Y=2.155 $X2=0 $Y2=0
cc_197 N_VPWR_c_277_n N_A_217_367#_c_321_n 0.0196832f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_198 N_VPWR_c_272_n N_A_217_367#_c_321_n 0.0118828f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
