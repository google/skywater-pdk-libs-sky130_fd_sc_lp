* File: sky130_fd_sc_lp__a21boi_4.pxi.spice
* Created: Fri Aug 28 09:50:15 2020
* 
x_PM_SKY130_FD_SC_LP__A21BOI_4%B1_N N_B1_N_M1007_g N_B1_N_c_103_n N_B1_N_M1014_g
+ B1_N B1_N N_B1_N_c_105_n PM_SKY130_FD_SC_LP__A21BOI_4%B1_N
x_PM_SKY130_FD_SC_LP__A21BOI_4%A_33_367# N_A_33_367#_M1014_s N_A_33_367#_M1007_s
+ N_A_33_367#_M1000_g N_A_33_367#_M1002_g N_A_33_367#_M1005_g
+ N_A_33_367#_M1009_g N_A_33_367#_M1017_g N_A_33_367#_M1016_g
+ N_A_33_367#_M1018_g N_A_33_367#_M1022_g N_A_33_367#_c_154_n
+ N_A_33_367#_c_155_n N_A_33_367#_c_144_n N_A_33_367#_c_156_n
+ N_A_33_367#_c_164_n N_A_33_367#_c_145_n N_A_33_367#_c_146_n
+ N_A_33_367#_c_147_n N_A_33_367#_c_219_p N_A_33_367#_c_148_n
+ N_A_33_367#_c_149_n PM_SKY130_FD_SC_LP__A21BOI_4%A_33_367#
x_PM_SKY130_FD_SC_LP__A21BOI_4%A2 N_A2_M1001_g N_A2_M1004_g N_A2_c_266_n
+ N_A2_M1010_g N_A2_M1011_g N_A2_c_268_n N_A2_M1015_g N_A2_M1013_g N_A2_c_270_n
+ N_A2_M1023_g N_A2_M1025_g N_A2_c_272_n N_A2_c_273_n A2 A2 A2 N_A2_c_276_n
+ N_A2_c_277_n N_A2_c_278_n PM_SKY130_FD_SC_LP__A21BOI_4%A2
x_PM_SKY130_FD_SC_LP__A21BOI_4%A1 N_A1_M1003_g N_A1_M1006_g N_A1_M1008_g
+ N_A1_M1012_g N_A1_M1020_g N_A1_M1019_g N_A1_M1021_g N_A1_M1024_g A1 A1 A1 A1
+ N_A1_c_382_n PM_SKY130_FD_SC_LP__A21BOI_4%A1
x_PM_SKY130_FD_SC_LP__A21BOI_4%VPWR N_VPWR_M1007_d N_VPWR_M1001_s N_VPWR_M1012_d
+ N_VPWR_M1024_d N_VPWR_M1013_s N_VPWR_c_456_n N_VPWR_c_488_n N_VPWR_c_457_n
+ N_VPWR_c_506_n N_VPWR_c_458_n N_VPWR_c_459_n N_VPWR_c_460_n N_VPWR_c_461_n
+ VPWR N_VPWR_c_462_n N_VPWR_c_463_n N_VPWR_c_464_n N_VPWR_c_465_n
+ N_VPWR_c_455_n N_VPWR_c_467_n N_VPWR_c_468_n N_VPWR_c_469_n
+ PM_SKY130_FD_SC_LP__A21BOI_4%VPWR
x_PM_SKY130_FD_SC_LP__A21BOI_4%A_223_367# N_A_223_367#_M1002_d
+ N_A_223_367#_M1009_d N_A_223_367#_M1022_d N_A_223_367#_M1006_s
+ N_A_223_367#_M1019_s N_A_223_367#_M1011_d N_A_223_367#_M1025_d
+ N_A_223_367#_c_559_n N_A_223_367#_c_560_n N_A_223_367#_c_570_n
+ N_A_223_367#_c_572_n N_A_223_367#_c_575_n N_A_223_367#_c_627_n
+ N_A_223_367#_c_577_n N_A_223_367#_c_582_n N_A_223_367#_c_578_n
+ N_A_223_367#_c_603_n N_A_223_367#_c_637_n N_A_223_367#_c_588_n
+ N_A_223_367#_c_641_n N_A_223_367#_c_561_n N_A_223_367#_c_562_n
+ N_A_223_367#_c_579_n N_A_223_367#_c_607_n N_A_223_367#_c_563_n
+ PM_SKY130_FD_SC_LP__A21BOI_4%A_223_367#
x_PM_SKY130_FD_SC_LP__A21BOI_4%Y N_Y_M1000_s N_Y_M1017_s N_Y_M1003_s N_Y_M1020_s
+ N_Y_M1002_s N_Y_M1016_s N_Y_c_666_n N_Y_c_658_n N_Y_c_662_n N_Y_c_729_p
+ N_Y_c_696_n N_Y_c_677_n N_Y_c_663_n Y Y Y Y N_Y_c_660_n N_Y_c_661_n
+ PM_SKY130_FD_SC_LP__A21BOI_4%Y
x_PM_SKY130_FD_SC_LP__A21BOI_4%VGND N_VGND_M1014_d N_VGND_M1005_d N_VGND_M1018_d
+ N_VGND_M1010_d N_VGND_M1023_d N_VGND_c_745_n N_VGND_c_746_n N_VGND_c_747_n
+ N_VGND_c_748_n N_VGND_c_749_n N_VGND_c_750_n N_VGND_c_751_n N_VGND_c_752_n
+ VGND N_VGND_c_753_n N_VGND_c_754_n N_VGND_c_755_n N_VGND_c_756_n
+ N_VGND_c_757_n N_VGND_c_758_n N_VGND_c_759_n PM_SKY130_FD_SC_LP__A21BOI_4%VGND
x_PM_SKY130_FD_SC_LP__A21BOI_4%A_658_47# N_A_658_47#_M1004_s N_A_658_47#_M1008_d
+ N_A_658_47#_M1021_d N_A_658_47#_M1015_s N_A_658_47#_c_840_n
+ N_A_658_47#_c_842_n N_A_658_47#_c_843_n N_A_658_47#_c_846_n
+ N_A_658_47#_c_851_n N_A_658_47#_c_875_n PM_SKY130_FD_SC_LP__A21BOI_4%A_658_47#
cc_1 VNB N_B1_N_M1007_g 0.00910877f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.465
cc_2 VNB N_B1_N_c_103_n 0.0222299f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=1.185
cc_3 VNB B1_N 0.030329f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_4 VNB N_B1_N_c_105_n 0.0373213f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=1.35
cc_5 VNB N_A_33_367#_M1000_g 0.0199775f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_6 VNB N_A_33_367#_M1002_g 0.00162055f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_A_33_367#_M1005_g 0.0194532f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_33_367#_M1009_g 0.00147374f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=1.35
cc_9 VNB N_A_33_367#_M1017_g 0.0194411f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_33_367#_M1016_g 0.00146748f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_33_367#_M1018_g 0.0226963f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_33_367#_M1022_g 0.00126884f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_33_367#_c_144_n 0.0235964f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_33_367#_c_145_n 0.00753748f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_33_367#_c_146_n 0.00231769f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_33_367#_c_147_n 0.00104164f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_33_367#_c_148_n 0.00107567f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_33_367#_c_149_n 0.109945f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A2_M1001_g 0.007686f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.465
cc_20 VNB N_A2_c_266_n 0.0153283f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_21 VNB N_A2_M1011_g 0.00726311f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A2_c_268_n 0.0161573f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A2_M1013_g 0.00706537f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=1.35
cc_24 VNB N_A2_c_270_n 0.0220609f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A2_M1025_g 0.0111859f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=1.48
cc_26 VNB N_A2_c_272_n 0.00278935f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A2_c_273_n 0.034992f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB A2 0.00274088f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB A2 0.0152949f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A2_c_276_n 0.0176974f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A2_c_277_n 0.0738534f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A2_c_278_n 0.0264324f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A1_M1003_g 0.0226607f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.465
cc_34 VNB N_A1_M1008_g 0.0229017f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A1_M1020_g 0.0229027f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=1.35
cc_36 VNB N_A1_M1021_g 0.0231059f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=1.48
cc_37 VNB A1 0.00638505f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A1_c_382_n 0.0630975f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_VPWR_c_455_n 0.283096f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_Y_c_658_n 0.00204712f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB Y 0.00704793f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_Y_c_660_n 0.00285879f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_Y_c_661_n 0.00426665f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_745_n 4.02668e-19 $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=1.35
cc_45 VNB N_VGND_c_746_n 0.0137825f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=1.35
cc_46 VNB N_VGND_c_747_n 3.19421e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_748_n 0.00438797f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.48
cc_48 VNB N_VGND_c_749_n 0.0116397f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_750_n 0.035768f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_751_n 0.0231432f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_752_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_753_n 0.0547364f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_754_n 0.0156625f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_755_n 0.00412824f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_756_n 0.0142001f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_VGND_c_757_n 0.016982f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_VGND_c_758_n 0.00439334f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_759_n 0.338061f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VPB N_B1_N_M1007_g 0.029639f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=2.465
cc_60 VPB B1_N 0.00962124f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_61 VPB N_A_33_367#_M1002_g 0.0228505f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_62 VPB N_A_33_367#_M1009_g 0.0187589f $X=-0.19 $Y=1.655 $X2=0.705 $Y2=1.35
cc_63 VPB N_A_33_367#_M1016_g 0.018746f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_64 VPB N_A_33_367#_M1022_g 0.0191689f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_65 VPB N_A_33_367#_c_154_n 0.00849091f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_66 VPB N_A_33_367#_c_155_n 0.0373194f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_67 VPB N_A_33_367#_c_156_n 0.0140011f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_68 VPB N_A_33_367#_c_147_n 0.00484149f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_69 VPB N_A2_M1001_g 0.020769f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=2.465
cc_70 VPB N_A2_M1011_g 0.019239f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_71 VPB N_A2_M1013_g 0.0183279f $X=-0.19 $Y=1.655 $X2=0.595 $Y2=1.35
cc_72 VPB N_A2_M1025_g 0.0241666f $X=-0.19 $Y=1.655 $X2=0.595 $Y2=1.48
cc_73 VPB N_A1_M1006_g 0.0182143f $X=-0.19 $Y=1.655 $X2=0.705 $Y2=0.655
cc_74 VPB N_A1_M1012_g 0.0181378f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_75 VPB N_A1_M1019_g 0.0181378f $X=-0.19 $Y=1.655 $X2=0.24 $Y2=1.48
cc_76 VPB N_A1_M1024_g 0.0180751f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_77 VPB A1 0.0116988f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_78 VPB N_A1_c_382_n 0.0121733f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_79 VPB N_VPWR_c_456_n 0.0107662f $X=-0.19 $Y=1.655 $X2=0.595 $Y2=1.35
cc_80 VPB N_VPWR_c_457_n 4.89148e-19 $X=-0.19 $Y=1.655 $X2=0.705 $Y2=1.35
cc_81 VPB N_VPWR_c_458_n 3.99129e-19 $X=-0.19 $Y=1.655 $X2=0.72 $Y2=1.48
cc_82 VPB N_VPWR_c_459_n 3.99129e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_83 VPB N_VPWR_c_460_n 0.0550875f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_84 VPB N_VPWR_c_461_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_85 VPB N_VPWR_c_462_n 0.0163305f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_86 VPB N_VPWR_c_463_n 0.0324039f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_87 VPB N_VPWR_c_464_n 0.0130339f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_88 VPB N_VPWR_c_465_n 0.0160123f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_89 VPB N_VPWR_c_455_n 0.0554878f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_90 VPB N_VPWR_c_467_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_91 VPB N_VPWR_c_468_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_92 VPB N_VPWR_c_469_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_93 VPB N_A_223_367#_c_559_n 0.00400003f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_94 VPB N_A_223_367#_c_560_n 0.00389786f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_95 VPB N_A_223_367#_c_561_n 0.0160029f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_96 VPB N_A_223_367#_c_562_n 0.0435297f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_97 VPB N_A_223_367#_c_563_n 0.00205147f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_98 VPB N_Y_c_662_n 0.00323168f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_99 VPB N_Y_c_663_n 0.00186402f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_100 VPB Y 0.0012151f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_101 VPB Y 0.00296597f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_102 N_B1_N_c_103_n N_A_33_367#_M1000_g 0.0312014f $X=0.705 $Y=1.185 $X2=0
+ $Y2=0
cc_103 B1_N N_A_33_367#_M1000_g 2.00078e-19 $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_104 B1_N N_A_33_367#_c_154_n 0.0201608f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_105 N_B1_N_M1007_g N_A_33_367#_c_156_n 0.0141776f $X=0.505 $Y=2.465 $X2=0
+ $Y2=0
cc_106 B1_N N_A_33_367#_c_156_n 0.0293291f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_107 N_B1_N_c_105_n N_A_33_367#_c_156_n 7.36615e-19 $X=0.705 $Y=1.35 $X2=0
+ $Y2=0
cc_108 N_B1_N_c_103_n N_A_33_367#_c_164_n 0.0127813f $X=0.705 $Y=1.185 $X2=0
+ $Y2=0
cc_109 B1_N N_A_33_367#_c_164_n 0.0132509f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_110 B1_N N_A_33_367#_c_145_n 0.0230438f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_111 N_B1_N_c_105_n N_A_33_367#_c_145_n 0.00470677f $X=0.705 $Y=1.35 $X2=0
+ $Y2=0
cc_112 N_B1_N_c_103_n N_A_33_367#_c_146_n 0.0034633f $X=0.705 $Y=1.185 $X2=0
+ $Y2=0
cc_113 B1_N N_A_33_367#_c_146_n 0.0137578f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_114 N_B1_N_c_105_n N_A_33_367#_c_146_n 4.74271e-19 $X=0.705 $Y=1.35 $X2=0
+ $Y2=0
cc_115 N_B1_N_M1007_g N_A_33_367#_c_147_n 0.00545546f $X=0.505 $Y=2.465 $X2=0
+ $Y2=0
cc_116 B1_N N_A_33_367#_c_147_n 0.0174328f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_117 B1_N N_A_33_367#_c_148_n 0.01587f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_118 N_B1_N_c_105_n N_A_33_367#_c_148_n 5.11719e-19 $X=0.705 $Y=1.35 $X2=0
+ $Y2=0
cc_119 N_B1_N_M1007_g N_A_33_367#_c_149_n 0.00258497f $X=0.505 $Y=2.465 $X2=0
+ $Y2=0
cc_120 B1_N N_A_33_367#_c_149_n 0.00124324f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_121 N_B1_N_c_105_n N_A_33_367#_c_149_n 0.0129255f $X=0.705 $Y=1.35 $X2=0
+ $Y2=0
cc_122 N_B1_N_M1007_g N_VPWR_c_456_n 0.0198657f $X=0.505 $Y=2.465 $X2=0 $Y2=0
cc_123 N_B1_N_M1007_g N_VPWR_c_462_n 0.00486043f $X=0.505 $Y=2.465 $X2=0 $Y2=0
cc_124 N_B1_N_M1007_g N_VPWR_c_455_n 0.00920706f $X=0.505 $Y=2.465 $X2=0 $Y2=0
cc_125 N_B1_N_M1007_g N_A_223_367#_c_559_n 9.71886e-19 $X=0.505 $Y=2.465 $X2=0
+ $Y2=0
cc_126 N_B1_N_M1007_g N_A_223_367#_c_560_n 8.87949e-19 $X=0.505 $Y=2.465 $X2=0
+ $Y2=0
cc_127 N_B1_N_c_103_n N_VGND_c_745_n 0.010472f $X=0.705 $Y=1.185 $X2=0 $Y2=0
cc_128 N_B1_N_c_103_n N_VGND_c_751_n 0.00564095f $X=0.705 $Y=1.185 $X2=0 $Y2=0
cc_129 N_B1_N_c_103_n N_VGND_c_759_n 0.0105725f $X=0.705 $Y=1.185 $X2=0 $Y2=0
cc_130 N_A_33_367#_c_149_n N_A2_M1001_g 0.0234516f $X=2.445 $Y=1.45 $X2=0 $Y2=0
cc_131 N_A_33_367#_M1018_g N_A2_c_272_n 2.9646e-19 $X=2.445 $Y=0.655 $X2=0 $Y2=0
cc_132 N_A_33_367#_M1018_g N_A2_c_273_n 0.00446003f $X=2.445 $Y=0.655 $X2=0
+ $Y2=0
cc_133 N_A_33_367#_c_149_n N_A2_c_273_n 0.00376649f $X=2.445 $Y=1.45 $X2=0 $Y2=0
cc_134 N_A_33_367#_M1018_g N_A2_c_276_n 0.0118876f $X=2.445 $Y=0.655 $X2=0 $Y2=0
cc_135 N_A_33_367#_c_156_n N_VPWR_M1007_d 0.00610475f $X=0.975 $Y=2.005
+ $X2=-0.19 $Y2=-0.245
cc_136 N_A_33_367#_M1002_g N_VPWR_c_456_n 0.0036914f $X=1.455 $Y=2.465 $X2=0
+ $Y2=0
cc_137 N_A_33_367#_c_156_n N_VPWR_c_456_n 0.0220026f $X=0.975 $Y=2.005 $X2=0
+ $Y2=0
cc_138 N_A_33_367#_M1022_g N_VPWR_c_457_n 0.00102873f $X=2.745 $Y=2.465 $X2=0
+ $Y2=0
cc_139 N_A_33_367#_M1002_g N_VPWR_c_460_n 0.00357877f $X=1.455 $Y=2.465 $X2=0
+ $Y2=0
cc_140 N_A_33_367#_M1009_g N_VPWR_c_460_n 0.00357842f $X=1.885 $Y=2.465 $X2=0
+ $Y2=0
cc_141 N_A_33_367#_M1016_g N_VPWR_c_460_n 0.00357842f $X=2.315 $Y=2.465 $X2=0
+ $Y2=0
cc_142 N_A_33_367#_M1022_g N_VPWR_c_460_n 0.00357877f $X=2.745 $Y=2.465 $X2=0
+ $Y2=0
cc_143 N_A_33_367#_c_155_n N_VPWR_c_462_n 0.0178111f $X=0.29 $Y=2.455 $X2=0
+ $Y2=0
cc_144 N_A_33_367#_M1007_s N_VPWR_c_455_n 0.00371702f $X=0.165 $Y=1.835 $X2=0
+ $Y2=0
cc_145 N_A_33_367#_M1002_g N_VPWR_c_455_n 0.00665089f $X=1.455 $Y=2.465 $X2=0
+ $Y2=0
cc_146 N_A_33_367#_M1009_g N_VPWR_c_455_n 0.00535118f $X=1.885 $Y=2.465 $X2=0
+ $Y2=0
cc_147 N_A_33_367#_M1016_g N_VPWR_c_455_n 0.00535118f $X=2.315 $Y=2.465 $X2=0
+ $Y2=0
cc_148 N_A_33_367#_M1022_g N_VPWR_c_455_n 0.00544745f $X=2.745 $Y=2.465 $X2=0
+ $Y2=0
cc_149 N_A_33_367#_c_155_n N_VPWR_c_455_n 0.0100304f $X=0.29 $Y=2.455 $X2=0
+ $Y2=0
cc_150 N_A_33_367#_c_156_n N_A_223_367#_M1002_d 0.00352261f $X=0.975 $Y=2.005
+ $X2=-0.19 $Y2=-0.245
cc_151 N_A_33_367#_c_147_n N_A_223_367#_M1002_d 0.00127666f $X=1.085 $Y=1.92
+ $X2=-0.19 $Y2=-0.245
cc_152 N_A_33_367#_c_156_n N_A_223_367#_c_560_n 0.0108386f $X=0.975 $Y=2.005
+ $X2=0 $Y2=0
cc_153 N_A_33_367#_c_149_n N_A_223_367#_c_560_n 0.004344f $X=2.445 $Y=1.45 $X2=0
+ $Y2=0
cc_154 N_A_33_367#_M1002_g N_A_223_367#_c_570_n 0.0193953f $X=1.455 $Y=2.465
+ $X2=0 $Y2=0
cc_155 N_A_33_367#_M1009_g N_A_223_367#_c_570_n 0.014321f $X=1.885 $Y=2.465
+ $X2=0 $Y2=0
cc_156 N_A_33_367#_M1002_g N_A_223_367#_c_572_n 4.79434e-19 $X=1.455 $Y=2.465
+ $X2=0 $Y2=0
cc_157 N_A_33_367#_M1009_g N_A_223_367#_c_572_n 0.00648293f $X=1.885 $Y=2.465
+ $X2=0 $Y2=0
cc_158 N_A_33_367#_M1016_g N_A_223_367#_c_572_n 0.00497151f $X=2.315 $Y=2.465
+ $X2=0 $Y2=0
cc_159 N_A_33_367#_M1016_g N_A_223_367#_c_575_n 0.0123313f $X=2.315 $Y=2.465
+ $X2=0 $Y2=0
cc_160 N_A_33_367#_M1022_g N_A_223_367#_c_575_n 0.0125861f $X=2.745 $Y=2.465
+ $X2=0 $Y2=0
cc_161 N_A_33_367#_M1022_g N_A_223_367#_c_577_n 0.00309738f $X=2.745 $Y=2.465
+ $X2=0 $Y2=0
cc_162 N_A_33_367#_M1022_g N_A_223_367#_c_578_n 8.25902e-19 $X=2.745 $Y=2.465
+ $X2=0 $Y2=0
cc_163 N_A_33_367#_M1009_g N_A_223_367#_c_579_n 0.00113216f $X=1.885 $Y=2.465
+ $X2=0 $Y2=0
cc_164 N_A_33_367#_M1016_g N_A_223_367#_c_579_n 0.00398489f $X=2.315 $Y=2.465
+ $X2=0 $Y2=0
cc_165 N_A_33_367#_M1022_g N_A_223_367#_c_579_n 4.53726e-19 $X=2.745 $Y=2.465
+ $X2=0 $Y2=0
cc_166 N_A_33_367#_M1000_g N_Y_c_666_n 0.00484678f $X=1.155 $Y=0.655 $X2=0 $Y2=0
cc_167 N_A_33_367#_c_164_n N_Y_c_666_n 0.0129322f $X=0.975 $Y=0.955 $X2=0 $Y2=0
cc_168 N_A_33_367#_M1000_g N_Y_c_658_n 0.00129003f $X=1.155 $Y=0.655 $X2=0 $Y2=0
cc_169 N_A_33_367#_c_164_n N_Y_c_658_n 4.37016e-19 $X=0.975 $Y=0.955 $X2=0 $Y2=0
cc_170 N_A_33_367#_c_146_n N_Y_c_658_n 0.0132161f $X=1.06 $Y=1.375 $X2=0 $Y2=0
cc_171 N_A_33_367#_c_219_p N_Y_c_658_n 0.0137165f $X=2.21 $Y=1.46 $X2=0 $Y2=0
cc_172 N_A_33_367#_c_149_n N_Y_c_658_n 0.00282613f $X=2.445 $Y=1.45 $X2=0 $Y2=0
cc_173 N_A_33_367#_M1009_g N_Y_c_662_n 0.0157024f $X=1.885 $Y=2.465 $X2=0 $Y2=0
cc_174 N_A_33_367#_M1016_g N_Y_c_662_n 0.018219f $X=2.315 $Y=2.465 $X2=0 $Y2=0
cc_175 N_A_33_367#_c_219_p N_Y_c_662_n 0.0447411f $X=2.21 $Y=1.46 $X2=0 $Y2=0
cc_176 N_A_33_367#_c_149_n N_Y_c_662_n 0.00293498f $X=2.445 $Y=1.45 $X2=0 $Y2=0
cc_177 N_A_33_367#_c_219_p N_Y_c_677_n 8.15674e-19 $X=2.21 $Y=1.46 $X2=0 $Y2=0
cc_178 N_A_33_367#_M1002_g N_Y_c_663_n 0.0170614f $X=1.455 $Y=2.465 $X2=0 $Y2=0
cc_179 N_A_33_367#_c_156_n N_Y_c_663_n 0.00911007f $X=0.975 $Y=2.005 $X2=0 $Y2=0
cc_180 N_A_33_367#_c_147_n N_Y_c_663_n 0.0104713f $X=1.085 $Y=1.92 $X2=0 $Y2=0
cc_181 N_A_33_367#_c_219_p N_Y_c_663_n 0.0208668f $X=2.21 $Y=1.46 $X2=0 $Y2=0
cc_182 N_A_33_367#_c_149_n N_Y_c_663_n 0.00299787f $X=2.445 $Y=1.45 $X2=0 $Y2=0
cc_183 N_A_33_367#_M1016_g Y 0.0021138f $X=2.315 $Y=2.465 $X2=0 $Y2=0
cc_184 N_A_33_367#_M1018_g Y 0.00668549f $X=2.445 $Y=0.655 $X2=0 $Y2=0
cc_185 N_A_33_367#_M1022_g Y 0.00226751f $X=2.745 $Y=2.465 $X2=0 $Y2=0
cc_186 N_A_33_367#_c_219_p Y 0.0136858f $X=2.21 $Y=1.46 $X2=0 $Y2=0
cc_187 N_A_33_367#_c_149_n Y 0.0162769f $X=2.445 $Y=1.45 $X2=0 $Y2=0
cc_188 N_A_33_367#_M1022_g Y 0.0217415f $X=2.745 $Y=2.465 $X2=0 $Y2=0
cc_189 N_A_33_367#_c_149_n Y 0.0021371f $X=2.445 $Y=1.45 $X2=0 $Y2=0
cc_190 N_A_33_367#_M1005_g N_Y_c_660_n 0.0142223f $X=1.585 $Y=0.655 $X2=0 $Y2=0
cc_191 N_A_33_367#_M1017_g N_Y_c_660_n 0.0137676f $X=2.015 $Y=0.655 $X2=0 $Y2=0
cc_192 N_A_33_367#_c_219_p N_Y_c_660_n 0.0640761f $X=2.21 $Y=1.46 $X2=0 $Y2=0
cc_193 N_A_33_367#_c_149_n N_Y_c_660_n 0.002964f $X=2.445 $Y=1.45 $X2=0 $Y2=0
cc_194 N_A_33_367#_M1018_g N_Y_c_661_n 0.0252189f $X=2.445 $Y=0.655 $X2=0 $Y2=0
cc_195 N_A_33_367#_c_149_n N_Y_c_661_n 0.00467596f $X=2.445 $Y=1.45 $X2=0 $Y2=0
cc_196 N_A_33_367#_c_164_n N_VGND_M1014_d 0.00726321f $X=0.975 $Y=0.955
+ $X2=-0.19 $Y2=-0.245
cc_197 N_A_33_367#_c_146_n N_VGND_M1014_d 4.01256e-19 $X=1.06 $Y=1.375 $X2=-0.19
+ $Y2=-0.245
cc_198 N_A_33_367#_M1000_g N_VGND_c_745_n 0.0113327f $X=1.155 $Y=0.655 $X2=0
+ $Y2=0
cc_199 N_A_33_367#_M1005_g N_VGND_c_745_n 8.61353e-19 $X=1.585 $Y=0.655 $X2=0
+ $Y2=0
cc_200 N_A_33_367#_c_164_n N_VGND_c_745_n 0.017018f $X=0.975 $Y=0.955 $X2=0
+ $Y2=0
cc_201 N_A_33_367#_M1000_g N_VGND_c_746_n 0.00486043f $X=1.155 $Y=0.655 $X2=0
+ $Y2=0
cc_202 N_A_33_367#_M1005_g N_VGND_c_746_n 0.00564095f $X=1.585 $Y=0.655 $X2=0
+ $Y2=0
cc_203 N_A_33_367#_M1000_g N_VGND_c_747_n 8.67983e-19 $X=1.155 $Y=0.655 $X2=0
+ $Y2=0
cc_204 N_A_33_367#_M1005_g N_VGND_c_747_n 0.00958615f $X=1.585 $Y=0.655 $X2=0
+ $Y2=0
cc_205 N_A_33_367#_M1017_g N_VGND_c_747_n 0.0105579f $X=2.015 $Y=0.655 $X2=0
+ $Y2=0
cc_206 N_A_33_367#_M1018_g N_VGND_c_747_n 6.59124e-19 $X=2.445 $Y=0.655 $X2=0
+ $Y2=0
cc_207 N_A_33_367#_c_144_n N_VGND_c_751_n 0.0185207f $X=0.49 $Y=0.42 $X2=0 $Y2=0
cc_208 N_A_33_367#_M1017_g N_VGND_c_756_n 0.00486043f $X=2.015 $Y=0.655 $X2=0
+ $Y2=0
cc_209 N_A_33_367#_M1018_g N_VGND_c_756_n 0.00433717f $X=2.445 $Y=0.655 $X2=0
+ $Y2=0
cc_210 N_A_33_367#_M1018_g N_VGND_c_757_n 0.00215947f $X=2.445 $Y=0.655 $X2=0
+ $Y2=0
cc_211 N_A_33_367#_M1014_s N_VGND_c_759_n 0.00302127f $X=0.365 $Y=0.235 $X2=0
+ $Y2=0
cc_212 N_A_33_367#_M1000_g N_VGND_c_759_n 0.00835506f $X=1.155 $Y=0.655 $X2=0
+ $Y2=0
cc_213 N_A_33_367#_M1005_g N_VGND_c_759_n 0.00959071f $X=1.585 $Y=0.655 $X2=0
+ $Y2=0
cc_214 N_A_33_367#_M1017_g N_VGND_c_759_n 0.00824727f $X=2.015 $Y=0.655 $X2=0
+ $Y2=0
cc_215 N_A_33_367#_M1018_g N_VGND_c_759_n 0.00642938f $X=2.445 $Y=0.655 $X2=0
+ $Y2=0
cc_216 N_A_33_367#_c_144_n N_VGND_c_759_n 0.010808f $X=0.49 $Y=0.42 $X2=0 $Y2=0
cc_217 N_A2_c_272_n N_A1_M1003_g 0.00120506f $X=3.172 $Y=1.16 $X2=0 $Y2=0
cc_218 N_A2_c_273_n N_A1_M1003_g 0.0216015f $X=3.195 $Y=1.35 $X2=0 $Y2=0
cc_219 N_A2_c_276_n N_A1_M1003_g 0.0336978f $X=3.195 $Y=1.185 $X2=0 $Y2=0
cc_220 N_A2_c_278_n N_A1_M1003_g 0.0101265f $X=5.335 $Y=1.295 $X2=0 $Y2=0
cc_221 N_A2_c_278_n N_A1_M1008_g 0.0105237f $X=5.335 $Y=1.295 $X2=0 $Y2=0
cc_222 N_A2_c_278_n N_A1_M1020_g 0.0105539f $X=5.335 $Y=1.295 $X2=0 $Y2=0
cc_223 N_A2_c_266_n N_A1_M1021_g 0.0259019f $X=5.365 $Y=1.185 $X2=0 $Y2=0
cc_224 A2 N_A1_M1021_g 0.0010397f $X=5.435 $Y=1.21 $X2=0 $Y2=0
cc_225 N_A2_c_278_n N_A1_M1021_g 0.0120038f $X=5.335 $Y=1.295 $X2=0 $Y2=0
cc_226 N_A2_M1011_g N_A1_M1024_g 0.0259019f $X=5.365 $Y=2.465 $X2=0 $Y2=0
cc_227 N_A2_M1001_g A1 0.00281783f $X=3.205 $Y=2.465 $X2=0 $Y2=0
cc_228 N_A2_c_272_n A1 0.00826557f $X=3.172 $Y=1.16 $X2=0 $Y2=0
cc_229 N_A2_c_273_n A1 6.64607e-19 $X=3.195 $Y=1.35 $X2=0 $Y2=0
cc_230 A2 A1 0.0087366f $X=5.435 $Y=1.21 $X2=0 $Y2=0
cc_231 N_A2_c_277_n A1 0.00625276f $X=6.28 $Y=1.35 $X2=0 $Y2=0
cc_232 N_A2_c_278_n A1 0.125162f $X=5.335 $Y=1.295 $X2=0 $Y2=0
cc_233 N_A2_M1001_g N_A1_c_382_n 0.0403046f $X=3.205 $Y=2.465 $X2=0 $Y2=0
cc_234 N_A2_c_277_n N_A1_c_382_n 0.0259019f $X=6.28 $Y=1.35 $X2=0 $Y2=0
cc_235 N_A2_c_278_n N_A1_c_382_n 0.00730626f $X=5.335 $Y=1.295 $X2=0 $Y2=0
cc_236 N_A2_M1001_g N_VPWR_c_488_n 0.00243873f $X=3.205 $Y=2.465 $X2=0 $Y2=0
cc_237 N_A2_M1001_g N_VPWR_c_457_n 0.0119987f $X=3.205 $Y=2.465 $X2=0 $Y2=0
cc_238 N_A2_M1011_g N_VPWR_c_458_n 0.0146917f $X=5.365 $Y=2.465 $X2=0 $Y2=0
cc_239 N_A2_M1013_g N_VPWR_c_458_n 6.80491e-19 $X=5.795 $Y=2.465 $X2=0 $Y2=0
cc_240 N_A2_M1011_g N_VPWR_c_459_n 7.39387e-19 $X=5.365 $Y=2.465 $X2=0 $Y2=0
cc_241 N_A2_M1013_g N_VPWR_c_459_n 0.0143508f $X=5.795 $Y=2.465 $X2=0 $Y2=0
cc_242 N_A2_M1025_g N_VPWR_c_459_n 0.0161027f $X=6.225 $Y=2.465 $X2=0 $Y2=0
cc_243 N_A2_M1001_g N_VPWR_c_460_n 0.00525069f $X=3.205 $Y=2.465 $X2=0 $Y2=0
cc_244 N_A2_M1011_g N_VPWR_c_464_n 0.00486043f $X=5.365 $Y=2.465 $X2=0 $Y2=0
cc_245 N_A2_M1013_g N_VPWR_c_464_n 0.00486043f $X=5.795 $Y=2.465 $X2=0 $Y2=0
cc_246 N_A2_M1025_g N_VPWR_c_465_n 0.00486043f $X=6.225 $Y=2.465 $X2=0 $Y2=0
cc_247 N_A2_M1001_g N_VPWR_c_455_n 0.00896134f $X=3.205 $Y=2.465 $X2=0 $Y2=0
cc_248 N_A2_M1011_g N_VPWR_c_455_n 0.00824727f $X=5.365 $Y=2.465 $X2=0 $Y2=0
cc_249 N_A2_M1013_g N_VPWR_c_455_n 0.00824727f $X=5.795 $Y=2.465 $X2=0 $Y2=0
cc_250 N_A2_M1025_g N_VPWR_c_455_n 0.00919827f $X=6.225 $Y=2.465 $X2=0 $Y2=0
cc_251 N_A2_M1001_g N_A_223_367#_c_582_n 0.0142506f $X=3.205 $Y=2.465 $X2=0
+ $Y2=0
cc_252 N_A2_c_272_n N_A_223_367#_c_582_n 0.00680714f $X=3.172 $Y=1.16 $X2=0
+ $Y2=0
cc_253 N_A2_c_273_n N_A_223_367#_c_582_n 8.34881e-19 $X=3.195 $Y=1.35 $X2=0
+ $Y2=0
cc_254 N_A2_c_278_n N_A_223_367#_c_582_n 0.00417719f $X=5.335 $Y=1.295 $X2=0
+ $Y2=0
cc_255 N_A2_c_272_n N_A_223_367#_c_578_n 0.00224645f $X=3.172 $Y=1.16 $X2=0
+ $Y2=0
cc_256 N_A2_c_273_n N_A_223_367#_c_578_n 3.55062e-19 $X=3.195 $Y=1.35 $X2=0
+ $Y2=0
cc_257 N_A2_M1011_g N_A_223_367#_c_588_n 0.00620501f $X=5.365 $Y=2.465 $X2=0
+ $Y2=0
cc_258 N_A2_c_278_n N_A_223_367#_c_588_n 0.00362077f $X=5.335 $Y=1.295 $X2=0
+ $Y2=0
cc_259 N_A2_M1013_g N_A_223_367#_c_561_n 0.0150775f $X=5.795 $Y=2.465 $X2=0
+ $Y2=0
cc_260 N_A2_M1025_g N_A_223_367#_c_561_n 0.0173007f $X=6.225 $Y=2.465 $X2=0
+ $Y2=0
cc_261 A2 N_A_223_367#_c_561_n 0.0734267f $X=6.395 $Y=1.21 $X2=0 $Y2=0
cc_262 N_A2_c_277_n N_A_223_367#_c_561_n 0.00560448f $X=6.28 $Y=1.35 $X2=0 $Y2=0
cc_263 N_A2_M1011_g N_A_223_367#_c_563_n 0.0151699f $X=5.365 $Y=2.465 $X2=0
+ $Y2=0
cc_264 N_A2_M1013_g N_A_223_367#_c_563_n 2.95608e-19 $X=5.795 $Y=2.465 $X2=0
+ $Y2=0
cc_265 A2 N_A_223_367#_c_563_n 0.0270977f $X=5.435 $Y=1.21 $X2=0 $Y2=0
cc_266 N_A2_c_277_n N_A_223_367#_c_563_n 0.00232957f $X=6.28 $Y=1.35 $X2=0 $Y2=0
cc_267 N_A2_c_272_n N_Y_c_696_n 0.0178722f $X=3.172 $Y=1.16 $X2=0 $Y2=0
cc_268 N_A2_c_273_n N_Y_c_696_n 6.57528e-19 $X=3.195 $Y=1.35 $X2=0 $Y2=0
cc_269 N_A2_c_276_n N_Y_c_696_n 0.0145231f $X=3.195 $Y=1.185 $X2=0 $Y2=0
cc_270 N_A2_c_278_n N_Y_c_696_n 0.0942903f $X=5.335 $Y=1.295 $X2=0 $Y2=0
cc_271 N_A2_M1001_g Y 0.00189296f $X=3.205 $Y=2.465 $X2=0 $Y2=0
cc_272 N_A2_c_272_n Y 0.0241844f $X=3.172 $Y=1.16 $X2=0 $Y2=0
cc_273 N_A2_c_273_n Y 0.00263941f $X=3.195 $Y=1.35 $X2=0 $Y2=0
cc_274 N_A2_M1001_g Y 0.00130782f $X=3.205 $Y=2.465 $X2=0 $Y2=0
cc_275 N_A2_c_272_n N_Y_c_661_n 0.0112153f $X=3.172 $Y=1.16 $X2=0 $Y2=0
cc_276 N_A2_c_276_n N_Y_c_661_n 0.0052476f $X=3.195 $Y=1.185 $X2=0 $Y2=0
cc_277 N_A2_c_272_n N_VGND_M1018_d 0.00122233f $X=3.172 $Y=1.16 $X2=0 $Y2=0
cc_278 N_A2_c_266_n N_VGND_c_748_n 0.00285858f $X=5.365 $Y=1.185 $X2=0 $Y2=0
cc_279 N_A2_c_268_n N_VGND_c_748_n 0.00162573f $X=5.795 $Y=1.185 $X2=0 $Y2=0
cc_280 N_A2_c_270_n N_VGND_c_750_n 0.0055868f $X=6.225 $Y=1.185 $X2=0 $Y2=0
cc_281 A2 N_VGND_c_750_n 0.0229011f $X=6.395 $Y=1.21 $X2=0 $Y2=0
cc_282 N_A2_c_277_n N_VGND_c_750_n 0.00317373f $X=6.28 $Y=1.35 $X2=0 $Y2=0
cc_283 N_A2_c_266_n N_VGND_c_753_n 0.00425616f $X=5.365 $Y=1.185 $X2=0 $Y2=0
cc_284 N_A2_c_276_n N_VGND_c_753_n 0.00421077f $X=3.195 $Y=1.185 $X2=0 $Y2=0
cc_285 N_A2_c_268_n N_VGND_c_754_n 0.00439206f $X=5.795 $Y=1.185 $X2=0 $Y2=0
cc_286 N_A2_c_270_n N_VGND_c_754_n 0.00585385f $X=6.225 $Y=1.185 $X2=0 $Y2=0
cc_287 N_A2_c_276_n N_VGND_c_757_n 0.0035885f $X=3.195 $Y=1.185 $X2=0 $Y2=0
cc_288 N_A2_c_266_n N_VGND_c_759_n 0.00586053f $X=5.365 $Y=1.185 $X2=0 $Y2=0
cc_289 N_A2_c_268_n N_VGND_c_759_n 0.00586174f $X=5.795 $Y=1.185 $X2=0 $Y2=0
cc_290 N_A2_c_270_n N_VGND_c_759_n 0.0114597f $X=6.225 $Y=1.185 $X2=0 $Y2=0
cc_291 N_A2_c_276_n N_VGND_c_759_n 0.00641677f $X=3.195 $Y=1.185 $X2=0 $Y2=0
cc_292 N_A2_c_272_n N_A_658_47#_M1004_s 2.69137e-19 $X=3.172 $Y=1.16 $X2=-0.19
+ $Y2=-0.245
cc_293 N_A2_c_276_n N_A_658_47#_c_840_n 0.00340138f $X=3.195 $Y=1.185 $X2=0
+ $Y2=0
cc_294 N_A2_c_278_n N_A_658_47#_c_840_n 0.004087f $X=5.335 $Y=1.295 $X2=0 $Y2=0
cc_295 N_A2_c_266_n N_A_658_47#_c_842_n 0.00294618f $X=5.365 $Y=1.185 $X2=0
+ $Y2=0
cc_296 N_A2_c_266_n N_A_658_47#_c_843_n 0.00418274f $X=5.365 $Y=1.185 $X2=0
+ $Y2=0
cc_297 N_A2_c_268_n N_A_658_47#_c_843_n 4.55047e-19 $X=5.795 $Y=1.185 $X2=0
+ $Y2=0
cc_298 N_A2_c_278_n N_A_658_47#_c_843_n 0.0181409f $X=5.335 $Y=1.295 $X2=0 $Y2=0
cc_299 N_A2_c_266_n N_A_658_47#_c_846_n 0.00879064f $X=5.365 $Y=1.185 $X2=0
+ $Y2=0
cc_300 N_A2_c_268_n N_A_658_47#_c_846_n 0.010928f $X=5.795 $Y=1.185 $X2=0 $Y2=0
cc_301 A2 N_A_658_47#_c_846_n 0.0110149f $X=6.395 $Y=1.21 $X2=0 $Y2=0
cc_302 N_A2_c_277_n N_A_658_47#_c_846_n 9.24773e-19 $X=6.28 $Y=1.35 $X2=0 $Y2=0
cc_303 N_A2_c_278_n N_A_658_47#_c_846_n 0.0200607f $X=5.335 $Y=1.295 $X2=0 $Y2=0
cc_304 A2 N_A_658_47#_c_851_n 0.0160173f $X=6.395 $Y=1.21 $X2=0 $Y2=0
cc_305 N_A2_c_277_n N_A_658_47#_c_851_n 0.00240082f $X=6.28 $Y=1.35 $X2=0 $Y2=0
cc_306 N_A1_M1006_g N_VPWR_c_488_n 8.78991e-19 $X=3.645 $Y=2.465 $X2=0 $Y2=0
cc_307 N_A1_M1006_g N_VPWR_c_457_n 0.0141507f $X=3.645 $Y=2.465 $X2=0 $Y2=0
cc_308 N_A1_M1012_g N_VPWR_c_457_n 0.0020759f $X=4.075 $Y=2.465 $X2=0 $Y2=0
cc_309 N_A1_M1006_g N_VPWR_c_506_n 0.0103094f $X=3.645 $Y=2.465 $X2=0 $Y2=0
cc_310 N_A1_M1012_g N_VPWR_c_506_n 0.0101831f $X=4.075 $Y=2.465 $X2=0 $Y2=0
cc_311 N_A1_M1019_g N_VPWR_c_506_n 0.00303044f $X=4.505 $Y=2.465 $X2=0 $Y2=0
cc_312 N_A1_M1019_g N_VPWR_c_458_n 0.0012362f $X=4.505 $Y=2.465 $X2=0 $Y2=0
cc_313 N_A1_M1024_g N_VPWR_c_458_n 0.015933f $X=4.935 $Y=2.465 $X2=0 $Y2=0
cc_314 N_A1_M1006_g N_VPWR_c_463_n 0.00486043f $X=3.645 $Y=2.465 $X2=0 $Y2=0
cc_315 N_A1_M1012_g N_VPWR_c_463_n 0.00359964f $X=4.075 $Y=2.465 $X2=0 $Y2=0
cc_316 N_A1_M1019_g N_VPWR_c_463_n 0.00359964f $X=4.505 $Y=2.465 $X2=0 $Y2=0
cc_317 N_A1_M1024_g N_VPWR_c_463_n 0.00486043f $X=4.935 $Y=2.465 $X2=0 $Y2=0
cc_318 N_A1_M1006_g N_VPWR_c_455_n 0.00459245f $X=3.645 $Y=2.465 $X2=0 $Y2=0
cc_319 N_A1_M1012_g N_VPWR_c_455_n 0.00542362f $X=4.075 $Y=2.465 $X2=0 $Y2=0
cc_320 N_A1_M1019_g N_VPWR_c_455_n 0.00535287f $X=4.505 $Y=2.465 $X2=0 $Y2=0
cc_321 N_A1_M1024_g N_VPWR_c_455_n 0.00824727f $X=4.935 $Y=2.465 $X2=0 $Y2=0
cc_322 N_A1_M1006_g N_A_223_367#_c_582_n 0.0105035f $X=3.645 $Y=2.465 $X2=0
+ $Y2=0
cc_323 N_A1_M1012_g N_A_223_367#_c_582_n 0.0104926f $X=4.075 $Y=2.465 $X2=0
+ $Y2=0
cc_324 N_A1_M1019_g N_A_223_367#_c_582_n 0.00997577f $X=4.505 $Y=2.465 $X2=0
+ $Y2=0
cc_325 A1 N_A_223_367#_c_582_n 0.0740081f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_326 N_A1_c_382_n N_A_223_367#_c_582_n 0.00115661f $X=4.935 $Y=1.51 $X2=0
+ $Y2=0
cc_327 N_A1_M1012_g N_A_223_367#_c_603_n 0.0140695f $X=4.075 $Y=2.465 $X2=0
+ $Y2=0
cc_328 N_A1_M1019_g N_A_223_367#_c_603_n 0.0152575f $X=4.505 $Y=2.465 $X2=0
+ $Y2=0
cc_329 N_A1_M1024_g N_A_223_367#_c_588_n 0.0122129f $X=4.935 $Y=2.465 $X2=0
+ $Y2=0
cc_330 A1 N_A_223_367#_c_588_n 0.022596f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_331 A1 N_A_223_367#_c_607_n 0.0154121f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_332 N_A1_c_382_n N_A_223_367#_c_607_n 6.52992e-19 $X=4.935 $Y=1.51 $X2=0
+ $Y2=0
cc_333 N_A1_M1024_g N_A_223_367#_c_563_n 0.00113534f $X=4.935 $Y=2.465 $X2=0
+ $Y2=0
cc_334 A1 N_A_223_367#_c_563_n 0.00539698f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_335 N_A1_M1003_g N_Y_c_696_n 0.00924124f $X=3.645 $Y=0.655 $X2=0 $Y2=0
cc_336 N_A1_M1008_g N_Y_c_696_n 0.00929613f $X=4.075 $Y=0.655 $X2=0 $Y2=0
cc_337 N_A1_M1020_g N_Y_c_696_n 0.00929613f $X=4.505 $Y=0.655 $X2=0 $Y2=0
cc_338 N_A1_M1021_g N_Y_c_696_n 0.0026751f $X=4.935 $Y=0.655 $X2=0 $Y2=0
cc_339 A1 Y 0.00700835f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_340 A1 Y 0.00126545f $X=4.955 $Y=1.58 $X2=0 $Y2=0
cc_341 N_A1_M1003_g N_VGND_c_753_n 0.00357877f $X=3.645 $Y=0.655 $X2=0 $Y2=0
cc_342 N_A1_M1008_g N_VGND_c_753_n 0.00357877f $X=4.075 $Y=0.655 $X2=0 $Y2=0
cc_343 N_A1_M1020_g N_VGND_c_753_n 0.00357877f $X=4.505 $Y=0.655 $X2=0 $Y2=0
cc_344 N_A1_M1021_g N_VGND_c_753_n 0.00357877f $X=4.935 $Y=0.655 $X2=0 $Y2=0
cc_345 N_A1_M1003_g N_VGND_c_759_n 0.00537654f $X=3.645 $Y=0.655 $X2=0 $Y2=0
cc_346 N_A1_M1008_g N_VGND_c_759_n 0.0053512f $X=4.075 $Y=0.655 $X2=0 $Y2=0
cc_347 N_A1_M1020_g N_VGND_c_759_n 0.0053512f $X=4.505 $Y=0.655 $X2=0 $Y2=0
cc_348 N_A1_M1021_g N_VGND_c_759_n 0.00537654f $X=4.935 $Y=0.655 $X2=0 $Y2=0
cc_349 N_A1_M1003_g N_A_658_47#_c_840_n 0.0103254f $X=3.645 $Y=0.655 $X2=0 $Y2=0
cc_350 N_A1_M1008_g N_A_658_47#_c_840_n 0.0103254f $X=4.075 $Y=0.655 $X2=0 $Y2=0
cc_351 N_A1_M1020_g N_A_658_47#_c_840_n 0.0103254f $X=4.505 $Y=0.655 $X2=0 $Y2=0
cc_352 N_A1_M1021_g N_A_658_47#_c_840_n 0.0118957f $X=4.935 $Y=0.655 $X2=0 $Y2=0
cc_353 N_VPWR_c_455_n N_A_223_367#_M1002_d 0.00215161f $X=6.48 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_354 N_VPWR_c_455_n N_A_223_367#_M1009_d 0.00223559f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_355 N_VPWR_c_455_n N_A_223_367#_M1022_d 0.00365966f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_356 N_VPWR_c_506_n N_A_223_367#_M1006_s 0.0034524f $X=4.29 $Y=2.375 $X2=0
+ $Y2=0
cc_357 N_VPWR_c_455_n N_A_223_367#_M1006_s 0.00254929f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_358 N_VPWR_c_455_n N_A_223_367#_M1019_s 0.00376849f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_359 N_VPWR_c_455_n N_A_223_367#_M1011_d 0.00571434f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_360 N_VPWR_c_455_n N_A_223_367#_M1025_d 0.00371702f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_361 N_VPWR_c_456_n N_A_223_367#_c_559_n 0.0335235f $X=0.72 $Y=2.345 $X2=0
+ $Y2=0
cc_362 N_VPWR_c_460_n N_A_223_367#_c_559_n 0.0179183f $X=3.265 $Y=3.33 $X2=0
+ $Y2=0
cc_363 N_VPWR_c_455_n N_A_223_367#_c_559_n 0.0101082f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_364 N_VPWR_c_456_n N_A_223_367#_c_560_n 0.0305961f $X=0.72 $Y=2.345 $X2=0
+ $Y2=0
cc_365 N_VPWR_c_460_n N_A_223_367#_c_570_n 0.0346841f $X=3.265 $Y=3.33 $X2=0
+ $Y2=0
cc_366 N_VPWR_c_455_n N_A_223_367#_c_570_n 0.0216765f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_367 N_VPWR_c_460_n N_A_223_367#_c_575_n 0.035191f $X=3.265 $Y=3.33 $X2=0
+ $Y2=0
cc_368 N_VPWR_c_455_n N_A_223_367#_c_575_n 0.0225315f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_369 N_VPWR_c_460_n N_A_223_367#_c_627_n 0.0132962f $X=3.265 $Y=3.33 $X2=0
+ $Y2=0
cc_370 N_VPWR_c_455_n N_A_223_367#_c_627_n 0.00777554f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_371 N_VPWR_M1001_s N_A_223_367#_c_582_n 0.00519998f $X=3.28 $Y=1.835 $X2=0
+ $Y2=0
cc_372 N_VPWR_M1012_d N_A_223_367#_c_582_n 0.00333266f $X=4.15 $Y=1.835 $X2=0
+ $Y2=0
cc_373 N_VPWR_c_488_n N_A_223_367#_c_582_n 0.0172819f $X=3.43 $Y=2.495 $X2=0
+ $Y2=0
cc_374 N_VPWR_c_506_n N_A_223_367#_c_582_n 0.0454597f $X=4.29 $Y=2.375 $X2=0
+ $Y2=0
cc_375 N_VPWR_M1012_d N_A_223_367#_c_603_n 0.00345221f $X=4.15 $Y=1.835 $X2=0
+ $Y2=0
cc_376 N_VPWR_c_506_n N_A_223_367#_c_603_n 0.0382912f $X=4.29 $Y=2.375 $X2=0
+ $Y2=0
cc_377 N_VPWR_c_463_n N_A_223_367#_c_603_n 0.0469096f $X=4.985 $Y=3.33 $X2=0
+ $Y2=0
cc_378 N_VPWR_c_455_n N_A_223_367#_c_603_n 0.031338f $X=6.48 $Y=3.33 $X2=0 $Y2=0
cc_379 N_VPWR_c_463_n N_A_223_367#_c_637_n 0.0117708f $X=4.985 $Y=3.33 $X2=0
+ $Y2=0
cc_380 N_VPWR_c_455_n N_A_223_367#_c_637_n 0.0073517f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_381 N_VPWR_M1024_d N_A_223_367#_c_588_n 0.00424963f $X=5.01 $Y=1.835 $X2=0
+ $Y2=0
cc_382 N_VPWR_c_458_n N_A_223_367#_c_588_n 0.0170777f $X=5.15 $Y=2.375 $X2=0
+ $Y2=0
cc_383 N_VPWR_c_464_n N_A_223_367#_c_641_n 0.0120977f $X=5.845 $Y=3.33 $X2=0
+ $Y2=0
cc_384 N_VPWR_c_455_n N_A_223_367#_c_641_n 0.00691495f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_385 N_VPWR_M1013_s N_A_223_367#_c_561_n 0.00182684f $X=5.87 $Y=1.835 $X2=0
+ $Y2=0
cc_386 N_VPWR_c_459_n N_A_223_367#_c_561_n 0.016744f $X=6.01 $Y=2.19 $X2=0 $Y2=0
cc_387 N_VPWR_c_465_n N_A_223_367#_c_562_n 0.0178111f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_388 N_VPWR_c_455_n N_A_223_367#_c_562_n 0.0100304f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_389 N_VPWR_c_460_n N_A_223_367#_c_579_n 0.01906f $X=3.265 $Y=3.33 $X2=0 $Y2=0
cc_390 N_VPWR_c_455_n N_A_223_367#_c_579_n 0.0124545f $X=6.48 $Y=3.33 $X2=0
+ $Y2=0
cc_391 N_VPWR_c_455_n N_Y_M1002_s 0.00225186f $X=6.48 $Y=3.33 $X2=0 $Y2=0
cc_392 N_VPWR_c_455_n N_Y_M1016_s 0.00225186f $X=6.48 $Y=3.33 $X2=0 $Y2=0
cc_393 N_A_223_367#_c_570_n N_Y_M1002_s 0.00345885f $X=1.935 $Y=2.87 $X2=0 $Y2=0
cc_394 N_A_223_367#_c_575_n N_Y_M1016_s 0.00335895f $X=2.895 $Y=2.955 $X2=0
+ $Y2=0
cc_395 N_A_223_367#_M1009_d N_Y_c_662_n 0.0017993f $X=1.96 $Y=1.835 $X2=0 $Y2=0
cc_396 N_A_223_367#_c_570_n N_Y_c_662_n 0.0031796f $X=1.935 $Y=2.87 $X2=0 $Y2=0
cc_397 N_A_223_367#_c_572_n N_Y_c_662_n 0.0178454f $X=2.1 $Y=2.29 $X2=0 $Y2=0
cc_398 N_A_223_367#_c_570_n N_Y_c_663_n 0.0151158f $X=1.935 $Y=2.87 $X2=0 $Y2=0
cc_399 N_A_223_367#_c_575_n Y 0.0170993f $X=2.895 $Y=2.955 $X2=0 $Y2=0
cc_400 N_A_223_367#_c_577_n Y 0.042511f $X=2.99 $Y=2.16 $X2=0 $Y2=0
cc_401 N_A_223_367#_c_578_n Y 0.0145156f $X=3.095 $Y=2.005 $X2=0 $Y2=0
cc_402 N_Y_c_660_n N_VGND_M1005_d 0.00176461f $X=2.135 $Y=0.95 $X2=0 $Y2=0
cc_403 N_Y_c_696_n N_VGND_M1018_d 0.0104757f $X=4.72 $Y=0.79 $X2=0 $Y2=0
cc_404 N_Y_c_661_n N_VGND_M1018_d 0.00903703f $X=2.86 $Y=0.95 $X2=0 $Y2=0
cc_405 N_Y_c_677_n N_VGND_c_746_n 0.00750381f $X=1.37 $Y=0.535 $X2=0 $Y2=0
cc_406 N_Y_c_660_n N_VGND_c_747_n 0.0155542f $X=2.135 $Y=0.95 $X2=0 $Y2=0
cc_407 N_Y_c_696_n N_VGND_c_753_n 0.00216965f $X=4.72 $Y=0.79 $X2=0 $Y2=0
cc_408 N_Y_c_729_p N_VGND_c_756_n 0.0135102f $X=2.23 $Y=0.42 $X2=0 $Y2=0
cc_409 N_Y_c_661_n N_VGND_c_756_n 0.0024769f $X=2.86 $Y=0.95 $X2=0 $Y2=0
cc_410 N_Y_c_661_n N_VGND_c_757_n 0.0408876f $X=2.86 $Y=0.95 $X2=0 $Y2=0
cc_411 N_Y_M1000_s N_VGND_c_759_n 0.0048535f $X=1.23 $Y=0.235 $X2=0 $Y2=0
cc_412 N_Y_M1017_s N_VGND_c_759_n 0.00378052f $X=2.09 $Y=0.235 $X2=0 $Y2=0
cc_413 N_Y_M1003_s N_VGND_c_759_n 0.00225186f $X=3.72 $Y=0.235 $X2=0 $Y2=0
cc_414 N_Y_M1020_s N_VGND_c_759_n 0.00225186f $X=4.58 $Y=0.235 $X2=0 $Y2=0
cc_415 N_Y_c_729_p N_VGND_c_759_n 0.00876635f $X=2.23 $Y=0.42 $X2=0 $Y2=0
cc_416 N_Y_c_696_n N_VGND_c_759_n 0.00675786f $X=4.72 $Y=0.79 $X2=0 $Y2=0
cc_417 N_Y_c_677_n N_VGND_c_759_n 0.00755479f $X=1.37 $Y=0.535 $X2=0 $Y2=0
cc_418 N_Y_c_661_n N_VGND_c_759_n 0.00646558f $X=2.86 $Y=0.95 $X2=0 $Y2=0
cc_419 N_Y_c_696_n N_A_658_47#_M1004_s 0.00352135f $X=4.72 $Y=0.79 $X2=-0.19
+ $Y2=-0.245
cc_420 N_Y_c_696_n N_A_658_47#_M1008_d 0.00340729f $X=4.72 $Y=0.79 $X2=0 $Y2=0
cc_421 N_Y_M1003_s N_A_658_47#_c_840_n 0.00337551f $X=3.72 $Y=0.235 $X2=0 $Y2=0
cc_422 N_Y_M1020_s N_A_658_47#_c_840_n 0.00337551f $X=4.58 $Y=0.235 $X2=0 $Y2=0
cc_423 N_Y_c_696_n N_A_658_47#_c_840_n 0.0822888f $X=4.72 $Y=0.79 $X2=0 $Y2=0
cc_424 N_VGND_c_759_n N_A_658_47#_M1004_s 0.00223577f $X=6.48 $Y=0 $X2=-0.19
+ $Y2=-0.245
cc_425 N_VGND_c_759_n N_A_658_47#_M1008_d 0.00223577f $X=6.48 $Y=0 $X2=0 $Y2=0
cc_426 N_VGND_c_759_n N_A_658_47#_M1021_d 0.00223562f $X=6.48 $Y=0 $X2=0 $Y2=0
cc_427 N_VGND_c_759_n N_A_658_47#_M1015_s 0.0028202f $X=6.48 $Y=0 $X2=0 $Y2=0
cc_428 N_VGND_c_753_n N_A_658_47#_c_840_n 0.100607f $X=5.485 $Y=0 $X2=0 $Y2=0
cc_429 N_VGND_c_759_n N_A_658_47#_c_840_n 0.0647738f $X=6.48 $Y=0 $X2=0 $Y2=0
cc_430 N_VGND_c_753_n N_A_658_47#_c_842_n 0.0157478f $X=5.485 $Y=0 $X2=0 $Y2=0
cc_431 N_VGND_c_759_n N_A_658_47#_c_842_n 0.00990873f $X=6.48 $Y=0 $X2=0 $Y2=0
cc_432 N_VGND_M1010_d N_A_658_47#_c_846_n 0.00346687f $X=5.44 $Y=0.235 $X2=0
+ $Y2=0
cc_433 N_VGND_c_748_n N_A_658_47#_c_846_n 0.0130182f $X=5.58 $Y=0.4 $X2=0 $Y2=0
cc_434 N_VGND_c_753_n N_A_658_47#_c_846_n 0.00196209f $X=5.485 $Y=0 $X2=0 $Y2=0
cc_435 N_VGND_c_754_n N_A_658_47#_c_846_n 0.00210007f $X=6.305 $Y=0 $X2=0 $Y2=0
cc_436 N_VGND_c_759_n N_A_658_47#_c_846_n 0.00833451f $X=6.48 $Y=0 $X2=0 $Y2=0
cc_437 N_VGND_c_754_n N_A_658_47#_c_875_n 0.0145813f $X=6.305 $Y=0 $X2=0 $Y2=0
cc_438 N_VGND_c_759_n N_A_658_47#_c_875_n 0.00964079f $X=6.48 $Y=0 $X2=0 $Y2=0
