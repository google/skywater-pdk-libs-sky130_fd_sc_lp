* File: sky130_fd_sc_lp__nand3_m.pxi.spice
* Created: Wed Sep  2 10:04:37 2020
* 
x_PM_SKY130_FD_SC_LP__NAND3_M%C N_C_c_44_n N_C_M1001_g N_C_M1000_g N_C_c_46_n
+ N_C_c_47_n N_C_c_52_n C C C C N_C_c_49_n PM_SKY130_FD_SC_LP__NAND3_M%C
x_PM_SKY130_FD_SC_LP__NAND3_M%B N_B_M1004_g N_B_M1003_g B B B N_B_c_83_n
+ PM_SKY130_FD_SC_LP__NAND3_M%B
x_PM_SKY130_FD_SC_LP__NAND3_M%A N_A_M1005_g N_A_M1002_g N_A_c_120_n N_A_c_121_n
+ A A A N_A_c_123_n PM_SKY130_FD_SC_LP__NAND3_M%A
x_PM_SKY130_FD_SC_LP__NAND3_M%VPWR N_VPWR_M1001_s N_VPWR_M1003_d N_VPWR_c_153_n
+ N_VPWR_c_154_n N_VPWR_c_155_n N_VPWR_c_156_n N_VPWR_c_157_n VPWR
+ N_VPWR_c_158_n N_VPWR_c_152_n PM_SKY130_FD_SC_LP__NAND3_M%VPWR
x_PM_SKY130_FD_SC_LP__NAND3_M%Y N_Y_M1005_d N_Y_M1001_d N_Y_M1002_d N_Y_c_179_n
+ Y Y Y N_Y_c_183_n N_Y_c_184_n N_Y_c_185_n PM_SKY130_FD_SC_LP__NAND3_M%Y
x_PM_SKY130_FD_SC_LP__NAND3_M%VGND N_VGND_M1000_s N_VGND_c_218_n N_VGND_c_219_n
+ VGND N_VGND_c_220_n N_VGND_c_221_n PM_SKY130_FD_SC_LP__NAND3_M%VGND
cc_1 VNB N_C_c_44_n 0.00968547f $X=-0.19 $Y=-0.245 $X2=0.36 $Y2=1.77
cc_2 VNB N_C_M1000_g 0.0271117f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.445
cc_3 VNB N_C_c_46_n 0.0364702f $X=-0.19 $Y=-0.245 $X2=0.345 $Y2=0.99
cc_4 VNB N_C_c_47_n 0.0236201f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.51
cc_5 VNB C 0.00741547f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_6 VNB N_C_c_49_n 0.0377822f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.005
cc_7 VNB N_B_M1004_g 0.0371034f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=1.92
cc_8 VNB N_B_M1003_g 0.0065655f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.84
cc_9 VNB B 0.00977786f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.445
cc_10 VNB N_B_c_83_n 0.0319905f $X=-0.19 $Y=-0.245 $X2=0.36 $Y2=1.845
cc_11 VNB N_A_M1005_g 0.0237277f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=1.92
cc_12 VNB N_A_M1002_g 0.00834029f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=0.84
cc_13 VNB N_A_c_120_n 0.0234523f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=0.99
cc_14 VNB N_A_c_121_n 0.0166897f $X=-0.19 $Y=-0.245 $X2=0.345 $Y2=0.84
cc_15 VNB A 0.00940341f $X=-0.19 $Y=-0.245 $X2=0.345 $Y2=0.99
cc_16 VNB N_A_c_123_n 0.0165521f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_17 VNB N_VPWR_c_152_n 0.0840719f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_Y_c_179_n 0.0117597f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB Y 0.0493865f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_VGND_c_218_n 0.0114503f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=2.52
cc_21 VNB N_VGND_c_219_n 0.0127275f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_VGND_c_220_n 0.0442298f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.51
cc_23 VNB N_VGND_c_221_n 0.130556f $X=-0.19 $Y=-0.245 $X2=0.36 $Y2=1.845
cc_24 VPB N_C_c_44_n 0.00776977f $X=-0.19 $Y=1.655 $X2=0.36 $Y2=1.77
cc_25 VPB N_C_M1001_g 0.0383356f $X=-0.19 $Y=1.655 $X2=0.5 $Y2=2.52
cc_26 VPB N_C_c_52_n 0.0245949f $X=-0.19 $Y=1.655 $X2=0.5 $Y2=1.845
cc_27 VPB C 0.0205076f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_28 VPB N_B_M1003_g 0.0449759f $X=-0.19 $Y=1.655 $X2=0.51 $Y2=0.84
cc_29 VPB B 0.00292132f $X=-0.19 $Y=1.655 $X2=0.51 $Y2=0.445
cc_30 VPB N_A_M1002_g 0.0524995f $X=-0.19 $Y=1.655 $X2=0.51 $Y2=0.84
cc_31 VPB A 0.00345348f $X=-0.19 $Y=1.655 $X2=0.345 $Y2=0.99
cc_32 VPB N_VPWR_c_153_n 0.0119561f $X=-0.19 $Y=1.655 $X2=0.51 $Y2=0.84
cc_33 VPB N_VPWR_c_154_n 0.0268267f $X=-0.19 $Y=1.655 $X2=0.51 $Y2=0.445
cc_34 VPB N_VPWR_c_155_n 0.0231558f $X=-0.19 $Y=1.655 $X2=0.345 $Y2=0.99
cc_35 VPB N_VPWR_c_156_n 0.0196081f $X=-0.19 $Y=1.655 $X2=0.36 $Y2=1.845
cc_36 VPB N_VPWR_c_157_n 0.00401341f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_37 VPB N_VPWR_c_158_n 0.0217943f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_38 VPB N_VPWR_c_152_n 0.0698947f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_39 VPB Y 0.00407097f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.51
cc_40 VPB Y 0.0278176f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_41 VPB N_Y_c_183_n 0.0125568f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_42 VPB N_Y_c_184_n 0.00657466f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.005
cc_43 VPB N_Y_c_185_n 0.032447f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_44 N_C_M1000_g N_B_M1004_g 0.049849f $X=0.51 $Y=0.445 $X2=0 $Y2=0
cc_45 C N_B_M1004_g 2.95886e-19 $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_46 N_C_c_49_n N_B_M1004_g 0.00565872f $X=0.27 $Y=1.005 $X2=0 $Y2=0
cc_47 N_C_c_44_n N_B_M1003_g 0.00560455f $X=0.36 $Y=1.77 $X2=0 $Y2=0
cc_48 N_C_c_52_n N_B_M1003_g 0.0285379f $X=0.5 $Y=1.845 $X2=0 $Y2=0
cc_49 C N_B_M1003_g 9.08905e-19 $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_50 N_C_c_46_n B 0.00147008f $X=0.345 $Y=0.99 $X2=0 $Y2=0
cc_51 C B 0.0473869f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_52 N_C_c_49_n B 0.00590534f $X=0.27 $Y=1.005 $X2=0 $Y2=0
cc_53 C N_B_c_83_n 3.51773e-19 $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_54 N_C_c_49_n N_B_c_83_n 0.0173752f $X=0.27 $Y=1.005 $X2=0 $Y2=0
cc_55 N_C_M1001_g N_VPWR_c_154_n 0.00452747f $X=0.5 $Y=2.52 $X2=0 $Y2=0
cc_56 N_C_c_52_n N_VPWR_c_154_n 0.00169694f $X=0.5 $Y=1.845 $X2=0 $Y2=0
cc_57 C N_VPWR_c_154_n 0.0155616f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_58 N_C_M1001_g N_VPWR_c_156_n 0.00428744f $X=0.5 $Y=2.52 $X2=0 $Y2=0
cc_59 N_C_M1001_g N_VPWR_c_152_n 0.00476395f $X=0.5 $Y=2.52 $X2=0 $Y2=0
cc_60 N_C_M1001_g Y 0.0017351f $X=0.5 $Y=2.52 $X2=0 $Y2=0
cc_61 C Y 0.0109123f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_62 N_C_M1001_g N_Y_c_184_n 0.00485489f $X=0.5 $Y=2.52 $X2=0 $Y2=0
cc_63 N_C_M1000_g N_VGND_c_219_n 0.0114059f $X=0.51 $Y=0.445 $X2=0 $Y2=0
cc_64 N_C_c_46_n N_VGND_c_219_n 0.0043931f $X=0.345 $Y=0.99 $X2=0 $Y2=0
cc_65 C N_VGND_c_219_n 0.00860018f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_66 N_C_M1000_g N_VGND_c_220_n 0.00486043f $X=0.51 $Y=0.445 $X2=0 $Y2=0
cc_67 N_C_M1000_g N_VGND_c_221_n 0.00827383f $X=0.51 $Y=0.445 $X2=0 $Y2=0
cc_68 N_C_c_46_n N_VGND_c_221_n 6.57488e-19 $X=0.345 $Y=0.99 $X2=0 $Y2=0
cc_69 C N_VGND_c_221_n 9.40005e-19 $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_70 N_B_M1004_g N_A_M1005_g 0.0593139f $X=0.9 $Y=0.445 $X2=0 $Y2=0
cc_71 B N_A_M1002_g 2.0812e-19 $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_72 N_B_c_83_n N_A_M1002_g 0.0402462f $X=0.84 $Y=1.365 $X2=0 $Y2=0
cc_73 N_B_c_83_n N_A_c_120_n 0.0191949f $X=0.84 $Y=1.365 $X2=0 $Y2=0
cc_74 N_B_M1004_g A 0.00220429f $X=0.9 $Y=0.445 $X2=0 $Y2=0
cc_75 B A 0.0658797f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_76 N_B_c_83_n A 0.00377198f $X=0.84 $Y=1.365 $X2=0 $Y2=0
cc_77 B N_A_c_123_n 6.36138e-19 $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_78 N_B_M1003_g N_VPWR_c_155_n 0.00194442f $X=0.93 $Y=2.52 $X2=0 $Y2=0
cc_79 N_B_M1003_g N_VPWR_c_156_n 0.00428744f $X=0.93 $Y=2.52 $X2=0 $Y2=0
cc_80 N_B_M1003_g N_VPWR_c_152_n 0.00476395f $X=0.93 $Y=2.52 $X2=0 $Y2=0
cc_81 N_B_M1004_g N_Y_c_179_n 0.0010274f $X=0.9 $Y=0.445 $X2=0 $Y2=0
cc_82 B Y 0.0153605f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_83 N_B_c_83_n Y 7.03267e-19 $X=0.84 $Y=1.365 $X2=0 $Y2=0
cc_84 N_B_M1003_g N_Y_c_183_n 0.017164f $X=0.93 $Y=2.52 $X2=0 $Y2=0
cc_85 B N_Y_c_183_n 0.00721341f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_86 N_B_M1003_g N_Y_c_184_n 0.00276293f $X=0.93 $Y=2.52 $X2=0 $Y2=0
cc_87 N_B_M1004_g N_VGND_c_219_n 0.00232702f $X=0.9 $Y=0.445 $X2=0 $Y2=0
cc_88 N_B_M1004_g N_VGND_c_220_n 0.00585385f $X=0.9 $Y=0.445 $X2=0 $Y2=0
cc_89 N_B_M1004_g N_VGND_c_221_n 0.00788151f $X=0.9 $Y=0.445 $X2=0 $Y2=0
cc_90 B N_VGND_c_221_n 0.0105931f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_91 N_A_M1002_g N_VPWR_c_155_n 0.00334685f $X=1.36 $Y=2.52 $X2=0 $Y2=0
cc_92 N_A_M1002_g N_VPWR_c_158_n 0.00428744f $X=1.36 $Y=2.52 $X2=0 $Y2=0
cc_93 N_A_M1002_g N_VPWR_c_152_n 0.00476395f $X=1.36 $Y=2.52 $X2=0 $Y2=0
cc_94 N_A_M1005_g N_Y_c_179_n 0.00458248f $X=1.29 $Y=0.445 $X2=0 $Y2=0
cc_95 A N_Y_c_179_n 0.00570189f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_96 N_A_c_123_n N_Y_c_179_n 0.00371573f $X=1.38 $Y=1.005 $X2=0 $Y2=0
cc_97 N_A_M1005_g Y 0.00621641f $X=1.29 $Y=0.445 $X2=0 $Y2=0
cc_98 N_A_M1002_g Y 0.00810018f $X=1.36 $Y=2.52 $X2=0 $Y2=0
cc_99 N_A_c_121_n Y 0.00270727f $X=1.38 $Y=1.51 $X2=0 $Y2=0
cc_100 A Y 0.0667312f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_101 N_A_c_123_n Y 0.0163648f $X=1.38 $Y=1.005 $X2=0 $Y2=0
cc_102 N_A_M1002_g N_Y_c_183_n 0.0167659f $X=1.36 $Y=2.52 $X2=0 $Y2=0
cc_103 N_A_c_121_n N_Y_c_183_n 5.71022e-19 $X=1.38 $Y=1.51 $X2=0 $Y2=0
cc_104 A N_Y_c_183_n 0.0249351f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_105 N_A_M1002_g N_Y_c_185_n 0.00646963f $X=1.36 $Y=2.52 $X2=0 $Y2=0
cc_106 N_A_M1005_g N_VGND_c_220_n 0.00552362f $X=1.29 $Y=0.445 $X2=0 $Y2=0
cc_107 N_A_M1005_g N_VGND_c_221_n 0.00741684f $X=1.29 $Y=0.445 $X2=0 $Y2=0
cc_108 A N_VGND_c_221_n 0.00810987f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_109 N_VPWR_c_155_n N_Y_c_183_n 0.0168699f $X=1.145 $Y=2.535 $X2=0 $Y2=0
cc_110 N_VPWR_c_154_n N_Y_c_184_n 0.00116713f $X=0.285 $Y=2.535 $X2=0 $Y2=0
cc_111 N_VPWR_c_155_n N_Y_c_184_n 0.00116713f $X=1.145 $Y=2.535 $X2=0 $Y2=0
cc_112 N_VPWR_c_156_n N_Y_c_184_n 0.00463811f $X=1.04 $Y=3.33 $X2=0 $Y2=0
cc_113 N_VPWR_c_152_n N_Y_c_184_n 0.00652376f $X=1.68 $Y=3.33 $X2=0 $Y2=0
cc_114 N_VPWR_c_155_n N_Y_c_185_n 0.00121271f $X=1.145 $Y=2.535 $X2=0 $Y2=0
cc_115 N_VPWR_c_158_n N_Y_c_185_n 0.00764843f $X=1.68 $Y=3.33 $X2=0 $Y2=0
cc_116 N_VPWR_c_152_n N_Y_c_185_n 0.0107579f $X=1.68 $Y=3.33 $X2=0 $Y2=0
cc_117 N_Y_c_179_n N_VGND_c_220_n 0.0153283f $X=1.645 $Y=0.51 $X2=0 $Y2=0
cc_118 N_Y_M1005_d N_VGND_c_221_n 0.00236056f $X=1.365 $Y=0.235 $X2=0 $Y2=0
cc_119 N_Y_c_179_n N_VGND_c_221_n 0.0163711f $X=1.645 $Y=0.51 $X2=0 $Y2=0
cc_120 N_VGND_c_221_n A_117_47# 0.00495496f $X=1.68 $Y=0 $X2=-0.19 $Y2=-0.245
cc_121 N_VGND_c_221_n A_195_47# 0.00749022f $X=1.68 $Y=0 $X2=-0.19 $Y2=-0.245
