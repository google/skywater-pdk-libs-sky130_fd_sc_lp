* File: sky130_fd_sc_lp__a2bb2oi_m.pex.spice
* Created: Fri Aug 28 09:57:08 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A2BB2OI_M%A1_N 2 3 4 5 6 9 11 13 16 17 18 19 20 21
+ 22 30
c46 11 0 1.07239e-19 $X=0.935 $Y=0.765
r47 21 22 20.5182 $w=1.98e-07 $l=3.7e-07 $layer=LI1_cond $X=0.255 $Y=2.035
+ $X2=0.255 $Y2=2.405
r48 20 21 20.5182 $w=1.98e-07 $l=3.7e-07 $layer=LI1_cond $X=0.255 $Y=1.665
+ $X2=0.255 $Y2=2.035
r49 19 20 20.5182 $w=1.98e-07 $l=3.7e-07 $layer=LI1_cond $X=0.255 $Y=1.295
+ $X2=0.255 $Y2=1.665
r50 18 19 20.5182 $w=1.98e-07 $l=3.7e-07 $layer=LI1_cond $X=0.255 $Y=0.925
+ $X2=0.255 $Y2=1.295
r51 18 30 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.27
+ $Y=0.93 $X2=0.27 $Y2=0.93
r52 17 18 20.5182 $w=1.98e-07 $l=3.7e-07 $layer=LI1_cond $X=0.255 $Y=0.555
+ $X2=0.255 $Y2=0.925
r53 15 30 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.27 $Y=1.27
+ $X2=0.27 $Y2=0.93
r54 15 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.27 $Y=1.27
+ $X2=0.27 $Y2=1.435
r55 14 30 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=0.27 $Y=0.915
+ $X2=0.27 $Y2=0.93
r56 11 13 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.935 $Y=0.765
+ $X2=0.935 $Y2=0.445
r57 7 9 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=0.585 $Y=2.215
+ $X2=0.585 $Y2=2.795
r58 6 14 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=0.435 $Y=0.84
+ $X2=0.27 $Y2=0.915
r59 5 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.86 $Y=0.84
+ $X2=0.935 $Y2=0.765
r60 5 6 217.926 $w=1.5e-07 $l=4.25e-07 $layer=POLY_cond $X=0.86 $Y=0.84
+ $X2=0.435 $Y2=0.84
r61 3 7 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.51 $Y=2.14
+ $X2=0.585 $Y2=2.215
r62 3 4 130.755 $w=1.5e-07 $l=2.55e-07 $layer=POLY_cond $X=0.51 $Y=2.14
+ $X2=0.255 $Y2=2.14
r63 2 4 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.18 $Y=2.065
+ $X2=0.255 $Y2=2.14
r64 2 16 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=0.18 $Y=2.065
+ $X2=0.18 $Y2=1.435
.ends

.subckt PM_SKY130_FD_SC_LP__A2BB2OI_M%A2_N 3 5 6 9 13 14 15 16 17 18 19 27
c51 9 0 1.04721e-19 $X=1.365 $Y=0.445
r52 27 28 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.81
+ $Y=1.32 $X2=0.81 $Y2=1.32
r53 18 19 16.4002 $w=2.58e-07 $l=3.7e-07 $layer=LI1_cond $X=0.765 $Y=2.405
+ $X2=0.765 $Y2=2.775
r54 17 18 16.4002 $w=2.58e-07 $l=3.7e-07 $layer=LI1_cond $X=0.765 $Y=2.035
+ $X2=0.765 $Y2=2.405
r55 16 17 16.4002 $w=2.58e-07 $l=3.7e-07 $layer=LI1_cond $X=0.765 $Y=1.665
+ $X2=0.765 $Y2=2.035
r56 16 28 15.292 $w=2.58e-07 $l=3.45e-07 $layer=LI1_cond $X=0.765 $Y=1.665
+ $X2=0.765 $Y2=1.32
r57 15 28 1.10812 $w=2.58e-07 $l=2.5e-08 $layer=LI1_cond $X=0.765 $Y=1.295
+ $X2=0.765 $Y2=1.32
r58 14 15 16.4002 $w=2.58e-07 $l=3.7e-07 $layer=LI1_cond $X=0.765 $Y=0.925
+ $X2=0.765 $Y2=1.295
r59 12 27 47.1618 $w=3.75e-07 $l=3.18e-07 $layer=POLY_cond $X=0.832 $Y=1.638
+ $X2=0.832 $Y2=1.32
r60 12 13 48.4185 $w=3.75e-07 $l=1.87e-07 $layer=POLY_cond $X=0.832 $Y=1.638
+ $X2=0.832 $Y2=1.825
r61 11 27 2.22462 $w=3.75e-07 $l=1.5e-08 $layer=POLY_cond $X=0.832 $Y=1.305
+ $X2=0.832 $Y2=1.32
r62 7 9 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=1.365 $Y=1.155
+ $X2=1.365 $Y2=0.445
r63 6 11 33.9315 $w=1.5e-07 $l=2.2236e-07 $layer=POLY_cond $X=1.02 $Y=1.23
+ $X2=0.832 $Y2=1.305
r64 5 7 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.29 $Y=1.23
+ $X2=1.365 $Y2=1.155
r65 5 6 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=1.29 $Y=1.23 $X2=1.02
+ $Y2=1.23
r66 3 13 497.383 $w=1.5e-07 $l=9.7e-07 $layer=POLY_cond $X=0.945 $Y=2.795
+ $X2=0.945 $Y2=1.825
.ends

.subckt PM_SKY130_FD_SC_LP__A2BB2OI_M%A_202_47# 1 2 8 9 10 11 12 15 17 19 21 23
+ 25 33 34
c65 25 0 1.07239e-19 $X=1.15 $Y=0.495
c66 17 0 7.39264e-20 $X=1.94 $Y=1.825
r67 34 36 27.9778 $w=3.3e-07 $l=1.6e-07 $layer=POLY_cond $X=1.61 $Y=2.86
+ $X2=1.45 $Y2=2.86
r68 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.61
+ $Y=2.86 $X2=1.61 $Y2=2.86
r69 31 33 15.3659 $w=3.28e-07 $l=4.4e-07 $layer=LI1_cond $X=1.17 $Y=2.86
+ $X2=1.61 $Y2=2.86
r70 29 31 0.349225 $w=3.28e-07 $l=1e-08 $layer=LI1_cond $X=1.16 $Y=2.86 $X2=1.17
+ $Y2=2.86
r71 25 27 8.88925 $w=2.18e-07 $l=1.65e-07 $layer=LI1_cond $X=1.155 $Y=0.495
+ $X2=1.155 $Y2=0.66
r72 23 31 3.96751 $w=1.9e-07 $l=1.65e-07 $layer=LI1_cond $X=1.17 $Y=2.695
+ $X2=1.17 $Y2=2.86
r73 23 27 118.789 $w=1.88e-07 $l=2.035e-06 $layer=LI1_cond $X=1.17 $Y=2.695
+ $X2=1.17 $Y2=0.66
r74 17 21 18.8402 $w=1.65e-07 $l=1.04283e-07 $layer=POLY_cond $X=1.94 $Y=1.825
+ $X2=1.87 $Y2=1.75
r75 17 19 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.94 $Y=1.825
+ $X2=1.94 $Y2=2.145
r76 15 20 507.638 $w=1.5e-07 $l=9.9e-07 $layer=POLY_cond $X=1.83 $Y=0.445
+ $X2=1.83 $Y2=1.435
r77 12 21 18.8402 $w=1.65e-07 $l=9.87421e-08 $layer=POLY_cond $X=1.815 $Y=1.675
+ $X2=1.87 $Y2=1.75
r78 11 20 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=1.815 $Y=1.525
+ $X2=1.815 $Y2=1.435
r79 11 12 58.3064 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=1.815 $Y=1.525
+ $X2=1.815 $Y2=1.675
r80 9 21 6.66866 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=1.725 $Y=1.75
+ $X2=1.87 $Y2=1.75
r81 9 10 102.553 $w=1.5e-07 $l=2e-07 $layer=POLY_cond $X=1.725 $Y=1.75 $X2=1.525
+ $Y2=1.75
r82 8 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.45 $Y=2.695
+ $X2=1.45 $Y2=2.86
r83 7 10 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.45 $Y=1.825
+ $X2=1.525 $Y2=1.75
r84 7 8 446.106 $w=1.5e-07 $l=8.7e-07 $layer=POLY_cond $X=1.45 $Y=1.825 $X2=1.45
+ $Y2=2.695
r85 2 29 600 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=1 $X=1.02
+ $Y=2.585 $X2=1.16 $Y2=2.86
r86 1 25 182 $w=1.7e-07 $l=3.2249e-07 $layer=licon1_NDIFF $count=1 $X=1.01
+ $Y=0.235 $X2=1.15 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__A2BB2OI_M%B2 3 6 9 10 11 12 13 17
c44 11 0 1.97996e-19 $X=2.28 $Y=1.435
r45 17 18 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.28
+ $Y=0.93 $X2=2.28 $Y2=0.93
r46 13 18 8.23714 $w=5.28e-07 $l=3.65e-07 $layer=LI1_cond $X=2.46 $Y=1.295
+ $X2=2.46 $Y2=0.93
r47 12 18 0.112838 $w=5.28e-07 $l=5e-09 $layer=LI1_cond $X=2.46 $Y=0.925
+ $X2=2.46 $Y2=0.93
r48 10 17 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.28 $Y=1.27
+ $X2=2.28 $Y2=0.93
r49 10 11 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.28 $Y=1.27
+ $X2=2.28 $Y2=1.435
r50 9 17 38.6168 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.28 $Y=0.765
+ $X2=2.28 $Y2=0.93
r51 6 11 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=2.37 $Y=2.145
+ $X2=2.37 $Y2=1.435
r52 3 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.26 $Y=0.445 $X2=2.26
+ $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_LP__A2BB2OI_M%B1 3 6 9 10 13 14 15 19
c31 10 0 1.50666e-19 $X=2.905 $Y=0.915
r32 19 20 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.99
+ $Y=0.93 $X2=2.99 $Y2=0.93
r33 15 20 14.0214 $w=2.98e-07 $l=3.65e-07 $layer=LI1_cond $X=3.055 $Y=1.295
+ $X2=3.055 $Y2=0.93
r34 14 20 0.192074 $w=2.98e-07 $l=5e-09 $layer=LI1_cond $X=3.055 $Y=0.925
+ $X2=3.055 $Y2=0.93
r35 12 19 58.5286 $w=3.5e-07 $l=3.55e-07 $layer=POLY_cond $X=2.98 $Y=1.285
+ $X2=2.98 $Y2=0.93
r36 12 13 43.9584 $w=3.5e-07 $l=1.5e-07 $layer=POLY_cond $X=2.94 $Y=1.285
+ $X2=2.94 $Y2=1.435
r37 10 19 2.47304 $w=3.5e-07 $l=1.5e-08 $layer=POLY_cond $X=2.98 $Y=0.915
+ $X2=2.98 $Y2=0.93
r38 9 10 43.9584 $w=3.5e-07 $l=1.5e-07 $layer=POLY_cond $X=2.905 $Y=0.765
+ $X2=2.905 $Y2=0.915
r39 6 13 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=2.8 $Y=2.145 $X2=2.8
+ $Y2=1.435
r40 3 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.73 $Y=0.445 $X2=2.73
+ $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_LP__A2BB2OI_M%VPWR 1 2 7 9 13 15 17 27 28 34
r32 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r33 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r34 28 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.64 $Y2=3.33
r35 27 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r36 25 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.75 $Y=3.33
+ $X2=2.585 $Y2=3.33
r37 25 27 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=2.75 $Y=3.33 $X2=3.12
+ $Y2=3.33
r38 24 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r39 23 24 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r40 21 32 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r41 20 23 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=0.72 $Y=3.33
+ $X2=2.16 $Y2=3.33
r42 20 21 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r43 18 31 4.70928 $w=1.7e-07 $l=2.28e-07 $layer=LI1_cond $X=0.455 $Y=3.33
+ $X2=0.227 $Y2=3.33
r44 18 20 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.455 $Y=3.33
+ $X2=0.72 $Y2=3.33
r45 17 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.42 $Y=3.33
+ $X2=2.585 $Y2=3.33
r46 17 23 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=2.42 $Y=3.33
+ $X2=2.16 $Y2=3.33
r47 15 24 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r48 15 21 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.72 $Y2=3.33
r49 11 34 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.585 $Y=3.245
+ $X2=2.585 $Y2=3.33
r50 11 13 36.1448 $w=3.28e-07 $l=1.035e-06 $layer=LI1_cond $X=2.585 $Y=3.245
+ $X2=2.585 $Y2=2.21
r51 7 31 3.0569 $w=3.3e-07 $l=1.12161e-07 $layer=LI1_cond $X=0.29 $Y=3.245
+ $X2=0.227 $Y2=3.33
r52 7 9 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=0.29 $Y=3.245
+ $X2=0.29 $Y2=2.86
r53 2 13 600 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=1 $X=2.445
+ $Y=1.935 $X2=2.585 $Y2=2.21
r54 1 9 600 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_PDIFF $count=1 $X=0.165
+ $Y=2.585 $X2=0.29 $Y2=2.86
.ends

.subckt PM_SKY130_FD_SC_LP__A2BB2OI_M%Y 1 2 8 12 17 19
c39 17 0 1.04721e-19 $X=2.045 $Y=0.48
c40 12 0 1.97996e-19 $X=1.93 $Y=1.49
r41 14 17 6.07359 $w=2.08e-07 $l=1.15e-07 $layer=LI1_cond $X=1.93 $Y=0.48
+ $X2=2.045 $Y2=0.48
r42 10 19 22.5585 $w=2.33e-07 $l=4.6e-07 $layer=LI1_cond $X=1.712 $Y=1.575
+ $X2=1.712 $Y2=2.035
r43 10 12 14.2225 $w=1.68e-07 $l=2.18e-07 $layer=LI1_cond $X=1.712 $Y=1.49
+ $X2=1.93 $Y2=1.49
r44 8 12 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.93 $Y=1.405
+ $X2=1.93 $Y2=1.49
r45 7 14 1.9771 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.93 $Y=0.585 $X2=1.93
+ $Y2=0.48
r46 7 8 53.4973 $w=1.68e-07 $l=8.2e-07 $layer=LI1_cond $X=1.93 $Y=0.585 $X2=1.93
+ $Y2=1.405
r47 2 19 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=1.6
+ $Y=1.935 $X2=1.725 $Y2=2.08
r48 1 17 182 $w=1.7e-07 $l=3.07124e-07 $layer=licon1_NDIFF $count=1 $X=1.905
+ $Y=0.235 $X2=2.045 $Y2=0.48
.ends

.subckt PM_SKY130_FD_SC_LP__A2BB2OI_M%A_403_387# 1 2 9 11 12 15
c17 9 0 2.18254e-19 $X=2.155 $Y=2.08
r18 13 15 9.04785 $w=1.88e-07 $l=1.55e-07 $layer=LI1_cond $X=3.025 $Y=1.925
+ $X2=3.025 $Y2=2.08
r19 11 13 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=2.93 $Y=1.84
+ $X2=3.025 $Y2=1.925
r20 11 12 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.93 $Y=1.84 $X2=2.24
+ $Y2=1.84
r21 7 12 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=2.145 $Y=1.925
+ $X2=2.24 $Y2=1.84
r22 7 9 9.04785 $w=1.88e-07 $l=1.55e-07 $layer=LI1_cond $X=2.145 $Y=1.925
+ $X2=2.145 $Y2=2.08
r23 2 15 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.875
+ $Y=1.935 $X2=3.015 $Y2=2.08
r24 1 9 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.015
+ $Y=1.935 $X2=2.155 $Y2=2.08
.ends

.subckt PM_SKY130_FD_SC_LP__A2BB2OI_M%VGND 1 2 3 12 16 18 20 23 24 25 27 36 44
+ 48
c49 18 0 1.50666e-19 $X=2.945 $Y=0.085
r50 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r51 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r52 42 48 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r53 41 42 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r54 38 41 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r55 36 47 4.50438 $w=1.7e-07 $l=2.9e-07 $layer=LI1_cond $X=2.78 $Y=0 $X2=3.07
+ $Y2=0
r56 36 41 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=2.78 $Y=0 $X2=2.64
+ $Y2=0
r57 35 45 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r58 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r59 32 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.865 $Y=0 $X2=0.7
+ $Y2=0
r60 32 34 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=0.865 $Y=0 $X2=1.2
+ $Y2=0
r61 30 45 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r62 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r63 27 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.535 $Y=0 $X2=0.7
+ $Y2=0
r64 27 29 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.535 $Y=0 $X2=0.24
+ $Y2=0
r65 25 42 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r66 25 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r67 25 38 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r68 23 34 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=1.475 $Y=0 $X2=1.2
+ $Y2=0
r69 23 24 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.475 $Y=0 $X2=1.57
+ $Y2=0
r70 22 38 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=1.665 $Y=0 $X2=1.68
+ $Y2=0
r71 22 24 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.665 $Y=0 $X2=1.57
+ $Y2=0
r72 18 47 3.26179 $w=3.3e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.945 $Y=0.085
+ $X2=3.07 $Y2=0
r73 18 20 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.945 $Y=0.085
+ $X2=2.945 $Y2=0.38
r74 14 24 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.57 $Y=0.085
+ $X2=1.57 $Y2=0
r75 14 16 17.2201 $w=1.88e-07 $l=2.95e-07 $layer=LI1_cond $X=1.57 $Y=0.085
+ $X2=1.57 $Y2=0.38
r76 10 44 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.7 $Y=0.085 $X2=0.7
+ $Y2=0
r77 10 12 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.7 $Y=0.085
+ $X2=0.7 $Y2=0.38
r78 3 20 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=2.805
+ $Y=0.235 $X2=2.945 $Y2=0.38
r79 2 16 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=1.44
+ $Y=0.235 $X2=1.58 $Y2=0.38
r80 1 12 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.575
+ $Y=0.235 $X2=0.7 $Y2=0.38
.ends

