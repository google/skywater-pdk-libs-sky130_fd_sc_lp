* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__nor4bb_m A B C_N D_N VGND VNB VPB VPWR Y
X0 a_27_507# D_N VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 VGND C_N a_284_99# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 a_454_397# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X3 Y A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 VGND a_27_507# Y VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 Y a_284_99# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 Y a_27_507# a_310_397# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X7 a_310_397# a_284_99# a_382_397# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X8 a_27_507# D_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X9 a_382_397# B a_454_397# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X10 VPWR C_N a_284_99# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X11 VGND B Y VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
