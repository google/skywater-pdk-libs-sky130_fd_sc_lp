* File: sky130_fd_sc_lp__buf_4.pex.spice
* Created: Fri Aug 28 10:10:27 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__BUF_4%A_122_23# 1 2 9 13 17 21 25 29 33 37 39 48 50
+ 51 52 53 54 57 61 65 72
r104 69 70 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=1.115 $Y=1.51
+ $X2=1.545 $Y2=1.51
r105 61 63 41.222 $w=2.58e-07 $l=9.3e-07 $layer=LI1_cond $X=2.655 $Y=1.98
+ $X2=2.655 $Y2=2.91
r106 59 61 2.43786 $w=2.58e-07 $l=5.5e-08 $layer=LI1_cond $X=2.655 $Y=1.925
+ $X2=2.655 $Y2=1.98
r107 55 57 19.5029 $w=2.58e-07 $l=4.4e-07 $layer=LI1_cond $X=2.655 $Y=0.86
+ $X2=2.655 $Y2=0.42
r108 53 59 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=2.525 $Y=1.84
+ $X2=2.655 $Y2=1.925
r109 53 54 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.525 $Y=1.84
+ $X2=2.22 $Y2=1.84
r110 51 55 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=2.525 $Y=0.945
+ $X2=2.655 $Y2=0.86
r111 51 52 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.525 $Y=0.945
+ $X2=2.22 $Y2=0.945
r112 50 54 6.85817 $w=1.7e-07 $l=1.33918e-07 $layer=LI1_cond $X=2.122 $Y=1.755
+ $X2=2.22 $Y2=1.84
r113 49 65 5.05528 $w=1.95e-07 $l=9.5e-08 $layer=LI1_cond $X=2.122 $Y=1.605
+ $X2=2.122 $Y2=1.51
r114 49 50 8.53147 $w=1.93e-07 $l=1.5e-07 $layer=LI1_cond $X=2.122 $Y=1.605
+ $X2=2.122 $Y2=1.755
r115 48 65 5.05528 $w=1.95e-07 $l=9.5e-08 $layer=LI1_cond $X=2.122 $Y=1.415
+ $X2=2.122 $Y2=1.51
r116 47 52 6.85817 $w=1.7e-07 $l=1.33918e-07 $layer=LI1_cond $X=2.122 $Y=1.03
+ $X2=2.22 $Y2=0.945
r117 47 48 21.8974 $w=1.93e-07 $l=3.85e-07 $layer=LI1_cond $X=2.122 $Y=1.03
+ $X2=2.122 $Y2=1.415
r118 46 72 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=1.885 $Y=1.51
+ $X2=1.975 $Y2=1.51
r119 46 70 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.885 $Y=1.51
+ $X2=1.545 $Y2=1.51
r120 45 46 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.885
+ $Y=1.51 $X2=1.885 $Y2=1.51
r121 42 69 43.7153 $w=3.3e-07 $l=2.5e-07 $layer=POLY_cond $X=0.865 $Y=1.51
+ $X2=1.115 $Y2=1.51
r122 42 66 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=0.865 $Y=1.51
+ $X2=0.685 $Y2=1.51
r123 41 45 59.5407 $w=1.88e-07 $l=1.02e-06 $layer=LI1_cond $X=0.865 $Y=1.51
+ $X2=1.885 $Y2=1.51
r124 41 42 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.865
+ $Y=1.51 $X2=0.865 $Y2=1.51
r125 39 65 1.43626 $w=1.9e-07 $l=9.7e-08 $layer=LI1_cond $X=2.025 $Y=1.51
+ $X2=2.122 $Y2=1.51
r126 39 45 8.17225 $w=1.88e-07 $l=1.4e-07 $layer=LI1_cond $X=2.025 $Y=1.51
+ $X2=1.885 $Y2=1.51
r127 35 72 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.975 $Y=1.675
+ $X2=1.975 $Y2=1.51
r128 35 37 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.975 $Y=1.675
+ $X2=1.975 $Y2=2.465
r129 31 72 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.975 $Y=1.345
+ $X2=1.975 $Y2=1.51
r130 31 33 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=1.975 $Y=1.345
+ $X2=1.975 $Y2=0.665
r131 27 70 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.545 $Y=1.675
+ $X2=1.545 $Y2=1.51
r132 27 29 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.545 $Y=1.675
+ $X2=1.545 $Y2=2.465
r133 23 70 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.545 $Y=1.345
+ $X2=1.545 $Y2=1.51
r134 23 25 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=1.545 $Y=1.345
+ $X2=1.545 $Y2=0.665
r135 19 69 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.115 $Y=1.675
+ $X2=1.115 $Y2=1.51
r136 19 21 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.115 $Y=1.675
+ $X2=1.115 $Y2=2.465
r137 15 69 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.115 $Y=1.345
+ $X2=1.115 $Y2=1.51
r138 15 17 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=1.115 $Y=1.345
+ $X2=1.115 $Y2=0.665
r139 11 66 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.685 $Y=1.675
+ $X2=0.685 $Y2=1.51
r140 11 13 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=0.685 $Y=1.675
+ $X2=0.685 $Y2=2.465
r141 7 66 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.685 $Y=1.345
+ $X2=0.685 $Y2=1.51
r142 7 9 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=0.685 $Y=1.345
+ $X2=0.685 $Y2=0.665
r143 2 63 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=2.48
+ $Y=1.835 $X2=2.62 $Y2=2.91
r144 2 61 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.48
+ $Y=1.835 $X2=2.62 $Y2=1.98
r145 1 57 91 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=2 $X=2.48
+ $Y=0.245 $X2=2.62 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__BUF_4%A 3 6 8 11 13
r26 11 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.495 $Y=1.375
+ $X2=2.495 $Y2=1.54
r27 11 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.495 $Y=1.375
+ $X2=2.495 $Y2=1.21
r28 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.495
+ $Y=1.375 $X2=2.495 $Y2=1.375
r29 8 12 4.91483 $w=3.38e-07 $l=1.45e-07 $layer=LI1_cond $X=2.64 $Y=1.37
+ $X2=2.495 $Y2=1.37
r30 6 14 474.309 $w=1.5e-07 $l=9.25e-07 $layer=POLY_cond $X=2.405 $Y=2.465
+ $X2=2.405 $Y2=1.54
r31 3 13 175.127 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=2.405 $Y=0.665
+ $X2=2.405 $Y2=1.21
.ends

.subckt PM_SKY130_FD_SC_LP__BUF_4%VPWR 1 2 3 12 16 20 26 30 31 32 37 44 45 48 51
r50 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r51 48 49 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r52 45 52 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r53 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r54 42 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.355 $Y=3.33
+ $X2=2.19 $Y2=3.33
r55 42 44 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=2.355 $Y=3.33
+ $X2=2.64 $Y2=3.33
r56 41 52 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r57 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r58 38 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.495 $Y=3.33
+ $X2=1.33 $Y2=3.33
r59 38 40 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=1.495 $Y=3.33
+ $X2=1.68 $Y2=3.33
r60 37 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.025 $Y=3.33
+ $X2=2.19 $Y2=3.33
r61 37 40 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=2.025 $Y=3.33
+ $X2=1.68 $Y2=3.33
r62 36 49 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.2 $Y2=3.33
r63 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r64 32 41 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=1.68 $Y2=3.33
r65 32 49 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=1.2 $Y2=3.33
r66 30 35 4.66471 $w=1.7e-07 $l=6.5e-08 $layer=LI1_cond $X=0.305 $Y=3.33
+ $X2=0.24 $Y2=3.33
r67 30 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.305 $Y=3.33
+ $X2=0.47 $Y2=3.33
r68 26 29 26.8903 $w=3.28e-07 $l=7.7e-07 $layer=LI1_cond $X=2.19 $Y=2.18
+ $X2=2.19 $Y2=2.95
r69 24 51 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.19 $Y=3.245
+ $X2=2.19 $Y2=3.33
r70 24 29 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.19 $Y=3.245
+ $X2=2.19 $Y2=2.95
r71 20 23 26.8903 $w=3.28e-07 $l=7.7e-07 $layer=LI1_cond $X=1.33 $Y=2.2 $X2=1.33
+ $Y2=2.97
r72 18 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.33 $Y=3.245
+ $X2=1.33 $Y2=3.33
r73 18 23 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=1.33 $Y=3.245
+ $X2=1.33 $Y2=2.97
r74 17 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.635 $Y=3.33
+ $X2=0.47 $Y2=3.33
r75 16 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.165 $Y=3.33
+ $X2=1.33 $Y2=3.33
r76 16 17 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=1.165 $Y=3.33
+ $X2=0.635 $Y2=3.33
r77 12 15 26.8903 $w=3.28e-07 $l=7.7e-07 $layer=LI1_cond $X=0.47 $Y=2.2 $X2=0.47
+ $Y2=2.97
r78 10 31 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.47 $Y=3.245
+ $X2=0.47 $Y2=3.33
r79 10 15 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=0.47 $Y=3.245
+ $X2=0.47 $Y2=2.97
r80 3 29 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=2.05
+ $Y=1.835 $X2=2.19 $Y2=2.95
r81 3 26 400 $w=1.7e-07 $l=4.09054e-07 $layer=licon1_PDIFF $count=1 $X=2.05
+ $Y=1.835 $X2=2.19 $Y2=2.18
r82 2 23 400 $w=1.7e-07 $l=1.20297e-06 $layer=licon1_PDIFF $count=1 $X=1.19
+ $Y=1.835 $X2=1.33 $Y2=2.97
r83 2 20 400 $w=1.7e-07 $l=4.29331e-07 $layer=licon1_PDIFF $count=1 $X=1.19
+ $Y=1.835 $X2=1.33 $Y2=2.2
r84 1 15 400 $w=1.7e-07 $l=1.20532e-06 $layer=licon1_PDIFF $count=1 $X=0.325
+ $Y=1.835 $X2=0.47 $Y2=2.97
r85 1 12 400 $w=1.7e-07 $l=4.31451e-07 $layer=licon1_PDIFF $count=1 $X=0.325
+ $Y=1.835 $X2=0.47 $Y2=2.2
.ends

.subckt PM_SKY130_FD_SC_LP__BUF_4%X 1 2 3 4 13 15 16 19 23 27 29 33 37 42 43 44
+ 45 49 51
r56 49 51 1.38849 $w=4.13e-07 $l=5e-08 $layer=LI1_cond $X=0.302 $Y=1.245
+ $X2=0.302 $Y2=1.295
r57 44 49 2.46632 $w=4.15e-07 $l=8.5e-08 $layer=LI1_cond $X=0.302 $Y=1.16
+ $X2=0.302 $Y2=1.245
r58 44 45 9.80271 $w=4.13e-07 $l=3.53e-07 $layer=LI1_cond $X=0.302 $Y=1.312
+ $X2=0.302 $Y2=1.665
r59 44 51 0.472085 $w=4.13e-07 $l=1.7e-08 $layer=LI1_cond $X=0.302 $Y=1.312
+ $X2=0.302 $Y2=1.295
r60 41 45 3.05467 $w=4.13e-07 $l=1.1e-07 $layer=LI1_cond $X=0.302 $Y=1.775
+ $X2=0.302 $Y2=1.665
r61 37 39 54.2871 $w=1.88e-07 $l=9.3e-07 $layer=LI1_cond $X=1.76 $Y=1.98
+ $X2=1.76 $Y2=2.91
r62 35 37 2.04306 $w=1.88e-07 $l=3.5e-08 $layer=LI1_cond $X=1.76 $Y=1.945
+ $X2=1.76 $Y2=1.98
r63 31 33 38.2345 $w=1.88e-07 $l=6.55e-07 $layer=LI1_cond $X=1.76 $Y=1.075
+ $X2=1.76 $Y2=0.42
r64 30 43 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=0.995 $Y=1.86 $X2=0.9
+ $Y2=1.86
r65 29 35 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=1.665 $Y=1.86
+ $X2=1.76 $Y2=1.945
r66 29 30 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.665 $Y=1.86
+ $X2=0.995 $Y2=1.86
r67 28 42 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=0.995 $Y=1.16 $X2=0.9
+ $Y2=1.16
r68 27 31 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=1.665 $Y=1.16
+ $X2=1.76 $Y2=1.075
r69 27 28 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.665 $Y=1.16
+ $X2=0.995 $Y2=1.16
r70 23 25 54.2871 $w=1.88e-07 $l=9.3e-07 $layer=LI1_cond $X=0.9 $Y=1.98 $X2=0.9
+ $Y2=2.91
r71 21 43 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=0.9 $Y=1.945 $X2=0.9
+ $Y2=1.86
r72 21 23 2.04306 $w=1.88e-07 $l=3.5e-08 $layer=LI1_cond $X=0.9 $Y=1.945 $X2=0.9
+ $Y2=1.98
r73 17 42 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=0.9 $Y=1.075 $X2=0.9
+ $Y2=1.16
r74 17 19 38.2345 $w=1.88e-07 $l=6.55e-07 $layer=LI1_cond $X=0.9 $Y=1.075
+ $X2=0.9 $Y2=0.42
r75 16 41 8.50155 $w=1.7e-07 $l=2.46868e-07 $layer=LI1_cond $X=0.51 $Y=1.86
+ $X2=0.302 $Y2=1.775
r76 15 43 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=0.805 $Y=1.86 $X2=0.9
+ $Y2=1.86
r77 15 16 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.805 $Y=1.86
+ $X2=0.51 $Y2=1.86
r78 14 44 6.03523 $w=1.7e-07 $l=2.08e-07 $layer=LI1_cond $X=0.51 $Y=1.16
+ $X2=0.302 $Y2=1.16
r79 13 42 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=0.805 $Y=1.16 $X2=0.9
+ $Y2=1.16
r80 13 14 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.805 $Y=1.16
+ $X2=0.51 $Y2=1.16
r81 4 39 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=1.62
+ $Y=1.835 $X2=1.76 $Y2=2.91
r82 4 37 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.62
+ $Y=1.835 $X2=1.76 $Y2=1.98
r83 3 25 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=0.76
+ $Y=1.835 $X2=0.9 $Y2=2.91
r84 3 23 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.76
+ $Y=1.835 $X2=0.9 $Y2=1.98
r85 2 33 91 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=2 $X=1.62
+ $Y=0.245 $X2=1.76 $Y2=0.42
r86 1 19 91 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=2 $X=0.76
+ $Y=0.245 $X2=0.9 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__BUF_4%VGND 1 2 3 12 14 18 22 24 25 26 31 38 39 42 45
r52 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r53 42 43 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r54 39 46 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=2.16
+ $Y2=0
r55 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r56 36 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.355 $Y=0 $X2=2.19
+ $Y2=0
r57 36 38 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=2.355 $Y=0 $X2=2.64
+ $Y2=0
r58 35 46 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r59 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r60 32 42 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.495 $Y=0 $X2=1.33
+ $Y2=0
r61 32 34 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=1.495 $Y=0 $X2=1.68
+ $Y2=0
r62 31 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.025 $Y=0 $X2=2.19
+ $Y2=0
r63 31 34 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=2.025 $Y=0 $X2=1.68
+ $Y2=0
r64 30 43 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r65 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r66 26 35 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=1.68
+ $Y2=0
r67 26 43 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=1.2
+ $Y2=0
r68 24 29 4.66471 $w=1.7e-07 $l=6.5e-08 $layer=LI1_cond $X=0.305 $Y=0 $X2=0.24
+ $Y2=0
r69 24 25 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.305 $Y=0 $X2=0.47
+ $Y2=0
r70 20 45 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.19 $Y=0.085
+ $X2=2.19 $Y2=0
r71 20 22 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=2.19 $Y=0.085
+ $X2=2.19 $Y2=0.565
r72 16 42 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.33 $Y=0.085
+ $X2=1.33 $Y2=0
r73 16 18 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=1.33 $Y=0.085
+ $X2=1.33 $Y2=0.39
r74 15 25 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.635 $Y=0 $X2=0.47
+ $Y2=0
r75 14 42 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.165 $Y=0 $X2=1.33
+ $Y2=0
r76 14 15 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=1.165 $Y=0 $X2=0.635
+ $Y2=0
r77 10 25 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.47 $Y=0.085
+ $X2=0.47 $Y2=0
r78 10 12 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=0.47 $Y=0.085
+ $X2=0.47 $Y2=0.39
r79 3 22 182 $w=1.7e-07 $l=3.83667e-07 $layer=licon1_NDIFF $count=1 $X=2.05
+ $Y=0.245 $X2=2.19 $Y2=0.565
r80 2 18 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.19
+ $Y=0.245 $X2=1.33 $Y2=0.39
r81 1 12 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.345
+ $Y=0.245 $X2=0.47 $Y2=0.39
.ends

