* File: sky130_fd_sc_lp__clkdlybuf4s25_1.spice
* Created: Fri Aug 28 10:16:50 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__clkdlybuf4s25_1.pex.spice"
.subckt sky130_fd_sc_lp__clkdlybuf4s25_1  VNB VPB A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* VPB	VPB
* VNB	VNB
MM1003 N_VGND_M1003_d N_A_M1003_g N_A_27_52#_M1003_s VNB NSHORT L=0.15 W=0.42
+ AD=0.161552 AS=0.1113 PD=0.952394 PS=1.37 NRD=15.708 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1004 N_A_282_52#_M1004_d N_A_27_52#_M1004_g N_VGND_M1003_d VNB NSHORT L=0.25
+ W=1 AD=0.265 AS=0.384648 PD=2.53 PS=2.26761 NRD=0 NRS=32.988 M=1 R=4 SA=125001
+ SB=125000 A=0.25 P=2.5 MULT=1
MM1006 N_VGND_M1006_d N_A_282_52#_M1006_g N_A_394_52#_M1006_s VNB NSHORT L=0.25
+ W=1 AD=0.384648 AS=0.265 PD=2.26761 PS=2.53 NRD=29.988 NRS=0 M=1 R=4 SA=125000
+ SB=125001 A=0.25 P=2.5 MULT=1
MM1005 N_X_M1005_d N_A_394_52#_M1005_g N_VGND_M1006_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.161552 PD=1.37 PS=0.952394 NRD=0 NRS=22.848 M=1 R=2.8
+ SA=75001.1 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1007 N_VPWR_M1007_d N_A_M1007_g N_A_27_52#_M1007_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.376327 AS=0.3339 PD=2.08513 PS=3.05 NRD=10.9335 NRS=0 M=1 R=8.4
+ SA=75000.2 SB=75000.9 A=0.189 P=2.82 MULT=1
MM1002 N_A_282_52#_M1002_d N_A_27_52#_M1002_g N_VPWR_M1007_d VPB PHIGHVT L=0.25
+ W=1 AD=0.265 AS=0.298673 PD=2.53 PS=1.65487 NRD=0 NRS=51.2003 M=1 R=4
+ SA=125001 SB=125000 A=0.25 P=2.5 MULT=1
MM1001 N_VPWR_M1001_d N_A_282_52#_M1001_g N_A_394_52#_M1001_s VPB PHIGHVT L=0.25
+ W=1 AD=0.298673 AS=0.265 PD=1.65487 PS=2.53 NRD=49.2303 NRS=0 M=1 R=4
+ SA=125000 SB=125001 A=0.25 P=2.5 MULT=1
MM1000 N_X_M1000_d N_A_394_52#_M1000_g N_VPWR_M1001_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.376327 PD=3.05 PS=2.08513 NRD=0 NRS=12.4898 M=1 R=8.4
+ SA=75000.9 SB=75000.2 A=0.189 P=2.82 MULT=1
DX8_noxref VNB VPB NWDIODE A=7.8703 P=12.17
*
.include "sky130_fd_sc_lp__clkdlybuf4s25_1.pxi.spice"
*
.ends
*
*
