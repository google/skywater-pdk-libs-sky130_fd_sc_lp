* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__ha_4 A B VGND VNB VPB VPWR COUT SUM
X0 VPWR a_454_263# COUT VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X1 a_851_47# B a_454_263# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X2 VPWR a_110_263# SUM VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X3 VPWR B a_454_263# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X4 VGND A a_1284_65# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X5 a_1284_65# A VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X6 VGND a_110_263# SUM VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X7 a_1284_65# B VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X8 COUT a_454_263# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X9 VPWR a_454_263# COUT VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X10 SUM a_110_263# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X11 VGND a_454_263# COUT VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X12 a_110_263# B a_1367_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X13 VPWR a_454_263# a_110_263# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X14 a_454_263# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X15 VGND B a_1284_65# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X16 VPWR A a_454_263# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X17 VGND a_110_263# SUM VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X18 a_1284_65# a_454_263# a_110_263# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X19 SUM a_110_263# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X20 SUM a_110_263# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X21 COUT a_454_263# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X22 a_454_263# B a_851_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X23 a_454_263# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X24 COUT a_454_263# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X25 VGND a_454_263# COUT VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X26 a_1367_367# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X27 a_110_263# a_454_263# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X28 VGND A a_851_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X29 a_110_263# a_454_263# a_1284_65# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X30 SUM a_110_263# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X31 a_851_47# A VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X32 VPWR a_110_263# SUM VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X33 COUT a_454_263# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X34 a_1367_367# B a_110_263# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X35 VPWR A a_1367_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
.ends
