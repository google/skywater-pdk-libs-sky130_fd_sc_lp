* File: sky130_fd_sc_lp__o21bai_m.spice
* Created: Wed Sep  2 10:17:58 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__o21bai_m.pex.spice"
.subckt sky130_fd_sc_lp__o21bai_m  VNB VPB B1_N A2 A1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A1	A1
* A2	A2
* B1_N	B1_N
* VPB	VPB
* VNB	VNB
MM1002 N_VGND_M1002_d N_B1_N_M1002_g N_A_32_62#_M1002_s VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.1113 PD=1.37 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1001 N_A_320_78#_M1001_d N_A_32_62#_M1001_g N_Y_M1001_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1006 N_VGND_M1006_d N_A2_M1006_g N_A_320_78#_M1001_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1000 N_A_320_78#_M1000_d N_A1_M1000_g N_VGND_M1006_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.1 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1005 N_VPWR_M1005_d N_B1_N_M1005_g N_A_32_62#_M1005_s VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0819 AS=0.1113 PD=0.81 PS=1.37 NRD=37.5088 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.5 A=0.063 P=1.14 MULT=1
MM1007 N_Y_M1007_d N_A_32_62#_M1007_g N_VPWR_M1005_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0588 AS=0.0819 PD=0.7 PS=0.81 NRD=0 NRS=14.0658 M=1 R=2.8 SA=75000.7
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1003 A_315_535# N_A2_M1003_g N_Y_M1007_d VPB PHIGHVT L=0.15 W=0.42 AD=0.0441
+ AS=0.0588 PD=0.63 PS=0.7 NRD=23.443 NRS=0 M=1 R=2.8 SA=75001.2 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1004 N_VPWR_M1004_d N_A1_M1004_g A_315_535# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=23.443 M=1 R=2.8 SA=75001.5
+ SB=75000.2 A=0.063 P=1.14 MULT=1
DX8_noxref VNB VPB NWDIODE A=6.0799 P=10.25
*
.include "sky130_fd_sc_lp__o21bai_m.pxi.spice"
*
.ends
*
*
