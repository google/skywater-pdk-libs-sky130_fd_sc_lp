* File: sky130_fd_sc_lp__o31ai_2.spice
* Created: Wed Sep  2 10:25:21 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__o31ai_2.pex.spice"
.subckt sky130_fd_sc_lp__o31ai_2  VNB VPB A1 A2 A3 B1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B1	B1
* A3	A3
* A2	A2
* A1	A1
* VPB	VPB
* VNB	VNB
MM1000 N_A_58_65#_M1000_d N_A1_M1000_g N_VGND_M1000_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75003.7 A=0.126 P=1.98 MULT=1
MM1010 N_A_58_65#_M1010_d N_A1_M1010_g N_VGND_M1000_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75003.3 A=0.126 P=1.98 MULT=1
MM1003 N_VGND_M1003_d N_A2_M1003_g N_A_58_65#_M1010_d VNB NSHORT L=0.15 W=0.84
+ AD=0.294 AS=0.1176 PD=1.54 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.1 SB=75002.8
+ A=0.126 P=1.98 MULT=1
MM1014 N_VGND_M1003_d N_A2_M1014_g N_A_58_65#_M1014_s VNB NSHORT L=0.15 W=0.84
+ AD=0.294 AS=0.1176 PD=1.54 PS=1.12 NRD=4.992 NRS=0 M=1 R=5.6 SA=75001.9
+ SB=75002 A=0.126 P=1.98 MULT=1
MM1008 N_VGND_M1008_d N_A3_M1008_g N_A_58_65#_M1014_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002.3
+ SB=75001.6 A=0.126 P=1.98 MULT=1
MM1013 N_VGND_M1008_d N_A3_M1013_g N_A_58_65#_M1013_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.147 PD=1.12 PS=1.19 NRD=0 NRS=0 M=1 R=5.6 SA=75002.8 SB=75001.1
+ A=0.126 P=1.98 MULT=1
MM1001 N_A_58_65#_M1013_s N_B1_M1001_g N_Y_M1001_s VNB NSHORT L=0.15 W=0.84
+ AD=0.147 AS=0.1176 PD=1.19 PS=1.12 NRD=9.996 NRS=0 M=1 R=5.6 SA=75003.3
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1011 N_A_58_65#_M1011_d N_B1_M1011_g N_Y_M1001_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75003.7
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1002 N_VPWR_M1002_d N_A1_M1002_g N_A_44_367#_M1002_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75001.5 A=0.189 P=2.82 MULT=1
MM1009 N_VPWR_M1002_d N_A1_M1009_g N_A_44_367#_M1009_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1004 N_A_299_367#_M1004_d N_A2_M1004_g N_A_44_367#_M1009_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1015 N_A_299_367#_M1004_d N_A2_M1015_g N_A_44_367#_M1015_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75001.5
+ SB=75000.2 A=0.189 P=2.82 MULT=1
MM1005 N_A_299_367#_M1005_d N_A3_M1005_g N_Y_M1005_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.2268 AS=0.3339 PD=1.62 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75001.7 A=0.189 P=2.82 MULT=1
MM1006 N_A_299_367#_M1005_d N_A3_M1006_g N_Y_M1006_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.2268 AS=0.27405 PD=1.62 PS=1.695 NRD=12.4898 NRS=8.5892 M=1 R=8.4
+ SA=75000.7 SB=75001.2 A=0.189 P=2.82 MULT=1
MM1007 N_Y_M1006_s N_B1_M1007_g N_VPWR_M1007_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.27405 AS=0.1764 PD=1.695 PS=1.54 NRD=15.6221 NRS=0 M=1 R=8.4 SA=75001.3
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1012 N_Y_M1012_d N_B1_M1012_g N_VPWR_M1007_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.7
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX16_noxref VNB VPB NWDIODE A=9.6607 P=14.09
*
.include "sky130_fd_sc_lp__o31ai_2.pxi.spice"
*
.ends
*
*
