* File: sky130_fd_sc_lp__o311ai_0.spice
* Created: Wed Sep  2 10:23:37 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__o311ai_0.pex.spice"
.subckt sky130_fd_sc_lp__o311ai_0  VNB VPB A1 A2 A3 B1 C1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* C1	C1
* B1	B1
* A3	A3
* A2	A2
* A1	A1
* VPB	VPB
* VNB	VNB
MM1005 N_A_193_48#_M1005_d N_A1_M1005_g N_VGND_M1005_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75001.9
+ A=0.063 P=1.14 MULT=1
MM1000 N_VGND_M1000_d N_A2_M1000_g N_A_193_48#_M1005_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0714 AS=0.0588 PD=0.76 PS=0.7 NRD=9.996 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75001.5 A=0.063 P=1.14 MULT=1
MM1006 N_A_193_48#_M1006_d N_A3_M1006_g N_VGND_M1000_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0714 PD=0.7 PS=0.76 NRD=0 NRS=7.14 M=1 R=2.8 SA=75001.1
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1009 A_463_48# N_B1_M1009_g N_A_193_48#_M1006_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.0588 PD=0.66 PS=0.7 NRD=18.564 NRS=0 M=1 R=2.8 SA=75001.5
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1008 N_Y_M1008_d N_C1_M1008_g A_463_48# VNB NSHORT L=0.15 W=0.42 AD=0.1113
+ AS=0.0504 PD=1.37 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75001.9 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1001 A_193_466# N_A1_M1001_g N_VPWR_M1001_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0672 AS=0.1696 PD=0.85 PS=1.81 NRD=15.3857 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75001.9 A=0.096 P=1.58 MULT=1
MM1002 A_265_466# N_A2_M1002_g A_193_466# VPB PHIGHVT L=0.15 W=0.64 AD=0.0672
+ AS=0.0672 PD=0.85 PS=0.85 NRD=15.3857 NRS=15.3857 M=1 R=4.26667 SA=75000.6
+ SB=75001.6 A=0.096 P=1.58 MULT=1
MM1004 N_Y_M1004_d N_A3_M1004_g A_265_466# VPB PHIGHVT L=0.15 W=0.64 AD=0.1088
+ AS=0.0672 PD=0.98 PS=0.85 NRD=13.8491 NRS=15.3857 M=1 R=4.26667 SA=75000.9
+ SB=75001.2 A=0.096 P=1.58 MULT=1
MM1007 N_VPWR_M1007_d N_B1_M1007_g N_Y_M1004_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1216 AS=0.1088 PD=1.02 PS=0.98 NRD=16.9223 NRS=4.6098 M=1 R=4.26667
+ SA=75001.4 SB=75000.7 A=0.096 P=1.58 MULT=1
MM1003 N_Y_M1003_d N_C1_M1003_g N_VPWR_M1007_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1696 AS=0.1216 PD=1.81 PS=1.02 NRD=0 NRS=13.8491 M=1 R=4.26667 SA=75001.9
+ SB=75000.2 A=0.096 P=1.58 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9751 P=11.21
*
.include "sky130_fd_sc_lp__o311ai_0.pxi.spice"
*
.ends
*
*
