* NGSPICE file created from sky130_fd_sc_lp__maj3_0.ext - technology: sky130A

.subckt sky130_fd_sc_lp__maj3_0 A B C VGND VNB VPB VPWR X
M1000 a_149_57# C a_28_431# VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=2.373e+11p ps=2.81e+06u
M1001 a_313_57# A VGND VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=2.352e+11p ps=2.8e+06u
M1002 a_28_431# B a_313_57# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 X a_28_431# VGND VNB nshort w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=0p ps=0u
M1004 a_477_431# B a_28_431# VPB phighvt w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=2.373e+11p ps=2.81e+06u
M1005 VPWR C a_477_431# VPB phighvt w=420000u l=150000u
+  ad=4.449e+11p pd=3.94e+06u as=0p ps=0u
M1006 a_28_431# B a_319_431# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1007 a_477_57# B a_28_431# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1008 a_319_431# A VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 X a_28_431# VPWR VPB phighvt w=640000u l=150000u
+  ad=2.56e+11p pd=2.08e+06u as=0p ps=0u
M1010 VGND A a_149_57# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND C a_477_57# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VPWR A a_115_431# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1013 a_115_431# C a_28_431# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

