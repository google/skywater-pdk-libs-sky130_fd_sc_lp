* NGSPICE file created from sky130_fd_sc_lp__sdlclkp_4.ext - technology: sky130A

.subckt sky130_fd_sc_lp__sdlclkp_4 CLK GATE SCE VGND VNB VPB VPWR GCLK
M1000 VPWR a_762_107# a_720_463# VPB phighvt w=420000u l=150000u
+  ad=2.5484e+12p pd=2.049e+07u as=8.82e+10p ps=1.26e+06u
M1001 GCLK a_1275_367# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=7.056e+11p pd=6.16e+06u as=0p ps=0u
M1002 a_1216_47# CLK VGND VNB nshort w=840000u l=150000u
+  ad=1.764e+11p pd=2.1e+06u as=1.6132e+12p ps=1.495e+07u
M1003 a_1275_367# a_762_107# a_1216_47# VNB nshort w=840000u l=150000u
+  ad=2.226e+11p pd=2.21e+06u as=0p ps=0u
M1004 a_762_107# a_634_133# VGND VNB nshort w=840000u l=150000u
+  ad=2.394e+11p pd=2.25e+06u as=0p ps=0u
M1005 a_762_107# a_634_133# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=3.339e+11p pd=3.05e+06u as=0p ps=0u
M1006 GCLK a_1275_367# VGND VNB nshort w=840000u l=150000u
+  ad=4.704e+11p pd=4.48e+06u as=0p ps=0u
M1007 VPWR a_762_107# a_1275_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=3.528e+11p ps=3.08e+06u
M1008 VPWR a_1275_367# GCLK VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND a_762_107# a_720_133# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1010 GCLK a_1275_367# VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_634_133# a_252_361# a_134_70# VNB nshort w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=2.436e+11p ps=2.84e+06u
M1012 VGND GATE a_134_70# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VPWR a_1275_367# GCLK VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_134_70# SCE VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_335_70# a_252_361# VPWR VPB phighvt w=640000u l=150000u
+  ad=2.112e+11p pd=1.94e+06u as=0p ps=0u
M1016 a_720_133# a_335_70# a_634_133# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VGND CLK a_252_361# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1018 a_1275_367# CLK VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_134_70# GATE a_110_468# VPB phighvt w=640000u l=150000u
+  ad=2.809e+11p pd=3.18e+06u as=1.344e+11p ps=1.7e+06u
M1020 a_634_133# a_335_70# a_134_70# VPB phighvt w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=0p ps=0u
M1021 VGND a_1275_367# GCLK VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_110_468# SCE VPWR VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 GCLK a_1275_367# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 VGND a_1275_367# GCLK VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_720_463# a_252_361# a_634_133# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 VPWR CLK a_252_361# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.696e+11p ps=1.81e+06u
M1027 a_335_70# a_252_361# VGND VNB nshort w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
.ends

