* File: sky130_fd_sc_lp__o2111ai_lp.pxi.spice
* Created: Wed Sep  2 10:13:22 2020
* 
x_PM_SKY130_FD_SC_LP__O2111AI_LP%D1 N_D1_M1008_g N_D1_M1002_g N_D1_c_67_n
+ N_D1_c_68_n D1 N_D1_c_69_n N_D1_c_70_n PM_SKY130_FD_SC_LP__O2111AI_LP%D1
x_PM_SKY130_FD_SC_LP__O2111AI_LP%C1 N_C1_M1003_g N_C1_c_103_n N_C1_M1004_g
+ N_C1_c_105_n C1 C1 C1 N_C1_c_107_n PM_SKY130_FD_SC_LP__O2111AI_LP%C1
x_PM_SKY130_FD_SC_LP__O2111AI_LP%B1 N_B1_M1007_g N_B1_M1006_g N_B1_c_152_n
+ N_B1_c_153_n B1 B1 N_B1_c_155_n PM_SKY130_FD_SC_LP__O2111AI_LP%B1
x_PM_SKY130_FD_SC_LP__O2111AI_LP%A2 N_A2_M1009_g N_A2_c_194_n N_A2_M1000_g
+ N_A2_c_195_n A2 A2 N_A2_c_196_n N_A2_c_197_n PM_SKY130_FD_SC_LP__O2111AI_LP%A2
x_PM_SKY130_FD_SC_LP__O2111AI_LP%A1 N_A1_M1001_g N_A1_M1005_g A1 A1 N_A1_c_237_n
+ PM_SKY130_FD_SC_LP__O2111AI_LP%A1
x_PM_SKY130_FD_SC_LP__O2111AI_LP%VPWR N_VPWR_M1008_s N_VPWR_M1004_d
+ N_VPWR_M1001_d N_VPWR_c_264_n N_VPWR_c_265_n N_VPWR_c_266_n N_VPWR_c_267_n
+ N_VPWR_c_268_n N_VPWR_c_269_n N_VPWR_c_270_n VPWR N_VPWR_c_271_n
+ N_VPWR_c_263_n PM_SKY130_FD_SC_LP__O2111AI_LP%VPWR
x_PM_SKY130_FD_SC_LP__O2111AI_LP%Y N_Y_M1002_s N_Y_M1008_d N_Y_M1006_d
+ N_Y_c_306_n N_Y_c_307_n N_Y_c_308_n N_Y_c_309_n N_Y_c_310_n N_Y_c_311_n Y Y Y
+ Y N_Y_c_305_n PM_SKY130_FD_SC_LP__O2111AI_LP%Y
x_PM_SKY130_FD_SC_LP__O2111AI_LP%A_347_57# N_A_347_57#_M1007_d
+ N_A_347_57#_M1005_d N_A_347_57#_c_363_n N_A_347_57#_c_364_n
+ N_A_347_57#_c_365_n N_A_347_57#_c_366_n
+ PM_SKY130_FD_SC_LP__O2111AI_LP%A_347_57#
x_PM_SKY130_FD_SC_LP__O2111AI_LP%VGND N_VGND_M1009_d N_VGND_c_390_n
+ N_VGND_c_391_n N_VGND_c_392_n VGND N_VGND_c_393_n N_VGND_c_394_n
+ PM_SKY130_FD_SC_LP__O2111AI_LP%VGND
cc_1 VNB N_D1_M1008_g 0.00553126f $X=-0.19 $Y=-0.245 $X2=0.68 $Y2=2.545
cc_2 VNB N_D1_M1002_g 0.0251878f $X=-0.19 $Y=-0.245 $X2=0.76 $Y2=0.495
cc_3 VNB N_D1_c_67_n 0.025617f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.41
cc_4 VNB N_D1_c_68_n 0.0147354f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.575
cc_5 VNB N_D1_c_69_n 0.0176283f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.07
cc_6 VNB N_D1_c_70_n 0.0022808f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.07
cc_7 VNB N_C1_M1003_g 0.020488f $X=-0.19 $Y=-0.245 $X2=0.68 $Y2=2.545
cc_8 VNB N_C1_c_103_n 0.0134953f $X=-0.19 $Y=-0.245 $X2=0.76 $Y2=0.905
cc_9 VNB N_C1_M1004_g 0.00442139f $X=-0.19 $Y=-0.245 $X2=0.76 $Y2=0.495
cc_10 VNB N_C1_c_105_n 0.023062f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.41
cc_11 VNB C1 0.00483595f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.575
cc_12 VNB N_C1_c_107_n 0.0163579f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_B1_M1007_g 0.0367131f $X=-0.19 $Y=-0.245 $X2=0.68 $Y2=2.545
cc_14 VNB N_B1_c_152_n 0.0209702f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.41
cc_15 VNB N_B1_c_153_n 0.0015918f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.575
cc_16 VNB B1 0.00809434f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_17 VNB N_B1_c_155_n 0.0153071f $X=-0.19 $Y=-0.245 $X2=0.675 $Y2=1.07
cc_18 VNB N_A2_M1009_g 0.0366539f $X=-0.19 $Y=-0.245 $X2=0.68 $Y2=2.545
cc_19 VNB N_A2_c_194_n 0.0015451f $X=-0.19 $Y=-0.245 $X2=0.76 $Y2=0.905
cc_20 VNB N_A2_c_195_n 0.0208897f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.41
cc_21 VNB N_A2_c_196_n 0.0152706f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.07
cc_22 VNB N_A2_c_197_n 0.00397284f $X=-0.19 $Y=-0.245 $X2=0.675 $Y2=1.07
cc_23 VNB N_A1_M1001_g 0.00849569f $X=-0.19 $Y=-0.245 $X2=0.68 $Y2=2.545
cc_24 VNB N_A1_M1005_g 0.0488934f $X=-0.19 $Y=-0.245 $X2=0.76 $Y2=0.495
cc_25 VNB A1 0.0127941f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.07
cc_26 VNB N_A1_c_237_n 0.0640223f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.07
cc_27 VNB N_VPWR_c_263_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB Y 0.047495f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_Y_c_305_n 0.0356539f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_347_57#_c_363_n 0.00465134f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.07
cc_31 VNB N_A_347_57#_c_364_n 0.0179167f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.41
cc_32 VNB N_A_347_57#_c_365_n 0.0119839f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.575
cc_33 VNB N_A_347_57#_c_366_n 0.0219254f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.07
cc_34 VNB N_VGND_c_390_n 0.00712414f $X=-0.19 $Y=-0.245 $X2=0.76 $Y2=0.495
cc_35 VNB N_VGND_c_391_n 0.0650376f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=1.07
cc_36 VNB N_VGND_c_392_n 0.00632158f $X=-0.19 $Y=-0.245 $X2=0.67 $Y2=0.905
cc_37 VNB N_VGND_c_393_n 0.0220291f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_394_n 0.224795f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VPB N_D1_M1008_g 0.0465431f $X=-0.19 $Y=1.655 $X2=0.68 $Y2=2.545
cc_40 VPB N_C1_M1004_g 0.0388167f $X=-0.19 $Y=1.655 $X2=0.76 $Y2=0.495
cc_41 VPB N_B1_M1006_g 0.0310667f $X=-0.19 $Y=1.655 $X2=0.76 $Y2=0.495
cc_42 VPB N_B1_c_153_n 0.0111706f $X=-0.19 $Y=1.655 $X2=0.67 $Y2=1.575
cc_43 VPB B1 0.00231208f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_44 VPB N_A2_c_194_n 0.0109074f $X=-0.19 $Y=1.655 $X2=0.76 $Y2=0.905
cc_45 VPB N_A2_M1000_g 0.0312512f $X=-0.19 $Y=1.655 $X2=0.76 $Y2=0.495
cc_46 VPB N_A2_c_197_n 0.0105362f $X=-0.19 $Y=1.655 $X2=0.675 $Y2=1.07
cc_47 VPB N_A1_M1001_g 0.0491548f $X=-0.19 $Y=1.655 $X2=0.68 $Y2=2.545
cc_48 VPB A1 0.0110329f $X=-0.19 $Y=1.655 $X2=0.67 $Y2=1.07
cc_49 VPB N_VPWR_c_264_n 0.0156631f $X=-0.19 $Y=1.655 $X2=0.67 $Y2=0.905
cc_50 VPB N_VPWR_c_265_n 0.0408332f $X=-0.19 $Y=1.655 $X2=0.67 $Y2=1.575
cc_51 VPB N_VPWR_c_266_n 0.00177638f $X=-0.19 $Y=1.655 $X2=0.67 $Y2=1.07
cc_52 VPB N_VPWR_c_267_n 0.0121543f $X=-0.19 $Y=1.655 $X2=0.675 $Y2=1.07
cc_53 VPB N_VPWR_c_268_n 0.0467569f $X=-0.19 $Y=1.655 $X2=0.675 $Y2=1.295
cc_54 VPB N_VPWR_c_269_n 0.0187052f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_55 VPB N_VPWR_c_270_n 0.00497896f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_56 VPB N_VPWR_c_271_n 0.0352526f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_57 VPB N_VPWR_c_263_n 0.0656967f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_58 VPB N_Y_c_306_n 0.0084465f $X=-0.19 $Y=1.655 $X2=0.67 $Y2=0.905
cc_59 VPB N_Y_c_307_n 0.0140157f $X=-0.19 $Y=1.655 $X2=0.67 $Y2=1.41
cc_60 VPB N_Y_c_308_n 0.00207453f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_61 VPB N_Y_c_309_n 0.0165171f $X=-0.19 $Y=1.655 $X2=0.675 $Y2=1.07
cc_62 VPB N_Y_c_310_n 0.00207453f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_63 VPB N_Y_c_311_n 0.00906423f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_64 VPB Y 0.00579578f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_65 N_D1_M1002_g N_C1_M1003_g 0.0396059f $X=0.76 $Y=0.495 $X2=0 $Y2=0
cc_66 N_D1_M1008_g N_C1_c_103_n 5.52405e-19 $X=0.68 $Y=2.545 $X2=0 $Y2=0
cc_67 N_D1_c_68_n N_C1_c_103_n 0.0133663f $X=0.67 $Y=1.575 $X2=0 $Y2=0
cc_68 N_D1_M1008_g N_C1_M1004_g 0.0289416f $X=0.68 $Y=2.545 $X2=0 $Y2=0
cc_69 N_D1_c_67_n N_C1_c_105_n 0.0133663f $X=0.67 $Y=1.41 $X2=0 $Y2=0
cc_70 N_D1_M1002_g C1 0.00488832f $X=0.76 $Y=0.495 $X2=0 $Y2=0
cc_71 N_D1_c_69_n C1 0.00229175f $X=0.67 $Y=1.07 $X2=0 $Y2=0
cc_72 N_D1_c_70_n C1 0.042276f $X=0.67 $Y=1.07 $X2=0 $Y2=0
cc_73 N_D1_c_69_n N_C1_c_107_n 0.0133663f $X=0.67 $Y=1.07 $X2=0 $Y2=0
cc_74 N_D1_c_70_n N_C1_c_107_n 0.00229208f $X=0.67 $Y=1.07 $X2=0 $Y2=0
cc_75 N_D1_M1008_g N_VPWR_c_265_n 0.0264607f $X=0.68 $Y=2.545 $X2=0 $Y2=0
cc_76 N_D1_M1008_g N_VPWR_c_266_n 8.61967e-19 $X=0.68 $Y=2.545 $X2=0 $Y2=0
cc_77 N_D1_M1008_g N_VPWR_c_269_n 0.00769046f $X=0.68 $Y=2.545 $X2=0 $Y2=0
cc_78 N_D1_M1008_g N_VPWR_c_263_n 0.0134474f $X=0.68 $Y=2.545 $X2=0 $Y2=0
cc_79 N_D1_M1008_g N_Y_c_306_n 0.0202065f $X=0.68 $Y=2.545 $X2=0 $Y2=0
cc_80 N_D1_c_68_n N_Y_c_306_n 7.0787e-19 $X=0.67 $Y=1.575 $X2=0 $Y2=0
cc_81 N_D1_c_70_n N_Y_c_306_n 0.0185116f $X=0.67 $Y=1.07 $X2=0 $Y2=0
cc_82 N_D1_M1008_g N_Y_c_308_n 0.0164995f $X=0.68 $Y=2.545 $X2=0 $Y2=0
cc_83 N_D1_M1008_g N_Y_c_311_n 0.0131612f $X=0.68 $Y=2.545 $X2=0 $Y2=0
cc_84 N_D1_c_68_n N_Y_c_311_n 2.23711e-19 $X=0.67 $Y=1.575 $X2=0 $Y2=0
cc_85 N_D1_c_70_n N_Y_c_311_n 0.00422809f $X=0.67 $Y=1.07 $X2=0 $Y2=0
cc_86 N_D1_M1008_g Y 0.00666089f $X=0.68 $Y=2.545 $X2=0 $Y2=0
cc_87 N_D1_M1002_g Y 0.00520357f $X=0.76 $Y=0.495 $X2=0 $Y2=0
cc_88 N_D1_c_69_n Y 0.0151382f $X=0.67 $Y=1.07 $X2=0 $Y2=0
cc_89 N_D1_c_70_n Y 0.0488376f $X=0.67 $Y=1.07 $X2=0 $Y2=0
cc_90 N_D1_M1002_g N_Y_c_305_n 0.00930927f $X=0.76 $Y=0.495 $X2=0 $Y2=0
cc_91 N_D1_c_69_n N_Y_c_305_n 0.00175544f $X=0.67 $Y=1.07 $X2=0 $Y2=0
cc_92 N_D1_c_70_n N_Y_c_305_n 0.0158642f $X=0.67 $Y=1.07 $X2=0 $Y2=0
cc_93 N_D1_M1002_g N_VGND_c_391_n 0.00501304f $X=0.76 $Y=0.495 $X2=0 $Y2=0
cc_94 N_D1_M1002_g N_VGND_c_394_n 0.0102203f $X=0.76 $Y=0.495 $X2=0 $Y2=0
cc_95 N_C1_M1003_g N_B1_M1007_g 0.0242392f $X=1.15 $Y=0.495 $X2=0 $Y2=0
cc_96 C1 N_B1_M1007_g 0.00567023f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_97 N_C1_c_107_n N_B1_M1007_g 0.0140242f $X=1.21 $Y=1.08 $X2=0 $Y2=0
cc_98 N_C1_M1004_g N_B1_M1006_g 0.0280117f $X=1.21 $Y=2.545 $X2=0 $Y2=0
cc_99 N_C1_c_103_n N_B1_c_152_n 0.0140242f $X=1.21 $Y=1.585 $X2=0 $Y2=0
cc_100 N_C1_M1004_g N_B1_c_152_n 0.0103561f $X=1.21 $Y=2.545 $X2=0 $Y2=0
cc_101 N_C1_M1004_g B1 0.00422732f $X=1.21 $Y=2.545 $X2=0 $Y2=0
cc_102 N_C1_c_105_n B1 0.00261922f $X=1.21 $Y=1.42 $X2=0 $Y2=0
cc_103 C1 B1 0.0335368f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_104 N_C1_c_105_n N_B1_c_155_n 0.0140242f $X=1.21 $Y=1.42 $X2=0 $Y2=0
cc_105 C1 N_B1_c_155_n 5.55455e-19 $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_106 N_C1_M1004_g N_VPWR_c_265_n 9.15489e-19 $X=1.21 $Y=2.545 $X2=0 $Y2=0
cc_107 N_C1_M1004_g N_VPWR_c_266_n 0.0175325f $X=1.21 $Y=2.545 $X2=0 $Y2=0
cc_108 N_C1_M1004_g N_VPWR_c_269_n 0.00769046f $X=1.21 $Y=2.545 $X2=0 $Y2=0
cc_109 N_C1_M1004_g N_VPWR_c_263_n 0.0134474f $X=1.21 $Y=2.545 $X2=0 $Y2=0
cc_110 N_C1_M1004_g N_Y_c_308_n 0.0165272f $X=1.21 $Y=2.545 $X2=0 $Y2=0
cc_111 N_C1_c_103_n N_Y_c_309_n 2.2693e-19 $X=1.21 $Y=1.585 $X2=0 $Y2=0
cc_112 N_C1_M1004_g N_Y_c_309_n 0.0202254f $X=1.21 $Y=2.545 $X2=0 $Y2=0
cc_113 C1 N_Y_c_309_n 0.01043f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_114 N_C1_M1004_g N_Y_c_310_n 9.16915e-19 $X=1.21 $Y=2.545 $X2=0 $Y2=0
cc_115 N_C1_c_103_n N_Y_c_311_n 3.03059e-19 $X=1.21 $Y=1.585 $X2=0 $Y2=0
cc_116 N_C1_M1004_g N_Y_c_311_n 0.00881339f $X=1.21 $Y=2.545 $X2=0 $Y2=0
cc_117 C1 N_Y_c_311_n 0.00526868f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_118 N_C1_M1003_g N_Y_c_305_n 0.00114658f $X=1.15 $Y=0.495 $X2=0 $Y2=0
cc_119 C1 N_Y_c_305_n 0.0072428f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_120 C1 A_245_57# 0.0046535f $X=1.115 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_121 C1 N_A_347_57#_c_363_n 0.0138553f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_122 C1 N_A_347_57#_c_365_n 0.00779855f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_123 N_C1_M1003_g N_VGND_c_391_n 0.00357038f $X=1.15 $Y=0.495 $X2=0 $Y2=0
cc_124 C1 N_VGND_c_391_n 0.00887369f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_125 N_C1_M1003_g N_VGND_c_394_n 0.00514204f $X=1.15 $Y=0.495 $X2=0 $Y2=0
cc_126 C1 N_VGND_c_394_n 0.0106888f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_127 N_B1_M1007_g N_A2_M1009_g 0.0195403f $X=1.66 $Y=0.495 $X2=0 $Y2=0
cc_128 N_B1_c_153_n N_A2_c_194_n 0.0135932f $X=1.75 $Y=1.795 $X2=0 $Y2=0
cc_129 N_B1_M1006_g N_A2_M1000_g 0.0195065f $X=1.76 $Y=2.545 $X2=0 $Y2=0
cc_130 N_B1_c_152_n N_A2_c_195_n 0.0135932f $X=1.75 $Y=1.63 $X2=0 $Y2=0
cc_131 B1 N_A2_c_196_n 0.00229184f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_132 N_B1_c_155_n N_A2_c_196_n 0.0135932f $X=1.75 $Y=1.29 $X2=0 $Y2=0
cc_133 B1 N_A2_c_197_n 0.0429487f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_134 N_B1_c_155_n N_A2_c_197_n 0.00233801f $X=1.75 $Y=1.29 $X2=0 $Y2=0
cc_135 N_B1_M1006_g N_VPWR_c_266_n 0.0157399f $X=1.76 $Y=2.545 $X2=0 $Y2=0
cc_136 N_B1_M1006_g N_VPWR_c_271_n 0.00840515f $X=1.76 $Y=2.545 $X2=0 $Y2=0
cc_137 N_B1_M1006_g N_VPWR_c_263_n 0.0146909f $X=1.76 $Y=2.545 $X2=0 $Y2=0
cc_138 N_B1_M1006_g N_Y_c_309_n 0.0200895f $X=1.76 $Y=2.545 $X2=0 $Y2=0
cc_139 N_B1_c_153_n N_Y_c_309_n 0.00101348f $X=1.75 $Y=1.795 $X2=0 $Y2=0
cc_140 B1 N_Y_c_309_n 0.0253127f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_141 N_B1_M1006_g N_Y_c_310_n 0.0170706f $X=1.76 $Y=2.545 $X2=0 $Y2=0
cc_142 N_B1_M1006_g N_Y_c_311_n 0.00154414f $X=1.76 $Y=2.545 $X2=0 $Y2=0
cc_143 B1 N_Y_c_311_n 0.00113935f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_144 N_B1_M1007_g N_A_347_57#_c_363_n 0.00930011f $X=1.66 $Y=0.495 $X2=0 $Y2=0
cc_145 N_B1_M1007_g N_A_347_57#_c_365_n 0.0024319f $X=1.66 $Y=0.495 $X2=0 $Y2=0
cc_146 B1 N_A_347_57#_c_365_n 0.00886827f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_147 N_B1_c_155_n N_A_347_57#_c_365_n 0.00132232f $X=1.75 $Y=1.29 $X2=0 $Y2=0
cc_148 N_B1_M1007_g N_VGND_c_391_n 0.0053602f $X=1.66 $Y=0.495 $X2=0 $Y2=0
cc_149 N_B1_M1007_g N_VGND_c_394_n 0.010796f $X=1.66 $Y=0.495 $X2=0 $Y2=0
cc_150 N_A2_M1000_g N_A1_M1001_g 0.074134f $X=2.29 $Y=2.545 $X2=0 $Y2=0
cc_151 N_A2_c_195_n N_A1_M1001_g 0.0199228f $X=2.29 $Y=1.63 $X2=0 $Y2=0
cc_152 N_A2_c_197_n N_A1_M1001_g 0.0120906f $X=2.29 $Y=1.29 $X2=0 $Y2=0
cc_153 N_A2_M1009_g N_A1_M1005_g 0.0234983f $X=2.23 $Y=0.495 $X2=0 $Y2=0
cc_154 N_A2_c_196_n N_A1_M1005_g 0.00298571f $X=2.29 $Y=1.29 $X2=0 $Y2=0
cc_155 N_A2_c_197_n N_A1_M1005_g 0.00390516f $X=2.29 $Y=1.29 $X2=0 $Y2=0
cc_156 N_A2_c_197_n A1 0.0462577f $X=2.29 $Y=1.29 $X2=0 $Y2=0
cc_157 N_A2_c_196_n N_A1_c_237_n 0.0199228f $X=2.29 $Y=1.29 $X2=0 $Y2=0
cc_158 N_A2_c_197_n N_A1_c_237_n 0.0108506f $X=2.29 $Y=1.29 $X2=0 $Y2=0
cc_159 N_A2_M1000_g N_VPWR_c_266_n 8.4511e-19 $X=2.29 $Y=2.545 $X2=0 $Y2=0
cc_160 N_A2_M1000_g N_VPWR_c_268_n 0.00518086f $X=2.29 $Y=2.545 $X2=0 $Y2=0
cc_161 N_A2_M1000_g N_VPWR_c_271_n 0.0086001f $X=2.29 $Y=2.545 $X2=0 $Y2=0
cc_162 N_A2_M1000_g N_VPWR_c_263_n 0.0157455f $X=2.29 $Y=2.545 $X2=0 $Y2=0
cc_163 N_A2_c_194_n N_Y_c_309_n 3.03059e-19 $X=2.29 $Y=1.795 $X2=0 $Y2=0
cc_164 N_A2_M1000_g N_Y_c_309_n 0.00483326f $X=2.29 $Y=2.545 $X2=0 $Y2=0
cc_165 N_A2_c_197_n N_Y_c_309_n 0.00534367f $X=2.29 $Y=1.29 $X2=0 $Y2=0
cc_166 N_A2_M1000_g N_Y_c_310_n 0.0186168f $X=2.29 $Y=2.545 $X2=0 $Y2=0
cc_167 N_A2_M1009_g N_A_347_57#_c_363_n 0.00243751f $X=2.23 $Y=0.495 $X2=0 $Y2=0
cc_168 N_A2_M1009_g N_A_347_57#_c_364_n 0.012656f $X=2.23 $Y=0.495 $X2=0 $Y2=0
cc_169 N_A2_c_196_n N_A_347_57#_c_364_n 0.00120075f $X=2.29 $Y=1.29 $X2=0 $Y2=0
cc_170 N_A2_c_197_n N_A_347_57#_c_364_n 0.0472367f $X=2.29 $Y=1.29 $X2=0 $Y2=0
cc_171 N_A2_M1009_g N_A_347_57#_c_366_n 8.33917e-19 $X=2.23 $Y=0.495 $X2=0 $Y2=0
cc_172 N_A2_M1009_g N_VGND_c_390_n 0.00308327f $X=2.23 $Y=0.495 $X2=0 $Y2=0
cc_173 N_A2_M1009_g N_VGND_c_391_n 0.0053602f $X=2.23 $Y=0.495 $X2=0 $Y2=0
cc_174 N_A2_M1009_g N_VGND_c_394_n 0.00597178f $X=2.23 $Y=0.495 $X2=0 $Y2=0
cc_175 N_A1_M1001_g N_VPWR_c_268_n 0.0277664f $X=2.79 $Y=2.545 $X2=0 $Y2=0
cc_176 A1 N_VPWR_c_268_n 0.0210234f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_177 N_A1_c_237_n N_VPWR_c_268_n 0.00165559f $X=3.09 $Y=1.345 $X2=0 $Y2=0
cc_178 N_A1_M1001_g N_VPWR_c_271_n 0.00802402f $X=2.79 $Y=2.545 $X2=0 $Y2=0
cc_179 N_A1_M1001_g N_VPWR_c_263_n 0.0142844f $X=2.79 $Y=2.545 $X2=0 $Y2=0
cc_180 N_A1_M1001_g N_Y_c_309_n 7.27634e-19 $X=2.79 $Y=2.545 $X2=0 $Y2=0
cc_181 N_A1_M1001_g N_Y_c_310_n 0.0039712f $X=2.79 $Y=2.545 $X2=0 $Y2=0
cc_182 N_A1_M1005_g N_A_347_57#_c_364_n 0.0162895f $X=2.77 $Y=0.495 $X2=0 $Y2=0
cc_183 A1 N_A_347_57#_c_364_n 0.0155077f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_184 N_A1_c_237_n N_A_347_57#_c_364_n 0.00546259f $X=3.09 $Y=1.345 $X2=0 $Y2=0
cc_185 N_A1_M1005_g N_A_347_57#_c_366_n 0.0096335f $X=2.77 $Y=0.495 $X2=0 $Y2=0
cc_186 N_A1_M1005_g N_VGND_c_390_n 0.00454763f $X=2.77 $Y=0.495 $X2=0 $Y2=0
cc_187 N_A1_M1005_g N_VGND_c_393_n 0.00502664f $X=2.77 $Y=0.495 $X2=0 $Y2=0
cc_188 N_A1_M1005_g N_VGND_c_394_n 0.00642538f $X=2.77 $Y=0.495 $X2=0 $Y2=0
cc_189 N_VPWR_c_265_n N_Y_c_306_n 0.0166661f $X=0.415 $Y=2.28 $X2=0 $Y2=0
cc_190 N_VPWR_c_265_n N_Y_c_307_n 0.00739446f $X=0.415 $Y=2.28 $X2=0 $Y2=0
cc_191 N_VPWR_c_266_n N_Y_c_308_n 0.0487591f $X=1.475 $Y=2.49 $X2=0 $Y2=0
cc_192 N_VPWR_c_269_n N_Y_c_308_n 0.021949f $X=1.31 $Y=3.33 $X2=0 $Y2=0
cc_193 N_VPWR_c_263_n N_Y_c_308_n 0.0124703f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_194 N_VPWR_M1004_d N_Y_c_309_n 0.00202522f $X=1.335 $Y=2.045 $X2=0 $Y2=0
cc_195 N_VPWR_c_266_n N_Y_c_309_n 0.0164557f $X=1.475 $Y=2.49 $X2=0 $Y2=0
cc_196 N_VPWR_c_266_n N_Y_c_310_n 0.0451886f $X=1.475 $Y=2.49 $X2=0 $Y2=0
cc_197 N_VPWR_c_271_n N_Y_c_310_n 0.021949f $X=2.89 $Y=3.33 $X2=0 $Y2=0
cc_198 N_VPWR_c_263_n N_Y_c_310_n 0.0124703f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_199 N_VPWR_c_265_n N_Y_c_311_n 0.0625632f $X=0.415 $Y=2.28 $X2=0 $Y2=0
cc_200 N_Y_c_305_n N_VGND_c_391_n 0.0379902f $X=0.545 $Y=0.495 $X2=0 $Y2=0
cc_201 N_Y_c_305_n N_VGND_c_394_n 0.0222729f $X=0.545 $Y=0.495 $X2=0 $Y2=0
cc_202 N_A_347_57#_c_363_n N_VGND_c_390_n 0.00151838f $X=1.965 $Y=0.495 $X2=0
+ $Y2=0
cc_203 N_A_347_57#_c_364_n N_VGND_c_390_n 0.0229108f $X=2.82 $Y=0.86 $X2=0 $Y2=0
cc_204 N_A_347_57#_c_366_n N_VGND_c_390_n 0.0125869f $X=2.985 $Y=0.495 $X2=0
+ $Y2=0
cc_205 N_A_347_57#_c_363_n N_VGND_c_391_n 0.0221152f $X=1.965 $Y=0.495 $X2=0
+ $Y2=0
cc_206 N_A_347_57#_c_366_n N_VGND_c_393_n 0.0220321f $X=2.985 $Y=0.495 $X2=0
+ $Y2=0
cc_207 N_A_347_57#_c_363_n N_VGND_c_394_n 0.0126914f $X=1.965 $Y=0.495 $X2=0
+ $Y2=0
cc_208 N_A_347_57#_c_364_n N_VGND_c_394_n 0.0124074f $X=2.82 $Y=0.86 $X2=0 $Y2=0
cc_209 N_A_347_57#_c_366_n N_VGND_c_394_n 0.0125808f $X=2.985 $Y=0.495 $X2=0
+ $Y2=0
