* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
X0 a_115_367# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X1 VGND A1 a_32_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X2 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X3 Y B1 a_32_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X4 a_115_367# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X5 Y B1 a_32_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X6 a_32_47# B1 Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X7 a_32_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X8 VGND A2 a_32_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X9 Y A2 a_115_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X10 VPWR A1 a_115_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X11 VPWR A1 a_115_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X12 a_32_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X13 a_115_367# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X14 a_32_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X15 VGND A2 a_32_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X16 a_32_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X17 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X18 Y B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X19 VPWR B1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X20 VGND A1 a_32_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X21 a_115_367# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X22 Y A2 a_115_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X23 a_32_47# B1 Y VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
.ends
