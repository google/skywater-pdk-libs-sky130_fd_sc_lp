* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__dlybuf4s50kapwr_1 A KAPWR VGND VNB VPB VPWR X
X0 KAPWR a_27_52# a_282_52# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=500000u
X1 a_394_52# a_282_52# VGND VNB sky130_fd_pr__nfet_01v8 w=1e+06u l=500000u
X2 a_27_52# A KAPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X3 a_27_52# A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 VGND a_394_52# X VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 KAPWR a_394_52# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X6 a_394_52# a_282_52# KAPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=500000u
X7 VGND a_27_52# a_282_52# VNB sky130_fd_pr__nfet_01v8 w=1e+06u l=500000u
.ends
