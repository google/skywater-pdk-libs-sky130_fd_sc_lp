* File: sky130_fd_sc_lp__o41a_1.pex.spice
* Created: Wed Sep  2 10:27:26 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O41A_1%A_155_23# 1 2 7 9 12 15 18 20 21 22 24 29 36
c53 36 0 1.35206e-19 $X=1.035 $Y=1.36
r54 28 36 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=0.945 $Y=1.36
+ $X2=1.035 $Y2=1.36
r55 28 33 16.6118 $w=3.3e-07 $l=9.5e-08 $layer=POLY_cond $X=0.945 $Y=1.36
+ $X2=0.85 $Y2=1.36
r56 27 29 11.8695 $w=4.06e-07 $l=3.95e-07 $layer=LI1_cond $X=0.945 $Y=1.26
+ $X2=1.34 $Y2=1.26
r57 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.945
+ $Y=1.36 $X2=0.945 $Y2=1.36
r58 22 32 2.93179 $w=2.5e-07 $l=8.8e-08 $layer=LI1_cond $X=1.78 $Y=2.1 $X2=1.78
+ $Y2=2.012
r59 22 24 37.3392 $w=2.48e-07 $l=8.1e-07 $layer=LI1_cond $X=1.78 $Y=2.1 $X2=1.78
+ $Y2=2.91
r60 20 32 4.16448 $w=1.75e-07 $l=1.25e-07 $layer=LI1_cond $X=1.655 $Y=2.012
+ $X2=1.78 $Y2=2.012
r61 20 21 14.5766 $w=1.73e-07 $l=2.3e-07 $layer=LI1_cond $X=1.655 $Y=2.012
+ $X2=1.425 $Y2=2.012
r62 16 29 6.76108 $w=4.06e-07 $l=3.60347e-07 $layer=LI1_cond $X=1.565 $Y=0.995
+ $X2=1.34 $Y2=1.26
r63 16 18 22.8502 $w=2.88e-07 $l=5.75e-07 $layer=LI1_cond $X=1.565 $Y=0.995
+ $X2=1.565 $Y2=0.42
r64 15 21 6.81835 $w=1.75e-07 $l=1.22327e-07 $layer=LI1_cond $X=1.34 $Y=1.925
+ $X2=1.425 $Y2=2.012
r65 14 29 5.869 $w=1.7e-07 $l=2.65e-07 $layer=LI1_cond $X=1.34 $Y=1.525 $X2=1.34
+ $Y2=1.26
r66 14 15 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=1.34 $Y=1.525 $X2=1.34
+ $Y2=1.925
r67 10 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.035 $Y=1.525
+ $X2=1.035 $Y2=1.36
r68 10 12 482 $w=1.5e-07 $l=9.4e-07 $layer=POLY_cond $X=1.035 $Y=1.525 $X2=1.035
+ $Y2=2.465
r69 7 33 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.85 $Y=1.195
+ $X2=0.85 $Y2=1.36
r70 7 9 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.85 $Y=1.195 $X2=0.85
+ $Y2=0.665
r71 2 32 400 $w=1.7e-07 $l=3.17372e-07 $layer=licon1_PDIFF $count=1 $X=1.68
+ $Y=1.835 $X2=1.82 $Y2=2.09
r72 2 24 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=1.68
+ $Y=1.835 $X2=1.82 $Y2=2.91
r73 1 18 91 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_NDIFF $count=2 $X=1.46
+ $Y=0.245 $X2=1.585 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__O41A_1%B1 3 7 9 15 16
c35 15 0 1.35206e-19 $X=1.71 $Y=1.51
r36 14 16 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=1.71 $Y=1.51 $X2=1.8
+ $Y2=1.51
r37 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.71
+ $Y=1.51 $X2=1.71 $Y2=1.51
r38 11 14 18.3604 $w=3.3e-07 $l=1.05e-07 $layer=POLY_cond $X=1.605 $Y=1.51
+ $X2=1.71 $Y2=1.51
r39 9 15 5.76222 $w=3.08e-07 $l=1.55e-07 $layer=LI1_cond $X=1.75 $Y=1.665
+ $X2=1.75 $Y2=1.51
r40 5 16 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.8 $Y=1.345 $X2=1.8
+ $Y2=1.51
r41 5 7 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=1.8 $Y=1.345 $X2=1.8
+ $Y2=0.665
r42 1 11 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.605 $Y=1.675
+ $X2=1.605 $Y2=1.51
r43 1 3 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.605 $Y=1.675
+ $X2=1.605 $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__O41A_1%A4 3 7 9 10 11 12 18 19
r38 18 21 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.25 $Y=1.51
+ $X2=2.25 $Y2=1.675
r39 18 20 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.25 $Y=1.51
+ $X2=2.25 $Y2=1.345
r40 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.25
+ $Y=1.51 $X2=2.25 $Y2=1.51
r41 11 12 16.4002 $w=2.58e-07 $l=3.7e-07 $layer=LI1_cond $X=2.205 $Y=2.405
+ $X2=2.205 $Y2=2.775
r42 10 11 16.4002 $w=2.58e-07 $l=3.7e-07 $layer=LI1_cond $X=2.205 $Y=2.035
+ $X2=2.205 $Y2=2.405
r43 9 10 16.4002 $w=2.58e-07 $l=3.7e-07 $layer=LI1_cond $X=2.205 $Y=1.665
+ $X2=2.205 $Y2=2.035
r44 9 19 6.87033 $w=2.58e-07 $l=1.55e-07 $layer=LI1_cond $X=2.205 $Y=1.665
+ $X2=2.205 $Y2=1.51
r45 7 20 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=2.23 $Y=0.665
+ $X2=2.23 $Y2=1.345
r46 3 21 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.16 $Y=2.465
+ $X2=2.16 $Y2=1.675
.ends

.subckt PM_SKY130_FD_SC_LP__O41A_1%A3 3 7 9 10 11 12 18 19
r39 18 20 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.79 $Y=1.51
+ $X2=2.79 $Y2=1.345
r40 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.79
+ $Y=1.51 $X2=2.79 $Y2=1.51
r41 11 12 9.83442 $w=4.48e-07 $l=3.7e-07 $layer=LI1_cond $X=2.73 $Y=2.405
+ $X2=2.73 $Y2=2.775
r42 10 11 9.83442 $w=4.48e-07 $l=3.7e-07 $layer=LI1_cond $X=2.73 $Y=2.035
+ $X2=2.73 $Y2=2.405
r43 9 10 9.83442 $w=4.48e-07 $l=3.7e-07 $layer=LI1_cond $X=2.73 $Y=1.665
+ $X2=2.73 $Y2=2.035
r44 9 19 4.11983 $w=4.48e-07 $l=1.55e-07 $layer=LI1_cond $X=2.73 $Y=1.665
+ $X2=2.73 $Y2=1.51
r45 7 20 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=2.81 $Y=0.665
+ $X2=2.81 $Y2=1.345
r46 1 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.79 $Y=1.675
+ $X2=2.79 $Y2=1.51
r47 1 3 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.79 $Y=1.675 $X2=2.79
+ $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__O41A_1%A2 3 7 9 10 11 12 19 20 36
c36 20 0 1.17498e-19 $X=3.33 $Y=1.51
r37 36 37 0.77464 $w=5.28e-07 $l=1e-08 $layer=LI1_cond $X=3.43 $Y=1.665 $X2=3.43
+ $Y2=1.675
r38 19 22 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.33 $Y=1.51
+ $X2=3.33 $Y2=1.675
r39 19 21 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.33 $Y=1.51
+ $X2=3.33 $Y2=1.345
r40 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.33
+ $Y=1.51 $X2=3.33 $Y2=1.51
r41 11 12 10.1525 $w=4.18e-07 $l=3.7e-07 $layer=LI1_cond $X=3.485 $Y=2.405
+ $X2=3.485 $Y2=2.775
r42 10 11 10.1525 $w=4.18e-07 $l=3.7e-07 $layer=LI1_cond $X=3.485 $Y=2.035
+ $X2=3.485 $Y2=2.405
r43 9 36 0.857566 $w=5.28e-07 $l=3.8e-08 $layer=LI1_cond $X=3.43 $Y=1.627
+ $X2=3.43 $Y2=1.665
r44 9 20 2.6404 $w=5.28e-07 $l=1.17e-07 $layer=LI1_cond $X=3.43 $Y=1.627
+ $X2=3.43 $Y2=1.51
r45 9 10 8.86284 $w=4.18e-07 $l=3.23e-07 $layer=LI1_cond $X=3.485 $Y=1.712
+ $X2=3.485 $Y2=2.035
r46 9 37 1.01525 $w=4.18e-07 $l=3.7e-08 $layer=LI1_cond $X=3.485 $Y=1.712
+ $X2=3.485 $Y2=1.675
r47 7 22 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.24 $Y=2.465
+ $X2=3.24 $Y2=1.675
r48 3 21 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=3.24 $Y=0.665
+ $X2=3.24 $Y2=1.345
.ends

.subckt PM_SKY130_FD_SC_LP__O41A_1%A1 3 7 9 14 15
r25 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.03
+ $Y=1.46 $X2=4.03 $Y2=1.46
r26 11 14 43.7153 $w=3.3e-07 $l=2.5e-07 $layer=POLY_cond $X=3.78 $Y=1.46
+ $X2=4.03 $Y2=1.46
r27 9 15 6.38516 $w=3.68e-07 $l=2.05e-07 $layer=LI1_cond $X=4.05 $Y=1.665
+ $X2=4.05 $Y2=1.46
r28 5 11 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.78 $Y=1.625
+ $X2=3.78 $Y2=1.46
r29 5 7 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=3.78 $Y=1.625 $X2=3.78
+ $Y2=2.465
r30 1 11 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.78 $Y=1.295
+ $X2=3.78 $Y2=1.46
r31 1 3 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=3.78 $Y=1.295 $X2=3.78
+ $Y2=0.665
.ends

.subckt PM_SKY130_FD_SC_LP__O41A_1%X 1 2 7 8 9 10 11 12 13 30
r16 13 49 2.17569 $w=7.57e-07 $l=1.35e-07 $layer=LI1_cond $X=0.505 $Y=2.775
+ $X2=0.505 $Y2=2.91
r17 12 13 5.96301 $w=7.57e-07 $l=3.7e-07 $layer=LI1_cond $X=0.505 $Y=2.405
+ $X2=0.505 $Y2=2.775
r18 11 12 5.96301 $w=7.57e-07 $l=3.7e-07 $layer=LI1_cond $X=0.505 $Y=2.035
+ $X2=0.505 $Y2=2.405
r19 11 41 0.886394 $w=7.57e-07 $l=5.5e-08 $layer=LI1_cond $X=0.505 $Y=2.035
+ $X2=0.505 $Y2=1.98
r20 10 41 5.07662 $w=7.57e-07 $l=3.15e-07 $layer=LI1_cond $X=0.505 $Y=1.665
+ $X2=0.505 $Y2=1.98
r21 10 23 6.41412 $w=7.57e-07 $l=3.30454e-07 $layer=LI1_cond $X=0.505 $Y=1.665
+ $X2=0.29 $Y2=1.425
r22 9 23 3.65409 $w=4.08e-07 $l=1.3e-07 $layer=LI1_cond $X=0.29 $Y=1.295
+ $X2=0.29 $Y2=1.425
r23 8 9 10.4001 $w=4.08e-07 $l=3.7e-07 $layer=LI1_cond $X=0.29 $Y=0.925 $X2=0.29
+ $Y2=1.295
r24 7 8 6.06384 $w=6.43e-07 $l=3.27e-07 $layer=LI1_cond $X=0.407 $Y=0.555
+ $X2=0.407 $Y2=0.882
r25 7 30 2.8743 $w=6.43e-07 $l=1.55e-07 $layer=LI1_cond $X=0.407 $Y=0.555
+ $X2=0.407 $Y2=0.4
r26 2 49 200 $w=1.7e-07 $l=1.13578e-06 $layer=licon1_PDIFF $count=3 $X=0.355
+ $Y=1.835 $X2=0.48 $Y2=2.91
r27 2 41 200 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=3 $X=0.355
+ $Y=1.835 $X2=0.48 $Y2=1.98
r28 1 30 91 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=2 $X=0.17
+ $Y=0.245 $X2=0.295 $Y2=0.4
r29 1 8 91 $w=1.7e-07 $l=7.54917e-07 $layer=licon1_NDIFF $count=2 $X=0.17
+ $Y=0.245 $X2=0.295 $Y2=0.94
.ends

.subckt PM_SKY130_FD_SC_LP__O41A_1%VPWR 1 2 9 11 13 17 19 24 33 37
r45 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r46 33 34 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r47 31 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r48 30 31 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r49 28 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r50 27 30 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=1.68 $Y=3.33
+ $X2=3.6 $Y2=3.33
r51 27 28 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r52 25 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.485 $Y=3.33
+ $X2=1.32 $Y2=3.33
r53 25 27 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=1.485 $Y=3.33
+ $X2=1.68 $Y2=3.33
r54 24 36 4.3301 $w=1.7e-07 $l=2.27e-07 $layer=LI1_cond $X=3.865 $Y=3.33
+ $X2=4.092 $Y2=3.33
r55 24 30 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=3.865 $Y=3.33
+ $X2=3.6 $Y2=3.33
r56 22 34 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.2 $Y2=3.33
r57 21 22 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r58 19 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.155 $Y=3.33
+ $X2=1.32 $Y2=3.33
r59 19 21 59.6952 $w=1.68e-07 $l=9.15e-07 $layer=LI1_cond $X=1.155 $Y=3.33
+ $X2=0.24 $Y2=3.33
r60 17 31 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.6 $Y2=3.33
r61 17 28 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r62 13 16 33.792 $w=2.93e-07 $l=8.65e-07 $layer=LI1_cond $X=4.012 $Y=2.085
+ $X2=4.012 $Y2=2.95
r63 11 36 3.14743 $w=2.95e-07 $l=1.18427e-07 $layer=LI1_cond $X=4.012 $Y=3.245
+ $X2=4.092 $Y2=3.33
r64 11 16 11.5244 $w=2.93e-07 $l=2.95e-07 $layer=LI1_cond $X=4.012 $Y=3.245
+ $X2=4.012 $Y2=2.95
r65 7 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.32 $Y=3.245 $X2=1.32
+ $Y2=3.33
r66 7 9 29.8588 $w=3.28e-07 $l=8.55e-07 $layer=LI1_cond $X=1.32 $Y=3.245
+ $X2=1.32 $Y2=2.39
r67 2 16 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=3.855
+ $Y=1.835 $X2=3.995 $Y2=2.95
r68 2 13 400 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_PDIFF $count=1 $X=3.855
+ $Y=1.835 $X2=3.995 $Y2=2.085
r69 1 9 300 $w=1.7e-07 $l=6.51594e-07 $layer=licon1_PDIFF $count=2 $X=1.11
+ $Y=1.835 $X2=1.32 $Y2=2.39
.ends

.subckt PM_SKY130_FD_SC_LP__O41A_1%VGND 1 2 3 12 16 20 23 24 25 27 36 42 43 46
+ 49
r52 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r53 46 47 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r54 43 50 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.6
+ $Y2=0
r55 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r56 40 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.69 $Y=0 $X2=3.525
+ $Y2=0
r57 40 42 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=3.69 $Y=0 $X2=4.08
+ $Y2=0
r58 39 50 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r59 38 39 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r60 36 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.36 $Y=0 $X2=3.525
+ $Y2=0
r61 36 38 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=3.36 $Y=0 $X2=3.12
+ $Y2=0
r62 32 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.23 $Y=0 $X2=1.065
+ $Y2=0
r63 32 34 60.6738 $w=1.68e-07 $l=9.3e-07 $layer=LI1_cond $X=1.23 $Y=0 $X2=2.16
+ $Y2=0
r64 30 47 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r65 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r66 27 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.9 $Y=0 $X2=1.065
+ $Y2=0
r67 27 29 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=0.9 $Y=0 $X2=0.72
+ $Y2=0
r68 25 39 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r69 25 47 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.2
+ $Y2=0
r70 25 34 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r71 23 34 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=2.35 $Y=0 $X2=2.16
+ $Y2=0
r72 23 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.35 $Y=0 $X2=2.515
+ $Y2=0
r73 22 38 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=2.68 $Y=0 $X2=3.12
+ $Y2=0
r74 22 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.68 $Y=0 $X2=2.515
+ $Y2=0
r75 18 49 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.525 $Y=0.085
+ $X2=3.525 $Y2=0
r76 18 20 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=3.525 $Y=0.085
+ $X2=3.525 $Y2=0.37
r77 14 24 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.515 $Y=0.085
+ $X2=2.515 $Y2=0
r78 14 16 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=2.515 $Y=0.085
+ $X2=2.515 $Y2=0.37
r79 10 46 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.065 $Y=0.085
+ $X2=1.065 $Y2=0
r80 10 12 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=1.065 $Y=0.085
+ $X2=1.065 $Y2=0.39
r81 3 20 91 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=2 $X=3.315
+ $Y=0.245 $X2=3.525 $Y2=0.37
r82 2 16 91 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=2 $X=2.305
+ $Y=0.245 $X2=2.515 $Y2=0.37
r83 1 12 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=0.925
+ $Y=0.245 $X2=1.065 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_LP__O41A_1%A_375_49# 1 2 3 12 14 15 18 20 24 26
r44 22 24 22.4726 $w=2.98e-07 $l=5.85e-07 $layer=LI1_cond $X=4.01 $Y=1.005
+ $X2=4.01 $Y2=0.42
r45 21 26 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.19 $Y=1.09
+ $X2=3.025 $Y2=1.09
r46 20 22 7.51767 $w=1.7e-07 $l=1.8775e-07 $layer=LI1_cond $X=3.86 $Y=1.09
+ $X2=4.01 $Y2=1.005
r47 20 21 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.86 $Y=1.09
+ $X2=3.19 $Y2=1.09
r48 16 26 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.025 $Y=1.005
+ $X2=3.025 $Y2=1.09
r49 16 18 20.4297 $w=3.28e-07 $l=5.85e-07 $layer=LI1_cond $X=3.025 $Y=1.005
+ $X2=3.025 $Y2=0.42
r50 14 26 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.86 $Y=1.09
+ $X2=3.025 $Y2=1.09
r51 14 15 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=2.86 $Y=1.09
+ $X2=2.15 $Y2=1.09
r52 10 15 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=2.015 $Y=1.005
+ $X2=2.15 $Y2=1.09
r53 10 12 24.9696 $w=2.68e-07 $l=5.85e-07 $layer=LI1_cond $X=2.015 $Y=1.005
+ $X2=2.015 $Y2=0.42
r54 3 24 91 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=2 $X=3.855
+ $Y=0.245 $X2=3.995 $Y2=0.42
r55 2 18 91 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=2 $X=2.885
+ $Y=0.245 $X2=3.025 $Y2=0.42
r56 1 12 91 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=2 $X=1.875
+ $Y=0.245 $X2=2.015 $Y2=0.42
.ends

