* File: sky130_fd_sc_lp__nor3b_lp.pex.spice
* Created: Wed Sep  2 10:09:56 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__NOR3B_LP%A 1 3 7 8 12 14 16 17 18 19 21 28 30
c43 28 0 1.89242e-19 $X=0.695 $Y=1.34
c44 8 0 7.83201e-20 $X=0.89 $Y=0.855
r45 28 30 45.9078 $w=4.1e-07 $l=1.65e-07 $layer=POLY_cond $X=0.735 $Y=1.34
+ $X2=0.735 $Y2=1.175
r46 21 28 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.695
+ $Y=1.34 $X2=0.695 $Y2=1.34
r47 19 21 8.12262 $w=6.68e-07 $l=4.55e-07 $layer=LI1_cond $X=0.24 $Y=1.51
+ $X2=0.695 $Y2=1.51
r48 14 16 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.965 $Y=0.78
+ $X2=0.965 $Y2=0.495
r49 12 18 173.918 $w=2.5e-07 $l=7e-07 $layer=POLY_cond $X=0.815 $Y=2.545
+ $X2=0.815 $Y2=1.845
r50 9 17 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.68 $Y=0.855
+ $X2=0.605 $Y2=0.855
r51 8 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.89 $Y=0.855
+ $X2=0.965 $Y2=0.78
r52 8 9 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=0.89 $Y=0.855 $X2=0.68
+ $Y2=0.855
r53 7 18 36.2176 $w=4.1e-07 $l=2.05e-07 $layer=POLY_cond $X=0.735 $Y=1.64
+ $X2=0.735 $Y2=1.845
r54 6 28 5.42589 $w=4.1e-07 $l=4e-08 $layer=POLY_cond $X=0.735 $Y=1.38 $X2=0.735
+ $Y2=1.34
r55 6 7 35.2683 $w=4.1e-07 $l=2.6e-07 $layer=POLY_cond $X=0.735 $Y=1.38
+ $X2=0.735 $Y2=1.64
r56 4 17 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.605 $Y=0.93
+ $X2=0.605 $Y2=0.855
r57 4 30 125.628 $w=1.5e-07 $l=2.45e-07 $layer=POLY_cond $X=0.605 $Y=0.93
+ $X2=0.605 $Y2=1.175
r58 1 17 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.605 $Y=0.78
+ $X2=0.605 $Y2=0.855
r59 1 3 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.605 $Y=0.78 $X2=0.605
+ $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__NOR3B_LP%B 3 5 7 10 12 14 16 17 18 19 20 21 22 23 24
+ 41
c63 16 0 1.89242e-19 $X=1.345 $Y=1.18
c64 10 0 6.10152e-20 $X=1.68 $Y=0.855
r65 41 42 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.345
+ $Y=1.345 $X2=1.345 $Y2=1.345
r66 23 24 6.23308 $w=7.08e-07 $l=3.7e-07 $layer=LI1_cond $X=1.44 $Y=2.405
+ $X2=1.44 $Y2=2.775
r67 22 23 6.23308 $w=7.08e-07 $l=3.7e-07 $layer=LI1_cond $X=1.44 $Y=2.035
+ $X2=1.44 $Y2=2.405
r68 21 22 6.23308 $w=7.08e-07 $l=3.7e-07 $layer=LI1_cond $X=1.44 $Y=1.665
+ $X2=1.44 $Y2=2.035
r69 21 42 5.39078 $w=7.08e-07 $l=3.2e-07 $layer=LI1_cond $X=1.44 $Y=1.665
+ $X2=1.44 $Y2=1.345
r70 20 42 0.842309 $w=7.08e-07 $l=5e-08 $layer=LI1_cond $X=1.44 $Y=1.295
+ $X2=1.44 $Y2=1.345
r71 17 41 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.345 $Y=1.685
+ $X2=1.345 $Y2=1.345
r72 17 18 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.345 $Y=1.685
+ $X2=1.345 $Y2=1.85
r73 16 41 40.8701 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.345 $Y=1.18
+ $X2=1.345 $Y2=1.345
r74 12 14 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=1.755 $Y=0.78
+ $X2=1.755 $Y2=0.495
r75 11 19 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.47 $Y=0.855
+ $X2=1.395 $Y2=0.855
r76 10 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.68 $Y=0.855
+ $X2=1.755 $Y2=0.78
r77 10 11 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=1.68 $Y=0.855
+ $X2=1.47 $Y2=0.855
r78 8 19 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.395 $Y=0.93
+ $X2=1.395 $Y2=0.855
r79 8 16 128.191 $w=1.5e-07 $l=2.5e-07 $layer=POLY_cond $X=1.395 $Y=0.93
+ $X2=1.395 $Y2=1.18
r80 5 19 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.395 $Y=0.78
+ $X2=1.395 $Y2=0.855
r81 5 7 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=1.395 $Y=0.78 $X2=1.395
+ $Y2=0.495
r82 3 18 172.675 $w=2.5e-07 $l=6.95e-07 $layer=POLY_cond $X=1.305 $Y=2.545
+ $X2=1.305 $Y2=1.85
.ends

.subckt PM_SKY130_FD_SC_LP__NOR3B_LP%A_350_269# 1 2 9 11 13 14 16 19 23 27 29 34
+ 35 36 37
c67 34 0 6.10152e-20 $X=2.49 $Y=0.99
r68 35 41 5.7257 $w=4.63e-07 $l=5.5e-08 $layer=POLY_cond $X=2.49 $Y=1.16
+ $X2=2.545 $Y2=1.16
r69 35 39 31.7516 $w=4.63e-07 $l=3.05e-07 $layer=POLY_cond $X=2.49 $Y=1.16
+ $X2=2.185 $Y2=1.16
r70 34 35 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.49
+ $Y=0.99 $X2=2.49 $Y2=0.99
r71 31 36 3.70735 $w=2.5e-07 $l=1.18427e-07 $layer=LI1_cond $X=3.63 $Y=0.995
+ $X2=3.55 $Y2=0.91
r72 31 37 67.1979 $w=1.68e-07 $l=1.03e-06 $layer=LI1_cond $X=3.63 $Y=0.995
+ $X2=3.63 $Y2=2.025
r73 27 37 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=3.55 $Y=2.19
+ $X2=3.55 $Y2=2.025
r74 27 29 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=3.55 $Y=2.19 $X2=3.55
+ $Y2=2.9
r75 21 36 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.55 $Y=0.825
+ $X2=3.55 $Y2=0.91
r76 21 23 11.5244 $w=3.28e-07 $l=3.3e-07 $layer=LI1_cond $X=3.55 $Y=0.825
+ $X2=3.55 $Y2=0.495
r77 20 34 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.655 $Y=0.91
+ $X2=2.49 $Y2=0.91
r78 19 36 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.385 $Y=0.91
+ $X2=3.55 $Y2=0.91
r79 19 20 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=3.385 $Y=0.91
+ $X2=2.655 $Y2=0.91
r80 14 41 29.4766 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=2.545 $Y=0.825
+ $X2=2.545 $Y2=1.16
r81 14 16 106.04 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=2.545 $Y=0.825
+ $X2=2.545 $Y2=0.495
r82 11 39 29.4766 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=2.185 $Y=0.825
+ $X2=2.185 $Y2=1.16
r83 11 13 106.04 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=2.185 $Y=0.825
+ $X2=2.185 $Y2=0.495
r84 7 39 32.2721 $w=4.63e-07 $l=4.64839e-07 $layer=POLY_cond $X=1.875 $Y=1.495
+ $X2=2.185 $Y2=1.16
r85 7 9 260.876 $w=2.5e-07 $l=1.05e-06 $layer=POLY_cond $X=1.875 $Y=1.495
+ $X2=1.875 $Y2=2.545
r86 2 29 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=3.41
+ $Y=2.045 $X2=3.55 $Y2=2.9
r87 2 27 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=3.41
+ $Y=2.045 $X2=3.55 $Y2=2.19
r88 1 23 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=3.41
+ $Y=0.285 $X2=3.55 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__NOR3B_LP%C_N 3 7 11 13 14 18
r34 18 20 66.9034 $w=5.1e-07 $l=5.05e-07 $layer=POLY_cond $X=3.155 $Y=1.34
+ $X2=3.155 $Y2=1.845
r35 13 14 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=3.07 $Y=1.295
+ $X2=3.07 $Y2=1.665
r36 13 18 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.07
+ $Y=1.34 $X2=3.07 $Y2=1.34
r37 9 18 32.933 $w=2.55e-07 $l=2.49199e-07 $layer=POLY_cond $X=3.335 $Y=1.175
+ $X2=3.155 $Y2=1.34
r38 9 11 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=3.335 $Y=1.175
+ $X2=3.335 $Y2=0.495
r39 7 20 173.918 $w=2.5e-07 $l=7e-07 $layer=POLY_cond $X=3.285 $Y=2.545
+ $X2=3.285 $Y2=1.845
r40 1 18 32.933 $w=2.55e-07 $l=2.49199e-07 $layer=POLY_cond $X=2.975 $Y=1.175
+ $X2=3.155 $Y2=1.34
r41 1 3 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=2.975 $Y=1.175
+ $X2=2.975 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__NOR3B_LP%VPWR 1 2 9 15 20 21 23 24 25 38 39
r33 38 39 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r34 36 39 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r35 35 36 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r36 32 35 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=0.72 $Y=3.33
+ $X2=2.64 $Y2=3.33
r37 32 33 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r38 29 33 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r39 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r40 25 36 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=2.64 $Y2=3.33
r41 25 33 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=0.72 $Y2=3.33
r42 23 35 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=2.855 $Y=3.33
+ $X2=2.64 $Y2=3.33
r43 23 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.855 $Y=3.33
+ $X2=3.02 $Y2=3.33
r44 22 38 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=3.185 $Y=3.33
+ $X2=3.6 $Y2=3.33
r45 22 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.185 $Y=3.33
+ $X2=3.02 $Y2=3.33
r46 20 28 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=0.385 $Y=3.33
+ $X2=0.24 $Y2=3.33
r47 20 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.385 $Y=3.33
+ $X2=0.55 $Y2=3.33
r48 19 32 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=0.715 $Y=3.33
+ $X2=0.72 $Y2=3.33
r49 19 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.715 $Y=3.33
+ $X2=0.55 $Y2=3.33
r50 15 18 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=3.02 $Y=2.19 $X2=3.02
+ $Y2=2.9
r51 13 24 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.02 $Y=3.245
+ $X2=3.02 $Y2=3.33
r52 13 18 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=3.02 $Y=3.245
+ $X2=3.02 $Y2=2.9
r53 9 12 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=0.55 $Y=2.19 $X2=0.55
+ $Y2=2.9
r54 7 21 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.55 $Y=3.245 $X2=0.55
+ $Y2=3.33
r55 7 12 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=0.55 $Y=3.245
+ $X2=0.55 $Y2=2.9
r56 2 18 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=2.875
+ $Y=2.045 $X2=3.02 $Y2=2.9
r57 2 15 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=2.875
+ $Y=2.045 $X2=3.02 $Y2=2.19
r58 1 12 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.405
+ $Y=2.045 $X2=0.55 $Y2=2.9
r59 1 9 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.405
+ $Y=2.045 $X2=0.55 $Y2=2.19
.ends

.subckt PM_SKY130_FD_SC_LP__NOR3B_LP%Y 1 2 3 10 14 20 22 24 25 26
r58 26 35 6.74611 $w=6.42e-07 $l=3.55e-07 $layer=LI1_cond $X=0.48 $Y=0.555
+ $X2=0.48 $Y2=0.91
r59 26 31 1.14019 $w=6.42e-07 $l=6e-08 $layer=LI1_cond $X=0.48 $Y=0.555 $X2=0.48
+ $Y2=0.495
r60 20 25 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=2.14 $Y=2.19
+ $X2=2.14 $Y2=2.025
r61 20 22 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=2.14 $Y=2.19 $X2=2.14
+ $Y2=2.9
r62 16 24 3.64284 $w=2.55e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.06 $Y=0.995
+ $X2=1.975 $Y2=0.91
r63 16 25 67.1979 $w=1.68e-07 $l=1.03e-06 $layer=LI1_cond $X=2.06 $Y=0.995
+ $X2=2.06 $Y2=2.025
r64 12 24 3.64284 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=1.975 $Y=0.825
+ $X2=1.975 $Y2=0.91
r65 12 14 11.1855 $w=3.38e-07 $l=3.3e-07 $layer=LI1_cond $X=1.975 $Y=0.825
+ $X2=1.975 $Y2=0.495
r66 11 35 8.75512 $w=1.7e-07 $l=3.55e-07 $layer=LI1_cond $X=0.835 $Y=0.91
+ $X2=0.48 $Y2=0.91
r67 10 24 2.83584 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=1.805 $Y=0.91
+ $X2=1.975 $Y2=0.91
r68 10 11 63.2834 $w=1.68e-07 $l=9.7e-07 $layer=LI1_cond $X=1.805 $Y=0.91
+ $X2=0.835 $Y2=0.91
r69 3 22 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=2
+ $Y=2.045 $X2=2.14 $Y2=2.9
r70 3 20 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2
+ $Y=2.045 $X2=2.14 $Y2=2.19
r71 2 14 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.83
+ $Y=0.285 $X2=1.97 $Y2=0.495
r72 1 31 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.245
+ $Y=0.285 $X2=0.39 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__NOR3B_LP%VGND 1 2 9 13 15 17 22 29 30 33 36
c50 17 0 7.83201e-20 $X=1.015 $Y=0
r51 36 37 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r52 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r53 30 37 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=2.64
+ $Y2=0
r54 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r55 27 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.925 $Y=0 $X2=2.76
+ $Y2=0
r56 27 29 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=2.925 $Y=0 $X2=3.6
+ $Y2=0
r57 26 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r58 25 26 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r59 23 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.345 $Y=0 $X2=1.18
+ $Y2=0
r60 23 25 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.345 $Y=0 $X2=1.68
+ $Y2=0
r61 22 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.595 $Y=0 $X2=2.76
+ $Y2=0
r62 22 25 59.6952 $w=1.68e-07 $l=9.15e-07 $layer=LI1_cond $X=2.595 $Y=0 $X2=1.68
+ $Y2=0
r63 20 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r64 19 20 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r65 17 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.015 $Y=0 $X2=1.18
+ $Y2=0
r66 17 19 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.015 $Y=0 $X2=0.72
+ $Y2=0
r67 15 37 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=2.64
+ $Y2=0
r68 15 26 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=1.68
+ $Y2=0
r69 11 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.76 $Y=0.085
+ $X2=2.76 $Y2=0
r70 11 13 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=2.76 $Y=0.085
+ $X2=2.76 $Y2=0.455
r71 7 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.18 $Y=0.085 $X2=1.18
+ $Y2=0
r72 7 9 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.18 $Y=0.085 $X2=1.18
+ $Y2=0.455
r73 2 13 182 $w=1.7e-07 $l=2.29565e-07 $layer=licon1_NDIFF $count=1 $X=2.62
+ $Y=0.285 $X2=2.76 $Y2=0.455
r74 1 9 182 $w=1.7e-07 $l=2.29565e-07 $layer=licon1_NDIFF $count=1 $X=1.04
+ $Y=0.285 $X2=1.18 $Y2=0.455
.ends

