* File: sky130_fd_sc_lp__srdlstp_1.spice
* Created: Fri Aug 28 11:33:10 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__srdlstp_1.pex.spice"
.subckt sky130_fd_sc_lp__srdlstp_1  VNB VPB D SET_B GATE SLEEP_B VPWR KAPWR Q
+ VGND
* 
* VGND	VGND
* Q	Q
* KAPWR	KAPWR
* VPWR	VPWR
* SLEEP_B	SLEEP_B
* GATE	GATE
* SET_B	SET_B
* D	D
* VPB	VPB
* VNB	VNB
MM1024 N_A_27_400#_M1024_d N_D_M1024_g N_VGND_M1024_s VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.1113 PD=1.37 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1031 A_300_130# N_A_27_400#_M1031_g N_A_217_130#_M1031_s VNB NSHORT L=0.15
+ W=0.64 AD=0.0672 AS=0.1696 PD=0.85 PS=1.81 NRD=9.372 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75000.9 A=0.096 P=1.58 MULT=1
MM1025 N_VGND_M1025_d N_SET_B_M1025_g A_300_130# VNB NSHORT L=0.15 W=0.64
+ AD=0.130294 AS=0.0672 PD=1.22566 PS=0.85 NRD=0 NRS=9.372 M=1 R=4.26667
+ SA=75000.6 SB=75000.5 A=0.096 P=1.58 MULT=1
MM1034 N_A_434_405#_M1034_d N_A_404_353#_M1034_g N_VGND_M1025_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.1113 AS=0.0855057 PD=1.37 PS=0.80434 NRD=0 NRS=27.132 M=1
+ R=2.8 SA=75001.1 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1019 A_667_47# N_A_434_405#_M1019_g N_A_217_130#_M1019_s VNB NSHORT L=0.15
+ W=0.64 AD=0.0672 AS=0.1696 PD=0.85 PS=1.81 NRD=9.372 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75001.4 A=0.096 P=1.58 MULT=1
MM1021 N_A_700_451#_M1021_d N_A_434_405#_M1021_g A_667_47# VNB NSHORT L=0.15
+ W=0.64 AD=0.130294 AS=0.0672 PD=1.22566 PS=0.85 NRD=0 NRS=9.372 M=1 R=4.26667
+ SA=75000.6 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1029 A_844_47# N_A_404_353#_M1029_g N_A_700_451#_M1021_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.0855057 PD=0.63 PS=0.80434 NRD=14.28 NRS=28.56 M=1 R=2.8
+ SA=75001.1 SB=75001 A=0.063 P=1.14 MULT=1
MM1012 A_916_47# N_A_878_357#_M1012_g A_844_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0441 PD=0.63 PS=0.63 NRD=14.28 NRS=14.28 M=1 R=2.8 SA=75001.4
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1016 N_A_988_47#_M1016_d N_A_878_357#_M1016_g A_916_47# VNB NSHORT L=0.15
+ W=0.42 AD=0.23045 AS=0.0441 PD=2.11 PS=0.63 NRD=141.048 NRS=14.28 M=1 R=2.8
+ SA=75001.8 SB=75000.3 A=0.063 P=1.14 MULT=1
MM1011 N_A_988_47#_M1011_d N_SET_B_M1011_g N_VGND_M1011_s VNB NSHORT L=0.15
+ W=0.42 AD=0.08085 AS=0.1155 PD=0.805 PS=1.39 NRD=30 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.8 A=0.063 P=1.14 MULT=1
MM1020 N_VGND_M1020_d N_A_1294_315#_M1020_g N_A_988_47#_M1011_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.0588 AS=0.08085 PD=0.7 PS=0.805 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.7 SB=75001.3 A=0.063 P=1.14 MULT=1
MM1022 A_1455_127# N_A_700_451#_M1022_g N_VGND_M1020_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0756 AS=0.0588 PD=0.78 PS=0.7 NRD=35.712 NRS=0 M=1 R=2.8 SA=75001.2
+ SB=75000.8 A=0.063 P=1.14 MULT=1
MM1006 N_A_878_357#_M1006_d N_A_700_451#_M1006_g A_1455_127# VNB NSHORT L=0.15
+ W=0.42 AD=0.244275 AS=0.0756 PD=2.18 PS=0.78 NRD=34.284 NRS=35.712 M=1 R=2.8
+ SA=75001.7 SB=75000.3 A=0.063 P=1.14 MULT=1
MM1013 A_1798_174# N_GATE_M1013_g N_A_404_353#_M1013_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.1638 PD=0.66 PS=1.62 NRD=18.564 NRS=31.428 M=1 R=2.8 SA=75000.3
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1004 A_1876_174# N_SLEEP_B_M1004_g A_1798_174# VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0504 PD=0.63 PS=0.66 NRD=14.28 NRS=18.564 M=1 R=2.8 SA=75000.7
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1032 N_VGND_M1032_d N_SLEEP_B_M1032_g A_1876_174# VNB NSHORT L=0.15 W=0.42
+ AD=0.1176 AS=0.0441 PD=1.4 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.1
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1023 A_2144_131# N_SLEEP_B_M1023_g N_A_1294_315#_M1023_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.1176 PD=0.63 PS=1.4 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1015 N_VGND_M1015_d N_SLEEP_B_M1015_g A_2144_131# VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1017 N_A_2266_367#_M1017_d N_A_700_451#_M1017_g N_VGND_M1015_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.1176 AS=0.0588 PD=1.4 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1008 N_Q_M1008_d N_A_2266_367#_M1008_g N_VGND_M1008_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2352 AS=0.2352 PD=2.24 PS=2.24 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1028 N_VPWR_M1028_d N_D_M1028_g N_A_27_400#_M1028_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.130335 AS=0.176 PD=1.05946 PS=1.83 NRD=33.8446 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75000.7 A=0.096 P=1.58 MULT=1
MM1005 N_A_217_130#_M1005_d N_A_27_400#_M1005_g N_VPWR_M1028_d VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.231 AS=0.171065 PD=2.23 PS=1.39054 NRD=0 NRS=0 M=1 R=5.6
+ SA=75000.6 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1010 N_A_434_405#_M1010_d N_A_404_353#_M1010_g N_VPWR_M1010_s VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.176 AS=0.3755 PD=1.83 PS=3.02 NRD=0 NRS=163.668 M=1
+ R=4.26667 SA=75000.3 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1033 A_628_451# N_A_404_353#_M1033_g N_A_217_130#_M1033_s VPB PHIGHVT L=0.15
+ W=0.84 AD=0.0882 AS=0.231 PD=1.05 PS=2.23 NRD=11.7215 NRS=0 M=1 R=5.6
+ SA=75000.2 SB=75001.7 A=0.126 P=1.98 MULT=1
MM1030 N_A_700_451#_M1030_d N_A_404_353#_M1030_g A_628_451# VPB PHIGHVT L=0.15
+ W=0.84 AD=0.174574 AS=0.0882 PD=1.27826 PS=1.05 NRD=26.9693 NRS=11.7215 M=1
+ R=5.6 SA=75000.6 SB=75001.3 A=0.126 P=1.98 MULT=1
MM1014 A_830_419# N_A_434_405#_M1014_g N_A_700_451#_M1030_d VPB PHIGHVT L=0.25
+ W=1 AD=0.12 AS=0.207826 PD=1.24 PS=1.52174 NRD=12.7853 NRS=0.9653 M=1 R=4
+ SA=125001 SB=125001 A=0.25 P=2.5 MULT=1
MM1000 N_KAPWR_M1000_d N_A_878_357#_M1000_g A_830_419# VPB PHIGHVT L=0.25 W=1
+ AD=0.28 AS=0.12 PD=2.56 PS=1.24 NRD=0 NRS=12.7853 M=1 R=4 SA=125001 SB=125000
+ A=0.25 P=2.5 MULT=1
MM1026 A_1246_341# N_SET_B_M1026_g N_A_700_451#_M1026_s VPB PHIGHVT L=0.25 W=1
+ AD=0.12 AS=0.4377 PD=1.24 PS=3.06 NRD=12.7853 NRS=23.6203 M=1 R=4 SA=125000
+ SB=125001 A=0.25 P=2.5 MULT=1
MM1002 N_KAPWR_M1002_d N_A_1294_315#_M1002_g A_1246_341# VPB PHIGHVT L=0.25 W=1
+ AD=0.2752 AS=0.12 PD=1.735 PS=1.24 NRD=43.3597 NRS=12.7853 M=1 R=4 SA=125001
+ SB=125001 A=0.25 P=2.5 MULT=1
MM1009 N_A_878_357#_M1009_d N_A_700_451#_M1009_g N_KAPWR_M1002_d VPB PHIGHVT
+ L=0.25 W=1 AD=0.285 AS=0.2752 PD=2.57 PS=1.735 NRD=0 NRS=43.3597 M=1 R=4
+ SA=125001 SB=125000 A=0.25 P=2.5 MULT=1
MM1007 N_A_404_353#_M1007_d N_GATE_M1007_g N_KAPWR_M1007_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1607 AS=0.1824 PD=1.525 PS=1.85 NRD=60.3411 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75000.5 A=0.096 P=1.58 MULT=1
MM1003 N_KAPWR_M1003_d N_SLEEP_B_M1003_g N_A_404_353#_M1007_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.198283 AS=0.1607 PD=1.28 PS=1.525 NRD=78.4257 NRS=0 M=1 R=4.26667
+ SA=75000.3 SB=75001 A=0.096 P=1.58 MULT=1
MM1001 N_A_1294_315#_M1001_d N_SLEEP_B_M1001_g N_KAPWR_M1003_d VPB PHIGHVT
+ L=0.25 W=1 AD=0.285 AS=0.309817 PD=2.57 PS=2 NRD=0 NRS=23.6203 M=1 R=4
+ SA=125001 SB=125000 A=0.25 P=2.5 MULT=1
MM1027 N_VPWR_M1027_d N_A_700_451#_M1027_g N_A_2266_367#_M1027_s VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.20672 AS=0.1824 PD=1.26316 PS=1.85 NRD=82.3263 NRS=0 M=1
+ R=4.26667 SA=75000.2 SB=75001 A=0.096 P=1.58 MULT=1
MM1018 N_Q_M1018_d N_A_2266_367#_M1018_g N_VPWR_M1027_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3591 AS=0.40698 PD=3.09 PS=2.48684 NRD=0 NRS=10.9335 M=1 R=8.4
+ SA=75000.6 SB=75000.2 A=0.189 P=2.82 MULT=1
DX35_noxref VNB VPB NWDIODE A=25.5811 P=30.93
c_142 VNB 0 1.06489e-19 $X=0 $Y=0
c_230 VPB 0 1.01441e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_lp__srdlstp_1.pxi.spice"
*
.ends
*
*
