* File: sky130_fd_sc_lp__o21bai_m.pxi.spice
* Created: Fri Aug 28 11:07:08 2020
* 
x_PM_SKY130_FD_SC_LP__O21BAI_M%B1_N N_B1_N_M1002_g N_B1_N_M1005_g N_B1_N_c_64_n
+ N_B1_N_c_65_n N_B1_N_c_66_n B1_N B1_N N_B1_N_c_68_n
+ PM_SKY130_FD_SC_LP__O21BAI_M%B1_N
x_PM_SKY130_FD_SC_LP__O21BAI_M%A_32_62# N_A_32_62#_M1002_s N_A_32_62#_M1005_s
+ N_A_32_62#_M1007_g N_A_32_62#_c_99_n N_A_32_62#_c_100_n N_A_32_62#_c_101_n
+ N_A_32_62#_M1001_g N_A_32_62#_c_102_n N_A_32_62#_c_107_n N_A_32_62#_c_108_n
+ N_A_32_62#_c_103_n N_A_32_62#_c_110_n N_A_32_62#_c_111_n N_A_32_62#_c_104_n
+ N_A_32_62#_c_112_n N_A_32_62#_c_113_n N_A_32_62#_c_114_n
+ PM_SKY130_FD_SC_LP__O21BAI_M%A_32_62#
x_PM_SKY130_FD_SC_LP__O21BAI_M%A2 N_A2_M1003_g N_A2_M1006_g A2 A2 A2
+ N_A2_c_160_n PM_SKY130_FD_SC_LP__O21BAI_M%A2
x_PM_SKY130_FD_SC_LP__O21BAI_M%A1 N_A1_M1004_g N_A1_c_196_n N_A1_c_197_n
+ N_A1_M1000_g N_A1_c_198_n A1 A1 A1 A1 N_A1_c_194_n
+ PM_SKY130_FD_SC_LP__O21BAI_M%A1
x_PM_SKY130_FD_SC_LP__O21BAI_M%VPWR N_VPWR_M1005_d N_VPWR_M1004_d N_VPWR_c_224_n
+ N_VPWR_c_225_n N_VPWR_c_226_n N_VPWR_c_227_n VPWR N_VPWR_c_228_n
+ N_VPWR_c_223_n N_VPWR_c_230_n PM_SKY130_FD_SC_LP__O21BAI_M%VPWR
x_PM_SKY130_FD_SC_LP__O21BAI_M%Y N_Y_M1001_s N_Y_M1007_d N_Y_c_253_n N_Y_c_254_n
+ Y Y PM_SKY130_FD_SC_LP__O21BAI_M%Y
x_PM_SKY130_FD_SC_LP__O21BAI_M%VGND N_VGND_M1002_d N_VGND_M1006_d N_VGND_c_286_n
+ N_VGND_c_287_n VGND N_VGND_c_288_n N_VGND_c_289_n N_VGND_c_290_n
+ N_VGND_c_291_n N_VGND_c_292_n N_VGND_c_293_n PM_SKY130_FD_SC_LP__O21BAI_M%VGND
x_PM_SKY130_FD_SC_LP__O21BAI_M%A_320_78# N_A_320_78#_M1001_d N_A_320_78#_M1000_d
+ N_A_320_78#_c_320_n N_A_320_78#_c_321_n N_A_320_78#_c_322_n
+ N_A_320_78#_c_323_n PM_SKY130_FD_SC_LP__O21BAI_M%A_320_78#
cc_1 VNB N_B1_N_M1005_g 0.00876313f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=2.885
cc_2 VNB N_B1_N_c_64_n 0.0234519f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=0.84
cc_3 VNB N_B1_N_c_65_n 0.0236725f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.345
cc_4 VNB N_B1_N_c_66_n 0.016658f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.51
cc_5 VNB B1_N 0.0106861f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.84
cc_6 VNB N_B1_N_c_68_n 0.0176617f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.005
cc_7 VNB N_A_32_62#_c_99_n 0.0335062f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_8 VNB N_A_32_62#_c_100_n 0.0133967f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_32_62#_c_101_n 0.019221f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_32_62#_c_102_n 0.0319415f $X=-0.19 $Y=-0.245 $X2=0.655 $Y2=0.925
cc_11 VNB N_A_32_62#_c_103_n 0.0461855f $X=-0.19 $Y=-0.245 $X2=0.655 $Y2=1.295
cc_12 VNB N_A_32_62#_c_104_n 0.0120122f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A2_M1006_g 0.0374171f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB A2 0.00447387f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=0.84
cc_15 VNB N_A2_c_160_n 0.0468191f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.005
cc_16 VNB N_A1_M1000_g 0.0651909f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=0.84
cc_17 VNB A1 0.0203058f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A1_c_194_n 0.011792f $X=-0.19 $Y=-0.245 $X2=0.655 $Y2=1.295
cc_19 VNB N_VPWR_c_223_n 0.123877f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_Y_c_253_n 0.0134221f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.005
cc_21 VNB N_Y_c_254_n 8.02662e-19 $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.345
cc_22 VNB N_VGND_c_286_n 0.00766036f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=0.84
cc_23 VNB N_VGND_c_287_n 0.00986829f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_24 VNB N_VGND_c_288_n 0.0196212f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.005
cc_25 VNB N_VGND_c_289_n 0.037182f $X=-0.19 $Y=-0.245 $X2=0.655 $Y2=1.005
cc_26 VNB N_VGND_c_290_n 0.0201858f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_291_n 0.211025f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_292_n 0.00401418f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_293_n 0.0040393f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_320_78#_c_320_n 8.22023e-19 $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=0.84
cc_31 VNB N_A_320_78#_c_321_n 0.0235686f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=1.51
cc_32 VNB N_A_320_78#_c_322_n 0.00329621f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.84
cc_33 VNB N_A_320_78#_c_323_n 0.00224906f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VPB N_B1_N_M1005_g 0.0765443f $X=-0.19 $Y=1.655 $X2=0.53 $Y2=2.885
cc_35 VPB N_A_32_62#_M1007_g 0.0259526f $X=-0.19 $Y=1.655 $X2=0.59 $Y2=1.51
cc_36 VPB N_A_32_62#_c_102_n 0.00543532f $X=-0.19 $Y=1.655 $X2=0.655 $Y2=0.925
cc_37 VPB N_A_32_62#_c_107_n 0.0239201f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_38 VPB N_A_32_62#_c_108_n 0.0170574f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_39 VPB N_A_32_62#_c_103_n 0.00454308f $X=-0.19 $Y=1.655 $X2=0.655 $Y2=1.295
cc_40 VPB N_A_32_62#_c_110_n 0.0416034f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_41 VPB N_A_32_62#_c_111_n 0.0091426f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_42 VPB N_A_32_62#_c_112_n 0.0123457f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_43 VPB N_A_32_62#_c_113_n 0.00554676f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_44 VPB N_A_32_62#_c_114_n 0.017872f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_45 VPB N_A2_M1003_g 0.0453611f $X=-0.19 $Y=1.655 $X2=0.5 $Y2=0.52
cc_46 VPB A2 0.00417338f $X=-0.19 $Y=1.655 $X2=0.59 $Y2=0.84
cc_47 VPB N_A2_c_160_n 0.0447445f $X=-0.19 $Y=1.655 $X2=0.59 $Y2=1.005
cc_48 VPB N_A1_M1004_g 0.0346884f $X=-0.19 $Y=1.655 $X2=0.5 $Y2=0.52
cc_49 VPB N_A1_c_196_n 0.0552156f $X=-0.19 $Y=1.655 $X2=0.53 $Y2=2.885
cc_50 VPB N_A1_c_197_n 0.00769697f $X=-0.19 $Y=1.655 $X2=0.53 $Y2=2.885
cc_51 VPB N_A1_c_198_n 0.0445567f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_52 VPB A1 0.039369f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_53 VPB N_A1_c_194_n 0.00707094f $X=-0.19 $Y=1.655 $X2=0.655 $Y2=1.295
cc_54 VPB N_VPWR_c_224_n 0.00561589f $X=-0.19 $Y=1.655 $X2=0.59 $Y2=1.51
cc_55 VPB N_VPWR_c_225_n 0.00495479f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_56 VPB N_VPWR_c_226_n 0.0269971f $X=-0.19 $Y=1.655 $X2=0.59 $Y2=1.005
cc_57 VPB N_VPWR_c_227_n 0.00401108f $X=-0.19 $Y=1.655 $X2=0.655 $Y2=0.925
cc_58 VPB N_VPWR_c_228_n 0.0244187f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_59 VPB N_VPWR_c_223_n 0.0607894f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_60 VPB N_VPWR_c_230_n 0.0271613f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_61 VPB N_Y_c_253_n 0.0117824f $X=-0.19 $Y=1.655 $X2=0.59 $Y2=1.005
cc_62 VPB Y 0.0111339f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_63 N_B1_N_M1005_g N_A_32_62#_M1007_g 0.0178952f $X=0.53 $Y=2.885 $X2=0 $Y2=0
cc_64 B1_N N_A_32_62#_c_100_n 0.00509978f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_65 N_B1_N_c_68_n N_A_32_62#_c_100_n 0.0151144f $X=0.59 $Y=1.005 $X2=0 $Y2=0
cc_66 N_B1_N_c_68_n N_A_32_62#_c_101_n 7.1714e-19 $X=0.59 $Y=1.005 $X2=0 $Y2=0
cc_67 N_B1_N_M1005_g N_A_32_62#_c_102_n 0.00702148f $X=0.53 $Y=2.885 $X2=0 $Y2=0
cc_68 N_B1_N_c_65_n N_A_32_62#_c_102_n 0.0151144f $X=0.59 $Y=1.345 $X2=0 $Y2=0
cc_69 N_B1_N_M1005_g N_A_32_62#_c_103_n 0.00849887f $X=0.53 $Y=2.885 $X2=0 $Y2=0
cc_70 N_B1_N_c_64_n N_A_32_62#_c_103_n 0.0223447f $X=0.59 $Y=0.84 $X2=0 $Y2=0
cc_71 B1_N N_A_32_62#_c_103_n 0.0468337f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_72 N_B1_N_M1005_g N_A_32_62#_c_110_n 0.0324563f $X=0.53 $Y=2.885 $X2=0 $Y2=0
cc_73 N_B1_N_M1005_g N_A_32_62#_c_111_n 0.0116809f $X=0.53 $Y=2.885 $X2=0 $Y2=0
cc_74 N_B1_N_c_66_n N_A_32_62#_c_111_n 9.72924e-19 $X=0.59 $Y=1.51 $X2=0 $Y2=0
cc_75 B1_N N_A_32_62#_c_111_n 0.0181851f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_76 N_B1_N_M1005_g N_A_32_62#_c_112_n 0.00513266f $X=0.53 $Y=2.885 $X2=0 $Y2=0
cc_77 N_B1_N_c_66_n N_A_32_62#_c_112_n 0.00134641f $X=0.59 $Y=1.51 $X2=0 $Y2=0
cc_78 N_B1_N_M1005_g N_A_32_62#_c_113_n 0.00146872f $X=0.53 $Y=2.885 $X2=0 $Y2=0
cc_79 N_B1_N_M1005_g N_A_32_62#_c_114_n 0.0407954f $X=0.53 $Y=2.885 $X2=0 $Y2=0
cc_80 N_B1_N_M1005_g N_VPWR_c_224_n 0.00445728f $X=0.53 $Y=2.885 $X2=0 $Y2=0
cc_81 N_B1_N_M1005_g N_VPWR_c_223_n 0.0113354f $X=0.53 $Y=2.885 $X2=0 $Y2=0
cc_82 N_B1_N_M1005_g N_VPWR_c_230_n 0.00553654f $X=0.53 $Y=2.885 $X2=0 $Y2=0
cc_83 B1_N N_Y_c_253_n 0.0266373f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_84 N_B1_N_c_68_n N_Y_c_253_n 4.22453e-19 $X=0.59 $Y=1.005 $X2=0 $Y2=0
cc_85 N_B1_N_c_64_n N_Y_c_254_n 0.00452173f $X=0.59 $Y=0.84 $X2=0 $Y2=0
cc_86 N_B1_N_c_64_n N_VGND_c_286_n 0.00488761f $X=0.59 $Y=0.84 $X2=0 $Y2=0
cc_87 B1_N N_VGND_c_286_n 0.0126177f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_88 N_B1_N_c_68_n N_VGND_c_286_n 0.00101807f $X=0.59 $Y=1.005 $X2=0 $Y2=0
cc_89 N_B1_N_c_64_n N_VGND_c_288_n 0.00512921f $X=0.59 $Y=0.84 $X2=0 $Y2=0
cc_90 N_B1_N_c_64_n N_VGND_c_291_n 0.00905395f $X=0.59 $Y=0.84 $X2=0 $Y2=0
cc_91 B1_N N_VGND_c_291_n 0.00419633f $X=0.635 $Y=0.84 $X2=0 $Y2=0
cc_92 N_A_32_62#_c_107_n N_A2_M1003_g 0.0316808f $X=0.98 $Y=2.255 $X2=0 $Y2=0
cc_93 N_A_32_62#_c_101_n N_A2_M1006_g 0.0216683f $X=1.525 $Y=0.92 $X2=0 $Y2=0
cc_94 N_A_32_62#_c_99_n N_A2_c_160_n 0.0126877f $X=1.45 $Y=0.995 $X2=0 $Y2=0
cc_95 N_A_32_62#_c_102_n N_A2_c_160_n 0.0316808f $X=0.98 $Y=1.75 $X2=0 $Y2=0
cc_96 N_A_32_62#_M1007_g N_VPWR_c_224_n 0.0033813f $X=1.07 $Y=2.885 $X2=0 $Y2=0
cc_97 N_A_32_62#_c_108_n N_VPWR_c_224_n 0.00330369f $X=0.98 $Y=2.42 $X2=0 $Y2=0
cc_98 N_A_32_62#_c_113_n N_VPWR_c_224_n 0.00279683f $X=0.98 $Y=1.915 $X2=0 $Y2=0
cc_99 N_A_32_62#_M1007_g N_VPWR_c_226_n 0.00585385f $X=1.07 $Y=2.885 $X2=0 $Y2=0
cc_100 N_A_32_62#_M1005_s N_VPWR_c_223_n 0.00235821f $X=0.19 $Y=2.675 $X2=0
+ $Y2=0
cc_101 N_A_32_62#_M1007_g N_VPWR_c_223_n 0.0109113f $X=1.07 $Y=2.885 $X2=0 $Y2=0
cc_102 N_A_32_62#_c_110_n N_VPWR_c_223_n 0.0115728f $X=0.315 $Y=2.82 $X2=0 $Y2=0
cc_103 N_A_32_62#_c_110_n N_VPWR_c_230_n 0.010662f $X=0.315 $Y=2.82 $X2=0 $Y2=0
cc_104 N_A_32_62#_c_99_n N_Y_c_253_n 0.0143311f $X=1.45 $Y=0.995 $X2=0 $Y2=0
cc_105 N_A_32_62#_c_102_n N_Y_c_253_n 0.0172208f $X=0.98 $Y=1.75 $X2=0 $Y2=0
cc_106 N_A_32_62#_c_113_n N_Y_c_253_n 0.0402692f $X=0.98 $Y=1.915 $X2=0 $Y2=0
cc_107 N_A_32_62#_c_99_n N_Y_c_254_n 0.00158117f $X=1.45 $Y=0.995 $X2=0 $Y2=0
cc_108 N_A_32_62#_c_101_n N_Y_c_254_n 0.00170825f $X=1.525 $Y=0.92 $X2=0 $Y2=0
cc_109 N_A_32_62#_c_108_n Y 0.00782126f $X=0.98 $Y=2.42 $X2=0 $Y2=0
cc_110 N_A_32_62#_c_113_n Y 0.00755153f $X=0.98 $Y=1.915 $X2=0 $Y2=0
cc_111 N_A_32_62#_c_101_n N_VGND_c_286_n 0.00517595f $X=1.525 $Y=0.92 $X2=0
+ $Y2=0
cc_112 N_A_32_62#_c_104_n N_VGND_c_288_n 0.0106787f $X=0.285 $Y=0.495 $X2=0
+ $Y2=0
cc_113 N_A_32_62#_c_101_n N_VGND_c_289_n 0.00563421f $X=1.525 $Y=0.92 $X2=0
+ $Y2=0
cc_114 N_A_32_62#_c_101_n N_VGND_c_291_n 0.00539454f $X=1.525 $Y=0.92 $X2=0
+ $Y2=0
cc_115 N_A_32_62#_c_104_n N_VGND_c_291_n 0.00883735f $X=0.285 $Y=0.495 $X2=0
+ $Y2=0
cc_116 N_A_32_62#_c_101_n N_A_320_78#_c_320_n 4.03889e-19 $X=1.525 $Y=0.92 $X2=0
+ $Y2=0
cc_117 N_A_32_62#_c_101_n N_A_320_78#_c_322_n 0.00178997f $X=1.525 $Y=0.92 $X2=0
+ $Y2=0
cc_118 N_A2_M1003_g N_A1_c_197_n 0.0616377f $X=1.5 $Y=2.885 $X2=0 $Y2=0
cc_119 N_A2_c_160_n N_A1_c_197_n 0.0173313f $X=1.68 $Y=1.475 $X2=0 $Y2=0
cc_120 N_A2_M1006_g N_A1_M1000_g 0.0317436f $X=1.955 $Y=0.6 $X2=0 $Y2=0
cc_121 A2 N_A1_M1000_g 0.0017067f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_122 A2 N_A1_c_198_n 0.00241165f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_123 N_A2_M1006_g A1 0.00316396f $X=1.955 $Y=0.6 $X2=0 $Y2=0
cc_124 A2 A1 0.0228966f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_125 N_A2_c_160_n N_A1_c_194_n 0.0317436f $X=1.68 $Y=1.475 $X2=0 $Y2=0
cc_126 N_A2_M1003_g N_VPWR_c_226_n 0.00398598f $X=1.5 $Y=2.885 $X2=0 $Y2=0
cc_127 N_A2_M1003_g N_VPWR_c_223_n 0.00551814f $X=1.5 $Y=2.885 $X2=0 $Y2=0
cc_128 N_A2_M1006_g N_Y_c_253_n 0.00390296f $X=1.955 $Y=0.6 $X2=0 $Y2=0
cc_129 A2 N_Y_c_253_n 0.0632484f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_130 N_A2_c_160_n N_Y_c_253_n 0.0125494f $X=1.68 $Y=1.475 $X2=0 $Y2=0
cc_131 N_A2_M1003_g Y 0.0241788f $X=1.5 $Y=2.885 $X2=0 $Y2=0
cc_132 A2 Y 0.0137852f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_133 N_A2_c_160_n Y 0.00172823f $X=1.68 $Y=1.475 $X2=0 $Y2=0
cc_134 N_A2_M1006_g N_VGND_c_287_n 0.00329204f $X=1.955 $Y=0.6 $X2=0 $Y2=0
cc_135 N_A2_M1006_g N_VGND_c_289_n 0.00563421f $X=1.955 $Y=0.6 $X2=0 $Y2=0
cc_136 N_A2_M1006_g N_VGND_c_291_n 0.00539454f $X=1.955 $Y=0.6 $X2=0 $Y2=0
cc_137 N_A2_M1006_g N_A_320_78#_c_320_n 6.71115e-19 $X=1.955 $Y=0.6 $X2=0 $Y2=0
cc_138 N_A2_M1006_g N_A_320_78#_c_321_n 0.0160784f $X=1.955 $Y=0.6 $X2=0 $Y2=0
cc_139 N_A2_c_160_n N_A_320_78#_c_321_n 0.00126371f $X=1.68 $Y=1.475 $X2=0 $Y2=0
cc_140 A2 N_A_320_78#_c_322_n 0.011359f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_141 N_A2_c_160_n N_A_320_78#_c_322_n 0.00408552f $X=1.68 $Y=1.475 $X2=0 $Y2=0
cc_142 N_A1_M1004_g N_VPWR_c_225_n 0.00460896f $X=1.86 $Y=2.885 $X2=0 $Y2=0
cc_143 N_A1_c_196_n N_VPWR_c_225_n 0.00595338f $X=2.31 $Y=2.295 $X2=0 $Y2=0
cc_144 N_A1_M1004_g N_VPWR_c_226_n 0.00585385f $X=1.86 $Y=2.885 $X2=0 $Y2=0
cc_145 N_A1_M1004_g N_VPWR_c_223_n 0.0118303f $X=1.86 $Y=2.885 $X2=0 $Y2=0
cc_146 A1 N_VPWR_c_223_n 0.0131302f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_147 N_A1_c_197_n Y 0.00881454f $X=1.935 $Y=2.295 $X2=0 $Y2=0
cc_148 A1 Y 0.00566818f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_149 N_A1_M1000_g N_VGND_c_287_n 0.00329204f $X=2.385 $Y=0.6 $X2=0 $Y2=0
cc_150 N_A1_M1000_g N_VGND_c_290_n 0.00563421f $X=2.385 $Y=0.6 $X2=0 $Y2=0
cc_151 N_A1_M1000_g N_VGND_c_291_n 0.00539454f $X=2.385 $Y=0.6 $X2=0 $Y2=0
cc_152 N_A1_M1000_g N_A_320_78#_c_321_n 0.0156361f $X=2.385 $Y=0.6 $X2=0 $Y2=0
cc_153 A1 N_A_320_78#_c_321_n 0.0263675f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_154 N_A1_c_194_n N_A_320_78#_c_321_n 6.30257e-19 $X=2.475 $Y=1.74 $X2=0 $Y2=0
cc_155 N_A1_M1000_g N_A_320_78#_c_323_n 0.00143084f $X=2.385 $Y=0.6 $X2=0 $Y2=0
cc_156 N_VPWR_c_223_n N_Y_M1007_d 0.00353471f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_157 N_VPWR_c_226_n Y 0.0178384f $X=1.97 $Y=3.33 $X2=0 $Y2=0
cc_158 N_VPWR_c_223_n Y 0.0198105f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_159 N_VPWR_c_223_n A_315_535# 0.00265196f $X=2.64 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_160 Y A_315_535# 0.00138834f $X=1.595 $Y=2.69 $X2=-0.19 $Y2=-0.245
cc_161 N_Y_c_254_n N_VGND_c_286_n 0.00493081f $X=1.31 $Y=0.665 $X2=0 $Y2=0
cc_162 N_Y_c_254_n N_VGND_c_289_n 0.00522733f $X=1.31 $Y=0.665 $X2=0 $Y2=0
cc_163 N_Y_c_254_n N_VGND_c_291_n 0.00692154f $X=1.31 $Y=0.665 $X2=0 $Y2=0
cc_164 N_Y_c_254_n N_A_320_78#_c_320_n 0.00308263f $X=1.31 $Y=0.665 $X2=0 $Y2=0
cc_165 N_Y_c_253_n N_A_320_78#_c_322_n 0.0115411f $X=1.33 $Y=2.32 $X2=0 $Y2=0
cc_166 N_VGND_c_289_n N_A_320_78#_c_320_n 0.00467386f $X=2.065 $Y=0 $X2=0 $Y2=0
cc_167 N_VGND_c_291_n N_A_320_78#_c_320_n 0.00677835f $X=2.64 $Y=0 $X2=0 $Y2=0
cc_168 N_VGND_c_287_n N_A_320_78#_c_321_n 0.0142847f $X=2.17 $Y=0.515 $X2=0
+ $Y2=0
cc_169 N_VGND_c_291_n N_A_320_78#_c_321_n 0.0146356f $X=2.64 $Y=0 $X2=0 $Y2=0
cc_170 N_VGND_c_290_n N_A_320_78#_c_323_n 0.00519224f $X=2.64 $Y=0 $X2=0 $Y2=0
cc_171 N_VGND_c_291_n N_A_320_78#_c_323_n 0.00688714f $X=2.64 $Y=0 $X2=0 $Y2=0
