* File: sky130_fd_sc_lp__dlrtp_lp2.pex.spice
* Created: Wed Sep  2 09:47:37 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__DLRTP_LP2%D 1 3 6 8 10 15 18 19 22 23
c42 22 0 7.69048e-20 $X=0.605 $Y=1.36
c43 18 0 6.58912e-21 $X=0.595 $Y=1.865
r44 22 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.605
+ $Y=1.36 $X2=0.605 $Y2=1.36
r45 19 23 9.63 $w=3.63e-07 $l=3.05e-07 $layer=LI1_cond $X=0.622 $Y=1.665
+ $X2=0.622 $Y2=1.36
r46 17 22 54.4068 $w=3.5e-07 $l=3.3e-07 $layer=POLY_cond $X=0.595 $Y=1.69
+ $X2=0.595 $Y2=1.36
r47 17 18 33.6482 $w=3.5e-07 $l=1.75e-07 $layer=POLY_cond $X=0.595 $Y=1.69
+ $X2=0.595 $Y2=1.865
r48 14 22 17.3113 $w=3.5e-07 $l=1.05e-07 $layer=POLY_cond $X=0.595 $Y=1.255
+ $X2=0.595 $Y2=1.36
r49 14 15 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=0.595 $Y=1.18
+ $X2=0.885 $Y2=1.18
r50 11 14 51.2766 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=0.495 $Y=1.18
+ $X2=0.595 $Y2=1.18
r51 8 15 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.885 $Y=1.105
+ $X2=0.885 $Y2=1.18
r52 8 10 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.885 $Y=1.105
+ $X2=0.885 $Y2=0.82
r53 6 18 181.371 $w=2.5e-07 $l=7.3e-07 $layer=POLY_cond $X=0.545 $Y=2.595
+ $X2=0.545 $Y2=1.865
r54 1 11 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.495 $Y=1.105
+ $X2=0.495 $Y2=1.18
r55 1 3 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.495 $Y=1.105
+ $X2=0.495 $Y2=0.82
.ends

.subckt PM_SKY130_FD_SC_LP__DLRTP_LP2%GATE 3 7 9 13 15 23
c47 13 0 1.53302e-19 $X=1.755 $Y=1.135
c48 9 0 8.75658e-20 $X=1.68 $Y=1.57
r49 22 23 30.474 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=1.395 $Y=1.66
+ $X2=1.47 $Y2=1.66
r50 21 22 41.9667 $w=3.3e-07 $l=2.4e-07 $layer=POLY_cond $X=1.155 $Y=1.66
+ $X2=1.395 $Y2=1.66
r51 18 21 1.74861 $w=3.3e-07 $l=1e-08 $layer=POLY_cond $X=1.145 $Y=1.66
+ $X2=1.155 $Y2=1.66
r52 15 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.145
+ $Y=1.66 $X2=1.145 $Y2=1.66
r53 11 13 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=1.755 $Y=1.495
+ $X2=1.755 $Y2=1.135
r54 9 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.68 $Y=1.57
+ $X2=1.755 $Y2=1.495
r55 9 23 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=1.68 $Y=1.57 $X2=1.47
+ $Y2=1.57
r56 5 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.395 $Y=1.495
+ $X2=1.395 $Y2=1.66
r57 5 7 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=1.395 $Y=1.495
+ $X2=1.395 $Y2=1.135
r58 1 21 9.34494 $w=2.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.155 $Y=1.825
+ $X2=1.155 $Y2=1.66
r59 1 3 173.918 $w=2.5e-07 $l=7e-07 $layer=POLY_cond $X=1.155 $Y=1.825 $X2=1.155
+ $Y2=2.525
.ends

.subckt PM_SKY130_FD_SC_LP__DLRTP_LP2%A_256_405# 1 2 7 9 14 16 17 19 21 22 24 27
+ 30 31 32 33 34 36 39 42 43 44 47 53 60 61 63 68
c150 68 0 3.54748e-20 $X=2.375 $Y=1.455
c151 63 0 1.22967e-19 $X=3.305 $Y=1.16
c152 61 0 7.69048e-20 $X=2.455 $Y=1.62
c153 60 0 6.60829e-20 $X=2.375 $Y=1.62
c154 53 0 4.59989e-21 $X=1.55 $Y=2.13
c155 42 0 3.46887e-19 $X=2.455 $Y=1.455
c156 36 0 6.58912e-21 $X=1.55 $Y=2.005
c157 34 0 1.03048e-19 $X=4.16 $Y=0.88
c158 33 0 1.07613e-19 $X=4.16 $Y=0.73
c159 31 0 1.97745e-19 $X=2.425 $Y=0.805
c160 27 0 1.08516e-19 $X=4.145 $Y=1.335
c161 22 0 7.00182e-20 $X=4.065 $Y=1.85
c162 17 0 1.06646e-19 $X=2.71 $Y=0.805
r163 60 69 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.375 $Y=1.62
+ $X2=2.375 $Y2=1.785
r164 60 68 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.375 $Y=1.62
+ $X2=2.375 $Y2=1.455
r165 59 61 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=2.375 $Y=1.62
+ $X2=2.455 $Y2=1.62
r166 59 60 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.375
+ $Y=1.62 $X2=2.375 $Y2=1.62
r167 57 59 14.1436 $w=3.28e-07 $l=4.05e-07 $layer=LI1_cond $X=1.97 $Y=1.62
+ $X2=2.375 $Y2=1.62
r168 55 57 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=1.55 $Y=1.62
+ $X2=1.97 $Y2=1.62
r169 51 53 5.9927 $w=2.48e-07 $l=1.3e-07 $layer=LI1_cond $X=1.42 $Y=2.13
+ $X2=1.55 $Y2=2.13
r170 47 48 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.005
+ $Y=1.5 $X2=4.005 $Y2=1.5
r171 45 63 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=3.305 $Y=1.5
+ $X2=3.305 $Y2=1.16
r172 45 47 21.4773 $w=3.28e-07 $l=6.15e-07 $layer=LI1_cond $X=3.39 $Y=1.5
+ $X2=4.005 $Y2=1.5
r173 43 63 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.22 $Y=1.16
+ $X2=3.305 $Y2=1.16
r174 43 44 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=3.22 $Y=1.16
+ $X2=2.54 $Y2=1.16
r175 42 61 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.455 $Y=1.455
+ $X2=2.455 $Y2=1.62
r176 41 44 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.455 $Y=1.245
+ $X2=2.54 $Y2=1.16
r177 41 42 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=2.455 $Y=1.245
+ $X2=2.455 $Y2=1.455
r178 37 57 0.716491 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=1.97 $Y=1.455
+ $X2=1.97 $Y2=1.62
r179 37 39 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=1.97 $Y=1.455
+ $X2=1.97 $Y2=1.09
r180 36 53 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.55 $Y=2.005
+ $X2=1.55 $Y2=2.13
r181 35 55 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.55 $Y=1.785
+ $X2=1.55 $Y2=1.62
r182 35 36 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=1.55 $Y=1.785
+ $X2=1.55 $Y2=2.005
r183 33 34 58.3064 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=4.16 $Y=0.73
+ $X2=4.16 $Y2=0.88
r184 32 69 92.2979 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=2.465 $Y=1.965
+ $X2=2.465 $Y2=1.785
r185 30 33 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=4.175 $Y=0.445
+ $X2=4.175 $Y2=0.73
r186 27 48 38.5334 $w=3.13e-07 $l=2.14942e-07 $layer=POLY_cond $X=4.145 $Y=1.335
+ $X2=4.03 $Y2=1.5
r187 27 34 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=4.145 $Y=1.335
+ $X2=4.145 $Y2=0.88
r188 22 48 55.9888 $w=3.13e-07 $l=3.67083e-07 $layer=POLY_cond $X=4.065 $Y=1.85
+ $X2=4.03 $Y2=1.5
r189 22 24 185.098 $w=2.5e-07 $l=7.45e-07 $layer=POLY_cond $X=4.065 $Y=1.85
+ $X2=4.065 $Y2=2.595
r190 19 21 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.785 $Y=0.73
+ $X2=2.785 $Y2=0.445
r191 18 31 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.5 $Y=0.805
+ $X2=2.425 $Y2=0.805
r192 17 19 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.71 $Y=0.805
+ $X2=2.785 $Y2=0.73
r193 17 18 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=2.71 $Y=0.805
+ $X2=2.5 $Y2=0.805
r194 14 32 40.9178 $w=2.5e-07 $l=1.25e-07 $layer=POLY_cond $X=2.515 $Y=2.09
+ $X2=2.515 $Y2=1.965
r195 14 16 97.364 $w=2.5e-07 $l=5.05e-07 $layer=POLY_cond $X=2.515 $Y=2.09
+ $X2=2.515 $Y2=2.595
r196 10 31 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.425 $Y=0.88
+ $X2=2.425 $Y2=0.805
r197 10 68 294.84 $w=1.5e-07 $l=5.75e-07 $layer=POLY_cond $X=2.425 $Y=0.88
+ $X2=2.425 $Y2=1.455
r198 7 31 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.425 $Y=0.73
+ $X2=2.425 $Y2=0.805
r199 7 9 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.425 $Y=0.73
+ $X2=2.425 $Y2=0.445
r200 2 51 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.28
+ $Y=2.025 $X2=1.42 $Y2=2.17
r201 1 39 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=1.83
+ $Y=0.925 $X2=1.97 $Y2=1.09
.ends

.subckt PM_SKY130_FD_SC_LP__DLRTP_LP2%A_27_122# 1 2 9 13 15 16 18 20 24 27 30 31
+ 32 35 39 43 44 45
c104 35 0 3.54748e-20 $X=2.915 $Y=1.59
c105 32 0 8.29659e-20 $X=1.985 $Y=2.05
c106 18 0 3.20827e-20 $X=3.525 $Y=1.59
c107 16 0 1.93585e-19 $X=3.14 $Y=1.59
c108 13 0 6.05954e-20 $X=3.575 $Y=2.03
r109 43 44 8.49906 $w=3.53e-07 $l=1.65e-07 $layer=LI1_cond $X=0.267 $Y=2.24
+ $X2=0.267 $Y2=2.075
r110 41 44 69.1551 $w=1.68e-07 $l=1.06e-06 $layer=LI1_cond $X=0.175 $Y=1.015
+ $X2=0.175 $Y2=2.075
r111 39 41 10.1222 $w=3.53e-07 $l=2.15e-07 $layer=LI1_cond $X=0.267 $Y=0.8
+ $X2=0.267 $Y2=1.015
r112 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.915
+ $Y=1.59 $X2=2.915 $Y2=1.59
r113 33 35 14.9023 $w=2.88e-07 $l=3.75e-07 $layer=LI1_cond $X=2.895 $Y=1.965
+ $X2=2.895 $Y2=1.59
r114 31 33 7.43784 $w=1.7e-07 $l=1.8262e-07 $layer=LI1_cond $X=2.75 $Y=2.05
+ $X2=2.895 $Y2=1.965
r115 31 32 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=2.75 $Y=2.05
+ $X2=1.985 $Y2=2.05
r116 29 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.9 $Y=2.135
+ $X2=1.985 $Y2=2.05
r117 29 30 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=1.9 $Y=2.135 $X2=1.9
+ $Y2=2.435
r118 28 45 4.08752 $w=1.7e-07 $l=1.78e-07 $layer=LI1_cond $X=0.445 $Y=2.52
+ $X2=0.267 $Y2=2.52
r119 27 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.815 $Y=2.52
+ $X2=1.9 $Y2=2.435
r120 27 28 89.3797 $w=1.68e-07 $l=1.37e-06 $layer=LI1_cond $X=1.815 $Y=2.52
+ $X2=0.445 $Y2=2.52
r121 24 45 2.70057 $w=3.55e-07 $l=8.5e-08 $layer=LI1_cond $X=0.267 $Y=2.435
+ $X2=0.267 $Y2=2.52
r122 23 43 0.389558 $w=3.53e-07 $l=1.2e-08 $layer=LI1_cond $X=0.267 $Y=2.252
+ $X2=0.267 $Y2=2.24
r123 23 24 5.94076 $w=3.53e-07 $l=1.83e-07 $layer=LI1_cond $X=0.267 $Y=2.252
+ $X2=0.267 $Y2=2.435
r124 17 18 54.207 $w=3.3e-07 $l=3.1e-07 $layer=POLY_cond $X=3.215 $Y=1.59
+ $X2=3.525 $Y2=1.59
r125 16 36 39.3438 $w=3.3e-07 $l=2.25e-07 $layer=POLY_cond $X=3.14 $Y=1.59
+ $X2=2.915 $Y2=1.59
r126 16 17 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=3.14 $Y=1.59
+ $X2=3.215 $Y2=1.59
r127 13 20 40.9178 $w=2.5e-07 $l=1.25e-07 $layer=POLY_cond $X=3.575 $Y=2.03
+ $X2=3.575 $Y2=1.905
r128 13 15 108.932 $w=2.5e-07 $l=5.65e-07 $layer=POLY_cond $X=3.575 $Y=2.03
+ $X2=3.575 $Y2=2.595
r129 11 18 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.525 $Y=1.755
+ $X2=3.525 $Y2=1.59
r130 11 20 76.9149 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=3.525 $Y=1.755
+ $X2=3.525 $Y2=1.905
r131 7 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.215 $Y=1.425
+ $X2=3.215 $Y2=1.59
r132 7 9 502.511 $w=1.5e-07 $l=9.8e-07 $layer=POLY_cond $X=3.215 $Y=1.425
+ $X2=3.215 $Y2=0.445
r133 2 43 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.095 $X2=0.28 $Y2=2.24
r134 1 39 182 $w=1.7e-07 $l=2.5229e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.61 $X2=0.28 $Y2=0.8
.ends

.subckt PM_SKY130_FD_SC_LP__DLRTP_LP2%A_413_47# 1 2 9 10 12 17 19 22 23 25 26 30
+ 32 35 36 40 44 45 46 50
c141 45 0 1.94025e-19 $X=4.595 $Y=1.43
c142 44 0 7.34056e-20 $X=4.595 $Y=1.43
c143 40 0 1.22967e-19 $X=3.695 $Y=0.93
c144 36 0 3.1823e-19 $X=3.715 $Y=0.81
c145 19 0 2.63828e-19 $X=3.57 $Y=0.81
r146 44 46 8.69073 $w=4.08e-07 $l=1.65e-07 $layer=LI1_cond $X=4.555 $Y=1.43
+ $X2=4.555 $Y2=1.265
r147 44 45 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.595
+ $Y=1.43 $X2=4.595 $Y2=1.43
r148 40 50 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.695 $Y=0.93
+ $X2=3.695 $Y2=0.765
r149 39 41 3.17915 $w=2.88e-07 $l=8e-08 $layer=LI1_cond $X=3.715 $Y=0.93
+ $X2=3.715 $Y2=1.01
r150 39 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.695
+ $Y=0.93 $X2=3.695 $Y2=0.93
r151 36 39 4.76873 $w=2.88e-07 $l=1.2e-07 $layer=LI1_cond $X=3.715 $Y=0.81
+ $X2=3.715 $Y2=0.93
r152 29 44 1.12433 $w=4.08e-07 $l=4e-08 $layer=LI1_cond $X=4.555 $Y=1.47
+ $X2=4.555 $Y2=1.43
r153 29 30 10.5406 $w=4.08e-07 $l=3.75e-07 $layer=LI1_cond $X=4.555 $Y=1.47
+ $X2=4.555 $Y2=1.845
r154 27 46 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=4.435 $Y=1.095
+ $X2=4.435 $Y2=1.265
r155 25 30 8.45803 $w=1.7e-07 $l=2.43824e-07 $layer=LI1_cond $X=4.35 $Y=1.93
+ $X2=4.555 $Y2=1.845
r156 25 26 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=4.35 $Y=1.93
+ $X2=3.985 $Y2=1.93
r157 24 41 3.86198 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=3.86 $Y=1.01
+ $X2=3.715 $Y2=1.01
r158 23 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.35 $Y=1.01
+ $X2=4.435 $Y2=1.095
r159 23 24 31.9679 $w=1.68e-07 $l=4.9e-07 $layer=LI1_cond $X=4.35 $Y=1.01
+ $X2=3.86 $Y2=1.01
r160 21 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.9 $Y=2.015
+ $X2=3.985 $Y2=1.93
r161 21 22 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=3.9 $Y=2.015 $X2=3.9
+ $Y2=2.315
r162 20 32 12.0232 $w=3.45e-07 $l=4.36348e-07 $layer=LI1_cond $X=2.485 $Y=0.81
+ $X2=2.265 $Y2=0.47
r163 19 36 3.86198 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=3.57 $Y=0.81
+ $X2=3.715 $Y2=0.81
r164 19 20 70.7861 $w=1.68e-07 $l=1.085e-06 $layer=LI1_cond $X=3.57 $Y=0.81
+ $X2=2.485 $Y2=0.81
r165 18 35 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.415 $Y=2.4
+ $X2=2.29 $Y2=2.4
r166 17 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.815 $Y=2.4
+ $X2=3.9 $Y2=2.315
r167 17 18 91.3369 $w=1.68e-07 $l=1.4e-06 $layer=LI1_cond $X=3.815 $Y=2.4
+ $X2=2.415 $Y2=2.4
r168 14 45 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=4.595 $Y=1.77
+ $X2=4.595 $Y2=1.43
r169 10 14 30.6163 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.595 $Y=1.935
+ $X2=4.595 $Y2=1.77
r170 10 12 163.979 $w=2.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.595 $Y=1.935
+ $X2=4.595 $Y2=2.595
r171 9 50 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=3.605 $Y=0.445
+ $X2=3.605 $Y2=0.765
r172 2 35 300 $w=1.7e-07 $l=4.51719e-07 $layer=licon1_PDIFF $count=2 $X=2.105
+ $Y=2.095 $X2=2.25 $Y2=2.48
r173 1 32 182 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_NDIFF $count=1 $X=2.065
+ $Y=0.235 $X2=2.21 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_LP__DLRTP_LP2%A_898_21# 1 2 9 11 12 15 17 21 25 29 32 33
+ 36 42 44 45 50 53 55 56
c125 45 0 1.2537e-19 $X=6.07 $Y=0.96
c126 11 0 7.34056e-20 $X=4.97 $Y=0.93
r127 56 60 66.9034 $w=5.1e-07 $l=5.05e-07 $layer=POLY_cond $X=7.005 $Y=1.04
+ $X2=7.005 $Y2=1.545
r128 55 56 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.94
+ $Y=1.04 $X2=6.94 $Y2=1.04
r129 49 50 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.455
+ $Y=1.02 $X2=5.455 $Y2=1.02
r130 44 55 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.775 $Y=0.96
+ $X2=6.94 $Y2=0.96
r131 44 45 45.9947 $w=1.68e-07 $l=7.05e-07 $layer=LI1_cond $X=6.775 $Y=0.96
+ $X2=6.07 $Y2=0.96
r132 42 53 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=6.065 $Y=2.24
+ $X2=6.065 $Y2=2.075
r133 38 45 5.3796 $w=2.42e-07 $l=1.11018e-07 $layer=LI1_cond $X=5.985 $Y=1.02
+ $X2=6.07 $Y2=0.96
r134 38 53 67.1979 $w=1.68e-07 $l=1.03e-06 $layer=LI1_cond $X=5.985 $Y=1.045
+ $X2=5.985 $Y2=2.075
r135 34 38 6.95702 $w=2.42e-07 $l=1.38e-07 $layer=LI1_cond $X=5.847 $Y=1.02
+ $X2=5.985 $Y2=1.02
r136 34 49 19.762 $w=2.42e-07 $l=3.92e-07 $layer=LI1_cond $X=5.847 $Y=1.02
+ $X2=5.455 $Y2=1.02
r137 34 36 9.32313 $w=4.43e-07 $l=3.6e-07 $layer=LI1_cond $X=5.847 $Y=0.855
+ $X2=5.847 $Y2=0.495
r138 31 50 58.5785 $w=3.3e-07 $l=3.35e-07 $layer=POLY_cond $X=5.12 $Y=1.02
+ $X2=5.455 $Y2=1.02
r139 31 32 13.5877 $w=2.4e-07 $l=7.5e-08 $layer=POLY_cond $X=5.12 $Y=1.02
+ $X2=5.045 $Y2=1.02
r140 27 56 32.933 $w=2.55e-07 $l=2.49199e-07 $layer=POLY_cond $X=7.185 $Y=0.875
+ $X2=7.005 $Y2=1.04
r141 27 29 194.851 $w=1.5e-07 $l=3.8e-07 $layer=POLY_cond $X=7.185 $Y=0.875
+ $X2=7.185 $Y2=0.495
r142 25 60 260.876 $w=2.5e-07 $l=1.05e-06 $layer=POLY_cond $X=6.905 $Y=2.595
+ $X2=6.905 $Y2=1.545
r143 19 56 32.933 $w=2.55e-07 $l=2.49199e-07 $layer=POLY_cond $X=6.825 $Y=0.875
+ $X2=7.005 $Y2=1.04
r144 19 21 194.851 $w=1.5e-07 $l=3.8e-07 $layer=POLY_cond $X=6.825 $Y=0.875
+ $X2=6.825 $Y2=0.495
r145 15 33 40.9178 $w=2.5e-07 $l=1.25e-07 $layer=POLY_cond $X=5.095 $Y=1.55
+ $X2=5.095 $Y2=1.425
r146 15 17 259.634 $w=2.5e-07 $l=1.045e-06 $layer=POLY_cond $X=5.095 $Y=1.55
+ $X2=5.095 $Y2=2.595
r147 13 32 12.1617 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.045 $Y=1.185
+ $X2=5.045 $Y2=1.02
r148 13 33 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=5.045 $Y=1.185
+ $X2=5.045 $Y2=1.425
r149 11 32 13.5877 $w=2.4e-07 $l=1.21861e-07 $layer=POLY_cond $X=4.97 $Y=0.93
+ $X2=5.045 $Y2=1.02
r150 11 12 169.213 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=4.97 $Y=0.93
+ $X2=4.64 $Y2=0.93
r151 7 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.565 $Y=0.855
+ $X2=4.64 $Y2=0.93
r152 7 9 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=4.565 $Y=0.855
+ $X2=4.565 $Y2=0.445
r153 2 42 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=5.925
+ $Y=2.095 $X2=6.065 $Y2=2.24
r154 1 36 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=5.645
+ $Y=0.285 $X2=5.79 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__DLRTP_LP2%A_736_47# 1 2 9 12 15 19 21 27 30 32 34 37
+ 41 44 46 50
c109 44 0 2.97072e-19 $X=5.025 $Y=0.94
c110 41 0 6.05954e-20 $X=4.33 $Y=2.36
c111 9 0 1.30515e-19 $X=5.8 $Y=2.595
r112 49 50 18.3604 $w=3.3e-07 $l=1.05e-07 $layer=POLY_cond $X=5.8 $Y=1.59
+ $X2=5.905 $Y2=1.59
r113 42 44 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=4.785 $Y=0.94
+ $X2=5.025 $Y2=0.94
r114 38 49 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=5.595 $Y=1.59
+ $X2=5.8 $Y2=1.59
r115 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.595
+ $Y=1.59 $X2=5.595 $Y2=1.59
r116 35 46 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.11 $Y=1.59
+ $X2=5.025 $Y2=1.59
r117 35 37 16.9374 $w=3.28e-07 $l=4.85e-07 $layer=LI1_cond $X=5.11 $Y=1.59
+ $X2=5.595 $Y2=1.59
r118 33 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.025 $Y=1.755
+ $X2=5.025 $Y2=1.59
r119 33 34 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=5.025 $Y=1.755
+ $X2=5.025 $Y2=2.195
r120 32 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.025 $Y=1.425
+ $X2=5.025 $Y2=1.59
r121 31 44 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.025 $Y=1.025
+ $X2=5.025 $Y2=0.94
r122 31 32 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=5.025 $Y=1.025
+ $X2=5.025 $Y2=1.425
r123 30 42 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.785 $Y=0.855
+ $X2=4.785 $Y2=0.94
r124 29 30 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=4.785 $Y=0.545
+ $X2=4.785 $Y2=0.855
r125 28 41 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.495 $Y=2.28
+ $X2=4.33 $Y2=2.28
r126 27 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.94 $Y=2.28
+ $X2=5.025 $Y2=2.195
r127 27 28 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=4.94 $Y=2.28
+ $X2=4.495 $Y2=2.28
r128 21 29 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=4.7 $Y=0.42
+ $X2=4.785 $Y2=0.545
r129 21 23 34.1123 $w=2.48e-07 $l=7.4e-07 $layer=LI1_cond $X=4.7 $Y=0.42
+ $X2=3.96 $Y2=0.42
r130 17 19 51.2766 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=5.905 $Y=0.91
+ $X2=6.005 $Y2=0.91
r131 13 19 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.005 $Y=0.835
+ $X2=6.005 $Y2=0.91
r132 13 15 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=6.005 $Y=0.835
+ $X2=6.005 $Y2=0.495
r133 12 50 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.905 $Y=1.425
+ $X2=5.905 $Y2=1.59
r134 11 17 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.905 $Y=0.985
+ $X2=5.905 $Y2=0.91
r135 11 12 225.617 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=5.905 $Y=0.985
+ $X2=5.905 $Y2=1.425
r136 7 49 9.34494 $w=2.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.8 $Y=1.755
+ $X2=5.8 $Y2=1.59
r137 7 9 208.701 $w=2.5e-07 $l=8.4e-07 $layer=POLY_cond $X=5.8 $Y=1.755 $X2=5.8
+ $Y2=2.595
r138 2 41 300 $w=1.7e-07 $l=3.27605e-07 $layer=licon1_PDIFF $count=2 $X=4.19
+ $Y=2.095 $X2=4.33 $Y2=2.36
r139 1 23 182 $w=1.7e-07 $l=3.44964e-07 $layer=licon1_NDIFF $count=1 $X=3.68
+ $Y=0.235 $X2=3.96 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_LP__DLRTP_LP2%RESET_B 2 5 9 11 12 15 16
c40 16 0 1.30515e-19 $X=6.375 $Y=1.39
c41 9 0 1.2537e-19 $X=6.395 $Y=0.495
r42 15 17 46.255 $w=3.35e-07 $l=1.65e-07 $layer=POLY_cond $X=6.372 $Y=1.39
+ $X2=6.372 $Y2=1.225
r43 15 16 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.375
+ $Y=1.39 $X2=6.375 $Y2=1.39
r44 12 16 9.18614 $w=3.43e-07 $l=2.75e-07 $layer=LI1_cond $X=6.422 $Y=1.665
+ $X2=6.422 $Y2=1.39
r45 9 17 374.319 $w=1.5e-07 $l=7.3e-07 $layer=POLY_cond $X=6.395 $Y=0.495
+ $X2=6.395 $Y2=1.225
r46 5 11 173.918 $w=2.5e-07 $l=7e-07 $layer=POLY_cond $X=6.33 $Y=2.595 $X2=6.33
+ $Y2=1.895
r47 2 11 32.6064 $w=3.35e-07 $l=1.67e-07 $layer=POLY_cond $X=6.372 $Y=1.728
+ $X2=6.372 $Y2=1.895
r48 1 15 0.344503 $w=3.35e-07 $l=2e-09 $layer=POLY_cond $X=6.372 $Y=1.392
+ $X2=6.372 $Y2=1.39
r49 1 2 57.8765 $w=3.35e-07 $l=3.36e-07 $layer=POLY_cond $X=6.372 $Y=1.392
+ $X2=6.372 $Y2=1.728
.ends

.subckt PM_SKY130_FD_SC_LP__DLRTP_LP2%VPWR 1 2 3 4 17 21 25 29 33 37 39 44 54 55
+ 58 61 64 67
r81 67 68 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r82 65 68 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=6.48 $Y2=3.33
r83 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r84 61 62 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r85 58 59 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r86 55 68 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=6.48 $Y2=3.33
r87 54 55 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r88 52 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.76 $Y=3.33
+ $X2=6.595 $Y2=3.33
r89 52 54 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=6.76 $Y=3.33
+ $X2=7.44 $Y2=3.33
r90 51 65 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=5.52 $Y2=3.33
r91 50 51 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r92 48 62 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.64 $Y2=3.33
r93 47 50 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=3.12 $Y=3.33
+ $X2=5.04 $Y2=3.33
r94 47 48 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r95 45 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.945 $Y=3.33
+ $X2=2.78 $Y2=3.33
r96 45 47 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=2.945 $Y=3.33
+ $X2=3.12 $Y2=3.33
r97 44 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.29 $Y=3.33
+ $X2=5.455 $Y2=3.33
r98 44 50 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=5.29 $Y=3.33
+ $X2=5.04 $Y2=3.33
r99 43 62 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r100 43 59 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r101 42 43 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r102 40 58 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.975 $Y=3.33
+ $X2=0.81 $Y2=3.33
r103 40 42 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=0.975 $Y=3.33
+ $X2=1.2 $Y2=3.33
r104 39 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.615 $Y=3.33
+ $X2=2.78 $Y2=3.33
r105 39 42 92.3155 $w=1.68e-07 $l=1.415e-06 $layer=LI1_cond $X=2.615 $Y=3.33
+ $X2=1.2 $Y2=3.33
r106 37 51 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=3.84 $Y=3.33
+ $X2=5.04 $Y2=3.33
r107 37 48 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=3.84 $Y=3.33
+ $X2=3.12 $Y2=3.33
r108 33 36 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=6.595 $Y=2.24
+ $X2=6.595 $Y2=2.95
r109 31 67 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.595 $Y=3.245
+ $X2=6.595 $Y2=3.33
r110 31 36 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=6.595 $Y=3.245
+ $X2=6.595 $Y2=2.95
r111 30 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.62 $Y=3.33
+ $X2=5.455 $Y2=3.33
r112 29 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.43 $Y=3.33
+ $X2=6.595 $Y2=3.33
r113 29 30 52.8449 $w=1.68e-07 $l=8.1e-07 $layer=LI1_cond $X=6.43 $Y=3.33
+ $X2=5.62 $Y2=3.33
r114 25 28 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=5.455 $Y=2.24
+ $X2=5.455 $Y2=2.95
r115 23 64 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.455 $Y=3.245
+ $X2=5.455 $Y2=3.33
r116 23 28 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=5.455 $Y=3.245
+ $X2=5.455 $Y2=2.95
r117 19 61 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.78 $Y=3.245
+ $X2=2.78 $Y2=3.33
r118 19 21 13.7944 $w=3.28e-07 $l=3.95e-07 $layer=LI1_cond $X=2.78 $Y=3.245
+ $X2=2.78 $Y2=2.85
r119 15 58 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.81 $Y=3.245
+ $X2=0.81 $Y2=3.33
r120 15 17 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.81 $Y=3.245
+ $X2=0.81 $Y2=2.95
r121 4 36 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=6.455
+ $Y=2.095 $X2=6.595 $Y2=2.95
r122 4 33 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=6.455
+ $Y=2.095 $X2=6.595 $Y2=2.24
r123 3 28 400 $w=1.7e-07 $l=9.65376e-07 $layer=licon1_PDIFF $count=1 $X=5.22
+ $Y=2.095 $X2=5.455 $Y2=2.95
r124 3 25 400 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_PDIFF $count=1 $X=5.22
+ $Y=2.095 $X2=5.455 $Y2=2.24
r125 2 21 600 $w=1.7e-07 $l=8.22025e-07 $layer=licon1_PDIFF $count=1 $X=2.64
+ $Y=2.095 $X2=2.78 $Y2=2.85
r126 1 17 600 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=0.67
+ $Y=2.095 $X2=0.81 $Y2=2.95
.ends

.subckt PM_SKY130_FD_SC_LP__DLRTP_LP2%Q 1 2 7 8 9 10 11 12 13 36 39
r19 37 39 1.06793 $w=5.58e-07 $l=5e-08 $layer=LI1_cond $X=7.285 $Y=2.355
+ $X2=7.285 $Y2=2.405
r20 36 45 1.84391 $w=2.48e-07 $l=4e-08 $layer=LI1_cond $X=7.44 $Y=2.035 $X2=7.44
+ $Y2=2.075
r21 12 37 0.384454 $w=5.58e-07 $l=1.8e-08 $layer=LI1_cond $X=7.285 $Y=2.337
+ $X2=7.285 $Y2=2.355
r22 12 47 2.07178 $w=5.58e-07 $l=9.7e-08 $layer=LI1_cond $X=7.285 $Y=2.337
+ $X2=7.285 $Y2=2.24
r23 12 13 7.53957 $w=5.58e-07 $l=3.53e-07 $layer=LI1_cond $X=7.285 $Y=2.422
+ $X2=7.285 $Y2=2.775
r24 12 39 0.363095 $w=5.58e-07 $l=1.7e-08 $layer=LI1_cond $X=7.285 $Y=2.422
+ $X2=7.285 $Y2=2.405
r25 11 47 3.05427 $w=5.58e-07 $l=1.43e-07 $layer=LI1_cond $X=7.285 $Y=2.097
+ $X2=7.285 $Y2=2.24
r26 11 45 4.18591 $w=5.58e-07 $l=2.2e-08 $layer=LI1_cond $X=7.285 $Y=2.097
+ $X2=7.285 $Y2=2.075
r27 11 36 1.06025 $w=2.48e-07 $l=2.3e-08 $layer=LI1_cond $X=7.44 $Y=2.012
+ $X2=7.44 $Y2=2.035
r28 10 11 15.9959 $w=2.48e-07 $l=3.47e-07 $layer=LI1_cond $X=7.44 $Y=1.665
+ $X2=7.44 $Y2=2.012
r29 9 10 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=7.44 $Y=1.295
+ $X2=7.44 $Y2=1.665
r30 8 9 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=7.44 $Y=0.925 $X2=7.44
+ $Y2=1.295
r31 7 8 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=7.44 $Y=0.495 $X2=7.44
+ $Y2=0.925
r32 2 47 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=7.03
+ $Y=2.095 $X2=7.17 $Y2=2.24
r33 1 7 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=7.26
+ $Y=0.285 $X2=7.4 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__DLRTP_LP2%VGND 1 2 3 4 15 19 23 27 30 31 32 34 39 48
+ 54 55 58 61 64
c96 39 0 1.06646e-19 $X=2.835 $Y=0
r97 64 65 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r98 61 62 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r99 58 59 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r100 55 65 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.44 $Y=0 $X2=6.48
+ $Y2=0
r101 54 55 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r102 52 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.775 $Y=0 $X2=6.61
+ $Y2=0
r103 52 54 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=6.775 $Y=0 $X2=7.44
+ $Y2=0
r104 51 65 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=6.48
+ $Y2=0
r105 50 51 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r106 48 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.445 $Y=0 $X2=6.61
+ $Y2=0
r107 48 50 60.3476 $w=1.68e-07 $l=9.25e-07 $layer=LI1_cond $X=6.445 $Y=0
+ $X2=5.52 $Y2=0
r108 47 51 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=5.52
+ $Y2=0
r109 46 47 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.04 $Y=0
+ $X2=5.04 $Y2=0
r110 44 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.165 $Y=0 $X2=3
+ $Y2=0
r111 44 46 122.326 $w=1.68e-07 $l=1.875e-06 $layer=LI1_cond $X=3.165 $Y=0
+ $X2=5.04 $Y2=0
r112 43 62 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r113 43 59 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=2.64 $Y=0 $X2=1.2
+ $Y2=0
r114 42 43 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r115 40 58 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.265 $Y=0 $X2=1.1
+ $Y2=0
r116 40 42 89.7059 $w=1.68e-07 $l=1.375e-06 $layer=LI1_cond $X=1.265 $Y=0
+ $X2=2.64 $Y2=0
r117 39 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.835 $Y=0 $X2=3
+ $Y2=0
r118 39 42 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=2.835 $Y=0
+ $X2=2.64 $Y2=0
r119 37 59 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r120 36 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r121 34 58 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.935 $Y=0 $X2=1.1
+ $Y2=0
r122 34 36 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=0.935 $Y=0
+ $X2=0.72 $Y2=0
r123 32 47 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=3.84 $Y=0 $X2=5.04
+ $Y2=0
r124 32 62 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=3.84 $Y=0 $X2=3.12
+ $Y2=0
r125 30 46 0.652406 $w=1.68e-07 $l=1e-08 $layer=LI1_cond $X=5.05 $Y=0 $X2=5.04
+ $Y2=0
r126 30 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.05 $Y=0 $X2=5.215
+ $Y2=0
r127 29 50 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=5.38 $Y=0 $X2=5.52
+ $Y2=0
r128 29 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.38 $Y=0 $X2=5.215
+ $Y2=0
r129 25 64 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.61 $Y=0.085
+ $X2=6.61 $Y2=0
r130 25 27 13.7944 $w=3.28e-07 $l=3.95e-07 $layer=LI1_cond $X=6.61 $Y=0.085
+ $X2=6.61 $Y2=0.48
r131 21 31 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.215 $Y=0.085
+ $X2=5.215 $Y2=0
r132 21 23 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=5.215 $Y=0.085
+ $X2=5.215 $Y2=0.445
r133 17 61 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3 $Y=0.085 $X2=3
+ $Y2=0
r134 17 19 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=3 $Y=0.085 $X2=3
+ $Y2=0.38
r135 13 58 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.1 $Y=0.085 $X2=1.1
+ $Y2=0
r136 13 15 24.9696 $w=3.28e-07 $l=7.15e-07 $layer=LI1_cond $X=1.1 $Y=0.085
+ $X2=1.1 $Y2=0.8
r137 4 27 182 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_NDIFF $count=1 $X=6.47
+ $Y=0.285 $X2=6.61 $Y2=0.48
r138 3 23 182 $w=1.7e-07 $l=6.71844e-07 $layer=licon1_NDIFF $count=1 $X=4.64
+ $Y=0.235 $X2=5.215 $Y2=0.445
r139 2 19 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=2.86
+ $Y=0.235 $X2=3 $Y2=0.38
r140 1 15 182 $w=1.7e-07 $l=2.504e-07 $layer=licon1_NDIFF $count=1 $X=0.96
+ $Y=0.61 $X2=1.1 $Y2=0.8
.ends

