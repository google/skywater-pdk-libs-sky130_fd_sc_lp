* NGSPICE file created from sky130_fd_sc_lp__dlrtp_2.ext - technology: sky130A

.subckt sky130_fd_sc_lp__dlrtp_2 D GATE RESET_B VGND VNB VPB VPWR Q
M1000 VPWR a_796_21# a_785_479# VPB phighvt w=420000u l=150000u
+  ad=2.2398e+12p pd=1.537e+07u as=1.008e+11p ps=1.32e+06u
M1001 VPWR a_796_21# Q VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=3.528e+11p ps=3.08e+06u
M1002 VGND RESET_B a_1043_73# VNB nshort w=840000u l=150000u
+  ad=1.1025e+12p pd=9.76e+06u as=1.764e+11p ps=2.1e+06u
M1003 a_251_475# GATE VPWR VPB phighvt w=640000u l=150000u
+  ad=2.08e+11p pd=1.93e+06u as=0p ps=0u
M1004 a_574_47# a_40_54# VGND VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1005 VGND a_796_21# a_754_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1006 Q a_796_21# VGND VNB nshort w=840000u l=150000u
+  ad=3.318e+11p pd=2.47e+06u as=0p ps=0u
M1007 a_646_47# a_383_479# a_574_47# VNB nshort w=420000u l=150000u
+  ad=1.638e+11p pd=1.62e+06u as=0p ps=0u
M1008 a_1043_73# a_646_47# a_796_21# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=2.226e+11p ps=2.21e+06u
M1009 Q a_796_21# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_611_479# a_40_54# VPWR VPB phighvt w=640000u l=150000u
+  ad=1.344e+11p pd=1.7e+06u as=0p ps=0u
M1011 VGND D a_40_54# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1012 a_796_21# a_646_47# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=3.528e+11p pd=3.08e+06u as=0p ps=0u
M1013 a_646_47# a_251_475# a_611_479# VPB phighvt w=640000u l=150000u
+  ad=2.062e+11p pd=2e+06u as=0p ps=0u
M1014 a_785_479# a_383_479# a_646_47# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_754_47# a_251_475# a_646_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VGND a_796_21# Q VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VPWR D a_40_54# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.696e+11p ps=1.81e+06u
M1018 VPWR RESET_B a_796_21# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_251_475# GATE VGND VNB nshort w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=0p ps=0u
M1020 VPWR a_251_475# a_383_479# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.696e+11p ps=1.81e+06u
M1021 VGND a_251_475# a_383_479# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
.ends

