* File: sky130_fd_sc_lp__and2_4.pxi.spice
* Created: Fri Aug 28 10:04:30 2020
* 
x_PM_SKY130_FD_SC_LP__AND2_4%A N_A_c_64_n N_A_M1004_g N_A_c_65_n N_A_M1011_g A
+ N_A_c_67_n PM_SKY130_FD_SC_LP__AND2_4%A
x_PM_SKY130_FD_SC_LP__AND2_4%B N_B_M1000_g N_B_M1005_g B N_B_c_89_n N_B_c_90_n
+ PM_SKY130_FD_SC_LP__AND2_4%B
x_PM_SKY130_FD_SC_LP__AND2_4%A_27_47# N_A_27_47#_M1004_s N_A_27_47#_M1011_d
+ N_A_27_47#_M1002_g N_A_27_47#_M1001_g N_A_27_47#_M1003_g N_A_27_47#_M1006_g
+ N_A_27_47#_M1007_g N_A_27_47#_M1008_g N_A_27_47#_M1009_g N_A_27_47#_M1010_g
+ N_A_27_47#_c_133_n N_A_27_47#_c_134_n N_A_27_47#_c_135_n N_A_27_47#_c_160_n
+ N_A_27_47#_c_188_p N_A_27_47#_c_161_n N_A_27_47#_c_136_n N_A_27_47#_c_137_n
+ N_A_27_47#_c_197_p N_A_27_47#_c_138_n N_A_27_47#_c_139_n
+ PM_SKY130_FD_SC_LP__AND2_4%A_27_47#
x_PM_SKY130_FD_SC_LP__AND2_4%VPWR N_VPWR_M1011_s N_VPWR_M1005_d N_VPWR_M1006_d
+ N_VPWR_M1010_d N_VPWR_c_244_n N_VPWR_c_245_n N_VPWR_c_246_n N_VPWR_c_247_n
+ N_VPWR_c_248_n N_VPWR_c_249_n N_VPWR_c_250_n N_VPWR_c_251_n N_VPWR_c_252_n
+ N_VPWR_c_253_n VPWR N_VPWR_c_254_n N_VPWR_c_243_n N_VPWR_c_256_n
+ PM_SKY130_FD_SC_LP__AND2_4%VPWR
x_PM_SKY130_FD_SC_LP__AND2_4%X N_X_M1002_d N_X_M1007_d N_X_M1001_s N_X_M1008_s
+ N_X_c_350_p N_X_c_336_n N_X_c_296_n N_X_c_297_n N_X_c_302_n N_X_c_303_n
+ N_X_c_351_p N_X_c_340_n N_X_c_298_n N_X_c_304_n N_X_c_299_n N_X_c_305_n X X
+ N_X_c_300_n X PM_SKY130_FD_SC_LP__AND2_4%X
x_PM_SKY130_FD_SC_LP__AND2_4%VGND N_VGND_M1000_d N_VGND_M1003_s N_VGND_M1009_s
+ N_VGND_c_358_n N_VGND_c_359_n N_VGND_c_360_n N_VGND_c_361_n N_VGND_c_362_n
+ N_VGND_c_363_n N_VGND_c_364_n N_VGND_c_365_n VGND N_VGND_c_366_n
+ N_VGND_c_367_n N_VGND_c_368_n PM_SKY130_FD_SC_LP__AND2_4%VGND
cc_1 VNB N_A_c_64_n 0.0195908f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.185
cc_2 VNB N_A_c_65_n 0.0614254f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.725
cc_3 VNB N_B_M1000_g 0.0249601f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.655
cc_4 VNB N_B_c_89_n 0.0253822f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.46
cc_5 VNB N_B_c_90_n 0.00434342f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_6 VNB N_A_27_47#_M1002_g 0.0246709f $X=-0.19 $Y=-0.245 $X2=0.337 $Y2=1.46
cc_7 VNB N_A_27_47#_M1003_g 0.0222554f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_27_47#_M1007_g 0.0222417f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_27_47#_M1009_g 0.0270419f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_27_47#_c_133_n 0.0285043f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_27_47#_c_134_n 0.00900767f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_27_47#_c_135_n 0.0102153f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_27_47#_c_136_n 0.00224589f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_27_47#_c_137_n 2.8618e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_27_47#_c_138_n 0.00119389f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_27_47#_c_139_n 0.0677742f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_VPWR_c_243_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_X_c_296_n 0.00304705f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_X_c_297_n 0.00262701f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_X_c_298_n 0.0014502f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_X_c_299_n 0.00144314f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_X_c_300_n 0.0165544f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB X 0.0247464f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_VGND_c_358_n 0.00501393f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.46
cc_25 VNB N_VGND_c_359_n 3.21684e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_360_n 0.0280468f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_361_n 0.0163732f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_362_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_363_n 0.0110534f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_364_n 0.0129398f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_365_n 0.00513431f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_366_n 0.0293201f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_367_n 0.19553f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_368_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VPB N_A_c_65_n 0.0369534f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=1.725
cc_36 VPB N_A_c_67_n 0.00347908f $X=-0.19 $Y=1.655 $X2=0.29 $Y2=1.46
cc_37 VPB N_B_M1005_g 0.019316f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_38 VPB N_B_c_89_n 0.00619162f $X=-0.19 $Y=1.655 $X2=0.29 $Y2=1.46
cc_39 VPB N_B_c_90_n 0.00328307f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_40 VPB N_A_27_47#_M1001_g 0.0193736f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_41 VPB N_A_27_47#_M1006_g 0.0185138f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_42 VPB N_A_27_47#_M1008_g 0.0185005f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_43 VPB N_A_27_47#_M1010_g 0.0218053f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_44 VPB N_A_27_47#_c_137_n 0.00141893f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_45 VPB N_A_27_47#_c_139_n 0.00893444f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_46 VPB N_VPWR_c_244_n 0.0103398f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_47 VPB N_VPWR_c_245_n 0.0492812f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_48 VPB N_VPWR_c_246_n 0.00431378f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_49 VPB N_VPWR_c_247_n 3.16049e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_50 VPB N_VPWR_c_248_n 0.0408143f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_51 VPB N_VPWR_c_249_n 0.0152595f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_52 VPB N_VPWR_c_250_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_53 VPB N_VPWR_c_251_n 0.0110534f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_54 VPB N_VPWR_c_252_n 0.0129398f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_55 VPB N_VPWR_c_253_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_56 VPB N_VPWR_c_254_n 0.0151004f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_57 VPB N_VPWR_c_243_n 0.0511401f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_58 VPB N_VPWR_c_256_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_59 VPB N_X_c_302_n 0.00304888f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_60 VPB N_X_c_303_n 0.00187836f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_61 VPB N_X_c_304_n 0.0176422f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_62 VPB N_X_c_305_n 0.00144499f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_63 VPB X 0.00709707f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_64 N_A_c_64_n N_B_M1000_g 0.0759723f $X=0.475 $Y=1.185 $X2=0 $Y2=0
cc_65 N_A_c_65_n N_B_M1000_g 0.00920199f $X=0.475 $Y=1.725 $X2=0 $Y2=0
cc_66 N_A_c_67_n N_B_M1000_g 3.4125e-19 $X=0.29 $Y=1.46 $X2=0 $Y2=0
cc_67 N_A_c_65_n N_B_M1005_g 0.0180283f $X=0.475 $Y=1.725 $X2=0 $Y2=0
cc_68 N_A_c_65_n N_B_c_89_n 0.00630129f $X=0.475 $Y=1.725 $X2=0 $Y2=0
cc_69 N_A_c_65_n N_B_c_90_n 0.00304452f $X=0.475 $Y=1.725 $X2=0 $Y2=0
cc_70 N_A_c_67_n N_B_c_90_n 0.0325794f $X=0.29 $Y=1.46 $X2=0 $Y2=0
cc_71 N_A_c_64_n N_A_27_47#_c_133_n 0.0151188f $X=0.475 $Y=1.185 $X2=0 $Y2=0
cc_72 N_A_c_64_n N_A_27_47#_c_134_n 0.0107927f $X=0.475 $Y=1.185 $X2=0 $Y2=0
cc_73 N_A_c_65_n N_A_27_47#_c_134_n 5.02965e-19 $X=0.475 $Y=1.725 $X2=0 $Y2=0
cc_74 N_A_c_67_n N_A_27_47#_c_134_n 0.00209071f $X=0.29 $Y=1.46 $X2=0 $Y2=0
cc_75 N_A_c_64_n N_A_27_47#_c_135_n 0.0023491f $X=0.475 $Y=1.185 $X2=0 $Y2=0
cc_76 N_A_c_65_n N_A_27_47#_c_135_n 0.00839838f $X=0.475 $Y=1.725 $X2=0 $Y2=0
cc_77 N_A_c_67_n N_A_27_47#_c_135_n 0.0256673f $X=0.29 $Y=1.46 $X2=0 $Y2=0
cc_78 N_A_c_65_n N_VPWR_c_245_n 0.0223827f $X=0.475 $Y=1.725 $X2=0 $Y2=0
cc_79 N_A_c_67_n N_VPWR_c_245_n 0.0236779f $X=0.29 $Y=1.46 $X2=0 $Y2=0
cc_80 N_A_c_65_n N_VPWR_c_254_n 0.00486043f $X=0.475 $Y=1.725 $X2=0 $Y2=0
cc_81 N_A_c_65_n N_VPWR_c_243_n 0.0082726f $X=0.475 $Y=1.725 $X2=0 $Y2=0
cc_82 N_A_c_64_n N_VGND_c_366_n 0.0054895f $X=0.475 $Y=1.185 $X2=0 $Y2=0
cc_83 N_A_c_64_n N_VGND_c_367_n 0.0107853f $X=0.475 $Y=1.185 $X2=0 $Y2=0
cc_84 N_B_M1000_g N_A_27_47#_M1002_g 0.0287785f $X=0.835 $Y=0.655 $X2=0 $Y2=0
cc_85 N_B_M1005_g N_A_27_47#_M1001_g 0.0255037f $X=0.905 $Y=2.465 $X2=0 $Y2=0
cc_86 N_B_c_90_n N_A_27_47#_M1001_g 2.01698e-19 $X=0.925 $Y=1.51 $X2=0 $Y2=0
cc_87 N_B_M1000_g N_A_27_47#_c_133_n 0.00243322f $X=0.835 $Y=0.655 $X2=0 $Y2=0
cc_88 N_B_M1000_g N_A_27_47#_c_134_n 0.0152408f $X=0.835 $Y=0.655 $X2=0 $Y2=0
cc_89 N_B_c_89_n N_A_27_47#_c_134_n 0.00330061f $X=0.925 $Y=1.51 $X2=0 $Y2=0
cc_90 N_B_c_90_n N_A_27_47#_c_134_n 0.029946f $X=0.925 $Y=1.51 $X2=0 $Y2=0
cc_91 N_B_c_90_n N_A_27_47#_c_160_n 0.0121915f $X=0.925 $Y=1.51 $X2=0 $Y2=0
cc_92 N_B_M1005_g N_A_27_47#_c_161_n 0.0134115f $X=0.905 $Y=2.465 $X2=0 $Y2=0
cc_93 N_B_c_89_n N_A_27_47#_c_161_n 0.0021314f $X=0.925 $Y=1.51 $X2=0 $Y2=0
cc_94 N_B_c_90_n N_A_27_47#_c_161_n 0.0139435f $X=0.925 $Y=1.51 $X2=0 $Y2=0
cc_95 N_B_M1000_g N_A_27_47#_c_136_n 0.00333998f $X=0.835 $Y=0.655 $X2=0 $Y2=0
cc_96 N_B_c_89_n N_A_27_47#_c_136_n 3.93074e-19 $X=0.925 $Y=1.51 $X2=0 $Y2=0
cc_97 N_B_c_90_n N_A_27_47#_c_136_n 0.00607903f $X=0.925 $Y=1.51 $X2=0 $Y2=0
cc_98 N_B_M1005_g N_A_27_47#_c_137_n 0.00390422f $X=0.905 $Y=2.465 $X2=0 $Y2=0
cc_99 N_B_c_89_n N_A_27_47#_c_137_n 4.59005e-19 $X=0.925 $Y=1.51 $X2=0 $Y2=0
cc_100 N_B_c_90_n N_A_27_47#_c_137_n 0.0112771f $X=0.925 $Y=1.51 $X2=0 $Y2=0
cc_101 N_B_c_89_n N_A_27_47#_c_138_n 0.00151598f $X=0.925 $Y=1.51 $X2=0 $Y2=0
cc_102 N_B_c_90_n N_A_27_47#_c_138_n 0.0171273f $X=0.925 $Y=1.51 $X2=0 $Y2=0
cc_103 N_B_c_89_n N_A_27_47#_c_139_n 0.0168015f $X=0.925 $Y=1.51 $X2=0 $Y2=0
cc_104 N_B_c_90_n N_A_27_47#_c_139_n 2.90095e-19 $X=0.925 $Y=1.51 $X2=0 $Y2=0
cc_105 N_B_M1005_g N_VPWR_c_245_n 7.40257e-19 $X=0.905 $Y=2.465 $X2=0 $Y2=0
cc_106 N_B_M1005_g N_VPWR_c_246_n 0.00273042f $X=0.905 $Y=2.465 $X2=0 $Y2=0
cc_107 N_B_M1005_g N_VPWR_c_254_n 0.00585385f $X=0.905 $Y=2.465 $X2=0 $Y2=0
cc_108 N_B_M1005_g N_VPWR_c_243_n 0.0107434f $X=0.905 $Y=2.465 $X2=0 $Y2=0
cc_109 N_B_M1000_g N_VGND_c_358_n 0.00672265f $X=0.835 $Y=0.655 $X2=0 $Y2=0
cc_110 N_B_M1000_g N_VGND_c_366_n 0.00585385f $X=0.835 $Y=0.655 $X2=0 $Y2=0
cc_111 N_B_M1000_g N_VGND_c_367_n 0.011026f $X=0.835 $Y=0.655 $X2=0 $Y2=0
cc_112 N_A_27_47#_c_161_n N_VPWR_M1005_d 0.00701161f $X=1.19 $Y=2.015 $X2=0
+ $Y2=0
cc_113 N_A_27_47#_c_137_n N_VPWR_M1005_d 0.00112177f $X=1.275 $Y=1.93 $X2=0
+ $Y2=0
cc_114 N_A_27_47#_M1001_g N_VPWR_c_246_n 0.0027042f $X=1.41 $Y=2.465 $X2=0 $Y2=0
cc_115 N_A_27_47#_c_161_n N_VPWR_c_246_n 0.0203005f $X=1.19 $Y=2.015 $X2=0 $Y2=0
cc_116 N_A_27_47#_M1001_g N_VPWR_c_247_n 7.37737e-19 $X=1.41 $Y=2.465 $X2=0
+ $Y2=0
cc_117 N_A_27_47#_M1006_g N_VPWR_c_247_n 0.0141689f $X=1.84 $Y=2.465 $X2=0 $Y2=0
cc_118 N_A_27_47#_M1008_g N_VPWR_c_247_n 0.014077f $X=2.27 $Y=2.465 $X2=0 $Y2=0
cc_119 N_A_27_47#_M1010_g N_VPWR_c_247_n 7.21513e-19 $X=2.7 $Y=2.465 $X2=0 $Y2=0
cc_120 N_A_27_47#_M1008_g N_VPWR_c_248_n 7.21513e-19 $X=2.27 $Y=2.465 $X2=0
+ $Y2=0
cc_121 N_A_27_47#_M1010_g N_VPWR_c_248_n 0.0150803f $X=2.7 $Y=2.465 $X2=0 $Y2=0
cc_122 N_A_27_47#_M1001_g N_VPWR_c_249_n 0.00585385f $X=1.41 $Y=2.465 $X2=0
+ $Y2=0
cc_123 N_A_27_47#_M1006_g N_VPWR_c_249_n 0.00486043f $X=1.84 $Y=2.465 $X2=0
+ $Y2=0
cc_124 N_A_27_47#_M1008_g N_VPWR_c_252_n 0.00486043f $X=2.27 $Y=2.465 $X2=0
+ $Y2=0
cc_125 N_A_27_47#_M1010_g N_VPWR_c_252_n 0.00486043f $X=2.7 $Y=2.465 $X2=0 $Y2=0
cc_126 N_A_27_47#_c_188_p N_VPWR_c_254_n 0.0124525f $X=0.69 $Y=2.91 $X2=0 $Y2=0
cc_127 N_A_27_47#_M1011_d N_VPWR_c_243_n 0.00536646f $X=0.55 $Y=1.835 $X2=0
+ $Y2=0
cc_128 N_A_27_47#_M1001_g N_VPWR_c_243_n 0.0107317f $X=1.41 $Y=2.465 $X2=0 $Y2=0
cc_129 N_A_27_47#_M1006_g N_VPWR_c_243_n 0.00824727f $X=1.84 $Y=2.465 $X2=0
+ $Y2=0
cc_130 N_A_27_47#_M1008_g N_VPWR_c_243_n 0.00824727f $X=2.27 $Y=2.465 $X2=0
+ $Y2=0
cc_131 N_A_27_47#_M1010_g N_VPWR_c_243_n 0.00824727f $X=2.7 $Y=2.465 $X2=0 $Y2=0
cc_132 N_A_27_47#_c_188_p N_VPWR_c_243_n 0.00730901f $X=0.69 $Y=2.91 $X2=0 $Y2=0
cc_133 N_A_27_47#_M1003_g N_X_c_296_n 0.0137623f $X=1.84 $Y=0.655 $X2=0 $Y2=0
cc_134 N_A_27_47#_M1007_g N_X_c_296_n 0.0141385f $X=2.27 $Y=0.655 $X2=0 $Y2=0
cc_135 N_A_27_47#_c_197_p N_X_c_296_n 0.0473014f $X=2.52 $Y=1.5 $X2=0 $Y2=0
cc_136 N_A_27_47#_c_139_n N_X_c_296_n 0.00243542f $X=2.7 $Y=1.5 $X2=0 $Y2=0
cc_137 N_A_27_47#_M1002_g N_X_c_297_n 0.00131418f $X=1.41 $Y=0.655 $X2=0 $Y2=0
cc_138 N_A_27_47#_c_134_n N_X_c_297_n 0.00750776f $X=1.19 $Y=1.07 $X2=0 $Y2=0
cc_139 N_A_27_47#_c_136_n N_X_c_297_n 0.00641961f $X=1.275 $Y=1.405 $X2=0 $Y2=0
cc_140 N_A_27_47#_c_197_p N_X_c_297_n 0.0154947f $X=2.52 $Y=1.5 $X2=0 $Y2=0
cc_141 N_A_27_47#_c_139_n N_X_c_297_n 0.00253619f $X=2.7 $Y=1.5 $X2=0 $Y2=0
cc_142 N_A_27_47#_M1006_g N_X_c_302_n 0.0128162f $X=1.84 $Y=2.465 $X2=0 $Y2=0
cc_143 N_A_27_47#_M1008_g N_X_c_302_n 0.0129249f $X=2.27 $Y=2.465 $X2=0 $Y2=0
cc_144 N_A_27_47#_c_197_p N_X_c_302_n 0.0473015f $X=2.52 $Y=1.5 $X2=0 $Y2=0
cc_145 N_A_27_47#_c_139_n N_X_c_302_n 0.00240656f $X=2.7 $Y=1.5 $X2=0 $Y2=0
cc_146 N_A_27_47#_M1001_g N_X_c_303_n 4.90985e-19 $X=1.41 $Y=2.465 $X2=0 $Y2=0
cc_147 N_A_27_47#_c_137_n N_X_c_303_n 0.00799443f $X=1.275 $Y=1.93 $X2=0 $Y2=0
cc_148 N_A_27_47#_c_197_p N_X_c_303_n 0.0154948f $X=2.52 $Y=1.5 $X2=0 $Y2=0
cc_149 N_A_27_47#_c_139_n N_X_c_303_n 0.00250529f $X=2.7 $Y=1.5 $X2=0 $Y2=0
cc_150 N_A_27_47#_M1009_g N_X_c_298_n 0.0169662f $X=2.7 $Y=0.655 $X2=0 $Y2=0
cc_151 N_A_27_47#_c_197_p N_X_c_298_n 0.00733859f $X=2.52 $Y=1.5 $X2=0 $Y2=0
cc_152 N_A_27_47#_M1010_g N_X_c_304_n 0.0157525f $X=2.7 $Y=2.465 $X2=0 $Y2=0
cc_153 N_A_27_47#_c_197_p N_X_c_304_n 0.00733859f $X=2.52 $Y=1.5 $X2=0 $Y2=0
cc_154 N_A_27_47#_c_197_p N_X_c_299_n 0.0154947f $X=2.52 $Y=1.5 $X2=0 $Y2=0
cc_155 N_A_27_47#_c_139_n N_X_c_299_n 0.00253619f $X=2.7 $Y=1.5 $X2=0 $Y2=0
cc_156 N_A_27_47#_c_197_p N_X_c_305_n 0.0154948f $X=2.52 $Y=1.5 $X2=0 $Y2=0
cc_157 N_A_27_47#_c_139_n N_X_c_305_n 0.00250529f $X=2.7 $Y=1.5 $X2=0 $Y2=0
cc_158 N_A_27_47#_M1009_g X 0.0212446f $X=2.7 $Y=0.655 $X2=0 $Y2=0
cc_159 N_A_27_47#_c_197_p X 0.0168735f $X=2.52 $Y=1.5 $X2=0 $Y2=0
cc_160 N_A_27_47#_c_134_n A_110_47# 0.00366293f $X=1.19 $Y=1.07 $X2=-0.19
+ $Y2=-0.245
cc_161 N_A_27_47#_c_134_n N_VGND_M1000_d 0.00365393f $X=1.19 $Y=1.07 $X2=-0.19
+ $Y2=-0.245
cc_162 N_A_27_47#_M1002_g N_VGND_c_358_n 0.0052226f $X=1.41 $Y=0.655 $X2=0 $Y2=0
cc_163 N_A_27_47#_c_134_n N_VGND_c_358_n 0.0260407f $X=1.19 $Y=1.07 $X2=0 $Y2=0
cc_164 N_A_27_47#_M1002_g N_VGND_c_359_n 6.58238e-19 $X=1.41 $Y=0.655 $X2=0
+ $Y2=0
cc_165 N_A_27_47#_M1003_g N_VGND_c_359_n 0.0112224f $X=1.84 $Y=0.655 $X2=0 $Y2=0
cc_166 N_A_27_47#_M1007_g N_VGND_c_359_n 0.0110534f $X=2.27 $Y=0.655 $X2=0 $Y2=0
cc_167 N_A_27_47#_M1009_g N_VGND_c_359_n 6.28154e-19 $X=2.7 $Y=0.655 $X2=0 $Y2=0
cc_168 N_A_27_47#_M1007_g N_VGND_c_360_n 6.28154e-19 $X=2.27 $Y=0.655 $X2=0
+ $Y2=0
cc_169 N_A_27_47#_M1009_g N_VGND_c_360_n 0.0123642f $X=2.7 $Y=0.655 $X2=0 $Y2=0
cc_170 N_A_27_47#_M1002_g N_VGND_c_361_n 0.00585385f $X=1.41 $Y=0.655 $X2=0
+ $Y2=0
cc_171 N_A_27_47#_M1003_g N_VGND_c_361_n 0.00486043f $X=1.84 $Y=0.655 $X2=0
+ $Y2=0
cc_172 N_A_27_47#_M1007_g N_VGND_c_364_n 0.00486043f $X=2.27 $Y=0.655 $X2=0
+ $Y2=0
cc_173 N_A_27_47#_M1009_g N_VGND_c_364_n 0.00486043f $X=2.7 $Y=0.655 $X2=0 $Y2=0
cc_174 N_A_27_47#_c_133_n N_VGND_c_366_n 0.0210467f $X=0.26 $Y=0.42 $X2=0 $Y2=0
cc_175 N_A_27_47#_M1004_s N_VGND_c_367_n 0.00215158f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_176 N_A_27_47#_M1002_g N_VGND_c_367_n 0.0110998f $X=1.41 $Y=0.655 $X2=0 $Y2=0
cc_177 N_A_27_47#_M1003_g N_VGND_c_367_n 0.00824727f $X=1.84 $Y=0.655 $X2=0
+ $Y2=0
cc_178 N_A_27_47#_M1007_g N_VGND_c_367_n 0.00824727f $X=2.27 $Y=0.655 $X2=0
+ $Y2=0
cc_179 N_A_27_47#_M1009_g N_VGND_c_367_n 0.00824727f $X=2.7 $Y=0.655 $X2=0 $Y2=0
cc_180 N_A_27_47#_c_133_n N_VGND_c_367_n 0.0125689f $X=0.26 $Y=0.42 $X2=0 $Y2=0
cc_181 N_VPWR_c_243_n N_X_M1001_s 0.00536646f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_182 N_VPWR_c_243_n N_X_M1008_s 0.00536646f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_183 N_VPWR_c_249_n N_X_c_336_n 0.0124525f $X=1.89 $Y=3.33 $X2=0 $Y2=0
cc_184 N_VPWR_c_243_n N_X_c_336_n 0.00730901f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_185 N_VPWR_M1006_d N_X_c_302_n 0.00176461f $X=1.915 $Y=1.835 $X2=0 $Y2=0
cc_186 N_VPWR_c_247_n N_X_c_302_n 0.0170777f $X=2.055 $Y=2.2 $X2=0 $Y2=0
cc_187 N_VPWR_c_252_n N_X_c_340_n 0.0124525f $X=2.75 $Y=3.33 $X2=0 $Y2=0
cc_188 N_VPWR_c_243_n N_X_c_340_n 0.00730901f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_189 N_VPWR_M1010_d N_X_c_304_n 0.00279864f $X=2.775 $Y=1.835 $X2=0 $Y2=0
cc_190 N_VPWR_c_248_n N_X_c_304_n 0.023955f $X=2.915 $Y=2.2 $X2=0 $Y2=0
cc_191 N_X_c_296_n N_VGND_M1003_s 0.00180746f $X=2.39 $Y=1.15 $X2=0 $Y2=0
cc_192 N_X_c_298_n N_VGND_M1009_s 2.39543e-19 $X=2.855 $Y=1.15 $X2=0 $Y2=0
cc_193 N_X_c_300_n N_VGND_M1009_s 0.00214448f $X=3.057 $Y=1.235 $X2=0 $Y2=0
cc_194 N_X_c_296_n N_VGND_c_359_n 0.0163515f $X=2.39 $Y=1.15 $X2=0 $Y2=0
cc_195 N_X_c_298_n N_VGND_c_360_n 0.00346358f $X=2.855 $Y=1.15 $X2=0 $Y2=0
cc_196 N_X_c_300_n N_VGND_c_360_n 0.0194858f $X=3.057 $Y=1.235 $X2=0 $Y2=0
cc_197 N_X_c_350_p N_VGND_c_361_n 0.0124525f $X=1.625 $Y=0.42 $X2=0 $Y2=0
cc_198 N_X_c_351_p N_VGND_c_364_n 0.0124525f $X=2.485 $Y=0.42 $X2=0 $Y2=0
cc_199 N_X_M1002_d N_VGND_c_367_n 0.00536646f $X=1.485 $Y=0.235 $X2=0 $Y2=0
cc_200 N_X_M1007_d N_VGND_c_367_n 0.00536646f $X=2.345 $Y=0.235 $X2=0 $Y2=0
cc_201 N_X_c_350_p N_VGND_c_367_n 0.00730901f $X=1.625 $Y=0.42 $X2=0 $Y2=0
cc_202 N_X_c_351_p N_VGND_c_367_n 0.00730901f $X=2.485 $Y=0.42 $X2=0 $Y2=0
cc_203 A_110_47# N_VGND_c_367_n 0.00899413f $X=0.55 $Y=0.235 $X2=0.425 $Y2=1.07
