* File: sky130_fd_sc_lp__einvp_m.pex.spice
* Created: Wed Sep  2 09:52:56 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__EINVP_M%TE 2 6 7 9 10 12 14 17 21 23 24 32
r53 30 32 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.64 $Y=0.37
+ $X2=0.805 $Y2=0.37
r54 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.64
+ $Y=0.37 $X2=0.64 $Y2=0.37
r55 27 30 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=0.55 $Y=0.37 $X2=0.64
+ $Y2=0.37
r56 24 31 2.59705 $w=3.53e-07 $l=8e-08 $layer=LI1_cond $X=0.72 $Y=0.462 $X2=0.64
+ $Y2=0.462
r57 23 31 12.9853 $w=3.53e-07 $l=4e-07 $layer=LI1_cond $X=0.24 $Y=0.462 $X2=0.64
+ $Y2=0.462
r58 19 21 87.1702 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=0.46 $Y=2.49
+ $X2=0.63 $Y2=2.49
r59 15 17 46.1489 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=0.46 $Y=1.25 $X2=0.55
+ $Y2=1.25
r60 12 14 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.06 $Y=0.535
+ $X2=1.06 $Y2=0.855
r61 10 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.985 $Y=0.46
+ $X2=1.06 $Y2=0.535
r62 10 32 92.2979 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=0.985 $Y=0.46
+ $X2=0.805 $Y2=0.46
r63 7 21 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.63 $Y=2.565
+ $X2=0.63 $Y2=2.49
r64 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.63 $Y=2.565 $X2=0.63
+ $Y2=2.885
r65 4 17 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.55 $Y=1.175
+ $X2=0.55 $Y2=1.25
r66 4 6 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.55 $Y=1.175 $X2=0.55
+ $Y2=0.855
r67 3 27 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.55 $Y=0.535
+ $X2=0.55 $Y2=0.37
r68 3 6 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.55 $Y=0.535 $X2=0.55
+ $Y2=0.855
r69 2 19 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.46 $Y=2.415
+ $X2=0.46 $Y2=2.49
r70 1 15 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.46 $Y=1.325
+ $X2=0.46 $Y2=1.25
r71 1 2 558.915 $w=1.5e-07 $l=1.09e-06 $layer=POLY_cond $X=0.46 $Y=1.325
+ $X2=0.46 $Y2=2.415
.ends

.subckt PM_SKY130_FD_SC_LP__EINVP_M%A_42_129# 1 2 9 13 16 20 22 26 28 29
r46 28 29 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.94 $Y=1.7
+ $X2=0.94 $Y2=1.7
r47 23 26 3.9231 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=0.52 $Y=1.62
+ $X2=0.345 $Y2=1.62
r48 22 28 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.855 $Y=1.62
+ $X2=0.94 $Y2=1.62
r49 22 23 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=0.855 $Y=1.62
+ $X2=0.52 $Y2=1.62
r50 18 26 2.80976 $w=3.4e-07 $l=8.5e-08 $layer=LI1_cond $X=0.345 $Y=1.705
+ $X2=0.345 $Y2=1.62
r51 18 20 36.7135 $w=3.48e-07 $l=1.115e-06 $layer=LI1_cond $X=0.345 $Y=1.705
+ $X2=0.345 $Y2=2.82
r52 14 26 2.80976 $w=3.4e-07 $l=8.9861e-08 $layer=LI1_cond $X=0.335 $Y=1.535
+ $X2=0.345 $Y2=1.62
r53 14 16 21.4773 $w=3.28e-07 $l=6.15e-07 $layer=LI1_cond $X=0.335 $Y=1.535
+ $X2=0.335 $Y2=0.92
r54 12 29 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=0.94 $Y=2.055
+ $X2=0.94 $Y2=1.7
r55 12 13 43.5886 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=0.955 $Y=2.055
+ $X2=0.955 $Y2=2.205
r56 9 13 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=1.06 $Y=2.885
+ $X2=1.06 $Y2=2.205
r57 2 20 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.29
+ $Y=2.675 $X2=0.415 $Y2=2.82
r58 1 16 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=0.21
+ $Y=0.645 $X2=0.335 $Y2=0.92
.ends

.subckt PM_SKY130_FD_SC_LP__EINVP_M%A 3 5 7 10 11
r24 10 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.51 $Y=0.37
+ $X2=1.51 $Y2=0.535
r25 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.51
+ $Y=0.37 $X2=1.51 $Y2=0.37
r26 7 11 4.8455 $w=4.38e-07 $l=1.85e-07 $layer=LI1_cond $X=1.545 $Y=0.555
+ $X2=1.545 $Y2=0.37
r27 3 5 1040.91 $w=1.5e-07 $l=2.03e-06 $layer=POLY_cond $X=1.42 $Y=0.855
+ $X2=1.42 $Y2=2.885
r28 3 13 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.42 $Y=0.855
+ $X2=1.42 $Y2=0.535
.ends

.subckt PM_SKY130_FD_SC_LP__EINVP_M%VPWR 1 6 9 10 11 18 19
r25 18 19 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r26 14 15 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r27 11 19 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=0.96 $Y=3.33
+ $X2=1.68 $Y2=3.33
r28 11 15 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=0.96 $Y=3.33
+ $X2=0.72 $Y2=3.33
r29 9 14 1.30481 $w=1.68e-07 $l=2e-08 $layer=LI1_cond $X=0.74 $Y=3.33 $X2=0.72
+ $Y2=3.33
r30 9 10 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=0.74 $Y=3.33
+ $X2=0.845 $Y2=3.33
r31 8 18 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=0.95 $Y=3.33 $X2=1.68
+ $Y2=3.33
r32 8 10 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=0.95 $Y=3.33
+ $X2=0.845 $Y2=3.33
r33 4 10 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=0.845 $Y=3.245
+ $X2=0.845 $Y2=3.33
r34 4 6 15.5801 $w=2.08e-07 $l=2.95e-07 $layer=LI1_cond $X=0.845 $Y=3.245
+ $X2=0.845 $Y2=2.95
r35 1 6 600 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=1 $X=0.705
+ $Y=2.675 $X2=0.845 $Y2=2.95
.ends

.subckt PM_SKY130_FD_SC_LP__EINVP_M%Z 1 2 7 8 9 10 11 12
r13 11 12 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.635 $Y=2.405
+ $X2=1.635 $Y2=2.775
r14 10 11 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.635 $Y=2.035
+ $X2=1.635 $Y2=2.405
r15 9 10 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.635 $Y=1.665
+ $X2=1.635 $Y2=2.035
r16 8 9 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.635 $Y=1.295
+ $X2=1.635 $Y2=1.665
r17 7 8 13.6198 $w=3.28e-07 $l=3.9e-07 $layer=LI1_cond $X=1.635 $Y=0.905
+ $X2=1.635 $Y2=1.295
r18 2 12 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.495
+ $Y=2.675 $X2=1.635 $Y2=2.82
r19 1 7 182 $w=1.7e-07 $l=3.2249e-07 $layer=licon1_NDIFF $count=1 $X=1.495
+ $Y=0.645 $X2=1.635 $Y2=0.905
.ends

.subckt PM_SKY130_FD_SC_LP__EINVP_M%VGND 1 4 9 11 12 13 20 21
r31 20 21 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r32 16 17 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r33 13 21 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=0.96 $Y=0 $X2=1.68
+ $Y2=0
r34 13 17 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=0.96 $Y=0 $X2=0.72
+ $Y2=0
r35 11 16 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.985 $Y=0 $X2=0.72
+ $Y2=0
r36 11 12 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.985 $Y=0 $X2=1.07
+ $Y2=0
r37 10 20 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=1.155 $Y=0 $X2=1.68
+ $Y2=0
r38 10 12 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.155 $Y=0 $X2=1.07
+ $Y2=0
r39 8 12 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.07 $Y=0.085 $X2=1.07
+ $Y2=0
r40 8 9 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=1.07 $Y=0.085
+ $X2=1.07 $Y2=0.82
r41 4 9 6.91519 $w=2.1e-07 $l=1.41244e-07 $layer=LI1_cond $X=0.985 $Y=0.925
+ $X2=1.07 $Y2=0.82
r42 4 6 7.39394 $w=2.08e-07 $l=1.4e-07 $layer=LI1_cond $X=0.985 $Y=0.925
+ $X2=0.845 $Y2=0.925
r43 1 6 182 $w=1.7e-07 $l=3.74166e-07 $layer=licon1_NDIFF $count=1 $X=0.625
+ $Y=0.645 $X2=0.845 $Y2=0.925
.ends

