* File: sky130_fd_sc_lp__sdfrbp_2.pex.spice
* Created: Wed Sep  2 10:34:13 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__SDFRBP_2%SCE 3 6 7 9 10 12 14 17 19 20 23 25 26 29
+ 30 38 44 50 52
c88 26 0 9.66853e-20 $X=2.35 $Y=1.23
c89 3 0 1.84245e-19 $X=0.475 $Y=0.615
r90 44 50 0.69845 $w=3.28e-07 $l=2e-08 $layer=LI1_cond $X=1.18 $Y=1.68 $X2=1.2
+ $Y2=1.68
r91 36 38 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=0.93 $Y=1.68
+ $X2=1.14 $Y2=1.68
r92 34 36 79.5619 $w=3.3e-07 $l=4.55e-07 $layer=POLY_cond $X=0.475 $Y=1.68
+ $X2=0.93 $Y2=1.68
r93 30 52 6.64621 $w=3.28e-07 $l=1.13e-07 $layer=LI1_cond $X=1.232 $Y=1.68
+ $X2=1.345 $Y2=1.68
r94 30 50 1.11752 $w=3.28e-07 $l=3.2e-08 $layer=LI1_cond $X=1.232 $Y=1.68
+ $X2=1.2 $Y2=1.68
r95 30 44 1.3969 $w=3.28e-07 $l=4e-08 $layer=LI1_cond $X=1.14 $Y=1.68 $X2=1.18
+ $Y2=1.68
r96 30 38 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.14
+ $Y=1.68 $X2=1.14 $Y2=1.68
r97 29 30 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=0.72 $Y=1.68
+ $X2=1.14 $Y2=1.68
r98 26 42 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.35 $Y=1.23
+ $X2=2.35 $Y2=1.065
r99 25 28 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=2.35 $Y=1.23
+ $X2=2.35 $Y2=1.395
r100 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.35
+ $Y=1.23 $X2=2.35 $Y2=1.23
r101 23 28 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=2.27 $Y=1.675
+ $X2=2.27 $Y2=1.395
r102 20 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.185 $Y=1.76
+ $X2=2.27 $Y2=1.675
r103 20 52 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=2.185 $Y=1.76
+ $X2=1.345 $Y2=1.76
r104 17 42 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=2.355 $Y=0.615
+ $X2=2.355 $Y2=1.065
r105 12 14 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=1.36 $Y=2.335
+ $X2=1.36 $Y2=2.765
r106 11 19 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.005 $Y=2.26
+ $X2=0.93 $Y2=2.26
r107 10 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.285 $Y=2.26
+ $X2=1.36 $Y2=2.335
r108 10 11 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=1.285 $Y=2.26
+ $X2=1.005 $Y2=2.26
r109 7 19 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.93 $Y=2.335
+ $X2=0.93 $Y2=2.26
r110 7 9 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=0.93 $Y=2.335
+ $X2=0.93 $Y2=2.765
r111 6 19 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.93 $Y=2.185
+ $X2=0.93 $Y2=2.26
r112 5 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.93 $Y=1.845
+ $X2=0.93 $Y2=1.68
r113 5 6 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=0.93 $Y=1.845 $X2=0.93
+ $Y2=2.185
r114 1 34 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=1.515
+ $X2=0.475 $Y2=1.68
r115 1 3 461.489 $w=1.5e-07 $l=9e-07 $layer=POLY_cond $X=0.475 $Y=1.515
+ $X2=0.475 $Y2=0.615
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRBP_2%A_27_81# 1 2 8 9 10 11 13 16 20 23 26 27 31
+ 33 35 36 38
c86 35 0 9.66853e-20 $X=2.17 $Y=2.11
r87 36 47 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.17 $Y=2.11
+ $X2=2.17 $Y2=2.275
r88 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.17
+ $Y=2.11 $X2=2.17 $Y2=2.11
r89 33 35 59.4661 $w=2.48e-07 $l=1.29e-06 $layer=LI1_cond $X=0.88 $Y=2.14
+ $X2=2.17 $Y2=2.14
r90 29 33 8.87234 $w=2.5e-07 $l=1.75e-07 $layer=LI1_cond $X=0.705 $Y=2.14
+ $X2=0.88 $Y2=2.14
r91 29 31 10.7013 $w=3.48e-07 $l=3.25e-07 $layer=LI1_cond $X=0.705 $Y=2.265
+ $X2=0.705 $Y2=2.59
r92 27 41 14.5135 $w=3.3e-07 $l=8.3e-08 $layer=POLY_cond $X=1.09 $Y=1.1
+ $X2=1.007 $Y2=1.1
r93 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.09
+ $Y=1.1 $X2=1.09 $Y2=1.1
r94 24 38 0.565906 $w=3.3e-07 $l=1.35e-07 $layer=LI1_cond $X=0.365 $Y=1.1
+ $X2=0.23 $Y2=1.1
r95 24 26 25.3188 $w=3.28e-07 $l=7.25e-07 $layer=LI1_cond $X=0.365 $Y=1.1
+ $X2=1.09 $Y2=1.1
r96 23 29 27.4645 $w=2.11e-07 $l=4.75e-07 $layer=LI1_cond $X=0.23 $Y=2.14
+ $X2=0.705 $Y2=2.14
r97 22 38 6.17543 $w=2.65e-07 $l=1.65e-07 $layer=LI1_cond $X=0.23 $Y=1.265
+ $X2=0.23 $Y2=1.1
r98 22 23 32.0123 $w=2.68e-07 $l=7.5e-07 $layer=LI1_cond $X=0.23 $Y=1.265
+ $X2=0.23 $Y2=2.015
r99 18 38 6.17543 $w=2.65e-07 $l=1.67481e-07 $layer=LI1_cond $X=0.225 $Y=0.935
+ $X2=0.23 $Y2=1.1
r100 18 20 13.519 $w=2.58e-07 $l=3.05e-07 $layer=LI1_cond $X=0.225 $Y=0.935
+ $X2=0.225 $Y2=0.63
r101 16 47 251.255 $w=1.5e-07 $l=4.9e-07 $layer=POLY_cond $X=2.15 $Y=2.765
+ $X2=2.15 $Y2=2.275
r102 11 13 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.54 $Y=0.295
+ $X2=1.54 $Y2=0.615
r103 9 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.465 $Y=0.22
+ $X2=1.54 $Y2=0.295
r104 9 10 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=1.465 $Y=0.22
+ $X2=1.125 $Y2=0.22
r105 8 41 10.8439 $w=2.35e-07 $l=1.65e-07 $layer=POLY_cond $X=1.007 $Y=0.935
+ $X2=1.007 $Y2=1.1
r106 7 10 28.6741 $w=1.5e-07 $l=1.50911e-07 $layer=POLY_cond $X=1.007 $Y=0.295
+ $X2=1.125 $Y2=0.22
r107 7 8 169.16 $w=2.35e-07 $l=6.4e-07 $layer=POLY_cond $X=1.007 $Y=0.295
+ $X2=1.007 $Y2=0.935
r108 2 31 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.59
+ $Y=2.445 $X2=0.715 $Y2=2.59
r109 1 20 182 $w=1.7e-07 $l=2.80624e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.405 $X2=0.26 $Y2=0.63
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRBP_2%D 3 7 9 10 16
r43 14 16 1.67361 $w=2.88e-07 $l=1e-08 $layer=POLY_cond $X=1.71 $Y=1.33 $X2=1.72
+ $Y2=1.33
r44 10 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.71
+ $Y=1.33 $X2=1.71 $Y2=1.33
r45 9 10 18.1448 $w=2.33e-07 $l=3.7e-07 $layer=LI1_cond $X=1.687 $Y=0.925
+ $X2=1.687 $Y2=1.295
r46 5 16 30.125 $w=2.88e-07 $l=2.49199e-07 $layer=POLY_cond $X=1.9 $Y=1.165
+ $X2=1.72 $Y2=1.33
r47 5 7 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=1.9 $Y=1.165 $X2=1.9
+ $Y2=0.615
r48 1 16 18.0107 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.72 $Y=1.495
+ $X2=1.72 $Y2=1.33
r49 1 3 651.213 $w=1.5e-07 $l=1.27e-06 $layer=POLY_cond $X=1.72 $Y=1.495
+ $X2=1.72 $Y2=2.765
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRBP_2%SCD 3 7 11 12 13 14 18
c44 7 0 1.81067e-19 $X=2.8 $Y=0.615
r45 18 19 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.71
+ $Y=1.77 $X2=2.71 $Y2=1.77
r46 14 19 10.9071 $w=2.78e-07 $l=2.65e-07 $layer=LI1_cond $X=2.665 $Y=2.035
+ $X2=2.665 $Y2=1.77
r47 13 19 4.32166 $w=2.78e-07 $l=1.05e-07 $layer=LI1_cond $X=2.665 $Y=1.665
+ $X2=2.665 $Y2=1.77
r48 11 18 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.71 $Y=2.11
+ $X2=2.71 $Y2=1.77
r49 11 12 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.71 $Y=2.11
+ $X2=2.71 $Y2=2.275
r50 10 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.71 $Y=1.605
+ $X2=2.71 $Y2=1.77
r51 7 10 507.638 $w=1.5e-07 $l=9.9e-07 $layer=POLY_cond $X=2.8 $Y=0.615 $X2=2.8
+ $Y2=1.605
r52 3 12 251.255 $w=1.5e-07 $l=4.9e-07 $layer=POLY_cond $X=2.62 $Y=2.765
+ $X2=2.62 $Y2=2.275
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRBP_2%CLK 1 3 4 6 9 11 13 25
c53 25 0 1.94544e-19 $X=4.165 $Y=1.35
c54 9 0 1.42869e-19 $X=4.165 $Y=2.465
c55 4 0 8.81973e-20 $X=4.15 $Y=1.09
r56 24 25 1.54335 $w=5.2e-07 $l=1.5e-08 $layer=POLY_cond $X=4.15 $Y=1.35
+ $X2=4.165 $Y2=1.35
r57 22 24 15.4335 $w=5.2e-07 $l=1.5e-07 $layer=POLY_cond $X=4 $Y=1.35 $X2=4.15
+ $Y2=1.35
r58 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4 $Y=1.445
+ $X2=4 $Y2=1.445
r59 19 22 28.8093 $w=5.2e-07 $l=2.8e-07 $layer=POLY_cond $X=3.72 $Y=1.35 $X2=4
+ $Y2=1.35
r60 13 23 1.77197 $w=5.38e-07 $l=8e-08 $layer=LI1_cond $X=4.08 $Y=1.48 $X2=4
+ $Y2=1.48
r61 11 23 8.85984 $w=5.38e-07 $l=4e-07 $layer=LI1_cond $X=3.6 $Y=1.48 $X2=4
+ $Y2=1.48
r62 7 25 32.4018 $w=1.5e-07 $l=2.6e-07 $layer=POLY_cond $X=4.165 $Y=1.61
+ $X2=4.165 $Y2=1.35
r63 7 9 438.415 $w=1.5e-07 $l=8.55e-07 $layer=POLY_cond $X=4.165 $Y=1.61
+ $X2=4.165 $Y2=2.465
r64 4 24 32.4018 $w=1.5e-07 $l=2.6e-07 $layer=POLY_cond $X=4.15 $Y=1.09 $X2=4.15
+ $Y2=1.35
r65 4 6 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=4.15 $Y=1.09 $X2=4.15
+ $Y2=0.805
r66 1 19 32.4018 $w=1.5e-07 $l=2.6e-07 $layer=POLY_cond $X=3.72 $Y=1.09 $X2=3.72
+ $Y2=1.35
r67 1 3 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.72 $Y=1.09 $X2=3.72
+ $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRBP_2%A_934_367# 1 2 9 11 15 19 22 25 27 31 32 34
+ 35 36 40 41 42 43 45 50 53 57 59
c187 59 0 1.37841e-19 $X=8.87 $Y=1.09
c188 57 0 1.77925e-19 $X=5.81 $Y=1.615
c189 41 0 1.71577e-19 $X=8.87 $Y=1.255
c190 40 0 1.19898e-19 $X=8.87 $Y=1.255
c191 11 0 1.67327e-19 $X=6.42 $Y=1.525
r192 56 57 30.474 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=5.735 $Y=1.615
+ $X2=5.81 $Y2=1.615
r193 53 63 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=9.44 $Y=2.155
+ $X2=9.44 $Y2=2.32
r194 52 53 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.44
+ $Y=2.155 $X2=9.44 $Y2=2.155
r195 50 52 15.3582 $w=2.82e-07 $l=3.55e-07 $layer=LI1_cond $X=9.435 $Y=1.8
+ $X2=9.435 $Y2=2.155
r196 46 56 34.9723 $w=3.3e-07 $l=2e-07 $layer=POLY_cond $X=5.535 $Y=1.615
+ $X2=5.735 $Y2=1.615
r197 45 48 10.1667 $w=6.42e-07 $l=7.13667e-07 $layer=LI1_cond $X=5.227 $Y=1.615
+ $X2=4.81 $Y2=2.15
r198 45 46 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.535
+ $Y=1.615 $X2=5.535 $Y2=1.615
r199 42 50 2.75002 $w=2e-07 $l=1.6e-07 $layer=LI1_cond $X=9.275 $Y=1.8 $X2=9.435
+ $Y2=1.8
r200 42 43 11.3682 $w=1.98e-07 $l=2.05e-07 $layer=LI1_cond $X=9.275 $Y=1.8
+ $X2=9.07 $Y2=1.8
r201 41 59 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.87 $Y=1.255
+ $X2=8.87 $Y2=1.09
r202 40 41 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.87
+ $Y=1.255 $X2=8.87 $Y2=1.255
r203 38 43 7.42997 $w=2e-07 $l=2.14243e-07 $layer=LI1_cond $X=8.9 $Y=1.7
+ $X2=9.07 $Y2=1.8
r204 38 40 15.0834 $w=3.38e-07 $l=4.45e-07 $layer=LI1_cond $X=8.9 $Y=1.7 $X2=8.9
+ $Y2=1.255
r205 37 40 9.82966 $w=3.38e-07 $l=2.9e-07 $layer=LI1_cond $X=8.9 $Y=0.965
+ $X2=8.9 $Y2=1.255
r206 35 37 14.8046 $w=1.92e-07 $l=2.4781e-07 $layer=LI1_cond $X=8.67 $Y=0.805
+ $X2=8.9 $Y2=0.842
r207 35 36 81.2246 $w=1.68e-07 $l=1.245e-06 $layer=LI1_cond $X=8.67 $Y=0.805
+ $X2=7.425 $Y2=0.805
r208 34 36 6.82373 $w=1.7e-07 $l=1.25499e-07 $layer=LI1_cond $X=7.335 $Y=0.72
+ $X2=7.425 $Y2=0.805
r209 33 34 14.7879 $w=1.78e-07 $l=2.4e-07 $layer=LI1_cond $X=7.335 $Y=0.48
+ $X2=7.335 $Y2=0.72
r210 31 33 6.82373 $w=1.7e-07 $l=1.25499e-07 $layer=LI1_cond $X=7.245 $Y=0.395
+ $X2=7.335 $Y2=0.48
r211 31 32 96.2299 $w=1.68e-07 $l=1.475e-06 $layer=LI1_cond $X=7.245 $Y=0.395
+ $X2=5.77 $Y2=0.395
r212 29 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.685 $Y=0.48
+ $X2=5.77 $Y2=0.395
r213 25 45 17.7646 $w=6.42e-07 $l=7.34112e-07 $layer=LI1_cond $X=5.685 $Y=1.075
+ $X2=5.227 $Y2=1.615
r214 25 29 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=5.685 $Y=1.075
+ $X2=5.685 $Y2=0.48
r215 25 27 9.54367 $w=3.18e-07 $l=2.65e-07 $layer=LI1_cond $X=4.93 $Y=1.05
+ $X2=4.93 $Y2=0.785
r216 22 63 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=9.35 $Y=2.69
+ $X2=9.35 $Y2=2.32
r217 19 59 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=8.82 $Y=0.66
+ $X2=8.82 $Y2=1.09
r218 13 24 6.7465 $w=1.5e-07 $l=1.02e-07 $layer=POLY_cond $X=6.67 $Y=1.395
+ $X2=6.67 $Y2=1.497
r219 13 15 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=6.67 $Y=1.395
+ $X2=6.67 $Y2=0.805
r220 11 24 69.3397 $w=1.77e-07 $l=2.63629e-07 $layer=POLY_cond $X=6.42 $Y=1.525
+ $X2=6.67 $Y2=1.497
r221 11 57 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=6.42 $Y=1.525
+ $X2=5.81 $Y2=1.525
r222 7 56 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.735 $Y=1.78
+ $X2=5.735 $Y2=1.615
r223 7 9 382.011 $w=1.5e-07 $l=7.45e-07 $layer=POLY_cond $X=5.735 $Y=1.78
+ $X2=5.735 $Y2=2.525
r224 2 48 600 $w=1.7e-07 $l=3.78583e-07 $layer=licon1_PDIFF $count=1 $X=4.67
+ $Y=1.835 $X2=4.81 $Y2=2.15
r225 1 27 182 $w=1.7e-07 $l=2.504e-07 $layer=licon1_NDIFF $count=1 $X=4.775
+ $Y=0.595 $X2=4.915 $Y2=0.785
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRBP_2%A_1290_365# 1 2 9 13 17 18 20 21 22 24 26
+ 30
c77 22 0 1.37841e-19 $X=8.435 $Y=1.235
c78 21 0 1.66848e-19 $X=6.79 $Y=1.147
c79 17 0 1.24056e-20 $X=6.705 $Y=1.99
r80 24 30 6.3449 $w=3.18e-07 $l=1.6e-07 $layer=LI1_cond $X=8.47 $Y=2.24 $X2=8.47
+ $Y2=2.08
r81 24 26 1.08042 $w=3.18e-07 $l=3e-08 $layer=LI1_cond $X=8.47 $Y=2.24 $X2=8.47
+ $Y2=2.27
r82 22 29 2.93179 $w=2.5e-07 $l=8.8e-08 $layer=LI1_cond $X=8.435 $Y=1.235
+ $X2=8.435 $Y2=1.147
r83 22 30 38.9526 $w=2.48e-07 $l=8.45e-07 $layer=LI1_cond $X=8.435 $Y=1.235
+ $X2=8.435 $Y2=2.08
r84 20 29 4.16448 $w=1.75e-07 $l=1.25e-07 $layer=LI1_cond $X=8.31 $Y=1.147
+ $X2=8.435 $Y2=1.147
r85 20 21 96.3325 $w=1.73e-07 $l=1.52e-06 $layer=LI1_cond $X=8.31 $Y=1.147
+ $X2=6.79 $Y2=1.147
r86 18 31 27.9871 $w=3.1e-07 $l=1.8e-07 $layer=POLY_cond $X=6.705 $Y=1.917
+ $X2=6.525 $Y2=1.917
r87 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.705
+ $Y=1.99 $X2=6.705 $Y2=1.99
r88 15 21 6.81835 $w=1.75e-07 $l=1.23386e-07 $layer=LI1_cond $X=6.705 $Y=1.235
+ $X2=6.79 $Y2=1.147
r89 15 17 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=6.705 $Y=1.235
+ $X2=6.705 $Y2=1.99
r90 11 18 50.5323 $w=3.1e-07 $l=4.27376e-07 $layer=POLY_cond $X=7.03 $Y=1.68
+ $X2=6.705 $Y2=1.917
r91 11 13 448.67 $w=1.5e-07 $l=8.75e-07 $layer=POLY_cond $X=7.03 $Y=1.68
+ $X2=7.03 $Y2=0.805
r92 7 31 19.7411 $w=1.5e-07 $l=2.38e-07 $layer=POLY_cond $X=6.525 $Y=2.155
+ $X2=6.525 $Y2=1.917
r93 7 9 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=6.525 $Y=2.155
+ $X2=6.525 $Y2=2.525
r94 2 26 300 $w=1.7e-07 $l=4.3946e-07 $layer=licon1_PDIFF $count=2 $X=8.275
+ $Y=1.895 $X2=8.415 $Y2=2.27
r95 1 29 182 $w=1.7e-07 $l=9.08364e-07 $layer=licon1_NDIFF $count=1 $X=8.175
+ $Y=0.34 $X2=8.395 $Y2=1.145
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRBP_2%RESET_B 3 8 9 10 11 13 17 20 24 26 27 28 29
+ 36 37 43 44 47 56 65
c205 47 0 7.96132e-21 $X=7.39 $Y=2.03
c206 44 0 3.22223e-19 $X=3.49 $Y=2.035
c207 28 0 1.97958e-19 $X=10.145 $Y=2.035
c208 27 0 1.42869e-19 $X=3.745 $Y=2.035
c209 20 0 1.47958e-19 $X=10.26 $Y=0.55
c210 8 0 1.07392e-19 $X=3.23 $Y=0.615
r211 54 56 30.6007 $w=3.3e-07 $l=1.75e-07 $layer=POLY_cond $X=10.34 $Y=2.155
+ $X2=10.515 $Y2=2.155
r212 54 65 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.34
+ $Y=2.155 $X2=10.34 $Y2=2.155
r213 51 54 13.9889 $w=3.3e-07 $l=8e-08 $layer=POLY_cond $X=10.26 $Y=2.155
+ $X2=10.34 $Y2=2.155
r214 47 49 15.3016 $w=3.15e-07 $l=1e-07 $layer=POLY_cond $X=7.39 $Y=2.03
+ $X2=7.49 $Y2=2.03
r215 43 44 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.49
+ $Y=2.035 $X2=3.49 $Y2=2.035
r216 41 43 45.4639 $w=3.3e-07 $l=2.6e-07 $layer=POLY_cond $X=3.23 $Y=2.035
+ $X2=3.49 $Y2=2.035
r217 39 41 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=3.16 $Y=2.035
+ $X2=3.23 $Y2=2.035
r218 37 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.29 $Y=2.035
+ $X2=10.29 $Y2=2.035
r219 36 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.49
+ $Y=1.99 $X2=7.49 $Y2=1.99
r220 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=2.035
+ $X2=7.44 $Y2=2.035
r221 31 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=2.035
+ $X2=3.6 $Y2=2.035
r222 29 35 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.585 $Y=2.035
+ $X2=7.44 $Y2=2.035
r223 28 37 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=10.145 $Y=2.035
+ $X2=10.29 $Y2=2.035
r224 28 29 3.16831 $w=1.4e-07 $l=2.56e-06 $layer=MET1_cond $X=10.145 $Y=2.035
+ $X2=7.585 $Y2=2.035
r225 27 31 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.745 $Y=2.035
+ $X2=3.6 $Y2=2.035
r226 26 35 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.295 $Y=2.035
+ $X2=7.44 $Y2=2.035
r227 26 27 4.39356 $w=1.4e-07 $l=3.55e-06 $layer=MET1_cond $X=7.295 $Y=2.035
+ $X2=3.745 $Y2=2.035
r228 22 56 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.515 $Y=2.32
+ $X2=10.515 $Y2=2.155
r229 22 24 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=10.515 $Y=2.32
+ $X2=10.515 $Y2=2.69
r230 18 51 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.26 $Y=1.99
+ $X2=10.26 $Y2=2.155
r231 18 20 738.383 $w=1.5e-07 $l=1.44e-06 $layer=POLY_cond $X=10.26 $Y=1.99
+ $X2=10.26 $Y2=0.55
r232 15 47 20.1192 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=7.39 $Y=1.82
+ $X2=7.39 $Y2=2.03
r233 15 17 520.457 $w=1.5e-07 $l=1.015e-06 $layer=POLY_cond $X=7.39 $Y=1.82
+ $X2=7.39 $Y2=0.805
r234 14 17 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=7.39 $Y=0.255
+ $X2=7.39 $Y2=0.805
r235 11 47 31.3683 $w=3.15e-07 $l=2.95212e-07 $layer=POLY_cond $X=7.185 $Y=2.24
+ $X2=7.39 $Y2=2.03
r236 11 13 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=7.185 $Y=2.24
+ $X2=7.185 $Y2=2.525
r237 9 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.315 $Y=0.18
+ $X2=7.39 $Y2=0.255
r238 9 10 2056.19 $w=1.5e-07 $l=4.01e-06 $layer=POLY_cond $X=7.315 $Y=0.18
+ $X2=3.305 $Y2=0.18
r239 6 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.23 $Y=1.87
+ $X2=3.23 $Y2=2.035
r240 6 8 643.521 $w=1.5e-07 $l=1.255e-06 $layer=POLY_cond $X=3.23 $Y=1.87
+ $X2=3.23 $Y2=0.615
r241 5 10 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.23 $Y=0.255
+ $X2=3.305 $Y2=0.18
r242 5 8 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=3.23 $Y=0.255
+ $X2=3.23 $Y2=0.615
r243 1 39 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.16 $Y=2.2
+ $X2=3.16 $Y2=2.035
r244 1 3 289.713 $w=1.5e-07 $l=5.65e-07 $layer=POLY_cond $X=3.16 $Y=2.2 $X2=3.16
+ $Y2=2.765
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRBP_2%A_1162_463# 1 2 3 12 16 18 23 24 27 29 33
+ 35 40 41 42
c113 29 0 1.67327e-19 $X=7.13 $Y=1.525
c114 27 0 8.72856e-20 $X=7.045 $Y=2.335
c115 18 0 1.69168e-19 $X=6.28 $Y=2.492
r116 41 46 45.456 $w=3.9e-07 $l=1.65e-07 $layer=POLY_cond $X=8.08 $Y=1.57
+ $X2=8.08 $Y2=1.735
r117 41 45 45.456 $w=3.9e-07 $l=1.65e-07 $layer=POLY_cond $X=8.08 $Y=1.57
+ $X2=8.08 $Y2=1.405
r118 40 42 3.84614 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=8.05 $Y=1.57
+ $X2=7.965 $Y2=1.57
r119 40 41 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.05
+ $Y=1.57 $X2=8.05 $Y2=1.57
r120 30 33 4.32166 $w=2.38e-07 $l=9e-08 $layer=LI1_cond $X=6.365 $Y=0.77
+ $X2=6.455 $Y2=0.77
r121 29 42 40.0954 $w=2.38e-07 $l=8.35e-07 $layer=LI1_cond $X=7.13 $Y=1.525
+ $X2=7.965 $Y2=1.525
r122 27 38 15.0906 $w=2.87e-07 $l=4.35804e-07 $layer=LI1_cond $X=7.045 $Y=2.335
+ $X2=7.4 $Y2=2.515
r123 26 29 7.07814 $w=2.4e-07 $l=1.56844e-07 $layer=LI1_cond $X=7.045 $Y=1.645
+ $X2=7.13 $Y2=1.525
r124 26 27 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=7.045 $Y=1.645
+ $X2=7.045 $Y2=2.335
r125 25 35 3.27229 $w=2.87e-07 $l=2.97993e-07 $layer=LI1_cond $X=6.52 $Y=2.42
+ $X2=6.28 $Y2=2.29
r126 24 27 5.6243 $w=2.87e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.96 $Y=2.42
+ $X2=7.045 $Y2=2.335
r127 24 25 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=6.96 $Y=2.42
+ $X2=6.52 $Y2=2.42
r128 23 35 3.2872 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.365 $Y=2.29
+ $X2=6.28 $Y2=2.29
r129 22 30 2.75731 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=6.365 $Y=0.89
+ $X2=6.365 $Y2=0.77
r130 22 23 91.3369 $w=1.68e-07 $l=1.4e-06 $layer=LI1_cond $X=6.365 $Y=0.89
+ $X2=6.365 $Y2=2.29
r131 18 35 3.27229 $w=2.87e-07 $l=2.02e-07 $layer=LI1_cond $X=6.28 $Y=2.492
+ $X2=6.28 $Y2=2.29
r132 18 20 9.39028 $w=4.03e-07 $l=3.3e-07 $layer=LI1_cond $X=6.28 $Y=2.492
+ $X2=5.95 $Y2=2.492
r133 16 46 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=8.2 $Y=2.315
+ $X2=8.2 $Y2=1.735
r134 12 45 382.011 $w=1.5e-07 $l=7.45e-07 $layer=POLY_cond $X=8.1 $Y=0.66
+ $X2=8.1 $Y2=1.405
r135 3 38 600 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_PDIFF $count=1 $X=7.26
+ $Y=2.315 $X2=7.4 $Y2=2.53
r136 2 20 600 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_PDIFF $count=1 $X=5.81
+ $Y=2.315 $X2=5.95 $Y2=2.53
r137 1 33 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=6.315
+ $Y=0.595 $X2=6.455 $Y2=0.775
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRBP_2%A_759_119# 1 2 9 11 13 15 16 18 19 20 21 22
+ 25 27 29 30 35 36 37 40 42 43 45 48 50 52 56 64
c184 64 0 6.19004e-20 $X=4.685 $Y=1.445
c185 52 0 8.81973e-20 $X=3.935 $Y=0.82
c186 50 0 1.27679e-19 $X=4.43 $Y=1.93
c187 36 0 1.44931e-19 $X=9.245 $Y=1.705
c188 35 0 4.11935e-20 $X=8.775 $Y=2.48
c189 27 0 1.66848e-19 $X=6.24 $Y=1.09
c190 21 0 4.44429e-21 $X=6.165 $Y=1.165
c191 15 0 1.69168e-19 $X=5.085 $Y=3.075
r192 70 71 4.65451 $w=4.66e-07 $l=4.5e-08 $layer=POLY_cond $X=5.085 $Y=1.35
+ $X2=5.13 $Y2=1.35
r193 69 70 39.8219 $w=4.66e-07 $l=3.85e-07 $layer=POLY_cond $X=4.7 $Y=1.35
+ $X2=5.085 $Y2=1.35
r194 65 69 1.5515 $w=4.66e-07 $l=1.5e-08 $layer=POLY_cond $X=4.685 $Y=1.35
+ $X2=4.7 $Y2=1.35
r195 65 67 9.30901 $w=4.66e-07 $l=9e-08 $layer=POLY_cond $X=4.685 $Y=1.35
+ $X2=4.595 $Y2=1.35
r196 64 65 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.685
+ $Y=1.445 $X2=4.685 $Y2=1.445
r197 61 64 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=4.43 $Y=1.445
+ $X2=4.685 $Y2=1.445
r198 56 59 6.22319 $w=2.48e-07 $l=1.35e-07 $layer=LI1_cond $X=3.99 $Y=2.015
+ $X2=3.99 $Y2=2.15
r199 52 54 5.76222 $w=2.58e-07 $l=1.3e-07 $layer=LI1_cond $X=3.93 $Y=0.82
+ $X2=3.93 $Y2=0.95
r200 49 61 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.43 $Y=1.61
+ $X2=4.43 $Y2=1.445
r201 49 50 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=4.43 $Y=1.61
+ $X2=4.43 $Y2=1.93
r202 48 61 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.43 $Y=1.28
+ $X2=4.43 $Y2=1.445
r203 47 48 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=4.43 $Y=1.04
+ $X2=4.43 $Y2=1.28
r204 46 56 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.115 $Y=2.015
+ $X2=3.99 $Y2=2.015
r205 45 50 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.345 $Y=2.015
+ $X2=4.43 $Y2=1.93
r206 45 46 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=4.345 $Y=2.015
+ $X2=4.115 $Y2=2.015
r207 44 54 2.89065 $w=1.8e-07 $l=1.3e-07 $layer=LI1_cond $X=4.06 $Y=0.95
+ $X2=3.93 $Y2=0.95
r208 43 47 6.82373 $w=1.8e-07 $l=1.25499e-07 $layer=LI1_cond $X=4.345 $Y=0.95
+ $X2=4.43 $Y2=1.04
r209 43 44 17.5606 $w=1.78e-07 $l=2.85e-07 $layer=LI1_cond $X=4.345 $Y=0.95
+ $X2=4.06 $Y2=0.95
r210 38 40 553.787 $w=1.5e-07 $l=1.08e-06 $layer=POLY_cond $X=9.32 $Y=1.63
+ $X2=9.32 $Y2=0.55
r211 36 38 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.245 $Y=1.705
+ $X2=9.32 $Y2=1.63
r212 36 37 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=9.245 $Y=1.705
+ $X2=8.85 $Y2=1.705
r213 33 35 305.096 $w=1.5e-07 $l=5.95e-07 $layer=POLY_cond $X=8.775 $Y=3.075
+ $X2=8.775 $Y2=2.48
r214 32 37 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.775 $Y=1.78
+ $X2=8.85 $Y2=1.705
r215 32 35 358.936 $w=1.5e-07 $l=7e-07 $layer=POLY_cond $X=8.775 $Y=1.78
+ $X2=8.775 $Y2=2.48
r216 31 42 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.24 $Y=3.15
+ $X2=6.165 $Y2=3.15
r217 30 33 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.7 $Y=3.15
+ $X2=8.775 $Y2=3.075
r218 30 31 1261.4 $w=1.5e-07 $l=2.46e-06 $layer=POLY_cond $X=8.7 $Y=3.15
+ $X2=6.24 $Y2=3.15
r219 27 29 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=6.24 $Y=1.09
+ $X2=6.24 $Y2=0.805
r220 23 42 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.165 $Y=3.075
+ $X2=6.165 $Y2=3.15
r221 23 25 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=6.165 $Y=3.075
+ $X2=6.165 $Y2=2.525
r222 22 71 31.7582 $w=4.66e-07 $l=2.19317e-07 $layer=POLY_cond $X=5.205 $Y=1.165
+ $X2=5.13 $Y2=1.35
r223 21 27 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.165 $Y=1.165
+ $X2=6.24 $Y2=1.09
r224 21 22 492.255 $w=1.5e-07 $l=9.6e-07 $layer=POLY_cond $X=6.165 $Y=1.165
+ $X2=5.205 $Y2=1.165
r225 19 42 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.09 $Y=3.15
+ $X2=6.165 $Y2=3.15
r226 19 20 476.872 $w=1.5e-07 $l=9.3e-07 $layer=POLY_cond $X=6.09 $Y=3.15
+ $X2=5.16 $Y2=3.15
r227 16 71 29.638 $w=1.5e-07 $l=2.6e-07 $layer=POLY_cond $X=5.13 $Y=1.09
+ $X2=5.13 $Y2=1.35
r228 16 18 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=5.13 $Y=1.09
+ $X2=5.13 $Y2=0.805
r229 15 20 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.085 $Y=3.075
+ $X2=5.16 $Y2=3.15
r230 14 70 29.638 $w=1.5e-07 $l=2.6e-07 $layer=POLY_cond $X=5.085 $Y=1.61
+ $X2=5.085 $Y2=1.35
r231 14 15 751.202 $w=1.5e-07 $l=1.465e-06 $layer=POLY_cond $X=5.085 $Y=1.61
+ $X2=5.085 $Y2=3.075
r232 11 69 29.638 $w=1.5e-07 $l=2.6e-07 $layer=POLY_cond $X=4.7 $Y=1.09 $X2=4.7
+ $Y2=1.35
r233 11 13 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=4.7 $Y=1.09 $X2=4.7
+ $Y2=0.805
r234 7 67 29.638 $w=1.5e-07 $l=2.6e-07 $layer=POLY_cond $X=4.595 $Y=1.61
+ $X2=4.595 $Y2=1.35
r235 7 9 438.415 $w=1.5e-07 $l=8.55e-07 $layer=POLY_cond $X=4.595 $Y=1.61
+ $X2=4.595 $Y2=2.465
r236 2 59 600 $w=1.7e-07 $l=3.7229e-07 $layer=licon1_PDIFF $count=1 $X=3.825
+ $Y=1.835 $X2=3.95 $Y2=2.15
r237 1 52 182 $w=1.7e-07 $l=2.86575e-07 $layer=licon1_NDIFF $count=1 $X=3.795
+ $Y=0.595 $X2=3.935 $Y2=0.82
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRBP_2%A_1923_174# 1 2 9 12 17 19 20 23 28 29 31
+ 32 34 38 41
c95 38 0 1.47958e-19 $X=11.15 $Y=2.025
c96 34 0 1.87138e-19 $X=10.835 $Y=1.06
c97 12 0 7.25196e-20 $X=9.89 $Y=2.69
r98 31 32 9.81945 $w=2.68e-07 $l=2.2e-07 $layer=LI1_cond $X=10.76 $Y=2.69
+ $X2=10.76 $Y2=2.47
r99 28 38 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.15 $Y=1.94
+ $X2=11.15 $Y2=2.025
r100 27 34 12.3173 $w=3.12e-07 $l=4.02772e-07 $layer=LI1_cond $X=11.15 $Y=1.26
+ $X2=10.835 $Y2=1.06
r101 27 28 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=11.15 $Y=1.26
+ $X2=11.15 $Y2=1.94
r102 25 38 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=10.785 $Y=2.025
+ $X2=11.15 $Y2=2.025
r103 25 32 18.8582 $w=2.18e-07 $l=3.6e-07 $layer=LI1_cond $X=10.785 $Y=2.11
+ $X2=10.785 $Y2=2.47
r104 21 34 0.37154 $w=3.3e-07 $l=2e-07 $layer=LI1_cond $X=10.835 $Y=0.86
+ $X2=10.835 $Y2=1.06
r105 21 23 10.826 $w=3.28e-07 $l=3.1e-07 $layer=LI1_cond $X=10.835 $Y=0.86
+ $X2=10.835 $Y2=0.55
r106 20 29 6.14925 $w=3.98e-07 $l=2e-07 $layer=LI1_cond $X=10.325 $Y=1.06
+ $X2=10.125 $Y2=1.06
r107 19 34 5.65586 $w=4e-07 $l=1.65e-07 $layer=LI1_cond $X=10.67 $Y=1.06
+ $X2=10.835 $Y2=1.06
r108 19 20 9.93982 $w=3.98e-07 $l=3.45e-07 $layer=LI1_cond $X=10.67 $Y=1.06
+ $X2=10.325 $Y2=1.06
r109 17 42 46.4315 $w=3.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.79 $Y=1.035
+ $X2=9.79 $Y2=1.2
r110 17 41 46.4315 $w=3.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.79 $Y=1.035
+ $X2=9.79 $Y2=0.87
r111 16 29 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=9.78 $Y=1.025
+ $X2=10.125 $Y2=1.025
r112 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.78
+ $Y=1.035 $X2=9.78 $Y2=1.035
r113 12 42 764.021 $w=1.5e-07 $l=1.49e-06 $layer=POLY_cond $X=9.89 $Y=2.69
+ $X2=9.89 $Y2=1.2
r114 9 41 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=9.83 $Y=0.55
+ $X2=9.83 $Y2=0.87
r115 2 31 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=10.59
+ $Y=2.48 $X2=10.73 $Y2=2.69
r116 1 23 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=10.695
+ $Y=0.34 $X2=10.835 $Y2=0.55
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRBP_2%A_1770_412# 1 2 9 13 15 19 23 25 29 33 35
+ 39 43 45 46 47 50 52 55 56 57 59 62 65 73 75 80
c188 73 0 6.20701e-20 $X=9.342 $Y=0.452
c189 65 0 7.25196e-20 $X=8.99 $Y=2.58
c190 59 0 5.43578e-20 $X=9.85 $Y=2.49
c191 57 0 9.05736e-20 $X=9.445 $Y=1.445
c192 52 0 4.11935e-20 $X=9.765 $Y=2.58
c193 50 0 1.40547e-20 $X=8.99 $Y=2.27
c194 29 0 8.72905e-20 $X=11.98 $Y=2.465
c195 2 0 1.02506e-19 $X=8.85 $Y=2.06
c196 1 0 1.19898e-19 $X=8.895 $Y=0.34
r197 79 80 33.1619 $w=4e-07 $l=7.5e-08 $layer=POLY_cond $X=10.945 $Y=1.58
+ $X2=11.02 $Y2=1.58
r198 71 73 6.91466 $w=3.93e-07 $l=2.37e-07 $layer=LI1_cond $X=9.105 $Y=0.452
+ $X2=9.342 $Y2=0.452
r199 65 68 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=8.99 $Y=2.58
+ $X2=8.99 $Y2=2.73
r200 65 66 3.44076 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=8.99 $Y=2.58 $X2=8.99
+ $Y2=2.49
r201 63 79 32.674 $w=4e-07 $l=2.35e-07 $layer=POLY_cond $X=10.71 $Y=1.58
+ $X2=10.945 $Y2=1.58
r202 63 76 12.5135 $w=4e-07 $l=9e-08 $layer=POLY_cond $X=10.71 $Y=1.58 $X2=10.62
+ $Y2=1.58
r203 62 63 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.71
+ $Y=1.595 $X2=10.71 $Y2=1.595
r204 60 75 3.70735 $w=2.5e-07 $l=1.11131e-07 $layer=LI1_cond $X=9.955 $Y=1.595
+ $X2=9.86 $Y2=1.56
r205 60 62 26.3665 $w=3.28e-07 $l=7.55e-07 $layer=LI1_cond $X=9.955 $Y=1.595
+ $X2=10.71 $Y2=1.595
r206 58 75 2.76166 $w=1.7e-07 $l=2.04939e-07 $layer=LI1_cond $X=9.85 $Y=1.76
+ $X2=9.86 $Y2=1.56
r207 58 59 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=9.85 $Y=1.76
+ $X2=9.85 $Y2=2.49
r208 56 75 3.70735 $w=2.5e-07 $l=1.55403e-07 $layer=LI1_cond $X=9.765 $Y=1.445
+ $X2=9.86 $Y2=1.56
r209 56 57 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=9.765 $Y=1.445
+ $X2=9.445 $Y2=1.445
r210 55 57 6.89401 $w=1.7e-07 $l=1.39155e-07 $layer=LI1_cond $X=9.342 $Y=1.36
+ $X2=9.445 $Y2=1.445
r211 54 73 4.5952 $w=2.05e-07 $l=1.98e-07 $layer=LI1_cond $X=9.342 $Y=0.65
+ $X2=9.342 $Y2=0.452
r212 54 55 38.4124 $w=2.03e-07 $l=7.1e-07 $layer=LI1_cond $X=9.342 $Y=0.65
+ $X2=9.342 $Y2=1.36
r213 53 65 4.28565 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=9.155 $Y=2.58
+ $X2=8.99 $Y2=2.58
r214 52 59 6.82373 $w=1.8e-07 $l=1.25499e-07 $layer=LI1_cond $X=9.765 $Y=2.58
+ $X2=9.85 $Y2=2.49
r215 52 53 37.5859 $w=1.78e-07 $l=6.1e-07 $layer=LI1_cond $X=9.765 $Y=2.58
+ $X2=9.155 $Y2=2.58
r216 50 66 9.05491 $w=2.78e-07 $l=2.2e-07 $layer=LI1_cond $X=8.965 $Y=2.27
+ $X2=8.965 $Y2=2.49
r217 41 47 20.4101 $w=1.5e-07 $l=7.98436e-08 $layer=POLY_cond $X=12.525 $Y=1.38
+ $X2=12.515 $Y2=1.455
r218 41 43 476.872 $w=1.5e-07 $l=9.3e-07 $layer=POLY_cond $X=12.525 $Y=1.38
+ $X2=12.525 $Y2=0.45
r219 37 47 20.4101 $w=1.5e-07 $l=7.98436e-08 $layer=POLY_cond $X=12.505 $Y=1.53
+ $X2=12.515 $Y2=1.455
r220 37 39 320.479 $w=1.5e-07 $l=6.25e-07 $layer=POLY_cond $X=12.505 $Y=1.53
+ $X2=12.505 $Y2=2.155
r221 36 46 12.05 $w=1.5e-07 $l=8.5e-08 $layer=POLY_cond $X=12.075 $Y=1.455
+ $X2=11.99 $Y2=1.455
r222 35 47 5.30422 $w=1.5e-07 $l=8.5e-08 $layer=POLY_cond $X=12.43 $Y=1.455
+ $X2=12.515 $Y2=1.455
r223 35 36 182.032 $w=1.5e-07 $l=3.55e-07 $layer=POLY_cond $X=12.43 $Y=1.455
+ $X2=12.075 $Y2=1.455
r224 31 46 12.05 $w=1.5e-07 $l=7.98436e-08 $layer=POLY_cond $X=12 $Y=1.38
+ $X2=11.99 $Y2=1.455
r225 31 33 369.191 $w=1.5e-07 $l=7.2e-07 $layer=POLY_cond $X=12 $Y=1.38 $X2=12
+ $Y2=0.66
r226 27 46 12.05 $w=1.5e-07 $l=7.98436e-08 $layer=POLY_cond $X=11.98 $Y=1.53
+ $X2=11.99 $Y2=1.455
r227 27 29 479.436 $w=1.5e-07 $l=9.35e-07 $layer=POLY_cond $X=11.98 $Y=1.53
+ $X2=11.98 $Y2=2.465
r228 26 45 12.05 $w=1.5e-07 $l=8.5e-08 $layer=POLY_cond $X=11.645 $Y=1.455
+ $X2=11.56 $Y2=1.455
r229 25 46 12.05 $w=1.5e-07 $l=8.5e-08 $layer=POLY_cond $X=11.905 $Y=1.455
+ $X2=11.99 $Y2=1.455
r230 25 26 133.319 $w=1.5e-07 $l=2.6e-07 $layer=POLY_cond $X=11.905 $Y=1.455
+ $X2=11.645 $Y2=1.455
r231 21 45 12.05 $w=1.5e-07 $l=7.98436e-08 $layer=POLY_cond $X=11.57 $Y=1.38
+ $X2=11.56 $Y2=1.455
r232 21 23 369.191 $w=1.5e-07 $l=7.2e-07 $layer=POLY_cond $X=11.57 $Y=1.38
+ $X2=11.57 $Y2=0.66
r233 17 45 12.05 $w=1.5e-07 $l=7.98436e-08 $layer=POLY_cond $X=11.55 $Y=1.53
+ $X2=11.56 $Y2=1.455
r234 17 19 479.436 $w=1.5e-07 $l=9.35e-07 $layer=POLY_cond $X=11.55 $Y=1.53
+ $X2=11.55 $Y2=2.465
r235 15 45 12.05 $w=1.5e-07 $l=8.5e-08 $layer=POLY_cond $X=11.475 $Y=1.455
+ $X2=11.56 $Y2=1.455
r236 15 80 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=11.475 $Y=1.455
+ $X2=11.02 $Y2=1.455
r237 11 79 25.8619 $w=1.5e-07 $l=2e-07 $layer=POLY_cond $X=10.945 $Y=1.78
+ $X2=10.945 $Y2=1.58
r238 11 13 466.617 $w=1.5e-07 $l=9.1e-07 $layer=POLY_cond $X=10.945 $Y=1.78
+ $X2=10.945 $Y2=2.69
r239 7 76 25.8619 $w=1.5e-07 $l=2e-07 $layer=POLY_cond $X=10.62 $Y=1.38
+ $X2=10.62 $Y2=1.58
r240 7 9 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=10.62 $Y=1.38
+ $X2=10.62 $Y2=0.55
r241 2 68 600 $w=1.7e-07 $l=7.36682e-07 $layer=licon1_PDIFF $count=1 $X=8.85
+ $Y=2.06 $X2=8.99 $Y2=2.73
r242 2 50 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=8.85
+ $Y=2.06 $X2=8.99 $Y2=2.27
r243 1 71 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=8.895
+ $Y=0.34 $X2=9.105 $Y2=0.485
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRBP_2%A_2516_367# 1 2 7 9 12 14 16 19 23 27 31 34
+ 38
c58 34 0 8.72905e-20 $X=12.74 $Y=1.395
r59 37 38 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=13.475 $Y=1.395
+ $X2=13.905 $Y2=1.395
r60 32 37 27.1035 $w=3.3e-07 $l=1.55e-07 $layer=POLY_cond $X=13.32 $Y=1.395
+ $X2=13.475 $Y2=1.395
r61 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=13.32
+ $Y=1.395 $X2=13.32 $Y2=1.395
r62 29 34 1.23199 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=12.905 $Y=1.395
+ $X2=12.74 $Y2=1.395
r63 29 31 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=12.905 $Y=1.395
+ $X2=13.32 $Y2=1.395
r64 25 34 5.29963 $w=3.2e-07 $l=1.69926e-07 $layer=LI1_cond $X=12.73 $Y=1.56
+ $X2=12.74 $Y2=1.395
r65 25 27 15.6137 $w=3.08e-07 $l=4.2e-07 $layer=LI1_cond $X=12.73 $Y=1.56
+ $X2=12.73 $Y2=1.98
r66 21 34 5.29963 $w=3.2e-07 $l=1.65e-07 $layer=LI1_cond $X=12.74 $Y=1.23
+ $X2=12.74 $Y2=1.395
r67 21 23 27.2396 $w=3.28e-07 $l=7.8e-07 $layer=LI1_cond $X=12.74 $Y=1.23
+ $X2=12.74 $Y2=0.45
r68 17 38 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=13.905 $Y=1.56
+ $X2=13.905 $Y2=1.395
r69 17 19 464.053 $w=1.5e-07 $l=9.05e-07 $layer=POLY_cond $X=13.905 $Y=1.56
+ $X2=13.905 $Y2=2.465
r70 14 38 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=13.905 $Y=1.23
+ $X2=13.905 $Y2=1.395
r71 14 16 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=13.905 $Y=1.23
+ $X2=13.905 $Y2=0.7
r72 10 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=13.475 $Y=1.56
+ $X2=13.475 $Y2=1.395
r73 10 12 464.053 $w=1.5e-07 $l=9.05e-07 $layer=POLY_cond $X=13.475 $Y=1.56
+ $X2=13.475 $Y2=2.465
r74 7 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=13.475 $Y=1.23
+ $X2=13.475 $Y2=1.395
r75 7 9 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=13.475 $Y=1.23
+ $X2=13.475 $Y2=0.7
r76 2 27 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=12.58
+ $Y=1.835 $X2=12.72 $Y2=1.98
r77 1 23 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=12.6
+ $Y=0.24 $X2=12.74 $Y2=0.45
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRBP_2%VPWR 1 2 3 4 5 6 7 8 9 10 33 37 41 45 49 53
+ 57 63 67 69 74 75 77 78 80 81 82 84 108 112 120 125 130 135 141 144 149 152
+ 155 158 162
r200 161 162 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.16 $Y=3.33
+ $X2=14.16 $Y2=3.33
r201 158 159 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.2 $Y=3.33
+ $X2=13.2 $Y2=3.33
r202 155 156 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.24 $Y=3.33
+ $X2=12.24 $Y2=3.33
r203 152 153 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.28 $Y=3.33
+ $X2=11.28 $Y2=3.33
r204 149 150 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.32 $Y=3.33
+ $X2=10.32 $Y2=3.33
r205 147 149 13.0133 $w=6e-07 $l=6.91896e-07 $layer=LI1_cond $X=10.19 $Y=2.69
+ $X2=10.082 $Y2=3.33
r206 144 145 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r207 141 142 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r208 139 162 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.68 $Y=3.33
+ $X2=14.16 $Y2=3.33
r209 139 159 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.68 $Y=3.33
+ $X2=13.2 $Y2=3.33
r210 138 139 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.68 $Y=3.33
+ $X2=13.68 $Y2=3.33
r211 136 158 8.23795 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=13.405 $Y=3.33
+ $X2=13.25 $Y2=3.33
r212 136 138 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=13.405 $Y=3.33
+ $X2=13.68 $Y2=3.33
r213 135 161 4.4964 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=13.98 $Y=3.33
+ $X2=14.19 $Y2=3.33
r214 135 138 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=13.98 $Y=3.33
+ $X2=13.68 $Y2=3.33
r215 134 159 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.72 $Y=3.33
+ $X2=13.2 $Y2=3.33
r216 134 156 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.72 $Y=3.33
+ $X2=12.24 $Y2=3.33
r217 133 134 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.72 $Y=3.33
+ $X2=12.72 $Y2=3.33
r218 131 155 8.42608 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=12.405 $Y=3.33
+ $X2=12.245 $Y2=3.33
r219 131 133 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=12.405 $Y=3.33
+ $X2=12.72 $Y2=3.33
r220 130 158 8.23795 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=13.095 $Y=3.33
+ $X2=13.25 $Y2=3.33
r221 130 133 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=13.095 $Y=3.33
+ $X2=12.72 $Y2=3.33
r222 129 156 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.76 $Y=3.33
+ $X2=12.24 $Y2=3.33
r223 129 153 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.76 $Y=3.33
+ $X2=11.28 $Y2=3.33
r224 128 129 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.76 $Y=3.33
+ $X2=11.76 $Y2=3.33
r225 126 152 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.48 $Y=3.33
+ $X2=11.315 $Y2=3.33
r226 126 128 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=11.48 $Y=3.33
+ $X2=11.76 $Y2=3.33
r227 125 155 8.42608 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=12.085 $Y=3.33
+ $X2=12.245 $Y2=3.33
r228 125 128 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=12.085 $Y=3.33
+ $X2=11.76 $Y2=3.33
r229 124 153 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.8 $Y=3.33
+ $X2=11.28 $Y2=3.33
r230 124 150 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.8 $Y=3.33
+ $X2=10.32 $Y2=3.33
r231 123 124 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=3.33
+ $X2=10.8 $Y2=3.33
r232 121 149 8.31678 $w=1.7e-07 $l=3.73e-07 $layer=LI1_cond $X=10.455 $Y=3.33
+ $X2=10.082 $Y2=3.33
r233 121 123 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=10.455 $Y=3.33
+ $X2=10.8 $Y2=3.33
r234 120 152 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.15 $Y=3.33
+ $X2=11.315 $Y2=3.33
r235 120 123 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=11.15 $Y=3.33
+ $X2=10.8 $Y2=3.33
r236 119 150 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=10.32 $Y2=3.33
r237 118 119 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r238 116 119 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=9.36 $Y2=3.33
r239 116 145 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=7.92 $Y2=3.33
r240 115 118 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=8.4 $Y=3.33
+ $X2=9.36 $Y2=3.33
r241 115 116 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r242 113 144 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.025 $Y=3.33
+ $X2=7.9 $Y2=3.33
r243 113 115 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=8.025 $Y=3.33
+ $X2=8.4 $Y2=3.33
r244 112 149 8.31678 $w=1.7e-07 $l=3.72e-07 $layer=LI1_cond $X=9.71 $Y=3.33
+ $X2=10.082 $Y2=3.33
r245 112 118 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=9.71 $Y=3.33
+ $X2=9.36 $Y2=3.33
r246 111 145 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=7.92 $Y2=3.33
r247 110 111 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r248 108 144 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.775 $Y=3.33
+ $X2=7.9 $Y2=3.33
r249 108 110 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=7.775 $Y=3.33
+ $X2=7.44 $Y2=3.33
r250 106 107 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r251 104 107 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=6.48 $Y2=3.33
r252 103 106 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=4.56 $Y=3.33
+ $X2=6.48 $Y2=3.33
r253 103 104 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r254 101 104 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r255 100 101 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r256 98 101 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=4.08 $Y2=3.33
r257 97 100 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=3.12 $Y=3.33
+ $X2=4.08 $Y2=3.33
r258 97 98 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r259 95 98 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r260 94 95 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r261 92 95 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r262 92 142 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r263 91 94 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r264 91 92 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r265 89 141 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.31 $Y=3.33
+ $X2=1.18 $Y2=3.33
r266 89 91 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=1.31 $Y=3.33
+ $X2=1.68 $Y2=3.33
r267 87 142 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r268 86 87 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r269 84 141 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.05 $Y=3.33
+ $X2=1.18 $Y2=3.33
r270 84 86 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=1.05 $Y=3.33
+ $X2=0.72 $Y2=3.33
r271 82 111 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=7.2 $Y=3.33
+ $X2=7.44 $Y2=3.33
r272 82 107 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=7.2 $Y=3.33
+ $X2=6.48 $Y2=3.33
r273 80 106 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=6.69 $Y=3.33
+ $X2=6.48 $Y2=3.33
r274 80 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.69 $Y=3.33
+ $X2=6.855 $Y2=3.33
r275 79 110 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=7.02 $Y=3.33
+ $X2=7.44 $Y2=3.33
r276 79 81 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.02 $Y=3.33
+ $X2=6.855 $Y2=3.33
r277 77 100 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=4.215 $Y=3.33
+ $X2=4.08 $Y2=3.33
r278 77 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.215 $Y=3.33
+ $X2=4.38 $Y2=3.33
r279 76 103 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=4.545 $Y=3.33
+ $X2=4.56 $Y2=3.33
r280 76 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.545 $Y=3.33
+ $X2=4.38 $Y2=3.33
r281 74 94 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=2.67 $Y=3.33 $X2=2.64
+ $Y2=3.33
r282 74 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.67 $Y=3.33
+ $X2=2.835 $Y2=3.33
r283 73 97 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=3 $Y=3.33 $X2=3.12
+ $Y2=3.33
r284 73 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3 $Y=3.33 $X2=2.835
+ $Y2=3.33
r285 69 72 36.6515 $w=3.03e-07 $l=9.7e-07 $layer=LI1_cond $X=14.132 $Y=1.98
+ $X2=14.132 $Y2=2.95
r286 67 161 3.06184 $w=3.05e-07 $l=1.1025e-07 $layer=LI1_cond $X=14.132 $Y=3.245
+ $X2=14.19 $Y2=3.33
r287 67 72 11.1466 $w=3.03e-07 $l=2.95e-07 $layer=LI1_cond $X=14.132 $Y=3.245
+ $X2=14.132 $Y2=2.95
r288 63 66 36.0603 $w=3.08e-07 $l=9.7e-07 $layer=LI1_cond $X=13.25 $Y=1.98
+ $X2=13.25 $Y2=2.95
r289 61 158 0.701276 $w=3.1e-07 $l=8.5e-08 $layer=LI1_cond $X=13.25 $Y=3.245
+ $X2=13.25 $Y2=3.33
r290 61 66 10.9668 $w=3.08e-07 $l=2.95e-07 $layer=LI1_cond $X=13.25 $Y=3.245
+ $X2=13.25 $Y2=2.95
r291 57 60 18.0069 $w=3.18e-07 $l=5e-07 $layer=LI1_cond $X=12.245 $Y=1.96
+ $X2=12.245 $Y2=2.46
r292 55 155 0.800721 $w=3.2e-07 $l=8.5e-08 $layer=LI1_cond $X=12.245 $Y=3.245
+ $X2=12.245 $Y2=3.33
r293 55 60 28.2709 $w=3.18e-07 $l=7.85e-07 $layer=LI1_cond $X=12.245 $Y=3.245
+ $X2=12.245 $Y2=2.46
r294 51 152 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=11.315 $Y=3.245
+ $X2=11.315 $Y2=3.33
r295 51 53 30.7318 $w=3.28e-07 $l=8.8e-07 $layer=LI1_cond $X=11.315 $Y=3.245
+ $X2=11.315 $Y2=2.365
r296 47 144 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.9 $Y=3.245
+ $X2=7.9 $Y2=3.33
r297 47 49 45.8672 $w=2.48e-07 $l=9.95e-07 $layer=LI1_cond $X=7.9 $Y=3.245
+ $X2=7.9 $Y2=2.25
r298 43 81 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.855 $Y=3.245
+ $X2=6.855 $Y2=3.33
r299 43 45 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=6.855 $Y=3.245
+ $X2=6.855 $Y2=2.765
r300 39 78 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.38 $Y=3.245
+ $X2=4.38 $Y2=3.33
r301 39 41 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=4.38 $Y=3.245
+ $X2=4.38 $Y2=2.93
r302 35 75 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.835 $Y=3.245
+ $X2=2.835 $Y2=3.33
r303 35 37 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=2.835 $Y=3.245
+ $X2=2.835 $Y2=2.94
r304 31 141 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=1.18 $Y=3.245
+ $X2=1.18 $Y2=3.33
r305 31 33 28.5895 $w=2.58e-07 $l=6.45e-07 $layer=LI1_cond $X=1.18 $Y=3.245
+ $X2=1.18 $Y2=2.6
r306 10 72 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=13.98
+ $Y=1.835 $X2=14.12 $Y2=2.95
r307 10 69 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=13.98
+ $Y=1.835 $X2=14.12 $Y2=1.98
r308 9 66 400 $w=1.7e-07 $l=1.17584e-06 $layer=licon1_PDIFF $count=1 $X=13.135
+ $Y=1.835 $X2=13.26 $Y2=2.95
r309 9 63 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=13.135
+ $Y=1.835 $X2=13.26 $Y2=1.98
r310 8 60 300 $w=1.7e-07 $l=6.91466e-07 $layer=licon1_PDIFF $count=2 $X=12.055
+ $Y=1.835 $X2=12.195 $Y2=2.46
r311 8 57 600 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_PDIFF $count=1 $X=12.055
+ $Y=1.835 $X2=12.24 $Y2=1.96
r312 7 53 300 $w=1.7e-07 $l=3.47779e-07 $layer=licon1_PDIFF $count=2 $X=11.02
+ $Y=2.48 $X2=11.315 $Y2=2.365
r313 6 147 600 $w=1.7e-07 $l=3.1285e-07 $layer=licon1_PDIFF $count=1 $X=9.965
+ $Y=2.48 $X2=10.19 $Y2=2.69
r314 5 49 300 $w=1.7e-07 $l=4.12795e-07 $layer=licon1_PDIFF $count=2 $X=7.815
+ $Y=1.895 $X2=7.94 $Y2=2.25
r315 4 45 600 $w=1.7e-07 $l=5.6325e-07 $layer=licon1_PDIFF $count=1 $X=6.6
+ $Y=2.315 $X2=6.855 $Y2=2.765
r316 3 41 600 $w=1.7e-07 $l=1.1629e-06 $layer=licon1_PDIFF $count=1 $X=4.24
+ $Y=1.835 $X2=4.38 $Y2=2.93
r317 2 37 600 $w=1.7e-07 $l=5.60647e-07 $layer=licon1_PDIFF $count=1 $X=2.695
+ $Y=2.445 $X2=2.835 $Y2=2.94
r318 1 33 300 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_PDIFF $count=2 $X=1.005
+ $Y=2.445 $X2=1.145 $Y2=2.6
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRBP_2%A_359_489# 1 2 3 4 5 18 20 23 26 27 30 31
+ 34 37 39 45 47 48
c136 47 0 1.16025e-19 $X=5.52 $Y=2.49
r137 47 49 3.41465 $w=2.68e-07 $l=8e-08 $layer=LI1_cond $X=5.49 $Y=2.49 $X2=5.49
+ $Y2=2.57
r138 47 48 7.26708 $w=2.68e-07 $l=1.65e-07 $layer=LI1_cond $X=5.49 $Y=2.49
+ $X2=5.49 $Y2=2.325
r139 43 45 21.1154 $w=1.82e-07 $l=3.15e-07 $layer=LI1_cond $X=3.06 $Y=2.55
+ $X2=3.375 $Y2=2.55
r140 39 41 6.28605 $w=3.28e-07 $l=1.8e-07 $layer=LI1_cond $X=2.14 $Y=0.7
+ $X2=2.14 $Y2=0.88
r141 32 34 74.0481 $w=1.68e-07 $l=1.135e-06 $layer=LI1_cond $X=6.025 $Y=1.95
+ $X2=6.025 $Y2=0.815
r142 30 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.94 $Y=2.035
+ $X2=6.025 $Y2=1.95
r143 30 31 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=5.94 $Y=2.035
+ $X2=5.625 $Y2=2.035
r144 28 31 7.04737 $w=1.7e-07 $l=1.54771e-07 $layer=LI1_cond $X=5.507 $Y=2.12
+ $X2=5.625 $Y2=2.035
r145 28 48 10.0532 $w=2.33e-07 $l=2.05e-07 $layer=LI1_cond $X=5.507 $Y=2.12
+ $X2=5.507 $Y2=2.325
r146 27 45 11.1305 $w=1.82e-07 $l=1.74714e-07 $layer=LI1_cond $X=3.54 $Y=2.57
+ $X2=3.375 $Y2=2.55
r147 26 49 3.44395 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=5.355 $Y=2.57
+ $X2=5.49 $Y2=2.57
r148 26 27 118.412 $w=1.68e-07 $l=1.815e-06 $layer=LI1_cond $X=5.355 $Y=2.57
+ $X2=3.54 $Y2=2.57
r149 23 43 1.129 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=3.06 $Y=2.445
+ $X2=3.06 $Y2=2.55
r150 22 23 96.5562 $w=1.68e-07 $l=1.48e-06 $layer=LI1_cond $X=3.06 $Y=0.965
+ $X2=3.06 $Y2=2.445
r151 21 41 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.305 $Y=0.88
+ $X2=2.14 $Y2=0.88
r152 20 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.975 $Y=0.88
+ $X2=3.06 $Y2=0.965
r153 20 21 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.975 $Y=0.88
+ $X2=2.305 $Y2=0.88
r154 19 37 4.43891 $w=2.1e-07 $l=1.65e-07 $layer=LI1_cond $X=2.1 $Y=2.55
+ $X2=1.935 $Y2=2.55
r155 18 43 5.18805 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=2.975 $Y=2.55
+ $X2=3.06 $Y2=2.55
r156 18 19 46.2121 $w=2.08e-07 $l=8.75e-07 $layer=LI1_cond $X=2.975 $Y=2.55
+ $X2=2.1 $Y2=2.55
r157 5 47 600 $w=1.7e-07 $l=2.38485e-07 $layer=licon1_PDIFF $count=1 $X=5.37
+ $Y=2.315 $X2=5.52 $Y2=2.49
r158 4 45 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=3.235
+ $Y=2.445 $X2=3.375 $Y2=2.59
r159 3 37 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=1.795
+ $Y=2.445 $X2=1.935 $Y2=2.59
r160 2 34 182 $w=1.7e-07 $l=2.755e-07 $layer=licon1_NDIFF $count=1 $X=5.9
+ $Y=0.595 $X2=6.025 $Y2=0.815
r161 1 39 182 $w=1.7e-07 $l=3.68375e-07 $layer=licon1_NDIFF $count=1 $X=1.975
+ $Y=0.405 $X2=2.14 $Y2=0.7
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRBP_2%Q_N 1 2 7 8 9 10 11 12 13 22
r22 13 40 5.87094 $w=2.63e-07 $l=1.35e-07 $layer=LI1_cond $X=11.782 $Y=2.775
+ $X2=11.782 $Y2=2.91
r23 12 13 16.0907 $w=2.63e-07 $l=3.7e-07 $layer=LI1_cond $X=11.782 $Y=2.405
+ $X2=11.782 $Y2=2.775
r24 11 12 19.3523 $w=2.63e-07 $l=4.45e-07 $layer=LI1_cond $X=11.782 $Y=1.96
+ $X2=11.782 $Y2=2.405
r25 10 11 12.8291 $w=2.63e-07 $l=2.95e-07 $layer=LI1_cond $X=11.782 $Y=1.665
+ $X2=11.782 $Y2=1.96
r26 9 10 16.0907 $w=2.63e-07 $l=3.7e-07 $layer=LI1_cond $X=11.782 $Y=1.295
+ $X2=11.782 $Y2=1.665
r27 8 9 16.0907 $w=2.63e-07 $l=3.7e-07 $layer=LI1_cond $X=11.782 $Y=0.925
+ $X2=11.782 $Y2=1.295
r28 7 8 16.0907 $w=2.63e-07 $l=3.7e-07 $layer=LI1_cond $X=11.782 $Y=0.555
+ $X2=11.782 $Y2=0.925
r29 7 22 5.87094 $w=2.63e-07 $l=1.35e-07 $layer=LI1_cond $X=11.782 $Y=0.555
+ $X2=11.782 $Y2=0.42
r30 2 40 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=11.625
+ $Y=1.835 $X2=11.765 $Y2=2.91
r31 2 11 400 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=11.625
+ $Y=1.835 $X2=11.765 $Y2=1.96
r32 1 22 91 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=2 $X=11.645 $Y=0.24
+ $X2=11.785 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRBP_2%Q 1 2 7 8 9 10 11 12 13 22
r18 13 40 6.62042 $w=2.33e-07 $l=1.35e-07 $layer=LI1_cond $X=13.692 $Y=2.775
+ $X2=13.692 $Y2=2.91
r19 12 13 18.1448 $w=2.33e-07 $l=3.7e-07 $layer=LI1_cond $X=13.692 $Y=2.405
+ $X2=13.692 $Y2=2.775
r20 11 12 20.8421 $w=2.33e-07 $l=4.25e-07 $layer=LI1_cond $X=13.692 $Y=1.98
+ $X2=13.692 $Y2=2.405
r21 10 11 15.4476 $w=2.33e-07 $l=3.15e-07 $layer=LI1_cond $X=13.692 $Y=1.665
+ $X2=13.692 $Y2=1.98
r22 9 10 18.1448 $w=2.33e-07 $l=3.7e-07 $layer=LI1_cond $X=13.692 $Y=1.295
+ $X2=13.692 $Y2=1.665
r23 8 9 18.1448 $w=2.33e-07 $l=3.7e-07 $layer=LI1_cond $X=13.692 $Y=0.925
+ $X2=13.692 $Y2=1.295
r24 7 8 18.1448 $w=2.33e-07 $l=3.7e-07 $layer=LI1_cond $X=13.692 $Y=0.555
+ $X2=13.692 $Y2=0.925
r25 7 22 6.62042 $w=2.33e-07 $l=1.35e-07 $layer=LI1_cond $X=13.692 $Y=0.555
+ $X2=13.692 $Y2=0.42
r26 2 40 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=13.55
+ $Y=1.835 $X2=13.69 $Y2=2.91
r27 2 11 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=13.55
+ $Y=1.835 $X2=13.69 $Y2=1.98
r28 1 22 91 $w=1.7e-07 $l=1.9799e-07 $layer=licon1_NDIFF $count=2 $X=13.55
+ $Y=0.28 $X2=13.69 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRBP_2%VGND 1 2 3 4 5 6 7 8 9 10 33 37 41 45 49 53
+ 57 61 67 69 71 74 75 77 78 80 81 83 84 85 87 105 116 120 125 130 136 139 142
+ 145 148 152
c162 152 0 3.56444e-20 $X=14.16 $Y=0
c163 37 0 1.45423e-19 $X=3.445 $Y=0.615
c164 7 0 1.87138e-19 $X=11.23 $Y=0.24
r165 151 152 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.16 $Y=0
+ $X2=14.16 $Y2=0
r166 148 149 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.2 $Y=0
+ $X2=13.2 $Y2=0
r167 145 146 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.24 $Y=0
+ $X2=12.24 $Y2=0
r168 142 143 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.28 $Y=0
+ $X2=11.28 $Y2=0
r169 139 140 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=7.92 $Y=0
+ $X2=7.92 $Y2=0
r170 136 137 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0
+ $X2=0.72 $Y2=0
r171 134 152 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.68 $Y=0
+ $X2=14.16 $Y2=0
r172 134 149 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.68 $Y=0
+ $X2=13.2 $Y2=0
r173 133 134 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.68 $Y=0
+ $X2=13.68 $Y2=0
r174 131 148 8.23795 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=13.405 $Y=0
+ $X2=13.25 $Y2=0
r175 131 133 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=13.405 $Y=0
+ $X2=13.68 $Y2=0
r176 130 151 4.4964 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=13.98 $Y=0
+ $X2=14.19 $Y2=0
r177 130 133 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=13.98 $Y=0
+ $X2=13.68 $Y2=0
r178 129 149 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.72 $Y=0
+ $X2=13.2 $Y2=0
r179 129 146 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.72 $Y=0
+ $X2=12.24 $Y2=0
r180 128 129 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.72 $Y=0
+ $X2=12.72 $Y2=0
r181 126 145 8.42608 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=12.405 $Y=0
+ $X2=12.245 $Y2=0
r182 126 128 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=12.405 $Y=0
+ $X2=12.72 $Y2=0
r183 125 148 8.23795 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=13.095 $Y=0
+ $X2=13.25 $Y2=0
r184 125 128 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=13.095 $Y=0
+ $X2=12.72 $Y2=0
r185 124 146 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.76 $Y=0
+ $X2=12.24 $Y2=0
r186 124 143 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.76 $Y=0
+ $X2=11.28 $Y2=0
r187 123 124 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.76 $Y=0
+ $X2=11.76 $Y2=0
r188 121 142 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=11.48 $Y=0
+ $X2=11.335 $Y2=0
r189 121 123 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=11.48 $Y=0
+ $X2=11.76 $Y2=0
r190 120 145 8.42608 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=12.085 $Y=0
+ $X2=12.245 $Y2=0
r191 120 123 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=12.085 $Y=0
+ $X2=11.76 $Y2=0
r192 119 143 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.8 $Y=0
+ $X2=11.28 $Y2=0
r193 118 119 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.8 $Y=0
+ $X2=10.8 $Y2=0
r194 116 142 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=11.19 $Y=0
+ $X2=11.335 $Y2=0
r195 116 118 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=11.19 $Y=0
+ $X2=10.8 $Y2=0
r196 115 119 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=9.84 $Y=0
+ $X2=10.8 $Y2=0
r197 115 140 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=9.84 $Y=0
+ $X2=7.92 $Y2=0
r198 114 115 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=9.84 $Y=0
+ $X2=9.84 $Y2=0
r199 112 139 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.925 $Y=0
+ $X2=7.76 $Y2=0
r200 112 114 124.936 $w=1.68e-07 $l=1.915e-06 $layer=LI1_cond $X=7.925 $Y=0
+ $X2=9.84 $Y2=0
r201 111 140 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0
+ $X2=7.92 $Y2=0
r202 110 111 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=7.44 $Y=0
+ $X2=7.44 $Y2=0
r203 107 110 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=5.52 $Y=0
+ $X2=7.44 $Y2=0
r204 107 108 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.52 $Y=0
+ $X2=5.52 $Y2=0
r205 105 139 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.595 $Y=0
+ $X2=7.76 $Y2=0
r206 105 110 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=7.595 $Y=0
+ $X2=7.44 $Y2=0
r207 104 108 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0
+ $X2=5.52 $Y2=0
r208 103 104 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=0
+ $X2=5.04 $Y2=0
r209 101 104 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=0
+ $X2=5.04 $Y2=0
r210 100 101 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=0
+ $X2=4.08 $Y2=0
r211 98 101 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=0
+ $X2=4.08 $Y2=0
r212 97 98 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=0
+ $X2=3.12 $Y2=0
r213 95 98 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=1.2 $Y=0 $X2=3.12
+ $Y2=0
r214 95 137 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r215 94 97 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=3.12
+ $Y2=0
r216 94 95 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r217 92 136 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.855 $Y=0
+ $X2=0.69 $Y2=0
r218 92 94 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.855 $Y=0 $X2=1.2
+ $Y2=0
r219 90 137 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0
+ $X2=0.72 $Y2=0
r220 89 90 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r221 87 136 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.525 $Y=0
+ $X2=0.69 $Y2=0
r222 87 89 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.525 $Y=0
+ $X2=0.24 $Y2=0
r223 85 111 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=7.2 $Y=0
+ $X2=7.44 $Y2=0
r224 85 108 0.468274 $w=4.9e-07 $l=1.68e-06 $layer=MET1_cond $X=7.2 $Y=0
+ $X2=5.52 $Y2=0
r225 83 114 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=9.88 $Y=0 $X2=9.84
+ $Y2=0
r226 83 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.88 $Y=0
+ $X2=10.045 $Y2=0
r227 82 118 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=10.21 $Y=0 $X2=10.8
+ $Y2=0
r228 82 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.21 $Y=0
+ $X2=10.045 $Y2=0
r229 80 103 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=5.26 $Y=0 $X2=5.04
+ $Y2=0
r230 80 81 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.26 $Y=0 $X2=5.345
+ $Y2=0
r231 79 107 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=5.43 $Y=0 $X2=5.52
+ $Y2=0
r232 79 81 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.43 $Y=0 $X2=5.345
+ $Y2=0
r233 77 100 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=4.26 $Y=0 $X2=4.08
+ $Y2=0
r234 77 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.26 $Y=0 $X2=4.425
+ $Y2=0
r235 76 103 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=4.59 $Y=0 $X2=5.04
+ $Y2=0
r236 76 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.59 $Y=0 $X2=4.425
+ $Y2=0
r237 74 97 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=3.35 $Y=0 $X2=3.12
+ $Y2=0
r238 74 75 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.35 $Y=0 $X2=3.48
+ $Y2=0
r239 73 100 30.6631 $w=1.68e-07 $l=4.7e-07 $layer=LI1_cond $X=3.61 $Y=0 $X2=4.08
+ $Y2=0
r240 73 75 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.61 $Y=0 $X2=3.48
+ $Y2=0
r241 69 151 3.06184 $w=3.05e-07 $l=1.1025e-07 $layer=LI1_cond $X=14.132 $Y=0.085
+ $X2=14.19 $Y2=0
r242 69 71 12.8469 $w=3.03e-07 $l=3.4e-07 $layer=LI1_cond $X=14.132 $Y=0.085
+ $X2=14.132 $Y2=0.425
r243 65 148 0.701276 $w=3.1e-07 $l=8.5e-08 $layer=LI1_cond $X=13.25 $Y=0.085
+ $X2=13.25 $Y2=0
r244 65 67 12.6397 $w=3.08e-07 $l=3.4e-07 $layer=LI1_cond $X=13.25 $Y=0.085
+ $X2=13.25 $Y2=0.425
r245 61 63 19.6275 $w=3.18e-07 $l=5.45e-07 $layer=LI1_cond $X=12.245 $Y=0.385
+ $X2=12.245 $Y2=0.93
r246 59 145 0.800721 $w=3.2e-07 $l=8.5e-08 $layer=LI1_cond $X=12.245 $Y=0.085
+ $X2=12.245 $Y2=0
r247 59 61 10.8042 $w=3.18e-07 $l=3e-07 $layer=LI1_cond $X=12.245 $Y=0.085
+ $X2=12.245 $Y2=0.385
r248 55 142 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=11.335 $Y=0.085
+ $X2=11.335 $Y2=0
r249 55 57 11.9218 $w=2.88e-07 $l=3e-07 $layer=LI1_cond $X=11.335 $Y=0.085
+ $X2=11.335 $Y2=0.385
r250 51 84 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.045 $Y=0.085
+ $X2=10.045 $Y2=0
r251 51 53 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=10.045 $Y=0.085
+ $X2=10.045 $Y2=0.505
r252 47 139 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.76 $Y=0.085
+ $X2=7.76 $Y2=0
r253 47 49 13.2706 $w=3.28e-07 $l=3.8e-07 $layer=LI1_cond $X=7.76 $Y=0.085
+ $X2=7.76 $Y2=0.465
r254 43 81 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.345 $Y=0.085
+ $X2=5.345 $Y2=0
r255 43 45 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=5.345 $Y=0.085
+ $X2=5.345 $Y2=0.74
r256 39 78 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.425 $Y=0.085
+ $X2=4.425 $Y2=0
r257 39 41 18.1597 $w=3.28e-07 $l=5.2e-07 $layer=LI1_cond $X=4.425 $Y=0.085
+ $X2=4.425 $Y2=0.605
r258 35 75 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=3.48 $Y=0.085
+ $X2=3.48 $Y2=0
r259 35 37 23.4921 $w=2.58e-07 $l=5.3e-07 $layer=LI1_cond $X=3.48 $Y=0.085
+ $X2=3.48 $Y2=0.615
r260 31 136 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=0.085
+ $X2=0.69 $Y2=0
r261 31 33 17.9851 $w=3.28e-07 $l=5.15e-07 $layer=LI1_cond $X=0.69 $Y=0.085
+ $X2=0.69 $Y2=0.6
r262 10 71 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=13.98
+ $Y=0.28 $X2=14.12 $Y2=0.425
r263 9 67 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=13.135
+ $Y=0.28 $X2=13.26 $Y2=0.425
r264 8 63 182 $w=1.7e-07 $l=7.56769e-07 $layer=licon1_NDIFF $count=1 $X=12.075
+ $Y=0.24 $X2=12.215 $Y2=0.93
r265 8 61 182 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_NDIFF $count=1 $X=12.075
+ $Y=0.24 $X2=12.31 $Y2=0.385
r266 7 57 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=11.23
+ $Y=0.24 $X2=11.355 $Y2=0.385
r267 6 53 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=9.905
+ $Y=0.34 $X2=10.045 $Y2=0.505
r268 5 49 182 $w=1.7e-07 $l=3.54083e-07 $layer=licon1_NDIFF $count=1 $X=7.465
+ $Y=0.595 $X2=7.76 $Y2=0.465
r269 4 45 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=5.205
+ $Y=0.595 $X2=5.345 $Y2=0.74
r270 3 41 182 $w=1.7e-07 $l=2.04939e-07 $layer=licon1_NDIFF $count=1 $X=4.225
+ $Y=0.595 $X2=4.425 $Y2=0.605
r271 2 37 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=3.305
+ $Y=0.405 $X2=3.445 $Y2=0.615
r272 1 33 182 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.405 $X2=0.69 $Y2=0.6
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRBP_2%noxref_25 1 2 7 9 12
c36 9 0 1.84245e-19 $X=1.302 $Y=0.35
c37 7 0 1.07392e-19 $X=2.85 $Y=0.35
r38 12 15 6.28605 $w=3.28e-07 $l=1.8e-07 $layer=LI1_cond $X=3.015 $Y=0.35
+ $X2=3.015 $Y2=0.53
r39 9 11 8.4022 $w=3.63e-07 $l=2.5e-07 $layer=LI1_cond $X=1.302 $Y=0.35
+ $X2=1.302 $Y2=0.6
r40 8 9 5.19232 $w=1.7e-07 $l=1.88e-07 $layer=LI1_cond $X=1.49 $Y=0.35 $X2=1.302
+ $Y2=0.35
r41 7 12 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.85 $Y=0.35
+ $X2=3.015 $Y2=0.35
r42 7 8 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=2.85 $Y=0.35 $X2=1.49
+ $Y2=0.35
r43 2 15 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=2.875
+ $Y=0.405 $X2=3.015 $Y2=0.53
r44 1 11 182 $w=1.7e-07 $l=2.498e-07 $layer=licon1_NDIFF $count=1 $X=1.2
+ $Y=0.405 $X2=1.325 $Y2=0.6
.ends

