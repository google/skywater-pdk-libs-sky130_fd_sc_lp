* File: sky130_fd_sc_lp__xnor2_4.pxi.spice
* Created: Fri Aug 28 11:35:15 2020
* 
x_PM_SKY130_FD_SC_LP__XNOR2_4%A N_A_M1019_g N_A_M1006_g N_A_M1031_g N_A_M1017_g
+ N_A_M1024_g N_A_M1036_g N_A_M1037_g N_A_M1027_g N_A_M1018_g N_A_M1008_g
+ N_A_M1014_g N_A_M1030_g N_A_M1026_g N_A_M1032_g N_A_M1039_g N_A_M1034_g
+ N_A_c_169_n N_A_c_185_n N_A_c_198_p N_A_c_286_p N_A_c_186_n N_A_c_170_n
+ N_A_c_188_n N_A_c_171_n N_A_c_172_n N_A_c_173_n N_A_c_190_n A A N_A_c_174_n
+ N_A_c_175_n PM_SKY130_FD_SC_LP__XNOR2_4%A
x_PM_SKY130_FD_SC_LP__XNOR2_4%B N_B_M1000_g N_B_M1002_g N_B_M1003_g N_B_M1012_g
+ N_B_M1011_g N_B_M1013_g N_B_M1023_g N_B_M1022_g N_B_c_440_n N_B_M1007_g
+ N_B_M1004_g N_B_c_441_n N_B_M1016_g N_B_M1015_g N_B_c_442_n N_B_M1021_g
+ N_B_M1025_g N_B_c_443_n N_B_M1035_g N_B_M1028_g N_B_c_431_n N_B_c_445_n
+ N_B_c_432_n N_B_c_447_n B N_B_c_433_n N_B_c_434_n N_B_c_435_n
+ PM_SKY130_FD_SC_LP__XNOR2_4%B
x_PM_SKY130_FD_SC_LP__XNOR2_4%A_808_39# N_A_808_39#_M1004_d N_A_808_39#_M1025_d
+ N_A_808_39#_M1008_s N_A_808_39#_M1026_s N_A_808_39#_M1007_d
+ N_A_808_39#_M1021_d N_A_808_39#_M1001_g N_A_808_39#_M1005_g
+ N_A_808_39#_M1009_g N_A_808_39#_M1020_g N_A_808_39#_M1010_g
+ N_A_808_39#_c_640_n N_A_808_39#_c_641_n N_A_808_39#_M1029_g
+ N_A_808_39#_M1033_g N_A_808_39#_M1038_g N_A_808_39#_c_643_n
+ N_A_808_39#_c_780_p N_A_808_39#_c_658_n N_A_808_39#_c_659_n
+ N_A_808_39#_c_774_p N_A_808_39#_c_694_n N_A_808_39#_c_696_n
+ N_A_808_39#_c_783_p N_A_808_39#_c_729_n N_A_808_39#_c_644_n
+ N_A_808_39#_c_737_n N_A_808_39#_c_784_p N_A_808_39#_c_660_n
+ N_A_808_39#_c_645_n N_A_808_39#_c_646_n N_A_808_39#_c_647_n
+ N_A_808_39#_c_648_n N_A_808_39#_c_662_n N_A_808_39#_c_649_n
+ N_A_808_39#_c_755_n N_A_808_39#_c_650_n N_A_808_39#_c_762_n
+ N_A_808_39#_c_651_n PM_SKY130_FD_SC_LP__XNOR2_4%A_808_39#
x_PM_SKY130_FD_SC_LP__XNOR2_4%VPWR N_VPWR_M1019_d N_VPWR_M1031_d N_VPWR_M1037_d
+ N_VPWR_M1020_d N_VPWR_M1038_d N_VPWR_M1014_d N_VPWR_M1039_d N_VPWR_M1016_s
+ N_VPWR_M1035_s N_VPWR_c_869_n N_VPWR_c_870_n N_VPWR_c_871_n N_VPWR_c_872_n
+ N_VPWR_c_873_n N_VPWR_c_874_n N_VPWR_c_875_n N_VPWR_c_876_n N_VPWR_c_877_n
+ N_VPWR_c_878_n N_VPWR_c_879_n N_VPWR_c_880_n N_VPWR_c_881_n N_VPWR_c_882_n
+ N_VPWR_c_883_n N_VPWR_c_884_n VPWR N_VPWR_c_885_n N_VPWR_c_886_n
+ N_VPWR_c_887_n N_VPWR_c_888_n N_VPWR_c_889_n N_VPWR_c_890_n N_VPWR_c_891_n
+ N_VPWR_c_892_n N_VPWR_c_868_n PM_SKY130_FD_SC_LP__XNOR2_4%VPWR
x_PM_SKY130_FD_SC_LP__XNOR2_4%A_110_367# N_A_110_367#_M1019_s
+ N_A_110_367#_M1036_s N_A_110_367#_M1012_d N_A_110_367#_M1022_d
+ N_A_110_367#_c_1030_n N_A_110_367#_c_1037_n N_A_110_367#_c_1032_n
+ N_A_110_367#_c_1034_n PM_SKY130_FD_SC_LP__XNOR2_4%A_110_367#
x_PM_SKY130_FD_SC_LP__XNOR2_4%Y N_Y_M1001_d N_Y_M1010_d N_Y_M1002_s N_Y_M1013_s
+ N_Y_M1005_s N_Y_M1033_s N_Y_c_1063_n N_Y_c_1064_n N_Y_c_1065_n N_Y_c_1087_n
+ N_Y_c_1069_n N_Y_c_1094_n N_Y_c_1098_n N_Y_c_1107_n N_Y_c_1193_p N_Y_c_1066_n
+ N_Y_c_1109_n N_Y_c_1138_n N_Y_c_1110_n N_Y_c_1140_n N_Y_c_1067_n Y Y
+ N_Y_c_1111_n Y PM_SKY130_FD_SC_LP__XNOR2_4%Y
x_PM_SKY130_FD_SC_LP__XNOR2_4%A_31_65# N_A_31_65#_M1006_d N_A_31_65#_M1017_d
+ N_A_31_65#_M1000_d N_A_31_65#_M1011_d N_A_31_65#_M1027_d N_A_31_65#_M1009_s
+ N_A_31_65#_M1029_s N_A_31_65#_c_1206_n N_A_31_65#_c_1218_n N_A_31_65#_c_1207_n
+ N_A_31_65#_c_1208_n N_A_31_65#_c_1223_n N_A_31_65#_c_1209_n
+ N_A_31_65#_c_1231_n N_A_31_65#_c_1210_n N_A_31_65#_c_1224_n
+ N_A_31_65#_c_1225_n N_A_31_65#_c_1211_n N_A_31_65#_c_1212_n
+ N_A_31_65#_c_1244_n N_A_31_65#_c_1213_n N_A_31_65#_c_1214_n
+ N_A_31_65#_c_1276_n N_A_31_65#_c_1277_n N_A_31_65#_c_1278_n
+ N_A_31_65#_c_1215_n PM_SKY130_FD_SC_LP__XNOR2_4%A_31_65#
x_PM_SKY130_FD_SC_LP__XNOR2_4%VGND N_VGND_M1006_s N_VGND_M1024_s N_VGND_M1003_s
+ N_VGND_M1023_s N_VGND_M1018_d N_VGND_M1032_d N_VGND_c_1326_n N_VGND_c_1327_n
+ N_VGND_c_1328_n N_VGND_c_1329_n N_VGND_c_1330_n N_VGND_c_1331_n
+ N_VGND_c_1332_n N_VGND_c_1333_n N_VGND_c_1334_n N_VGND_c_1335_n
+ N_VGND_c_1336_n N_VGND_c_1337_n N_VGND_c_1338_n N_VGND_c_1339_n VGND
+ N_VGND_c_1340_n N_VGND_c_1341_n N_VGND_c_1342_n N_VGND_c_1343_n
+ N_VGND_c_1344_n N_VGND_c_1345_n PM_SKY130_FD_SC_LP__XNOR2_4%VGND
x_PM_SKY130_FD_SC_LP__XNOR2_4%A_1235_65# N_A_1235_65#_M1018_s
+ N_A_1235_65#_M1030_s N_A_1235_65#_M1034_s N_A_1235_65#_M1015_s
+ N_A_1235_65#_M1028_s N_A_1235_65#_c_1483_n N_A_1235_65#_c_1493_n
+ N_A_1235_65#_c_1484_n N_A_1235_65#_c_1485_n N_A_1235_65#_c_1498_n
+ N_A_1235_65#_c_1514_n N_A_1235_65#_c_1486_n N_A_1235_65#_c_1487_n
+ N_A_1235_65#_c_1519_n N_A_1235_65#_c_1488_n N_A_1235_65#_c_1489_n
+ N_A_1235_65#_c_1525_n N_A_1235_65#_c_1490_n
+ PM_SKY130_FD_SC_LP__XNOR2_4%A_1235_65#
cc_1 VNB N_A_M1006_g 0.0250755f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=0.745
cc_2 VNB N_A_M1017_g 0.0201423f $X=-0.19 $Y=-0.245 $X2=1.025 $Y2=0.745
cc_3 VNB N_A_M1024_g 0.0193564f $X=-0.19 $Y=-0.245 $X2=1.455 $Y2=0.745
cc_4 VNB N_A_M1027_g 0.0208081f $X=-0.19 $Y=-0.245 $X2=3.685 $Y2=0.745
cc_5 VNB N_A_M1018_g 0.0244634f $X=-0.19 $Y=-0.245 $X2=6.515 $Y2=0.745
cc_6 VNB N_A_M1030_g 0.0200802f $X=-0.19 $Y=-0.245 $X2=7.025 $Y2=0.745
cc_7 VNB N_A_M1032_g 0.0190877f $X=-0.19 $Y=-0.245 $X2=7.455 $Y2=0.745
cc_8 VNB N_A_M1034_g 0.0193946f $X=-0.19 $Y=-0.245 $X2=7.885 $Y2=0.745
cc_9 VNB N_A_c_169_n 0.00174495f $X=-0.19 $Y=-0.245 $X2=1.427 $Y2=1.75
cc_10 VNB N_A_c_170_n 0.0250704f $X=-0.19 $Y=-0.245 $X2=3.665 $Y2=1.51
cc_11 VNB N_A_c_171_n 7.55444e-19 $X=-0.19 $Y=-0.245 $X2=6.39 $Y2=1.765
cc_12 VNB N_A_c_172_n 0.00232352f $X=-0.19 $Y=-0.245 $X2=6.475 $Y2=1.51
cc_13 VNB N_A_c_173_n 0.00123532f $X=-0.19 $Y=-0.245 $X2=7.705 $Y2=1.51
cc_14 VNB N_A_c_174_n 0.0592876f $X=-0.19 $Y=-0.245 $X2=1.495 $Y2=1.51
cc_15 VNB N_A_c_175_n 0.0674048f $X=-0.19 $Y=-0.245 $X2=7.885 $Y2=1.51
cc_16 VNB N_B_M1000_g 0.0193562f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.465
cc_17 VNB N_B_M1003_g 0.0191712f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=2.465
cc_18 VNB N_B_M1011_g 0.0191712f $X=-0.19 $Y=-0.245 $X2=1.455 $Y2=0.745
cc_19 VNB N_B_M1023_g 0.0202608f $X=-0.19 $Y=-0.245 $X2=3.645 $Y2=2.465
cc_20 VNB N_B_M1004_g 0.019205f $X=-0.19 $Y=-0.245 $X2=6.56 $Y2=2.465
cc_21 VNB N_B_M1015_g 0.0190024f $X=-0.19 $Y=-0.245 $X2=7.025 $Y2=1.345
cc_22 VNB N_B_M1025_g 0.0189994f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_B_M1028_g 0.0230814f $X=-0.19 $Y=-0.245 $X2=7.85 $Y2=2.465
cc_24 VNB N_B_c_431_n 0.00127856f $X=-0.19 $Y=-0.245 $X2=7.885 $Y2=1.345
cc_25 VNB N_B_c_432_n 0.00629445f $X=-0.19 $Y=-0.245 $X2=3.665 $Y2=1.765
cc_26 VNB N_B_c_433_n 0.0659705f $X=-0.19 $Y=-0.245 $X2=3.665 $Y2=2.015
cc_27 VNB N_B_c_434_n 0.00114442f $X=-0.19 $Y=-0.245 $X2=1.025 $Y2=1.51
cc_28 VNB N_B_c_435_n 0.0684576f $X=-0.19 $Y=-0.245 $X2=1.29 $Y2=1.51
cc_29 VNB N_A_808_39#_M1001_g 0.0187781f $X=-0.19 $Y=-0.245 $X2=1.495 $Y2=1.675
cc_30 VNB N_A_808_39#_M1009_g 0.0187f $X=-0.19 $Y=-0.245 $X2=3.685 $Y2=1.345
cc_31 VNB N_A_808_39#_M1010_g 0.0195012f $X=-0.19 $Y=-0.245 $X2=6.56 $Y2=1.675
cc_32 VNB N_A_808_39#_c_640_n 0.015776f $X=-0.19 $Y=-0.245 $X2=6.56 $Y2=2.465
cc_33 VNB N_A_808_39#_c_641_n 0.0434854f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_808_39#_M1029_g 0.0227784f $X=-0.19 $Y=-0.245 $X2=6.99 $Y2=2.465
cc_35 VNB N_A_808_39#_c_643_n 0.0126811f $X=-0.19 $Y=-0.245 $X2=7.885 $Y2=1.345
cc_36 VNB N_A_808_39#_c_644_n 0.00224127f $X=-0.19 $Y=-0.245 $X2=3.665 $Y2=2.015
cc_37 VNB N_A_808_39#_c_645_n 0.010294f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=1.51
cc_38 VNB N_A_808_39#_c_646_n 0.0197549f $X=-0.19 $Y=-0.245 $X2=1.29 $Y2=1.51
cc_39 VNB N_A_808_39#_c_647_n 0.00112395f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_808_39#_c_648_n 0.011145f $X=-0.19 $Y=-0.245 $X2=3.665 $Y2=1.51
cc_41 VNB N_A_808_39#_c_649_n 0.00211339f $X=-0.19 $Y=-0.245 $X2=6.99 $Y2=1.51
cc_42 VNB N_A_808_39#_c_650_n 0.00228422f $X=-0.19 $Y=-0.245 $X2=7.455 $Y2=1.51
cc_43 VNB N_A_808_39#_c_651_n 0.0529446f $X=-0.19 $Y=-0.245 $X2=1.427 $Y2=1.582
cc_44 VNB N_VPWR_c_868_n 0.422413f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_Y_c_1063_n 0.0197038f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_Y_c_1064_n 0.0284631f $X=-0.19 $Y=-0.245 $X2=1.495 $Y2=1.675
cc_47 VNB N_Y_c_1065_n 0.00942816f $X=-0.19 $Y=-0.245 $X2=1.495 $Y2=2.465
cc_48 VNB N_Y_c_1066_n 0.00466212f $X=-0.19 $Y=-0.245 $X2=6.56 $Y2=1.675
cc_49 VNB N_Y_c_1067_n 0.00133697f $X=-0.19 $Y=-0.245 $X2=7.42 $Y2=1.675
cc_50 VNB N_A_31_65#_c_1206_n 0.0191545f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_31_65#_c_1207_n 0.00722716f $X=-0.19 $Y=-0.245 $X2=3.645 $Y2=2.465
cc_52 VNB N_A_31_65#_c_1208_n 0.0020741f $X=-0.19 $Y=-0.245 $X2=3.685 $Y2=0.745
cc_53 VNB N_A_31_65#_c_1209_n 0.00214592f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_31_65#_c_1210_n 0.00214592f $X=-0.19 $Y=-0.245 $X2=6.99 $Y2=2.465
cc_55 VNB N_A_31_65#_c_1211_n 0.0019956f $X=-0.19 $Y=-0.245 $X2=7.42 $Y2=2.465
cc_56 VNB N_A_31_65#_c_1212_n 0.00203674f $X=-0.19 $Y=-0.245 $X2=7.42 $Y2=2.465
cc_57 VNB N_A_31_65#_c_1213_n 0.00749893f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_31_65#_c_1214_n 0.00446793f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_31_65#_c_1215_n 0.00210948f $X=-0.19 $Y=-0.245 $X2=1.57 $Y2=2.015
cc_60 VNB N_VGND_c_1326_n 0.00472689f $X=-0.19 $Y=-0.245 $X2=1.495 $Y2=1.675
cc_61 VNB N_VGND_c_1327_n 0.00178357f $X=-0.19 $Y=-0.245 $X2=3.645 $Y2=1.675
cc_62 VNB N_VGND_c_1328_n 0.00177331f $X=-0.19 $Y=-0.245 $X2=3.685 $Y2=1.345
cc_63 VNB N_VGND_c_1329_n 0.00453825f $X=-0.19 $Y=-0.245 $X2=6.515 $Y2=1.345
cc_64 VNB N_VGND_c_1330_n 0.00476969f $X=-0.19 $Y=-0.245 $X2=6.56 $Y2=1.675
cc_65 VNB N_VGND_c_1331_n 0.00229999f $X=-0.19 $Y=-0.245 $X2=6.99 $Y2=1.675
cc_66 VNB N_VGND_c_1332_n 0.0129698f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_1333_n 0.00546567f $X=-0.19 $Y=-0.245 $X2=7.025 $Y2=1.345
cc_68 VNB N_VGND_c_1334_n 0.0129698f $X=-0.19 $Y=-0.245 $X2=7.025 $Y2=0.745
cc_69 VNB N_VGND_c_1335_n 0.0057893f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_VGND_c_1336_n 0.0725107f $X=-0.19 $Y=-0.245 $X2=7.42 $Y2=2.465
cc_71 VNB N_VGND_c_1337_n 0.0058157f $X=-0.19 $Y=-0.245 $X2=7.42 $Y2=2.465
cc_72 VNB N_VGND_c_1338_n 0.0132237f $X=-0.19 $Y=-0.245 $X2=7.455 $Y2=1.345
cc_73 VNB N_VGND_c_1339_n 0.00546618f $X=-0.19 $Y=-0.245 $X2=7.455 $Y2=0.745
cc_74 VNB N_VGND_c_1340_n 0.0188687f $X=-0.19 $Y=-0.245 $X2=7.85 $Y2=1.675
cc_75 VNB N_VGND_c_1341_n 0.0133039f $X=-0.19 $Y=-0.245 $X2=7.885 $Y2=0.745
cc_76 VNB N_VGND_c_1342_n 0.0533913f $X=-0.19 $Y=-0.245 $X2=3.665 $Y2=2.015
cc_77 VNB N_VGND_c_1343_n 0.514694f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_78 VNB N_VGND_c_1344_n 0.00581519f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_VGND_c_1345_n 0.00546567f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_A_1235_65#_c_1483_n 0.00656764f $X=-0.19 $Y=-0.245 $X2=1.455
+ $Y2=0.745
cc_81 VNB N_A_1235_65#_c_1484_n 0.0018836f $X=-0.19 $Y=-0.245 $X2=1.495
+ $Y2=1.675
cc_82 VNB N_A_1235_65#_c_1485_n 0.00223748f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_A_1235_65#_c_1486_n 0.00262279f $X=-0.19 $Y=-0.245 $X2=3.685
+ $Y2=0.745
cc_84 VNB N_A_1235_65#_c_1487_n 0.00190905f $X=-0.19 $Y=-0.245 $X2=3.685
+ $Y2=0.745
cc_85 VNB N_A_1235_65#_c_1488_n 0.0118917f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_A_1235_65#_c_1489_n 0.0180172f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_A_1235_65#_c_1490_n 0.00136716f $X=-0.19 $Y=-0.245 $X2=7.025
+ $Y2=0.745
cc_88 VPB N_A_M1019_g 0.0209109f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.465
cc_89 VPB N_A_M1031_g 0.0197283f $X=-0.19 $Y=1.655 $X2=0.905 $Y2=2.465
cc_90 VPB N_A_M1036_g 0.0195088f $X=-0.19 $Y=1.655 $X2=1.495 $Y2=2.465
cc_91 VPB N_A_M1037_g 0.0176798f $X=-0.19 $Y=1.655 $X2=3.645 $Y2=2.465
cc_92 VPB N_A_M1008_g 0.0184626f $X=-0.19 $Y=1.655 $X2=6.56 $Y2=2.465
cc_93 VPB N_A_M1014_g 0.0175335f $X=-0.19 $Y=1.655 $X2=6.99 $Y2=2.465
cc_94 VPB N_A_M1026_g 0.0175359f $X=-0.19 $Y=1.655 $X2=7.42 $Y2=2.465
cc_95 VPB N_A_M1039_g 0.0179929f $X=-0.19 $Y=1.655 $X2=7.85 $Y2=2.465
cc_96 VPB N_A_c_169_n 7.92397e-19 $X=-0.19 $Y=1.655 $X2=1.427 $Y2=1.75
cc_97 VPB N_A_c_185_n 9.5877e-19 $X=-0.19 $Y=1.655 $X2=1.427 $Y2=1.93
cc_98 VPB N_A_c_186_n 0.00171885f $X=-0.19 $Y=1.655 $X2=3.665 $Y2=1.51
cc_99 VPB N_A_c_170_n 0.00622015f $X=-0.19 $Y=1.655 $X2=3.665 $Y2=1.51
cc_100 VPB N_A_c_188_n 0.0138651f $X=-0.19 $Y=1.655 $X2=6.305 $Y2=1.85
cc_101 VPB N_A_c_171_n 0.00232169f $X=-0.19 $Y=1.655 $X2=6.39 $Y2=1.765
cc_102 VPB N_A_c_190_n 8.19341e-19 $X=-0.19 $Y=1.655 $X2=3.665 $Y2=1.85
cc_103 VPB A 0.00638985f $X=-0.19 $Y=1.655 $X2=1.115 $Y2=1.58
cc_104 VPB N_A_c_174_n 0.0134798f $X=-0.19 $Y=1.655 $X2=1.495 $Y2=1.51
cc_105 VPB N_A_c_175_n 0.0164028f $X=-0.19 $Y=1.655 $X2=7.885 $Y2=1.51
cc_106 VPB N_B_M1002_g 0.0190224f $X=-0.19 $Y=1.655 $X2=0.515 $Y2=0.745
cc_107 VPB N_B_M1012_g 0.0180123f $X=-0.19 $Y=1.655 $X2=1.025 $Y2=0.745
cc_108 VPB N_B_M1013_g 0.0181366f $X=-0.19 $Y=1.655 $X2=1.495 $Y2=2.465
cc_109 VPB N_B_M1022_g 0.0184286f $X=-0.19 $Y=1.655 $X2=3.685 $Y2=0.745
cc_110 VPB N_B_c_440_n 0.0159075f $X=-0.19 $Y=1.655 $X2=6.515 $Y2=1.345
cc_111 VPB N_B_c_441_n 0.0158138f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_112 VPB N_B_c_442_n 0.0158117f $X=-0.19 $Y=1.655 $X2=7.025 $Y2=0.745
cc_113 VPB N_B_c_443_n 0.0183612f $X=-0.19 $Y=1.655 $X2=7.455 $Y2=0.745
cc_114 VPB N_B_c_431_n 0.00133468f $X=-0.19 $Y=1.655 $X2=7.885 $Y2=1.345
cc_115 VPB N_B_c_445_n 0.00530689f $X=-0.19 $Y=1.655 $X2=1.427 $Y2=1.93
cc_116 VPB N_B_c_432_n 0.0210011f $X=-0.19 $Y=1.655 $X2=3.665 $Y2=1.765
cc_117 VPB N_B_c_447_n 0.00299325f $X=-0.19 $Y=1.655 $X2=3.665 $Y2=1.51
cc_118 VPB B 0.00178588f $X=-0.19 $Y=1.655 $X2=3.83 $Y2=1.85
cc_119 VPB N_B_c_433_n 0.0133993f $X=-0.19 $Y=1.655 $X2=3.665 $Y2=2.015
cc_120 VPB N_B_c_434_n 0.00668211f $X=-0.19 $Y=1.655 $X2=1.025 $Y2=1.51
cc_121 VPB N_B_c_435_n 0.023023f $X=-0.19 $Y=1.655 $X2=1.29 $Y2=1.51
cc_122 VPB N_A_808_39#_M1005_g 0.0183619f $X=-0.19 $Y=1.655 $X2=3.645 $Y2=1.675
cc_123 VPB N_A_808_39#_M1020_g 0.0240761f $X=-0.19 $Y=1.655 $X2=6.515 $Y2=1.345
cc_124 VPB N_A_808_39#_c_640_n 0.0121883f $X=-0.19 $Y=1.655 $X2=6.56 $Y2=2.465
cc_125 VPB N_A_808_39#_c_641_n 0.0164749f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_126 VPB N_A_808_39#_M1033_g 0.0232092f $X=-0.19 $Y=1.655 $X2=7.025 $Y2=0.745
cc_127 VPB N_A_808_39#_M1038_g 0.0181721f $X=-0.19 $Y=1.655 $X2=7.42 $Y2=2.465
cc_128 VPB N_A_808_39#_c_658_n 0.00253078f $X=-0.19 $Y=1.655 $X2=3.665 $Y2=1.765
cc_129 VPB N_A_808_39#_c_659_n 0.00192526f $X=-0.19 $Y=1.655 $X2=3.665 $Y2=1.51
cc_130 VPB N_A_808_39#_c_660_n 0.00942129f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=1.51
cc_131 VPB N_A_808_39#_c_646_n 0.012264f $X=-0.19 $Y=1.655 $X2=1.29 $Y2=1.51
cc_132 VPB N_A_808_39#_c_662_n 0.00157076f $X=-0.19 $Y=1.655 $X2=3.665 $Y2=1.345
cc_133 VPB N_A_808_39#_c_651_n 0.00946866f $X=-0.19 $Y=1.655 $X2=1.427 $Y2=1.582
cc_134 VPB N_VPWR_c_869_n 0.0103398f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_135 VPB N_VPWR_c_870_n 0.0352145f $X=-0.19 $Y=1.655 $X2=3.685 $Y2=0.745
cc_136 VPB N_VPWR_c_871_n 4.89148e-19 $X=-0.19 $Y=1.655 $X2=6.515 $Y2=0.745
cc_137 VPB N_VPWR_c_872_n 0.0037094f $X=-0.19 $Y=1.655 $X2=6.56 $Y2=2.465
cc_138 VPB N_VPWR_c_873_n 3.16049e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_139 VPB N_VPWR_c_874_n 0.0129398f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_140 VPB N_VPWR_c_875_n 3.0911e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_141 VPB N_VPWR_c_876_n 3.0911e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_142 VPB N_VPWR_c_877_n 0.0114562f $X=-0.19 $Y=1.655 $X2=7.85 $Y2=2.465
cc_143 VPB N_VPWR_c_878_n 0.0352012f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_144 VPB N_VPWR_c_879_n 0.0579909f $X=-0.19 $Y=1.655 $X2=7.885 $Y2=0.745
cc_145 VPB N_VPWR_c_880_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_146 VPB N_VPWR_c_881_n 0.0154574f $X=-0.19 $Y=1.655 $X2=1.427 $Y2=1.93
cc_147 VPB N_VPWR_c_882_n 0.00420242f $X=-0.19 $Y=1.655 $X2=3.5 $Y2=2.015
cc_148 VPB N_VPWR_c_883_n 0.0149302f $X=-0.19 $Y=1.655 $X2=1.57 $Y2=2.015
cc_149 VPB N_VPWR_c_884_n 0.00436868f $X=-0.19 $Y=1.655 $X2=3.665 $Y2=1.765
cc_150 VPB N_VPWR_c_885_n 0.0157043f $X=-0.19 $Y=1.655 $X2=3.665 $Y2=1.51
cc_151 VPB N_VPWR_c_886_n 0.0192284f $X=-0.19 $Y=1.655 $X2=7.705 $Y2=1.51
cc_152 VPB N_VPWR_c_887_n 0.0129398f $X=-0.19 $Y=1.655 $X2=0.515 $Y2=1.51
cc_153 VPB N_VPWR_c_888_n 0.0129398f $X=-0.19 $Y=1.655 $X2=1.025 $Y2=1.51
cc_154 VPB N_VPWR_c_889_n 0.0103178f $X=-0.19 $Y=1.655 $X2=3.665 $Y2=1.675
cc_155 VPB N_VPWR_c_890_n 0.0204351f $X=-0.19 $Y=1.655 $X2=7.42 $Y2=1.51
cc_156 VPB N_VPWR_c_891_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=1.582
cc_157 VPB N_VPWR_c_892_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_158 VPB N_VPWR_c_868_n 0.0458569f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_159 VPB N_Y_c_1063_n 0.0115862f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_160 VPB N_Y_c_1069_n 0.00754068f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_161 N_A_M1024_g N_B_M1000_g 0.0386035f $X=1.455 $Y=0.745 $X2=0 $Y2=0
cc_162 N_A_M1036_g N_B_M1002_g 0.0544899f $X=1.495 $Y=2.465 $X2=0 $Y2=0
cc_163 N_A_c_169_n N_B_M1002_g 2.78861e-19 $X=1.427 $Y=1.75 $X2=0 $Y2=0
cc_164 N_A_c_185_n N_B_M1002_g 0.00112333f $X=1.427 $Y=1.93 $X2=0 $Y2=0
cc_165 N_A_c_198_p N_B_M1002_g 0.0113592f $X=3.5 $Y=2.015 $X2=0 $Y2=0
cc_166 N_A_c_198_p N_B_M1012_g 0.0104705f $X=3.5 $Y=2.015 $X2=0 $Y2=0
cc_167 N_A_c_198_p N_B_M1013_g 0.0104777f $X=3.5 $Y=2.015 $X2=0 $Y2=0
cc_168 N_A_M1027_g N_B_M1023_g 0.0327867f $X=3.685 $Y=0.745 $X2=0 $Y2=0
cc_169 N_A_M1037_g N_B_M1022_g 0.0542152f $X=3.645 $Y=2.465 $X2=0 $Y2=0
cc_170 N_A_c_198_p N_B_M1022_g 0.0106983f $X=3.5 $Y=2.015 $X2=0 $Y2=0
cc_171 N_A_c_186_n N_B_M1022_g 7.74286e-19 $X=3.665 $Y=1.51 $X2=0 $Y2=0
cc_172 N_A_c_190_n N_B_M1022_g 0.00433446f $X=3.665 $Y=1.85 $X2=0 $Y2=0
cc_173 N_A_M1034_g N_B_M1004_g 0.0224768f $X=7.885 $Y=0.745 $X2=0 $Y2=0
cc_174 N_A_c_169_n N_B_c_431_n 0.0142789f $X=1.427 $Y=1.75 $X2=0 $Y2=0
cc_175 N_A_c_198_p N_B_c_431_n 0.027187f $X=3.5 $Y=2.015 $X2=0 $Y2=0
cc_176 N_A_c_174_n N_B_c_431_n 3.66386e-19 $X=1.495 $Y=1.51 $X2=0 $Y2=0
cc_177 N_A_c_198_p N_B_c_445_n 0.0434451f $X=3.5 $Y=2.015 $X2=0 $Y2=0
cc_178 N_A_c_186_n N_B_c_445_n 0.0131562f $X=3.665 $Y=1.51 $X2=0 $Y2=0
cc_179 N_A_c_170_n N_B_c_445_n 7.95579e-19 $X=3.665 $Y=1.51 $X2=0 $Y2=0
cc_180 N_A_M1008_g N_B_c_432_n 0.00705804f $X=6.56 $Y=2.465 $X2=0 $Y2=0
cc_181 N_A_M1014_g N_B_c_432_n 0.00233988f $X=6.99 $Y=2.465 $X2=0 $Y2=0
cc_182 N_A_M1026_g N_B_c_432_n 0.00233988f $X=7.42 $Y=2.465 $X2=0 $Y2=0
cc_183 N_A_M1039_g N_B_c_432_n 0.00246119f $X=7.85 $Y=2.465 $X2=0 $Y2=0
cc_184 N_A_c_198_p N_B_c_432_n 0.0202764f $X=3.5 $Y=2.015 $X2=0 $Y2=0
cc_185 N_A_c_186_n N_B_c_432_n 0.0221483f $X=3.665 $Y=1.51 $X2=0 $Y2=0
cc_186 N_A_c_170_n N_B_c_432_n 7.93769e-19 $X=3.665 $Y=1.51 $X2=0 $Y2=0
cc_187 N_A_c_188_n N_B_c_432_n 0.0734108f $X=6.305 $Y=1.85 $X2=0 $Y2=0
cc_188 N_A_c_171_n N_B_c_432_n 0.014126f $X=6.39 $Y=1.765 $X2=0 $Y2=0
cc_189 N_A_c_172_n N_B_c_432_n 0.00230187f $X=6.475 $Y=1.51 $X2=0 $Y2=0
cc_190 N_A_c_173_n N_B_c_432_n 0.0432217f $X=7.705 $Y=1.51 $X2=0 $Y2=0
cc_191 N_A_c_175_n N_B_c_432_n 0.0201941f $X=7.885 $Y=1.51 $X2=0 $Y2=0
cc_192 N_A_c_169_n N_B_c_447_n 0.00425878f $X=1.427 $Y=1.75 $X2=0 $Y2=0
cc_193 N_A_c_185_n N_B_c_447_n 0.00105246f $X=1.427 $Y=1.93 $X2=0 $Y2=0
cc_194 N_A_c_198_p N_B_c_447_n 0.00822789f $X=3.5 $Y=2.015 $X2=0 $Y2=0
cc_195 N_A_c_173_n B 3.2027e-19 $X=7.705 $Y=1.51 $X2=0 $Y2=0
cc_196 N_A_c_169_n N_B_c_433_n 6.13387e-19 $X=1.427 $Y=1.75 $X2=0 $Y2=0
cc_197 N_A_c_198_p N_B_c_433_n 0.00171452f $X=3.5 $Y=2.015 $X2=0 $Y2=0
cc_198 N_A_c_186_n N_B_c_433_n 0.0011525f $X=3.665 $Y=1.51 $X2=0 $Y2=0
cc_199 N_A_c_170_n N_B_c_433_n 0.0209654f $X=3.665 $Y=1.51 $X2=0 $Y2=0
cc_200 N_A_c_174_n N_B_c_433_n 0.0197105f $X=1.495 $Y=1.51 $X2=0 $Y2=0
cc_201 N_A_M1039_g N_B_c_434_n 6.70067e-19 $X=7.85 $Y=2.465 $X2=0 $Y2=0
cc_202 N_A_c_173_n N_B_c_434_n 0.00913702f $X=7.705 $Y=1.51 $X2=0 $Y2=0
cc_203 N_A_c_175_n N_B_c_434_n 0.00106839f $X=7.885 $Y=1.51 $X2=0 $Y2=0
cc_204 N_A_M1039_g N_B_c_435_n 0.0380572f $X=7.85 $Y=2.465 $X2=0 $Y2=0
cc_205 N_A_c_173_n N_B_c_435_n 2.71349e-19 $X=7.705 $Y=1.51 $X2=0 $Y2=0
cc_206 N_A_c_175_n N_B_c_435_n 0.0284877f $X=7.885 $Y=1.51 $X2=0 $Y2=0
cc_207 N_A_M1027_g N_A_808_39#_M1001_g 0.021669f $X=3.685 $Y=0.745 $X2=0 $Y2=0
cc_208 N_A_M1037_g N_A_808_39#_M1005_g 0.0447738f $X=3.645 $Y=2.465 $X2=0 $Y2=0
cc_209 N_A_c_186_n N_A_808_39#_M1005_g 0.00165571f $X=3.665 $Y=1.51 $X2=0 $Y2=0
cc_210 N_A_c_188_n N_A_808_39#_M1005_g 0.0113135f $X=6.305 $Y=1.85 $X2=0 $Y2=0
cc_211 N_A_c_190_n N_A_808_39#_M1005_g 9.01012e-19 $X=3.665 $Y=1.85 $X2=0 $Y2=0
cc_212 N_A_c_188_n N_A_808_39#_M1020_g 0.0124709f $X=6.305 $Y=1.85 $X2=0 $Y2=0
cc_213 N_A_c_186_n N_A_808_39#_c_641_n 0.00119154f $X=3.665 $Y=1.51 $X2=0 $Y2=0
cc_214 N_A_c_170_n N_A_808_39#_c_641_n 0.0226938f $X=3.665 $Y=1.51 $X2=0 $Y2=0
cc_215 N_A_c_188_n N_A_808_39#_c_641_n 0.0188613f $X=6.305 $Y=1.85 $X2=0 $Y2=0
cc_216 N_A_c_188_n N_A_808_39#_M1033_g 0.0124305f $X=6.305 $Y=1.85 $X2=0 $Y2=0
cc_217 N_A_M1008_g N_A_808_39#_M1038_g 0.0247242f $X=6.56 $Y=2.465 $X2=0 $Y2=0
cc_218 N_A_c_188_n N_A_808_39#_M1038_g 0.0143409f $X=6.305 $Y=1.85 $X2=0 $Y2=0
cc_219 N_A_c_171_n N_A_808_39#_M1038_g 0.00195518f $X=6.39 $Y=1.765 $X2=0 $Y2=0
cc_220 N_A_c_175_n N_A_808_39#_M1038_g 5.59183e-19 $X=7.885 $Y=1.51 $X2=0 $Y2=0
cc_221 N_A_M1018_g N_A_808_39#_c_643_n 0.0129276f $X=6.515 $Y=0.745 $X2=0 $Y2=0
cc_222 N_A_M1030_g N_A_808_39#_c_643_n 0.0109029f $X=7.025 $Y=0.745 $X2=0 $Y2=0
cc_223 N_A_M1032_g N_A_808_39#_c_643_n 0.0104593f $X=7.455 $Y=0.745 $X2=0 $Y2=0
cc_224 N_A_M1034_g N_A_808_39#_c_643_n 0.0104127f $X=7.885 $Y=0.745 $X2=0 $Y2=0
cc_225 N_A_c_188_n N_A_808_39#_c_643_n 0.00256707f $X=6.305 $Y=1.85 $X2=0 $Y2=0
cc_226 N_A_c_172_n N_A_808_39#_c_643_n 0.0129903f $X=6.475 $Y=1.51 $X2=0 $Y2=0
cc_227 N_A_c_173_n N_A_808_39#_c_643_n 0.0975251f $X=7.705 $Y=1.51 $X2=0 $Y2=0
cc_228 N_A_c_175_n N_A_808_39#_c_643_n 0.0100107f $X=7.885 $Y=1.51 $X2=0 $Y2=0
cc_229 N_A_M1014_g N_A_808_39#_c_658_n 0.0127613f $X=6.99 $Y=2.465 $X2=0 $Y2=0
cc_230 N_A_M1026_g N_A_808_39#_c_658_n 0.0124425f $X=7.42 $Y=2.465 $X2=0 $Y2=0
cc_231 N_A_c_173_n N_A_808_39#_c_658_n 0.0338255f $X=7.705 $Y=1.51 $X2=0 $Y2=0
cc_232 N_A_c_175_n N_A_808_39#_c_658_n 0.00200268f $X=7.885 $Y=1.51 $X2=0 $Y2=0
cc_233 N_A_M1008_g N_A_808_39#_c_659_n 5.2759e-19 $X=6.56 $Y=2.465 $X2=0 $Y2=0
cc_234 N_A_c_188_n N_A_808_39#_c_659_n 0.00552416f $X=6.305 $Y=1.85 $X2=0 $Y2=0
cc_235 N_A_c_173_n N_A_808_39#_c_659_n 0.0131837f $X=7.705 $Y=1.51 $X2=0 $Y2=0
cc_236 N_A_c_175_n N_A_808_39#_c_659_n 0.00205036f $X=7.885 $Y=1.51 $X2=0 $Y2=0
cc_237 N_A_M1039_g N_A_808_39#_c_694_n 0.011933f $X=7.85 $Y=2.465 $X2=0 $Y2=0
cc_238 N_A_c_173_n N_A_808_39#_c_694_n 0.00323873f $X=7.705 $Y=1.51 $X2=0 $Y2=0
cc_239 N_A_M1034_g N_A_808_39#_c_696_n 6.64188e-19 $X=7.885 $Y=0.745 $X2=0 $Y2=0
cc_240 N_A_c_186_n N_A_808_39#_c_647_n 0.0113144f $X=3.665 $Y=1.51 $X2=0 $Y2=0
cc_241 N_A_c_170_n N_A_808_39#_c_647_n 5.83919e-19 $X=3.665 $Y=1.51 $X2=0 $Y2=0
cc_242 N_A_c_188_n N_A_808_39#_c_647_n 0.109113f $X=6.305 $Y=1.85 $X2=0 $Y2=0
cc_243 N_A_M1018_g N_A_808_39#_c_648_n 0.00326483f $X=6.515 $Y=0.745 $X2=0 $Y2=0
cc_244 N_A_c_172_n N_A_808_39#_c_648_n 0.0141739f $X=6.475 $Y=1.51 $X2=0 $Y2=0
cc_245 N_A_M1039_g N_A_808_39#_c_662_n 0.00539797f $X=7.85 $Y=2.465 $X2=0 $Y2=0
cc_246 N_A_c_173_n N_A_808_39#_c_662_n 0.0147861f $X=7.705 $Y=1.51 $X2=0 $Y2=0
cc_247 N_A_c_175_n N_A_808_39#_c_662_n 0.00210954f $X=7.885 $Y=1.51 $X2=0 $Y2=0
cc_248 N_A_M1018_g N_A_808_39#_c_651_n 0.0228714f $X=6.515 $Y=0.745 $X2=0 $Y2=0
cc_249 N_A_c_188_n N_A_808_39#_c_651_n 0.00252705f $X=6.305 $Y=1.85 $X2=0 $Y2=0
cc_250 N_A_c_171_n N_A_808_39#_c_651_n 0.00133779f $X=6.39 $Y=1.765 $X2=0 $Y2=0
cc_251 N_A_c_172_n N_A_808_39#_c_651_n 0.00164025f $X=6.475 $Y=1.51 $X2=0 $Y2=0
cc_252 N_A_c_185_n N_VPWR_M1031_d 0.00124912f $X=1.427 $Y=1.93 $X2=0 $Y2=0
cc_253 N_A_c_286_p N_VPWR_M1031_d 0.00241064f $X=1.57 $Y=2.015 $X2=0 $Y2=0
cc_254 N_A_c_188_n N_VPWR_M1037_d 0.00222395f $X=6.305 $Y=1.85 $X2=0 $Y2=0
cc_255 N_A_c_190_n N_VPWR_M1037_d 7.87838e-19 $X=3.665 $Y=1.85 $X2=0 $Y2=0
cc_256 N_A_c_188_n N_VPWR_M1020_d 0.013029f $X=6.305 $Y=1.85 $X2=0 $Y2=0
cc_257 N_A_c_188_n N_VPWR_M1038_d 0.00207349f $X=6.305 $Y=1.85 $X2=0 $Y2=0
cc_258 N_A_M1019_g N_VPWR_c_870_n 0.0215771f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_259 N_A_M1031_g N_VPWR_c_870_n 0.00217805f $X=0.905 $Y=2.465 $X2=0 $Y2=0
cc_260 N_A_M1037_g N_VPWR_c_871_n 0.0115759f $X=3.645 $Y=2.465 $X2=0 $Y2=0
cc_261 N_A_M1008_g N_VPWR_c_872_n 0.00155004f $X=6.56 $Y=2.465 $X2=0 $Y2=0
cc_262 N_A_c_188_n N_VPWR_c_872_n 0.0122851f $X=6.305 $Y=1.85 $X2=0 $Y2=0
cc_263 N_A_M1008_g N_VPWR_c_873_n 7.34908e-19 $X=6.56 $Y=2.465 $X2=0 $Y2=0
cc_264 N_A_M1014_g N_VPWR_c_873_n 0.0140134f $X=6.99 $Y=2.465 $X2=0 $Y2=0
cc_265 N_A_M1026_g N_VPWR_c_873_n 0.0139215f $X=7.42 $Y=2.465 $X2=0 $Y2=0
cc_266 N_A_M1039_g N_VPWR_c_873_n 7.18684e-19 $X=7.85 $Y=2.465 $X2=0 $Y2=0
cc_267 N_A_M1026_g N_VPWR_c_874_n 0.00486043f $X=7.42 $Y=2.465 $X2=0 $Y2=0
cc_268 N_A_M1039_g N_VPWR_c_874_n 0.00486043f $X=7.85 $Y=2.465 $X2=0 $Y2=0
cc_269 N_A_M1026_g N_VPWR_c_875_n 6.80491e-19 $X=7.42 $Y=2.465 $X2=0 $Y2=0
cc_270 N_A_M1039_g N_VPWR_c_875_n 0.0150429f $X=7.85 $Y=2.465 $X2=0 $Y2=0
cc_271 N_A_M1036_g N_VPWR_c_879_n 0.00461823f $X=1.495 $Y=2.465 $X2=0 $Y2=0
cc_272 N_A_M1037_g N_VPWR_c_879_n 0.00564095f $X=3.645 $Y=2.465 $X2=0 $Y2=0
cc_273 N_A_M1008_g N_VPWR_c_883_n 0.00585385f $X=6.56 $Y=2.465 $X2=0 $Y2=0
cc_274 N_A_M1014_g N_VPWR_c_883_n 0.00486043f $X=6.99 $Y=2.465 $X2=0 $Y2=0
cc_275 N_A_M1019_g N_VPWR_c_885_n 0.00486043f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_276 N_A_M1031_g N_VPWR_c_885_n 0.00462261f $X=0.905 $Y=2.465 $X2=0 $Y2=0
cc_277 N_A_M1031_g N_VPWR_c_889_n 0.00253916f $X=0.905 $Y=2.465 $X2=0 $Y2=0
cc_278 N_A_M1036_g N_VPWR_c_889_n 0.00395787f $X=1.495 $Y=2.465 $X2=0 $Y2=0
cc_279 N_A_M1019_g N_VPWR_c_868_n 0.00835506f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_280 N_A_M1031_g N_VPWR_c_868_n 0.00772963f $X=0.905 $Y=2.465 $X2=0 $Y2=0
cc_281 N_A_M1036_g N_VPWR_c_868_n 0.00775396f $X=1.495 $Y=2.465 $X2=0 $Y2=0
cc_282 N_A_M1037_g N_VPWR_c_868_n 0.00961799f $X=3.645 $Y=2.465 $X2=0 $Y2=0
cc_283 N_A_M1008_g N_VPWR_c_868_n 0.0105614f $X=6.56 $Y=2.465 $X2=0 $Y2=0
cc_284 N_A_M1014_g N_VPWR_c_868_n 0.00824727f $X=6.99 $Y=2.465 $X2=0 $Y2=0
cc_285 N_A_M1026_g N_VPWR_c_868_n 0.00824727f $X=7.42 $Y=2.465 $X2=0 $Y2=0
cc_286 N_A_M1039_g N_VPWR_c_868_n 0.00824727f $X=7.85 $Y=2.465 $X2=0 $Y2=0
cc_287 N_A_c_198_p N_A_110_367#_M1036_s 0.00810274f $X=3.5 $Y=2.015 $X2=0 $Y2=0
cc_288 N_A_c_198_p N_A_110_367#_M1012_d 0.00323209f $X=3.5 $Y=2.015 $X2=0 $Y2=0
cc_289 N_A_c_198_p N_A_110_367#_M1022_d 0.00363947f $X=3.5 $Y=2.015 $X2=0 $Y2=0
cc_290 N_A_c_190_n N_A_110_367#_M1022_d 0.0014725f $X=3.665 $Y=1.85 $X2=0 $Y2=0
cc_291 N_A_M1031_g N_A_110_367#_c_1030_n 5.49162e-19 $X=0.905 $Y=2.465 $X2=0
+ $Y2=0
cc_292 N_A_M1036_g N_A_110_367#_c_1030_n 0.00508048f $X=1.495 $Y=2.465 $X2=0
+ $Y2=0
cc_293 N_A_M1031_g N_A_110_367#_c_1032_n 0.00527951f $X=0.905 $Y=2.465 $X2=0
+ $Y2=0
cc_294 N_A_M1036_g N_A_110_367#_c_1032_n 5.06159e-19 $X=1.495 $Y=2.465 $X2=0
+ $Y2=0
cc_295 N_A_M1031_g N_A_110_367#_c_1034_n 0.00848239f $X=0.905 $Y=2.465 $X2=0
+ $Y2=0
cc_296 N_A_M1036_g N_A_110_367#_c_1034_n 0.00750559f $X=1.495 $Y=2.465 $X2=0
+ $Y2=0
cc_297 N_A_c_198_p N_Y_M1002_s 0.00326293f $X=3.5 $Y=2.015 $X2=0 $Y2=0
cc_298 N_A_c_198_p N_Y_M1013_s 0.00323209f $X=3.5 $Y=2.015 $X2=0 $Y2=0
cc_299 N_A_c_188_n N_Y_M1005_s 0.00176461f $X=6.305 $Y=1.85 $X2=0 $Y2=0
cc_300 N_A_c_188_n N_Y_M1033_s 0.00176461f $X=6.305 $Y=1.85 $X2=0 $Y2=0
cc_301 N_A_M1006_g N_Y_c_1063_n 0.00343071f $X=0.515 $Y=0.745 $X2=0 $Y2=0
cc_302 A N_Y_c_1063_n 0.0266782f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_303 N_A_c_174_n N_Y_c_1063_n 0.0179552f $X=1.495 $Y=1.51 $X2=0 $Y2=0
cc_304 N_A_M1006_g N_Y_c_1064_n 0.0124948f $X=0.515 $Y=0.745 $X2=0 $Y2=0
cc_305 N_A_M1017_g N_Y_c_1064_n 0.0109362f $X=1.025 $Y=0.745 $X2=0 $Y2=0
cc_306 N_A_M1024_g N_Y_c_1064_n 0.0104398f $X=1.455 $Y=0.745 $X2=0 $Y2=0
cc_307 N_A_M1027_g N_Y_c_1064_n 0.010789f $X=3.685 $Y=0.745 $X2=0 $Y2=0
cc_308 N_A_c_169_n N_Y_c_1064_n 0.0222295f $X=1.427 $Y=1.75 $X2=0 $Y2=0
cc_309 N_A_c_186_n N_Y_c_1064_n 0.0240115f $X=3.665 $Y=1.51 $X2=0 $Y2=0
cc_310 N_A_c_170_n N_Y_c_1064_n 0.00458374f $X=3.665 $Y=1.51 $X2=0 $Y2=0
cc_311 N_A_c_188_n N_Y_c_1064_n 0.00325319f $X=6.305 $Y=1.85 $X2=0 $Y2=0
cc_312 A N_Y_c_1064_n 0.0620646f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_313 N_A_c_174_n N_Y_c_1064_n 0.00984183f $X=1.495 $Y=1.51 $X2=0 $Y2=0
cc_314 N_A_M1019_g N_Y_c_1087_n 0.0162717f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_315 N_A_M1031_g N_Y_c_1087_n 0.0110854f $X=0.905 $Y=2.465 $X2=0 $Y2=0
cc_316 N_A_M1036_g N_Y_c_1087_n 5.53723e-19 $X=1.495 $Y=2.465 $X2=0 $Y2=0
cc_317 N_A_c_185_n N_Y_c_1087_n 8.035e-19 $X=1.427 $Y=1.93 $X2=0 $Y2=0
cc_318 N_A_c_286_p N_Y_c_1087_n 0.0144257f $X=1.57 $Y=2.015 $X2=0 $Y2=0
cc_319 A N_Y_c_1087_n 0.0451815f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_320 N_A_c_174_n N_Y_c_1087_n 8.57757e-19 $X=1.495 $Y=1.51 $X2=0 $Y2=0
cc_321 N_A_M1019_g N_Y_c_1094_n 8.79042e-19 $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_322 N_A_M1031_g N_Y_c_1094_n 0.00500789f $X=0.905 $Y=2.465 $X2=0 $Y2=0
cc_323 N_A_M1036_g N_Y_c_1094_n 0.00321615f $X=1.495 $Y=2.465 $X2=0 $Y2=0
cc_324 N_A_c_286_p N_Y_c_1094_n 7.77101e-19 $X=1.57 $Y=2.015 $X2=0 $Y2=0
cc_325 N_A_M1036_g N_Y_c_1098_n 0.0116766f $X=1.495 $Y=2.465 $X2=0 $Y2=0
cc_326 N_A_M1037_g N_Y_c_1098_n 0.01575f $X=3.645 $Y=2.465 $X2=0 $Y2=0
cc_327 N_A_c_198_p N_Y_c_1098_n 0.0977584f $X=3.5 $Y=2.015 $X2=0 $Y2=0
cc_328 N_A_c_286_p N_Y_c_1098_n 0.0178078f $X=1.57 $Y=2.015 $X2=0 $Y2=0
cc_329 N_A_c_170_n N_Y_c_1098_n 4.568e-19 $X=3.665 $Y=1.51 $X2=0 $Y2=0
cc_330 N_A_c_188_n N_Y_c_1098_n 0.010272f $X=6.305 $Y=1.85 $X2=0 $Y2=0
cc_331 N_A_c_190_n N_Y_c_1098_n 0.0126842f $X=3.665 $Y=1.85 $X2=0 $Y2=0
cc_332 A N_Y_c_1098_n 0.00595256f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_333 N_A_c_174_n N_Y_c_1098_n 9.51513e-19 $X=1.495 $Y=1.51 $X2=0 $Y2=0
cc_334 N_A_M1019_g N_Y_c_1107_n 5.36358e-19 $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_335 N_A_M1031_g N_Y_c_1107_n 0.00676893f $X=0.905 $Y=2.465 $X2=0 $Y2=0
cc_336 N_A_c_188_n N_Y_c_1109_n 0.0707086f $X=6.305 $Y=1.85 $X2=0 $Y2=0
cc_337 N_A_c_188_n N_Y_c_1110_n 0.0144401f $X=6.305 $Y=1.85 $X2=0 $Y2=0
cc_338 N_A_M1037_g N_Y_c_1111_n 8.73981e-19 $X=3.645 $Y=2.465 $X2=0 $Y2=0
cc_339 N_A_c_188_n N_Y_c_1111_n 0.02498f $X=6.305 $Y=1.85 $X2=0 $Y2=0
cc_340 N_A_M1006_g N_A_31_65#_c_1206_n 0.00683735f $X=0.515 $Y=0.745 $X2=0 $Y2=0
cc_341 N_A_M1017_g N_A_31_65#_c_1206_n 6.84198e-19 $X=1.025 $Y=0.745 $X2=0 $Y2=0
cc_342 N_A_M1006_g N_A_31_65#_c_1218_n 0.00920546f $X=0.515 $Y=0.745 $X2=0 $Y2=0
cc_343 N_A_M1017_g N_A_31_65#_c_1218_n 0.0103828f $X=1.025 $Y=0.745 $X2=0 $Y2=0
cc_344 N_A_M1006_g N_A_31_65#_c_1207_n 6.58326e-19 $X=0.515 $Y=0.745 $X2=0 $Y2=0
cc_345 N_A_M1017_g N_A_31_65#_c_1208_n 2.89865e-19 $X=1.025 $Y=0.745 $X2=0 $Y2=0
cc_346 N_A_M1024_g N_A_31_65#_c_1208_n 2.8404e-19 $X=1.455 $Y=0.745 $X2=0 $Y2=0
cc_347 N_A_M1024_g N_A_31_65#_c_1223_n 0.00977853f $X=1.455 $Y=0.745 $X2=0 $Y2=0
cc_348 N_A_M1027_g N_A_31_65#_c_1224_n 0.00987455f $X=3.685 $Y=0.745 $X2=0 $Y2=0
cc_349 N_A_M1027_g N_A_31_65#_c_1225_n 0.00463764f $X=3.685 $Y=0.745 $X2=0 $Y2=0
cc_350 N_A_M1027_g N_A_31_65#_c_1212_n 0.00286088f $X=3.685 $Y=0.745 $X2=0 $Y2=0
cc_351 N_A_M1018_g N_A_31_65#_c_1213_n 0.00172249f $X=6.515 $Y=0.745 $X2=0 $Y2=0
cc_352 N_A_M1006_g N_VGND_c_1326_n 0.0041164f $X=0.515 $Y=0.745 $X2=0 $Y2=0
cc_353 N_A_M1017_g N_VGND_c_1326_n 0.00613738f $X=1.025 $Y=0.745 $X2=0 $Y2=0
cc_354 N_A_M1024_g N_VGND_c_1326_n 3.61965e-19 $X=1.455 $Y=0.745 $X2=0 $Y2=0
cc_355 N_A_M1017_g N_VGND_c_1327_n 3.61976e-19 $X=1.025 $Y=0.745 $X2=0 $Y2=0
cc_356 N_A_M1024_g N_VGND_c_1327_n 0.00651658f $X=1.455 $Y=0.745 $X2=0 $Y2=0
cc_357 N_A_M1027_g N_VGND_c_1329_n 0.00326924f $X=3.685 $Y=0.745 $X2=0 $Y2=0
cc_358 N_A_M1018_g N_VGND_c_1330_n 0.00436824f $X=6.515 $Y=0.745 $X2=0 $Y2=0
cc_359 N_A_M1030_g N_VGND_c_1330_n 0.00610259f $X=7.025 $Y=0.745 $X2=0 $Y2=0
cc_360 N_A_M1032_g N_VGND_c_1330_n 3.56287e-19 $X=7.455 $Y=0.745 $X2=0 $Y2=0
cc_361 N_A_M1030_g N_VGND_c_1331_n 3.64805e-19 $X=7.025 $Y=0.745 $X2=0 $Y2=0
cc_362 N_A_M1032_g N_VGND_c_1331_n 0.00665361f $X=7.455 $Y=0.745 $X2=0 $Y2=0
cc_363 N_A_M1034_g N_VGND_c_1331_n 0.00683027f $X=7.885 $Y=0.745 $X2=0 $Y2=0
cc_364 N_A_M1027_g N_VGND_c_1336_n 0.0035672f $X=3.685 $Y=0.745 $X2=0 $Y2=0
cc_365 N_A_M1018_g N_VGND_c_1336_n 0.0036024f $X=6.515 $Y=0.745 $X2=0 $Y2=0
cc_366 N_A_M1030_g N_VGND_c_1338_n 0.00331181f $X=7.025 $Y=0.745 $X2=0 $Y2=0
cc_367 N_A_M1032_g N_VGND_c_1338_n 0.00306601f $X=7.455 $Y=0.745 $X2=0 $Y2=0
cc_368 N_A_M1006_g N_VGND_c_1340_n 0.00359072f $X=0.515 $Y=0.745 $X2=0 $Y2=0
cc_369 N_A_M1017_g N_VGND_c_1341_n 0.003302f $X=1.025 $Y=0.745 $X2=0 $Y2=0
cc_370 N_A_M1024_g N_VGND_c_1341_n 0.00305694f $X=1.455 $Y=0.745 $X2=0 $Y2=0
cc_371 N_A_M1034_g N_VGND_c_1342_n 0.00306601f $X=7.885 $Y=0.745 $X2=0 $Y2=0
cc_372 N_A_M1006_g N_VGND_c_1343_n 0.00537318f $X=0.515 $Y=0.745 $X2=0 $Y2=0
cc_373 N_A_M1017_g N_VGND_c_1343_n 0.00422442f $X=1.025 $Y=0.745 $X2=0 $Y2=0
cc_374 N_A_M1024_g N_VGND_c_1343_n 0.00391883f $X=1.455 $Y=0.745 $X2=0 $Y2=0
cc_375 N_A_M1027_g N_VGND_c_1343_n 0.00504476f $X=3.685 $Y=0.745 $X2=0 $Y2=0
cc_376 N_A_M1018_g N_VGND_c_1343_n 0.00552236f $X=6.515 $Y=0.745 $X2=0 $Y2=0
cc_377 N_A_M1030_g N_VGND_c_1343_n 0.00424707f $X=7.025 $Y=0.745 $X2=0 $Y2=0
cc_378 N_A_M1032_g N_VGND_c_1343_n 0.00393982f $X=7.455 $Y=0.745 $X2=0 $Y2=0
cc_379 N_A_M1034_g N_VGND_c_1343_n 0.00394956f $X=7.885 $Y=0.745 $X2=0 $Y2=0
cc_380 N_A_M1018_g N_A_1235_65#_c_1483_n 0.00674466f $X=6.515 $Y=0.745 $X2=0
+ $Y2=0
cc_381 N_A_M1030_g N_A_1235_65#_c_1483_n 4.39148e-19 $X=7.025 $Y=0.745 $X2=0
+ $Y2=0
cc_382 N_A_M1018_g N_A_1235_65#_c_1493_n 0.00923879f $X=6.515 $Y=0.745 $X2=0
+ $Y2=0
cc_383 N_A_M1030_g N_A_1235_65#_c_1493_n 0.0104189f $X=7.025 $Y=0.745 $X2=0
+ $Y2=0
cc_384 N_A_M1018_g N_A_1235_65#_c_1484_n 7.16038e-19 $X=6.515 $Y=0.745 $X2=0
+ $Y2=0
cc_385 N_A_M1030_g N_A_1235_65#_c_1485_n 2.92907e-19 $X=7.025 $Y=0.745 $X2=0
+ $Y2=0
cc_386 N_A_M1032_g N_A_1235_65#_c_1485_n 2.86798e-19 $X=7.455 $Y=0.745 $X2=0
+ $Y2=0
cc_387 N_A_M1032_g N_A_1235_65#_c_1498_n 0.00981198f $X=7.455 $Y=0.745 $X2=0
+ $Y2=0
cc_388 N_A_M1034_g N_A_1235_65#_c_1498_n 0.00985855f $X=7.885 $Y=0.745 $X2=0
+ $Y2=0
cc_389 N_A_M1034_g N_A_1235_65#_c_1487_n 0.00104712f $X=7.885 $Y=0.745 $X2=0
+ $Y2=0
cc_390 N_B_c_432_n N_A_808_39#_M1005_g 0.00256215f $X=8.255 $Y=1.665 $X2=0 $Y2=0
cc_391 N_B_c_432_n N_A_808_39#_M1020_g 0.00321596f $X=8.255 $Y=1.665 $X2=0 $Y2=0
cc_392 N_B_c_432_n N_A_808_39#_c_640_n 0.00694764f $X=8.255 $Y=1.665 $X2=0 $Y2=0
cc_393 N_B_c_432_n N_A_808_39#_c_641_n 0.0157441f $X=8.255 $Y=1.665 $X2=0 $Y2=0
cc_394 N_B_c_432_n N_A_808_39#_M1033_g 0.00321596f $X=8.255 $Y=1.665 $X2=0 $Y2=0
cc_395 N_B_c_432_n N_A_808_39#_M1038_g 0.00253168f $X=8.255 $Y=1.665 $X2=0 $Y2=0
cc_396 N_B_M1004_g N_A_808_39#_c_643_n 0.00911078f $X=8.315 $Y=0.745 $X2=0 $Y2=0
cc_397 N_B_c_432_n N_A_808_39#_c_643_n 0.0148652f $X=8.255 $Y=1.665 $X2=0 $Y2=0
cc_398 B N_A_808_39#_c_643_n 5.66826e-19 $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_399 N_B_c_434_n N_A_808_39#_c_643_n 0.00830555f $X=9.425 $Y=1.51 $X2=0 $Y2=0
cc_400 N_B_c_435_n N_A_808_39#_c_643_n 9.10663e-19 $X=9.57 $Y=1.535 $X2=0 $Y2=0
cc_401 N_B_c_432_n N_A_808_39#_c_658_n 0.0184461f $X=8.255 $Y=1.665 $X2=0 $Y2=0
cc_402 N_B_c_432_n N_A_808_39#_c_659_n 0.00691665f $X=8.255 $Y=1.665 $X2=0 $Y2=0
cc_403 N_B_c_440_n N_A_808_39#_c_694_n 0.012412f $X=8.28 $Y=1.725 $X2=0 $Y2=0
cc_404 N_B_c_432_n N_A_808_39#_c_694_n 0.012411f $X=8.255 $Y=1.665 $X2=0 $Y2=0
cc_405 B N_A_808_39#_c_694_n 0.00367942f $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_406 N_B_c_434_n N_A_808_39#_c_694_n 0.00854305f $X=9.425 $Y=1.51 $X2=0 $Y2=0
cc_407 N_B_M1004_g N_A_808_39#_c_696_n 0.00607153f $X=8.315 $Y=0.745 $X2=0 $Y2=0
cc_408 N_B_M1015_g N_A_808_39#_c_696_n 0.00611576f $X=8.745 $Y=0.745 $X2=0 $Y2=0
cc_409 N_B_M1025_g N_A_808_39#_c_696_n 5.14064e-19 $X=9.175 $Y=0.745 $X2=0 $Y2=0
cc_410 N_B_c_441_n N_A_808_39#_c_729_n 0.0122595f $X=8.71 $Y=1.725 $X2=0 $Y2=0
cc_411 N_B_c_442_n N_A_808_39#_c_729_n 0.0122595f $X=9.14 $Y=1.725 $X2=0 $Y2=0
cc_412 N_B_c_434_n N_A_808_39#_c_729_n 0.0427275f $X=9.425 $Y=1.51 $X2=0 $Y2=0
cc_413 N_B_c_435_n N_A_808_39#_c_729_n 6.53383e-19 $X=9.57 $Y=1.535 $X2=0 $Y2=0
cc_414 N_B_M1015_g N_A_808_39#_c_644_n 0.00963507f $X=8.745 $Y=0.745 $X2=0 $Y2=0
cc_415 N_B_M1025_g N_A_808_39#_c_644_n 0.00966333f $X=9.175 $Y=0.745 $X2=0 $Y2=0
cc_416 N_B_c_434_n N_A_808_39#_c_644_n 0.0391098f $X=9.425 $Y=1.51 $X2=0 $Y2=0
cc_417 N_B_c_435_n N_A_808_39#_c_644_n 0.00266877f $X=9.57 $Y=1.535 $X2=0 $Y2=0
cc_418 N_B_M1015_g N_A_808_39#_c_737_n 5.14064e-19 $X=8.745 $Y=0.745 $X2=0 $Y2=0
cc_419 N_B_M1025_g N_A_808_39#_c_737_n 0.00612526f $X=9.175 $Y=0.745 $X2=0 $Y2=0
cc_420 N_B_M1028_g N_A_808_39#_c_737_n 0.0106545f $X=9.605 $Y=0.745 $X2=0 $Y2=0
cc_421 N_B_c_443_n N_A_808_39#_c_660_n 0.0145491f $X=9.57 $Y=1.725 $X2=0 $Y2=0
cc_422 N_B_c_434_n N_A_808_39#_c_660_n 0.00861123f $X=9.425 $Y=1.51 $X2=0 $Y2=0
cc_423 N_B_M1028_g N_A_808_39#_c_645_n 0.012425f $X=9.605 $Y=0.745 $X2=0 $Y2=0
cc_424 N_B_c_434_n N_A_808_39#_c_645_n 0.00248238f $X=9.425 $Y=1.51 $X2=0 $Y2=0
cc_425 N_B_M1028_g N_A_808_39#_c_646_n 0.0144684f $X=9.605 $Y=0.745 $X2=0 $Y2=0
cc_426 N_B_c_434_n N_A_808_39#_c_646_n 0.0251396f $X=9.425 $Y=1.51 $X2=0 $Y2=0
cc_427 N_B_c_435_n N_A_808_39#_c_646_n 0.00819324f $X=9.57 $Y=1.535 $X2=0 $Y2=0
cc_428 N_B_c_432_n N_A_808_39#_c_647_n 0.0552874f $X=8.255 $Y=1.665 $X2=0 $Y2=0
cc_429 N_B_c_440_n N_A_808_39#_c_662_n 7.90905e-19 $X=8.28 $Y=1.725 $X2=0 $Y2=0
cc_430 N_B_c_432_n N_A_808_39#_c_662_n 0.00777635f $X=8.255 $Y=1.665 $X2=0 $Y2=0
cc_431 N_B_M1004_g N_A_808_39#_c_649_n 0.00219079f $X=8.315 $Y=0.745 $X2=0 $Y2=0
cc_432 N_B_M1015_g N_A_808_39#_c_649_n 0.00184788f $X=8.745 $Y=0.745 $X2=0 $Y2=0
cc_433 B N_A_808_39#_c_649_n 0.00111726f $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_434 N_B_c_434_n N_A_808_39#_c_649_n 0.0263082f $X=9.425 $Y=1.51 $X2=0 $Y2=0
cc_435 N_B_c_435_n N_A_808_39#_c_649_n 0.00275564f $X=9.57 $Y=1.535 $X2=0 $Y2=0
cc_436 B N_A_808_39#_c_755_n 0.00426309f $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_437 N_B_c_434_n N_A_808_39#_c_755_n 0.013394f $X=9.425 $Y=1.51 $X2=0 $Y2=0
cc_438 N_B_c_435_n N_A_808_39#_c_755_n 7.3596e-19 $X=9.57 $Y=1.535 $X2=0 $Y2=0
cc_439 N_B_M1025_g N_A_808_39#_c_650_n 0.00184788f $X=9.175 $Y=0.745 $X2=0 $Y2=0
cc_440 N_B_M1028_g N_A_808_39#_c_650_n 0.00184788f $X=9.605 $Y=0.745 $X2=0 $Y2=0
cc_441 N_B_c_434_n N_A_808_39#_c_650_n 0.0274411f $X=9.425 $Y=1.51 $X2=0 $Y2=0
cc_442 N_B_c_435_n N_A_808_39#_c_650_n 0.00275564f $X=9.57 $Y=1.535 $X2=0 $Y2=0
cc_443 N_B_c_434_n N_A_808_39#_c_762_n 0.0153756f $X=9.425 $Y=1.51 $X2=0 $Y2=0
cc_444 N_B_c_435_n N_A_808_39#_c_762_n 7.3596e-19 $X=9.57 $Y=1.535 $X2=0 $Y2=0
cc_445 N_B_c_432_n N_A_808_39#_c_651_n 0.0113989f $X=8.255 $Y=1.665 $X2=0 $Y2=0
cc_446 N_B_M1022_g N_VPWR_c_871_n 0.00156628f $X=3.215 $Y=2.465 $X2=0 $Y2=0
cc_447 N_B_c_432_n N_VPWR_c_872_n 0.00108767f $X=8.255 $Y=1.665 $X2=0 $Y2=0
cc_448 N_B_c_440_n N_VPWR_c_875_n 0.0150429f $X=8.28 $Y=1.725 $X2=0 $Y2=0
cc_449 N_B_c_441_n N_VPWR_c_875_n 6.80491e-19 $X=8.71 $Y=1.725 $X2=0 $Y2=0
cc_450 N_B_c_440_n N_VPWR_c_876_n 6.80491e-19 $X=8.28 $Y=1.725 $X2=0 $Y2=0
cc_451 N_B_c_441_n N_VPWR_c_876_n 0.0151398f $X=8.71 $Y=1.725 $X2=0 $Y2=0
cc_452 N_B_c_442_n N_VPWR_c_876_n 0.0151398f $X=9.14 $Y=1.725 $X2=0 $Y2=0
cc_453 N_B_c_443_n N_VPWR_c_876_n 6.80491e-19 $X=9.57 $Y=1.725 $X2=0 $Y2=0
cc_454 N_B_c_442_n N_VPWR_c_878_n 6.80491e-19 $X=9.14 $Y=1.725 $X2=0 $Y2=0
cc_455 N_B_c_443_n N_VPWR_c_878_n 0.0175702f $X=9.57 $Y=1.725 $X2=0 $Y2=0
cc_456 N_B_M1002_g N_VPWR_c_879_n 0.00380755f $X=1.925 $Y=2.465 $X2=0 $Y2=0
cc_457 N_B_M1012_g N_VPWR_c_879_n 0.00380755f $X=2.355 $Y=2.465 $X2=0 $Y2=0
cc_458 N_B_M1013_g N_VPWR_c_879_n 0.00380755f $X=2.785 $Y=2.465 $X2=0 $Y2=0
cc_459 N_B_M1022_g N_VPWR_c_879_n 0.00380755f $X=3.215 $Y=2.465 $X2=0 $Y2=0
cc_460 N_B_c_440_n N_VPWR_c_887_n 0.00486043f $X=8.28 $Y=1.725 $X2=0 $Y2=0
cc_461 N_B_c_441_n N_VPWR_c_887_n 0.00486043f $X=8.71 $Y=1.725 $X2=0 $Y2=0
cc_462 N_B_c_442_n N_VPWR_c_888_n 0.00486043f $X=9.14 $Y=1.725 $X2=0 $Y2=0
cc_463 N_B_c_443_n N_VPWR_c_888_n 0.00486043f $X=9.57 $Y=1.725 $X2=0 $Y2=0
cc_464 N_B_M1002_g N_VPWR_c_868_n 0.005529f $X=1.925 $Y=2.465 $X2=0 $Y2=0
cc_465 N_B_M1012_g N_VPWR_c_868_n 0.00550172f $X=2.355 $Y=2.465 $X2=0 $Y2=0
cc_466 N_B_M1013_g N_VPWR_c_868_n 0.00550172f $X=2.785 $Y=2.465 $X2=0 $Y2=0
cc_467 N_B_M1022_g N_VPWR_c_868_n 0.005529f $X=3.215 $Y=2.465 $X2=0 $Y2=0
cc_468 N_B_c_440_n N_VPWR_c_868_n 0.00824727f $X=8.28 $Y=1.725 $X2=0 $Y2=0
cc_469 N_B_c_441_n N_VPWR_c_868_n 0.00824727f $X=8.71 $Y=1.725 $X2=0 $Y2=0
cc_470 N_B_c_442_n N_VPWR_c_868_n 0.00824727f $X=9.14 $Y=1.725 $X2=0 $Y2=0
cc_471 N_B_c_443_n N_VPWR_c_868_n 0.00824727f $X=9.57 $Y=1.725 $X2=0 $Y2=0
cc_472 N_B_M1002_g N_A_110_367#_c_1030_n 0.00142813f $X=1.925 $Y=2.465 $X2=0
+ $Y2=0
cc_473 N_B_M1002_g N_A_110_367#_c_1037_n 0.0114157f $X=1.925 $Y=2.465 $X2=0
+ $Y2=0
cc_474 N_B_M1012_g N_A_110_367#_c_1037_n 0.0129034f $X=2.355 $Y=2.465 $X2=0
+ $Y2=0
cc_475 N_B_M1013_g N_A_110_367#_c_1037_n 0.0128097f $X=2.785 $Y=2.465 $X2=0
+ $Y2=0
cc_476 N_B_M1022_g N_A_110_367#_c_1037_n 0.0129034f $X=3.215 $Y=2.465 $X2=0
+ $Y2=0
cc_477 N_B_M1000_g N_Y_c_1064_n 0.0104398f $X=1.885 $Y=0.745 $X2=0 $Y2=0
cc_478 N_B_M1003_g N_Y_c_1064_n 0.0104512f $X=2.315 $Y=0.745 $X2=0 $Y2=0
cc_479 N_B_M1011_g N_Y_c_1064_n 0.0104613f $X=2.745 $Y=0.745 $X2=0 $Y2=0
cc_480 N_B_M1023_g N_Y_c_1064_n 0.0113345f $X=3.175 $Y=0.745 $X2=0 $Y2=0
cc_481 N_B_c_431_n N_Y_c_1064_n 0.0414865f $X=2.41 $Y=1.582 $X2=0 $Y2=0
cc_482 N_B_c_445_n N_Y_c_1064_n 0.0523751f $X=2.995 $Y=1.51 $X2=0 $Y2=0
cc_483 N_B_c_432_n N_Y_c_1064_n 0.0235128f $X=8.255 $Y=1.665 $X2=0 $Y2=0
cc_484 N_B_c_447_n N_Y_c_1064_n 0.00155525f $X=2.305 $Y=1.665 $X2=0 $Y2=0
cc_485 N_B_c_433_n N_Y_c_1064_n 0.0092909f $X=3.175 $Y=1.51 $X2=0 $Y2=0
cc_486 N_B_M1002_g N_Y_c_1098_n 0.00866338f $X=1.925 $Y=2.465 $X2=0 $Y2=0
cc_487 N_B_M1012_g N_Y_c_1098_n 0.00870325f $X=2.355 $Y=2.465 $X2=0 $Y2=0
cc_488 N_B_M1013_g N_Y_c_1098_n 0.0087038f $X=2.785 $Y=2.465 $X2=0 $Y2=0
cc_489 N_B_M1022_g N_Y_c_1098_n 0.00865446f $X=3.215 $Y=2.465 $X2=0 $Y2=0
cc_490 N_B_c_432_n N_Y_c_1098_n 0.00280171f $X=8.255 $Y=1.665 $X2=0 $Y2=0
cc_491 N_B_M1000_g N_A_31_65#_c_1223_n 0.00977853f $X=1.885 $Y=0.745 $X2=0 $Y2=0
cc_492 N_B_M1000_g N_A_31_65#_c_1209_n 2.85448e-19 $X=1.885 $Y=0.745 $X2=0 $Y2=0
cc_493 N_B_M1003_g N_A_31_65#_c_1209_n 2.85448e-19 $X=2.315 $Y=0.745 $X2=0 $Y2=0
cc_494 N_B_M1003_g N_A_31_65#_c_1231_n 0.00982509f $X=2.315 $Y=0.745 $X2=0 $Y2=0
cc_495 N_B_M1011_g N_A_31_65#_c_1231_n 0.00982509f $X=2.745 $Y=0.745 $X2=0 $Y2=0
cc_496 N_B_M1011_g N_A_31_65#_c_1210_n 2.85448e-19 $X=2.745 $Y=0.745 $X2=0 $Y2=0
cc_497 N_B_M1023_g N_A_31_65#_c_1210_n 2.85448e-19 $X=3.175 $Y=0.745 $X2=0 $Y2=0
cc_498 N_B_M1023_g N_A_31_65#_c_1224_n 0.0102064f $X=3.175 $Y=0.745 $X2=0 $Y2=0
cc_499 N_B_M1023_g N_A_31_65#_c_1225_n 6.08169e-19 $X=3.175 $Y=0.745 $X2=0 $Y2=0
cc_500 N_B_M1000_g N_VGND_c_1327_n 0.00650228f $X=1.885 $Y=0.745 $X2=0 $Y2=0
cc_501 N_B_M1003_g N_VGND_c_1327_n 3.60064e-19 $X=2.315 $Y=0.745 $X2=0 $Y2=0
cc_502 N_B_M1000_g N_VGND_c_1328_n 3.60064e-19 $X=1.885 $Y=0.745 $X2=0 $Y2=0
cc_503 N_B_M1003_g N_VGND_c_1328_n 0.00653804f $X=2.315 $Y=0.745 $X2=0 $Y2=0
cc_504 N_B_M1011_g N_VGND_c_1328_n 0.00653804f $X=2.745 $Y=0.745 $X2=0 $Y2=0
cc_505 N_B_M1023_g N_VGND_c_1328_n 3.60064e-19 $X=3.175 $Y=0.745 $X2=0 $Y2=0
cc_506 N_B_M1011_g N_VGND_c_1329_n 3.60064e-19 $X=2.745 $Y=0.745 $X2=0 $Y2=0
cc_507 N_B_M1023_g N_VGND_c_1329_n 0.00657168f $X=3.175 $Y=0.745 $X2=0 $Y2=0
cc_508 N_B_M1004_g N_VGND_c_1331_n 6.09758e-19 $X=8.315 $Y=0.745 $X2=0 $Y2=0
cc_509 N_B_M1000_g N_VGND_c_1332_n 0.00305694f $X=1.885 $Y=0.745 $X2=0 $Y2=0
cc_510 N_B_M1003_g N_VGND_c_1332_n 0.00305694f $X=2.315 $Y=0.745 $X2=0 $Y2=0
cc_511 N_B_M1011_g N_VGND_c_1334_n 0.00305694f $X=2.745 $Y=0.745 $X2=0 $Y2=0
cc_512 N_B_M1023_g N_VGND_c_1334_n 0.00305694f $X=3.175 $Y=0.745 $X2=0 $Y2=0
cc_513 N_B_M1004_g N_VGND_c_1342_n 0.00302501f $X=8.315 $Y=0.745 $X2=0 $Y2=0
cc_514 N_B_M1015_g N_VGND_c_1342_n 0.00302501f $X=8.745 $Y=0.745 $X2=0 $Y2=0
cc_515 N_B_M1025_g N_VGND_c_1342_n 0.00302501f $X=9.175 $Y=0.745 $X2=0 $Y2=0
cc_516 N_B_M1028_g N_VGND_c_1342_n 0.00302501f $X=9.605 $Y=0.745 $X2=0 $Y2=0
cc_517 N_B_M1000_g N_VGND_c_1343_n 0.00391883f $X=1.885 $Y=0.745 $X2=0 $Y2=0
cc_518 N_B_M1003_g N_VGND_c_1343_n 0.00391883f $X=2.315 $Y=0.745 $X2=0 $Y2=0
cc_519 N_B_M1011_g N_VGND_c_1343_n 0.00391883f $X=2.745 $Y=0.745 $X2=0 $Y2=0
cc_520 N_B_M1023_g N_VGND_c_1343_n 0.00391883f $X=3.175 $Y=0.745 $X2=0 $Y2=0
cc_521 N_B_M1004_g N_VGND_c_1343_n 0.00435646f $X=8.315 $Y=0.745 $X2=0 $Y2=0
cc_522 N_B_M1015_g N_VGND_c_1343_n 0.00434671f $X=8.745 $Y=0.745 $X2=0 $Y2=0
cc_523 N_B_M1025_g N_VGND_c_1343_n 0.00434671f $X=9.175 $Y=0.745 $X2=0 $Y2=0
cc_524 N_B_M1028_g N_VGND_c_1343_n 0.00470541f $X=9.605 $Y=0.745 $X2=0 $Y2=0
cc_525 N_B_M1004_g N_A_1235_65#_c_1486_n 0.0111391f $X=8.315 $Y=0.745 $X2=0
+ $Y2=0
cc_526 N_B_M1015_g N_A_1235_65#_c_1486_n 0.0114881f $X=8.745 $Y=0.745 $X2=0
+ $Y2=0
cc_527 N_B_M1025_g N_A_1235_65#_c_1488_n 0.0112092f $X=9.175 $Y=0.745 $X2=0
+ $Y2=0
cc_528 N_B_M1028_g N_A_1235_65#_c_1488_n 0.0125968f $X=9.605 $Y=0.745 $X2=0
+ $Y2=0
cc_529 N_A_808_39#_c_658_n N_VPWR_M1014_d 0.00180746f $X=7.54 $Y=1.86 $X2=0
+ $Y2=0
cc_530 N_A_808_39#_c_694_n N_VPWR_M1039_d 0.00448889f $X=8.4 $Y=2.005 $X2=0
+ $Y2=0
cc_531 N_A_808_39#_c_729_n N_VPWR_M1016_s 0.00331217f $X=9.26 $Y=2.005 $X2=0
+ $Y2=0
cc_532 N_A_808_39#_c_660_n N_VPWR_M1035_s 0.00438662f $X=9.77 $Y=2.005 $X2=0
+ $Y2=0
cc_533 N_A_808_39#_c_646_n N_VPWR_M1035_s 0.00137373f $X=9.88 $Y=1.92 $X2=0
+ $Y2=0
cc_534 N_A_808_39#_M1005_g N_VPWR_c_871_n 0.0106578f $X=4.115 $Y=2.465 $X2=0
+ $Y2=0
cc_535 N_A_808_39#_M1020_g N_VPWR_c_871_n 0.00105111f $X=4.545 $Y=2.465 $X2=0
+ $Y2=0
cc_536 N_A_808_39#_M1038_g N_VPWR_c_872_n 0.00146828f $X=6.13 $Y=2.465 $X2=0
+ $Y2=0
cc_537 N_A_808_39#_c_658_n N_VPWR_c_873_n 0.0153048f $X=7.54 $Y=1.86 $X2=0 $Y2=0
cc_538 N_A_808_39#_c_774_p N_VPWR_c_874_n 0.0124525f $X=7.635 $Y=2.45 $X2=0
+ $Y2=0
cc_539 N_A_808_39#_c_694_n N_VPWR_c_875_n 0.0164785f $X=8.4 $Y=2.005 $X2=0 $Y2=0
cc_540 N_A_808_39#_c_729_n N_VPWR_c_876_n 0.0170777f $X=9.26 $Y=2.005 $X2=0
+ $Y2=0
cc_541 N_A_808_39#_c_660_n N_VPWR_c_878_n 0.0235138f $X=9.77 $Y=2.005 $X2=0
+ $Y2=0
cc_542 N_A_808_39#_M1033_g N_VPWR_c_881_n 0.00487821f $X=5.7 $Y=2.465 $X2=0
+ $Y2=0
cc_543 N_A_808_39#_M1038_g N_VPWR_c_881_n 0.0054895f $X=6.13 $Y=2.465 $X2=0
+ $Y2=0
cc_544 N_A_808_39#_c_780_p N_VPWR_c_883_n 0.0136943f $X=6.775 $Y=1.96 $X2=0
+ $Y2=0
cc_545 N_A_808_39#_M1005_g N_VPWR_c_886_n 0.00564095f $X=4.115 $Y=2.465 $X2=0
+ $Y2=0
cc_546 N_A_808_39#_M1020_g N_VPWR_c_886_n 0.00357668f $X=4.545 $Y=2.465 $X2=0
+ $Y2=0
cc_547 N_A_808_39#_c_783_p N_VPWR_c_887_n 0.0124525f $X=8.495 $Y=2.45 $X2=0
+ $Y2=0
cc_548 N_A_808_39#_c_784_p N_VPWR_c_888_n 0.0124525f $X=9.355 $Y=2.45 $X2=0
+ $Y2=0
cc_549 N_A_808_39#_M1020_g N_VPWR_c_890_n 0.00911637f $X=4.545 $Y=2.465 $X2=0
+ $Y2=0
cc_550 N_A_808_39#_M1033_g N_VPWR_c_890_n 0.0136165f $X=5.7 $Y=2.465 $X2=0 $Y2=0
cc_551 N_A_808_39#_M1038_g N_VPWR_c_890_n 4.98916e-19 $X=6.13 $Y=2.465 $X2=0
+ $Y2=0
cc_552 N_A_808_39#_M1008_s N_VPWR_c_868_n 0.0041489f $X=6.635 $Y=1.835 $X2=0
+ $Y2=0
cc_553 N_A_808_39#_M1026_s N_VPWR_c_868_n 0.00536646f $X=7.495 $Y=1.835 $X2=0
+ $Y2=0
cc_554 N_A_808_39#_M1007_d N_VPWR_c_868_n 0.00536646f $X=8.355 $Y=1.835 $X2=0
+ $Y2=0
cc_555 N_A_808_39#_M1021_d N_VPWR_c_868_n 0.00536646f $X=9.215 $Y=1.835 $X2=0
+ $Y2=0
cc_556 N_A_808_39#_M1005_g N_VPWR_c_868_n 0.00948291f $X=4.115 $Y=2.465 $X2=0
+ $Y2=0
cc_557 N_A_808_39#_M1020_g N_VPWR_c_868_n 0.00675076f $X=4.545 $Y=2.465 $X2=0
+ $Y2=0
cc_558 N_A_808_39#_M1033_g N_VPWR_c_868_n 0.00824731f $X=5.7 $Y=2.465 $X2=0
+ $Y2=0
cc_559 N_A_808_39#_M1038_g N_VPWR_c_868_n 0.00979102f $X=6.13 $Y=2.465 $X2=0
+ $Y2=0
cc_560 N_A_808_39#_c_780_p N_VPWR_c_868_n 0.00866972f $X=6.775 $Y=1.96 $X2=0
+ $Y2=0
cc_561 N_A_808_39#_c_774_p N_VPWR_c_868_n 0.00730901f $X=7.635 $Y=2.45 $X2=0
+ $Y2=0
cc_562 N_A_808_39#_c_783_p N_VPWR_c_868_n 0.00730901f $X=8.495 $Y=2.45 $X2=0
+ $Y2=0
cc_563 N_A_808_39#_c_784_p N_VPWR_c_868_n 0.00730901f $X=9.355 $Y=2.45 $X2=0
+ $Y2=0
cc_564 N_A_808_39#_M1001_g N_Y_c_1064_n 0.0122297f $X=4.115 $Y=0.745 $X2=0 $Y2=0
cc_565 N_A_808_39#_c_647_n N_Y_c_1064_n 0.0125536f $X=5.625 $Y=1.335 $X2=0 $Y2=0
cc_566 N_A_808_39#_M1005_g N_Y_c_1098_n 0.0127827f $X=4.115 $Y=2.465 $X2=0 $Y2=0
cc_567 N_A_808_39#_M1009_g N_Y_c_1066_n 0.0124691f $X=4.545 $Y=0.745 $X2=0 $Y2=0
cc_568 N_A_808_39#_M1010_g N_Y_c_1066_n 0.0127446f $X=4.985 $Y=0.745 $X2=0 $Y2=0
cc_569 N_A_808_39#_c_640_n N_Y_c_1066_n 0.00435084f $X=5.41 $Y=1.5 $X2=0 $Y2=0
cc_570 N_A_808_39#_c_641_n N_Y_c_1066_n 0.00271119f $X=5.06 $Y=1.5 $X2=0 $Y2=0
cc_571 N_A_808_39#_M1029_g N_Y_c_1066_n 0.0037746f $X=5.485 $Y=0.745 $X2=0 $Y2=0
cc_572 N_A_808_39#_c_647_n N_Y_c_1066_n 0.0684624f $X=5.625 $Y=1.335 $X2=0 $Y2=0
cc_573 N_A_808_39#_c_648_n N_Y_c_1066_n 0.0128849f $X=6.135 $Y=1.335 $X2=0 $Y2=0
cc_574 N_A_808_39#_M1033_g N_Y_c_1109_n 0.0142726f $X=5.7 $Y=2.465 $X2=0 $Y2=0
cc_575 N_A_808_39#_M1029_g N_Y_c_1138_n 0.0106276f $X=5.485 $Y=0.745 $X2=0 $Y2=0
cc_576 N_A_808_39#_M1038_g N_Y_c_1110_n 0.00222705f $X=6.13 $Y=2.465 $X2=0 $Y2=0
cc_577 N_A_808_39#_M1038_g N_Y_c_1140_n 0.00827074f $X=6.13 $Y=2.465 $X2=0 $Y2=0
cc_578 N_A_808_39#_c_641_n N_Y_c_1067_n 0.00255808f $X=5.06 $Y=1.5 $X2=0 $Y2=0
cc_579 N_A_808_39#_c_647_n N_Y_c_1067_n 0.0149737f $X=5.625 $Y=1.335 $X2=0 $Y2=0
cc_580 N_A_808_39#_M1020_g Y 0.0189913f $X=4.545 $Y=2.465 $X2=0 $Y2=0
cc_581 N_A_808_39#_M1005_g N_Y_c_1111_n 0.0056065f $X=4.115 $Y=2.465 $X2=0 $Y2=0
cc_582 N_A_808_39#_M1020_g N_Y_c_1111_n 0.0119108f $X=4.545 $Y=2.465 $X2=0 $Y2=0
cc_583 N_A_808_39#_c_648_n N_A_31_65#_M1029_s 0.00484404f $X=6.135 $Y=1.335
+ $X2=0 $Y2=0
cc_584 N_A_808_39#_M1001_g N_A_31_65#_c_1224_n 0.00207279f $X=4.115 $Y=0.745
+ $X2=0 $Y2=0
cc_585 N_A_808_39#_M1001_g N_A_31_65#_c_1225_n 0.00427993f $X=4.115 $Y=0.745
+ $X2=0 $Y2=0
cc_586 N_A_808_39#_M1009_g N_A_31_65#_c_1225_n 4.73428e-19 $X=4.545 $Y=0.745
+ $X2=0 $Y2=0
cc_587 N_A_808_39#_M1001_g N_A_31_65#_c_1211_n 0.00849712f $X=4.115 $Y=0.745
+ $X2=0 $Y2=0
cc_588 N_A_808_39#_M1009_g N_A_31_65#_c_1211_n 0.00901092f $X=4.545 $Y=0.745
+ $X2=0 $Y2=0
cc_589 N_A_808_39#_M1001_g N_A_31_65#_c_1212_n 0.00137527f $X=4.115 $Y=0.745
+ $X2=0 $Y2=0
cc_590 N_A_808_39#_M1001_g N_A_31_65#_c_1244_n 5.10831e-19 $X=4.115 $Y=0.745
+ $X2=0 $Y2=0
cc_591 N_A_808_39#_M1009_g N_A_31_65#_c_1244_n 0.0058748f $X=4.545 $Y=0.745
+ $X2=0 $Y2=0
cc_592 N_A_808_39#_M1010_g N_A_31_65#_c_1244_n 0.0066764f $X=4.985 $Y=0.745
+ $X2=0 $Y2=0
cc_593 N_A_808_39#_M1029_g N_A_31_65#_c_1244_n 2.43858e-19 $X=5.485 $Y=0.745
+ $X2=0 $Y2=0
cc_594 N_A_808_39#_M1010_g N_A_31_65#_c_1213_n 0.00867251f $X=4.985 $Y=0.745
+ $X2=0 $Y2=0
cc_595 N_A_808_39#_M1029_g N_A_31_65#_c_1213_n 0.015181f $X=5.485 $Y=0.745 $X2=0
+ $Y2=0
cc_596 N_A_808_39#_c_647_n N_A_31_65#_c_1214_n 4.13799e-19 $X=5.625 $Y=1.335
+ $X2=0 $Y2=0
cc_597 N_A_808_39#_c_648_n N_A_31_65#_c_1214_n 0.0271488f $X=6.135 $Y=1.335
+ $X2=0 $Y2=0
cc_598 N_A_808_39#_c_651_n N_A_31_65#_c_1214_n 0.00177372f $X=6.13 $Y=1.5 $X2=0
+ $Y2=0
cc_599 N_A_808_39#_M1009_g N_A_31_65#_c_1215_n 0.00118084f $X=4.545 $Y=0.745
+ $X2=0 $Y2=0
cc_600 N_A_808_39#_M1010_g N_A_31_65#_c_1215_n 0.00159077f $X=4.985 $Y=0.745
+ $X2=0 $Y2=0
cc_601 N_A_808_39#_c_643_n N_VGND_M1018_d 0.0026214f $X=8.365 $Y=1.17 $X2=0
+ $Y2=0
cc_602 N_A_808_39#_c_643_n N_VGND_M1032_d 0.00176891f $X=8.365 $Y=1.17 $X2=0
+ $Y2=0
cc_603 N_A_808_39#_M1001_g N_VGND_c_1336_n 0.00302473f $X=4.115 $Y=0.745 $X2=0
+ $Y2=0
cc_604 N_A_808_39#_M1009_g N_VGND_c_1336_n 0.00302484f $X=4.545 $Y=0.745 $X2=0
+ $Y2=0
cc_605 N_A_808_39#_M1010_g N_VGND_c_1336_n 0.00302473f $X=4.985 $Y=0.745 $X2=0
+ $Y2=0
cc_606 N_A_808_39#_M1029_g N_VGND_c_1336_n 0.00302501f $X=5.485 $Y=0.745 $X2=0
+ $Y2=0
cc_607 N_A_808_39#_M1001_g N_VGND_c_1343_n 0.00435644f $X=4.115 $Y=0.745 $X2=0
+ $Y2=0
cc_608 N_A_808_39#_M1009_g N_VGND_c_1343_n 0.00435666f $X=4.545 $Y=0.745 $X2=0
+ $Y2=0
cc_609 N_A_808_39#_M1010_g N_VGND_c_1343_n 0.00442246f $X=4.985 $Y=0.745 $X2=0
+ $Y2=0
cc_610 N_A_808_39#_M1029_g N_VGND_c_1343_n 0.00491241f $X=5.485 $Y=0.745 $X2=0
+ $Y2=0
cc_611 N_A_808_39#_c_643_n N_A_1235_65#_M1018_s 0.00253571f $X=8.365 $Y=1.17
+ $X2=-0.19 $Y2=-0.245
cc_612 N_A_808_39#_c_643_n N_A_1235_65#_M1030_s 0.00176461f $X=8.365 $Y=1.17
+ $X2=0 $Y2=0
cc_613 N_A_808_39#_c_643_n N_A_1235_65#_M1034_s 0.00176461f $X=8.365 $Y=1.17
+ $X2=0 $Y2=0
cc_614 N_A_808_39#_c_644_n N_A_1235_65#_M1015_s 0.00177068f $X=9.225 $Y=1.16
+ $X2=0 $Y2=0
cc_615 N_A_808_39#_c_645_n N_A_1235_65#_M1028_s 0.00274841f $X=9.77 $Y=1.16
+ $X2=0 $Y2=0
cc_616 N_A_808_39#_M1029_g N_A_1235_65#_c_1483_n 8.79814e-19 $X=5.485 $Y=0.745
+ $X2=0 $Y2=0
cc_617 N_A_808_39#_c_643_n N_A_1235_65#_c_1493_n 0.0364396f $X=8.365 $Y=1.17
+ $X2=0 $Y2=0
cc_618 N_A_808_39#_c_643_n N_A_1235_65#_c_1484_n 0.0219308f $X=8.365 $Y=1.17
+ $X2=0 $Y2=0
cc_619 N_A_808_39#_c_643_n N_A_1235_65#_c_1498_n 0.0323235f $X=8.365 $Y=1.17
+ $X2=0 $Y2=0
cc_620 N_A_808_39#_c_643_n N_A_1235_65#_c_1514_n 0.0134726f $X=8.365 $Y=1.17
+ $X2=0 $Y2=0
cc_621 N_A_808_39#_M1004_d N_A_1235_65#_c_1486_n 0.00181066f $X=8.39 $Y=0.325
+ $X2=0 $Y2=0
cc_622 N_A_808_39#_c_643_n N_A_1235_65#_c_1486_n 0.00277205f $X=8.365 $Y=1.17
+ $X2=0 $Y2=0
cc_623 N_A_808_39#_c_696_n N_A_1235_65#_c_1486_n 0.0152308f $X=8.53 $Y=0.7 $X2=0
+ $Y2=0
cc_624 N_A_808_39#_c_644_n N_A_1235_65#_c_1486_n 0.00287913f $X=9.225 $Y=1.16
+ $X2=0 $Y2=0
cc_625 N_A_808_39#_c_644_n N_A_1235_65#_c_1519_n 0.0135407f $X=9.225 $Y=1.16
+ $X2=0 $Y2=0
cc_626 N_A_808_39#_M1025_d N_A_1235_65#_c_1488_n 0.00184993f $X=9.25 $Y=0.325
+ $X2=0 $Y2=0
cc_627 N_A_808_39#_c_644_n N_A_1235_65#_c_1488_n 0.0028245f $X=9.225 $Y=1.16
+ $X2=0 $Y2=0
cc_628 N_A_808_39#_c_737_n N_A_1235_65#_c_1488_n 0.014436f $X=9.39 $Y=0.7 $X2=0
+ $Y2=0
cc_629 N_A_808_39#_c_645_n N_A_1235_65#_c_1488_n 0.0028245f $X=9.77 $Y=1.16
+ $X2=0 $Y2=0
cc_630 N_A_808_39#_c_645_n N_A_1235_65#_c_1489_n 0.0220001f $X=9.77 $Y=1.16
+ $X2=0 $Y2=0
cc_631 N_A_808_39#_c_643_n N_A_1235_65#_c_1525_n 0.0134216f $X=8.365 $Y=1.17
+ $X2=0 $Y2=0
cc_632 N_VPWR_c_868_n N_A_110_367#_M1019_s 0.00394625f $X=9.84 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_633 N_VPWR_c_868_n N_A_110_367#_M1036_s 0.00238445f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_634 N_VPWR_c_868_n N_A_110_367#_M1012_d 0.00238445f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_635 N_VPWR_c_868_n N_A_110_367#_M1022_d 0.00324228f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_636 N_VPWR_c_879_n N_A_110_367#_c_1030_n 0.0663374f $X=3.715 $Y=3.33 $X2=0
+ $Y2=0
cc_637 N_VPWR_c_868_n N_A_110_367#_c_1030_n 0.068452f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_638 N_VPWR_c_885_n N_A_110_367#_c_1032_n 0.00871781f $X=1.035 $Y=3.33 $X2=0
+ $Y2=0
cc_639 N_VPWR_c_868_n N_A_110_367#_c_1032_n 0.00936171f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_640 N_VPWR_M1031_d N_A_110_367#_c_1034_n 0.00746518f $X=0.98 $Y=1.835 $X2=0
+ $Y2=0
cc_641 N_VPWR_c_879_n N_A_110_367#_c_1034_n 0.00203583f $X=3.715 $Y=3.33 $X2=0
+ $Y2=0
cc_642 N_VPWR_c_885_n N_A_110_367#_c_1034_n 0.00203583f $X=1.035 $Y=3.33 $X2=0
+ $Y2=0
cc_643 N_VPWR_c_889_n N_A_110_367#_c_1034_n 0.0240398f $X=1.2 $Y=3.065 $X2=0
+ $Y2=0
cc_644 N_VPWR_c_868_n N_A_110_367#_c_1034_n 0.00849449f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_645 N_VPWR_c_868_n N_Y_M1002_s 0.00238445f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_646 N_VPWR_c_868_n N_Y_M1013_s 0.00238445f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_647 N_VPWR_c_868_n N_Y_M1005_s 0.00310528f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_648 N_VPWR_c_868_n N_Y_M1033_s 0.00380103f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_649 N_VPWR_M1019_d N_Y_c_1063_n 0.00135026f $X=0.135 $Y=1.835 $X2=0 $Y2=0
cc_650 N_VPWR_M1019_d N_Y_c_1087_n 0.00206092f $X=0.135 $Y=1.835 $X2=0 $Y2=0
cc_651 N_VPWR_M1031_d N_Y_c_1087_n 0.00231953f $X=0.98 $Y=1.835 $X2=0 $Y2=0
cc_652 N_VPWR_c_870_n N_Y_c_1087_n 0.00728199f $X=0.26 $Y=2.365 $X2=0 $Y2=0
cc_653 N_VPWR_M1019_d N_Y_c_1069_n 0.00233802f $X=0.135 $Y=1.835 $X2=0 $Y2=0
cc_654 N_VPWR_c_870_n N_Y_c_1069_n 0.0162318f $X=0.26 $Y=2.365 $X2=0 $Y2=0
cc_655 N_VPWR_M1031_d N_Y_c_1094_n 0.00226212f $X=0.98 $Y=1.835 $X2=0 $Y2=0
cc_656 N_VPWR_c_870_n N_Y_c_1094_n 2.72595e-19 $X=0.26 $Y=2.365 $X2=0 $Y2=0
cc_657 N_VPWR_M1031_d N_Y_c_1098_n 0.00692369f $X=0.98 $Y=1.835 $X2=0 $Y2=0
cc_658 N_VPWR_M1037_d N_Y_c_1098_n 0.00502871f $X=3.72 $Y=1.835 $X2=0 $Y2=0
cc_659 N_VPWR_c_871_n N_Y_c_1098_n 0.0173521f $X=3.88 $Y=2.745 $X2=0 $Y2=0
cc_660 N_VPWR_M1031_d N_Y_c_1107_n 8.58736e-19 $X=0.98 $Y=1.835 $X2=0 $Y2=0
cc_661 N_VPWR_c_870_n N_Y_c_1107_n 0.00574049f $X=0.26 $Y=2.365 $X2=0 $Y2=0
cc_662 N_VPWR_M1020_d N_Y_c_1109_n 0.0272988f $X=4.62 $Y=1.835 $X2=0 $Y2=0
cc_663 N_VPWR_c_890_n N_Y_c_1109_n 0.0629677f $X=5.485 $Y=2.53 $X2=0 $Y2=0
cc_664 N_VPWR_c_881_n N_Y_c_1140_n 0.015688f $X=6.25 $Y=3.33 $X2=0 $Y2=0
cc_665 N_VPWR_c_868_n N_Y_c_1140_n 0.00984745f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_666 N_VPWR_c_886_n Y 0.0258389f $X=4.815 $Y=3.33 $X2=0 $Y2=0
cc_667 N_VPWR_c_868_n Y 0.0158801f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_668 N_A_110_367#_c_1037_n N_Y_M1002_s 0.0038093f $X=3.43 $Y=2.795 $X2=0.475
+ $Y2=2.465
cc_669 N_A_110_367#_c_1037_n N_Y_M1013_s 0.0038093f $X=3.43 $Y=2.795 $X2=0 $Y2=0
cc_670 N_A_110_367#_M1019_s N_Y_c_1087_n 0.00465691f $X=0.55 $Y=1.835 $X2=1.495
+ $Y2=2.465
cc_671 N_A_110_367#_c_1032_n N_Y_c_1087_n 0.0086898f $X=0.865 $Y=2.785 $X2=1.495
+ $Y2=2.465
cc_672 N_A_110_367#_M1036_s N_Y_c_1098_n 0.00354408f $X=1.57 $Y=1.835 $X2=3.645
+ $Y2=2.465
cc_673 N_A_110_367#_M1012_d N_Y_c_1098_n 0.00341991f $X=2.43 $Y=1.835 $X2=3.645
+ $Y2=2.465
cc_674 N_A_110_367#_M1022_d N_Y_c_1098_n 0.00348918f $X=3.29 $Y=1.835 $X2=3.645
+ $Y2=2.465
cc_675 N_A_110_367#_c_1034_n N_Y_c_1098_n 0.135365f $X=1.535 $Y=2.79 $X2=3.645
+ $Y2=2.465
cc_676 N_A_110_367#_c_1034_n N_Y_c_1107_n 0.0088302f $X=1.535 $Y=2.79 $X2=0
+ $Y2=0
cc_677 N_Y_c_1064_n N_A_31_65#_M1006_d 0.00113743f $X=4.235 $Y=1.16 $X2=-0.19
+ $Y2=-0.245
cc_678 N_Y_c_1065_n N_A_31_65#_M1006_d 0.00185101f $X=0.275 $Y=1.16 $X2=-0.19
+ $Y2=-0.245
cc_679 N_Y_c_1064_n N_A_31_65#_M1017_d 0.00176461f $X=4.235 $Y=1.16 $X2=0 $Y2=0
cc_680 N_Y_c_1064_n N_A_31_65#_M1000_d 0.00176461f $X=4.235 $Y=1.16 $X2=0 $Y2=0
cc_681 N_Y_c_1064_n N_A_31_65#_M1011_d 0.00176461f $X=4.235 $Y=1.16 $X2=0 $Y2=0
cc_682 N_Y_c_1064_n N_A_31_65#_M1027_d 0.00176461f $X=4.235 $Y=1.16 $X2=0 $Y2=0
cc_683 N_Y_c_1066_n N_A_31_65#_M1009_s 0.00187091f $X=5.105 $Y=1.16 $X2=0 $Y2=0
cc_684 N_Y_c_1064_n N_A_31_65#_c_1218_n 0.0364396f $X=4.235 $Y=1.16 $X2=0 $Y2=0
cc_685 N_Y_c_1064_n N_A_31_65#_c_1207_n 0.0105191f $X=4.235 $Y=1.16 $X2=0 $Y2=0
cc_686 N_Y_c_1065_n N_A_31_65#_c_1207_n 0.0125925f $X=0.275 $Y=1.16 $X2=0 $Y2=0
cc_687 N_Y_c_1064_n N_A_31_65#_c_1223_n 0.0323235f $X=4.235 $Y=1.16 $X2=0 $Y2=0
cc_688 N_Y_c_1064_n N_A_31_65#_c_1231_n 0.0323235f $X=4.235 $Y=1.16 $X2=0 $Y2=0
cc_689 N_Y_c_1064_n N_A_31_65#_c_1224_n 0.0536061f $X=4.235 $Y=1.16 $X2=0 $Y2=0
cc_690 N_Y_M1001_d N_A_31_65#_c_1211_n 0.00176773f $X=4.19 $Y=0.325 $X2=0 $Y2=0
cc_691 N_Y_c_1064_n N_A_31_65#_c_1211_n 0.00281275f $X=4.235 $Y=1.16 $X2=0 $Y2=0
cc_692 N_Y_c_1193_p N_A_31_65#_c_1211_n 0.012655f $X=4.33 $Y=0.77 $X2=0 $Y2=0
cc_693 N_Y_c_1066_n N_A_31_65#_c_1211_n 0.00303868f $X=5.105 $Y=1.16 $X2=0 $Y2=0
cc_694 N_Y_c_1066_n N_A_31_65#_c_1244_n 0.0170664f $X=5.105 $Y=1.16 $X2=0 $Y2=0
cc_695 N_Y_M1010_d N_A_31_65#_c_1213_n 0.00250873f $X=5.06 $Y=0.325 $X2=0 $Y2=0
cc_696 N_Y_c_1066_n N_A_31_65#_c_1213_n 0.00275981f $X=5.105 $Y=1.16 $X2=0 $Y2=0
cc_697 N_Y_c_1138_n N_A_31_65#_c_1213_n 0.0195673f $X=5.27 $Y=0.68 $X2=0 $Y2=0
cc_698 N_Y_c_1064_n N_A_31_65#_c_1276_n 0.0134041f $X=4.235 $Y=1.16 $X2=0 $Y2=0
cc_699 N_Y_c_1064_n N_A_31_65#_c_1277_n 0.0134041f $X=4.235 $Y=1.16 $X2=0 $Y2=0
cc_700 N_Y_c_1064_n N_A_31_65#_c_1278_n 0.0134041f $X=4.235 $Y=1.16 $X2=0 $Y2=0
cc_701 N_Y_c_1064_n N_VGND_M1006_s 0.0026214f $X=4.235 $Y=1.16 $X2=-0.19
+ $Y2=-0.245
cc_702 N_Y_c_1064_n N_VGND_M1024_s 0.00176891f $X=4.235 $Y=1.16 $X2=0 $Y2=0
cc_703 N_Y_c_1064_n N_VGND_M1003_s 0.00176891f $X=4.235 $Y=1.16 $X2=0 $Y2=0
cc_704 N_Y_c_1064_n N_VGND_M1023_s 0.0026214f $X=4.235 $Y=1.16 $X2=0 $Y2=0
cc_705 N_A_31_65#_c_1218_n N_VGND_M1006_s 0.00492724f $X=1.155 $Y=0.82 $X2=-0.19
+ $Y2=-0.245
cc_706 N_A_31_65#_c_1223_n N_VGND_M1024_s 0.00349176f $X=2.005 $Y=0.82 $X2=0
+ $Y2=0
cc_707 N_A_31_65#_c_1231_n N_VGND_M1003_s 0.00335437f $X=2.865 $Y=0.82 $X2=0
+ $Y2=0
cc_708 N_A_31_65#_c_1224_n N_VGND_M1023_s 0.00509244f $X=3.735 $Y=0.82 $X2=0
+ $Y2=0
cc_709 N_A_31_65#_c_1206_n N_VGND_c_1326_n 0.0113376f $X=0.3 $Y=0.46 $X2=0 $Y2=0
cc_710 N_A_31_65#_c_1218_n N_VGND_c_1326_n 0.0202782f $X=1.155 $Y=0.82 $X2=0
+ $Y2=0
cc_711 N_A_31_65#_c_1208_n N_VGND_c_1326_n 0.0109791f $X=1.24 $Y=0.48 $X2=0
+ $Y2=0
cc_712 N_A_31_65#_c_1208_n N_VGND_c_1327_n 0.0119864f $X=1.24 $Y=0.48 $X2=0
+ $Y2=0
cc_713 N_A_31_65#_c_1223_n N_VGND_c_1327_n 0.016459f $X=2.005 $Y=0.82 $X2=0
+ $Y2=0
cc_714 N_A_31_65#_c_1209_n N_VGND_c_1327_n 0.0119986f $X=2.1 $Y=0.48 $X2=0 $Y2=0
cc_715 N_A_31_65#_c_1209_n N_VGND_c_1328_n 0.0119986f $X=2.1 $Y=0.48 $X2=0 $Y2=0
cc_716 N_A_31_65#_c_1231_n N_VGND_c_1328_n 0.016459f $X=2.865 $Y=0.82 $X2=0
+ $Y2=0
cc_717 N_A_31_65#_c_1210_n N_VGND_c_1328_n 0.0119986f $X=2.96 $Y=0.45 $X2=0
+ $Y2=0
cc_718 N_A_31_65#_c_1210_n N_VGND_c_1329_n 0.0119986f $X=2.96 $Y=0.45 $X2=0
+ $Y2=0
cc_719 N_A_31_65#_c_1224_n N_VGND_c_1329_n 0.0210125f $X=3.735 $Y=0.82 $X2=0
+ $Y2=0
cc_720 N_A_31_65#_c_1212_n N_VGND_c_1329_n 0.0100087f $X=4.065 $Y=0.345 $X2=0
+ $Y2=0
cc_721 N_A_31_65#_c_1223_n N_VGND_c_1332_n 0.00196209f $X=2.005 $Y=0.82 $X2=0
+ $Y2=0
cc_722 N_A_31_65#_c_1209_n N_VGND_c_1332_n 0.0112458f $X=2.1 $Y=0.48 $X2=0 $Y2=0
cc_723 N_A_31_65#_c_1231_n N_VGND_c_1332_n 0.00196209f $X=2.865 $Y=0.82 $X2=0
+ $Y2=0
cc_724 N_A_31_65#_c_1231_n N_VGND_c_1334_n 0.00196209f $X=2.865 $Y=0.82 $X2=0
+ $Y2=0
cc_725 N_A_31_65#_c_1210_n N_VGND_c_1334_n 0.0112458f $X=2.96 $Y=0.45 $X2=0
+ $Y2=0
cc_726 N_A_31_65#_c_1224_n N_VGND_c_1334_n 0.00196209f $X=3.735 $Y=0.82 $X2=0
+ $Y2=0
cc_727 N_A_31_65#_c_1224_n N_VGND_c_1336_n 0.00203769f $X=3.735 $Y=0.82 $X2=0
+ $Y2=0
cc_728 N_A_31_65#_c_1211_n N_VGND_c_1336_n 0.0341076f $X=4.605 $Y=0.345 $X2=0
+ $Y2=0
cc_729 N_A_31_65#_c_1212_n N_VGND_c_1336_n 0.0234012f $X=4.065 $Y=0.345 $X2=0
+ $Y2=0
cc_730 N_A_31_65#_c_1213_n N_VGND_c_1336_n 0.0659078f $X=5.605 $Y=0.34 $X2=0
+ $Y2=0
cc_731 N_A_31_65#_c_1215_n N_VGND_c_1336_n 0.0234366f $X=4.77 $Y=0.345 $X2=0
+ $Y2=0
cc_732 N_A_31_65#_c_1206_n N_VGND_c_1340_n 0.0185237f $X=0.3 $Y=0.46 $X2=0 $Y2=0
cc_733 N_A_31_65#_c_1218_n N_VGND_c_1340_n 0.00196209f $X=1.155 $Y=0.82 $X2=0
+ $Y2=0
cc_734 N_A_31_65#_c_1218_n N_VGND_c_1341_n 0.00216849f $X=1.155 $Y=0.82 $X2=0
+ $Y2=0
cc_735 N_A_31_65#_c_1208_n N_VGND_c_1341_n 0.0106476f $X=1.24 $Y=0.48 $X2=0
+ $Y2=0
cc_736 N_A_31_65#_c_1223_n N_VGND_c_1341_n 0.00196209f $X=2.005 $Y=0.82 $X2=0
+ $Y2=0
cc_737 N_A_31_65#_c_1206_n N_VGND_c_1343_n 0.0123459f $X=0.3 $Y=0.46 $X2=0 $Y2=0
cc_738 N_A_31_65#_c_1218_n N_VGND_c_1343_n 0.00950092f $X=1.155 $Y=0.82 $X2=0
+ $Y2=0
cc_739 N_A_31_65#_c_1208_n N_VGND_c_1343_n 0.00680041f $X=1.24 $Y=0.48 $X2=0
+ $Y2=0
cc_740 N_A_31_65#_c_1223_n N_VGND_c_1343_n 0.00899218f $X=2.005 $Y=0.82 $X2=0
+ $Y2=0
cc_741 N_A_31_65#_c_1209_n N_VGND_c_1343_n 0.00718246f $X=2.1 $Y=0.48 $X2=0
+ $Y2=0
cc_742 N_A_31_65#_c_1231_n N_VGND_c_1343_n 0.00899218f $X=2.865 $Y=0.82 $X2=0
+ $Y2=0
cc_743 N_A_31_65#_c_1210_n N_VGND_c_1343_n 0.00718246f $X=2.96 $Y=0.45 $X2=0
+ $Y2=0
cc_744 N_A_31_65#_c_1224_n N_VGND_c_1343_n 0.00928306f $X=3.735 $Y=0.82 $X2=0
+ $Y2=0
cc_745 N_A_31_65#_c_1211_n N_VGND_c_1343_n 0.0191369f $X=4.605 $Y=0.345 $X2=0
+ $Y2=0
cc_746 N_A_31_65#_c_1212_n N_VGND_c_1343_n 0.0125856f $X=4.065 $Y=0.345 $X2=0
+ $Y2=0
cc_747 N_A_31_65#_c_1213_n N_VGND_c_1343_n 0.0367512f $X=5.605 $Y=0.34 $X2=0
+ $Y2=0
cc_748 N_A_31_65#_c_1215_n N_VGND_c_1343_n 0.0126315f $X=4.77 $Y=0.345 $X2=0
+ $Y2=0
cc_749 N_A_31_65#_c_1213_n N_A_1235_65#_c_1483_n 0.00946438f $X=5.605 $Y=0.34
+ $X2=0 $Y2=0
cc_750 N_A_31_65#_c_1214_n N_A_1235_65#_c_1483_n 0.0236988f $X=5.77 $Y=0.47
+ $X2=0 $Y2=0
cc_751 N_A_31_65#_c_1214_n N_A_1235_65#_c_1484_n 0.0134079f $X=5.77 $Y=0.47
+ $X2=0 $Y2=0
cc_752 N_VGND_c_1330_n N_A_1235_65#_c_1483_n 0.0109215f $X=6.8 $Y=0.45 $X2=0
+ $Y2=0
cc_753 N_VGND_c_1336_n N_A_1235_65#_c_1483_n 0.0176244f $X=6.635 $Y=0 $X2=0
+ $Y2=0
cc_754 N_VGND_c_1343_n N_A_1235_65#_c_1483_n 0.0122772f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_755 N_VGND_M1018_d N_A_1235_65#_c_1493_n 0.00492443f $X=6.59 $Y=0.325 $X2=0
+ $Y2=0
cc_756 N_VGND_c_1330_n N_A_1235_65#_c_1493_n 0.0203287f $X=6.8 $Y=0.45 $X2=0
+ $Y2=0
cc_757 N_VGND_c_1336_n N_A_1235_65#_c_1493_n 0.00191958f $X=6.635 $Y=0 $X2=0
+ $Y2=0
cc_758 N_VGND_c_1338_n N_A_1235_65#_c_1493_n 0.00197392f $X=7.505 $Y=0 $X2=0
+ $Y2=0
cc_759 N_VGND_c_1343_n N_A_1235_65#_c_1493_n 0.00888322f $X=9.84 $Y=0 $X2=0
+ $Y2=0
cc_760 N_VGND_c_1330_n N_A_1235_65#_c_1485_n 0.0123855f $X=6.8 $Y=0.45 $X2=0
+ $Y2=0
cc_761 N_VGND_c_1331_n N_A_1235_65#_c_1485_n 0.0123855f $X=7.67 $Y=0.45 $X2=0
+ $Y2=0
cc_762 N_VGND_c_1338_n N_A_1235_65#_c_1485_n 0.0118581f $X=7.505 $Y=0 $X2=0
+ $Y2=0
cc_763 N_VGND_c_1343_n N_A_1235_65#_c_1485_n 0.00756799f $X=9.84 $Y=0 $X2=0
+ $Y2=0
cc_764 N_VGND_M1032_d N_A_1235_65#_c_1498_n 0.00335318f $X=7.53 $Y=0.325 $X2=0
+ $Y2=0
cc_765 N_VGND_c_1331_n N_A_1235_65#_c_1498_n 0.0165001f $X=7.67 $Y=0.45 $X2=0
+ $Y2=0
cc_766 N_VGND_c_1338_n N_A_1235_65#_c_1498_n 0.00191958f $X=7.505 $Y=0 $X2=0
+ $Y2=0
cc_767 N_VGND_c_1342_n N_A_1235_65#_c_1498_n 0.00191958f $X=9.84 $Y=0 $X2=0
+ $Y2=0
cc_768 N_VGND_c_1343_n N_A_1235_65#_c_1498_n 0.00890342f $X=9.84 $Y=0 $X2=0
+ $Y2=0
cc_769 N_VGND_c_1342_n N_A_1235_65#_c_1486_n 0.0423919f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_770 N_VGND_c_1343_n N_A_1235_65#_c_1486_n 0.0238473f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_771 N_VGND_c_1331_n N_A_1235_65#_c_1487_n 0.0100029f $X=7.67 $Y=0.45 $X2=0
+ $Y2=0
cc_772 N_VGND_c_1342_n N_A_1235_65#_c_1487_n 0.0135897f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_773 N_VGND_c_1343_n N_A_1235_65#_c_1487_n 0.00738095f $X=9.84 $Y=0 $X2=0
+ $Y2=0
cc_774 N_VGND_c_1342_n N_A_1235_65#_c_1488_n 0.0607825f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_775 N_VGND_c_1343_n N_A_1235_65#_c_1488_n 0.0339095f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_776 N_VGND_c_1342_n N_A_1235_65#_c_1490_n 0.0135587f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_777 N_VGND_c_1343_n N_A_1235_65#_c_1490_n 0.00737512f $X=9.84 $Y=0 $X2=0
+ $Y2=0
