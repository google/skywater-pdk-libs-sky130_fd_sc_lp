* File: sky130_fd_sc_lp__a211o_4.spice
* Created: Wed Sep  2 09:17:39 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__a211o_4.pex.spice"
.subckt sky130_fd_sc_lp__a211o_4  VNB VPB B1 C1 A2 A1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A1	A1
* A2	A2
* C1	C1
* B1	B1
* VPB	VPB
* VNB	VNB
MM1007 N_X_M1007_d N_A_103_263#_M1007_g N_VGND_M1007_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75005.3 A=0.126 P=1.98 MULT=1
MM1008 N_X_M1007_d N_A_103_263#_M1008_g N_VGND_M1008_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75004.9 A=0.126 P=1.98 MULT=1
MM1013 N_X_M1013_d N_A_103_263#_M1013_g N_VGND_M1008_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1239 AS=0.1176 PD=1.135 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.1
+ SB=75004.4 A=0.126 P=1.98 MULT=1
MM1023 N_X_M1013_d N_A_103_263#_M1023_g N_VGND_M1023_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1239 AS=0.1176 PD=1.135 PS=1.12 NRD=2.136 NRS=0 M=1 R=5.6 SA=75001.5
+ SB=75004 A=0.126 P=1.98 MULT=1
MM1002 N_VGND_M1023_s N_B1_M1002_g N_A_103_263#_M1002_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1239 PD=1.12 PS=1.135 NRD=0 NRS=0 M=1 R=5.6 SA=75001.9
+ SB=75003.6 A=0.126 P=1.98 MULT=1
MM1004 N_VGND_M1004_d N_C1_M1004_g N_A_103_263#_M1002_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1239 PD=1.12 PS=1.135 NRD=0 NRS=2.136 M=1 R=5.6 SA=75002.4
+ SB=75003.1 A=0.126 P=1.98 MULT=1
MM1019 N_VGND_M1004_d N_C1_M1019_g N_A_103_263#_M1019_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002.8
+ SB=75002.7 A=0.126 P=1.98 MULT=1
MM1016 N_VGND_M1016_d N_B1_M1016_g N_A_103_263#_M1019_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2604 AS=0.1176 PD=1.46 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75003.2
+ SB=75002.2 A=0.126 P=1.98 MULT=1
MM1012 N_A_1006_47#_M1012_d N_A2_M1012_g N_VGND_M1016_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2604 PD=1.12 PS=1.46 NRD=0 NRS=0 M=1 R=5.6 SA=75004 SB=75001.5
+ A=0.126 P=1.98 MULT=1
MM1009 N_A_1006_47#_M1012_d N_A1_M1009_g N_A_103_263#_M1009_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75004.4
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1020 N_A_1006_47#_M1020_d N_A1_M1020_g N_A_103_263#_M1009_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75004.9
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1017 N_A_1006_47#_M1020_d N_A2_M1017_g N_VGND_M1017_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75005.3
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1001 N_VPWR_M1001_d N_A_103_263#_M1001_g N_X_M1001_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75001.5 A=0.189 P=2.82 MULT=1
MM1006 N_VPWR_M1006_d N_A_103_263#_M1006_g N_X_M1001_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1014 N_VPWR_M1006_d N_A_103_263#_M1014_g N_X_M1014_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1021 N_VPWR_M1021_d N_A_103_263#_M1021_g N_X_M1014_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.5
+ SB=75000.2 A=0.189 P=2.82 MULT=1
MM1015 N_A_610_367#_M1015_d N_B1_M1015_g N_A_527_367#_M1015_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75003.5 A=0.189 P=2.82 MULT=1
MM1000 N_A_610_367#_M1015_d N_C1_M1000_g N_A_103_263#_M1000_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75003 A=0.189 P=2.82 MULT=1
MM1010 N_A_610_367#_M1010_d N_C1_M1010_g N_A_103_263#_M1000_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.2016 AS=0.1764 PD=1.58 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75002.6 A=0.189 P=2.82 MULT=1
MM1022 N_A_610_367#_M1010_d N_B1_M1022_g N_A_527_367#_M1022_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.2016 AS=0.2457 PD=1.58 PS=1.65 NRD=6.2449 NRS=7.0329 M=1 R=8.4
+ SA=75001.5 SB=75002.1 A=0.189 P=2.82 MULT=1
MM1005 N_VPWR_M1005_d N_A2_M1005_g N_A_527_367#_M1022_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.2457 AS=0.2457 PD=1.65 PS=1.65 NRD=0 NRS=10.1455 M=1 R=8.4
+ SA=75002.1 SB=75001.6 A=0.189 P=2.82 MULT=1
MM1003 N_VPWR_M1005_d N_A1_M1003_g N_A_527_367#_M1003_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.2457 AS=0.1764 PD=1.65 PS=1.54 NRD=17.1981 NRS=0 M=1 R=8.4
+ SA=75002.6 SB=75001.1 A=0.189 P=2.82 MULT=1
MM1011 N_VPWR_M1011_d N_A1_M1011_g N_A_527_367#_M1003_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75003
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1018 N_VPWR_M1011_d N_A2_M1018_g N_A_527_367#_M1018_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75003.5
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX24_noxref VNB VPB NWDIODE A=13.2415 P=17.93
*
.include "sky130_fd_sc_lp__a211o_4.pxi.spice"
*
.ends
*
*
