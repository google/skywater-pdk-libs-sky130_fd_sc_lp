* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__nor3b_lp A B C_N VGND VNB VPB VPWR Y
X0 a_610_57# C_N a_350_269# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 a_286_409# a_350_269# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X2 a_294_57# B Y VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 Y a_350_269# a_452_57# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 a_452_57# a_350_269# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 VPWR C_N a_350_269# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X6 VGND C_N a_610_57# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 Y A a_136_57# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 a_136_57# A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 VPWR A a_188_409# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X10 VGND B a_294_57# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X11 a_188_409# B a_286_409# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
.ends
