* File: sky130_fd_sc_lp__inputiso1p_lp.pxi.spice
* Created: Wed Sep  2 09:55:18 2020
* 
x_PM_SKY130_FD_SC_LP__INPUTISO1P_LP%A N_A_c_43_n N_A_M1007_g N_A_c_44_n
+ N_A_M1005_g N_A_c_46_n N_A_M1008_g A A PM_SKY130_FD_SC_LP__INPUTISO1P_LP%A
x_PM_SKY130_FD_SC_LP__INPUTISO1P_LP%SLEEP N_SLEEP_M1000_g N_SLEEP_M1001_g
+ N_SLEEP_M1009_g SLEEP N_SLEEP_c_83_n N_SLEEP_c_81_n
+ PM_SKY130_FD_SC_LP__INPUTISO1P_LP%SLEEP
x_PM_SKY130_FD_SC_LP__INPUTISO1P_LP%A_161_489# N_A_161_489#_M1008_d
+ N_A_161_489#_M1005_s N_A_161_489#_c_118_n N_A_161_489#_M1002_g
+ N_A_161_489#_M1003_g N_A_161_489#_c_119_n N_A_161_489#_M1004_g
+ N_A_161_489#_M1006_g N_A_161_489#_c_126_n N_A_161_489#_c_127_n
+ N_A_161_489#_c_128_n N_A_161_489#_c_120_n N_A_161_489#_c_121_n
+ N_A_161_489#_c_122_n N_A_161_489#_c_169_p N_A_161_489#_c_151_n
+ N_A_161_489#_c_123_n PM_SKY130_FD_SC_LP__INPUTISO1P_LP%A_161_489#
x_PM_SKY130_FD_SC_LP__INPUTISO1P_LP%VPWR N_VPWR_M1000_d N_VPWR_c_183_n VPWR
+ N_VPWR_c_184_n N_VPWR_c_185_n N_VPWR_c_182_n N_VPWR_c_187_n
+ PM_SKY130_FD_SC_LP__INPUTISO1P_LP%VPWR
x_PM_SKY130_FD_SC_LP__INPUTISO1P_LP%X N_X_M1004_d N_X_M1006_d X X X X X
+ N_X_c_211_n X X X X X PM_SKY130_FD_SC_LP__INPUTISO1P_LP%X
x_PM_SKY130_FD_SC_LP__INPUTISO1P_LP%VGND N_VGND_M1007_s N_VGND_M1009_d
+ N_VGND_c_221_n N_VGND_c_222_n VGND N_VGND_c_223_n N_VGND_c_224_n
+ N_VGND_c_225_n N_VGND_c_226_n N_VGND_c_227_n N_VGND_c_228_n
+ PM_SKY130_FD_SC_LP__INPUTISO1P_LP%VGND
cc_1 VNB N_A_c_43_n 0.0174937f $X=-0.19 $Y=-0.245 $X2=0.81 $Y2=0.96
cc_2 VNB N_A_c_44_n 0.100216f $X=-0.19 $Y=-0.245 $X2=1.15 $Y2=1.645
cc_3 VNB N_A_M1005_g 4.92816e-19 $X=-0.19 $Y=-0.245 $X2=1.15 $Y2=2.655
cc_4 VNB N_A_c_46_n 0.0141934f $X=-0.19 $Y=-0.245 $X2=1.17 $Y2=0.96
cc_5 VNB A 0.0235969f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_6 VNB N_SLEEP_M1000_g 5.47148e-19 $X=-0.19 $Y=-0.245 $X2=0.81 $Y2=0.675
cc_7 VNB N_SLEEP_M1001_g 0.0301649f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_SLEEP_M1009_g 0.0292713f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_9 VNB N_SLEEP_c_81_n 0.054154f $X=-0.19 $Y=-0.245 $X2=0.89 $Y2=1.665
cc_10 VNB N_A_161_489#_c_118_n 0.0156843f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_161_489#_c_119_n 0.020326f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_161_489#_c_120_n 0.00525468f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_161_489#_c_121_n 0.0206002f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_161_489#_c_122_n 0.00879765f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_161_489#_c_123_n 0.0632971f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_VPWR_c_182_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_X_c_211_n 0.0692912f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.295
cc_18 VNB N_VGND_c_221_n 0.0316526f $X=-0.19 $Y=-0.245 $X2=1.17 $Y2=0.675
cc_19 VNB N_VGND_c_222_n 0.0116388f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_VGND_c_223_n 0.0167814f $X=-0.19 $Y=-0.245 $X2=1.06 $Y2=1.48
cc_21 VNB N_VGND_c_224_n 0.0383522f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_VGND_c_225_n 0.0319968f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_VGND_c_226_n 0.252491f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_VGND_c_227_n 0.00577043f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_228_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VPB N_A_M1005_g 0.0646632f $X=-0.19 $Y=1.655 $X2=1.15 $Y2=2.655
cc_27 VPB A 0.0161359f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_28 VPB N_SLEEP_M1000_g 0.0659857f $X=-0.19 $Y=1.655 $X2=0.81 $Y2=0.675
cc_29 VPB N_SLEEP_c_83_n 0.00582997f $X=-0.19 $Y=1.655 $X2=0.89 $Y2=1.48
cc_30 VPB N_A_161_489#_M1003_g 0.0216969f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_31 VPB N_A_161_489#_M1006_g 0.0203893f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_32 VPB N_A_161_489#_c_126_n 0.0281772f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_33 VPB N_A_161_489#_c_127_n 0.0236459f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_34 VPB N_A_161_489#_c_128_n 0.00984468f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_35 VPB N_A_161_489#_c_123_n 0.00293676f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_36 VPB N_VPWR_c_183_n 0.0161717f $X=-0.19 $Y=1.655 $X2=1.15 $Y2=2.655
cc_37 VPB N_VPWR_c_184_n 0.0499151f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_38 VPB N_VPWR_c_185_n 0.028827f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_39 VPB N_VPWR_c_182_n 0.0894076f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_40 VPB N_VPWR_c_187_n 0.014097f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_41 VPB N_X_c_211_n 0.0680606f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=1.295
cc_42 N_A_M1005_g N_SLEEP_M1000_g 0.0519587f $X=1.15 $Y=2.655 $X2=0 $Y2=0
cc_43 N_A_c_44_n N_SLEEP_M1001_g 0.00938378f $X=1.15 $Y=1.645 $X2=0 $Y2=0
cc_44 N_A_c_46_n N_SLEEP_M1001_g 0.0171659f $X=1.17 $Y=0.96 $X2=0 $Y2=0
cc_45 A N_SLEEP_M1001_g 4.46117e-19 $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_46 N_A_c_44_n N_SLEEP_c_83_n 4.97555e-19 $X=1.15 $Y=1.645 $X2=0 $Y2=0
cc_47 A N_SLEEP_c_83_n 0.0282905f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_48 N_A_c_44_n N_SLEEP_c_81_n 0.0519587f $X=1.15 $Y=1.645 $X2=0 $Y2=0
cc_49 A N_SLEEP_c_81_n 0.00161646f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_50 N_A_M1005_g N_A_161_489#_c_126_n 0.0184025f $X=1.15 $Y=2.655 $X2=0 $Y2=0
cc_51 N_A_M1005_g N_A_161_489#_c_127_n 0.010818f $X=1.15 $Y=2.655 $X2=0 $Y2=0
cc_52 A N_A_161_489#_c_127_n 0.00780975f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_53 N_A_c_44_n N_A_161_489#_c_128_n 0.00183499f $X=1.15 $Y=1.645 $X2=0 $Y2=0
cc_54 N_A_M1005_g N_A_161_489#_c_128_n 0.00423371f $X=1.15 $Y=2.655 $X2=0 $Y2=0
cc_55 A N_A_161_489#_c_128_n 0.0260029f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_56 N_A_c_46_n N_A_161_489#_c_120_n 0.00377352f $X=1.17 $Y=0.96 $X2=0 $Y2=0
cc_57 N_A_c_44_n N_A_161_489#_c_122_n 0.00533946f $X=1.15 $Y=1.645 $X2=0 $Y2=0
cc_58 A N_A_161_489#_c_122_n 8.46245e-19 $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_59 N_A_M1005_g N_VPWR_c_183_n 0.00228737f $X=1.15 $Y=2.655 $X2=0 $Y2=0
cc_60 N_A_M1005_g N_VPWR_c_184_n 0.00489592f $X=1.15 $Y=2.655 $X2=0 $Y2=0
cc_61 N_A_M1005_g N_VPWR_c_182_n 0.00515964f $X=1.15 $Y=2.655 $X2=0 $Y2=0
cc_62 N_A_c_43_n N_VGND_c_221_n 0.0124306f $X=0.81 $Y=0.96 $X2=0 $Y2=0
cc_63 N_A_c_44_n N_VGND_c_221_n 8.10401e-19 $X=1.15 $Y=1.645 $X2=0 $Y2=0
cc_64 N_A_c_46_n N_VGND_c_221_n 0.0016536f $X=1.17 $Y=0.96 $X2=0 $Y2=0
cc_65 A N_VGND_c_221_n 0.00995469f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_66 N_A_c_43_n N_VGND_c_224_n 0.00424179f $X=0.81 $Y=0.96 $X2=0 $Y2=0
cc_67 N_A_c_46_n N_VGND_c_224_n 0.00510437f $X=1.17 $Y=0.96 $X2=0 $Y2=0
cc_68 N_A_c_43_n N_VGND_c_226_n 0.0043341f $X=0.81 $Y=0.96 $X2=0 $Y2=0
cc_69 N_A_c_46_n N_VGND_c_226_n 0.00515964f $X=1.17 $Y=0.96 $X2=0 $Y2=0
cc_70 N_SLEEP_M1009_g N_A_161_489#_c_118_n 0.0280814f $X=1.96 $Y=0.675 $X2=0
+ $Y2=0
cc_71 N_SLEEP_M1000_g N_A_161_489#_c_126_n 0.00227848f $X=1.51 $Y=2.655 $X2=0
+ $Y2=0
cc_72 N_SLEEP_M1000_g N_A_161_489#_c_127_n 0.0160247f $X=1.51 $Y=2.655 $X2=0
+ $Y2=0
cc_73 N_SLEEP_c_83_n N_A_161_489#_c_127_n 0.0460501f $X=1.94 $Y=1.48 $X2=0 $Y2=0
cc_74 N_SLEEP_c_81_n N_A_161_489#_c_127_n 0.0027233f $X=1.96 $Y=1.48 $X2=0 $Y2=0
cc_75 N_SLEEP_M1001_g N_A_161_489#_c_120_n 0.00370726f $X=1.6 $Y=0.675 $X2=0
+ $Y2=0
cc_76 N_SLEEP_M1001_g N_A_161_489#_c_121_n 0.0140103f $X=1.6 $Y=0.675 $X2=0
+ $Y2=0
cc_77 N_SLEEP_M1009_g N_A_161_489#_c_121_n 0.01362f $X=1.96 $Y=0.675 $X2=0 $Y2=0
cc_78 N_SLEEP_c_83_n N_A_161_489#_c_121_n 0.0459044f $X=1.94 $Y=1.48 $X2=0 $Y2=0
cc_79 N_SLEEP_c_81_n N_A_161_489#_c_121_n 0.00330876f $X=1.96 $Y=1.48 $X2=0
+ $Y2=0
cc_80 N_SLEEP_c_83_n N_A_161_489#_c_122_n 0.00463681f $X=1.94 $Y=1.48 $X2=0
+ $Y2=0
cc_81 N_SLEEP_c_81_n N_A_161_489#_c_122_n 0.00158276f $X=1.96 $Y=1.48 $X2=0
+ $Y2=0
cc_82 N_SLEEP_M1009_g N_A_161_489#_c_151_n 7.7944e-19 $X=1.96 $Y=0.675 $X2=0
+ $Y2=0
cc_83 N_SLEEP_c_83_n N_A_161_489#_c_151_n 0.0241847f $X=1.94 $Y=1.48 $X2=0 $Y2=0
cc_84 N_SLEEP_c_81_n N_A_161_489#_c_151_n 0.0013583f $X=1.96 $Y=1.48 $X2=0 $Y2=0
cc_85 N_SLEEP_c_83_n N_A_161_489#_c_123_n 0.00338649f $X=1.94 $Y=1.48 $X2=0
+ $Y2=0
cc_86 N_SLEEP_c_81_n N_A_161_489#_c_123_n 0.0223211f $X=1.96 $Y=1.48 $X2=0 $Y2=0
cc_87 N_SLEEP_M1000_g N_VPWR_c_183_n 0.0199846f $X=1.51 $Y=2.655 $X2=0 $Y2=0
cc_88 N_SLEEP_M1000_g N_VPWR_c_184_n 0.00424179f $X=1.51 $Y=2.655 $X2=0 $Y2=0
cc_89 N_SLEEP_M1000_g N_VPWR_c_182_n 0.0043341f $X=1.51 $Y=2.655 $X2=0 $Y2=0
cc_90 N_SLEEP_M1001_g N_VGND_c_222_n 0.00165191f $X=1.6 $Y=0.675 $X2=0 $Y2=0
cc_91 N_SLEEP_M1009_g N_VGND_c_222_n 0.0111446f $X=1.96 $Y=0.675 $X2=0 $Y2=0
cc_92 N_SLEEP_M1001_g N_VGND_c_224_n 0.00510437f $X=1.6 $Y=0.675 $X2=0 $Y2=0
cc_93 N_SLEEP_M1009_g N_VGND_c_224_n 0.00424179f $X=1.96 $Y=0.675 $X2=0 $Y2=0
cc_94 N_SLEEP_M1001_g N_VGND_c_226_n 0.00515964f $X=1.6 $Y=0.675 $X2=0 $Y2=0
cc_95 N_SLEEP_M1009_g N_VGND_c_226_n 0.0043341f $X=1.96 $Y=0.675 $X2=0 $Y2=0
cc_96 N_A_161_489#_c_127_n N_VPWR_M1000_d 0.00938962f $X=2.35 $Y=2.04 $X2=-0.19
+ $Y2=-0.245
cc_97 N_A_161_489#_M1003_g N_VPWR_c_183_n 0.0266547f $X=2.39 $Y=2.465 $X2=0
+ $Y2=0
cc_98 N_A_161_489#_M1006_g N_VPWR_c_183_n 0.00363785f $X=2.75 $Y=2.465 $X2=0
+ $Y2=0
cc_99 N_A_161_489#_c_126_n N_VPWR_c_183_n 0.0185956f $X=0.935 $Y=2.655 $X2=0
+ $Y2=0
cc_100 N_A_161_489#_c_127_n N_VPWR_c_183_n 0.0617576f $X=2.35 $Y=2.04 $X2=0
+ $Y2=0
cc_101 N_A_161_489#_c_126_n N_VPWR_c_184_n 0.00780098f $X=0.935 $Y=2.655 $X2=0
+ $Y2=0
cc_102 N_A_161_489#_M1003_g N_VPWR_c_185_n 0.00388479f $X=2.39 $Y=2.465 $X2=0
+ $Y2=0
cc_103 N_A_161_489#_M1006_g N_VPWR_c_185_n 0.00585385f $X=2.75 $Y=2.465 $X2=0
+ $Y2=0
cc_104 N_A_161_489#_M1003_g N_VPWR_c_182_n 0.006597f $X=2.39 $Y=2.465 $X2=0
+ $Y2=0
cc_105 N_A_161_489#_M1006_g N_VPWR_c_182_n 0.0116999f $X=2.75 $Y=2.465 $X2=0
+ $Y2=0
cc_106 N_A_161_489#_c_126_n N_VPWR_c_182_n 0.0108571f $X=0.935 $Y=2.655 $X2=0
+ $Y2=0
cc_107 N_A_161_489#_c_127_n A_493_367# 0.00433061f $X=2.35 $Y=2.04 $X2=-0.19
+ $Y2=-0.245
cc_108 N_A_161_489#_c_119_n N_X_c_211_n 0.0325138f $X=2.75 $Y=1.005 $X2=0 $Y2=0
cc_109 N_A_161_489#_c_169_p N_X_c_211_n 0.0145272f $X=2.517 $Y=1.18 $X2=0 $Y2=0
cc_110 N_A_161_489#_c_151_n N_X_c_211_n 0.0572537f $X=2.517 $Y=1.955 $X2=0 $Y2=0
cc_111 N_A_161_489#_c_120_n N_VGND_c_221_n 0.00635101f $X=1.385 $Y=0.72 $X2=0
+ $Y2=0
cc_112 N_A_161_489#_c_118_n N_VGND_c_222_n 0.0111236f $X=2.39 $Y=1.17 $X2=0
+ $Y2=0
cc_113 N_A_161_489#_c_119_n N_VGND_c_222_n 0.00170417f $X=2.75 $Y=1.005 $X2=0
+ $Y2=0
cc_114 N_A_161_489#_c_120_n N_VGND_c_222_n 0.00643814f $X=1.385 $Y=0.72 $X2=0
+ $Y2=0
cc_115 N_A_161_489#_c_121_n N_VGND_c_222_n 0.0216087f $X=2.35 $Y=1.095 $X2=0
+ $Y2=0
cc_116 N_A_161_489#_c_120_n N_VGND_c_224_n 0.00680149f $X=1.385 $Y=0.72 $X2=0
+ $Y2=0
cc_117 N_A_161_489#_c_118_n N_VGND_c_225_n 0.00424179f $X=2.39 $Y=1.17 $X2=0
+ $Y2=0
cc_118 N_A_161_489#_c_119_n N_VGND_c_225_n 0.00510437f $X=2.75 $Y=1.005 $X2=0
+ $Y2=0
cc_119 N_A_161_489#_c_118_n N_VGND_c_226_n 0.0043341f $X=2.39 $Y=1.17 $X2=0
+ $Y2=0
cc_120 N_A_161_489#_c_119_n N_VGND_c_226_n 0.00515964f $X=2.75 $Y=1.005 $X2=0
+ $Y2=0
cc_121 N_A_161_489#_c_120_n N_VGND_c_226_n 0.00725225f $X=1.385 $Y=0.72 $X2=0
+ $Y2=0
cc_122 N_VPWR_c_182_n A_493_367# 0.00899413f $X=3.12 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_123 N_VPWR_c_182_n N_X_M1006_d 0.00319521f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_124 N_VPWR_c_185_n N_X_c_211_n 0.0287379f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_125 N_VPWR_c_182_n N_X_c_211_n 0.0162509f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_126 N_X_c_211_n N_VGND_c_225_n 0.0121076f $X=2.965 $Y=0.72 $X2=0 $Y2=0
cc_127 N_X_c_211_n N_VGND_c_226_n 0.0143287f $X=2.965 $Y=0.72 $X2=0 $Y2=0
