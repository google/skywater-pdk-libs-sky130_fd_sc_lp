* File: sky130_fd_sc_lp__and4_lp.pxi.spice
* Created: Fri Aug 28 10:08:01 2020
* 
x_PM_SKY130_FD_SC_LP__AND4_LP%D N_D_M1005_g N_D_c_88_n N_D_c_89_n N_D_M1004_g
+ N_D_M1000_g N_D_c_95_n D D D N_D_c_92_n PM_SKY130_FD_SC_LP__AND4_LP%D
x_PM_SKY130_FD_SC_LP__AND4_LP%C N_C_M1011_g N_C_M1014_g N_C_M1015_g N_C_c_131_n
+ N_C_c_132_n C C C C N_C_c_134_n PM_SKY130_FD_SC_LP__AND4_LP%C
x_PM_SKY130_FD_SC_LP__AND4_LP%B N_B_M1001_g N_B_c_185_n N_B_M1007_g N_B_M1003_g
+ N_B_c_191_n B B B B N_B_c_187_n PM_SKY130_FD_SC_LP__AND4_LP%B
x_PM_SKY130_FD_SC_LP__AND4_LP%A N_A_c_239_n N_A_M1002_g N_A_c_240_n N_A_c_241_n
+ N_A_c_246_n N_A_c_247_n N_A_M1013_g N_A_c_248_n N_A_c_249_n N_A_M1012_g
+ N_A_c_242_n N_A_c_243_n N_A_c_251_n N_A_c_252_n A A N_A_c_245_n
+ PM_SKY130_FD_SC_LP__AND4_LP%A
x_PM_SKY130_FD_SC_LP__AND4_LP%A_186_485# N_A_186_485#_M1002_d
+ N_A_186_485#_M1004_d N_A_186_485#_M1003_d N_A_186_485#_M1006_g
+ N_A_186_485#_M1008_g N_A_186_485#_M1010_g N_A_186_485#_M1009_g
+ N_A_186_485#_c_325_n N_A_186_485#_c_326_n N_A_186_485#_c_315_n
+ N_A_186_485#_c_327_n N_A_186_485#_c_316_n N_A_186_485#_c_317_n
+ N_A_186_485#_c_328_n N_A_186_485#_c_318_n N_A_186_485#_c_319_n
+ N_A_186_485#_c_320_n N_A_186_485#_c_330_n N_A_186_485#_c_331_n
+ N_A_186_485#_c_332_n N_A_186_485#_c_321_n N_A_186_485#_c_322_n
+ PM_SKY130_FD_SC_LP__AND4_LP%A_186_485#
x_PM_SKY130_FD_SC_LP__AND4_LP%VPWR N_VPWR_M1005_s N_VPWR_M1015_d N_VPWR_M1012_d
+ N_VPWR_c_433_n N_VPWR_c_434_n N_VPWR_c_435_n N_VPWR_c_436_n N_VPWR_c_437_n
+ N_VPWR_c_438_n VPWR N_VPWR_c_439_n N_VPWR_c_440_n N_VPWR_c_432_n
+ N_VPWR_c_442_n PM_SKY130_FD_SC_LP__AND4_LP%VPWR
x_PM_SKY130_FD_SC_LP__AND4_LP%X N_X_M1010_d N_X_M1009_d X X X X X X X
+ N_X_c_488_n PM_SKY130_FD_SC_LP__AND4_LP%X
x_PM_SKY130_FD_SC_LP__AND4_LP%VGND N_VGND_M1000_s N_VGND_M1006_s N_VGND_c_507_n
+ N_VGND_c_508_n N_VGND_c_509_n N_VGND_c_510_n VGND N_VGND_c_511_n
+ N_VGND_c_512_n N_VGND_c_513_n N_VGND_c_514_n PM_SKY130_FD_SC_LP__AND4_LP%VGND
cc_1 VNB N_D_c_88_n 0.0295887f $X=-0.19 $Y=-0.245 $X2=1 $Y2=1.315
cc_2 VNB N_D_c_89_n 0.0189522f $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=1.315
cc_3 VNB N_D_M1000_g 0.0515411f $X=-0.19 $Y=-0.245 $X2=1.075 $Y2=0.485
cc_4 VNB D 0.0464177f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_5 VNB N_D_c_92_n 0.0227429f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.405
cc_6 VNB N_C_M1014_g 0.0303919f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=1.91
cc_7 VNB N_C_c_131_n 0.0232486f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.835
cc_8 VNB N_C_c_132_n 0.00725972f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB C 0.00849603f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_C_c_134_n 0.0147433f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_B_M1001_g 0.0392588f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.635
cc_12 VNB N_B_c_185_n 0.0232429f $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=1.315
cc_13 VNB B 0.0042636f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=1.835
cc_14 VNB N_B_c_187_n 0.0185675f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_c_239_n 0.0198632f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.91
cc_16 VNB N_A_c_240_n 0.0332627f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_c_241_n 0.0127142f $X=-0.19 $Y=-0.245 $X2=1 $Y2=1.315
cc_18 VNB N_A_c_242_n 0.0181159f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.76
cc_19 VNB N_A_c_243_n 0.0189688f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=1.835
cc_20 VNB A 0.00987627f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.95
cc_21 VNB N_A_c_245_n 0.0162489f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_186_485#_M1006_g 0.0237572f $X=-0.19 $Y=-0.245 $X2=1.075 $Y2=0.485
cc_23 VNB N_A_186_485#_M1008_g 0.00553415f $X=-0.19 $Y=-0.245 $X2=0.495
+ $Y2=1.835
cc_24 VNB N_A_186_485#_M1010_g 0.0245438f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=1.835
cc_25 VNB N_A_186_485#_M1009_g 0.00555131f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.95
cc_26 VNB N_A_186_485#_c_315_n 0.00853486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_186_485#_c_316_n 0.0182736f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_186_485#_c_317_n 0.00440257f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_186_485#_c_318_n 0.00286098f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=1.665
cc_30 VNB N_A_186_485#_c_319_n 0.00322403f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_186_485#_c_320_n 0.00139017f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=2.035
cc_32 VNB N_A_186_485#_c_321_n 0.09109f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_186_485#_c_322_n 0.00140986f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VPWR_c_432_n 0.203486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB X 0.0478938f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=2.635
cc_36 VNB N_X_c_488_n 0.032864f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.405
cc_37 VNB N_VGND_c_507_n 0.0287737f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=2.635
cc_38 VNB N_VGND_c_508_n 0.0116374f $X=-0.19 $Y=-0.245 $X2=1.075 $Y2=0.485
cc_39 VNB N_VGND_c_509_n 0.0609039f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.835
cc_40 VNB N_VGND_c_510_n 0.0054376f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_511_n 0.0207592f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=1.835
cc_42 VNB N_VGND_c_512_n 0.0378037f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.405
cc_43 VNB N_VGND_c_513_n 0.314364f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=1.295
cc_44 VNB N_VGND_c_514_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VPB N_D_M1005_g 0.0457572f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=2.635
cc_46 VPB N_D_M1004_g 0.0346642f $X=-0.19 $Y=1.655 $X2=0.855 $Y2=2.635
cc_47 VPB N_D_c_95_n 0.0196429f $X=-0.19 $Y=1.655 $X2=0.855 $Y2=1.835
cc_48 VPB D 0.0349274f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_49 VPB N_D_c_92_n 0.00861426f $X=-0.19 $Y=1.655 $X2=0.585 $Y2=1.405
cc_50 VPB N_C_M1011_g 0.0394837f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=2.635
cc_51 VPB N_C_M1015_g 0.0397231f $X=-0.19 $Y=1.655 $X2=1.075 $Y2=1.24
cc_52 VPB N_C_c_132_n 0.0113521f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_53 VPB C 0.00431719f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_54 VPB N_B_c_185_n 0.00469634f $X=-0.19 $Y=1.655 $X2=0.75 $Y2=1.315
cc_55 VPB N_B_M1007_g 0.0356563f $X=-0.19 $Y=1.655 $X2=0.855 $Y2=2.635
cc_56 VPB N_B_M1003_g 0.0353059f $X=-0.19 $Y=1.655 $X2=1.075 $Y2=0.485
cc_57 VPB N_B_c_191_n 0.027631f $X=-0.19 $Y=1.655 $X2=0.585 $Y2=1.835
cc_58 VPB B 6.36302e-19 $X=-0.19 $Y=1.655 $X2=0.855 $Y2=1.835
cc_59 VPB N_A_c_246_n 0.0160862f $X=-0.19 $Y=1.655 $X2=0.855 $Y2=2.635
cc_60 VPB N_A_c_247_n 0.0152383f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_61 VPB N_A_c_248_n 0.0170484f $X=-0.19 $Y=1.655 $X2=1.075 $Y2=0.485
cc_62 VPB N_A_c_249_n 0.0151025f $X=-0.19 $Y=1.655 $X2=0.585 $Y2=1.39
cc_63 VPB N_A_c_243_n 0.00540481f $X=-0.19 $Y=1.655 $X2=0.855 $Y2=1.835
cc_64 VPB N_A_c_251_n 0.0141458f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_65 VPB N_A_c_252_n 0.00437176f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_66 VPB A 0.00727184f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.95
cc_67 VPB N_A_186_485#_M1008_g 0.0525914f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=1.835
cc_68 VPB N_A_186_485#_M1009_g 0.0564712f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.95
cc_69 VPB N_A_186_485#_c_325_n 0.0296005f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_70 VPB N_A_186_485#_c_326_n 0.00317422f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_71 VPB N_A_186_485#_c_327_n 0.00290479f $X=-0.19 $Y=1.655 $X2=0.585 $Y2=1.405
cc_72 VPB N_A_186_485#_c_328_n 0.0123746f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_73 VPB N_A_186_485#_c_320_n 0.0085894f $X=-0.19 $Y=1.655 $X2=0.48 $Y2=2.035
cc_74 VPB N_A_186_485#_c_330_n 0.00813668f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_75 VPB N_A_186_485#_c_331_n 0.00157764f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_76 VPB N_A_186_485#_c_332_n 0.00309939f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_77 VPB N_VPWR_c_433_n 0.0121909f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_78 VPB N_VPWR_c_434_n 0.0400385f $X=-0.19 $Y=1.655 $X2=1.075 $Y2=0.485
cc_79 VPB N_VPWR_c_435_n 0.0159245f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=1.835
cc_80 VPB N_VPWR_c_436_n 0.0161363f $X=-0.19 $Y=1.655 $X2=0.855 $Y2=1.835
cc_81 VPB N_VPWR_c_437_n 0.0376698f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_82 VPB N_VPWR_c_438_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.95
cc_83 VPB N_VPWR_c_439_n 0.0376698f $X=-0.19 $Y=1.655 $X2=0.585 $Y2=1.405
cc_84 VPB N_VPWR_c_440_n 0.0355107f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_85 VPB N_VPWR_c_432_n 0.122531f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_86 VPB N_VPWR_c_442_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_87 VPB X 0.0790269f $X=-0.19 $Y=1.655 $X2=0.855 $Y2=2.635
cc_88 N_D_M1004_g N_C_M1011_g 0.0184472f $X=0.855 $Y=2.635 $X2=0 $Y2=0
cc_89 D N_C_M1011_g 0.00152595f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_90 N_D_M1000_g N_C_M1014_g 0.0342341f $X=1.075 $Y=0.485 $X2=0 $Y2=0
cc_91 D N_C_c_131_n 6.70584e-19 $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_92 N_D_c_92_n N_C_c_131_n 0.00284682f $X=0.585 $Y=1.405 $X2=0 $Y2=0
cc_93 N_D_c_95_n N_C_c_132_n 0.0184472f $X=0.855 $Y=1.835 $X2=0 $Y2=0
cc_94 D N_C_c_132_n 4.97845e-19 $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_95 N_D_c_92_n N_C_c_132_n 0.00290169f $X=0.585 $Y=1.405 $X2=0 $Y2=0
cc_96 N_D_c_88_n C 0.00652285f $X=1 $Y=1.315 $X2=0 $Y2=0
cc_97 N_D_M1000_g C 0.0372319f $X=1.075 $Y=0.485 $X2=0 $Y2=0
cc_98 D C 0.0410367f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_99 N_D_c_92_n C 0.00154428f $X=0.585 $Y=1.405 $X2=0 $Y2=0
cc_100 N_D_c_88_n N_C_c_134_n 0.0342341f $X=1 $Y=1.315 $X2=0 $Y2=0
cc_101 N_D_c_88_n N_A_186_485#_c_326_n 8.4008e-19 $X=1 $Y=1.315 $X2=0 $Y2=0
cc_102 N_D_M1004_g N_A_186_485#_c_326_n 0.00311199f $X=0.855 $Y=2.635 $X2=0
+ $Y2=0
cc_103 D N_A_186_485#_c_326_n 0.00602937f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_104 N_D_M1005_g N_A_186_485#_c_330_n 0.00125204f $X=0.495 $Y=2.635 $X2=0
+ $Y2=0
cc_105 N_D_M1004_g N_A_186_485#_c_330_n 0.00959421f $X=0.855 $Y=2.635 $X2=0
+ $Y2=0
cc_106 N_D_M1004_g N_A_186_485#_c_331_n 0.00363396f $X=0.855 $Y=2.635 $X2=0
+ $Y2=0
cc_107 N_D_M1005_g N_VPWR_c_434_n 0.013834f $X=0.495 $Y=2.635 $X2=0 $Y2=0
cc_108 N_D_M1004_g N_VPWR_c_434_n 0.00180376f $X=0.855 $Y=2.635 $X2=0 $Y2=0
cc_109 D N_VPWR_c_434_n 0.0221756f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_110 N_D_M1005_g N_VPWR_c_437_n 0.00413255f $X=0.495 $Y=2.635 $X2=0 $Y2=0
cc_111 N_D_M1004_g N_VPWR_c_437_n 0.00476381f $X=0.855 $Y=2.635 $X2=0 $Y2=0
cc_112 N_D_M1005_g N_VPWR_c_432_n 0.00428305f $X=0.495 $Y=2.635 $X2=0 $Y2=0
cc_113 N_D_M1004_g N_VPWR_c_432_n 0.00509887f $X=0.855 $Y=2.635 $X2=0 $Y2=0
cc_114 N_D_c_88_n N_VGND_c_507_n 0.00226844f $X=1 $Y=1.315 $X2=0 $Y2=0
cc_115 N_D_c_89_n N_VGND_c_507_n 0.00152148f $X=0.75 $Y=1.315 $X2=0 $Y2=0
cc_116 N_D_M1000_g N_VGND_c_507_n 0.017151f $X=1.075 $Y=0.485 $X2=0 $Y2=0
cc_117 D N_VGND_c_507_n 0.0115263f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_118 N_D_M1000_g N_VGND_c_509_n 0.00468089f $X=1.075 $Y=0.485 $X2=0 $Y2=0
cc_119 N_D_M1000_g N_VGND_c_513_n 0.0091487f $X=1.075 $Y=0.485 $X2=0 $Y2=0
cc_120 N_C_M1014_g N_B_M1001_g 0.0252224f $X=1.465 $Y=0.485 $X2=0 $Y2=0
cc_121 C N_B_M1001_g 0.0096672f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_122 N_C_c_134_n N_B_M1001_g 0.0100096f $X=1.555 $Y=1.275 $X2=0 $Y2=0
cc_123 N_C_c_132_n N_B_c_185_n 0.0100096f $X=1.645 $Y=1.705 $X2=0 $Y2=0
cc_124 N_C_M1015_g N_B_M1007_g 0.0345393f $X=1.645 $Y=2.635 $X2=0 $Y2=0
cc_125 N_C_M1015_g N_B_c_191_n 0.0100096f $X=1.645 $Y=2.635 $X2=0 $Y2=0
cc_126 N_C_M1014_g B 5.93888e-19 $X=1.465 $Y=0.485 $X2=0 $Y2=0
cc_127 N_C_M1015_g B 5.41769e-19 $X=1.645 $Y=2.635 $X2=0 $Y2=0
cc_128 C B 0.112322f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_129 N_C_c_134_n B 7.25073e-19 $X=1.555 $Y=1.275 $X2=0 $Y2=0
cc_130 N_C_c_131_n N_B_c_187_n 0.0100096f $X=1.555 $Y=1.63 $X2=0 $Y2=0
cc_131 N_C_M1011_g N_A_186_485#_c_325_n 0.0112168f $X=1.285 $Y=2.635 $X2=0 $Y2=0
cc_132 N_C_M1015_g N_A_186_485#_c_325_n 0.0144463f $X=1.645 $Y=2.635 $X2=0 $Y2=0
cc_133 C N_A_186_485#_c_325_n 0.0295493f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_134 N_C_M1011_g N_A_186_485#_c_326_n 0.00211986f $X=1.285 $Y=2.635 $X2=0
+ $Y2=0
cc_135 C N_A_186_485#_c_326_n 0.0094831f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_136 N_C_M1011_g N_A_186_485#_c_330_n 0.00844904f $X=1.285 $Y=2.635 $X2=0
+ $Y2=0
cc_137 N_C_M1011_g N_A_186_485#_c_331_n 0.00395284f $X=1.285 $Y=2.635 $X2=0
+ $Y2=0
cc_138 N_C_M1015_g N_A_186_485#_c_331_n 0.00210733f $X=1.645 $Y=2.635 $X2=0
+ $Y2=0
cc_139 N_C_M1011_g N_VPWR_c_435_n 0.00180376f $X=1.285 $Y=2.635 $X2=0 $Y2=0
cc_140 N_C_M1015_g N_VPWR_c_435_n 0.0122162f $X=1.645 $Y=2.635 $X2=0 $Y2=0
cc_141 N_C_M1011_g N_VPWR_c_437_n 0.00476381f $X=1.285 $Y=2.635 $X2=0 $Y2=0
cc_142 N_C_M1015_g N_VPWR_c_437_n 0.00413255f $X=1.645 $Y=2.635 $X2=0 $Y2=0
cc_143 N_C_M1011_g N_VPWR_c_432_n 0.00509887f $X=1.285 $Y=2.635 $X2=0 $Y2=0
cc_144 N_C_M1015_g N_VPWR_c_432_n 0.00428305f $X=1.645 $Y=2.635 $X2=0 $Y2=0
cc_145 C N_VGND_c_507_n 0.0226587f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_146 N_C_M1014_g N_VGND_c_509_n 0.00364003f $X=1.465 $Y=0.485 $X2=0 $Y2=0
cc_147 C N_VGND_c_509_n 0.0195413f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_148 N_C_M1014_g N_VGND_c_513_n 0.00535522f $X=1.465 $Y=0.485 $X2=0 $Y2=0
cc_149 C N_VGND_c_513_n 0.0236192f $X=1.115 $Y=0.47 $X2=0 $Y2=0
cc_150 C A_230_55# 0.00175001f $X=1.115 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_151 C A_308_55# 0.00589388f $X=1.115 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_152 N_B_M1001_g N_A_c_239_n 0.0423846f $X=2.035 $Y=0.485 $X2=-0.19 $Y2=-0.245
cc_153 B N_A_c_239_n 0.00296994f $X=2.075 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_154 N_B_M1003_g N_A_c_246_n 0.0202114f $X=2.435 $Y=2.635 $X2=0 $Y2=0
cc_155 N_B_M1001_g N_A_c_242_n 0.00254917f $X=2.035 $Y=0.485 $X2=0 $Y2=0
cc_156 B N_A_c_242_n 0.00296068f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_157 N_B_c_187_n N_A_c_242_n 0.00498947f $X=2.13 $Y=1.36 $X2=0 $Y2=0
cc_158 N_B_c_191_n N_A_c_243_n 0.0202114f $X=2.435 $Y=1.79 $X2=0 $Y2=0
cc_159 N_B_c_191_n A 0.00270914f $X=2.435 $Y=1.79 $X2=0 $Y2=0
cc_160 B A 0.0430835f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_161 N_B_c_187_n A 0.00460162f $X=2.13 $Y=1.36 $X2=0 $Y2=0
cc_162 N_B_c_185_n N_A_c_245_n 0.00498947f $X=2.127 $Y=1.715 $X2=0 $Y2=0
cc_163 B N_A_c_245_n 5.28372e-19 $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_164 N_B_M1007_g N_A_186_485#_c_325_n 0.0139944f $X=2.075 $Y=2.635 $X2=0 $Y2=0
cc_165 N_B_M1003_g N_A_186_485#_c_325_n 0.0140031f $X=2.435 $Y=2.635 $X2=0 $Y2=0
cc_166 N_B_c_191_n N_A_186_485#_c_325_n 6.71602e-19 $X=2.435 $Y=1.79 $X2=0 $Y2=0
cc_167 B N_A_186_485#_c_325_n 0.0226028f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_168 N_B_M1001_g N_A_186_485#_c_315_n 0.00126053f $X=2.035 $Y=0.485 $X2=0
+ $Y2=0
cc_169 B N_A_186_485#_c_315_n 0.02343f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_170 N_B_M1007_g N_A_186_485#_c_327_n 0.00210156f $X=2.075 $Y=2.635 $X2=0
+ $Y2=0
cc_171 N_B_M1003_g N_A_186_485#_c_327_n 0.0133586f $X=2.435 $Y=2.635 $X2=0 $Y2=0
cc_172 N_B_M1001_g N_A_186_485#_c_317_n 3.84419e-19 $X=2.035 $Y=0.485 $X2=0
+ $Y2=0
cc_173 N_B_c_191_n N_A_186_485#_c_317_n 0.00102146f $X=2.435 $Y=1.79 $X2=0 $Y2=0
cc_174 B N_A_186_485#_c_317_n 0.0141182f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_175 N_B_M1003_g N_A_186_485#_c_332_n 0.00357037f $X=2.435 $Y=2.635 $X2=0
+ $Y2=0
cc_176 N_B_M1007_g N_VPWR_c_435_n 0.0122162f $X=2.075 $Y=2.635 $X2=0 $Y2=0
cc_177 N_B_M1003_g N_VPWR_c_435_n 0.00180376f $X=2.435 $Y=2.635 $X2=0 $Y2=0
cc_178 N_B_M1007_g N_VPWR_c_439_n 0.00413255f $X=2.075 $Y=2.635 $X2=0 $Y2=0
cc_179 N_B_M1003_g N_VPWR_c_439_n 0.00476381f $X=2.435 $Y=2.635 $X2=0 $Y2=0
cc_180 N_B_M1007_g N_VPWR_c_432_n 0.00428305f $X=2.075 $Y=2.635 $X2=0 $Y2=0
cc_181 N_B_M1003_g N_VPWR_c_432_n 0.00509887f $X=2.435 $Y=2.635 $X2=0 $Y2=0
cc_182 N_B_M1001_g N_VGND_c_509_n 0.00371265f $X=2.035 $Y=0.485 $X2=0 $Y2=0
cc_183 B N_VGND_c_509_n 0.00929408f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_184 N_B_M1001_g N_VGND_c_513_n 0.00557027f $X=2.035 $Y=0.485 $X2=0 $Y2=0
cc_185 B N_VGND_c_513_n 0.0107116f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_186 B A_422_55# 0.00179236f $X=2.075 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_187 N_A_c_240_n N_A_186_485#_M1006_g 0.00427478f $X=2.79 $Y=0.88 $X2=0 $Y2=0
cc_188 N_A_c_246_n N_A_186_485#_M1008_g 0.00291108f $X=2.865 $Y=2.165 $X2=0
+ $Y2=0
cc_189 N_A_c_248_n N_A_186_485#_M1008_g 0.0193856f $X=3.15 $Y=2.24 $X2=0 $Y2=0
cc_190 N_A_c_243_n N_A_186_485#_M1008_g 0.00656604f $X=2.955 $Y=1.73 $X2=0 $Y2=0
cc_191 N_A_c_239_n N_A_186_485#_c_315_n 0.0104165f $X=2.425 $Y=0.805 $X2=0 $Y2=0
cc_192 N_A_c_240_n N_A_186_485#_c_315_n 0.0107318f $X=2.79 $Y=0.88 $X2=0 $Y2=0
cc_193 N_A_c_241_n N_A_186_485#_c_315_n 8.17915e-19 $X=2.5 $Y=0.88 $X2=0 $Y2=0
cc_194 N_A_c_247_n N_A_186_485#_c_327_n 0.0110345f $X=2.865 $Y=2.315 $X2=0 $Y2=0
cc_195 N_A_c_249_n N_A_186_485#_c_327_n 0.00169843f $X=3.225 $Y=2.315 $X2=0
+ $Y2=0
cc_196 N_A_c_252_n N_A_186_485#_c_327_n 0.00466277f $X=2.865 $Y=2.24 $X2=0 $Y2=0
cc_197 N_A_c_240_n N_A_186_485#_c_316_n 0.00715309f $X=2.79 $Y=0.88 $X2=0 $Y2=0
cc_198 N_A_c_242_n N_A_186_485#_c_316_n 0.00481178f $X=2.955 $Y=1.225 $X2=0
+ $Y2=0
cc_199 A N_A_186_485#_c_316_n 0.0341444f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_200 N_A_c_245_n N_A_186_485#_c_316_n 0.00467405f $X=2.955 $Y=1.39 $X2=0 $Y2=0
cc_201 N_A_c_240_n N_A_186_485#_c_317_n 0.00667524f $X=2.79 $Y=0.88 $X2=0 $Y2=0
cc_202 N_A_c_241_n N_A_186_485#_c_317_n 0.00113402f $X=2.5 $Y=0.88 $X2=0 $Y2=0
cc_203 N_A_c_242_n N_A_186_485#_c_317_n 0.00203373f $X=2.955 $Y=1.225 $X2=0
+ $Y2=0
cc_204 A N_A_186_485#_c_317_n 0.0259524f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_205 N_A_c_246_n N_A_186_485#_c_328_n 0.00477433f $X=2.865 $Y=2.165 $X2=0
+ $Y2=0
cc_206 N_A_c_248_n N_A_186_485#_c_328_n 0.0218626f $X=3.15 $Y=2.24 $X2=0 $Y2=0
cc_207 N_A_c_251_n N_A_186_485#_c_328_n 0.00121357f $X=2.955 $Y=1.895 $X2=0
+ $Y2=0
cc_208 N_A_c_252_n N_A_186_485#_c_328_n 0.00629013f $X=2.865 $Y=2.24 $X2=0 $Y2=0
cc_209 A N_A_186_485#_c_328_n 0.0333863f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_210 N_A_c_242_n N_A_186_485#_c_319_n 0.00313734f $X=2.955 $Y=1.225 $X2=0
+ $Y2=0
cc_211 A N_A_186_485#_c_319_n 0.0581159f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_212 N_A_c_245_n N_A_186_485#_c_319_n 6.15659e-19 $X=2.955 $Y=1.39 $X2=0 $Y2=0
cc_213 N_A_c_246_n N_A_186_485#_c_320_n 0.0028256f $X=2.865 $Y=2.165 $X2=0 $Y2=0
cc_214 N_A_c_251_n N_A_186_485#_c_320_n 6.15659e-19 $X=2.955 $Y=1.895 $X2=0
+ $Y2=0
cc_215 N_A_c_246_n N_A_186_485#_c_332_n 0.00175047f $X=2.865 $Y=2.165 $X2=0
+ $Y2=0
cc_216 N_A_c_252_n N_A_186_485#_c_332_n 9.97332e-19 $X=2.865 $Y=2.24 $X2=0 $Y2=0
cc_217 A N_A_186_485#_c_332_n 0.0267962f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_218 N_A_c_242_n N_A_186_485#_c_321_n 0.00427478f $X=2.955 $Y=1.225 $X2=0
+ $Y2=0
cc_219 A N_A_186_485#_c_321_n 0.00122026f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_220 N_A_c_245_n N_A_186_485#_c_321_n 0.0121241f $X=2.955 $Y=1.39 $X2=0 $Y2=0
cc_221 N_A_c_243_n N_A_186_485#_c_322_n 6.15659e-19 $X=2.955 $Y=1.73 $X2=0 $Y2=0
cc_222 N_A_c_247_n N_VPWR_c_436_n 0.00180376f $X=2.865 $Y=2.315 $X2=0 $Y2=0
cc_223 N_A_c_249_n N_VPWR_c_436_n 0.0122162f $X=3.225 $Y=2.315 $X2=0 $Y2=0
cc_224 N_A_c_247_n N_VPWR_c_439_n 0.00476381f $X=2.865 $Y=2.315 $X2=0 $Y2=0
cc_225 N_A_c_249_n N_VPWR_c_439_n 0.00413255f $X=3.225 $Y=2.315 $X2=0 $Y2=0
cc_226 N_A_c_247_n N_VPWR_c_432_n 0.00509887f $X=2.865 $Y=2.315 $X2=0 $Y2=0
cc_227 N_A_c_249_n N_VPWR_c_432_n 0.00428305f $X=3.225 $Y=2.315 $X2=0 $Y2=0
cc_228 N_A_c_239_n N_VGND_c_508_n 0.002534f $X=2.425 $Y=0.805 $X2=0 $Y2=0
cc_229 N_A_c_239_n N_VGND_c_509_n 0.00511358f $X=2.425 $Y=0.805 $X2=0 $Y2=0
cc_230 N_A_c_239_n N_VGND_c_513_n 0.0105915f $X=2.425 $Y=0.805 $X2=0 $Y2=0
cc_231 N_A_c_240_n N_VGND_c_513_n 0.00355095f $X=2.79 $Y=0.88 $X2=0 $Y2=0
cc_232 N_A_186_485#_c_330_n N_VPWR_c_434_n 0.0153904f $X=1.07 $Y=2.635 $X2=0
+ $Y2=0
cc_233 N_A_186_485#_c_325_n N_VPWR_c_435_n 0.0273053f $X=2.485 $Y=2.15 $X2=0
+ $Y2=0
cc_234 N_A_186_485#_c_327_n N_VPWR_c_435_n 0.0153904f $X=2.65 $Y=2.635 $X2=0
+ $Y2=0
cc_235 N_A_186_485#_c_330_n N_VPWR_c_435_n 0.0153904f $X=1.07 $Y=2.635 $X2=0
+ $Y2=0
cc_236 N_A_186_485#_M1008_g N_VPWR_c_436_n 0.0122661f $X=3.655 $Y=2.635 $X2=0
+ $Y2=0
cc_237 N_A_186_485#_M1009_g N_VPWR_c_436_n 9.38339e-19 $X=4.045 $Y=2.635 $X2=0
+ $Y2=0
cc_238 N_A_186_485#_c_327_n N_VPWR_c_436_n 0.0153904f $X=2.65 $Y=2.635 $X2=0
+ $Y2=0
cc_239 N_A_186_485#_c_328_n N_VPWR_c_436_n 0.0264936f $X=3.405 $Y=2.15 $X2=0
+ $Y2=0
cc_240 N_A_186_485#_c_330_n N_VPWR_c_437_n 0.00971891f $X=1.07 $Y=2.635 $X2=0
+ $Y2=0
cc_241 N_A_186_485#_c_327_n N_VPWR_c_439_n 0.00984895f $X=2.65 $Y=2.635 $X2=0
+ $Y2=0
cc_242 N_A_186_485#_M1008_g N_VPWR_c_440_n 0.00413255f $X=3.655 $Y=2.635 $X2=0
+ $Y2=0
cc_243 N_A_186_485#_M1009_g N_VPWR_c_440_n 0.00364307f $X=4.045 $Y=2.635 $X2=0
+ $Y2=0
cc_244 N_A_186_485#_M1008_g N_VPWR_c_432_n 0.00428305f $X=3.655 $Y=2.635 $X2=0
+ $Y2=0
cc_245 N_A_186_485#_M1009_g N_VPWR_c_432_n 0.00509887f $X=4.045 $Y=2.635 $X2=0
+ $Y2=0
cc_246 N_A_186_485#_c_327_n N_VPWR_c_432_n 0.0111949f $X=2.65 $Y=2.635 $X2=0
+ $Y2=0
cc_247 N_A_186_485#_c_330_n N_VPWR_c_432_n 0.0111118f $X=1.07 $Y=2.635 $X2=0
+ $Y2=0
cc_248 N_A_186_485#_M1006_g X 4.33282e-19 $X=3.525 $Y=0.485 $X2=0 $Y2=0
cc_249 N_A_186_485#_M1008_g X 0.0114066f $X=3.655 $Y=2.635 $X2=0 $Y2=0
cc_250 N_A_186_485#_M1010_g X 0.00378204f $X=3.915 $Y=0.485 $X2=0 $Y2=0
cc_251 N_A_186_485#_M1009_g X 0.0448339f $X=4.045 $Y=2.635 $X2=0 $Y2=0
cc_252 N_A_186_485#_c_328_n X 0.00890613f $X=3.405 $Y=2.15 $X2=0 $Y2=0
cc_253 N_A_186_485#_c_318_n X 0.0134196f $X=3.592 $Y=1.055 $X2=0 $Y2=0
cc_254 N_A_186_485#_c_319_n X 0.0375163f $X=3.592 $Y=1.368 $X2=0 $Y2=0
cc_255 N_A_186_485#_c_320_n X 0.0241114f $X=3.49 $Y=2.065 $X2=0 $Y2=0
cc_256 N_A_186_485#_c_321_n X 0.0383338f $X=3.615 $Y=1.05 $X2=0 $Y2=0
cc_257 N_A_186_485#_M1006_g N_X_c_488_n 0.00169259f $X=3.525 $Y=0.485 $X2=0
+ $Y2=0
cc_258 N_A_186_485#_M1010_g N_X_c_488_n 0.012829f $X=3.915 $Y=0.485 $X2=0 $Y2=0
cc_259 N_A_186_485#_M1006_g N_VGND_c_508_n 0.014393f $X=3.525 $Y=0.485 $X2=0
+ $Y2=0
cc_260 N_A_186_485#_M1010_g N_VGND_c_508_n 0.00216336f $X=3.915 $Y=0.485 $X2=0
+ $Y2=0
cc_261 N_A_186_485#_c_315_n N_VGND_c_508_n 0.0237131f $X=2.64 $Y=0.485 $X2=0
+ $Y2=0
cc_262 N_A_186_485#_c_316_n N_VGND_c_508_n 0.0218374f $X=3.405 $Y=0.97 $X2=0
+ $Y2=0
cc_263 N_A_186_485#_c_318_n N_VGND_c_508_n 0.00624801f $X=3.592 $Y=1.055 $X2=0
+ $Y2=0
cc_264 N_A_186_485#_c_315_n N_VGND_c_509_n 0.0234289f $X=2.64 $Y=0.485 $X2=0
+ $Y2=0
cc_265 N_A_186_485#_M1006_g N_VGND_c_512_n 0.00452967f $X=3.525 $Y=0.485 $X2=0
+ $Y2=0
cc_266 N_A_186_485#_M1010_g N_VGND_c_512_n 0.00509933f $X=3.915 $Y=0.485 $X2=0
+ $Y2=0
cc_267 N_A_186_485#_M1006_g N_VGND_c_513_n 0.00806665f $X=3.525 $Y=0.485 $X2=0
+ $Y2=0
cc_268 N_A_186_485#_M1010_g N_VGND_c_513_n 0.0105289f $X=3.915 $Y=0.485 $X2=0
+ $Y2=0
cc_269 N_A_186_485#_c_315_n N_VGND_c_513_n 0.0126421f $X=2.64 $Y=0.485 $X2=0
+ $Y2=0
cc_270 N_VPWR_c_436_n X 0.0117133f $X=3.44 $Y=2.635 $X2=0 $Y2=0
cc_271 N_VPWR_c_440_n X 0.0227539f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_272 N_VPWR_c_432_n X 0.0245391f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_273 N_X_c_488_n N_VGND_c_508_n 0.0151459f $X=4.32 $Y=0.795 $X2=0 $Y2=0
cc_274 N_X_c_488_n N_VGND_c_512_n 0.0359946f $X=4.32 $Y=0.795 $X2=0 $Y2=0
cc_275 N_X_c_488_n N_VGND_c_513_n 0.0259646f $X=4.32 $Y=0.795 $X2=0 $Y2=0
