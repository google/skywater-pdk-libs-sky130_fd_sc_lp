* File: sky130_fd_sc_lp__a22oi_1.pex.spice
* Created: Fri Aug 28 09:54:52 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A22OI_1%B2 1 3 6 8 9 16
r26 13 16 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=0.45 $Y=1.46
+ $X2=0.665 $Y2=1.46
r27 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.45
+ $Y=1.46 $X2=0.45 $Y2=1.46
r28 9 14 5.4488 $w=4.48e-07 $l=2.05e-07 $layer=LI1_cond $X=0.31 $Y=1.665
+ $X2=0.31 $Y2=1.46
r29 8 14 4.38562 $w=4.48e-07 $l=1.65e-07 $layer=LI1_cond $X=0.31 $Y=1.295
+ $X2=0.31 $Y2=1.46
r30 4 16 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.665 $Y=1.625
+ $X2=0.665 $Y2=1.46
r31 4 6 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=0.665 $Y=1.625
+ $X2=0.665 $Y2=2.465
r32 1 16 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.665 $Y=1.295
+ $X2=0.665 $Y2=1.46
r33 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.665 $Y=1.295
+ $X2=0.665 $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_LP__A22OI_1%B1 3 6 8 9 13 15
c37 13 0 5.1293e-20 $X=1.13 $Y=1.46
c38 6 0 1.18028e-19 $X=1.095 $Y=2.465
r39 13 16 46.3655 $w=3.45e-07 $l=1.65e-07 $layer=POLY_cond $X=1.122 $Y=1.46
+ $X2=1.122 $Y2=1.625
r40 13 15 46.3655 $w=3.45e-07 $l=1.65e-07 $layer=POLY_cond $X=1.122 $Y=1.46
+ $X2=1.122 $Y2=1.295
r41 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.13
+ $Y=1.46 $X2=1.13 $Y2=1.46
r42 9 14 7.74593 $w=3.03e-07 $l=2.05e-07 $layer=LI1_cond $X=1.197 $Y=1.665
+ $X2=1.197 $Y2=1.46
r43 8 14 6.23453 $w=3.03e-07 $l=1.65e-07 $layer=LI1_cond $X=1.197 $Y=1.295
+ $X2=1.197 $Y2=1.46
r44 6 16 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=1.095 $Y=2.465
+ $X2=1.095 $Y2=1.625
r45 3 15 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.025 $Y=0.765
+ $X2=1.025 $Y2=1.295
.ends

.subckt PM_SKY130_FD_SC_LP__A22OI_1%A1 3 6 8 9 10 11 18 20 28 36
c48 28 0 5.1293e-20 $X=1.682 $Y=1.342
c49 10 0 1.18028e-19 $X=1.595 $Y=1.21
r50 28 36 1.83781 $w=3.25e-07 $l=4.7e-08 $layer=LI1_cond $X=1.682 $Y=1.342
+ $X2=1.682 $Y2=1.295
r51 18 21 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.67 $Y=1.46
+ $X2=1.67 $Y2=1.625
r52 18 20 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.67 $Y=1.46
+ $X2=1.67 $Y2=1.295
r53 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.67
+ $Y=1.46 $X2=1.67 $Y2=1.46
r54 11 19 7.26926 $w=3.23e-07 $l=2.05e-07 $layer=LI1_cond $X=1.682 $Y=1.665
+ $X2=1.682 $Y2=1.46
r55 10 36 0.765016 $w=3.03e-07 $l=1.9e-08 $layer=LI1_cond $X=1.682 $Y=1.276
+ $X2=1.682 $Y2=1.295
r56 10 22 7.92059 $w=3.03e-07 $l=1.83347e-07 $layer=LI1_cond $X=1.682 $Y=1.276
+ $X2=1.697 $Y2=1.1
r57 10 19 3.51052 $w=3.23e-07 $l=9.9e-08 $layer=LI1_cond $X=1.682 $Y=1.361
+ $X2=1.682 $Y2=1.46
r58 10 28 0.673736 $w=3.23e-07 $l=1.9e-08 $layer=LI1_cond $X=1.682 $Y=1.361
+ $X2=1.682 $Y2=1.342
r59 9 22 8.96345 $w=2.23e-07 $l=1.75e-07 $layer=LI1_cond $X=1.697 $Y=0.925
+ $X2=1.697 $Y2=1.1
r60 8 9 18.9513 $w=2.23e-07 $l=3.7e-07 $layer=LI1_cond $X=1.697 $Y=0.555
+ $X2=1.697 $Y2=0.925
r61 6 21 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=1.58 $Y=2.465
+ $X2=1.58 $Y2=1.625
r62 3 20 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.58 $Y=0.765
+ $X2=1.58 $Y2=1.295
.ends

.subckt PM_SKY130_FD_SC_LP__A22OI_1%A2 1 3 6 8 10 20
r35 20 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.55
+ $Y=1.46 $X2=2.55 $Y2=1.46
r36 18 20 34.9723 $w=3.3e-07 $l=2e-07 $layer=POLY_cond $X=2.35 $Y=1.46 $X2=2.55
+ $Y2=1.46
r37 16 18 40.2181 $w=3.3e-07 $l=2.3e-07 $layer=POLY_cond $X=2.12 $Y=1.46
+ $X2=2.35 $Y2=1.46
r38 10 21 1.99346 $w=5.38e-07 $l=9e-08 $layer=LI1_cond $X=2.64 $Y=1.48 $X2=2.55
+ $Y2=1.48
r39 8 21 8.63834 $w=5.38e-07 $l=3.9e-07 $layer=LI1_cond $X=2.16 $Y=1.48 $X2=2.55
+ $Y2=1.48
r40 4 18 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.35 $Y=1.625
+ $X2=2.35 $Y2=1.46
r41 4 6 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=2.35 $Y=1.625 $X2=2.35
+ $Y2=2.465
r42 1 16 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.12 $Y=1.295
+ $X2=2.12 $Y2=1.46
r43 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.12 $Y=1.295 $X2=2.12
+ $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_LP__A22OI_1%A_65_367# 1 2 3 10 12 14 16 18 22 26 32
r35 24 32 3.27229 $w=2.87e-07 $l=9.80051e-08 $layer=LI1_cond $X=2.6 $Y=2.47
+ $X2=2.572 $Y2=2.385
r36 24 26 1.55137 $w=2.58e-07 $l=3.5e-08 $layer=LI1_cond $X=2.6 $Y=2.47 $X2=2.6
+ $Y2=2.505
r37 20 32 3.27229 $w=2.87e-07 $l=8.5e-08 $layer=LI1_cond $X=2.572 $Y=2.3
+ $X2=2.572 $Y2=2.385
r38 20 22 7.50003 $w=3.13e-07 $l=2.05e-07 $layer=LI1_cond $X=2.572 $Y=2.3
+ $X2=2.572 $Y2=2.095
r39 19 31 4.20453 $w=1.7e-07 $l=1.23e-07 $layer=LI1_cond $X=1.46 $Y=2.385
+ $X2=1.337 $Y2=2.385
r40 18 32 3.2872 $w=1.7e-07 $l=1.57e-07 $layer=LI1_cond $X=2.415 $Y=2.385
+ $X2=2.572 $Y2=2.385
r41 18 19 62.3048 $w=1.68e-07 $l=9.55e-07 $layer=LI1_cond $X=2.415 $Y=2.385
+ $X2=1.46 $Y2=2.385
r42 16 31 2.90557 $w=2.45e-07 $l=8.5e-08 $layer=LI1_cond $X=1.337 $Y=2.47
+ $X2=1.337 $Y2=2.385
r43 16 17 20.4617 $w=2.43e-07 $l=4.35e-07 $layer=LI1_cond $X=1.337 $Y=2.47
+ $X2=1.337 $Y2=2.905
r44 15 29 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.535 $Y=2.99
+ $X2=0.41 $Y2=2.99
r45 14 17 7.11011 $w=1.7e-07 $l=1.58915e-07 $layer=LI1_cond $X=1.215 $Y=2.99
+ $X2=1.337 $Y2=2.905
r46 14 15 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.215 $Y=2.99
+ $X2=0.535 $Y2=2.99
r47 10 29 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.41 $Y=2.905
+ $X2=0.41 $Y2=2.99
r48 10 12 37.8001 $w=2.48e-07 $l=8.2e-07 $layer=LI1_cond $X=0.41 $Y=2.905
+ $X2=0.41 $Y2=2.085
r49 3 26 300 $w=1.7e-07 $l=7.36682e-07 $layer=licon1_PDIFF $count=2 $X=2.425
+ $Y=1.835 $X2=2.565 $Y2=2.505
r50 3 22 600 $w=1.7e-07 $l=3.2249e-07 $layer=licon1_PDIFF $count=1 $X=2.425
+ $Y=1.835 $X2=2.565 $Y2=2.095
r51 2 31 300 $w=1.7e-07 $l=7.0993e-07 $layer=licon1_PDIFF $count=2 $X=1.17
+ $Y=1.835 $X2=1.34 $Y2=2.465
r52 1 29 400 $w=1.7e-07 $l=1.13578e-06 $layer=licon1_PDIFF $count=1 $X=0.325
+ $Y=1.835 $X2=0.45 $Y2=2.91
r53 1 12 400 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_PDIFF $count=1 $X=0.325
+ $Y=1.835 $X2=0.45 $Y2=2.085
.ends

.subckt PM_SKY130_FD_SC_LP__A22OI_1%Y 1 2 8 11 12 15 19 20 21 22
r46 21 22 25.3506 $w=2.08e-07 $l=4.8e-07 $layer=LI1_cond $X=1.68 $Y=2.025
+ $X2=2.16 $Y2=2.025
r47 20 21 25.3506 $w=2.08e-07 $l=4.8e-07 $layer=LI1_cond $X=1.2 $Y=2.025
+ $X2=1.68 $Y2=2.025
r48 17 20 8.18615 $w=2.08e-07 $l=1.55e-07 $layer=LI1_cond $X=1.045 $Y=2.025
+ $X2=1.2 $Y2=2.025
r49 17 19 2.05017 $w=2.1e-07 $l=1.7e-07 $layer=LI1_cond $X=1.045 $Y=2.025
+ $X2=0.875 $Y2=2.025
r50 13 15 19.5411 $w=2.08e-07 $l=3.7e-07 $layer=LI1_cond $X=1.31 $Y=0.86
+ $X2=1.31 $Y2=0.49
r51 11 13 6.86909 $w=1.8e-07 $l=1.43091e-07 $layer=LI1_cond $X=1.205 $Y=0.95
+ $X2=1.31 $Y2=0.86
r52 11 12 20.3333 $w=1.78e-07 $l=3.3e-07 $layer=LI1_cond $X=1.205 $Y=0.95
+ $X2=0.875 $Y2=0.95
r53 8 19 4.38255 $w=2.55e-07 $l=1.41244e-07 $layer=LI1_cond $X=0.79 $Y=1.92
+ $X2=0.875 $Y2=2.025
r54 7 12 6.82373 $w=1.8e-07 $l=1.25499e-07 $layer=LI1_cond $X=0.79 $Y=1.04
+ $X2=0.875 $Y2=0.95
r55 7 8 57.4118 $w=1.68e-07 $l=8.8e-07 $layer=LI1_cond $X=0.79 $Y=1.04 $X2=0.79
+ $Y2=1.92
r56 2 19 300 $w=1.7e-07 $l=2.60768e-07 $layer=licon1_PDIFF $count=2 $X=0.74
+ $Y=1.835 $X2=0.88 $Y2=2.035
r57 1 15 91 $w=1.7e-07 $l=2.93684e-07 $layer=licon1_NDIFF $count=2 $X=1.1
+ $Y=0.345 $X2=1.33 $Y2=0.49
.ends

.subckt PM_SKY130_FD_SC_LP__A22OI_1%VPWR 1 4 6 13 14 17
r31 21 23 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r32 20 23 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r33 20 21 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r34 17 20 10.0863 $w=6.68e-07 $l=5.65e-07 $layer=LI1_cond $X=1.965 $Y=2.765
+ $X2=1.965 $Y2=3.33
r35 14 23 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r36 13 14 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r37 11 20 9.03384 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=2.3 $Y=3.33
+ $X2=1.965 $Y2=3.33
r38 11 13 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=2.3 $Y=3.33 $X2=2.64
+ $Y2=3.33
r39 8 9 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.24 $Y=3.33 $X2=0.24
+ $Y2=3.33
r40 6 20 9.03384 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=1.63 $Y=3.33
+ $X2=1.965 $Y2=3.33
r41 6 8 90.6845 $w=1.68e-07 $l=1.39e-06 $layer=LI1_cond $X=1.63 $Y=3.33 $X2=0.24
+ $Y2=3.33
r42 4 21 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=1.68 $Y2=3.33
r43 4 9 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=1.44 $Y=3.33 $X2=0.24
+ $Y2=3.33
r44 1 17 300 $w=1.7e-07 $l=1.14512e-06 $layer=licon1_PDIFF $count=2 $X=1.655
+ $Y=1.835 $X2=2.135 $Y2=2.765
.ends

.subckt PM_SKY130_FD_SC_LP__A22OI_1%VGND 1 2 9 13 16 17 19 20 21 33 34
r31 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r32 31 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r33 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r34 27 30 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=0.72 $Y=0 $X2=2.16
+ $Y2=0
r35 27 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r36 25 28 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r37 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r38 21 31 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=2.16
+ $Y2=0
r39 21 28 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=0.72
+ $Y2=0
r40 19 30 0.652406 $w=1.68e-07 $l=1e-08 $layer=LI1_cond $X=2.17 $Y=0 $X2=2.16
+ $Y2=0
r41 19 20 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.17 $Y=0 $X2=2.335
+ $Y2=0
r42 18 33 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=2.5 $Y=0 $X2=2.64
+ $Y2=0
r43 18 20 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.5 $Y=0 $X2=2.335
+ $Y2=0
r44 16 24 3.22941 $w=1.7e-07 $l=4.5e-08 $layer=LI1_cond $X=0.285 $Y=0 $X2=0.24
+ $Y2=0
r45 16 17 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.285 $Y=0 $X2=0.41
+ $Y2=0
r46 15 27 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=0.535 $Y=0 $X2=0.72
+ $Y2=0
r47 15 17 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.535 $Y=0 $X2=0.41
+ $Y2=0
r48 11 20 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.335 $Y=0.085
+ $X2=2.335 $Y2=0
r49 11 13 14.1436 $w=3.28e-07 $l=4.05e-07 $layer=LI1_cond $X=2.335 $Y=0.085
+ $X2=2.335 $Y2=0.49
r50 7 17 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.41 $Y=0.085
+ $X2=0.41 $Y2=0
r51 7 9 18.6696 $w=2.48e-07 $l=4.05e-07 $layer=LI1_cond $X=0.41 $Y=0.085
+ $X2=0.41 $Y2=0.49
r52 2 13 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.195
+ $Y=0.345 $X2=2.335 $Y2=0.49
r53 1 9 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.325
+ $Y=0.345 $X2=0.45 $Y2=0.49
.ends

