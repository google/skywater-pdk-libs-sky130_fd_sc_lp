# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__nand3b_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_lp__nand3b_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.200000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A_N
    ANTENNAGATEAREA  0.315000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.600000 1.210000 0.805000 1.750000 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.385000 1.405000 4.735000 1.760000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.950000 1.405000 7.045000 1.760000 ;
    END
  END C
  PIN Y
    ANTENNADIFFAREA  2.587200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.355000 1.690000 3.205000 1.930000 ;
        RECT 1.355000 1.930000 6.190000 1.945000 ;
        RECT 1.355000 1.945000 1.595000 3.075000 ;
        RECT 1.515000 0.595000 1.775000 0.975000 ;
        RECT 1.515000 0.975000 3.090000 1.145000 ;
        RECT 2.265000 1.945000 6.190000 2.100000 ;
        RECT 2.265000 2.100000 3.380000 2.490000 ;
        RECT 2.265000 2.490000 2.455000 3.075000 ;
        RECT 2.445000 0.595000 2.635000 0.975000 ;
        RECT 2.920000 1.145000 3.090000 1.210000 ;
        RECT 2.920000 1.210000 3.205000 1.690000 ;
        RECT 3.145000 2.490000 3.380000 3.075000 ;
        RECT 4.050000 2.100000 4.365000 3.075000 ;
        RECT 5.035000 2.100000 5.330000 3.075000 ;
        RECT 6.000000 2.100000 6.190000 3.075000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 7.200000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 7.200000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.200000 0.085000 ;
      RECT 0.000000  3.245000 7.200000 3.415000 ;
      RECT 0.135000  0.360000 0.395000 0.870000 ;
      RECT 0.135000  0.870000 1.320000 1.040000 ;
      RECT 0.135000  1.040000 0.405000 1.920000 ;
      RECT 0.135000  1.920000 0.740000 3.075000 ;
      RECT 0.565000  0.085000 0.895000 0.700000 ;
      RECT 0.910000  1.885000 1.185000 3.245000 ;
      RECT 0.975000  1.040000 1.320000 1.315000 ;
      RECT 0.975000  1.315000 2.750000 1.520000 ;
      RECT 1.085000  0.255000 4.855000 0.425000 ;
      RECT 1.085000  0.425000 1.345000 0.700000 ;
      RECT 1.765000  2.115000 2.095000 3.245000 ;
      RECT 1.945000  0.425000 2.275000 0.805000 ;
      RECT 2.625000  2.660000 2.955000 3.245000 ;
      RECT 2.805000  0.425000 4.855000 0.445000 ;
      RECT 2.805000  0.445000 3.135000 0.805000 ;
      RECT 3.305000  0.615000 3.495000 0.955000 ;
      RECT 3.305000  0.955000 4.355000 1.065000 ;
      RECT 3.330000  1.065000 6.630000 1.085000 ;
      RECT 3.375000  1.085000 6.630000 1.235000 ;
      RECT 3.550000  2.270000 3.880000 3.245000 ;
      RECT 3.665000  0.445000 3.995000 0.785000 ;
      RECT 4.165000  0.615000 4.355000 0.955000 ;
      RECT 4.525000  0.445000 4.855000 0.895000 ;
      RECT 4.535000  2.270000 4.865000 3.245000 ;
      RECT 5.045000  0.085000 5.375000 0.885000 ;
      RECT 5.500000  2.270000 5.830000 3.245000 ;
      RECT 5.545000  0.255000 5.735000 1.065000 ;
      RECT 5.905000  0.085000 6.235000 0.895000 ;
      RECT 6.360000  1.930000 6.690000 3.245000 ;
      RECT 6.405000  0.255000 6.630000 1.065000 ;
      RECT 6.800000  0.085000 7.095000 1.095000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
  END
END sky130_fd_sc_lp__nand3b_4
END LIBRARY
