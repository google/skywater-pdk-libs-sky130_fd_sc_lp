* NGSPICE file created from sky130_fd_sc_lp__busdrivernovlp2_20.ext - technology: sky130A

.subckt sky130_fd_sc_lp__busdrivernovlp2_20 A TE_B VGND VNB VPB VPWR Z
M1000 a_1238_47# a_726_47# a_1260_373# VPB pshort w=840000u l=150000u
+  ad=2.394e+11p pd=2.25e+06u as=2.016e+11p ps=2.16e+06u
M1001 a_726_47# A VGND VNB nshort w=840000u l=150000u
+  ad=6.774e+11p pd=5.18e+06u as=3.1757e+12p ps=2.682e+07u
M1002 VGND A a_1451_47# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=8.022e+11p ps=6.95e+06u
M1003 a_1451_47# A VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VPWR a_217_367# Z VPB pshort w=1.26e+06u l=150000u
+  ad=6.6423e+12p pd=5.222e+07u as=3.528e+12p ps=3.08e+07u
M1005 VGND a_726_47# Z VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=1.44e+12p ps=1.474e+07u
M1006 VGND a_726_47# Z VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_658_367# a_381_85# a_726_47# VPB pshort w=1.26e+06u l=150000u
+  ad=1.4049e+12p pd=9.79e+06u as=3.528e+11p ps=3.08e+06u
M1008 VPWR a_217_367# Z VPB pshort w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR a_217_367# Z VPB pshort w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND A a_726_47# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND a_726_47# a_1238_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.47e+11p ps=1.54e+06u
M1012 Z a_217_367# VPWR VPB pshort w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VGND a_726_47# Z VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 Z a_217_367# VPWR VPB pshort w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_217_367# a_27_367# VPWR VPB pshort w=1.26e+06u l=150000u
+  ad=7.056e+11p pd=6.16e+06u as=0p ps=0u
M1016 VPWR a_217_367# Z VPB pshort w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VPWR a_217_367# Z VPB pshort w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_1238_47# TE_B VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VPWR a_27_367# a_217_367# VPB pshort w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_217_367# a_1238_47# a_1451_47# VNB nshort w=840000u l=150000u
+  ad=3.024e+11p pd=2.4e+06u as=0p ps=0u
M1021 Z a_726_47# VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 Z a_217_367# VPWR VPB pshort w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_726_47# a_381_85# a_658_367# VPB pshort w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_726_47# TE_B VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 Z a_217_367# VPWR VPB pshort w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 VPWR a_217_367# Z VPB pshort w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 Z a_217_367# VPWR VPB pshort w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_217_367# A VPWR VPB pshort w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 VGND a_726_47# Z VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 VPWR A a_658_367# VPB pshort w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 VPWR A a_217_367# VPB pshort w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 Z a_217_367# VPWR VPB pshort w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 VPWR a_217_367# Z VPB pshort w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1034 VGND a_726_47# Z VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1035 a_381_85# a_27_367# VPWR VPB pshort w=840000u l=150000u
+  ad=2.352e+11p pd=2.24e+06u as=0p ps=0u
M1036 VPWR a_217_367# Z VPB pshort w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1037 VPWR a_217_367# Z VPB pshort w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1038 VPWR a_217_367# a_381_85# VPB pshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1039 a_1451_47# a_1238_47# a_217_367# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1040 Z a_726_47# VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1041 VGND TE_B a_27_367# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1042 Z a_217_367# VPWR VPB pshort w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1043 Z a_726_47# VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1044 a_1260_373# TE_B VPWR VPB pshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1045 a_658_367# A VPWR VPB pshort w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1046 Z a_726_47# VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1047 VGND a_726_47# Z VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1048 Z a_217_367# VPWR VPB pshort w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1049 VGND TE_B a_726_47# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1050 Z a_217_367# VPWR VPB pshort w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1051 Z a_217_367# VPWR VPB pshort w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1052 VPWR TE_B a_27_367# VPB pshort w=840000u l=150000u
+  ad=0p pd=0u as=2.268e+11p ps=2.22e+06u
M1053 VPWR a_217_367# Z VPB pshort w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1054 Z a_726_47# VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1055 a_381_85# a_217_367# a_303_85# VNB nshort w=420000u l=150000u
+  ad=1.912e+11p pd=1.8e+06u as=1.008e+11p ps=1.32e+06u
M1056 Z a_726_47# VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1057 a_303_85# a_27_367# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1058 VGND a_726_47# Z VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1059 Z a_726_47# VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

