* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__srdlrtp_1 D GATE RESET_B SLEEP_B KAPWR VGND VNB VPB VPWR
+ Q
X0 a_570_97# a_612_71# a_642_97# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 VPWR a_2120_55# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X2 a_336_71# a_393_335# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X3 a_366_97# a_336_71# a_438_97# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 a_642_97# a_612_71# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 VPWR D a_27_97# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X6 KAPWR a_1324_394# a_1765_419# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X7 a_2120_55# a_438_97# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X8 VGND a_27_97# a_280_97# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 a_1624_47# a_438_97# a_1917_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 VGND a_393_335# a_336_71# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X11 a_27_97# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X12 a_1565_419# a_612_71# KAPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X13 a_438_97# a_393_335# a_570_97# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X14 a_280_97# a_393_335# a_423_487# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X15 a_423_487# a_393_335# a_438_97# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X16 VGND a_2120_55# Q VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X17 a_280_97# a_336_71# a_366_97# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X18 a_1069_97# SLEEP_B a_1147_97# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X19 a_393_335# SLEEP_B KAPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X20 a_1147_97# SLEEP_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X21 a_1624_47# a_1324_394# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X22 a_2120_55# a_438_97# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X23 VPWR a_27_97# a_280_97# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X24 a_438_97# a_336_71# a_1565_419# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X25 a_1765_419# RESET_B a_612_71# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X26 KAPWR SLEEP_B a_1324_394# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X27 a_114_97# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X28 VGND SLEEP_B a_1344_97# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X29 VGND RESET_B a_1624_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X30 a_27_97# D a_114_97# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X31 a_1344_97# SLEEP_B a_1324_394# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X32 a_1917_47# a_438_97# a_612_71# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X33 a_612_71# a_438_97# KAPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X34 a_393_335# GATE a_1069_97# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X35 KAPWR GATE a_393_335# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
.ends
