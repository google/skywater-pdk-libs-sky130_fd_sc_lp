* NGSPICE file created from sky130_fd_sc_lp__a2bb2o_1.ext - technology: sky130A

.subckt sky130_fd_sc_lp__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
M1000 a_271_367# A1_N VPWR VPB phighvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=5.271e+11p ps=4.81e+06u
M1001 a_505_529# B1 VPWR VPB phighvt w=420000u l=150000u
+  ad=2.289e+11p pd=2.77e+06u as=0p ps=0u
M1002 a_571_47# B2 a_91_269# VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=1.176e+11p ps=1.4e+06u
M1003 VGND B1 a_571_47# VNB nshort w=420000u l=150000u
+  ad=6.762e+11p pd=6.05e+06u as=0p ps=0u
M1004 VPWR B2 a_505_529# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_271_47# A1_N VGND VNB nshort w=420000u l=150000u
+  ad=1.407e+11p pd=1.51e+06u as=0p ps=0u
M1006 VGND A2_N a_271_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_271_47# A2_N a_271_367# VPB phighvt w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1008 a_91_269# a_271_47# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR a_91_269# X VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=3.339e+11p ps=3.05e+06u
M1010 a_505_529# a_271_47# a_91_269# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1011 VGND a_91_269# X VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=2.226e+11p ps=2.21e+06u
.ends

