* File: sky130_fd_sc_lp__a2111o_4.pxi.spice
* Created: Fri Aug 28 09:46:04 2020
* 
x_PM_SKY130_FD_SC_LP__A2111O_4%D1 N_D1_M1006_g N_D1_M1004_g N_D1_c_144_n
+ N_D1_M1018_g N_D1_M1022_g N_D1_c_147_n N_D1_c_148_n N_D1_c_149_n D1
+ N_D1_c_150_n PM_SKY130_FD_SC_LP__A2111O_4%D1
x_PM_SKY130_FD_SC_LP__A2111O_4%C1 N_C1_M1000_g N_C1_M1002_g N_C1_M1013_g
+ N_C1_M1012_g C1 C1 C1 C1 N_C1_c_193_n PM_SKY130_FD_SC_LP__A2111O_4%C1
x_PM_SKY130_FD_SC_LP__A2111O_4%B1 N_B1_M1005_g N_B1_c_247_n N_B1_M1009_g
+ N_B1_M1025_g N_B1_M1014_g B1 B1 N_B1_c_250_n N_B1_c_251_n N_B1_c_262_n
+ PM_SKY130_FD_SC_LP__A2111O_4%B1
x_PM_SKY130_FD_SC_LP__A2111O_4%A1 N_A1_c_313_n N_A1_M1003_g N_A1_M1015_g
+ N_A1_c_315_n N_A1_c_316_n N_A1_M1016_g N_A1_M1023_g N_A1_c_318_n N_A1_c_319_n
+ A1 N_A1_c_321_n PM_SKY130_FD_SC_LP__A2111O_4%A1
x_PM_SKY130_FD_SC_LP__A2111O_4%A2 N_A2_c_374_n N_A2_M1010_g N_A2_M1001_g
+ N_A2_c_376_n N_A2_M1021_g N_A2_M1020_g A2 N_A2_c_381_n N_A2_c_378_n
+ PM_SKY130_FD_SC_LP__A2111O_4%A2
x_PM_SKY130_FD_SC_LP__A2111O_4%A_77_47# N_A_77_47#_M1004_s N_A_77_47#_M1022_s
+ N_A_77_47#_M1012_s N_A_77_47#_M1014_d N_A_77_47#_M1016_d N_A_77_47#_M1006_s
+ N_A_77_47#_M1007_g N_A_77_47#_M1011_g N_A_77_47#_M1008_g N_A_77_47#_M1017_g
+ N_A_77_47#_M1019_g N_A_77_47#_M1024_g N_A_77_47#_M1027_g N_A_77_47#_M1026_g
+ N_A_77_47#_c_425_n N_A_77_47#_c_426_n N_A_77_47#_c_427_n N_A_77_47#_c_570_p
+ N_A_77_47#_c_428_n N_A_77_47#_c_591_p N_A_77_47#_c_429_n N_A_77_47#_c_585_p
+ N_A_77_47#_c_430_n N_A_77_47#_c_431_n N_A_77_47#_c_432_n N_A_77_47#_c_433_n
+ N_A_77_47#_c_446_n N_A_77_47#_c_523_p N_A_77_47#_c_455_n N_A_77_47#_c_434_n
+ N_A_77_47#_c_435_n N_A_77_47#_c_436_n N_A_77_47#_c_437_n N_A_77_47#_c_438_n
+ N_A_77_47#_c_439_n PM_SKY130_FD_SC_LP__A2111O_4%A_77_47#
x_PM_SKY130_FD_SC_LP__A2111O_4%A_63_367# N_A_63_367#_M1006_d N_A_63_367#_M1018_d
+ N_A_63_367#_M1013_d N_A_63_367#_c_614_n N_A_63_367#_c_615_n
+ N_A_63_367#_c_620_n N_A_63_367#_c_622_n N_A_63_367#_c_616_n
+ N_A_63_367#_c_617_n N_A_63_367#_c_638_p PM_SKY130_FD_SC_LP__A2111O_4%A_63_367#
x_PM_SKY130_FD_SC_LP__A2111O_4%A_318_367# N_A_318_367#_M1000_s
+ N_A_318_367#_M1009_d N_A_318_367#_c_646_n N_A_318_367#_c_670_p
+ N_A_318_367#_c_651_n N_A_318_367#_c_647_n
+ PM_SKY130_FD_SC_LP__A2111O_4%A_318_367#
x_PM_SKY130_FD_SC_LP__A2111O_4%A_511_349# N_A_511_349#_M1009_s
+ N_A_511_349#_M1025_s N_A_511_349#_M1023_d N_A_511_349#_M1001_d
+ N_A_511_349#_c_672_n N_A_511_349#_c_673_n N_A_511_349#_c_674_n
+ N_A_511_349#_c_685_n N_A_511_349#_c_688_n N_A_511_349#_c_689_n
+ N_A_511_349#_c_675_n N_A_511_349#_c_676_n N_A_511_349#_c_719_p
+ N_A_511_349#_c_677_n PM_SKY130_FD_SC_LP__A2111O_4%A_511_349#
x_PM_SKY130_FD_SC_LP__A2111O_4%VPWR N_VPWR_M1015_s N_VPWR_M1001_s N_VPWR_M1020_s
+ N_VPWR_M1017_s N_VPWR_M1026_s N_VPWR_c_726_n N_VPWR_c_727_n N_VPWR_c_728_n
+ N_VPWR_c_729_n N_VPWR_c_730_n N_VPWR_c_731_n N_VPWR_c_732_n VPWR
+ N_VPWR_c_733_n N_VPWR_c_734_n N_VPWR_c_735_n N_VPWR_c_736_n N_VPWR_c_737_n
+ N_VPWR_c_738_n N_VPWR_c_739_n N_VPWR_c_740_n N_VPWR_c_725_n
+ PM_SKY130_FD_SC_LP__A2111O_4%VPWR
x_PM_SKY130_FD_SC_LP__A2111O_4%X N_X_M1007_s N_X_M1019_s N_X_M1011_d N_X_M1024_d
+ N_X_c_888_p N_X_c_872_n N_X_c_832_n N_X_c_833_n N_X_c_838_n N_X_c_839_n
+ N_X_c_889_p N_X_c_876_n N_X_c_834_n N_X_c_840_n N_X_c_835_n N_X_c_841_n X X
+ N_X_c_836_n N_X_c_842_n X X PM_SKY130_FD_SC_LP__A2111O_4%X
x_PM_SKY130_FD_SC_LP__A2111O_4%VGND N_VGND_M1004_d N_VGND_M1002_d N_VGND_M1005_s
+ N_VGND_M1010_s N_VGND_M1021_s N_VGND_M1008_d N_VGND_M1027_d N_VGND_c_894_n
+ N_VGND_c_895_n N_VGND_c_896_n N_VGND_c_897_n N_VGND_c_898_n N_VGND_c_899_n
+ N_VGND_c_900_n N_VGND_c_901_n N_VGND_c_902_n N_VGND_c_903_n VGND
+ N_VGND_c_904_n N_VGND_c_905_n N_VGND_c_906_n N_VGND_c_907_n N_VGND_c_908_n
+ N_VGND_c_909_n N_VGND_c_910_n N_VGND_c_911_n N_VGND_c_912_n N_VGND_c_913_n
+ N_VGND_c_914_n PM_SKY130_FD_SC_LP__A2111O_4%VGND
x_PM_SKY130_FD_SC_LP__A2111O_4%A_813_47# N_A_813_47#_M1003_s N_A_813_47#_M1010_d
+ N_A_813_47#_c_1014_n N_A_813_47#_c_1024_n N_A_813_47#_c_1041_n
+ N_A_813_47#_c_1016_n N_A_813_47#_c_1015_n
+ PM_SKY130_FD_SC_LP__A2111O_4%A_813_47#
cc_1 VNB N_D1_M1004_g 0.0306293f $X=-0.19 $Y=-0.245 $X2=0.725 $Y2=0.655
cc_2 VNB N_D1_c_144_n 0.0116648f $X=-0.19 $Y=-0.245 $X2=1.01 $Y2=1.42
cc_3 VNB N_D1_M1018_g 0.00692255f $X=-0.19 $Y=-0.245 $X2=1.085 $Y2=2.465
cc_4 VNB N_D1_M1022_g 0.0229769f $X=-0.19 $Y=-0.245 $X2=1.155 $Y2=0.655
cc_5 VNB N_D1_c_147_n 0.0359041f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=1.51
cc_6 VNB N_D1_c_148_n 0.0106252f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=1.51
cc_7 VNB N_D1_c_149_n 0.00758588f $X=-0.19 $Y=-0.245 $X2=1.12 $Y2=1.42
cc_8 VNB N_D1_c_150_n 0.0133334f $X=-0.19 $Y=-0.245 $X2=0.37 $Y2=1.51
cc_9 VNB N_C1_M1002_g 0.0252029f $X=-0.19 $Y=-0.245 $X2=0.725 $Y2=0.655
cc_10 VNB N_C1_M1012_g 0.0252278f $X=-0.19 $Y=-0.245 $X2=1.155 $Y2=1.345
cc_11 VNB C1 0.0106955f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=1.51
cc_12 VNB N_C1_c_193_n 0.041915f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_B1_M1005_g 0.0252601f $X=-0.19 $Y=-0.245 $X2=0.655 $Y2=2.465
cc_14 VNB N_B1_c_247_n 0.00912187f $X=-0.19 $Y=-0.245 $X2=0.725 $Y2=0.655
cc_15 VNB N_B1_M1014_g 0.0252601f $X=-0.19 $Y=-0.245 $X2=1.155 $Y2=0.655
cc_16 VNB B1 0.00435131f $X=-0.19 $Y=-0.245 $X2=0.37 $Y2=1.51
cc_17 VNB N_B1_c_250_n 0.0113791f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_B1_c_251_n 0.0536335f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A1_c_313_n 0.0155902f $X=-0.19 $Y=-0.245 $X2=0.655 $Y2=1.675
cc_20 VNB N_A1_M1015_g 0.00902388f $X=-0.19 $Y=-0.245 $X2=0.725 $Y2=0.655
cc_21 VNB N_A1_c_315_n 0.00950625f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A1_c_316_n 0.0196497f $X=-0.19 $Y=-0.245 $X2=0.8 $Y2=1.42
cc_23 VNB N_A1_M1023_g 0.00302787f $X=-0.19 $Y=-0.245 $X2=1.155 $Y2=1.345
cc_24 VNB N_A1_c_318_n 0.00515988f $X=-0.19 $Y=-0.245 $X2=1.155 $Y2=0.655
cc_25 VNB N_A1_c_319_n 0.0083384f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=1.51
cc_26 VNB A1 0.00409524f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=1.51
cc_27 VNB N_A1_c_321_n 0.0497705f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A2_c_374_n 0.0212151f $X=-0.19 $Y=-0.245 $X2=0.655 $Y2=1.675
cc_29 VNB N_A2_M1001_g 0.0103004f $X=-0.19 $Y=-0.245 $X2=0.725 $Y2=0.655
cc_30 VNB N_A2_c_376_n 0.0161955f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A2_M1020_g 0.00688395f $X=-0.19 $Y=-0.245 $X2=1.085 $Y2=2.465
cc_32 VNB N_A2_c_378_n 0.0384348f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_33 VNB N_A_77_47#_M1007_g 0.0234946f $X=-0.19 $Y=-0.245 $X2=1.12 $Y2=1.42
cc_34 VNB N_A_77_47#_M1008_g 0.0217542f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_77_47#_M1019_g 0.0217335f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_77_47#_M1027_g 0.0264939f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_77_47#_c_425_n 0.0308502f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_77_47#_c_426_n 0.00401221f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_77_47#_c_427_n 0.0102628f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_77_47#_c_428_n 0.00323641f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_77_47#_c_429_n 0.00893822f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_77_47#_c_430_n 0.00219402f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_77_47#_c_431_n 0.00840189f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_77_47#_c_432_n 0.00271393f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_77_47#_c_433_n 0.00858526f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_77_47#_c_434_n 0.00239411f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_77_47#_c_435_n 0.002926f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_77_47#_c_436_n 0.0025736f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_77_47#_c_437_n 0.00173208f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_77_47#_c_438_n 0.00410226f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_77_47#_c_439_n 0.0706322f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_VPWR_c_725_n 0.342803f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_X_c_832_n 0.00304538f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_X_c_833_n 0.00336604f $X=-0.19 $Y=-0.245 $X2=0.37 $Y2=1.51
cc_55 VNB N_X_c_834_n 0.00141236f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_X_c_835_n 0.00144145f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_X_c_836_n 0.0144315f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB X 0.0238099f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_894_n 4.06069e-19 $X=-0.19 $Y=-0.245 $X2=0.37 $Y2=1.51
cc_60 VNB N_VGND_c_895_n 0.0148832f $X=-0.19 $Y=-0.245 $X2=0.37 $Y2=1.51
cc_61 VNB N_VGND_c_896_n 0.00431919f $X=-0.19 $Y=-0.245 $X2=0.31 $Y2=1.665
cc_62 VNB N_VGND_c_897_n 0.0069711f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_VGND_c_898_n 3.0911e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_VGND_c_899_n 3.0911e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_VGND_c_900_n 0.014353f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_VGND_c_901_n 0.0284267f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_902_n 0.0233314f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_VGND_c_903_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_VGND_c_904_n 0.0356045f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_VGND_c_905_n 0.012342f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_VGND_c_906_n 0.0129398f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_VGND_c_907_n 0.0129398f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_VGND_c_908_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_VGND_c_909_n 0.0148773f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_VGND_c_910_n 0.0188651f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_VGND_c_911_n 0.00510817f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_VGND_c_912_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_VGND_c_913_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_VGND_c_914_n 0.406298f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_A_813_47#_c_1014_n 0.00579851f $X=-0.19 $Y=-0.245 $X2=1.085
+ $Y2=1.495
cc_81 VNB N_A_813_47#_c_1015_n 0.00393963f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VPB N_D1_M1006_g 0.0235111f $X=-0.19 $Y=1.655 $X2=0.655 $Y2=2.465
cc_83 VPB N_D1_M1018_g 0.0193998f $X=-0.19 $Y=1.655 $X2=1.085 $Y2=2.465
cc_84 VPB N_D1_c_147_n 0.0130672f $X=-0.19 $Y=1.655 $X2=0.58 $Y2=1.51
cc_85 VPB N_D1_c_148_n 0.00266576f $X=-0.19 $Y=1.655 $X2=0.69 $Y2=1.51
cc_86 VPB N_D1_c_150_n 0.013579f $X=-0.19 $Y=1.655 $X2=0.37 $Y2=1.51
cc_87 VPB N_C1_M1000_g 0.0181399f $X=-0.19 $Y=1.655 $X2=0.655 $Y2=2.465
cc_88 VPB N_C1_M1013_g 0.0240007f $X=-0.19 $Y=1.655 $X2=1.085 $Y2=1.495
cc_89 VPB C1 0.0172841f $X=-0.19 $Y=1.655 $X2=0.69 $Y2=1.51
cc_90 VPB N_C1_c_193_n 0.0094119f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_91 VPB N_B1_M1009_g 0.022194f $X=-0.19 $Y=1.655 $X2=1.01 $Y2=1.42
cc_92 VPB N_B1_M1025_g 0.0202196f $X=-0.19 $Y=1.655 $X2=1.085 $Y2=2.465
cc_93 VPB B1 0.00112826f $X=-0.19 $Y=1.655 $X2=0.37 $Y2=1.51
cc_94 VPB N_B1_c_251_n 0.0137429f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_95 VPB N_A1_M1015_g 0.0205609f $X=-0.19 $Y=1.655 $X2=0.725 $Y2=0.655
cc_96 VPB N_A1_M1023_g 0.0230909f $X=-0.19 $Y=1.655 $X2=1.155 $Y2=1.345
cc_97 VPB N_A2_M1001_g 0.0240097f $X=-0.19 $Y=1.655 $X2=0.725 $Y2=0.655
cc_98 VPB N_A2_M1020_g 0.0186413f $X=-0.19 $Y=1.655 $X2=1.085 $Y2=2.465
cc_99 VPB N_A_77_47#_M1011_g 0.0190885f $X=-0.19 $Y=1.655 $X2=0.37 $Y2=1.51
cc_100 VPB N_A_77_47#_M1017_g 0.0187605f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_101 VPB N_A_77_47#_M1024_g 0.0187589f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_102 VPB N_A_77_47#_M1026_g 0.0224447f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_103 VPB N_A_77_47#_c_432_n 0.00168332f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_104 VPB N_A_77_47#_c_433_n 0.015699f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_105 VPB N_A_77_47#_c_446_n 8.5146e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_106 VPB N_A_77_47#_c_434_n 0.00129067f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_107 VPB N_A_77_47#_c_438_n 0.00185869f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_108 VPB N_A_77_47#_c_439_n 0.00698451f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_109 VPB N_A_63_367#_c_614_n 0.00746637f $X=-0.19 $Y=1.655 $X2=0.8 $Y2=1.42
cc_110 VPB N_A_63_367#_c_615_n 0.0372837f $X=-0.19 $Y=1.655 $X2=1.085 $Y2=2.465
cc_111 VPB N_A_63_367#_c_616_n 0.0018268f $X=-0.19 $Y=1.655 $X2=0.69 $Y2=1.51
cc_112 VPB N_A_63_367#_c_617_n 0.00591924f $X=-0.19 $Y=1.655 $X2=0.37 $Y2=1.51
cc_113 VPB N_A_318_367#_c_646_n 0.0112697f $X=-0.19 $Y=1.655 $X2=1.01 $Y2=1.42
cc_114 VPB N_A_318_367#_c_647_n 0.00213431f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_115 VPB N_A_511_349#_c_672_n 0.0059387f $X=-0.19 $Y=1.655 $X2=1.155 $Y2=1.345
cc_116 VPB N_A_511_349#_c_673_n 0.00614905f $X=-0.19 $Y=1.655 $X2=1.155
+ $Y2=0.655
cc_117 VPB N_A_511_349#_c_674_n 0.00396087f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_118 VPB N_A_511_349#_c_675_n 0.0118892f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_119 VPB N_A_511_349#_c_676_n 0.0119005f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_120 VPB N_A_511_349#_c_677_n 5.3557e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_121 VPB N_VPWR_c_726_n 0.00240833f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_122 VPB N_VPWR_c_727_n 0.0182835f $X=-0.19 $Y=1.655 $X2=0.69 $Y2=1.51
cc_123 VPB N_VPWR_c_728_n 0.0104336f $X=-0.19 $Y=1.655 $X2=0.37 $Y2=1.51
cc_124 VPB N_VPWR_c_729_n 3.0911e-19 $X=-0.19 $Y=1.655 $X2=0.31 $Y2=1.51
cc_125 VPB N_VPWR_c_730_n 3.0911e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_126 VPB N_VPWR_c_731_n 0.0143271f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_127 VPB N_VPWR_c_732_n 0.0412086f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_128 VPB N_VPWR_c_733_n 0.0978523f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_129 VPB N_VPWR_c_734_n 0.0129398f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_130 VPB N_VPWR_c_735_n 0.0129398f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_131 VPB N_VPWR_c_736_n 0.0129398f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_132 VPB N_VPWR_c_737_n 0.00546719f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_133 VPB N_VPWR_c_738_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_134 VPB N_VPWR_c_739_n 0.00435574f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_135 VPB N_VPWR_c_740_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_136 VPB N_VPWR_c_725_n 0.0902605f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_137 VPB N_X_c_838_n 0.0030484f $X=-0.19 $Y=1.655 $X2=0.37 $Y2=1.51
cc_138 VPB N_X_c_839_n 0.00235076f $X=-0.19 $Y=1.655 $X2=0.37 $Y2=1.51
cc_139 VPB N_X_c_840_n 0.00141276f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_140 VPB N_X_c_841_n 0.00144145f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_141 VPB N_X_c_842_n 0.0146499f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_142 VPB X 0.00509812f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_143 N_D1_M1022_g N_C1_M1002_g 0.0226656f $X=1.155 $Y=0.655 $X2=0 $Y2=0
cc_144 N_D1_M1018_g C1 0.00915472f $X=1.085 $Y=2.465 $X2=0 $Y2=0
cc_145 N_D1_c_149_n C1 0.00569498f $X=1.12 $Y=1.42 $X2=0 $Y2=0
cc_146 N_D1_M1018_g N_C1_c_193_n 0.0270296f $X=1.085 $Y=2.465 $X2=0 $Y2=0
cc_147 N_D1_c_149_n N_C1_c_193_n 0.0109718f $X=1.12 $Y=1.42 $X2=0 $Y2=0
cc_148 N_D1_M1022_g N_A_77_47#_c_426_n 0.0147574f $X=1.155 $Y=0.655 $X2=0 $Y2=0
cc_149 N_D1_M1004_g N_A_77_47#_c_427_n 0.0161882f $X=0.725 $Y=0.655 $X2=0 $Y2=0
cc_150 N_D1_c_144_n N_A_77_47#_c_427_n 0.00230653f $X=1.01 $Y=1.42 $X2=0 $Y2=0
cc_151 N_D1_c_147_n N_A_77_47#_c_427_n 0.00951993f $X=0.58 $Y=1.51 $X2=0 $Y2=0
cc_152 N_D1_c_150_n N_A_77_47#_c_427_n 0.0131054f $X=0.37 $Y=1.51 $X2=0 $Y2=0
cc_153 N_D1_M1006_g N_A_77_47#_c_455_n 0.0113007f $X=0.655 $Y=2.465 $X2=0 $Y2=0
cc_154 N_D1_c_144_n N_A_77_47#_c_455_n 0.00138011f $X=1.01 $Y=1.42 $X2=0 $Y2=0
cc_155 N_D1_M1018_g N_A_77_47#_c_455_n 0.0121359f $X=1.085 $Y=2.465 $X2=0 $Y2=0
cc_156 N_D1_M1006_g N_A_77_47#_c_434_n 0.00934402f $X=0.655 $Y=2.465 $X2=0 $Y2=0
cc_157 N_D1_M1004_g N_A_77_47#_c_434_n 0.00622794f $X=0.725 $Y=0.655 $X2=0 $Y2=0
cc_158 N_D1_c_144_n N_A_77_47#_c_434_n 0.00824334f $X=1.01 $Y=1.42 $X2=0 $Y2=0
cc_159 N_D1_M1018_g N_A_77_47#_c_434_n 0.00528155f $X=1.085 $Y=2.465 $X2=0 $Y2=0
cc_160 N_D1_M1022_g N_A_77_47#_c_434_n 0.00248345f $X=1.155 $Y=0.655 $X2=0 $Y2=0
cc_161 N_D1_c_148_n N_A_77_47#_c_434_n 0.0125509f $X=0.69 $Y=1.51 $X2=0 $Y2=0
cc_162 N_D1_c_150_n N_A_77_47#_c_434_n 0.0246093f $X=0.37 $Y=1.51 $X2=0 $Y2=0
cc_163 N_D1_c_147_n N_A_63_367#_c_615_n 0.00165221f $X=0.58 $Y=1.51 $X2=0 $Y2=0
cc_164 N_D1_c_150_n N_A_63_367#_c_615_n 0.0220204f $X=0.37 $Y=1.51 $X2=0 $Y2=0
cc_165 N_D1_M1006_g N_A_63_367#_c_620_n 0.0115031f $X=0.655 $Y=2.465 $X2=0 $Y2=0
cc_166 N_D1_M1018_g N_A_63_367#_c_620_n 0.0115031f $X=1.085 $Y=2.465 $X2=0 $Y2=0
cc_167 N_D1_M1006_g N_VPWR_c_733_n 0.00357877f $X=0.655 $Y=2.465 $X2=0 $Y2=0
cc_168 N_D1_M1018_g N_VPWR_c_733_n 0.00357877f $X=1.085 $Y=2.465 $X2=0 $Y2=0
cc_169 N_D1_M1006_g N_VPWR_c_725_n 0.00641531f $X=0.655 $Y=2.465 $X2=0 $Y2=0
cc_170 N_D1_M1018_g N_VPWR_c_725_n 0.00537654f $X=1.085 $Y=2.465 $X2=0 $Y2=0
cc_171 N_D1_M1004_g N_VGND_c_894_n 0.0128419f $X=0.725 $Y=0.655 $X2=0 $Y2=0
cc_172 N_D1_M1022_g N_VGND_c_894_n 0.0111453f $X=1.155 $Y=0.655 $X2=0 $Y2=0
cc_173 N_D1_M1022_g N_VGND_c_895_n 0.00486043f $X=1.155 $Y=0.655 $X2=0 $Y2=0
cc_174 N_D1_M1004_g N_VGND_c_902_n 0.00486043f $X=0.725 $Y=0.655 $X2=0 $Y2=0
cc_175 N_D1_M1004_g N_VGND_c_914_n 0.00934593f $X=0.725 $Y=0.655 $X2=0 $Y2=0
cc_176 N_D1_M1022_g N_VGND_c_914_n 0.0082726f $X=1.155 $Y=0.655 $X2=0 $Y2=0
cc_177 N_C1_M1012_g N_B1_M1005_g 0.0142043f $X=2.095 $Y=0.655 $X2=0 $Y2=0
cc_178 C1 N_B1_c_247_n 0.0107351f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_179 N_C1_c_193_n N_B1_c_247_n 0.0142043f $X=2.095 $Y=1.51 $X2=0 $Y2=0
cc_180 C1 B1 0.00590724f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_181 C1 N_B1_c_251_n 0.00729958f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_182 N_C1_c_193_n N_B1_c_251_n 0.0033964f $X=2.095 $Y=1.51 $X2=0 $Y2=0
cc_183 C1 N_B1_c_262_n 0.00962719f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_184 C1 N_A_77_47#_c_426_n 0.0114711f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_185 N_C1_M1002_g N_A_77_47#_c_428_n 0.0149477f $X=1.585 $Y=0.655 $X2=0 $Y2=0
cc_186 N_C1_M1012_g N_A_77_47#_c_428_n 0.0149477f $X=2.095 $Y=0.655 $X2=0 $Y2=0
cc_187 C1 N_A_77_47#_c_428_n 0.0345758f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_188 N_C1_c_193_n N_A_77_47#_c_428_n 0.0048507f $X=2.095 $Y=1.51 $X2=0 $Y2=0
cc_189 C1 N_A_77_47#_c_429_n 0.0218601f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_190 C1 N_A_77_47#_c_434_n 0.0277067f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_191 N_C1_c_193_n N_A_77_47#_c_434_n 3.78945e-19 $X=2.095 $Y=1.51 $X2=0 $Y2=0
cc_192 N_C1_M1002_g N_A_77_47#_c_435_n 0.00253148f $X=1.585 $Y=0.655 $X2=0 $Y2=0
cc_193 C1 N_A_77_47#_c_435_n 0.0176969f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_194 N_C1_c_193_n N_A_77_47#_c_435_n 0.00185184f $X=2.095 $Y=1.51 $X2=0 $Y2=0
cc_195 C1 N_A_77_47#_c_436_n 0.0147742f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_196 C1 N_A_63_367#_c_622_n 0.0153635f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_197 N_C1_M1000_g N_A_63_367#_c_616_n 0.0115031f $X=1.515 $Y=2.465 $X2=0 $Y2=0
cc_198 N_C1_M1013_g N_A_63_367#_c_616_n 0.0115031f $X=1.945 $Y=2.465 $X2=0 $Y2=0
cc_199 N_C1_M1013_g N_A_318_367#_c_646_n 0.0131906f $X=1.945 $Y=2.465 $X2=0
+ $Y2=0
cc_200 C1 N_A_318_367#_c_646_n 0.0650203f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_201 N_C1_c_193_n N_A_318_367#_c_646_n 7.12775e-19 $X=2.095 $Y=1.51 $X2=0
+ $Y2=0
cc_202 N_C1_M1000_g N_A_318_367#_c_651_n 0.0109342f $X=1.515 $Y=2.465 $X2=0
+ $Y2=0
cc_203 N_C1_M1013_g N_A_318_367#_c_651_n 0.0154589f $X=1.945 $Y=2.465 $X2=0
+ $Y2=0
cc_204 C1 N_A_318_367#_c_651_n 0.0231556f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_205 N_C1_c_193_n N_A_318_367#_c_651_n 6.18419e-19 $X=2.095 $Y=1.51 $X2=0
+ $Y2=0
cc_206 C1 N_A_318_367#_c_647_n 0.00411603f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_207 C1 N_A_511_349#_M1009_s 0.00248713f $X=2.555 $Y=1.58 $X2=-0.19 $Y2=-0.245
cc_208 N_C1_M1000_g N_VPWR_c_733_n 0.00357877f $X=1.515 $Y=2.465 $X2=0 $Y2=0
cc_209 N_C1_M1013_g N_VPWR_c_733_n 0.00357877f $X=1.945 $Y=2.465 $X2=0 $Y2=0
cc_210 N_C1_M1000_g N_VPWR_c_725_n 0.00537654f $X=1.515 $Y=2.465 $X2=0 $Y2=0
cc_211 N_C1_M1013_g N_VPWR_c_725_n 0.00665089f $X=1.945 $Y=2.465 $X2=0 $Y2=0
cc_212 N_C1_M1002_g N_VGND_c_894_n 6.44378e-19 $X=1.585 $Y=0.655 $X2=0 $Y2=0
cc_213 N_C1_M1002_g N_VGND_c_895_n 0.00585385f $X=1.585 $Y=0.655 $X2=0 $Y2=0
cc_214 N_C1_M1002_g N_VGND_c_896_n 0.00172953f $X=1.585 $Y=0.655 $X2=0 $Y2=0
cc_215 N_C1_M1012_g N_VGND_c_896_n 0.0017281f $X=2.095 $Y=0.655 $X2=0 $Y2=0
cc_216 N_C1_M1012_g N_VGND_c_909_n 0.00585385f $X=2.095 $Y=0.655 $X2=0 $Y2=0
cc_217 N_C1_M1012_g N_VGND_c_910_n 6.41557e-19 $X=2.095 $Y=0.655 $X2=0 $Y2=0
cc_218 N_C1_M1002_g N_VGND_c_914_n 0.0107551f $X=1.585 $Y=0.655 $X2=0 $Y2=0
cc_219 N_C1_M1012_g N_VGND_c_914_n 0.0107551f $X=2.095 $Y=0.655 $X2=0 $Y2=0
cc_220 N_B1_M1014_g N_A1_c_313_n 0.0198426f $X=3.56 $Y=0.655 $X2=-0.19
+ $Y2=-0.245
cc_221 N_B1_M1025_g N_A1_M1015_g 0.0262825f $X=3.325 $Y=2.375 $X2=0 $Y2=0
cc_222 B1 N_A1_M1015_g 0.0191941f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_223 B1 N_A1_c_315_n 2.44763e-19 $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_224 B1 N_A1_M1023_g 6.89199e-19 $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_225 N_B1_c_251_n N_A1_c_318_n 0.0226739f $X=3.56 $Y=1.42 $X2=0 $Y2=0
cc_226 B1 N_A1_c_319_n 0.00203292f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_227 N_B1_M1005_g N_A_77_47#_c_429_n 0.0152237f $X=2.525 $Y=0.655 $X2=0 $Y2=0
cc_228 N_B1_M1014_g N_A_77_47#_c_429_n 0.0152629f $X=3.56 $Y=0.655 $X2=0 $Y2=0
cc_229 N_B1_c_250_n N_A_77_47#_c_429_n 0.0216507f $X=2.82 $Y=1.42 $X2=0 $Y2=0
cc_230 N_B1_c_251_n N_A_77_47#_c_429_n 0.0010994f $X=3.56 $Y=1.42 $X2=0 $Y2=0
cc_231 N_B1_c_262_n N_A_77_47#_c_429_n 0.0502783f $X=3.375 $Y=1.56 $X2=0 $Y2=0
cc_232 B1 N_A_77_47#_c_431_n 0.0217771f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_233 B1 N_A_77_47#_c_432_n 0.0215004f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_234 N_B1_c_251_n N_A_77_47#_c_432_n 2.77945e-19 $X=3.56 $Y=1.42 $X2=0 $Y2=0
cc_235 B1 N_A_77_47#_c_446_n 0.0143571f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_236 B1 N_A_77_47#_c_437_n 0.0163972f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_237 N_B1_c_251_n N_A_77_47#_c_437_n 6.38802e-19 $X=3.56 $Y=1.42 $X2=0 $Y2=0
cc_238 N_B1_M1009_g N_A_63_367#_c_616_n 4.78188e-19 $X=2.895 $Y=2.375 $X2=0
+ $Y2=0
cc_239 N_B1_M1009_g N_A_63_367#_c_617_n 0.00111808f $X=2.895 $Y=2.375 $X2=0
+ $Y2=0
cc_240 N_B1_M1009_g N_A_318_367#_c_646_n 0.0194052f $X=2.895 $Y=2.375 $X2=0
+ $Y2=0
cc_241 N_B1_c_250_n N_A_318_367#_c_646_n 6.28671e-19 $X=2.82 $Y=1.42 $X2=0 $Y2=0
cc_242 N_B1_M1009_g N_A_318_367#_c_647_n 0.00844828f $X=2.895 $Y=2.375 $X2=0
+ $Y2=0
cc_243 N_B1_M1025_g N_A_318_367#_c_647_n 2.9108e-19 $X=3.325 $Y=2.375 $X2=0
+ $Y2=0
cc_244 B1 N_A_318_367#_c_647_n 0.00488049f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_245 N_B1_c_251_n N_A_318_367#_c_647_n 0.00247486f $X=3.56 $Y=1.42 $X2=0 $Y2=0
cc_246 N_B1_c_262_n N_A_318_367#_c_647_n 0.0192218f $X=3.375 $Y=1.56 $X2=0 $Y2=0
cc_247 B1 N_A_511_349#_M1025_s 0.00577051f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_248 N_B1_M1009_g N_A_511_349#_c_672_n 0.00991161f $X=2.895 $Y=2.375 $X2=0
+ $Y2=0
cc_249 N_B1_M1025_g N_A_511_349#_c_672_n 5.87701e-19 $X=3.325 $Y=2.375 $X2=0
+ $Y2=0
cc_250 N_B1_M1009_g N_A_511_349#_c_673_n 0.0102372f $X=2.895 $Y=2.375 $X2=0
+ $Y2=0
cc_251 N_B1_M1025_g N_A_511_349#_c_673_n 0.0147228f $X=3.325 $Y=2.375 $X2=0
+ $Y2=0
cc_252 N_B1_M1009_g N_A_511_349#_c_674_n 0.00194169f $X=2.895 $Y=2.375 $X2=0
+ $Y2=0
cc_253 N_B1_M1025_g N_A_511_349#_c_685_n 0.00208301f $X=3.325 $Y=2.375 $X2=0
+ $Y2=0
cc_254 B1 N_A_511_349#_c_685_n 0.0287331f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_255 N_B1_c_251_n N_A_511_349#_c_685_n 0.00104244f $X=3.56 $Y=1.42 $X2=0 $Y2=0
cc_256 N_B1_M1025_g N_A_511_349#_c_688_n 0.00956635f $X=3.325 $Y=2.375 $X2=0
+ $Y2=0
cc_257 B1 N_A_511_349#_c_689_n 0.0169014f $X=3.995 $Y=1.58 $X2=0 $Y2=0
cc_258 B1 N_VPWR_M1015_s 8.19824e-19 $X=3.995 $Y=1.58 $X2=-0.19 $Y2=-0.245
cc_259 N_B1_M1025_g N_VPWR_c_726_n 5.57444e-19 $X=3.325 $Y=2.375 $X2=0 $Y2=0
cc_260 N_B1_M1009_g N_VPWR_c_733_n 0.00302473f $X=2.895 $Y=2.375 $X2=0 $Y2=0
cc_261 N_B1_M1025_g N_VPWR_c_733_n 0.00302501f $X=3.325 $Y=2.375 $X2=0 $Y2=0
cc_262 N_B1_M1009_g N_VPWR_c_725_n 0.00484658f $X=2.895 $Y=2.375 $X2=0 $Y2=0
cc_263 N_B1_M1025_g N_VPWR_c_725_n 0.00453511f $X=3.325 $Y=2.375 $X2=0 $Y2=0
cc_264 N_B1_M1014_g N_VGND_c_904_n 0.00486043f $X=3.56 $Y=0.655 $X2=0 $Y2=0
cc_265 N_B1_M1005_g N_VGND_c_909_n 0.00486043f $X=2.525 $Y=0.655 $X2=0 $Y2=0
cc_266 N_B1_M1005_g N_VGND_c_910_n 0.0116906f $X=2.525 $Y=0.655 $X2=0 $Y2=0
cc_267 N_B1_M1014_g N_VGND_c_910_n 0.0127907f $X=3.56 $Y=0.655 $X2=0 $Y2=0
cc_268 N_B1_M1005_g N_VGND_c_914_n 0.00822376f $X=2.525 $Y=0.655 $X2=0 $Y2=0
cc_269 N_B1_M1014_g N_VGND_c_914_n 0.00822376f $X=3.56 $Y=0.655 $X2=0 $Y2=0
cc_270 A1 N_A2_c_381_n 0.0197774f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_271 N_A1_c_321_n N_A2_c_381_n 2.28319e-19 $X=4.86 $Y=1.35 $X2=0 $Y2=0
cc_272 A1 N_A2_c_378_n 0.00182191f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_273 N_A1_c_321_n N_A2_c_378_n 0.0147198f $X=4.86 $Y=1.35 $X2=0 $Y2=0
cc_274 N_A1_c_313_n N_A_77_47#_c_430_n 0.0100732f $X=3.99 $Y=1.185 $X2=0 $Y2=0
cc_275 N_A1_c_316_n N_A_77_47#_c_430_n 0.0086866f $X=4.42 $Y=1.185 $X2=0 $Y2=0
cc_276 N_A1_c_313_n N_A_77_47#_c_431_n 0.0107334f $X=3.99 $Y=1.185 $X2=0 $Y2=0
cc_277 N_A1_c_315_n N_A_77_47#_c_431_n 0.00381847f $X=4.345 $Y=1.26 $X2=0 $Y2=0
cc_278 N_A1_c_316_n N_A_77_47#_c_431_n 0.00902926f $X=4.42 $Y=1.185 $X2=0 $Y2=0
cc_279 N_A1_M1015_g N_A_77_47#_c_432_n 3.0349e-19 $X=3.99 $Y=2.375 $X2=0 $Y2=0
cc_280 N_A1_c_316_n N_A_77_47#_c_432_n 0.00114834f $X=4.42 $Y=1.185 $X2=0 $Y2=0
cc_281 N_A1_M1023_g N_A_77_47#_c_432_n 0.00321319f $X=4.42 $Y=2.375 $X2=0 $Y2=0
cc_282 N_A1_c_319_n N_A_77_47#_c_432_n 0.00989839f $X=4.42 $Y=1.35 $X2=0 $Y2=0
cc_283 A1 N_A_77_47#_c_432_n 0.016451f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_284 N_A1_c_321_n N_A_77_47#_c_432_n 0.00857804f $X=4.86 $Y=1.35 $X2=0 $Y2=0
cc_285 A1 N_A_77_47#_c_433_n 0.0353654f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_286 N_A1_c_321_n N_A_77_47#_c_433_n 0.0151996f $X=4.86 $Y=1.35 $X2=0 $Y2=0
cc_287 N_A1_M1023_g N_A_77_47#_c_446_n 0.00866676f $X=4.42 $Y=2.375 $X2=0 $Y2=0
cc_288 N_A1_M1015_g N_A_511_349#_c_673_n 0.00187224f $X=3.99 $Y=2.375 $X2=0
+ $Y2=0
cc_289 N_A1_M1015_g N_A_511_349#_c_688_n 0.0111042f $X=3.99 $Y=2.375 $X2=0 $Y2=0
cc_290 N_A1_M1015_g N_A_511_349#_c_689_n 0.0150835f $X=3.99 $Y=2.375 $X2=0 $Y2=0
cc_291 N_A1_c_315_n N_A_511_349#_c_689_n 0.00194301f $X=4.345 $Y=1.26 $X2=0
+ $Y2=0
cc_292 N_A1_M1023_g N_A_511_349#_c_689_n 0.012226f $X=4.42 $Y=2.375 $X2=0 $Y2=0
cc_293 N_A1_M1023_g N_A_511_349#_c_675_n 0.0012215f $X=4.42 $Y=2.375 $X2=0 $Y2=0
cc_294 N_A1_M1015_g N_VPWR_c_726_n 0.0132163f $X=3.99 $Y=2.375 $X2=0 $Y2=0
cc_295 N_A1_M1023_g N_VPWR_c_726_n 0.0128134f $X=4.42 $Y=2.375 $X2=0 $Y2=0
cc_296 N_A1_M1023_g N_VPWR_c_727_n 0.00414769f $X=4.42 $Y=2.375 $X2=0 $Y2=0
cc_297 N_A1_M1023_g N_VPWR_c_728_n 0.00270101f $X=4.42 $Y=2.375 $X2=0 $Y2=0
cc_298 N_A1_M1015_g N_VPWR_c_733_n 0.00414769f $X=3.99 $Y=2.375 $X2=0 $Y2=0
cc_299 N_A1_M1015_g N_VPWR_c_725_n 0.00806345f $X=3.99 $Y=2.375 $X2=0 $Y2=0
cc_300 N_A1_M1023_g N_VPWR_c_725_n 0.00837493f $X=4.42 $Y=2.375 $X2=0 $Y2=0
cc_301 N_A1_c_316_n N_VGND_c_897_n 0.00418794f $X=4.42 $Y=1.185 $X2=0 $Y2=0
cc_302 N_A1_c_313_n N_VGND_c_904_n 0.00357877f $X=3.99 $Y=1.185 $X2=0 $Y2=0
cc_303 N_A1_c_316_n N_VGND_c_904_n 0.00357877f $X=4.42 $Y=1.185 $X2=0 $Y2=0
cc_304 N_A1_c_313_n N_VGND_c_910_n 0.00116005f $X=3.99 $Y=1.185 $X2=0 $Y2=0
cc_305 N_A1_c_313_n N_VGND_c_914_n 0.00537654f $X=3.99 $Y=1.185 $X2=0 $Y2=0
cc_306 N_A1_c_316_n N_VGND_c_914_n 0.00665089f $X=4.42 $Y=1.185 $X2=0 $Y2=0
cc_307 N_A1_c_313_n N_A_813_47#_c_1016_n 0.00246154f $X=3.99 $Y=1.185 $X2=0
+ $Y2=0
cc_308 N_A1_c_316_n N_A_813_47#_c_1016_n 0.0104679f $X=4.42 $Y=1.185 $X2=0 $Y2=0
cc_309 N_A1_c_321_n N_A_813_47#_c_1016_n 0.00467265f $X=4.86 $Y=1.35 $X2=0 $Y2=0
cc_310 N_A1_c_316_n N_A_813_47#_c_1015_n 0.00724828f $X=4.42 $Y=1.185 $X2=0
+ $Y2=0
cc_311 A1 N_A_813_47#_c_1015_n 0.0368057f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_312 N_A1_c_321_n N_A_813_47#_c_1015_n 0.00803572f $X=4.86 $Y=1.35 $X2=0 $Y2=0
cc_313 N_A2_c_376_n N_A_77_47#_M1007_g 0.0205086f $X=5.84 $Y=1.185 $X2=0 $Y2=0
cc_314 N_A2_c_381_n N_A_77_47#_M1007_g 0.00108724f $X=5.685 $Y=1.35 $X2=0 $Y2=0
cc_315 N_A2_M1020_g N_A_77_47#_M1011_g 0.0205086f $X=5.84 $Y=2.465 $X2=0 $Y2=0
cc_316 N_A2_c_374_n N_A_77_47#_c_430_n 4.6165e-19 $X=5.41 $Y=1.185 $X2=0 $Y2=0
cc_317 N_A2_M1001_g N_A_77_47#_c_433_n 0.0125516f $X=5.41 $Y=2.465 $X2=0 $Y2=0
cc_318 N_A2_M1020_g N_A_77_47#_c_433_n 0.0149455f $X=5.84 $Y=2.465 $X2=0 $Y2=0
cc_319 N_A2_c_381_n N_A_77_47#_c_433_n 0.0365006f $X=5.685 $Y=1.35 $X2=0 $Y2=0
cc_320 N_A2_c_378_n N_A_77_47#_c_433_n 0.00243542f $X=5.84 $Y=1.35 $X2=0 $Y2=0
cc_321 N_A2_M1020_g N_A_77_47#_c_438_n 2.30627e-19 $X=5.84 $Y=2.465 $X2=0 $Y2=0
cc_322 N_A2_c_381_n N_A_77_47#_c_438_n 0.00305897f $X=5.685 $Y=1.35 $X2=0 $Y2=0
cc_323 N_A2_c_378_n N_A_77_47#_c_438_n 0.00429049f $X=5.84 $Y=1.35 $X2=0 $Y2=0
cc_324 N_A2_c_378_n N_A_77_47#_c_439_n 0.0205086f $X=5.84 $Y=1.35 $X2=0 $Y2=0
cc_325 N_A2_M1001_g N_A_511_349#_c_675_n 0.00486687f $X=5.41 $Y=2.465 $X2=0
+ $Y2=0
cc_326 N_A2_M1001_g N_A_511_349#_c_676_n 0.0144916f $X=5.41 $Y=2.465 $X2=0 $Y2=0
cc_327 N_A2_M1001_g N_VPWR_c_728_n 0.016101f $X=5.41 $Y=2.465 $X2=0 $Y2=0
cc_328 N_A2_M1020_g N_VPWR_c_728_n 7.06778e-19 $X=5.84 $Y=2.465 $X2=0 $Y2=0
cc_329 N_A2_M1001_g N_VPWR_c_729_n 8.11048e-19 $X=5.41 $Y=2.465 $X2=0 $Y2=0
cc_330 N_A2_M1020_g N_VPWR_c_729_n 0.017107f $X=5.84 $Y=2.465 $X2=0 $Y2=0
cc_331 N_A2_M1001_g N_VPWR_c_734_n 0.00486043f $X=5.41 $Y=2.465 $X2=0 $Y2=0
cc_332 N_A2_M1020_g N_VPWR_c_734_n 0.00486043f $X=5.84 $Y=2.465 $X2=0 $Y2=0
cc_333 N_A2_M1001_g N_VPWR_c_725_n 0.00835506f $X=5.41 $Y=2.465 $X2=0 $Y2=0
cc_334 N_A2_M1020_g N_VPWR_c_725_n 0.00835506f $X=5.84 $Y=2.465 $X2=0 $Y2=0
cc_335 N_A2_c_381_n N_X_c_833_n 8.6987e-19 $X=5.685 $Y=1.35 $X2=0 $Y2=0
cc_336 N_A2_c_374_n N_VGND_c_897_n 0.00943681f $X=5.41 $Y=1.185 $X2=0 $Y2=0
cc_337 N_A2_c_376_n N_VGND_c_897_n 5.44696e-19 $X=5.84 $Y=1.185 $X2=0 $Y2=0
cc_338 N_A2_c_374_n N_VGND_c_898_n 5.93071e-19 $X=5.41 $Y=1.185 $X2=0 $Y2=0
cc_339 N_A2_c_376_n N_VGND_c_898_n 0.014628f $X=5.84 $Y=1.185 $X2=0 $Y2=0
cc_340 N_A2_c_374_n N_VGND_c_905_n 0.00367954f $X=5.41 $Y=1.185 $X2=0 $Y2=0
cc_341 N_A2_c_376_n N_VGND_c_905_n 0.00486043f $X=5.84 $Y=1.185 $X2=0 $Y2=0
cc_342 N_A2_c_374_n N_VGND_c_914_n 0.00437452f $X=5.41 $Y=1.185 $X2=0 $Y2=0
cc_343 N_A2_c_376_n N_VGND_c_914_n 0.00824727f $X=5.84 $Y=1.185 $X2=0 $Y2=0
cc_344 N_A2_c_374_n N_A_813_47#_c_1014_n 0.01621f $X=5.41 $Y=1.185 $X2=0 $Y2=0
cc_345 N_A2_c_381_n N_A_813_47#_c_1014_n 0.0120367f $X=5.685 $Y=1.35 $X2=0 $Y2=0
cc_346 N_A2_c_381_n N_A_813_47#_c_1024_n 0.01425f $X=5.685 $Y=1.35 $X2=0 $Y2=0
cc_347 N_A2_c_378_n N_A_813_47#_c_1024_n 0.00240082f $X=5.84 $Y=1.35 $X2=0 $Y2=0
cc_348 N_A2_c_374_n N_A_813_47#_c_1015_n 0.00195518f $X=5.41 $Y=1.185 $X2=0
+ $Y2=0
cc_349 N_A_77_47#_M1006_s N_A_63_367#_c_620_n 0.00332344f $X=0.73 $Y=1.835 $X2=0
+ $Y2=0
cc_350 N_A_77_47#_c_455_n N_A_63_367#_c_620_n 0.0159805f $X=0.87 $Y=2.03 $X2=0
+ $Y2=0
cc_351 N_A_77_47#_c_433_n N_A_511_349#_M1023_d 0.00239457f $X=6.02 $Y=1.7 $X2=0
+ $Y2=0
cc_352 N_A_77_47#_c_446_n N_A_511_349#_c_689_n 0.0113161f $X=4.515 $Y=1.7 $X2=0
+ $Y2=0
cc_353 N_A_77_47#_c_433_n N_A_511_349#_c_676_n 0.0643198f $X=6.02 $Y=1.7 $X2=0
+ $Y2=0
cc_354 N_A_77_47#_c_433_n N_A_511_349#_c_677_n 0.0203009f $X=6.02 $Y=1.7 $X2=0
+ $Y2=0
cc_355 N_A_77_47#_M1011_g N_VPWR_c_729_n 0.0172227f $X=6.27 $Y=2.465 $X2=0 $Y2=0
cc_356 N_A_77_47#_M1017_g N_VPWR_c_729_n 7.66778e-19 $X=6.7 $Y=2.465 $X2=0 $Y2=0
cc_357 N_A_77_47#_c_433_n N_VPWR_c_729_n 0.00791023f $X=6.02 $Y=1.7 $X2=0 $Y2=0
cc_358 N_A_77_47#_c_523_p N_VPWR_c_729_n 7.56038e-19 $X=7.38 $Y=1.49 $X2=0 $Y2=0
cc_359 N_A_77_47#_c_438_n N_VPWR_c_729_n 0.0130252f $X=6.11 $Y=1.49 $X2=0 $Y2=0
cc_360 N_A_77_47#_M1011_g N_VPWR_c_730_n 7.27171e-19 $X=6.27 $Y=2.465 $X2=0
+ $Y2=0
cc_361 N_A_77_47#_M1017_g N_VPWR_c_730_n 0.0143393f $X=6.7 $Y=2.465 $X2=0 $Y2=0
cc_362 N_A_77_47#_M1024_g N_VPWR_c_730_n 0.0143393f $X=7.13 $Y=2.465 $X2=0 $Y2=0
cc_363 N_A_77_47#_M1026_g N_VPWR_c_730_n 7.27171e-19 $X=7.56 $Y=2.465 $X2=0
+ $Y2=0
cc_364 N_A_77_47#_M1024_g N_VPWR_c_732_n 7.24342e-19 $X=7.13 $Y=2.465 $X2=0
+ $Y2=0
cc_365 N_A_77_47#_M1026_g N_VPWR_c_732_n 0.0151914f $X=7.56 $Y=2.465 $X2=0 $Y2=0
cc_366 N_A_77_47#_M1011_g N_VPWR_c_735_n 0.00486043f $X=6.27 $Y=2.465 $X2=0
+ $Y2=0
cc_367 N_A_77_47#_M1017_g N_VPWR_c_735_n 0.00486043f $X=6.7 $Y=2.465 $X2=0 $Y2=0
cc_368 N_A_77_47#_M1024_g N_VPWR_c_736_n 0.00486043f $X=7.13 $Y=2.465 $X2=0
+ $Y2=0
cc_369 N_A_77_47#_M1026_g N_VPWR_c_736_n 0.00486043f $X=7.56 $Y=2.465 $X2=0
+ $Y2=0
cc_370 N_A_77_47#_M1006_s N_VPWR_c_725_n 0.00225186f $X=0.73 $Y=1.835 $X2=0
+ $Y2=0
cc_371 N_A_77_47#_M1011_g N_VPWR_c_725_n 0.00824727f $X=6.27 $Y=2.465 $X2=0
+ $Y2=0
cc_372 N_A_77_47#_M1017_g N_VPWR_c_725_n 0.00824727f $X=6.7 $Y=2.465 $X2=0 $Y2=0
cc_373 N_A_77_47#_M1024_g N_VPWR_c_725_n 0.00824727f $X=7.13 $Y=2.465 $X2=0
+ $Y2=0
cc_374 N_A_77_47#_M1026_g N_VPWR_c_725_n 0.00824727f $X=7.56 $Y=2.465 $X2=0
+ $Y2=0
cc_375 N_A_77_47#_M1008_g N_X_c_832_n 0.0137525f $X=6.7 $Y=0.655 $X2=0 $Y2=0
cc_376 N_A_77_47#_M1019_g N_X_c_832_n 0.0141287f $X=7.13 $Y=0.655 $X2=0 $Y2=0
cc_377 N_A_77_47#_c_523_p N_X_c_832_n 0.0467265f $X=7.38 $Y=1.49 $X2=0 $Y2=0
cc_378 N_A_77_47#_c_439_n N_X_c_832_n 0.00246472f $X=7.56 $Y=1.49 $X2=0 $Y2=0
cc_379 N_A_77_47#_M1007_g N_X_c_833_n 0.00468797f $X=6.27 $Y=0.655 $X2=0 $Y2=0
cc_380 N_A_77_47#_c_523_p N_X_c_833_n 0.0153308f $X=7.38 $Y=1.49 $X2=0 $Y2=0
cc_381 N_A_77_47#_c_439_n N_X_c_833_n 0.00256759f $X=7.56 $Y=1.49 $X2=0 $Y2=0
cc_382 N_A_77_47#_M1017_g N_X_c_838_n 0.0133903f $X=6.7 $Y=2.465 $X2=0 $Y2=0
cc_383 N_A_77_47#_M1024_g N_X_c_838_n 0.0135857f $X=7.13 $Y=2.465 $X2=0 $Y2=0
cc_384 N_A_77_47#_c_523_p N_X_c_838_n 0.0469373f $X=7.38 $Y=1.49 $X2=0 $Y2=0
cc_385 N_A_77_47#_c_439_n N_X_c_838_n 0.00246815f $X=7.56 $Y=1.49 $X2=0 $Y2=0
cc_386 N_A_77_47#_M1011_g N_X_c_839_n 0.00192093f $X=6.27 $Y=2.465 $X2=0 $Y2=0
cc_387 N_A_77_47#_c_523_p N_X_c_839_n 0.0153308f $X=7.38 $Y=1.49 $X2=0 $Y2=0
cc_388 N_A_77_47#_c_438_n N_X_c_839_n 0.0029796f $X=6.11 $Y=1.49 $X2=0 $Y2=0
cc_389 N_A_77_47#_c_439_n N_X_c_839_n 0.00256759f $X=7.56 $Y=1.49 $X2=0 $Y2=0
cc_390 N_A_77_47#_M1027_g N_X_c_834_n 0.0168048f $X=7.56 $Y=0.655 $X2=0 $Y2=0
cc_391 N_A_77_47#_c_523_p N_X_c_834_n 0.0072485f $X=7.38 $Y=1.49 $X2=0 $Y2=0
cc_392 N_A_77_47#_M1026_g N_X_c_840_n 0.0163713f $X=7.56 $Y=2.465 $X2=0 $Y2=0
cc_393 N_A_77_47#_c_523_p N_X_c_840_n 0.00728094f $X=7.38 $Y=1.49 $X2=0 $Y2=0
cc_394 N_A_77_47#_c_523_p N_X_c_835_n 0.0153308f $X=7.38 $Y=1.49 $X2=0 $Y2=0
cc_395 N_A_77_47#_c_439_n N_X_c_835_n 0.00256759f $X=7.56 $Y=1.49 $X2=0 $Y2=0
cc_396 N_A_77_47#_c_523_p N_X_c_841_n 0.0153308f $X=7.38 $Y=1.49 $X2=0 $Y2=0
cc_397 N_A_77_47#_c_439_n N_X_c_841_n 0.00256759f $X=7.56 $Y=1.49 $X2=0 $Y2=0
cc_398 N_A_77_47#_M1027_g X 0.0203636f $X=7.56 $Y=0.655 $X2=0 $Y2=0
cc_399 N_A_77_47#_c_523_p X 0.0141892f $X=7.38 $Y=1.49 $X2=0 $Y2=0
cc_400 N_A_77_47#_c_426_n N_VGND_M1004_d 9.47283e-19 $X=1.275 $Y=1.15 $X2=-0.19
+ $Y2=-0.245
cc_401 N_A_77_47#_c_427_n N_VGND_M1004_d 8.49288e-19 $X=0.935 $Y=1.15 $X2=-0.19
+ $Y2=-0.245
cc_402 N_A_77_47#_c_428_n N_VGND_M1002_d 0.00261503f $X=2.175 $Y=1.07 $X2=0
+ $Y2=0
cc_403 N_A_77_47#_c_429_n N_VGND_M1005_s 0.0108021f $X=3.68 $Y=1.07 $X2=0 $Y2=0
cc_404 N_A_77_47#_c_427_n N_VGND_c_894_n 0.0163165f $X=0.935 $Y=1.15 $X2=0 $Y2=0
cc_405 N_A_77_47#_c_570_p N_VGND_c_895_n 0.0138717f $X=1.37 $Y=0.42 $X2=0 $Y2=0
cc_406 N_A_77_47#_c_428_n N_VGND_c_896_n 0.0200142f $X=2.175 $Y=1.07 $X2=0 $Y2=0
cc_407 N_A_77_47#_c_430_n N_VGND_c_897_n 0.0148801f $X=4.635 $Y=0.37 $X2=0 $Y2=0
cc_408 N_A_77_47#_M1007_g N_VGND_c_898_n 0.014416f $X=6.27 $Y=0.655 $X2=0 $Y2=0
cc_409 N_A_77_47#_M1008_g N_VGND_c_898_n 6.72004e-19 $X=6.7 $Y=0.655 $X2=0 $Y2=0
cc_410 N_A_77_47#_c_433_n N_VGND_c_898_n 0.0032168f $X=6.02 $Y=1.7 $X2=0 $Y2=0
cc_411 N_A_77_47#_c_523_p N_VGND_c_898_n 7.81623e-19 $X=7.38 $Y=1.49 $X2=0 $Y2=0
cc_412 N_A_77_47#_c_438_n N_VGND_c_898_n 0.00752936f $X=6.11 $Y=1.49 $X2=0 $Y2=0
cc_413 N_A_77_47#_M1007_g N_VGND_c_899_n 6.30983e-19 $X=6.27 $Y=0.655 $X2=0
+ $Y2=0
cc_414 N_A_77_47#_M1008_g N_VGND_c_899_n 0.0115056f $X=6.7 $Y=0.655 $X2=0 $Y2=0
cc_415 N_A_77_47#_M1019_g N_VGND_c_899_n 0.0115056f $X=7.13 $Y=0.655 $X2=0 $Y2=0
cc_416 N_A_77_47#_M1027_g N_VGND_c_899_n 6.30983e-19 $X=7.56 $Y=0.655 $X2=0
+ $Y2=0
cc_417 N_A_77_47#_M1019_g N_VGND_c_901_n 6.30983e-19 $X=7.13 $Y=0.655 $X2=0
+ $Y2=0
cc_418 N_A_77_47#_M1027_g N_VGND_c_901_n 0.0126581f $X=7.56 $Y=0.655 $X2=0 $Y2=0
cc_419 N_A_77_47#_c_425_n N_VGND_c_902_n 0.0178111f $X=0.51 $Y=0.42 $X2=0 $Y2=0
cc_420 N_A_77_47#_c_585_p N_VGND_c_904_n 0.0125234f $X=3.775 $Y=0.465 $X2=0
+ $Y2=0
cc_421 N_A_77_47#_c_430_n N_VGND_c_904_n 0.0529145f $X=4.635 $Y=0.37 $X2=0 $Y2=0
cc_422 N_A_77_47#_M1007_g N_VGND_c_906_n 0.00486043f $X=6.27 $Y=0.655 $X2=0
+ $Y2=0
cc_423 N_A_77_47#_M1008_g N_VGND_c_906_n 0.00486043f $X=6.7 $Y=0.655 $X2=0 $Y2=0
cc_424 N_A_77_47#_M1019_g N_VGND_c_907_n 0.00486043f $X=7.13 $Y=0.655 $X2=0
+ $Y2=0
cc_425 N_A_77_47#_M1027_g N_VGND_c_907_n 0.00486043f $X=7.56 $Y=0.655 $X2=0
+ $Y2=0
cc_426 N_A_77_47#_c_591_p N_VGND_c_909_n 0.0138717f $X=2.31 $Y=0.42 $X2=0 $Y2=0
cc_427 N_A_77_47#_c_429_n N_VGND_c_910_n 0.0661592f $X=3.68 $Y=1.07 $X2=0 $Y2=0
cc_428 N_A_77_47#_M1004_s N_VGND_c_914_n 0.00371702f $X=0.385 $Y=0.235 $X2=0
+ $Y2=0
cc_429 N_A_77_47#_M1022_s N_VGND_c_914_n 0.00397496f $X=1.23 $Y=0.235 $X2=0
+ $Y2=0
cc_430 N_A_77_47#_M1012_s N_VGND_c_914_n 0.00397496f $X=2.17 $Y=0.235 $X2=0
+ $Y2=0
cc_431 N_A_77_47#_M1014_d N_VGND_c_914_n 0.00376627f $X=3.635 $Y=0.235 $X2=0
+ $Y2=0
cc_432 N_A_77_47#_M1016_d N_VGND_c_914_n 0.00231933f $X=4.495 $Y=0.235 $X2=0
+ $Y2=0
cc_433 N_A_77_47#_M1007_g N_VGND_c_914_n 0.00824727f $X=6.27 $Y=0.655 $X2=0
+ $Y2=0
cc_434 N_A_77_47#_M1008_g N_VGND_c_914_n 0.00824727f $X=6.7 $Y=0.655 $X2=0 $Y2=0
cc_435 N_A_77_47#_M1019_g N_VGND_c_914_n 0.00824727f $X=7.13 $Y=0.655 $X2=0
+ $Y2=0
cc_436 N_A_77_47#_M1027_g N_VGND_c_914_n 0.00824727f $X=7.56 $Y=0.655 $X2=0
+ $Y2=0
cc_437 N_A_77_47#_c_425_n N_VGND_c_914_n 0.0100304f $X=0.51 $Y=0.42 $X2=0 $Y2=0
cc_438 N_A_77_47#_c_570_p N_VGND_c_914_n 0.00886411f $X=1.37 $Y=0.42 $X2=0 $Y2=0
cc_439 N_A_77_47#_c_591_p N_VGND_c_914_n 0.00886411f $X=2.31 $Y=0.42 $X2=0 $Y2=0
cc_440 N_A_77_47#_c_585_p N_VGND_c_914_n 0.00738676f $X=3.775 $Y=0.465 $X2=0
+ $Y2=0
cc_441 N_A_77_47#_c_430_n N_VGND_c_914_n 0.033612f $X=4.635 $Y=0.37 $X2=0 $Y2=0
cc_442 N_A_77_47#_c_430_n N_A_813_47#_M1003_s 0.0033495f $X=4.635 $Y=0.37
+ $X2=-0.19 $Y2=-0.245
cc_443 N_A_77_47#_c_431_n N_A_813_47#_M1003_s 0.00176891f $X=4.345 $Y=1.07
+ $X2=-0.19 $Y2=-0.245
cc_444 N_A_77_47#_M1016_d N_A_813_47#_c_1016_n 0.00326365f $X=4.495 $Y=0.235
+ $X2=0 $Y2=0
cc_445 N_A_77_47#_c_430_n N_A_813_47#_c_1016_n 0.0410142f $X=4.635 $Y=0.37 $X2=0
+ $Y2=0
cc_446 N_A_77_47#_c_431_n N_A_813_47#_c_1016_n 0.0252139f $X=4.345 $Y=1.07 $X2=0
+ $Y2=0
cc_447 N_A_77_47#_M1016_d N_A_813_47#_c_1015_n 0.00675588f $X=4.495 $Y=0.235
+ $X2=0 $Y2=0
cc_448 N_A_77_47#_c_433_n N_A_813_47#_c_1015_n 0.00482382f $X=6.02 $Y=1.7 $X2=0
+ $Y2=0
cc_449 N_A_63_367#_c_616_n N_A_318_367#_M1000_s 0.00332344f $X=2.065 $Y=2.99
+ $X2=-0.19 $Y2=1.655
cc_450 N_A_63_367#_M1013_d N_A_318_367#_c_646_n 0.00503353f $X=2.02 $Y=1.835
+ $X2=0 $Y2=0
cc_451 N_A_63_367#_c_617_n N_A_318_367#_c_646_n 0.0202165f $X=2.16 $Y=2.445
+ $X2=0 $Y2=0
cc_452 N_A_63_367#_c_616_n N_A_318_367#_c_651_n 0.0159805f $X=2.065 $Y=2.99
+ $X2=0 $Y2=0
cc_453 N_A_63_367#_c_617_n N_A_511_349#_c_672_n 0.0471978f $X=2.16 $Y=2.445
+ $X2=0 $Y2=0
cc_454 N_A_63_367#_c_616_n N_A_511_349#_c_674_n 0.0147157f $X=2.065 $Y=2.99
+ $X2=0 $Y2=0
cc_455 N_A_63_367#_c_614_n N_VPWR_c_733_n 0.0179183f $X=0.405 $Y=2.905 $X2=0
+ $Y2=0
cc_456 N_A_63_367#_c_620_n N_VPWR_c_733_n 0.0361172f $X=1.205 $Y=2.99 $X2=0
+ $Y2=0
cc_457 N_A_63_367#_c_616_n N_VPWR_c_733_n 0.0540354f $X=2.065 $Y=2.99 $X2=0
+ $Y2=0
cc_458 N_A_63_367#_c_638_p N_VPWR_c_733_n 0.0125234f $X=1.3 $Y=2.91 $X2=0 $Y2=0
cc_459 N_A_63_367#_M1006_d N_VPWR_c_725_n 0.00215161f $X=0.315 $Y=1.835 $X2=0
+ $Y2=0
cc_460 N_A_63_367#_M1018_d N_VPWR_c_725_n 0.00223565f $X=1.16 $Y=1.835 $X2=0
+ $Y2=0
cc_461 N_A_63_367#_M1013_d N_VPWR_c_725_n 0.00215161f $X=2.02 $Y=1.835 $X2=0
+ $Y2=0
cc_462 N_A_63_367#_c_614_n N_VPWR_c_725_n 0.0101082f $X=0.405 $Y=2.905 $X2=0
+ $Y2=0
cc_463 N_A_63_367#_c_620_n N_VPWR_c_725_n 0.023676f $X=1.205 $Y=2.99 $X2=0 $Y2=0
cc_464 N_A_63_367#_c_616_n N_VPWR_c_725_n 0.0337842f $X=2.065 $Y=2.99 $X2=0
+ $Y2=0
cc_465 N_A_63_367#_c_638_p N_VPWR_c_725_n 0.00738676f $X=1.3 $Y=2.91 $X2=0 $Y2=0
cc_466 N_A_318_367#_c_646_n N_A_511_349#_M1009_s 0.00499247f $X=2.965 $Y=2.025
+ $X2=-0.19 $Y2=1.655
cc_467 N_A_318_367#_c_646_n N_A_511_349#_c_672_n 0.0220026f $X=2.965 $Y=2.025
+ $X2=0 $Y2=0
cc_468 N_A_318_367#_M1009_d N_A_511_349#_c_673_n 0.00176461f $X=2.97 $Y=1.745
+ $X2=0 $Y2=0
cc_469 N_A_318_367#_c_670_p N_A_511_349#_c_673_n 0.0126348f $X=3.11 $Y=2.21
+ $X2=0 $Y2=0
cc_470 N_A_318_367#_M1000_s N_VPWR_c_725_n 0.00225186f $X=1.59 $Y=1.835 $X2=0
+ $Y2=0
cc_471 N_A_511_349#_c_689_n N_VPWR_M1015_s 0.00500673f $X=4.54 $Y=2.04 $X2=-0.19
+ $Y2=1.655
cc_472 N_A_511_349#_c_676_n N_VPWR_M1001_s 0.00521795f $X=5.53 $Y=2.04 $X2=0
+ $Y2=0
cc_473 N_A_511_349#_c_673_n N_VPWR_c_726_n 0.0118397f $X=3.495 $Y=2.99 $X2=0
+ $Y2=0
cc_474 N_A_511_349#_c_688_n N_VPWR_c_726_n 0.0394963f $X=3.66 $Y=2.445 $X2=0
+ $Y2=0
cc_475 N_A_511_349#_c_689_n N_VPWR_c_726_n 0.0170436f $X=4.54 $Y=2.04 $X2=0
+ $Y2=0
cc_476 N_A_511_349#_c_675_n N_VPWR_c_726_n 0.0281538f $X=4.635 $Y=2.46 $X2=0
+ $Y2=0
cc_477 N_A_511_349#_c_675_n N_VPWR_c_727_n 0.0140356f $X=4.635 $Y=2.46 $X2=0
+ $Y2=0
cc_478 N_A_511_349#_c_675_n N_VPWR_c_728_n 0.0483431f $X=4.635 $Y=2.46 $X2=0
+ $Y2=0
cc_479 N_A_511_349#_c_676_n N_VPWR_c_728_n 0.0220026f $X=5.53 $Y=2.04 $X2=0
+ $Y2=0
cc_480 N_A_511_349#_c_673_n N_VPWR_c_733_n 0.0646726f $X=3.495 $Y=2.99 $X2=0
+ $Y2=0
cc_481 N_A_511_349#_c_674_n N_VPWR_c_733_n 0.0235688f $X=2.845 $Y=2.99 $X2=0
+ $Y2=0
cc_482 N_A_511_349#_c_719_p N_VPWR_c_734_n 0.0124525f $X=5.625 $Y=2.17 $X2=0
+ $Y2=0
cc_483 N_A_511_349#_M1001_d N_VPWR_c_725_n 0.00545212f $X=5.485 $Y=1.835 $X2=0
+ $Y2=0
cc_484 N_A_511_349#_c_673_n N_VPWR_c_725_n 0.0360093f $X=3.495 $Y=2.99 $X2=0
+ $Y2=0
cc_485 N_A_511_349#_c_674_n N_VPWR_c_725_n 0.0127152f $X=2.845 $Y=2.99 $X2=0
+ $Y2=0
cc_486 N_A_511_349#_c_675_n N_VPWR_c_725_n 0.00977851f $X=4.635 $Y=2.46 $X2=0
+ $Y2=0
cc_487 N_A_511_349#_c_719_p N_VPWR_c_725_n 0.00730901f $X=5.625 $Y=2.17 $X2=0
+ $Y2=0
cc_488 N_VPWR_c_725_n N_X_M1011_d 0.00536646f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_489 N_VPWR_c_725_n N_X_M1024_d 0.00536646f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_490 N_VPWR_c_735_n N_X_c_872_n 0.0124525f $X=6.75 $Y=3.33 $X2=0 $Y2=0
cc_491 N_VPWR_c_725_n N_X_c_872_n 0.00730901f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_492 N_VPWR_M1017_s N_X_c_838_n 0.00176773f $X=6.775 $Y=1.835 $X2=0 $Y2=0
cc_493 N_VPWR_c_730_n N_X_c_838_n 0.0171443f $X=6.915 $Y=2.18 $X2=0 $Y2=0
cc_494 N_VPWR_c_736_n N_X_c_876_n 0.0124525f $X=7.61 $Y=3.33 $X2=0 $Y2=0
cc_495 N_VPWR_c_725_n N_X_c_876_n 0.00730901f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_496 N_VPWR_M1026_s N_X_c_840_n 2.39967e-19 $X=7.635 $Y=1.835 $X2=0 $Y2=0
cc_497 N_VPWR_c_732_n N_X_c_840_n 0.00347709f $X=7.775 $Y=2.19 $X2=0 $Y2=0
cc_498 N_VPWR_M1026_s N_X_c_842_n 0.00252087f $X=7.635 $Y=1.835 $X2=0 $Y2=0
cc_499 N_VPWR_c_732_n N_X_c_842_n 0.0194858f $X=7.775 $Y=2.19 $X2=0 $Y2=0
cc_500 N_X_c_832_n N_VGND_M1008_d 0.00176461f $X=7.25 $Y=1.15 $X2=0 $Y2=0
cc_501 N_X_c_834_n N_VGND_M1027_d 2.33864e-19 $X=7.715 $Y=1.15 $X2=0 $Y2=0
cc_502 N_X_c_836_n N_VGND_M1027_d 0.0020943f $X=7.895 $Y=1.235 $X2=0 $Y2=0
cc_503 N_X_c_832_n N_VGND_c_899_n 0.0170777f $X=7.25 $Y=1.15 $X2=0 $Y2=0
cc_504 N_X_c_834_n N_VGND_c_901_n 0.00362085f $X=7.715 $Y=1.15 $X2=0 $Y2=0
cc_505 N_X_c_836_n N_VGND_c_901_n 0.0203341f $X=7.895 $Y=1.235 $X2=0 $Y2=0
cc_506 N_X_c_888_p N_VGND_c_906_n 0.0124525f $X=6.485 $Y=0.42 $X2=0 $Y2=0
cc_507 N_X_c_889_p N_VGND_c_907_n 0.0124525f $X=7.345 $Y=0.42 $X2=0 $Y2=0
cc_508 N_X_M1007_s N_VGND_c_914_n 0.00536646f $X=6.345 $Y=0.235 $X2=0 $Y2=0
cc_509 N_X_M1019_s N_VGND_c_914_n 0.00536646f $X=7.205 $Y=0.235 $X2=0 $Y2=0
cc_510 N_X_c_888_p N_VGND_c_914_n 0.00730901f $X=6.485 $Y=0.42 $X2=0 $Y2=0
cc_511 N_X_c_889_p N_VGND_c_914_n 0.00730901f $X=7.345 $Y=0.42 $X2=0 $Y2=0
cc_512 N_VGND_c_914_n N_A_813_47#_M1003_s 0.00225186f $X=7.92 $Y=0 $X2=-0.19
+ $Y2=-0.245
cc_513 N_VGND_c_914_n N_A_813_47#_M1010_d 0.00403208f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_514 N_VGND_M1010_s N_A_813_47#_c_1014_n 0.00741677f $X=5.05 $Y=0.235 $X2=0
+ $Y2=0
cc_515 N_VGND_c_897_n N_A_813_47#_c_1014_n 0.0219934f $X=5.195 $Y=0.465 $X2=0
+ $Y2=0
cc_516 N_VGND_c_904_n N_A_813_47#_c_1014_n 0.00250018f $X=5.03 $Y=0 $X2=0 $Y2=0
cc_517 N_VGND_c_905_n N_A_813_47#_c_1014_n 0.0019105f $X=5.89 $Y=0 $X2=0 $Y2=0
cc_518 N_VGND_c_914_n N_A_813_47#_c_1014_n 0.00962135f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_519 N_VGND_c_905_n N_A_813_47#_c_1041_n 0.0124525f $X=5.89 $Y=0 $X2=0 $Y2=0
cc_520 N_VGND_c_914_n N_A_813_47#_c_1041_n 0.00730901f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_521 N_VGND_c_914_n N_A_813_47#_c_1016_n 0.00325124f $X=7.92 $Y=0 $X2=0 $Y2=0
cc_522 N_VGND_c_904_n N_A_813_47#_c_1015_n 0.00116529f $X=5.03 $Y=0 $X2=0 $Y2=0
