* NGSPICE file created from sky130_fd_sc_lp__a22oi_lp.ext - technology: sky130A

.subckt sky130_fd_sc_lp__a22oi_lp A1 A2 B1 B2 VGND VNB VPB VPWR Y
M1000 a_357_47# A1 Y VNB nshort w=420000u l=150000u
+  ad=1.764e+11p pd=1.68e+06u as=1.638e+11p ps=1.62e+06u
M1001 a_64_409# A2 VPWR VPB phighvt w=1e+06u l=250000u
+  ad=8.5e+11p pd=7.7e+06u as=2.9e+11p ps=2.58e+06u
M1002 a_64_409# B1 Y VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=2.8e+11p ps=2.56e+06u
M1003 VGND A2 a_357_47# VNB nshort w=420000u l=150000u
+  ad=2.394e+11p pd=2.82e+06u as=0p ps=0u
M1004 Y B2 a_64_409# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_171_47# B2 VGND VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1006 VPWR A1 a_64_409# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1007 Y B1 a_171_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

