* File: sky130_fd_sc_lp__dlxtp_lp.pxi.spice
* Created: Wed Sep  2 09:48:58 2020
* 
x_PM_SKY130_FD_SC_LP__DLXTP_LP%GATE N_GATE_M1010_g N_GATE_M1022_g N_GATE_M1001_g
+ N_GATE_M1000_g GATE GATE N_GATE_c_146_n PM_SKY130_FD_SC_LP__DLXTP_LP%GATE
x_PM_SKY130_FD_SC_LP__DLXTP_LP%D N_D_M1012_g N_D_M1019_g N_D_M1020_g N_D_M1017_g
+ D N_D_c_188_n N_D_c_189_n PM_SKY130_FD_SC_LP__DLXTP_LP%D
x_PM_SKY130_FD_SC_LP__DLXTP_LP%A_27_102# N_A_27_102#_M1010_s N_A_27_102#_M1022_s
+ N_A_27_102#_c_228_n N_A_27_102#_M1021_g N_A_27_102#_c_230_n
+ N_A_27_102#_M1003_g N_A_27_102#_M1024_g N_A_27_102#_M1002_g
+ N_A_27_102#_M1016_g N_A_27_102#_c_233_n N_A_27_102#_M1009_g
+ N_A_27_102#_c_235_n N_A_27_102#_c_236_n N_A_27_102#_c_237_n
+ N_A_27_102#_c_238_n N_A_27_102#_c_239_n N_A_27_102#_c_240_n
+ N_A_27_102#_c_241_n N_A_27_102#_c_242_n N_A_27_102#_c_243_n
+ N_A_27_102#_c_244_n N_A_27_102#_c_245_n N_A_27_102#_c_246_n
+ N_A_27_102#_c_247_n PM_SKY130_FD_SC_LP__DLXTP_LP%A_27_102#
x_PM_SKY130_FD_SC_LP__DLXTP_LP%A_350_102# N_A_350_102#_M1020_d
+ N_A_350_102#_M1017_d N_A_350_102#_M1014_g N_A_350_102#_M1023_g
+ N_A_350_102#_c_383_n N_A_350_102#_c_390_n N_A_350_102#_c_384_n
+ N_A_350_102#_c_385_n N_A_350_102#_c_391_n N_A_350_102#_c_392_n
+ N_A_350_102#_c_393_n N_A_350_102#_c_394_n N_A_350_102#_c_395_n
+ N_A_350_102#_c_386_n N_A_350_102#_c_387_n N_A_350_102#_c_388_n
+ PM_SKY130_FD_SC_LP__DLXTP_LP%A_350_102#
x_PM_SKY130_FD_SC_LP__DLXTP_LP%A_463_491# N_A_463_491#_M1003_s
+ N_A_463_491#_M1021_s N_A_463_491#_M1004_g N_A_463_491#_M1008_g
+ N_A_463_491#_c_491_n N_A_463_491#_c_484_n N_A_463_491#_c_492_n
+ N_A_463_491#_c_493_n N_A_463_491#_c_485_n N_A_463_491#_c_486_n
+ N_A_463_491#_c_487_n N_A_463_491#_c_488_n N_A_463_491#_c_494_n
+ N_A_463_491#_c_495_n N_A_463_491#_c_489_n
+ PM_SKY130_FD_SC_LP__DLXTP_LP%A_463_491#
x_PM_SKY130_FD_SC_LP__DLXTP_LP%A_1027_407# N_A_1027_407#_M1026_d
+ N_A_1027_407#_M1013_d N_A_1027_407#_M1027_g N_A_1027_407#_M1005_g
+ N_A_1027_407#_M1015_g N_A_1027_407#_M1006_g N_A_1027_407#_M1018_g
+ N_A_1027_407#_M1007_g N_A_1027_407#_c_600_n N_A_1027_407#_c_615_n
+ N_A_1027_407#_c_601_n N_A_1027_407#_c_602_n N_A_1027_407#_c_603_n
+ N_A_1027_407#_c_604_n N_A_1027_407#_c_605_n N_A_1027_407#_c_606_n
+ N_A_1027_407#_c_607_n N_A_1027_407#_c_608_n N_A_1027_407#_c_609_n
+ N_A_1027_407#_c_610_n PM_SKY130_FD_SC_LP__DLXTP_LP%A_1027_407#
x_PM_SKY130_FD_SC_LP__DLXTP_LP%A_824_491# N_A_824_491#_M1004_d
+ N_A_824_491#_M1016_d N_A_824_491#_M1025_g N_A_824_491#_M1011_g
+ N_A_824_491#_M1026_g N_A_824_491#_M1013_g N_A_824_491#_c_719_n
+ N_A_824_491#_c_709_n N_A_824_491#_c_710_n N_A_824_491#_c_711_n
+ N_A_824_491#_c_712_n N_A_824_491#_c_713_n N_A_824_491#_c_714_n
+ N_A_824_491#_c_715_n PM_SKY130_FD_SC_LP__DLXTP_LP%A_824_491#
x_PM_SKY130_FD_SC_LP__DLXTP_LP%VPWR N_VPWR_M1000_d N_VPWR_M1024_d N_VPWR_M1027_d
+ N_VPWR_M1006_s N_VPWR_c_807_n N_VPWR_c_808_n N_VPWR_c_809_n N_VPWR_c_810_n
+ N_VPWR_c_811_n N_VPWR_c_812_n N_VPWR_c_813_n N_VPWR_c_814_n VPWR
+ N_VPWR_c_815_n N_VPWR_c_816_n N_VPWR_c_817_n N_VPWR_c_806_n N_VPWR_c_819_n
+ N_VPWR_c_820_n PM_SKY130_FD_SC_LP__DLXTP_LP%VPWR
x_PM_SKY130_FD_SC_LP__DLXTP_LP%Q N_Q_M1018_d N_Q_M1007_d Q Q Q Q Q Q Q
+ N_Q_c_910_n PM_SKY130_FD_SC_LP__DLXTP_LP%Q
x_PM_SKY130_FD_SC_LP__DLXTP_LP%VGND N_VGND_M1001_d N_VGND_M1002_d N_VGND_M1005_d
+ N_VGND_M1015_s N_VGND_c_925_n N_VGND_c_926_n N_VGND_c_927_n N_VGND_c_928_n
+ VGND N_VGND_c_929_n N_VGND_c_930_n N_VGND_c_931_n N_VGND_c_932_n
+ N_VGND_c_933_n N_VGND_c_934_n N_VGND_c_935_n N_VGND_c_936_n N_VGND_c_937_n
+ N_VGND_c_938_n PM_SKY130_FD_SC_LP__DLXTP_LP%VGND
cc_1 VNB N_GATE_M1010_g 0.0442009f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.72
cc_2 VNB N_GATE_M1001_g 0.0359725f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=0.72
cc_3 VNB GATE 2.87194e-19 $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_4 VNB N_GATE_c_146_n 0.0193702f $X=-0.19 $Y=-0.245 $X2=0.74 $Y2=1.645
cc_5 VNB N_D_M1012_g 0.0442646f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.72
cc_6 VNB N_D_M1020_g 0.0602997f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=0.72
cc_7 VNB N_A_27_102#_c_228_n 0.0189958f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_27_102#_M1021_g 0.00577161f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=0.72
cc_9 VNB N_A_27_102#_c_230_n 0.0127219f $X=-0.19 $Y=-0.245 $X2=0.885 $Y2=2.15
cc_10 VNB N_A_27_102#_M1003_g 0.0377378f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_11 VNB N_A_27_102#_M1002_g 0.0506486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_27_102#_c_233_n 0.0161071f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_27_102#_M1009_g 0.0590464f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_27_102#_c_235_n 0.0191471f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_27_102#_c_236_n 0.00664034f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_27_102#_c_237_n 0.0283939f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_27_102#_c_238_n 0.0179711f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_27_102#_c_239_n 0.0191533f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_27_102#_c_240_n 0.0302601f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_27_102#_c_241_n 0.00475157f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_27_102#_c_242_n 0.00994965f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_27_102#_c_243_n 0.0101082f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_27_102#_c_244_n 8.41671e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_27_102#_c_245_n 0.00841726f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_27_102#_c_246_n 0.0154976f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_27_102#_c_247_n 0.0089424f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_350_102#_M1023_g 0.0343652f $X=-0.19 $Y=-0.245 $X2=0.885 $Y2=2.67
cc_28 VNB N_A_350_102#_c_383_n 0.0155104f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_350_102#_c_384_n 0.0331502f $X=-0.19 $Y=-0.245 $X2=0.74 $Y2=2.035
cc_30 VNB N_A_350_102#_c_385_n 0.00370651f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_350_102#_c_386_n 0.00399298f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_350_102#_c_387_n 0.0181743f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_350_102#_c_388_n 0.0414637f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_463_491#_M1004_g 0.0218328f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=1.48
cc_35 VNB N_A_463_491#_c_484_n 0.0122385f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_463_491#_c_485_n 0.0227043f $X=-0.19 $Y=-0.245 $X2=0.74 $Y2=1.645
cc_37 VNB N_A_463_491#_c_486_n 0.00541394f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_463_491#_c_487_n 0.0136679f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_463_491#_c_488_n 0.0306837f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_463_491#_c_489_n 0.0126855f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_1027_407#_M1005_g 0.0275732f $X=-0.19 $Y=-0.245 $X2=0.885 $Y2=2.15
cc_42 VNB N_A_1027_407#_M1015_g 0.0238669f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_1027_407#_M1006_g 0.0011252f $X=-0.19 $Y=-0.245 $X2=0.74 $Y2=1.645
cc_44 VNB N_A_1027_407#_M1018_g 0.0249073f $X=-0.19 $Y=-0.245 $X2=0.74 $Y2=2.035
cc_45 VNB N_A_1027_407#_M1007_g 0.00112085f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_1027_407#_c_600_n 0.0219019f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_1027_407#_c_601_n 0.00908276f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_1027_407#_c_602_n 0.00597105f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_1027_407#_c_603_n 0.00376039f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_1027_407#_c_604_n 3.5996e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_1027_407#_c_605_n 0.0264113f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_1027_407#_c_606_n 0.00360454f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_1027_407#_c_607_n 0.0340419f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_1027_407#_c_608_n 0.00160334f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_1027_407#_c_609_n 0.0015257f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_1027_407#_c_610_n 0.041805f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_824_491#_M1025_g 0.022059f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=1.48
cc_58 VNB N_A_824_491#_M1011_g 0.00286875f $X=-0.19 $Y=-0.245 $X2=0.885 $Y2=2.15
cc_59 VNB N_A_824_491#_M1026_g 0.0249238f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_60 VNB N_A_824_491#_M1013_g 0.00286199f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=1.645
cc_61 VNB N_A_824_491#_c_709_n 0.00633431f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_A_824_491#_c_710_n 6.36335e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_A_824_491#_c_711_n 0.018411f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_A_824_491#_c_712_n 0.0122908f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_A_824_491#_c_713_n 0.00716838f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_A_824_491#_c_714_n 0.00197566f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_A_824_491#_c_715_n 0.0398646f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_VPWR_c_806_n 0.342803f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_Q_c_910_n 0.0567461f $X=-0.19 $Y=-0.245 $X2=0.74 $Y2=1.645
cc_70 VNB N_VGND_c_925_n 0.0212986f $X=-0.19 $Y=-0.245 $X2=0.885 $Y2=2.67
cc_71 VNB N_VGND_c_926_n 0.00284591f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_VGND_c_927_n 0.00544418f $X=-0.19 $Y=-0.245 $X2=0.74 $Y2=1.645
cc_73 VNB N_VGND_c_928_n 0.0142982f $X=-0.19 $Y=-0.245 $X2=0.74 $Y2=2.035
cc_74 VNB N_VGND_c_929_n 0.0289964f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_VGND_c_930_n 0.0572732f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_VGND_c_931_n 0.0453151f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_VGND_c_932_n 0.0384381f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_VGND_c_933_n 0.0273851f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_VGND_c_934_n 0.46053f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_VGND_c_935_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_VGND_c_936_n 0.00510584f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_VGND_c_937_n 0.0051639f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_VGND_c_938_n 0.00536178f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VPB N_GATE_M1022_g 0.0247511f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=2.67
cc_85 VPB N_GATE_M1000_g 0.0206145f $X=-0.19 $Y=1.655 $X2=0.885 $Y2=2.67
cc_86 VPB GATE 0.00243924f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_87 VPB N_GATE_c_146_n 0.0517849f $X=-0.19 $Y=1.655 $X2=0.74 $Y2=1.645
cc_88 VPB N_D_M1012_g 0.00810144f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=0.72
cc_89 VPB N_D_M1019_g 0.0201757f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=2.67
cc_90 VPB N_D_M1020_g 0.0126995f $X=-0.19 $Y=1.655 $X2=0.855 $Y2=0.72
cc_91 VPB N_D_M1017_g 0.0236641f $X=-0.19 $Y=1.655 $X2=0.885 $Y2=2.67
cc_92 VPB N_D_c_188_n 0.00579238f $X=-0.19 $Y=1.655 $X2=0.74 $Y2=1.645
cc_93 VPB N_D_c_189_n 0.0368333f $X=-0.19 $Y=1.655 $X2=0.74 $Y2=1.645
cc_94 VPB N_A_27_102#_M1021_g 0.0663648f $X=-0.19 $Y=1.655 $X2=0.855 $Y2=0.72
cc_95 VPB N_A_27_102#_M1024_g 0.046589f $X=-0.19 $Y=1.655 $X2=0.69 $Y2=1.645
cc_96 VPB N_A_27_102#_M1016_g 0.0385009f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_97 VPB N_A_27_102#_c_233_n 0.0285496f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_98 VPB N_A_27_102#_c_238_n 0.0629748f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_99 VPB N_A_27_102#_c_241_n 0.00930159f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_100 VPB N_A_27_102#_c_244_n 0.00177921f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_101 VPB N_A_27_102#_c_245_n 0.00262429f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_102 VPB N_A_27_102#_c_246_n 0.0112639f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_103 VPB N_A_27_102#_c_247_n 0.0257619f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_104 VPB N_A_350_102#_M1014_g 0.0205209f $X=-0.19 $Y=1.655 $X2=0.855 $Y2=0.72
cc_105 VPB N_A_350_102#_c_390_n 0.0148954f $X=-0.19 $Y=1.655 $X2=0.74 $Y2=1.645
cc_106 VPB N_A_350_102#_c_391_n 0.0309098f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_107 VPB N_A_350_102#_c_392_n 0.00448003f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_108 VPB N_A_350_102#_c_393_n 0.00525711f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_109 VPB N_A_350_102#_c_394_n 0.00341323f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_110 VPB N_A_350_102#_c_395_n 0.0326084f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_111 VPB N_A_350_102#_c_387_n 0.0158483f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_112 VPB N_A_463_491#_M1008_g 0.020863f $X=-0.19 $Y=1.655 $X2=0.885 $Y2=2.15
cc_113 VPB N_A_463_491#_c_491_n 0.00425587f $X=-0.19 $Y=1.655 $X2=0.885 $Y2=2.67
cc_114 VPB N_A_463_491#_c_492_n 0.00137094f $X=-0.19 $Y=1.655 $X2=0.74 $Y2=1.645
cc_115 VPB N_A_463_491#_c_493_n 0.00554693f $X=-0.19 $Y=1.655 $X2=0.74 $Y2=1.645
cc_116 VPB N_A_463_491#_c_494_n 0.010704f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_117 VPB N_A_463_491#_c_495_n 0.0380297f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_118 VPB N_A_463_491#_c_489_n 0.00764203f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_119 VPB N_A_1027_407#_M1027_g 0.0411095f $X=-0.19 $Y=1.655 $X2=0.855 $Y2=1.48
cc_120 VPB N_A_1027_407#_M1006_g 0.0226588f $X=-0.19 $Y=1.655 $X2=0.74 $Y2=1.645
cc_121 VPB N_A_1027_407#_M1007_g 0.0234886f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_122 VPB N_A_1027_407#_c_600_n 0.025078f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_123 VPB N_A_1027_407#_c_615_n 0.0123193f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_124 VPB N_A_1027_407#_c_604_n 0.0143086f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_125 VPB N_A_824_491#_M1011_g 0.0215593f $X=-0.19 $Y=1.655 $X2=0.885 $Y2=2.15
cc_126 VPB N_A_824_491#_M1013_g 0.0234886f $X=-0.19 $Y=1.655 $X2=0.69 $Y2=1.645
cc_127 VPB N_A_824_491#_c_710_n 0.00986511f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_128 VPB N_VPWR_c_807_n 0.00976748f $X=-0.19 $Y=1.655 $X2=0.885 $Y2=2.67
cc_129 VPB N_VPWR_c_808_n 0.0051887f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_130 VPB N_VPWR_c_809_n 0.0133431f $X=-0.19 $Y=1.655 $X2=0.74 $Y2=1.645
cc_131 VPB N_VPWR_c_810_n 0.017248f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_132 VPB N_VPWR_c_811_n 0.0529526f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_133 VPB N_VPWR_c_812_n 0.00631679f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_134 VPB N_VPWR_c_813_n 0.052568f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_135 VPB N_VPWR_c_814_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_136 VPB N_VPWR_c_815_n 0.0294867f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_137 VPB N_VPWR_c_816_n 0.028322f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_138 VPB N_VPWR_c_817_n 0.0271876f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_139 VPB N_VPWR_c_806_n 0.0918341f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_140 VPB N_VPWR_c_819_n 0.00565027f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_141 VPB N_VPWR_c_820_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_142 VPB N_Q_c_910_n 0.0543794f $X=-0.19 $Y=1.655 $X2=0.74 $Y2=1.645
cc_143 N_GATE_M1001_g N_D_M1012_g 0.0287144f $X=0.855 $Y=0.72 $X2=0 $Y2=0
cc_144 GATE N_D_M1012_g 0.00164079f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_145 N_GATE_c_146_n N_D_M1012_g 0.0234541f $X=0.74 $Y=1.645 $X2=0 $Y2=0
cc_146 GATE N_D_c_188_n 0.0258926f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_147 N_GATE_c_146_n N_D_c_188_n 0.00267572f $X=0.74 $Y=1.645 $X2=0 $Y2=0
cc_148 N_GATE_M1000_g N_D_c_189_n 0.0234541f $X=0.885 $Y=2.67 $X2=0 $Y2=0
cc_149 GATE N_D_c_189_n 2.94447e-19 $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_150 N_GATE_M1010_g N_A_27_102#_c_237_n 0.0157852f $X=0.495 $Y=0.72 $X2=0
+ $Y2=0
cc_151 N_GATE_M1001_g N_A_27_102#_c_237_n 0.00215172f $X=0.855 $Y=0.72 $X2=0
+ $Y2=0
cc_152 N_GATE_M1010_g N_A_27_102#_c_238_n 0.0353151f $X=0.495 $Y=0.72 $X2=0
+ $Y2=0
cc_153 GATE N_A_27_102#_c_238_n 0.0442702f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_154 N_GATE_M1010_g N_A_27_102#_c_239_n 0.0144626f $X=0.495 $Y=0.72 $X2=0
+ $Y2=0
cc_155 N_GATE_M1001_g N_A_27_102#_c_239_n 0.0147236f $X=0.855 $Y=0.72 $X2=0
+ $Y2=0
cc_156 GATE N_A_27_102#_c_239_n 0.0246023f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_157 N_GATE_c_146_n N_A_27_102#_c_239_n 0.0014382f $X=0.74 $Y=1.645 $X2=0
+ $Y2=0
cc_158 N_GATE_M1010_g N_A_27_102#_c_242_n 0.00513266f $X=0.495 $Y=0.72 $X2=0
+ $Y2=0
cc_159 N_GATE_M1001_g N_A_27_102#_c_243_n 9.36765e-19 $X=0.855 $Y=0.72 $X2=0
+ $Y2=0
cc_160 GATE N_A_27_102#_c_243_n 0.00359454f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_161 N_GATE_c_146_n N_A_27_102#_c_243_n 4.07611e-19 $X=0.74 $Y=1.645 $X2=0
+ $Y2=0
cc_162 N_GATE_M1022_g N_VPWR_c_807_n 0.0026553f $X=0.495 $Y=2.67 $X2=0 $Y2=0
cc_163 N_GATE_M1000_g N_VPWR_c_807_n 0.0176964f $X=0.885 $Y=2.67 $X2=0 $Y2=0
cc_164 N_GATE_M1022_g N_VPWR_c_815_n 0.00486513f $X=0.495 $Y=2.67 $X2=0 $Y2=0
cc_165 N_GATE_M1000_g N_VPWR_c_815_n 0.0040395f $X=0.885 $Y=2.67 $X2=0 $Y2=0
cc_166 N_GATE_M1022_g N_VPWR_c_806_n 0.00986222f $X=0.495 $Y=2.67 $X2=0 $Y2=0
cc_167 N_GATE_M1000_g N_VPWR_c_806_n 0.00774838f $X=0.885 $Y=2.67 $X2=0 $Y2=0
cc_168 N_GATE_M1010_g N_VGND_c_925_n 0.00180376f $X=0.495 $Y=0.72 $X2=0 $Y2=0
cc_169 N_GATE_M1001_g N_VGND_c_925_n 0.0121401f $X=0.855 $Y=0.72 $X2=0 $Y2=0
cc_170 N_GATE_M1010_g N_VGND_c_929_n 0.00461605f $X=0.495 $Y=0.72 $X2=0 $Y2=0
cc_171 N_GATE_M1001_g N_VGND_c_929_n 0.00400048f $X=0.855 $Y=0.72 $X2=0 $Y2=0
cc_172 N_GATE_M1010_g N_VGND_c_934_n 0.00502397f $X=0.495 $Y=0.72 $X2=0 $Y2=0
cc_173 N_GATE_M1001_g N_VGND_c_934_n 0.00422014f $X=0.855 $Y=0.72 $X2=0 $Y2=0
cc_174 N_D_M1012_g N_A_27_102#_c_239_n 0.0142937f $X=1.315 $Y=0.72 $X2=0 $Y2=0
cc_175 N_D_c_188_n N_A_27_102#_c_239_n 0.0095317f $X=1.435 $Y=1.985 $X2=0 $Y2=0
cc_176 N_D_M1020_g N_A_27_102#_c_240_n 0.0194362f $X=1.675 $Y=0.72 $X2=0 $Y2=0
cc_177 N_D_c_188_n N_A_27_102#_c_240_n 0.0033518f $X=1.435 $Y=1.985 $X2=0 $Y2=0
cc_178 N_D_M1012_g N_A_27_102#_c_243_n 0.0091938f $X=1.315 $Y=0.72 $X2=0 $Y2=0
cc_179 N_D_M1020_g N_A_27_102#_c_243_n 0.00511336f $X=1.675 $Y=0.72 $X2=0 $Y2=0
cc_180 N_D_c_188_n N_A_27_102#_c_243_n 0.0110721f $X=1.435 $Y=1.985 $X2=0 $Y2=0
cc_181 N_D_c_189_n N_A_27_102#_c_243_n 6.68747e-19 $X=1.675 $Y=1.985 $X2=0 $Y2=0
cc_182 N_D_M1012_g N_A_350_102#_c_383_n 0.00189708f $X=1.315 $Y=0.72 $X2=0 $Y2=0
cc_183 N_D_M1020_g N_A_350_102#_c_383_n 0.0139544f $X=1.675 $Y=0.72 $X2=0 $Y2=0
cc_184 N_D_M1019_g N_A_350_102#_c_390_n 0.00185f $X=1.315 $Y=2.67 $X2=0 $Y2=0
cc_185 N_D_M1017_g N_A_350_102#_c_390_n 0.0130453f $X=1.675 $Y=2.67 $X2=0 $Y2=0
cc_186 N_D_M1012_g N_A_350_102#_c_385_n 3.6289e-19 $X=1.315 $Y=0.72 $X2=0 $Y2=0
cc_187 N_D_M1020_g N_A_350_102#_c_385_n 0.00668379f $X=1.675 $Y=0.72 $X2=0 $Y2=0
cc_188 N_D_c_188_n N_A_350_102#_c_392_n 0.0100803f $X=1.435 $Y=1.985 $X2=0 $Y2=0
cc_189 N_D_c_189_n N_A_350_102#_c_392_n 0.00483418f $X=1.675 $Y=1.985 $X2=0
+ $Y2=0
cc_190 N_D_c_188_n N_A_350_102#_c_393_n 7.15467e-19 $X=1.435 $Y=1.985 $X2=0
+ $Y2=0
cc_191 N_D_c_189_n N_A_350_102#_c_393_n 0.00677995f $X=1.675 $Y=1.985 $X2=0
+ $Y2=0
cc_192 N_D_M1017_g N_A_463_491#_c_491_n 0.00206871f $X=1.675 $Y=2.67 $X2=0 $Y2=0
cc_193 N_D_M1019_g N_VPWR_c_807_n 0.0154529f $X=1.315 $Y=2.67 $X2=0 $Y2=0
cc_194 N_D_M1017_g N_VPWR_c_807_n 0.00252244f $X=1.675 $Y=2.67 $X2=0 $Y2=0
cc_195 N_D_c_188_n N_VPWR_c_807_n 0.0149963f $X=1.435 $Y=1.985 $X2=0 $Y2=0
cc_196 N_D_M1019_g N_VPWR_c_811_n 0.0040395f $X=1.315 $Y=2.67 $X2=0 $Y2=0
cc_197 N_D_M1017_g N_VPWR_c_811_n 0.00457319f $X=1.675 $Y=2.67 $X2=0 $Y2=0
cc_198 N_D_M1019_g N_VPWR_c_806_n 0.00772493f $X=1.315 $Y=2.67 $X2=0 $Y2=0
cc_199 N_D_M1017_g N_VPWR_c_806_n 0.00904779f $X=1.675 $Y=2.67 $X2=0 $Y2=0
cc_200 N_D_M1012_g N_VGND_c_925_n 0.00392072f $X=1.315 $Y=0.72 $X2=0 $Y2=0
cc_201 N_D_M1012_g N_VGND_c_930_n 0.00481372f $X=1.315 $Y=0.72 $X2=0 $Y2=0
cc_202 N_D_M1020_g N_VGND_c_930_n 0.00461605f $X=1.675 $Y=0.72 $X2=0 $Y2=0
cc_203 N_D_M1012_g N_VGND_c_934_n 0.00502397f $X=1.315 $Y=0.72 $X2=0 $Y2=0
cc_204 N_D_M1020_g N_VGND_c_934_n 0.00502397f $X=1.675 $Y=0.72 $X2=0 $Y2=0
cc_205 N_A_27_102#_M1024_g N_A_350_102#_M1014_g 0.0249456f $X=3.065 $Y=2.775
+ $X2=0 $Y2=0
cc_206 N_A_27_102#_M1002_g N_A_350_102#_M1023_g 0.0193708f $X=3.235 $Y=0.445
+ $X2=0 $Y2=0
cc_207 N_A_27_102#_c_235_n N_A_350_102#_c_383_n 0.00107574f $X=2.845 $Y=1.11
+ $X2=0 $Y2=0
cc_208 N_A_27_102#_M1021_g N_A_350_102#_c_390_n 0.00141583f $X=2.675 $Y=2.775
+ $X2=0 $Y2=0
cc_209 N_A_27_102#_c_228_n N_A_350_102#_c_384_n 0.00525722f $X=2.675 $Y=1.425
+ $X2=0 $Y2=0
cc_210 N_A_27_102#_c_230_n N_A_350_102#_c_384_n 0.00156877f $X=2.98 $Y=1.5 $X2=0
+ $Y2=0
cc_211 N_A_27_102#_M1002_g N_A_350_102#_c_384_n 0.0103673f $X=3.235 $Y=0.445
+ $X2=0 $Y2=0
cc_212 N_A_27_102#_c_235_n N_A_350_102#_c_384_n 0.0119583f $X=2.845 $Y=1.11
+ $X2=0 $Y2=0
cc_213 N_A_27_102#_c_240_n N_A_350_102#_c_384_n 0.0647901f $X=2.98 $Y=1.51 $X2=0
+ $Y2=0
cc_214 N_A_27_102#_c_241_n N_A_350_102#_c_384_n 0.0111886f $X=3.94 $Y=1.67 $X2=0
+ $Y2=0
cc_215 N_A_27_102#_c_244_n N_A_350_102#_c_384_n 0.0231617f $X=3.145 $Y=1.51
+ $X2=0 $Y2=0
cc_216 N_A_27_102#_c_246_n N_A_350_102#_c_384_n 6.12359e-19 $X=3.145 $Y=1.5
+ $X2=0 $Y2=0
cc_217 N_A_27_102#_c_240_n N_A_350_102#_c_385_n 0.0265557f $X=2.98 $Y=1.51 $X2=0
+ $Y2=0
cc_218 N_A_27_102#_c_243_n N_A_350_102#_c_385_n 0.00879787f $X=1.46 $Y=1.215
+ $X2=0 $Y2=0
cc_219 N_A_27_102#_M1021_g N_A_350_102#_c_391_n 0.0141952f $X=2.675 $Y=2.775
+ $X2=0 $Y2=0
cc_220 N_A_27_102#_c_230_n N_A_350_102#_c_391_n 0.00131698f $X=2.98 $Y=1.5 $X2=0
+ $Y2=0
cc_221 N_A_27_102#_M1024_g N_A_350_102#_c_391_n 0.0112421f $X=3.065 $Y=2.775
+ $X2=0 $Y2=0
cc_222 N_A_27_102#_c_240_n N_A_350_102#_c_391_n 0.039512f $X=2.98 $Y=1.51 $X2=0
+ $Y2=0
cc_223 N_A_27_102#_c_241_n N_A_350_102#_c_391_n 0.0058444f $X=3.94 $Y=1.67 $X2=0
+ $Y2=0
cc_224 N_A_27_102#_c_244_n N_A_350_102#_c_391_n 0.0205475f $X=3.145 $Y=1.51
+ $X2=0 $Y2=0
cc_225 N_A_27_102#_c_246_n N_A_350_102#_c_391_n 0.00118556f $X=3.145 $Y=1.5
+ $X2=0 $Y2=0
cc_226 N_A_27_102#_c_240_n N_A_350_102#_c_392_n 0.00836921f $X=2.98 $Y=1.51
+ $X2=0 $Y2=0
cc_227 N_A_27_102#_M1021_g N_A_350_102#_c_393_n 0.0071235f $X=2.675 $Y=2.775
+ $X2=0 $Y2=0
cc_228 N_A_27_102#_M1024_g N_A_350_102#_c_394_n 0.00113572f $X=3.065 $Y=2.775
+ $X2=0 $Y2=0
cc_229 N_A_27_102#_M1016_g N_A_350_102#_c_394_n 0.00207094f $X=4.045 $Y=2.775
+ $X2=0 $Y2=0
cc_230 N_A_27_102#_c_241_n N_A_350_102#_c_394_n 0.0205475f $X=3.94 $Y=1.67 $X2=0
+ $Y2=0
cc_231 N_A_27_102#_c_245_n N_A_350_102#_c_394_n 6.33735e-19 $X=4.105 $Y=1.67
+ $X2=0 $Y2=0
cc_232 N_A_27_102#_M1024_g N_A_350_102#_c_395_n 0.0166711f $X=3.065 $Y=2.775
+ $X2=0 $Y2=0
cc_233 N_A_27_102#_M1016_g N_A_350_102#_c_395_n 0.0695472f $X=4.045 $Y=2.775
+ $X2=0 $Y2=0
cc_234 N_A_27_102#_c_241_n N_A_350_102#_c_395_n 0.00111736f $X=3.94 $Y=1.67
+ $X2=0 $Y2=0
cc_235 N_A_27_102#_c_247_n N_A_350_102#_c_395_n 6.09406e-19 $X=4.105 $Y=1.72
+ $X2=0 $Y2=0
cc_236 N_A_27_102#_M1002_g N_A_350_102#_c_386_n 0.00115306f $X=3.235 $Y=0.445
+ $X2=0 $Y2=0
cc_237 N_A_27_102#_c_241_n N_A_350_102#_c_386_n 0.0231602f $X=3.94 $Y=1.67 $X2=0
+ $Y2=0
cc_238 N_A_27_102#_M1024_g N_A_350_102#_c_387_n 0.00751587f $X=3.065 $Y=2.775
+ $X2=0 $Y2=0
cc_239 N_A_27_102#_c_241_n N_A_350_102#_c_387_n 0.0107036f $X=3.94 $Y=1.67 $X2=0
+ $Y2=0
cc_240 N_A_27_102#_c_244_n N_A_350_102#_c_387_n 0.00115059f $X=3.145 $Y=1.51
+ $X2=0 $Y2=0
cc_241 N_A_27_102#_c_245_n N_A_350_102#_c_387_n 0.00167141f $X=4.105 $Y=1.67
+ $X2=0 $Y2=0
cc_242 N_A_27_102#_c_246_n N_A_350_102#_c_387_n 0.019203f $X=3.145 $Y=1.5 $X2=0
+ $Y2=0
cc_243 N_A_27_102#_c_247_n N_A_350_102#_c_387_n 0.0179314f $X=4.105 $Y=1.72
+ $X2=0 $Y2=0
cc_244 N_A_27_102#_M1002_g N_A_350_102#_c_388_n 0.019203f $X=3.235 $Y=0.445
+ $X2=0 $Y2=0
cc_245 N_A_27_102#_c_241_n N_A_350_102#_c_388_n 0.00365246f $X=3.94 $Y=1.67
+ $X2=0 $Y2=0
cc_246 N_A_27_102#_c_245_n N_A_350_102#_c_388_n 2.24039e-19 $X=4.105 $Y=1.67
+ $X2=0 $Y2=0
cc_247 N_A_27_102#_c_247_n N_A_350_102#_c_388_n 5.73335e-19 $X=4.105 $Y=1.72
+ $X2=0 $Y2=0
cc_248 N_A_27_102#_M1009_g N_A_463_491#_M1004_g 0.0140464f $X=4.835 $Y=0.445
+ $X2=0 $Y2=0
cc_249 N_A_27_102#_M1021_g N_A_463_491#_c_491_n 0.0101071f $X=2.675 $Y=2.775
+ $X2=0 $Y2=0
cc_250 N_A_27_102#_M1024_g N_A_463_491#_c_491_n 0.0015949f $X=3.065 $Y=2.775
+ $X2=0 $Y2=0
cc_251 N_A_27_102#_M1003_g N_A_463_491#_c_484_n 0.00960915f $X=2.845 $Y=0.445
+ $X2=0 $Y2=0
cc_252 N_A_27_102#_M1002_g N_A_463_491#_c_484_n 0.00168185f $X=3.235 $Y=0.445
+ $X2=0 $Y2=0
cc_253 N_A_27_102#_M1021_g N_A_463_491#_c_492_n 0.00919462f $X=2.675 $Y=2.775
+ $X2=0 $Y2=0
cc_254 N_A_27_102#_M1024_g N_A_463_491#_c_492_n 0.0134552f $X=3.065 $Y=2.775
+ $X2=0 $Y2=0
cc_255 N_A_27_102#_M1016_g N_A_463_491#_c_492_n 0.0134062f $X=4.045 $Y=2.775
+ $X2=0 $Y2=0
cc_256 N_A_27_102#_c_233_n N_A_463_491#_c_492_n 0.00363563f $X=4.76 $Y=1.72
+ $X2=0 $Y2=0
cc_257 N_A_27_102#_c_245_n N_A_463_491#_c_492_n 0.00887007f $X=4.105 $Y=1.67
+ $X2=0 $Y2=0
cc_258 N_A_27_102#_c_247_n N_A_463_491#_c_492_n 6.30355e-19 $X=4.105 $Y=1.72
+ $X2=0 $Y2=0
cc_259 N_A_27_102#_M1021_g N_A_463_491#_c_493_n 0.00400408f $X=2.675 $Y=2.775
+ $X2=0 $Y2=0
cc_260 N_A_27_102#_M1003_g N_A_463_491#_c_485_n 0.00854758f $X=2.845 $Y=0.445
+ $X2=0 $Y2=0
cc_261 N_A_27_102#_M1002_g N_A_463_491#_c_485_n 0.0126021f $X=3.235 $Y=0.445
+ $X2=0 $Y2=0
cc_262 N_A_27_102#_M1003_g N_A_463_491#_c_486_n 0.00419197f $X=2.845 $Y=0.445
+ $X2=0 $Y2=0
cc_263 N_A_27_102#_c_235_n N_A_463_491#_c_486_n 0.00466095f $X=2.845 $Y=1.11
+ $X2=0 $Y2=0
cc_264 N_A_27_102#_M1009_g N_A_463_491#_c_487_n 0.00250644f $X=4.835 $Y=0.445
+ $X2=0 $Y2=0
cc_265 N_A_27_102#_c_245_n N_A_463_491#_c_487_n 0.00753299f $X=4.105 $Y=1.67
+ $X2=0 $Y2=0
cc_266 N_A_27_102#_c_247_n N_A_463_491#_c_487_n 0.00159057f $X=4.105 $Y=1.72
+ $X2=0 $Y2=0
cc_267 N_A_27_102#_M1009_g N_A_463_491#_c_488_n 0.0163772f $X=4.835 $Y=0.445
+ $X2=0 $Y2=0
cc_268 N_A_27_102#_c_245_n N_A_463_491#_c_488_n 3.49744e-19 $X=4.105 $Y=1.67
+ $X2=0 $Y2=0
cc_269 N_A_27_102#_c_247_n N_A_463_491#_c_488_n 0.00724017f $X=4.105 $Y=1.72
+ $X2=0 $Y2=0
cc_270 N_A_27_102#_c_233_n N_A_463_491#_c_494_n 0.00157122f $X=4.76 $Y=1.72
+ $X2=0 $Y2=0
cc_271 N_A_27_102#_M1016_g N_A_463_491#_c_495_n 0.0258971f $X=4.045 $Y=2.775
+ $X2=0 $Y2=0
cc_272 N_A_27_102#_c_233_n N_A_463_491#_c_495_n 0.0109777f $X=4.76 $Y=1.72 $X2=0
+ $Y2=0
cc_273 N_A_27_102#_M1016_g N_A_463_491#_c_489_n 0.012319f $X=4.045 $Y=2.775
+ $X2=0 $Y2=0
cc_274 N_A_27_102#_c_233_n N_A_463_491#_c_489_n 0.0137693f $X=4.76 $Y=1.72 $X2=0
+ $Y2=0
cc_275 N_A_27_102#_M1009_g N_A_463_491#_c_489_n 0.00929147f $X=4.835 $Y=0.445
+ $X2=0 $Y2=0
cc_276 N_A_27_102#_c_245_n N_A_463_491#_c_489_n 0.0277591f $X=4.105 $Y=1.67
+ $X2=0 $Y2=0
cc_277 N_A_27_102#_c_247_n N_A_463_491#_c_489_n 0.00400978f $X=4.105 $Y=1.72
+ $X2=0 $Y2=0
cc_278 N_A_27_102#_M1009_g N_A_1027_407#_M1005_g 0.0438816f $X=4.835 $Y=0.445
+ $X2=0 $Y2=0
cc_279 N_A_27_102#_M1009_g N_A_1027_407#_c_606_n 3.77891e-19 $X=4.835 $Y=0.445
+ $X2=0 $Y2=0
cc_280 N_A_27_102#_c_233_n N_A_1027_407#_c_607_n 0.0438816f $X=4.76 $Y=1.72
+ $X2=0 $Y2=0
cc_281 N_A_27_102#_M1016_g N_A_824_491#_c_719_n 0.00431856f $X=4.045 $Y=2.775
+ $X2=0 $Y2=0
cc_282 N_A_27_102#_M1009_g N_A_824_491#_c_709_n 0.0173723f $X=4.835 $Y=0.445
+ $X2=0 $Y2=0
cc_283 N_A_27_102#_M1009_g N_A_824_491#_c_710_n 0.00174833f $X=4.835 $Y=0.445
+ $X2=0 $Y2=0
cc_284 N_A_27_102#_M1009_g N_A_824_491#_c_712_n 0.00718564f $X=4.835 $Y=0.445
+ $X2=0 $Y2=0
cc_285 N_A_27_102#_M1009_g N_A_824_491#_c_713_n 0.0118985f $X=4.835 $Y=0.445
+ $X2=0 $Y2=0
cc_286 N_A_27_102#_c_238_n N_VPWR_c_807_n 0.0100601f $X=0.28 $Y=2.495 $X2=0
+ $Y2=0
cc_287 N_A_27_102#_M1024_g N_VPWR_c_808_n 0.00479274f $X=3.065 $Y=2.775 $X2=0
+ $Y2=0
cc_288 N_A_27_102#_M1021_g N_VPWR_c_811_n 0.00421724f $X=2.675 $Y=2.775 $X2=0
+ $Y2=0
cc_289 N_A_27_102#_M1024_g N_VPWR_c_811_n 0.00432313f $X=3.065 $Y=2.775 $X2=0
+ $Y2=0
cc_290 N_A_27_102#_M1016_g N_VPWR_c_813_n 0.00421279f $X=4.045 $Y=2.775 $X2=0
+ $Y2=0
cc_291 N_A_27_102#_c_238_n N_VPWR_c_815_n 0.0125753f $X=0.28 $Y=2.495 $X2=0
+ $Y2=0
cc_292 N_A_27_102#_M1021_g N_VPWR_c_806_n 0.00729982f $X=2.675 $Y=2.775 $X2=0
+ $Y2=0
cc_293 N_A_27_102#_M1024_g N_VPWR_c_806_n 0.00629995f $X=3.065 $Y=2.775 $X2=0
+ $Y2=0
cc_294 N_A_27_102#_M1016_g N_VPWR_c_806_n 0.0061535f $X=4.045 $Y=2.775 $X2=0
+ $Y2=0
cc_295 N_A_27_102#_c_238_n N_VPWR_c_806_n 0.00932134f $X=0.28 $Y=2.495 $X2=0
+ $Y2=0
cc_296 N_A_27_102#_c_237_n N_VGND_c_925_n 0.0153904f $X=0.28 $Y=0.72 $X2=0 $Y2=0
cc_297 N_A_27_102#_c_239_n N_VGND_c_925_n 0.0264018f $X=1.375 $Y=1.215 $X2=0
+ $Y2=0
cc_298 N_A_27_102#_M1003_g N_VGND_c_926_n 0.00202904f $X=2.845 $Y=0.445 $X2=0
+ $Y2=0
cc_299 N_A_27_102#_M1002_g N_VGND_c_926_n 0.0106538f $X=3.235 $Y=0.445 $X2=0
+ $Y2=0
cc_300 N_A_27_102#_M1009_g N_VGND_c_927_n 0.00206354f $X=4.835 $Y=0.445 $X2=0
+ $Y2=0
cc_301 N_A_27_102#_c_237_n N_VGND_c_929_n 0.00925243f $X=0.28 $Y=0.72 $X2=0
+ $Y2=0
cc_302 N_A_27_102#_M1003_g N_VGND_c_930_n 0.00426341f $X=2.845 $Y=0.445 $X2=0
+ $Y2=0
cc_303 N_A_27_102#_M1002_g N_VGND_c_930_n 0.00364083f $X=3.235 $Y=0.445 $X2=0
+ $Y2=0
cc_304 N_A_27_102#_M1009_g N_VGND_c_931_n 0.00397065f $X=4.835 $Y=0.445 $X2=0
+ $Y2=0
cc_305 N_A_27_102#_M1003_g N_VGND_c_934_n 0.00738256f $X=2.845 $Y=0.445 $X2=0
+ $Y2=0
cc_306 N_A_27_102#_M1002_g N_VGND_c_934_n 0.0042609f $X=3.235 $Y=0.445 $X2=0
+ $Y2=0
cc_307 N_A_27_102#_M1009_g N_VGND_c_934_n 0.00594666f $X=4.835 $Y=0.445 $X2=0
+ $Y2=0
cc_308 N_A_27_102#_c_237_n N_VGND_c_934_n 0.0110254f $X=0.28 $Y=0.72 $X2=0 $Y2=0
cc_309 N_A_350_102#_M1023_g N_A_463_491#_M1004_g 0.0290094f $X=3.875 $Y=0.445
+ $X2=0 $Y2=0
cc_310 N_A_350_102#_c_390_n N_A_463_491#_c_491_n 0.0238622f $X=1.89 $Y=2.495
+ $X2=0 $Y2=0
cc_311 N_A_350_102#_c_383_n N_A_463_491#_c_484_n 0.01063f $X=1.89 $Y=0.72 $X2=0
+ $Y2=0
cc_312 N_A_350_102#_M1014_g N_A_463_491#_c_492_n 0.0125532f $X=3.655 $Y=2.775
+ $X2=0 $Y2=0
cc_313 N_A_350_102#_c_391_n N_A_463_491#_c_492_n 0.0295088f $X=3.4 $Y=2.05 $X2=0
+ $Y2=0
cc_314 N_A_350_102#_c_394_n N_A_463_491#_c_492_n 0.0209281f $X=3.565 $Y=2.05
+ $X2=0 $Y2=0
cc_315 N_A_350_102#_c_395_n N_A_463_491#_c_492_n 0.00111495f $X=3.565 $Y=2.13
+ $X2=0 $Y2=0
cc_316 N_A_350_102#_c_390_n N_A_463_491#_c_493_n 0.0144023f $X=1.89 $Y=2.495
+ $X2=0 $Y2=0
cc_317 N_A_350_102#_c_391_n N_A_463_491#_c_493_n 0.0184329f $X=3.4 $Y=2.05 $X2=0
+ $Y2=0
cc_318 N_A_350_102#_M1023_g N_A_463_491#_c_485_n 0.0148812f $X=3.875 $Y=0.445
+ $X2=0 $Y2=0
cc_319 N_A_350_102#_c_384_n N_A_463_491#_c_485_n 0.0524894f $X=3.55 $Y=1.16
+ $X2=0 $Y2=0
cc_320 N_A_350_102#_c_386_n N_A_463_491#_c_485_n 0.0234243f $X=3.715 $Y=1.16
+ $X2=0 $Y2=0
cc_321 N_A_350_102#_c_388_n N_A_463_491#_c_485_n 0.00172004f $X=3.875 $Y=1.24
+ $X2=0 $Y2=0
cc_322 N_A_350_102#_c_383_n N_A_463_491#_c_486_n 0.00816634f $X=1.89 $Y=0.72
+ $X2=0 $Y2=0
cc_323 N_A_350_102#_c_384_n N_A_463_491#_c_486_n 0.0257405f $X=3.55 $Y=1.16
+ $X2=0 $Y2=0
cc_324 N_A_350_102#_M1023_g N_A_463_491#_c_487_n 0.00546389f $X=3.875 $Y=0.445
+ $X2=0 $Y2=0
cc_325 N_A_350_102#_c_386_n N_A_463_491#_c_487_n 0.00734858f $X=3.715 $Y=1.16
+ $X2=0 $Y2=0
cc_326 N_A_350_102#_c_388_n N_A_463_491#_c_488_n 0.0290094f $X=3.875 $Y=1.24
+ $X2=0 $Y2=0
cc_327 N_A_350_102#_c_386_n N_A_463_491#_c_489_n 0.00660374f $X=3.715 $Y=1.16
+ $X2=0 $Y2=0
cc_328 N_A_350_102#_c_388_n N_A_463_491#_c_489_n 0.00406419f $X=3.875 $Y=1.24
+ $X2=0 $Y2=0
cc_329 N_A_350_102#_M1014_g N_A_824_491#_c_719_n 6.08765e-19 $X=3.655 $Y=2.775
+ $X2=0 $Y2=0
cc_330 N_A_350_102#_c_390_n N_VPWR_c_807_n 0.0227343f $X=1.89 $Y=2.495 $X2=0
+ $Y2=0
cc_331 N_A_350_102#_M1014_g N_VPWR_c_808_n 0.00479274f $X=3.655 $Y=2.775 $X2=0
+ $Y2=0
cc_332 N_A_350_102#_c_390_n N_VPWR_c_811_n 0.0165564f $X=1.89 $Y=2.495 $X2=0
+ $Y2=0
cc_333 N_A_350_102#_M1014_g N_VPWR_c_813_n 0.00432313f $X=3.655 $Y=2.775 $X2=0
+ $Y2=0
cc_334 N_A_350_102#_M1014_g N_VPWR_c_806_n 0.0063357f $X=3.655 $Y=2.775 $X2=0
+ $Y2=0
cc_335 N_A_350_102#_c_390_n N_VPWR_c_806_n 0.0122141f $X=1.89 $Y=2.495 $X2=0
+ $Y2=0
cc_336 N_A_350_102#_c_383_n N_VGND_c_925_n 0.00803878f $X=1.89 $Y=0.72 $X2=0
+ $Y2=0
cc_337 N_A_350_102#_M1023_g N_VGND_c_926_n 0.0101381f $X=3.875 $Y=0.445 $X2=0
+ $Y2=0
cc_338 N_A_350_102#_c_383_n N_VGND_c_930_n 0.00925243f $X=1.89 $Y=0.72 $X2=0
+ $Y2=0
cc_339 N_A_350_102#_M1023_g N_VGND_c_931_n 0.00437852f $X=3.875 $Y=0.445 $X2=0
+ $Y2=0
cc_340 N_A_350_102#_M1023_g N_VGND_c_934_n 0.00664875f $X=3.875 $Y=0.445 $X2=0
+ $Y2=0
cc_341 N_A_350_102#_c_383_n N_VGND_c_934_n 0.0110254f $X=1.89 $Y=0.72 $X2=0
+ $Y2=0
cc_342 N_A_463_491#_M1008_g N_A_1027_407#_M1027_g 0.0163661f $X=4.59 $Y=2.885
+ $X2=0 $Y2=0
cc_343 N_A_463_491#_c_494_n N_A_1027_407#_M1027_g 8.55913e-19 $X=4.73 $Y=2.35
+ $X2=0 $Y2=0
cc_344 N_A_463_491#_c_495_n N_A_1027_407#_M1027_g 0.0174966f $X=4.73 $Y=2.35
+ $X2=0 $Y2=0
cc_345 N_A_463_491#_c_489_n N_A_1027_407#_c_600_n 0.00131459f $X=4.672 $Y=2.185
+ $X2=0 $Y2=0
cc_346 N_A_463_491#_c_489_n N_A_1027_407#_c_615_n 7.63216e-19 $X=4.672 $Y=2.185
+ $X2=0 $Y2=0
cc_347 N_A_463_491#_c_492_n N_A_824_491#_M1016_d 0.00654576f $X=4.45 $Y=2.56
+ $X2=0 $Y2=0
cc_348 N_A_463_491#_M1008_g N_A_824_491#_c_719_n 0.0133076f $X=4.59 $Y=2.885
+ $X2=0 $Y2=0
cc_349 N_A_463_491#_c_492_n N_A_824_491#_c_719_n 0.0199446f $X=4.45 $Y=2.56
+ $X2=0 $Y2=0
cc_350 N_A_463_491#_c_494_n N_A_824_491#_c_719_n 0.0281346f $X=4.73 $Y=2.35
+ $X2=0 $Y2=0
cc_351 N_A_463_491#_c_495_n N_A_824_491#_c_719_n 0.00107667f $X=4.73 $Y=2.35
+ $X2=0 $Y2=0
cc_352 N_A_463_491#_M1004_g N_A_824_491#_c_709_n 7.16946e-19 $X=4.265 $Y=0.445
+ $X2=0 $Y2=0
cc_353 N_A_463_491#_c_487_n N_A_824_491#_c_709_n 0.0288813f $X=4.355 $Y=1.02
+ $X2=0 $Y2=0
cc_354 N_A_463_491#_c_488_n N_A_824_491#_c_709_n 3.28046e-19 $X=4.355 $Y=1.02
+ $X2=0 $Y2=0
cc_355 N_A_463_491#_c_489_n N_A_824_491#_c_709_n 0.0170925f $X=4.672 $Y=2.185
+ $X2=0 $Y2=0
cc_356 N_A_463_491#_M1008_g N_A_824_491#_c_710_n 0.00330151f $X=4.59 $Y=2.885
+ $X2=0 $Y2=0
cc_357 N_A_463_491#_c_494_n N_A_824_491#_c_710_n 0.0344482f $X=4.73 $Y=2.35
+ $X2=0 $Y2=0
cc_358 N_A_463_491#_c_495_n N_A_824_491#_c_710_n 0.00191077f $X=4.73 $Y=2.35
+ $X2=0 $Y2=0
cc_359 N_A_463_491#_c_489_n N_A_824_491#_c_710_n 0.0214978f $X=4.672 $Y=2.185
+ $X2=0 $Y2=0
cc_360 N_A_463_491#_c_494_n N_A_824_491#_c_712_n 0.00251056f $X=4.73 $Y=2.35
+ $X2=0 $Y2=0
cc_361 N_A_463_491#_c_489_n N_A_824_491#_c_712_n 0.0128538f $X=4.672 $Y=2.185
+ $X2=0 $Y2=0
cc_362 N_A_463_491#_M1004_g N_A_824_491#_c_713_n 0.0113744f $X=4.265 $Y=0.445
+ $X2=0 $Y2=0
cc_363 N_A_463_491#_c_487_n N_A_824_491#_c_713_n 0.0136156f $X=4.355 $Y=1.02
+ $X2=0 $Y2=0
cc_364 N_A_463_491#_c_488_n N_A_824_491#_c_713_n 4.86079e-19 $X=4.355 $Y=1.02
+ $X2=0 $Y2=0
cc_365 N_A_463_491#_c_492_n N_VPWR_M1024_d 0.00821965f $X=4.45 $Y=2.56 $X2=0
+ $Y2=0
cc_366 N_A_463_491#_c_492_n N_VPWR_c_808_n 0.0239947f $X=4.45 $Y=2.56 $X2=0
+ $Y2=0
cc_367 N_A_463_491#_c_491_n N_VPWR_c_811_n 0.019689f $X=2.46 $Y=2.645 $X2=0
+ $Y2=0
cc_368 N_A_463_491#_c_492_n N_VPWR_c_811_n 0.0074229f $X=4.45 $Y=2.56 $X2=0
+ $Y2=0
cc_369 N_A_463_491#_M1008_g N_VPWR_c_813_n 0.00366111f $X=4.59 $Y=2.885 $X2=0
+ $Y2=0
cc_370 N_A_463_491#_c_492_n N_VPWR_c_813_n 0.00742889f $X=4.45 $Y=2.56 $X2=0
+ $Y2=0
cc_371 N_A_463_491#_M1021_s N_VPWR_c_806_n 0.00232985f $X=2.315 $Y=2.455 $X2=0
+ $Y2=0
cc_372 N_A_463_491#_M1008_g N_VPWR_c_806_n 0.00618118f $X=4.59 $Y=2.885 $X2=0
+ $Y2=0
cc_373 N_A_463_491#_c_491_n N_VPWR_c_806_n 0.0125545f $X=2.46 $Y=2.645 $X2=0
+ $Y2=0
cc_374 N_A_463_491#_c_492_n N_VPWR_c_806_n 0.030613f $X=4.45 $Y=2.56 $X2=0 $Y2=0
cc_375 N_A_463_491#_c_492_n A_550_491# 0.00417663f $X=4.45 $Y=2.56 $X2=-0.19
+ $Y2=-0.245
cc_376 N_A_463_491#_c_492_n A_746_491# 0.00712663f $X=4.45 $Y=2.56 $X2=-0.19
+ $Y2=-0.245
cc_377 N_A_463_491#_c_484_n N_VGND_c_926_n 0.00887059f $X=2.63 $Y=0.47 $X2=0
+ $Y2=0
cc_378 N_A_463_491#_c_485_n N_VGND_c_926_n 0.0222125f $X=4.105 $Y=0.81 $X2=0
+ $Y2=0
cc_379 N_A_463_491#_c_484_n N_VGND_c_930_n 0.019689f $X=2.63 $Y=0.47 $X2=0 $Y2=0
cc_380 N_A_463_491#_c_485_n N_VGND_c_930_n 0.00697632f $X=4.105 $Y=0.81 $X2=0
+ $Y2=0
cc_381 N_A_463_491#_M1004_g N_VGND_c_931_n 0.00501706f $X=4.265 $Y=0.445 $X2=0
+ $Y2=0
cc_382 N_A_463_491#_c_485_n N_VGND_c_931_n 0.0071588f $X=4.105 $Y=0.81 $X2=0
+ $Y2=0
cc_383 N_A_463_491#_c_487_n N_VGND_c_931_n 0.00261587f $X=4.355 $Y=1.02 $X2=0
+ $Y2=0
cc_384 N_A_463_491#_M1003_s N_VGND_c_934_n 0.00232985f $X=2.485 $Y=0.235 $X2=0
+ $Y2=0
cc_385 N_A_463_491#_M1004_g N_VGND_c_934_n 0.00665371f $X=4.265 $Y=0.445 $X2=0
+ $Y2=0
cc_386 N_A_463_491#_c_484_n N_VGND_c_934_n 0.0125545f $X=2.63 $Y=0.47 $X2=0
+ $Y2=0
cc_387 N_A_463_491#_c_485_n N_VGND_c_934_n 0.0254529f $X=4.105 $Y=0.81 $X2=0
+ $Y2=0
cc_388 N_A_463_491#_c_487_n N_VGND_c_934_n 0.0102353f $X=4.355 $Y=1.02 $X2=0
+ $Y2=0
cc_389 N_A_1027_407#_M1005_g N_A_824_491#_M1025_g 0.0129895f $X=5.225 $Y=0.445
+ $X2=0 $Y2=0
cc_390 N_A_1027_407#_c_600_n N_A_824_491#_M1025_g 0.00749249f $X=5.217 $Y=2.035
+ $X2=0 $Y2=0
cc_391 N_A_1027_407#_c_601_n N_A_824_491#_M1025_g 0.0151998f $X=6.355 $Y=1.01
+ $X2=0 $Y2=0
cc_392 N_A_1027_407#_c_602_n N_A_824_491#_M1025_g 0.00326863f $X=6.52 $Y=0.43
+ $X2=0 $Y2=0
cc_393 N_A_1027_407#_c_603_n N_A_824_491#_M1025_g 8.84346e-19 $X=6.52 $Y=1.305
+ $X2=0 $Y2=0
cc_394 N_A_1027_407#_c_606_n N_A_824_491#_M1025_g 0.00105957f $X=5.315 $Y=1.01
+ $X2=0 $Y2=0
cc_395 N_A_1027_407#_c_607_n N_A_824_491#_M1025_g 0.0114028f $X=5.315 $Y=1.09
+ $X2=0 $Y2=0
cc_396 N_A_1027_407#_M1027_g N_A_824_491#_M1011_g 0.00922615f $X=5.21 $Y=2.885
+ $X2=0 $Y2=0
cc_397 N_A_1027_407#_c_600_n N_A_824_491#_M1011_g 0.00714936f $X=5.217 $Y=2.035
+ $X2=0 $Y2=0
cc_398 N_A_1027_407#_c_604_n N_A_824_491#_M1011_g 0.00430196f $X=6.52 $Y=1.98
+ $X2=0 $Y2=0
cc_399 N_A_1027_407#_c_601_n N_A_824_491#_M1026_g 0.0146769f $X=6.355 $Y=1.01
+ $X2=0 $Y2=0
cc_400 N_A_1027_407#_c_602_n N_A_824_491#_M1026_g 0.0141035f $X=6.52 $Y=0.43
+ $X2=0 $Y2=0
cc_401 N_A_1027_407#_c_603_n N_A_824_491#_M1026_g 0.00676102f $X=6.52 $Y=1.305
+ $X2=0 $Y2=0
cc_402 N_A_1027_407#_c_608_n N_A_824_491#_M1026_g 7.69939e-19 $X=6.52 $Y=1.01
+ $X2=0 $Y2=0
cc_403 N_A_1027_407#_c_604_n N_A_824_491#_M1013_g 0.0300568f $X=6.52 $Y=1.98
+ $X2=0 $Y2=0
cc_404 N_A_1027_407#_c_609_n N_A_824_491#_M1013_g 0.00124383f $X=6.52 $Y=1.47
+ $X2=0 $Y2=0
cc_405 N_A_1027_407#_M1027_g N_A_824_491#_c_719_n 0.00886129f $X=5.21 $Y=2.885
+ $X2=0 $Y2=0
cc_406 N_A_1027_407#_M1005_g N_A_824_491#_c_709_n 0.0104525f $X=5.225 $Y=0.445
+ $X2=0 $Y2=0
cc_407 N_A_1027_407#_c_606_n N_A_824_491#_c_709_n 0.0237562f $X=5.315 $Y=1.01
+ $X2=0 $Y2=0
cc_408 N_A_1027_407#_M1027_g N_A_824_491#_c_710_n 0.0165691f $X=5.21 $Y=2.885
+ $X2=0 $Y2=0
cc_409 N_A_1027_407#_c_600_n N_A_824_491#_c_710_n 0.0145243f $X=5.217 $Y=2.035
+ $X2=0 $Y2=0
cc_410 N_A_1027_407#_c_615_n N_A_824_491#_c_710_n 0.00565524f $X=5.217 $Y=2.185
+ $X2=0 $Y2=0
cc_411 N_A_1027_407#_c_600_n N_A_824_491#_c_711_n 0.00705157f $X=5.217 $Y=2.035
+ $X2=0 $Y2=0
cc_412 N_A_1027_407#_c_601_n N_A_824_491#_c_711_n 0.0167829f $X=6.355 $Y=1.01
+ $X2=0 $Y2=0
cc_413 N_A_1027_407#_c_607_n N_A_824_491#_c_711_n 0.00124625f $X=5.315 $Y=1.09
+ $X2=0 $Y2=0
cc_414 N_A_1027_407#_c_600_n N_A_824_491#_c_712_n 0.00483065f $X=5.217 $Y=2.035
+ $X2=0 $Y2=0
cc_415 N_A_1027_407#_c_606_n N_A_824_491#_c_712_n 0.0231277f $X=5.315 $Y=1.01
+ $X2=0 $Y2=0
cc_416 N_A_1027_407#_M1005_g N_A_824_491#_c_713_n 0.00197903f $X=5.225 $Y=0.445
+ $X2=0 $Y2=0
cc_417 N_A_1027_407#_c_600_n N_A_824_491#_c_714_n 9.35823e-19 $X=5.217 $Y=2.035
+ $X2=0 $Y2=0
cc_418 N_A_1027_407#_c_601_n N_A_824_491#_c_714_n 0.0231622f $X=6.355 $Y=1.01
+ $X2=0 $Y2=0
cc_419 N_A_1027_407#_c_603_n N_A_824_491#_c_714_n 0.00206876f $X=6.52 $Y=1.305
+ $X2=0 $Y2=0
cc_420 N_A_1027_407#_c_609_n N_A_824_491#_c_714_n 0.0223693f $X=6.52 $Y=1.47
+ $X2=0 $Y2=0
cc_421 N_A_1027_407#_c_601_n N_A_824_491#_c_715_n 4.15005e-19 $X=6.355 $Y=1.01
+ $X2=0 $Y2=0
cc_422 N_A_1027_407#_c_603_n N_A_824_491#_c_715_n 0.00107786f $X=6.52 $Y=1.305
+ $X2=0 $Y2=0
cc_423 N_A_1027_407#_c_609_n N_A_824_491#_c_715_n 0.0127182f $X=6.52 $Y=1.47
+ $X2=0 $Y2=0
cc_424 N_A_1027_407#_M1027_g N_VPWR_c_809_n 0.0108417f $X=5.21 $Y=2.885 $X2=0
+ $Y2=0
cc_425 N_A_1027_407#_c_600_n N_VPWR_c_809_n 0.00330804f $X=5.217 $Y=2.035 $X2=0
+ $Y2=0
cc_426 N_A_1027_407#_c_604_n N_VPWR_c_809_n 0.0418217f $X=6.52 $Y=1.98 $X2=0
+ $Y2=0
cc_427 N_A_1027_407#_M1006_g N_VPWR_c_810_n 0.0308985f $X=7.295 $Y=2.465 $X2=0
+ $Y2=0
cc_428 N_A_1027_407#_M1007_g N_VPWR_c_810_n 0.00468428f $X=7.655 $Y=2.465 $X2=0
+ $Y2=0
cc_429 N_A_1027_407#_c_604_n N_VPWR_c_810_n 0.0842731f $X=6.52 $Y=1.98 $X2=0
+ $Y2=0
cc_430 N_A_1027_407#_c_605_n N_VPWR_c_810_n 0.0275493f $X=7.36 $Y=1.47 $X2=0
+ $Y2=0
cc_431 N_A_1027_407#_c_610_n N_VPWR_c_810_n 5.79521e-19 $X=7.655 $Y=1.47 $X2=0
+ $Y2=0
cc_432 N_A_1027_407#_M1027_g N_VPWR_c_813_n 0.00424436f $X=5.21 $Y=2.885 $X2=0
+ $Y2=0
cc_433 N_A_1027_407#_c_604_n N_VPWR_c_816_n 0.019758f $X=6.52 $Y=1.98 $X2=0
+ $Y2=0
cc_434 N_A_1027_407#_M1006_g N_VPWR_c_817_n 0.00486043f $X=7.295 $Y=2.465 $X2=0
+ $Y2=0
cc_435 N_A_1027_407#_M1007_g N_VPWR_c_817_n 0.00549284f $X=7.655 $Y=2.465 $X2=0
+ $Y2=0
cc_436 N_A_1027_407#_M1013_d N_VPWR_c_806_n 0.0023218f $X=6.38 $Y=1.835 $X2=0
+ $Y2=0
cc_437 N_A_1027_407#_M1027_g N_VPWR_c_806_n 0.00800058f $X=5.21 $Y=2.885 $X2=0
+ $Y2=0
cc_438 N_A_1027_407#_M1006_g N_VPWR_c_806_n 0.00814425f $X=7.295 $Y=2.465 $X2=0
+ $Y2=0
cc_439 N_A_1027_407#_M1007_g N_VPWR_c_806_n 0.0107699f $X=7.655 $Y=2.465 $X2=0
+ $Y2=0
cc_440 N_A_1027_407#_c_604_n N_VPWR_c_806_n 0.012508f $X=6.52 $Y=1.98 $X2=0
+ $Y2=0
cc_441 N_A_1027_407#_M1015_g N_Q_c_910_n 0.00323857f $X=7.295 $Y=0.685 $X2=0
+ $Y2=0
cc_442 N_A_1027_407#_M1006_g N_Q_c_910_n 0.00430008f $X=7.295 $Y=2.465 $X2=0
+ $Y2=0
cc_443 N_A_1027_407#_M1018_g N_Q_c_910_n 0.0238324f $X=7.655 $Y=0.685 $X2=0
+ $Y2=0
cc_444 N_A_1027_407#_M1007_g N_Q_c_910_n 0.0300568f $X=7.655 $Y=2.465 $X2=0
+ $Y2=0
cc_445 N_A_1027_407#_c_605_n N_Q_c_910_n 0.0250026f $X=7.36 $Y=1.47 $X2=0 $Y2=0
cc_446 N_A_1027_407#_c_610_n N_Q_c_910_n 0.0121537f $X=7.655 $Y=1.47 $X2=0 $Y2=0
cc_447 N_A_1027_407#_c_601_n N_VGND_M1005_d 0.00687908f $X=6.355 $Y=1.01 $X2=0
+ $Y2=0
cc_448 N_A_1027_407#_M1005_g N_VGND_c_927_n 0.0128234f $X=5.225 $Y=0.445 $X2=0
+ $Y2=0
cc_449 N_A_1027_407#_c_601_n N_VGND_c_927_n 0.00825341f $X=6.355 $Y=1.01 $X2=0
+ $Y2=0
cc_450 N_A_1027_407#_c_606_n N_VGND_c_927_n 0.0124765f $X=5.315 $Y=1.01 $X2=0
+ $Y2=0
cc_451 N_A_1027_407#_c_607_n N_VGND_c_927_n 0.0013518f $X=5.315 $Y=1.09 $X2=0
+ $Y2=0
cc_452 N_A_1027_407#_M1015_g N_VGND_c_928_n 0.0234518f $X=7.295 $Y=0.685 $X2=0
+ $Y2=0
cc_453 N_A_1027_407#_M1018_g N_VGND_c_928_n 0.00336955f $X=7.655 $Y=0.685 $X2=0
+ $Y2=0
cc_454 N_A_1027_407#_c_602_n N_VGND_c_928_n 0.0444625f $X=6.52 $Y=0.43 $X2=0
+ $Y2=0
cc_455 N_A_1027_407#_c_603_n N_VGND_c_928_n 0.00198884f $X=6.52 $Y=1.305 $X2=0
+ $Y2=0
cc_456 N_A_1027_407#_c_605_n N_VGND_c_928_n 0.0275493f $X=7.36 $Y=1.47 $X2=0
+ $Y2=0
cc_457 N_A_1027_407#_c_608_n N_VGND_c_928_n 0.0121616f $X=6.52 $Y=1.01 $X2=0
+ $Y2=0
cc_458 N_A_1027_407#_c_610_n N_VGND_c_928_n 5.79521e-19 $X=7.655 $Y=1.47 $X2=0
+ $Y2=0
cc_459 N_A_1027_407#_M1005_g N_VGND_c_931_n 0.00505556f $X=5.225 $Y=0.445 $X2=0
+ $Y2=0
cc_460 N_A_1027_407#_c_602_n N_VGND_c_932_n 0.019758f $X=6.52 $Y=0.43 $X2=0
+ $Y2=0
cc_461 N_A_1027_407#_M1015_g N_VGND_c_933_n 0.00461019f $X=7.295 $Y=0.685 $X2=0
+ $Y2=0
cc_462 N_A_1027_407#_M1018_g N_VGND_c_933_n 0.00520813f $X=7.655 $Y=0.685 $X2=0
+ $Y2=0
cc_463 N_A_1027_407#_M1026_d N_VGND_c_934_n 0.0023218f $X=6.38 $Y=0.235 $X2=0
+ $Y2=0
cc_464 N_A_1027_407#_M1005_g N_VGND_c_934_n 0.00858274f $X=5.225 $Y=0.445 $X2=0
+ $Y2=0
cc_465 N_A_1027_407#_M1015_g N_VGND_c_934_n 0.00803623f $X=7.295 $Y=0.685 $X2=0
+ $Y2=0
cc_466 N_A_1027_407#_M1018_g N_VGND_c_934_n 0.0104074f $X=7.655 $Y=0.685 $X2=0
+ $Y2=0
cc_467 N_A_1027_407#_c_602_n N_VGND_c_934_n 0.012508f $X=6.52 $Y=0.43 $X2=0
+ $Y2=0
cc_468 N_A_1027_407#_c_601_n A_1198_47# 0.0048076f $X=6.355 $Y=1.01 $X2=-0.19
+ $Y2=-0.245
cc_469 N_A_824_491#_M1011_g N_VPWR_c_809_n 0.0294135f $X=5.945 $Y=2.465 $X2=0
+ $Y2=0
cc_470 N_A_824_491#_M1013_g N_VPWR_c_809_n 0.00468428f $X=6.305 $Y=2.465 $X2=0
+ $Y2=0
cc_471 N_A_824_491#_c_719_n N_VPWR_c_809_n 0.0106216f $X=5.075 $Y=2.93 $X2=0
+ $Y2=0
cc_472 N_A_824_491#_c_710_n N_VPWR_c_809_n 0.0474269f $X=5.16 $Y=2.825 $X2=0
+ $Y2=0
cc_473 N_A_824_491#_c_711_n N_VPWR_c_809_n 0.0199403f $X=5.84 $Y=1.52 $X2=0
+ $Y2=0
cc_474 N_A_824_491#_c_714_n N_VPWR_c_809_n 0.00371908f $X=6.005 $Y=1.44 $X2=0
+ $Y2=0
cc_475 N_A_824_491#_c_715_n N_VPWR_c_809_n 2.21141e-19 $X=6.305 $Y=1.44 $X2=0
+ $Y2=0
cc_476 N_A_824_491#_M1013_g N_VPWR_c_810_n 0.0048055f $X=6.305 $Y=2.465 $X2=0
+ $Y2=0
cc_477 N_A_824_491#_c_719_n N_VPWR_c_813_n 0.0536297f $X=5.075 $Y=2.93 $X2=0
+ $Y2=0
cc_478 N_A_824_491#_M1011_g N_VPWR_c_816_n 0.00486043f $X=5.945 $Y=2.465 $X2=0
+ $Y2=0
cc_479 N_A_824_491#_M1013_g N_VPWR_c_816_n 0.00549284f $X=6.305 $Y=2.465 $X2=0
+ $Y2=0
cc_480 N_A_824_491#_M1016_d N_VPWR_c_806_n 0.00320268f $X=4.12 $Y=2.455 $X2=0
+ $Y2=0
cc_481 N_A_824_491#_M1011_g N_VPWR_c_806_n 0.00814425f $X=5.945 $Y=2.465 $X2=0
+ $Y2=0
cc_482 N_A_824_491#_M1013_g N_VPWR_c_806_n 0.0111098f $X=6.305 $Y=2.465 $X2=0
+ $Y2=0
cc_483 N_A_824_491#_c_719_n N_VPWR_c_806_n 0.0411834f $X=5.075 $Y=2.93 $X2=0
+ $Y2=0
cc_484 N_A_824_491#_c_719_n A_933_535# 0.0134944f $X=5.075 $Y=2.93 $X2=-0.19
+ $Y2=-0.245
cc_485 N_A_824_491#_c_710_n A_933_535# 0.00211708f $X=5.16 $Y=2.825 $X2=-0.19
+ $Y2=-0.245
cc_486 N_A_824_491#_M1025_g N_VGND_c_927_n 0.01282f $X=5.915 $Y=0.655 $X2=0
+ $Y2=0
cc_487 N_A_824_491#_c_713_n N_VGND_c_927_n 0.0162395f $X=4.62 $Y=0.47 $X2=0
+ $Y2=0
cc_488 N_A_824_491#_M1026_g N_VGND_c_928_n 0.0041367f $X=6.305 $Y=0.655 $X2=0
+ $Y2=0
cc_489 N_A_824_491#_c_713_n N_VGND_c_931_n 0.0231974f $X=4.62 $Y=0.47 $X2=0
+ $Y2=0
cc_490 N_A_824_491#_M1025_g N_VGND_c_932_n 0.00585385f $X=5.915 $Y=0.655 $X2=0
+ $Y2=0
cc_491 N_A_824_491#_M1026_g N_VGND_c_932_n 0.00549284f $X=6.305 $Y=0.655 $X2=0
+ $Y2=0
cc_492 N_A_824_491#_M1004_d N_VGND_c_934_n 0.00418738f $X=4.34 $Y=0.235 $X2=0
+ $Y2=0
cc_493 N_A_824_491#_M1025_g N_VGND_c_934_n 0.0114331f $X=5.915 $Y=0.655 $X2=0
+ $Y2=0
cc_494 N_A_824_491#_M1026_g N_VGND_c_934_n 0.0112036f $X=6.305 $Y=0.655 $X2=0
+ $Y2=0
cc_495 N_A_824_491#_c_713_n N_VGND_c_934_n 0.0179959f $X=4.62 $Y=0.47 $X2=0
+ $Y2=0
cc_496 N_A_824_491#_c_713_n A_982_47# 0.00166536f $X=4.62 $Y=0.47 $X2=-0.19
+ $Y2=-0.245
cc_497 N_VPWR_c_806_n A_550_491# 0.00296601f $X=7.92 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_498 N_VPWR_c_806_n A_746_491# 0.00296601f $X=7.92 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_499 N_VPWR_c_806_n A_933_535# 0.00384478f $X=7.92 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_500 N_VPWR_c_806_n A_1204_367# 0.00899413f $X=7.92 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_501 N_VPWR_c_806_n A_1474_367# 0.00899413f $X=7.92 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_502 N_VPWR_c_806_n N_Q_M1007_d 0.0023218f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_503 N_VPWR_c_810_n N_Q_c_910_n 0.0418217f $X=7.08 $Y=1.98 $X2=0 $Y2=0
cc_504 N_VPWR_c_817_n N_Q_c_910_n 0.019758f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_505 N_VPWR_c_806_n N_Q_c_910_n 0.012508f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_506 N_Q_c_910_n N_VGND_c_928_n 0.0287733f $X=7.87 $Y=0.43 $X2=0 $Y2=0
cc_507 N_Q_c_910_n N_VGND_c_933_n 0.019758f $X=7.87 $Y=0.43 $X2=0 $Y2=0
cc_508 N_Q_c_910_n N_VGND_c_934_n 0.0125705f $X=7.87 $Y=0.43 $X2=0 $Y2=0
cc_509 N_VGND_c_934_n A_584_47# 0.0031085f $X=7.92 $Y=0 $X2=-0.19 $Y2=-0.245
cc_510 N_VGND_c_934_n A_790_47# 0.00310724f $X=7.92 $Y=0 $X2=-0.19 $Y2=-0.245
cc_511 N_VGND_c_934_n A_982_47# 0.00830093f $X=7.92 $Y=0 $X2=-0.19 $Y2=-0.245
cc_512 N_VGND_c_934_n A_1198_47# 0.010279f $X=7.92 $Y=0 $X2=-0.19 $Y2=-0.245
