* File: sky130_fd_sc_lp__nand2_lp.spice
* Created: Fri Aug 28 10:47:41 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__nand2_lp.pex.spice"
.subckt sky130_fd_sc_lp__nand2_lp  VNB VPB B A Y VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Y	Y
* A	A
* B	B
* VPB	VPB
* VNB	VNB
MM1000 A_121_57# N_B_M1000_g N_VGND_M1000_s VNB NSHORT L=0.15 W=0.42 AD=0.0504
+ AS=0.1197 PD=0.66 PS=1.41 NRD=18.564 NRS=0 M=1 R=2.8 SA=75000.2 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1004 N_Y_M1004_d N_A_M1004_g A_121_57# VNB NSHORT L=0.15 W=0.42 AD=0.1197
+ AS=0.0504 PD=1.41 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75000.6 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1003 N_Y_M1003_d N_B_M1003_g A_39_367# VPB PHIGHVT L=0.15 W=0.42 AD=0.0588
+ AS=0.134175 PD=0.7 PS=1.445 NRD=0 NRS=124.031 M=1 R=2.8 SA=75000.2 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1002 N_VPWR_M1002_d N_B_M1002_g A_39_367# VPB PHIGHVT L=0.15 W=0.42 AD=0.0588
+ AS=0.134175 PD=0.7 PS=1.445 NRD=0 NRS=124.031 M=1 R=2.8 SA=75000.2 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1001 A_207_367# N_A_M1001_g N_Y_M1003_d VPB PHIGHVT L=0.15 W=0.42 AD=0.134175
+ AS=0.0588 PD=1.445 PS=0.7 NRD=124.031 NRS=0 M=1 R=2.8 SA=75000.6 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1005 A_207_367# N_A_M1005_g N_VPWR_M1002_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.134175 AS=0.0588 PD=1.445 PS=0.7 NRD=124.031 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
DX6_noxref VNB VPB NWDIODE A=3.3943 P=7.37
*
.include "sky130_fd_sc_lp__nand2_lp.pxi.spice"
*
.ends
*
*
