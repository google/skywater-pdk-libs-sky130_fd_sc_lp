* File: sky130_fd_sc_lp__conb_1.pxi.spice
* Created: Wed Sep  2 09:41:39 2020
* 
x_PM_SKY130_FD_SC_LP__CONB_1%HI N_HI_M1002_d N_HI_M1001_g N_HI_M1002_g
+ N_HI_c_37_n N_HI_c_42_n HI HI HI N_HI_c_39_n N_HI_c_45_n
+ PM_SKY130_FD_SC_LP__CONB_1%HI
x_PM_SKY130_FD_SC_LP__CONB_1%LO N_LO_M1001_d N_LO_M1003_g N_LO_c_76_n
+ N_LO_M1000_g N_LO_c_78_n N_LO_c_79_n N_LO_c_80_n N_LO_c_81_n LO LO LO LO
+ N_LO_c_83_n N_LO_c_84_n N_LO_c_85_n PM_SKY130_FD_SC_LP__CONB_1%LO
x_PM_SKY130_FD_SC_LP__CONB_1%VPWR N_VPWR_M1002_s N_VPWR_M1000_d N_VPWR_c_117_n
+ N_VPWR_c_118_n N_VPWR_c_119_n N_VPWR_c_120_n VPWR N_VPWR_c_121_n
+ N_VPWR_c_116_n PM_SKY130_FD_SC_LP__CONB_1%VPWR
x_PM_SKY130_FD_SC_LP__CONB_1%VGND N_VGND_M1001_s N_VGND_M1003_d N_VGND_c_137_n
+ N_VGND_c_138_n N_VGND_c_139_n N_VGND_c_140_n VGND N_VGND_c_141_n
+ N_VGND_c_142_n PM_SKY130_FD_SC_LP__CONB_1%VGND
cc_1 VNB N_HI_M1001_g 0.0478609f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=0.56
cc_2 VNB N_HI_c_37_n 0.0277298f $X=-0.19 $Y=-0.245 $X2=0.445 $Y2=1.715
cc_3 VNB HI 0.0105848f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_4 VNB N_HI_c_39_n 0.0215086f $X=-0.19 $Y=-0.245 $X2=0.445 $Y2=1.375
cc_5 VNB N_LO_c_76_n 0.0246543f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=1.88
cc_6 VNB N_LO_M1000_g 0.00659088f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_LO_c_78_n 0.0246924f $X=-0.19 $Y=-0.245 $X2=0.445 $Y2=1.21
cc_8 VNB N_LO_c_79_n 0.00149799f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_9 VNB N_LO_c_80_n 0.00206843f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.95
cc_10 VNB N_LO_c_81_n 0.00443662f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB LO 0.00985671f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_LO_c_83_n 0.0239118f $X=-0.19 $Y=-0.245 $X2=0.567 $Y2=1.375
cc_13 VNB N_LO_c_84_n 0.0239107f $X=-0.19 $Y=-0.245 $X2=0.567 $Y2=1.665
cc_14 VNB N_LO_c_85_n 0.0210234f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_VPWR_c_116_n 0.0641695f $X=-0.19 $Y=-0.245 $X2=0.567 $Y2=1.295
cc_16 VNB N_VGND_c_137_n 0.0128195f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_VGND_c_138_n 0.0268384f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=2.63
cc_18 VNB N_VGND_c_139_n 0.0112376f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_VGND_c_140_n 0.0210568f $X=-0.19 $Y=-0.245 $X2=0.445 $Y2=1.21
cc_20 VNB N_VGND_c_141_n 0.0160313f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_21 VNB N_VGND_c_142_n 0.112687f $X=-0.19 $Y=-0.245 $X2=0.567 $Y2=1.295
cc_22 VPB N_HI_M1002_g 0.0388983f $X=-0.19 $Y=1.655 $X2=0.535 $Y2=2.63
cc_23 VPB N_HI_c_37_n 0.00586401f $X=-0.19 $Y=1.655 $X2=0.445 $Y2=1.715
cc_24 VPB N_HI_c_42_n 0.0214953f $X=-0.19 $Y=1.655 $X2=0.445 $Y2=1.88
cc_25 VPB HI 0.00148033f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_26 VPB HI 0.0147767f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.95
cc_27 VPB N_HI_c_45_n 0.00439212f $X=-0.19 $Y=1.655 $X2=0.75 $Y2=2.465
cc_28 VPB N_LO_M1000_g 0.0567796f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_29 VPB N_LO_c_84_n 0.022454f $X=-0.19 $Y=1.655 $X2=0.567 $Y2=1.665
cc_30 VPB N_VPWR_c_117_n 0.0123127f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_31 VPB N_VPWR_c_118_n 0.0435358f $X=-0.19 $Y=1.655 $X2=0.535 $Y2=2.63
cc_32 VPB N_VPWR_c_119_n 0.0112524f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_33 VPB N_VPWR_c_120_n 0.0382385f $X=-0.19 $Y=1.655 $X2=0.445 $Y2=1.21
cc_34 VPB N_VPWR_c_121_n 0.016961f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_35 VPB N_VPWR_c_116_n 0.0553055f $X=-0.19 $Y=1.655 $X2=0.567 $Y2=1.295
cc_36 N_HI_c_37_n N_LO_c_76_n 0.0151632f $X=0.445 $Y=1.715 $X2=0 $Y2=0
cc_37 HI N_LO_c_76_n 0.00436619f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_38 N_HI_M1002_g N_LO_M1000_g 0.0151632f $X=0.535 $Y=2.63 $X2=0 $Y2=0
cc_39 N_HI_c_45_n N_LO_M1000_g 0.00436619f $X=0.75 $Y=2.465 $X2=0 $Y2=0
cc_40 N_HI_c_42_n N_LO_c_78_n 0.0151632f $X=0.445 $Y=1.88 $X2=0 $Y2=0
cc_41 HI N_LO_c_78_n 0.00436619f $X=0.635 $Y=1.95 $X2=0 $Y2=0
cc_42 N_HI_M1001_g N_LO_c_79_n 0.00189162f $X=0.535 $Y=0.56 $X2=0 $Y2=0
cc_43 HI N_LO_c_80_n 7.22336e-19 $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_44 N_HI_M1001_g N_LO_c_81_n 0.00568793f $X=0.535 $Y=0.56 $X2=0 $Y2=0
cc_45 HI N_LO_c_81_n 0.0209253f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_46 N_HI_c_39_n N_LO_c_83_n 0.0151632f $X=0.445 $Y=1.375 $X2=0 $Y2=0
cc_47 N_HI_M1001_g N_LO_c_84_n 0.00145908f $X=0.535 $Y=0.56 $X2=0 $Y2=0
cc_48 HI N_LO_c_84_n 0.0742647f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_49 N_HI_M1001_g N_LO_c_85_n 0.0151632f $X=0.535 $Y=0.56 $X2=0 $Y2=0
cc_50 N_HI_M1002_g N_VPWR_c_118_n 0.0040936f $X=0.535 $Y=2.63 $X2=0 $Y2=0
cc_51 N_HI_c_42_n N_VPWR_c_118_n 6.54183e-19 $X=0.445 $Y=1.88 $X2=0 $Y2=0
cc_52 HI N_VPWR_c_118_n 0.0133984f $X=0.635 $Y=1.95 $X2=0 $Y2=0
cc_53 N_HI_c_45_n N_VPWR_c_118_n 0.0261336f $X=0.75 $Y=2.465 $X2=0 $Y2=0
cc_54 N_HI_M1002_g N_VPWR_c_120_n 5.31725e-19 $X=0.535 $Y=2.63 $X2=0 $Y2=0
cc_55 N_HI_c_45_n N_VPWR_c_120_n 0.0269202f $X=0.75 $Y=2.465 $X2=0 $Y2=0
cc_56 N_HI_M1002_g N_VPWR_c_121_n 0.0055545f $X=0.535 $Y=2.63 $X2=0 $Y2=0
cc_57 N_HI_c_45_n N_VPWR_c_121_n 0.0110266f $X=0.75 $Y=2.465 $X2=0 $Y2=0
cc_58 N_HI_M1002_g N_VPWR_c_116_n 0.00542671f $X=0.535 $Y=2.63 $X2=0 $Y2=0
cc_59 N_HI_c_45_n N_VPWR_c_116_n 0.00945959f $X=0.75 $Y=2.465 $X2=0 $Y2=0
cc_60 N_HI_M1001_g N_VGND_c_138_n 0.00406185f $X=0.535 $Y=0.56 $X2=0 $Y2=0
cc_61 HI N_VGND_c_138_n 0.00660914f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_62 N_HI_c_39_n N_VGND_c_138_n 8.94736e-19 $X=0.445 $Y=1.375 $X2=0 $Y2=0
cc_63 N_HI_M1001_g N_VGND_c_140_n 5.44985e-19 $X=0.535 $Y=0.56 $X2=0 $Y2=0
cc_64 N_HI_M1001_g N_VGND_c_141_n 0.00478016f $X=0.535 $Y=0.56 $X2=0 $Y2=0
cc_65 N_HI_M1001_g N_VGND_c_142_n 0.00954948f $X=0.535 $Y=0.56 $X2=0 $Y2=0
cc_66 N_LO_M1000_g N_VPWR_c_120_n 0.0121794f $X=0.965 $Y=2.63 $X2=0 $Y2=0
cc_67 N_LO_c_84_n N_VPWR_c_120_n 0.0288227f $X=1.12 $Y=1.045 $X2=0 $Y2=0
cc_68 N_LO_M1000_g N_VPWR_c_121_n 0.00512473f $X=0.965 $Y=2.63 $X2=0 $Y2=0
cc_69 N_LO_M1000_g N_VPWR_c_116_n 0.00492022f $X=0.965 $Y=2.63 $X2=0 $Y2=0
cc_70 N_LO_c_80_n N_VGND_c_140_n 0.00138333f $X=1.035 $Y=0.925 $X2=0 $Y2=0
cc_71 LO N_VGND_c_140_n 0.0251301f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_72 N_LO_c_83_n N_VGND_c_140_n 0.00156152f $X=1.12 $Y=1.045 $X2=0 $Y2=0
cc_73 N_LO_c_85_n N_VGND_c_140_n 0.00952f $X=1.087 $Y=0.88 $X2=0 $Y2=0
cc_74 N_LO_c_79_n N_VGND_c_141_n 0.00715561f $X=0.75 $Y=0.56 $X2=0 $Y2=0
cc_75 N_LO_c_85_n N_VGND_c_141_n 0.00396895f $X=1.087 $Y=0.88 $X2=0 $Y2=0
cc_76 N_LO_c_79_n N_VGND_c_142_n 0.00797928f $X=0.75 $Y=0.56 $X2=0 $Y2=0
cc_77 N_LO_c_80_n N_VGND_c_142_n 0.00504476f $X=1.035 $Y=0.925 $X2=0 $Y2=0
cc_78 LO N_VGND_c_142_n 0.00155659f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_79 N_LO_c_85_n N_VGND_c_142_n 0.00398153f $X=1.087 $Y=0.88 $X2=0 $Y2=0
