* File: sky130_fd_sc_lp__nand4b_1.pex.spice
* Created: Wed Sep  2 10:06:03 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__NAND4B_1%A_N 3 6 8 11 13
r26 11 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.605 $Y=1.35
+ $X2=0.605 $Y2=1.515
r27 11 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.605 $Y=1.35
+ $X2=0.605 $Y2=1.185
r28 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.605
+ $Y=1.35 $X2=0.605 $Y2=1.35
r29 8 12 4.01609 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=0.72 $Y=1.35
+ $X2=0.605 $Y2=1.35
r30 6 14 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.695 $Y=2.045
+ $X2=0.695 $Y2=1.515
r31 3 13 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.695 $Y=0.865
+ $X2=0.695 $Y2=1.185
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4B_1%D 3 6 8 11 13
r29 11 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.145 $Y=1.35
+ $X2=1.145 $Y2=1.515
r30 11 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.145 $Y=1.35
+ $X2=1.145 $Y2=1.185
r31 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.145
+ $Y=1.35 $X2=1.145 $Y2=1.35
r32 6 14 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=1.235 $Y=2.465
+ $X2=1.235 $Y2=1.515
r33 3 13 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.235 $Y=0.655
+ $X2=1.235 $Y2=1.185
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4B_1%C 3 6 8 9 10 15 17
r35 15 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.685 $Y=1.35
+ $X2=1.685 $Y2=1.515
r36 15 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.685 $Y=1.35
+ $X2=1.685 $Y2=1.185
r37 10 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.685
+ $Y=1.35 $X2=1.685 $Y2=1.35
r38 9 10 14.4544 $w=2.93e-07 $l=3.7e-07 $layer=LI1_cond $X=1.677 $Y=0.925
+ $X2=1.677 $Y2=1.295
r39 8 9 14.4544 $w=2.93e-07 $l=3.7e-07 $layer=LI1_cond $X=1.677 $Y=0.555
+ $X2=1.677 $Y2=0.925
r40 6 18 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=1.665 $Y=2.465
+ $X2=1.665 $Y2=1.515
r41 3 17 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.595 $Y=0.655
+ $X2=1.595 $Y2=1.185
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4B_1%B 3 6 8 9 10 15 17
r40 15 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.225 $Y=1.35
+ $X2=2.225 $Y2=1.515
r41 15 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.225 $Y=1.35
+ $X2=2.225 $Y2=1.185
r42 10 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.225
+ $Y=1.35 $X2=2.225 $Y2=1.35
r43 9 10 10.795 $w=3.93e-07 $l=3.7e-07 $layer=LI1_cond $X=2.192 $Y=0.925
+ $X2=2.192 $Y2=1.295
r44 8 9 10.795 $w=3.93e-07 $l=3.7e-07 $layer=LI1_cond $X=2.192 $Y=0.555
+ $X2=2.192 $Y2=0.925
r45 6 18 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=2.245 $Y=2.465
+ $X2=2.245 $Y2=1.515
r46 3 17 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.135 $Y=0.655
+ $X2=2.135 $Y2=1.185
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4B_1%A_71_131# 1 2 9 13 16 17 21 22 27 33
c64 21 0 1.75712e-19 $X=2.765 $Y=1.51
r65 32 33 7.88995 $w=5.03e-07 $l=9.5e-08 $layer=LI1_cond $X=0.48 $Y=1.947
+ $X2=0.575 $Y2=1.947
r66 24 27 9.18462 $w=3.28e-07 $l=2.63e-07 $layer=LI1_cond $X=0.217 $Y=0.85
+ $X2=0.48 $Y2=0.85
r67 22 36 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.765 $Y=1.51
+ $X2=2.765 $Y2=1.675
r68 22 35 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.765 $Y=1.51
+ $X2=2.765 $Y2=1.345
r69 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.765
+ $Y=1.51 $X2=2.765 $Y2=1.51
r70 19 21 8.52808 $w=2.48e-07 $l=1.85e-07 $layer=LI1_cond $X=2.725 $Y=1.695
+ $X2=2.725 $Y2=1.51
r71 17 19 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.6 $Y=1.78
+ $X2=2.725 $Y2=1.695
r72 17 33 132.112 $w=1.68e-07 $l=2.025e-06 $layer=LI1_cond $X=2.6 $Y=1.78
+ $X2=0.575 $Y2=1.78
r73 16 32 6.22908 $w=5.03e-07 $l=2.63e-07 $layer=LI1_cond $X=0.217 $Y=1.947
+ $X2=0.48 $Y2=1.947
r74 15 24 2.04284 $w=2.65e-07 $l=1.65e-07 $layer=LI1_cond $X=0.217 $Y=1.015
+ $X2=0.217 $Y2=0.85
r75 15 16 29.5721 $w=2.63e-07 $l=6.8e-07 $layer=LI1_cond $X=0.217 $Y=1.015
+ $X2=0.217 $Y2=1.695
r76 13 36 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.675 $Y=2.465
+ $X2=2.675 $Y2=1.675
r77 9 35 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.675 $Y=0.655
+ $X2=2.675 $Y2=1.345
r78 2 32 600 $w=1.7e-07 $l=2.54951e-07 $layer=licon1_PDIFF $count=1 $X=0.355
+ $Y=1.835 $X2=0.48 $Y2=2.035
r79 1 27 182 $w=1.7e-07 $l=2.498e-07 $layer=licon1_NDIFF $count=1 $X=0.355
+ $Y=0.655 $X2=0.48 $Y2=0.85
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4B_1%VPWR 1 2 3 12 18 22 25 26 28 29 30 31 32 33
+ 47
r41 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r42 44 47 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r43 43 44 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r44 36 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r45 33 44 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r46 33 37 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.72 $Y2=3.33
r47 33 40 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r48 31 43 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=2.725 $Y=3.33
+ $X2=2.64 $Y2=3.33
r49 31 32 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.725 $Y=3.33
+ $X2=2.89 $Y2=3.33
r50 30 46 4.66471 $w=1.7e-07 $l=6.5e-08 $layer=LI1_cond $X=3.055 $Y=3.33
+ $X2=3.12 $Y2=3.33
r51 30 32 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.055 $Y=3.33
+ $X2=2.89 $Y2=3.33
r52 28 40 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=1.785 $Y=3.33
+ $X2=1.68 $Y2=3.33
r53 28 29 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.785 $Y=3.33
+ $X2=1.95 $Y2=3.33
r54 27 43 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=2.115 $Y=3.33
+ $X2=2.64 $Y2=3.33
r55 27 29 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.115 $Y=3.33
+ $X2=1.95 $Y2=3.33
r56 25 36 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=0.745 $Y=3.33
+ $X2=0.72 $Y2=3.33
r57 25 26 10.0494 $w=1.7e-07 $l=2.07e-07 $layer=LI1_cond $X=0.745 $Y=3.33
+ $X2=0.952 $Y2=3.33
r58 24 40 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=1.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r59 24 26 10.0494 $w=1.7e-07 $l=2.08e-07 $layer=LI1_cond $X=1.16 $Y=3.33
+ $X2=0.952 $Y2=3.33
r60 20 32 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.89 $Y=3.245
+ $X2=2.89 $Y2=3.33
r61 20 22 26.5411 $w=3.28e-07 $l=7.6e-07 $layer=LI1_cond $X=2.89 $Y=3.245
+ $X2=2.89 $Y2=2.485
r62 16 29 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.95 $Y=3.245
+ $X2=1.95 $Y2=3.33
r63 16 18 26.7157 $w=3.28e-07 $l=7.65e-07 $layer=LI1_cond $X=1.95 $Y=3.245
+ $X2=1.95 $Y2=2.48
r64 12 15 11.8021 $w=4.13e-07 $l=4.25e-07 $layer=LI1_cond $X=0.952 $Y=2.12
+ $X2=0.952 $Y2=2.545
r65 10 26 1.57254 $w=4.15e-07 $l=8.5e-08 $layer=LI1_cond $X=0.952 $Y=3.245
+ $X2=0.952 $Y2=3.33
r66 10 15 19.4388 $w=4.13e-07 $l=7e-07 $layer=LI1_cond $X=0.952 $Y=3.245
+ $X2=0.952 $Y2=2.545
r67 3 22 300 $w=1.7e-07 $l=7.16589e-07 $layer=licon1_PDIFF $count=2 $X=2.75
+ $Y=1.835 $X2=2.89 $Y2=2.485
r68 2 18 300 $w=1.7e-07 $l=7.42614e-07 $layer=licon1_PDIFF $count=2 $X=1.74
+ $Y=1.835 $X2=1.95 $Y2=2.48
r69 1 15 300 $w=1.7e-07 $l=8.25591e-07 $layer=licon1_PDIFF $count=2 $X=0.77
+ $Y=1.835 $X2=1.02 $Y2=2.545
r70 1 12 600 $w=1.7e-07 $l=3.4803e-07 $layer=licon1_PDIFF $count=1 $X=0.77
+ $Y=1.835 $X2=0.91 $Y2=2.12
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4B_1%Y 1 2 3 10 12 14 18 20 25 26 27 28 29 30 39
c47 20 0 2.4855e-20 $X=3.02 $Y=2.12
r48 29 30 14.7784 $w=2.53e-07 $l=3.27e-07 $layer=LI1_cond $X=3.147 $Y=1.665
+ $X2=3.147 $Y2=1.992
r49 28 29 16.7217 $w=2.53e-07 $l=3.7e-07 $layer=LI1_cond $X=3.147 $Y=1.295
+ $X2=3.147 $Y2=1.665
r50 28 54 9.03877 $w=2.53e-07 $l=2e-07 $layer=LI1_cond $X=3.147 $Y=1.295
+ $X2=3.147 $Y2=1.095
r51 27 54 7.16656 $w=5.48e-07 $l=1.7e-07 $layer=LI1_cond $X=3 $Y=0.925 $X2=3
+ $Y2=1.095
r52 27 37 2.28342 $w=5.48e-07 $l=1.05e-07 $layer=LI1_cond $X=3 $Y=0.925 $X2=3
+ $Y2=0.82
r53 26 37 5.76292 $w=5.48e-07 $l=2.65e-07 $layer=LI1_cond $X=3 $Y=0.555 $X2=3
+ $Y2=0.82
r54 26 39 2.93583 $w=5.48e-07 $l=1.35e-07 $layer=LI1_cond $X=3 $Y=0.555 $X2=3
+ $Y2=0.42
r55 21 25 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.555 $Y=2.12
+ $X2=2.425 $Y2=2.12
r56 20 30 4.29957 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=3.02 $Y=2.12
+ $X2=3.147 $Y2=2.12
r57 20 21 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=3.02 $Y=2.12
+ $X2=2.555 $Y2=2.12
r58 16 25 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=2.425 $Y=2.205
+ $X2=2.425 $Y2=2.12
r59 16 18 14.8488 $w=2.58e-07 $l=3.35e-07 $layer=LI1_cond $X=2.425 $Y=2.205
+ $X2=2.425 $Y2=2.54
r60 15 23 4.64039 $w=1.7e-07 $l=1.43e-07 $layer=LI1_cond $X=1.615 $Y=2.12
+ $X2=1.472 $Y2=2.12
r61 14 25 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.295 $Y=2.12
+ $X2=2.425 $Y2=2.12
r62 14 15 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=2.295 $Y=2.12
+ $X2=1.615 $Y2=2.12
r63 10 23 2.75828 $w=2.85e-07 $l=8.5e-08 $layer=LI1_cond $X=1.472 $Y=2.205
+ $X2=1.472 $Y2=2.12
r64 10 12 28.5078 $w=2.83e-07 $l=7.05e-07 $layer=LI1_cond $X=1.472 $Y=2.205
+ $X2=1.472 $Y2=2.91
r65 3 25 600 $w=1.7e-07 $l=3.4803e-07 $layer=licon1_PDIFF $count=1 $X=2.32
+ $Y=1.835 $X2=2.46 $Y2=2.12
r66 3 18 300 $w=1.7e-07 $l=7.71832e-07 $layer=licon1_PDIFF $count=2 $X=2.32
+ $Y=1.835 $X2=2.46 $Y2=2.54
r67 2 23 400 $w=1.7e-07 $l=4.29331e-07 $layer=licon1_PDIFF $count=1 $X=1.31
+ $Y=1.835 $X2=1.45 $Y2=2.2
r68 2 12 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=1.31
+ $Y=1.835 $X2=1.45 $Y2=2.91
r69 1 39 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=2.75
+ $Y=0.235 $X2=2.89 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4B_1%VGND 1 6 11 12 13 23 24
r32 23 24 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r33 20 23 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=3.12
+ $Y2=0
r34 20 21 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r35 17 21 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r36 16 17 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r37 13 24 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.68 $Y=0 $X2=3.12
+ $Y2=0
r38 13 21 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r39 11 16 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=0.795 $Y=0 $X2=0.72
+ $Y2=0
r40 11 12 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.795 $Y=0 $X2=0.96
+ $Y2=0
r41 10 20 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=1.125 $Y=0 $X2=1.2
+ $Y2=0
r42 10 12 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.125 $Y=0 $X2=0.96
+ $Y2=0
r43 6 8 17.9851 $w=3.28e-07 $l=5.15e-07 $layer=LI1_cond $X=0.96 $Y=0.38 $X2=0.96
+ $Y2=0.895
r44 4 12 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.96 $Y=0.085 $X2=0.96
+ $Y2=0
r45 4 6 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.96 $Y=0.085
+ $X2=0.96 $Y2=0.38
r46 1 8 182 $w=1.7e-07 $l=3.21248e-07 $layer=licon1_NDIFF $count=1 $X=0.77
+ $Y=0.655 $X2=0.96 $Y2=0.895
r47 1 6 182 $w=1.7e-07 $l=3.745e-07 $layer=licon1_NDIFF $count=1 $X=0.77
+ $Y=0.655 $X2=1.005 $Y2=0.38
.ends

