* File: sky130_fd_sc_lp__einvn_2.pex.spice
* Created: Wed Sep  2 09:51:39 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__EINVN_2%TE_B 3 5 6 8 9 11 12 13 14 16 21 22 26 28
r58 26 28 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=0.612 $Y=1.005
+ $X2=0.612 $Y2=0.84
r59 21 22 10.795 $w=3.93e-07 $l=3.7e-07 $layer=LI1_cond $X=0.747 $Y=0.925
+ $X2=0.747 $Y2=1.295
r60 21 26 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.635
+ $Y=1.005 $X2=0.635 $Y2=1.005
r61 14 16 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=1.455 $Y=1.725
+ $X2=1.455 $Y2=2.465
r62 13 20 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.1 $Y=1.65
+ $X2=1.025 $Y2=1.65
r63 12 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.38 $Y=1.65
+ $X2=1.455 $Y2=1.725
r64 12 13 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=1.38 $Y=1.65 $X2=1.1
+ $Y2=1.65
r65 9 20 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.025 $Y=1.725
+ $X2=1.025 $Y2=1.65
r66 9 11 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=1.025 $Y=1.725
+ $X2=1.025 $Y2=2.465
r67 6 17 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.5 $Y=1.725 $X2=0.5
+ $Y2=1.65
r68 6 8 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=0.5 $Y=1.725 $X2=0.5
+ $Y2=2.155
r69 5 20 211.772 $w=1.5e-07 $l=4.13e-07 $layer=POLY_cond $X=0.612 $Y=1.65
+ $X2=1.025 $Y2=1.65
r70 5 17 57.4298 $w=1.5e-07 $l=1.12e-07 $layer=POLY_cond $X=0.612 $Y=1.65
+ $X2=0.5 $Y2=1.65
r71 4 26 3.26277 $w=3.75e-07 $l=2.2e-08 $layer=POLY_cond $X=0.612 $Y=1.027
+ $X2=0.612 $Y2=1.005
r72 4 5 81.2726 $w=3.75e-07 $l=5.48e-07 $layer=POLY_cond $X=0.612 $Y=1.027
+ $X2=0.612 $Y2=1.575
r73 3 28 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.5 $Y=0.52 $X2=0.5
+ $Y2=0.84
.ends

.subckt PM_SKY130_FD_SC_LP__EINVN_2%A_28_62# 1 2 7 9 10 12 15 19 21 24 25 29 30
r62 30 34 14.3168 $w=3.03e-07 $l=9e-08 $layer=POLY_cond $X=1.935 $Y=1.395
+ $X2=2.025 $Y2=1.395
r63 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.935
+ $Y=1.44 $X2=1.935 $Y2=1.44
r64 26 29 4.66986 $w=1.88e-07 $l=8e-08 $layer=LI1_cond $X=1.855 $Y=1.44
+ $X2=1.935 $Y2=1.44
r65 23 26 1.386 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.855 $Y=1.535
+ $X2=1.855 $Y2=1.44
r66 23 24 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=1.855 $Y=1.535
+ $X2=1.855 $Y2=1.68
r67 22 25 3.44808 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.43 $Y=1.765
+ $X2=0.265 $Y2=1.765
r68 21 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.77 $Y=1.765
+ $X2=1.855 $Y2=1.68
r69 21 22 87.4225 $w=1.68e-07 $l=1.34e-06 $layer=LI1_cond $X=1.77 $Y=1.765
+ $X2=0.43 $Y2=1.765
r70 17 25 3.14896 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.265 $Y=1.85 $X2=0.265
+ $Y2=1.765
r71 17 19 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=0.265 $Y=1.85
+ $X2=0.265 $Y2=1.98
r72 13 25 3.14896 $w=3e-07 $l=9.88686e-08 $layer=LI1_cond $X=0.235 $Y=1.68
+ $X2=0.265 $Y2=1.765
r73 13 15 49.5124 $w=2.68e-07 $l=1.16e-06 $layer=LI1_cond $X=0.235 $Y=1.68
+ $X2=0.235 $Y2=0.52
r74 10 34 19.2026 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=2.025 $Y=1.185
+ $X2=2.025 $Y2=1.395
r75 10 12 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.025 $Y=1.185
+ $X2=2.025 $Y2=0.655
r76 7 30 54.0858 $w=3.03e-07 $l=4.32435e-07 $layer=POLY_cond $X=1.595 $Y=1.185
+ $X2=1.935 $Y2=1.395
r77 7 9 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.595 $Y=1.185
+ $X2=1.595 $Y2=0.655
r78 2 19 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.16
+ $Y=1.835 $X2=0.285 $Y2=1.98
r79 1 15 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.14
+ $Y=0.31 $X2=0.265 $Y2=0.52
.ends

.subckt PM_SKY130_FD_SC_LP__EINVN_2%A 3 7 9 13 16 18 19 22 24
r47 22 24 46.3655 $w=3.45e-07 $l=1.65e-07 $layer=POLY_cond $X=2.982 $Y=1.36
+ $X2=2.982 $Y2=1.195
r48 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.99
+ $Y=1.36 $X2=2.99 $Y2=1.36
r49 19 23 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=3.12 $Y=1.36
+ $X2=2.99 $Y2=1.36
r50 16 26 482 $w=1.5e-07 $l=9.4e-07 $layer=POLY_cond $X=2.885 $Y=2.465 $X2=2.885
+ $Y2=1.525
r51 13 24 173.52 $w=1.5e-07 $l=5.4e-07 $layer=POLY_cond $X=2.885 $Y=0.655
+ $X2=2.885 $Y2=1.195
r52 10 18 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.53 $Y=1.45
+ $X2=2.455 $Y2=1.45
r53 9 26 31.3122 $w=3.45e-07 $l=7.5e-08 $layer=POLY_cond $X=2.982 $Y=1.45
+ $X2=2.982 $Y2=1.525
r54 9 22 15.0533 $w=3.45e-07 $l=9e-08 $layer=POLY_cond $X=2.982 $Y=1.45
+ $X2=2.982 $Y2=1.36
r55 9 10 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.81 $Y=1.45 $X2=2.53
+ $Y2=1.45
r56 5 18 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.455 $Y=1.525
+ $X2=2.455 $Y2=1.45
r57 5 7 482 $w=1.5e-07 $l=9.4e-07 $layer=POLY_cond $X=2.455 $Y=1.525 $X2=2.455
+ $Y2=2.465
r58 1 18 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.455 $Y=1.375
+ $X2=2.455 $Y2=1.45
r59 1 3 369.191 $w=1.5e-07 $l=7.2e-07 $layer=POLY_cond $X=2.455 $Y=1.375
+ $X2=2.455 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__EINVN_2%VPWR 1 2 9 15 17 19 24 34 35 38 41
r45 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r46 34 35 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r47 32 35 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r48 31 34 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.16 $Y=3.33 $X2=3.12
+ $Y2=3.33
r49 31 32 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r50 29 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.835 $Y=3.33
+ $X2=1.67 $Y2=3.33
r51 29 31 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=1.835 $Y=3.33
+ $X2=2.16 $Y2=3.33
r52 28 39 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r53 27 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r54 25 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.93 $Y=3.33
+ $X2=0.765 $Y2=3.33
r55 25 27 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=0.93 $Y=3.33 $X2=1.2
+ $Y2=3.33
r56 24 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.505 $Y=3.33
+ $X2=1.67 $Y2=3.33
r57 24 27 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.505 $Y=3.33
+ $X2=1.2 $Y2=3.33
r58 22 39 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r59 21 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r60 19 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.6 $Y=3.33
+ $X2=0.765 $Y2=3.33
r61 19 21 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=0.6 $Y=3.33 $X2=0.24
+ $Y2=3.33
r62 17 32 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r63 17 28 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r64 17 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r65 13 41 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.67 $Y=3.245
+ $X2=1.67 $Y2=3.33
r66 13 15 15.8897 $w=3.28e-07 $l=4.55e-07 $layer=LI1_cond $X=1.67 $Y=3.245
+ $X2=1.67 $Y2=2.79
r67 9 12 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=0.765 $Y=2.105
+ $X2=0.765 $Y2=2.525
r68 7 38 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.765 $Y=3.245
+ $X2=0.765 $Y2=3.33
r69 7 12 25.1442 $w=3.28e-07 $l=7.2e-07 $layer=LI1_cond $X=0.765 $Y=3.245
+ $X2=0.765 $Y2=2.525
r70 2 15 600 $w=1.7e-07 $l=1.02261e-06 $layer=licon1_PDIFF $count=1 $X=1.53
+ $Y=1.835 $X2=1.67 $Y2=2.79
r71 1 12 300 $w=1.7e-07 $l=7.98906e-07 $layer=licon1_PDIFF $count=2 $X=0.575
+ $Y=1.835 $X2=0.81 $Y2=2.525
r72 1 9 600 $w=1.7e-07 $l=3.5242e-07 $layer=licon1_PDIFF $count=1 $X=0.575
+ $Y=1.835 $X2=0.765 $Y2=2.105
.ends

.subckt PM_SKY130_FD_SC_LP__EINVN_2%A_220_367# 1 2 9 11 15 19 22 26
c27 2 0 1.80713e-19 $X=2.53 $Y=1.835
r28 24 25 3.84843 $w=3.03e-07 $l=8.5e-08 $layer=LI1_cond $X=1.252 $Y=2.41
+ $X2=1.252 $Y2=2.495
r29 22 24 8.50163 $w=3.03e-07 $l=2.25e-07 $layer=LI1_cond $X=1.252 $Y=2.185
+ $X2=1.252 $Y2=2.41
r30 17 26 3.32435 $w=2.82e-07 $l=9.31128e-08 $layer=LI1_cond $X=2.672 $Y=2.325
+ $X2=2.655 $Y2=2.41
r31 17 19 5.00117 $w=2.63e-07 $l=1.15e-07 $layer=LI1_cond $X=2.672 $Y=2.325
+ $X2=2.672 $Y2=2.21
r32 13 26 3.32435 $w=2.82e-07 $l=8.5e-08 $layer=LI1_cond $X=2.655 $Y=2.495
+ $X2=2.655 $Y2=2.41
r33 13 15 2.49696 $w=2.98e-07 $l=6.5e-08 $layer=LI1_cond $X=2.655 $Y=2.495
+ $X2=2.655 $Y2=2.56
r34 12 24 4.15824 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=1.405 $Y=2.41
+ $X2=1.252 $Y2=2.41
r35 11 26 3.22099 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=2.505 $Y=2.41
+ $X2=2.655 $Y2=2.41
r36 11 12 71.7647 $w=1.68e-07 $l=1.1e-06 $layer=LI1_cond $X=2.505 $Y=2.41
+ $X2=1.405 $Y2=2.41
r37 9 25 2.45201 $w=2.33e-07 $l=5e-08 $layer=LI1_cond $X=1.217 $Y=2.545
+ $X2=1.217 $Y2=2.495
r38 2 19 600 $w=1.7e-07 $l=4.3946e-07 $layer=licon1_PDIFF $count=1 $X=2.53
+ $Y=1.835 $X2=2.67 $Y2=2.21
r39 2 15 300 $w=1.7e-07 $l=7.91912e-07 $layer=licon1_PDIFF $count=2 $X=2.53
+ $Y=1.835 $X2=2.67 $Y2=2.56
r40 1 22 600 $w=1.7e-07 $l=4.14126e-07 $layer=licon1_PDIFF $count=1 $X=1.1
+ $Y=1.835 $X2=1.24 $Y2=2.185
r41 1 9 300 $w=1.7e-07 $l=7.76853e-07 $layer=licon1_PDIFF $count=2 $X=1.1
+ $Y=1.835 $X2=1.24 $Y2=2.545
.ends

.subckt PM_SKY130_FD_SC_LP__EINVN_2%Z 1 2 3 12 14 15 18 22 23 24 33 39 41
c44 14 0 1.80713e-19 $X=2.975 $Y=1.79
r45 33 44 1.92074 $w=2.38e-07 $l=4e-08 $layer=LI1_cond $X=2.615 $Y=0.925
+ $X2=2.615 $Y2=0.885
r46 31 39 1.92074 $w=2.38e-07 $l=4e-08 $layer=LI1_cond $X=2.615 $Y=1.705
+ $X2=2.615 $Y2=1.665
r47 24 31 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=2.64 $Y=1.79
+ $X2=2.615 $Y2=1.79
r48 24 39 1.10442 $w=2.38e-07 $l=2.3e-08 $layer=LI1_cond $X=2.615 $Y=1.642
+ $X2=2.615 $Y2=1.665
r49 23 24 16.6624 $w=2.38e-07 $l=3.47e-07 $layer=LI1_cond $X=2.615 $Y=1.295
+ $X2=2.615 $Y2=1.642
r50 22 44 1.79124 $w=3.38e-07 $l=2.3e-08 $layer=LI1_cond $X=2.665 $Y=0.862
+ $X2=2.665 $Y2=0.885
r51 22 41 4.81314 $w=3.38e-07 $l=1.42e-07 $layer=LI1_cond $X=2.665 $Y=0.862
+ $X2=2.665 $Y2=0.72
r52 22 23 16.7104 $w=2.38e-07 $l=3.48e-07 $layer=LI1_cond $X=2.615 $Y=0.947
+ $X2=2.615 $Y2=1.295
r53 22 33 1.05641 $w=2.38e-07 $l=2.2e-08 $layer=LI1_cond $X=2.615 $Y=0.947
+ $X2=2.615 $Y2=0.925
r54 18 20 36.9577 $w=2.88e-07 $l=9.3e-07 $layer=LI1_cond $X=3.12 $Y=1.98
+ $X2=3.12 $Y2=2.91
r55 16 18 4.17264 $w=2.88e-07 $l=1.05e-07 $layer=LI1_cond $X=3.12 $Y=1.875
+ $X2=3.12 $Y2=1.98
r56 15 24 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=2.735 $Y=1.79
+ $X2=2.64 $Y2=1.79
r57 14 16 7.43784 $w=1.7e-07 $l=1.8262e-07 $layer=LI1_cond $X=2.975 $Y=1.79
+ $X2=3.12 $Y2=1.875
r58 14 15 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=2.975 $Y=1.79
+ $X2=2.735 $Y2=1.79
r59 10 31 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=2.24 $Y=1.79
+ $X2=2.615 $Y2=1.79
r60 10 12 5.09734 $w=2.58e-07 $l=1.15e-07 $layer=LI1_cond $X=2.24 $Y=1.875
+ $X2=2.24 $Y2=1.99
r61 3 20 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=2.96
+ $Y=1.835 $X2=3.1 $Y2=2.91
r62 3 18 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.96
+ $Y=1.835 $X2=3.1 $Y2=1.98
r63 2 12 600 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_PDIFF $count=1 $X=2.115
+ $Y=1.835 $X2=2.24 $Y2=1.99
r64 1 41 182 $w=1.7e-07 $l=5.50568e-07 $layer=licon1_NDIFF $count=1 $X=2.53
+ $Y=0.235 $X2=2.67 $Y2=0.72
.ends

.subckt PM_SKY130_FD_SC_LP__EINVN_2%VGND 1 2 9 11 15 17 19 29 30 33 36
r43 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r44 29 30 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r45 27 30 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r46 26 29 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r47 26 27 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r48 24 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.975 $Y=0 $X2=1.81
+ $Y2=0
r49 24 26 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=1.975 $Y=0 $X2=2.16
+ $Y2=0
r50 22 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r51 21 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r52 19 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.55 $Y=0 $X2=0.715
+ $Y2=0
r53 19 21 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=0.55 $Y=0 $X2=0.24
+ $Y2=0
r54 17 27 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r55 17 34 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=0.72
+ $Y2=0
r56 17 36 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r57 13 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.81 $Y=0.085
+ $X2=1.81 $Y2=0
r58 13 15 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.81 $Y=0.085
+ $X2=1.81 $Y2=0.38
r59 12 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.88 $Y=0 $X2=0.715
+ $Y2=0
r60 11 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.645 $Y=0 $X2=1.81
+ $Y2=0
r61 11 12 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=1.645 $Y=0 $X2=0.88
+ $Y2=0
r62 7 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.715 $Y=0.085
+ $X2=0.715 $Y2=0
r63 7 9 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.715 $Y=0.085
+ $X2=0.715 $Y2=0.455
r64 2 15 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.67
+ $Y=0.235 $X2=1.81 $Y2=0.38
r65 1 9 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=0.575
+ $Y=0.31 $X2=0.715 $Y2=0.455
.ends

.subckt PM_SKY130_FD_SC_LP__EINVN_2%A_251_47# 1 2 3 12 14 15 16 18 25
r40 19 23 3.50935 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=2.325 $Y=0.34 $X2=2.235
+ $Y2=0.34
r41 18 25 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.005 $Y=0.34
+ $X2=3.135 $Y2=0.34
r42 18 19 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=3.005 $Y=0.34
+ $X2=2.325 $Y2=0.34
r43 16 23 3.31438 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.235 $Y=0.425
+ $X2=2.235 $Y2=0.34
r44 16 17 35.7374 $w=1.78e-07 $l=5.8e-07 $layer=LI1_cond $X=2.235 $Y=0.425
+ $X2=2.235 $Y2=1.005
r45 14 17 6.82373 $w=1.7e-07 $l=1.25499e-07 $layer=LI1_cond $X=2.145 $Y=1.09
+ $X2=2.235 $Y2=1.005
r46 14 15 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.145 $Y=1.09
+ $X2=1.475 $Y2=1.09
r47 10 15 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=1.345 $Y=1.005
+ $X2=1.475 $Y2=1.09
r48 10 12 25.93 $w=2.58e-07 $l=5.85e-07 $layer=LI1_cond $X=1.345 $Y=1.005
+ $X2=1.345 $Y2=0.42
r49 3 25 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=2.96
+ $Y=0.235 $X2=3.1 $Y2=0.42
r50 2 23 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=2.1
+ $Y=0.235 $X2=2.24 $Y2=0.42
r51 1 12 91 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=2 $X=1.255
+ $Y=0.235 $X2=1.38 $Y2=0.42
.ends

