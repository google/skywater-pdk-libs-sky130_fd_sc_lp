* File: sky130_fd_sc_lp__o2bb2ai_1.pxi.spice
* Created: Wed Sep  2 10:22:09 2020
* 
x_PM_SKY130_FD_SC_LP__O2BB2AI_1%A1_N N_A1_N_M1003_g N_A1_N_M1005_g A1_N A1_N
+ N_A1_N_c_67_n N_A1_N_c_68_n PM_SKY130_FD_SC_LP__O2BB2AI_1%A1_N
x_PM_SKY130_FD_SC_LP__O2BB2AI_1%A2_N N_A2_N_M1009_g N_A2_N_M1007_g A2_N
+ N_A2_N_c_92_n N_A2_N_c_93_n N_A2_N_c_94_n PM_SKY130_FD_SC_LP__O2BB2AI_1%A2_N
x_PM_SKY130_FD_SC_LP__O2BB2AI_1%A_115_367# N_A_115_367#_M1009_d
+ N_A_115_367#_M1005_d N_A_115_367#_M1004_g N_A_115_367#_M1001_g
+ N_A_115_367#_c_126_n N_A_115_367#_c_127_n N_A_115_367#_c_171_p
+ N_A_115_367#_c_136_n N_A_115_367#_c_137_n N_A_115_367#_c_128_n
+ N_A_115_367#_c_129_n N_A_115_367#_c_130_n N_A_115_367#_c_131_n
+ N_A_115_367#_c_132_n PM_SKY130_FD_SC_LP__O2BB2AI_1%A_115_367#
x_PM_SKY130_FD_SC_LP__O2BB2AI_1%B2 N_B2_M1006_g N_B2_M1002_g B2 B2 B2 B2
+ N_B2_c_202_n B2 PM_SKY130_FD_SC_LP__O2BB2AI_1%B2
x_PM_SKY130_FD_SC_LP__O2BB2AI_1%B1 N_B1_M1008_g N_B1_M1000_g B1 B1 N_B1_c_246_n
+ PM_SKY130_FD_SC_LP__O2BB2AI_1%B1
x_PM_SKY130_FD_SC_LP__O2BB2AI_1%VPWR N_VPWR_M1005_s N_VPWR_M1007_d
+ N_VPWR_M1000_d N_VPWR_c_271_n N_VPWR_c_272_n N_VPWR_c_273_n N_VPWR_c_274_n
+ N_VPWR_c_275_n VPWR N_VPWR_c_276_n N_VPWR_c_277_n N_VPWR_c_278_n
+ N_VPWR_c_270_n PM_SKY130_FD_SC_LP__O2BB2AI_1%VPWR
x_PM_SKY130_FD_SC_LP__O2BB2AI_1%Y N_Y_M1004_s N_Y_M1001_d N_Y_c_316_n
+ N_Y_c_317_n N_Y_c_321_n Y Y Y Y Y N_Y_c_319_n PM_SKY130_FD_SC_LP__O2BB2AI_1%Y
x_PM_SKY130_FD_SC_LP__O2BB2AI_1%VGND N_VGND_M1003_s N_VGND_M1006_d
+ N_VGND_c_357_n N_VGND_c_358_n N_VGND_c_359_n VGND N_VGND_c_360_n
+ N_VGND_c_361_n N_VGND_c_362_n N_VGND_c_363_n
+ PM_SKY130_FD_SC_LP__O2BB2AI_1%VGND
x_PM_SKY130_FD_SC_LP__O2BB2AI_1%A_396_47# N_A_396_47#_M1004_d
+ N_A_396_47#_M1008_d N_A_396_47#_c_401_n N_A_396_47#_c_398_n
+ N_A_396_47#_c_399_n N_A_396_47#_c_400_n
+ PM_SKY130_FD_SC_LP__O2BB2AI_1%A_396_47#
cc_1 VNB N_A1_N_M1005_g 0.00726307f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=2.465
cc_2 VNB A1_N 0.0210144f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_3 VNB N_A1_N_c_67_n 0.0408688f $X=-0.19 $Y=-0.245 $X2=0.365 $Y2=1.375
cc_4 VNB N_A1_N_c_68_n 0.0208407f $X=-0.19 $Y=-0.245 $X2=0.387 $Y2=1.21
cc_5 VNB N_A2_N_M1007_g 0.00668675f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=2.465
cc_6 VNB N_A2_N_c_92_n 0.0352178f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_A2_N_c_93_n 0.00951551f $X=-0.19 $Y=-0.245 $X2=0.387 $Y2=1.375
cc_8 VNB N_A2_N_c_94_n 0.0192405f $X=-0.19 $Y=-0.245 $X2=0.365 $Y2=1.375
cc_9 VNB N_A_115_367#_M1004_g 0.0252453f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_10 VNB N_A_115_367#_c_126_n 0.0341923f $X=-0.19 $Y=-0.245 $X2=0.387 $Y2=1.21
cc_11 VNB N_A_115_367#_c_127_n 0.0121053f $X=-0.19 $Y=-0.245 $X2=0.387 $Y2=1.54
cc_12 VNB N_A_115_367#_c_128_n 0.00770517f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_115_367#_c_129_n 0.00425982f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_115_367#_c_130_n 0.00106797f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_115_367#_c_131_n 0.00355209f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_115_367#_c_132_n 0.00638668f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_B2_M1006_g 0.0188208f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=0.68
cc_18 VNB N_B2_M1002_g 0.0055253f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB B2 0.00782114f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_20 VNB N_B2_c_202_n 0.033349f $X=-0.19 $Y=-0.245 $X2=0.267 $Y2=1.665
cc_21 VNB B2 9.59021e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_B1_M1008_g 0.0248658f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=0.68
cc_23 VNB N_B1_M1000_g 0.00716568f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB B1 0.0217681f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_25 VNB N_B1_c_246_n 0.0399602f $X=-0.19 $Y=-0.245 $X2=0.365 $Y2=1.375
cc_26 VNB N_VPWR_c_270_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_Y_c_316_n 0.00564492f $X=-0.19 $Y=-0.245 $X2=0.387 $Y2=1.375
cc_28 VNB N_Y_c_317_n 0.00322053f $X=-0.19 $Y=-0.245 $X2=0.387 $Y2=1.21
cc_29 VNB Y 0.00360025f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_Y_c_319_n 0.00433849f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_357_n 0.0113527f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_358_n 0.0345158f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_33 VNB N_VGND_c_359_n 0.00557258f $X=-0.19 $Y=-0.245 $X2=0.365 $Y2=1.375
cc_34 VNB N_VGND_c_360_n 0.0537891f $X=-0.19 $Y=-0.245 $X2=0.267 $Y2=1.295
cc_35 VNB N_VGND_c_361_n 0.0172175f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_362_n 0.210385f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_363_n 0.00631953f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_396_47#_c_398_n 0.0126149f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_39 VNB N_A_396_47#_c_399_n 0.0176418f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VPB N_A1_N_M1005_g 0.0255057f $X=-0.19 $Y=1.655 $X2=0.5 $Y2=2.465
cc_41 VPB A1_N 0.00798479f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_42 VPB N_A2_N_M1007_g 0.0228385f $X=-0.19 $Y=1.655 $X2=0.5 $Y2=2.465
cc_43 VPB N_A_115_367#_M1001_g 0.0231482f $X=-0.19 $Y=1.655 $X2=0.365 $Y2=1.375
cc_44 VPB N_A_115_367#_c_126_n 0.0131316f $X=-0.19 $Y=1.655 $X2=0.387 $Y2=1.21
cc_45 VPB N_A_115_367#_c_127_n 0.0023656f $X=-0.19 $Y=1.655 $X2=0.387 $Y2=1.54
cc_46 VPB N_A_115_367#_c_136_n 0.0038924f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_47 VPB N_A_115_367#_c_137_n 0.00296539f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_48 VPB N_A_115_367#_c_129_n 0.00316862f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_49 VPB N_A_115_367#_c_130_n 2.43024e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_50 VPB N_B2_M1002_g 0.0201778f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_51 VPB B2 0.00145512f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_52 VPB N_B1_M1000_g 0.0253554f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_53 VPB B1 0.00779597f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_54 VPB N_VPWR_c_271_n 0.0111372f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_55 VPB N_VPWR_c_272_n 0.0483629f $X=-0.19 $Y=1.655 $X2=0.387 $Y2=1.375
cc_56 VPB N_VPWR_c_273_n 0.00552031f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_57 VPB N_VPWR_c_274_n 0.0109777f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_58 VPB N_VPWR_c_275_n 0.0484529f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_59 VPB N_VPWR_c_276_n 0.0129398f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_60 VPB N_VPWR_c_277_n 0.0285511f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_61 VPB N_VPWR_c_278_n 0.0149019f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_62 VPB N_VPWR_c_270_n 0.0453059f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_63 VPB N_Y_c_317_n 8.50753e-19 $X=-0.19 $Y=1.655 $X2=0.387 $Y2=1.21
cc_64 VPB N_Y_c_321_n 0.00699933f $X=-0.19 $Y=1.655 $X2=0.387 $Y2=1.54
cc_65 N_A1_N_M1005_g N_A2_N_M1007_g 0.0240654f $X=0.5 $Y=2.465 $X2=0 $Y2=0
cc_66 A1_N N_A2_N_M1007_g 0.0010177f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_67 A1_N N_A2_N_c_92_n 2.51383e-19 $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_68 N_A1_N_c_67_n N_A2_N_c_92_n 0.0424883f $X=0.365 $Y=1.375 $X2=0 $Y2=0
cc_69 A1_N N_A2_N_c_93_n 0.0261495f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_70 N_A1_N_c_67_n N_A2_N_c_93_n 0.00248716f $X=0.365 $Y=1.375 $X2=0 $Y2=0
cc_71 N_A1_N_c_68_n N_A2_N_c_94_n 0.0424883f $X=0.387 $Y=1.21 $X2=0 $Y2=0
cc_72 N_A1_N_M1005_g N_A_115_367#_c_137_n 0.00243507f $X=0.5 $Y=2.465 $X2=0
+ $Y2=0
cc_73 N_A1_N_c_68_n N_A_115_367#_c_129_n 5.21768e-19 $X=0.387 $Y=1.21 $X2=0
+ $Y2=0
cc_74 N_A1_N_M1005_g N_VPWR_c_272_n 0.0203566f $X=0.5 $Y=2.465 $X2=0 $Y2=0
cc_75 A1_N N_VPWR_c_272_n 0.026915f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_76 N_A1_N_c_67_n N_VPWR_c_272_n 9.85169e-19 $X=0.365 $Y=1.375 $X2=0 $Y2=0
cc_77 N_A1_N_M1005_g N_VPWR_c_273_n 7.40603e-19 $X=0.5 $Y=2.465 $X2=0 $Y2=0
cc_78 N_A1_N_M1005_g N_VPWR_c_276_n 0.00486043f $X=0.5 $Y=2.465 $X2=0 $Y2=0
cc_79 N_A1_N_M1005_g N_VPWR_c_270_n 0.0082726f $X=0.5 $Y=2.465 $X2=0 $Y2=0
cc_80 A1_N N_VGND_c_358_n 0.0259278f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_81 N_A1_N_c_67_n N_VGND_c_358_n 0.00160808f $X=0.365 $Y=1.375 $X2=0 $Y2=0
cc_82 N_A1_N_c_68_n N_VGND_c_358_n 0.0221448f $X=0.387 $Y=1.21 $X2=0 $Y2=0
cc_83 N_A1_N_c_68_n N_VGND_c_360_n 0.00465098f $X=0.387 $Y=1.21 $X2=0 $Y2=0
cc_84 N_A1_N_c_68_n N_VGND_c_362_n 0.00808963f $X=0.387 $Y=1.21 $X2=0 $Y2=0
cc_85 N_A2_N_c_92_n N_A_115_367#_M1004_g 7.57158e-19 $X=0.95 $Y=1.375 $X2=0
+ $Y2=0
cc_86 N_A2_N_M1007_g N_A_115_367#_c_126_n 0.0030583f $X=0.93 $Y=2.465 $X2=0
+ $Y2=0
cc_87 N_A2_N_c_92_n N_A_115_367#_c_126_n 0.0104662f $X=0.95 $Y=1.375 $X2=0 $Y2=0
cc_88 N_A2_N_M1007_g N_A_115_367#_c_136_n 0.0143552f $X=0.93 $Y=2.465 $X2=0
+ $Y2=0
cc_89 N_A2_N_c_92_n N_A_115_367#_c_136_n 0.00573545f $X=0.95 $Y=1.375 $X2=0
+ $Y2=0
cc_90 N_A2_N_c_93_n N_A_115_367#_c_136_n 0.0135725f $X=0.95 $Y=1.375 $X2=0 $Y2=0
cc_91 N_A2_N_c_92_n N_A_115_367#_c_137_n 6.62823e-19 $X=0.95 $Y=1.375 $X2=0
+ $Y2=0
cc_92 N_A2_N_c_93_n N_A_115_367#_c_137_n 0.0137652f $X=0.95 $Y=1.375 $X2=0 $Y2=0
cc_93 N_A2_N_c_94_n N_A_115_367#_c_128_n 0.0151547f $X=0.965 $Y=1.21 $X2=0 $Y2=0
cc_94 N_A2_N_M1007_g N_A_115_367#_c_129_n 0.0064995f $X=0.93 $Y=2.465 $X2=0
+ $Y2=0
cc_95 N_A2_N_c_92_n N_A_115_367#_c_131_n 0.00608668f $X=0.95 $Y=1.375 $X2=0
+ $Y2=0
cc_96 N_A2_N_c_93_n N_A_115_367#_c_131_n 0.00377717f $X=0.95 $Y=1.375 $X2=0
+ $Y2=0
cc_97 N_A2_N_c_92_n N_A_115_367#_c_132_n 0.00306048f $X=0.95 $Y=1.375 $X2=0
+ $Y2=0
cc_98 N_A2_N_c_93_n N_A_115_367#_c_132_n 0.0253128f $X=0.95 $Y=1.375 $X2=0 $Y2=0
cc_99 N_A2_N_c_94_n N_A_115_367#_c_132_n 0.00519821f $X=0.965 $Y=1.21 $X2=0
+ $Y2=0
cc_100 N_A2_N_M1007_g N_VPWR_c_272_n 7.75547e-19 $X=0.93 $Y=2.465 $X2=0 $Y2=0
cc_101 N_A2_N_M1007_g N_VPWR_c_273_n 0.0161485f $X=0.93 $Y=2.465 $X2=0 $Y2=0
cc_102 N_A2_N_M1007_g N_VPWR_c_276_n 0.00486043f $X=0.93 $Y=2.465 $X2=0 $Y2=0
cc_103 N_A2_N_M1007_g N_VPWR_c_270_n 0.0082726f $X=0.93 $Y=2.465 $X2=0 $Y2=0
cc_104 N_A2_N_c_94_n N_VGND_c_358_n 0.00324664f $X=0.965 $Y=1.21 $X2=0 $Y2=0
cc_105 N_A2_N_c_94_n N_VGND_c_360_n 0.00560159f $X=0.965 $Y=1.21 $X2=0 $Y2=0
cc_106 N_A2_N_c_94_n N_VGND_c_362_n 0.0117172f $X=0.965 $Y=1.21 $X2=0 $Y2=0
cc_107 N_A_115_367#_M1004_g N_B2_M1006_g 0.0183171f $X=1.905 $Y=0.655 $X2=0
+ $Y2=0
cc_108 N_A_115_367#_c_127_n N_B2_M1002_g 0.0312909f $X=1.83 $Y=1.285 $X2=0 $Y2=0
cc_109 N_A_115_367#_M1004_g B2 2.20288e-19 $X=1.905 $Y=0.655 $X2=0 $Y2=0
cc_110 N_A_115_367#_c_127_n B2 2.42453e-19 $X=1.83 $Y=1.285 $X2=0 $Y2=0
cc_111 N_A_115_367#_M1004_g N_B2_c_202_n 0.011827f $X=1.905 $Y=0.655 $X2=0 $Y2=0
cc_112 N_A_115_367#_c_127_n N_B2_c_202_n 0.00658093f $X=1.83 $Y=1.285 $X2=0
+ $Y2=0
cc_113 N_A_115_367#_c_127_n B2 5.47237e-19 $X=1.83 $Y=1.285 $X2=0 $Y2=0
cc_114 N_A_115_367#_c_136_n N_VPWR_M1007_d 0.00186704f $X=1.205 $Y=1.84 $X2=0
+ $Y2=0
cc_115 N_A_115_367#_c_129_n N_VPWR_M1007_d 0.00474727f $X=1.415 $Y=1.54 $X2=0
+ $Y2=0
cc_116 N_A_115_367#_M1001_g N_VPWR_c_273_n 0.00495914f $X=1.935 $Y=2.465 $X2=0
+ $Y2=0
cc_117 N_A_115_367#_c_126_n N_VPWR_c_273_n 0.00851455f $X=1.83 $Y=1.48 $X2=0
+ $Y2=0
cc_118 N_A_115_367#_c_136_n N_VPWR_c_273_n 0.0134204f $X=1.205 $Y=1.84 $X2=0
+ $Y2=0
cc_119 N_A_115_367#_c_129_n N_VPWR_c_273_n 0.0186851f $X=1.415 $Y=1.54 $X2=0
+ $Y2=0
cc_120 N_A_115_367#_c_130_n N_VPWR_c_273_n 0.0140517f $X=1.595 $Y=1.51 $X2=0
+ $Y2=0
cc_121 N_A_115_367#_c_171_p N_VPWR_c_276_n 0.0124525f $X=0.715 $Y=1.98 $X2=0
+ $Y2=0
cc_122 N_A_115_367#_M1001_g N_VPWR_c_277_n 0.0055654f $X=1.935 $Y=2.465 $X2=0
+ $Y2=0
cc_123 N_A_115_367#_M1005_d N_VPWR_c_270_n 0.00536646f $X=0.575 $Y=1.835 $X2=0
+ $Y2=0
cc_124 N_A_115_367#_M1001_g N_VPWR_c_270_n 0.0114432f $X=1.935 $Y=2.465 $X2=0
+ $Y2=0
cc_125 N_A_115_367#_c_171_p N_VPWR_c_270_n 0.00730901f $X=0.715 $Y=1.98 $X2=0
+ $Y2=0
cc_126 N_A_115_367#_M1004_g N_Y_c_316_n 0.0168876f $X=1.905 $Y=0.655 $X2=0 $Y2=0
cc_127 N_A_115_367#_c_126_n N_Y_c_316_n 0.00878963f $X=1.83 $Y=1.48 $X2=0 $Y2=0
cc_128 N_A_115_367#_c_130_n N_Y_c_316_n 0.0159122f $X=1.595 $Y=1.51 $X2=0 $Y2=0
cc_129 N_A_115_367#_c_132_n N_Y_c_316_n 0.0139533f $X=1.31 $Y=1.405 $X2=0 $Y2=0
cc_130 N_A_115_367#_M1004_g N_Y_c_317_n 0.00150192f $X=1.905 $Y=0.655 $X2=0
+ $Y2=0
cc_131 N_A_115_367#_M1001_g N_Y_c_317_n 0.00237946f $X=1.935 $Y=2.465 $X2=0
+ $Y2=0
cc_132 N_A_115_367#_c_127_n N_Y_c_317_n 0.0118133f $X=1.83 $Y=1.285 $X2=0 $Y2=0
cc_133 N_A_115_367#_c_129_n N_Y_c_317_n 0.00815923f $X=1.415 $Y=1.54 $X2=0 $Y2=0
cc_134 N_A_115_367#_c_130_n N_Y_c_317_n 0.0193074f $X=1.595 $Y=1.51 $X2=0 $Y2=0
cc_135 N_A_115_367#_c_132_n N_Y_c_317_n 0.0049394f $X=1.31 $Y=1.405 $X2=0 $Y2=0
cc_136 N_A_115_367#_M1001_g N_Y_c_321_n 0.0079581f $X=1.935 $Y=2.465 $X2=0 $Y2=0
cc_137 N_A_115_367#_c_128_n Y 0.0111256f $X=1.15 $Y=0.405 $X2=0 $Y2=0
cc_138 N_A_115_367#_c_131_n Y 0.0200176f $X=1.18 $Y=1.04 $X2=0 $Y2=0
cc_139 N_A_115_367#_M1001_g Y 0.0194399f $X=1.935 $Y=2.465 $X2=0 $Y2=0
cc_140 N_A_115_367#_c_126_n N_Y_c_319_n 4.94824e-19 $X=1.83 $Y=1.48 $X2=0 $Y2=0
cc_141 N_A_115_367#_c_128_n N_Y_c_319_n 0.0278617f $X=1.15 $Y=0.405 $X2=0 $Y2=0
cc_142 N_A_115_367#_c_128_n N_VGND_c_358_n 0.0115796f $X=1.15 $Y=0.405 $X2=0
+ $Y2=0
cc_143 N_A_115_367#_M1004_g N_VGND_c_360_n 0.00548467f $X=1.905 $Y=0.655 $X2=0
+ $Y2=0
cc_144 N_A_115_367#_c_128_n N_VGND_c_360_n 0.0235133f $X=1.15 $Y=0.405 $X2=0
+ $Y2=0
cc_145 N_A_115_367#_M1004_g N_VGND_c_362_n 0.0112021f $X=1.905 $Y=0.655 $X2=0
+ $Y2=0
cc_146 N_A_115_367#_c_128_n N_VGND_c_362_n 0.0127519f $X=1.15 $Y=0.405 $X2=0
+ $Y2=0
cc_147 N_A_115_367#_c_131_n N_VGND_c_362_n 0.00236759f $X=1.18 $Y=1.04 $X2=0
+ $Y2=0
cc_148 N_A_115_367#_M1004_g N_A_396_47#_c_400_n 0.00746708f $X=1.905 $Y=0.655
+ $X2=0 $Y2=0
cc_149 N_B2_M1006_g N_B1_M1008_g 0.0275214f $X=2.335 $Y=0.655 $X2=0 $Y2=0
cc_150 B2 N_B1_M1008_g 0.00296649f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_151 N_B2_M1002_g N_B1_M1000_g 0.0722606f $X=2.445 $Y=2.465 $X2=0 $Y2=0
cc_152 B2 N_B1_M1000_g 0.00800845f $X=2.64 $Y=1.665 $X2=0 $Y2=0
cc_153 B2 B1 0.0323572f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_154 N_B2_c_202_n B1 2.57343e-19 $X=2.415 $Y=1.375 $X2=0 $Y2=0
cc_155 B2 B1 0.0128002f $X=2.64 $Y=1.665 $X2=0 $Y2=0
cc_156 N_B2_c_202_n N_B1_c_246_n 0.0205292f $X=2.415 $Y=1.375 $X2=0 $Y2=0
cc_157 N_B2_M1002_g N_VPWR_c_275_n 0.00219712f $X=2.445 $Y=2.465 $X2=0 $Y2=0
cc_158 N_B2_M1002_g N_VPWR_c_277_n 0.00565642f $X=2.445 $Y=2.465 $X2=0 $Y2=0
cc_159 B2 N_VPWR_c_277_n 0.0092441f $X=2.64 $Y=1.665 $X2=0 $Y2=0
cc_160 N_B2_M1002_g N_VPWR_c_270_n 0.0106888f $X=2.445 $Y=2.465 $X2=0 $Y2=0
cc_161 B2 N_VPWR_c_270_n 0.00842255f $X=2.64 $Y=1.665 $X2=0 $Y2=0
cc_162 N_B2_M1006_g N_Y_c_316_n 0.00334594f $X=2.335 $Y=0.655 $X2=0 $Y2=0
cc_163 B2 N_Y_c_316_n 0.00320024f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_164 N_B2_M1002_g N_Y_c_317_n 0.00141255f $X=2.445 $Y=2.465 $X2=0 $Y2=0
cc_165 B2 N_Y_c_317_n 0.0215085f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_166 N_B2_c_202_n N_Y_c_317_n 0.00211956f $X=2.415 $Y=1.375 $X2=0 $Y2=0
cc_167 B2 N_Y_c_317_n 0.0064823f $X=2.64 $Y=1.665 $X2=0 $Y2=0
cc_168 N_B2_M1002_g N_Y_c_321_n 0.00747352f $X=2.445 $Y=2.465 $X2=0 $Y2=0
cc_169 N_B2_c_202_n N_Y_c_321_n 0.00492039f $X=2.415 $Y=1.375 $X2=0 $Y2=0
cc_170 B2 N_Y_c_321_n 0.0474129f $X=2.64 $Y=1.665 $X2=0 $Y2=0
cc_171 B2 A_504_367# 0.00388106f $X=2.64 $Y=1.665 $X2=-0.19 $Y2=-0.245
cc_172 N_B2_M1006_g N_VGND_c_359_n 0.00489332f $X=2.335 $Y=0.655 $X2=0 $Y2=0
cc_173 N_B2_M1006_g N_VGND_c_360_n 0.00425523f $X=2.335 $Y=0.655 $X2=0 $Y2=0
cc_174 N_B2_M1006_g N_VGND_c_362_n 0.0061834f $X=2.335 $Y=0.655 $X2=0 $Y2=0
cc_175 N_B2_M1006_g N_A_396_47#_c_401_n 0.0138372f $X=2.335 $Y=0.655 $X2=0 $Y2=0
cc_176 B2 N_A_396_47#_c_401_n 0.0304292f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_177 N_B2_c_202_n N_A_396_47#_c_401_n 0.00101998f $X=2.415 $Y=1.375 $X2=0
+ $Y2=0
cc_178 N_B2_M1006_g N_A_396_47#_c_400_n 0.00946263f $X=2.335 $Y=0.655 $X2=0
+ $Y2=0
cc_179 N_B1_M1000_g N_VPWR_c_275_n 0.0224615f $X=2.865 $Y=2.465 $X2=0 $Y2=0
cc_180 B1 N_VPWR_c_275_n 0.0270157f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_181 N_B1_c_246_n N_VPWR_c_275_n 9.3623e-19 $X=2.99 $Y=1.375 $X2=0 $Y2=0
cc_182 N_B1_M1000_g N_VPWR_c_277_n 0.00486043f $X=2.865 $Y=2.465 $X2=0 $Y2=0
cc_183 N_B1_M1000_g N_VPWR_c_270_n 0.00835595f $X=2.865 $Y=2.465 $X2=0 $Y2=0
cc_184 N_B1_M1008_g N_VGND_c_359_n 0.00336601f $X=2.865 $Y=0.655 $X2=0 $Y2=0
cc_185 N_B1_M1008_g N_VGND_c_361_n 0.00437852f $X=2.865 $Y=0.655 $X2=0 $Y2=0
cc_186 N_B1_M1008_g N_VGND_c_362_n 0.00703555f $X=2.865 $Y=0.655 $X2=0 $Y2=0
cc_187 N_B1_M1008_g N_A_396_47#_c_401_n 0.0181948f $X=2.865 $Y=0.655 $X2=0 $Y2=0
cc_188 B1 N_A_396_47#_c_401_n 0.00420013f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_189 B1 N_A_396_47#_c_398_n 0.0235522f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_190 N_B1_c_246_n N_A_396_47#_c_398_n 0.00126577f $X=2.99 $Y=1.375 $X2=0 $Y2=0
cc_191 N_B1_M1008_g N_A_396_47#_c_400_n 6.83828e-19 $X=2.865 $Y=0.655 $X2=0
+ $Y2=0
cc_192 N_VPWR_c_270_n N_Y_M1001_d 0.00413932f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_193 N_VPWR_c_277_n Y 0.021327f $X=2.915 $Y=3.33 $X2=0 $Y2=0
cc_194 N_VPWR_c_270_n Y 0.0131749f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_195 N_VPWR_c_270_n A_504_367# 0.0041718f $X=3.12 $Y=3.33 $X2=-0.19 $Y2=-0.245
cc_196 N_Y_c_319_n N_VGND_c_360_n 0.0177571f $X=1.69 $Y=0.42 $X2=0 $Y2=0
cc_197 N_Y_M1004_s N_VGND_c_362_n 0.00371702f $X=1.565 $Y=0.235 $X2=0 $Y2=0
cc_198 N_Y_c_319_n N_VGND_c_362_n 0.0100204f $X=1.69 $Y=0.42 $X2=0 $Y2=0
cc_199 N_Y_c_316_n N_A_396_47#_M1004_d 7.89293e-19 $X=2.015 $Y=1.15 $X2=-0.19
+ $Y2=-0.245
cc_200 N_Y_c_316_n N_A_396_47#_c_400_n 0.00692608f $X=2.015 $Y=1.15 $X2=0 $Y2=0
cc_201 N_VGND_c_362_n N_A_396_47#_M1004_d 0.00224858f $X=3.12 $Y=0 $X2=-0.19
+ $Y2=-0.245
cc_202 N_VGND_c_362_n N_A_396_47#_M1008_d 0.00231264f $X=3.12 $Y=0 $X2=0 $Y2=0
cc_203 N_VGND_M1006_d N_A_396_47#_c_401_n 0.00574897f $X=2.41 $Y=0.235 $X2=0
+ $Y2=0
cc_204 N_VGND_c_359_n N_A_396_47#_c_401_n 0.0215546f $X=2.62 $Y=0.43 $X2=0 $Y2=0
cc_205 N_VGND_c_360_n N_A_396_47#_c_401_n 0.00206528f $X=2.455 $Y=0 $X2=0 $Y2=0
cc_206 N_VGND_c_361_n N_A_396_47#_c_401_n 0.00237862f $X=3.12 $Y=0 $X2=0 $Y2=0
cc_207 N_VGND_c_362_n N_A_396_47#_c_401_n 0.00964661f $X=3.12 $Y=0 $X2=0 $Y2=0
cc_208 N_VGND_c_361_n N_A_396_47#_c_399_n 0.0170745f $X=3.12 $Y=0 $X2=0 $Y2=0
cc_209 N_VGND_c_362_n N_A_396_47#_c_399_n 0.0103698f $X=3.12 $Y=0 $X2=0 $Y2=0
cc_210 N_VGND_c_360_n N_A_396_47#_c_400_n 0.0159203f $X=2.455 $Y=0 $X2=0 $Y2=0
cc_211 N_VGND_c_362_n N_A_396_47#_c_400_n 0.0122269f $X=3.12 $Y=0 $X2=0 $Y2=0
