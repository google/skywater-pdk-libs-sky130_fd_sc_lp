* File: sky130_fd_sc_lp__dfstp_lp.spice
* Created: Wed Sep  2 09:44:41 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__dfstp_lp.pex.spice"
.subckt sky130_fd_sc_lp__dfstp_lp  VNB VPB D CLK SET_B VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* SET_B	SET_B
* CLK	CLK
* D	D
* VPB	VPB
* VNB	VNB
MM1022 A_110_57# N_D_M1022_g N_VGND_M1022_s VNB NSHORT L=0.15 W=0.42 AD=0.0441
+ AS=0.1113 PD=0.63 PS=1.37 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1010 N_A_135_409#_M1010_d N_D_M1010_g A_110_57# VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.0441 PD=1.37 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1023 A_373_109# N_CLK_M1023_g N_A_266_409#_M1023_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1134 PD=0.63 PS=1.38 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.3 A=0.063 P=1.14 MULT=1
MM1013 N_VGND_M1013_d N_CLK_M1013_g A_373_109# VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1014 A_531_109# N_A_266_409#_M1014_g N_VGND_M1013_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75001
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1011 N_A_479_409#_M1011_d N_A_266_409#_M1011_g A_531_109# VNB NSHORT L=0.15
+ W=0.42 AD=0.1113 AS=0.0441 PD=1.37 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8
+ SA=75001.3 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1028 N_A_709_419#_M1028_d N_A_266_409#_M1028_g N_A_135_409#_M1028_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.08505 AS=0.1113 PD=0.825 PS=1.37 NRD=18.564 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.2 A=0.063 P=1.14 MULT=1
MM1017 A_904_125# N_A_479_409#_M1017_g N_A_709_419#_M1028_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.08505 PD=0.63 PS=0.825 NRD=14.28 NRS=17.136 M=1 R=2.8
+ SA=75000.7 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1008 N_VGND_M1008_d N_A_943_321#_M1008_g A_904_125# VNB NSHORT L=0.15 W=0.42
+ AD=0.2097 AS=0.0441 PD=2.01 PS=0.63 NRD=126.936 NRS=14.28 M=1 R=2.8 SA=75001.1
+ SB=75000.3 A=0.063 P=1.14 MULT=1
MM1019 A_1256_125# N_A_709_419#_M1019_g N_A_943_321#_M1019_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0504 AS=0.1197 PD=0.66 PS=1.41 NRD=18.564 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75003.4 A=0.063 P=1.14 MULT=1
MM1007 N_VGND_M1007_d N_SET_B_M1007_g A_1256_125# VNB NSHORT L=0.15 W=0.42
+ AD=0.0882 AS=0.0504 PD=0.84 PS=0.66 NRD=11.424 NRS=18.564 M=1 R=2.8 SA=75000.6
+ SB=75003 A=0.063 P=1.14 MULT=1
MM1002 A_1448_125# N_A_709_419#_M1002_g N_VGND_M1007_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.0882 PD=0.66 PS=0.84 NRD=18.564 NRS=28.56 M=1 R=2.8 SA=75001.2
+ SB=75002.4 A=0.063 P=1.14 MULT=1
MM1030 N_A_1526_125#_M1030_d N_A_479_409#_M1030_g A_1448_125# VNB NSHORT L=0.15
+ W=0.42 AD=0.13335 AS=0.0504 PD=1.055 PS=0.66 NRD=101.424 NRS=18.564 M=1 R=2.8
+ SA=75001.6 SB=75002 A=0.063 P=1.14 MULT=1
MM1032 A_1683_125# N_A_266_409#_M1032_g N_A_1526_125#_M1030_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0504 AS=0.13335 PD=0.66 PS=1.055 NRD=18.564 NRS=0 M=1 R=2.8
+ SA=75002.3 SB=75001.3 A=0.063 P=1.14 MULT=1
MM1020 A_1761_125# N_A_1731_99#_M1020_g A_1683_125# VNB NSHORT L=0.15 W=0.42
+ AD=0.10605 AS=0.0504 PD=0.925 PS=0.66 NRD=56.424 NRS=18.564 M=1 R=2.8
+ SA=75002.7 SB=75000.9 A=0.063 P=1.14 MULT=1
MM1036 N_VGND_M1036_d N_SET_B_M1036_g A_1761_125# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.10605 PD=1.41 PS=0.925 NRD=0 NRS=56.424 M=1 R=2.8 SA=75003.4
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1035 A_2104_47# N_A_1526_125#_M1035_g N_A_1731_99#_M1035_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.1197 PD=0.63 PS=1.41 NRD=14.28 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1037 N_VGND_M1037_d N_A_1526_125#_M1037_g A_2104_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1001 A_2374_74# N_A_1526_125#_M1001_g N_A_2287_74#_M1001_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.1197 PD=0.63 PS=1.41 NRD=14.28 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.4 A=0.063 P=1.14 MULT=1
MM1003 N_VGND_M1003_d N_A_1526_125#_M1003_g A_2374_74# VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1015 A_2532_74# N_A_2287_74#_M1015_g N_VGND_M1003_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75001
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1006 N_Q_M1006_d N_A_2287_74#_M1006_g A_2532_74# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.4
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1005 N_A_135_409#_M1005_d N_D_M1005_g N_VPWR_M1005_s VPB PHIGHVT L=0.25 W=1
+ AD=0.285 AS=0.285 PD=2.57 PS=2.57 NRD=0 NRS=0 M=1 R=4 SA=125000 SB=125000
+ A=0.25 P=2.5 MULT=1
MM1029 N_VPWR_M1029_d N_CLK_M1029_g N_A_266_409#_M1029_s VPB PHIGHVT L=0.25 W=1
+ AD=0.14 AS=0.285 PD=1.28 PS=2.57 NRD=0 NRS=0 M=1 R=4 SA=125000 SB=125001
+ A=0.25 P=2.5 MULT=1
MM1018 N_A_479_409#_M1018_d N_A_266_409#_M1018_g N_VPWR_M1029_d VPB PHIGHVT
+ L=0.25 W=1 AD=0.285 AS=0.14 PD=2.57 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125001
+ SB=125000 A=0.25 P=2.5 MULT=1
MM1021 N_A_709_419#_M1021_d N_A_479_409#_M1021_g N_A_135_409#_M1021_s VPB
+ PHIGHVT L=0.25 W=1 AD=0.305 AS=0.285 PD=1.61 PS=2.57 NRD=65.01 NRS=0 M=1 R=4
+ SA=125000 SB=125007 A=0.25 P=2.5 MULT=1
MM1026 A_881_419# N_A_266_409#_M1026_g N_A_709_419#_M1021_d VPB PHIGHVT L=0.25
+ W=1 AD=0.155 AS=0.305 PD=1.31 PS=1.61 NRD=19.6803 NRS=0 M=1 R=4 SA=125001
+ SB=125006 A=0.25 P=2.5 MULT=1
MM1027 N_VPWR_M1027_d N_A_943_321#_M1027_g A_881_419# VPB PHIGHVT L=0.25 W=1
+ AD=0.3175 AS=0.155 PD=1.635 PS=1.31 NRD=0 NRS=19.6803 M=1 R=4 SA=125002
+ SB=125005 A=0.25 P=2.5 MULT=1
MM1012 N_A_943_321#_M1012_d N_A_709_419#_M1012_g N_VPWR_M1027_d VPB PHIGHVT
+ L=0.25 W=1 AD=0.1475 AS=0.3175 PD=1.295 PS=1.635 NRD=0 NRS=69.9153 M=1 R=4
+ SA=125002 SB=125004 A=0.25 P=2.5 MULT=1
MM1025 N_VPWR_M1025_d N_SET_B_M1025_g N_A_943_321#_M1012_d VPB PHIGHVT L=0.25
+ W=1 AD=0.2975 AS=0.1475 PD=1.595 PS=1.295 NRD=62.0353 NRS=2.9353 M=1 R=4
+ SA=125003 SB=125004 A=0.25 P=2.5 MULT=1
MM1031 A_1448_419# N_A_709_419#_M1031_g N_VPWR_M1025_d VPB PHIGHVT L=0.25 W=1
+ AD=0.12 AS=0.2975 PD=1.24 PS=1.595 NRD=12.7853 NRS=0 M=1 R=4 SA=125004
+ SB=125003 A=0.25 P=2.5 MULT=1
MM1009 N_A_1526_125#_M1009_d N_A_266_409#_M1009_g A_1448_419# VPB PHIGHVT L=0.25
+ W=1 AD=0.325 AS=0.12 PD=1.65 PS=1.24 NRD=66.98 NRS=12.7853 M=1 R=4 SA=125004
+ SB=125002 A=0.25 P=2.5 MULT=1
MM1024 A_1726_419# N_A_479_409#_M1024_g N_A_1526_125#_M1009_d VPB PHIGHVT L=0.25
+ W=1 AD=0.145 AS=0.325 PD=1.29 PS=1.65 NRD=17.7103 NRS=5.8903 M=1 R=4 SA=125005
+ SB=125001 A=0.25 P=2.5 MULT=1
MM1000 N_VPWR_M1000_d N_A_1731_99#_M1000_g A_1726_419# VPB PHIGHVT L=0.25 W=1
+ AD=0.265 AS=0.145 PD=1.53 PS=1.29 NRD=0 NRS=17.7103 M=1 R=4 SA=125006
+ SB=125001 A=0.25 P=2.5 MULT=1
MM1033 N_A_1526_125#_M1033_d N_SET_B_M1033_g N_VPWR_M1000_d VPB PHIGHVT L=0.25
+ W=1 AD=0.285 AS=0.265 PD=2.57 PS=1.53 NRD=0 NRS=49.2303 M=1 R=4 SA=125007
+ SB=125000 A=0.25 P=2.5 MULT=1
MM1034 N_VPWR_M1034_d N_A_1526_125#_M1034_g N_A_1731_99#_M1034_s VPB PHIGHVT
+ L=0.25 W=1 AD=0.455 AS=0.285 PD=2.91 PS=2.57 NRD=33.4703 NRS=0 M=1 R=4
+ SA=125000 SB=125000 A=0.25 P=2.5 MULT=1
MM1016 N_VPWR_M1016_d N_A_1526_125#_M1016_g N_A_2287_74#_M1016_s VPB PHIGHVT
+ L=0.25 W=1 AD=0.14 AS=0.285 PD=1.28 PS=2.57 NRD=0 NRS=0 M=1 R=4 SA=125000
+ SB=125001 A=0.25 P=2.5 MULT=1
MM1004 N_Q_M1004_d N_A_2287_74#_M1004_g N_VPWR_M1016_d VPB PHIGHVT L=0.25 W=1
+ AD=0.285 AS=0.14 PD=2.57 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125001 SB=125000
+ A=0.25 P=2.5 MULT=1
DX38_noxref VNB VPB NWDIODE A=25.9633 P=31.65
c_269 VPB 0 1.2513e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_lp__dfstp_lp.pxi.spice"
*
.ends
*
*
