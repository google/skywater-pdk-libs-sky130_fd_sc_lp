* File: sky130_fd_sc_lp__a32oi_4.pxi.spice
* Created: Fri Aug 28 10:02:01 2020
* 
x_PM_SKY130_FD_SC_LP__A32OI_4%B2 N_B2_c_134_n N_B2_M1002_g N_B2_M1006_g
+ N_B2_c_136_n N_B2_M1013_g N_B2_M1020_g N_B2_c_138_n N_B2_M1016_g N_B2_M1021_g
+ N_B2_c_140_n N_B2_M1025_g N_B2_M1032_g B2 B2 B2 B2 N_B2_c_143_n
+ PM_SKY130_FD_SC_LP__A32OI_4%B2
x_PM_SKY130_FD_SC_LP__A32OI_4%B1 N_B1_c_217_n N_B1_M1010_g N_B1_M1001_g
+ N_B1_c_219_n N_B1_M1023_g N_B1_M1015_g N_B1_c_221_n N_B1_M1024_g N_B1_M1019_g
+ N_B1_c_223_n N_B1_M1038_g N_B1_M1033_g B1 B1 B1 B1 N_B1_c_226_n
+ PM_SKY130_FD_SC_LP__A32OI_4%B1
x_PM_SKY130_FD_SC_LP__A32OI_4%A1 N_A1_M1003_g N_A1_M1012_g N_A1_c_300_n
+ N_A1_M1005_g N_A1_M1034_g N_A1_c_301_n N_A1_M1014_g N_A1_c_302_n N_A1_M1027_g
+ N_A1_M1039_g N_A1_c_303_n N_A1_M1037_g A1 A1 A1 A1 N_A1_c_305_n
+ PM_SKY130_FD_SC_LP__A32OI_4%A1
x_PM_SKY130_FD_SC_LP__A32OI_4%A2 N_A2_c_381_n N_A2_M1004_g N_A2_c_372_n
+ N_A2_M1009_g N_A2_c_373_n N_A2_M1028_g N_A2_M1017_g N_A2_c_375_n N_A2_M1030_g
+ N_A2_M1022_g N_A2_c_377_n N_A2_M1035_g N_A2_M1029_g A2 A2 A2 A2 N_A2_c_380_n
+ PM_SKY130_FD_SC_LP__A32OI_4%A2
x_PM_SKY130_FD_SC_LP__A32OI_4%A3 N_A3_M1000_g N_A3_c_453_n N_A3_M1008_g
+ N_A3_M1007_g N_A3_c_454_n N_A3_M1011_g N_A3_M1018_g N_A3_c_455_n N_A3_M1031_g
+ N_A3_M1026_g N_A3_c_456_n N_A3_M1036_g A3 A3 A3 A3 A3 N_A3_c_458_n
+ N_A3_c_459_n PM_SKY130_FD_SC_LP__A32OI_4%A3
x_PM_SKY130_FD_SC_LP__A32OI_4%A_42_367# N_A_42_367#_M1006_d N_A_42_367#_M1020_d
+ N_A_42_367#_M1032_d N_A_42_367#_M1015_s N_A_42_367#_M1033_s
+ N_A_42_367#_M1012_s N_A_42_367#_M1039_s N_A_42_367#_M1017_d
+ N_A_42_367#_M1029_d N_A_42_367#_M1007_s N_A_42_367#_M1026_s
+ N_A_42_367#_c_534_n N_A_42_367#_c_535_n N_A_42_367#_c_546_n
+ N_A_42_367#_c_598_p N_A_42_367#_c_548_n N_A_42_367#_c_602_p
+ N_A_42_367#_c_550_n N_A_42_367#_c_605_p N_A_42_367#_c_552_n
+ N_A_42_367#_c_610_p N_A_42_367#_c_632_p N_A_42_367#_c_554_n
+ N_A_42_367#_c_620_p N_A_42_367#_c_557_n N_A_42_367#_c_636_p
+ N_A_42_367#_c_561_n N_A_42_367#_c_536_n N_A_42_367#_c_623_p
+ N_A_42_367#_c_529_n N_A_42_367#_c_530_n N_A_42_367#_c_538_n
+ N_A_42_367#_c_531_n N_A_42_367#_c_540_n N_A_42_367#_c_532_n
+ N_A_42_367#_c_542_n N_A_42_367#_c_633_p N_A_42_367#_c_634_p
+ N_A_42_367#_c_635_p N_A_42_367#_c_560_n N_A_42_367#_c_615_p
+ N_A_42_367#_c_575_n N_A_42_367#_c_533_n N_A_42_367#_c_590_n
+ PM_SKY130_FD_SC_LP__A32OI_4%A_42_367#
x_PM_SKY130_FD_SC_LP__A32OI_4%Y N_Y_M1010_d N_Y_M1024_d N_Y_M1005_d N_Y_M1027_d
+ N_Y_M1006_s N_Y_M1021_s N_Y_M1001_d N_Y_M1019_d N_Y_c_678_n N_Y_c_668_n
+ N_Y_c_669_n N_Y_c_689_n N_Y_c_670_n N_Y_c_694_n N_Y_c_671_n N_Y_c_710_n
+ N_Y_c_672_n N_Y_c_737_n N_Y_c_673_n N_Y_c_674_n N_Y_c_675_n N_Y_c_676_n Y Y Y
+ Y Y N_Y_c_677_n PM_SKY130_FD_SC_LP__A32OI_4%Y
x_PM_SKY130_FD_SC_LP__A32OI_4%VPWR N_VPWR_M1003_d N_VPWR_M1034_d N_VPWR_M1004_s
+ N_VPWR_M1022_s N_VPWR_M1000_d N_VPWR_M1018_d N_VPWR_c_805_n N_VPWR_c_806_n
+ N_VPWR_c_807_n N_VPWR_c_808_n N_VPWR_c_809_n N_VPWR_c_810_n N_VPWR_c_811_n
+ N_VPWR_c_812_n N_VPWR_c_813_n N_VPWR_c_814_n VPWR N_VPWR_c_815_n
+ N_VPWR_c_816_n N_VPWR_c_817_n N_VPWR_c_818_n N_VPWR_c_804_n N_VPWR_c_820_n
+ N_VPWR_c_821_n N_VPWR_c_822_n N_VPWR_c_823_n N_VPWR_c_824_n
+ PM_SKY130_FD_SC_LP__A32OI_4%VPWR
x_PM_SKY130_FD_SC_LP__A32OI_4%A_28_47# N_A_28_47#_M1002_s N_A_28_47#_M1013_s
+ N_A_28_47#_M1025_s N_A_28_47#_M1023_s N_A_28_47#_M1038_s N_A_28_47#_c_946_n
+ N_A_28_47#_c_949_n N_A_28_47#_c_947_n N_A_28_47#_c_980_p N_A_28_47#_c_955_n
+ N_A_28_47#_c_977_p N_A_28_47#_c_959_n N_A_28_47#_c_948_n N_A_28_47#_c_960_n
+ PM_SKY130_FD_SC_LP__A32OI_4%A_28_47#
x_PM_SKY130_FD_SC_LP__A32OI_4%VGND N_VGND_M1002_d N_VGND_M1016_d N_VGND_M1008_d
+ N_VGND_M1011_d N_VGND_M1036_d N_VGND_c_991_n N_VGND_c_992_n N_VGND_c_993_n
+ N_VGND_c_994_n N_VGND_c_995_n N_VGND_c_996_n N_VGND_c_997_n N_VGND_c_998_n
+ N_VGND_c_999_n N_VGND_c_1000_n VGND N_VGND_c_1001_n N_VGND_c_1002_n
+ N_VGND_c_1003_n N_VGND_c_1004_n N_VGND_c_1005_n N_VGND_c_1006_n
+ N_VGND_c_1007_n PM_SKY130_FD_SC_LP__A32OI_4%VGND
x_PM_SKY130_FD_SC_LP__A32OI_4%A_840_47# N_A_840_47#_M1005_s N_A_840_47#_M1014_s
+ N_A_840_47#_M1037_s N_A_840_47#_M1028_d N_A_840_47#_M1035_d
+ N_A_840_47#_c_1110_n PM_SKY130_FD_SC_LP__A32OI_4%A_840_47#
x_PM_SKY130_FD_SC_LP__A32OI_4%A_1267_47# N_A_1267_47#_M1009_s
+ N_A_1267_47#_M1030_s N_A_1267_47#_M1008_s N_A_1267_47#_M1031_s
+ N_A_1267_47#_c_1143_n N_A_1267_47#_c_1170_n N_A_1267_47#_c_1154_n
+ N_A_1267_47#_c_1175_n N_A_1267_47#_c_1158_n
+ PM_SKY130_FD_SC_LP__A32OI_4%A_1267_47#
cc_1 VNB N_B2_c_134_n 0.0218823f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=1.185
cc_2 VNB N_B2_M1006_g 0.0109769f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=2.465
cc_3 VNB N_B2_c_136_n 0.0160063f $X=-0.19 $Y=-0.245 $X2=0.91 $Y2=1.185
cc_4 VNB N_B2_M1020_g 0.00665511f $X=-0.19 $Y=-0.245 $X2=0.98 $Y2=2.465
cc_5 VNB N_B2_c_138_n 0.0160063f $X=-0.19 $Y=-0.245 $X2=1.34 $Y2=1.185
cc_6 VNB N_B2_M1021_g 0.00665511f $X=-0.19 $Y=-0.245 $X2=1.41 $Y2=2.465
cc_7 VNB N_B2_c_140_n 0.0162447f $X=-0.19 $Y=-0.245 $X2=1.77 $Y2=1.185
cc_8 VNB N_B2_M1032_g 0.0068117f $X=-0.19 $Y=-0.245 $X2=1.84 $Y2=2.465
cc_9 VNB B2 0.0101842f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.21
cc_10 VNB N_B2_c_143_n 0.110923f $X=-0.19 $Y=-0.245 $X2=1.77 $Y2=1.35
cc_11 VNB N_B1_c_217_n 0.0164438f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=1.185
cc_12 VNB N_B1_M1001_g 0.0068117f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=2.465
cc_13 VNB N_B1_c_219_n 0.0162054f $X=-0.19 $Y=-0.245 $X2=0.91 $Y2=1.185
cc_14 VNB N_B1_M1015_g 0.00665511f $X=-0.19 $Y=-0.245 $X2=0.98 $Y2=2.465
cc_15 VNB N_B1_c_221_n 0.0162054f $X=-0.19 $Y=-0.245 $X2=1.34 $Y2=1.185
cc_16 VNB N_B1_M1019_g 0.00665511f $X=-0.19 $Y=-0.245 $X2=1.41 $Y2=2.465
cc_17 VNB N_B1_c_223_n 0.0220814f $X=-0.19 $Y=-0.245 $X2=1.77 $Y2=1.185
cc_18 VNB N_B1_M1033_g 0.00735693f $X=-0.19 $Y=-0.245 $X2=1.84 $Y2=2.465
cc_19 VNB B1 0.00418971f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.21
cc_20 VNB N_B1_c_226_n 0.0949524f $X=-0.19 $Y=-0.245 $X2=1.84 $Y2=1.35
cc_21 VNB N_A1_c_300_n 0.0220814f $X=-0.19 $Y=-0.245 $X2=0.91 $Y2=0.655
cc_22 VNB N_A1_c_301_n 0.0162054f $X=-0.19 $Y=-0.245 $X2=1.34 $Y2=0.655
cc_23 VNB N_A1_c_302_n 0.0161977f $X=-0.19 $Y=-0.245 $X2=1.41 $Y2=2.465
cc_24 VNB N_A1_c_303_n 0.0157951f $X=-0.19 $Y=-0.245 $X2=1.84 $Y2=2.465
cc_25 VNB A1 0.00195099f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.21
cc_26 VNB N_A1_c_305_n 0.127904f $X=-0.19 $Y=-0.245 $X2=1.77 $Y2=1.35
cc_27 VNB N_A2_c_372_n 0.016408f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=1.515
cc_28 VNB N_A2_c_373_n 0.0162018f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A2_M1017_g 0.00812411f $X=-0.19 $Y=-0.245 $X2=0.98 $Y2=2.465
cc_30 VNB N_A2_c_375_n 0.0162054f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A2_M1022_g 0.00665929f $X=-0.19 $Y=-0.245 $X2=1.41 $Y2=2.465
cc_32 VNB N_A2_c_377_n 0.0220814f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A2_M1029_g 0.00681588f $X=-0.19 $Y=-0.245 $X2=1.84 $Y2=2.465
cc_34 VNB A2 0.00285297f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.21
cc_35 VNB N_A2_c_380_n 0.125239f $X=-0.19 $Y=-0.245 $X2=1.68 $Y2=1.35
cc_36 VNB N_A3_c_453_n 0.0212151f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=2.465
cc_37 VNB N_A3_c_454_n 0.0160063f $X=-0.19 $Y=-0.245 $X2=0.98 $Y2=2.465
cc_38 VNB N_A3_c_455_n 0.0160063f $X=-0.19 $Y=-0.245 $X2=1.41 $Y2=2.465
cc_39 VNB N_A3_c_456_n 0.0212151f $X=-0.19 $Y=-0.245 $X2=1.84 $Y2=2.465
cc_40 VNB A3 0.0126061f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A3_c_458_n 0.109735f $X=-0.19 $Y=-0.245 $X2=0.32 $Y2=1.35
cc_42 VNB N_A3_c_459_n 0.0835631f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=1.35
cc_43 VNB N_A_42_367#_c_529_n 0.00289786f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_42_367#_c_530_n 0.00186335f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_42_367#_c_531_n 6.77852e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_42_367#_c_532_n 0.00403301f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_42_367#_c_533_n 0.00244474f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_Y_c_668_n 0.00225492f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.21
cc_49 VNB N_Y_c_669_n 0.00228659f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.21
cc_50 VNB N_Y_c_670_n 0.00336316f $X=-0.19 $Y=-0.245 $X2=0.32 $Y2=1.35
cc_51 VNB N_Y_c_671_n 0.00225492f $X=-0.19 $Y=-0.245 $X2=1.68 $Y2=1.35
cc_52 VNB N_Y_c_672_n 0.00452108f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_Y_c_673_n 0.00608928f $X=-0.19 $Y=-0.245 $X2=1.68 $Y2=1.322
cc_54 VNB N_Y_c_674_n 0.00228659f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_Y_c_675_n 0.00228659f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_Y_c_676_n 0.00228659f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_Y_c_677_n 0.0128441f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_VPWR_c_804_n 0.442315f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_28_47#_c_946_n 0.0233935f $X=-0.19 $Y=-0.245 $X2=1.41 $Y2=1.515
cc_60 VNB N_A_28_47#_c_947_n 0.00879096f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_A_28_47#_c_948_n 0.00434881f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_991_n 3.99129e-19 $X=-0.19 $Y=-0.245 $X2=1.41 $Y2=1.515
cc_63 VNB N_VGND_c_992_n 3.99129e-19 $X=-0.19 $Y=-0.245 $X2=1.77 $Y2=1.185
cc_64 VNB N_VGND_c_993_n 0.0065129f $X=-0.19 $Y=-0.245 $X2=1.84 $Y2=2.465
cc_65 VNB N_VGND_c_994_n 3.0911e-19 $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_66 VNB N_VGND_c_995_n 0.0129398f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.21
cc_67 VNB N_VGND_c_996_n 0.0338983f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_VGND_c_997_n 0.148711f $X=-0.19 $Y=-0.245 $X2=0.32 $Y2=1.35
cc_69 VNB N_VGND_c_998_n 0.00510842f $X=-0.19 $Y=-0.245 $X2=0.48 $Y2=1.35
cc_70 VNB N_VGND_c_999_n 0.0129398f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=1.35
cc_71 VNB N_VGND_c_1000_n 0.00436868f $X=-0.19 $Y=-0.245 $X2=0.91 $Y2=1.35
cc_72 VNB N_VGND_c_1001_n 0.015535f $X=-0.19 $Y=-0.245 $X2=1.41 $Y2=1.35
cc_73 VNB N_VGND_c_1002_n 0.0129398f $X=-0.19 $Y=-0.245 $X2=1.84 $Y2=1.35
cc_74 VNB N_VGND_c_1003_n 0.0145539f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_VGND_c_1004_n 0.507607f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_VGND_c_1005_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_VGND_c_1006_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_VGND_c_1007_n 0.00513431f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_A_840_47#_c_1110_n 0.00766655f $X=-0.19 $Y=-0.245 $X2=1.84 $Y2=2.465
cc_80 VNB N_A_1267_47#_c_1143_n 0.00986158f $X=-0.19 $Y=-0.245 $X2=0.98
+ $Y2=2.465
cc_81 VPB N_B2_M1006_g 0.0267679f $X=-0.19 $Y=1.655 $X2=0.55 $Y2=2.465
cc_82 VPB N_B2_M1020_g 0.0182686f $X=-0.19 $Y=1.655 $X2=0.98 $Y2=2.465
cc_83 VPB N_B2_M1021_g 0.0182686f $X=-0.19 $Y=1.655 $X2=1.41 $Y2=2.465
cc_84 VPB N_B2_M1032_g 0.0183346f $X=-0.19 $Y=1.655 $X2=1.84 $Y2=2.465
cc_85 VPB N_B1_M1001_g 0.0183346f $X=-0.19 $Y=1.655 $X2=0.55 $Y2=2.465
cc_86 VPB N_B1_M1015_g 0.0182686f $X=-0.19 $Y=1.655 $X2=0.98 $Y2=2.465
cc_87 VPB N_B1_M1019_g 0.0182686f $X=-0.19 $Y=1.655 $X2=1.41 $Y2=2.465
cc_88 VPB N_B1_M1033_g 0.0195511f $X=-0.19 $Y=1.655 $X2=1.84 $Y2=2.465
cc_89 VPB N_A1_M1003_g 0.0188406f $X=-0.19 $Y=1.655 $X2=0.48 $Y2=0.655
cc_90 VPB N_A1_M1012_g 0.017602f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_91 VPB N_A1_M1034_g 0.020365f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_92 VPB N_A1_M1039_g 0.0204302f $X=-0.19 $Y=1.655 $X2=1.77 $Y2=0.655
cc_93 VPB N_A1_c_305_n 0.0204667f $X=-0.19 $Y=1.655 $X2=1.77 $Y2=1.35
cc_94 VPB N_A2_c_381_n 0.0181291f $X=-0.19 $Y=1.655 $X2=0.48 $Y2=1.185
cc_95 VPB N_A2_M1017_g 0.0220157f $X=-0.19 $Y=1.655 $X2=0.98 $Y2=2.465
cc_96 VPB N_A2_M1022_g 0.0185652f $X=-0.19 $Y=1.655 $X2=1.41 $Y2=2.465
cc_97 VPB N_A2_M1029_g 0.018727f $X=-0.19 $Y=1.655 $X2=1.84 $Y2=2.465
cc_98 VPB N_A2_c_380_n 0.00754403f $X=-0.19 $Y=1.655 $X2=1.68 $Y2=1.35
cc_99 VPB N_A3_M1000_g 0.0182588f $X=-0.19 $Y=1.655 $X2=0.48 $Y2=0.655
cc_100 VPB N_A3_M1007_g 0.0180978f $X=-0.19 $Y=1.655 $X2=0.91 $Y2=0.655
cc_101 VPB N_A3_M1018_g 0.0180978f $X=-0.19 $Y=1.655 $X2=1.34 $Y2=0.655
cc_102 VPB N_A3_M1026_g 0.0226484f $X=-0.19 $Y=1.655 $X2=1.77 $Y2=0.655
cc_103 VPB N_A3_c_458_n 0.0105104f $X=-0.19 $Y=1.655 $X2=0.32 $Y2=1.35
cc_104 VPB N_A_42_367#_c_534_n 0.00746637f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_105 VPB N_A_42_367#_c_535_n 0.0430376f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_106 VPB N_A_42_367#_c_536_n 4.98048e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_107 VPB N_A_42_367#_c_529_n 0.00559032f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_108 VPB N_A_42_367#_c_538_n 9.96097e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_109 VPB N_A_42_367#_c_531_n 0.00559032f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_110 VPB N_A_42_367#_c_540_n 9.96097e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_111 VPB N_A_42_367#_c_532_n 0.0110324f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_112 VPB N_A_42_367#_c_542_n 0.0498589f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_113 VPB N_VPWR_c_805_n 3.99129e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_114 VPB N_VPWR_c_806_n 0.0129398f $X=-0.19 $Y=1.655 $X2=1.77 $Y2=0.655
cc_115 VPB N_VPWR_c_807_n 0.00174197f $X=-0.19 $Y=1.655 $X2=1.84 $Y2=2.465
cc_116 VPB N_VPWR_c_808_n 0.00185219f $X=-0.19 $Y=1.655 $X2=1.115 $Y2=1.21
cc_117 VPB N_VPWR_c_809_n 0.0129398f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_118 VPB N_VPWR_c_810_n 3.0911e-19 $X=-0.19 $Y=1.655 $X2=0.32 $Y2=1.35
cc_119 VPB N_VPWR_c_811_n 3.0911e-19 $X=-0.19 $Y=1.655 $X2=0.98 $Y2=1.35
cc_120 VPB N_VPWR_c_812_n 3.99129e-19 $X=-0.19 $Y=1.655 $X2=1.77 $Y2=1.35
cc_121 VPB N_VPWR_c_813_n 0.0963228f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_122 VPB N_VPWR_c_814_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=1.322
cc_123 VPB N_VPWR_c_815_n 0.0129398f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_124 VPB N_VPWR_c_816_n 0.0129398f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_125 VPB N_VPWR_c_817_n 0.0129398f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_126 VPB N_VPWR_c_818_n 0.0330243f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_127 VPB N_VPWR_c_804_n 0.0719349f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_128 VPB N_VPWR_c_820_n 0.0104351f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_129 VPB N_VPWR_c_821_n 0.0108198f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_130 VPB N_VPWR_c_822_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_131 VPB N_VPWR_c_823_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_132 VPB N_VPWR_c_824_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_133 N_B2_c_140_n N_B1_c_217_n 0.0116609f $X=1.77 $Y=1.185 $X2=-0.19
+ $Y2=-0.245
cc_134 N_B2_M1032_g N_B1_M1001_g 0.0288895f $X=1.84 $Y=2.465 $X2=0 $Y2=0
cc_135 B2 B1 0.0158272f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_136 N_B2_c_143_n B1 0.00120583f $X=1.77 $Y=1.35 $X2=0 $Y2=0
cc_137 B2 N_B1_c_226_n 2.48316e-19 $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_138 N_B2_c_143_n N_B1_c_226_n 0.0230167f $X=1.77 $Y=1.35 $X2=0 $Y2=0
cc_139 N_B2_M1006_g N_A_42_367#_c_535_n 0.0029331f $X=0.55 $Y=2.465 $X2=0 $Y2=0
cc_140 B2 N_A_42_367#_c_535_n 0.0114434f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_141 N_B2_c_143_n N_A_42_367#_c_535_n 0.00585523f $X=1.77 $Y=1.35 $X2=0 $Y2=0
cc_142 N_B2_M1006_g N_A_42_367#_c_546_n 0.0115031f $X=0.55 $Y=2.465 $X2=0 $Y2=0
cc_143 N_B2_M1020_g N_A_42_367#_c_546_n 0.0115031f $X=0.98 $Y=2.465 $X2=0 $Y2=0
cc_144 N_B2_M1021_g N_A_42_367#_c_548_n 0.0115031f $X=1.41 $Y=2.465 $X2=0 $Y2=0
cc_145 N_B2_M1032_g N_A_42_367#_c_548_n 0.0115031f $X=1.84 $Y=2.465 $X2=0 $Y2=0
cc_146 N_B2_M1006_g N_Y_c_678_n 0.00947894f $X=0.55 $Y=2.465 $X2=0 $Y2=0
cc_147 N_B2_M1020_g N_Y_c_678_n 0.0102493f $X=0.98 $Y=2.465 $X2=0 $Y2=0
cc_148 N_B2_M1021_g N_Y_c_678_n 6.30056e-19 $X=1.41 $Y=2.465 $X2=0 $Y2=0
cc_149 N_B2_M1020_g N_Y_c_668_n 0.0138481f $X=0.98 $Y=2.465 $X2=0 $Y2=0
cc_150 N_B2_M1021_g N_Y_c_668_n 0.0138481f $X=1.41 $Y=2.465 $X2=0 $Y2=0
cc_151 B2 N_Y_c_668_n 0.0390831f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_152 N_B2_c_143_n N_Y_c_668_n 0.00279461f $X=1.77 $Y=1.35 $X2=0 $Y2=0
cc_153 N_B2_M1006_g N_Y_c_669_n 0.0140106f $X=0.55 $Y=2.465 $X2=0 $Y2=0
cc_154 N_B2_M1020_g N_Y_c_669_n 0.00372942f $X=0.98 $Y=2.465 $X2=0 $Y2=0
cc_155 B2 N_Y_c_669_n 0.0268977f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_156 N_B2_c_143_n N_Y_c_669_n 0.00286879f $X=1.77 $Y=1.35 $X2=0 $Y2=0
cc_157 N_B2_M1020_g N_Y_c_689_n 6.30056e-19 $X=0.98 $Y=2.465 $X2=0 $Y2=0
cc_158 N_B2_M1021_g N_Y_c_689_n 0.0102493f $X=1.41 $Y=2.465 $X2=0 $Y2=0
cc_159 N_B2_M1032_g N_Y_c_689_n 0.0102493f $X=1.84 $Y=2.465 $X2=0 $Y2=0
cc_160 N_B2_M1032_g N_Y_c_670_n 0.0142293f $X=1.84 $Y=2.465 $X2=0 $Y2=0
cc_161 B2 N_Y_c_670_n 0.00391091f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_162 N_B2_M1032_g N_Y_c_694_n 6.30056e-19 $X=1.84 $Y=2.465 $X2=0 $Y2=0
cc_163 N_B2_M1021_g N_Y_c_674_n 0.00372942f $X=1.41 $Y=2.465 $X2=0 $Y2=0
cc_164 N_B2_M1032_g N_Y_c_674_n 0.00372942f $X=1.84 $Y=2.465 $X2=0 $Y2=0
cc_165 B2 N_Y_c_674_n 0.0268977f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_166 N_B2_c_143_n N_Y_c_674_n 0.00286879f $X=1.77 $Y=1.35 $X2=0 $Y2=0
cc_167 N_B2_M1006_g N_VPWR_c_813_n 0.00357877f $X=0.55 $Y=2.465 $X2=0 $Y2=0
cc_168 N_B2_M1020_g N_VPWR_c_813_n 0.00357877f $X=0.98 $Y=2.465 $X2=0 $Y2=0
cc_169 N_B2_M1021_g N_VPWR_c_813_n 0.00357877f $X=1.41 $Y=2.465 $X2=0 $Y2=0
cc_170 N_B2_M1032_g N_VPWR_c_813_n 0.00357877f $X=1.84 $Y=2.465 $X2=0 $Y2=0
cc_171 N_B2_M1006_g N_VPWR_c_804_n 0.00634741f $X=0.55 $Y=2.465 $X2=0 $Y2=0
cc_172 N_B2_M1020_g N_VPWR_c_804_n 0.0053512f $X=0.98 $Y=2.465 $X2=0 $Y2=0
cc_173 N_B2_M1021_g N_VPWR_c_804_n 0.0053512f $X=1.41 $Y=2.465 $X2=0 $Y2=0
cc_174 N_B2_M1032_g N_VPWR_c_804_n 0.00537654f $X=1.84 $Y=2.465 $X2=0 $Y2=0
cc_175 N_B2_c_134_n N_A_28_47#_c_949_n 0.0122595f $X=0.48 $Y=1.185 $X2=0 $Y2=0
cc_176 N_B2_c_136_n N_A_28_47#_c_949_n 0.0122595f $X=0.91 $Y=1.185 $X2=0 $Y2=0
cc_177 B2 N_A_28_47#_c_949_n 0.039834f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_178 N_B2_c_143_n N_A_28_47#_c_949_n 0.0025922f $X=1.77 $Y=1.35 $X2=0 $Y2=0
cc_179 B2 N_A_28_47#_c_947_n 0.0159497f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_180 N_B2_c_143_n N_A_28_47#_c_947_n 0.00488323f $X=1.77 $Y=1.35 $X2=0 $Y2=0
cc_181 N_B2_c_138_n N_A_28_47#_c_955_n 0.0122129f $X=1.34 $Y=1.185 $X2=0 $Y2=0
cc_182 N_B2_c_140_n N_A_28_47#_c_955_n 0.0122595f $X=1.77 $Y=1.185 $X2=0 $Y2=0
cc_183 B2 N_A_28_47#_c_955_n 0.0382418f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_184 N_B2_c_143_n N_A_28_47#_c_955_n 0.0025922f $X=1.77 $Y=1.35 $X2=0 $Y2=0
cc_185 N_B2_c_143_n N_A_28_47#_c_959_n 5.98225e-19 $X=1.77 $Y=1.35 $X2=0 $Y2=0
cc_186 B2 N_A_28_47#_c_960_n 0.0142048f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_187 N_B2_c_143_n N_A_28_47#_c_960_n 0.00268449f $X=1.77 $Y=1.35 $X2=0 $Y2=0
cc_188 N_B2_c_134_n N_VGND_c_991_n 0.0120769f $X=0.48 $Y=1.185 $X2=0 $Y2=0
cc_189 N_B2_c_136_n N_VGND_c_991_n 0.0103898f $X=0.91 $Y=1.185 $X2=0 $Y2=0
cc_190 N_B2_c_138_n N_VGND_c_991_n 5.75816e-19 $X=1.34 $Y=1.185 $X2=0 $Y2=0
cc_191 N_B2_c_136_n N_VGND_c_992_n 5.75816e-19 $X=0.91 $Y=1.185 $X2=0 $Y2=0
cc_192 N_B2_c_138_n N_VGND_c_992_n 0.0103898f $X=1.34 $Y=1.185 $X2=0 $Y2=0
cc_193 N_B2_c_140_n N_VGND_c_992_n 0.0115588f $X=1.77 $Y=1.185 $X2=0 $Y2=0
cc_194 N_B2_c_140_n N_VGND_c_997_n 0.00486043f $X=1.77 $Y=1.185 $X2=0 $Y2=0
cc_195 N_B2_c_134_n N_VGND_c_1001_n 0.00486043f $X=0.48 $Y=1.185 $X2=0 $Y2=0
cc_196 N_B2_c_136_n N_VGND_c_1002_n 0.00486043f $X=0.91 $Y=1.185 $X2=0 $Y2=0
cc_197 N_B2_c_138_n N_VGND_c_1002_n 0.00486043f $X=1.34 $Y=1.185 $X2=0 $Y2=0
cc_198 N_B2_c_134_n N_VGND_c_1004_n 0.00918457f $X=0.48 $Y=1.185 $X2=0 $Y2=0
cc_199 N_B2_c_136_n N_VGND_c_1004_n 0.00824727f $X=0.91 $Y=1.185 $X2=0 $Y2=0
cc_200 N_B2_c_138_n N_VGND_c_1004_n 0.00824727f $X=1.34 $Y=1.185 $X2=0 $Y2=0
cc_201 N_B2_c_140_n N_VGND_c_1004_n 0.0082726f $X=1.77 $Y=1.185 $X2=0 $Y2=0
cc_202 B1 A1 0.0190359f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_203 N_B1_c_226_n A1 8.5474e-19 $X=3.65 $Y=1.35 $X2=0 $Y2=0
cc_204 N_B1_M1033_g N_A1_c_305_n 0.0206357f $X=3.56 $Y=2.465 $X2=0 $Y2=0
cc_205 B1 N_A1_c_305_n 2.5821e-19 $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_206 N_B1_c_226_n N_A1_c_305_n 0.0235325f $X=3.65 $Y=1.35 $X2=0 $Y2=0
cc_207 N_B1_M1001_g N_A_42_367#_c_550_n 0.0115031f $X=2.27 $Y=2.465 $X2=0 $Y2=0
cc_208 N_B1_M1015_g N_A_42_367#_c_550_n 0.0115031f $X=2.7 $Y=2.465 $X2=0 $Y2=0
cc_209 N_B1_M1019_g N_A_42_367#_c_552_n 0.0115031f $X=3.13 $Y=2.465 $X2=0 $Y2=0
cc_210 N_B1_M1033_g N_A_42_367#_c_552_n 0.0115031f $X=3.56 $Y=2.465 $X2=0 $Y2=0
cc_211 N_B1_M1001_g N_Y_c_689_n 6.30056e-19 $X=2.27 $Y=2.465 $X2=0 $Y2=0
cc_212 N_B1_M1001_g N_Y_c_670_n 0.0137739f $X=2.27 $Y=2.465 $X2=0 $Y2=0
cc_213 B1 N_Y_c_670_n 0.0182209f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_214 N_B1_c_226_n N_Y_c_670_n 0.00204649f $X=3.65 $Y=1.35 $X2=0 $Y2=0
cc_215 N_B1_M1001_g N_Y_c_694_n 0.0102493f $X=2.27 $Y=2.465 $X2=0 $Y2=0
cc_216 N_B1_M1015_g N_Y_c_694_n 0.0102493f $X=2.7 $Y=2.465 $X2=0 $Y2=0
cc_217 N_B1_M1019_g N_Y_c_694_n 6.30056e-19 $X=3.13 $Y=2.465 $X2=0 $Y2=0
cc_218 N_B1_M1015_g N_Y_c_671_n 0.0138481f $X=2.7 $Y=2.465 $X2=0 $Y2=0
cc_219 N_B1_M1019_g N_Y_c_671_n 0.0138481f $X=3.13 $Y=2.465 $X2=0 $Y2=0
cc_220 B1 N_Y_c_671_n 0.0390831f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_221 N_B1_c_226_n N_Y_c_671_n 0.00279461f $X=3.65 $Y=1.35 $X2=0 $Y2=0
cc_222 N_B1_M1015_g N_Y_c_710_n 6.30056e-19 $X=2.7 $Y=2.465 $X2=0 $Y2=0
cc_223 N_B1_M1019_g N_Y_c_710_n 0.0102493f $X=3.13 $Y=2.465 $X2=0 $Y2=0
cc_224 N_B1_M1033_g N_Y_c_710_n 0.0107612f $X=3.56 $Y=2.465 $X2=0 $Y2=0
cc_225 N_B1_M1033_g N_Y_c_672_n 0.0146778f $X=3.56 $Y=2.465 $X2=0 $Y2=0
cc_226 B1 N_Y_c_672_n 0.0225691f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_227 N_B1_c_226_n N_Y_c_672_n 0.00448874f $X=3.65 $Y=1.35 $X2=0 $Y2=0
cc_228 N_B1_M1001_g N_Y_c_675_n 0.00372942f $X=2.27 $Y=2.465 $X2=0 $Y2=0
cc_229 N_B1_M1015_g N_Y_c_675_n 0.00372942f $X=2.7 $Y=2.465 $X2=0 $Y2=0
cc_230 B1 N_Y_c_675_n 0.0268977f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_231 N_B1_c_226_n N_Y_c_675_n 0.00286879f $X=3.65 $Y=1.35 $X2=0 $Y2=0
cc_232 N_B1_M1019_g N_Y_c_676_n 0.00372942f $X=3.13 $Y=2.465 $X2=0 $Y2=0
cc_233 N_B1_M1033_g N_Y_c_676_n 0.00372942f $X=3.56 $Y=2.465 $X2=0 $Y2=0
cc_234 B1 N_Y_c_676_n 0.0268977f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_235 N_B1_c_226_n N_Y_c_676_n 0.00286879f $X=3.65 $Y=1.35 $X2=0 $Y2=0
cc_236 N_B1_c_217_n N_Y_c_677_n 0.00342863f $X=2.2 $Y=1.185 $X2=0 $Y2=0
cc_237 N_B1_c_219_n N_Y_c_677_n 0.0112464f $X=2.63 $Y=1.185 $X2=0 $Y2=0
cc_238 N_B1_c_221_n N_Y_c_677_n 0.0112464f $X=3.06 $Y=1.185 $X2=0 $Y2=0
cc_239 N_B1_c_223_n N_Y_c_677_n 0.0145623f $X=3.49 $Y=1.185 $X2=0 $Y2=0
cc_240 B1 N_Y_c_677_n 0.0995276f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_241 N_B1_c_226_n N_Y_c_677_n 0.0138338f $X=3.65 $Y=1.35 $X2=0 $Y2=0
cc_242 N_B1_M1033_g N_VPWR_c_805_n 9.37752e-19 $X=3.56 $Y=2.465 $X2=0 $Y2=0
cc_243 N_B1_M1001_g N_VPWR_c_813_n 0.00357877f $X=2.27 $Y=2.465 $X2=0 $Y2=0
cc_244 N_B1_M1015_g N_VPWR_c_813_n 0.00357877f $X=2.7 $Y=2.465 $X2=0 $Y2=0
cc_245 N_B1_M1019_g N_VPWR_c_813_n 0.00357877f $X=3.13 $Y=2.465 $X2=0 $Y2=0
cc_246 N_B1_M1033_g N_VPWR_c_813_n 0.00357877f $X=3.56 $Y=2.465 $X2=0 $Y2=0
cc_247 N_B1_M1001_g N_VPWR_c_804_n 0.00537654f $X=2.27 $Y=2.465 $X2=0 $Y2=0
cc_248 N_B1_M1015_g N_VPWR_c_804_n 0.0053512f $X=2.7 $Y=2.465 $X2=0 $Y2=0
cc_249 N_B1_M1019_g N_VPWR_c_804_n 0.0053512f $X=3.13 $Y=2.465 $X2=0 $Y2=0
cc_250 N_B1_M1033_g N_VPWR_c_804_n 0.0056187f $X=3.56 $Y=2.465 $X2=0 $Y2=0
cc_251 N_B1_c_217_n N_A_28_47#_c_948_n 0.0139555f $X=2.2 $Y=1.185 $X2=0 $Y2=0
cc_252 N_B1_c_219_n N_A_28_47#_c_948_n 0.0120709f $X=2.63 $Y=1.185 $X2=0 $Y2=0
cc_253 N_B1_c_221_n N_A_28_47#_c_948_n 0.0121645f $X=3.06 $Y=1.185 $X2=0 $Y2=0
cc_254 N_B1_c_223_n N_A_28_47#_c_948_n 0.0121645f $X=3.49 $Y=1.185 $X2=0 $Y2=0
cc_255 B1 N_A_28_47#_c_948_n 0.0038559f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_256 N_B1_c_217_n N_VGND_c_992_n 0.00109252f $X=2.2 $Y=1.185 $X2=0 $Y2=0
cc_257 N_B1_c_217_n N_VGND_c_997_n 0.00357877f $X=2.2 $Y=1.185 $X2=0 $Y2=0
cc_258 N_B1_c_219_n N_VGND_c_997_n 0.00357877f $X=2.63 $Y=1.185 $X2=0 $Y2=0
cc_259 N_B1_c_221_n N_VGND_c_997_n 0.00357877f $X=3.06 $Y=1.185 $X2=0 $Y2=0
cc_260 N_B1_c_223_n N_VGND_c_997_n 0.00357877f $X=3.49 $Y=1.185 $X2=0 $Y2=0
cc_261 N_B1_c_217_n N_VGND_c_1004_n 0.00537654f $X=2.2 $Y=1.185 $X2=0 $Y2=0
cc_262 N_B1_c_219_n N_VGND_c_1004_n 0.0053512f $X=2.63 $Y=1.185 $X2=0 $Y2=0
cc_263 N_B1_c_221_n N_VGND_c_1004_n 0.0053512f $X=3.06 $Y=1.185 $X2=0 $Y2=0
cc_264 N_B1_c_223_n N_VGND_c_1004_n 0.00665089f $X=3.49 $Y=1.185 $X2=0 $Y2=0
cc_265 N_A1_M1039_g N_A2_c_381_n 0.0135818f $X=5.73 $Y=2.465 $X2=-0.19
+ $Y2=-0.245
cc_266 N_A1_c_303_n N_A2_c_372_n 0.0186199f $X=5.83 $Y=1.185 $X2=0 $Y2=0
cc_267 N_A1_c_305_n N_A2_c_380_n 0.0388247f $X=5.73 $Y=1.425 $X2=0 $Y2=0
cc_268 N_A1_M1003_g N_A_42_367#_c_554_n 0.0125619f $X=4.1 $Y=2.465 $X2=0 $Y2=0
cc_269 N_A1_M1012_g N_A_42_367#_c_554_n 0.0125619f $X=4.53 $Y=2.465 $X2=0 $Y2=0
cc_270 N_A1_c_305_n N_A_42_367#_c_554_n 4.31989e-19 $X=5.73 $Y=1.425 $X2=0 $Y2=0
cc_271 N_A1_M1034_g N_A_42_367#_c_557_n 0.0140656f $X=4.96 $Y=2.465 $X2=0 $Y2=0
cc_272 N_A1_M1039_g N_A_42_367#_c_557_n 0.0140656f $X=5.73 $Y=2.465 $X2=0 $Y2=0
cc_273 N_A1_c_305_n N_A_42_367#_c_557_n 0.00189104f $X=5.73 $Y=1.425 $X2=0 $Y2=0
cc_274 N_A1_c_305_n N_A_42_367#_c_560_n 4.8757e-19 $X=5.73 $Y=1.425 $X2=0 $Y2=0
cc_275 N_A1_M1003_g N_Y_c_710_n 7.13394e-19 $X=4.1 $Y=2.465 $X2=0 $Y2=0
cc_276 N_A1_M1003_g N_Y_c_672_n 0.0106456f $X=4.1 $Y=2.465 $X2=0 $Y2=0
cc_277 N_A1_M1012_g N_Y_c_672_n 0.0100017f $X=4.53 $Y=2.465 $X2=0 $Y2=0
cc_278 N_A1_M1034_g N_Y_c_672_n 0.0117027f $X=4.96 $Y=2.465 $X2=0 $Y2=0
cc_279 N_A1_M1039_g N_Y_c_672_n 0.011645f $X=5.73 $Y=2.465 $X2=0 $Y2=0
cc_280 A1 N_Y_c_672_n 0.12368f $X=5.435 $Y=1.21 $X2=0 $Y2=0
cc_281 N_A1_c_305_n N_Y_c_672_n 0.0514992f $X=5.73 $Y=1.425 $X2=0 $Y2=0
cc_282 N_A1_c_303_n N_Y_c_737_n 0.00308541f $X=5.83 $Y=1.185 $X2=0 $Y2=0
cc_283 N_A1_c_302_n N_Y_c_673_n 6.22434e-19 $X=5.4 $Y=1.185 $X2=0 $Y2=0
cc_284 N_A1_c_303_n N_Y_c_673_n 0.0036441f $X=5.83 $Y=1.185 $X2=0 $Y2=0
cc_285 A1 N_Y_c_673_n 0.0176181f $X=5.435 $Y=1.21 $X2=0 $Y2=0
cc_286 N_A1_c_305_n N_Y_c_673_n 0.0104827f $X=5.73 $Y=1.425 $X2=0 $Y2=0
cc_287 N_A1_c_300_n N_Y_c_677_n 0.0145623f $X=4.54 $Y=1.185 $X2=0 $Y2=0
cc_288 N_A1_c_301_n N_Y_c_677_n 0.0112464f $X=4.97 $Y=1.185 $X2=0 $Y2=0
cc_289 N_A1_c_302_n N_Y_c_677_n 0.0112464f $X=5.4 $Y=1.185 $X2=0 $Y2=0
cc_290 N_A1_c_303_n N_Y_c_677_n 0.0080264f $X=5.83 $Y=1.185 $X2=0 $Y2=0
cc_291 A1 N_Y_c_677_n 0.113138f $X=5.435 $Y=1.21 $X2=0 $Y2=0
cc_292 N_A1_c_305_n N_Y_c_677_n 0.0194978f $X=5.73 $Y=1.425 $X2=0 $Y2=0
cc_293 N_A1_M1003_g N_VPWR_c_805_n 0.0132143f $X=4.1 $Y=2.465 $X2=0 $Y2=0
cc_294 N_A1_M1012_g N_VPWR_c_805_n 0.0119098f $X=4.53 $Y=2.465 $X2=0 $Y2=0
cc_295 N_A1_M1034_g N_VPWR_c_805_n 6.42299e-19 $X=4.96 $Y=2.465 $X2=0 $Y2=0
cc_296 N_A1_M1012_g N_VPWR_c_806_n 0.00486043f $X=4.53 $Y=2.465 $X2=0 $Y2=0
cc_297 N_A1_M1034_g N_VPWR_c_806_n 0.00486043f $X=4.96 $Y=2.465 $X2=0 $Y2=0
cc_298 N_A1_M1012_g N_VPWR_c_807_n 6.41962e-19 $X=4.53 $Y=2.465 $X2=0 $Y2=0
cc_299 N_A1_M1034_g N_VPWR_c_807_n 0.0120894f $X=4.96 $Y=2.465 $X2=0 $Y2=0
cc_300 N_A1_M1039_g N_VPWR_c_807_n 0.0120894f $X=5.73 $Y=2.465 $X2=0 $Y2=0
cc_301 N_A1_M1039_g N_VPWR_c_808_n 6.56457e-19 $X=5.73 $Y=2.465 $X2=0 $Y2=0
cc_302 N_A1_M1003_g N_VPWR_c_813_n 0.00486043f $X=4.1 $Y=2.465 $X2=0 $Y2=0
cc_303 N_A1_M1039_g N_VPWR_c_815_n 0.00486043f $X=5.73 $Y=2.465 $X2=0 $Y2=0
cc_304 N_A1_M1003_g N_VPWR_c_804_n 0.00851476f $X=4.1 $Y=2.465 $X2=0 $Y2=0
cc_305 N_A1_M1012_g N_VPWR_c_804_n 0.00824727f $X=4.53 $Y=2.465 $X2=0 $Y2=0
cc_306 N_A1_M1034_g N_VPWR_c_804_n 0.00824727f $X=4.96 $Y=2.465 $X2=0 $Y2=0
cc_307 N_A1_M1039_g N_VPWR_c_804_n 0.0082726f $X=5.73 $Y=2.465 $X2=0 $Y2=0
cc_308 N_A1_c_300_n N_VGND_c_997_n 0.00359964f $X=4.54 $Y=1.185 $X2=0 $Y2=0
cc_309 N_A1_c_301_n N_VGND_c_997_n 0.00359964f $X=4.97 $Y=1.185 $X2=0 $Y2=0
cc_310 N_A1_c_302_n N_VGND_c_997_n 0.00359964f $X=5.4 $Y=1.185 $X2=0 $Y2=0
cc_311 N_A1_c_303_n N_VGND_c_997_n 0.00359964f $X=5.83 $Y=1.185 $X2=0 $Y2=0
cc_312 N_A1_c_300_n N_VGND_c_1004_n 0.00665257f $X=4.54 $Y=1.185 $X2=0 $Y2=0
cc_313 N_A1_c_301_n N_VGND_c_1004_n 0.00535287f $X=4.97 $Y=1.185 $X2=0 $Y2=0
cc_314 N_A1_c_302_n N_VGND_c_1004_n 0.00535287f $X=5.4 $Y=1.185 $X2=0 $Y2=0
cc_315 N_A1_c_303_n N_VGND_c_1004_n 0.00537821f $X=5.83 $Y=1.185 $X2=0 $Y2=0
cc_316 N_A1_c_300_n N_A_840_47#_c_1110_n 0.0119698f $X=4.54 $Y=1.185 $X2=0 $Y2=0
cc_317 N_A1_c_301_n N_A_840_47#_c_1110_n 0.0119698f $X=4.97 $Y=1.185 $X2=0 $Y2=0
cc_318 N_A1_c_302_n N_A_840_47#_c_1110_n 0.0119698f $X=5.4 $Y=1.185 $X2=0 $Y2=0
cc_319 N_A1_c_303_n N_A_840_47#_c_1110_n 0.011969f $X=5.83 $Y=1.185 $X2=0 $Y2=0
cc_320 N_A1_c_303_n N_A_1267_47#_c_1143_n 2.17945e-19 $X=5.83 $Y=1.185 $X2=0
+ $Y2=0
cc_321 A2 A3 0.0137205f $X=7.835 $Y=1.21 $X2=0 $Y2=0
cc_322 N_A2_c_380_n A3 9.94636e-19 $X=7.79 $Y=1.35 $X2=0 $Y2=0
cc_323 N_A2_M1029_g N_A3_c_458_n 0.0273985f $X=7.81 $Y=2.465 $X2=0 $Y2=0
cc_324 A2 N_A3_c_458_n 8.86223e-19 $X=7.835 $Y=1.21 $X2=0 $Y2=0
cc_325 N_A2_c_380_n N_A3_c_458_n 0.0091505f $X=7.79 $Y=1.35 $X2=0 $Y2=0
cc_326 N_A2_c_381_n N_A_42_367#_c_561_n 0.0181224f $X=6.16 $Y=1.725 $X2=0 $Y2=0
cc_327 N_A2_M1017_g N_A_42_367#_c_561_n 0.0139144f $X=6.95 $Y=2.465 $X2=0 $Y2=0
cc_328 A2 N_A_42_367#_c_561_n 0.0178983f $X=7.835 $Y=1.21 $X2=0 $Y2=0
cc_329 N_A2_c_380_n N_A_42_367#_c_561_n 0.00928151f $X=7.79 $Y=1.35 $X2=0 $Y2=0
cc_330 N_A2_M1017_g N_A_42_367#_c_536_n 0.0118539f $X=6.95 $Y=2.465 $X2=0 $Y2=0
cc_331 N_A2_M1022_g N_A_42_367#_c_536_n 8.32811e-19 $X=7.38 $Y=2.465 $X2=0 $Y2=0
cc_332 N_A2_M1022_g N_A_42_367#_c_529_n 0.0143398f $X=7.38 $Y=2.465 $X2=0 $Y2=0
cc_333 N_A2_M1029_g N_A_42_367#_c_529_n 0.0142932f $X=7.81 $Y=2.465 $X2=0 $Y2=0
cc_334 A2 N_A_42_367#_c_529_n 0.0477254f $X=7.835 $Y=1.21 $X2=0 $Y2=0
cc_335 N_A2_c_380_n N_A_42_367#_c_529_n 0.00391511f $X=7.79 $Y=1.35 $X2=0 $Y2=0
cc_336 N_A2_M1017_g N_A_42_367#_c_530_n 0.0076428f $X=6.95 $Y=2.465 $X2=0 $Y2=0
cc_337 A2 N_A_42_367#_c_530_n 0.0212131f $X=7.835 $Y=1.21 $X2=0 $Y2=0
cc_338 N_A2_c_380_n N_A_42_367#_c_530_n 0.00354402f $X=7.79 $Y=1.35 $X2=0 $Y2=0
cc_339 N_A2_M1029_g N_A_42_367#_c_538_n 0.00152323f $X=7.81 $Y=2.465 $X2=0 $Y2=0
cc_340 N_A2_M1017_g N_A_42_367#_c_575_n 0.00234635f $X=6.95 $Y=2.465 $X2=0 $Y2=0
cc_341 A2 N_A_42_367#_c_533_n 0.00635961f $X=7.835 $Y=1.21 $X2=0 $Y2=0
cc_342 N_A2_c_380_n N_A_42_367#_c_533_n 6.41898e-19 $X=7.79 $Y=1.35 $X2=0 $Y2=0
cc_343 N_A2_c_381_n N_Y_c_672_n 0.00873161f $X=6.16 $Y=1.725 $X2=0 $Y2=0
cc_344 N_A2_c_380_n N_Y_c_672_n 0.00707792f $X=7.79 $Y=1.35 $X2=0 $Y2=0
cc_345 N_A2_c_372_n N_Y_c_737_n 0.00234085f $X=6.26 $Y=1.185 $X2=0 $Y2=0
cc_346 N_A2_c_372_n N_Y_c_673_n 0.00980241f $X=6.26 $Y=1.185 $X2=0 $Y2=0
cc_347 A2 N_Y_c_673_n 0.0180945f $X=7.835 $Y=1.21 $X2=0 $Y2=0
cc_348 N_A2_c_380_n N_Y_c_673_n 0.00167014f $X=7.79 $Y=1.35 $X2=0 $Y2=0
cc_349 N_A2_c_381_n N_VPWR_c_807_n 6.41962e-19 $X=6.16 $Y=1.725 $X2=0 $Y2=0
cc_350 N_A2_c_381_n N_VPWR_c_808_n 0.0135096f $X=6.16 $Y=1.725 $X2=0 $Y2=0
cc_351 N_A2_M1017_g N_VPWR_c_808_n 0.0135096f $X=6.95 $Y=2.465 $X2=0 $Y2=0
cc_352 N_A2_M1022_g N_VPWR_c_808_n 6.56457e-19 $X=7.38 $Y=2.465 $X2=0 $Y2=0
cc_353 N_A2_M1017_g N_VPWR_c_809_n 0.00486043f $X=6.95 $Y=2.465 $X2=0 $Y2=0
cc_354 N_A2_M1022_g N_VPWR_c_809_n 0.00486043f $X=7.38 $Y=2.465 $X2=0 $Y2=0
cc_355 N_A2_M1017_g N_VPWR_c_810_n 8.01113e-19 $X=6.95 $Y=2.465 $X2=0 $Y2=0
cc_356 N_A2_M1022_g N_VPWR_c_810_n 0.0174f $X=7.38 $Y=2.465 $X2=0 $Y2=0
cc_357 N_A2_M1029_g N_VPWR_c_810_n 0.01742f $X=7.81 $Y=2.465 $X2=0 $Y2=0
cc_358 N_A2_M1029_g N_VPWR_c_811_n 7.69607e-19 $X=7.81 $Y=2.465 $X2=0 $Y2=0
cc_359 N_A2_c_381_n N_VPWR_c_815_n 0.00486043f $X=6.16 $Y=1.725 $X2=0 $Y2=0
cc_360 N_A2_M1029_g N_VPWR_c_816_n 0.00486043f $X=7.81 $Y=2.465 $X2=0 $Y2=0
cc_361 N_A2_c_381_n N_VPWR_c_804_n 0.0082726f $X=6.16 $Y=1.725 $X2=0 $Y2=0
cc_362 N_A2_M1017_g N_VPWR_c_804_n 0.00824727f $X=6.95 $Y=2.465 $X2=0 $Y2=0
cc_363 N_A2_M1022_g N_VPWR_c_804_n 0.00824727f $X=7.38 $Y=2.465 $X2=0 $Y2=0
cc_364 N_A2_M1029_g N_VPWR_c_804_n 0.0082726f $X=7.81 $Y=2.465 $X2=0 $Y2=0
cc_365 N_A2_c_377_n N_VGND_c_993_n 0.00245808f $X=7.55 $Y=1.185 $X2=0 $Y2=0
cc_366 N_A2_c_372_n N_VGND_c_997_n 0.00359964f $X=6.26 $Y=1.185 $X2=0 $Y2=0
cc_367 N_A2_c_373_n N_VGND_c_997_n 0.00359964f $X=6.69 $Y=1.185 $X2=0 $Y2=0
cc_368 N_A2_c_375_n N_VGND_c_997_n 0.00359964f $X=7.12 $Y=1.185 $X2=0 $Y2=0
cc_369 N_A2_c_377_n N_VGND_c_997_n 0.00359964f $X=7.55 $Y=1.185 $X2=0 $Y2=0
cc_370 N_A2_c_372_n N_VGND_c_1004_n 0.00537821f $X=6.26 $Y=1.185 $X2=0 $Y2=0
cc_371 N_A2_c_373_n N_VGND_c_1004_n 0.00535287f $X=6.69 $Y=1.185 $X2=0 $Y2=0
cc_372 N_A2_c_375_n N_VGND_c_1004_n 0.00535287f $X=7.12 $Y=1.185 $X2=0 $Y2=0
cc_373 N_A2_c_377_n N_VGND_c_1004_n 0.00665257f $X=7.55 $Y=1.185 $X2=0 $Y2=0
cc_374 N_A2_c_372_n N_A_840_47#_c_1110_n 0.0152783f $X=6.26 $Y=1.185 $X2=0 $Y2=0
cc_375 N_A2_c_373_n N_A_840_47#_c_1110_n 0.0119698f $X=6.69 $Y=1.185 $X2=0 $Y2=0
cc_376 N_A2_c_375_n N_A_840_47#_c_1110_n 0.0119698f $X=7.12 $Y=1.185 $X2=0 $Y2=0
cc_377 N_A2_c_377_n N_A_840_47#_c_1110_n 0.0119698f $X=7.55 $Y=1.185 $X2=0 $Y2=0
cc_378 A2 N_A_840_47#_c_1110_n 0.00113001f $X=7.835 $Y=1.21 $X2=0 $Y2=0
cc_379 N_A2_c_372_n N_A_1267_47#_c_1143_n 0.00371663f $X=6.26 $Y=1.185 $X2=0
+ $Y2=0
cc_380 N_A2_c_373_n N_A_1267_47#_c_1143_n 0.0112464f $X=6.69 $Y=1.185 $X2=0
+ $Y2=0
cc_381 N_A2_c_375_n N_A_1267_47#_c_1143_n 0.0112464f $X=7.12 $Y=1.185 $X2=0
+ $Y2=0
cc_382 N_A2_c_377_n N_A_1267_47#_c_1143_n 0.0145623f $X=7.55 $Y=1.185 $X2=0
+ $Y2=0
cc_383 A2 N_A_1267_47#_c_1143_n 0.109564f $X=7.835 $Y=1.21 $X2=0 $Y2=0
cc_384 N_A2_c_380_n N_A_1267_47#_c_1143_n 0.0163501f $X=7.79 $Y=1.35 $X2=0 $Y2=0
cc_385 N_A3_M1000_g N_A_42_367#_c_538_n 0.00152323f $X=8.24 $Y=2.465 $X2=0 $Y2=0
cc_386 N_A3_M1000_g N_A_42_367#_c_531_n 0.00997588f $X=8.24 $Y=2.465 $X2=0 $Y2=0
cc_387 N_A3_M1007_g N_A_42_367#_c_531_n 0.0100058f $X=8.67 $Y=2.465 $X2=0 $Y2=0
cc_388 A3 N_A_42_367#_c_531_n 0.0332975f $X=10.235 $Y=1.21 $X2=0 $Y2=0
cc_389 N_A3_c_458_n N_A_42_367#_c_531_n 0.014209f $X=9.865 $Y=1.35 $X2=0 $Y2=0
cc_390 N_A3_M1007_g N_A_42_367#_c_540_n 0.0014373f $X=8.67 $Y=2.465 $X2=0 $Y2=0
cc_391 N_A3_M1018_g N_A_42_367#_c_540_n 0.0014373f $X=9.1 $Y=2.465 $X2=0 $Y2=0
cc_392 N_A3_M1018_g N_A_42_367#_c_532_n 0.0100058f $X=9.1 $Y=2.465 $X2=0 $Y2=0
cc_393 N_A3_M1026_g N_A_42_367#_c_532_n 0.0108978f $X=9.53 $Y=2.465 $X2=0 $Y2=0
cc_394 A3 N_A_42_367#_c_532_n 0.0678391f $X=10.235 $Y=1.21 $X2=0 $Y2=0
cc_395 N_A3_c_458_n N_A_42_367#_c_532_n 0.0236381f $X=9.865 $Y=1.35 $X2=0 $Y2=0
cc_396 N_A3_M1026_g N_A_42_367#_c_542_n 0.0046421f $X=9.53 $Y=2.465 $X2=0 $Y2=0
cc_397 A3 N_A_42_367#_c_590_n 0.0147582f $X=10.235 $Y=1.21 $X2=0 $Y2=0
cc_398 N_A3_c_458_n N_A_42_367#_c_590_n 0.00634147f $X=9.865 $Y=1.35 $X2=0 $Y2=0
cc_399 N_A3_M1000_g N_VPWR_c_810_n 7.69607e-19 $X=8.24 $Y=2.465 $X2=0 $Y2=0
cc_400 N_A3_M1000_g N_VPWR_c_811_n 0.01742f $X=8.24 $Y=2.465 $X2=0 $Y2=0
cc_401 N_A3_M1007_g N_VPWR_c_811_n 0.01742f $X=8.67 $Y=2.465 $X2=0 $Y2=0
cc_402 N_A3_M1018_g N_VPWR_c_811_n 7.69607e-19 $X=9.1 $Y=2.465 $X2=0 $Y2=0
cc_403 N_A3_c_458_n N_VPWR_c_811_n 5.98711e-19 $X=9.865 $Y=1.35 $X2=0 $Y2=0
cc_404 N_A3_M1007_g N_VPWR_c_812_n 7.69607e-19 $X=8.67 $Y=2.465 $X2=0 $Y2=0
cc_405 N_A3_M1018_g N_VPWR_c_812_n 0.01742f $X=9.1 $Y=2.465 $X2=0 $Y2=0
cc_406 N_A3_M1026_g N_VPWR_c_812_n 0.0194824f $X=9.53 $Y=2.465 $X2=0 $Y2=0
cc_407 N_A3_c_458_n N_VPWR_c_812_n 5.95909e-19 $X=9.865 $Y=1.35 $X2=0 $Y2=0
cc_408 N_A3_M1000_g N_VPWR_c_816_n 0.00486043f $X=8.24 $Y=2.465 $X2=0 $Y2=0
cc_409 N_A3_M1007_g N_VPWR_c_817_n 0.00486043f $X=8.67 $Y=2.465 $X2=0 $Y2=0
cc_410 N_A3_M1018_g N_VPWR_c_817_n 0.00486043f $X=9.1 $Y=2.465 $X2=0 $Y2=0
cc_411 N_A3_M1026_g N_VPWR_c_818_n 0.00486043f $X=9.53 $Y=2.465 $X2=0 $Y2=0
cc_412 N_A3_M1000_g N_VPWR_c_804_n 0.0082726f $X=8.24 $Y=2.465 $X2=0 $Y2=0
cc_413 N_A3_M1007_g N_VPWR_c_804_n 0.00824727f $X=8.67 $Y=2.465 $X2=0 $Y2=0
cc_414 N_A3_M1018_g N_VPWR_c_804_n 0.00824727f $X=9.1 $Y=2.465 $X2=0 $Y2=0
cc_415 N_A3_M1026_g N_VPWR_c_804_n 0.00954696f $X=9.53 $Y=2.465 $X2=0 $Y2=0
cc_416 N_A3_c_453_n N_VGND_c_993_n 0.00946465f $X=8.5 $Y=1.185 $X2=0 $Y2=0
cc_417 N_A3_c_454_n N_VGND_c_993_n 5.4611e-19 $X=8.93 $Y=1.185 $X2=0 $Y2=0
cc_418 N_A3_c_453_n N_VGND_c_994_n 5.4611e-19 $X=8.5 $Y=1.185 $X2=0 $Y2=0
cc_419 N_A3_c_454_n N_VGND_c_994_n 0.00823407f $X=8.93 $Y=1.185 $X2=0 $Y2=0
cc_420 N_A3_c_455_n N_VGND_c_994_n 0.00823407f $X=9.36 $Y=1.185 $X2=0 $Y2=0
cc_421 N_A3_c_456_n N_VGND_c_994_n 5.4611e-19 $X=9.79 $Y=1.185 $X2=0 $Y2=0
cc_422 N_A3_c_455_n N_VGND_c_995_n 0.00486043f $X=9.36 $Y=1.185 $X2=0 $Y2=0
cc_423 N_A3_c_456_n N_VGND_c_995_n 0.00486043f $X=9.79 $Y=1.185 $X2=0 $Y2=0
cc_424 N_A3_c_455_n N_VGND_c_996_n 6.08631e-19 $X=9.36 $Y=1.185 $X2=0 $Y2=0
cc_425 N_A3_c_456_n N_VGND_c_996_n 0.0165361f $X=9.79 $Y=1.185 $X2=0 $Y2=0
cc_426 A3 N_VGND_c_996_n 0.0237475f $X=10.235 $Y=1.21 $X2=0 $Y2=0
cc_427 N_A3_c_459_n N_VGND_c_996_n 0.00709505f $X=10.29 $Y=1.35 $X2=0 $Y2=0
cc_428 N_A3_c_453_n N_VGND_c_999_n 0.00486043f $X=8.5 $Y=1.185 $X2=0 $Y2=0
cc_429 N_A3_c_454_n N_VGND_c_999_n 0.00486043f $X=8.93 $Y=1.185 $X2=0 $Y2=0
cc_430 N_A3_c_453_n N_VGND_c_1004_n 0.00438495f $X=8.5 $Y=1.185 $X2=0 $Y2=0
cc_431 N_A3_c_454_n N_VGND_c_1004_n 0.00448921f $X=8.93 $Y=1.185 $X2=0 $Y2=0
cc_432 N_A3_c_455_n N_VGND_c_1004_n 0.00448921f $X=9.36 $Y=1.185 $X2=0 $Y2=0
cc_433 N_A3_c_456_n N_VGND_c_1004_n 0.00824727f $X=9.79 $Y=1.185 $X2=0 $Y2=0
cc_434 N_A3_c_453_n N_A_840_47#_c_1110_n 6.17781e-19 $X=8.5 $Y=1.185 $X2=0 $Y2=0
cc_435 N_A3_c_453_n N_A_1267_47#_c_1143_n 0.0156969f $X=8.5 $Y=1.185 $X2=0 $Y2=0
cc_436 A3 N_A_1267_47#_c_1143_n 0.0187267f $X=10.235 $Y=1.21 $X2=0 $Y2=0
cc_437 N_A3_c_458_n N_A_1267_47#_c_1143_n 0.00331754f $X=9.865 $Y=1.35 $X2=0
+ $Y2=0
cc_438 N_A3_c_454_n N_A_1267_47#_c_1154_n 0.0112011f $X=8.93 $Y=1.185 $X2=0
+ $Y2=0
cc_439 N_A3_c_455_n N_A_1267_47#_c_1154_n 0.0112768f $X=9.36 $Y=1.185 $X2=0
+ $Y2=0
cc_440 A3 N_A_1267_47#_c_1154_n 0.0547422f $X=10.235 $Y=1.21 $X2=0 $Y2=0
cc_441 N_A3_c_458_n N_A_1267_47#_c_1154_n 0.00545404f $X=9.865 $Y=1.35 $X2=0
+ $Y2=0
cc_442 A3 N_A_1267_47#_c_1158_n 0.0142048f $X=10.235 $Y=1.21 $X2=0 $Y2=0
cc_443 N_A3_c_458_n N_A_1267_47#_c_1158_n 0.00280606f $X=9.865 $Y=1.35 $X2=0
+ $Y2=0
cc_444 N_A_42_367#_c_546_n N_Y_M1006_s 0.00332344f $X=1.1 $Y=2.99 $X2=0 $Y2=0
cc_445 N_A_42_367#_c_548_n N_Y_M1021_s 0.00332344f $X=1.96 $Y=2.99 $X2=0 $Y2=0
cc_446 N_A_42_367#_c_550_n N_Y_M1001_d 0.00332344f $X=2.82 $Y=2.99 $X2=0 $Y2=0
cc_447 N_A_42_367#_c_552_n N_Y_M1019_d 0.00332344f $X=3.68 $Y=2.99 $X2=0 $Y2=0
cc_448 N_A_42_367#_c_546_n N_Y_c_678_n 0.0159805f $X=1.1 $Y=2.99 $X2=0 $Y2=0
cc_449 N_A_42_367#_M1020_d N_Y_c_668_n 0.00178994f $X=1.055 $Y=1.835 $X2=0 $Y2=0
cc_450 N_A_42_367#_c_598_p N_Y_c_668_n 0.0139398f $X=1.195 $Y=2.21 $X2=0 $Y2=0
cc_451 N_A_42_367#_c_535_n N_Y_c_669_n 0.00246889f $X=0.335 $Y=1.99 $X2=0 $Y2=0
cc_452 N_A_42_367#_c_548_n N_Y_c_689_n 0.0159805f $X=1.96 $Y=2.99 $X2=0 $Y2=0
cc_453 N_A_42_367#_M1032_d N_Y_c_670_n 0.00178994f $X=1.915 $Y=1.835 $X2=0 $Y2=0
cc_454 N_A_42_367#_c_602_p N_Y_c_670_n 0.0139398f $X=2.055 $Y=2.21 $X2=0 $Y2=0
cc_455 N_A_42_367#_c_550_n N_Y_c_694_n 0.0159805f $X=2.82 $Y=2.99 $X2=0 $Y2=0
cc_456 N_A_42_367#_M1015_s N_Y_c_671_n 0.00178994f $X=2.775 $Y=1.835 $X2=0 $Y2=0
cc_457 N_A_42_367#_c_605_p N_Y_c_671_n 0.0139398f $X=2.915 $Y=2.21 $X2=0 $Y2=0
cc_458 N_A_42_367#_c_552_n N_Y_c_710_n 0.0159805f $X=3.68 $Y=2.99 $X2=0 $Y2=0
cc_459 N_A_42_367#_M1033_s N_Y_c_672_n 0.0030408f $X=3.635 $Y=1.835 $X2=0 $Y2=0
cc_460 N_A_42_367#_M1012_s N_Y_c_672_n 0.00178994f $X=4.605 $Y=1.835 $X2=0 $Y2=0
cc_461 N_A_42_367#_M1039_s N_Y_c_672_n 0.00181969f $X=5.805 $Y=1.835 $X2=0 $Y2=0
cc_462 N_A_42_367#_c_610_p N_Y_c_672_n 0.023177f $X=3.83 $Y=2.225 $X2=0 $Y2=0
cc_463 N_A_42_367#_c_554_n N_Y_c_672_n 0.0336459f $X=4.65 $Y=2.135 $X2=0 $Y2=0
cc_464 N_A_42_367#_c_557_n N_Y_c_672_n 0.0593331f $X=5.85 $Y=2.135 $X2=0 $Y2=0
cc_465 N_A_42_367#_c_561_n N_Y_c_672_n 7.3041e-19 $X=7 $Y=2.135 $X2=0 $Y2=0
cc_466 N_A_42_367#_c_560_n N_Y_c_672_n 0.0139398f $X=4.745 $Y=2.21 $X2=0 $Y2=0
cc_467 N_A_42_367#_c_615_p N_Y_c_672_n 0.0147855f $X=5.945 $Y=2.21 $X2=0 $Y2=0
cc_468 N_A_42_367#_c_554_n N_VPWR_M1003_d 0.0033818f $X=4.65 $Y=2.135 $X2=-0.19
+ $Y2=-0.245
cc_469 N_A_42_367#_c_557_n N_VPWR_M1034_d 0.0132993f $X=5.85 $Y=2.135 $X2=0
+ $Y2=0
cc_470 N_A_42_367#_c_561_n N_VPWR_M1004_s 0.0175711f $X=7 $Y=2.135 $X2=0 $Y2=0
cc_471 N_A_42_367#_c_554_n N_VPWR_c_805_n 0.0171443f $X=4.65 $Y=2.135 $X2=0
+ $Y2=0
cc_472 N_A_42_367#_c_620_p N_VPWR_c_806_n 0.0124525f $X=4.745 $Y=2.91 $X2=0
+ $Y2=0
cc_473 N_A_42_367#_c_557_n N_VPWR_c_807_n 0.0370354f $X=5.85 $Y=2.135 $X2=0
+ $Y2=0
cc_474 N_A_42_367#_c_561_n N_VPWR_c_808_n 0.0465465f $X=7 $Y=2.135 $X2=0 $Y2=0
cc_475 N_A_42_367#_c_623_p N_VPWR_c_809_n 0.0124525f $X=7.165 $Y=2.465 $X2=0
+ $Y2=0
cc_476 N_A_42_367#_c_529_n N_VPWR_c_810_n 0.0216087f $X=7.93 $Y=1.69 $X2=0 $Y2=0
cc_477 N_A_42_367#_c_531_n N_VPWR_c_811_n 0.0216087f $X=8.79 $Y=1.69 $X2=0 $Y2=0
cc_478 N_A_42_367#_c_532_n N_VPWR_c_812_n 0.0216087f $X=9.65 $Y=1.69 $X2=0 $Y2=0
cc_479 N_A_42_367#_c_534_n N_VPWR_c_813_n 0.0179183f $X=0.3 $Y=2.905 $X2=0 $Y2=0
cc_480 N_A_42_367#_c_546_n N_VPWR_c_813_n 0.0361172f $X=1.1 $Y=2.99 $X2=0 $Y2=0
cc_481 N_A_42_367#_c_548_n N_VPWR_c_813_n 0.0361172f $X=1.96 $Y=2.99 $X2=0 $Y2=0
cc_482 N_A_42_367#_c_550_n N_VPWR_c_813_n 0.0361172f $X=2.82 $Y=2.99 $X2=0 $Y2=0
cc_483 N_A_42_367#_c_552_n N_VPWR_c_813_n 0.0361172f $X=3.68 $Y=2.99 $X2=0 $Y2=0
cc_484 N_A_42_367#_c_632_p N_VPWR_c_813_n 0.0202578f $X=3.83 $Y=2.905 $X2=0
+ $Y2=0
cc_485 N_A_42_367#_c_633_p N_VPWR_c_813_n 0.0125234f $X=1.195 $Y=2.91 $X2=0
+ $Y2=0
cc_486 N_A_42_367#_c_634_p N_VPWR_c_813_n 0.0125234f $X=2.055 $Y=2.91 $X2=0
+ $Y2=0
cc_487 N_A_42_367#_c_635_p N_VPWR_c_813_n 0.0125234f $X=2.915 $Y=2.91 $X2=0
+ $Y2=0
cc_488 N_A_42_367#_c_636_p N_VPWR_c_815_n 0.0124525f $X=5.945 $Y=2.91 $X2=0
+ $Y2=0
cc_489 N_A_42_367#_c_538_n N_VPWR_c_816_n 0.0124525f $X=8.025 $Y=1.96 $X2=0
+ $Y2=0
cc_490 N_A_42_367#_c_540_n N_VPWR_c_817_n 0.0124525f $X=8.885 $Y=1.98 $X2=0
+ $Y2=0
cc_491 N_A_42_367#_c_542_n N_VPWR_c_818_n 0.0178111f $X=9.745 $Y=1.98 $X2=0
+ $Y2=0
cc_492 N_A_42_367#_M1006_d N_VPWR_c_804_n 0.00215161f $X=0.21 $Y=1.835 $X2=0
+ $Y2=0
cc_493 N_A_42_367#_M1020_d N_VPWR_c_804_n 0.00223565f $X=1.055 $Y=1.835 $X2=0
+ $Y2=0
cc_494 N_A_42_367#_M1032_d N_VPWR_c_804_n 0.00223565f $X=1.915 $Y=1.835 $X2=0
+ $Y2=0
cc_495 N_A_42_367#_M1015_s N_VPWR_c_804_n 0.00223565f $X=2.775 $Y=1.835 $X2=0
+ $Y2=0
cc_496 N_A_42_367#_M1033_s N_VPWR_c_804_n 0.00466094f $X=3.635 $Y=1.835 $X2=0
+ $Y2=0
cc_497 N_A_42_367#_M1012_s N_VPWR_c_804_n 0.00536646f $X=4.605 $Y=1.835 $X2=0
+ $Y2=0
cc_498 N_A_42_367#_M1039_s N_VPWR_c_804_n 0.00536646f $X=5.805 $Y=1.835 $X2=0
+ $Y2=0
cc_499 N_A_42_367#_M1017_d N_VPWR_c_804_n 0.00536646f $X=7.025 $Y=1.835 $X2=0
+ $Y2=0
cc_500 N_A_42_367#_M1029_d N_VPWR_c_804_n 0.00536646f $X=7.885 $Y=1.835 $X2=0
+ $Y2=0
cc_501 N_A_42_367#_M1007_s N_VPWR_c_804_n 0.00536646f $X=8.745 $Y=1.835 $X2=0
+ $Y2=0
cc_502 N_A_42_367#_M1026_s N_VPWR_c_804_n 0.00371702f $X=9.605 $Y=1.835 $X2=0
+ $Y2=0
cc_503 N_A_42_367#_c_534_n N_VPWR_c_804_n 0.0101029f $X=0.3 $Y=2.905 $X2=0 $Y2=0
cc_504 N_A_42_367#_c_546_n N_VPWR_c_804_n 0.023676f $X=1.1 $Y=2.99 $X2=0 $Y2=0
cc_505 N_A_42_367#_c_548_n N_VPWR_c_804_n 0.023676f $X=1.96 $Y=2.99 $X2=0 $Y2=0
cc_506 N_A_42_367#_c_550_n N_VPWR_c_804_n 0.023676f $X=2.82 $Y=2.99 $X2=0 $Y2=0
cc_507 N_A_42_367#_c_552_n N_VPWR_c_804_n 0.023676f $X=3.68 $Y=2.99 $X2=0 $Y2=0
cc_508 N_A_42_367#_c_632_p N_VPWR_c_804_n 0.0116633f $X=3.83 $Y=2.905 $X2=0
+ $Y2=0
cc_509 N_A_42_367#_c_620_p N_VPWR_c_804_n 0.00730901f $X=4.745 $Y=2.91 $X2=0
+ $Y2=0
cc_510 N_A_42_367#_c_636_p N_VPWR_c_804_n 0.00730901f $X=5.945 $Y=2.91 $X2=0
+ $Y2=0
cc_511 N_A_42_367#_c_623_p N_VPWR_c_804_n 0.00730901f $X=7.165 $Y=2.465 $X2=0
+ $Y2=0
cc_512 N_A_42_367#_c_538_n N_VPWR_c_804_n 0.00730901f $X=8.025 $Y=1.96 $X2=0
+ $Y2=0
cc_513 N_A_42_367#_c_540_n N_VPWR_c_804_n 0.00730901f $X=8.885 $Y=1.98 $X2=0
+ $Y2=0
cc_514 N_A_42_367#_c_542_n N_VPWR_c_804_n 0.0100304f $X=9.745 $Y=1.98 $X2=0
+ $Y2=0
cc_515 N_A_42_367#_c_633_p N_VPWR_c_804_n 0.00738676f $X=1.195 $Y=2.91 $X2=0
+ $Y2=0
cc_516 N_A_42_367#_c_634_p N_VPWR_c_804_n 0.00738676f $X=2.055 $Y=2.91 $X2=0
+ $Y2=0
cc_517 N_A_42_367#_c_635_p N_VPWR_c_804_n 0.00738676f $X=2.915 $Y=2.91 $X2=0
+ $Y2=0
cc_518 N_A_42_367#_c_531_n N_A_1267_47#_c_1143_n 0.00578749f $X=8.79 $Y=1.69
+ $X2=0 $Y2=0
cc_519 N_A_42_367#_c_533_n N_A_1267_47#_c_1143_n 0.00435179f $X=8.025 $Y=1.69
+ $X2=0 $Y2=0
cc_520 N_Y_c_672_n N_VPWR_M1003_d 0.00179431f $X=5.885 $Y=1.74 $X2=-0.19
+ $Y2=-0.245
cc_521 N_Y_c_672_n N_VPWR_M1034_d 0.00588674f $X=5.885 $Y=1.74 $X2=0 $Y2=0
cc_522 N_Y_M1006_s N_VPWR_c_804_n 0.00225186f $X=0.625 $Y=1.835 $X2=0 $Y2=0
cc_523 N_Y_M1021_s N_VPWR_c_804_n 0.00225186f $X=1.485 $Y=1.835 $X2=0 $Y2=0
cc_524 N_Y_M1001_d N_VPWR_c_804_n 0.00225186f $X=2.345 $Y=1.835 $X2=0 $Y2=0
cc_525 N_Y_M1019_d N_VPWR_c_804_n 0.00225186f $X=3.205 $Y=1.835 $X2=0 $Y2=0
cc_526 N_Y_c_677_n N_A_28_47#_M1023_s 0.00331529f $X=5.885 $Y=0.902 $X2=0 $Y2=0
cc_527 N_Y_c_677_n N_A_28_47#_M1038_s 0.00534708f $X=5.885 $Y=0.902 $X2=0 $Y2=0
cc_528 N_Y_c_670_n N_A_28_47#_c_959_n 0.00618711f $X=2.32 $Y=1.74 $X2=0 $Y2=0
cc_529 N_Y_M1010_d N_A_28_47#_c_948_n 0.00330375f $X=2.275 $Y=0.235 $X2=0 $Y2=0
cc_530 N_Y_M1024_d N_A_28_47#_c_948_n 0.00330375f $X=3.135 $Y=0.235 $X2=0 $Y2=0
cc_531 N_Y_c_677_n N_A_28_47#_c_948_n 0.0912146f $X=5.885 $Y=0.902 $X2=0 $Y2=0
cc_532 N_Y_M1010_d N_VGND_c_1004_n 0.00225186f $X=2.275 $Y=0.235 $X2=0 $Y2=0
cc_533 N_Y_M1024_d N_VGND_c_1004_n 0.00225186f $X=3.135 $Y=0.235 $X2=0 $Y2=0
cc_534 N_Y_M1005_d N_VGND_c_1004_n 0.00225465f $X=4.615 $Y=0.235 $X2=0 $Y2=0
cc_535 N_Y_M1027_d N_VGND_c_1004_n 0.00225465f $X=5.475 $Y=0.235 $X2=0 $Y2=0
cc_536 N_Y_c_677_n N_VGND_c_1004_n 0.0166261f $X=5.885 $Y=0.902 $X2=0 $Y2=0
cc_537 N_Y_c_677_n N_A_840_47#_M1005_s 0.00520331f $X=5.885 $Y=0.902 $X2=-0.19
+ $Y2=-0.245
cc_538 N_Y_c_677_n N_A_840_47#_M1014_s 0.00331529f $X=5.885 $Y=0.902 $X2=0 $Y2=0
cc_539 N_Y_c_737_n N_A_840_47#_M1037_s 0.0041329f $X=5.99 $Y=1.04 $X2=0 $Y2=0
cc_540 N_Y_c_673_n N_A_840_47#_M1037_s 3.87548e-19 $X=5.99 $Y=1.605 $X2=0 $Y2=0
cc_541 N_Y_M1005_d N_A_840_47#_c_1110_n 0.00333618f $X=4.615 $Y=0.235 $X2=0
+ $Y2=0
cc_542 N_Y_M1027_d N_A_840_47#_c_1110_n 0.00333618f $X=5.475 $Y=0.235 $X2=0
+ $Y2=0
cc_543 N_Y_c_737_n N_A_840_47#_c_1110_n 0.0124428f $X=5.99 $Y=1.04 $X2=0 $Y2=0
cc_544 N_Y_c_677_n N_A_840_47#_c_1110_n 0.0984845f $X=5.885 $Y=0.902 $X2=0 $Y2=0
cc_545 N_Y_c_737_n N_A_1267_47#_c_1143_n 0.0198799f $X=5.99 $Y=1.04 $X2=0 $Y2=0
cc_546 N_A_28_47#_c_949_n N_VGND_M1002_d 0.00329816f $X=1.03 $Y=0.955 $X2=-0.19
+ $Y2=-0.245
cc_547 N_A_28_47#_c_955_n N_VGND_M1016_d 0.00329816f $X=1.89 $Y=0.955 $X2=0
+ $Y2=0
cc_548 N_A_28_47#_c_949_n N_VGND_c_991_n 0.0170777f $X=1.03 $Y=0.955 $X2=0 $Y2=0
cc_549 N_A_28_47#_c_955_n N_VGND_c_992_n 0.0170777f $X=1.89 $Y=0.955 $X2=0 $Y2=0
cc_550 N_A_28_47#_c_977_p N_VGND_c_997_n 0.0125234f $X=1.985 $Y=0.595 $X2=0
+ $Y2=0
cc_551 N_A_28_47#_c_948_n N_VGND_c_997_n 0.10384f $X=3.705 $Y=0.43 $X2=0 $Y2=0
cc_552 N_A_28_47#_c_946_n N_VGND_c_1001_n 0.0178111f $X=0.265 $Y=0.42 $X2=0
+ $Y2=0
cc_553 N_A_28_47#_c_980_p N_VGND_c_1002_n 0.0124525f $X=1.125 $Y=0.42 $X2=0
+ $Y2=0
cc_554 N_A_28_47#_M1002_s N_VGND_c_1004_n 0.00371702f $X=0.14 $Y=0.235 $X2=0
+ $Y2=0
cc_555 N_A_28_47#_M1013_s N_VGND_c_1004_n 0.00536646f $X=0.985 $Y=0.235 $X2=0
+ $Y2=0
cc_556 N_A_28_47#_M1025_s N_VGND_c_1004_n 0.00376627f $X=1.845 $Y=0.235 $X2=0
+ $Y2=0
cc_557 N_A_28_47#_M1023_s N_VGND_c_1004_n 0.00223577f $X=2.705 $Y=0.235 $X2=0
+ $Y2=0
cc_558 N_A_28_47#_M1038_s N_VGND_c_1004_n 0.00215176f $X=3.565 $Y=0.235 $X2=0
+ $Y2=0
cc_559 N_A_28_47#_c_946_n N_VGND_c_1004_n 0.0100304f $X=0.265 $Y=0.42 $X2=0
+ $Y2=0
cc_560 N_A_28_47#_c_980_p N_VGND_c_1004_n 0.00730901f $X=1.125 $Y=0.42 $X2=0
+ $Y2=0
cc_561 N_A_28_47#_c_977_p N_VGND_c_1004_n 0.00738676f $X=1.985 $Y=0.595 $X2=0
+ $Y2=0
cc_562 N_A_28_47#_c_948_n N_VGND_c_1004_n 0.0653197f $X=3.705 $Y=0.43 $X2=0
+ $Y2=0
cc_563 N_A_28_47#_c_948_n N_A_840_47#_c_1110_n 0.0211385f $X=3.705 $Y=0.43 $X2=0
+ $Y2=0
cc_564 N_VGND_c_1004_n N_A_840_47#_M1005_s 0.00215439f $X=10.32 $Y=0 $X2=-0.19
+ $Y2=-0.245
cc_565 N_VGND_c_1004_n N_A_840_47#_M1014_s 0.00223855f $X=10.32 $Y=0 $X2=0 $Y2=0
cc_566 N_VGND_c_1004_n N_A_840_47#_M1037_s 0.00223855f $X=10.32 $Y=0 $X2=0 $Y2=0
cc_567 N_VGND_c_1004_n N_A_840_47#_M1028_d 0.00223855f $X=10.32 $Y=0 $X2=0 $Y2=0
cc_568 N_VGND_c_1004_n N_A_840_47#_M1035_d 0.00215439f $X=10.32 $Y=0 $X2=0 $Y2=0
cc_569 N_VGND_c_993_n N_A_840_47#_c_1110_n 0.0268188f $X=8.285 $Y=0.465 $X2=0
+ $Y2=0
cc_570 N_VGND_c_997_n N_A_840_47#_c_1110_n 0.206111f $X=8.12 $Y=0 $X2=0 $Y2=0
cc_571 N_VGND_c_1004_n N_A_840_47#_c_1110_n 0.136992f $X=10.32 $Y=0 $X2=0 $Y2=0
cc_572 N_VGND_c_1004_n N_A_1267_47#_M1009_s 0.00225465f $X=10.32 $Y=0 $X2=-0.19
+ $Y2=-0.245
cc_573 N_VGND_c_1004_n N_A_1267_47#_M1030_s 0.00225465f $X=10.32 $Y=0 $X2=0
+ $Y2=0
cc_574 N_VGND_c_1004_n N_A_1267_47#_M1008_s 0.00273727f $X=10.32 $Y=0 $X2=0
+ $Y2=0
cc_575 N_VGND_c_1004_n N_A_1267_47#_M1031_s 0.00406837f $X=10.32 $Y=0 $X2=0
+ $Y2=0
cc_576 N_VGND_M1008_d N_A_1267_47#_c_1143_n 0.00651576f $X=8.16 $Y=0.235 $X2=0
+ $Y2=0
cc_577 N_VGND_c_993_n N_A_1267_47#_c_1143_n 0.0220556f $X=8.285 $Y=0.465 $X2=0
+ $Y2=0
cc_578 N_VGND_c_1004_n N_A_1267_47#_c_1143_n 0.016802f $X=10.32 $Y=0 $X2=0 $Y2=0
cc_579 N_VGND_c_999_n N_A_1267_47#_c_1170_n 0.0124525f $X=8.98 $Y=0 $X2=0 $Y2=0
cc_580 N_VGND_c_1004_n N_A_1267_47#_c_1170_n 0.00730901f $X=10.32 $Y=0 $X2=0
+ $Y2=0
cc_581 N_VGND_M1011_d N_A_1267_47#_c_1154_n 0.00350298f $X=9.005 $Y=0.235 $X2=0
+ $Y2=0
cc_582 N_VGND_c_994_n N_A_1267_47#_c_1154_n 0.0136397f $X=9.145 $Y=0.465 $X2=0
+ $Y2=0
cc_583 N_VGND_c_1004_n N_A_1267_47#_c_1154_n 0.0116172f $X=10.32 $Y=0 $X2=0
+ $Y2=0
cc_584 N_VGND_c_995_n N_A_1267_47#_c_1175_n 0.0124525f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_585 N_VGND_c_1004_n N_A_1267_47#_c_1175_n 0.00730901f $X=10.32 $Y=0 $X2=0
+ $Y2=0
cc_586 N_A_840_47#_c_1110_n N_A_1267_47#_M1009_s 0.00333618f $X=7.765 $Y=0.43
+ $X2=-0.19 $Y2=-0.245
cc_587 N_A_840_47#_c_1110_n N_A_1267_47#_M1030_s 0.00333618f $X=7.765 $Y=0.43
+ $X2=0 $Y2=0
cc_588 N_A_840_47#_M1028_d N_A_1267_47#_c_1143_n 0.00331529f $X=6.765 $Y=0.235
+ $X2=0 $Y2=0
cc_589 N_A_840_47#_M1035_d N_A_1267_47#_c_1143_n 0.00520331f $X=7.625 $Y=0.235
+ $X2=0 $Y2=0
cc_590 N_A_840_47#_c_1110_n N_A_1267_47#_c_1143_n 0.0909995f $X=7.765 $Y=0.43
+ $X2=0 $Y2=0
