* File: sky130_fd_sc_lp__or4bb_2.spice
* Created: Wed Sep  2 10:33:12 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__or4bb_2.pex.spice"
.subckt sky130_fd_sc_lp__or4bb_2  VNB VPB C_N A B D_N VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* D_N	D_N
* B	B
* A	A
* C_N	C_N
* VPB	VPB
* VNB	VNB
MM1003 N_VGND_M1003_d N_C_N_M1003_g N_A_40_47#_M1003_s VNB NSHORT L=0.15 W=0.42
+ AD=0.12915 AS=0.1113 PD=1.035 PS=1.37 NRD=95.712 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75003.4 A=0.063 P=1.14 MULT=1
MM1000 N_A_276_47#_M1000_d N_A_M1000_g N_VGND_M1003_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.12915 PD=0.7 PS=1.035 NRD=0 NRS=0 M=1 R=2.8 SA=75001 SB=75002.6
+ A=0.063 P=1.14 MULT=1
MM1006 N_VGND_M1006_d N_B_M1006_g N_A_276_47#_M1000_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1108 AS=0.0588 PD=0.96 PS=0.7 NRD=24.276 NRS=0 M=1 R=2.8 SA=75001.4
+ SB=75002.2 A=0.063 P=1.14 MULT=1
MM1010 N_A_276_47#_M1010_d N_A_40_47#_M1010_g N_VGND_M1006_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0588 AS=0.1108 PD=0.7 PS=0.96 NRD=0 NRS=41.424 M=1 R=2.8 SA=75002
+ SB=75001.6 A=0.063 P=1.14 MULT=1
MM1001 N_VGND_M1001_d N_A_462_351#_M1001_g N_A_276_47#_M1010_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0882 AS=0.0588 PD=0.803333 PS=0.7 NRD=24.276 NRS=0 M=1 R=2.8
+ SA=75002.5 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1008 N_VGND_M1001_d N_A_276_47#_M1008_g N_X_M1008_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1764 AS=0.1176 PD=1.60667 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.6
+ SB=75000.9 A=0.126 P=1.98 MULT=1
MM1014 N_VGND_M1014_d N_A_276_47#_M1014_g N_X_M1008_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1792 AS=0.1176 PD=1.62 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002 SB=75000.5
+ A=0.126 P=1.98 MULT=1
MM1009 N_A_462_351#_M1009_d N_D_N_M1009_g N_VGND_M1014_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1113 AS=0.0896 PD=1.37 PS=0.81 NRD=0 NRS=28.56 M=1 R=2.8
+ SA=75001.1 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1007 N_VPWR_M1007_d N_C_N_M1007_g N_A_40_47#_M1007_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75001.7
+ A=0.063 P=1.14 MULT=1
MM1002 A_276_403# N_A_M1002_g N_VPWR_M1007_d VPB PHIGHVT L=0.15 W=0.42 AD=0.0441
+ AS=0.0588 PD=0.63 PS=0.7 NRD=23.443 NRS=0 M=1 R=2.8 SA=75000.6 SB=75001.3
+ A=0.063 P=1.14 MULT=1
MM1004 A_348_403# N_B_M1004_g A_276_403# VPB PHIGHVT L=0.15 W=0.42 AD=0.0441
+ AS=0.0441 PD=0.63 PS=0.63 NRD=23.443 NRS=23.443 M=1 R=2.8 SA=75001 SB=75000.9
+ A=0.063 P=1.14 MULT=1
MM1012 A_420_403# N_A_40_47#_M1012_g A_348_403# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0441 AS=0.0441 PD=0.63 PS=0.63 NRD=23.443 NRS=23.443 M=1 R=2.8 SA=75001.3
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1015 N_A_276_47#_M1015_d N_A_462_351#_M1015_g A_420_403# VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1113 AS=0.0441 PD=1.37 PS=0.63 NRD=0 NRS=23.443 M=1 R=2.8
+ SA=75001.7 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1005 N_X_M1005_d N_A_276_47#_M1005_g N_VPWR_M1005_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75000.8 A=0.189 P=2.82 MULT=1
MM1013 N_X_M1005_d N_A_276_47#_M1013_g N_VPWR_M1013_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.285075 PD=1.54 PS=2.4525 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75000.4 A=0.189 P=2.82 MULT=1
MM1011 N_A_462_351#_M1011_d N_D_N_M1011_g N_VPWR_M1013_s VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1113 AS=0.095025 PD=1.37 PS=0.8175 NRD=0 NRS=80.3169 M=1 R=2.8
+ SA=75001.1 SB=75000.2 A=0.063 P=1.14 MULT=1
DX16_noxref VNB VPB NWDIODE A=9.6607 P=14.09
*
.include "sky130_fd_sc_lp__or4bb_2.pxi.spice"
*
.ends
*
*
