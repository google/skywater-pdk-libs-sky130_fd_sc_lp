* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__dlygate4s18_1 A VGND VNB VPB VPWR X
X0 VGND a_27_52# a_288_52# VNB sky130_fd_pr__nfet_01v8 w=420000u l=180000u
X1 a_405_136# a_288_52# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X2 VGND a_405_136# X VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X3 VPWR a_405_136# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X4 a_405_136# a_288_52# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=180000u
X5 a_27_52# A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 a_27_52# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X7 VPWR a_27_52# a_288_52# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
.ends
