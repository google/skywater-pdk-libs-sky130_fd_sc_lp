* File: sky130_fd_sc_lp__a2111oi_lp.pxi.spice
* Created: Fri Aug 28 09:47:04 2020
* 
x_PM_SKY130_FD_SC_LP__A2111OI_LP%A1 N_A1_M1006_g N_A1_M1008_g N_A1_c_89_n
+ N_A1_c_94_n A1 A1 N_A1_c_91_n PM_SKY130_FD_SC_LP__A2111OI_LP%A1
x_PM_SKY130_FD_SC_LP__A2111OI_LP%A2 N_A2_M1005_g N_A2_M1012_g A2 A2 N_A2_c_123_n
+ PM_SKY130_FD_SC_LP__A2111OI_LP%A2
x_PM_SKY130_FD_SC_LP__A2111OI_LP%B1 N_B1_c_160_n N_B1_M1000_g N_B1_c_161_n
+ N_B1_c_162_n N_B1_c_163_n N_B1_M1009_g N_B1_c_164_n N_B1_c_165_n N_B1_c_166_n
+ N_B1_c_170_n N_B1_M1004_g N_B1_c_167_n N_B1_c_171_n B1 B1 N_B1_c_169_n
+ PM_SKY130_FD_SC_LP__A2111OI_LP%B1
x_PM_SKY130_FD_SC_LP__A2111OI_LP%C1 N_C1_c_222_n N_C1_M1001_g N_C1_c_223_n
+ N_C1_c_224_n N_C1_M1007_g N_C1_c_225_n N_C1_M1010_g N_C1_c_226_n N_C1_c_227_n
+ N_C1_c_233_n N_C1_c_228_n C1 C1 C1 C1 C1 N_C1_c_230_n
+ PM_SKY130_FD_SC_LP__A2111OI_LP%C1
x_PM_SKY130_FD_SC_LP__A2111OI_LP%D1 N_D1_c_288_n N_D1_M1002_g N_D1_M1011_g
+ N_D1_c_289_n N_D1_M1003_g N_D1_c_290_n N_D1_c_291_n N_D1_c_292_n N_D1_c_297_n
+ D1 D1 N_D1_c_294_n PM_SKY130_FD_SC_LP__A2111OI_LP%D1
x_PM_SKY130_FD_SC_LP__A2111OI_LP%VPWR N_VPWR_M1006_s N_VPWR_M1012_d
+ N_VPWR_c_337_n N_VPWR_c_338_n N_VPWR_c_339_n N_VPWR_c_340_n VPWR
+ N_VPWR_c_341_n N_VPWR_c_336_n N_VPWR_c_343_n
+ PM_SKY130_FD_SC_LP__A2111OI_LP%VPWR
x_PM_SKY130_FD_SC_LP__A2111OI_LP%A_131_409# N_A_131_409#_M1006_d
+ N_A_131_409#_M1004_s N_A_131_409#_c_374_n N_A_131_409#_c_375_n
+ N_A_131_409#_c_376_n N_A_131_409#_c_377_n N_A_131_409#_c_378_n
+ PM_SKY130_FD_SC_LP__A2111OI_LP%A_131_409#
x_PM_SKY130_FD_SC_LP__A2111OI_LP%Y N_Y_M1008_s N_Y_M1009_d N_Y_M1010_d
+ N_Y_M1011_d N_Y_c_409_n N_Y_c_410_n N_Y_c_411_n N_Y_c_412_n N_Y_c_413_n
+ N_Y_c_414_n N_Y_c_418_n N_Y_c_415_n N_Y_c_416_n N_Y_c_419_n N_Y_c_417_n Y
+ N_Y_c_459_n PM_SKY130_FD_SC_LP__A2111OI_LP%Y
x_PM_SKY130_FD_SC_LP__A2111OI_LP%VGND N_VGND_M1005_d N_VGND_M1001_s
+ N_VGND_M1003_d N_VGND_c_498_n N_VGND_c_499_n N_VGND_c_500_n N_VGND_c_501_n
+ N_VGND_c_502_n N_VGND_c_503_n VGND N_VGND_c_504_n N_VGND_c_505_n
+ N_VGND_c_506_n N_VGND_c_507_n PM_SKY130_FD_SC_LP__A2111OI_LP%VGND
cc_1 VNB N_A1_M1008_g 0.0448828f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=0.495
cc_2 VNB N_A1_c_89_n 0.0231689f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=1.68
cc_3 VNB A1 0.0278758f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_4 VNB N_A1_c_91_n 0.0168566f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=1.34
cc_5 VNB N_A2_M1005_g 0.0358192f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=2.545
cc_6 VNB A2 0.00621905f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=1.68
cc_7 VNB N_A2_c_123_n 0.0523032f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_B1_c_160_n 0.0138901f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=1.845
cc_9 VNB N_B1_c_161_n 0.0102086f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_B1_c_162_n 0.00812973f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=1.175
cc_11 VNB N_B1_c_163_n 0.0171565f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=0.495
cc_12 VNB N_B1_c_164_n 0.0210019f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=1.175
cc_13 VNB N_B1_c_165_n 0.0512484f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=1.68
cc_14 VNB N_B1_c_166_n 0.00909426f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=1.845
cc_15 VNB N_B1_c_167_n 0.00664349f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB B1 0.00733255f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=1.34
cc_17 VNB N_B1_c_169_n 0.0260638f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=1.51
cc_18 VNB N_C1_c_222_n 0.0163717f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=1.845
cc_19 VNB N_C1_c_223_n 0.00960421f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_C1_c_224_n 0.0112613f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=1.175
cc_21 VNB N_C1_c_225_n 0.0135165f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=1.175
cc_22 VNB N_C1_c_226_n 0.022534f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_C1_c_227_n 0.0229706f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_C1_c_228_n 0.00437176f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB C1 0.00160428f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_C1_c_230_n 0.0167832f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_D1_c_288_n 0.0135266f $X=-0.19 $Y=-0.245 $X2=0.53 $Y2=1.845
cc_28 VNB N_D1_c_289_n 0.0177624f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=1.175
cc_29 VNB N_D1_c_290_n 0.0253496f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_D1_c_291_n 0.0184734f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_D1_c_292_n 0.0222717f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB D1 0.00459407f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=1.34
cc_33 VNB N_D1_c_294_n 0.0142188f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VPWR_c_336_n 0.183584f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_Y_c_409_n 0.0240181f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_36 VNB N_Y_c_410_n 0.0143904f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_Y_c_411_n 0.0101352f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_Y_c_412_n 0.00882835f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=1.34
cc_39 VNB N_Y_c_413_n 0.0190356f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=1.34
cc_40 VNB N_Y_c_414_n 0.0192522f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_Y_c_415_n 0.00394169f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_Y_c_416_n 0.00764113f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_Y_c_417_n 0.0315111f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_498_n 0.00177638f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=1.845
cc_45 VNB N_VGND_c_499_n 0.00693483f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_500_n 0.0105251f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_501_n 0.0197824f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_502_n 0.0276965f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=1.34
cc_49 VNB N_VGND_c_503_n 0.00513431f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.51
cc_50 VNB N_VGND_c_504_n 0.0299034f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_505_n 0.0337178f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_506_n 0.00500486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_507_n 0.24372f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VPB N_A1_M1006_g 0.0357919f $X=-0.19 $Y=1.655 $X2=0.53 $Y2=2.545
cc_55 VPB N_A1_c_89_n 0.00177087f $X=-0.19 $Y=1.655 $X2=0.49 $Y2=1.68
cc_56 VPB N_A1_c_94_n 0.0142253f $X=-0.19 $Y=1.655 $X2=0.49 $Y2=1.845
cc_57 VPB A1 0.0126484f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_58 VPB N_A2_M1012_g 0.0357919f $X=-0.19 $Y=1.655 $X2=0.55 $Y2=0.495
cc_59 VPB A2 0.00775354f $X=-0.19 $Y=1.655 $X2=0.49 $Y2=1.68
cc_60 VPB N_A2_c_123_n 0.0242554f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_61 VPB N_B1_c_170_n 0.0248365f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_62 VPB N_B1_c_171_n 0.0319413f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_63 VPB B1 0.00879768f $X=-0.19 $Y=1.655 $X2=0.49 $Y2=1.34
cc_64 VPB N_B1_c_169_n 0.00190131f $X=-0.19 $Y=1.655 $X2=0.49 $Y2=1.51
cc_65 VPB N_C1_M1007_g 0.0274235f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_66 VPB N_C1_c_227_n 0.00215581f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_67 VPB N_C1_c_233_n 0.0144827f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_68 VPB C1 0.00210243f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_69 VPB N_D1_M1011_g 0.0330709f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_70 VPB N_D1_c_292_n 0.00170229f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_71 VPB N_D1_c_297_n 0.0139582f $X=-0.19 $Y=1.655 $X2=0.49 $Y2=1.34
cc_72 VPB D1 0.00281229f $X=-0.19 $Y=1.655 $X2=0.49 $Y2=1.34
cc_73 VPB N_VPWR_c_337_n 0.0108784f $X=-0.19 $Y=1.655 $X2=0.55 $Y2=0.495
cc_74 VPB N_VPWR_c_338_n 0.0480962f $X=-0.19 $Y=1.655 $X2=0.49 $Y2=1.34
cc_75 VPB N_VPWR_c_339_n 0.0187052f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_76 VPB N_VPWR_c_340_n 0.0168378f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_77 VPB N_VPWR_c_341_n 0.0828343f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_78 VPB N_VPWR_c_336_n 0.10019f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_79 VPB N_VPWR_c_343_n 0.00548753f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_80 VPB N_A_131_409#_c_374_n 0.00374687f $X=-0.19 $Y=1.655 $X2=0.55 $Y2=0.495
cc_81 VPB N_A_131_409#_c_375_n 0.00207453f $X=-0.19 $Y=1.655 $X2=0.49 $Y2=1.34
cc_82 VPB N_A_131_409#_c_376_n 0.0414037f $X=-0.19 $Y=1.655 $X2=0.49 $Y2=1.68
cc_83 VPB N_A_131_409#_c_377_n 0.00234699f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_84 VPB N_A_131_409#_c_378_n 0.0212039f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_85 VPB N_Y_c_418_n 0.0390561f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=1.51
cc_86 VPB N_Y_c_419_n 0.0179524f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_87 VPB N_Y_c_417_n 0.0179785f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_88 N_A1_M1008_g N_A2_M1005_g 0.0542058f $X=0.55 $Y=0.495 $X2=0 $Y2=0
cc_89 N_A1_M1006_g N_A2_M1012_g 0.0171479f $X=0.53 $Y=2.545 $X2=0 $Y2=0
cc_90 A1 A2 0.0572071f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_91 N_A1_c_91_n A2 4.78066e-19 $X=0.49 $Y=1.34 $X2=0 $Y2=0
cc_92 A1 N_A2_c_123_n 0.00583555f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_93 N_A1_c_91_n N_A2_c_123_n 0.0424156f $X=0.49 $Y=1.34 $X2=0 $Y2=0
cc_94 N_A1_M1006_g N_VPWR_c_338_n 0.0236969f $X=0.53 $Y=2.545 $X2=0 $Y2=0
cc_95 N_A1_c_94_n N_VPWR_c_338_n 0.00213543f $X=0.49 $Y=1.845 $X2=0 $Y2=0
cc_96 A1 N_VPWR_c_338_n 0.0266157f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_97 N_A1_M1006_g N_VPWR_c_339_n 0.00769046f $X=0.53 $Y=2.545 $X2=0 $Y2=0
cc_98 N_A1_M1006_g N_VPWR_c_340_n 8.49223e-19 $X=0.53 $Y=2.545 $X2=0 $Y2=0
cc_99 N_A1_M1006_g N_VPWR_c_336_n 0.0134474f $X=0.53 $Y=2.545 $X2=0 $Y2=0
cc_100 N_A1_M1006_g N_A_131_409#_c_374_n 0.0036669f $X=0.53 $Y=2.545 $X2=0 $Y2=0
cc_101 A1 N_A_131_409#_c_374_n 0.0181148f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_102 N_A1_M1006_g N_A_131_409#_c_375_n 0.0156243f $X=0.53 $Y=2.545 $X2=0 $Y2=0
cc_103 N_A1_M1008_g N_Y_c_409_n 0.0130843f $X=0.55 $Y=0.495 $X2=0 $Y2=0
cc_104 N_A1_M1008_g N_Y_c_410_n 0.0082765f $X=0.55 $Y=0.495 $X2=0 $Y2=0
cc_105 A1 N_Y_c_410_n 0.0258094f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_106 N_A1_c_91_n N_Y_c_410_n 7.85225e-19 $X=0.49 $Y=1.34 $X2=0 $Y2=0
cc_107 N_A1_M1008_g N_Y_c_411_n 0.00420809f $X=0.55 $Y=0.495 $X2=0 $Y2=0
cc_108 A1 N_Y_c_411_n 0.0286122f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_109 N_A1_c_91_n N_Y_c_411_n 0.00403122f $X=0.49 $Y=1.34 $X2=0 $Y2=0
cc_110 N_A1_M1008_g N_VGND_c_498_n 0.0019059f $X=0.55 $Y=0.495 $X2=0 $Y2=0
cc_111 N_A1_M1008_g N_VGND_c_504_n 0.00502664f $X=0.55 $Y=0.495 $X2=0 $Y2=0
cc_112 N_A1_M1008_g N_VGND_c_507_n 0.00639278f $X=0.55 $Y=0.495 $X2=0 $Y2=0
cc_113 N_A2_M1005_g N_B1_c_160_n 0.0197172f $X=0.94 $Y=0.495 $X2=-0.19
+ $Y2=-0.245
cc_114 A2 N_B1_c_162_n 0.00208265f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_115 N_A2_c_123_n N_B1_c_162_n 0.00271936f $X=1.18 $Y=1.34 $X2=0 $Y2=0
cc_116 N_A2_M1005_g N_B1_c_164_n 0.00501416f $X=0.94 $Y=0.495 $X2=0 $Y2=0
cc_117 A2 N_B1_c_166_n 0.0118236f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_118 N_A2_c_123_n N_B1_c_166_n 0.00602469f $X=1.18 $Y=1.34 $X2=0 $Y2=0
cc_119 A2 B1 0.0464561f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_120 N_A2_c_123_n B1 0.00179847f $X=1.18 $Y=1.34 $X2=0 $Y2=0
cc_121 A2 N_B1_c_169_n 0.00253761f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_122 N_A2_M1012_g N_VPWR_c_338_n 9.45181e-19 $X=1.06 $Y=2.545 $X2=0 $Y2=0
cc_123 N_A2_M1012_g N_VPWR_c_339_n 0.00769046f $X=1.06 $Y=2.545 $X2=0 $Y2=0
cc_124 N_A2_M1012_g N_VPWR_c_340_n 0.0174419f $X=1.06 $Y=2.545 $X2=0 $Y2=0
cc_125 N_A2_M1012_g N_VPWR_c_336_n 0.0134474f $X=1.06 $Y=2.545 $X2=0 $Y2=0
cc_126 N_A2_M1012_g N_A_131_409#_c_374_n 0.00190741f $X=1.06 $Y=2.545 $X2=0
+ $Y2=0
cc_127 N_A2_c_123_n N_A_131_409#_c_374_n 0.00335061f $X=1.18 $Y=1.34 $X2=0 $Y2=0
cc_128 N_A2_M1012_g N_A_131_409#_c_375_n 0.0204671f $X=1.06 $Y=2.545 $X2=0 $Y2=0
cc_129 N_A2_M1012_g N_A_131_409#_c_376_n 0.0216154f $X=1.06 $Y=2.545 $X2=0 $Y2=0
cc_130 A2 N_A_131_409#_c_376_n 0.0607674f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_131 N_A2_c_123_n N_A_131_409#_c_376_n 0.00412558f $X=1.18 $Y=1.34 $X2=0 $Y2=0
cc_132 N_A2_M1005_g N_Y_c_409_n 0.0019649f $X=0.94 $Y=0.495 $X2=0 $Y2=0
cc_133 N_A2_M1005_g N_Y_c_410_n 0.0164432f $X=0.94 $Y=0.495 $X2=0 $Y2=0
cc_134 A2 N_Y_c_410_n 0.059118f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_135 N_A2_c_123_n N_Y_c_410_n 0.00760358f $X=1.18 $Y=1.34 $X2=0 $Y2=0
cc_136 A2 N_Y_c_415_n 0.00120514f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_137 N_A2_M1005_g N_VGND_c_498_n 0.0109044f $X=0.94 $Y=0.495 $X2=0 $Y2=0
cc_138 N_A2_M1005_g N_VGND_c_504_n 0.00445056f $X=0.94 $Y=0.495 $X2=0 $Y2=0
cc_139 N_A2_M1005_g N_VGND_c_507_n 0.0042789f $X=0.94 $Y=0.495 $X2=0 $Y2=0
cc_140 B1 N_C1_c_224_n 8.19797e-19 $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_141 N_B1_c_170_n N_C1_M1007_g 0.0360568f $X=2.57 $Y=1.97 $X2=0 $Y2=0
cc_142 N_B1_c_169_n N_C1_c_227_n 0.00731454f $X=2.43 $Y=1.34 $X2=0 $Y2=0
cc_143 N_B1_c_171_n N_C1_c_233_n 0.0433713f $X=2.43 $Y=1.68 $X2=0 $Y2=0
cc_144 N_B1_c_165_n C1 6.55083e-19 $X=2.265 $Y=1.25 $X2=0 $Y2=0
cc_145 N_B1_c_171_n C1 0.00467433f $X=2.43 $Y=1.68 $X2=0 $Y2=0
cc_146 B1 C1 0.0537598f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_147 N_B1_c_165_n N_C1_c_230_n 0.00731454f $X=2.265 $Y=1.25 $X2=0 $Y2=0
cc_148 B1 N_C1_c_230_n 0.00517248f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_149 N_B1_c_170_n N_VPWR_c_341_n 0.0086001f $X=2.57 $Y=1.97 $X2=0 $Y2=0
cc_150 N_B1_c_170_n N_VPWR_c_336_n 0.0166232f $X=2.57 $Y=1.97 $X2=0 $Y2=0
cc_151 B1 N_A_131_409#_c_376_n 0.00762737f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_152 N_B1_c_165_n N_A_131_409#_c_377_n 3.66268e-19 $X=2.265 $Y=1.25 $X2=0
+ $Y2=0
cc_153 N_B1_c_170_n N_A_131_409#_c_377_n 0.00400521f $X=2.57 $Y=1.97 $X2=0 $Y2=0
cc_154 N_B1_c_171_n N_A_131_409#_c_377_n 0.00480473f $X=2.43 $Y=1.68 $X2=0 $Y2=0
cc_155 B1 N_A_131_409#_c_377_n 0.0284747f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_156 N_B1_c_170_n N_A_131_409#_c_378_n 0.0168999f $X=2.57 $Y=1.97 $X2=0 $Y2=0
cc_157 N_B1_c_161_n N_Y_c_410_n 0.0100615f $X=1.655 $Y=0.855 $X2=0 $Y2=0
cc_158 N_B1_c_162_n N_Y_c_410_n 0.00769153f $X=1.445 $Y=0.855 $X2=0 $Y2=0
cc_159 N_B1_c_164_n N_Y_c_410_n 0.00373707f $X=1.73 $Y=1.175 $X2=0 $Y2=0
cc_160 N_B1_c_167_n N_Y_c_410_n 0.00407103f $X=1.73 $Y=0.855 $X2=0 $Y2=0
cc_161 N_B1_c_160_n N_Y_c_412_n 0.00170639f $X=1.37 $Y=0.78 $X2=0 $Y2=0
cc_162 N_B1_c_163_n N_Y_c_412_n 0.0110693f $X=1.73 $Y=0.78 $X2=0 $Y2=0
cc_163 N_B1_c_167_n N_Y_c_412_n 0.00296195f $X=1.73 $Y=0.855 $X2=0 $Y2=0
cc_164 N_B1_c_165_n N_Y_c_413_n 0.0114907f $X=2.265 $Y=1.25 $X2=0 $Y2=0
cc_165 B1 N_Y_c_413_n 0.0497312f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_166 N_B1_c_164_n N_Y_c_415_n 0.00238911f $X=1.73 $Y=1.175 $X2=0 $Y2=0
cc_167 N_B1_c_165_n N_Y_c_415_n 0.0110357f $X=2.265 $Y=1.25 $X2=0 $Y2=0
cc_168 N_B1_c_167_n N_Y_c_415_n 0.00286205f $X=1.73 $Y=0.855 $X2=0 $Y2=0
cc_169 B1 N_Y_c_415_n 0.00551823f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_170 N_B1_c_160_n N_VGND_c_498_n 0.0106307f $X=1.37 $Y=0.78 $X2=0 $Y2=0
cc_171 N_B1_c_163_n N_VGND_c_498_n 0.00189426f $X=1.73 $Y=0.78 $X2=0 $Y2=0
cc_172 N_B1_c_163_n N_VGND_c_499_n 0.00262237f $X=1.73 $Y=0.78 $X2=0 $Y2=0
cc_173 N_B1_c_160_n N_VGND_c_502_n 0.00445056f $X=1.37 $Y=0.78 $X2=0 $Y2=0
cc_174 N_B1_c_161_n N_VGND_c_502_n 4.57848e-19 $X=1.655 $Y=0.855 $X2=0 $Y2=0
cc_175 N_B1_c_163_n N_VGND_c_502_n 0.00502664f $X=1.73 $Y=0.78 $X2=0 $Y2=0
cc_176 N_B1_c_160_n N_VGND_c_507_n 0.0041956f $X=1.37 $Y=0.78 $X2=0 $Y2=0
cc_177 N_B1_c_161_n N_VGND_c_507_n 6.33118e-19 $X=1.655 $Y=0.855 $X2=0 $Y2=0
cc_178 N_B1_c_163_n N_VGND_c_507_n 0.00651958f $X=1.73 $Y=0.78 $X2=0 $Y2=0
cc_179 N_C1_c_225_n N_D1_c_288_n 0.0093481f $X=3.05 $Y=0.73 $X2=-0.19 $Y2=-0.245
cc_180 N_C1_M1007_g N_D1_M1011_g 0.0497549f $X=3.06 $Y=2.545 $X2=0 $Y2=0
cc_181 C1 N_D1_M1011_g 0.0118681f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_182 N_C1_c_228_n N_D1_c_290_n 0.0093481f $X=3.05 $Y=0.805 $X2=0 $Y2=0
cc_183 N_C1_c_226_n N_D1_c_291_n 0.0104505f $X=3.1 $Y=1.18 $X2=0 $Y2=0
cc_184 N_C1_c_227_n N_D1_c_292_n 0.0118393f $X=3.1 $Y=1.685 $X2=0 $Y2=0
cc_185 N_C1_c_233_n N_D1_c_297_n 0.0118393f $X=3.1 $Y=1.85 $X2=0 $Y2=0
cc_186 C1 D1 0.0435539f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_187 N_C1_c_230_n D1 0.00407139f $X=3.1 $Y=1.345 $X2=0 $Y2=0
cc_188 C1 N_D1_c_294_n 8.17099e-19 $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_189 N_C1_c_230_n N_D1_c_294_n 0.0118393f $X=3.1 $Y=1.345 $X2=0 $Y2=0
cc_190 N_C1_M1007_g N_VPWR_c_341_n 0.00596257f $X=3.06 $Y=2.545 $X2=0 $Y2=0
cc_191 C1 N_VPWR_c_341_n 0.00914393f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_192 N_C1_M1007_g N_VPWR_c_336_n 0.00771107f $X=3.06 $Y=2.545 $X2=0 $Y2=0
cc_193 C1 N_VPWR_c_336_n 0.0101955f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_194 N_C1_M1007_g N_A_131_409#_c_377_n 4.23425e-19 $X=3.06 $Y=2.545 $X2=0
+ $Y2=0
cc_195 C1 N_A_131_409#_c_377_n 0.00597643f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_196 N_C1_M1007_g N_A_131_409#_c_378_n 0.0024926f $X=3.06 $Y=2.545 $X2=0 $Y2=0
cc_197 C1 N_A_131_409#_c_378_n 0.0230193f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_198 C1 A_637_409# 0.0116484f $X=3.035 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_199 N_C1_c_222_n N_Y_c_412_n 0.00569354f $X=2.69 $Y=0.73 $X2=0 $Y2=0
cc_200 N_C1_c_223_n N_Y_c_413_n 0.00895817f $X=2.975 $Y=0.805 $X2=0 $Y2=0
cc_201 N_C1_c_224_n N_Y_c_413_n 0.00792219f $X=2.765 $Y=0.805 $X2=0 $Y2=0
cc_202 N_C1_c_226_n N_Y_c_413_n 0.00344427f $X=3.1 $Y=1.18 $X2=0 $Y2=0
cc_203 N_C1_c_228_n N_Y_c_413_n 8.36434e-19 $X=3.05 $Y=0.805 $X2=0 $Y2=0
cc_204 C1 N_Y_c_413_n 0.00502555f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_205 N_C1_M1007_g N_Y_c_418_n 7.44155e-19 $X=3.06 $Y=2.545 $X2=0 $Y2=0
cc_206 N_C1_c_226_n N_Y_c_416_n 0.00478475f $X=3.1 $Y=1.18 $X2=0 $Y2=0
cc_207 N_C1_c_228_n N_Y_c_416_n 0.00127563f $X=3.05 $Y=0.805 $X2=0 $Y2=0
cc_208 C1 N_Y_c_416_n 0.0211064f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_209 N_C1_c_230_n N_Y_c_416_n 0.00107634f $X=3.1 $Y=1.345 $X2=0 $Y2=0
cc_210 N_C1_M1007_g N_Y_c_419_n 7.35394e-19 $X=3.06 $Y=2.545 $X2=0 $Y2=0
cc_211 C1 N_Y_c_419_n 0.0315475f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_212 N_C1_c_222_n N_Y_c_459_n 0.00172293f $X=2.69 $Y=0.73 $X2=0 $Y2=0
cc_213 N_C1_c_225_n N_Y_c_459_n 0.0119213f $X=3.05 $Y=0.73 $X2=0 $Y2=0
cc_214 N_C1_c_228_n N_Y_c_459_n 0.00643468f $X=3.05 $Y=0.805 $X2=0 $Y2=0
cc_215 N_C1_c_222_n N_VGND_c_499_n 0.0125463f $X=2.69 $Y=0.73 $X2=0 $Y2=0
cc_216 N_C1_c_225_n N_VGND_c_499_n 0.00225836f $X=3.05 $Y=0.73 $X2=0 $Y2=0
cc_217 N_C1_c_222_n N_VGND_c_505_n 0.00486043f $X=2.69 $Y=0.73 $X2=0 $Y2=0
cc_218 N_C1_c_223_n N_VGND_c_505_n 4.87571e-19 $X=2.975 $Y=0.805 $X2=0 $Y2=0
cc_219 N_C1_c_225_n N_VGND_c_505_n 0.00406386f $X=3.05 $Y=0.73 $X2=0 $Y2=0
cc_220 N_C1_c_222_n N_VGND_c_507_n 0.00437711f $X=2.69 $Y=0.73 $X2=0 $Y2=0
cc_221 N_C1_c_223_n N_VGND_c_507_n 6.51792e-19 $X=2.975 $Y=0.805 $X2=0 $Y2=0
cc_222 N_C1_c_225_n N_VGND_c_507_n 0.00544533f $X=3.05 $Y=0.73 $X2=0 $Y2=0
cc_223 N_D1_M1011_g N_VPWR_c_341_n 0.0086001f $X=3.63 $Y=2.545 $X2=0 $Y2=0
cc_224 N_D1_M1011_g N_VPWR_c_336_n 0.0165732f $X=3.63 $Y=2.545 $X2=0 $Y2=0
cc_225 N_D1_c_290_n N_Y_c_414_n 0.0184565f $X=3.84 $Y=0.805 $X2=0 $Y2=0
cc_226 N_D1_c_291_n N_Y_c_414_n 0.00794702f $X=3.67 $Y=1.175 $X2=0 $Y2=0
cc_227 D1 N_Y_c_414_n 0.0261167f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_228 N_D1_c_294_n N_Y_c_414_n 5.73473e-19 $X=3.67 $Y=1.34 $X2=0 $Y2=0
cc_229 N_D1_M1011_g N_Y_c_418_n 0.01643f $X=3.63 $Y=2.545 $X2=0 $Y2=0
cc_230 N_D1_c_290_n N_Y_c_416_n 0.00119835f $X=3.84 $Y=0.805 $X2=0 $Y2=0
cc_231 N_D1_M1011_g N_Y_c_419_n 0.00506601f $X=3.63 $Y=2.545 $X2=0 $Y2=0
cc_232 N_D1_c_297_n N_Y_c_419_n 6.14058e-19 $X=3.67 $Y=1.845 $X2=0 $Y2=0
cc_233 D1 N_Y_c_419_n 0.00867382f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_234 N_D1_M1011_g N_Y_c_417_n 0.00590404f $X=3.63 $Y=2.545 $X2=0 $Y2=0
cc_235 N_D1_c_291_n N_Y_c_417_n 0.00500796f $X=3.67 $Y=1.175 $X2=0 $Y2=0
cc_236 D1 N_Y_c_417_n 0.0483772f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_237 N_D1_c_294_n N_Y_c_417_n 0.0148853f $X=3.67 $Y=1.34 $X2=0 $Y2=0
cc_238 N_D1_c_288_n N_Y_c_459_n 0.00873255f $X=3.48 $Y=0.73 $X2=0 $Y2=0
cc_239 N_D1_c_289_n N_Y_c_459_n 0.0014519f $X=3.84 $Y=0.73 $X2=0 $Y2=0
cc_240 N_D1_c_290_n N_Y_c_459_n 0.00566982f $X=3.84 $Y=0.805 $X2=0 $Y2=0
cc_241 N_D1_c_288_n N_VGND_c_501_n 0.00231629f $X=3.48 $Y=0.73 $X2=0 $Y2=0
cc_242 N_D1_c_289_n N_VGND_c_501_n 0.0132154f $X=3.84 $Y=0.73 $X2=0 $Y2=0
cc_243 N_D1_c_288_n N_VGND_c_505_n 0.00549284f $X=3.48 $Y=0.73 $X2=0 $Y2=0
cc_244 N_D1_c_289_n N_VGND_c_505_n 0.00486043f $X=3.84 $Y=0.73 $X2=0 $Y2=0
cc_245 N_D1_c_290_n N_VGND_c_505_n 5.32072e-19 $X=3.84 $Y=0.805 $X2=0 $Y2=0
cc_246 N_D1_c_288_n N_VGND_c_507_n 0.00612472f $X=3.48 $Y=0.73 $X2=0 $Y2=0
cc_247 N_D1_c_289_n N_VGND_c_507_n 0.00437711f $X=3.84 $Y=0.73 $X2=0 $Y2=0
cc_248 N_D1_c_290_n N_VGND_c_507_n 7.07256e-19 $X=3.84 $Y=0.805 $X2=0 $Y2=0
cc_249 N_VPWR_c_338_n N_A_131_409#_c_374_n 0.0119061f $X=0.265 $Y=2.19 $X2=0
+ $Y2=0
cc_250 N_VPWR_c_338_n N_A_131_409#_c_375_n 0.0572919f $X=0.265 $Y=2.19 $X2=0
+ $Y2=0
cc_251 N_VPWR_c_339_n N_A_131_409#_c_375_n 0.021949f $X=1.16 $Y=3.33 $X2=0 $Y2=0
cc_252 N_VPWR_c_340_n N_A_131_409#_c_375_n 0.0454646f $X=1.325 $Y=2.54 $X2=0
+ $Y2=0
cc_253 N_VPWR_c_336_n N_A_131_409#_c_375_n 0.0124703f $X=4.08 $Y=3.33 $X2=0
+ $Y2=0
cc_254 N_VPWR_M1012_d N_A_131_409#_c_376_n 0.00334849f $X=1.185 $Y=2.045 $X2=0
+ $Y2=0
cc_255 N_VPWR_c_340_n N_A_131_409#_c_376_n 0.02102f $X=1.325 $Y=2.54 $X2=0 $Y2=0
cc_256 N_VPWR_c_340_n N_A_131_409#_c_378_n 0.0225453f $X=1.325 $Y=2.54 $X2=0
+ $Y2=0
cc_257 N_VPWR_c_341_n N_A_131_409#_c_378_n 0.0220321f $X=4.08 $Y=3.33 $X2=0
+ $Y2=0
cc_258 N_VPWR_c_336_n N_A_131_409#_c_378_n 0.0125808f $X=4.08 $Y=3.33 $X2=0
+ $Y2=0
cc_259 N_VPWR_c_341_n N_Y_c_418_n 0.0304602f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_260 N_VPWR_c_336_n N_Y_c_418_n 0.0174175f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_261 N_Y_c_409_n N_VGND_c_498_n 0.0120387f $X=0.335 $Y=0.495 $X2=0 $Y2=0
cc_262 N_Y_c_410_n N_VGND_c_498_n 0.0200008f $X=1.78 $Y=0.91 $X2=0 $Y2=0
cc_263 N_Y_c_412_n N_VGND_c_498_n 0.0127138f $X=1.945 $Y=0.495 $X2=0 $Y2=0
cc_264 N_Y_c_412_n N_VGND_c_499_n 0.0282303f $X=1.945 $Y=0.495 $X2=0 $Y2=0
cc_265 N_Y_c_413_n N_VGND_c_499_n 0.0227455f $X=3.005 $Y=0.91 $X2=0 $Y2=0
cc_266 N_Y_c_459_n N_VGND_c_499_n 0.0157411f $X=3.265 $Y=0.47 $X2=0 $Y2=0
cc_267 N_Y_c_414_n N_VGND_c_501_n 0.0214493f $X=4.015 $Y=0.91 $X2=0 $Y2=0
cc_268 N_Y_c_459_n N_VGND_c_501_n 0.0129647f $X=3.265 $Y=0.47 $X2=0 $Y2=0
cc_269 N_Y_c_412_n N_VGND_c_502_n 0.0220321f $X=1.945 $Y=0.495 $X2=0 $Y2=0
cc_270 N_Y_c_409_n N_VGND_c_504_n 0.0220321f $X=0.335 $Y=0.495 $X2=0 $Y2=0
cc_271 N_Y_c_459_n N_VGND_c_505_n 0.0239324f $X=3.265 $Y=0.47 $X2=0 $Y2=0
cc_272 N_Y_M1010_d N_VGND_c_507_n 0.0022543f $X=3.125 $Y=0.235 $X2=0 $Y2=0
cc_273 N_Y_c_409_n N_VGND_c_507_n 0.0125808f $X=0.335 $Y=0.495 $X2=0 $Y2=0
cc_274 N_Y_c_410_n N_VGND_c_507_n 0.0300466f $X=1.78 $Y=0.91 $X2=0 $Y2=0
cc_275 N_Y_c_412_n N_VGND_c_507_n 0.0125808f $X=1.945 $Y=0.495 $X2=0 $Y2=0
cc_276 N_Y_c_413_n N_VGND_c_507_n 0.0190593f $X=3.005 $Y=0.91 $X2=0 $Y2=0
cc_277 N_Y_c_414_n N_VGND_c_507_n 0.0146689f $X=4.015 $Y=0.91 $X2=0 $Y2=0
cc_278 N_Y_c_459_n N_VGND_c_507_n 0.0157085f $X=3.265 $Y=0.47 $X2=0 $Y2=0
cc_279 N_VGND_c_507_n A_553_47# 0.00303453f $X=4.08 $Y=0 $X2=-0.19 $Y2=-0.245
cc_280 N_VGND_c_507_n A_711_47# 0.00303453f $X=4.08 $Y=0 $X2=-0.19 $Y2=-0.245
