* File: sky130_fd_sc_lp__bushold_1.pxi.spice
* Created: Wed Sep  2 09:37:34 2020
* 
x_PM_SKY130_FD_SC_LP__BUSHOLD_1%X N_X_M1003_d N_X_M1001_d N_X_M1005_g
+ N_X_M1002_g N_X_c_56_n N_X_c_57_n N_X_c_52_n N_X_c_53_n N_X_c_54_n N_X_c_60_n
+ N_X_c_61_n X X X X X X X N_X_c_64_n N_X_c_55_n PM_SKY130_FD_SC_LP__BUSHOLD_1%X
x_PM_SKY130_FD_SC_LP__BUSHOLD_1%RESET N_RESET_M1000_g N_RESET_M1004_g RESET
+ RESET RESET N_RESET_c_117_n N_RESET_c_118_n N_RESET_c_122_n
+ PM_SKY130_FD_SC_LP__BUSHOLD_1%RESET
x_PM_SKY130_FD_SC_LP__BUSHOLD_1%A_89_535# N_A_89_535#_M1005_d
+ N_A_89_535#_M1002_s N_A_89_535#_c_157_n N_A_89_535#_M1003_g
+ N_A_89_535#_c_166_n N_A_89_535#_M1001_g N_A_89_535#_c_158_n
+ N_A_89_535#_c_159_n N_A_89_535#_c_160_n N_A_89_535#_c_161_n
+ N_A_89_535#_c_162_n N_A_89_535#_c_163_n N_A_89_535#_c_184_n
+ N_A_89_535#_c_164_n N_A_89_535#_c_169_n N_A_89_535#_c_165_n
+ PM_SKY130_FD_SC_LP__BUSHOLD_1%A_89_535#
x_PM_SKY130_FD_SC_LP__BUSHOLD_1%VPWR N_VPWR_M1004_d N_VPWR_c_231_n VPWR
+ N_VPWR_c_232_n N_VPWR_c_233_n N_VPWR_c_230_n N_VPWR_c_235_n VPWR
+ PM_SKY130_FD_SC_LP__BUSHOLD_1%VPWR
x_PM_SKY130_FD_SC_LP__BUSHOLD_1%VGND N_VGND_M1005_s N_VGND_M1000_d
+ N_VGND_c_256_n N_VGND_c_257_n N_VGND_c_258_n N_VGND_c_259_n N_VGND_c_260_n
+ N_VGND_c_261_n VGND N_VGND_c_262_n N_VGND_c_263_n VGND
+ PM_SKY130_FD_SC_LP__BUSHOLD_1%VGND
cc_1 VNB N_X_M1005_g 0.0457531f $X=-0.19 $Y=-0.245 $X2=0.715 $Y2=0.445
cc_2 VNB N_X_c_52_n 0.00247473f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=1.35
cc_3 VNB N_X_c_53_n 0.0175853f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=1.35
cc_4 VNB N_X_c_54_n 0.0230401f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=2.03
cc_5 VNB N_X_c_55_n 0.0688121f $X=-0.19 $Y=-0.245 $X2=2.14 $Y2=0.445
cc_6 VNB N_RESET_M1000_g 0.0364367f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB RESET 0.00235741f $X=-0.19 $Y=-0.245 $X2=0.74 $Y2=2.195
cc_8 VNB N_RESET_c_117_n 0.0163407f $X=-0.19 $Y=-0.245 $X2=0.762 $Y2=2.555
cc_9 VNB N_RESET_c_118_n 0.020747f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=1.35
cc_10 VNB N_A_89_535#_c_157_n 0.0364793f $X=-0.19 $Y=-0.245 $X2=0.715 $Y2=1.185
cc_11 VNB N_A_89_535#_c_158_n 0.0262454f $X=-0.19 $Y=-0.245 $X2=0.785 $Y2=2.885
cc_12 VNB N_A_89_535#_c_159_n 0.0352638f $X=-0.19 $Y=-0.245 $X2=0.762 $Y2=2.405
cc_13 VNB N_A_89_535#_c_160_n 0.0113319f $X=-0.19 $Y=-0.245 $X2=0.762 $Y2=2.555
cc_14 VNB N_A_89_535#_c_161_n 0.0156584f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=2.365
cc_15 VNB N_A_89_535#_c_162_n 0.00110238f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=1.35
cc_16 VNB N_A_89_535#_c_163_n 0.00877659f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=2.03
cc_17 VNB N_A_89_535#_c_164_n 0.0598669f $X=-0.19 $Y=-0.245 $X2=2.075 $Y2=0.47
cc_18 VNB N_A_89_535#_c_165_n 0.00895372f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_VPWR_c_230_n 0.103974f $X=-0.19 $Y=-0.245 $X2=0.762 $Y2=2.405
cc_20 VNB N_VGND_c_256_n 0.0167439f $X=-0.19 $Y=-0.245 $X2=0.715 $Y2=0.445
cc_21 VNB N_VGND_c_257_n 0.0020563f $X=-0.19 $Y=-0.245 $X2=0.785 $Y2=2.555
cc_22 VNB N_VGND_c_258_n 0.0118587f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=1.35
cc_23 VNB N_VGND_c_259_n 0.00554993f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=1.185
cc_24 VNB N_VGND_c_260_n 0.0153073f $X=-0.19 $Y=-0.245 $X2=0.762 $Y2=2.555
cc_25 VNB N_VGND_c_261_n 0.00452904f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=2.365
cc_26 VNB N_VGND_c_262_n 0.0249832f $X=-0.19 $Y=-0.245 $X2=2.075 $Y2=0.84
cc_27 VNB N_VGND_c_263_n 0.150307f $X=-0.19 $Y=-0.245 $X2=2.075 $Y2=1.21
cc_28 VPB N_X_c_56_n 0.0127944f $X=-0.19 $Y=1.655 $X2=0.762 $Y2=2.405
cc_29 VPB N_X_c_57_n 0.0313627f $X=-0.19 $Y=1.655 $X2=0.762 $Y2=2.555
cc_30 VPB N_X_c_52_n 0.00157041f $X=-0.19 $Y=1.655 $X2=0.65 $Y2=1.35
cc_31 VPB N_X_c_54_n 0.0283454f $X=-0.19 $Y=1.655 $X2=0.65 $Y2=2.03
cc_32 VPB N_X_c_60_n 0.0227117f $X=-0.19 $Y=1.655 $X2=2.025 $Y2=2.45
cc_33 VPB N_X_c_61_n 0.00323215f $X=-0.19 $Y=1.655 $X2=0.815 $Y2=2.45
cc_34 VPB X 0.00777251f $X=-0.19 $Y=1.655 $X2=2.075 $Y2=2.32
cc_35 VPB X 0.0219272f $X=-0.19 $Y=1.655 $X2=2.075 $Y2=2.69
cc_36 VPB N_X_c_64_n 0.0176138f $X=-0.19 $Y=1.655 $X2=0.65 $Y2=2.195
cc_37 VPB N_X_c_55_n 0.0371619f $X=-0.19 $Y=1.655 $X2=2.14 $Y2=0.445
cc_38 VPB N_RESET_M1004_g 0.0336208f $X=-0.19 $Y=1.655 $X2=0.715 $Y2=1.185
cc_39 VPB RESET 0.00167151f $X=-0.19 $Y=1.655 $X2=0.74 $Y2=2.195
cc_40 VPB N_RESET_c_118_n 0.0255243f $X=-0.19 $Y=1.655 $X2=0.65 $Y2=1.35
cc_41 VPB N_RESET_c_122_n 0.0163407f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_42 VPB N_A_89_535#_c_166_n 0.0575103f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_43 VPB N_A_89_535#_c_159_n 0.0550794f $X=-0.19 $Y=1.655 $X2=0.762 $Y2=2.405
cc_44 VPB N_A_89_535#_c_164_n 0.0658598f $X=-0.19 $Y=1.655 $X2=2.075 $Y2=0.47
cc_45 VPB N_A_89_535#_c_169_n 0.0258866f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_46 VPB N_VPWR_c_231_n 4.89148e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_47 VPB N_VPWR_c_232_n 0.0333079f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_48 VPB N_VPWR_c_233_n 0.0263605f $X=-0.19 $Y=1.655 $X2=0.65 $Y2=1.185
cc_49 VPB N_VPWR_c_230_n 0.0465025f $X=-0.19 $Y=1.655 $X2=0.762 $Y2=2.405
cc_50 VPB N_VPWR_c_235_n 0.00436942f $X=-0.19 $Y=1.655 $X2=0.65 $Y2=1.35
cc_51 N_X_M1005_g N_RESET_M1000_g 0.031969f $X=0.715 $Y=0.445 $X2=0 $Y2=0
cc_52 N_X_c_56_n N_RESET_M1004_g 0.0102775f $X=0.762 $Y=2.405 $X2=0 $Y2=0
cc_53 N_X_c_57_n N_RESET_M1004_g 0.0511007f $X=0.762 $Y=2.555 $X2=0 $Y2=0
cc_54 N_X_c_52_n N_RESET_M1004_g 0.00107715f $X=0.65 $Y=1.35 $X2=0 $Y2=0
cc_55 N_X_c_60_n N_RESET_M1004_g 0.0112944f $X=2.025 $Y=2.45 $X2=0 $Y2=0
cc_56 N_X_c_52_n RESET 0.0674694f $X=0.65 $Y=1.35 $X2=0 $Y2=0
cc_57 N_X_c_53_n RESET 0.00351077f $X=0.65 $Y=1.35 $X2=0 $Y2=0
cc_58 N_X_c_60_n RESET 0.0256513f $X=2.025 $Y=2.45 $X2=0 $Y2=0
cc_59 N_X_c_52_n N_RESET_c_117_n 0.00351077f $X=0.65 $Y=1.35 $X2=0 $Y2=0
cc_60 N_X_c_53_n N_RESET_c_117_n 0.0204761f $X=0.65 $Y=1.35 $X2=0 $Y2=0
cc_61 N_X_c_54_n N_RESET_c_118_n 0.0204761f $X=0.65 $Y=2.03 $X2=0 $Y2=0
cc_62 N_X_c_60_n N_RESET_c_122_n 0.00123805f $X=2.025 $Y=2.45 $X2=0 $Y2=0
cc_63 N_X_c_64_n N_RESET_c_122_n 0.0204761f $X=0.65 $Y=2.195 $X2=0 $Y2=0
cc_64 N_X_c_55_n N_A_89_535#_c_157_n 0.0539579f $X=2.14 $Y=0.445 $X2=0 $Y2=0
cc_65 N_X_c_60_n N_A_89_535#_c_166_n 0.0225501f $X=2.025 $Y=2.45 $X2=0 $Y2=0
cc_66 X N_A_89_535#_c_166_n 0.00718359f $X=2.075 $Y=2.69 $X2=0 $Y2=0
cc_67 N_X_M1005_g N_A_89_535#_c_159_n 0.00534586f $X=0.715 $Y=0.445 $X2=0 $Y2=0
cc_68 N_X_c_56_n N_A_89_535#_c_159_n 0.00162067f $X=0.762 $Y=2.405 $X2=0 $Y2=0
cc_69 N_X_c_57_n N_A_89_535#_c_159_n 0.00480441f $X=0.762 $Y=2.555 $X2=0 $Y2=0
cc_70 N_X_c_52_n N_A_89_535#_c_159_n 0.0954087f $X=0.65 $Y=1.35 $X2=0 $Y2=0
cc_71 N_X_c_53_n N_A_89_535#_c_159_n 0.0227642f $X=0.65 $Y=1.35 $X2=0 $Y2=0
cc_72 N_X_c_61_n N_A_89_535#_c_159_n 0.0146597f $X=0.815 $Y=2.45 $X2=0 $Y2=0
cc_73 N_X_M1005_g N_A_89_535#_c_160_n 0.0179332f $X=0.715 $Y=0.445 $X2=0 $Y2=0
cc_74 N_X_c_52_n N_A_89_535#_c_160_n 0.0254879f $X=0.65 $Y=1.35 $X2=0 $Y2=0
cc_75 N_X_c_53_n N_A_89_535#_c_160_n 9.90912e-19 $X=0.65 $Y=1.35 $X2=0 $Y2=0
cc_76 N_X_M1005_g N_A_89_535#_c_162_n 0.00167927f $X=0.715 $Y=0.445 $X2=0 $Y2=0
cc_77 N_X_c_55_n N_A_89_535#_c_163_n 0.0207313f $X=2.14 $Y=0.445 $X2=0 $Y2=0
cc_78 N_X_c_60_n N_A_89_535#_c_184_n 0.0188915f $X=2.025 $Y=2.45 $X2=0 $Y2=0
cc_79 N_X_c_55_n N_A_89_535#_c_184_n 0.0943407f $X=2.14 $Y=0.445 $X2=0 $Y2=0
cc_80 N_X_c_60_n N_A_89_535#_c_164_n 0.0145178f $X=2.025 $Y=2.45 $X2=0 $Y2=0
cc_81 N_X_c_57_n N_A_89_535#_c_169_n 0.0058241f $X=0.762 $Y=2.555 $X2=0 $Y2=0
cc_82 N_X_c_61_n N_A_89_535#_c_169_n 0.0170817f $X=0.815 $Y=2.45 $X2=0 $Y2=0
cc_83 N_X_c_64_n N_A_89_535#_c_169_n 6.22595e-19 $X=0.65 $Y=2.195 $X2=0 $Y2=0
cc_84 N_X_c_52_n N_A_89_535#_c_165_n 0.00178367f $X=0.65 $Y=1.35 $X2=0 $Y2=0
cc_85 N_X_c_57_n N_VPWR_c_231_n 0.00225951f $X=0.762 $Y=2.555 $X2=0 $Y2=0
cc_86 N_X_c_60_n N_VPWR_c_231_n 0.0194922f $X=2.025 $Y=2.45 $X2=0 $Y2=0
cc_87 N_X_c_57_n N_VPWR_c_232_n 0.0054833f $X=0.762 $Y=2.555 $X2=0 $Y2=0
cc_88 X N_VPWR_c_233_n 0.0165867f $X=2.075 $Y=2.69 $X2=0 $Y2=0
cc_89 N_X_M1001_d N_VPWR_c_230_n 0.00230893f $X=2 $Y=2.675 $X2=0 $Y2=0
cc_90 N_X_c_57_n N_VPWR_c_230_n 0.00729566f $X=0.762 $Y=2.555 $X2=0 $Y2=0
cc_91 N_X_c_60_n N_VPWR_c_230_n 0.0281454f $X=2.025 $Y=2.45 $X2=0 $Y2=0
cc_92 N_X_c_61_n N_VPWR_c_230_n 0.00316817f $X=0.815 $Y=2.45 $X2=0 $Y2=0
cc_93 X N_VPWR_c_230_n 0.0110608f $X=2.075 $Y=2.69 $X2=0 $Y2=0
cc_94 N_X_M1005_g N_VGND_c_256_n 0.00340048f $X=0.715 $Y=0.445 $X2=0 $Y2=0
cc_95 N_X_M1005_g N_VGND_c_260_n 0.00436487f $X=0.715 $Y=0.445 $X2=0 $Y2=0
cc_96 N_X_c_55_n N_VGND_c_262_n 0.0192376f $X=2.14 $Y=0.445 $X2=0 $Y2=0
cc_97 N_X_M1003_d N_VGND_c_263_n 0.0030641f $X=2 $Y=0.235 $X2=0 $Y2=0
cc_98 N_X_M1005_g N_VGND_c_263_n 0.0070374f $X=0.715 $Y=0.445 $X2=0 $Y2=0
cc_99 N_X_c_55_n N_VGND_c_263_n 0.0111968f $X=2.14 $Y=0.445 $X2=0 $Y2=0
cc_100 N_RESET_M1000_g N_A_89_535#_c_157_n 0.0250761f $X=1.145 $Y=0.445 $X2=0
+ $Y2=0
cc_101 N_RESET_M1004_g N_A_89_535#_c_166_n 0.0210977f $X=1.145 $Y=2.885 $X2=0
+ $Y2=0
cc_102 N_RESET_M1000_g N_A_89_535#_c_162_n 0.00165727f $X=1.145 $Y=0.445 $X2=0
+ $Y2=0
cc_103 N_RESET_M1000_g N_A_89_535#_c_163_n 0.0151316f $X=1.145 $Y=0.445 $X2=0
+ $Y2=0
cc_104 RESET N_A_89_535#_c_163_n 0.0246206f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_105 N_RESET_c_117_n N_A_89_535#_c_163_n 9.28455e-19 $X=1.19 $Y=1.35 $X2=0
+ $Y2=0
cc_106 N_RESET_M1000_g N_A_89_535#_c_184_n 9.82596e-19 $X=1.145 $Y=0.445 $X2=0
+ $Y2=0
cc_107 RESET N_A_89_535#_c_184_n 0.0573914f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_108 N_RESET_c_117_n N_A_89_535#_c_184_n 0.00331304f $X=1.19 $Y=1.35 $X2=0
+ $Y2=0
cc_109 N_RESET_M1000_g N_A_89_535#_c_164_n 0.00797786f $X=1.145 $Y=0.445 $X2=0
+ $Y2=0
cc_110 N_RESET_M1004_g N_A_89_535#_c_164_n 0.00912501f $X=1.145 $Y=2.885 $X2=0
+ $Y2=0
cc_111 RESET N_A_89_535#_c_164_n 0.0042184f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_112 N_RESET_c_117_n N_A_89_535#_c_164_n 0.0632433f $X=1.19 $Y=1.35 $X2=0
+ $Y2=0
cc_113 N_RESET_M1004_g N_A_89_535#_c_169_n 8.89483e-19 $X=1.145 $Y=2.885 $X2=0
+ $Y2=0
cc_114 RESET N_A_89_535#_c_165_n 0.00272255f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_115 N_RESET_M1004_g N_VPWR_c_231_n 0.0113342f $X=1.145 $Y=2.885 $X2=0 $Y2=0
cc_116 N_RESET_M1004_g N_VPWR_c_232_n 0.00486043f $X=1.145 $Y=2.885 $X2=0 $Y2=0
cc_117 N_RESET_M1004_g N_VPWR_c_230_n 0.00435698f $X=1.145 $Y=2.885 $X2=0 $Y2=0
cc_118 N_RESET_M1000_g N_VGND_c_257_n 0.00167616f $X=1.145 $Y=0.445 $X2=0 $Y2=0
cc_119 N_RESET_M1000_g N_VGND_c_260_n 0.00436487f $X=1.145 $Y=0.445 $X2=0 $Y2=0
cc_120 N_RESET_M1000_g N_VGND_c_263_n 0.00594123f $X=1.145 $Y=0.445 $X2=0 $Y2=0
cc_121 N_A_89_535#_c_166_n N_VPWR_c_231_n 0.0157659f $X=1.75 $Y=2.655 $X2=0
+ $Y2=0
cc_122 N_A_89_535#_c_169_n N_VPWR_c_231_n 0.0115975f $X=0.57 $Y=2.885 $X2=0
+ $Y2=0
cc_123 N_A_89_535#_c_169_n N_VPWR_c_232_n 0.0359911f $X=0.57 $Y=2.885 $X2=0
+ $Y2=0
cc_124 N_A_89_535#_c_166_n N_VPWR_c_233_n 0.0185194f $X=1.75 $Y=2.655 $X2=0
+ $Y2=0
cc_125 N_A_89_535#_M1002_s N_VPWR_c_230_n 0.0021695f $X=0.445 $Y=2.675 $X2=0
+ $Y2=0
cc_126 N_A_89_535#_c_166_n N_VPWR_c_230_n 0.0165138f $X=1.75 $Y=2.655 $X2=0
+ $Y2=0
cc_127 N_A_89_535#_c_169_n N_VPWR_c_230_n 0.0243313f $X=0.57 $Y=2.885 $X2=0
+ $Y2=0
cc_128 N_A_89_535#_c_160_n N_VGND_c_256_n 0.0216778f $X=0.795 $Y=0.84 $X2=0
+ $Y2=0
cc_129 N_A_89_535#_c_157_n N_VGND_c_257_n 0.0131493f $X=1.75 $Y=0.725 $X2=0
+ $Y2=0
cc_130 N_A_89_535#_c_163_n N_VGND_c_257_n 0.0192551f $X=1.605 $Y=0.84 $X2=0
+ $Y2=0
cc_131 N_A_89_535#_c_160_n N_VGND_c_258_n 3.03177e-19 $X=0.795 $Y=0.84 $X2=0
+ $Y2=0
cc_132 N_A_89_535#_c_161_n N_VGND_c_258_n 0.00397886f $X=0.315 $Y=0.84 $X2=0
+ $Y2=0
cc_133 N_A_89_535#_c_160_n N_VGND_c_260_n 0.00240324f $X=0.795 $Y=0.84 $X2=0
+ $Y2=0
cc_134 N_A_89_535#_c_162_n N_VGND_c_260_n 0.0140722f $X=0.93 $Y=0.445 $X2=0
+ $Y2=0
cc_135 N_A_89_535#_c_163_n N_VGND_c_260_n 0.00240324f $X=1.605 $Y=0.84 $X2=0
+ $Y2=0
cc_136 N_A_89_535#_c_157_n N_VGND_c_262_n 0.0152513f $X=1.75 $Y=0.725 $X2=0
+ $Y2=0
cc_137 N_A_89_535#_c_163_n N_VGND_c_262_n 0.0048648f $X=1.605 $Y=0.84 $X2=0
+ $Y2=0
cc_138 N_A_89_535#_M1005_d N_VGND_c_263_n 0.00233323f $X=0.79 $Y=0.235 $X2=0
+ $Y2=0
cc_139 N_A_89_535#_c_157_n N_VGND_c_263_n 0.0204761f $X=1.75 $Y=0.725 $X2=0
+ $Y2=0
cc_140 N_A_89_535#_c_160_n N_VGND_c_263_n 0.00557564f $X=0.795 $Y=0.84 $X2=0
+ $Y2=0
cc_141 N_A_89_535#_c_161_n N_VGND_c_263_n 0.00657838f $X=0.315 $Y=0.84 $X2=0
+ $Y2=0
cc_142 N_A_89_535#_c_162_n N_VGND_c_263_n 0.00999079f $X=0.93 $Y=0.445 $X2=0
+ $Y2=0
cc_143 N_A_89_535#_c_163_n N_VGND_c_263_n 0.0126957f $X=1.605 $Y=0.84 $X2=0
+ $Y2=0
cc_144 A_172_535# N_VPWR_c_230_n 0.0029401f $X=0.86 $Y=2.675 $X2=2.16 $Y2=3.33
