* File: sky130_fd_sc_lp__dfrtn_1.pxi.spice
* Created: Wed Sep  2 09:43:34 2020
* 
x_PM_SKY130_FD_SC_LP__DFRTN_1%D N_D_M1020_g N_D_M1004_g D D D N_D_c_230_n
+ N_D_c_231_n PM_SKY130_FD_SC_LP__DFRTN_1%D
x_PM_SKY130_FD_SC_LP__DFRTN_1%A_294_35# N_A_294_35#_M1016_s N_A_294_35#_M1008_s
+ N_A_294_35#_M1001_g N_A_294_35#_M1002_g N_A_294_35#_M1003_g
+ N_A_294_35#_M1018_g N_A_294_35#_c_272_n N_A_294_35#_c_273_n
+ N_A_294_35#_c_274_n N_A_294_35#_c_275_n N_A_294_35#_c_291_n
+ N_A_294_35#_c_276_n N_A_294_35#_c_292_n N_A_294_35#_c_293_n
+ N_A_294_35#_c_306_p N_A_294_35#_c_277_n N_A_294_35#_c_367_p
+ N_A_294_35#_c_278_n N_A_294_35#_c_279_n N_A_294_35#_c_280_n
+ N_A_294_35#_c_281_n N_A_294_35#_c_282_n N_A_294_35#_c_356_p
+ N_A_294_35#_c_283_n N_A_294_35#_c_284_n N_A_294_35#_c_285_n
+ N_A_294_35#_c_286_n N_A_294_35#_c_287_n PM_SKY130_FD_SC_LP__DFRTN_1%A_294_35#
x_PM_SKY130_FD_SC_LP__DFRTN_1%A_501_229# N_A_501_229#_M1028_d
+ N_A_501_229#_M1017_d N_A_501_229#_M1006_g N_A_501_229#_M1015_g
+ N_A_501_229#_c_469_n N_A_501_229#_c_470_n N_A_501_229#_c_491_n
+ N_A_501_229#_c_471_n N_A_501_229#_c_472_n N_A_501_229#_c_473_n
+ N_A_501_229#_c_474_n N_A_501_229#_c_475_n N_A_501_229#_c_504_n
+ N_A_501_229#_c_476_n PM_SKY130_FD_SC_LP__DFRTN_1%A_501_229#
x_PM_SKY130_FD_SC_LP__DFRTN_1%RESET_B N_RESET_B_M1029_g N_RESET_B_c_588_n
+ N_RESET_B_c_589_n N_RESET_B_M1023_g N_RESET_B_M1031_g N_RESET_B_c_590_n
+ N_RESET_B_M1022_g N_RESET_B_c_592_n N_RESET_B_M1000_g N_RESET_B_M1019_g
+ N_RESET_B_c_594_n N_RESET_B_c_595_n N_RESET_B_c_596_n N_RESET_B_c_597_n
+ N_RESET_B_c_576_n N_RESET_B_c_577_n N_RESET_B_c_578_n N_RESET_B_c_579_n
+ N_RESET_B_c_580_n RESET_B N_RESET_B_c_581_n N_RESET_B_c_582_n
+ N_RESET_B_c_583_n N_RESET_B_c_584_n N_RESET_B_c_585_n N_RESET_B_c_586_n
+ N_RESET_B_c_608_n PM_SKY130_FD_SC_LP__DFRTN_1%RESET_B
x_PM_SKY130_FD_SC_LP__DFRTN_1%A_306_277# N_A_306_277#_M1025_s
+ N_A_306_277#_M1009_d N_A_306_277#_M1030_g N_A_306_277#_c_775_n
+ N_A_306_277#_c_776_n N_A_306_277#_c_777_n N_A_306_277#_M1011_g
+ N_A_306_277#_c_779_n N_A_306_277#_c_780_n N_A_306_277#_c_781_n
+ N_A_306_277#_c_782_n N_A_306_277#_c_783_n N_A_306_277#_c_784_n
+ N_A_306_277#_M1016_g N_A_306_277#_M1008_g N_A_306_277#_M1007_g
+ N_A_306_277#_c_787_n N_A_306_277#_c_788_n N_A_306_277#_M1005_g
+ N_A_306_277#_c_789_n N_A_306_277#_c_798_n N_A_306_277#_c_850_n
+ N_A_306_277#_c_799_n N_A_306_277#_c_800_n N_A_306_277#_c_801_n
+ N_A_306_277#_c_802_n N_A_306_277#_c_895_n N_A_306_277#_c_803_n
+ N_A_306_277#_c_804_n N_A_306_277#_c_805_n N_A_306_277#_c_790_n
+ N_A_306_277#_c_791_n N_A_306_277#_c_792_n N_A_306_277#_c_793_n
+ N_A_306_277#_c_807_n N_A_306_277#_c_851_n N_A_306_277#_c_808_n
+ N_A_306_277#_c_809_n N_A_306_277#_c_810_n N_A_306_277#_c_811_n
+ N_A_306_277#_c_794_n PM_SKY130_FD_SC_LP__DFRTN_1%A_306_277#
x_PM_SKY130_FD_SC_LP__DFRTN_1%A_336_463# N_A_336_463#_M1001_d
+ N_A_336_463#_M1030_d N_A_336_463#_M1022_d N_A_336_463#_M1017_g
+ N_A_336_463#_M1028_g N_A_336_463#_c_1048_n N_A_336_463#_c_1053_n
+ N_A_336_463#_c_1054_n N_A_336_463#_c_1049_n N_A_336_463#_c_1056_n
+ N_A_336_463#_c_1050_n PM_SKY130_FD_SC_LP__DFRTN_1%A_336_463#
x_PM_SKY130_FD_SC_LP__DFRTN_1%A_1287_276# N_A_1287_276#_M1014_d
+ N_A_1287_276#_M1000_d N_A_1287_276#_M1027_g N_A_1287_276#_M1013_g
+ N_A_1287_276#_c_1142_n N_A_1287_276#_c_1151_n N_A_1287_276#_c_1152_n
+ N_A_1287_276#_c_1143_n N_A_1287_276#_c_1144_n N_A_1287_276#_c_1145_n
+ N_A_1287_276#_c_1146_n N_A_1287_276#_c_1147_n N_A_1287_276#_c_1148_n
+ PM_SKY130_FD_SC_LP__DFRTN_1%A_1287_276#
x_PM_SKY130_FD_SC_LP__DFRTN_1%CLK_N N_CLK_N_M1009_g N_CLK_N_M1025_g CLK_N CLK_N
+ N_CLK_N_c_1237_n PM_SKY130_FD_SC_LP__DFRTN_1%CLK_N
x_PM_SKY130_FD_SC_LP__DFRTN_1%A_1099_447# N_A_1099_447#_M1007_d
+ N_A_1099_447#_M1003_d N_A_1099_447#_c_1273_n N_A_1099_447#_M1014_g
+ N_A_1099_447#_M1021_g N_A_1099_447#_c_1275_n N_A_1099_447#_c_1276_n
+ N_A_1099_447#_c_1277_n N_A_1099_447#_c_1278_n N_A_1099_447#_c_1279_n
+ N_A_1099_447#_M1024_g N_A_1099_447#_c_1281_n N_A_1099_447#_M1026_g
+ N_A_1099_447#_c_1282_n N_A_1099_447#_c_1283_n N_A_1099_447#_c_1294_n
+ N_A_1099_447#_c_1284_n N_A_1099_447#_c_1285_n N_A_1099_447#_c_1286_n
+ N_A_1099_447#_c_1287_n N_A_1099_447#_c_1288_n N_A_1099_447#_c_1289_n
+ N_A_1099_447#_c_1296_n N_A_1099_447#_c_1290_n N_A_1099_447#_c_1291_n
+ PM_SKY130_FD_SC_LP__DFRTN_1%A_1099_447#
x_PM_SKY130_FD_SC_LP__DFRTN_1%A_1832_367# N_A_1832_367#_M1026_s
+ N_A_1832_367#_M1024_s N_A_1832_367#_M1010_g N_A_1832_367#_M1012_g
+ N_A_1832_367#_c_1441_n N_A_1832_367#_c_1435_n N_A_1832_367#_c_1436_n
+ N_A_1832_367#_c_1437_n N_A_1832_367#_c_1438_n N_A_1832_367#_c_1439_n
+ PM_SKY130_FD_SC_LP__DFRTN_1%A_1832_367#
x_PM_SKY130_FD_SC_LP__DFRTN_1%A_27_463# N_A_27_463#_M1020_d N_A_27_463#_M1029_s
+ N_A_27_463#_M1004_d N_A_27_463#_c_1497_n N_A_27_463#_c_1500_n
+ N_A_27_463#_c_1498_n N_A_27_463#_c_1502_n N_A_27_463#_c_1495_n
+ N_A_27_463#_c_1496_n PM_SKY130_FD_SC_LP__DFRTN_1%A_27_463#
x_PM_SKY130_FD_SC_LP__DFRTN_1%VPWR N_VPWR_M1029_d N_VPWR_M1015_d N_VPWR_M1008_d
+ N_VPWR_M1027_d N_VPWR_M1021_d N_VPWR_M1024_d N_VPWR_c_1555_n N_VPWR_c_1556_n
+ N_VPWR_c_1557_n N_VPWR_c_1558_n N_VPWR_c_1559_n N_VPWR_c_1560_n
+ N_VPWR_c_1561_n N_VPWR_c_1562_n N_VPWR_c_1563_n N_VPWR_c_1564_n VPWR
+ N_VPWR_c_1565_n N_VPWR_c_1566_n N_VPWR_c_1567_n N_VPWR_c_1554_n
+ N_VPWR_c_1569_n N_VPWR_c_1570_n N_VPWR_c_1571_n N_VPWR_c_1572_n
+ PM_SKY130_FD_SC_LP__DFRTN_1%VPWR
x_PM_SKY130_FD_SC_LP__DFRTN_1%Q N_Q_M1010_d N_Q_M1012_d Q Q Q Q Q Q Q
+ N_Q_c_1672_n Q Q PM_SKY130_FD_SC_LP__DFRTN_1%Q
x_PM_SKY130_FD_SC_LP__DFRTN_1%VGND N_VGND_M1023_s N_VGND_M1031_d N_VGND_M1016_d
+ N_VGND_M1013_d N_VGND_M1025_d N_VGND_M1026_d N_VGND_c_1688_n N_VGND_c_1689_n
+ N_VGND_c_1690_n N_VGND_c_1691_n N_VGND_c_1692_n N_VGND_c_1693_n
+ N_VGND_c_1694_n N_VGND_c_1695_n N_VGND_c_1696_n N_VGND_c_1697_n VGND
+ N_VGND_c_1698_n N_VGND_c_1699_n N_VGND_c_1700_n N_VGND_c_1701_n
+ N_VGND_c_1702_n N_VGND_c_1703_n N_VGND_c_1704_n N_VGND_c_1705_n
+ PM_SKY130_FD_SC_LP__DFRTN_1%VGND
cc_1 VNB N_D_M1004_g 0.0101621f $X=-0.19 $Y=-0.245 $X2=1.135 $Y2=2.525
cc_2 VNB D 0.0365669f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.21
cc_3 VNB N_D_c_230_n 0.0360858f $X=-0.19 $Y=-0.245 $X2=1.085 $Y2=1.3
cc_4 VNB N_D_c_231_n 0.0330512f $X=-0.19 $Y=-0.245 $X2=1.085 $Y2=1.135
cc_5 VNB N_A_294_35#_c_272_n 0.0167117f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_6 VNB N_A_294_35#_c_273_n 0.0392774f $X=-0.19 $Y=-0.245 $X2=1.085 $Y2=1.272
cc_7 VNB N_A_294_35#_c_274_n 0.0012986f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_294_35#_c_275_n 0.00724134f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_294_35#_c_276_n 0.00287557f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_294_35#_c_277_n 0.00210846f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_294_35#_c_278_n 0.00300949f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_294_35#_c_279_n 3.25977e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_294_35#_c_280_n 0.00394787f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_294_35#_c_281_n 0.00546405f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_294_35#_c_282_n 0.0425609f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_294_35#_c_283_n 0.00537658f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_294_35#_c_284_n 0.0180618f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_294_35#_c_285_n 0.00105555f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_294_35#_c_286_n 0.0166117f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_294_35#_c_287_n 0.0194192f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_501_229#_M1015_g 0.0105936f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_501_229#_c_469_n 0.0220029f $X=-0.19 $Y=-0.245 $X2=1.085 $Y2=1.3
cc_23 VNB N_A_501_229#_c_470_n 0.00413668f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.272
cc_24 VNB N_A_501_229#_c_471_n 0.00246094f $X=-0.19 $Y=-0.245 $X2=1.085
+ $Y2=1.272
cc_25 VNB N_A_501_229#_c_472_n 0.0336265f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_501_229#_c_473_n 0.00310927f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_501_229#_c_474_n 0.00435986f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_501_229#_c_475_n 0.00601882f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_501_229#_c_476_n 0.0157661f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_RESET_B_M1023_g 0.0587756f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_31 VNB N_RESET_B_M1031_g 0.0410991f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_RESET_B_M1019_g 0.0413713f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_RESET_B_c_576_n 0.0124797f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_RESET_B_c_577_n 0.00595384f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_RESET_B_c_578_n 0.0152122f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_RESET_B_c_579_n 0.00185747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_RESET_B_c_580_n 0.00264232f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_RESET_B_c_581_n 0.0222559f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_RESET_B_c_582_n 0.00227299f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_RESET_B_c_583_n 0.0105881f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_RESET_B_c_584_n 9.36892e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_RESET_B_c_585_n 0.0203298f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_RESET_B_c_586_n 0.00545353f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_306_277#_M1030_g 0.00696784f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_45 VNB N_A_306_277#_c_775_n 0.021515f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_306_277#_c_776_n 0.00762295f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_306_277#_c_777_n 0.0311244f $X=-0.19 $Y=-0.245 $X2=1.085 $Y2=1.3
cc_48 VNB N_A_306_277#_M1011_g 0.0232017f $X=-0.19 $Y=-0.245 $X2=1.085 $Y2=1.3
cc_49 VNB N_A_306_277#_c_779_n 0.11834f $X=-0.19 $Y=-0.245 $X2=1.085 $Y2=1.135
cc_50 VNB N_A_306_277#_c_780_n 0.0109058f $X=-0.19 $Y=-0.245 $X2=1.085 $Y2=1.465
cc_51 VNB N_A_306_277#_c_781_n 0.0538793f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_306_277#_c_782_n 0.0209237f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_306_277#_c_783_n 0.0128814f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.272
cc_54 VNB N_A_306_277#_c_784_n 0.0171428f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_306_277#_M1008_g 0.0328709f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_306_277#_M1007_g 0.0212018f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_306_277#_c_787_n 0.0232443f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_306_277#_c_788_n 0.00914604f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_306_277#_c_789_n 0.00558121f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_306_277#_c_790_n 0.00279977f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_A_306_277#_c_791_n 0.00130001f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_A_306_277#_c_792_n 0.00318643f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_A_306_277#_c_793_n 0.00497498f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_A_306_277#_c_794_n 0.0223006f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_A_336_463#_M1017_g 0.00241418f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_A_336_463#_M1028_g 0.0313684f $X=-0.19 $Y=-0.245 $X2=1.085 $Y2=1.3
cc_67 VNB N_A_336_463#_c_1048_n 0.00397872f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_A_336_463#_c_1049_n 0.00239763f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_336_463#_c_1050_n 0.0500508f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_A_1287_276#_M1013_g 0.0313759f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_A_1287_276#_c_1142_n 0.00801725f $X=-0.19 $Y=-0.245 $X2=1.085
+ $Y2=1.135
cc_72 VNB N_A_1287_276#_c_1143_n 0.0189137f $X=-0.19 $Y=-0.245 $X2=0.72
+ $Y2=1.272
cc_73 VNB N_A_1287_276#_c_1144_n 0.0123131f $X=-0.19 $Y=-0.245 $X2=1.085
+ $Y2=1.272
cc_74 VNB N_A_1287_276#_c_1145_n 0.00208892f $X=-0.19 $Y=-0.245 $X2=1.2
+ $Y2=1.272
cc_75 VNB N_A_1287_276#_c_1146_n 0.00482322f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_A_1287_276#_c_1147_n 0.00489447f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_A_1287_276#_c_1148_n 0.00961292f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_CLK_N_M1025_g 0.0251982f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB CLK_N 0.0022984f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_CLK_N_c_1237_n 0.0201645f $X=-0.19 $Y=-0.245 $X2=1.085 $Y2=1.465
cc_81 VNB N_A_1099_447#_c_1273_n 0.0157172f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_A_1099_447#_M1021_g 0.0210557f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_A_1099_447#_c_1275_n 0.0383129f $X=-0.19 $Y=-0.245 $X2=1.085 $Y2=1.3
cc_84 VNB N_A_1099_447#_c_1276_n 0.0519558f $X=-0.19 $Y=-0.245 $X2=1.085 $Y2=1.3
cc_85 VNB N_A_1099_447#_c_1277_n 0.0140525f $X=-0.19 $Y=-0.245 $X2=0.24
+ $Y2=1.272
cc_86 VNB N_A_1099_447#_c_1278_n 0.0162768f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_A_1099_447#_c_1279_n 0.00970515f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_A_1099_447#_M1024_g 0.0464401f $X=-0.19 $Y=-0.245 $X2=1.085
+ $Y2=1.272
cc_89 VNB N_A_1099_447#_c_1281_n 0.0196242f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_A_1099_447#_c_1282_n 0.0340431f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_A_1099_447#_c_1283_n 0.00867771f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_A_1099_447#_c_1284_n 0.00169848f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_93 VNB N_A_1099_447#_c_1285_n 0.0111912f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_94 VNB N_A_1099_447#_c_1286_n 0.00688092f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_95 VNB N_A_1099_447#_c_1287_n 0.00117709f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_96 VNB N_A_1099_447#_c_1288_n 0.00386238f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_97 VNB N_A_1099_447#_c_1289_n 0.0148949f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_98 VNB N_A_1099_447#_c_1290_n 0.00111377f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_99 VNB N_A_1099_447#_c_1291_n 0.0408874f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_100 VNB N_A_1832_367#_M1010_g 0.0304293f $X=-0.19 $Y=-0.245 $X2=0.635
+ $Y2=1.21
cc_101 VNB N_A_1832_367#_c_1435_n 0.00504709f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_102 VNB N_A_1832_367#_c_1436_n 0.00481073f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_103 VNB N_A_1832_367#_c_1437_n 0.0291131f $X=-0.19 $Y=-0.245 $X2=1.085
+ $Y2=1.272
cc_104 VNB N_A_1832_367#_c_1438_n 0.00795841f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_105 VNB N_A_1832_367#_c_1439_n 0.00386788f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_106 VNB N_A_27_463#_c_1495_n 0.00590875f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_107 VNB N_A_27_463#_c_1496_n 0.00302902f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_108 VNB N_VPWR_c_1554_n 0.442315f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_109 VNB Q 0.00811041f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_110 VNB Q 0.0292897f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_111 VNB N_Q_c_1672_n 0.0266027f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=1.272
cc_112 VNB N_VGND_c_1688_n 0.0163414f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.272
cc_113 VNB N_VGND_c_1689_n 0.0344316f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_114 VNB N_VGND_c_1690_n 0.012902f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=1.272
cc_115 VNB N_VGND_c_1691_n 0.0168151f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_116 VNB N_VGND_c_1692_n 0.0227886f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_117 VNB N_VGND_c_1693_n 0.0102098f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_118 VNB N_VGND_c_1694_n 0.0700839f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_119 VNB N_VGND_c_1695_n 0.00436584f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_120 VNB N_VGND_c_1696_n 0.0424496f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_121 VNB N_VGND_c_1697_n 0.00326991f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_122 VNB N_VGND_c_1698_n 0.0231222f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_123 VNB N_VGND_c_1699_n 0.0487342f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_124 VNB N_VGND_c_1700_n 0.0218779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_125 VNB N_VGND_c_1701_n 0.0173182f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_126 VNB N_VGND_c_1702_n 0.559499f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_127 VNB N_VGND_c_1703_n 0.0151894f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_128 VNB N_VGND_c_1704_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_129 VNB N_VGND_c_1705_n 0.00499771f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_130 VPB N_D_M1004_g 0.0458461f $X=-0.19 $Y=1.655 $X2=1.135 $Y2=2.525
cc_131 VPB N_A_294_35#_M1002_g 0.0247889f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_132 VPB N_A_294_35#_M1003_g 0.0355946f $X=-0.19 $Y=1.655 $X2=1.085 $Y2=1.3
cc_133 VPB N_A_294_35#_c_275_n 7.414e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_134 VPB N_A_294_35#_c_291_n 0.03819f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_135 VPB N_A_294_35#_c_292_n 9.29659e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_136 VPB N_A_294_35#_c_293_n 0.0231463f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_137 VPB N_A_294_35#_c_283_n 0.00284159f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_138 VPB N_A_294_35#_c_284_n 0.0146096f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_139 VPB N_A_501_229#_M1015_g 0.0438862f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_140 VPB N_A_501_229#_c_470_n 0.00417494f $X=-0.19 $Y=1.655 $X2=0.24 $Y2=1.272
cc_141 VPB N_RESET_B_M1029_g 0.0413667f $X=-0.19 $Y=1.655 $X2=1.135 $Y2=1.465
cc_142 VPB N_RESET_B_c_588_n 0.205199f $X=-0.19 $Y=1.655 $X2=1.135 $Y2=2.525
cc_143 VPB N_RESET_B_c_589_n 0.012806f $X=-0.19 $Y=1.655 $X2=1.135 $Y2=2.525
cc_144 VPB N_RESET_B_c_590_n 0.0227958f $X=-0.19 $Y=1.655 $X2=1.085 $Y2=1.3
cc_145 VPB N_RESET_B_M1022_g 0.0285504f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_146 VPB N_RESET_B_c_592_n 0.0191808f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_147 VPB N_RESET_B_M1000_g 0.0398711f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_148 VPB N_RESET_B_c_594_n 0.0281128f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_149 VPB N_RESET_B_c_595_n 0.0193388f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_150 VPB N_RESET_B_c_596_n 0.02033f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_151 VPB N_RESET_B_c_597_n 0.0260617f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_152 VPB N_RESET_B_c_576_n 0.00988275f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_153 VPB N_RESET_B_c_577_n 0.00495812f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_154 VPB N_RESET_B_c_578_n 0.0248017f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_155 VPB N_RESET_B_c_579_n 0.00177885f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_156 VPB N_RESET_B_c_580_n 0.00180715f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_157 VPB N_RESET_B_c_582_n 0.0235066f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_158 VPB N_RESET_B_c_583_n 0.00650089f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_159 VPB N_RESET_B_c_584_n 0.00377849f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_160 VPB N_RESET_B_c_585_n 0.0143238f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_161 VPB N_RESET_B_c_586_n 0.00467533f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_162 VPB N_RESET_B_c_608_n 9.95493e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_163 VPB N_A_306_277#_M1030_g 0.0466189f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_164 VPB N_A_306_277#_M1008_g 0.0331871f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_165 VPB N_A_306_277#_M1005_g 0.0207044f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_166 VPB N_A_306_277#_c_798_n 0.00323482f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_167 VPB N_A_306_277#_c_799_n 0.0012114f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_168 VPB N_A_306_277#_c_800_n 0.0245299f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_169 VPB N_A_306_277#_c_801_n 6.22938e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_170 VPB N_A_306_277#_c_802_n 0.00708469f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_171 VPB N_A_306_277#_c_803_n 3.27367e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_172 VPB N_A_306_277#_c_804_n 0.00317221f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_173 VPB N_A_306_277#_c_805_n 2.92632e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_174 VPB N_A_306_277#_c_793_n 0.0158068f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_175 VPB N_A_306_277#_c_807_n 0.0035542f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_176 VPB N_A_306_277#_c_808_n 0.00106894f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_177 VPB N_A_306_277#_c_809_n 0.0419979f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_178 VPB N_A_306_277#_c_810_n 0.0255336f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_179 VPB N_A_306_277#_c_811_n 0.0500163f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_180 VPB N_A_306_277#_c_794_n 0.0281506f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_181 VPB N_A_336_463#_M1017_g 0.0447623f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_182 VPB N_A_336_463#_c_1048_n 0.00702505f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_183 VPB N_A_336_463#_c_1053_n 0.0169819f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=1.272
cc_184 VPB N_A_336_463#_c_1054_n 0.0133779f $X=-0.19 $Y=1.655 $X2=1.085
+ $Y2=1.272
cc_185 VPB N_A_336_463#_c_1049_n 0.00769549f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_186 VPB N_A_336_463#_c_1056_n 0.00834648f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_187 VPB N_A_1287_276#_M1027_g 0.0473476f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_188 VPB N_A_1287_276#_c_1142_n 0.0172228f $X=-0.19 $Y=1.655 $X2=1.085
+ $Y2=1.135
cc_189 VPB N_A_1287_276#_c_1151_n 0.0184793f $X=-0.19 $Y=1.655 $X2=1.085
+ $Y2=1.465
cc_190 VPB N_A_1287_276#_c_1152_n 2.47789e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_191 VPB N_A_1287_276#_c_1146_n 0.0146376f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_192 VPB N_CLK_N_M1009_g 0.028766f $X=-0.19 $Y=1.655 $X2=0.995 $Y2=0.815
cc_193 VPB CLK_N 0.00205079f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_194 VPB N_CLK_N_c_1237_n 0.0593405f $X=-0.19 $Y=1.655 $X2=1.085 $Y2=1.465
cc_195 VPB N_A_1099_447#_M1021_g 0.0530258f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_196 VPB N_A_1099_447#_M1024_g 0.0264879f $X=-0.19 $Y=1.655 $X2=1.085
+ $Y2=1.272
cc_197 VPB N_A_1099_447#_c_1294_n 0.00164671f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_198 VPB N_A_1099_447#_c_1285_n 0.00401141f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_199 VPB N_A_1099_447#_c_1296_n 0.0102246f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_200 VPB N_A_1832_367#_M1012_g 0.0257516f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_201 VPB N_A_1832_367#_c_1441_n 0.0148903f $X=-0.19 $Y=1.655 $X2=1.085
+ $Y2=1.135
cc_202 VPB N_A_1832_367#_c_1436_n 0.00281539f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_203 VPB N_A_1832_367#_c_1437_n 0.00785779f $X=-0.19 $Y=1.655 $X2=1.085
+ $Y2=1.272
cc_204 VPB N_A_1832_367#_c_1438_n 2.60844e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_205 VPB N_A_27_463#_c_1497_n 0.00858256f $X=-0.19 $Y=1.655 $X2=1.115 $Y2=1.21
cc_206 VPB N_A_27_463#_c_1498_n 0.0228957f $X=-0.19 $Y=1.655 $X2=1.085 $Y2=1.3
cc_207 VPB N_VPWR_c_1555_n 0.00928684f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_208 VPB N_VPWR_c_1556_n 0.0133721f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_209 VPB N_VPWR_c_1557_n 0.0368773f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_210 VPB N_VPWR_c_1558_n 0.00549813f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_211 VPB N_VPWR_c_1559_n 0.00610746f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_212 VPB N_VPWR_c_1560_n 0.0284125f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_213 VPB N_VPWR_c_1561_n 0.048229f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_214 VPB N_VPWR_c_1562_n 0.0038195f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_215 VPB N_VPWR_c_1563_n 0.0295512f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_216 VPB N_VPWR_c_1564_n 0.0036251f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_217 VPB N_VPWR_c_1565_n 0.0536192f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_218 VPB N_VPWR_c_1566_n 0.0364423f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_219 VPB N_VPWR_c_1567_n 0.0175526f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_220 VPB N_VPWR_c_1554_n 0.112094f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_221 VPB N_VPWR_c_1569_n 0.0240575f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_222 VPB N_VPWR_c_1570_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_223 VPB N_VPWR_c_1571_n 0.0122641f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_224 VPB N_VPWR_c_1572_n 0.00708764f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_225 VPB Q 0.0094786f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_226 VPB Q 0.0483872f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_227 N_D_c_231_n N_A_294_35#_c_272_n 0.00127107f $X=1.085 $Y=1.135 $X2=0 $Y2=0
cc_228 N_D_c_231_n N_A_294_35#_c_273_n 0.00814529f $X=1.085 $Y=1.135 $X2=0 $Y2=0
cc_229 N_D_c_230_n N_A_294_35#_c_286_n 0.00131767f $X=1.085 $Y=1.3 $X2=0 $Y2=0
cc_230 N_D_c_231_n N_A_294_35#_c_286_n 0.0117119f $X=1.085 $Y=1.135 $X2=0 $Y2=0
cc_231 N_D_M1004_g N_RESET_B_M1029_g 0.0127063f $X=1.135 $Y=2.525 $X2=0 $Y2=0
cc_232 N_D_M1004_g N_RESET_B_c_588_n 0.00996588f $X=1.135 $Y=2.525 $X2=0 $Y2=0
cc_233 N_D_M1004_g N_RESET_B_M1023_g 0.007503f $X=1.135 $Y=2.525 $X2=0 $Y2=0
cc_234 D N_RESET_B_M1023_g 0.0192116f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_235 N_D_c_231_n N_RESET_B_M1023_g 0.0775755f $X=1.085 $Y=1.135 $X2=0 $Y2=0
cc_236 N_D_M1004_g N_RESET_B_c_594_n 0.0153418f $X=1.135 $Y=2.525 $X2=0 $Y2=0
cc_237 N_D_M1004_g N_RESET_B_c_576_n 0.00335926f $X=1.135 $Y=2.525 $X2=0 $Y2=0
cc_238 D N_RESET_B_c_576_n 0.0235465f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_239 N_D_c_230_n N_RESET_B_c_576_n 0.0039933f $X=1.085 $Y=1.3 $X2=0 $Y2=0
cc_240 D N_RESET_B_c_577_n 0.00803612f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_241 D N_RESET_B_c_581_n 0.00610826f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_242 N_D_M1004_g N_RESET_B_c_582_n 0.0020763f $X=1.135 $Y=2.525 $X2=0 $Y2=0
cc_243 D N_RESET_B_c_582_n 0.0410206f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_244 N_D_M1004_g N_A_306_277#_c_776_n 0.039379f $X=1.135 $Y=2.525 $X2=0 $Y2=0
cc_245 N_D_c_230_n N_A_306_277#_c_776_n 0.00350448f $X=1.085 $Y=1.3 $X2=0 $Y2=0
cc_246 N_D_c_230_n N_A_306_277#_c_777_n 0.00190028f $X=1.085 $Y=1.3 $X2=0 $Y2=0
cc_247 N_D_M1004_g N_A_27_463#_c_1497_n 0.0178078f $X=1.135 $Y=2.525 $X2=0 $Y2=0
cc_248 N_D_M1004_g N_A_27_463#_c_1500_n 0.0156765f $X=1.135 $Y=2.525 $X2=0 $Y2=0
cc_249 N_D_M1004_g N_A_27_463#_c_1498_n 8.98407e-19 $X=1.135 $Y=2.525 $X2=0
+ $Y2=0
cc_250 D N_A_27_463#_c_1502_n 0.0109229f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_251 N_D_c_230_n N_A_27_463#_c_1502_n 0.00255937f $X=1.085 $Y=1.3 $X2=0 $Y2=0
cc_252 N_D_c_231_n N_A_27_463#_c_1502_n 0.00533795f $X=1.085 $Y=1.135 $X2=0
+ $Y2=0
cc_253 N_D_M1004_g N_A_27_463#_c_1495_n 0.00188365f $X=1.135 $Y=2.525 $X2=0
+ $Y2=0
cc_254 D N_A_27_463#_c_1495_n 0.0205207f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_255 N_D_c_230_n N_A_27_463#_c_1495_n 0.00265631f $X=1.085 $Y=1.3 $X2=0 $Y2=0
cc_256 N_D_c_231_n N_A_27_463#_c_1495_n 0.0027112f $X=1.085 $Y=1.135 $X2=0 $Y2=0
cc_257 N_D_M1004_g N_A_27_463#_c_1496_n 0.00812563f $X=1.135 $Y=2.525 $X2=0
+ $Y2=0
cc_258 D N_A_27_463#_c_1496_n 0.0101521f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_259 N_D_c_230_n N_A_27_463#_c_1496_n 0.00101448f $X=1.085 $Y=1.3 $X2=0 $Y2=0
cc_260 N_D_M1004_g N_VPWR_c_1555_n 0.00474243f $X=1.135 $Y=2.525 $X2=0 $Y2=0
cc_261 N_D_M1004_g N_VPWR_c_1554_n 9.39239e-19 $X=1.135 $Y=2.525 $X2=0 $Y2=0
cc_262 D N_VGND_c_1689_n 0.0245369f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_263 N_D_c_231_n N_VGND_c_1689_n 0.0031963f $X=1.085 $Y=1.135 $X2=0 $Y2=0
cc_264 N_D_c_231_n N_VGND_c_1694_n 0.00478016f $X=1.085 $Y=1.135 $X2=0 $Y2=0
cc_265 N_D_c_231_n N_VGND_c_1702_n 0.00948019f $X=1.085 $Y=1.135 $X2=0 $Y2=0
cc_266 N_A_294_35#_c_278_n N_A_501_229#_M1028_d 0.00511607f $X=5.66 $Y=0.34
+ $X2=-0.19 $Y2=-0.245
cc_267 N_A_294_35#_M1002_g N_A_501_229#_M1015_g 0.024745f $X=2.16 $Y=2.525 $X2=0
+ $Y2=0
cc_268 N_A_294_35#_c_275_n N_A_501_229#_M1015_g 0.00394325f $X=2.25 $Y=1.91
+ $X2=0 $Y2=0
cc_269 N_A_294_35#_c_291_n N_A_501_229#_M1015_g 0.0215646f $X=2.25 $Y=1.91 $X2=0
+ $Y2=0
cc_270 N_A_294_35#_c_293_n N_A_501_229#_M1015_g 0.0102963f $X=4.035 $Y=2.015
+ $X2=0 $Y2=0
cc_271 N_A_294_35#_c_276_n N_A_501_229#_c_469_n 0.0733194f $X=3.915 $Y=0.795
+ $X2=0 $Y2=0
cc_272 N_A_294_35#_c_306_p N_A_501_229#_c_469_n 0.00403163f $X=4.97 $Y=0.675
+ $X2=0 $Y2=0
cc_273 N_A_294_35#_c_277_n N_A_501_229#_c_469_n 0.020945f $X=4.245 $Y=0.675
+ $X2=0 $Y2=0
cc_274 N_A_294_35#_M1003_g N_A_501_229#_c_470_n 0.00480154f $X=5.42 $Y=2.655
+ $X2=0 $Y2=0
cc_275 N_A_294_35#_c_280_n N_A_501_229#_c_470_n 0.0102613f $X=5.745 $Y=1.48
+ $X2=0 $Y2=0
cc_276 N_A_294_35#_c_283_n N_A_501_229#_c_470_n 0.022756f $X=5.47 $Y=1.645 $X2=0
+ $Y2=0
cc_277 N_A_294_35#_c_284_n N_A_501_229#_c_470_n 0.00199174f $X=5.47 $Y=1.645
+ $X2=0 $Y2=0
cc_278 N_A_294_35#_c_278_n N_A_501_229#_c_491_n 0.0120642f $X=5.66 $Y=0.34 $X2=0
+ $Y2=0
cc_279 N_A_294_35#_c_275_n N_A_501_229#_c_471_n 0.026433f $X=2.25 $Y=1.91 $X2=0
+ $Y2=0
cc_280 N_A_294_35#_c_276_n N_A_501_229#_c_471_n 0.0211138f $X=3.915 $Y=0.795
+ $X2=0 $Y2=0
cc_281 N_A_294_35#_c_293_n N_A_501_229#_c_471_n 6.54133e-19 $X=4.035 $Y=2.015
+ $X2=0 $Y2=0
cc_282 N_A_294_35#_c_275_n N_A_501_229#_c_472_n 0.00360786f $X=2.25 $Y=1.91
+ $X2=0 $Y2=0
cc_283 N_A_294_35#_c_276_n N_A_501_229#_c_472_n 6.29107e-19 $X=3.915 $Y=0.795
+ $X2=0 $Y2=0
cc_284 N_A_294_35#_c_293_n N_A_501_229#_c_472_n 0.00105705f $X=4.035 $Y=2.015
+ $X2=0 $Y2=0
cc_285 N_A_294_35#_c_306_p N_A_501_229#_c_473_n 0.00821848f $X=4.97 $Y=0.675
+ $X2=0 $Y2=0
cc_286 N_A_294_35#_c_306_p N_A_501_229#_c_474_n 0.039044f $X=4.97 $Y=0.675 $X2=0
+ $Y2=0
cc_287 N_A_294_35#_c_278_n N_A_501_229#_c_475_n 0.00529894f $X=5.66 $Y=0.34
+ $X2=0 $Y2=0
cc_288 N_A_294_35#_c_280_n N_A_501_229#_c_475_n 0.019076f $X=5.745 $Y=1.48 $X2=0
+ $Y2=0
cc_289 N_A_294_35#_c_283_n N_A_501_229#_c_475_n 0.00451812f $X=5.47 $Y=1.645
+ $X2=0 $Y2=0
cc_290 N_A_294_35#_c_284_n N_A_501_229#_c_475_n 0.00359411f $X=5.47 $Y=1.645
+ $X2=0 $Y2=0
cc_291 N_A_294_35#_M1003_g N_A_501_229#_c_504_n 0.00300044f $X=5.42 $Y=2.655
+ $X2=0 $Y2=0
cc_292 N_A_294_35#_c_274_n N_A_501_229#_c_476_n 0.00460994f $X=2.245 $Y=0.71
+ $X2=0 $Y2=0
cc_293 N_A_294_35#_c_275_n N_A_501_229#_c_476_n 0.00376846f $X=2.25 $Y=1.91
+ $X2=0 $Y2=0
cc_294 N_A_294_35#_c_276_n N_A_501_229#_c_476_n 0.0118504f $X=3.915 $Y=0.795
+ $X2=0 $Y2=0
cc_295 N_A_294_35#_M1002_g N_RESET_B_c_588_n 0.0101001f $X=2.16 $Y=2.525 $X2=0
+ $Y2=0
cc_296 N_A_294_35#_c_276_n N_RESET_B_M1031_g 0.0122037f $X=3.915 $Y=0.795 $X2=0
+ $Y2=0
cc_297 N_A_294_35#_c_293_n N_RESET_B_c_590_n 0.0146408f $X=4.035 $Y=2.015 $X2=0
+ $Y2=0
cc_298 N_A_294_35#_c_293_n N_RESET_B_c_596_n 0.00480714f $X=4.035 $Y=2.015 $X2=0
+ $Y2=0
cc_299 N_A_294_35#_c_275_n N_RESET_B_c_576_n 0.0177979f $X=2.25 $Y=1.91 $X2=0
+ $Y2=0
cc_300 N_A_294_35#_c_291_n N_RESET_B_c_576_n 0.00333701f $X=2.25 $Y=1.91 $X2=0
+ $Y2=0
cc_301 N_A_294_35#_c_293_n N_RESET_B_c_576_n 0.00685766f $X=4.035 $Y=2.015 $X2=0
+ $Y2=0
cc_302 N_A_294_35#_c_286_n N_RESET_B_c_576_n 2.16771e-19 $X=1.635 $Y=0.505 $X2=0
+ $Y2=0
cc_303 N_A_294_35#_c_293_n N_RESET_B_c_578_n 0.0444817f $X=4.035 $Y=2.015 $X2=0
+ $Y2=0
cc_304 N_A_294_35#_c_283_n N_RESET_B_c_578_n 0.0291915f $X=5.47 $Y=1.645 $X2=0
+ $Y2=0
cc_305 N_A_294_35#_c_284_n N_RESET_B_c_578_n 0.00368395f $X=5.47 $Y=1.645 $X2=0
+ $Y2=0
cc_306 N_A_294_35#_c_287_n N_RESET_B_c_578_n 0.0036078f $X=6.21 $Y=0.515 $X2=0
+ $Y2=0
cc_307 N_A_294_35#_c_275_n N_RESET_B_c_579_n 0.00349019f $X=2.25 $Y=1.91 $X2=0
+ $Y2=0
cc_308 N_A_294_35#_c_291_n N_RESET_B_c_579_n 5.68001e-19 $X=2.25 $Y=1.91 $X2=0
+ $Y2=0
cc_309 N_A_294_35#_c_293_n N_RESET_B_c_579_n 0.00808928f $X=4.035 $Y=2.015 $X2=0
+ $Y2=0
cc_310 N_A_294_35#_c_293_n N_RESET_B_c_585_n 2.42426e-19 $X=4.035 $Y=2.015 $X2=0
+ $Y2=0
cc_311 N_A_294_35#_c_275_n N_RESET_B_c_586_n 0.0100909f $X=2.25 $Y=1.91 $X2=0
+ $Y2=0
cc_312 N_A_294_35#_c_293_n N_RESET_B_c_586_n 0.0527834f $X=4.035 $Y=2.015 $X2=0
+ $Y2=0
cc_313 N_A_294_35#_c_291_n N_A_306_277#_M1030_g 0.021441f $X=2.25 $Y=1.91 $X2=0
+ $Y2=0
cc_314 N_A_294_35#_c_286_n N_A_306_277#_c_776_n 0.0111194f $X=1.635 $Y=0.505
+ $X2=0 $Y2=0
cc_315 N_A_294_35#_c_272_n N_A_306_277#_c_777_n 0.00143082f $X=2.155 $Y=0.367
+ $X2=0 $Y2=0
cc_316 N_A_294_35#_c_275_n N_A_306_277#_c_777_n 0.00715279f $X=2.25 $Y=1.91
+ $X2=0 $Y2=0
cc_317 N_A_294_35#_c_291_n N_A_306_277#_c_777_n 0.00455573f $X=2.25 $Y=1.91
+ $X2=0 $Y2=0
cc_318 N_A_294_35#_c_286_n N_A_306_277#_c_777_n 0.00357022f $X=1.635 $Y=0.505
+ $X2=0 $Y2=0
cc_319 N_A_294_35#_c_272_n N_A_306_277#_M1011_g 0.0154575f $X=2.155 $Y=0.367
+ $X2=0 $Y2=0
cc_320 N_A_294_35#_c_274_n N_A_306_277#_M1011_g 0.00589014f $X=2.245 $Y=0.71
+ $X2=0 $Y2=0
cc_321 N_A_294_35#_c_275_n N_A_306_277#_M1011_g 0.00451923f $X=2.25 $Y=1.91
+ $X2=0 $Y2=0
cc_322 N_A_294_35#_c_356_p N_A_306_277#_M1011_g 0.00427676f $X=2.245 $Y=0.795
+ $X2=0 $Y2=0
cc_323 N_A_294_35#_c_286_n N_A_306_277#_M1011_g 0.00860374f $X=1.635 $Y=0.505
+ $X2=0 $Y2=0
cc_324 N_A_294_35#_c_272_n N_A_306_277#_c_779_n 0.00255845f $X=2.155 $Y=0.367
+ $X2=0 $Y2=0
cc_325 N_A_294_35#_c_276_n N_A_306_277#_c_779_n 0.0104567f $X=3.915 $Y=0.795
+ $X2=0 $Y2=0
cc_326 N_A_294_35#_c_272_n N_A_306_277#_c_780_n 2.99808e-19 $X=2.155 $Y=0.367
+ $X2=0 $Y2=0
cc_327 N_A_294_35#_c_273_n N_A_306_277#_c_780_n 0.0187484f $X=1.635 $Y=0.34
+ $X2=0 $Y2=0
cc_328 N_A_294_35#_c_276_n N_A_306_277#_c_781_n 0.0172408f $X=3.915 $Y=0.795
+ $X2=0 $Y2=0
cc_329 N_A_294_35#_c_277_n N_A_306_277#_c_781_n 0.00518403f $X=4.245 $Y=0.675
+ $X2=0 $Y2=0
cc_330 N_A_294_35#_c_277_n N_A_306_277#_c_782_n 0.00384172f $X=4.245 $Y=0.675
+ $X2=0 $Y2=0
cc_331 N_A_294_35#_c_306_p N_A_306_277#_c_784_n 0.0102773f $X=4.97 $Y=0.675
+ $X2=0 $Y2=0
cc_332 N_A_294_35#_c_277_n N_A_306_277#_c_784_n 0.00120481f $X=4.245 $Y=0.675
+ $X2=0 $Y2=0
cc_333 N_A_294_35#_c_367_p N_A_306_277#_c_784_n 7.89798e-19 $X=5.055 $Y=0.585
+ $X2=0 $Y2=0
cc_334 N_A_294_35#_c_293_n N_A_306_277#_M1008_g 0.00850276f $X=4.035 $Y=2.015
+ $X2=0 $Y2=0
cc_335 N_A_294_35#_c_278_n N_A_306_277#_M1007_g 0.0109656f $X=5.66 $Y=0.34 $X2=0
+ $Y2=0
cc_336 N_A_294_35#_c_280_n N_A_306_277#_M1007_g 0.0164033f $X=5.745 $Y=1.48
+ $X2=0 $Y2=0
cc_337 N_A_294_35#_c_282_n N_A_306_277#_M1007_g 0.0106413f $X=6.21 $Y=0.35 $X2=0
+ $Y2=0
cc_338 N_A_294_35#_c_285_n N_A_306_277#_M1007_g 0.00328101f $X=5.745 $Y=0.345
+ $X2=0 $Y2=0
cc_339 N_A_294_35#_c_287_n N_A_306_277#_M1007_g 0.00702265f $X=6.21 $Y=0.515
+ $X2=0 $Y2=0
cc_340 N_A_294_35#_c_280_n N_A_306_277#_c_787_n 0.0100231f $X=5.745 $Y=1.48
+ $X2=0 $Y2=0
cc_341 N_A_294_35#_c_281_n N_A_306_277#_c_787_n 0.00396962f $X=6.21 $Y=0.35
+ $X2=0 $Y2=0
cc_342 N_A_294_35#_c_287_n N_A_306_277#_c_787_n 0.00275836f $X=6.21 $Y=0.515
+ $X2=0 $Y2=0
cc_343 N_A_294_35#_c_280_n N_A_306_277#_c_788_n 0.00252429f $X=5.745 $Y=1.48
+ $X2=0 $Y2=0
cc_344 N_A_294_35#_c_283_n N_A_306_277#_c_788_n 0.00180959f $X=5.47 $Y=1.645
+ $X2=0 $Y2=0
cc_345 N_A_294_35#_c_284_n N_A_306_277#_c_788_n 0.00667168f $X=5.47 $Y=1.645
+ $X2=0 $Y2=0
cc_346 N_A_294_35#_M1003_g N_A_306_277#_M1005_g 0.0147196f $X=5.42 $Y=2.655
+ $X2=0 $Y2=0
cc_347 N_A_294_35#_M1003_g N_A_306_277#_c_850_n 0.0127368f $X=5.42 $Y=2.655
+ $X2=0 $Y2=0
cc_348 N_A_294_35#_M1003_g N_A_306_277#_c_851_n 0.00646619f $X=5.42 $Y=2.655
+ $X2=0 $Y2=0
cc_349 N_A_294_35#_M1003_g N_A_306_277#_c_808_n 0.0019166f $X=5.42 $Y=2.655
+ $X2=0 $Y2=0
cc_350 N_A_294_35#_M1003_g N_A_306_277#_c_794_n 0.0161625f $X=5.42 $Y=2.655
+ $X2=0 $Y2=0
cc_351 N_A_294_35#_c_280_n N_A_306_277#_c_794_n 0.00481687f $X=5.745 $Y=1.48
+ $X2=0 $Y2=0
cc_352 N_A_294_35#_c_283_n N_A_306_277#_c_794_n 0.00192149f $X=5.47 $Y=1.645
+ $X2=0 $Y2=0
cc_353 N_A_294_35#_c_284_n N_A_306_277#_c_794_n 0.0206036f $X=5.47 $Y=1.645
+ $X2=0 $Y2=0
cc_354 N_A_294_35#_M1003_g N_A_336_463#_M1017_g 0.0469934f $X=5.42 $Y=2.655
+ $X2=0 $Y2=0
cc_355 N_A_294_35#_c_306_p N_A_336_463#_M1028_g 0.00982196f $X=4.97 $Y=0.675
+ $X2=0 $Y2=0
cc_356 N_A_294_35#_c_367_p N_A_336_463#_M1028_g 0.00569505f $X=5.055 $Y=0.585
+ $X2=0 $Y2=0
cc_357 N_A_294_35#_c_279_n N_A_336_463#_M1028_g 0.00663757f $X=5.14 $Y=0.34
+ $X2=0 $Y2=0
cc_358 N_A_294_35#_c_280_n N_A_336_463#_M1028_g 0.00144297f $X=5.745 $Y=1.48
+ $X2=0 $Y2=0
cc_359 N_A_294_35#_c_272_n N_A_336_463#_c_1048_n 0.0126346f $X=2.155 $Y=0.367
+ $X2=0 $Y2=0
cc_360 N_A_294_35#_c_275_n N_A_336_463#_c_1048_n 0.0682685f $X=2.25 $Y=1.91
+ $X2=0 $Y2=0
cc_361 N_A_294_35#_c_291_n N_A_336_463#_c_1048_n 0.00299963f $X=2.25 $Y=1.91
+ $X2=0 $Y2=0
cc_362 N_A_294_35#_c_292_n N_A_336_463#_c_1048_n 0.0131592f $X=2.335 $Y=2.01
+ $X2=0 $Y2=0
cc_363 N_A_294_35#_c_286_n N_A_336_463#_c_1048_n 9.37404e-19 $X=1.635 $Y=0.505
+ $X2=0 $Y2=0
cc_364 N_A_294_35#_M1002_g N_A_336_463#_c_1053_n 0.0110651f $X=2.16 $Y=2.525
+ $X2=0 $Y2=0
cc_365 N_A_294_35#_c_291_n N_A_336_463#_c_1053_n 0.00119747f $X=2.25 $Y=1.91
+ $X2=0 $Y2=0
cc_366 N_A_294_35#_c_292_n N_A_336_463#_c_1053_n 0.0140936f $X=2.335 $Y=2.01
+ $X2=0 $Y2=0
cc_367 N_A_294_35#_c_293_n N_A_336_463#_c_1053_n 0.0947914f $X=4.035 $Y=2.015
+ $X2=0 $Y2=0
cc_368 N_A_294_35#_M1008_s N_A_336_463#_c_1054_n 0.00996611f $X=3.91 $Y=1.835
+ $X2=0 $Y2=0
cc_369 N_A_294_35#_c_293_n N_A_336_463#_c_1054_n 0.0410027f $X=4.035 $Y=2.015
+ $X2=0 $Y2=0
cc_370 N_A_294_35#_c_293_n N_A_336_463#_c_1049_n 0.00725836f $X=4.035 $Y=2.015
+ $X2=0 $Y2=0
cc_371 N_A_294_35#_M1002_g N_A_336_463#_c_1056_n 0.00450632f $X=2.16 $Y=2.525
+ $X2=0 $Y2=0
cc_372 N_A_294_35#_c_292_n N_A_336_463#_c_1056_n 0.00123909f $X=2.335 $Y=2.01
+ $X2=0 $Y2=0
cc_373 N_A_294_35#_c_283_n N_A_336_463#_c_1050_n 3.6011e-19 $X=5.47 $Y=1.645
+ $X2=0 $Y2=0
cc_374 N_A_294_35#_c_284_n N_A_336_463#_c_1050_n 0.0183704f $X=5.47 $Y=1.645
+ $X2=0 $Y2=0
cc_375 N_A_294_35#_c_282_n N_A_1287_276#_M1013_g 0.04212f $X=6.21 $Y=0.35 $X2=0
+ $Y2=0
cc_376 N_A_294_35#_c_280_n N_A_1099_447#_M1007_d 0.00621293f $X=5.745 $Y=1.48
+ $X2=-0.19 $Y2=-0.245
cc_377 N_A_294_35#_c_281_n N_A_1099_447#_M1007_d 0.00187632f $X=6.21 $Y=0.35
+ $X2=-0.19 $Y2=-0.245
cc_378 N_A_294_35#_M1003_g N_A_1099_447#_c_1294_n 8.26397e-19 $X=5.42 $Y=2.655
+ $X2=0 $Y2=0
cc_379 N_A_294_35#_c_280_n N_A_1099_447#_c_1284_n 0.0203928f $X=5.745 $Y=1.48
+ $X2=0 $Y2=0
cc_380 N_A_294_35#_c_281_n N_A_1099_447#_c_1284_n 0.0169172f $X=6.21 $Y=0.35
+ $X2=0 $Y2=0
cc_381 N_A_294_35#_c_282_n N_A_1099_447#_c_1284_n 0.00457674f $X=6.21 $Y=0.35
+ $X2=0 $Y2=0
cc_382 N_A_294_35#_c_287_n N_A_1099_447#_c_1284_n 3.29708e-19 $X=6.21 $Y=0.515
+ $X2=0 $Y2=0
cc_383 N_A_294_35#_c_280_n N_A_1099_447#_c_1285_n 0.0309707f $X=5.745 $Y=1.48
+ $X2=0 $Y2=0
cc_384 N_A_294_35#_c_283_n N_A_1099_447#_c_1285_n 0.0220759f $X=5.47 $Y=1.645
+ $X2=0 $Y2=0
cc_385 N_A_294_35#_c_287_n N_A_1099_447#_c_1285_n 0.00287214f $X=6.21 $Y=0.515
+ $X2=0 $Y2=0
cc_386 N_A_294_35#_c_281_n N_A_1099_447#_c_1286_n 0.00469004f $X=6.21 $Y=0.35
+ $X2=0 $Y2=0
cc_387 N_A_294_35#_c_287_n N_A_1099_447#_c_1286_n 0.0105032f $X=6.21 $Y=0.515
+ $X2=0 $Y2=0
cc_388 N_A_294_35#_M1003_g N_A_1099_447#_c_1296_n 0.00284411f $X=5.42 $Y=2.655
+ $X2=0 $Y2=0
cc_389 N_A_294_35#_c_283_n N_A_1099_447#_c_1296_n 0.0180207f $X=5.47 $Y=1.645
+ $X2=0 $Y2=0
cc_390 N_A_294_35#_c_284_n N_A_1099_447#_c_1296_n 0.00206688f $X=5.47 $Y=1.645
+ $X2=0 $Y2=0
cc_391 N_A_294_35#_c_280_n N_A_1099_447#_c_1290_n 0.0146909f $X=5.745 $Y=1.48
+ $X2=0 $Y2=0
cc_392 N_A_294_35#_c_287_n N_A_1099_447#_c_1290_n 0.00129385f $X=6.21 $Y=0.515
+ $X2=0 $Y2=0
cc_393 N_A_294_35#_c_272_n N_A_27_463#_c_1502_n 0.00966059f $X=2.155 $Y=0.367
+ $X2=0 $Y2=0
cc_394 N_A_294_35#_c_273_n N_A_27_463#_c_1502_n 0.00289777f $X=1.635 $Y=0.34
+ $X2=0 $Y2=0
cc_395 N_A_294_35#_c_274_n N_A_27_463#_c_1502_n 7.13058e-19 $X=2.245 $Y=0.71
+ $X2=0 $Y2=0
cc_396 N_A_294_35#_c_286_n N_A_27_463#_c_1502_n 0.00989803f $X=1.635 $Y=0.505
+ $X2=0 $Y2=0
cc_397 N_A_294_35#_c_286_n N_A_27_463#_c_1495_n 0.00467544f $X=1.635 $Y=0.505
+ $X2=0 $Y2=0
cc_398 N_A_294_35#_M1003_g N_VPWR_c_1561_n 0.00372091f $X=5.42 $Y=2.655 $X2=0
+ $Y2=0
cc_399 N_A_294_35#_M1002_g N_VPWR_c_1554_n 9.39239e-19 $X=2.16 $Y=2.525 $X2=0
+ $Y2=0
cc_400 N_A_294_35#_M1003_g N_VPWR_c_1554_n 0.00575806f $X=5.42 $Y=2.655 $X2=0
+ $Y2=0
cc_401 N_A_294_35#_c_276_n N_VGND_M1031_d 0.00672482f $X=3.915 $Y=0.795 $X2=0
+ $Y2=0
cc_402 N_A_294_35#_c_306_p N_VGND_M1016_d 0.0116066f $X=4.97 $Y=0.675 $X2=0
+ $Y2=0
cc_403 N_A_294_35#_c_276_n N_VGND_c_1690_n 0.0256127f $X=3.915 $Y=0.795 $X2=0
+ $Y2=0
cc_404 N_A_294_35#_c_281_n N_VGND_c_1691_n 0.00764423f $X=6.21 $Y=0.35 $X2=0
+ $Y2=0
cc_405 N_A_294_35#_c_282_n N_VGND_c_1691_n 0.0048738f $X=6.21 $Y=0.35 $X2=0
+ $Y2=0
cc_406 N_A_294_35#_c_272_n N_VGND_c_1694_n 0.0558605f $X=2.155 $Y=0.367 $X2=0
+ $Y2=0
cc_407 N_A_294_35#_c_273_n N_VGND_c_1694_n 0.00659816f $X=1.635 $Y=0.34 $X2=0
+ $Y2=0
cc_408 N_A_294_35#_c_276_n N_VGND_c_1694_n 0.0117357f $X=3.915 $Y=0.795 $X2=0
+ $Y2=0
cc_409 N_A_294_35#_c_276_n N_VGND_c_1698_n 0.00481146f $X=3.915 $Y=0.795 $X2=0
+ $Y2=0
cc_410 N_A_294_35#_c_306_p N_VGND_c_1698_n 0.0037653f $X=4.97 $Y=0.675 $X2=0
+ $Y2=0
cc_411 N_A_294_35#_c_277_n N_VGND_c_1698_n 0.00677348f $X=4.245 $Y=0.675 $X2=0
+ $Y2=0
cc_412 N_A_294_35#_c_306_p N_VGND_c_1699_n 0.00282015f $X=4.97 $Y=0.675 $X2=0
+ $Y2=0
cc_413 N_A_294_35#_c_278_n N_VGND_c_1699_n 0.0330783f $X=5.66 $Y=0.34 $X2=0
+ $Y2=0
cc_414 N_A_294_35#_c_279_n N_VGND_c_1699_n 0.0115034f $X=5.14 $Y=0.34 $X2=0
+ $Y2=0
cc_415 N_A_294_35#_c_281_n N_VGND_c_1699_n 0.0342492f $X=6.21 $Y=0.35 $X2=0
+ $Y2=0
cc_416 N_A_294_35#_c_282_n N_VGND_c_1699_n 0.00647615f $X=6.21 $Y=0.35 $X2=0
+ $Y2=0
cc_417 N_A_294_35#_c_285_n N_VGND_c_1699_n 0.0120989f $X=5.745 $Y=0.345 $X2=0
+ $Y2=0
cc_418 N_A_294_35#_c_272_n N_VGND_c_1702_n 0.0300189f $X=2.155 $Y=0.367 $X2=0
+ $Y2=0
cc_419 N_A_294_35#_c_273_n N_VGND_c_1702_n 0.00946248f $X=1.635 $Y=0.34 $X2=0
+ $Y2=0
cc_420 N_A_294_35#_c_276_n N_VGND_c_1702_n 0.0297987f $X=3.915 $Y=0.795 $X2=0
+ $Y2=0
cc_421 N_A_294_35#_c_306_p N_VGND_c_1702_n 0.0131873f $X=4.97 $Y=0.675 $X2=0
+ $Y2=0
cc_422 N_A_294_35#_c_277_n N_VGND_c_1702_n 0.0102743f $X=4.245 $Y=0.675 $X2=0
+ $Y2=0
cc_423 N_A_294_35#_c_278_n N_VGND_c_1702_n 0.0189745f $X=5.66 $Y=0.34 $X2=0
+ $Y2=0
cc_424 N_A_294_35#_c_279_n N_VGND_c_1702_n 0.00598876f $X=5.14 $Y=0.34 $X2=0
+ $Y2=0
cc_425 N_A_294_35#_c_281_n N_VGND_c_1702_n 0.0190094f $X=6.21 $Y=0.35 $X2=0
+ $Y2=0
cc_426 N_A_294_35#_c_282_n N_VGND_c_1702_n 0.00966139f $X=6.21 $Y=0.35 $X2=0
+ $Y2=0
cc_427 N_A_294_35#_c_285_n N_VGND_c_1702_n 0.00649482f $X=5.745 $Y=0.345 $X2=0
+ $Y2=0
cc_428 N_A_294_35#_c_306_p N_VGND_c_1703_n 0.0247132f $X=4.97 $Y=0.675 $X2=0
+ $Y2=0
cc_429 N_A_294_35#_c_279_n N_VGND_c_1703_n 0.0132902f $X=5.14 $Y=0.34 $X2=0
+ $Y2=0
cc_430 N_A_294_35#_c_274_n A_438_123# 0.00113389f $X=2.245 $Y=0.71 $X2=-0.19
+ $Y2=-0.245
cc_431 N_A_294_35#_c_275_n A_438_123# 0.00185765f $X=2.25 $Y=1.91 $X2=-0.19
+ $Y2=-0.245
cc_432 N_A_294_35#_c_276_n A_438_123# 0.00839362f $X=3.915 $Y=0.795 $X2=-0.19
+ $Y2=-0.245
cc_433 N_A_294_35#_c_276_n A_540_123# 0.00583264f $X=3.915 $Y=0.795 $X2=-0.19
+ $Y2=-0.245
cc_434 N_A_501_229#_M1015_g N_RESET_B_c_588_n 0.0101001f $X=2.7 $Y=2.525 $X2=0
+ $Y2=0
cc_435 N_A_501_229#_M1015_g N_RESET_B_M1031_g 0.039348f $X=2.7 $Y=2.525 $X2=0
+ $Y2=0
cc_436 N_A_501_229#_c_469_n N_RESET_B_M1031_g 0.0119503f $X=4.335 $Y=1.135 $X2=0
+ $Y2=0
cc_437 N_A_501_229#_c_471_n N_RESET_B_M1031_g 0.00131701f $X=2.67 $Y=1.135 $X2=0
+ $Y2=0
cc_438 N_A_501_229#_c_472_n N_RESET_B_M1031_g 0.0216916f $X=2.67 $Y=1.31 $X2=0
+ $Y2=0
cc_439 N_A_501_229#_c_476_n N_RESET_B_M1031_g 0.0254331f $X=2.67 $Y=1.145 $X2=0
+ $Y2=0
cc_440 N_A_501_229#_M1015_g N_RESET_B_M1022_g 0.0144319f $X=2.7 $Y=2.525 $X2=0
+ $Y2=0
cc_441 N_A_501_229#_c_469_n N_RESET_B_c_578_n 0.0384802f $X=4.335 $Y=1.135 $X2=0
+ $Y2=0
cc_442 N_A_501_229#_c_470_n N_RESET_B_c_578_n 0.0116543f $X=5.115 $Y=2.245 $X2=0
+ $Y2=0
cc_443 N_A_501_229#_c_471_n N_RESET_B_c_578_n 3.44377e-19 $X=2.67 $Y=1.135 $X2=0
+ $Y2=0
cc_444 N_A_501_229#_c_473_n N_RESET_B_c_578_n 0.00623901f $X=4.42 $Y=1.02 $X2=0
+ $Y2=0
cc_445 N_A_501_229#_c_474_n N_RESET_B_c_578_n 0.011244f $X=5.025 $Y=1.07 $X2=0
+ $Y2=0
cc_446 N_A_501_229#_c_475_n N_RESET_B_c_578_n 0.00774726f $X=5.395 $Y=1.07 $X2=0
+ $Y2=0
cc_447 N_A_501_229#_c_504_n N_RESET_B_c_578_n 0.00562515f $X=5.205 $Y=2.36 $X2=0
+ $Y2=0
cc_448 N_A_501_229#_M1015_g N_RESET_B_c_579_n 0.00285523f $X=2.7 $Y=2.525 $X2=0
+ $Y2=0
cc_449 N_A_501_229#_c_471_n N_RESET_B_c_579_n 0.00745627f $X=2.67 $Y=1.135 $X2=0
+ $Y2=0
cc_450 N_A_501_229#_c_472_n N_RESET_B_c_579_n 0.00385318f $X=2.67 $Y=1.31 $X2=0
+ $Y2=0
cc_451 N_A_501_229#_c_469_n N_RESET_B_c_585_n 0.00451626f $X=4.335 $Y=1.135
+ $X2=0 $Y2=0
cc_452 N_A_501_229#_M1015_g N_RESET_B_c_586_n 0.00969248f $X=2.7 $Y=2.525 $X2=0
+ $Y2=0
cc_453 N_A_501_229#_c_469_n N_RESET_B_c_586_n 0.0192516f $X=4.335 $Y=1.135 $X2=0
+ $Y2=0
cc_454 N_A_501_229#_c_471_n N_RESET_B_c_586_n 0.018207f $X=2.67 $Y=1.135 $X2=0
+ $Y2=0
cc_455 N_A_501_229#_c_472_n N_RESET_B_c_586_n 0.00348938f $X=2.67 $Y=1.31 $X2=0
+ $Y2=0
cc_456 N_A_501_229#_M1015_g N_A_306_277#_c_777_n 9.90593e-19 $X=2.7 $Y=2.525
+ $X2=0 $Y2=0
cc_457 N_A_501_229#_c_472_n N_A_306_277#_c_777_n 0.00951197f $X=2.67 $Y=1.31
+ $X2=0 $Y2=0
cc_458 N_A_501_229#_c_471_n N_A_306_277#_M1011_g 2.52457e-19 $X=2.67 $Y=1.135
+ $X2=0 $Y2=0
cc_459 N_A_501_229#_c_476_n N_A_306_277#_M1011_g 0.0199582f $X=2.67 $Y=1.145
+ $X2=0 $Y2=0
cc_460 N_A_501_229#_c_476_n N_A_306_277#_c_779_n 0.0088955f $X=2.67 $Y=1.145
+ $X2=0 $Y2=0
cc_461 N_A_501_229#_c_473_n N_A_306_277#_c_781_n 5.36282e-19 $X=4.42 $Y=1.02
+ $X2=0 $Y2=0
cc_462 N_A_501_229#_c_469_n N_A_306_277#_c_782_n 0.0140129f $X=4.335 $Y=1.135
+ $X2=0 $Y2=0
cc_463 N_A_501_229#_c_469_n N_A_306_277#_c_783_n 0.0116057f $X=4.335 $Y=1.135
+ $X2=0 $Y2=0
cc_464 N_A_501_229#_c_473_n N_A_306_277#_c_784_n 0.00399646f $X=4.42 $Y=1.02
+ $X2=0 $Y2=0
cc_465 N_A_501_229#_c_474_n N_A_306_277#_c_784_n 3.7338e-19 $X=5.025 $Y=1.07
+ $X2=0 $Y2=0
cc_466 N_A_501_229#_c_469_n N_A_306_277#_M1008_g 0.00229709f $X=4.335 $Y=1.135
+ $X2=0 $Y2=0
cc_467 N_A_501_229#_c_470_n N_A_306_277#_M1008_g 5.19963e-19 $X=5.115 $Y=2.245
+ $X2=0 $Y2=0
cc_468 N_A_501_229#_c_473_n N_A_306_277#_M1008_g 0.00155987f $X=4.42 $Y=1.02
+ $X2=0 $Y2=0
cc_469 N_A_501_229#_c_475_n N_A_306_277#_M1007_g 0.00261653f $X=5.395 $Y=1.07
+ $X2=0 $Y2=0
cc_470 N_A_501_229#_c_470_n N_A_306_277#_c_788_n 5.66581e-19 $X=5.115 $Y=2.245
+ $X2=0 $Y2=0
cc_471 N_A_501_229#_c_469_n N_A_306_277#_c_789_n 0.00354752f $X=4.335 $Y=1.135
+ $X2=0 $Y2=0
cc_472 N_A_501_229#_c_473_n N_A_306_277#_c_789_n 0.00334836f $X=4.42 $Y=1.02
+ $X2=0 $Y2=0
cc_473 N_A_501_229#_M1017_d N_A_306_277#_c_798_n 0.00243029f $X=5.065 $Y=2.235
+ $X2=0 $Y2=0
cc_474 N_A_501_229#_c_504_n N_A_306_277#_c_798_n 0.00844254f $X=5.205 $Y=2.36
+ $X2=0 $Y2=0
cc_475 N_A_501_229#_M1017_d N_A_306_277#_c_851_n 0.00396689f $X=5.065 $Y=2.235
+ $X2=0 $Y2=0
cc_476 N_A_501_229#_c_504_n N_A_306_277#_c_851_n 0.00845703f $X=5.205 $Y=2.36
+ $X2=0 $Y2=0
cc_477 N_A_501_229#_c_470_n N_A_306_277#_c_794_n 6.65272e-19 $X=5.115 $Y=2.245
+ $X2=0 $Y2=0
cc_478 N_A_501_229#_c_470_n N_A_336_463#_M1017_g 0.0114591f $X=5.115 $Y=2.245
+ $X2=0 $Y2=0
cc_479 N_A_501_229#_c_504_n N_A_336_463#_M1017_g 0.00322732f $X=5.205 $Y=2.36
+ $X2=0 $Y2=0
cc_480 N_A_501_229#_c_470_n N_A_336_463#_M1028_g 0.00248343f $X=5.115 $Y=2.245
+ $X2=0 $Y2=0
cc_481 N_A_501_229#_c_491_n N_A_336_463#_M1028_g 0.00412662f $X=5.395 $Y=0.76
+ $X2=0 $Y2=0
cc_482 N_A_501_229#_c_473_n N_A_336_463#_M1028_g 0.00100111f $X=4.42 $Y=1.02
+ $X2=0 $Y2=0
cc_483 N_A_501_229#_c_474_n N_A_336_463#_M1028_g 0.00694645f $X=5.025 $Y=1.07
+ $X2=0 $Y2=0
cc_484 N_A_501_229#_c_475_n N_A_336_463#_M1028_g 0.00840546f $X=5.395 $Y=1.07
+ $X2=0 $Y2=0
cc_485 N_A_501_229#_M1015_g N_A_336_463#_c_1053_n 0.0134975f $X=2.7 $Y=2.525
+ $X2=0 $Y2=0
cc_486 N_A_501_229#_c_504_n N_A_336_463#_c_1054_n 0.0135357f $X=5.205 $Y=2.36
+ $X2=0 $Y2=0
cc_487 N_A_501_229#_c_470_n N_A_336_463#_c_1049_n 0.0647845f $X=5.115 $Y=2.245
+ $X2=0 $Y2=0
cc_488 N_A_501_229#_c_474_n N_A_336_463#_c_1049_n 0.012967f $X=5.025 $Y=1.07
+ $X2=0 $Y2=0
cc_489 N_A_501_229#_c_504_n N_A_336_463#_c_1049_n 0.00167448f $X=5.205 $Y=2.36
+ $X2=0 $Y2=0
cc_490 N_A_501_229#_c_470_n N_A_336_463#_c_1050_n 0.0112118f $X=5.115 $Y=2.245
+ $X2=0 $Y2=0
cc_491 N_A_501_229#_c_474_n N_A_336_463#_c_1050_n 0.00813957f $X=5.025 $Y=1.07
+ $X2=0 $Y2=0
cc_492 N_A_501_229#_c_470_n N_A_1099_447#_c_1294_n 0.00396295f $X=5.115 $Y=2.245
+ $X2=0 $Y2=0
cc_493 N_A_501_229#_c_470_n N_A_1099_447#_c_1296_n 0.0119518f $X=5.115 $Y=2.245
+ $X2=0 $Y2=0
cc_494 N_A_501_229#_M1015_g N_VPWR_c_1556_n 0.00453079f $X=2.7 $Y=2.525 $X2=0
+ $Y2=0
cc_495 N_A_501_229#_M1015_g N_VPWR_c_1554_n 9.39239e-19 $X=2.7 $Y=2.525 $X2=0
+ $Y2=0
cc_496 N_A_501_229#_c_473_n N_VGND_M1016_d 7.46626e-19 $X=4.42 $Y=1.02 $X2=0
+ $Y2=0
cc_497 N_A_501_229#_c_474_n N_VGND_M1016_d 0.00447145f $X=5.025 $Y=1.07 $X2=0
+ $Y2=0
cc_498 N_A_501_229#_c_476_n N_VGND_c_1702_n 9.46663e-19 $X=2.67 $Y=1.145 $X2=0
+ $Y2=0
cc_499 N_RESET_B_c_588_n N_A_306_277#_M1030_g 0.010259f $X=3.215 $Y=3.15 $X2=0
+ $Y2=0
cc_500 N_RESET_B_c_576_n N_A_306_277#_M1030_g 0.00491761f $X=2.495 $Y=1.665
+ $X2=0 $Y2=0
cc_501 N_RESET_B_c_576_n N_A_306_277#_c_775_n 0.00618561f $X=2.495 $Y=1.665
+ $X2=0 $Y2=0
cc_502 N_RESET_B_c_576_n N_A_306_277#_c_777_n 5.01403e-19 $X=2.495 $Y=1.665
+ $X2=0 $Y2=0
cc_503 N_RESET_B_M1031_g N_A_306_277#_c_779_n 0.0088955f $X=3.12 $Y=0.825 $X2=0
+ $Y2=0
cc_504 N_RESET_B_M1031_g N_A_306_277#_c_781_n 0.0203057f $X=3.12 $Y=0.825 $X2=0
+ $Y2=0
cc_505 N_RESET_B_c_578_n N_A_306_277#_M1008_g 0.00814325f $X=6.815 $Y=1.665
+ $X2=0 $Y2=0
cc_506 N_RESET_B_c_578_n N_A_306_277#_c_788_n 3.05922e-19 $X=6.815 $Y=1.665
+ $X2=0 $Y2=0
cc_507 N_RESET_B_c_592_n N_A_306_277#_c_800_n 6.46241e-19 $X=7.21 $Y=2.25 $X2=0
+ $Y2=0
cc_508 N_RESET_B_M1000_g N_A_306_277#_c_800_n 0.00771082f $X=7.21 $Y=2.865 $X2=0
+ $Y2=0
cc_509 N_RESET_B_c_584_n N_A_306_277#_c_800_n 0.00620864f $X=7.21 $Y=1.745 $X2=0
+ $Y2=0
cc_510 N_RESET_B_c_608_n N_A_306_277#_c_800_n 0.016575f $X=7.17 $Y=1.707 $X2=0
+ $Y2=0
cc_511 N_RESET_B_M1000_g N_A_306_277#_c_801_n 0.0087683f $X=7.21 $Y=2.865 $X2=0
+ $Y2=0
cc_512 N_RESET_B_c_592_n N_A_306_277#_c_802_n 0.00153654f $X=7.21 $Y=2.25 $X2=0
+ $Y2=0
cc_513 N_RESET_B_M1000_g N_A_306_277#_c_802_n 0.00478301f $X=7.21 $Y=2.865 $X2=0
+ $Y2=0
cc_514 N_RESET_B_c_608_n N_A_306_277#_c_802_n 7.0458e-19 $X=7.17 $Y=1.707 $X2=0
+ $Y2=0
cc_515 N_RESET_B_M1000_g N_A_306_277#_c_895_n 0.00439379f $X=7.21 $Y=2.865 $X2=0
+ $Y2=0
cc_516 N_RESET_B_M1000_g N_A_306_277#_c_803_n 6.50273e-19 $X=7.21 $Y=2.865 $X2=0
+ $Y2=0
cc_517 N_RESET_B_M1022_g N_A_306_277#_c_807_n 0.00230604f $X=3.29 $Y=2.525 $X2=0
+ $Y2=0
cc_518 N_RESET_B_c_578_n N_A_306_277#_c_808_n 0.00353542f $X=6.815 $Y=1.665
+ $X2=0 $Y2=0
cc_519 N_RESET_B_c_578_n N_A_306_277#_c_809_n 0.00167546f $X=6.815 $Y=1.665
+ $X2=0 $Y2=0
cc_520 N_RESET_B_M1022_g N_A_306_277#_c_811_n 0.00667767f $X=3.29 $Y=2.525 $X2=0
+ $Y2=0
cc_521 N_RESET_B_c_578_n N_A_306_277#_c_794_n 0.00885802f $X=6.815 $Y=1.665
+ $X2=0 $Y2=0
cc_522 N_RESET_B_c_578_n N_A_336_463#_M1017_g 0.00585951f $X=6.815 $Y=1.665
+ $X2=0 $Y2=0
cc_523 N_RESET_B_c_576_n N_A_336_463#_c_1048_n 0.0197342f $X=2.495 $Y=1.665
+ $X2=0 $Y2=0
cc_524 N_RESET_B_c_588_n N_A_336_463#_c_1053_n 0.00874783f $X=3.215 $Y=3.15
+ $X2=0 $Y2=0
cc_525 N_RESET_B_M1022_g N_A_336_463#_c_1053_n 0.0204879f $X=3.29 $Y=2.525 $X2=0
+ $Y2=0
cc_526 N_RESET_B_c_596_n N_A_336_463#_c_1053_n 0.00528575f $X=3.205 $Y=2.24
+ $X2=0 $Y2=0
cc_527 N_RESET_B_c_576_n N_A_336_463#_c_1053_n 0.00434742f $X=2.495 $Y=1.665
+ $X2=0 $Y2=0
cc_528 N_RESET_B_c_578_n N_A_336_463#_c_1054_n 0.013022f $X=6.815 $Y=1.665 $X2=0
+ $Y2=0
cc_529 N_RESET_B_c_578_n N_A_336_463#_c_1049_n 0.0206576f $X=6.815 $Y=1.665
+ $X2=0 $Y2=0
cc_530 N_RESET_B_c_588_n N_A_336_463#_c_1056_n 0.00598542f $X=3.215 $Y=3.15
+ $X2=0 $Y2=0
cc_531 N_RESET_B_c_576_n N_A_336_463#_c_1056_n 0.00503928f $X=2.495 $Y=1.665
+ $X2=0 $Y2=0
cc_532 N_RESET_B_c_578_n N_A_336_463#_c_1050_n 0.00477965f $X=6.815 $Y=1.665
+ $X2=0 $Y2=0
cc_533 N_RESET_B_M1000_g N_A_1287_276#_M1027_g 0.0205381f $X=7.21 $Y=2.865 $X2=0
+ $Y2=0
cc_534 N_RESET_B_c_597_n N_A_1287_276#_M1027_g 0.00731858f $X=7.21 $Y=2.085
+ $X2=0 $Y2=0
cc_535 N_RESET_B_c_608_n N_A_1287_276#_M1027_g 0.00117963f $X=7.17 $Y=1.707
+ $X2=0 $Y2=0
cc_536 N_RESET_B_M1019_g N_A_1287_276#_M1013_g 0.022304f $X=7.25 $Y=0.835 $X2=0
+ $Y2=0
cc_537 N_RESET_B_c_578_n N_A_1287_276#_c_1142_n 0.00972765f $X=6.815 $Y=1.665
+ $X2=0 $Y2=0
cc_538 N_RESET_B_c_580_n N_A_1287_276#_c_1142_n 0.00159717f $X=6.96 $Y=1.665
+ $X2=0 $Y2=0
cc_539 N_RESET_B_c_583_n N_A_1287_276#_c_1142_n 0.0105236f $X=7.21 $Y=1.745
+ $X2=0 $Y2=0
cc_540 N_RESET_B_c_584_n N_A_1287_276#_c_1142_n 0.00169221f $X=7.21 $Y=1.745
+ $X2=0 $Y2=0
cc_541 N_RESET_B_c_608_n N_A_1287_276#_c_1142_n 8.68484e-19 $X=7.17 $Y=1.707
+ $X2=0 $Y2=0
cc_542 N_RESET_B_c_597_n N_A_1287_276#_c_1151_n 0.0105236f $X=7.21 $Y=2.085
+ $X2=0 $Y2=0
cc_543 N_RESET_B_M1019_g N_A_1287_276#_c_1152_n 8.90694e-19 $X=7.25 $Y=0.835
+ $X2=0 $Y2=0
cc_544 N_RESET_B_c_597_n N_A_1287_276#_c_1152_n 7.46323e-19 $X=7.21 $Y=2.085
+ $X2=0 $Y2=0
cc_545 N_RESET_B_c_578_n N_A_1287_276#_c_1152_n 0.0171672f $X=6.815 $Y=1.665
+ $X2=0 $Y2=0
cc_546 N_RESET_B_c_580_n N_A_1287_276#_c_1152_n 0.00319427f $X=6.96 $Y=1.665
+ $X2=0 $Y2=0
cc_547 N_RESET_B_c_583_n N_A_1287_276#_c_1152_n 2.59625e-19 $X=7.21 $Y=1.745
+ $X2=0 $Y2=0
cc_548 N_RESET_B_c_584_n N_A_1287_276#_c_1152_n 0.0176502f $X=7.21 $Y=1.745
+ $X2=0 $Y2=0
cc_549 N_RESET_B_c_608_n N_A_1287_276#_c_1152_n 0.00820365f $X=7.17 $Y=1.707
+ $X2=0 $Y2=0
cc_550 N_RESET_B_M1019_g N_A_1287_276#_c_1143_n 0.00629629f $X=7.25 $Y=0.835
+ $X2=0 $Y2=0
cc_551 N_RESET_B_M1019_g N_A_1287_276#_c_1144_n 0.0123938f $X=7.25 $Y=0.835
+ $X2=0 $Y2=0
cc_552 N_RESET_B_c_578_n N_A_1287_276#_c_1144_n 0.00512563f $X=6.815 $Y=1.665
+ $X2=0 $Y2=0
cc_553 N_RESET_B_c_580_n N_A_1287_276#_c_1144_n 0.0090132f $X=6.96 $Y=1.665
+ $X2=0 $Y2=0
cc_554 N_RESET_B_c_583_n N_A_1287_276#_c_1144_n 0.00494356f $X=7.21 $Y=1.745
+ $X2=0 $Y2=0
cc_555 N_RESET_B_c_584_n N_A_1287_276#_c_1144_n 0.0283032f $X=7.21 $Y=1.745
+ $X2=0 $Y2=0
cc_556 N_RESET_B_M1000_g N_A_1287_276#_c_1146_n 0.0064365f $X=7.21 $Y=2.865
+ $X2=0 $Y2=0
cc_557 N_RESET_B_M1019_g N_A_1287_276#_c_1146_n 0.0041958f $X=7.25 $Y=0.835
+ $X2=0 $Y2=0
cc_558 N_RESET_B_c_580_n N_A_1287_276#_c_1146_n 0.00217491f $X=6.96 $Y=1.665
+ $X2=0 $Y2=0
cc_559 N_RESET_B_c_583_n N_A_1287_276#_c_1146_n 0.00619796f $X=7.21 $Y=1.745
+ $X2=0 $Y2=0
cc_560 N_RESET_B_c_584_n N_A_1287_276#_c_1146_n 0.0186457f $X=7.21 $Y=1.745
+ $X2=0 $Y2=0
cc_561 N_RESET_B_c_608_n N_A_1287_276#_c_1146_n 0.0305022f $X=7.17 $Y=1.707
+ $X2=0 $Y2=0
cc_562 N_RESET_B_M1019_g N_A_1287_276#_c_1147_n 0.00115508f $X=7.25 $Y=0.835
+ $X2=0 $Y2=0
cc_563 N_RESET_B_M1019_g N_A_1099_447#_c_1273_n 0.0487111f $X=7.25 $Y=0.835
+ $X2=0 $Y2=0
cc_564 N_RESET_B_M1000_g N_A_1099_447#_M1021_g 0.011565f $X=7.21 $Y=2.865 $X2=0
+ $Y2=0
cc_565 N_RESET_B_M1019_g N_A_1099_447#_M1021_g 0.00497514f $X=7.25 $Y=0.835
+ $X2=0 $Y2=0
cc_566 N_RESET_B_c_583_n N_A_1099_447#_M1021_g 0.0138178f $X=7.21 $Y=1.745 $X2=0
+ $Y2=0
cc_567 N_RESET_B_c_578_n N_A_1099_447#_c_1285_n 0.0184062f $X=6.815 $Y=1.665
+ $X2=0 $Y2=0
cc_568 N_RESET_B_M1019_g N_A_1099_447#_c_1286_n 0.0140302f $X=7.25 $Y=0.835
+ $X2=0 $Y2=0
cc_569 N_RESET_B_c_578_n N_A_1099_447#_c_1286_n 0.00936463f $X=6.815 $Y=1.665
+ $X2=0 $Y2=0
cc_570 N_RESET_B_M1019_g N_A_1099_447#_c_1287_n 0.0079323f $X=7.25 $Y=0.835
+ $X2=0 $Y2=0
cc_571 N_RESET_B_c_578_n N_A_1099_447#_c_1296_n 0.00900975f $X=6.815 $Y=1.665
+ $X2=0 $Y2=0
cc_572 N_RESET_B_c_578_n N_A_1099_447#_c_1290_n 0.0019604f $X=6.815 $Y=1.665
+ $X2=0 $Y2=0
cc_573 N_RESET_B_M1029_g N_A_27_463#_c_1497_n 0.0102793f $X=0.475 $Y=2.525 $X2=0
+ $Y2=0
cc_574 N_RESET_B_c_588_n N_A_27_463#_c_1497_n 0.00855576f $X=3.215 $Y=3.15 $X2=0
+ $Y2=0
cc_575 N_RESET_B_c_595_n N_A_27_463#_c_1497_n 0.00362941f $X=0.515 $Y=2.17 $X2=0
+ $Y2=0
cc_576 N_RESET_B_c_576_n N_A_27_463#_c_1497_n 0.0151832f $X=2.495 $Y=1.665 $X2=0
+ $Y2=0
cc_577 N_RESET_B_c_581_n N_A_27_463#_c_1497_n 5.33861e-19 $X=0.515 $Y=1.65 $X2=0
+ $Y2=0
cc_578 N_RESET_B_c_582_n N_A_27_463#_c_1497_n 0.015695f $X=0.515 $Y=1.65 $X2=0
+ $Y2=0
cc_579 N_RESET_B_M1029_g N_A_27_463#_c_1500_n 5.40796e-19 $X=0.475 $Y=2.525
+ $X2=0 $Y2=0
cc_580 N_RESET_B_c_595_n N_A_27_463#_c_1500_n 5.59306e-19 $X=0.515 $Y=2.17 $X2=0
+ $Y2=0
cc_581 N_RESET_B_M1029_g N_A_27_463#_c_1498_n 0.0109107f $X=0.475 $Y=2.525 $X2=0
+ $Y2=0
cc_582 N_RESET_B_c_595_n N_A_27_463#_c_1498_n 0.00141368f $X=0.515 $Y=2.17 $X2=0
+ $Y2=0
cc_583 N_RESET_B_c_576_n N_A_27_463#_c_1498_n 3.00994e-19 $X=2.495 $Y=1.665
+ $X2=0 $Y2=0
cc_584 N_RESET_B_c_577_n N_A_27_463#_c_1498_n 0.0011655f $X=0.385 $Y=1.665 $X2=0
+ $Y2=0
cc_585 N_RESET_B_c_582_n N_A_27_463#_c_1498_n 0.0308986f $X=0.515 $Y=1.65 $X2=0
+ $Y2=0
cc_586 N_RESET_B_c_576_n N_A_27_463#_c_1502_n 0.00168624f $X=2.495 $Y=1.665
+ $X2=0 $Y2=0
cc_587 N_RESET_B_c_594_n N_A_27_463#_c_1496_n 2.86836e-19 $X=0.515 $Y=2.005
+ $X2=0 $Y2=0
cc_588 N_RESET_B_c_576_n N_A_27_463#_c_1496_n 0.0443763f $X=2.495 $Y=1.665 $X2=0
+ $Y2=0
cc_589 N_RESET_B_c_581_n N_A_27_463#_c_1496_n 2.92583e-19 $X=0.515 $Y=1.65 $X2=0
+ $Y2=0
cc_590 N_RESET_B_c_582_n N_A_27_463#_c_1496_n 0.0165522f $X=0.515 $Y=1.65 $X2=0
+ $Y2=0
cc_591 N_RESET_B_M1029_g N_VPWR_c_1555_n 0.0131885f $X=0.475 $Y=2.525 $X2=0
+ $Y2=0
cc_592 N_RESET_B_c_588_n N_VPWR_c_1555_n 0.0249986f $X=3.215 $Y=3.15 $X2=0 $Y2=0
cc_593 N_RESET_B_c_588_n N_VPWR_c_1556_n 0.0242455f $X=3.215 $Y=3.15 $X2=0 $Y2=0
cc_594 N_RESET_B_M1022_g N_VPWR_c_1556_n 0.0133427f $X=3.29 $Y=2.525 $X2=0 $Y2=0
cc_595 N_RESET_B_c_588_n N_VPWR_c_1557_n 0.00758391f $X=3.215 $Y=3.15 $X2=0
+ $Y2=0
cc_596 N_RESET_B_M1000_g N_VPWR_c_1558_n 0.0033399f $X=7.21 $Y=2.865 $X2=0 $Y2=0
cc_597 N_RESET_B_M1000_g N_VPWR_c_1563_n 0.00346518f $X=7.21 $Y=2.865 $X2=0
+ $Y2=0
cc_598 N_RESET_B_c_588_n N_VPWR_c_1565_n 0.0577631f $X=3.215 $Y=3.15 $X2=0 $Y2=0
cc_599 N_RESET_B_c_588_n N_VPWR_c_1554_n 0.088427f $X=3.215 $Y=3.15 $X2=0 $Y2=0
cc_600 N_RESET_B_c_589_n N_VPWR_c_1554_n 0.00877912f $X=0.55 $Y=3.15 $X2=0 $Y2=0
cc_601 N_RESET_B_M1000_g N_VPWR_c_1554_n 0.00675432f $X=7.21 $Y=2.865 $X2=0
+ $Y2=0
cc_602 N_RESET_B_c_589_n N_VPWR_c_1569_n 0.0085614f $X=0.55 $Y=3.15 $X2=0 $Y2=0
cc_603 N_RESET_B_M1023_g N_VGND_c_1689_n 0.0222634f $X=0.635 $Y=0.815 $X2=0
+ $Y2=0
cc_604 N_RESET_B_M1031_g N_VGND_c_1690_n 0.00159951f $X=3.12 $Y=0.825 $X2=0
+ $Y2=0
cc_605 N_RESET_B_M1019_g N_VGND_c_1691_n 0.0017917f $X=7.25 $Y=0.835 $X2=0 $Y2=0
cc_606 N_RESET_B_M1023_g N_VGND_c_1694_n 0.00396895f $X=0.635 $Y=0.815 $X2=0
+ $Y2=0
cc_607 N_RESET_B_M1019_g N_VGND_c_1696_n 0.00380818f $X=7.25 $Y=0.835 $X2=0
+ $Y2=0
cc_608 N_RESET_B_M1023_g N_VGND_c_1702_n 0.0076824f $X=0.635 $Y=0.815 $X2=0
+ $Y2=0
cc_609 N_RESET_B_M1031_g N_VGND_c_1702_n 9.46663e-19 $X=3.12 $Y=0.825 $X2=0
+ $Y2=0
cc_610 N_RESET_B_M1019_g N_VGND_c_1702_n 0.00424146f $X=7.25 $Y=0.835 $X2=0
+ $Y2=0
cc_611 N_A_306_277#_M1008_g N_A_336_463#_M1017_g 0.0272815f $X=4.31 $Y=2.28
+ $X2=0 $Y2=0
cc_612 N_A_306_277#_c_798_n N_A_336_463#_M1017_g 0.0149263f $X=5.2 $Y=2.71 $X2=0
+ $Y2=0
cc_613 N_A_306_277#_c_807_n N_A_336_463#_M1017_g 9.64506e-19 $X=4.19 $Y=2.71
+ $X2=0 $Y2=0
cc_614 N_A_306_277#_c_851_n N_A_336_463#_M1017_g 0.00324017f $X=5.285 $Y=2.71
+ $X2=0 $Y2=0
cc_615 N_A_306_277#_c_784_n N_A_336_463#_M1028_g 0.016719f $X=4.31 $Y=1.04 $X2=0
+ $Y2=0
cc_616 N_A_306_277#_M1007_g N_A_336_463#_M1028_g 0.0201687f $X=5.61 $Y=0.645
+ $X2=0 $Y2=0
cc_617 N_A_306_277#_M1030_g N_A_336_463#_c_1048_n 0.00647971f $X=1.605 $Y=2.525
+ $X2=0 $Y2=0
cc_618 N_A_306_277#_c_775_n N_A_336_463#_c_1048_n 0.0120987f $X=1.97 $Y=1.46
+ $X2=0 $Y2=0
cc_619 N_A_306_277#_c_777_n N_A_336_463#_c_1048_n 0.00895496f $X=2.115 $Y=1.11
+ $X2=0 $Y2=0
cc_620 N_A_306_277#_M1011_g N_A_336_463#_c_1048_n 5.29542e-19 $X=2.115 $Y=0.825
+ $X2=0 $Y2=0
cc_621 N_A_306_277#_M1008_g N_A_336_463#_c_1053_n 0.00497221f $X=4.31 $Y=2.28
+ $X2=0 $Y2=0
cc_622 N_A_306_277#_c_807_n N_A_336_463#_c_1053_n 0.00523551f $X=4.19 $Y=2.71
+ $X2=0 $Y2=0
cc_623 N_A_306_277#_M1008_g N_A_336_463#_c_1054_n 0.0142751f $X=4.31 $Y=2.28
+ $X2=0 $Y2=0
cc_624 N_A_306_277#_c_798_n N_A_336_463#_c_1054_n 0.0328222f $X=5.2 $Y=2.71
+ $X2=0 $Y2=0
cc_625 N_A_306_277#_c_807_n N_A_336_463#_c_1054_n 0.0219053f $X=4.19 $Y=2.71
+ $X2=0 $Y2=0
cc_626 N_A_306_277#_c_811_n N_A_336_463#_c_1054_n 9.46513e-19 $X=4.31 $Y=2.925
+ $X2=0 $Y2=0
cc_627 N_A_306_277#_M1008_g N_A_336_463#_c_1049_n 0.012326f $X=4.31 $Y=2.28
+ $X2=0 $Y2=0
cc_628 N_A_306_277#_M1030_g N_A_336_463#_c_1056_n 0.00449259f $X=1.605 $Y=2.525
+ $X2=0 $Y2=0
cc_629 N_A_306_277#_c_775_n N_A_336_463#_c_1056_n 0.0019093f $X=1.97 $Y=1.46
+ $X2=0 $Y2=0
cc_630 N_A_306_277#_M1008_g N_A_336_463#_c_1050_n 0.0222836f $X=4.31 $Y=2.28
+ $X2=0 $Y2=0
cc_631 N_A_306_277#_c_802_n N_A_1287_276#_M1000_d 0.0124647f $X=7.805 $Y=2.98
+ $X2=0 $Y2=0
cc_632 N_A_306_277#_M1005_g N_A_1287_276#_M1027_g 0.020896f $X=6.07 $Y=2.865
+ $X2=0 $Y2=0
cc_633 N_A_306_277#_c_850_n N_A_1287_276#_M1027_g 0.00194265f $X=5.92 $Y=2.85
+ $X2=0 $Y2=0
cc_634 N_A_306_277#_c_799_n N_A_1287_276#_M1027_g 0.00347446f $X=6.082 $Y=2.765
+ $X2=0 $Y2=0
cc_635 N_A_306_277#_c_800_n N_A_1287_276#_M1027_g 0.0141649f $X=7.09 $Y=2.515
+ $X2=0 $Y2=0
cc_636 N_A_306_277#_c_801_n N_A_1287_276#_M1027_g 0.00122748f $X=7.175 $Y=2.895
+ $X2=0 $Y2=0
cc_637 N_A_306_277#_c_808_n N_A_1287_276#_M1027_g 0.00129436f $X=6.085 $Y=2.33
+ $X2=0 $Y2=0
cc_638 N_A_306_277#_c_809_n N_A_1287_276#_M1027_g 0.0160183f $X=6.085 $Y=2.33
+ $X2=0 $Y2=0
cc_639 N_A_306_277#_c_794_n N_A_1287_276#_M1027_g 0.00288477f $X=6.047 $Y=2.165
+ $X2=0 $Y2=0
cc_640 N_A_306_277#_c_787_n N_A_1287_276#_M1013_g 0.00261881f $X=5.845 $Y=1.195
+ $X2=0 $Y2=0
cc_641 N_A_306_277#_c_800_n N_A_1287_276#_c_1151_n 0.00542451f $X=7.09 $Y=2.515
+ $X2=0 $Y2=0
cc_642 N_A_306_277#_c_800_n N_A_1287_276#_c_1152_n 0.00675773f $X=7.09 $Y=2.515
+ $X2=0 $Y2=0
cc_643 N_A_306_277#_c_794_n N_A_1287_276#_c_1143_n 0.0151239f $X=6.047 $Y=2.165
+ $X2=0 $Y2=0
cc_644 N_A_306_277#_c_800_n N_A_1287_276#_c_1146_n 0.0115533f $X=7.09 $Y=2.515
+ $X2=0 $Y2=0
cc_645 N_A_306_277#_c_801_n N_A_1287_276#_c_1146_n 0.00756935f $X=7.175 $Y=2.895
+ $X2=0 $Y2=0
cc_646 N_A_306_277#_c_802_n N_A_1287_276#_c_1146_n 0.0128145f $X=7.805 $Y=2.98
+ $X2=0 $Y2=0
cc_647 N_A_306_277#_c_803_n N_A_1287_276#_c_1146_n 0.0104969f $X=7.89 $Y=2.895
+ $X2=0 $Y2=0
cc_648 N_A_306_277#_c_805_n N_A_1287_276#_c_1146_n 0.0133882f $X=7.975 $Y=2.49
+ $X2=0 $Y2=0
cc_649 N_A_306_277#_c_790_n N_A_1287_276#_c_1147_n 0.0190956f $X=8.38 $Y=1.105
+ $X2=0 $Y2=0
cc_650 N_A_306_277#_c_792_n N_A_1287_276#_c_1148_n 0.0126348f $X=8.475 $Y=1.315
+ $X2=0 $Y2=0
cc_651 N_A_306_277#_c_803_n N_CLK_N_M1009_g 5.47663e-19 $X=7.89 $Y=2.895 $X2=0
+ $Y2=0
cc_652 N_A_306_277#_c_804_n N_CLK_N_M1009_g 0.00968684f $X=8.505 $Y=2.49 $X2=0
+ $Y2=0
cc_653 N_A_306_277#_c_793_n N_CLK_N_M1009_g 0.00664828f $X=8.76 $Y=2.405 $X2=0
+ $Y2=0
cc_654 N_A_306_277#_c_810_n N_CLK_N_M1009_g 0.00889698f $X=8.67 $Y=2.57 $X2=0
+ $Y2=0
cc_655 N_A_306_277#_c_791_n N_CLK_N_M1025_g 0.0196452f $X=8.675 $Y=1.315 $X2=0
+ $Y2=0
cc_656 N_A_306_277#_c_793_n N_CLK_N_M1025_g 0.0264162f $X=8.76 $Y=2.405 $X2=0
+ $Y2=0
cc_657 N_A_306_277#_c_804_n CLK_N 0.0388841f $X=8.505 $Y=2.49 $X2=0 $Y2=0
cc_658 N_A_306_277#_c_805_n CLK_N 0.0132842f $X=7.975 $Y=2.49 $X2=0 $Y2=0
cc_659 N_A_306_277#_c_791_n CLK_N 0.00233841f $X=8.675 $Y=1.315 $X2=0 $Y2=0
cc_660 N_A_306_277#_c_792_n CLK_N 0.0222965f $X=8.475 $Y=1.315 $X2=0 $Y2=0
cc_661 N_A_306_277#_c_793_n CLK_N 0.0514981f $X=8.76 $Y=2.405 $X2=0 $Y2=0
cc_662 N_A_306_277#_c_804_n N_CLK_N_c_1237_n 0.00576039f $X=8.505 $Y=2.49 $X2=0
+ $Y2=0
cc_663 N_A_306_277#_c_791_n N_CLK_N_c_1237_n 0.00145146f $X=8.675 $Y=1.315 $X2=0
+ $Y2=0
cc_664 N_A_306_277#_c_792_n N_CLK_N_c_1237_n 0.00714865f $X=8.475 $Y=1.315 $X2=0
+ $Y2=0
cc_665 N_A_306_277#_c_810_n N_CLK_N_c_1237_n 0.00657539f $X=8.67 $Y=2.57 $X2=0
+ $Y2=0
cc_666 N_A_306_277#_c_850_n N_A_1099_447#_M1003_d 0.0116194f $X=5.92 $Y=2.85
+ $X2=0 $Y2=0
cc_667 N_A_306_277#_c_799_n N_A_1099_447#_M1003_d 0.00156338f $X=6.082 $Y=2.765
+ $X2=0 $Y2=0
cc_668 N_A_306_277#_c_801_n N_A_1099_447#_M1021_g 6.3291e-19 $X=7.175 $Y=2.895
+ $X2=0 $Y2=0
cc_669 N_A_306_277#_c_802_n N_A_1099_447#_M1021_g 0.00586912f $X=7.805 $Y=2.98
+ $X2=0 $Y2=0
cc_670 N_A_306_277#_c_803_n N_A_1099_447#_M1021_g 0.00933533f $X=7.89 $Y=2.895
+ $X2=0 $Y2=0
cc_671 N_A_306_277#_c_805_n N_A_1099_447#_M1021_g 0.00795745f $X=7.975 $Y=2.49
+ $X2=0 $Y2=0
cc_672 N_A_306_277#_c_792_n N_A_1099_447#_M1021_g 4.16867e-19 $X=8.475 $Y=1.315
+ $X2=0 $Y2=0
cc_673 N_A_306_277#_c_810_n N_A_1099_447#_M1021_g 2.15264e-19 $X=8.67 $Y=2.57
+ $X2=0 $Y2=0
cc_674 N_A_306_277#_c_790_n N_A_1099_447#_c_1275_n 0.00284459f $X=8.38 $Y=1.105
+ $X2=0 $Y2=0
cc_675 N_A_306_277#_c_791_n N_A_1099_447#_M1024_g 6.18221e-19 $X=8.675 $Y=1.315
+ $X2=0 $Y2=0
cc_676 N_A_306_277#_c_793_n N_A_1099_447#_M1024_g 0.00266576f $X=8.76 $Y=2.405
+ $X2=0 $Y2=0
cc_677 N_A_306_277#_c_810_n N_A_1099_447#_M1024_g 0.00310748f $X=8.67 $Y=2.57
+ $X2=0 $Y2=0
cc_678 N_A_306_277#_c_792_n N_A_1099_447#_c_1282_n 9.20737e-19 $X=8.475 $Y=1.315
+ $X2=0 $Y2=0
cc_679 N_A_306_277#_M1005_g N_A_1099_447#_c_1294_n 2.87704e-19 $X=6.07 $Y=2.865
+ $X2=0 $Y2=0
cc_680 N_A_306_277#_c_850_n N_A_1099_447#_c_1294_n 0.0123568f $X=5.92 $Y=2.85
+ $X2=0 $Y2=0
cc_681 N_A_306_277#_c_808_n N_A_1099_447#_c_1294_n 0.0226192f $X=6.085 $Y=2.33
+ $X2=0 $Y2=0
cc_682 N_A_306_277#_c_794_n N_A_1099_447#_c_1294_n 0.00422533f $X=6.047 $Y=2.165
+ $X2=0 $Y2=0
cc_683 N_A_306_277#_M1007_g N_A_1099_447#_c_1284_n 7.70741e-19 $X=5.61 $Y=0.645
+ $X2=0 $Y2=0
cc_684 N_A_306_277#_c_787_n N_A_1099_447#_c_1285_n 0.0100893f $X=5.845 $Y=1.195
+ $X2=0 $Y2=0
cc_685 N_A_306_277#_c_790_n N_A_1099_447#_c_1289_n 0.00535487f $X=8.38 $Y=1.105
+ $X2=0 $Y2=0
cc_686 N_A_306_277#_c_787_n N_A_1099_447#_c_1296_n 6.95202e-19 $X=5.845 $Y=1.195
+ $X2=0 $Y2=0
cc_687 N_A_306_277#_c_850_n N_A_1099_447#_c_1296_n 0.00321541f $X=5.92 $Y=2.85
+ $X2=0 $Y2=0
cc_688 N_A_306_277#_c_808_n N_A_1099_447#_c_1296_n 0.0205003f $X=6.085 $Y=2.33
+ $X2=0 $Y2=0
cc_689 N_A_306_277#_c_809_n N_A_1099_447#_c_1296_n 0.00512672f $X=6.085 $Y=2.33
+ $X2=0 $Y2=0
cc_690 N_A_306_277#_c_794_n N_A_1099_447#_c_1296_n 0.0148312f $X=6.047 $Y=2.165
+ $X2=0 $Y2=0
cc_691 N_A_306_277#_M1007_g N_A_1099_447#_c_1290_n 6.02377e-19 $X=5.61 $Y=0.645
+ $X2=0 $Y2=0
cc_692 N_A_306_277#_c_790_n N_A_1099_447#_c_1291_n 0.00494201f $X=8.38 $Y=1.105
+ $X2=0 $Y2=0
cc_693 N_A_306_277#_c_793_n N_A_1832_367#_c_1441_n 0.0412248f $X=8.76 $Y=2.405
+ $X2=0 $Y2=0
cc_694 N_A_306_277#_c_810_n N_A_1832_367#_c_1441_n 0.0056714f $X=8.67 $Y=2.57
+ $X2=0 $Y2=0
cc_695 N_A_306_277#_c_791_n N_A_1832_367#_c_1435_n 9.21963e-19 $X=8.675 $Y=1.315
+ $X2=0 $Y2=0
cc_696 N_A_306_277#_c_791_n N_A_1832_367#_c_1438_n 0.00227871f $X=8.675 $Y=1.315
+ $X2=0 $Y2=0
cc_697 N_A_306_277#_c_793_n N_A_1832_367#_c_1438_n 0.0141984f $X=8.76 $Y=2.405
+ $X2=0 $Y2=0
cc_698 N_A_306_277#_M1030_g N_A_27_463#_c_1497_n 0.0064356f $X=1.605 $Y=2.525
+ $X2=0 $Y2=0
cc_699 N_A_306_277#_M1030_g N_A_27_463#_c_1500_n 0.0117036f $X=1.605 $Y=2.525
+ $X2=0 $Y2=0
cc_700 N_A_306_277#_M1030_g N_A_27_463#_c_1495_n 6.14495e-19 $X=1.605 $Y=2.525
+ $X2=0 $Y2=0
cc_701 N_A_306_277#_c_776_n N_A_27_463#_c_1495_n 0.00615898f $X=1.68 $Y=1.46
+ $X2=0 $Y2=0
cc_702 N_A_306_277#_c_777_n N_A_27_463#_c_1495_n 6.45401e-19 $X=2.115 $Y=1.11
+ $X2=0 $Y2=0
cc_703 N_A_306_277#_M1030_g N_A_27_463#_c_1496_n 0.0103692f $X=1.605 $Y=2.525
+ $X2=0 $Y2=0
cc_704 N_A_306_277#_c_798_n N_VPWR_M1008_d 0.00836508f $X=5.2 $Y=2.71 $X2=0
+ $Y2=0
cc_705 N_A_306_277#_c_804_n N_VPWR_M1021_d 0.00528156f $X=8.505 $Y=2.49 $X2=0
+ $Y2=0
cc_706 N_A_306_277#_c_798_n N_VPWR_c_1557_n 0.00383366f $X=5.2 $Y=2.71 $X2=0
+ $Y2=0
cc_707 N_A_306_277#_c_807_n N_VPWR_c_1557_n 0.020339f $X=4.19 $Y=2.71 $X2=0
+ $Y2=0
cc_708 N_A_306_277#_c_811_n N_VPWR_c_1557_n 0.00648328f $X=4.31 $Y=2.925 $X2=0
+ $Y2=0
cc_709 N_A_306_277#_c_800_n N_VPWR_c_1558_n 0.0137841f $X=7.09 $Y=2.515 $X2=0
+ $Y2=0
cc_710 N_A_306_277#_c_802_n N_VPWR_c_1559_n 0.0142358f $X=7.805 $Y=2.98 $X2=0
+ $Y2=0
cc_711 N_A_306_277#_c_803_n N_VPWR_c_1559_n 0.00734609f $X=7.89 $Y=2.895 $X2=0
+ $Y2=0
cc_712 N_A_306_277#_c_804_n N_VPWR_c_1559_n 0.0139492f $X=8.505 $Y=2.49 $X2=0
+ $Y2=0
cc_713 N_A_306_277#_c_810_n N_VPWR_c_1559_n 0.0127835f $X=8.67 $Y=2.57 $X2=0
+ $Y2=0
cc_714 N_A_306_277#_M1005_g N_VPWR_c_1561_n 0.00370648f $X=6.07 $Y=2.865 $X2=0
+ $Y2=0
cc_715 N_A_306_277#_c_798_n N_VPWR_c_1561_n 0.00638684f $X=5.2 $Y=2.71 $X2=0
+ $Y2=0
cc_716 N_A_306_277#_c_850_n N_VPWR_c_1561_n 0.0270354f $X=5.92 $Y=2.85 $X2=0
+ $Y2=0
cc_717 N_A_306_277#_c_800_n N_VPWR_c_1561_n 0.00679452f $X=7.09 $Y=2.515 $X2=0
+ $Y2=0
cc_718 N_A_306_277#_c_851_n N_VPWR_c_1561_n 0.00493724f $X=5.285 $Y=2.71 $X2=0
+ $Y2=0
cc_719 N_A_306_277#_c_800_n N_VPWR_c_1563_n 0.00254515f $X=7.09 $Y=2.515 $X2=0
+ $Y2=0
cc_720 N_A_306_277#_c_802_n N_VPWR_c_1563_n 0.0424499f $X=7.805 $Y=2.98 $X2=0
+ $Y2=0
cc_721 N_A_306_277#_c_895_n N_VPWR_c_1563_n 0.0094633f $X=7.26 $Y=2.98 $X2=0
+ $Y2=0
cc_722 N_A_306_277#_c_804_n N_VPWR_c_1563_n 0.00213323f $X=8.505 $Y=2.49 $X2=0
+ $Y2=0
cc_723 N_A_306_277#_c_804_n N_VPWR_c_1566_n 0.00187826f $X=8.505 $Y=2.49 $X2=0
+ $Y2=0
cc_724 N_A_306_277#_c_810_n N_VPWR_c_1566_n 0.0241323f $X=8.67 $Y=2.57 $X2=0
+ $Y2=0
cc_725 N_A_306_277#_M1030_g N_VPWR_c_1554_n 9.39239e-19 $X=1.605 $Y=2.525 $X2=0
+ $Y2=0
cc_726 N_A_306_277#_M1005_g N_VPWR_c_1554_n 0.00599025f $X=6.07 $Y=2.865 $X2=0
+ $Y2=0
cc_727 N_A_306_277#_c_798_n N_VPWR_c_1554_n 0.0168824f $X=5.2 $Y=2.71 $X2=0
+ $Y2=0
cc_728 N_A_306_277#_c_850_n N_VPWR_c_1554_n 0.0291602f $X=5.92 $Y=2.85 $X2=0
+ $Y2=0
cc_729 N_A_306_277#_c_800_n N_VPWR_c_1554_n 0.0170891f $X=7.09 $Y=2.515 $X2=0
+ $Y2=0
cc_730 N_A_306_277#_c_802_n N_VPWR_c_1554_n 0.0268186f $X=7.805 $Y=2.98 $X2=0
+ $Y2=0
cc_731 N_A_306_277#_c_895_n N_VPWR_c_1554_n 0.00598452f $X=7.26 $Y=2.98 $X2=0
+ $Y2=0
cc_732 N_A_306_277#_c_804_n N_VPWR_c_1554_n 0.00897947f $X=8.505 $Y=2.49 $X2=0
+ $Y2=0
cc_733 N_A_306_277#_c_807_n N_VPWR_c_1554_n 0.0110374f $X=4.19 $Y=2.71 $X2=0
+ $Y2=0
cc_734 N_A_306_277#_c_851_n N_VPWR_c_1554_n 0.0057536f $X=5.285 $Y=2.71 $X2=0
+ $Y2=0
cc_735 N_A_306_277#_c_810_n N_VPWR_c_1554_n 0.0130283f $X=8.67 $Y=2.57 $X2=0
+ $Y2=0
cc_736 N_A_306_277#_c_811_n N_VPWR_c_1554_n 0.00826958f $X=4.31 $Y=2.925 $X2=0
+ $Y2=0
cc_737 N_A_306_277#_c_798_n N_VPWR_c_1571_n 0.0241934f $X=5.2 $Y=2.71 $X2=0
+ $Y2=0
cc_738 N_A_306_277#_c_807_n N_VPWR_c_1571_n 0.00791361f $X=4.19 $Y=2.71 $X2=0
+ $Y2=0
cc_739 N_A_306_277#_c_811_n N_VPWR_c_1571_n 0.00168733f $X=4.31 $Y=2.925 $X2=0
+ $Y2=0
cc_740 N_A_306_277#_c_850_n A_1229_531# 0.00297074f $X=5.92 $Y=2.85 $X2=-0.19
+ $Y2=-0.245
cc_741 N_A_306_277#_c_799_n A_1229_531# 0.00150261f $X=6.082 $Y=2.765 $X2=-0.19
+ $Y2=-0.245
cc_742 N_A_306_277#_c_791_n N_VGND_M1025_d 0.00328293f $X=8.675 $Y=1.315 $X2=0
+ $Y2=0
cc_743 N_A_306_277#_c_779_n N_VGND_c_1690_n 0.0236978f $X=3.635 $Y=0.18 $X2=0
+ $Y2=0
cc_744 N_A_306_277#_c_781_n N_VGND_c_1690_n 0.0117106f $X=3.747 $Y=1.04 $X2=0
+ $Y2=0
cc_745 N_A_306_277#_c_791_n N_VGND_c_1692_n 0.0150747f $X=8.675 $Y=1.315 $X2=0
+ $Y2=0
cc_746 N_A_306_277#_c_780_n N_VGND_c_1694_n 0.0299753f $X=2.19 $Y=0.18 $X2=0
+ $Y2=0
cc_747 N_A_306_277#_c_779_n N_VGND_c_1698_n 0.00810586f $X=3.635 $Y=0.18 $X2=0
+ $Y2=0
cc_748 N_A_306_277#_c_784_n N_VGND_c_1698_n 0.00350154f $X=4.31 $Y=1.04 $X2=0
+ $Y2=0
cc_749 N_A_306_277#_M1007_g N_VGND_c_1699_n 0.00302473f $X=5.61 $Y=0.645 $X2=0
+ $Y2=0
cc_750 N_A_306_277#_c_779_n N_VGND_c_1702_n 0.0390385f $X=3.635 $Y=0.18 $X2=0
+ $Y2=0
cc_751 N_A_306_277#_c_780_n N_VGND_c_1702_n 0.0052711f $X=2.19 $Y=0.18 $X2=0
+ $Y2=0
cc_752 N_A_306_277#_c_784_n N_VGND_c_1702_n 0.00492109f $X=4.31 $Y=1.04 $X2=0
+ $Y2=0
cc_753 N_A_306_277#_M1007_g N_VGND_c_1702_n 0.00456544f $X=5.61 $Y=0.645 $X2=0
+ $Y2=0
cc_754 N_A_306_277#_c_779_n N_VGND_c_1703_n 0.00620368f $X=3.635 $Y=0.18 $X2=0
+ $Y2=0
cc_755 N_A_336_463#_c_1048_n N_A_27_463#_c_1500_n 0.0156326f $X=1.89 $Y=0.84
+ $X2=0 $Y2=0
cc_756 N_A_336_463#_c_1056_n N_A_27_463#_c_1500_n 0.0347179f $X=1.887 $Y=2.355
+ $X2=0 $Y2=0
cc_757 N_A_336_463#_c_1048_n N_A_27_463#_c_1495_n 0.0585208f $X=1.89 $Y=0.84
+ $X2=0 $Y2=0
cc_758 N_A_336_463#_c_1053_n N_VPWR_M1015_d 0.00377249f $X=3.33 $Y=2.355 $X2=0
+ $Y2=0
cc_759 N_A_336_463#_c_1054_n N_VPWR_M1008_d 0.0121459f $X=4.675 $Y=2.355 $X2=0
+ $Y2=0
cc_760 N_A_336_463#_c_1049_n N_VPWR_M1008_d 0.00699957f $X=4.76 $Y=1.44 $X2=0
+ $Y2=0
cc_761 N_A_336_463#_c_1053_n N_VPWR_c_1556_n 0.0265229f $X=3.33 $Y=2.355 $X2=0
+ $Y2=0
cc_762 N_A_336_463#_c_1053_n N_VPWR_c_1557_n 0.00584059f $X=3.33 $Y=2.355 $X2=0
+ $Y2=0
cc_763 N_A_336_463#_M1017_g N_VPWR_c_1561_n 0.00393847f $X=4.99 $Y=2.655 $X2=0
+ $Y2=0
cc_764 N_A_336_463#_c_1056_n N_VPWR_c_1565_n 0.00625105f $X=1.887 $Y=2.355 $X2=0
+ $Y2=0
cc_765 N_A_336_463#_M1017_g N_VPWR_c_1554_n 0.00665989f $X=4.99 $Y=2.655 $X2=0
+ $Y2=0
cc_766 N_A_336_463#_c_1053_n N_VPWR_c_1554_n 0.00944361f $X=3.33 $Y=2.355 $X2=0
+ $Y2=0
cc_767 N_A_336_463#_c_1056_n N_VPWR_c_1554_n 0.0082772f $X=1.887 $Y=2.355 $X2=0
+ $Y2=0
cc_768 N_A_336_463#_M1017_g N_VPWR_c_1571_n 0.00765242f $X=4.99 $Y=2.655 $X2=0
+ $Y2=0
cc_769 N_A_336_463#_c_1053_n A_447_463# 0.00496461f $X=3.33 $Y=2.355 $X2=-0.19
+ $Y2=-0.245
cc_770 N_A_336_463#_M1028_g N_VGND_c_1699_n 0.00310277f $X=5.02 $Y=0.645 $X2=0
+ $Y2=0
cc_771 N_A_336_463#_M1028_g N_VGND_c_1702_n 0.00506666f $X=5.02 $Y=0.645 $X2=0
+ $Y2=0
cc_772 N_A_336_463#_M1028_g N_VGND_c_1703_n 0.0050636f $X=5.02 $Y=0.645 $X2=0
+ $Y2=0
cc_773 N_A_1287_276#_c_1148_n N_CLK_N_M1025_g 2.72057e-19 $X=7.727 $Y=1.315
+ $X2=0 $Y2=0
cc_774 N_A_1287_276#_c_1146_n CLK_N 0.051505f $X=7.55 $Y=2.55 $X2=0 $Y2=0
cc_775 N_A_1287_276#_c_1148_n CLK_N 0.0159255f $X=7.727 $Y=1.315 $X2=0 $Y2=0
cc_776 N_A_1287_276#_c_1147_n N_A_1099_447#_c_1273_n 0.00743317f $X=7.825
+ $Y=0.825 $X2=0 $Y2=0
cc_777 N_A_1287_276#_c_1146_n N_A_1099_447#_M1021_g 0.0153793f $X=7.55 $Y=2.55
+ $X2=0 $Y2=0
cc_778 N_A_1287_276#_c_1148_n N_A_1099_447#_M1021_g 0.00637617f $X=7.727
+ $Y=1.315 $X2=0 $Y2=0
cc_779 N_A_1287_276#_c_1147_n N_A_1099_447#_c_1275_n 0.010014f $X=7.825 $Y=0.825
+ $X2=0 $Y2=0
cc_780 N_A_1287_276#_c_1147_n N_A_1099_447#_c_1282_n 0.00792042f $X=7.825
+ $Y=0.825 $X2=0 $Y2=0
cc_781 N_A_1287_276#_c_1148_n N_A_1099_447#_c_1282_n 0.0168207f $X=7.727
+ $Y=1.315 $X2=0 $Y2=0
cc_782 N_A_1287_276#_M1013_g N_A_1099_447#_c_1285_n 0.00166927f $X=6.66 $Y=0.835
+ $X2=0 $Y2=0
cc_783 N_A_1287_276#_c_1152_n N_A_1099_447#_c_1285_n 0.0197434f $X=6.6 $Y=1.545
+ $X2=0 $Y2=0
cc_784 N_A_1287_276#_c_1143_n N_A_1099_447#_c_1285_n 0.00406144f $X=6.6 $Y=1.545
+ $X2=0 $Y2=0
cc_785 N_A_1287_276#_c_1145_n N_A_1099_447#_c_1285_n 0.00868435f $X=6.685
+ $Y=1.315 $X2=0 $Y2=0
cc_786 N_A_1287_276#_M1013_g N_A_1099_447#_c_1286_n 0.0152037f $X=6.66 $Y=0.835
+ $X2=0 $Y2=0
cc_787 N_A_1287_276#_c_1143_n N_A_1099_447#_c_1286_n 0.00330263f $X=6.6 $Y=1.545
+ $X2=0 $Y2=0
cc_788 N_A_1287_276#_c_1144_n N_A_1099_447#_c_1286_n 0.0575868f $X=7.465
+ $Y=1.315 $X2=0 $Y2=0
cc_789 N_A_1287_276#_c_1145_n N_A_1099_447#_c_1286_n 0.0132086f $X=6.685
+ $Y=1.315 $X2=0 $Y2=0
cc_790 N_A_1287_276#_c_1147_n N_A_1099_447#_c_1286_n 0.00743877f $X=7.825
+ $Y=0.825 $X2=0 $Y2=0
cc_791 N_A_1287_276#_c_1148_n N_A_1099_447#_c_1286_n 0.00234244f $X=7.727
+ $Y=1.315 $X2=0 $Y2=0
cc_792 N_A_1287_276#_M1013_g N_A_1099_447#_c_1287_n 8.03334e-19 $X=6.66 $Y=0.835
+ $X2=0 $Y2=0
cc_793 N_A_1287_276#_c_1147_n N_A_1099_447#_c_1289_n 0.0239189f $X=7.825
+ $Y=0.825 $X2=0 $Y2=0
cc_794 N_A_1287_276#_M1027_g N_A_1099_447#_c_1296_n 5.75984e-19 $X=6.61 $Y=2.865
+ $X2=0 $Y2=0
cc_795 N_A_1287_276#_c_1151_n N_A_1099_447#_c_1296_n 0.00138011f $X=6.6 $Y=2.05
+ $X2=0 $Y2=0
cc_796 N_A_1287_276#_c_1152_n N_A_1099_447#_c_1296_n 0.00680369f $X=6.6 $Y=1.545
+ $X2=0 $Y2=0
cc_797 N_A_1287_276#_M1027_g N_VPWR_c_1558_n 0.00305857f $X=6.61 $Y=2.865 $X2=0
+ $Y2=0
cc_798 N_A_1287_276#_M1027_g N_VPWR_c_1561_n 0.00421441f $X=6.61 $Y=2.865 $X2=0
+ $Y2=0
cc_799 N_A_1287_276#_M1027_g N_VPWR_c_1554_n 0.00646169f $X=6.61 $Y=2.865 $X2=0
+ $Y2=0
cc_800 N_A_1287_276#_M1013_g N_VGND_c_1691_n 0.00402018f $X=6.66 $Y=0.835 $X2=0
+ $Y2=0
cc_801 N_A_1287_276#_M1013_g N_VGND_c_1699_n 0.00415323f $X=6.66 $Y=0.835 $X2=0
+ $Y2=0
cc_802 N_A_1287_276#_M1013_g N_VGND_c_1702_n 0.00469432f $X=6.66 $Y=0.835 $X2=0
+ $Y2=0
cc_803 N_CLK_N_M1009_g N_A_1099_447#_M1021_g 0.0170851f $X=8.455 $Y=2.745 $X2=0
+ $Y2=0
cc_804 N_CLK_N_M1025_g N_A_1099_447#_M1021_g 0.00519642f $X=8.595 $Y=1.105 $X2=0
+ $Y2=0
cc_805 CLK_N N_A_1099_447#_M1021_g 0.0214495f $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_806 N_CLK_N_c_1237_n N_A_1099_447#_M1021_g 0.0435206f $X=8.32 $Y=1.71 $X2=0
+ $Y2=0
cc_807 N_CLK_N_M1025_g N_A_1099_447#_c_1275_n 0.0107281f $X=8.595 $Y=1.105 $X2=0
+ $Y2=0
cc_808 N_CLK_N_M1025_g N_A_1099_447#_c_1276_n 0.009099f $X=8.595 $Y=1.105 $X2=0
+ $Y2=0
cc_809 N_CLK_N_M1025_g N_A_1099_447#_c_1279_n 0.00478955f $X=8.595 $Y=1.105
+ $X2=0 $Y2=0
cc_810 CLK_N N_A_1099_447#_c_1282_n 0.00756238f $X=8.315 $Y=1.58 $X2=0 $Y2=0
cc_811 N_CLK_N_c_1237_n N_A_1099_447#_c_1282_n 0.00165136f $X=8.32 $Y=1.71 $X2=0
+ $Y2=0
cc_812 N_CLK_N_M1009_g N_A_1832_367#_c_1441_n 2.05787e-19 $X=8.455 $Y=2.745
+ $X2=0 $Y2=0
cc_813 N_CLK_N_M1009_g N_VPWR_c_1559_n 0.00435904f $X=8.455 $Y=2.745 $X2=0 $Y2=0
cc_814 N_CLK_N_M1009_g N_VPWR_c_1566_n 0.00404714f $X=8.455 $Y=2.745 $X2=0 $Y2=0
cc_815 N_CLK_N_M1009_g N_VPWR_c_1554_n 0.00788322f $X=8.455 $Y=2.745 $X2=0 $Y2=0
cc_816 N_CLK_N_M1025_g N_VGND_c_1692_n 0.0111006f $X=8.595 $Y=1.105 $X2=0 $Y2=0
cc_817 N_A_1099_447#_M1024_g N_A_1832_367#_M1010_g 0.00779624f $X=9.5 $Y=2.155
+ $X2=0 $Y2=0
cc_818 N_A_1099_447#_c_1281_n N_A_1832_367#_M1010_g 0.0146958f $X=9.56 $Y=0.765
+ $X2=0 $Y2=0
cc_819 N_A_1099_447#_M1024_g N_A_1832_367#_M1012_g 0.011655f $X=9.5 $Y=2.155
+ $X2=0 $Y2=0
cc_820 N_A_1099_447#_M1024_g N_A_1832_367#_c_1441_n 0.0131281f $X=9.5 $Y=2.155
+ $X2=0 $Y2=0
cc_821 N_A_1099_447#_c_1277_n N_A_1832_367#_c_1435_n 0.0012466f $X=9.07 $Y=0.765
+ $X2=0 $Y2=0
cc_822 N_A_1099_447#_c_1278_n N_A_1832_367#_c_1435_n 0.00453792f $X=9.425
+ $Y=0.84 $X2=0 $Y2=0
cc_823 N_A_1099_447#_M1024_g N_A_1832_367#_c_1435_n 0.0161997f $X=9.5 $Y=2.155
+ $X2=0 $Y2=0
cc_824 N_A_1099_447#_c_1281_n N_A_1832_367#_c_1435_n 0.00339055f $X=9.56
+ $Y=0.765 $X2=0 $Y2=0
cc_825 N_A_1099_447#_c_1283_n N_A_1832_367#_c_1435_n 0.00285322f $X=9.53 $Y=0.84
+ $X2=0 $Y2=0
cc_826 N_A_1099_447#_M1024_g N_A_1832_367#_c_1436_n 0.00533951f $X=9.5 $Y=2.155
+ $X2=0 $Y2=0
cc_827 N_A_1099_447#_c_1283_n N_A_1832_367#_c_1436_n 0.00202298f $X=9.53 $Y=0.84
+ $X2=0 $Y2=0
cc_828 N_A_1099_447#_M1024_g N_A_1832_367#_c_1437_n 0.0213482f $X=9.5 $Y=2.155
+ $X2=0 $Y2=0
cc_829 N_A_1099_447#_c_1278_n N_A_1832_367#_c_1438_n 0.00461057f $X=9.425
+ $Y=0.84 $X2=0 $Y2=0
cc_830 N_A_1099_447#_c_1279_n N_A_1832_367#_c_1438_n 3.26906e-19 $X=9.145
+ $Y=0.84 $X2=0 $Y2=0
cc_831 N_A_1099_447#_M1024_g N_A_1832_367#_c_1438_n 0.0160158f $X=9.5 $Y=2.155
+ $X2=0 $Y2=0
cc_832 N_A_1099_447#_c_1276_n N_A_1832_367#_c_1439_n 0.00280018f $X=8.995
+ $Y=0.44 $X2=0 $Y2=0
cc_833 N_A_1099_447#_c_1278_n N_A_1832_367#_c_1439_n 0.00574037f $X=9.425
+ $Y=0.84 $X2=0 $Y2=0
cc_834 N_A_1099_447#_c_1281_n N_A_1832_367#_c_1439_n 0.00525535f $X=9.56
+ $Y=0.765 $X2=0 $Y2=0
cc_835 N_A_1099_447#_M1021_g N_VPWR_c_1559_n 7.83384e-19 $X=7.87 $Y=2.635 $X2=0
+ $Y2=0
cc_836 N_A_1099_447#_M1024_g N_VPWR_c_1560_n 0.00549518f $X=9.5 $Y=2.155 $X2=0
+ $Y2=0
cc_837 N_A_1099_447#_M1021_g N_VPWR_c_1563_n 7.63364e-19 $X=7.87 $Y=2.635 $X2=0
+ $Y2=0
cc_838 N_A_1099_447#_M1024_g N_VPWR_c_1566_n 0.00312414f $X=9.5 $Y=2.155 $X2=0
+ $Y2=0
cc_839 N_A_1099_447#_M1024_g N_VPWR_c_1554_n 0.00410284f $X=9.5 $Y=2.155 $X2=0
+ $Y2=0
cc_840 N_A_1099_447#_c_1286_n N_VGND_M1013_d 0.00419776f $X=7.31 $Y=0.97 $X2=0
+ $Y2=0
cc_841 N_A_1099_447#_c_1284_n N_VGND_c_1691_n 0.00208878f $X=6.085 $Y=0.77 $X2=0
+ $Y2=0
cc_842 N_A_1099_447#_c_1286_n N_VGND_c_1691_n 0.0266253f $X=7.31 $Y=0.97 $X2=0
+ $Y2=0
cc_843 N_A_1099_447#_c_1287_n N_VGND_c_1691_n 0.0120194f $X=7.4 $Y=0.88 $X2=0
+ $Y2=0
cc_844 N_A_1099_447#_c_1288_n N_VGND_c_1691_n 0.0183975f $X=7.49 $Y=0.377 $X2=0
+ $Y2=0
cc_845 N_A_1099_447#_c_1275_n N_VGND_c_1692_n 0.00581612f $X=8.105 $Y=1.155
+ $X2=0 $Y2=0
cc_846 N_A_1099_447#_c_1276_n N_VGND_c_1692_n 0.0150361f $X=8.995 $Y=0.44 $X2=0
+ $Y2=0
cc_847 N_A_1099_447#_c_1277_n N_VGND_c_1692_n 0.0076862f $X=9.07 $Y=0.765 $X2=0
+ $Y2=0
cc_848 N_A_1099_447#_c_1278_n N_VGND_c_1692_n 0.00433238f $X=9.425 $Y=0.84 $X2=0
+ $Y2=0
cc_849 N_A_1099_447#_c_1279_n N_VGND_c_1692_n 0.0106481f $X=9.145 $Y=0.84 $X2=0
+ $Y2=0
cc_850 N_A_1099_447#_M1024_g N_VGND_c_1692_n 0.00268626f $X=9.5 $Y=2.155 $X2=0
+ $Y2=0
cc_851 N_A_1099_447#_c_1281_n N_VGND_c_1692_n 0.00239967f $X=9.56 $Y=0.765 $X2=0
+ $Y2=0
cc_852 N_A_1099_447#_c_1289_n N_VGND_c_1692_n 0.00888104f $X=8.195 $Y=0.35 $X2=0
+ $Y2=0
cc_853 N_A_1099_447#_c_1291_n N_VGND_c_1692_n 0.00233438f $X=8.36 $Y=0.35 $X2=0
+ $Y2=0
cc_854 N_A_1099_447#_M1024_g N_VGND_c_1693_n 0.0013257f $X=9.5 $Y=2.155 $X2=0
+ $Y2=0
cc_855 N_A_1099_447#_c_1281_n N_VGND_c_1693_n 0.00915502f $X=9.56 $Y=0.765 $X2=0
+ $Y2=0
cc_856 N_A_1099_447#_c_1276_n N_VGND_c_1696_n 0.0104781f $X=8.995 $Y=0.44 $X2=0
+ $Y2=0
cc_857 N_A_1099_447#_c_1288_n N_VGND_c_1696_n 0.0121364f $X=7.49 $Y=0.377 $X2=0
+ $Y2=0
cc_858 N_A_1099_447#_c_1289_n N_VGND_c_1696_n 0.0527754f $X=8.195 $Y=0.35 $X2=0
+ $Y2=0
cc_859 N_A_1099_447#_c_1291_n N_VGND_c_1696_n 0.00666509f $X=8.36 $Y=0.35 $X2=0
+ $Y2=0
cc_860 N_A_1099_447#_c_1276_n N_VGND_c_1700_n 0.0068107f $X=8.995 $Y=0.44 $X2=0
+ $Y2=0
cc_861 N_A_1099_447#_c_1281_n N_VGND_c_1700_n 0.00481633f $X=9.56 $Y=0.765 $X2=0
+ $Y2=0
cc_862 N_A_1099_447#_c_1276_n N_VGND_c_1702_n 0.0178506f $X=8.995 $Y=0.44 $X2=0
+ $Y2=0
cc_863 N_A_1099_447#_c_1281_n N_VGND_c_1702_n 0.010011f $X=9.56 $Y=0.765 $X2=0
+ $Y2=0
cc_864 N_A_1099_447#_c_1288_n N_VGND_c_1702_n 0.00696477f $X=7.49 $Y=0.377 $X2=0
+ $Y2=0
cc_865 N_A_1099_447#_c_1289_n N_VGND_c_1702_n 0.0312017f $X=8.195 $Y=0.35 $X2=0
+ $Y2=0
cc_866 N_A_1099_447#_c_1291_n N_VGND_c_1702_n 0.0102095f $X=8.36 $Y=0.35 $X2=0
+ $Y2=0
cc_867 N_A_1099_447#_c_1286_n A_1275_125# 0.00368839f $X=7.31 $Y=0.97 $X2=-0.19
+ $Y2=-0.245
cc_868 N_A_1832_367#_M1012_g N_VPWR_c_1560_n 0.00941964f $X=10.085 $Y=2.465
+ $X2=0 $Y2=0
cc_869 N_A_1832_367#_c_1441_n N_VPWR_c_1560_n 0.0250207f $X=9.285 $Y=1.98 $X2=0
+ $Y2=0
cc_870 N_A_1832_367#_c_1436_n N_VPWR_c_1560_n 0.029016f $X=9.95 $Y=1.51 $X2=0
+ $Y2=0
cc_871 N_A_1832_367#_c_1437_n N_VPWR_c_1560_n 0.00433889f $X=9.95 $Y=1.51 $X2=0
+ $Y2=0
cc_872 N_A_1832_367#_M1012_g N_VPWR_c_1567_n 0.00564131f $X=10.085 $Y=2.465
+ $X2=0 $Y2=0
cc_873 N_A_1832_367#_M1012_g N_VPWR_c_1554_n 0.0123412f $X=10.085 $Y=2.465 $X2=0
+ $Y2=0
cc_874 N_A_1832_367#_c_1441_n N_VPWR_c_1554_n 0.0123605f $X=9.285 $Y=1.98 $X2=0
+ $Y2=0
cc_875 N_A_1832_367#_M1010_g Q 0.00171858f $X=10.085 $Y=0.655 $X2=0 $Y2=0
cc_876 N_A_1832_367#_M1010_g Q 0.0229496f $X=10.085 $Y=0.655 $X2=0 $Y2=0
cc_877 N_A_1832_367#_c_1435_n Q 0.00675703f $X=9.47 $Y=1.345 $X2=0 $Y2=0
cc_878 N_A_1832_367#_c_1436_n Q 0.0270645f $X=9.95 $Y=1.51 $X2=0 $Y2=0
cc_879 N_A_1832_367#_M1012_g Q 0.0152416f $X=10.085 $Y=2.465 $X2=0 $Y2=0
cc_880 N_A_1832_367#_M1010_g N_Q_c_1672_n 0.00842648f $X=10.085 $Y=0.655 $X2=0
+ $Y2=0
cc_881 N_A_1832_367#_c_1435_n N_VGND_c_1692_n 0.043208f $X=9.47 $Y=1.345 $X2=0
+ $Y2=0
cc_882 N_A_1832_367#_c_1438_n N_VGND_c_1692_n 0.00810162f $X=9.12 $Y=1.505 $X2=0
+ $Y2=0
cc_883 N_A_1832_367#_c_1439_n N_VGND_c_1692_n 0.0215005f $X=9.47 $Y=0.445 $X2=0
+ $Y2=0
cc_884 N_A_1832_367#_M1010_g N_VGND_c_1693_n 0.00419028f $X=10.085 $Y=0.655
+ $X2=0 $Y2=0
cc_885 N_A_1832_367#_c_1435_n N_VGND_c_1693_n 0.0354001f $X=9.47 $Y=1.345 $X2=0
+ $Y2=0
cc_886 N_A_1832_367#_c_1436_n N_VGND_c_1693_n 0.0163331f $X=9.95 $Y=1.51 $X2=0
+ $Y2=0
cc_887 N_A_1832_367#_c_1437_n N_VGND_c_1693_n 0.0044244f $X=9.95 $Y=1.51 $X2=0
+ $Y2=0
cc_888 N_A_1832_367#_c_1439_n N_VGND_c_1693_n 0.0253698f $X=9.47 $Y=0.445 $X2=0
+ $Y2=0
cc_889 N_A_1832_367#_c_1439_n N_VGND_c_1700_n 0.0198336f $X=9.47 $Y=0.445 $X2=0
+ $Y2=0
cc_890 N_A_1832_367#_M1010_g N_VGND_c_1701_n 0.00579312f $X=10.085 $Y=0.655
+ $X2=0 $Y2=0
cc_891 N_A_1832_367#_M1026_s N_VGND_c_1702_n 0.0021695f $X=9.22 $Y=0.235 $X2=0
+ $Y2=0
cc_892 N_A_1832_367#_M1010_g N_VGND_c_1702_n 0.0115948f $X=10.085 $Y=0.655 $X2=0
+ $Y2=0
cc_893 N_A_1832_367#_c_1439_n N_VGND_c_1702_n 0.0137784f $X=9.47 $Y=0.445 $X2=0
+ $Y2=0
cc_894 N_A_27_463#_c_1497_n N_VPWR_M1029_d 0.00627032f $X=1.16 $Y=2.375
+ $X2=-0.19 $Y2=-0.245
cc_895 N_A_27_463#_c_1497_n N_VPWR_c_1555_n 0.0342813f $X=1.16 $Y=2.375 $X2=0
+ $Y2=0
cc_896 N_A_27_463#_c_1498_n N_VPWR_c_1555_n 0.0082202f $X=0.285 $Y=2.375 $X2=0
+ $Y2=0
cc_897 N_A_27_463#_c_1497_n N_VPWR_c_1565_n 0.00719673f $X=1.16 $Y=2.375 $X2=0
+ $Y2=0
cc_898 N_A_27_463#_c_1497_n N_VPWR_c_1554_n 0.0108756f $X=1.16 $Y=2.375 $X2=0
+ $Y2=0
cc_899 N_A_27_463#_c_1498_n N_VPWR_c_1554_n 0.010934f $X=0.285 $Y=2.375 $X2=0
+ $Y2=0
cc_900 N_A_27_463#_c_1498_n N_VPWR_c_1569_n 0.00692187f $X=0.285 $Y=2.375 $X2=0
+ $Y2=0
cc_901 N_A_27_463#_c_1502_n N_VGND_c_1689_n 0.0102508f $X=1.55 $Y=0.815 $X2=0
+ $Y2=0
cc_902 N_A_27_463#_c_1502_n N_VGND_c_1694_n 0.00565819f $X=1.55 $Y=0.815 $X2=0
+ $Y2=0
cc_903 N_A_27_463#_c_1502_n N_VGND_c_1702_n 0.00963258f $X=1.55 $Y=0.815 $X2=0
+ $Y2=0
cc_904 N_VPWR_c_1554_n N_Q_M1012_d 0.00215158f $X=10.32 $Y=3.33 $X2=0 $Y2=0
cc_905 N_VPWR_c_1567_n Q 0.0210818f $X=10.32 $Y=3.33 $X2=0 $Y2=0
cc_906 N_VPWR_c_1554_n Q 0.0126146f $X=10.32 $Y=3.33 $X2=0 $Y2=0
cc_907 N_Q_c_1672_n N_VGND_c_1693_n 0.0317084f $X=10.3 $Y=0.42 $X2=0 $Y2=0
cc_908 N_Q_c_1672_n N_VGND_c_1701_n 0.0204001f $X=10.3 $Y=0.42 $X2=0 $Y2=0
cc_909 N_Q_M1010_d N_VGND_c_1702_n 0.00215158f $X=10.16 $Y=0.235 $X2=0 $Y2=0
cc_910 N_Q_c_1672_n N_VGND_c_1702_n 0.0122716f $X=10.3 $Y=0.42 $X2=0 $Y2=0
