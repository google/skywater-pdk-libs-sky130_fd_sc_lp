* File: sky130_fd_sc_lp__decapkapwr_3.spice
* Created: Wed Sep  2 09:42:27 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__decapkapwr_3.pex.spice"
.subckt sky130_fd_sc_lp__decapkapwr_3  VNB VPB VGND KAPWR VPWR
* 
* KAPWR	KAPWR
* VGND	VGND
* VPB	VPB
* VNB	VNB
MM1001 N_VGND_M1001_s N_KAPWR_M1001_g N_VGND_M1001_s VNB NSHORT L=0.5 W=0.55
+ AD=0.15675 AS=0.14575 PD=1.67 PS=1.63 NRD=0 NRS=0 M=1 R=1.1 SA=250000
+ SB=250000 A=0.275 P=2.1 MULT=1
MM1000 N_KAPWR_M1000_s N_VGND_M1000_g N_KAPWR_M1000_s VPB PHIGHVT L=0.5 W=1
+ AD=0.285 AS=0.275 PD=2.57 PS=2.55 NRD=0 NRS=1.9503 M=1 R=2 SA=250000 SB=250000
+ A=0.5 P=3 MULT=1
DX2_noxref VNB VPB NWDIODE A=3.3943 P=7.37
*
.include "sky130_fd_sc_lp__decapkapwr_3.pxi.spice"
*
.ends
*
*
