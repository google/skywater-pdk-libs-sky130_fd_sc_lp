# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_lp__invkapwr_8
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.760000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  2.772000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515000 1.210000 5.265000 1.540000 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  2.587200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.175000 0.840000 5.620000 1.040000 ;
        RECT 0.175000 1.040000 0.345000 1.710000 ;
        RECT 0.175000 1.710000 5.620000 1.885000 ;
        RECT 0.635000 1.885000 0.890000 3.045000 ;
        RECT 1.490000 0.395000 1.750000 0.840000 ;
        RECT 1.495000 1.885000 1.750000 3.045000 ;
        RECT 2.350000 0.395000 2.610000 0.840000 ;
        RECT 2.355000 1.885000 2.610000 3.045000 ;
        RECT 3.210000 0.395000 3.470000 0.840000 ;
        RECT 3.215000 1.885000 3.470000 3.045000 ;
        RECT 4.070000 0.395000 4.330000 0.840000 ;
        RECT 4.075000 1.885000 4.330000 3.045000 ;
        RECT 4.930000 1.885000 5.190000 3.045000 ;
        RECT 5.435000 1.040000 5.620000 1.710000 ;
    END
  END Y
  PIN KAPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.070000 2.690000 5.690000 2.945000 ;
    END
  END KAPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 5.760000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.500000 0.500000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.800000 0.500000 3.300000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 5.760000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.760000 0.085000 ;
      RECT 0.000000  3.245000 5.760000 3.415000 ;
      RECT 0.200000  2.055000 0.460000 3.075000 ;
      RECT 1.025000  0.085000 1.320000 0.670000 ;
      RECT 1.060000  2.055000 1.320000 3.075000 ;
      RECT 1.920000  0.085000 2.180000 0.670000 ;
      RECT 1.920000  2.055000 2.180000 3.075000 ;
      RECT 2.780000  0.085000 3.040000 0.670000 ;
      RECT 2.780000  2.055000 3.040000 3.075000 ;
      RECT 3.640000  0.085000 3.900000 0.670000 ;
      RECT 3.640000  2.055000 3.900000 3.075000 ;
      RECT 4.500000  0.085000 4.795000 0.670000 ;
      RECT 4.500000  2.055000 4.760000 3.075000 ;
      RECT 5.360000  2.055000 5.615000 3.075000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.245000  2.725000 0.415000 2.895000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.100000  2.725000 1.270000 2.895000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 1.970000  2.725000 2.140000 2.895000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 2.825000  2.725000 2.995000 2.895000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.690000  2.725000 3.860000 2.895000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.550000  2.725000 4.720000 2.895000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.410000  2.725000 5.580000 2.895000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
  END
END sky130_fd_sc_lp__invkapwr_8
END LIBRARY
