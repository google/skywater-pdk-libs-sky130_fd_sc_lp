* File: sky130_fd_sc_lp__dlrtp_4.pex.spice
* Created: Fri Aug 28 10:27:19 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__DLRTP_4%D 3 5 8 10 11 12 13 14 15 24 26 44
c40 26 0 1.01808e-19 $X=0.697 $Y=0.88
c41 12 0 1.08714e-19 $X=0.635 $Y=0.84
r42 32 44 1.84391 $w=2.48e-07 $l=4e-08 $layer=LI1_cond $X=0.75 $Y=0.965 $X2=0.75
+ $Y2=0.925
r43 24 26 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=0.697 $Y=1.045
+ $X2=0.697 $Y2=0.88
r44 14 15 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=0.75 $Y=1.665
+ $X2=0.75 $Y2=2.035
r45 13 14 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=0.75 $Y=1.295
+ $X2=0.75 $Y2=1.665
r46 12 44 1.06025 $w=2.48e-07 $l=2.3e-08 $layer=LI1_cond $X=0.75 $Y=0.902
+ $X2=0.75 $Y2=0.925
r47 12 13 14.1981 $w=2.48e-07 $l=3.08e-07 $layer=LI1_cond $X=0.75 $Y=0.987
+ $X2=0.75 $Y2=1.295
r48 12 32 1.01415 $w=2.48e-07 $l=2.2e-08 $layer=LI1_cond $X=0.75 $Y=0.987
+ $X2=0.75 $Y2=0.965
r49 12 24 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.72
+ $Y=1.045 $X2=0.72 $Y2=1.045
r50 11 12 12.0942 $w=3.48e-07 $l=2.85e-07 $layer=LI1_cond $X=0.715 $Y=0.555
+ $X2=0.715 $Y2=0.84
r51 8 10 558.915 $w=1.5e-07 $l=1.09e-06 $layer=POLY_cond $X=0.585 $Y=2.64
+ $X2=0.585 $Y2=1.55
r52 5 10 48.4185 $w=3.75e-07 $l=1.87e-07 $layer=POLY_cond $X=0.697 $Y=1.363
+ $X2=0.697 $Y2=1.55
r53 4 24 3.26277 $w=3.75e-07 $l=2.2e-08 $layer=POLY_cond $X=0.697 $Y=1.067
+ $X2=0.697 $Y2=1.045
r54 4 5 43.8991 $w=3.75e-07 $l=2.96e-07 $layer=POLY_cond $X=0.697 $Y=1.067
+ $X2=0.697 $Y2=1.363
r55 3 26 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.585 $Y=0.56
+ $X2=0.585 $Y2=0.88
.ends

.subckt PM_SKY130_FD_SC_LP__DLRTP_4%GATE 1 3 7 9 10 11 12 13 14 20
c48 11 0 1.01808e-19 $X=1.2 $Y=0.925
c49 9 0 1.08714e-19 $X=1.26 $Y=0.88
r50 20 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.26
+ $Y=1.045 $X2=1.26 $Y2=1.045
r51 13 14 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.21 $Y=1.665
+ $X2=1.21 $Y2=2.035
r52 12 13 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.21 $Y=1.295
+ $X2=1.21 $Y2=1.665
r53 12 21 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=1.21 $Y=1.295
+ $X2=1.21 $Y2=1.045
r54 11 21 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=1.21 $Y=0.925
+ $X2=1.21 $Y2=1.045
r55 10 20 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.26 $Y=1.385
+ $X2=1.26 $Y2=1.045
r56 9 20 38.9318 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.26 $Y=0.88
+ $X2=1.26 $Y2=1.045
r57 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.285 $Y=0.56
+ $X2=1.285 $Y2=0.88
r58 1 10 37.5318 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.26 $Y=1.55
+ $X2=1.26 $Y2=1.385
r59 1 3 558.915 $w=1.5e-07 $l=1.09e-06 $layer=POLY_cond $X=1.26 $Y=1.55 $X2=1.26
+ $Y2=2.64
.ends

.subckt PM_SKY130_FD_SC_LP__DLRTP_4%A_267_464# 1 2 7 8 9 11 13 16 20 24 27 29 32
+ 37 38 41 45 53 54 55 57 61 66 67
c159 61 0 3.63245e-19 $X=2.41 $Y=0.93
c160 38 0 1.84641e-19 $X=3.745 $Y=0.74
r161 67 74 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.91 $Y=1.16
+ $X2=3.91 $Y2=1.325
r162 67 73 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.91 $Y=1.16
+ $X2=3.91 $Y2=0.995
r163 66 67 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.91
+ $Y=1.16 $X2=3.91 $Y2=1.16
r164 63 66 3.84148 $w=2.38e-07 $l=8e-08 $layer=LI1_cond $X=3.83 $Y=1.185
+ $X2=3.91 $Y2=1.185
r165 60 61 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.41
+ $Y=0.93 $X2=2.41 $Y2=0.93
r166 57 60 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=2.41 $Y=0.74
+ $X2=2.41 $Y2=0.93
r167 53 56 17.9287 $w=4.18e-07 $l=5e-07 $layer=LI1_cond $X=1.755 $Y=1.655
+ $X2=1.755 $Y2=2.155
r168 53 55 7.50184 $w=4.18e-07 $l=1.2e-07 $layer=LI1_cond $X=1.755 $Y=1.655
+ $X2=1.755 $Y2=1.535
r169 53 54 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.8
+ $Y=1.655 $X2=1.8 $Y2=1.655
r170 43 45 5.44791 $w=2.73e-07 $l=1.3e-07 $layer=LI1_cond $X=1.5 $Y=0.532
+ $X2=1.63 $Y2=0.532
r171 41 63 2.75731 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=3.83 $Y=1.065
+ $X2=3.83 $Y2=1.185
r172 40 41 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=3.83 $Y=0.825
+ $X2=3.83 $Y2=1.065
r173 39 57 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.575 $Y=0.74
+ $X2=2.41 $Y2=0.74
r174 38 40 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.745 $Y=0.74
+ $X2=3.83 $Y2=0.825
r175 38 39 76.3316 $w=1.68e-07 $l=1.17e-06 $layer=LI1_cond $X=3.745 $Y=0.74
+ $X2=2.575 $Y2=0.74
r176 37 48 4.10459 $w=3.63e-07 $l=1.3e-07 $layer=LI1_cond $X=1.63 $Y=2.482
+ $X2=1.5 $Y2=2.482
r177 37 56 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=1.63 $Y=2.3
+ $X2=1.63 $Y2=2.155
r178 34 45 3.55113 $w=1.7e-07 $l=1.38e-07 $layer=LI1_cond $X=1.63 $Y=0.67
+ $X2=1.63 $Y2=0.532
r179 34 55 56.4332 $w=1.68e-07 $l=8.65e-07 $layer=LI1_cond $X=1.63 $Y=0.67
+ $X2=1.63 $Y2=1.535
r180 30 32 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=3.54 $Y=1.54
+ $X2=3.82 $Y2=1.54
r181 28 54 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=1.8 $Y=1.64 $X2=1.8
+ $Y2=1.655
r182 27 32 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.82 $Y=1.465
+ $X2=3.82 $Y2=1.54
r183 27 74 71.7872 $w=1.5e-07 $l=1.4e-07 $layer=POLY_cond $X=3.82 $Y=1.465
+ $X2=3.82 $Y2=1.325
r184 24 73 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=3.82 $Y=0.445
+ $X2=3.82 $Y2=0.995
r185 18 30 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.54 $Y=1.615
+ $X2=3.54 $Y2=1.54
r186 18 20 538.404 $w=1.5e-07 $l=1.05e-06 $layer=POLY_cond $X=3.54 $Y=1.615
+ $X2=3.54 $Y2=2.665
r187 14 29 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.41 $Y=1.64
+ $X2=2.41 $Y2=1.565
r188 14 16 525.585 $w=1.5e-07 $l=1.025e-06 $layer=POLY_cond $X=2.41 $Y=1.64
+ $X2=2.41 $Y2=2.665
r189 13 29 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.41 $Y=1.49
+ $X2=2.41 $Y2=1.565
r190 12 61 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.41 $Y=1.095
+ $X2=2.41 $Y2=0.93
r191 12 13 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=2.41 $Y=1.095
+ $X2=2.41 $Y2=1.49
r192 9 61 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.41 $Y=0.765
+ $X2=2.41 $Y2=0.93
r193 9 11 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.41 $Y=0.765
+ $X2=2.41 $Y2=0.445
r194 8 28 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=1.965 $Y=1.565
+ $X2=1.8 $Y2=1.64
r195 7 29 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.335 $Y=1.565
+ $X2=2.41 $Y2=1.565
r196 7 8 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=2.335 $Y=1.565
+ $X2=1.965 $Y2=1.565
r197 2 48 600 $w=1.7e-07 $l=2.49199e-07 $layer=licon1_PDIFF $count=1 $X=1.335
+ $Y=2.32 $X2=1.5 $Y2=2.5
r198 1 43 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.36
+ $Y=0.35 $X2=1.5 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_LP__DLRTP_4%A_49_70# 1 2 7 11 15 20 24 27 28 29 31 33 35
+ 36 40
c95 40 0 2.08111e-20 $X=2.975 $Y=1.495
c96 36 0 1.45014e-19 $X=2.86 $Y=1.66
c97 7 0 1.67315e-19 $X=2.905 $Y=1.315
r98 36 41 80.7798 $w=5.6e-07 $l=5.05e-07 $layer=POLY_cond $X=2.975 $Y=1.66
+ $X2=2.975 $Y2=2.165
r99 36 40 42.4508 $w=5.6e-07 $l=1.65e-07 $layer=POLY_cond $X=2.975 $Y=1.66
+ $X2=2.975 $Y2=1.495
r100 35 38 17.3773 $w=5.28e-07 $l=5.05e-07 $layer=LI1_cond $X=2.76 $Y=1.66
+ $X2=2.76 $Y2=2.165
r101 35 36 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.86
+ $Y=1.66 $X2=2.86 $Y2=1.66
r102 31 38 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=2.58 $Y=2.905
+ $X2=2.58 $Y2=2.165
r103 28 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.495 $Y=2.99
+ $X2=2.58 $Y2=2.905
r104 28 29 82.2032 $w=1.68e-07 $l=1.26e-06 $layer=LI1_cond $X=2.495 $Y=2.99
+ $X2=1.235 $Y2=2.99
r105 27 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.15 $Y=2.905
+ $X2=1.235 $Y2=2.99
r106 26 27 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=1.15 $Y=2.47
+ $X2=1.15 $Y2=2.905
r107 25 33 2.90867 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=0.475 $Y=2.385
+ $X2=0.34 $Y2=2.385
r108 24 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.065 $Y=2.385
+ $X2=1.15 $Y2=2.47
r109 24 25 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=1.065 $Y=2.385
+ $X2=0.475 $Y2=2.385
r110 18 33 3.58051 $w=2.6e-07 $l=8.9861e-08 $layer=LI1_cond $X=0.33 $Y=2.3
+ $X2=0.34 $Y2=2.385
r111 18 20 80.21 $w=2.48e-07 $l=1.74e-06 $layer=LI1_cond $X=0.33 $Y=2.3 $X2=0.33
+ $Y2=0.56
r112 15 41 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=3.18 $Y=2.665
+ $X2=3.18 $Y2=2.165
r113 11 17 399.957 $w=1.5e-07 $l=7.8e-07 $layer=POLY_cond $X=2.92 $Y=0.445
+ $X2=2.92 $Y2=1.225
r114 7 17 37.1337 $w=1.8e-07 $l=9e-08 $layer=POLY_cond $X=2.905 $Y=1.315
+ $X2=2.905 $Y2=1.225
r115 7 40 69.9677 $w=1.8e-07 $l=1.8e-07 $layer=POLY_cond $X=2.905 $Y=1.315
+ $X2=2.905 $Y2=1.495
r116 2 33 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.245
+ $Y=2.32 $X2=0.37 $Y2=2.465
r117 1 20 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.245
+ $Y=0.35 $X2=0.37 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_LP__DLRTP_4%A_414_47# 1 2 9 13 16 17 19 23 24 25 26 27
+ 28 30 35 36 40 44 46
c132 36 0 2.08111e-20 $X=2.177 $Y=2.405
c133 19 0 2.92934e-20 $X=2.195 $Y=0.39
c134 13 0 2.94792e-19 $X=4.065 $Y=2.555
r135 44 53 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.99 $Y=2.02
+ $X2=3.99 $Y2=2.185
r136 43 46 4.71454 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=3.99 $Y=2.02
+ $X2=4.125 $Y2=2.02
r137 43 44 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.99
+ $Y=2.02 $X2=3.99 $Y2=2.02
r138 40 49 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.37 $Y=1.09
+ $X2=3.37 $Y2=0.925
r139 39 41 8.21986 $w=2.82e-07 $l=1.9e-07 $layer=LI1_cond $X=3.37 $Y=1.09
+ $X2=3.37 $Y2=1.28
r140 39 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.37
+ $Y=1.09 $X2=3.37 $Y2=1.09
r141 35 36 8.1849 $w=2.93e-07 $l=1.65e-07 $layer=LI1_cond $X=2.177 $Y=2.57
+ $X2=2.177 $Y2=2.405
r142 31 33 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=1.98 $Y=1.28
+ $X2=2.235 $Y2=1.28
r143 29 46 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.125 $Y=2.185
+ $X2=4.125 $Y2=2.02
r144 29 30 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=4.125 $Y=2.185
+ $X2=4.125 $Y2=2.885
r145 27 30 6.84389 $w=1.9e-07 $l=1.30767e-07 $layer=LI1_cond $X=4.04 $Y=2.98
+ $X2=4.125 $Y2=2.885
r146 27 28 38.8182 $w=1.88e-07 $l=6.65e-07 $layer=LI1_cond $X=4.04 $Y=2.98
+ $X2=3.375 $Y2=2.98
r147 26 28 6.84389 $w=1.9e-07 $l=1.30767e-07 $layer=LI1_cond $X=3.29 $Y=2.885
+ $X2=3.375 $Y2=2.98
r148 25 41 5.58713 $w=2.82e-07 $l=1.18427e-07 $layer=LI1_cond $X=3.29 $Y=1.365
+ $X2=3.37 $Y2=1.28
r149 25 26 99.1658 $w=1.68e-07 $l=1.52e-06 $layer=LI1_cond $X=3.29 $Y=1.365
+ $X2=3.29 $Y2=2.885
r150 24 33 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=2.325 $Y=1.28
+ $X2=2.235 $Y2=1.28
r151 23 41 3.69812 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.205 $Y=1.28
+ $X2=3.37 $Y2=1.28
r152 23 24 57.4118 $w=1.68e-07 $l=8.8e-07 $layer=LI1_cond $X=3.205 $Y=1.28
+ $X2=2.325 $Y2=1.28
r153 21 33 0.364908 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.235 $Y=1.365
+ $X2=2.235 $Y2=1.28
r154 21 36 64.0808 $w=1.78e-07 $l=1.04e-06 $layer=LI1_cond $X=2.235 $Y=1.365
+ $X2=2.235 $Y2=2.405
r155 17 19 7.20909 $w=1.98e-07 $l=1.3e-07 $layer=LI1_cond $X=2.065 $Y=0.385
+ $X2=2.195 $Y2=0.385
r156 16 31 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.98 $Y=1.195
+ $X2=1.98 $Y2=1.28
r157 15 17 6.87494 $w=2e-07 $l=1.36015e-07 $layer=LI1_cond $X=1.98 $Y=0.485
+ $X2=2.065 $Y2=0.385
r158 15 16 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=1.98 $Y=0.485
+ $X2=1.98 $Y2=1.195
r159 13 53 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=4.065 $Y=2.555
+ $X2=4.065 $Y2=2.185
r160 9 49 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=3.28 $Y=0.445
+ $X2=3.28 $Y2=0.925
r161 2 35 600 $w=1.7e-07 $l=2.80624e-07 $layer=licon1_PDIFF $count=1 $X=2.07
+ $Y=2.345 $X2=2.195 $Y2=2.57
r162 1 19 182 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=1 $X=2.07
+ $Y=0.235 $X2=2.195 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_LP__DLRTP_4%A_857_21# 1 2 7 9 14 16 18 19 21 22 24 25 27
+ 28 30 31 33 34 36 37 39 42 46 47 49 50 53 55 56 59 61 64 66 72 75 76 78 88
c177 75 0 7.97575e-20 $X=5.56 $Y=2.375
c178 53 0 6.44416e-20 $X=5.125 $Y=0.525
c179 50 0 1.8265e-19 $X=4.695 $Y=2.375
c180 46 0 1.65159e-19 $X=4.53 $Y=2.02
c181 19 0 1.05921e-19 $X=6.28 $Y=1.325
r182 88 89 0.607053 $w=3.97e-07 $l=5e-09 $layer=POLY_cond $X=7.565 $Y=1.525
+ $X2=7.57 $Y2=1.525
r183 87 88 51.5995 $w=3.97e-07 $l=4.25e-07 $layer=POLY_cond $X=7.14 $Y=1.525
+ $X2=7.565 $Y2=1.525
r184 86 87 0.607053 $w=3.97e-07 $l=5e-09 $layer=POLY_cond $X=7.135 $Y=1.525
+ $X2=7.14 $Y2=1.525
r185 83 84 0.607053 $w=3.97e-07 $l=5e-09 $layer=POLY_cond $X=6.705 $Y=1.525
+ $X2=6.71 $Y2=1.525
r186 80 81 0.607053 $w=3.97e-07 $l=5e-09 $layer=POLY_cond $X=6.275 $Y=1.525
+ $X2=6.28 $Y2=1.525
r187 73 86 15.1763 $w=3.97e-07 $l=1.25e-07 $layer=POLY_cond $X=7.01 $Y=1.525
+ $X2=7.135 $Y2=1.525
r188 73 84 36.4232 $w=3.97e-07 $l=3e-07 $layer=POLY_cond $X=7.01 $Y=1.525
+ $X2=6.71 $Y2=1.525
r189 72 73 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=7.01
+ $Y=1.49 $X2=7.01 $Y2=1.49
r190 70 83 45.529 $w=3.97e-07 $l=3.75e-07 $layer=POLY_cond $X=6.33 $Y=1.525
+ $X2=6.705 $Y2=1.525
r191 70 81 6.07053 $w=3.97e-07 $l=5e-08 $layer=POLY_cond $X=6.33 $Y=1.525
+ $X2=6.28 $Y2=1.525
r192 69 72 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=6.33 $Y=1.49
+ $X2=7.01 $Y2=1.49
r193 69 70 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=6.33
+ $Y=1.49 $X2=6.33 $Y2=1.49
r194 67 76 1.39518 $w=1.7e-07 $l=8.8e-08 $layer=LI1_cond $X=6.23 $Y=1.49
+ $X2=6.142 $Y2=1.49
r195 67 69 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=6.23 $Y=1.49 $X2=6.33
+ $Y2=1.49
r196 65 76 5.10356 $w=1.72e-07 $l=8.59942e-08 $layer=LI1_cond $X=6.14 $Y=1.575
+ $X2=6.142 $Y2=1.49
r197 65 66 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=6.14 $Y=1.575
+ $X2=6.14 $Y2=2.29
r198 64 76 5.10356 $w=1.72e-07 $l=8.5e-08 $layer=LI1_cond $X=6.142 $Y=1.405
+ $X2=6.142 $Y2=1.49
r199 63 64 23.1325 $w=1.73e-07 $l=3.65e-07 $layer=LI1_cond $X=6.142 $Y=1.04
+ $X2=6.142 $Y2=1.405
r200 62 75 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=5.66 $Y=2.375 $X2=5.56
+ $Y2=2.375
r201 61 66 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.055 $Y=2.375
+ $X2=6.14 $Y2=2.29
r202 61 62 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=6.055 $Y=2.375
+ $X2=5.66 $Y2=2.375
r203 57 75 0.764409 $w=2e-07 $l=8.5e-08 $layer=LI1_cond $X=5.56 $Y=2.46 $X2=5.56
+ $Y2=2.375
r204 57 59 0.277273 $w=1.98e-07 $l=5e-09 $layer=LI1_cond $X=5.56 $Y=2.46
+ $X2=5.56 $Y2=2.465
r205 55 63 6.81835 $w=1.7e-07 $l=1.22327e-07 $layer=LI1_cond $X=6.055 $Y=0.955
+ $X2=6.142 $Y2=1.04
r206 55 56 53.8235 $w=1.68e-07 $l=8.25e-07 $layer=LI1_cond $X=6.055 $Y=0.955
+ $X2=5.23 $Y2=0.955
r207 51 56 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=5.125 $Y=0.87
+ $X2=5.23 $Y2=0.955
r208 51 53 18.2208 $w=2.08e-07 $l=3.45e-07 $layer=LI1_cond $X=5.125 $Y=0.87
+ $X2=5.125 $Y2=0.525
r209 49 75 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=5.46 $Y=2.375 $X2=5.56
+ $Y2=2.375
r210 49 50 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=5.46 $Y=2.375
+ $X2=4.695 $Y2=2.375
r211 47 79 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.53 $Y=2.02
+ $X2=4.53 $Y2=2.185
r212 47 78 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.53 $Y=2.02
+ $X2=4.53 $Y2=1.855
r213 46 47 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.53
+ $Y=2.02 $X2=4.53 $Y2=2.02
r214 44 50 7.64049 $w=1.7e-07 $l=1.95944e-07 $layer=LI1_cond $X=4.537 $Y=2.29
+ $X2=4.695 $Y2=2.375
r215 44 46 9.87808 $w=3.13e-07 $l=2.7e-07 $layer=LI1_cond $X=4.537 $Y=2.29
+ $X2=4.537 $Y2=2.02
r216 40 42 41.0213 $w=1.5e-07 $l=8e-08 $layer=POLY_cond $X=4.36 $Y=0.84 $X2=4.44
+ $Y2=0.84
r217 37 89 25.678 $w=1.5e-07 $l=2e-07 $layer=POLY_cond $X=7.57 $Y=1.325 $X2=7.57
+ $Y2=1.525
r218 37 39 173.52 $w=1.5e-07 $l=5.4e-07 $layer=POLY_cond $X=7.57 $Y=1.325
+ $X2=7.57 $Y2=0.785
r219 34 88 25.678 $w=1.5e-07 $l=2e-07 $layer=POLY_cond $X=7.565 $Y=1.725
+ $X2=7.565 $Y2=1.525
r220 34 36 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=7.565 $Y=1.725
+ $X2=7.565 $Y2=2.465
r221 31 87 25.678 $w=1.5e-07 $l=2e-07 $layer=POLY_cond $X=7.14 $Y=1.325 $X2=7.14
+ $Y2=1.525
r222 31 33 173.52 $w=1.5e-07 $l=5.4e-07 $layer=POLY_cond $X=7.14 $Y=1.325
+ $X2=7.14 $Y2=0.785
r223 28 86 25.678 $w=1.5e-07 $l=2e-07 $layer=POLY_cond $X=7.135 $Y=1.725
+ $X2=7.135 $Y2=1.525
r224 28 30 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=7.135 $Y=1.725
+ $X2=7.135 $Y2=2.465
r225 25 84 25.678 $w=1.5e-07 $l=2e-07 $layer=POLY_cond $X=6.71 $Y=1.325 $X2=6.71
+ $Y2=1.525
r226 25 27 173.52 $w=1.5e-07 $l=5.4e-07 $layer=POLY_cond $X=6.71 $Y=1.325
+ $X2=6.71 $Y2=0.785
r227 22 83 25.678 $w=1.5e-07 $l=2e-07 $layer=POLY_cond $X=6.705 $Y=1.725
+ $X2=6.705 $Y2=1.525
r228 22 24 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=6.705 $Y=1.725
+ $X2=6.705 $Y2=2.465
r229 19 81 25.678 $w=1.5e-07 $l=2e-07 $layer=POLY_cond $X=6.28 $Y=1.325 $X2=6.28
+ $Y2=1.525
r230 19 21 173.52 $w=1.5e-07 $l=5.4e-07 $layer=POLY_cond $X=6.28 $Y=1.325
+ $X2=6.28 $Y2=0.785
r231 16 80 25.678 $w=1.5e-07 $l=2e-07 $layer=POLY_cond $X=6.275 $Y=1.725
+ $X2=6.275 $Y2=1.525
r232 16 18 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=6.275 $Y=1.725
+ $X2=6.275 $Y2=2.465
r233 14 79 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=4.44 $Y=2.555
+ $X2=4.44 $Y2=2.185
r234 10 42 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.44 $Y=0.915
+ $X2=4.44 $Y2=0.84
r235 10 78 482 $w=1.5e-07 $l=9.4e-07 $layer=POLY_cond $X=4.44 $Y=0.915 $X2=4.44
+ $Y2=1.855
r236 7 40 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.36 $Y=0.765
+ $X2=4.36 $Y2=0.84
r237 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=4.36 $Y=0.765
+ $X2=4.36 $Y2=0.445
r238 2 59 300 $w=1.7e-07 $l=6.96491e-07 $layer=licon1_PDIFF $count=2 $X=5.415
+ $Y=1.835 $X2=5.555 $Y2=2.465
r239 1 53 91 $w=1.7e-07 $l=2.13542e-07 $layer=licon1_NDIFF $count=2 $X=5
+ $Y=0.365 $X2=5.125 $Y2=0.525
.ends

.subckt PM_SKY130_FD_SC_LP__DLRTP_4%A_671_47# 1 2 8 9 10 11 13 15 16 18 19 24 25
+ 26 28 30 33 34 39 43 45
c115 26 0 1.27688e-19 $X=3.725 $Y=1.56
c116 24 0 1.83205e-19 $X=3.64 $Y=2.385
c117 13 0 6.44416e-20 $X=5.34 $Y=0.255
r118 41 43 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=4.175 $Y=0.81
+ $X2=4.34 $Y2=0.81
r119 36 39 4.01609 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=3.64 $Y=2.55
+ $X2=3.755 $Y2=2.55
r120 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.89
+ $Y=1.48 $X2=4.89 $Y2=1.48
r121 31 45 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.425 $Y=1.48
+ $X2=4.34 $Y2=1.48
r122 31 33 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=4.425 $Y=1.48
+ $X2=4.89 $Y2=1.48
r123 30 45 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.34 $Y=1.315
+ $X2=4.34 $Y2=1.48
r124 29 43 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.34 $Y=0.895
+ $X2=4.34 $Y2=0.81
r125 29 30 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=4.34 $Y=0.895
+ $X2=4.34 $Y2=1.315
r126 28 41 0.364908 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=4.175 $Y=0.725
+ $X2=4.175 $Y2=0.81
r127 27 28 14.7879 $w=1.78e-07 $l=2.4e-07 $layer=LI1_cond $X=4.175 $Y=0.485
+ $X2=4.175 $Y2=0.725
r128 25 45 3.70735 $w=2.5e-07 $l=1.18427e-07 $layer=LI1_cond $X=4.255 $Y=1.56
+ $X2=4.34 $Y2=1.48
r129 25 26 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=4.255 $Y=1.56
+ $X2=3.725 $Y2=1.56
r130 24 36 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.64 $Y=2.385
+ $X2=3.64 $Y2=2.55
r131 23 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.64 $Y=1.645
+ $X2=3.725 $Y2=1.56
r132 23 24 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=3.64 $Y=1.645
+ $X2=3.64 $Y2=2.385
r133 19 27 6.90553 $w=2.2e-07 $l=1.48324e-07 $layer=LI1_cond $X=4.085 $Y=0.375
+ $X2=4.175 $Y2=0.485
r134 19 21 25.1442 $w=2.18e-07 $l=4.8e-07 $layer=LI1_cond $X=4.085 $Y=0.375
+ $X2=3.605 $Y2=0.375
r135 16 18 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=5.34 $Y=1.725
+ $X2=5.34 $Y2=2.465
r136 13 15 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=5.34 $Y=0.255
+ $X2=5.34 $Y2=0.785
r137 12 34 27.8707 $w=2.94e-07 $l=2.38642e-07 $layer=POLY_cond $X=5.055 $Y=1.65
+ $X2=4.89 $Y2=1.48
r138 11 16 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.265 $Y=1.65
+ $X2=5.34 $Y2=1.725
r139 11 12 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=5.265 $Y=1.65
+ $X2=5.055 $Y2=1.65
r140 9 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.265 $Y=0.18
+ $X2=5.34 $Y2=0.255
r141 9 10 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=5.265 $Y=0.18
+ $X2=4.925 $Y2=0.18
r142 8 34 38.5845 $w=2.94e-07 $l=1.83916e-07 $layer=POLY_cond $X=4.85 $Y=1.315
+ $X2=4.89 $Y2=1.48
r143 7 10 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.85 $Y=0.255
+ $X2=4.925 $Y2=0.18
r144 7 8 543.532 $w=1.5e-07 $l=1.06e-06 $layer=POLY_cond $X=4.85 $Y=0.255
+ $X2=4.85 $Y2=1.315
r145 2 39 600 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=1 $X=3.615
+ $Y=2.345 $X2=3.755 $Y2=2.55
r146 1 21 182 $w=1.7e-07 $l=3.10242e-07 $layer=licon1_NDIFF $count=1 $X=3.355
+ $Y=0.235 $X2=3.605 $Y2=0.37
.ends

.subckt PM_SKY130_FD_SC_LP__DLRTP_4%RESET_B 3 7 8 9 10 15 17
c49 15 0 7.97575e-20 $X=5.79 $Y=1.48
c50 8 0 1.05921e-19 $X=5.52 $Y=1.295
r51 15 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.79 $Y=1.48
+ $X2=5.79 $Y2=1.645
r52 15 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.79 $Y=1.48
+ $X2=5.79 $Y2=1.315
r53 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.79
+ $Y=1.48 $X2=5.79 $Y2=1.48
r54 9 10 7.76402 $w=5.68e-07 $l=3.7e-07 $layer=LI1_cond $X=5.6 $Y=1.665 $X2=5.6
+ $Y2=2.035
r55 9 16 3.88201 $w=5.68e-07 $l=1.85e-07 $layer=LI1_cond $X=5.6 $Y=1.665 $X2=5.6
+ $Y2=1.48
r56 8 16 3.88201 $w=5.68e-07 $l=1.85e-07 $layer=LI1_cond $X=5.6 $Y=1.295 $X2=5.6
+ $Y2=1.48
r57 7 17 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=5.85 $Y=0.785
+ $X2=5.85 $Y2=1.315
r58 3 18 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=5.77 $Y=2.465
+ $X2=5.77 $Y2=1.645
.ends

.subckt PM_SKY130_FD_SC_LP__DLRTP_4%VPWR 1 2 3 4 5 6 23 27 31 35 39 43 45 50 51
+ 52 61 65 70 75 81 84 87 90 94
r104 93 94 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r105 90 91 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r106 87 88 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r107 84 85 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r108 81 82 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r109 79 94 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=7.92 $Y2=3.33
r110 79 91 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=6.96 $Y2=3.33
r111 78 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r112 76 90 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.085 $Y=3.33
+ $X2=6.92 $Y2=3.33
r113 76 78 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=7.085 $Y=3.33
+ $X2=7.44 $Y2=3.33
r114 75 93 4.55259 $w=1.7e-07 $l=2.72e-07 $layer=LI1_cond $X=7.615 $Y=3.33
+ $X2=7.887 $Y2=3.33
r115 75 78 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=7.615 $Y=3.33
+ $X2=7.44 $Y2=3.33
r116 74 91 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=6.96 $Y2=3.33
r117 74 88 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33 $X2=6
+ $Y2=3.33
r118 73 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r119 71 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.18 $Y=3.33
+ $X2=6.015 $Y2=3.33
r120 71 73 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=6.18 $Y=3.33 $X2=6.48
+ $Y2=3.33
r121 70 90 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.755 $Y=3.33
+ $X2=6.92 $Y2=3.33
r122 70 73 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=6.755 $Y=3.33
+ $X2=6.48 $Y2=3.33
r123 69 88 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33 $X2=6
+ $Y2=3.33
r124 69 85 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=5.04 $Y2=3.33
r125 68 69 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r126 66 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.29 $Y=3.33
+ $X2=5.125 $Y2=3.33
r127 66 68 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=5.29 $Y=3.33
+ $X2=5.52 $Y2=3.33
r128 65 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.85 $Y=3.33
+ $X2=6.015 $Y2=3.33
r129 65 68 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=5.85 $Y=3.33
+ $X2=5.52 $Y2=3.33
r130 63 64 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r131 61 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.96 $Y=3.33
+ $X2=5.125 $Y2=3.33
r132 61 63 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=4.96 $Y=3.33
+ $X2=3.12 $Y2=3.33
r133 60 64 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r134 59 60 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r135 57 60 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r136 57 82 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r137 56 59 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r138 56 57 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r139 54 81 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.895 $Y=3.33
+ $X2=0.77 $Y2=3.33
r140 54 56 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.895 $Y=3.33
+ $X2=1.2 $Y2=3.33
r141 52 85 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=5.04 $Y2=3.33
r142 52 64 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.12 $Y2=3.33
r143 50 59 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=2.835 $Y=3.33
+ $X2=2.64 $Y2=3.33
r144 50 51 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=2.835 $Y=3.33
+ $X2=2.935 $Y2=3.33
r145 49 63 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=3.035 $Y=3.33
+ $X2=3.12 $Y2=3.33
r146 49 51 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=3.035 $Y=3.33
+ $X2=2.935 $Y2=3.33
r147 45 48 27.2396 $w=3.28e-07 $l=7.8e-07 $layer=LI1_cond $X=7.78 $Y=2.17
+ $X2=7.78 $Y2=2.95
r148 43 93 3.21359 $w=3.3e-07 $l=1.43332e-07 $layer=LI1_cond $X=7.78 $Y=3.245
+ $X2=7.887 $Y2=3.33
r149 43 48 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=7.78 $Y=3.245
+ $X2=7.78 $Y2=2.95
r150 39 42 27.2396 $w=3.28e-07 $l=7.8e-07 $layer=LI1_cond $X=6.92 $Y=2.17
+ $X2=6.92 $Y2=2.95
r151 37 90 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.92 $Y=3.245
+ $X2=6.92 $Y2=3.33
r152 37 42 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=6.92 $Y=3.245
+ $X2=6.92 $Y2=2.95
r153 33 87 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.015 $Y=3.245
+ $X2=6.015 $Y2=3.33
r154 33 35 17.112 $w=3.28e-07 $l=4.9e-07 $layer=LI1_cond $X=6.015 $Y=3.245
+ $X2=6.015 $Y2=2.755
r155 29 84 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.125 $Y=3.245
+ $X2=5.125 $Y2=3.33
r156 29 31 17.112 $w=3.28e-07 $l=4.9e-07 $layer=LI1_cond $X=5.125 $Y=3.245
+ $X2=5.125 $Y2=2.755
r157 25 51 0.764409 $w=2e-07 $l=8.5e-08 $layer=LI1_cond $X=2.935 $Y=3.245
+ $X2=2.935 $Y2=3.33
r158 25 27 41.3136 $w=1.98e-07 $l=7.45e-07 $layer=LI1_cond $X=2.935 $Y=3.245
+ $X2=2.935 $Y2=2.5
r159 21 81 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.77 $Y=3.245
+ $X2=0.77 $Y2=3.33
r160 21 23 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=0.77 $Y=3.245
+ $X2=0.77 $Y2=2.815
r161 6 48 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=7.64
+ $Y=1.835 $X2=7.78 $Y2=2.95
r162 6 45 400 $w=1.7e-07 $l=3.98905e-07 $layer=licon1_PDIFF $count=1 $X=7.64
+ $Y=1.835 $X2=7.78 $Y2=2.17
r163 5 42 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=6.78
+ $Y=1.835 $X2=6.92 $Y2=2.95
r164 5 39 400 $w=1.7e-07 $l=3.98905e-07 $layer=licon1_PDIFF $count=1 $X=6.78
+ $Y=1.835 $X2=6.92 $Y2=2.17
r165 4 35 600 $w=1.7e-07 $l=1.0014e-06 $layer=licon1_PDIFF $count=1 $X=5.845
+ $Y=1.835 $X2=6.015 $Y2=2.755
r166 3 31 600 $w=1.7e-07 $l=7.88797e-07 $layer=licon1_PDIFF $count=1 $X=4.515
+ $Y=2.345 $X2=5.125 $Y2=2.755
r167 2 27 300 $w=1.7e-07 $l=5.1672e-07 $layer=licon1_PDIFF $count=2 $X=2.485
+ $Y=2.345 $X2=2.93 $Y2=2.5
r168 1 23 600 $w=1.7e-07 $l=5.65044e-07 $layer=licon1_PDIFF $count=1 $X=0.66
+ $Y=2.32 $X2=0.81 $Y2=2.815
.ends

.subckt PM_SKY130_FD_SC_LP__DLRTP_4%Q 1 2 3 4 15 21 23 24 25 26 29 33 38 39 47
r62 45 47 0.983078 $w=7.28e-07 $l=6e-08 $layer=LI1_cond $X=7.71 $Y=1.235
+ $X2=7.71 $Y2=1.295
r63 39 45 2.04931 $w=4.77e-07 $l=5.67913e-07 $layer=LI1_cond $X=7.225 $Y=1.055
+ $X2=7.71 $Y2=1.235
r64 39 47 0.196616 $w=7.28e-07 $l=1.2e-08 $layer=LI1_cond $X=7.71 $Y=1.307
+ $X2=7.71 $Y2=1.295
r65 37 39 7.17647 $w=7.28e-07 $l=4.38e-07 $layer=LI1_cond $X=7.71 $Y=1.745
+ $X2=7.71 $Y2=1.307
r66 37 38 2.1225 $w=4.6e-07 $l=1.05119e-07 $layer=LI1_cond $X=7.71 $Y=1.745
+ $X2=7.665 $Y2=1.83
r67 33 35 54.2871 $w=1.88e-07 $l=9.3e-07 $layer=LI1_cond $X=7.35 $Y=1.98
+ $X2=7.35 $Y2=2.91
r68 31 38 2.1225 $w=4.6e-07 $l=3.54965e-07 $layer=LI1_cond $X=7.35 $Y=1.915
+ $X2=7.665 $Y2=1.83
r69 31 33 3.79426 $w=1.88e-07 $l=6.5e-08 $layer=LI1_cond $X=7.35 $Y=1.915
+ $X2=7.35 $Y2=1.98
r70 27 39 2.04931 $w=4.77e-07 $l=1.12e-07 $layer=LI1_cond $X=7.337 $Y=1.055
+ $X2=7.225 $Y2=1.055
r71 27 29 27.9147 $w=2.23e-07 $l=5.45e-07 $layer=LI1_cond $X=7.337 $Y=1.055
+ $X2=7.337 $Y2=0.51
r72 25 39 5.22257 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=7.225 $Y=1.15
+ $X2=7.225 $Y2=1.055
r73 25 26 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=7.225 $Y=1.15
+ $X2=6.625 $Y2=1.15
r74 23 38 5.07913 $w=1.7e-07 $l=4.1e-07 $layer=LI1_cond $X=7.255 $Y=1.83
+ $X2=7.665 $Y2=1.83
r75 23 24 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=7.255 $Y=1.83
+ $X2=6.585 $Y2=1.83
r76 19 26 6.9898 $w=1.7e-07 $l=1.49579e-07 $layer=LI1_cond $X=6.512 $Y=1.065
+ $X2=6.625 $Y2=1.15
r77 19 21 27.9147 $w=2.23e-07 $l=5.45e-07 $layer=LI1_cond $X=6.512 $Y=1.065
+ $X2=6.512 $Y2=0.52
r78 15 17 54.2871 $w=1.88e-07 $l=9.3e-07 $layer=LI1_cond $X=6.49 $Y=1.98
+ $X2=6.49 $Y2=2.91
r79 13 24 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=6.49 $Y=1.915
+ $X2=6.585 $Y2=1.83
r80 13 15 3.79426 $w=1.88e-07 $l=6.5e-08 $layer=LI1_cond $X=6.49 $Y=1.915
+ $X2=6.49 $Y2=1.98
r81 4 35 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=7.21
+ $Y=1.835 $X2=7.35 $Y2=2.91
r82 4 33 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=7.21
+ $Y=1.835 $X2=7.35 $Y2=1.98
r83 3 17 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=6.35
+ $Y=1.835 $X2=6.49 $Y2=2.91
r84 3 15 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=6.35
+ $Y=1.835 $X2=6.49 $Y2=1.98
r85 2 29 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=7.215
+ $Y=0.365 $X2=7.355 $Y2=0.51
r86 1 21 91 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=2 $X=6.355
+ $Y=0.365 $X2=6.495 $Y2=0.52
.ends

.subckt PM_SKY130_FD_SC_LP__DLRTP_4%VGND 1 2 3 4 5 6 21 25 29 33 37 39 41 44 45
+ 46 52 59 67 72 77 83 86 89 92 96
c114 52 0 1.71278e-19 $X=2.54 $Y=0
c115 25 0 1.91967e-19 $X=2.705 $Y=0.375
r116 95 96 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r117 92 93 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r118 89 90 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6 $Y2=0
r119 86 87 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r120 83 84 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r121 81 96 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0 $X2=7.92
+ $Y2=0
r122 81 93 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0 $X2=6.96
+ $Y2=0
r123 80 81 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r124 78 92 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=7.055 $Y=0 $X2=6.925
+ $Y2=0
r125 78 80 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=7.055 $Y=0
+ $X2=7.44 $Y2=0
r126 77 95 4.55841 $w=1.7e-07 $l=2.7e-07 $layer=LI1_cond $X=7.62 $Y=0 $X2=7.89
+ $Y2=0
r127 77 80 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=7.62 $Y=0 $X2=7.44
+ $Y2=0
r128 76 93 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6.96
+ $Y2=0
r129 76 90 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6
+ $Y2=0
r130 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r131 73 89 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.23 $Y=0 $X2=6.065
+ $Y2=0
r132 73 75 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=6.23 $Y=0 $X2=6.48
+ $Y2=0
r133 72 92 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=6.795 $Y=0 $X2=6.925
+ $Y2=0
r134 72 75 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=6.795 $Y=0
+ $X2=6.48 $Y2=0
r135 71 90 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=6
+ $Y2=0
r136 71 87 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=4.56
+ $Y2=0
r137 70 71 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r138 68 86 8.14251 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=4.74 $Y=0 $X2=4.587
+ $Y2=0
r139 68 70 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=4.74 $Y=0 $X2=5.52
+ $Y2=0
r140 67 89 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.9 $Y=0 $X2=6.065
+ $Y2=0
r141 67 70 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=5.9 $Y=0 $X2=5.52
+ $Y2=0
r142 63 84 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.64
+ $Y2=0
r143 62 65 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=3.12 $Y=0 $X2=4.08
+ $Y2=0
r144 62 63 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r145 60 83 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.87 $Y=0 $X2=2.705
+ $Y2=0
r146 60 62 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=2.87 $Y=0 $X2=3.12
+ $Y2=0
r147 59 86 8.14251 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=4.435 $Y=0
+ $X2=4.587 $Y2=0
r148 59 65 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=4.435 $Y=0
+ $X2=4.08 $Y2=0
r149 58 84 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r150 57 58 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r151 55 58 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r152 54 57 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r153 54 55 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r154 52 83 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.54 $Y=0 $X2=2.705
+ $Y2=0
r155 52 57 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=2.54 $Y=0 $X2=2.16
+ $Y2=0
r156 50 55 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r157 49 50 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r158 46 87 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=4.56
+ $Y2=0
r159 46 63 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.12
+ $Y2=0
r160 46 65 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r161 44 49 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.975 $Y=0
+ $X2=0.72 $Y2=0
r162 44 45 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=0.975 $Y=0 $X2=1.07
+ $Y2=0
r163 43 54 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=1.165 $Y=0 $X2=1.2
+ $Y2=0
r164 43 45 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.165 $Y=0 $X2=1.07
+ $Y2=0
r165 39 95 3.20777 $w=3.3e-07 $l=1.41244e-07 $layer=LI1_cond $X=7.785 $Y=0.085
+ $X2=7.89 $Y2=0
r166 39 41 14.8421 $w=3.28e-07 $l=4.25e-07 $layer=LI1_cond $X=7.785 $Y=0.085
+ $X2=7.785 $Y2=0.51
r167 35 92 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=6.925 $Y=0.085
+ $X2=6.925 $Y2=0
r168 35 37 28.5895 $w=2.58e-07 $l=6.45e-07 $layer=LI1_cond $X=6.925 $Y=0.085
+ $X2=6.925 $Y2=0.73
r169 31 89 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.065 $Y=0.085
+ $X2=6.065 $Y2=0
r170 31 33 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=6.065 $Y=0.085
+ $X2=6.065 $Y2=0.58
r171 27 86 0.649941 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=4.587 $Y=0.085
+ $X2=4.587 $Y2=0
r172 27 29 11.5244 $w=3.03e-07 $l=3.05e-07 $layer=LI1_cond $X=4.587 $Y=0.085
+ $X2=4.587 $Y2=0.39
r173 23 83 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.705 $Y=0.085
+ $X2=2.705 $Y2=0
r174 23 25 10.1275 $w=3.28e-07 $l=2.9e-07 $layer=LI1_cond $X=2.705 $Y=0.085
+ $X2=2.705 $Y2=0.375
r175 19 45 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.07 $Y=0.085
+ $X2=1.07 $Y2=0
r176 19 21 24.5167 $w=1.88e-07 $l=4.2e-07 $layer=LI1_cond $X=1.07 $Y=0.085
+ $X2=1.07 $Y2=0.505
r177 6 41 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=7.645
+ $Y=0.365 $X2=7.785 $Y2=0.51
r178 5 37 182 $w=1.7e-07 $l=4.29331e-07 $layer=licon1_NDIFF $count=1 $X=6.785
+ $Y=0.365 $X2=6.925 $Y2=0.73
r179 4 33 182 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_NDIFF $count=1 $X=5.925
+ $Y=0.365 $X2=6.065 $Y2=0.58
r180 3 29 182 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=1 $X=4.435
+ $Y=0.235 $X2=4.575 $Y2=0.39
r181 2 25 182 $w=1.7e-07 $l=2.81425e-07 $layer=licon1_NDIFF $count=1 $X=2.485
+ $Y=0.235 $X2=2.705 $Y2=0.375
r182 1 21 182 $w=1.7e-07 $l=4.813e-07 $layer=licon1_NDIFF $count=1 $X=0.66
+ $Y=0.35 $X2=1.07 $Y2=0.505
.ends

