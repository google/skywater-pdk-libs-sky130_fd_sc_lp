# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_sc_lp__dlrtp_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_lp__dlrtp_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.160000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.625000 0.470000 0.805000 0.840000 ;
        RECT 0.625000 0.840000 0.875000 2.130000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  1.176000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.395000 1.745000 8.075000 1.915000 ;
        RECT 6.395000 1.915000 6.585000 3.075000 ;
        RECT 6.400000 0.355000 6.625000 1.065000 ;
        RECT 6.400000 1.065000 7.495000 1.105000 ;
        RECT 6.400000 1.105000 8.075000 1.235000 ;
        RECT 7.225000 0.345000 7.450000 1.055000 ;
        RECT 7.225000 1.055000 7.495000 1.065000 ;
        RECT 7.255000 1.915000 7.445000 3.075000 ;
        RECT 7.345000 1.235000 8.075000 1.745000 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  0.315000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.315000 1.210000 5.885000 2.120000 ;
    END
  END RESET_B
  PIN GATE
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 1.045000 0.840000 1.375000 2.130000 ;
    END
  END GATE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 8.160000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.000000 0.000000 8.160000 0.245000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.655000 8.350000 3.520000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 8.160000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.160000 0.085000 ;
      RECT 0.000000  3.245000 8.160000 3.415000 ;
      RECT 0.205000  0.395000 0.455000 2.300000 ;
      RECT 0.205000  2.300000 1.235000 2.470000 ;
      RECT 0.205000  2.470000 0.475000 2.970000 ;
      RECT 0.645000  2.640000 0.895000 3.245000 ;
      RECT 0.975000  0.085000 1.165000 0.670000 ;
      RECT 1.065000  2.470000 1.235000 2.905000 ;
      RECT 1.065000  2.905000 2.665000 3.075000 ;
      RECT 1.335000  0.395000 1.715000 0.670000 ;
      RECT 1.405000  2.300000 1.715000 2.665000 ;
      RECT 1.545000  0.670000 1.715000 1.535000 ;
      RECT 1.545000  1.535000 1.965000 2.155000 ;
      RECT 1.545000  2.155000 1.715000 2.300000 ;
      RECT 1.895000  0.285000 2.360000 0.485000 ;
      RECT 1.895000  0.485000 2.065000 1.195000 ;
      RECT 1.895000  1.195000 3.535000 1.255000 ;
      RECT 1.895000  1.255000 3.375000 1.365000 ;
      RECT 2.030000  2.405000 2.325000 2.735000 ;
      RECT 2.145000  1.365000 2.325000 2.405000 ;
      RECT 2.245000  0.655000 3.915000 0.825000 ;
      RECT 2.245000  0.825000 2.575000 1.025000 ;
      RECT 2.495000  1.535000 3.025000 2.165000 ;
      RECT 2.495000  2.165000 2.665000 2.905000 ;
      RECT 2.540000  0.085000 2.870000 0.485000 ;
      RECT 2.835000  2.335000 3.035000 3.245000 ;
      RECT 3.205000  0.995000 3.535000 1.195000 ;
      RECT 3.205000  1.365000 3.375000 2.885000 ;
      RECT 3.205000  2.885000 4.210000 3.075000 ;
      RECT 3.440000  0.265000 4.265000 0.485000 ;
      RECT 3.555000  1.475000 5.055000 1.645000 ;
      RECT 3.555000  1.645000 3.725000 2.385000 ;
      RECT 3.555000  2.385000 3.870000 2.715000 ;
      RECT 3.745000  0.825000 3.915000 1.065000 ;
      RECT 3.745000  1.065000 4.075000 1.305000 ;
      RECT 3.895000  1.855000 4.210000 2.185000 ;
      RECT 4.040000  2.185000 4.210000 2.885000 ;
      RECT 4.085000  0.485000 4.265000 0.725000 ;
      RECT 4.085000  0.725000 4.425000 0.895000 ;
      RECT 4.255000  0.895000 4.425000 1.315000 ;
      RECT 4.255000  1.315000 5.055000 1.475000 ;
      RECT 4.380000  1.855000 4.695000 2.290000 ;
      RECT 4.380000  2.290000 6.225000 2.460000 ;
      RECT 4.435000  0.085000 4.740000 0.555000 ;
      RECT 4.960000  2.630000 5.290000 3.245000 ;
      RECT 5.020000  0.360000 5.230000 0.870000 ;
      RECT 5.020000  0.870000 6.230000 1.040000 ;
      RECT 5.460000  2.460000 5.660000 3.075000 ;
      RECT 5.850000  2.630000 6.180000 3.245000 ;
      RECT 5.900000  0.085000 6.230000 0.700000 ;
      RECT 6.055000  1.040000 6.230000 1.405000 ;
      RECT 6.055000  1.405000 7.175000 1.575000 ;
      RECT 6.055000  1.575000 6.225000 2.290000 ;
      RECT 6.755000  2.085000 7.085000 3.245000 ;
      RECT 6.795000  0.085000 7.055000 0.895000 ;
      RECT 7.615000  2.085000 7.945000 3.245000 ;
      RECT 7.620000  0.085000 7.950000 0.935000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
  END
END sky130_fd_sc_lp__dlrtp_4
END LIBRARY
