* File: sky130_fd_sc_lp__mux4_0.spice
* Created: Fri Aug 28 10:45:49 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__mux4_0.pex.spice"
.subckt sky130_fd_sc_lp__mux4_0  VNB VPB A2 S0 A3 A1 A0 S1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* S1	S1
* A0	A0
* A1	A1
* A3	A3
* S0	S0
* A2	A2
* VPB	VPB
* VNB	VNB
MM1014 N_VGND_M1014_d N_S0_M1014_g N_A_31_506#_M1014_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75003.6
+ A=0.063 P=1.14 MULT=1
MM1015 A_270_119# N_A2_M1015_g N_VGND_M1014_d VNB NSHORT L=0.15 W=0.42 AD=0.0441
+ AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.6 SB=75003.2
+ A=0.063 P=1.14 MULT=1
MM1009 N_A_294_506#_M1009_d N_A_31_506#_M1009_g A_270_119# VNB NSHORT L=0.15
+ W=0.42 AD=0.0735 AS=0.0441 PD=0.77 PS=0.63 NRD=19.992 NRS=14.28 M=1 R=2.8
+ SA=75001 SB=75002.8 A=0.063 P=1.14 MULT=1
MM1007 A_442_119# N_S0_M1007_g N_A_294_506#_M1009_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0735 PD=0.63 PS=0.77 NRD=14.28 NRS=0 M=1 R=2.8 SA=75001.5
+ SB=75002.3 A=0.063 P=1.14 MULT=1
MM1002 N_VGND_M1002_d N_A3_M1002_g A_442_119# VNB NSHORT L=0.15 W=0.42 AD=0.1029
+ AS=0.0441 PD=0.91 PS=0.63 NRD=31.428 NRS=14.28 M=1 R=2.8 SA=75001.8 SB=75002
+ A=0.063 P=1.14 MULT=1
MM1005 A_642_119# N_A1_M1005_g N_VGND_M1002_d VNB NSHORT L=0.15 W=0.42 AD=0.0441
+ AS=0.1029 PD=0.63 PS=0.91 NRD=14.28 NRS=28.56 M=1 R=2.8 SA=75002.5 SB=75001.3
+ A=0.063 P=1.14 MULT=1
MM1001 N_A_685_504#_M1001_d N_S0_M1001_g A_642_119# VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75002.8
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1003 A_800_119# N_A_31_506#_M1003_g N_A_685_504#_M1001_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75003.3
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1024 N_VGND_M1024_d N_A0_M1024_g A_800_119# VNB NSHORT L=0.15 W=0.42 AD=0.1113
+ AS=0.0441 PD=1.37 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75003.6 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1016 N_A_1075_493#_M1016_d N_A_1029_37#_M1016_g N_A_685_504#_M1016_s VNB
+ NSHORT L=0.15 W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1006 N_A_294_506#_M1006_d N_S1_M1006_g N_A_1075_493#_M1016_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1021 N_VGND_M1021_d N_S1_M1021_g N_A_1029_37#_M1021_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1008 N_X_M1008_d N_A_1075_493#_M1008_g N_VGND_M1021_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1012 N_VPWR_M1012_d N_S0_M1012_g N_A_31_506#_M1012_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0819 AS=0.1113 PD=0.81 PS=1.37 NRD=32.8202 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75003.9 A=0.063 P=1.14 MULT=1
MM1017 A_222_506# N_A2_M1017_g N_VPWR_M1012_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0441 AS=0.0819 PD=0.63 PS=0.81 NRD=23.443 NRS=18.7544 M=1 R=2.8
+ SA=75000.7 SB=75003.3 A=0.063 P=1.14 MULT=1
MM1020 N_A_294_506#_M1020_d N_S0_M1020_g A_222_506# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.110725 AS=0.0441 PD=0.955 PS=0.63 NRD=53.9386 NRS=23.443 M=1 R=2.8
+ SA=75001.1 SB=75003 A=0.063 P=1.14 MULT=1
MM1004 A_426_504# N_A_31_506#_M1004_g N_A_294_506#_M1020_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0441 AS=0.110725 PD=0.63 PS=0.955 NRD=23.443 NRS=53.9386 M=1 R=2.8
+ SA=75001.7 SB=75002.4 A=0.063 P=1.14 MULT=1
MM1010 N_VPWR_M1010_d N_A3_M1010_g A_426_504# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.08925 AS=0.0441 PD=0.845 PS=0.63 NRD=58.6272 NRS=23.443 M=1 R=2.8
+ SA=75002.1 SB=75002 A=0.063 P=1.14 MULT=1
MM1023 A_613_504# N_A1_M1023_g N_VPWR_M1010_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0441 AS=0.08925 PD=0.63 PS=0.845 NRD=23.443 NRS=9.3772 M=1 R=2.8
+ SA=75002.7 SB=75001.4 A=0.063 P=1.14 MULT=1
MM1025 N_A_685_504#_M1025_d N_A_31_506#_M1025_g A_613_504# VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0819 AS=0.0441 PD=0.81 PS=0.63 NRD=25.7873 NRS=23.443 M=1 R=2.8
+ SA=75003 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1011 A_793_504# N_S0_M1011_g N_A_685_504#_M1025_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0441 AS=0.0819 PD=0.63 PS=0.81 NRD=23.443 NRS=25.7873 M=1 R=2.8
+ SA=75003.6 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1013 N_VPWR_M1013_d N_A0_M1013_g A_793_504# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.1113 AS=0.0441 PD=1.37 PS=0.63 NRD=0 NRS=23.443 M=1 R=2.8 SA=75003.9
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1018 N_A_1075_493#_M1018_d N_S1_M1018_g N_A_685_504#_M1018_s VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1000 N_A_294_506#_M1000_d N_A_1029_37#_M1000_g N_A_1075_493#_M1018_d VPB
+ PHIGHVT L=0.15 W=0.42 AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.6 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1022 N_VPWR_M1022_d N_S1_M1022_g N_A_1029_37#_M1022_s VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0855057 AS=0.1113 PD=0.80434 PS=1.37 NRD=23.443 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1019 N_X_M1019_d N_A_1075_493#_M1019_g N_VPWR_M1022_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1696 AS=0.130294 PD=1.81 PS=1.22566 NRD=0 NRS=14.6174 M=1
+ R=4.26667 SA=75000.5 SB=75000.2 A=0.096 P=1.58 MULT=1
DX26_noxref VNB VPB NWDIODE A=15.0319 P=19.85
c_174 VPB 0 3.3911e-19 $X=0 $Y=3.085
c_1064 A_222_506# 0 9.03317e-20 $X=1.11 $Y=2.53
*
.include "sky130_fd_sc_lp__mux4_0.pxi.spice"
*
.ends
*
*
