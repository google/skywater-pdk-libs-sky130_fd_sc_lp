# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__mux2_lp
  CLASS CORE ;
  FOREIGN sky130_fd_sc_lp__mux2_lp ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.320000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A0
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.040000 1.535000 3.235000 1.865000 ;
    END
  END A0
  PIN A1
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.500000 1.195000 2.730000 1.365000 ;
        RECT 1.500000 1.365000 1.830000 1.780000 ;
        RECT 2.400000 0.965000 2.730000 1.195000 ;
    END
  END A1
  PIN S
    ANTENNAGATEAREA  0.378000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.405000 1.180000 3.735000 1.865000 ;
    END
  END S
  PIN X
    ANTENNADIFFAREA  0.239400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.115000 0.255000 0.445000 0.715000 ;
        RECT 0.115000 0.715000 0.355000 2.615000 ;
        RECT 0.115000 2.615000 0.490000 3.075000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.320000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.320000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.320000 0.085000 ;
      RECT 0.000000  3.245000 4.320000 3.415000 ;
      RECT 0.525000  0.885000 2.230000 1.025000 ;
      RECT 0.525000  1.025000 0.855000 1.555000 ;
      RECT 0.660000  1.555000 0.830000 2.375000 ;
      RECT 0.660000  2.375000 2.100000 2.545000 ;
      RECT 0.685000  0.855000 2.230000 0.885000 ;
      RECT 0.905000  0.085000 1.235000 0.685000 ;
      RECT 0.950000  2.715000 1.280000 3.245000 ;
      RECT 1.000000  1.835000 1.330000 2.035000 ;
      RECT 1.000000  2.035000 4.185000 2.205000 ;
      RECT 1.770000  2.545000 2.100000 3.075000 ;
      RECT 1.900000  0.255000 2.230000 0.855000 ;
      RECT 2.590000  2.615000 2.920000 3.245000 ;
      RECT 3.065000  0.085000 3.395000 0.715000 ;
      RECT 3.845000  2.205000 4.185000 3.075000 ;
      RECT 3.855000  0.255000 4.185000 0.715000 ;
      RECT 4.015000  0.715000 4.185000 2.035000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
  END
END sky130_fd_sc_lp__mux2_lp
END LIBRARY
