* File: sky130_fd_sc_lp__a32o_2.spice
* Created: Fri Aug 28 10:01:02 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__a32o_2.pex.spice"
.subckt sky130_fd_sc_lp__a32o_2  VNB VPB B2 B1 A1 A2 A3 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* A3	A3
* A2	A2
* A1	A1
* B1	B1
* B2	B2
* VPB	VPB
* VNB	VNB
MM1001 N_VGND_M1001_d N_A_108_267#_M1001_g N_X_M1001_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75003.6 A=0.126 P=1.98 MULT=1
MM1011 N_VGND_M1011_d N_A_108_267#_M1011_g N_X_M1001_s VNB NSHORT L=0.15 W=0.84
+ AD=0.3108 AS=0.1176 PD=1.58 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75003.2 A=0.126 P=1.98 MULT=1
MM1000 A_432_47# N_B2_M1000_g N_VGND_M1011_d VNB NSHORT L=0.15 W=0.84 AD=0.0882
+ AS=0.3108 PD=1.05 PS=1.58 NRD=7.14 NRS=0 M=1 R=5.6 SA=75001.5 SB=75002.3
+ A=0.126 P=1.98 MULT=1
MM1010 N_A_108_267#_M1010_d N_B1_M1010_g A_432_47# VNB NSHORT L=0.15 W=0.84
+ AD=0.2037 AS=0.0882 PD=1.325 PS=1.05 NRD=10.704 NRS=7.14 M=1 R=5.6 SA=75001.9
+ SB=75002 A=0.126 P=1.98 MULT=1
MM1002 A_631_47# N_A1_M1002_g N_A_108_267#_M1010_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1638 AS=0.2037 PD=1.23 PS=1.325 NRD=19.992 NRS=18.564 M=1 R=5.6
+ SA=75002.5 SB=75001.3 A=0.126 P=1.98 MULT=1
MM1009 A_739_47# N_A2_M1009_g A_631_47# VNB NSHORT L=0.15 W=0.84 AD=0.1638
+ AS=0.1638 PD=1.23 PS=1.23 NRD=19.992 NRS=19.992 M=1 R=5.6 SA=75003 SB=75000.8
+ A=0.126 P=1.98 MULT=1
MM1013 N_VGND_M1013_d N_A3_M1013_g A_739_47# VNB NSHORT L=0.15 W=0.84 AD=0.2646
+ AS=0.1638 PD=2.31 PS=1.23 NRD=7.14 NRS=19.992 M=1 R=5.6 SA=75003.6 SB=75000.2
+ A=0.126 P=1.98 MULT=1
MM1005 N_VPWR_M1005_d N_A_108_267#_M1005_g N_X_M1005_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1006 N_VPWR_M1005_d N_A_108_267#_M1006_g N_X_M1006_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75000.2 A=0.189 P=2.82 MULT=1
MM1008 N_A_108_267#_M1008_d N_B2_M1008_g N_A_345_367#_M1008_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75002.3 A=0.189 P=2.82 MULT=1
MM1003 N_A_345_367#_M1003_d N_B1_M1003_g N_A_108_267#_M1008_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3528 AS=0.1764 PD=1.82 PS=1.54 NRD=29.1757 NRS=0 M=1 R=8.4
+ SA=75000.6 SB=75001.9 A=0.189 P=2.82 MULT=1
MM1007 N_VPWR_M1007_d N_A1_M1007_g N_A_345_367#_M1003_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.23625 AS=0.3528 PD=1.635 PS=1.82 NRD=7.0329 NRS=14.578 M=1 R=8.4
+ SA=75001.3 SB=75001.1 A=0.189 P=2.82 MULT=1
MM1004 N_A_345_367#_M1004_d N_A2_M1004_g N_VPWR_M1007_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.23625 PD=1.54 PS=1.635 NRD=0 NRS=7.8012 M=1 R=8.4
+ SA=75001.9 SB=75000.6 A=0.189 P=2.82 MULT=1
MM1012 N_VPWR_M1012_d N_A3_M1012_g N_A_345_367#_M1004_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.3
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX14_noxref VNB VPB NWDIODE A=9.6607 P=14.09
*
.include "sky130_fd_sc_lp__a32o_2.pxi.spice"
*
.ends
*
*
