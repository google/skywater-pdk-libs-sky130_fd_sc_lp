* File: sky130_fd_sc_lp__ha_4.pxi.spice
* Created: Wed Sep  2 09:54:37 2020
* 
x_PM_SKY130_FD_SC_LP__HA_4%A_110_263# N_A_110_263#_M1005_d N_A_110_263#_M1008_d
+ N_A_110_263#_M1028_d N_A_110_263#_M1015_d N_A_110_263#_M1003_g
+ N_A_110_263#_M1009_g N_A_110_263#_M1014_g N_A_110_263#_M1021_g
+ N_A_110_263#_M1025_g N_A_110_263#_M1022_g N_A_110_263#_M1035_g
+ N_A_110_263#_M1034_g N_A_110_263#_c_197_n N_A_110_263#_c_206_n
+ N_A_110_263#_c_207_n N_A_110_263#_c_222_p N_A_110_263#_c_208_n
+ N_A_110_263#_c_209_n N_A_110_263#_c_198_n N_A_110_263#_c_211_n
+ N_A_110_263#_c_212_n N_A_110_263#_c_225_p N_A_110_263#_c_250_p
+ N_A_110_263#_c_226_p N_A_110_263#_c_292_p N_A_110_263#_c_199_n
+ N_A_110_263#_c_217_p N_A_110_263#_c_200_n N_A_110_263#_c_414_p
+ N_A_110_263#_c_201_n N_A_110_263#_c_229_p PM_SKY130_FD_SC_LP__HA_4%A_110_263#
x_PM_SKY130_FD_SC_LP__HA_4%A_454_263# N_A_454_263#_M1001_d N_A_454_263#_M1000_s
+ N_A_454_263#_M1027_s N_A_454_263#_M1006_g N_A_454_263#_M1016_g
+ N_A_454_263#_M1012_g N_A_454_263#_M1019_g N_A_454_263#_M1023_g
+ N_A_454_263#_M1030_g N_A_454_263#_M1032_g N_A_454_263#_M1033_g
+ N_A_454_263#_M1004_g N_A_454_263#_M1005_g N_A_454_263#_c_437_n
+ N_A_454_263#_M1026_g N_A_454_263#_M1015_g N_A_454_263#_c_440_n
+ N_A_454_263#_c_441_n N_A_454_263#_c_492_n N_A_454_263#_c_442_n
+ N_A_454_263#_c_443_n N_A_454_263#_c_444_n N_A_454_263#_c_494_n
+ N_A_454_263#_c_525_p N_A_454_263#_c_586_p N_A_454_263#_c_526_p
+ N_A_454_263#_c_527_p N_A_454_263#_c_536_p N_A_454_263#_c_495_n
+ N_A_454_263#_c_612_p N_A_454_263#_c_459_n N_A_454_263#_c_496_n
+ N_A_454_263#_c_445_n N_A_454_263#_c_446_n N_A_454_263#_c_447_n
+ N_A_454_263#_c_448_n N_A_454_263#_c_551_p N_A_454_263#_c_461_n
+ N_A_454_263#_c_449_n N_A_454_263#_c_450_n N_A_454_263#_c_451_n
+ PM_SKY130_FD_SC_LP__HA_4%A_454_263#
x_PM_SKY130_FD_SC_LP__HA_4%A N_A_M1020_g N_A_M1000_g N_A_M1031_g N_A_M1017_g
+ N_A_M1013_g N_A_M1011_g N_A_M1024_g N_A_M1018_g N_A_c_699_n N_A_c_700_n
+ N_A_c_713_n N_A_c_714_n N_A_c_701_n A A A N_A_c_717_n N_A_c_703_n N_A_c_704_n
+ N_A_c_705_n A N_A_c_706_n A PM_SKY130_FD_SC_LP__HA_4%A
x_PM_SKY130_FD_SC_LP__HA_4%B N_B_M1001_g N_B_M1007_g N_B_c_867_n N_B_M1002_g
+ N_B_M1027_g N_B_c_870_n N_B_c_871_n N_B_M1010_g N_B_M1008_g N_B_M1028_g
+ N_B_M1029_g N_B_c_874_n N_B_c_875_n N_B_c_876_n N_B_c_877_n N_B_c_878_n
+ N_B_c_879_n N_B_c_880_n B N_B_c_881_n N_B_c_882_n B PM_SKY130_FD_SC_LP__HA_4%B
x_PM_SKY130_FD_SC_LP__HA_4%VPWR N_VPWR_M1003_s N_VPWR_M1014_s N_VPWR_M1035_s
+ N_VPWR_M1012_d N_VPWR_M1032_d N_VPWR_M1007_d N_VPWR_M1017_d N_VPWR_M1013_d
+ N_VPWR_M1004_s N_VPWR_c_1031_n N_VPWR_c_1032_n N_VPWR_c_1033_n N_VPWR_c_1034_n
+ N_VPWR_c_1035_n N_VPWR_c_1036_n N_VPWR_c_1037_n N_VPWR_c_1038_n
+ N_VPWR_c_1074_n N_VPWR_c_1039_n N_VPWR_c_1076_n N_VPWR_c_1040_n
+ N_VPWR_c_1041_n N_VPWR_c_1042_n N_VPWR_c_1043_n N_VPWR_c_1044_n
+ N_VPWR_c_1045_n N_VPWR_c_1046_n N_VPWR_c_1047_n VPWR N_VPWR_c_1048_n
+ N_VPWR_c_1049_n N_VPWR_c_1050_n N_VPWR_c_1051_n N_VPWR_c_1052_n
+ N_VPWR_c_1030_n N_VPWR_c_1054_n N_VPWR_c_1055_n N_VPWR_c_1056_n
+ N_VPWR_c_1057_n PM_SKY130_FD_SC_LP__HA_4%VPWR
x_PM_SKY130_FD_SC_LP__HA_4%SUM N_SUM_M1009_d N_SUM_M1022_d N_SUM_M1003_d
+ N_SUM_M1025_d N_SUM_c_1204_n N_SUM_c_1209_n N_SUM_c_1210_n N_SUM_c_1244_n
+ N_SUM_c_1257_p N_SUM_c_1211_n N_SUM_c_1205_n N_SUM_c_1249_n N_SUM_c_1230_n
+ N_SUM_c_1212_n N_SUM_c_1206_n SUM SUM N_SUM_c_1207_n SUM
+ PM_SKY130_FD_SC_LP__HA_4%SUM
x_PM_SKY130_FD_SC_LP__HA_4%COUT N_COUT_M1016_s N_COUT_M1030_s N_COUT_M1006_s
+ N_COUT_M1023_s N_COUT_c_1264_n N_COUT_c_1274_n N_COUT_c_1265_n N_COUT_c_1268_n
+ N_COUT_c_1316_n N_COUT_c_1278_n N_COUT_c_1266_n N_COUT_c_1269_n COUT COUT COUT
+ PM_SKY130_FD_SC_LP__HA_4%COUT
x_PM_SKY130_FD_SC_LP__HA_4%A_1367_367# N_A_1367_367#_M1008_s
+ N_A_1367_367#_M1018_s N_A_1367_367#_c_1334_n N_A_1367_367#_c_1335_n
+ N_A_1367_367#_c_1337_n PM_SKY130_FD_SC_LP__HA_4%A_1367_367#
x_PM_SKY130_FD_SC_LP__HA_4%VGND N_VGND_M1009_s N_VGND_M1021_s N_VGND_M1034_s
+ N_VGND_M1019_d N_VGND_M1033_d N_VGND_M1031_s N_VGND_M1010_d N_VGND_M1024_s
+ N_VGND_c_1361_n N_VGND_c_1362_n N_VGND_c_1363_n N_VGND_c_1364_n
+ N_VGND_c_1365_n N_VGND_c_1366_n N_VGND_c_1367_n N_VGND_c_1368_n
+ N_VGND_c_1369_n N_VGND_c_1370_n N_VGND_c_1371_n N_VGND_c_1372_n
+ N_VGND_c_1373_n N_VGND_c_1374_n N_VGND_c_1375_n N_VGND_c_1376_n VGND
+ N_VGND_c_1377_n N_VGND_c_1378_n N_VGND_c_1379_n N_VGND_c_1380_n
+ N_VGND_c_1381_n N_VGND_c_1382_n N_VGND_c_1383_n N_VGND_c_1384_n
+ N_VGND_c_1385_n PM_SKY130_FD_SC_LP__HA_4%VGND
x_PM_SKY130_FD_SC_LP__HA_4%A_851_47# N_A_851_47#_M1020_d N_A_851_47#_M1002_s
+ N_A_851_47#_c_1526_n N_A_851_47#_c_1527_n N_A_851_47#_c_1528_n
+ PM_SKY130_FD_SC_LP__HA_4%A_851_47#
x_PM_SKY130_FD_SC_LP__HA_4%A_1284_65# N_A_1284_65#_M1010_s N_A_1284_65#_M1011_d
+ N_A_1284_65#_M1029_s N_A_1284_65#_M1026_s N_A_1284_65#_c_1552_n
+ N_A_1284_65#_c_1561_n N_A_1284_65#_c_1553_n N_A_1284_65#_c_1554_n
+ N_A_1284_65#_c_1563_n N_A_1284_65#_c_1564_n N_A_1284_65#_c_1567_n
+ N_A_1284_65#_c_1555_n N_A_1284_65#_c_1556_n N_A_1284_65#_c_1557_n
+ N_A_1284_65#_c_1577_n N_A_1284_65#_c_1578_n
+ PM_SKY130_FD_SC_LP__HA_4%A_1284_65#
cc_1 VNB N_A_110_263#_M1003_g 4.98466e-19 $X=-0.19 $Y=-0.245 $X2=0.625 $Y2=2.465
cc_2 VNB N_A_110_263#_M1009_g 0.0259851f $X=-0.19 $Y=-0.245 $X2=0.66 $Y2=0.655
cc_3 VNB N_A_110_263#_M1014_g 4.57504e-19 $X=-0.19 $Y=-0.245 $X2=1.055 $Y2=2.465
cc_4 VNB N_A_110_263#_M1021_g 0.0213937f $X=-0.19 $Y=-0.245 $X2=1.09 $Y2=0.655
cc_5 VNB N_A_110_263#_M1025_g 4.57707e-19 $X=-0.19 $Y=-0.245 $X2=1.485 $Y2=2.465
cc_6 VNB N_A_110_263#_M1022_g 0.0214084f $X=-0.19 $Y=-0.245 $X2=1.52 $Y2=0.655
cc_7 VNB N_A_110_263#_M1035_g 4.72413e-19 $X=-0.19 $Y=-0.245 $X2=1.915 $Y2=2.465
cc_8 VNB N_A_110_263#_M1034_g 0.0229053f $X=-0.19 $Y=-0.245 $X2=1.95 $Y2=0.655
cc_9 VNB N_A_110_263#_c_197_n 0.00425932f $X=-0.19 $Y=-0.245 $X2=2.075 $Y2=1.48
cc_10 VNB N_A_110_263#_c_198_n 0.00794445f $X=-0.19 $Y=-0.245 $X2=9.425
+ $Y2=1.755
cc_11 VNB N_A_110_263#_c_199_n 0.0221093f $X=-0.19 $Y=-0.245 $X2=9.215 $Y2=0.925
cc_12 VNB N_A_110_263#_c_200_n 0.00552246f $X=-0.19 $Y=-0.245 $X2=2.16 $Y2=0.925
cc_13 VNB N_A_110_263#_c_201_n 0.081704f $X=-0.19 $Y=-0.245 $X2=1.95 $Y2=1.48
cc_14 VNB N_A_454_263#_M1006_g 0.00959882f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_454_263#_M1016_g 0.0219219f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_454_263#_M1012_g 4.55097e-19 $X=-0.19 $Y=-0.245 $X2=1.055
+ $Y2=2.465
cc_17 VNB N_A_454_263#_M1019_g 0.0213691f $X=-0.19 $Y=-0.245 $X2=1.09 $Y2=0.655
cc_18 VNB N_A_454_263#_M1023_g 4.56909e-19 $X=-0.19 $Y=-0.245 $X2=1.485
+ $Y2=2.465
cc_19 VNB N_A_454_263#_M1030_g 0.0213857f $X=-0.19 $Y=-0.245 $X2=1.52 $Y2=0.655
cc_20 VNB N_A_454_263#_M1032_g 4.71393e-19 $X=-0.19 $Y=-0.245 $X2=1.915
+ $Y2=2.465
cc_21 VNB N_A_454_263#_M1033_g 0.0226565f $X=-0.19 $Y=-0.245 $X2=1.95 $Y2=0.655
cc_22 VNB N_A_454_263#_M1005_g 0.0191654f $X=-0.19 $Y=-0.245 $X2=1.86 $Y2=1.48
cc_23 VNB N_A_454_263#_c_437_n 0.00884591f $X=-0.19 $Y=-0.245 $X2=1.86 $Y2=1.48
cc_24 VNB N_A_454_263#_M1026_g 0.0231046f $X=-0.19 $Y=-0.245 $X2=6.82 $Y2=2.355
cc_25 VNB N_A_454_263#_M1015_g 0.0148695f $X=-0.19 $Y=-0.245 $X2=9.04 $Y2=2.27
cc_26 VNB N_A_454_263#_c_440_n 0.00696733f $X=-0.19 $Y=-0.245 $X2=9.125 $Y2=1.84
cc_27 VNB N_A_454_263#_c_441_n 0.0286887f $X=-0.19 $Y=-0.245 $X2=9.425 $Y2=1.755
cc_28 VNB N_A_454_263#_c_442_n 0.00206355f $X=-0.19 $Y=-0.245 $X2=6.545 $Y2=2.56
cc_29 VNB N_A_454_263#_c_443_n 6.24225e-19 $X=-0.19 $Y=-0.245 $X2=8.615
+ $Y2=2.405
cc_30 VNB N_A_454_263#_c_444_n 0.0102285f $X=-0.19 $Y=-0.245 $X2=8.45 $Y2=2.36
cc_31 VNB N_A_454_263#_c_445_n 0.00117459f $X=-0.19 $Y=-0.245 $X2=1.915 $Y2=1.48
cc_32 VNB N_A_454_263#_c_446_n 0.00200204f $X=-0.19 $Y=-0.245 $X2=1.95 $Y2=1.48
cc_33 VNB N_A_454_263#_c_447_n 0.003525f $X=-0.19 $Y=-0.245 $X2=2.16 $Y2=0.925
cc_34 VNB N_A_454_263#_c_448_n 0.00104295f $X=-0.19 $Y=-0.245 $X2=9.2 $Y2=0.7
cc_35 VNB N_A_454_263#_c_449_n 0.00924492f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_454_263#_c_450_n 0.0575381f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_454_263#_c_451_n 0.0231053f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_M1020_g 0.0253265f $X=-0.19 $Y=-0.245 $X2=8.395 $Y2=1.835
cc_39 VNB N_A_M1031_g 0.0276626f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_M1011_g 0.0213314f $X=-0.19 $Y=-0.245 $X2=1.055 $Y2=2.465
cc_41 VNB N_A_M1024_g 0.0225575f $X=-0.19 $Y=-0.245 $X2=1.09 $Y2=0.655
cc_42 VNB N_A_c_699_n 0.00377352f $X=-0.19 $Y=-0.245 $X2=1.52 $Y2=1.315
cc_43 VNB N_A_c_700_n 0.0235337f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_c_701_n 0.0320941f $X=-0.19 $Y=-0.245 $X2=0.84 $Y2=1.48
cc_45 VNB A 0.00526709f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_c_703_n 0.0472936f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_c_704_n 0.00232022f $X=-0.19 $Y=-0.245 $X2=6.51 $Y2=2.417
cc_48 VNB N_A_c_705_n 0.00296105f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_c_706_n 0.00136288f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_B_M1001_g 0.0196887f $X=-0.19 $Y=-0.245 $X2=8.395 $Y2=1.835
cc_51 VNB N_B_M1007_g 0.00893442f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_B_c_867_n 0.0108887f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_B_M1002_g 0.0200738f $X=-0.19 $Y=-0.245 $X2=0.625 $Y2=1.645
cc_54 VNB N_B_M1027_g 0.00317493f $X=-0.19 $Y=-0.245 $X2=0.66 $Y2=1.315
cc_55 VNB N_B_c_870_n 0.0220573f $X=-0.19 $Y=-0.245 $X2=0.66 $Y2=0.655
cc_56 VNB N_B_c_871_n 0.0212396f $X=-0.19 $Y=-0.245 $X2=1.055 $Y2=1.645
cc_57 VNB N_B_M1008_g 0.0163062f $X=-0.19 $Y=-0.245 $X2=1.09 $Y2=0.655
cc_58 VNB N_B_M1029_g 0.0243713f $X=-0.19 $Y=-0.245 $X2=1.52 $Y2=0.655
cc_59 VNB N_B_c_874_n 0.00468939f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_B_c_875_n 0.00556806f $X=-0.19 $Y=-0.245 $X2=1.915 $Y2=1.645
cc_61 VNB N_B_c_876_n 0.00923264f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_B_c_877_n 0.00445092f $X=-0.19 $Y=-0.245 $X2=1.95 $Y2=0.655
cc_63 VNB N_B_c_878_n 0.0376007f $X=-0.19 $Y=-0.245 $X2=0.84 $Y2=1.48
cc_64 VNB N_B_c_879_n 0.0107349f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_B_c_880_n 0.00496049f $X=-0.19 $Y=-0.245 $X2=1.86 $Y2=1.48
cc_66 VNB N_B_c_881_n 0.0251386f $X=-0.19 $Y=-0.245 $X2=6.51 $Y2=2.565
cc_67 VNB N_B_c_882_n 0.0345865f $X=-0.19 $Y=-0.245 $X2=9.425 $Y2=1.145
cc_68 VNB B 0.00626431f $X=-0.19 $Y=-0.245 $X2=9.837 $Y2=1.925
cc_69 VNB N_VPWR_c_1030_n 0.422413f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_SUM_c_1204_n 0.00259121f $X=-0.19 $Y=-0.245 $X2=0.625 $Y2=1.645
cc_71 VNB N_SUM_c_1205_n 0.00578413f $X=-0.19 $Y=-0.245 $X2=1.485 $Y2=1.645
cc_72 VNB N_SUM_c_1206_n 0.00147023f $X=-0.19 $Y=-0.245 $X2=1.95 $Y2=0.655
cc_73 VNB N_SUM_c_1207_n 0.0167448f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB SUM 0.025209f $X=-0.19 $Y=-0.245 $X2=1.86 $Y2=1.48
cc_75 VNB N_COUT_c_1264_n 0.0037883f $X=-0.19 $Y=-0.245 $X2=0.625 $Y2=2.465
cc_76 VNB N_COUT_c_1265_n 0.00579255f $X=-0.19 $Y=-0.245 $X2=0.66 $Y2=0.655
cc_77 VNB N_COUT_c_1266_n 9.82815e-19 $X=-0.19 $Y=-0.245 $X2=1.52 $Y2=1.315
cc_78 VNB N_VGND_c_1361_n 0.0269916f $X=-0.19 $Y=-0.245 $X2=1.09 $Y2=0.655
cc_79 VNB N_VGND_c_1362_n 0.0129398f $X=-0.19 $Y=-0.245 $X2=1.485 $Y2=1.645
cc_80 VNB N_VGND_c_1363_n 3.0911e-19 $X=-0.19 $Y=-0.245 $X2=1.52 $Y2=1.315
cc_81 VNB N_VGND_c_1364_n 3.0911e-19 $X=-0.19 $Y=-0.245 $X2=1.915 $Y2=1.645
cc_82 VNB N_VGND_c_1365_n 3.0911e-19 $X=-0.19 $Y=-0.245 $X2=1.95 $Y2=1.315
cc_83 VNB N_VGND_c_1366_n 0.00274891f $X=-0.19 $Y=-0.245 $X2=2.075 $Y2=1.48
cc_84 VNB N_VGND_c_1367_n 0.0185889f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_VGND_c_1368_n 0.00768835f $X=-0.19 $Y=-0.245 $X2=6.51 $Y2=2.565
cc_86 VNB N_VGND_c_1369_n 0.0110534f $X=-0.19 $Y=-0.245 $X2=8.45 $Y2=2.355
cc_87 VNB N_VGND_c_1370_n 0.00513431f $X=-0.19 $Y=-0.245 $X2=6.82 $Y2=2.355
cc_88 VNB N_VGND_c_1371_n 0.0129398f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_VGND_c_1372_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=9.04 $Y2=1.925
cc_90 VNB N_VGND_c_1373_n 0.0129398f $X=-0.19 $Y=-0.245 $X2=9.34 $Y2=1.84
cc_91 VNB N_VGND_c_1374_n 0.00532666f $X=-0.19 $Y=-0.245 $X2=9.125 $Y2=1.84
cc_92 VNB N_VGND_c_1375_n 0.0379942f $X=-0.19 $Y=-0.245 $X2=9.425 $Y2=1.755
cc_93 VNB N_VGND_c_1376_n 0.00548191f $X=-0.19 $Y=-0.245 $X2=9.69 $Y2=1.84
cc_94 VNB N_VGND_c_1377_n 0.0129398f $X=-0.19 $Y=-0.245 $X2=9.82 $Y2=2.91
cc_95 VNB N_VGND_c_1378_n 0.0285929f $X=-0.19 $Y=-0.245 $X2=9.36 $Y2=0.925
cc_96 VNB N_VGND_c_1379_n 0.0152967f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_97 VNB N_VGND_c_1380_n 0.0425166f $X=-0.19 $Y=-0.245 $X2=1.86 $Y2=1.48
cc_98 VNB N_VGND_c_1381_n 0.513091f $X=-0.19 $Y=-0.245 $X2=1.915 $Y2=1.48
cc_99 VNB N_VGND_c_1382_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=2.16 $Y2=0.925
cc_100 VNB N_VGND_c_1383_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=9.2 $Y2=0.7
cc_101 VNB N_VGND_c_1384_n 0.00631846f $X=-0.19 $Y=-0.245 $X2=9.272 $Y2=1.145
cc_102 VNB N_VGND_c_1385_n 0.0185583f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_103 VNB N_A_1284_65#_c_1552_n 0.00608525f $X=-0.19 $Y=-0.245 $X2=0.625
+ $Y2=2.465
cc_104 VNB N_A_1284_65#_c_1553_n 0.002805f $X=-0.19 $Y=-0.245 $X2=0.66 $Y2=0.655
cc_105 VNB N_A_1284_65#_c_1554_n 0.00208605f $X=-0.19 $Y=-0.245 $X2=1.055
+ $Y2=1.645
cc_106 VNB N_A_1284_65#_c_1555_n 0.013221f $X=-0.19 $Y=-0.245 $X2=1.485
+ $Y2=2.465
cc_107 VNB N_A_1284_65#_c_1556_n 0.00192831f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_108 VNB N_A_1284_65#_c_1557_n 0.0317446f $X=-0.19 $Y=-0.245 $X2=1.52
+ $Y2=0.655
cc_109 VPB N_A_110_263#_M1003_g 0.0225273f $X=-0.19 $Y=1.655 $X2=0.625 $Y2=2.465
cc_110 VPB N_A_110_263#_M1014_g 0.0188943f $X=-0.19 $Y=1.655 $X2=1.055 $Y2=2.465
cc_111 VPB N_A_110_263#_M1025_g 0.018914f $X=-0.19 $Y=1.655 $X2=1.485 $Y2=2.465
cc_112 VPB N_A_110_263#_M1035_g 0.02013f $X=-0.19 $Y=1.655 $X2=1.915 $Y2=2.465
cc_113 VPB N_A_110_263#_c_206_n 0.00838926f $X=-0.19 $Y=1.655 $X2=6.51 $Y2=2.565
cc_114 VPB N_A_110_263#_c_207_n 0.0031179f $X=-0.19 $Y=1.655 $X2=6.82 $Y2=2.355
cc_115 VPB N_A_110_263#_c_208_n 0.00229096f $X=-0.19 $Y=1.655 $X2=9.34 $Y2=1.84
cc_116 VPB N_A_110_263#_c_209_n 8.11403e-19 $X=-0.19 $Y=1.655 $X2=9.125 $Y2=1.84
cc_117 VPB N_A_110_263#_c_198_n 0.00191374f $X=-0.19 $Y=1.655 $X2=9.425
+ $Y2=1.755
cc_118 VPB N_A_110_263#_c_211_n 0.0138391f $X=-0.19 $Y=1.655 $X2=9.69 $Y2=1.84
cc_119 VPB N_A_110_263#_c_212_n 0.0441787f $X=-0.19 $Y=1.655 $X2=9.82 $Y2=1.98
cc_120 VPB N_A_454_263#_M1006_g 0.0201041f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_121 VPB N_A_454_263#_M1012_g 0.01908f $X=-0.19 $Y=1.655 $X2=1.055 $Y2=2.465
cc_122 VPB N_A_454_263#_M1023_g 0.0190693f $X=-0.19 $Y=1.655 $X2=1.485 $Y2=2.465
cc_123 VPB N_A_454_263#_M1032_g 0.0209516f $X=-0.19 $Y=1.655 $X2=1.915 $Y2=2.465
cc_124 VPB N_A_454_263#_M1004_g 0.0234937f $X=-0.19 $Y=1.655 $X2=0.84 $Y2=1.48
cc_125 VPB N_A_454_263#_M1015_g 0.0284167f $X=-0.19 $Y=1.655 $X2=9.04 $Y2=2.27
cc_126 VPB N_A_454_263#_c_443_n 0.00316024f $X=-0.19 $Y=1.655 $X2=8.615
+ $Y2=2.405
cc_127 VPB N_A_454_263#_c_459_n 0.0215394f $X=-0.19 $Y=1.655 $X2=1.055 $Y2=1.48
cc_128 VPB N_A_454_263#_c_445_n 0.00345006f $X=-0.19 $Y=1.655 $X2=1.915 $Y2=1.48
cc_129 VPB N_A_454_263#_c_461_n 0.00986601f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_130 VPB N_A_454_263#_c_451_n 0.00451573f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_131 VPB N_A_M1000_g 0.0204802f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_132 VPB N_A_M1017_g 0.0217638f $X=-0.19 $Y=1.655 $X2=0.625 $Y2=2.465
cc_133 VPB N_A_M1013_g 0.0208598f $X=-0.19 $Y=1.655 $X2=0.66 $Y2=0.655
cc_134 VPB N_A_M1018_g 0.0212309f $X=-0.19 $Y=1.655 $X2=1.485 $Y2=2.465
cc_135 VPB N_A_c_699_n 0.00325385f $X=-0.19 $Y=1.655 $X2=1.52 $Y2=1.315
cc_136 VPB N_A_c_700_n 0.00565746f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_137 VPB N_A_c_713_n 0.0057732f $X=-0.19 $Y=1.655 $X2=1.915 $Y2=2.465
cc_138 VPB N_A_c_714_n 4.56824e-19 $X=-0.19 $Y=1.655 $X2=2.075 $Y2=1.48
cc_139 VPB N_A_c_701_n 0.00693548f $X=-0.19 $Y=1.655 $X2=0.84 $Y2=1.48
cc_140 VPB A 0.00731372f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_141 VPB N_A_c_717_n 0.00253205f $X=-0.19 $Y=1.655 $X2=9.837 $Y2=2.91
cc_142 VPB N_A_c_703_n 0.0143978f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_143 VPB N_A_c_704_n 0.00169939f $X=-0.19 $Y=1.655 $X2=6.51 $Y2=2.417
cc_144 VPB N_A_c_705_n 0.0015344f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_145 VPB N_A_c_706_n 0.00439465f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_146 VPB N_B_M1007_g 0.0194906f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_147 VPB N_B_M1027_g 0.0189997f $X=-0.19 $Y=1.655 $X2=0.66 $Y2=1.315
cc_148 VPB N_B_M1008_g 0.0242684f $X=-0.19 $Y=1.655 $X2=1.09 $Y2=0.655
cc_149 VPB N_B_M1028_g 0.0201048f $X=-0.19 $Y=1.655 $X2=1.485 $Y2=2.465
cc_150 VPB N_B_c_882_n 0.00628305f $X=-0.19 $Y=1.655 $X2=9.425 $Y2=1.145
cc_151 VPB B 0.00347565f $X=-0.19 $Y=1.655 $X2=9.837 $Y2=1.925
cc_152 VPB N_VPWR_c_1031_n 0.0151245f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_153 VPB N_VPWR_c_1032_n 0.0415885f $X=-0.19 $Y=1.655 $X2=1.485 $Y2=2.465
cc_154 VPB N_VPWR_c_1033_n 3.15212e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_155 VPB N_VPWR_c_1034_n 0.00738827f $X=-0.19 $Y=1.655 $X2=1.95 $Y2=0.655
cc_156 VPB N_VPWR_c_1035_n 0.00373551f $X=-0.19 $Y=1.655 $X2=0.84 $Y2=1.48
cc_157 VPB N_VPWR_c_1036_n 0.00222527f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_158 VPB N_VPWR_c_1037_n 3.34013e-19 $X=-0.19 $Y=1.655 $X2=9.04 $Y2=2.27
cc_159 VPB N_VPWR_c_1038_n 0.0149194f $X=-0.19 $Y=1.655 $X2=9.425 $Y2=1.755
cc_160 VPB N_VPWR_c_1039_n 0.00408071f $X=-0.19 $Y=1.655 $X2=9.82 $Y2=1.98
cc_161 VPB N_VPWR_c_1040_n 0.0173748f $X=-0.19 $Y=1.655 $X2=6.545 $Y2=2.56
cc_162 VPB N_VPWR_c_1041_n 0.00410625f $X=-0.19 $Y=1.655 $X2=8.615 $Y2=2.36
cc_163 VPB N_VPWR_c_1042_n 0.0149824f $X=-0.19 $Y=1.655 $X2=8.45 $Y2=2.36
cc_164 VPB N_VPWR_c_1043_n 0.00510842f $X=-0.19 $Y=1.655 $X2=9.04 $Y2=2.36
cc_165 VPB N_VPWR_c_1044_n 0.0172194f $X=-0.19 $Y=1.655 $X2=9.425 $Y2=1.84
cc_166 VPB N_VPWR_c_1045_n 0.00436868f $X=-0.19 $Y=1.655 $X2=9.215 $Y2=0.925
cc_167 VPB N_VPWR_c_1046_n 0.0133881f $X=-0.19 $Y=1.655 $X2=2.16 $Y2=0.925
cc_168 VPB N_VPWR_c_1047_n 0.00510842f $X=-0.19 $Y=1.655 $X2=2.16 $Y2=0.925
cc_169 VPB N_VPWR_c_1048_n 0.0129398f $X=-0.19 $Y=1.655 $X2=9.36 $Y2=0.925
cc_170 VPB N_VPWR_c_1049_n 0.0147711f $X=-0.19 $Y=1.655 $X2=0.66 $Y2=1.48
cc_171 VPB N_VPWR_c_1050_n 0.0401112f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_172 VPB N_VPWR_c_1051_n 0.0322729f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_173 VPB N_VPWR_c_1052_n 0.0172072f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_174 VPB N_VPWR_c_1030_n 0.0721188f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_175 VPB N_VPWR_c_1054_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_176 VPB N_VPWR_c_1055_n 0.00487897f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_177 VPB N_VPWR_c_1056_n 0.0113436f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_178 VPB N_VPWR_c_1057_n 0.00963599f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_179 VPB N_SUM_c_1209_n 0.00232651f $X=-0.19 $Y=1.655 $X2=0.625 $Y2=2.465
cc_180 VPB N_SUM_c_1210_n 0.0150795f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_181 VPB N_SUM_c_1211_n 0.00592362f $X=-0.19 $Y=1.655 $X2=1.09 $Y2=0.655
cc_182 VPB N_SUM_c_1212_n 0.00149902f $X=-0.19 $Y=1.655 $X2=1.95 $Y2=0.655
cc_183 VPB SUM 0.00569894f $X=-0.19 $Y=1.655 $X2=1.86 $Y2=1.48
cc_184 VPB N_COUT_c_1264_n 0.00215235f $X=-0.19 $Y=1.655 $X2=0.625 $Y2=2.465
cc_185 VPB N_COUT_c_1268_n 0.00492294f $X=-0.19 $Y=1.655 $X2=1.055 $Y2=1.645
cc_186 VPB N_COUT_c_1269_n 0.00225024f $X=-0.19 $Y=1.655 $X2=1.52 $Y2=0.655
cc_187 N_A_110_263#_c_199_n N_A_454_263#_M1001_d 0.00135308f $X=9.215 $Y=0.925
+ $X2=-0.19 $Y2=-0.245
cc_188 N_A_110_263#_M1035_g N_A_454_263#_M1006_g 0.021484f $X=1.915 $Y=2.465
+ $X2=0 $Y2=0
cc_189 N_A_110_263#_M1034_g N_A_454_263#_M1016_g 0.0351183f $X=1.95 $Y=0.655
+ $X2=0 $Y2=0
cc_190 N_A_110_263#_c_199_n N_A_454_263#_M1016_g 0.0108286f $X=9.215 $Y=0.925
+ $X2=0 $Y2=0
cc_191 N_A_110_263#_c_217_p N_A_454_263#_M1016_g 0.00243785f $X=2.305 $Y=0.925
+ $X2=0 $Y2=0
cc_192 N_A_110_263#_c_200_n N_A_454_263#_M1016_g 0.00332633f $X=2.16 $Y=0.925
+ $X2=0 $Y2=0
cc_193 N_A_110_263#_c_199_n N_A_454_263#_M1019_g 0.00666595f $X=9.215 $Y=0.925
+ $X2=0 $Y2=0
cc_194 N_A_110_263#_c_199_n N_A_454_263#_M1030_g 0.00666595f $X=9.215 $Y=0.925
+ $X2=0 $Y2=0
cc_195 N_A_110_263#_c_199_n N_A_454_263#_M1033_g 0.00815201f $X=9.215 $Y=0.925
+ $X2=0 $Y2=0
cc_196 N_A_110_263#_c_222_p N_A_454_263#_M1004_g 0.00950023f $X=9.04 $Y=2.27
+ $X2=0 $Y2=0
cc_197 N_A_110_263#_c_209_n N_A_454_263#_M1004_g 0.00563752f $X=9.125 $Y=1.84
+ $X2=0 $Y2=0
cc_198 N_A_110_263#_c_198_n N_A_454_263#_M1004_g 8.66121e-19 $X=9.425 $Y=1.755
+ $X2=0 $Y2=0
cc_199 N_A_110_263#_c_225_p N_A_454_263#_M1004_g 0.00678733f $X=8.615 $Y=2.405
+ $X2=0 $Y2=0
cc_200 N_A_110_263#_c_226_p N_A_454_263#_M1004_g 0.0182767f $X=9.04 $Y=2.36
+ $X2=0 $Y2=0
cc_201 N_A_110_263#_c_198_n N_A_454_263#_M1005_g 0.00100605f $X=9.425 $Y=1.755
+ $X2=0 $Y2=0
cc_202 N_A_110_263#_c_199_n N_A_454_263#_M1005_g 0.00300773f $X=9.215 $Y=0.925
+ $X2=0 $Y2=0
cc_203 N_A_110_263#_c_229_p N_A_454_263#_M1005_g 0.00618083f $X=9.2 $Y=0.7 $X2=0
+ $Y2=0
cc_204 N_A_110_263#_c_208_n N_A_454_263#_c_437_n 0.00401553f $X=9.34 $Y=1.84
+ $X2=0 $Y2=0
cc_205 N_A_110_263#_c_198_n N_A_454_263#_M1026_g 0.00705783f $X=9.425 $Y=1.755
+ $X2=0 $Y2=0
cc_206 N_A_110_263#_c_229_p N_A_454_263#_M1026_g 0.0171703f $X=9.2 $Y=0.7 $X2=0
+ $Y2=0
cc_207 N_A_110_263#_c_222_p N_A_454_263#_M1015_g 0.0015459f $X=9.04 $Y=2.27
+ $X2=0 $Y2=0
cc_208 N_A_110_263#_c_198_n N_A_454_263#_M1015_g 0.0074869f $X=9.425 $Y=1.755
+ $X2=0 $Y2=0
cc_209 N_A_110_263#_c_211_n N_A_454_263#_M1015_g 0.0198738f $X=9.69 $Y=1.84
+ $X2=0 $Y2=0
cc_210 N_A_110_263#_c_197_n N_A_454_263#_c_440_n 0.00153174f $X=2.075 $Y=1.48
+ $X2=0 $Y2=0
cc_211 N_A_110_263#_c_217_p N_A_454_263#_c_440_n 9.73607e-19 $X=2.305 $Y=0.925
+ $X2=0 $Y2=0
cc_212 N_A_110_263#_c_200_n N_A_454_263#_c_440_n 7.02094e-19 $X=2.16 $Y=0.925
+ $X2=0 $Y2=0
cc_213 N_A_110_263#_c_201_n N_A_454_263#_c_440_n 0.01754f $X=1.95 $Y=1.48 $X2=0
+ $Y2=0
cc_214 N_A_110_263#_c_198_n N_A_454_263#_c_441_n 0.016556f $X=9.425 $Y=1.755
+ $X2=0 $Y2=0
cc_215 N_A_110_263#_c_211_n N_A_454_263#_c_441_n 5.93267e-19 $X=9.69 $Y=1.84
+ $X2=0 $Y2=0
cc_216 N_A_110_263#_c_199_n N_A_454_263#_c_492_n 0.00588371f $X=9.215 $Y=0.925
+ $X2=0 $Y2=0
cc_217 N_A_110_263#_c_199_n N_A_454_263#_c_444_n 0.0347526f $X=9.215 $Y=0.925
+ $X2=0 $Y2=0
cc_218 N_A_110_263#_c_199_n N_A_454_263#_c_494_n 0.00554859f $X=9.215 $Y=0.925
+ $X2=0 $Y2=0
cc_219 N_A_110_263#_c_199_n N_A_454_263#_c_495_n 0.0153382f $X=9.215 $Y=0.925
+ $X2=0 $Y2=0
cc_220 N_A_110_263#_M1008_d N_A_454_263#_c_496_n 0.00451902f $X=6.42 $Y=1.835
+ $X2=0 $Y2=0
cc_221 N_A_110_263#_M1028_d N_A_454_263#_c_496_n 0.00886509f $X=8.395 $Y=1.835
+ $X2=0 $Y2=0
cc_222 N_A_110_263#_c_207_n N_A_454_263#_c_496_n 0.0181599f $X=6.82 $Y=2.355
+ $X2=0 $Y2=0
cc_223 N_A_110_263#_c_222_p N_A_454_263#_c_496_n 0.0128377f $X=9.04 $Y=2.27
+ $X2=0 $Y2=0
cc_224 N_A_110_263#_c_250_p N_A_454_263#_c_496_n 0.0983908f $X=8.45 $Y=2.36
+ $X2=0 $Y2=0
cc_225 N_A_110_263#_c_226_p N_A_454_263#_c_496_n 0.013819f $X=9.04 $Y=2.36 $X2=0
+ $Y2=0
cc_226 N_A_110_263#_M1028_d N_A_454_263#_c_445_n 0.00274351f $X=8.395 $Y=1.835
+ $X2=0 $Y2=0
cc_227 N_A_110_263#_c_222_p N_A_454_263#_c_445_n 2.68697e-19 $X=9.04 $Y=2.27
+ $X2=0 $Y2=0
cc_228 N_A_110_263#_c_209_n N_A_454_263#_c_445_n 0.0128858f $X=9.125 $Y=1.84
+ $X2=0 $Y2=0
cc_229 N_A_110_263#_c_198_n N_A_454_263#_c_445_n 0.00579644f $X=9.425 $Y=1.755
+ $X2=0 $Y2=0
cc_230 N_A_110_263#_c_199_n N_A_454_263#_c_446_n 0.00116831f $X=9.215 $Y=0.925
+ $X2=0 $Y2=0
cc_231 N_A_110_263#_c_208_n N_A_454_263#_c_447_n 0.00304683f $X=9.34 $Y=1.84
+ $X2=0 $Y2=0
cc_232 N_A_110_263#_c_209_n N_A_454_263#_c_447_n 0.0126773f $X=9.125 $Y=1.84
+ $X2=0 $Y2=0
cc_233 N_A_110_263#_c_198_n N_A_454_263#_c_447_n 0.012971f $X=9.425 $Y=1.755
+ $X2=0 $Y2=0
cc_234 N_A_110_263#_c_199_n N_A_454_263#_c_447_n 0.00650085f $X=9.215 $Y=0.925
+ $X2=0 $Y2=0
cc_235 N_A_110_263#_c_229_p N_A_454_263#_c_447_n 0.00488374f $X=9.2 $Y=0.7 $X2=0
+ $Y2=0
cc_236 N_A_110_263#_M1008_d N_A_454_263#_c_461_n 0.00359741f $X=6.42 $Y=1.835
+ $X2=0 $Y2=0
cc_237 N_A_110_263#_c_207_n N_A_454_263#_c_461_n 0.00735348f $X=6.82 $Y=2.355
+ $X2=0 $Y2=0
cc_238 N_A_110_263#_c_208_n N_A_454_263#_c_451_n 0.00120568f $X=9.34 $Y=1.84
+ $X2=0 $Y2=0
cc_239 N_A_110_263#_c_209_n N_A_454_263#_c_451_n 0.00398757f $X=9.125 $Y=1.84
+ $X2=0 $Y2=0
cc_240 N_A_110_263#_c_198_n N_A_454_263#_c_451_n 0.00125523f $X=9.425 $Y=1.755
+ $X2=0 $Y2=0
cc_241 N_A_110_263#_c_199_n N_A_454_263#_c_451_n 0.00137534f $X=9.215 $Y=0.925
+ $X2=0 $Y2=0
cc_242 N_A_110_263#_c_229_p N_A_454_263#_c_451_n 0.00248134f $X=9.2 $Y=0.7 $X2=0
+ $Y2=0
cc_243 N_A_110_263#_c_199_n N_A_M1020_g 0.0091494f $X=9.215 $Y=0.925 $X2=0 $Y2=0
cc_244 N_A_110_263#_c_199_n N_A_M1031_g 0.0091438f $X=9.215 $Y=0.925 $X2=0 $Y2=0
cc_245 N_A_110_263#_c_207_n N_A_M1013_g 7.56926e-19 $X=6.82 $Y=2.355 $X2=0 $Y2=0
cc_246 N_A_110_263#_c_250_p N_A_M1013_g 0.0116272f $X=8.45 $Y=2.36 $X2=0 $Y2=0
cc_247 N_A_110_263#_c_199_n N_A_M1011_g 0.00194685f $X=9.215 $Y=0.925 $X2=0
+ $Y2=0
cc_248 N_A_110_263#_c_199_n N_A_M1024_g 0.00247742f $X=9.215 $Y=0.925 $X2=0
+ $Y2=0
cc_249 N_A_110_263#_c_250_p N_A_M1018_g 0.0116147f $X=8.45 $Y=2.36 $X2=0 $Y2=0
cc_250 N_A_110_263#_c_199_n N_B_M1001_g 0.00423273f $X=9.215 $Y=0.925 $X2=0
+ $Y2=0
cc_251 N_A_110_263#_c_199_n N_B_M1002_g 0.00468816f $X=9.215 $Y=0.925 $X2=0
+ $Y2=0
cc_252 N_A_110_263#_c_199_n N_B_c_871_n 0.00194685f $X=9.215 $Y=0.925 $X2=0
+ $Y2=0
cc_253 N_A_110_263#_c_207_n N_B_M1008_g 0.0118423f $X=6.82 $Y=2.355 $X2=0 $Y2=0
cc_254 N_A_110_263#_c_250_p N_B_M1008_g 0.00263572f $X=8.45 $Y=2.36 $X2=0 $Y2=0
cc_255 N_A_110_263#_c_222_p N_B_M1028_g 9.03645e-19 $X=9.04 $Y=2.27 $X2=0 $Y2=0
cc_256 N_A_110_263#_c_250_p N_B_M1028_g 0.0150411f $X=8.45 $Y=2.36 $X2=0 $Y2=0
cc_257 N_A_110_263#_c_199_n N_B_M1029_g 0.00688812f $X=9.215 $Y=0.925 $X2=0
+ $Y2=0
cc_258 N_A_110_263#_c_229_p N_B_M1029_g 3.63342e-19 $X=9.2 $Y=0.7 $X2=0 $Y2=0
cc_259 N_A_110_263#_c_199_n N_B_c_877_n 0.0106603f $X=9.215 $Y=0.925 $X2=0 $Y2=0
cc_260 N_A_110_263#_c_199_n N_B_c_879_n 0.0761721f $X=9.215 $Y=0.925 $X2=0 $Y2=0
cc_261 N_A_110_263#_c_199_n B 0.0116561f $X=9.215 $Y=0.925 $X2=0 $Y2=0
cc_262 N_A_110_263#_c_250_p N_VPWR_M1013_d 0.0107167f $X=8.45 $Y=2.36 $X2=0
+ $Y2=0
cc_263 N_A_110_263#_c_222_p N_VPWR_M1004_s 0.00432078f $X=9.04 $Y=2.27 $X2=0
+ $Y2=0
cc_264 N_A_110_263#_c_208_n N_VPWR_M1004_s 0.00778717f $X=9.34 $Y=1.84 $X2=0
+ $Y2=0
cc_265 N_A_110_263#_c_226_p N_VPWR_M1004_s 0.00276213f $X=9.04 $Y=2.36 $X2=0
+ $Y2=0
cc_266 N_A_110_263#_c_292_p N_VPWR_M1004_s 0.0015577f $X=9.425 $Y=1.84 $X2=0
+ $Y2=0
cc_267 N_A_110_263#_M1003_g N_VPWR_c_1032_n 0.0152824f $X=0.625 $Y=2.465 $X2=0
+ $Y2=0
cc_268 N_A_110_263#_M1014_g N_VPWR_c_1032_n 7.27171e-19 $X=1.055 $Y=2.465 $X2=0
+ $Y2=0
cc_269 N_A_110_263#_M1003_g N_VPWR_c_1033_n 7.27171e-19 $X=0.625 $Y=2.465 $X2=0
+ $Y2=0
cc_270 N_A_110_263#_M1014_g N_VPWR_c_1033_n 0.0142189f $X=1.055 $Y=2.465 $X2=0
+ $Y2=0
cc_271 N_A_110_263#_M1025_g N_VPWR_c_1033_n 0.0142995f $X=1.485 $Y=2.465 $X2=0
+ $Y2=0
cc_272 N_A_110_263#_M1035_g N_VPWR_c_1033_n 7.4139e-19 $X=1.915 $Y=2.465 $X2=0
+ $Y2=0
cc_273 N_A_110_263#_M1035_g N_VPWR_c_1034_n 0.00268082f $X=1.915 $Y=2.465 $X2=0
+ $Y2=0
cc_274 N_A_110_263#_c_197_n N_VPWR_c_1034_n 0.0170277f $X=2.075 $Y=1.48 $X2=0
+ $Y2=0
cc_275 N_A_110_263#_c_201_n N_VPWR_c_1034_n 6.87012e-19 $X=1.95 $Y=1.48 $X2=0
+ $Y2=0
cc_276 N_A_110_263#_c_206_n N_VPWR_c_1038_n 0.0200402f $X=6.51 $Y=2.565 $X2=0
+ $Y2=0
cc_277 N_A_110_263#_c_207_n N_VPWR_c_1038_n 0.00703466f $X=6.82 $Y=2.355 $X2=0
+ $Y2=0
cc_278 N_A_110_263#_c_225_p N_VPWR_c_1074_n 0.0359573f $X=8.615 $Y=2.405 $X2=0
+ $Y2=0
cc_279 N_A_110_263#_c_226_p N_VPWR_c_1074_n 0.00895202f $X=9.04 $Y=2.36 $X2=0
+ $Y2=0
cc_280 N_A_110_263#_c_222_p N_VPWR_c_1076_n 0.0122415f $X=9.04 $Y=2.27 $X2=0
+ $Y2=0
cc_281 N_A_110_263#_c_208_n N_VPWR_c_1076_n 0.003395f $X=9.34 $Y=1.84 $X2=0
+ $Y2=0
cc_282 N_A_110_263#_c_225_p N_VPWR_c_1076_n 0.00613218f $X=8.615 $Y=2.405 $X2=0
+ $Y2=0
cc_283 N_A_110_263#_c_226_p N_VPWR_c_1076_n 0.0147598f $X=9.04 $Y=2.36 $X2=0
+ $Y2=0
cc_284 N_A_110_263#_c_292_p N_VPWR_c_1076_n 0.0114866f $X=9.425 $Y=1.84 $X2=0
+ $Y2=0
cc_285 N_A_110_263#_M1003_g N_VPWR_c_1048_n 0.00486043f $X=0.625 $Y=2.465 $X2=0
+ $Y2=0
cc_286 N_A_110_263#_M1014_g N_VPWR_c_1048_n 0.00486043f $X=1.055 $Y=2.465 $X2=0
+ $Y2=0
cc_287 N_A_110_263#_M1025_g N_VPWR_c_1049_n 0.00486043f $X=1.485 $Y=2.465 $X2=0
+ $Y2=0
cc_288 N_A_110_263#_M1035_g N_VPWR_c_1049_n 0.00585385f $X=1.915 $Y=2.465 $X2=0
+ $Y2=0
cc_289 N_A_110_263#_c_206_n N_VPWR_c_1050_n 0.0178111f $X=6.51 $Y=2.565 $X2=0
+ $Y2=0
cc_290 N_A_110_263#_c_225_p N_VPWR_c_1051_n 0.0228861f $X=8.615 $Y=2.405 $X2=0
+ $Y2=0
cc_291 N_A_110_263#_c_212_n N_VPWR_c_1052_n 0.0190529f $X=9.82 $Y=1.98 $X2=0
+ $Y2=0
cc_292 N_A_110_263#_M1008_d N_VPWR_c_1030_n 0.00238527f $X=6.42 $Y=1.835 $X2=0
+ $Y2=0
cc_293 N_A_110_263#_M1028_d N_VPWR_c_1030_n 0.00767727f $X=8.395 $Y=1.835 $X2=0
+ $Y2=0
cc_294 N_A_110_263#_M1015_d N_VPWR_c_1030_n 0.00249946f $X=9.68 $Y=1.835 $X2=0
+ $Y2=0
cc_295 N_A_110_263#_M1003_g N_VPWR_c_1030_n 0.00824727f $X=0.625 $Y=2.465 $X2=0
+ $Y2=0
cc_296 N_A_110_263#_M1014_g N_VPWR_c_1030_n 0.00824727f $X=1.055 $Y=2.465 $X2=0
+ $Y2=0
cc_297 N_A_110_263#_M1025_g N_VPWR_c_1030_n 0.00824727f $X=1.485 $Y=2.465 $X2=0
+ $Y2=0
cc_298 N_A_110_263#_M1035_g N_VPWR_c_1030_n 0.0105477f $X=1.915 $Y=2.465 $X2=0
+ $Y2=0
cc_299 N_A_110_263#_c_206_n N_VPWR_c_1030_n 0.0100304f $X=6.51 $Y=2.565 $X2=0
+ $Y2=0
cc_300 N_A_110_263#_c_207_n N_VPWR_c_1030_n 0.00559745f $X=6.82 $Y=2.355 $X2=0
+ $Y2=0
cc_301 N_A_110_263#_c_212_n N_VPWR_c_1030_n 0.0113912f $X=9.82 $Y=1.98 $X2=0
+ $Y2=0
cc_302 N_A_110_263#_c_225_p N_VPWR_c_1030_n 0.0127185f $X=8.615 $Y=2.405 $X2=0
+ $Y2=0
cc_303 N_A_110_263#_M1009_g N_SUM_c_1204_n 0.0167554f $X=0.66 $Y=0.655 $X2=0
+ $Y2=0
cc_304 N_A_110_263#_c_197_n N_SUM_c_1204_n 0.00693257f $X=2.075 $Y=1.48 $X2=0
+ $Y2=0
cc_305 N_A_110_263#_c_201_n N_SUM_c_1204_n 0.00115314f $X=1.95 $Y=1.48 $X2=0
+ $Y2=0
cc_306 N_A_110_263#_M1003_g N_SUM_c_1209_n 0.0162939f $X=0.625 $Y=2.465 $X2=0
+ $Y2=0
cc_307 N_A_110_263#_c_197_n N_SUM_c_1209_n 0.00447707f $X=2.075 $Y=1.48 $X2=0
+ $Y2=0
cc_308 N_A_110_263#_M1014_g N_SUM_c_1211_n 0.0132876f $X=1.055 $Y=2.465 $X2=0
+ $Y2=0
cc_309 N_A_110_263#_M1025_g N_SUM_c_1211_n 0.0131749f $X=1.485 $Y=2.465 $X2=0
+ $Y2=0
cc_310 N_A_110_263#_M1035_g N_SUM_c_1211_n 0.00114834f $X=1.915 $Y=2.465 $X2=0
+ $Y2=0
cc_311 N_A_110_263#_c_197_n N_SUM_c_1211_n 0.0595851f $X=2.075 $Y=1.48 $X2=0
+ $Y2=0
cc_312 N_A_110_263#_c_201_n N_SUM_c_1211_n 0.00527005f $X=1.95 $Y=1.48 $X2=0
+ $Y2=0
cc_313 N_A_110_263#_M1021_g N_SUM_c_1205_n 0.0139591f $X=1.09 $Y=0.655 $X2=0
+ $Y2=0
cc_314 N_A_110_263#_M1022_g N_SUM_c_1205_n 0.0136364f $X=1.52 $Y=0.655 $X2=0
+ $Y2=0
cc_315 N_A_110_263#_M1034_g N_SUM_c_1205_n 0.00136599f $X=1.95 $Y=0.655 $X2=0
+ $Y2=0
cc_316 N_A_110_263#_c_197_n N_SUM_c_1205_n 0.0593934f $X=2.075 $Y=1.48 $X2=0
+ $Y2=0
cc_317 N_A_110_263#_c_200_n N_SUM_c_1205_n 0.00907245f $X=2.16 $Y=0.925 $X2=0
+ $Y2=0
cc_318 N_A_110_263#_c_201_n N_SUM_c_1205_n 0.00530199f $X=1.95 $Y=1.48 $X2=0
+ $Y2=0
cc_319 N_A_110_263#_c_217_p N_SUM_c_1230_n 0.00663498f $X=2.305 $Y=0.925 $X2=0
+ $Y2=0
cc_320 N_A_110_263#_c_197_n N_SUM_c_1212_n 0.014105f $X=2.075 $Y=1.48 $X2=0
+ $Y2=0
cc_321 N_A_110_263#_c_201_n N_SUM_c_1212_n 0.00268975f $X=1.95 $Y=1.48 $X2=0
+ $Y2=0
cc_322 N_A_110_263#_c_197_n N_SUM_c_1206_n 0.014687f $X=2.075 $Y=1.48 $X2=0
+ $Y2=0
cc_323 N_A_110_263#_c_201_n N_SUM_c_1206_n 0.00270417f $X=1.95 $Y=1.48 $X2=0
+ $Y2=0
cc_324 N_A_110_263#_M1009_g SUM 0.00361203f $X=0.66 $Y=0.655 $X2=0 $Y2=0
cc_325 N_A_110_263#_c_197_n SUM 0.00992202f $X=2.075 $Y=1.48 $X2=0 $Y2=0
cc_326 N_A_110_263#_c_201_n SUM 0.0163274f $X=1.95 $Y=1.48 $X2=0 $Y2=0
cc_327 N_A_110_263#_c_199_n N_COUT_M1016_s 0.00389099f $X=9.215 $Y=0.925
+ $X2=-0.19 $Y2=-0.245
cc_328 N_A_110_263#_c_199_n N_COUT_M1030_s 0.00403064f $X=9.215 $Y=0.925 $X2=0
+ $Y2=0
cc_329 N_A_110_263#_c_197_n N_COUT_c_1264_n 0.0135133f $X=2.075 $Y=1.48 $X2=0
+ $Y2=0
cc_330 N_A_110_263#_c_200_n N_COUT_c_1264_n 0.0122303f $X=2.16 $Y=0.925 $X2=0
+ $Y2=0
cc_331 N_A_110_263#_c_199_n N_COUT_c_1274_n 0.0252989f $X=9.215 $Y=0.925 $X2=0
+ $Y2=0
cc_332 N_A_110_263#_c_217_p N_COUT_c_1274_n 0.00243274f $X=2.305 $Y=0.925 $X2=0
+ $Y2=0
cc_333 N_A_110_263#_c_200_n N_COUT_c_1274_n 0.00633079f $X=2.16 $Y=0.925 $X2=0
+ $Y2=0
cc_334 N_A_110_263#_c_199_n N_COUT_c_1265_n 0.024707f $X=9.215 $Y=0.925 $X2=0
+ $Y2=0
cc_335 N_A_110_263#_c_199_n N_COUT_c_1278_n 0.0240827f $X=9.215 $Y=0.925 $X2=0
+ $Y2=0
cc_336 N_A_110_263#_c_199_n N_COUT_c_1266_n 0.00406406f $X=9.215 $Y=0.925 $X2=0
+ $Y2=0
cc_337 N_A_110_263#_c_200_n N_COUT_c_1266_n 0.0129657f $X=2.16 $Y=0.925 $X2=0
+ $Y2=0
cc_338 N_A_110_263#_c_250_p N_A_1367_367#_M1008_s 0.0038777f $X=8.45 $Y=2.36
+ $X2=-0.19 $Y2=-0.245
cc_339 N_A_110_263#_c_250_p N_A_1367_367#_M1018_s 0.0035215f $X=8.45 $Y=2.36
+ $X2=0 $Y2=0
cc_340 N_A_110_263#_c_250_p N_A_1367_367#_c_1334_n 0.0465459f $X=8.45 $Y=2.36
+ $X2=0 $Y2=0
cc_341 N_A_110_263#_c_207_n N_A_1367_367#_c_1335_n 6.67238e-19 $X=6.82 $Y=2.355
+ $X2=0 $Y2=0
cc_342 N_A_110_263#_c_250_p N_A_1367_367#_c_1335_n 0.0142411f $X=8.45 $Y=2.36
+ $X2=0 $Y2=0
cc_343 N_A_110_263#_c_250_p N_A_1367_367#_c_1337_n 0.0161925f $X=8.45 $Y=2.36
+ $X2=0 $Y2=0
cc_344 N_A_110_263#_c_217_p N_VGND_M1034_s 0.00438817f $X=2.305 $Y=0.925 $X2=0
+ $Y2=0
cc_345 N_A_110_263#_c_200_n N_VGND_M1034_s 0.00445181f $X=2.16 $Y=0.925 $X2=0
+ $Y2=0
cc_346 N_A_110_263#_c_199_n N_VGND_M1019_d 0.00201894f $X=9.215 $Y=0.925 $X2=0
+ $Y2=0
cc_347 N_A_110_263#_c_199_n N_VGND_M1033_d 0.00513355f $X=9.215 $Y=0.925 $X2=0
+ $Y2=0
cc_348 N_A_110_263#_c_199_n N_VGND_M1031_s 0.00262872f $X=9.215 $Y=0.925 $X2=0
+ $Y2=0
cc_349 N_A_110_263#_c_199_n N_VGND_M1010_d 0.00324014f $X=9.215 $Y=0.925 $X2=0
+ $Y2=0
cc_350 N_A_110_263#_c_199_n N_VGND_M1024_s 0.00484878f $X=9.215 $Y=0.925 $X2=0
+ $Y2=0
cc_351 N_A_110_263#_M1009_g N_VGND_c_1361_n 0.012456f $X=0.66 $Y=0.655 $X2=0
+ $Y2=0
cc_352 N_A_110_263#_M1021_g N_VGND_c_1361_n 6.25324e-19 $X=1.09 $Y=0.655 $X2=0
+ $Y2=0
cc_353 N_A_110_263#_M1009_g N_VGND_c_1362_n 0.00486043f $X=0.66 $Y=0.655 $X2=0
+ $Y2=0
cc_354 N_A_110_263#_M1021_g N_VGND_c_1362_n 0.00486043f $X=1.09 $Y=0.655 $X2=0
+ $Y2=0
cc_355 N_A_110_263#_M1009_g N_VGND_c_1363_n 6.22495e-19 $X=0.66 $Y=0.655 $X2=0
+ $Y2=0
cc_356 N_A_110_263#_M1021_g N_VGND_c_1363_n 0.0107911f $X=1.09 $Y=0.655 $X2=0
+ $Y2=0
cc_357 N_A_110_263#_M1022_g N_VGND_c_1363_n 0.0107894f $X=1.52 $Y=0.655 $X2=0
+ $Y2=0
cc_358 N_A_110_263#_M1034_g N_VGND_c_1363_n 6.22495e-19 $X=1.95 $Y=0.655 $X2=0
+ $Y2=0
cc_359 N_A_110_263#_M1022_g N_VGND_c_1364_n 5.67328e-19 $X=1.52 $Y=0.655 $X2=0
+ $Y2=0
cc_360 N_A_110_263#_M1034_g N_VGND_c_1364_n 0.0104508f $X=1.95 $Y=0.655 $X2=0
+ $Y2=0
cc_361 N_A_110_263#_c_199_n N_VGND_c_1364_n 0.00101532f $X=9.215 $Y=0.925 $X2=0
+ $Y2=0
cc_362 N_A_110_263#_c_217_p N_VGND_c_1364_n 0.0116773f $X=2.305 $Y=0.925 $X2=0
+ $Y2=0
cc_363 N_A_110_263#_c_200_n N_VGND_c_1364_n 0.0117735f $X=2.16 $Y=0.925 $X2=0
+ $Y2=0
cc_364 N_A_110_263#_c_199_n N_VGND_c_1365_n 0.0201619f $X=9.215 $Y=0.925 $X2=0
+ $Y2=0
cc_365 N_A_110_263#_c_199_n N_VGND_c_1366_n 0.0101857f $X=9.215 $Y=0.925 $X2=0
+ $Y2=0
cc_366 N_A_110_263#_c_199_n N_VGND_c_1367_n 0.0216342f $X=9.215 $Y=0.925 $X2=0
+ $Y2=0
cc_367 N_A_110_263#_c_199_n N_VGND_c_1368_n 0.00207933f $X=9.215 $Y=0.925 $X2=0
+ $Y2=0
cc_368 N_A_110_263#_M1022_g N_VGND_c_1377_n 0.00486043f $X=1.52 $Y=0.655 $X2=0
+ $Y2=0
cc_369 N_A_110_263#_M1034_g N_VGND_c_1377_n 0.00486043f $X=1.95 $Y=0.655 $X2=0
+ $Y2=0
cc_370 N_A_110_263#_M1009_g N_VGND_c_1381_n 0.00824727f $X=0.66 $Y=0.655 $X2=0
+ $Y2=0
cc_371 N_A_110_263#_M1021_g N_VGND_c_1381_n 0.00824727f $X=1.09 $Y=0.655 $X2=0
+ $Y2=0
cc_372 N_A_110_263#_M1022_g N_VGND_c_1381_n 0.00824727f $X=1.52 $Y=0.655 $X2=0
+ $Y2=0
cc_373 N_A_110_263#_M1034_g N_VGND_c_1381_n 0.00824727f $X=1.95 $Y=0.655 $X2=0
+ $Y2=0
cc_374 N_A_110_263#_c_200_n N_VGND_c_1381_n 3.29889e-19 $X=2.16 $Y=0.925 $X2=0
+ $Y2=0
cc_375 N_A_110_263#_c_199_n N_VGND_c_1385_n 0.0116609f $X=9.215 $Y=0.925 $X2=0
+ $Y2=0
cc_376 N_A_110_263#_c_199_n N_A_851_47#_M1020_d 0.00318191f $X=9.215 $Y=0.925
+ $X2=-0.19 $Y2=-0.245
cc_377 N_A_110_263#_c_199_n N_A_851_47#_M1002_s 0.00463382f $X=9.215 $Y=0.925
+ $X2=0 $Y2=0
cc_378 N_A_110_263#_c_199_n N_A_851_47#_c_1526_n 0.00956405f $X=9.215 $Y=0.925
+ $X2=0 $Y2=0
cc_379 N_A_110_263#_c_199_n N_A_851_47#_c_1527_n 0.00969048f $X=9.215 $Y=0.925
+ $X2=0 $Y2=0
cc_380 N_A_110_263#_c_199_n N_A_851_47#_c_1528_n 0.0106965f $X=9.215 $Y=0.925
+ $X2=0 $Y2=0
cc_381 N_A_110_263#_c_199_n N_A_1284_65#_M1010_s 0.00194409f $X=9.215 $Y=0.925
+ $X2=-0.19 $Y2=-0.245
cc_382 N_A_110_263#_c_199_n N_A_1284_65#_M1011_d 0.00204646f $X=9.215 $Y=0.925
+ $X2=0 $Y2=0
cc_383 N_A_110_263#_c_199_n N_A_1284_65#_M1029_s 0.00238396f $X=9.215 $Y=0.925
+ $X2=0 $Y2=0
cc_384 N_A_110_263#_c_199_n N_A_1284_65#_c_1561_n 0.0278568f $X=9.215 $Y=0.925
+ $X2=0 $Y2=0
cc_385 N_A_110_263#_c_199_n N_A_1284_65#_c_1553_n 0.0210601f $X=9.215 $Y=0.925
+ $X2=0 $Y2=0
cc_386 N_A_110_263#_c_199_n N_A_1284_65#_c_1563_n 0.0120832f $X=9.215 $Y=0.925
+ $X2=0 $Y2=0
cc_387 N_A_110_263#_c_199_n N_A_1284_65#_c_1564_n 0.0276175f $X=9.215 $Y=0.925
+ $X2=0 $Y2=0
cc_388 N_A_110_263#_c_414_p N_A_1284_65#_c_1564_n 2.53795e-19 $X=9.36 $Y=0.925
+ $X2=0 $Y2=0
cc_389 N_A_110_263#_c_229_p N_A_1284_65#_c_1564_n 0.0071942f $X=9.2 $Y=0.7 $X2=0
+ $Y2=0
cc_390 N_A_110_263#_c_199_n N_A_1284_65#_c_1567_n 0.0139157f $X=9.215 $Y=0.925
+ $X2=0 $Y2=0
cc_391 N_A_110_263#_c_414_p N_A_1284_65#_c_1567_n 2.25469e-19 $X=9.36 $Y=0.925
+ $X2=0 $Y2=0
cc_392 N_A_110_263#_c_229_p N_A_1284_65#_c_1567_n 0.0123978f $X=9.2 $Y=0.7 $X2=0
+ $Y2=0
cc_393 N_A_110_263#_M1005_d N_A_1284_65#_c_1555_n 0.0017389f $X=9.06 $Y=0.325
+ $X2=0 $Y2=0
cc_394 N_A_110_263#_c_199_n N_A_1284_65#_c_1555_n 0.00627201f $X=9.215 $Y=0.925
+ $X2=0 $Y2=0
cc_395 N_A_110_263#_c_414_p N_A_1284_65#_c_1555_n 0.00134844f $X=9.36 $Y=0.925
+ $X2=0 $Y2=0
cc_396 N_A_110_263#_c_229_p N_A_1284_65#_c_1555_n 0.0221927f $X=9.2 $Y=0.7 $X2=0
+ $Y2=0
cc_397 N_A_110_263#_c_198_n N_A_1284_65#_c_1557_n 0.0210163f $X=9.425 $Y=1.755
+ $X2=0 $Y2=0
cc_398 N_A_110_263#_c_211_n N_A_1284_65#_c_1557_n 0.00992576f $X=9.69 $Y=1.84
+ $X2=0 $Y2=0
cc_399 N_A_110_263#_c_414_p N_A_1284_65#_c_1557_n 0.00173565f $X=9.36 $Y=0.925
+ $X2=0 $Y2=0
cc_400 N_A_110_263#_c_199_n N_A_1284_65#_c_1577_n 0.0167748f $X=9.215 $Y=0.925
+ $X2=0 $Y2=0
cc_401 N_A_110_263#_c_199_n N_A_1284_65#_c_1578_n 0.0113958f $X=9.215 $Y=0.925
+ $X2=0 $Y2=0
cc_402 N_A_454_263#_M1033_g N_A_M1020_g 0.0266358f $X=3.67 $Y=0.655 $X2=0 $Y2=0
cc_403 N_A_454_263#_c_442_n N_A_M1020_g 0.00363063f $X=3.805 $Y=1.395 $X2=0
+ $Y2=0
cc_404 N_A_454_263#_c_444_n N_A_M1020_g 0.0109501f $X=4.73 $Y=1.08 $X2=0 $Y2=0
cc_405 N_A_454_263#_c_450_n N_A_M1020_g 0.00101956f $X=3.67 $Y=1.48 $X2=0 $Y2=0
cc_406 N_A_454_263#_M1032_g N_A_M1000_g 0.0247993f $X=3.635 $Y=2.465 $X2=0 $Y2=0
cc_407 N_A_454_263#_c_443_n N_A_M1000_g 0.00189608f $X=3.805 $Y=1.855 $X2=0
+ $Y2=0
cc_408 N_A_454_263#_c_525_p N_A_M1000_g 0.00895433f $X=4.195 $Y=1.94 $X2=0 $Y2=0
cc_409 N_A_454_263#_c_526_p N_A_M1000_g 0.00717762f $X=4.352 $Y=2.215 $X2=0
+ $Y2=0
cc_410 N_A_454_263#_c_527_p N_A_M1000_g 0.0113543f $X=4.395 $Y=2.89 $X2=0 $Y2=0
cc_411 N_A_454_263#_c_459_n N_A_M1017_g 0.0141866f $X=6.3 $Y=2.13 $X2=0 $Y2=0
cc_412 N_A_454_263#_c_496_n N_A_M1013_g 0.0116908f $X=8.605 $Y=2.015 $X2=0 $Y2=0
cc_413 N_A_454_263#_c_496_n N_A_M1018_g 0.0118361f $X=8.605 $Y=2.015 $X2=0 $Y2=0
cc_414 N_A_454_263#_c_442_n N_A_c_699_n 0.00353071f $X=3.805 $Y=1.395 $X2=0
+ $Y2=0
cc_415 N_A_454_263#_c_443_n N_A_c_699_n 0.0124655f $X=3.805 $Y=1.855 $X2=0 $Y2=0
cc_416 N_A_454_263#_c_444_n N_A_c_699_n 0.0429443f $X=4.73 $Y=1.08 $X2=0 $Y2=0
cc_417 N_A_454_263#_c_525_p N_A_c_699_n 0.00718205f $X=4.195 $Y=1.94 $X2=0 $Y2=0
cc_418 N_A_454_263#_c_526_p N_A_c_699_n 0.0188722f $X=4.352 $Y=2.215 $X2=0 $Y2=0
cc_419 N_A_454_263#_c_536_p N_A_c_699_n 0.0113427f $X=5.18 $Y=2.13 $X2=0 $Y2=0
cc_420 N_A_454_263#_c_448_n N_A_c_699_n 0.0138444f $X=3.805 $Y=1.48 $X2=0 $Y2=0
cc_421 N_A_454_263#_c_450_n N_A_c_699_n 2.7171e-19 $X=3.67 $Y=1.48 $X2=0 $Y2=0
cc_422 N_A_454_263#_M1032_g N_A_c_700_n 0.0010743f $X=3.635 $Y=2.465 $X2=0 $Y2=0
cc_423 N_A_454_263#_c_442_n N_A_c_700_n 3.12545e-19 $X=3.805 $Y=1.395 $X2=0
+ $Y2=0
cc_424 N_A_454_263#_c_443_n N_A_c_700_n 7.17913e-19 $X=3.805 $Y=1.855 $X2=0
+ $Y2=0
cc_425 N_A_454_263#_c_444_n N_A_c_700_n 0.00520069f $X=4.73 $Y=1.08 $X2=0 $Y2=0
cc_426 N_A_454_263#_c_525_p N_A_c_700_n 0.00311017f $X=4.195 $Y=1.94 $X2=0 $Y2=0
cc_427 N_A_454_263#_c_526_p N_A_c_700_n 0.00144312f $X=4.352 $Y=2.215 $X2=0
+ $Y2=0
cc_428 N_A_454_263#_c_448_n N_A_c_700_n 0.00123361f $X=3.805 $Y=1.48 $X2=0 $Y2=0
cc_429 N_A_454_263#_c_450_n N_A_c_700_n 0.0186796f $X=3.67 $Y=1.48 $X2=0 $Y2=0
cc_430 N_A_454_263#_M1027_s N_A_c_713_n 0.00176773f $X=5.155 $Y=1.835 $X2=0
+ $Y2=0
cc_431 N_A_454_263#_c_444_n N_A_c_713_n 0.00670675f $X=4.73 $Y=1.08 $X2=0 $Y2=0
cc_432 N_A_454_263#_c_536_p N_A_c_713_n 0.025205f $X=5.18 $Y=2.13 $X2=0 $Y2=0
cc_433 N_A_454_263#_c_459_n N_A_c_713_n 3.06509e-19 $X=6.3 $Y=2.13 $X2=0 $Y2=0
cc_434 N_A_454_263#_c_551_p N_A_c_713_n 0.0135577f $X=5.295 $Y=2.21 $X2=0 $Y2=0
cc_435 N_A_454_263#_c_459_n N_A_c_714_n 0.0205938f $X=6.3 $Y=2.13 $X2=0 $Y2=0
cc_436 N_A_454_263#_c_459_n N_A_c_701_n 7.25369e-19 $X=6.3 $Y=2.13 $X2=0 $Y2=0
cc_437 N_A_454_263#_c_459_n A 0.0092222f $X=6.3 $Y=2.13 $X2=0 $Y2=0
cc_438 N_A_454_263#_c_496_n A 0.056163f $X=8.605 $Y=2.015 $X2=0 $Y2=0
cc_439 N_A_454_263#_c_461_n A 0.0126292f $X=6.385 $Y=2.015 $X2=0 $Y2=0
cc_440 N_A_454_263#_c_496_n N_A_c_703_n 0.00957374f $X=8.605 $Y=2.015 $X2=0
+ $Y2=0
cc_441 N_A_454_263#_c_459_n N_A_c_704_n 0.0272375f $X=6.3 $Y=2.13 $X2=0 $Y2=0
cc_442 N_A_454_263#_c_444_n N_B_M1001_g 0.0111613f $X=4.73 $Y=1.08 $X2=0 $Y2=0
cc_443 N_A_454_263#_c_495_n N_B_M1001_g 0.00131003f $X=4.825 $Y=0.77 $X2=0 $Y2=0
cc_444 N_A_454_263#_c_526_p N_B_M1007_g 0.00448516f $X=4.352 $Y=2.215 $X2=0
+ $Y2=0
cc_445 N_A_454_263#_c_536_p N_B_M1007_g 0.013052f $X=5.18 $Y=2.13 $X2=0 $Y2=0
cc_446 N_A_454_263#_c_444_n N_B_c_867_n 0.00271657f $X=4.73 $Y=1.08 $X2=0 $Y2=0
cc_447 N_A_454_263#_c_444_n N_B_M1002_g 0.0012953f $X=4.73 $Y=1.08 $X2=0 $Y2=0
cc_448 N_A_454_263#_c_495_n N_B_M1002_g 0.00131003f $X=4.825 $Y=0.77 $X2=0 $Y2=0
cc_449 N_A_454_263#_c_536_p N_B_M1027_g 0.0130502f $X=5.18 $Y=2.13 $X2=0 $Y2=0
cc_450 N_A_454_263#_c_496_n N_B_M1008_g 0.0116317f $X=8.605 $Y=2.015 $X2=0 $Y2=0
cc_451 N_A_454_263#_c_461_n N_B_M1008_g 0.0045098f $X=6.385 $Y=2.015 $X2=0 $Y2=0
cc_452 N_A_454_263#_M1004_g N_B_M1028_g 0.0324645f $X=8.915 $Y=2.465 $X2=0 $Y2=0
cc_453 N_A_454_263#_c_496_n N_B_M1028_g 0.0109855f $X=8.605 $Y=2.015 $X2=0 $Y2=0
cc_454 N_A_454_263#_c_445_n N_B_M1028_g 0.00405802f $X=8.69 $Y=1.93 $X2=0 $Y2=0
cc_455 N_A_454_263#_M1005_g N_B_M1029_g 0.0208299f $X=8.985 $Y=0.745 $X2=0 $Y2=0
cc_456 N_A_454_263#_c_451_n N_B_M1029_g 0.0118881f $X=9.005 $Y=1.4 $X2=0 $Y2=0
cc_457 N_A_454_263#_c_496_n N_B_c_876_n 0.00467301f $X=8.605 $Y=2.015 $X2=0
+ $Y2=0
cc_458 N_A_454_263#_c_444_n N_B_c_877_n 0.00894054f $X=4.73 $Y=1.08 $X2=0 $Y2=0
cc_459 N_A_454_263#_c_496_n N_B_c_882_n 0.00582151f $X=8.605 $Y=2.015 $X2=0
+ $Y2=0
cc_460 N_A_454_263#_c_445_n N_B_c_882_n 8.00128e-19 $X=8.69 $Y=1.93 $X2=0 $Y2=0
cc_461 N_A_454_263#_c_446_n N_B_c_882_n 0.00413325f $X=8.775 $Y=1.49 $X2=0 $Y2=0
cc_462 N_A_454_263#_c_451_n N_B_c_882_n 0.00566101f $X=9.005 $Y=1.4 $X2=0 $Y2=0
cc_463 N_A_454_263#_c_496_n B 0.0473799f $X=8.605 $Y=2.015 $X2=0 $Y2=0
cc_464 N_A_454_263#_c_445_n B 0.0135392f $X=8.69 $Y=1.93 $X2=0 $Y2=0
cc_465 N_A_454_263#_c_446_n B 0.0138521f $X=8.775 $Y=1.49 $X2=0 $Y2=0
cc_466 N_A_454_263#_c_451_n B 4.48481e-19 $X=9.005 $Y=1.4 $X2=0 $Y2=0
cc_467 N_A_454_263#_c_443_n N_VPWR_M1032_d 4.12128e-19 $X=3.805 $Y=1.855 $X2=0
+ $Y2=0
cc_468 N_A_454_263#_c_525_p N_VPWR_M1032_d 0.00750802f $X=4.195 $Y=1.94 $X2=0
+ $Y2=0
cc_469 N_A_454_263#_c_586_p N_VPWR_M1032_d 0.00243993f $X=3.89 $Y=1.94 $X2=0
+ $Y2=0
cc_470 N_A_454_263#_c_536_p N_VPWR_M1007_d 0.00418526f $X=5.18 $Y=2.13 $X2=0
+ $Y2=0
cc_471 N_A_454_263#_c_459_n N_VPWR_M1017_d 0.00498939f $X=6.3 $Y=2.13 $X2=0
+ $Y2=0
cc_472 N_A_454_263#_c_496_n N_VPWR_M1013_d 0.0123975f $X=8.605 $Y=2.015 $X2=0
+ $Y2=0
cc_473 N_A_454_263#_M1006_g N_VPWR_c_1034_n 0.00274882f $X=2.345 $Y=2.465 $X2=0
+ $Y2=0
cc_474 N_A_454_263#_M1012_g N_VPWR_c_1035_n 0.00151382f $X=2.775 $Y=2.465 $X2=0
+ $Y2=0
cc_475 N_A_454_263#_M1023_g N_VPWR_c_1035_n 0.00153321f $X=3.205 $Y=2.465 $X2=0
+ $Y2=0
cc_476 N_A_454_263#_M1023_g N_VPWR_c_1036_n 7.17104e-19 $X=3.205 $Y=2.465 $X2=0
+ $Y2=0
cc_477 N_A_454_263#_M1032_g N_VPWR_c_1036_n 0.0137841f $X=3.635 $Y=2.465 $X2=0
+ $Y2=0
cc_478 N_A_454_263#_c_492_n N_VPWR_c_1036_n 7.02467e-19 $X=3.72 $Y=1.48 $X2=0
+ $Y2=0
cc_479 N_A_454_263#_c_525_p N_VPWR_c_1036_n 0.010052f $X=4.195 $Y=1.94 $X2=0
+ $Y2=0
cc_480 N_A_454_263#_c_586_p N_VPWR_c_1036_n 0.0110448f $X=3.89 $Y=1.94 $X2=0
+ $Y2=0
cc_481 N_A_454_263#_c_526_p N_VPWR_c_1036_n 0.00157637f $X=4.352 $Y=2.215 $X2=0
+ $Y2=0
cc_482 N_A_454_263#_c_527_p N_VPWR_c_1036_n 0.0621415f $X=4.395 $Y=2.89 $X2=0
+ $Y2=0
cc_483 N_A_454_263#_c_536_p N_VPWR_c_1037_n 0.017285f $X=5.18 $Y=2.13 $X2=0
+ $Y2=0
cc_484 N_A_454_263#_c_459_n N_VPWR_c_1038_n 0.0219213f $X=6.3 $Y=2.13 $X2=0
+ $Y2=0
cc_485 N_A_454_263#_M1004_g N_VPWR_c_1074_n 0.00605603f $X=8.915 $Y=2.465 $X2=0
+ $Y2=0
cc_486 N_A_454_263#_M1004_g N_VPWR_c_1039_n 0.00821858f $X=8.915 $Y=2.465 $X2=0
+ $Y2=0
cc_487 N_A_454_263#_M1015_g N_VPWR_c_1039_n 0.00604308f $X=9.605 $Y=2.465 $X2=0
+ $Y2=0
cc_488 N_A_454_263#_M1004_g N_VPWR_c_1076_n 0.00269338f $X=8.915 $Y=2.465 $X2=0
+ $Y2=0
cc_489 N_A_454_263#_c_441_n N_VPWR_c_1076_n 5.67722e-19 $X=9.605 $Y=1.4 $X2=0
+ $Y2=0
cc_490 N_A_454_263#_M1006_g N_VPWR_c_1040_n 0.00585385f $X=2.345 $Y=2.465 $X2=0
+ $Y2=0
cc_491 N_A_454_263#_M1012_g N_VPWR_c_1040_n 0.0054895f $X=2.775 $Y=2.465 $X2=0
+ $Y2=0
cc_492 N_A_454_263#_M1023_g N_VPWR_c_1042_n 0.00585385f $X=3.205 $Y=2.465 $X2=0
+ $Y2=0
cc_493 N_A_454_263#_M1032_g N_VPWR_c_1042_n 0.00486043f $X=3.635 $Y=2.465 $X2=0
+ $Y2=0
cc_494 N_A_454_263#_c_527_p N_VPWR_c_1044_n 0.0166585f $X=4.395 $Y=2.89 $X2=0
+ $Y2=0
cc_495 N_A_454_263#_c_612_p N_VPWR_c_1046_n 0.0131621f $X=5.295 $Y=2.91 $X2=0
+ $Y2=0
cc_496 N_A_454_263#_M1004_g N_VPWR_c_1051_n 0.00427505f $X=8.915 $Y=2.465 $X2=0
+ $Y2=0
cc_497 N_A_454_263#_M1015_g N_VPWR_c_1052_n 0.00585385f $X=9.605 $Y=2.465 $X2=0
+ $Y2=0
cc_498 N_A_454_263#_M1000_s N_VPWR_c_1030_n 0.00311159f $X=4.255 $Y=1.835 $X2=0
+ $Y2=0
cc_499 N_A_454_263#_M1027_s N_VPWR_c_1030_n 0.00467071f $X=5.155 $Y=1.835 $X2=0
+ $Y2=0
cc_500 N_A_454_263#_M1006_g N_VPWR_c_1030_n 0.0105614f $X=2.345 $Y=2.465 $X2=0
+ $Y2=0
cc_501 N_A_454_263#_M1012_g N_VPWR_c_1030_n 0.00976568f $X=2.775 $Y=2.465 $X2=0
+ $Y2=0
cc_502 N_A_454_263#_M1023_g N_VPWR_c_1030_n 0.0105497f $X=3.205 $Y=2.465 $X2=0
+ $Y2=0
cc_503 N_A_454_263#_M1032_g N_VPWR_c_1030_n 0.00824727f $X=3.635 $Y=2.465 $X2=0
+ $Y2=0
cc_504 N_A_454_263#_M1004_g N_VPWR_c_1030_n 0.00782849f $X=8.915 $Y=2.465 $X2=0
+ $Y2=0
cc_505 N_A_454_263#_M1015_g N_VPWR_c_1030_n 0.0121382f $X=9.605 $Y=2.465 $X2=0
+ $Y2=0
cc_506 N_A_454_263#_c_527_p N_VPWR_c_1030_n 0.0117055f $X=4.395 $Y=2.89 $X2=0
+ $Y2=0
cc_507 N_A_454_263#_c_612_p N_VPWR_c_1030_n 0.00808656f $X=5.295 $Y=2.91 $X2=0
+ $Y2=0
cc_508 N_A_454_263#_M1006_g N_COUT_c_1264_n 0.00560122f $X=2.345 $Y=2.465 $X2=0
+ $Y2=0
cc_509 N_A_454_263#_M1016_g N_COUT_c_1264_n 0.00175596f $X=2.38 $Y=0.655 $X2=0
+ $Y2=0
cc_510 N_A_454_263#_M1019_g N_COUT_c_1264_n 0.00212407f $X=2.81 $Y=0.655 $X2=0
+ $Y2=0
cc_511 N_A_454_263#_c_440_n N_COUT_c_1264_n 0.0017266f $X=2.362 $Y=1.39 $X2=0
+ $Y2=0
cc_512 N_A_454_263#_c_492_n N_COUT_c_1264_n 0.0125935f $X=3.72 $Y=1.48 $X2=0
+ $Y2=0
cc_513 N_A_454_263#_c_449_n N_COUT_c_1264_n 0.00974233f $X=2.7 $Y=1.48 $X2=0
+ $Y2=0
cc_514 N_A_454_263#_c_450_n N_COUT_c_1264_n 0.00518775f $X=3.67 $Y=1.48 $X2=0
+ $Y2=0
cc_515 N_A_454_263#_M1016_g N_COUT_c_1274_n 7.63874e-19 $X=2.38 $Y=0.655 $X2=0
+ $Y2=0
cc_516 N_A_454_263#_M1019_g N_COUT_c_1274_n 0.0010349f $X=2.81 $Y=0.655 $X2=0
+ $Y2=0
cc_517 N_A_454_263#_M1019_g N_COUT_c_1265_n 0.0106504f $X=2.81 $Y=0.655 $X2=0
+ $Y2=0
cc_518 N_A_454_263#_M1030_g N_COUT_c_1265_n 0.00988766f $X=3.24 $Y=0.655 $X2=0
+ $Y2=0
cc_519 N_A_454_263#_M1033_g N_COUT_c_1265_n 0.00114899f $X=3.67 $Y=0.655 $X2=0
+ $Y2=0
cc_520 N_A_454_263#_c_492_n N_COUT_c_1265_n 0.0509053f $X=3.72 $Y=1.48 $X2=0
+ $Y2=0
cc_521 N_A_454_263#_c_442_n N_COUT_c_1265_n 0.00399949f $X=3.805 $Y=1.395 $X2=0
+ $Y2=0
cc_522 N_A_454_263#_c_494_n N_COUT_c_1265_n 0.00924569f $X=3.89 $Y=1.08 $X2=0
+ $Y2=0
cc_523 N_A_454_263#_c_450_n N_COUT_c_1265_n 0.00530199f $X=3.67 $Y=1.48 $X2=0
+ $Y2=0
cc_524 N_A_454_263#_M1012_g N_COUT_c_1268_n 0.0117234f $X=2.775 $Y=2.465 $X2=0
+ $Y2=0
cc_525 N_A_454_263#_M1023_g N_COUT_c_1268_n 0.0137909f $X=3.205 $Y=2.465 $X2=0
+ $Y2=0
cc_526 N_A_454_263#_M1032_g N_COUT_c_1268_n 7.14036e-19 $X=3.635 $Y=2.465 $X2=0
+ $Y2=0
cc_527 N_A_454_263#_c_492_n N_COUT_c_1268_n 0.0497925f $X=3.72 $Y=1.48 $X2=0
+ $Y2=0
cc_528 N_A_454_263#_c_443_n N_COUT_c_1268_n 0.00584052f $X=3.805 $Y=1.855 $X2=0
+ $Y2=0
cc_529 N_A_454_263#_c_450_n N_COUT_c_1268_n 0.00527005f $X=3.67 $Y=1.48 $X2=0
+ $Y2=0
cc_530 N_A_454_263#_M1030_g N_COUT_c_1278_n 0.0010349f $X=3.24 $Y=0.655 $X2=0
+ $Y2=0
cc_531 N_A_454_263#_M1033_g N_COUT_c_1278_n 0.00172265f $X=3.67 $Y=0.655 $X2=0
+ $Y2=0
cc_532 N_A_454_263#_M1016_g N_COUT_c_1266_n 0.00398558f $X=2.38 $Y=0.655 $X2=0
+ $Y2=0
cc_533 N_A_454_263#_c_449_n N_COUT_c_1266_n 0.00166574f $X=2.7 $Y=1.48 $X2=0
+ $Y2=0
cc_534 N_A_454_263#_M1006_g N_COUT_c_1269_n 0.00116014f $X=2.345 $Y=2.465 $X2=0
+ $Y2=0
cc_535 N_A_454_263#_M1012_g N_COUT_c_1269_n 0.00180758f $X=2.775 $Y=2.465 $X2=0
+ $Y2=0
cc_536 N_A_454_263#_c_449_n N_COUT_c_1269_n 3.24172e-19 $X=2.7 $Y=1.48 $X2=0
+ $Y2=0
cc_537 N_A_454_263#_M1012_g COUT 0.0146269f $X=2.775 $Y=2.465 $X2=0 $Y2=0
cc_538 N_A_454_263#_M1023_g COUT 7.18277e-19 $X=3.205 $Y=2.465 $X2=0 $Y2=0
cc_539 N_A_454_263#_c_496_n N_A_1367_367#_M1008_s 0.00355352f $X=8.605 $Y=2.015
+ $X2=-0.19 $Y2=-0.245
cc_540 N_A_454_263#_c_496_n N_A_1367_367#_M1018_s 0.00354935f $X=8.605 $Y=2.015
+ $X2=0 $Y2=0
cc_541 N_A_454_263#_c_444_n N_VGND_M1033_d 0.00153475f $X=4.73 $Y=1.08 $X2=0
+ $Y2=0
cc_542 N_A_454_263#_c_494_n N_VGND_M1033_d 4.62606e-19 $X=3.89 $Y=1.08 $X2=0
+ $Y2=0
cc_543 N_A_454_263#_M1016_g N_VGND_c_1364_n 0.00999083f $X=2.38 $Y=0.655 $X2=0
+ $Y2=0
cc_544 N_A_454_263#_M1019_g N_VGND_c_1364_n 5.67328e-19 $X=2.81 $Y=0.655 $X2=0
+ $Y2=0
cc_545 N_A_454_263#_M1016_g N_VGND_c_1365_n 6.26181e-19 $X=2.38 $Y=0.655 $X2=0
+ $Y2=0
cc_546 N_A_454_263#_M1019_g N_VGND_c_1365_n 0.0105363f $X=2.81 $Y=0.655 $X2=0
+ $Y2=0
cc_547 N_A_454_263#_M1030_g N_VGND_c_1365_n 0.0105376f $X=3.24 $Y=0.655 $X2=0
+ $Y2=0
cc_548 N_A_454_263#_M1033_g N_VGND_c_1365_n 6.26181e-19 $X=3.67 $Y=0.655 $X2=0
+ $Y2=0
cc_549 N_A_454_263#_M1030_g N_VGND_c_1366_n 6.06088e-19 $X=3.24 $Y=0.655 $X2=0
+ $Y2=0
cc_550 N_A_454_263#_M1033_g N_VGND_c_1366_n 0.00992688f $X=3.67 $Y=0.655 $X2=0
+ $Y2=0
cc_551 N_A_454_263#_c_444_n N_VGND_c_1366_n 0.00872962f $X=4.73 $Y=1.08 $X2=0
+ $Y2=0
cc_552 N_A_454_263#_c_494_n N_VGND_c_1366_n 0.00782853f $X=3.89 $Y=1.08 $X2=0
+ $Y2=0
cc_553 N_A_454_263#_M1016_g N_VGND_c_1371_n 0.00486043f $X=2.38 $Y=0.655 $X2=0
+ $Y2=0
cc_554 N_A_454_263#_M1019_g N_VGND_c_1371_n 0.00486043f $X=2.81 $Y=0.655 $X2=0
+ $Y2=0
cc_555 N_A_454_263#_M1030_g N_VGND_c_1373_n 0.00486043f $X=3.24 $Y=0.655 $X2=0
+ $Y2=0
cc_556 N_A_454_263#_M1033_g N_VGND_c_1373_n 0.00486043f $X=3.67 $Y=0.655 $X2=0
+ $Y2=0
cc_557 N_A_454_263#_M1005_g N_VGND_c_1380_n 0.0030414f $X=8.985 $Y=0.745 $X2=0
+ $Y2=0
cc_558 N_A_454_263#_M1026_g N_VGND_c_1380_n 0.0030414f $X=9.415 $Y=0.745 $X2=0
+ $Y2=0
cc_559 N_A_454_263#_M1001_d N_VGND_c_1381_n 0.00225465f $X=4.685 $Y=0.235 $X2=0
+ $Y2=0
cc_560 N_A_454_263#_M1016_g N_VGND_c_1381_n 0.00824727f $X=2.38 $Y=0.655 $X2=0
+ $Y2=0
cc_561 N_A_454_263#_M1019_g N_VGND_c_1381_n 0.00824727f $X=2.81 $Y=0.655 $X2=0
+ $Y2=0
cc_562 N_A_454_263#_M1030_g N_VGND_c_1381_n 0.00824727f $X=3.24 $Y=0.655 $X2=0
+ $Y2=0
cc_563 N_A_454_263#_M1033_g N_VGND_c_1381_n 0.00824727f $X=3.67 $Y=0.655 $X2=0
+ $Y2=0
cc_564 N_A_454_263#_M1005_g N_VGND_c_1381_n 0.00435814f $X=8.985 $Y=0.745 $X2=0
+ $Y2=0
cc_565 N_A_454_263#_M1026_g N_VGND_c_1381_n 0.00475975f $X=9.415 $Y=0.745 $X2=0
+ $Y2=0
cc_566 N_A_454_263#_c_444_n N_A_851_47#_M1020_d 0.0015892f $X=4.73 $Y=1.08
+ $X2=-0.19 $Y2=-0.245
cc_567 N_A_454_263#_M1001_d N_A_851_47#_c_1526_n 0.00329871f $X=4.685 $Y=0.235
+ $X2=0 $Y2=0
cc_568 N_A_454_263#_c_444_n N_A_851_47#_c_1526_n 0.00139391f $X=4.73 $Y=1.08
+ $X2=0 $Y2=0
cc_569 N_A_454_263#_c_495_n N_A_851_47#_c_1526_n 0.0119144f $X=4.825 $Y=0.77
+ $X2=0 $Y2=0
cc_570 N_A_454_263#_c_444_n N_A_851_47#_c_1527_n 0.0121806f $X=4.73 $Y=1.08
+ $X2=0 $Y2=0
cc_571 N_A_454_263#_M1005_g N_A_1284_65#_c_1564_n 4.83482e-19 $X=8.985 $Y=0.745
+ $X2=0 $Y2=0
cc_572 N_A_454_263#_c_446_n N_A_1284_65#_c_1564_n 0.00678298f $X=8.775 $Y=1.49
+ $X2=0 $Y2=0
cc_573 N_A_454_263#_c_447_n N_A_1284_65#_c_1564_n 0.00362918f $X=9.005 $Y=1.49
+ $X2=0 $Y2=0
cc_574 N_A_454_263#_c_451_n N_A_1284_65#_c_1564_n 4.01098e-19 $X=9.005 $Y=1.4
+ $X2=0 $Y2=0
cc_575 N_A_454_263#_M1005_g N_A_1284_65#_c_1555_n 0.00882974f $X=8.985 $Y=0.745
+ $X2=0 $Y2=0
cc_576 N_A_454_263#_M1026_g N_A_1284_65#_c_1555_n 0.0111245f $X=9.415 $Y=0.745
+ $X2=0 $Y2=0
cc_577 N_A_454_263#_M1026_g N_A_1284_65#_c_1557_n 0.0102713f $X=9.415 $Y=0.745
+ $X2=0 $Y2=0
cc_578 N_A_M1020_g N_B_M1001_g 0.0277254f $X=4.18 $Y=0.655 $X2=0 $Y2=0
cc_579 N_A_M1000_g N_B_M1007_g 0.0209603f $X=4.18 $Y=2.465 $X2=0 $Y2=0
cc_580 N_A_c_699_n N_B_M1007_g 0.0167613f $X=4.545 $Y=1.51 $X2=0 $Y2=0
cc_581 N_A_c_713_n N_B_M1007_g 5.44548e-19 $X=5.44 $Y=1.785 $X2=0 $Y2=0
cc_582 N_A_c_699_n N_B_c_867_n 0.00219562f $X=4.545 $Y=1.51 $X2=0 $Y2=0
cc_583 N_A_c_713_n N_B_c_867_n 0.00408241f $X=5.44 $Y=1.785 $X2=0 $Y2=0
cc_584 N_A_M1031_g N_B_M1002_g 0.019507f $X=5.51 $Y=0.655 $X2=0 $Y2=0
cc_585 N_A_c_699_n N_B_M1027_g 0.00196881f $X=4.545 $Y=1.51 $X2=0 $Y2=0
cc_586 N_A_c_713_n N_B_M1027_g 0.0106924f $X=5.44 $Y=1.785 $X2=0 $Y2=0
cc_587 N_A_c_714_n N_B_M1027_g 7.35015e-19 $X=5.605 $Y=1.51 $X2=0 $Y2=0
cc_588 N_A_c_701_n N_B_M1027_g 0.0264264f $X=5.605 $Y=1.51 $X2=0 $Y2=0
cc_589 A N_B_c_870_n 0.00788237f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_590 N_A_M1011_g N_B_c_871_n 0.0284604f $X=7.35 $Y=0.745 $X2=0 $Y2=0
cc_591 N_A_M1013_g N_B_M1008_g 0.0543479f $X=7.19 $Y=2.465 $X2=0 $Y2=0
cc_592 A N_B_M1008_g 0.0131404f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_593 N_A_c_705_n N_B_M1008_g 0.00446935f $X=7.037 $Y=1.587 $X2=0 $Y2=0
cc_594 N_A_c_706_n N_B_M1008_g 0.00307599f $X=6.12 $Y=1.727 $X2=0 $Y2=0
cc_595 N_A_M1018_g N_B_M1028_g 0.0544203f $X=7.89 $Y=2.465 $X2=0 $Y2=0
cc_596 N_A_M1024_g N_B_M1029_g 0.0130454f $X=7.78 $Y=0.745 $X2=0 $Y2=0
cc_597 N_A_c_699_n N_B_c_874_n 0.00419604f $X=4.545 $Y=1.51 $X2=0 $Y2=0
cc_598 N_A_c_700_n N_B_c_874_n 0.0213439f $X=4.16 $Y=1.51 $X2=0 $Y2=0
cc_599 N_A_c_703_n N_B_c_875_n 0.0219291f $X=7.78 $Y=1.51 $X2=0 $Y2=0
cc_600 N_A_M1011_g N_B_c_876_n 0.0116824f $X=7.35 $Y=0.745 $X2=0 $Y2=0
cc_601 A N_B_c_876_n 0.0231768f $X=6.875 $Y=1.58 $X2=0 $Y2=0
cc_602 N_A_c_703_n N_B_c_876_n 0.00756285f $X=7.78 $Y=1.51 $X2=0 $Y2=0
cc_603 N_A_c_705_n N_B_c_876_n 0.0360615f $X=7.037 $Y=1.587 $X2=0 $Y2=0
cc_604 N_A_M1031_g N_B_c_877_n 0.00421195f $X=5.51 $Y=0.655 $X2=0 $Y2=0
cc_605 N_A_c_699_n N_B_c_877_n 0.0121257f $X=4.545 $Y=1.51 $X2=0 $Y2=0
cc_606 N_A_c_713_n N_B_c_877_n 0.0256704f $X=5.44 $Y=1.785 $X2=0 $Y2=0
cc_607 N_A_c_714_n N_B_c_877_n 0.00691026f $X=5.605 $Y=1.51 $X2=0 $Y2=0
cc_608 N_A_M1031_g N_B_c_878_n 0.00693925f $X=5.51 $Y=0.655 $X2=0 $Y2=0
cc_609 N_A_c_701_n N_B_c_878_n 0.00632341f $X=5.605 $Y=1.51 $X2=0 $Y2=0
cc_610 N_A_c_706_n N_B_c_878_n 0.00788237f $X=6.12 $Y=1.727 $X2=0 $Y2=0
cc_611 N_A_M1031_g N_B_c_879_n 0.0114672f $X=5.51 $Y=0.655 $X2=0 $Y2=0
cc_612 N_A_c_713_n N_B_c_879_n 0.00699939f $X=5.44 $Y=1.785 $X2=0 $Y2=0
cc_613 N_A_c_714_n N_B_c_879_n 0.0236675f $X=5.605 $Y=1.51 $X2=0 $Y2=0
cc_614 N_A_c_701_n N_B_c_879_n 0.0045735f $X=5.605 $Y=1.51 $X2=0 $Y2=0
cc_615 N_A_c_704_n N_B_c_879_n 0.00933782f $X=5.973 $Y=1.727 $X2=0 $Y2=0
cc_616 N_A_M1031_g N_B_c_880_n 5.13818e-19 $X=5.51 $Y=0.655 $X2=0 $Y2=0
cc_617 N_A_c_706_n N_B_c_880_n 0.0182621f $X=6.12 $Y=1.727 $X2=0 $Y2=0
cc_618 N_A_M1031_g N_B_c_881_n 0.02081f $X=5.51 $Y=0.655 $X2=0 $Y2=0
cc_619 N_A_c_699_n N_B_c_881_n 0.00191037f $X=4.545 $Y=1.51 $X2=0 $Y2=0
cc_620 N_A_c_713_n N_B_c_881_n 0.00487979f $X=5.44 $Y=1.785 $X2=0 $Y2=0
cc_621 N_A_c_714_n N_B_c_881_n 6.67797e-19 $X=5.605 $Y=1.51 $X2=0 $Y2=0
cc_622 N_A_c_703_n N_B_c_882_n 0.016682f $X=7.78 $Y=1.51 $X2=0 $Y2=0
cc_623 N_A_M1011_g B 0.0019582f $X=7.35 $Y=0.745 $X2=0 $Y2=0
cc_624 N_A_M1024_g B 0.0141101f $X=7.78 $Y=0.745 $X2=0 $Y2=0
cc_625 N_A_M1018_g B 0.00453547f $X=7.89 $Y=2.465 $X2=0 $Y2=0
cc_626 N_A_c_717_n B 0.0159858f $X=7.21 $Y=1.51 $X2=0 $Y2=0
cc_627 N_A_c_703_n B 0.0307959f $X=7.78 $Y=1.51 $X2=0 $Y2=0
cc_628 N_A_c_713_n N_VPWR_M1007_d 0.00219904f $X=5.44 $Y=1.785 $X2=0 $Y2=0
cc_629 N_A_c_714_n N_VPWR_M1017_d 0.00150655f $X=5.605 $Y=1.51 $X2=0 $Y2=0
cc_630 N_A_c_704_n N_VPWR_M1017_d 0.0010459f $X=5.973 $Y=1.727 $X2=0 $Y2=0
cc_631 N_A_M1000_g N_VPWR_c_1036_n 0.00936229f $X=4.18 $Y=2.465 $X2=0 $Y2=0
cc_632 N_A_M1000_g N_VPWR_c_1037_n 5.1077e-19 $X=4.18 $Y=2.465 $X2=0 $Y2=0
cc_633 N_A_M1017_g N_VPWR_c_1037_n 6.21053e-19 $X=5.51 $Y=2.465 $X2=0 $Y2=0
cc_634 N_A_M1017_g N_VPWR_c_1038_n 0.0137168f $X=5.51 $Y=2.465 $X2=0 $Y2=0
cc_635 N_A_M1000_g N_VPWR_c_1044_n 0.00497452f $X=4.18 $Y=2.465 $X2=0 $Y2=0
cc_636 N_A_M1017_g N_VPWR_c_1046_n 0.00486043f $X=5.51 $Y=2.465 $X2=0 $Y2=0
cc_637 N_A_M1013_g N_VPWR_c_1050_n 0.00400841f $X=7.19 $Y=2.465 $X2=0 $Y2=0
cc_638 N_A_M1018_g N_VPWR_c_1051_n 0.00408154f $X=7.89 $Y=2.465 $X2=0 $Y2=0
cc_639 N_A_M1000_g N_VPWR_c_1030_n 0.0090882f $X=4.18 $Y=2.465 $X2=0 $Y2=0
cc_640 N_A_M1017_g N_VPWR_c_1030_n 0.0082726f $X=5.51 $Y=2.465 $X2=0 $Y2=0
cc_641 N_A_M1013_g N_VPWR_c_1030_n 0.00626381f $X=7.19 $Y=2.465 $X2=0 $Y2=0
cc_642 N_A_M1018_g N_VPWR_c_1030_n 0.00638276f $X=7.89 $Y=2.465 $X2=0 $Y2=0
cc_643 N_A_M1013_g N_VPWR_c_1056_n 0.00722687f $X=7.19 $Y=2.465 $X2=0 $Y2=0
cc_644 N_A_M1018_g N_VPWR_c_1056_n 0.00653806f $X=7.89 $Y=2.465 $X2=0 $Y2=0
cc_645 N_A_M1013_g N_A_1367_367#_c_1334_n 0.00786328f $X=7.19 $Y=2.465 $X2=0
+ $Y2=0
cc_646 N_A_M1018_g N_A_1367_367#_c_1334_n 0.00990242f $X=7.89 $Y=2.465 $X2=0
+ $Y2=0
cc_647 N_A_M1013_g N_A_1367_367#_c_1335_n 0.00695426f $X=7.19 $Y=2.465 $X2=0
+ $Y2=0
cc_648 N_A_M1018_g N_A_1367_367#_c_1335_n 7.5635e-19 $X=7.89 $Y=2.465 $X2=0
+ $Y2=0
cc_649 N_A_M1013_g N_A_1367_367#_c_1337_n 8.01371e-19 $X=7.19 $Y=2.465 $X2=0
+ $Y2=0
cc_650 N_A_M1018_g N_A_1367_367#_c_1337_n 0.00546488f $X=7.89 $Y=2.465 $X2=0
+ $Y2=0
cc_651 N_A_M1020_g N_VGND_c_1366_n 0.00612989f $X=4.18 $Y=0.655 $X2=0 $Y2=0
cc_652 N_A_M1031_g N_VGND_c_1367_n 0.00539551f $X=5.51 $Y=0.655 $X2=0 $Y2=0
cc_653 N_A_M1011_g N_VGND_c_1368_n 0.00295453f $X=7.35 $Y=0.745 $X2=0 $Y2=0
cc_654 N_A_M1020_g N_VGND_c_1375_n 0.0054778f $X=4.18 $Y=0.655 $X2=0 $Y2=0
cc_655 N_A_M1031_g N_VGND_c_1375_n 0.00585385f $X=5.51 $Y=0.655 $X2=0 $Y2=0
cc_656 N_A_M1011_g N_VGND_c_1379_n 0.00357893f $X=7.35 $Y=0.745 $X2=0 $Y2=0
cc_657 N_A_M1024_g N_VGND_c_1379_n 0.00305694f $X=7.78 $Y=0.745 $X2=0 $Y2=0
cc_658 N_A_M1020_g N_VGND_c_1381_n 0.0100836f $X=4.18 $Y=0.655 $X2=0 $Y2=0
cc_659 N_A_M1031_g N_VGND_c_1381_n 0.0119685f $X=5.51 $Y=0.655 $X2=0 $Y2=0
cc_660 N_A_M1011_g N_VGND_c_1381_n 0.00506653f $X=7.35 $Y=0.745 $X2=0 $Y2=0
cc_661 N_A_M1024_g N_VGND_c_1381_n 0.00390184f $X=7.78 $Y=0.745 $X2=0 $Y2=0
cc_662 N_A_M1011_g N_VGND_c_1385_n 3.97749e-19 $X=7.35 $Y=0.745 $X2=0 $Y2=0
cc_663 N_A_M1024_g N_VGND_c_1385_n 0.00881205f $X=7.78 $Y=0.745 $X2=0 $Y2=0
cc_664 N_A_M1020_g N_A_851_47#_c_1527_n 0.00624684f $X=4.18 $Y=0.655 $X2=0 $Y2=0
cc_665 N_A_M1011_g N_A_1284_65#_c_1552_n 8.89871e-19 $X=7.35 $Y=0.745 $X2=0
+ $Y2=0
cc_666 N_A_M1011_g N_A_1284_65#_c_1561_n 0.00925479f $X=7.35 $Y=0.745 $X2=0
+ $Y2=0
cc_667 N_A_M1011_g N_A_1284_65#_c_1554_n 0.00700473f $X=7.35 $Y=0.745 $X2=0
+ $Y2=0
cc_668 N_A_M1024_g N_A_1284_65#_c_1554_n 2.93294e-19 $X=7.78 $Y=0.745 $X2=0
+ $Y2=0
cc_669 N_A_M1024_g N_A_1284_65#_c_1563_n 0.010042f $X=7.78 $Y=0.745 $X2=0 $Y2=0
cc_670 N_A_M1011_g N_A_1284_65#_c_1577_n 6.01152e-19 $X=7.35 $Y=0.745 $X2=0
+ $Y2=0
cc_671 N_A_c_703_n N_A_1284_65#_c_1577_n 2.17324e-19 $X=7.78 $Y=1.51 $X2=0 $Y2=0
cc_672 N_A_M1024_g N_A_1284_65#_c_1578_n 0.00279126f $X=7.78 $Y=0.745 $X2=0
+ $Y2=0
cc_673 N_A_c_703_n N_A_1284_65#_c_1578_n 2.70821e-19 $X=7.78 $Y=1.51 $X2=0 $Y2=0
cc_674 N_B_M1007_g N_VPWR_c_1037_n 0.0108795f $X=4.61 $Y=2.465 $X2=0 $Y2=0
cc_675 N_B_M1027_g N_VPWR_c_1037_n 0.0104525f $X=5.08 $Y=2.465 $X2=0 $Y2=0
cc_676 N_B_M1027_g N_VPWR_c_1038_n 6.53292e-19 $X=5.08 $Y=2.465 $X2=0 $Y2=0
cc_677 N_B_M1028_g N_VPWR_c_1074_n 0.00105185f $X=8.32 $Y=2.465 $X2=0 $Y2=0
cc_678 N_B_M1007_g N_VPWR_c_1044_n 0.00564095f $X=4.61 $Y=2.465 $X2=0 $Y2=0
cc_679 N_B_M1027_g N_VPWR_c_1046_n 0.00564095f $X=5.08 $Y=2.465 $X2=0 $Y2=0
cc_680 N_B_M1008_g N_VPWR_c_1050_n 0.00551405f $X=6.76 $Y=2.465 $X2=0 $Y2=0
cc_681 N_B_M1028_g N_VPWR_c_1051_n 0.00552614f $X=8.32 $Y=2.465 $X2=0 $Y2=0
cc_682 N_B_M1007_g N_VPWR_c_1030_n 0.00957184f $X=4.61 $Y=2.465 $X2=0 $Y2=0
cc_683 N_B_M1027_g N_VPWR_c_1030_n 0.00950825f $X=5.08 $Y=2.465 $X2=0 $Y2=0
cc_684 N_B_M1008_g N_VPWR_c_1030_n 0.00745417f $X=6.76 $Y=2.465 $X2=0 $Y2=0
cc_685 N_B_M1028_g N_VPWR_c_1030_n 0.0105314f $X=8.32 $Y=2.465 $X2=0 $Y2=0
cc_686 N_B_M1008_g N_A_1367_367#_c_1335_n 0.00395016f $X=6.76 $Y=2.465 $X2=0
+ $Y2=0
cc_687 N_B_M1028_g N_A_1367_367#_c_1337_n 0.00433966f $X=8.32 $Y=2.465 $X2=0
+ $Y2=0
cc_688 N_B_c_876_n N_VGND_M1010_d 0.00344049f $X=7.555 $Y=1.17 $X2=0 $Y2=0
cc_689 N_B_c_879_n N_VGND_c_1367_n 0.01793f $X=5.98 $Y=1.215 $X2=0 $Y2=0
cc_690 N_B_c_871_n N_VGND_c_1368_n 0.00477543f $X=6.76 $Y=1.275 $X2=0 $Y2=0
cc_691 N_B_M1001_g N_VGND_c_1375_n 0.0035993f $X=4.61 $Y=0.655 $X2=0 $Y2=0
cc_692 N_B_M1002_g N_VGND_c_1375_n 0.00359951f $X=5.04 $Y=0.655 $X2=0 $Y2=0
cc_693 N_B_c_871_n N_VGND_c_1378_n 0.00359883f $X=6.76 $Y=1.275 $X2=0 $Y2=0
cc_694 N_B_M1029_g N_VGND_c_1380_n 0.00499542f $X=8.555 $Y=0.745 $X2=0 $Y2=0
cc_695 N_B_M1001_g N_VGND_c_1381_n 0.00537818f $X=4.61 $Y=0.655 $X2=0 $Y2=0
cc_696 N_B_M1002_g N_VGND_c_1381_n 0.0054719f $X=5.04 $Y=0.655 $X2=0 $Y2=0
cc_697 N_B_c_871_n N_VGND_c_1381_n 0.00557678f $X=6.76 $Y=1.275 $X2=0 $Y2=0
cc_698 N_B_M1029_g N_VGND_c_1381_n 0.0100189f $X=8.555 $Y=0.745 $X2=0 $Y2=0
cc_699 N_B_M1029_g N_VGND_c_1385_n 0.00348887f $X=8.555 $Y=0.745 $X2=0 $Y2=0
cc_700 N_B_M1001_g N_A_851_47#_c_1526_n 0.00822721f $X=4.61 $Y=0.655 $X2=0 $Y2=0
cc_701 N_B_M1002_g N_A_851_47#_c_1526_n 0.00839656f $X=5.04 $Y=0.655 $X2=0 $Y2=0
cc_702 N_B_M1001_g N_A_851_47#_c_1527_n 0.00601143f $X=4.61 $Y=0.655 $X2=0 $Y2=0
cc_703 N_B_M1002_g N_A_851_47#_c_1527_n 4.97379e-19 $X=5.04 $Y=0.655 $X2=0 $Y2=0
cc_704 N_B_M1001_g N_A_851_47#_c_1528_n 4.89636e-19 $X=4.61 $Y=0.655 $X2=0 $Y2=0
cc_705 N_B_M1002_g N_A_851_47#_c_1528_n 0.00523994f $X=5.04 $Y=0.655 $X2=0 $Y2=0
cc_706 N_B_c_877_n N_A_851_47#_c_1528_n 0.00507407f $X=5.09 $Y=1.17 $X2=0 $Y2=0
cc_707 N_B_c_879_n N_A_851_47#_c_1528_n 0.0054497f $X=5.98 $Y=1.215 $X2=0 $Y2=0
cc_708 N_B_c_881_n N_A_851_47#_c_1528_n 4.14065e-19 $X=5.06 $Y=1.34 $X2=0 $Y2=0
cc_709 N_B_c_876_n N_A_1284_65#_M1010_s 0.0020332f $X=7.555 $Y=1.17 $X2=-0.19
+ $Y2=-0.245
cc_710 N_B_c_876_n N_A_1284_65#_M1011_d 6.81095e-19 $X=7.555 $Y=1.17 $X2=0 $Y2=0
cc_711 B N_A_1284_65#_M1011_d 9.03142e-19 $X=7.92 $Y=1.665 $X2=0 $Y2=0
cc_712 N_B_c_871_n N_A_1284_65#_c_1552_n 0.00596972f $X=6.76 $Y=1.275 $X2=0
+ $Y2=0
cc_713 N_B_c_871_n N_A_1284_65#_c_1561_n 0.00925479f $X=6.76 $Y=1.275 $X2=0
+ $Y2=0
cc_714 N_B_c_876_n N_A_1284_65#_c_1561_n 0.0372793f $X=7.555 $Y=1.17 $X2=0 $Y2=0
cc_715 N_B_c_871_n N_A_1284_65#_c_1553_n 6.0125e-19 $X=6.76 $Y=1.275 $X2=0 $Y2=0
cc_716 N_B_c_876_n N_A_1284_65#_c_1553_n 0.0185689f $X=7.555 $Y=1.17 $X2=0 $Y2=0
cc_717 N_B_c_871_n N_A_1284_65#_c_1554_n 9.0852e-19 $X=6.76 $Y=1.275 $X2=0 $Y2=0
cc_718 B N_A_1284_65#_c_1563_n 0.00560145f $X=7.92 $Y=1.665 $X2=0 $Y2=0
cc_719 N_B_M1029_g N_A_1284_65#_c_1564_n 0.0153335f $X=8.555 $Y=0.745 $X2=0
+ $Y2=0
cc_720 N_B_c_882_n N_A_1284_65#_c_1564_n 0.00160857f $X=8.34 $Y=1.51 $X2=0 $Y2=0
cc_721 B N_A_1284_65#_c_1564_n 0.0175561f $X=7.92 $Y=1.665 $X2=0 $Y2=0
cc_722 N_B_M1029_g N_A_1284_65#_c_1556_n 5.63048e-19 $X=8.555 $Y=0.745 $X2=0
+ $Y2=0
cc_723 N_B_c_876_n N_A_1284_65#_c_1577_n 0.00723093f $X=7.555 $Y=1.17 $X2=0
+ $Y2=0
cc_724 B N_A_1284_65#_c_1577_n 0.0066542f $X=7.92 $Y=1.665 $X2=0 $Y2=0
cc_725 N_B_M1029_g N_A_1284_65#_c_1578_n 0.00132882f $X=8.555 $Y=0.745 $X2=0
+ $Y2=0
cc_726 B N_A_1284_65#_c_1578_n 0.00925818f $X=7.92 $Y=1.665 $X2=0 $Y2=0
cc_727 N_VPWR_c_1030_n N_SUM_M1003_d 0.00536646f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_728 N_VPWR_c_1030_n N_SUM_M1025_d 0.0041489f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_729 N_VPWR_M1003_s N_SUM_c_1209_n 9.24827e-19 $X=0.285 $Y=1.835 $X2=0 $Y2=0
cc_730 N_VPWR_c_1032_n N_SUM_c_1209_n 0.00890916f $X=0.41 $Y=2.18 $X2=0 $Y2=0
cc_731 N_VPWR_M1003_s N_SUM_c_1210_n 0.00175138f $X=0.285 $Y=1.835 $X2=0 $Y2=0
cc_732 N_VPWR_c_1032_n N_SUM_c_1210_n 0.0144736f $X=0.41 $Y=2.18 $X2=0 $Y2=0
cc_733 N_VPWR_c_1048_n N_SUM_c_1244_n 0.0124525f $X=1.105 $Y=3.33 $X2=0 $Y2=0
cc_734 N_VPWR_c_1030_n N_SUM_c_1244_n 0.00730901f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_735 N_VPWR_M1014_s N_SUM_c_1211_n 0.00176461f $X=1.13 $Y=1.835 $X2=0 $Y2=0
cc_736 N_VPWR_c_1033_n N_SUM_c_1211_n 0.0170777f $X=1.27 $Y=2.18 $X2=0 $Y2=0
cc_737 N_VPWR_c_1034_n N_SUM_c_1211_n 0.00208313f $X=2.13 $Y=1.975 $X2=0 $Y2=0
cc_738 N_VPWR_c_1049_n N_SUM_c_1249_n 0.0136943f $X=2 $Y=3.33 $X2=0 $Y2=0
cc_739 N_VPWR_c_1030_n N_SUM_c_1249_n 0.00866972f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_740 N_VPWR_c_1030_n N_COUT_M1006_s 0.00240953f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_741 N_VPWR_c_1030_n N_COUT_M1023_s 0.00380103f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_742 N_VPWR_M1012_d N_COUT_c_1268_n 0.00176461f $X=2.85 $Y=1.835 $X2=0 $Y2=0
cc_743 N_VPWR_c_1035_n N_COUT_c_1268_n 0.0135055f $X=2.99 $Y=2.26 $X2=0 $Y2=0
cc_744 N_VPWR_c_1042_n N_COUT_c_1316_n 0.0140491f $X=3.685 $Y=3.33 $X2=0 $Y2=0
cc_745 N_VPWR_c_1030_n N_COUT_c_1316_n 0.0090585f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_746 N_VPWR_c_1034_n N_COUT_c_1269_n 0.00208313f $X=2.13 $Y=1.975 $X2=0 $Y2=0
cc_747 N_VPWR_c_1040_n COUT 0.0171073f $X=2.895 $Y=3.33 $X2=0 $Y2=0
cc_748 N_VPWR_c_1030_n COUT 0.0114026f $X=9.84 $Y=3.33 $X2=0 $Y2=0
cc_749 N_VPWR_c_1030_n N_A_1367_367#_M1008_s 0.00239272f $X=9.84 $Y=3.33
+ $X2=-0.19 $Y2=-0.245
cc_750 N_VPWR_c_1030_n N_A_1367_367#_M1018_s 0.00238241f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_751 N_VPWR_M1013_d N_A_1367_367#_c_1334_n 0.011276f $X=7.265 $Y=1.835 $X2=0
+ $Y2=0
cc_752 N_VPWR_c_1050_n N_A_1367_367#_c_1334_n 0.00298563f $X=7.34 $Y=3.33 $X2=0
+ $Y2=0
cc_753 N_VPWR_c_1051_n N_A_1367_367#_c_1334_n 0.00476773f $X=8.95 $Y=3.33 $X2=0
+ $Y2=0
cc_754 N_VPWR_c_1030_n N_A_1367_367#_c_1334_n 0.0137709f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_755 N_VPWR_c_1056_n N_A_1367_367#_c_1334_n 0.0253897f $X=7.52 $Y=3.065 $X2=0
+ $Y2=0
cc_756 N_VPWR_c_1050_n N_A_1367_367#_c_1335_n 0.0113302f $X=7.34 $Y=3.33 $X2=0
+ $Y2=0
cc_757 N_VPWR_c_1030_n N_A_1367_367#_c_1335_n 0.0122846f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_758 N_VPWR_c_1056_n N_A_1367_367#_c_1335_n 3.93927e-19 $X=7.52 $Y=3.065 $X2=0
+ $Y2=0
cc_759 N_VPWR_c_1051_n N_A_1367_367#_c_1337_n 0.0105325f $X=8.95 $Y=3.33 $X2=0
+ $Y2=0
cc_760 N_VPWR_c_1030_n N_A_1367_367#_c_1337_n 0.011448f $X=9.84 $Y=3.33 $X2=0
+ $Y2=0
cc_761 N_VPWR_c_1056_n N_A_1367_367#_c_1337_n 5.70781e-19 $X=7.52 $Y=3.065 $X2=0
+ $Y2=0
cc_762 N_SUM_c_1211_n N_COUT_c_1269_n 0.00210944f $X=1.605 $Y=1.84 $X2=0 $Y2=0
cc_763 N_SUM_c_1204_n N_VGND_M1009_s 0.00129688f $X=0.78 $Y=1.13 $X2=-0.19
+ $Y2=-0.245
cc_764 N_SUM_c_1207_n N_VGND_M1009_s 0.00133631f $X=0.247 $Y=1.215 $X2=-0.19
+ $Y2=-0.245
cc_765 N_SUM_c_1205_n N_VGND_M1021_s 0.00180746f $X=1.64 $Y=1.13 $X2=0 $Y2=0
cc_766 N_SUM_c_1204_n N_VGND_c_1361_n 0.0117567f $X=0.78 $Y=1.13 $X2=0 $Y2=0
cc_767 N_SUM_c_1207_n N_VGND_c_1361_n 0.0112472f $X=0.247 $Y=1.215 $X2=0 $Y2=0
cc_768 N_SUM_c_1257_p N_VGND_c_1362_n 0.0124525f $X=0.875 $Y=0.42 $X2=0 $Y2=0
cc_769 N_SUM_c_1205_n N_VGND_c_1363_n 0.0163515f $X=1.64 $Y=1.13 $X2=0 $Y2=0
cc_770 N_SUM_c_1230_n N_VGND_c_1377_n 0.0124525f $X=1.735 $Y=0.42 $X2=0 $Y2=0
cc_771 N_SUM_M1009_d N_VGND_c_1381_n 0.00536646f $X=0.735 $Y=0.235 $X2=0 $Y2=0
cc_772 N_SUM_M1022_d N_VGND_c_1381_n 0.00536646f $X=1.595 $Y=0.235 $X2=0 $Y2=0
cc_773 N_SUM_c_1257_p N_VGND_c_1381_n 0.00730901f $X=0.875 $Y=0.42 $X2=0 $Y2=0
cc_774 N_SUM_c_1230_n N_VGND_c_1381_n 0.00730901f $X=1.735 $Y=0.42 $X2=0 $Y2=0
cc_775 N_COUT_c_1265_n N_VGND_M1019_d 0.0015943f $X=3.36 $Y=1.13 $X2=0 $Y2=0
cc_776 N_COUT_c_1274_n N_VGND_c_1365_n 0.022919f $X=2.595 $Y=0.42 $X2=0 $Y2=0
cc_777 N_COUT_c_1265_n N_VGND_c_1365_n 0.0146797f $X=3.36 $Y=1.13 $X2=0 $Y2=0
cc_778 N_COUT_c_1278_n N_VGND_c_1365_n 0.0230167f $X=3.455 $Y=0.42 $X2=0 $Y2=0
cc_779 N_COUT_c_1274_n N_VGND_c_1371_n 0.0124525f $X=2.595 $Y=0.42 $X2=0 $Y2=0
cc_780 N_COUT_c_1278_n N_VGND_c_1373_n 0.0124525f $X=3.455 $Y=0.42 $X2=0 $Y2=0
cc_781 N_COUT_M1016_s N_VGND_c_1381_n 0.00536646f $X=2.455 $Y=0.235 $X2=0 $Y2=0
cc_782 N_COUT_M1030_s N_VGND_c_1381_n 0.00536646f $X=3.315 $Y=0.235 $X2=0 $Y2=0
cc_783 N_COUT_c_1274_n N_VGND_c_1381_n 0.00730901f $X=2.595 $Y=0.42 $X2=0 $Y2=0
cc_784 N_COUT_c_1278_n N_VGND_c_1381_n 0.00730901f $X=3.455 $Y=0.42 $X2=0 $Y2=0
cc_785 N_VGND_c_1381_n N_A_851_47#_M1020_d 0.00223819f $X=9.84 $Y=0 $X2=-0.19
+ $Y2=-0.245
cc_786 N_VGND_c_1381_n N_A_851_47#_M1002_s 0.00256024f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_787 N_VGND_c_1375_n N_A_851_47#_c_1526_n 0.0289534f $X=5.605 $Y=0 $X2=0 $Y2=0
cc_788 N_VGND_c_1381_n N_A_851_47#_c_1526_n 0.019148f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_789 N_VGND_c_1375_n N_A_851_47#_c_1527_n 0.0177111f $X=5.605 $Y=0 $X2=0 $Y2=0
cc_790 N_VGND_c_1381_n N_A_851_47#_c_1527_n 0.0123216f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_791 N_VGND_c_1375_n N_A_851_47#_c_1528_n 0.0178402f $X=5.605 $Y=0 $X2=0 $Y2=0
cc_792 N_VGND_c_1381_n N_A_851_47#_c_1528_n 0.0125454f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_793 N_VGND_c_1367_n N_A_1284_65#_c_1552_n 0.014237f $X=5.725 $Y=0.38 $X2=0
+ $Y2=0
cc_794 N_VGND_c_1378_n N_A_1284_65#_c_1552_n 0.0121482f $X=6.89 $Y=0 $X2=0 $Y2=0
cc_795 N_VGND_c_1381_n N_A_1284_65#_c_1552_n 0.011788f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_796 N_VGND_M1010_d N_A_1284_65#_c_1561_n 0.00592763f $X=6.835 $Y=0.325 $X2=0
+ $Y2=0
cc_797 N_VGND_c_1368_n N_A_1284_65#_c_1561_n 0.021205f $X=7.055 $Y=0.45 $X2=0
+ $Y2=0
cc_798 N_VGND_c_1378_n N_A_1284_65#_c_1561_n 0.0020954f $X=6.89 $Y=0 $X2=0 $Y2=0
cc_799 N_VGND_c_1379_n N_A_1284_65#_c_1561_n 0.0020954f $X=7.83 $Y=0 $X2=0 $Y2=0
cc_800 N_VGND_c_1381_n N_A_1284_65#_c_1561_n 0.0097839f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_801 N_VGND_c_1367_n N_A_1284_65#_c_1553_n 0.0068814f $X=5.725 $Y=0.38 $X2=0
+ $Y2=0
cc_802 N_VGND_c_1368_n N_A_1284_65#_c_1554_n 0.0101973f $X=7.055 $Y=0.45 $X2=0
+ $Y2=0
cc_803 N_VGND_c_1379_n N_A_1284_65#_c_1554_n 0.0153719f $X=7.83 $Y=0 $X2=0 $Y2=0
cc_804 N_VGND_c_1381_n N_A_1284_65#_c_1554_n 0.00974941f $X=9.84 $Y=0 $X2=0
+ $Y2=0
cc_805 N_VGND_c_1385_n N_A_1284_65#_c_1554_n 0.0131874f $X=7.995 $Y=0.45 $X2=0
+ $Y2=0
cc_806 N_VGND_c_1379_n N_A_1284_65#_c_1563_n 0.00196814f $X=7.83 $Y=0 $X2=0
+ $Y2=0
cc_807 N_VGND_c_1381_n N_A_1284_65#_c_1563_n 0.00414053f $X=9.84 $Y=0 $X2=0
+ $Y2=0
cc_808 N_VGND_c_1385_n N_A_1284_65#_c_1563_n 0.00166021f $X=7.995 $Y=0.45 $X2=0
+ $Y2=0
cc_809 N_VGND_M1024_s N_A_1284_65#_c_1564_n 0.00846951f $X=7.855 $Y=0.325 $X2=0
+ $Y2=0
cc_810 N_VGND_c_1385_n N_A_1284_65#_c_1564_n 0.0181316f $X=7.995 $Y=0.45 $X2=0
+ $Y2=0
cc_811 N_VGND_c_1380_n N_A_1284_65#_c_1555_n 0.0659657f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_812 N_VGND_c_1381_n N_A_1284_65#_c_1555_n 0.0391244f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_813 N_VGND_c_1380_n N_A_1284_65#_c_1556_n 0.0128106f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_814 N_VGND_c_1381_n N_A_1284_65#_c_1556_n 0.0073517f $X=9.84 $Y=0 $X2=0 $Y2=0
cc_815 N_VGND_c_1385_n N_A_1284_65#_c_1556_n 0.00456606f $X=7.995 $Y=0.45 $X2=0
+ $Y2=0
cc_816 N_VGND_M1024_s N_A_1284_65#_c_1578_n 0.00727847f $X=7.855 $Y=0.325 $X2=0
+ $Y2=0
cc_817 N_VGND_c_1381_n N_A_1284_65#_c_1578_n 6.77079e-19 $X=9.84 $Y=0 $X2=0
+ $Y2=0
cc_818 N_VGND_c_1385_n N_A_1284_65#_c_1578_n 0.0138995f $X=7.995 $Y=0.45 $X2=0
+ $Y2=0
