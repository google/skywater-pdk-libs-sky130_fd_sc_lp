* File: sky130_fd_sc_lp__nand4bb_m.pex.spice
* Created: Wed Sep  2 10:07:08 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__NAND4BB_M%B_N 3 6 8 9 13 15
r34 13 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.53 $Y=1.45
+ $X2=0.53 $Y2=1.615
r35 13 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.53 $Y=1.45
+ $X2=0.53 $Y2=1.285
r36 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.53
+ $Y=1.45 $X2=0.53 $Y2=1.45
r37 9 14 6.88265 $w=3.58e-07 $l=2.15e-07 $layer=LI1_cond $X=0.625 $Y=1.665
+ $X2=0.625 $Y2=1.45
r38 8 14 4.96191 $w=3.58e-07 $l=1.55e-07 $layer=LI1_cond $X=0.625 $Y=1.295
+ $X2=0.625 $Y2=1.45
r39 6 16 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=0.54 $Y=2.225
+ $X2=0.54 $Y2=1.615
r40 3 15 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.475 $Y=0.965
+ $X2=0.475 $Y2=1.285
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4BB_M%D 3 6 8 9 10 16 18
c40 18 0 1.32534e-19 $X=1.07 $Y=1.285
r41 16 19 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.07 $Y=1.45
+ $X2=1.07 $Y2=1.615
r42 16 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.07 $Y=1.45
+ $X2=1.07 $Y2=1.285
r43 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.07
+ $Y=1.45 $X2=1.07 $Y2=1.45
r44 10 17 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=1.2 $Y=1.45 $X2=1.07
+ $Y2=1.45
r45 10 20 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.2 $Y=1.45 $X2=1.2
+ $Y2=1.285
r46 10 20 2.47914 $w=1.68e-07 $l=3.8e-08 $layer=LI1_cond $X=1.2 $Y=1.247 $X2=1.2
+ $Y2=1.285
r47 9 10 21.0075 $w=1.68e-07 $l=3.22e-07 $layer=LI1_cond $X=1.2 $Y=0.925 $X2=1.2
+ $Y2=1.247
r48 8 9 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=1.2 $Y=0.555 $X2=1.2
+ $Y2=0.925
r49 6 19 333.298 $w=1.5e-07 $l=6.5e-07 $layer=POLY_cond $X=1.16 $Y=2.265
+ $X2=1.16 $Y2=1.615
r50 3 18 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.16 $Y=0.965
+ $X2=1.16 $Y2=1.285
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4BB_M%C 3 6 8 9 10 15 17
c37 17 0 2.16919e-19 $X=1.61 $Y=1.285
r38 15 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.61 $Y=1.45
+ $X2=1.61 $Y2=1.615
r39 15 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.61 $Y=1.45
+ $X2=1.61 $Y2=1.285
r40 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.61
+ $Y=1.45 $X2=1.61 $Y2=1.45
r41 10 16 7.44286 $w=2.38e-07 $l=1.55e-07 $layer=LI1_cond $X=1.645 $Y=1.295
+ $X2=1.645 $Y2=1.45
r42 9 10 17.7668 $w=2.38e-07 $l=3.7e-07 $layer=LI1_cond $X=1.645 $Y=0.925
+ $X2=1.645 $Y2=1.295
r43 8 9 17.7668 $w=2.38e-07 $l=3.7e-07 $layer=LI1_cond $X=1.645 $Y=0.555
+ $X2=1.645 $Y2=0.925
r44 6 18 333.298 $w=1.5e-07 $l=6.5e-07 $layer=POLY_cond $X=1.59 $Y=2.265
+ $X2=1.59 $Y2=1.615
r45 3 17 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.52 $Y=0.965
+ $X2=1.52 $Y2=1.285
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4BB_M%A_27_151# 1 2 7 11 14 18 22 25 26 31 32
c56 22 0 1.32534e-19 $X=0.26 $Y=0.925
c57 11 0 5.80257e-20 $X=2.06 $Y=0.965
r58 32 36 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=0.575 $Y=2.94
+ $X2=0.575 $Y2=3.03
r59 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.575
+ $Y=2.94 $X2=0.575 $Y2=2.94
r60 28 31 7.29881 $w=2.98e-07 $l=1.9e-07 $layer=LI1_cond $X=0.385 $Y=2.925
+ $X2=0.575 $Y2=2.925
r61 25 27 3.68369 $w=4.53e-07 $l=1.05e-07 $layer=LI1_cond $X=0.322 $Y=2.29
+ $X2=0.322 $Y2=2.395
r62 25 26 7.67467 $w=4.53e-07 $l=1.05e-07 $layer=LI1_cond $X=0.322 $Y=2.29
+ $X2=0.322 $Y2=2.185
r63 19 22 4.22511 $w=2.08e-07 $l=8e-08 $layer=LI1_cond $X=0.18 $Y=0.925 $X2=0.26
+ $Y2=0.925
r64 18 28 0.126616 $w=3.3e-07 $l=1.5e-07 $layer=LI1_cond $X=0.385 $Y=2.775
+ $X2=0.385 $Y2=2.925
r65 18 27 13.2706 $w=3.28e-07 $l=3.8e-07 $layer=LI1_cond $X=0.385 $Y=2.775
+ $X2=0.385 $Y2=2.395
r66 15 19 1.9771 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=0.18 $Y=1.03 $X2=0.18
+ $Y2=0.925
r67 15 26 75.3529 $w=1.68e-07 $l=1.155e-06 $layer=LI1_cond $X=0.18 $Y=1.03
+ $X2=0.18 $Y2=2.185
r68 11 14 666.596 $w=1.5e-07 $l=1.3e-06 $layer=POLY_cond $X=2.06 $Y=0.965
+ $X2=2.06 $Y2=2.265
r69 9 14 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.06 $Y=2.955
+ $X2=2.06 $Y2=2.265
r70 8 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.74 $Y=3.03
+ $X2=0.575 $Y2=3.03
r71 7 9 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.985 $Y=3.03
+ $X2=2.06 $Y2=2.955
r72 7 8 638.394 $w=1.5e-07 $l=1.245e-06 $layer=POLY_cond $X=1.985 $Y=3.03
+ $X2=0.74 $Y2=3.03
r73 2 25 600 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_PDIFF $count=1 $X=0.2
+ $Y=2.015 $X2=0.325 $Y2=2.29
r74 1 22 182 $w=1.7e-07 $l=2.23942e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.755 $X2=0.26 $Y2=0.925
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4BB_M%A_469_125# 1 2 9 11 13 15 22 26 28
c51 28 0 1.6639e-20 $X=3.44 $Y=1.725
c52 15 0 1.96656e-19 $X=3.205 $Y=1.725
r53 24 28 6.26932 $w=2.6e-07 $l=2.24332e-07 $layer=LI1_cond $X=3.58 $Y=1.56
+ $X2=3.44 $Y2=1.725
r54 24 26 62.4593 $w=1.88e-07 $l=1.07e-06 $layer=LI1_cond $X=3.58 $Y=1.56
+ $X2=3.58 $Y2=0.49
r55 20 28 6.26932 $w=2.6e-07 $l=1.96914e-07 $layer=LI1_cond $X=3.37 $Y=1.89
+ $X2=3.44 $Y2=1.725
r56 20 22 10.826 $w=3.28e-07 $l=3.1e-07 $layer=LI1_cond $X=3.37 $Y=1.89 $X2=3.37
+ $Y2=2.2
r57 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.625
+ $Y=1.725 $X2=2.625 $Y2=1.725
r58 15 28 0.499868 $w=3.3e-07 $l=2.35e-07 $layer=LI1_cond $X=3.205 $Y=1.725
+ $X2=3.44 $Y2=1.725
r59 15 17 20.2551 $w=3.28e-07 $l=5.8e-07 $layer=LI1_cond $X=3.205 $Y=1.725
+ $X2=2.625 $Y2=1.725
r60 11 18 39.5078 $w=3.96e-07 $l=1.99825e-07 $layer=POLY_cond $X=2.49 $Y=1.89
+ $X2=2.567 $Y2=1.725
r61 11 13 192.287 $w=1.5e-07 $l=3.75e-07 $layer=POLY_cond $X=2.49 $Y=1.89
+ $X2=2.49 $Y2=2.265
r62 7 18 58.374 $w=3.96e-07 $l=3.86575e-07 $layer=POLY_cond $X=2.42 $Y=1.405
+ $X2=2.567 $Y2=1.725
r63 7 9 225.617 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=2.42 $Y=1.405 $X2=2.42
+ $Y2=0.965
r64 2 22 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=3.23
+ $Y=2.055 $X2=3.37 $Y2=2.2
r65 1 26 182 $w=1.7e-07 $l=3.17372e-07 $layer=licon1_NDIFF $count=1 $X=3.43
+ $Y=0.235 $X2=3.57 $Y2=0.49
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4BB_M%A_N 3 7 10 13 15 16 20
c33 20 0 2.13295e-19 $X=3.22 $Y=1
r34 20 23 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=3.242 $Y=1
+ $X2=3.242 $Y2=1.165
r35 20 22 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=3.242 $Y=1
+ $X2=3.242 $Y2=0.835
r36 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.22 $Y=1
+ $X2=3.22 $Y2=1
r37 16 21 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=3.17 $Y=1.295
+ $X2=3.17 $Y2=1
r38 15 21 3.20123 $w=2.68e-07 $l=7.5e-08 $layer=LI1_cond $X=3.17 $Y=0.925
+ $X2=3.17 $Y2=1
r39 11 13 102.553 $w=1.5e-07 $l=2e-07 $layer=POLY_cond $X=3.155 $Y=1.46
+ $X2=3.355 $Y2=1.46
r40 10 13 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.355 $Y=1.385
+ $X2=3.355 $Y2=1.46
r41 10 23 112.809 $w=1.5e-07 $l=2.2e-07 $layer=POLY_cond $X=3.355 $Y=1.385
+ $X2=3.355 $Y2=1.165
r42 7 22 199.979 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=3.355 $Y=0.445
+ $X2=3.355 $Y2=0.835
r43 1 11 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.155 $Y=1.535
+ $X2=3.155 $Y2=1.46
r44 1 3 374.319 $w=1.5e-07 $l=7.3e-07 $layer=POLY_cond $X=3.155 $Y=1.535
+ $X2=3.155 $Y2=2.265
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4BB_M%VPWR 1 2 3 10 11 14 18 23 24 26 27 28 37
+ 43 44 47
r51 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r52 44 48 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=2.64 $Y2=3.33
r53 43 44 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r54 41 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.87 $Y=3.33
+ $X2=2.705 $Y2=3.33
r55 41 43 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=2.87 $Y=3.33 $X2=3.6
+ $Y2=3.33
r56 40 48 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r57 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r58 37 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.54 $Y=3.33
+ $X2=2.705 $Y2=3.33
r59 37 39 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=2.54 $Y=3.33
+ $X2=2.16 $Y2=3.33
r60 35 36 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r61 32 36 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r62 31 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r63 28 40 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=2.16 $Y2=3.33
r64 28 36 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=1.68 $Y2=3.33
r65 26 35 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=1.72 $Y=3.33 $X2=1.68
+ $Y2=3.33
r66 26 27 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.72 $Y=3.33
+ $X2=1.805 $Y2=3.33
r67 25 39 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=1.89 $Y=3.33 $X2=2.16
+ $Y2=3.33
r68 25 27 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.89 $Y=3.33
+ $X2=1.805 $Y2=3.33
r69 23 31 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=0.91 $Y=3.33
+ $X2=0.72 $Y2=3.33
r70 23 24 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=0.91 $Y=3.33
+ $X2=1.005 $Y2=3.33
r71 22 35 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=1.1 $Y=3.33 $X2=1.68
+ $Y2=3.33
r72 22 24 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.1 $Y=3.33 $X2=1.005
+ $Y2=3.33
r73 16 47 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.705 $Y=3.245
+ $X2=2.705 $Y2=3.33
r74 16 18 31.9541 $w=3.28e-07 $l=9.15e-07 $layer=LI1_cond $X=2.705 $Y=3.245
+ $X2=2.705 $Y2=2.33
r75 12 27 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.805 $Y=3.245
+ $X2=1.805 $Y2=3.33
r76 12 14 59.6952 $w=1.68e-07 $l=9.15e-07 $layer=LI1_cond $X=1.805 $Y=3.245
+ $X2=1.805 $Y2=2.33
r77 11 24 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.005 $Y=3.245
+ $X2=1.005 $Y2=3.33
r78 10 21 13.2743 $w=2.79e-07 $l=3.13767e-07 $layer=LI1_cond $X=1.005 $Y=2.605
+ $X2=0.922 $Y2=2.33
r79 10 11 37.3589 $w=1.88e-07 $l=6.4e-07 $layer=LI1_cond $X=1.005 $Y=2.605
+ $X2=1.005 $Y2=3.245
r80 3 18 600 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=1 $X=2.565
+ $Y=2.055 $X2=2.705 $Y2=2.33
r81 2 14 600 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=1 $X=1.665
+ $Y=2.055 $X2=1.805 $Y2=2.33
r82 1 21 600 $w=1.7e-07 $l=4.16233e-07 $layer=licon1_PDIFF $count=1 $X=0.615
+ $Y=2.015 $X2=0.85 $Y2=2.33
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4BB_M%Y 1 2 3 12 14 15 16 19 23 24 25 36
c47 23 0 6.29215e-20 $X=2.16 $Y=1.665
c48 19 0 5.80257e-20 $X=2.75 $Y=1.05
c49 15 0 1.53998e-19 $X=2.36 $Y=1.13
r50 34 36 2.02183 $w=2.83e-07 $l=5e-08 $layer=LI1_cond $X=2.217 $Y=1.985
+ $X2=2.217 $Y2=2.035
r51 25 39 3.03274 $w=2.83e-07 $l=7.5e-08 $layer=LI1_cond $X=2.217 $Y=2.405
+ $X2=2.217 $Y2=2.33
r52 24 31 3.29812 $w=2.85e-07 $l=8.5e-08 $layer=LI1_cond $X=2.217 $Y=1.9
+ $X2=2.217 $Y2=1.815
r53 24 34 3.29812 $w=2.85e-07 $l=8.5e-08 $layer=LI1_cond $X=2.217 $Y=1.9
+ $X2=2.217 $Y2=1.985
r54 24 39 11.2414 $w=2.83e-07 $l=2.78e-07 $layer=LI1_cond $X=2.217 $Y=2.052
+ $X2=2.217 $Y2=2.33
r55 24 36 0.687422 $w=2.83e-07 $l=1.7e-08 $layer=LI1_cond $X=2.217 $Y=2.052
+ $X2=2.217 $Y2=2.035
r56 23 31 6.06549 $w=2.83e-07 $l=1.5e-07 $layer=LI1_cond $X=2.217 $Y=1.665
+ $X2=2.217 $Y2=1.815
r57 19 21 4.22511 $w=2.08e-07 $l=8e-08 $layer=LI1_cond $X=2.75 $Y=1.05 $X2=2.75
+ $Y2=1.13
r58 17 23 18.1965 $w=2.83e-07 $l=4.5e-07 $layer=LI1_cond $X=2.217 $Y=1.215
+ $X2=2.217 $Y2=1.665
r59 16 24 32.5468 $w=2.03e-07 $l=5.95e-07 $layer=LI1_cond $X=1.48 $Y=1.9
+ $X2=2.075 $Y2=1.9
r60 15 17 7.39867 $w=1.7e-07 $l=1.80566e-07 $layer=LI1_cond $X=2.36 $Y=1.13
+ $X2=2.217 $Y2=1.215
r61 14 21 1.9771 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=2.645 $Y=1.13
+ $X2=2.75 $Y2=1.13
r62 14 15 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=2.645 $Y=1.13
+ $X2=2.36 $Y2=1.13
r63 10 16 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=1.375 $Y=1.985
+ $X2=1.48 $Y2=1.9
r64 10 12 11.355 $w=2.08e-07 $l=2.15e-07 $layer=LI1_cond $X=1.375 $Y=1.985
+ $X2=1.375 $Y2=2.2
r65 3 39 600 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=1 $X=2.135
+ $Y=2.055 $X2=2.275 $Y2=2.33
r66 2 12 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.235
+ $Y=2.055 $X2=1.375 $Y2=2.2
r67 1 19 182 $w=1.7e-07 $l=4.02803e-07 $layer=licon1_NDIFF $count=1 $X=2.495
+ $Y=0.755 $X2=2.75 $Y2=1.05
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4BB_M%VGND 1 2 9 13 15 17 22 32 33 36 39
r38 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r39 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r40 33 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=3.12
+ $Y2=0
r41 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r42 30 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.305 $Y=0 $X2=3.14
+ $Y2=0
r43 30 32 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=3.305 $Y=0 $X2=3.6
+ $Y2=0
r44 29 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r45 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r46 26 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r47 25 28 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.64
+ $Y2=0
r48 25 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r49 23 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.935 $Y=0 $X2=0.77
+ $Y2=0
r50 23 25 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.935 $Y=0 $X2=1.2
+ $Y2=0
r51 22 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.975 $Y=0 $X2=3.14
+ $Y2=0
r52 22 28 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=2.975 $Y=0 $X2=2.64
+ $Y2=0
r53 20 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r54 19 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r55 17 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.605 $Y=0 $X2=0.77
+ $Y2=0
r56 17 19 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.605 $Y=0 $X2=0.24
+ $Y2=0
r57 15 29 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=2.64
+ $Y2=0
r58 15 26 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=1.2
+ $Y2=0
r59 11 39 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.14 $Y=0.085
+ $X2=3.14 $Y2=0
r60 11 13 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=3.14 $Y=0.085
+ $X2=3.14 $Y2=0.38
r61 7 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.77 $Y=0.085 $X2=0.77
+ $Y2=0
r62 7 9 28.4618 $w=3.28e-07 $l=8.15e-07 $layer=LI1_cond $X=0.77 $Y=0.085
+ $X2=0.77 $Y2=0.9
r63 2 13 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=3.015
+ $Y=0.235 $X2=3.14 $Y2=0.38
r64 1 9 182 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.755 $X2=0.77 $Y2=0.9
.ends

