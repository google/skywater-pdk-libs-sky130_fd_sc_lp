* File: sky130_fd_sc_lp__o22ai_1.pxi.spice
* Created: Wed Sep  2 10:20:35 2020
* 
x_PM_SKY130_FD_SC_LP__O22AI_1%B1 N_B1_c_45_n N_B1_M1003_g N_B1_M1007_g B1 B1
+ N_B1_c_48_n PM_SKY130_FD_SC_LP__O22AI_1%B1
x_PM_SKY130_FD_SC_LP__O22AI_1%B2 N_B2_M1004_g N_B2_M1005_g B2 N_B2_c_74_n
+ PM_SKY130_FD_SC_LP__O22AI_1%B2
x_PM_SKY130_FD_SC_LP__O22AI_1%A2 N_A2_c_108_n N_A2_M1001_g N_A2_M1002_g A2 A2
+ N_A2_c_111_n PM_SKY130_FD_SC_LP__O22AI_1%A2
x_PM_SKY130_FD_SC_LP__O22AI_1%A1 N_A1_M1000_g N_A1_M1006_g N_A1_c_146_n
+ N_A1_c_147_n A1 A1 N_A1_c_149_n PM_SKY130_FD_SC_LP__O22AI_1%A1
x_PM_SKY130_FD_SC_LP__O22AI_1%VPWR N_VPWR_M1007_s N_VPWR_M1000_d N_VPWR_c_176_n
+ N_VPWR_c_177_n N_VPWR_c_178_n VPWR N_VPWR_c_179_n N_VPWR_c_180_n
+ N_VPWR_c_175_n N_VPWR_c_182_n PM_SKY130_FD_SC_LP__O22AI_1%VPWR
x_PM_SKY130_FD_SC_LP__O22AI_1%Y N_Y_M1003_d N_Y_M1004_d N_Y_c_209_n N_Y_c_210_n
+ Y Y Y N_Y_c_211_n N_Y_c_207_n PM_SKY130_FD_SC_LP__O22AI_1%Y
x_PM_SKY130_FD_SC_LP__O22AI_1%A_27_69# N_A_27_69#_M1003_s N_A_27_69#_M1005_d
+ N_A_27_69#_M1006_d N_A_27_69#_c_239_n N_A_27_69#_c_240_n N_A_27_69#_c_241_n
+ N_A_27_69#_c_251_n N_A_27_69#_c_248_n N_A_27_69#_c_242_n N_A_27_69#_c_243_n
+ PM_SKY130_FD_SC_LP__O22AI_1%A_27_69#
x_PM_SKY130_FD_SC_LP__O22AI_1%VGND N_VGND_M1001_d VGND N_VGND_c_272_n
+ N_VGND_c_273_n N_VGND_c_274_n N_VGND_c_275_n PM_SKY130_FD_SC_LP__O22AI_1%VGND
cc_1 VNB N_B1_c_45_n 0.0191457f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.295
cc_2 VNB N_B1_M1007_g 0.00137316f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.465
cc_3 VNB B1 0.019656f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_4 VNB N_B1_c_48_n 0.0474479f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.46
cc_5 VNB N_B2_M1005_g 0.0200321f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_6 VNB B2 0.00381107f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_7 VNB N_B2_c_74_n 0.0267215f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.46
cc_8 VNB N_A2_c_108_n 0.0192131f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.295
cc_9 VNB N_A2_M1002_g 0.00130053f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.465
cc_10 VNB A2 0.0062341f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_11 VNB N_A2_c_111_n 0.0355497f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A1_M1000_g 0.00154482f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.765
cc_13 VNB N_A1_c_146_n 0.027236f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_14 VNB N_A1_c_147_n 0.0231063f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB A1 0.0319634f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.46
cc_16 VNB N_A1_c_149_n 0.0494327f $X=-0.19 $Y=-0.245 $X2=0.22 $Y2=1.46
cc_17 VNB N_VPWR_c_175_n 0.123877f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_Y_c_207_n 0.00291572f $X=-0.19 $Y=-0.245 $X2=0.22 $Y2=1.665
cc_19 VNB N_A_27_69#_c_239_n 0.0233858f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.46
cc_20 VNB N_A_27_69#_c_240_n 0.00537169f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.46
cc_21 VNB N_A_27_69#_c_241_n 0.00935084f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_27_69#_c_242_n 0.00742531f $X=-0.19 $Y=-0.245 $X2=0.22 $Y2=1.665
cc_23 VNB N_A_27_69#_c_243_n 0.0228642f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_VGND_c_272_n 0.0365787f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.465
cc_25 VNB N_VGND_c_273_n 0.0239188f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.46
cc_26 VNB N_VGND_c_274_n 0.189401f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_275_n 0.0179862f $X=-0.19 $Y=-0.245 $X2=0.22 $Y2=1.46
cc_28 VPB N_B1_M1007_g 0.0236813f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.465
cc_29 VPB B1 0.00680654f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_30 VPB N_B2_M1004_g 0.0211166f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.765
cc_31 VPB B2 0.00416097f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_32 VPB N_B2_c_74_n 0.00731574f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.46
cc_33 VPB N_A2_M1002_g 0.0215979f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.465
cc_34 VPB A2 0.00465001f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_35 VPB N_A1_M1000_g 0.0239242f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.765
cc_36 VPB A1 0.0241466f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.46
cc_37 VPB N_VPWR_c_176_n 0.0102032f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_38 VPB N_VPWR_c_177_n 0.0494649f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_39 VPB N_VPWR_c_178_n 0.048343f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_40 VPB N_VPWR_c_179_n 0.0420371f $X=-0.19 $Y=1.655 $X2=0.22 $Y2=1.46
cc_41 VPB N_VPWR_c_180_n 0.0183725f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_42 VPB N_VPWR_c_175_n 0.0610419f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_43 VPB N_VPWR_c_182_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_44 VPB N_Y_c_207_n 0.00132737f $X=-0.19 $Y=1.655 $X2=0.22 $Y2=1.665
cc_45 N_B1_M1007_g N_B2_M1004_g 0.059804f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_46 N_B1_c_45_n N_B2_M1005_g 0.0194746f $X=0.475 $Y=1.295 $X2=0 $Y2=0
cc_47 N_B1_c_48_n B2 3.24211e-19 $X=0.475 $Y=1.46 $X2=0 $Y2=0
cc_48 N_B1_c_48_n N_B2_c_74_n 0.059804f $X=0.475 $Y=1.46 $X2=0 $Y2=0
cc_49 N_B1_M1007_g N_VPWR_c_177_n 0.00623768f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_50 B1 N_VPWR_c_177_n 0.0228788f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_51 N_B1_c_48_n N_VPWR_c_177_n 0.0014231f $X=0.475 $Y=1.46 $X2=0 $Y2=0
cc_52 N_B1_M1007_g N_VPWR_c_179_n 0.0054895f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_53 N_B1_M1007_g N_VPWR_c_175_n 0.0106011f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_54 N_B1_c_45_n N_Y_c_209_n 0.00473852f $X=0.475 $Y=1.295 $X2=0 $Y2=0
cc_55 N_B1_c_45_n N_Y_c_210_n 0.00617052f $X=0.475 $Y=1.295 $X2=0 $Y2=0
cc_56 N_B1_M1007_g N_Y_c_211_n 0.0227669f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_57 N_B1_c_45_n N_Y_c_207_n 0.00345977f $X=0.475 $Y=1.295 $X2=0 $Y2=0
cc_58 N_B1_M1007_g N_Y_c_207_n 0.0103984f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_59 B1 N_Y_c_207_n 0.0388366f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_60 N_B1_c_48_n N_Y_c_207_n 0.00716372f $X=0.475 $Y=1.46 $X2=0 $Y2=0
cc_61 B1 N_A_27_69#_c_239_n 0.0228787f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_62 N_B1_c_48_n N_A_27_69#_c_239_n 0.0015566f $X=0.475 $Y=1.46 $X2=0 $Y2=0
cc_63 N_B1_c_45_n N_A_27_69#_c_240_n 0.0128219f $X=0.475 $Y=1.295 $X2=0 $Y2=0
cc_64 N_B1_c_45_n N_VGND_c_272_n 0.0029147f $X=0.475 $Y=1.295 $X2=0 $Y2=0
cc_65 N_B1_c_45_n N_VGND_c_274_n 0.00420739f $X=0.475 $Y=1.295 $X2=0 $Y2=0
cc_66 N_B2_M1005_g N_A2_c_108_n 0.024313f $X=0.905 $Y=0.765 $X2=-0.19 $Y2=-0.245
cc_67 N_B2_M1004_g N_A2_M1002_g 0.00643395f $X=0.835 $Y=2.465 $X2=0 $Y2=0
cc_68 B2 N_A2_M1002_g 4.26661e-19 $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_69 N_B2_c_74_n N_A2_M1002_g 0.00118578f $X=0.95 $Y=1.51 $X2=0 $Y2=0
cc_70 N_B2_M1005_g A2 6.29711e-19 $X=0.905 $Y=0.765 $X2=0 $Y2=0
cc_71 B2 A2 0.0330309f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_72 N_B2_c_74_n A2 3.38776e-19 $X=0.95 $Y=1.51 $X2=0 $Y2=0
cc_73 B2 N_A2_c_111_n 0.0021435f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_74 N_B2_c_74_n N_A2_c_111_n 0.0174657f $X=0.95 $Y=1.51 $X2=0 $Y2=0
cc_75 N_B2_M1004_g N_VPWR_c_179_n 0.00357668f $X=0.835 $Y=2.465 $X2=0 $Y2=0
cc_76 N_B2_M1004_g N_VPWR_c_175_n 0.00585628f $X=0.835 $Y=2.465 $X2=0 $Y2=0
cc_77 N_B2_M1005_g N_Y_c_209_n 0.00454205f $X=0.905 $Y=0.765 $X2=0 $Y2=0
cc_78 N_B2_M1005_g N_Y_c_210_n 0.00406561f $X=0.905 $Y=0.765 $X2=0 $Y2=0
cc_79 N_B2_c_74_n N_Y_c_210_n 0.00199286f $X=0.95 $Y=1.51 $X2=0 $Y2=0
cc_80 N_B2_M1004_g N_Y_c_211_n 0.0358388f $X=0.835 $Y=2.465 $X2=0 $Y2=0
cc_81 B2 N_Y_c_211_n 0.0326455f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_82 N_B2_c_74_n N_Y_c_211_n 0.00117633f $X=0.95 $Y=1.51 $X2=0 $Y2=0
cc_83 N_B2_M1005_g N_Y_c_207_n 0.002587f $X=0.905 $Y=0.765 $X2=0 $Y2=0
cc_84 B2 N_Y_c_207_n 0.0309629f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_85 N_B2_c_74_n N_Y_c_207_n 0.00558565f $X=0.95 $Y=1.51 $X2=0 $Y2=0
cc_86 N_B2_M1005_g N_A_27_69#_c_240_n 0.0120858f $X=0.905 $Y=0.765 $X2=0 $Y2=0
cc_87 B2 N_A_27_69#_c_248_n 0.0136578f $X=1.115 $Y=1.58 $X2=0 $Y2=0
cc_88 N_B2_c_74_n N_A_27_69#_c_248_n 0.00189079f $X=0.95 $Y=1.51 $X2=0 $Y2=0
cc_89 N_B2_M1005_g N_VGND_c_272_n 0.0029147f $X=0.905 $Y=0.765 $X2=0 $Y2=0
cc_90 N_B2_M1005_g N_VGND_c_274_n 0.00403238f $X=0.905 $Y=0.765 $X2=0 $Y2=0
cc_91 N_B2_M1005_g N_VGND_c_275_n 3.53401e-19 $X=0.905 $Y=0.765 $X2=0 $Y2=0
cc_92 N_A2_M1002_g N_A1_M1000_g 0.057908f $X=1.63 $Y=2.465 $X2=0 $Y2=0
cc_93 A2 N_A1_c_146_n 0.00365516f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_94 N_A2_c_111_n N_A1_c_146_n 0.057908f $X=1.63 $Y=1.46 $X2=0 $Y2=0
cc_95 N_A2_c_108_n N_A1_c_147_n 0.0119266f $X=1.4 $Y=1.295 $X2=0 $Y2=0
cc_96 A2 N_A1_c_147_n 3.61226e-19 $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_97 N_A2_c_108_n A1 2.53397e-19 $X=1.4 $Y=1.295 $X2=0 $Y2=0
cc_98 A2 A1 0.0297204f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_99 N_A2_c_111_n A1 2.98809e-19 $X=1.63 $Y=1.46 $X2=0 $Y2=0
cc_100 N_A2_M1002_g N_VPWR_c_178_n 0.00436267f $X=1.63 $Y=2.465 $X2=0 $Y2=0
cc_101 N_A2_M1002_g N_VPWR_c_179_n 0.00518588f $X=1.63 $Y=2.465 $X2=0 $Y2=0
cc_102 N_A2_M1002_g N_VPWR_c_175_n 0.00978465f $X=1.63 $Y=2.465 $X2=0 $Y2=0
cc_103 N_A2_c_108_n N_Y_c_210_n 6.42044e-19 $X=1.4 $Y=1.295 $X2=0 $Y2=0
cc_104 N_A2_M1002_g N_Y_c_211_n 0.0226876f $X=1.63 $Y=2.465 $X2=0 $Y2=0
cc_105 A2 N_Y_c_211_n 0.00956873f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_106 N_A2_c_111_n N_Y_c_211_n 0.0059224f $X=1.63 $Y=1.46 $X2=0 $Y2=0
cc_107 N_A2_c_108_n N_A_27_69#_c_240_n 0.00122813f $X=1.4 $Y=1.295 $X2=0 $Y2=0
cc_108 N_A2_c_108_n N_A_27_69#_c_251_n 0.0191868f $X=1.4 $Y=1.295 $X2=0 $Y2=0
cc_109 A2 N_A_27_69#_c_251_n 0.0229055f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_110 N_A2_c_111_n N_A_27_69#_c_251_n 0.00118005f $X=1.63 $Y=1.46 $X2=0 $Y2=0
cc_111 N_A2_c_108_n N_VGND_c_272_n 0.00401871f $X=1.4 $Y=1.295 $X2=0 $Y2=0
cc_112 N_A2_c_108_n N_VGND_c_274_n 0.00778525f $X=1.4 $Y=1.295 $X2=0 $Y2=0
cc_113 N_A2_c_108_n N_VGND_c_275_n 0.00944302f $X=1.4 $Y=1.295 $X2=0 $Y2=0
cc_114 N_A1_M1000_g N_VPWR_c_178_n 0.028715f $X=1.99 $Y=2.465 $X2=0 $Y2=0
cc_115 N_A1_c_146_n N_VPWR_c_178_n 0.00158919f $X=2.08 $Y=1.46 $X2=0 $Y2=0
cc_116 A1 N_VPWR_c_178_n 0.0243957f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_117 N_A1_M1000_g N_VPWR_c_179_n 0.00486043f $X=1.99 $Y=2.465 $X2=0 $Y2=0
cc_118 N_A1_M1000_g N_VPWR_c_175_n 0.00818711f $X=1.99 $Y=2.465 $X2=0 $Y2=0
cc_119 N_A1_M1000_g N_Y_c_211_n 0.00319849f $X=1.99 $Y=2.465 $X2=0 $Y2=0
cc_120 N_A1_c_146_n N_A_27_69#_c_251_n 0.00544064f $X=2.08 $Y=1.46 $X2=0 $Y2=0
cc_121 N_A1_c_147_n N_A_27_69#_c_251_n 0.0133695f $X=2.08 $Y=1.295 $X2=0 $Y2=0
cc_122 A1 N_A_27_69#_c_251_n 0.0140335f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_123 A1 N_A_27_69#_c_242_n 0.0229944f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_124 N_A1_c_149_n N_A_27_69#_c_242_n 0.00162655f $X=2.5 $Y=1.46 $X2=0 $Y2=0
cc_125 N_A1_c_147_n N_A_27_69#_c_243_n 0.00189935f $X=2.08 $Y=1.295 $X2=0 $Y2=0
cc_126 N_A1_c_147_n N_VGND_c_273_n 0.00401871f $X=2.08 $Y=1.295 $X2=0 $Y2=0
cc_127 N_A1_c_147_n N_VGND_c_274_n 0.00799701f $X=2.08 $Y=1.295 $X2=0 $Y2=0
cc_128 N_A1_c_147_n N_VGND_c_275_n 0.0124591f $X=2.08 $Y=1.295 $X2=0 $Y2=0
cc_129 N_VPWR_c_175_n A_110_367# 0.00168875f $X=2.64 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_130 N_VPWR_c_175_n N_Y_M1004_d 0.00526662f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_131 N_VPWR_c_178_n N_Y_c_211_n 0.0421251f $X=2.205 $Y=2.005 $X2=0 $Y2=0
cc_132 N_VPWR_c_179_n N_Y_c_211_n 0.0669719f $X=2.04 $Y=3.33 $X2=0 $Y2=0
cc_133 N_VPWR_c_175_n N_Y_c_211_n 0.0405719f $X=2.64 $Y=3.33 $X2=0 $Y2=0
cc_134 N_VPWR_c_175_n A_341_367# 0.00899413f $X=2.64 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_135 A_110_367# N_Y_c_211_n 0.00129957f $X=0.55 $Y=1.835 $X2=2.04 $Y2=3.33
cc_136 A_110_367# N_Y_c_207_n 4.95691e-19 $X=0.55 $Y=1.835 $X2=0.355 $Y2=3.33
cc_137 N_Y_M1003_d N_A_27_69#_c_240_n 0.00176461f $X=0.55 $Y=0.345 $X2=0 $Y2=0
cc_138 N_Y_c_209_n N_A_27_69#_c_240_n 0.0158879f $X=0.69 $Y=0.695 $X2=0 $Y2=0
cc_139 N_A_27_69#_c_251_n N_VGND_M1001_d 0.017198f $X=2.29 $Y=0.955 $X2=-0.19
+ $Y2=-0.245
cc_140 N_A_27_69#_c_240_n N_VGND_c_272_n 0.0605088f $X=1.025 $Y=0.34 $X2=0 $Y2=0
cc_141 N_A_27_69#_c_241_n N_VGND_c_272_n 0.0186386f $X=0.355 $Y=0.34 $X2=0 $Y2=0
cc_142 N_A_27_69#_c_243_n N_VGND_c_273_n 0.0128398f $X=2.385 $Y=0.49 $X2=0 $Y2=0
cc_143 N_A_27_69#_c_240_n N_VGND_c_274_n 0.0337311f $X=1.025 $Y=0.34 $X2=0 $Y2=0
cc_144 N_A_27_69#_c_241_n N_VGND_c_274_n 0.0101082f $X=0.355 $Y=0.34 $X2=0 $Y2=0
cc_145 N_A_27_69#_c_243_n N_VGND_c_274_n 0.00968545f $X=2.385 $Y=0.49 $X2=0
+ $Y2=0
cc_146 N_A_27_69#_c_240_n N_VGND_c_275_n 0.0112909f $X=1.025 $Y=0.34 $X2=0 $Y2=0
cc_147 N_A_27_69#_c_251_n N_VGND_c_275_n 0.0447396f $X=2.29 $Y=0.955 $X2=0 $Y2=0
cc_148 N_A_27_69#_c_243_n N_VGND_c_275_n 0.0164418f $X=2.385 $Y=0.49 $X2=0 $Y2=0
