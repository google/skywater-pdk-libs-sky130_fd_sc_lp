* File: sky130_fd_sc_lp__o41ai_0.pex.spice
* Created: Fri Aug 28 11:20:01 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O41AI_0%B1 2 7 11 12 13 14 15 16 17 22 24
c44 14 0 2.76886e-21 $X=0.86 $Y=2.265
c45 13 0 7.63037e-20 $X=0.86 $Y=2.115
c46 2 0 4.48098e-20 $X=0.74 $Y=1.26
r47 22 25 4.07001 $w=5.75e-07 $l=1.5e-08 $layer=POLY_cond $X=0.802 $Y=0.98
+ $X2=0.802 $Y2=0.995
r48 22 24 48.7424 $w=5.75e-07 $l=1.65e-07 $layer=POLY_cond $X=0.802 $Y=0.98
+ $X2=0.802 $Y2=0.815
r49 16 17 14.2135 $w=2.98e-07 $l=3.7e-07 $layer=LI1_cond $X=0.745 $Y=1.295
+ $X2=0.745 $Y2=1.665
r50 15 16 14.2135 $w=2.98e-07 $l=3.7e-07 $layer=LI1_cond $X=0.745 $Y=0.925
+ $X2=0.745 $Y2=1.295
r51 15 22 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.68
+ $Y=0.98 $X2=0.68 $Y2=0.98
r52 13 14 45.0833 $w=2.7e-07 $l=1.5e-07 $layer=POLY_cond $X=0.86 $Y=2.115
+ $X2=0.86 $Y2=2.265
r53 12 13 139.969 $w=2.7e-07 $l=6.3e-07 $layer=POLY_cond $X=0.83 $Y=1.485
+ $X2=0.83 $Y2=2.115
r54 11 24 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.015 $Y=0.495
+ $X2=1.015 $Y2=0.815
r55 7 14 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=0.95 $Y=2.735 $X2=0.95
+ $Y2=2.265
r56 2 12 36.6371 $w=4.5e-07 $l=2.25e-07 $layer=POLY_cond $X=0.74 $Y=1.26
+ $X2=0.74 $Y2=1.485
r57 2 25 32.7513 $w=4.5e-07 $l=2.65e-07 $layer=POLY_cond $X=0.74 $Y=1.26
+ $X2=0.74 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_LP__O41AI_0%A4 2 5 9 11 12 16
c45 11 0 3.19103e-21 $X=1.2 $Y=1.295
r46 16 18 46.3655 $w=3.45e-07 $l=1.65e-07 $layer=POLY_cond $X=1.347 $Y=1.37
+ $X2=1.347 $Y2=1.205
r47 16 17 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.34
+ $Y=1.37 $X2=1.34 $Y2=1.37
r48 12 17 9.44363 $w=3.58e-07 $l=2.95e-07 $layer=LI1_cond $X=1.245 $Y=1.665
+ $X2=1.245 $Y2=1.37
r49 11 17 2.40092 $w=3.58e-07 $l=7.5e-08 $layer=LI1_cond $X=1.245 $Y=1.295
+ $X2=1.245 $Y2=1.37
r50 9 18 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=1.445 $Y=0.495
+ $X2=1.445 $Y2=1.205
r51 3 5 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.38 $Y=2.27 $X2=1.38
+ $Y2=2.735
r52 2 3 103.13 $w=2.65e-07 $l=5.83267e-07 $layer=POLY_cond $X=1.347 $Y=1.703
+ $X2=1.38 $Y2=2.27
r53 1 16 1.17081 $w=3.45e-07 $l=7e-09 $layer=POLY_cond $X=1.347 $Y=1.377
+ $X2=1.347 $Y2=1.37
r54 1 2 54.5263 $w=3.45e-07 $l=3.26e-07 $layer=POLY_cond $X=1.347 $Y=1.377
+ $X2=1.347 $Y2=1.703
.ends

.subckt PM_SKY130_FD_SC_LP__O41AI_0%A3 1 3 7 11 12 13 14 15 16 25 36 39
c50 25 0 9.77123e-20 $X=1.895 $Y=1.375
c51 14 0 7.90725e-20 $X=1.595 $Y=1.95
c52 7 0 5.16718e-20 $X=1.97 $Y=0.495
c53 3 0 1.12009e-19 $X=1.895 $Y=2.735
r54 37 39 1.70868 $w=5.58e-07 $l=8e-08 $layer=LI1_cond $X=1.78 $Y=2.325 $X2=1.78
+ $Y2=2.405
r55 36 45 0.257221 $w=4.63e-07 $l=1e-08 $layer=LI1_cond $X=1.827 $Y=2.035
+ $X2=1.827 $Y2=2.045
r56 25 26 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.895
+ $Y=1.375 $X2=1.895 $Y2=1.375
r57 15 37 0.0640756 $w=5.58e-07 $l=3e-09 $layer=LI1_cond $X=1.78 $Y=2.322
+ $X2=1.78 $Y2=2.325
r58 15 16 7.85994 $w=5.58e-07 $l=3.68e-07 $layer=LI1_cond $X=1.78 $Y=2.407
+ $X2=1.78 $Y2=2.775
r59 15 39 0.0427171 $w=5.58e-07 $l=2e-09 $layer=LI1_cond $X=1.78 $Y=2.407
+ $X2=1.78 $Y2=2.405
r60 14 15 5.12605 $w=5.58e-07 $l=2.4e-07 $layer=LI1_cond $X=1.78 $Y=2.082
+ $X2=1.78 $Y2=2.322
r61 14 45 1.16982 $w=5.58e-07 $l=3.7e-08 $layer=LI1_cond $X=1.78 $Y=2.082
+ $X2=1.78 $Y2=2.045
r62 14 36 0.97744 $w=4.63e-07 $l=3.8e-08 $layer=LI1_cond $X=1.827 $Y=1.997
+ $X2=1.827 $Y2=2.035
r63 13 14 8.53974 $w=4.63e-07 $l=3.32e-07 $layer=LI1_cond $X=1.827 $Y=1.665
+ $X2=1.827 $Y2=1.997
r64 13 26 7.45941 $w=4.63e-07 $l=2.9e-07 $layer=LI1_cond $X=1.827 $Y=1.665
+ $X2=1.827 $Y2=1.375
r65 12 26 2.05777 $w=4.63e-07 $l=8e-08 $layer=LI1_cond $X=1.827 $Y=1.295
+ $X2=1.827 $Y2=1.375
r66 11 25 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.895 $Y=1.715
+ $X2=1.895 $Y2=1.375
r67 10 25 43.7316 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.895 $Y=1.21
+ $X2=1.895 $Y2=1.375
r68 7 10 366.628 $w=1.5e-07 $l=7.15e-07 $layer=POLY_cond $X=1.97 $Y=0.495
+ $X2=1.97 $Y2=1.21
r69 1 11 37.5318 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.895 $Y=1.88
+ $X2=1.895 $Y2=1.715
r70 1 3 438.415 $w=1.5e-07 $l=8.55e-07 $layer=POLY_cond $X=1.895 $Y=1.88
+ $X2=1.895 $Y2=2.735
.ends

.subckt PM_SKY130_FD_SC_LP__O41AI_0%A2 1 5 9 13 14 15 16 17 18 23
c47 16 0 4.84808e-20 $X=2.64 $Y=1.295
c48 13 0 2.88954e-20 $X=2.435 $Y=1.21
r49 23 24 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.435
+ $Y=1.375 $X2=2.435 $Y2=1.375
r50 17 18 9.31682 $w=4.73e-07 $l=3.7e-07 $layer=LI1_cond $X=2.507 $Y=1.665
+ $X2=2.507 $Y2=2.035
r51 17 24 7.30237 $w=4.73e-07 $l=2.9e-07 $layer=LI1_cond $X=2.507 $Y=1.665
+ $X2=2.507 $Y2=1.375
r52 16 24 2.01445 $w=4.73e-07 $l=8e-08 $layer=LI1_cond $X=2.507 $Y=1.295
+ $X2=2.507 $Y2=1.375
r53 14 23 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.435 $Y=1.715
+ $X2=2.435 $Y2=1.375
r54 14 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.435 $Y=1.715
+ $X2=2.435 $Y2=1.88
r55 13 23 37.0826 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.435 $Y=1.21
+ $X2=2.435 $Y2=1.375
r56 9 11 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=2.4 $Y=0.495 $X2=2.4
+ $Y2=0.965
r57 5 15 438.415 $w=1.5e-07 $l=8.55e-07 $layer=POLY_cond $X=2.345 $Y=2.735
+ $X2=2.345 $Y2=1.88
r58 1 11 37.894 $w=2.05e-07 $l=1.02e-07 $layer=POLY_cond $X=2.372 $Y=1.067
+ $X2=2.372 $Y2=0.965
r59 1 13 46.2591 $w=2.05e-07 $l=1.43e-07 $layer=POLY_cond $X=2.372 $Y=1.067
+ $X2=2.372 $Y2=1.21
.ends

.subckt PM_SKY130_FD_SC_LP__O41AI_0%A1 3 7 10 12 15 17 18 19 20 25
c33 18 0 2.88954e-20 $X=3.12 $Y=1.295
c34 10 0 9.44548e-20 $X=3.032 $Y=1.658
r35 25 27 46.8028 $w=4.45e-07 $l=1.65e-07 $layer=POLY_cond $X=3.032 $Y=1.375
+ $X2=3.032 $Y2=1.21
r36 25 26 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3 $Y=1.375
+ $X2=3 $Y2=1.375
r37 19 20 11.8446 $w=3.58e-07 $l=3.7e-07 $layer=LI1_cond $X=3.095 $Y=1.665
+ $X2=3.095 $Y2=2.035
r38 19 26 9.28357 $w=3.58e-07 $l=2.9e-07 $layer=LI1_cond $X=3.095 $Y=1.665
+ $X2=3.095 $Y2=1.375
r39 18 26 2.56098 $w=3.58e-07 $l=8e-08 $layer=LI1_cond $X=3.095 $Y=1.295
+ $X2=3.095 $Y2=1.375
r40 13 15 92.2979 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=2.705 $Y=2.195
+ $X2=2.885 $Y2=2.195
r41 12 15 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.885 $Y=2.12
+ $X2=2.885 $Y2=2.195
r42 12 17 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=2.885 $Y=2.12
+ $X2=2.885 $Y2=1.88
r43 10 17 53.9265 $w=4.45e-07 $l=2.22e-07 $layer=POLY_cond $X=3.032 $Y=1.658
+ $X2=3.032 $Y2=1.88
r44 9 25 7.12377 $w=4.45e-07 $l=5.7e-08 $layer=POLY_cond $X=3.032 $Y=1.432
+ $X2=3.032 $Y2=1.375
r45 9 10 28.2451 $w=4.45e-07 $l=2.26e-07 $layer=POLY_cond $X=3.032 $Y=1.432
+ $X2=3.032 $Y2=1.658
r46 7 27 366.628 $w=1.5e-07 $l=7.15e-07 $layer=POLY_cond $X=2.885 $Y=0.495
+ $X2=2.885 $Y2=1.21
r47 1 13 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.705 $Y=2.27
+ $X2=2.705 $Y2=2.195
r48 1 3 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.705 $Y=2.27
+ $X2=2.705 $Y2=2.735
.ends

.subckt PM_SKY130_FD_SC_LP__O41AI_0%VPWR 1 2 9 13 15 16 17 18 20 34 36
r34 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r35 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r36 31 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r37 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r38 28 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r39 27 30 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r40 27 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r41 25 36 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=0.86 $Y=3.33
+ $X2=0.715 $Y2=3.33
r42 25 27 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=0.86 $Y=3.33 $X2=1.2
+ $Y2=3.33
r43 23 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r44 22 23 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r45 20 36 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=0.57 $Y=3.33
+ $X2=0.715 $Y2=3.33
r46 20 22 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=0.57 $Y=3.33
+ $X2=0.24 $Y2=3.33
r47 18 31 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r48 18 28 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r49 16 30 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=2.71 $Y=3.33 $X2=2.64
+ $Y2=3.33
r50 16 17 9.39981 $w=1.7e-07 $l=1.87e-07 $layer=LI1_cond $X=2.71 $Y=3.33
+ $X2=2.897 $Y2=3.33
r51 15 33 2.51176 $w=1.7e-07 $l=3.5e-08 $layer=LI1_cond $X=3.085 $Y=3.33
+ $X2=3.12 $Y2=3.33
r52 15 17 9.39981 $w=1.7e-07 $l=1.88e-07 $layer=LI1_cond $X=3.085 $Y=3.33
+ $X2=2.897 $Y2=3.33
r53 11 17 1.28102 $w=3.75e-07 $l=8.5e-08 $layer=LI1_cond $X=2.897 $Y=3.245
+ $X2=2.897 $Y2=3.33
r54 11 13 20.744 $w=3.73e-07 $l=6.75e-07 $layer=LI1_cond $X=2.897 $Y=3.245
+ $X2=2.897 $Y2=2.57
r55 7 36 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=0.715 $Y=3.245
+ $X2=0.715 $Y2=3.33
r56 7 9 26.8241 $w=2.88e-07 $l=6.75e-07 $layer=LI1_cond $X=0.715 $Y=3.245
+ $X2=0.715 $Y2=2.57
r57 2 13 300 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_PDIFF $count=2 $X=2.78
+ $Y=2.415 $X2=2.92 $Y2=2.57
r58 1 9 300 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_PDIFF $count=2 $X=0.61
+ $Y=2.415 $X2=0.735 $Y2=2.57
.ends

.subckt PM_SKY130_FD_SC_LP__O41AI_0%Y 1 2 7 11 13 14 15 16 17 18 26 27 36
c33 7 0 1.12009e-19 $X=1.03 $Y=2.14
r34 27 36 0.73171 $w=3.13e-07 $l=2e-08 $layer=LI1_cond $X=0.257 $Y=2.055
+ $X2=0.257 $Y2=2.035
r35 18 37 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=0.72 $Y=0.48
+ $X2=0.415 $Y2=0.48
r36 17 27 2.6726 $w=3.15e-07 $l=8.5e-08 $layer=LI1_cond $X=0.257 $Y=2.14
+ $X2=0.257 $Y2=2.055
r37 17 36 1.20732 $w=3.13e-07 $l=3.3e-08 $layer=LI1_cond $X=0.257 $Y=2.002
+ $X2=0.257 $Y2=2.035
r38 16 17 12.3293 $w=3.13e-07 $l=3.37e-07 $layer=LI1_cond $X=0.257 $Y=1.665
+ $X2=0.257 $Y2=2.002
r39 15 16 13.5366 $w=3.13e-07 $l=3.7e-07 $layer=LI1_cond $X=0.257 $Y=1.295
+ $X2=0.257 $Y2=1.665
r40 14 15 13.5366 $w=3.13e-07 $l=3.7e-07 $layer=LI1_cond $X=0.257 $Y=0.925
+ $X2=0.257 $Y2=1.295
r41 14 26 10.2439 $w=3.13e-07 $l=2.8e-07 $layer=LI1_cond $X=0.257 $Y=0.925
+ $X2=0.257 $Y2=0.645
r42 13 26 3.48456 $w=3.15e-07 $l=1.65e-07 $layer=LI1_cond $X=0.257 $Y=0.48
+ $X2=0.257 $Y2=0.645
r43 13 37 3.33673 $w=3.3e-07 $l=1.58e-07 $layer=LI1_cond $X=0.257 $Y=0.48
+ $X2=0.415 $Y2=0.48
r44 9 11 12.8689 $w=2.98e-07 $l=3.35e-07 $layer=LI1_cond $X=1.18 $Y=2.225
+ $X2=1.18 $Y2=2.56
r45 8 17 4.96789 $w=1.7e-07 $l=1.58e-07 $layer=LI1_cond $X=0.415 $Y=2.14
+ $X2=0.257 $Y2=2.14
r46 7 9 7.51767 $w=1.7e-07 $l=1.8775e-07 $layer=LI1_cond $X=1.03 $Y=2.14
+ $X2=1.18 $Y2=2.225
r47 7 8 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=1.03 $Y=2.14 $X2=0.415
+ $Y2=2.14
r48 2 11 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=1.025
+ $Y=2.415 $X2=1.165 $Y2=2.56
r49 1 13 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.205
+ $Y=0.285 $X2=0.33 $Y2=0.495
r50 1 18 182 $w=1.7e-07 $l=6.85602e-07 $layer=licon1_NDIFF $count=1 $X=0.205
+ $Y=0.285 $X2=0.8 $Y2=0.48
.ends

.subckt PM_SKY130_FD_SC_LP__O41AI_0%A_218_57# 1 2 3 12 14 15 18 20 24 26
c45 26 0 9.77123e-20 $X=2.175 $Y=0.915
c46 15 0 4.48098e-20 $X=1.37 $Y=0.915
r47 22 24 13.0871 $w=2.93e-07 $l=3.35e-07 $layer=LI1_cond $X=3.117 $Y=0.83
+ $X2=3.117 $Y2=0.495
r48 21 26 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=2.31 $Y=0.915
+ $X2=2.175 $Y2=0.915
r49 20 22 7.47753 $w=1.7e-07 $l=1.84673e-07 $layer=LI1_cond $X=2.97 $Y=0.915
+ $X2=3.117 $Y2=0.83
r50 20 21 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=2.97 $Y=0.915
+ $X2=2.31 $Y2=0.915
r51 16 26 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.175 $Y=0.83
+ $X2=2.175 $Y2=0.915
r52 16 18 14.2988 $w=2.68e-07 $l=3.35e-07 $layer=LI1_cond $X=2.175 $Y=0.83
+ $X2=2.175 $Y2=0.495
r53 14 26 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=2.04 $Y=0.915
+ $X2=2.175 $Y2=0.915
r54 14 15 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.04 $Y=0.915
+ $X2=1.37 $Y2=0.915
r55 10 15 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=1.235 $Y=0.83
+ $X2=1.37 $Y2=0.915
r56 10 12 14.2988 $w=2.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.235 $Y=0.83
+ $X2=1.235 $Y2=0.495
r57 3 24 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.96
+ $Y=0.285 $X2=3.1 $Y2=0.495
r58 2 18 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.045
+ $Y=0.285 $X2=2.185 $Y2=0.495
r59 1 12 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.09
+ $Y=0.285 $X2=1.23 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__O41AI_0%VGND 1 2 9 13 15 17 25 32 33 36 39
r37 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r38 33 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.64
+ $Y2=0
r39 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r40 30 39 8.42608 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=2.8 $Y=0 $X2=2.64
+ $Y2=0
r41 30 32 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=2.8 $Y=0 $X2=3.12
+ $Y2=0
r42 29 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r43 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r44 26 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.87 $Y=0 $X2=1.705
+ $Y2=0
r45 26 28 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=1.87 $Y=0 $X2=2.16
+ $Y2=0
r46 25 39 8.42608 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=2.48 $Y=0 $X2=2.64
+ $Y2=0
r47 25 28 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=2.48 $Y=0 $X2=2.16
+ $Y2=0
r48 23 24 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r49 20 24 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r50 19 23 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r51 19 20 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r52 17 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.54 $Y=0 $X2=1.705
+ $Y2=0
r53 17 23 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=1.54 $Y=0 $X2=1.2
+ $Y2=0
r54 15 29 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r55 15 24 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r56 15 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r57 11 39 0.800721 $w=3.2e-07 $l=8.5e-08 $layer=LI1_cond $X=2.64 $Y=0.085
+ $X2=2.64 $Y2=0
r58 11 13 14.7657 $w=3.18e-07 $l=4.1e-07 $layer=LI1_cond $X=2.64 $Y=0.085
+ $X2=2.64 $Y2=0.495
r59 7 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.705 $Y=0.085
+ $X2=1.705 $Y2=0
r60 7 9 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=1.705 $Y=0.085
+ $X2=1.705 $Y2=0.495
r61 2 13 182 $w=1.7e-07 $l=2.82489e-07 $layer=licon1_NDIFF $count=1 $X=2.475
+ $Y=0.285 $X2=2.645 $Y2=0.495
r62 1 9 182 $w=1.7e-07 $l=2.8801e-07 $layer=licon1_NDIFF $count=1 $X=1.52
+ $Y=0.285 $X2=1.705 $Y2=0.495
.ends

