* File: sky130_fd_sc_lp__busreceiver_1.pex.spice
* Created: Wed Sep  2 09:37:54 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__BUSRECEIVER_1%A_70_237# 1 2 9 12 14 17 18 21 22 23
+ 24 27 29 31 36
r56 31 33 2.88111 $w=3.18e-07 $l=8e-08 $layer=LI1_cond $X=1.185 $Y=0.855
+ $X2=1.185 $Y2=0.935
r57 25 27 7.38284 $w=3.18e-07 $l=2.05e-07 $layer=LI1_cond $X=1.185 $Y=1.775
+ $X2=1.185 $Y2=1.98
r58 23 25 7.68211 $w=1.7e-07 $l=1.9799e-07 $layer=LI1_cond $X=1.025 $Y=1.69
+ $X2=1.185 $Y2=1.775
r59 23 24 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=1.025 $Y=1.69
+ $X2=0.695 $Y2=1.69
r60 21 33 4.44149 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=1.025 $Y=0.935
+ $X2=1.185 $Y2=0.935
r61 21 22 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=1.025 $Y=0.935
+ $X2=0.695 $Y2=0.935
r62 19 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.61 $Y=1.02
+ $X2=0.695 $Y2=0.935
r63 19 29 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=0.61 $Y=1.02
+ $X2=0.61 $Y2=1.185
r64 18 37 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.515 $Y=1.35
+ $X2=0.515 $Y2=1.515
r65 18 36 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.515 $Y=1.35
+ $X2=0.515 $Y2=1.185
r66 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.515
+ $Y=1.35 $X2=0.515 $Y2=1.35
r67 15 24 12.7888 $w=1.23e-07 $l=1.70276e-07 $layer=LI1_cond $X=0.562 $Y=1.605
+ $X2=0.695 $Y2=1.69
r68 15 17 11.0895 $w=2.63e-07 $l=2.55e-07 $layer=LI1_cond $X=0.562 $Y=1.605
+ $X2=0.562 $Y2=1.35
r69 14 29 7.21712 $w=2.63e-07 $l=1.32e-07 $layer=LI1_cond $X=0.562 $Y=1.317
+ $X2=0.562 $Y2=1.185
r70 14 17 1.43512 $w=2.63e-07 $l=3.3e-08 $layer=LI1_cond $X=0.562 $Y=1.317
+ $X2=0.562 $Y2=1.35
r71 12 37 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=0.475 $Y=2.465
+ $X2=0.475 $Y2=1.515
r72 9 36 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.475 $Y=0.655
+ $X2=0.475 $Y2=1.185
r73 2 27 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=1.04
+ $Y=1.835 $X2=1.18 $Y2=1.98
r74 1 31 182 $w=1.7e-07 $l=2.60768e-07 $layer=licon1_NDIFF $count=1 $X=1.04
+ $Y=0.655 $X2=1.18 $Y2=0.855
.ends

.subckt PM_SKY130_FD_SC_LP__BUSRECEIVER_1%A 1 3 6 8 13
r28 10 13 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=0.965 $Y=1.35
+ $X2=1.17 $Y2=1.35
r29 8 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.17
+ $Y=1.35 $X2=1.17 $Y2=1.35
r30 4 10 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.965 $Y=1.515
+ $X2=0.965 $Y2=1.35
r31 4 6 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=0.965 $Y=1.515
+ $X2=0.965 $Y2=2.155
r32 1 10 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.965 $Y=1.185
+ $X2=0.965 $Y2=1.35
r33 1 3 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.965 $Y=1.185
+ $X2=0.965 $Y2=0.865
.ends

.subckt PM_SKY130_FD_SC_LP__BUSRECEIVER_1%X 1 2 9 10 11 12 13 23 31 41 45
r18 43 45 52.9195 $w=1.73e-07 $l=8.35e-07 $layer=LI1_cond $X=0.172 $Y=1.03
+ $X2=0.172 $Y2=1.865
r19 28 31 1.28049 $w=2.68e-07 $l=3e-08 $layer=LI1_cond $X=0.22 $Y=2 $X2=0.22
+ $Y2=2.03
r20 21 41 1.28049 $w=2.68e-07 $l=3e-08 $layer=LI1_cond $X=0.22 $Y=0.895 $X2=0.22
+ $Y2=0.925
r21 13 38 5.76222 $w=2.68e-07 $l=1.35e-07 $layer=LI1_cond $X=0.22 $Y=2.775
+ $X2=0.22 $Y2=2.91
r22 12 13 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.22 $Y=2.405
+ $X2=0.22 $Y2=2.775
r23 11 28 1.06708 $w=2.68e-07 $l=2.5e-08 $layer=LI1_cond $X=0.22 $Y=1.975
+ $X2=0.22 $Y2=2
r24 11 45 6.11934 $w=2.68e-07 $l=1.1e-07 $layer=LI1_cond $X=0.22 $Y=1.975
+ $X2=0.22 $Y2=1.865
r25 11 12 14.7257 $w=2.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.22 $Y=2.06
+ $X2=0.22 $Y2=2.405
r26 11 31 1.28049 $w=2.68e-07 $l=3e-08 $layer=LI1_cond $X=0.22 $Y=2.06 $X2=0.22
+ $Y2=2.03
r27 10 43 4.75348 $w=2.68e-07 $l=7.8e-08 $layer=LI1_cond $X=0.22 $Y=0.952
+ $X2=0.22 $Y2=1.03
r28 10 41 1.15244 $w=2.68e-07 $l=2.7e-08 $layer=LI1_cond $X=0.22 $Y=0.952
+ $X2=0.22 $Y2=0.925
r29 10 21 1.19513 $w=2.68e-07 $l=2.8e-08 $layer=LI1_cond $X=0.22 $Y=0.867
+ $X2=0.22 $Y2=0.895
r30 9 10 13.3171 $w=2.68e-07 $l=3.12e-07 $layer=LI1_cond $X=0.22 $Y=0.555
+ $X2=0.22 $Y2=0.867
r31 9 23 5.76222 $w=2.68e-07 $l=1.35e-07 $layer=LI1_cond $X=0.22 $Y=0.555
+ $X2=0.22 $Y2=0.42
r32 2 38 400 $w=1.7e-07 $l=1.13578e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.835 $X2=0.26 $Y2=2.91
r33 2 31 400 $w=1.7e-07 $l=2.498e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.835 $X2=0.26 $Y2=2.03
r34 1 23 91 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__BUSRECEIVER_1%VPWR 1 6 10 12 19 20 23
r20 19 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r21 17 23 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.855 $Y=3.33
+ $X2=0.69 $Y2=3.33
r22 17 19 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.855 $Y=3.33
+ $X2=1.2 $Y2=3.33
r23 14 15 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r24 12 23 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.525 $Y=3.33
+ $X2=0.69 $Y2=3.33
r25 12 14 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.525 $Y=3.33
+ $X2=0.24 $Y2=3.33
r26 10 20 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r27 10 15 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r28 10 23 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r29 6 9 15.3659 $w=3.28e-07 $l=4.4e-07 $layer=LI1_cond $X=0.69 $Y=2.055 $X2=0.69
+ $Y2=2.495
r30 4 23 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=3.245 $X2=0.69
+ $Y2=3.33
r31 4 9 26.1919 $w=3.28e-07 $l=7.5e-07 $layer=LI1_cond $X=0.69 $Y=3.245 $X2=0.69
+ $Y2=2.495
r32 1 9 300 $w=1.7e-07 $l=7.26636e-07 $layer=licon1_PDIFF $count=2 $X=0.55
+ $Y=1.835 $X2=0.69 $Y2=2.495
r33 1 6 600 $w=1.7e-07 $l=2.81425e-07 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=1.835 $X2=0.69 $Y2=2.055
.ends

.subckt PM_SKY130_FD_SC_LP__BUSRECEIVER_1%VGND 1 6 8 10 17 18 21
r24 17 18 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r25 15 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.855 $Y=0 $X2=0.69
+ $Y2=0
r26 15 17 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.855 $Y=0 $X2=1.2
+ $Y2=0
r27 12 13 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r28 10 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.525 $Y=0 $X2=0.69
+ $Y2=0
r29 10 12 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.525 $Y=0 $X2=0.24
+ $Y2=0
r30 8 18 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r31 8 13 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r32 8 21 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r33 4 21 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=0.085 $X2=0.69
+ $Y2=0
r34 4 6 16.4136 $w=3.28e-07 $l=4.7e-07 $layer=LI1_cond $X=0.69 $Y=0.085 $X2=0.69
+ $Y2=0.555
r35 1 6 182 $w=1.7e-07 $l=3.83667e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.235 $X2=0.69 $Y2=0.555
.ends

