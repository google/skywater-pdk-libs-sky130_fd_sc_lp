* File: sky130_fd_sc_lp__inv_m.pex.spice
* Created: Fri Aug 28 10:38:51 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__INV_M%A 3 7 9 10 11 12 18 19 22
r21 19 22 3.60455 $w=1.98e-07 $l=6.5e-08 $layer=LI1_cond $X=0.255 $Y=1.12
+ $X2=0.255 $Y2=1.055
r22 18 21 88.6355 $w=4.55e-07 $l=5.05e-07 $layer=POLY_cond $X=0.332 $Y=1.12
+ $X2=0.332 $Y2=1.625
r23 18 20 47.0767 $w=4.55e-07 $l=1.65e-07 $layer=POLY_cond $X=0.332 $Y=1.12
+ $X2=0.332 $Y2=0.955
r24 18 19 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.27
+ $Y=1.12 $X2=0.27 $Y2=1.12
r25 11 12 20.5182 $w=1.98e-07 $l=3.7e-07 $layer=LI1_cond $X=0.255 $Y=1.665
+ $X2=0.255 $Y2=2.035
r26 10 11 20.5182 $w=1.98e-07 $l=3.7e-07 $layer=LI1_cond $X=0.255 $Y=1.295
+ $X2=0.255 $Y2=1.665
r27 10 19 9.70455 $w=1.98e-07 $l=1.75e-07 $layer=LI1_cond $X=0.255 $Y=1.295
+ $X2=0.255 $Y2=1.12
r28 9 22 8.04083 $w=2e-07 $l=1.3e-07 $layer=LI1_cond $X=0.255 $Y=0.925 $X2=0.255
+ $Y2=1.055
r29 7 21 458.926 $w=1.5e-07 $l=8.95e-07 $layer=POLY_cond $X=0.485 $Y=2.52
+ $X2=0.485 $Y2=1.625
r30 3 20 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.485 $Y=0.56
+ $X2=0.485 $Y2=0.955
.ends

.subckt PM_SKY130_FD_SC_LP__INV_M%VPWR 1 4 6 8 12 13
r13 16 17 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r14 12 13 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r15 10 16 3.65184 $w=1.7e-07 $l=1.88e-07 $layer=LI1_cond $X=0.375 $Y=3.33
+ $X2=0.187 $Y2=3.33
r16 10 12 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.375 $Y=3.33
+ $X2=0.72 $Y2=3.33
r17 8 13 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=0.48 $Y=3.33
+ $X2=0.72 $Y2=3.33
r18 8 17 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=0.48 $Y=3.33
+ $X2=0.24 $Y2=3.33
r19 4 16 3.26335 $w=2.1e-07 $l=1.19499e-07 $layer=LI1_cond $X=0.27 $Y=3.245
+ $X2=0.187 $Y2=3.33
r20 4 6 38.026 $w=2.08e-07 $l=7.2e-07 $layer=LI1_cond $X=0.27 $Y=3.245 $X2=0.27
+ $Y2=2.525
r21 1 6 600 $w=1.7e-07 $l=2.7037e-07 $layer=licon1_PDIFF $count=1 $X=0.145
+ $Y=2.31 $X2=0.27 $Y2=2.525
.ends

.subckt PM_SKY130_FD_SC_LP__INV_M%Y 1 2 7 8 9 10 11 12 20
r10 12 33 13.7316 $w=2.08e-07 $l=2.6e-07 $layer=LI1_cond $X=0.7 $Y=2.775 $X2=0.7
+ $Y2=2.515
r11 11 33 5.80952 $w=2.08e-07 $l=1.1e-07 $layer=LI1_cond $X=0.7 $Y=2.405 $X2=0.7
+ $Y2=2.515
r12 10 11 19.5411 $w=2.08e-07 $l=3.7e-07 $layer=LI1_cond $X=0.7 $Y=2.035 $X2=0.7
+ $Y2=2.405
r13 9 10 19.5411 $w=2.08e-07 $l=3.7e-07 $layer=LI1_cond $X=0.7 $Y=1.665 $X2=0.7
+ $Y2=2.035
r14 8 9 19.5411 $w=2.08e-07 $l=3.7e-07 $layer=LI1_cond $X=0.7 $Y=1.295 $X2=0.7
+ $Y2=1.665
r15 7 8 19.5411 $w=2.08e-07 $l=3.7e-07 $layer=LI1_cond $X=0.7 $Y=0.925 $X2=0.7
+ $Y2=1.295
r16 7 20 16.6364 $w=2.08e-07 $l=3.15e-07 $layer=LI1_cond $X=0.7 $Y=0.925 $X2=0.7
+ $Y2=0.61
r17 2 33 600 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=1 $X=0.56
+ $Y=2.31 $X2=0.7 $Y2=2.515
r18 1 20 182 $w=1.7e-07 $l=3.2249e-07 $layer=licon1_NDIFF $count=1 $X=0.56
+ $Y=0.35 $X2=0.7 $Y2=0.61
.ends

.subckt PM_SKY130_FD_SC_LP__INV_M%VGND 1 4 6 8 12 13
r12 16 17 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r13 12 13 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r14 10 16 3.52085 $w=1.7e-07 $l=1.78e-07 $layer=LI1_cond $X=0.355 $Y=0 $X2=0.177
+ $Y2=0
r15 10 12 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.355 $Y=0 $X2=0.72
+ $Y2=0
r16 8 13 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=0.48 $Y=0 $X2=0.72
+ $Y2=0
r17 8 17 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=0.48 $Y=0 $X2=0.24
+ $Y2=0
r18 4 16 3.32305 $w=1.9e-07 $l=1.19499e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.177 $Y2=0
r19 4 6 23.933 $w=1.88e-07 $l=4.1e-07 $layer=LI1_cond $X=0.26 $Y=0.085 $X2=0.26
+ $Y2=0.495
r20 1 6 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.145
+ $Y=0.35 $X2=0.27 $Y2=0.495
.ends

