* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__o2bb2ai_m A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
X0 a_110_535# A2_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X1 VPWR A1_N a_110_535# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X2 Y B2 a_390_535# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X3 a_390_535# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X4 Y a_110_535# a_410_78# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 a_116_81# A2_N a_110_535# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 VGND A1_N a_116_81# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 a_410_78# B2 VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 VGND B1 a_410_78# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 VPWR a_110_535# Y VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
.ends
