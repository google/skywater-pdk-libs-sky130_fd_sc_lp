* File: sky130_fd_sc_lp__inv_16.pxi.spice
* Created: Wed Sep  2 09:55:38 2020
* 
x_PM_SKY130_FD_SC_LP__INV_16%A N_A_M1001_g N_A_c_147_n N_A_M1000_g N_A_M1002_g
+ N_A_c_148_n N_A_M1004_g N_A_M1003_g N_A_c_149_n N_A_M1006_g N_A_M1005_g
+ N_A_c_150_n N_A_M1007_g N_A_M1008_g N_A_c_151_n N_A_M1010_g N_A_M1009_g
+ N_A_c_152_n N_A_M1011_g N_A_M1012_g N_A_c_153_n N_A_M1013_g N_A_M1014_g
+ N_A_c_154_n N_A_M1015_g N_A_M1016_g N_A_c_155_n N_A_M1018_g N_A_M1017_g
+ N_A_c_156_n N_A_M1020_g N_A_M1019_g N_A_c_157_n N_A_M1022_g N_A_M1021_g
+ N_A_c_158_n N_A_M1025_g N_A_M1023_g N_A_c_159_n N_A_M1027_g N_A_M1024_g
+ N_A_c_160_n N_A_M1028_g N_A_M1026_g N_A_c_161_n N_A_M1030_g N_A_M1029_g
+ N_A_c_162_n N_A_M1031_g A N_A_c_139_n N_A_c_140_n N_A_c_141_n N_A_c_142_n
+ N_A_c_143_n N_A_c_144_n N_A_c_145_n N_A_c_146_n N_A_c_171_n
+ PM_SKY130_FD_SC_LP__INV_16%A
x_PM_SKY130_FD_SC_LP__INV_16%VPB N_VPB_M1000_s N_VPB_M1004_s N_VPB_M1007_s
+ N_VPB_M1011_s N_VPB_M1015_s N_VPB_M1020_s N_VPB_M1025_s N_VPB_M1028_s
+ N_VPB_M1031_s N_VPB_c_397_n N_VPB_c_398_n N_VPB_c_399_n N_VPB_c_400_n
+ N_VPB_c_401_n N_VPB_c_402_n N_VPB_c_403_n N_VPB_c_404_n N_VPB_c_405_n
+ N_VPB_c_406_n N_VPB_c_407_n N_VPB_c_408_n N_VPB_c_409_n N_VPB_c_410_n
+ N_VPB_c_411_n N_VPB_c_412_n N_VPB_c_413_n N_VPB_c_414_n N_VPB_c_415_n
+ N_VPB_c_416_n N_VPB_c_417_n N_VPB_c_418_n VPB N_VPB_c_419_n N_VPB_c_420_n
+ N_VPB_c_396_n N_VPB_c_422_n N_VPB_c_423_n N_VPB_c_424_n
+ PM_SKY130_FD_SC_LP__INV_16%VPB
x_PM_SKY130_FD_SC_LP__INV_16%Y N_Y_M1001_s N_Y_M1003_s N_Y_M1008_s N_Y_M1012_s
+ N_Y_M1016_s N_Y_M1019_s N_Y_M1023_s N_Y_M1026_s N_Y_M1000_d N_Y_M1006_d
+ N_Y_M1010_d N_Y_M1013_d N_Y_M1018_d N_Y_M1022_d N_Y_M1027_d N_Y_M1030_d Y
+ N_Y_c_548_n N_Y_c_549_n N_Y_c_550_n N_Y_c_551_n N_Y_c_552_n N_Y_c_553_n
+ N_Y_c_554_n N_Y_c_555_n N_Y_c_626_n PM_SKY130_FD_SC_LP__INV_16%Y
x_PM_SKY130_FD_SC_LP__INV_16%VGND N_VGND_M1001_d N_VGND_M1002_d N_VGND_M1005_d
+ N_VGND_M1009_d N_VGND_M1014_d N_VGND_M1017_d N_VGND_M1021_d N_VGND_M1024_d
+ N_VGND_M1029_d N_VGND_c_728_n N_VGND_c_729_n N_VGND_c_730_n N_VGND_c_731_n
+ N_VGND_c_732_n N_VGND_c_733_n N_VGND_c_734_n N_VGND_c_735_n N_VGND_c_736_n
+ N_VGND_c_737_n N_VGND_c_738_n N_VGND_c_739_n N_VGND_c_740_n N_VGND_c_741_n
+ N_VGND_c_742_n N_VGND_c_743_n N_VGND_c_744_n N_VGND_c_745_n N_VGND_c_746_n
+ N_VGND_c_747_n N_VGND_c_748_n N_VGND_c_749_n VGND N_VGND_c_750_n
+ N_VGND_c_751_n N_VGND_c_752_n N_VGND_c_753_n N_VGND_c_754_n N_VGND_c_755_n
+ PM_SKY130_FD_SC_LP__INV_16%VGND
cc_1 VNB N_A_M1001_g 0.034068f $X=-0.19 $Y=-0.245 $X2=0.55 $Y2=0.655
cc_2 VNB N_A_M1002_g 0.0237342f $X=-0.19 $Y=-0.245 $X2=0.98 $Y2=0.655
cc_3 VNB N_A_M1003_g 0.0237342f $X=-0.19 $Y=-0.245 $X2=1.41 $Y2=0.655
cc_4 VNB N_A_M1005_g 0.0237342f $X=-0.19 $Y=-0.245 $X2=1.84 $Y2=0.655
cc_5 VNB N_A_M1008_g 0.0237342f $X=-0.19 $Y=-0.245 $X2=2.27 $Y2=0.655
cc_6 VNB N_A_M1009_g 0.0237342f $X=-0.19 $Y=-0.245 $X2=2.7 $Y2=0.655
cc_7 VNB N_A_M1012_g 0.0237342f $X=-0.19 $Y=-0.245 $X2=3.13 $Y2=0.655
cc_8 VNB N_A_M1014_g 0.0237342f $X=-0.19 $Y=-0.245 $X2=3.56 $Y2=0.655
cc_9 VNB N_A_M1016_g 0.0237342f $X=-0.19 $Y=-0.245 $X2=3.99 $Y2=0.655
cc_10 VNB N_A_M1017_g 0.0237342f $X=-0.19 $Y=-0.245 $X2=4.42 $Y2=0.655
cc_11 VNB N_A_M1019_g 0.0237342f $X=-0.19 $Y=-0.245 $X2=4.85 $Y2=0.655
cc_12 VNB N_A_M1021_g 0.0237342f $X=-0.19 $Y=-0.245 $X2=5.28 $Y2=0.655
cc_13 VNB N_A_M1023_g 0.0237342f $X=-0.19 $Y=-0.245 $X2=5.71 $Y2=0.655
cc_14 VNB N_A_M1024_g 0.0237342f $X=-0.19 $Y=-0.245 $X2=6.14 $Y2=0.655
cc_15 VNB N_A_M1026_g 0.0237342f $X=-0.19 $Y=-0.245 $X2=6.57 $Y2=0.655
cc_16 VNB N_A_M1029_g 0.034068f $X=-0.19 $Y=-0.245 $X2=7 $Y2=0.655
cc_17 VNB N_A_c_139_n 0.00120838f $X=-0.19 $Y=-0.245 $X2=1.195 $Y2=1.5
cc_18 VNB N_A_c_140_n 0.00120838f $X=-0.19 $Y=-0.245 $X2=2.055 $Y2=1.5
cc_19 VNB N_A_c_141_n 0.00120838f $X=-0.19 $Y=-0.245 $X2=2.915 $Y2=1.5
cc_20 VNB N_A_c_142_n 0.00120838f $X=-0.19 $Y=-0.245 $X2=3.775 $Y2=1.5
cc_21 VNB N_A_c_143_n 0.00120838f $X=-0.19 $Y=-0.245 $X2=4.635 $Y2=1.5
cc_22 VNB N_A_c_144_n 0.00120838f $X=-0.19 $Y=-0.245 $X2=5.495 $Y2=1.5
cc_23 VNB N_A_c_145_n 0.00120838f $X=-0.19 $Y=-0.245 $X2=6.355 $Y2=1.5
cc_24 VNB N_A_c_146_n 0.302385f $X=-0.19 $Y=-0.245 $X2=7 $Y2=1.53
cc_25 VNB N_VPB_c_396_n 0.322901f $X=-0.19 $Y=-0.245 $X2=2.915 $Y2=1.5
cc_26 VNB N_Y_c_548_n 0.00531707f $X=-0.19 $Y=-0.245 $X2=3.56 $Y2=0.655
cc_27 VNB N_Y_c_549_n 0.00495171f $X=-0.19 $Y=-0.245 $X2=3.99 $Y2=2.465
cc_28 VNB N_Y_c_550_n 0.00495171f $X=-0.19 $Y=-0.245 $X2=4.85 $Y2=0.655
cc_29 VNB N_Y_c_551_n 0.00495171f $X=-0.19 $Y=-0.245 $X2=5.28 $Y2=1.725
cc_30 VNB N_Y_c_552_n 0.00495171f $X=-0.19 $Y=-0.245 $X2=6.14 $Y2=1.335
cc_31 VNB N_Y_c_553_n 0.00495171f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_Y_c_554_n 0.00495171f $X=-0.19 $Y=-0.245 $X2=7 $Y2=2.465
cc_33 VNB N_Y_c_555_n 0.00531707f $X=-0.19 $Y=-0.245 $X2=1.84 $Y2=1.53
cc_34 VNB N_VGND_c_728_n 0.013298f $X=-0.19 $Y=-0.245 $X2=1.84 $Y2=2.465
cc_35 VNB N_VGND_c_729_n 0.0355904f $X=-0.19 $Y=-0.245 $X2=2.27 $Y2=0.655
cc_36 VNB N_VGND_c_730_n 0.00400996f $X=-0.19 $Y=-0.245 $X2=2.27 $Y2=2.465
cc_37 VNB N_VGND_c_731_n 0.00400996f $X=-0.19 $Y=-0.245 $X2=2.7 $Y2=0.655
cc_38 VNB N_VGND_c_732_n 0.00400996f $X=-0.19 $Y=-0.245 $X2=2.7 $Y2=2.465
cc_39 VNB N_VGND_c_733_n 0.00400996f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_734_n 0.0168284f $X=-0.19 $Y=-0.245 $X2=3.13 $Y2=2.465
cc_41 VNB N_VGND_c_735_n 0.00400996f $X=-0.19 $Y=-0.245 $X2=3.56 $Y2=0.655
cc_42 VNB N_VGND_c_736_n 0.00400996f $X=-0.19 $Y=-0.245 $X2=3.56 $Y2=2.465
cc_43 VNB N_VGND_c_737_n 0.00400996f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_738_n 0.0355904f $X=-0.19 $Y=-0.245 $X2=4.42 $Y2=1.335
cc_45 VNB N_VGND_c_739_n 0.0168284f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_740_n 0.00500104f $X=-0.19 $Y=-0.245 $X2=4.42 $Y2=1.725
cc_47 VNB N_VGND_c_741_n 0.0168284f $X=-0.19 $Y=-0.245 $X2=4.42 $Y2=2.465
cc_48 VNB N_VGND_c_742_n 0.00500104f $X=-0.19 $Y=-0.245 $X2=4.85 $Y2=1.335
cc_49 VNB N_VGND_c_743_n 0.0168284f $X=-0.19 $Y=-0.245 $X2=4.85 $Y2=0.655
cc_50 VNB N_VGND_c_744_n 0.00500104f $X=-0.19 $Y=-0.245 $X2=4.85 $Y2=0.655
cc_51 VNB N_VGND_c_745_n 0.0168284f $X=-0.19 $Y=-0.245 $X2=4.85 $Y2=1.725
cc_52 VNB N_VGND_c_746_n 0.00500104f $X=-0.19 $Y=-0.245 $X2=4.85 $Y2=2.465
cc_53 VNB N_VGND_c_747_n 0.0116899f $X=-0.19 $Y=-0.245 $X2=4.85 $Y2=2.465
cc_54 VNB N_VGND_c_748_n 0.0168284f $X=-0.19 $Y=-0.245 $X2=5.28 $Y2=1.335
cc_55 VNB N_VGND_c_749_n 0.00567425f $X=-0.19 $Y=-0.245 $X2=5.28 $Y2=0.655
cc_56 VNB N_VGND_c_750_n 0.0168284f $X=-0.19 $Y=-0.245 $X2=5.28 $Y2=1.725
cc_57 VNB N_VGND_c_751_n 0.0168284f $X=-0.19 $Y=-0.245 $X2=6.14 $Y2=2.465
cc_58 VNB N_VGND_c_752_n 0.378599f $X=-0.19 $Y=-0.245 $X2=7 $Y2=2.465
cc_59 VNB N_VGND_c_753_n 0.00500104f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_754_n 0.00500104f $X=-0.19 $Y=-0.245 $X2=1.195 $Y2=1.5
cc_61 VNB N_VGND_c_755_n 0.00500104f $X=-0.19 $Y=-0.245 $X2=1.84 $Y2=1.53
cc_62 W_N38_331# N_A_c_147_n 0.0220458f $X=-0.19 $Y=1.655 $X2=0.55 $Y2=1.725
cc_63 W_N38_331# N_A_c_148_n 0.0159482f $X=-0.19 $Y=1.655 $X2=0.98 $Y2=1.725
cc_64 W_N38_331# N_A_c_149_n 0.0157473f $X=-0.19 $Y=1.655 $X2=1.41 $Y2=1.725
cc_65 W_N38_331# N_A_c_150_n 0.0157473f $X=-0.19 $Y=1.655 $X2=1.84 $Y2=1.725
cc_66 W_N38_331# N_A_c_151_n 0.0157473f $X=-0.19 $Y=1.655 $X2=2.27 $Y2=1.725
cc_67 W_N38_331# N_A_c_152_n 0.0157473f $X=-0.19 $Y=1.655 $X2=2.7 $Y2=1.725
cc_68 W_N38_331# N_A_c_153_n 0.0157473f $X=-0.19 $Y=1.655 $X2=3.13 $Y2=1.725
cc_69 W_N38_331# N_A_c_154_n 0.0157473f $X=-0.19 $Y=1.655 $X2=3.56 $Y2=1.725
cc_70 W_N38_331# N_A_c_155_n 0.0157473f $X=-0.19 $Y=1.655 $X2=3.99 $Y2=1.725
cc_71 W_N38_331# N_A_c_156_n 0.0157473f $X=-0.19 $Y=1.655 $X2=4.42 $Y2=1.725
cc_72 W_N38_331# N_A_c_157_n 0.0157473f $X=-0.19 $Y=1.655 $X2=4.85 $Y2=1.725
cc_73 W_N38_331# N_A_c_158_n 0.0157473f $X=-0.19 $Y=1.655 $X2=5.28 $Y2=1.725
cc_74 W_N38_331# N_A_c_159_n 0.0157473f $X=-0.19 $Y=1.655 $X2=5.71 $Y2=1.725
cc_75 W_N38_331# N_A_c_160_n 0.0157473f $X=-0.19 $Y=1.655 $X2=6.14 $Y2=1.725
cc_76 W_N38_331# N_A_c_161_n 0.0159482f $X=-0.19 $Y=1.655 $X2=6.57 $Y2=1.725
cc_77 W_N38_331# N_A_c_162_n 0.0220458f $X=-0.19 $Y=1.655 $X2=7 $Y2=1.725
cc_78 W_N38_331# N_A_c_139_n 0.00104594f $X=-0.19 $Y=1.655 $X2=1.195 $Y2=1.5
cc_79 W_N38_331# N_A_c_140_n 0.00104594f $X=-0.19 $Y=1.655 $X2=2.055 $Y2=1.5
cc_80 W_N38_331# N_A_c_141_n 0.00104594f $X=-0.19 $Y=1.655 $X2=2.915 $Y2=1.5
cc_81 W_N38_331# N_A_c_142_n 0.00104594f $X=-0.19 $Y=1.655 $X2=3.775 $Y2=1.5
cc_82 W_N38_331# N_A_c_143_n 0.00104594f $X=-0.19 $Y=1.655 $X2=4.635 $Y2=1.5
cc_83 W_N38_331# N_A_c_144_n 0.00104594f $X=-0.19 $Y=1.655 $X2=5.495 $Y2=1.5
cc_84 W_N38_331# N_A_c_145_n 0.00104594f $X=-0.19 $Y=1.655 $X2=6.355 $Y2=1.5
cc_85 W_N38_331# N_A_c_146_n 0.0996368f $X=-0.19 $Y=1.655 $X2=7 $Y2=1.53
cc_86 W_N38_331# N_A_c_171_n 0.00826739f $X=-0.19 $Y=1.655 $X2=6.355 $Y2=1.665
cc_87 W_N38_331# N_VPB_c_397_n 0.0132721f $X=-0.19 $Y=1.655 $X2=1.84 $Y2=2.465
cc_88 W_N38_331# N_VPB_c_398_n 0.0510625f $X=-0.19 $Y=1.655 $X2=2.27 $Y2=0.655
cc_89 W_N38_331# N_VPB_c_399_n 0.00400996f $X=-0.19 $Y=1.655 $X2=2.7 $Y2=1.335
cc_90 W_N38_331# N_VPB_c_400_n 0.00400996f $X=-0.19 $Y=1.655 $X2=2.7 $Y2=2.465
cc_91 W_N38_331# N_VPB_c_401_n 0.00400996f $X=-0.19 $Y=1.655 $X2=3.13 $Y2=2.465
cc_92 W_N38_331# N_VPB_c_402_n 0.00400996f $X=-0.19 $Y=1.655 $X2=3.56 $Y2=1.725
cc_93 W_N38_331# N_VPB_c_403_n 0.0167181f $X=-0.19 $Y=1.655 $X2=3.99 $Y2=0.655
cc_94 W_N38_331# N_VPB_c_404_n 0.00400996f $X=-0.19 $Y=1.655 $X2=3.99 $Y2=2.465
cc_95 W_N38_331# N_VPB_c_405_n 0.00400996f $X=-0.19 $Y=1.655 $X2=4.42 $Y2=1.725
cc_96 W_N38_331# N_VPB_c_406_n 0.00400996f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_97 W_N38_331# N_VPB_c_407_n 0.0493788f $X=-0.19 $Y=1.655 $X2=5.28 $Y2=0.655
cc_98 W_N38_331# N_VPB_c_408_n 0.0167181f $X=-0.19 $Y=1.655 $X2=5.71 $Y2=1.335
cc_99 W_N38_331# N_VPB_c_409_n 0.00497514f $X=-0.19 $Y=1.655 $X2=5.71 $Y2=0.655
cc_100 W_N38_331# N_VPB_c_410_n 0.0167181f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_101 W_N38_331# N_VPB_c_411_n 0.00497514f $X=-0.19 $Y=1.655 $X2=5.71 $Y2=1.725
cc_102 W_N38_331# N_VPB_c_412_n 0.0167181f $X=-0.19 $Y=1.655 $X2=5.71 $Y2=2.465
cc_103 W_N38_331# N_VPB_c_413_n 0.00497514f $X=-0.19 $Y=1.655 $X2=5.71 $Y2=2.465
cc_104 W_N38_331# N_VPB_c_414_n 0.0167181f $X=-0.19 $Y=1.655 $X2=6.14 $Y2=0.655
cc_105 W_N38_331# N_VPB_c_415_n 0.00497514f $X=-0.19 $Y=1.655 $X2=6.14 $Y2=0.655
cc_106 W_N38_331# N_VPB_c_416_n 0.0116899f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_107 W_N38_331# N_VPB_c_417_n 0.0167181f $X=-0.19 $Y=1.655 $X2=6.14 $Y2=1.725
cc_108 W_N38_331# N_VPB_c_418_n 0.00564836f $X=-0.19 $Y=1.655 $X2=6.14 $Y2=2.465
cc_109 W_N38_331# N_VPB_c_419_n 0.0167181f $X=-0.19 $Y=1.655 $X2=6.57 $Y2=0.655
cc_110 W_N38_331# N_VPB_c_420_n 0.0167181f $X=-0.19 $Y=1.655 $X2=0.55 $Y2=1.53
cc_111 W_N38_331# N_VPB_c_396_n 0.0556981f $X=-0.19 $Y=1.655 $X2=2.915 $Y2=1.5
cc_112 W_N38_331# N_VPB_c_422_n 0.00497514f $X=-0.19 $Y=1.655 $X2=3.775 $Y2=1.5
cc_113 W_N38_331# N_VPB_c_423_n 0.00497514f $X=-0.19 $Y=1.655 $X2=4.42 $Y2=1.53
cc_114 W_N38_331# N_VPB_c_424_n 0.00497514f $X=-0.19 $Y=1.655 $X2=4.635 $Y2=1.5
cc_115 W_N38_331# N_Y_c_548_n 0.0017675f $X=-0.19 $Y=1.655 $X2=3.56 $Y2=0.655
cc_116 W_N38_331# N_Y_c_549_n 0.00157031f $X=-0.19 $Y=1.655 $X2=3.99 $Y2=2.465
cc_117 W_N38_331# N_Y_c_550_n 0.00157031f $X=-0.19 $Y=1.655 $X2=4.85 $Y2=0.655
cc_118 W_N38_331# N_Y_c_551_n 0.00157031f $X=-0.19 $Y=1.655 $X2=5.28 $Y2=1.725
cc_119 W_N38_331# N_Y_c_552_n 0.00157031f $X=-0.19 $Y=1.655 $X2=6.14 $Y2=1.335
cc_120 W_N38_331# N_Y_c_553_n 0.00157031f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_121 W_N38_331# N_Y_c_554_n 0.00157031f $X=-0.19 $Y=1.655 $X2=7 $Y2=2.465
cc_122 W_N38_331# N_Y_c_555_n 0.0017675f $X=-0.19 $Y=1.655 $X2=1.84 $Y2=1.53
cc_123 N_A_c_147_n N_VPB_c_398_n 0.00413086f $X=0.55 $Y=1.725 $X2=0 $Y2=0
cc_124 N_A_c_148_n N_VPB_c_399_n 0.00211829f $X=0.98 $Y=1.725 $X2=0 $Y2=0
cc_125 N_A_c_149_n N_VPB_c_399_n 0.00211829f $X=1.41 $Y=1.725 $X2=0 $Y2=0
cc_126 N_A_c_139_n N_VPB_c_399_n 0.0171244f $X=1.195 $Y=1.5 $X2=0 $Y2=0
cc_127 N_A_c_146_n N_VPB_c_399_n 6.39733e-19 $X=7 $Y=1.53 $X2=0 $Y2=0
cc_128 N_A_c_171_n N_VPB_c_399_n 8.68506e-19 $X=6.355 $Y=1.665 $X2=0 $Y2=0
cc_129 N_A_c_150_n N_VPB_c_400_n 0.00211829f $X=1.84 $Y=1.725 $X2=0 $Y2=0
cc_130 N_A_c_151_n N_VPB_c_400_n 0.00211829f $X=2.27 $Y=1.725 $X2=0 $Y2=0
cc_131 N_A_c_140_n N_VPB_c_400_n 0.0171244f $X=2.055 $Y=1.5 $X2=0 $Y2=0
cc_132 N_A_c_146_n N_VPB_c_400_n 6.39733e-19 $X=7 $Y=1.53 $X2=0 $Y2=0
cc_133 N_A_c_171_n N_VPB_c_400_n 8.68506e-19 $X=6.355 $Y=1.665 $X2=0 $Y2=0
cc_134 N_A_c_152_n N_VPB_c_401_n 0.00211829f $X=2.7 $Y=1.725 $X2=0 $Y2=0
cc_135 N_A_c_153_n N_VPB_c_401_n 0.00211829f $X=3.13 $Y=1.725 $X2=0 $Y2=0
cc_136 N_A_c_141_n N_VPB_c_401_n 0.0171244f $X=2.915 $Y=1.5 $X2=0 $Y2=0
cc_137 N_A_c_146_n N_VPB_c_401_n 6.39733e-19 $X=7 $Y=1.53 $X2=0 $Y2=0
cc_138 N_A_c_171_n N_VPB_c_401_n 8.68506e-19 $X=6.355 $Y=1.665 $X2=0 $Y2=0
cc_139 N_A_c_154_n N_VPB_c_402_n 0.00211829f $X=3.56 $Y=1.725 $X2=0 $Y2=0
cc_140 N_A_c_155_n N_VPB_c_402_n 0.00211829f $X=3.99 $Y=1.725 $X2=0 $Y2=0
cc_141 N_A_c_142_n N_VPB_c_402_n 0.0171244f $X=3.775 $Y=1.5 $X2=0 $Y2=0
cc_142 N_A_c_146_n N_VPB_c_402_n 6.39733e-19 $X=7 $Y=1.53 $X2=0 $Y2=0
cc_143 N_A_c_171_n N_VPB_c_402_n 8.68506e-19 $X=6.355 $Y=1.665 $X2=0 $Y2=0
cc_144 N_A_c_155_n N_VPB_c_403_n 0.00585385f $X=3.99 $Y=1.725 $X2=0 $Y2=0
cc_145 N_A_c_156_n N_VPB_c_403_n 0.00585385f $X=4.42 $Y=1.725 $X2=0 $Y2=0
cc_146 N_A_c_156_n N_VPB_c_404_n 0.00211829f $X=4.42 $Y=1.725 $X2=0 $Y2=0
cc_147 N_A_c_157_n N_VPB_c_404_n 0.00211829f $X=4.85 $Y=1.725 $X2=0 $Y2=0
cc_148 N_A_c_143_n N_VPB_c_404_n 0.0171244f $X=4.635 $Y=1.5 $X2=0 $Y2=0
cc_149 N_A_c_146_n N_VPB_c_404_n 6.39733e-19 $X=7 $Y=1.53 $X2=0 $Y2=0
cc_150 N_A_c_171_n N_VPB_c_404_n 8.68506e-19 $X=6.355 $Y=1.665 $X2=0 $Y2=0
cc_151 N_A_c_158_n N_VPB_c_405_n 0.00211829f $X=5.28 $Y=1.725 $X2=0 $Y2=0
cc_152 N_A_c_159_n N_VPB_c_405_n 0.00211829f $X=5.71 $Y=1.725 $X2=0 $Y2=0
cc_153 N_A_c_144_n N_VPB_c_405_n 0.0171244f $X=5.495 $Y=1.5 $X2=0 $Y2=0
cc_154 N_A_c_146_n N_VPB_c_405_n 6.39733e-19 $X=7 $Y=1.53 $X2=0 $Y2=0
cc_155 N_A_c_171_n N_VPB_c_405_n 8.68506e-19 $X=6.355 $Y=1.665 $X2=0 $Y2=0
cc_156 N_A_c_160_n N_VPB_c_406_n 0.00211829f $X=6.14 $Y=1.725 $X2=0 $Y2=0
cc_157 N_A_c_161_n N_VPB_c_406_n 0.00211829f $X=6.57 $Y=1.725 $X2=0 $Y2=0
cc_158 N_A_c_145_n N_VPB_c_406_n 0.0171244f $X=6.355 $Y=1.5 $X2=0 $Y2=0
cc_159 N_A_c_146_n N_VPB_c_406_n 6.39733e-19 $X=7 $Y=1.53 $X2=0 $Y2=0
cc_160 N_A_c_171_n N_VPB_c_406_n 8.68506e-19 $X=6.355 $Y=1.665 $X2=0 $Y2=0
cc_161 N_A_c_162_n N_VPB_c_407_n 0.00413086f $X=7 $Y=1.725 $X2=0 $Y2=0
cc_162 N_A_c_149_n N_VPB_c_408_n 0.00585385f $X=1.41 $Y=1.725 $X2=0 $Y2=0
cc_163 N_A_c_150_n N_VPB_c_408_n 0.00585385f $X=1.84 $Y=1.725 $X2=0 $Y2=0
cc_164 N_A_c_151_n N_VPB_c_410_n 0.00585385f $X=2.27 $Y=1.725 $X2=0 $Y2=0
cc_165 N_A_c_152_n N_VPB_c_410_n 0.00585385f $X=2.7 $Y=1.725 $X2=0 $Y2=0
cc_166 N_A_c_153_n N_VPB_c_412_n 0.00585385f $X=3.13 $Y=1.725 $X2=0 $Y2=0
cc_167 N_A_c_154_n N_VPB_c_412_n 0.00585385f $X=3.56 $Y=1.725 $X2=0 $Y2=0
cc_168 N_A_c_159_n N_VPB_c_414_n 0.00585385f $X=5.71 $Y=1.725 $X2=0 $Y2=0
cc_169 N_A_c_160_n N_VPB_c_414_n 0.00585385f $X=6.14 $Y=1.725 $X2=0 $Y2=0
cc_170 N_A_c_161_n N_VPB_c_417_n 0.00585385f $X=6.57 $Y=1.725 $X2=0 $Y2=0
cc_171 N_A_c_162_n N_VPB_c_417_n 0.00585385f $X=7 $Y=1.725 $X2=0 $Y2=0
cc_172 N_A_c_147_n N_VPB_c_419_n 0.00585385f $X=0.55 $Y=1.725 $X2=0 $Y2=0
cc_173 N_A_c_148_n N_VPB_c_419_n 0.00585385f $X=0.98 $Y=1.725 $X2=0 $Y2=0
cc_174 N_A_c_157_n N_VPB_c_420_n 0.00585385f $X=4.85 $Y=1.725 $X2=0 $Y2=0
cc_175 N_A_c_158_n N_VPB_c_420_n 0.00585385f $X=5.28 $Y=1.725 $X2=0 $Y2=0
cc_176 N_A_c_147_n N_VPB_c_396_n 0.0116953f $X=0.55 $Y=1.725 $X2=0 $Y2=0
cc_177 N_A_c_148_n N_VPB_c_396_n 0.0104762f $X=0.98 $Y=1.725 $X2=0 $Y2=0
cc_178 N_A_c_149_n N_VPB_c_396_n 0.0106608f $X=1.41 $Y=1.725 $X2=0 $Y2=0
cc_179 N_A_c_150_n N_VPB_c_396_n 0.0106608f $X=1.84 $Y=1.725 $X2=0 $Y2=0
cc_180 N_A_c_151_n N_VPB_c_396_n 0.0106608f $X=2.27 $Y=1.725 $X2=0 $Y2=0
cc_181 N_A_c_152_n N_VPB_c_396_n 0.0106608f $X=2.7 $Y=1.725 $X2=0 $Y2=0
cc_182 N_A_c_153_n N_VPB_c_396_n 0.0106608f $X=3.13 $Y=1.725 $X2=0 $Y2=0
cc_183 N_A_c_154_n N_VPB_c_396_n 0.0106608f $X=3.56 $Y=1.725 $X2=0 $Y2=0
cc_184 N_A_c_155_n N_VPB_c_396_n 0.0106608f $X=3.99 $Y=1.725 $X2=0 $Y2=0
cc_185 N_A_c_156_n N_VPB_c_396_n 0.0106608f $X=4.42 $Y=1.725 $X2=0 $Y2=0
cc_186 N_A_c_157_n N_VPB_c_396_n 0.0106608f $X=4.85 $Y=1.725 $X2=0 $Y2=0
cc_187 N_A_c_158_n N_VPB_c_396_n 0.0106608f $X=5.28 $Y=1.725 $X2=0 $Y2=0
cc_188 N_A_c_159_n N_VPB_c_396_n 0.0106608f $X=5.71 $Y=1.725 $X2=0 $Y2=0
cc_189 N_A_c_160_n N_VPB_c_396_n 0.0106608f $X=6.14 $Y=1.725 $X2=0 $Y2=0
cc_190 N_A_c_161_n N_VPB_c_396_n 0.0104762f $X=6.57 $Y=1.725 $X2=0 $Y2=0
cc_191 N_A_c_162_n N_VPB_c_396_n 0.0117795f $X=7 $Y=1.725 $X2=0 $Y2=0
cc_192 N_A_M1001_g N_Y_c_548_n 0.00728339f $X=0.55 $Y=0.655 $X2=0 $Y2=0
cc_193 N_A_c_147_n N_Y_c_548_n 0.00365908f $X=0.55 $Y=1.725 $X2=0 $Y2=0
cc_194 N_A_M1002_g N_Y_c_548_n 0.00391701f $X=0.98 $Y=0.655 $X2=0 $Y2=0
cc_195 N_A_c_148_n N_Y_c_548_n 0.00208211f $X=0.98 $Y=1.725 $X2=0 $Y2=0
cc_196 N_A_c_139_n N_Y_c_548_n 0.0280537f $X=1.195 $Y=1.5 $X2=0 $Y2=0
cc_197 N_A_c_146_n N_Y_c_548_n 0.0355455f $X=7 $Y=1.53 $X2=0 $Y2=0
cc_198 N_A_c_171_n N_Y_c_548_n 0.00697809f $X=6.355 $Y=1.665 $X2=0 $Y2=0
cc_199 N_A_M1003_g N_Y_c_549_n 0.00391701f $X=1.41 $Y=0.655 $X2=0 $Y2=0
cc_200 N_A_c_149_n N_Y_c_549_n 0.00199205f $X=1.41 $Y=1.725 $X2=0 $Y2=0
cc_201 N_A_M1005_g N_Y_c_549_n 0.00391701f $X=1.84 $Y=0.655 $X2=0 $Y2=0
cc_202 N_A_c_150_n N_Y_c_549_n 0.00199205f $X=1.84 $Y=1.725 $X2=0 $Y2=0
cc_203 N_A_c_139_n N_Y_c_549_n 0.0287397f $X=1.195 $Y=1.5 $X2=0 $Y2=0
cc_204 N_A_c_140_n N_Y_c_549_n 0.0287397f $X=2.055 $Y=1.5 $X2=0 $Y2=0
cc_205 N_A_c_146_n N_Y_c_549_n 0.0230554f $X=7 $Y=1.53 $X2=0 $Y2=0
cc_206 N_A_c_171_n N_Y_c_549_n 0.0295778f $X=6.355 $Y=1.665 $X2=0 $Y2=0
cc_207 N_A_M1008_g N_Y_c_550_n 0.00391701f $X=2.27 $Y=0.655 $X2=0 $Y2=0
cc_208 N_A_c_151_n N_Y_c_550_n 0.00199205f $X=2.27 $Y=1.725 $X2=0 $Y2=0
cc_209 N_A_M1009_g N_Y_c_550_n 0.00391701f $X=2.7 $Y=0.655 $X2=0 $Y2=0
cc_210 N_A_c_152_n N_Y_c_550_n 0.00199205f $X=2.7 $Y=1.725 $X2=0 $Y2=0
cc_211 N_A_c_140_n N_Y_c_550_n 0.0287397f $X=2.055 $Y=1.5 $X2=0 $Y2=0
cc_212 N_A_c_141_n N_Y_c_550_n 0.0287397f $X=2.915 $Y=1.5 $X2=0 $Y2=0
cc_213 N_A_c_146_n N_Y_c_550_n 0.0230554f $X=7 $Y=1.53 $X2=0 $Y2=0
cc_214 N_A_c_171_n N_Y_c_550_n 0.0296325f $X=6.355 $Y=1.665 $X2=0 $Y2=0
cc_215 N_A_M1012_g N_Y_c_551_n 0.00391701f $X=3.13 $Y=0.655 $X2=0 $Y2=0
cc_216 N_A_c_153_n N_Y_c_551_n 0.00199205f $X=3.13 $Y=1.725 $X2=0 $Y2=0
cc_217 N_A_M1014_g N_Y_c_551_n 0.00391701f $X=3.56 $Y=0.655 $X2=0 $Y2=0
cc_218 N_A_c_154_n N_Y_c_551_n 0.00199205f $X=3.56 $Y=1.725 $X2=0 $Y2=0
cc_219 N_A_c_141_n N_Y_c_551_n 0.0287397f $X=2.915 $Y=1.5 $X2=0 $Y2=0
cc_220 N_A_c_142_n N_Y_c_551_n 0.0287397f $X=3.775 $Y=1.5 $X2=0 $Y2=0
cc_221 N_A_c_146_n N_Y_c_551_n 0.0230554f $X=7 $Y=1.53 $X2=0 $Y2=0
cc_222 N_A_c_171_n N_Y_c_551_n 0.0296325f $X=6.355 $Y=1.665 $X2=0 $Y2=0
cc_223 N_A_M1016_g N_Y_c_552_n 0.00391701f $X=3.99 $Y=0.655 $X2=0 $Y2=0
cc_224 N_A_c_155_n N_Y_c_552_n 0.00199205f $X=3.99 $Y=1.725 $X2=0 $Y2=0
cc_225 N_A_M1017_g N_Y_c_552_n 0.00391701f $X=4.42 $Y=0.655 $X2=0 $Y2=0
cc_226 N_A_c_156_n N_Y_c_552_n 0.00199205f $X=4.42 $Y=1.725 $X2=0 $Y2=0
cc_227 N_A_c_142_n N_Y_c_552_n 0.0287397f $X=3.775 $Y=1.5 $X2=0 $Y2=0
cc_228 N_A_c_143_n N_Y_c_552_n 0.0287397f $X=4.635 $Y=1.5 $X2=0 $Y2=0
cc_229 N_A_c_146_n N_Y_c_552_n 0.0230554f $X=7 $Y=1.53 $X2=0 $Y2=0
cc_230 N_A_c_171_n N_Y_c_552_n 0.0296325f $X=6.355 $Y=1.665 $X2=0 $Y2=0
cc_231 N_A_M1019_g N_Y_c_553_n 0.00391701f $X=4.85 $Y=0.655 $X2=0 $Y2=0
cc_232 N_A_c_157_n N_Y_c_553_n 0.00199205f $X=4.85 $Y=1.725 $X2=0 $Y2=0
cc_233 N_A_M1021_g N_Y_c_553_n 0.00391701f $X=5.28 $Y=0.655 $X2=0 $Y2=0
cc_234 N_A_c_158_n N_Y_c_553_n 0.00199205f $X=5.28 $Y=1.725 $X2=0 $Y2=0
cc_235 N_A_c_143_n N_Y_c_553_n 0.0287397f $X=4.635 $Y=1.5 $X2=0 $Y2=0
cc_236 N_A_c_144_n N_Y_c_553_n 0.0287397f $X=5.495 $Y=1.5 $X2=0 $Y2=0
cc_237 N_A_c_146_n N_Y_c_553_n 0.0230554f $X=7 $Y=1.53 $X2=0 $Y2=0
cc_238 N_A_c_171_n N_Y_c_553_n 0.0296325f $X=6.355 $Y=1.665 $X2=0 $Y2=0
cc_239 N_A_M1023_g N_Y_c_554_n 0.00391701f $X=5.71 $Y=0.655 $X2=0 $Y2=0
cc_240 N_A_c_159_n N_Y_c_554_n 0.00199205f $X=5.71 $Y=1.725 $X2=0 $Y2=0
cc_241 N_A_M1024_g N_Y_c_554_n 0.00391701f $X=6.14 $Y=0.655 $X2=0 $Y2=0
cc_242 N_A_c_160_n N_Y_c_554_n 0.00199205f $X=6.14 $Y=1.725 $X2=0 $Y2=0
cc_243 N_A_c_144_n N_Y_c_554_n 0.0287397f $X=5.495 $Y=1.5 $X2=0 $Y2=0
cc_244 N_A_c_145_n N_Y_c_554_n 0.0287397f $X=6.355 $Y=1.5 $X2=0 $Y2=0
cc_245 N_A_c_146_n N_Y_c_554_n 0.0230554f $X=7 $Y=1.53 $X2=0 $Y2=0
cc_246 N_A_c_171_n N_Y_c_554_n 0.0295778f $X=6.355 $Y=1.665 $X2=0 $Y2=0
cc_247 N_A_M1026_g N_Y_c_555_n 0.00391701f $X=6.57 $Y=0.655 $X2=0 $Y2=0
cc_248 N_A_c_161_n N_Y_c_555_n 0.00208211f $X=6.57 $Y=1.725 $X2=0 $Y2=0
cc_249 N_A_M1029_g N_Y_c_555_n 0.00728339f $X=7 $Y=0.655 $X2=0 $Y2=0
cc_250 N_A_c_162_n N_Y_c_555_n 0.00365908f $X=7 $Y=1.725 $X2=0 $Y2=0
cc_251 N_A_c_145_n N_Y_c_555_n 0.0280537f $X=6.355 $Y=1.5 $X2=0 $Y2=0
cc_252 N_A_c_146_n N_Y_c_555_n 0.0355455f $X=7 $Y=1.53 $X2=0 $Y2=0
cc_253 N_A_c_171_n N_Y_c_555_n 0.00697809f $X=6.355 $Y=1.665 $X2=0 $Y2=0
cc_254 N_A_c_147_n N_Y_c_626_n 0.00197372f $X=0.55 $Y=1.725 $X2=0 $Y2=0
cc_255 N_A_c_148_n N_Y_c_626_n 0.0123908f $X=0.98 $Y=1.725 $X2=0 $Y2=0
cc_256 N_A_c_149_n N_Y_c_626_n 0.00766908f $X=1.41 $Y=1.725 $X2=0 $Y2=0
cc_257 N_A_c_150_n N_Y_c_626_n 0.00766908f $X=1.84 $Y=1.725 $X2=0 $Y2=0
cc_258 N_A_c_151_n N_Y_c_626_n 0.00766908f $X=2.27 $Y=1.725 $X2=0 $Y2=0
cc_259 N_A_c_152_n N_Y_c_626_n 0.00766908f $X=2.7 $Y=1.725 $X2=0 $Y2=0
cc_260 N_A_c_153_n N_Y_c_626_n 0.00766908f $X=3.13 $Y=1.725 $X2=0 $Y2=0
cc_261 N_A_c_154_n N_Y_c_626_n 0.00766908f $X=3.56 $Y=1.725 $X2=0 $Y2=0
cc_262 N_A_c_155_n N_Y_c_626_n 0.00766908f $X=3.99 $Y=1.725 $X2=0 $Y2=0
cc_263 N_A_c_156_n N_Y_c_626_n 0.00766908f $X=4.42 $Y=1.725 $X2=0 $Y2=0
cc_264 N_A_c_157_n N_Y_c_626_n 0.00766908f $X=4.85 $Y=1.725 $X2=0 $Y2=0
cc_265 N_A_c_158_n N_Y_c_626_n 0.00766908f $X=5.28 $Y=1.725 $X2=0 $Y2=0
cc_266 N_A_c_159_n N_Y_c_626_n 0.00766908f $X=5.71 $Y=1.725 $X2=0 $Y2=0
cc_267 N_A_c_160_n N_Y_c_626_n 0.00766908f $X=6.14 $Y=1.725 $X2=0 $Y2=0
cc_268 N_A_c_161_n N_Y_c_626_n 0.0123908f $X=6.57 $Y=1.725 $X2=0 $Y2=0
cc_269 N_A_c_162_n N_Y_c_626_n 0.00197372f $X=7 $Y=1.725 $X2=0 $Y2=0
cc_270 N_A_c_139_n N_Y_c_626_n 2.76232e-19 $X=1.195 $Y=1.5 $X2=0 $Y2=0
cc_271 N_A_c_140_n N_Y_c_626_n 2.76232e-19 $X=2.055 $Y=1.5 $X2=0 $Y2=0
cc_272 N_A_c_141_n N_Y_c_626_n 2.76232e-19 $X=2.915 $Y=1.5 $X2=0 $Y2=0
cc_273 N_A_c_142_n N_Y_c_626_n 2.76232e-19 $X=3.775 $Y=1.5 $X2=0 $Y2=0
cc_274 N_A_c_143_n N_Y_c_626_n 2.76232e-19 $X=4.635 $Y=1.5 $X2=0 $Y2=0
cc_275 N_A_c_144_n N_Y_c_626_n 2.76232e-19 $X=5.495 $Y=1.5 $X2=0 $Y2=0
cc_276 N_A_c_145_n N_Y_c_626_n 2.76232e-19 $X=6.355 $Y=1.5 $X2=0 $Y2=0
cc_277 N_A_c_171_n N_Y_c_626_n 0.5279f $X=6.355 $Y=1.665 $X2=0 $Y2=0
cc_278 N_A_M1001_g N_VGND_c_729_n 0.00422005f $X=0.55 $Y=0.655 $X2=0 $Y2=0
cc_279 N_A_M1002_g N_VGND_c_730_n 0.00181392f $X=0.98 $Y=0.655 $X2=0 $Y2=0
cc_280 N_A_M1003_g N_VGND_c_730_n 0.00181392f $X=1.41 $Y=0.655 $X2=0 $Y2=0
cc_281 N_A_c_139_n N_VGND_c_730_n 0.00944516f $X=1.195 $Y=1.5 $X2=0 $Y2=0
cc_282 N_A_c_146_n N_VGND_c_730_n 7.26853e-19 $X=7 $Y=1.53 $X2=0 $Y2=0
cc_283 N_A_c_171_n N_VGND_c_730_n 0.00147804f $X=6.355 $Y=1.665 $X2=0 $Y2=0
cc_284 N_A_M1005_g N_VGND_c_731_n 0.00181392f $X=1.84 $Y=0.655 $X2=0 $Y2=0
cc_285 N_A_M1008_g N_VGND_c_731_n 0.00181392f $X=2.27 $Y=0.655 $X2=0 $Y2=0
cc_286 N_A_c_140_n N_VGND_c_731_n 0.00944516f $X=2.055 $Y=1.5 $X2=0 $Y2=0
cc_287 N_A_c_146_n N_VGND_c_731_n 7.26853e-19 $X=7 $Y=1.53 $X2=0 $Y2=0
cc_288 N_A_c_171_n N_VGND_c_731_n 0.00147804f $X=6.355 $Y=1.665 $X2=0 $Y2=0
cc_289 N_A_M1009_g N_VGND_c_732_n 0.00181392f $X=2.7 $Y=0.655 $X2=0 $Y2=0
cc_290 N_A_M1012_g N_VGND_c_732_n 0.00181392f $X=3.13 $Y=0.655 $X2=0 $Y2=0
cc_291 N_A_c_141_n N_VGND_c_732_n 0.00944516f $X=2.915 $Y=1.5 $X2=0 $Y2=0
cc_292 N_A_c_146_n N_VGND_c_732_n 7.26853e-19 $X=7 $Y=1.53 $X2=0 $Y2=0
cc_293 N_A_c_171_n N_VGND_c_732_n 0.00147804f $X=6.355 $Y=1.665 $X2=0 $Y2=0
cc_294 N_A_M1014_g N_VGND_c_733_n 0.00181392f $X=3.56 $Y=0.655 $X2=0 $Y2=0
cc_295 N_A_M1016_g N_VGND_c_733_n 0.00181392f $X=3.99 $Y=0.655 $X2=0 $Y2=0
cc_296 N_A_c_142_n N_VGND_c_733_n 0.00944516f $X=3.775 $Y=1.5 $X2=0 $Y2=0
cc_297 N_A_c_146_n N_VGND_c_733_n 7.26853e-19 $X=7 $Y=1.53 $X2=0 $Y2=0
cc_298 N_A_c_171_n N_VGND_c_733_n 0.00147804f $X=6.355 $Y=1.665 $X2=0 $Y2=0
cc_299 N_A_M1016_g N_VGND_c_734_n 0.00585385f $X=3.99 $Y=0.655 $X2=0 $Y2=0
cc_300 N_A_M1017_g N_VGND_c_734_n 0.00585385f $X=4.42 $Y=0.655 $X2=0 $Y2=0
cc_301 N_A_M1017_g N_VGND_c_735_n 0.00181392f $X=4.42 $Y=0.655 $X2=0 $Y2=0
cc_302 N_A_M1019_g N_VGND_c_735_n 0.00181392f $X=4.85 $Y=0.655 $X2=0 $Y2=0
cc_303 N_A_c_143_n N_VGND_c_735_n 0.00944516f $X=4.635 $Y=1.5 $X2=0 $Y2=0
cc_304 N_A_c_146_n N_VGND_c_735_n 7.26853e-19 $X=7 $Y=1.53 $X2=0 $Y2=0
cc_305 N_A_c_171_n N_VGND_c_735_n 0.00147804f $X=6.355 $Y=1.665 $X2=0 $Y2=0
cc_306 N_A_M1021_g N_VGND_c_736_n 0.00181392f $X=5.28 $Y=0.655 $X2=0 $Y2=0
cc_307 N_A_M1023_g N_VGND_c_736_n 0.00181392f $X=5.71 $Y=0.655 $X2=0 $Y2=0
cc_308 N_A_c_144_n N_VGND_c_736_n 0.00944516f $X=5.495 $Y=1.5 $X2=0 $Y2=0
cc_309 N_A_c_146_n N_VGND_c_736_n 7.26853e-19 $X=7 $Y=1.53 $X2=0 $Y2=0
cc_310 N_A_c_171_n N_VGND_c_736_n 0.00147804f $X=6.355 $Y=1.665 $X2=0 $Y2=0
cc_311 N_A_M1024_g N_VGND_c_737_n 0.00181392f $X=6.14 $Y=0.655 $X2=0 $Y2=0
cc_312 N_A_M1026_g N_VGND_c_737_n 0.00181392f $X=6.57 $Y=0.655 $X2=0 $Y2=0
cc_313 N_A_c_145_n N_VGND_c_737_n 0.00944516f $X=6.355 $Y=1.5 $X2=0 $Y2=0
cc_314 N_A_c_146_n N_VGND_c_737_n 7.26853e-19 $X=7 $Y=1.53 $X2=0 $Y2=0
cc_315 N_A_c_171_n N_VGND_c_737_n 0.00147804f $X=6.355 $Y=1.665 $X2=0 $Y2=0
cc_316 N_A_M1029_g N_VGND_c_738_n 0.00422005f $X=7 $Y=0.655 $X2=0 $Y2=0
cc_317 N_A_M1003_g N_VGND_c_739_n 0.00585385f $X=1.41 $Y=0.655 $X2=0 $Y2=0
cc_318 N_A_M1005_g N_VGND_c_739_n 0.00585385f $X=1.84 $Y=0.655 $X2=0 $Y2=0
cc_319 N_A_M1008_g N_VGND_c_741_n 0.00585385f $X=2.27 $Y=0.655 $X2=0 $Y2=0
cc_320 N_A_M1009_g N_VGND_c_741_n 0.00585385f $X=2.7 $Y=0.655 $X2=0 $Y2=0
cc_321 N_A_M1012_g N_VGND_c_743_n 0.00585385f $X=3.13 $Y=0.655 $X2=0 $Y2=0
cc_322 N_A_M1014_g N_VGND_c_743_n 0.00585385f $X=3.56 $Y=0.655 $X2=0 $Y2=0
cc_323 N_A_M1023_g N_VGND_c_745_n 0.00585385f $X=5.71 $Y=0.655 $X2=0 $Y2=0
cc_324 N_A_M1024_g N_VGND_c_745_n 0.00585385f $X=6.14 $Y=0.655 $X2=0 $Y2=0
cc_325 N_A_M1026_g N_VGND_c_748_n 0.00585385f $X=6.57 $Y=0.655 $X2=0 $Y2=0
cc_326 N_A_M1029_g N_VGND_c_748_n 0.00585385f $X=7 $Y=0.655 $X2=0 $Y2=0
cc_327 N_A_M1001_g N_VGND_c_750_n 0.00585385f $X=0.55 $Y=0.655 $X2=0 $Y2=0
cc_328 N_A_M1002_g N_VGND_c_750_n 0.00585385f $X=0.98 $Y=0.655 $X2=0 $Y2=0
cc_329 N_A_M1019_g N_VGND_c_751_n 0.00585385f $X=4.85 $Y=0.655 $X2=0 $Y2=0
cc_330 N_A_M1021_g N_VGND_c_751_n 0.00585385f $X=5.28 $Y=0.655 $X2=0 $Y2=0
cc_331 N_A_M1001_g N_VGND_c_752_n 0.0118104f $X=0.55 $Y=0.655 $X2=0 $Y2=0
cc_332 N_A_M1002_g N_VGND_c_752_n 0.0107375f $X=0.98 $Y=0.655 $X2=0 $Y2=0
cc_333 N_A_M1003_g N_VGND_c_752_n 0.0107375f $X=1.41 $Y=0.655 $X2=0 $Y2=0
cc_334 N_A_M1005_g N_VGND_c_752_n 0.0107375f $X=1.84 $Y=0.655 $X2=0 $Y2=0
cc_335 N_A_M1008_g N_VGND_c_752_n 0.0107375f $X=2.27 $Y=0.655 $X2=0 $Y2=0
cc_336 N_A_M1009_g N_VGND_c_752_n 0.0107375f $X=2.7 $Y=0.655 $X2=0 $Y2=0
cc_337 N_A_M1012_g N_VGND_c_752_n 0.0107375f $X=3.13 $Y=0.655 $X2=0 $Y2=0
cc_338 N_A_M1014_g N_VGND_c_752_n 0.0107375f $X=3.56 $Y=0.655 $X2=0 $Y2=0
cc_339 N_A_M1016_g N_VGND_c_752_n 0.0107375f $X=3.99 $Y=0.655 $X2=0 $Y2=0
cc_340 N_A_M1017_g N_VGND_c_752_n 0.0107375f $X=4.42 $Y=0.655 $X2=0 $Y2=0
cc_341 N_A_M1019_g N_VGND_c_752_n 0.0107375f $X=4.85 $Y=0.655 $X2=0 $Y2=0
cc_342 N_A_M1021_g N_VGND_c_752_n 0.0107375f $X=5.28 $Y=0.655 $X2=0 $Y2=0
cc_343 N_A_M1023_g N_VGND_c_752_n 0.0107375f $X=5.71 $Y=0.655 $X2=0 $Y2=0
cc_344 N_A_M1024_g N_VGND_c_752_n 0.0107375f $X=6.14 $Y=0.655 $X2=0 $Y2=0
cc_345 N_A_M1026_g N_VGND_c_752_n 0.0107375f $X=6.57 $Y=0.655 $X2=0 $Y2=0
cc_346 N_A_M1029_g N_VGND_c_752_n 0.0118977f $X=7 $Y=0.655 $X2=0 $Y2=0
cc_347 N_VPB_c_396_n N_Y_M1000_d 0.00302605f $X=7.44 $Y=3.33 $X2=0 $Y2=0
cc_348 N_VPB_c_396_n N_Y_M1006_d 0.00302605f $X=7.44 $Y=3.33 $X2=0 $Y2=0
cc_349 N_VPB_c_396_n N_Y_M1010_d 0.00302605f $X=7.44 $Y=3.33 $X2=0 $Y2=0
cc_350 N_VPB_c_396_n N_Y_M1013_d 0.00302605f $X=7.44 $Y=3.33 $X2=0 $Y2=0
cc_351 N_VPB_c_396_n N_Y_M1018_d 0.00302605f $X=7.44 $Y=3.33 $X2=0 $Y2=0
cc_352 N_VPB_c_396_n N_Y_M1022_d 0.00302605f $X=7.44 $Y=3.33 $X2=0 $Y2=0
cc_353 N_VPB_c_396_n N_Y_M1027_d 0.00302605f $X=7.44 $Y=3.33 $X2=0 $Y2=0
cc_354 N_VPB_c_396_n N_Y_M1030_d 0.00302605f $X=7.44 $Y=3.33 $X2=0 $Y2=0
cc_355 N_VPB_c_399_n N_Y_c_548_n 0.00822181f $X=1.195 $Y=2.085 $X2=0 $Y2=0
cc_356 N_VPB_c_419_n N_Y_c_548_n 0.0128989f $X=1.065 $Y=3.33 $X2=0 $Y2=0
cc_357 N_VPB_c_396_n N_Y_c_548_n 0.00990863f $X=7.44 $Y=3.33 $X2=0 $Y2=0
cc_358 N_VPB_c_399_n N_Y_c_549_n 0.00822181f $X=1.195 $Y=2.085 $X2=0 $Y2=0
cc_359 N_VPB_c_400_n N_Y_c_549_n 0.00822181f $X=2.055 $Y=2.085 $X2=0 $Y2=0
cc_360 N_VPB_c_408_n N_Y_c_549_n 0.0128989f $X=1.925 $Y=3.33 $X2=0 $Y2=0
cc_361 N_VPB_c_396_n N_Y_c_549_n 0.00990863f $X=7.44 $Y=3.33 $X2=0 $Y2=0
cc_362 N_VPB_c_400_n N_Y_c_550_n 0.00822181f $X=2.055 $Y=2.085 $X2=0 $Y2=0
cc_363 N_VPB_c_401_n N_Y_c_550_n 0.00822181f $X=2.915 $Y=2.085 $X2=0 $Y2=0
cc_364 N_VPB_c_410_n N_Y_c_550_n 0.0128989f $X=2.785 $Y=3.33 $X2=0 $Y2=0
cc_365 N_VPB_c_396_n N_Y_c_550_n 0.00990863f $X=7.44 $Y=3.33 $X2=0 $Y2=0
cc_366 N_VPB_c_401_n N_Y_c_551_n 0.00822181f $X=2.915 $Y=2.085 $X2=0 $Y2=0
cc_367 N_VPB_c_402_n N_Y_c_551_n 0.00822181f $X=3.775 $Y=2.085 $X2=0 $Y2=0
cc_368 N_VPB_c_412_n N_Y_c_551_n 0.0128989f $X=3.645 $Y=3.33 $X2=0 $Y2=0
cc_369 N_VPB_c_396_n N_Y_c_551_n 0.00990863f $X=7.44 $Y=3.33 $X2=0 $Y2=0
cc_370 N_VPB_c_402_n N_Y_c_552_n 0.00822181f $X=3.775 $Y=2.085 $X2=0 $Y2=0
cc_371 N_VPB_c_403_n N_Y_c_552_n 0.0128989f $X=4.505 $Y=3.33 $X2=0 $Y2=0
cc_372 N_VPB_c_404_n N_Y_c_552_n 0.00822181f $X=4.635 $Y=2.085 $X2=0 $Y2=0
cc_373 N_VPB_c_396_n N_Y_c_552_n 0.00990863f $X=7.44 $Y=3.33 $X2=0 $Y2=0
cc_374 N_VPB_c_404_n N_Y_c_553_n 0.00822181f $X=4.635 $Y=2.085 $X2=0 $Y2=0
cc_375 N_VPB_c_405_n N_Y_c_553_n 0.00822181f $X=5.495 $Y=2.085 $X2=0 $Y2=0
cc_376 N_VPB_c_420_n N_Y_c_553_n 0.0128989f $X=5.365 $Y=3.33 $X2=0 $Y2=0
cc_377 N_VPB_c_396_n N_Y_c_553_n 0.00990863f $X=7.44 $Y=3.33 $X2=0 $Y2=0
cc_378 N_VPB_c_405_n N_Y_c_554_n 0.00822181f $X=5.495 $Y=2.085 $X2=0 $Y2=0
cc_379 N_VPB_c_406_n N_Y_c_554_n 0.00822181f $X=6.355 $Y=2.085 $X2=0 $Y2=0
cc_380 N_VPB_c_414_n N_Y_c_554_n 0.0128989f $X=6.225 $Y=3.33 $X2=0 $Y2=0
cc_381 N_VPB_c_396_n N_Y_c_554_n 0.00990863f $X=7.44 $Y=3.33 $X2=0 $Y2=0
cc_382 N_VPB_c_406_n N_Y_c_555_n 0.00822181f $X=6.355 $Y=2.085 $X2=0 $Y2=0
cc_383 N_VPB_c_417_n N_Y_c_555_n 0.0128989f $X=7.085 $Y=3.33 $X2=0 $Y2=0
cc_384 N_VPB_c_396_n N_Y_c_555_n 0.00990863f $X=7.44 $Y=3.33 $X2=0 $Y2=0
cc_385 N_VPB_M1004_s N_Y_c_626_n 0.00149321f $X=1.055 $Y=1.835 $X2=0 $Y2=0
cc_386 N_VPB_M1007_s N_Y_c_626_n 0.00149321f $X=1.915 $Y=1.835 $X2=0 $Y2=0
cc_387 N_VPB_M1011_s N_Y_c_626_n 0.00149321f $X=2.775 $Y=1.835 $X2=0 $Y2=0
cc_388 N_VPB_M1015_s N_Y_c_626_n 0.00149321f $X=3.635 $Y=1.835 $X2=0 $Y2=0
cc_389 N_VPB_M1020_s N_Y_c_626_n 0.00149321f $X=4.495 $Y=1.835 $X2=0 $Y2=0
cc_390 N_VPB_M1025_s N_Y_c_626_n 0.00149321f $X=5.355 $Y=1.835 $X2=0 $Y2=0
cc_391 N_VPB_M1028_s N_Y_c_626_n 0.00149321f $X=6.215 $Y=1.835 $X2=0 $Y2=0
cc_392 N_VPB_c_398_n N_Y_c_626_n 0.00691659f $X=0.335 $Y=2.085 $X2=0 $Y2=0
cc_393 N_VPB_c_399_n N_Y_c_626_n 0.025736f $X=1.195 $Y=2.085 $X2=0 $Y2=0
cc_394 N_VPB_c_400_n N_Y_c_626_n 0.025736f $X=2.055 $Y=2.085 $X2=0 $Y2=0
cc_395 N_VPB_c_401_n N_Y_c_626_n 0.025736f $X=2.915 $Y=2.085 $X2=0 $Y2=0
cc_396 N_VPB_c_402_n N_Y_c_626_n 0.025736f $X=3.775 $Y=2.085 $X2=0 $Y2=0
cc_397 N_VPB_c_404_n N_Y_c_626_n 0.025736f $X=4.635 $Y=2.085 $X2=0 $Y2=0
cc_398 N_VPB_c_405_n N_Y_c_626_n 0.025736f $X=5.495 $Y=2.085 $X2=0 $Y2=0
cc_399 N_VPB_c_406_n N_Y_c_626_n 0.025736f $X=6.355 $Y=2.085 $X2=0 $Y2=0
cc_400 N_VPB_c_407_n N_Y_c_626_n 0.00691659f $X=7.215 $Y=2.085 $X2=0 $Y2=0
cc_401 N_Y_c_552_n N_VGND_c_734_n 0.0113476f $X=4.205 $Y=0.47 $X2=0 $Y2=0
cc_402 N_Y_c_549_n N_VGND_c_739_n 0.0113476f $X=1.625 $Y=0.47 $X2=0 $Y2=0
cc_403 N_Y_c_550_n N_VGND_c_741_n 0.0113476f $X=2.485 $Y=0.47 $X2=0 $Y2=0
cc_404 N_Y_c_551_n N_VGND_c_743_n 0.0113476f $X=3.345 $Y=0.47 $X2=0 $Y2=0
cc_405 N_Y_c_554_n N_VGND_c_745_n 0.0113476f $X=5.925 $Y=0.47 $X2=0 $Y2=0
cc_406 N_Y_c_555_n N_VGND_c_748_n 0.0113476f $X=6.785 $Y=0.47 $X2=0 $Y2=0
cc_407 N_Y_c_548_n N_VGND_c_750_n 0.0113476f $X=0.765 $Y=0.47 $X2=0 $Y2=0
cc_408 N_Y_c_553_n N_VGND_c_751_n 0.0113476f $X=5.065 $Y=0.47 $X2=0 $Y2=0
cc_409 N_Y_M1001_s N_VGND_c_752_n 0.00304497f $X=0.625 $Y=0.235 $X2=0 $Y2=0
cc_410 N_Y_M1003_s N_VGND_c_752_n 0.00304497f $X=1.485 $Y=0.235 $X2=0 $Y2=0
cc_411 N_Y_M1008_s N_VGND_c_752_n 0.00304497f $X=2.345 $Y=0.235 $X2=0 $Y2=0
cc_412 N_Y_M1012_s N_VGND_c_752_n 0.00304497f $X=3.205 $Y=0.235 $X2=0 $Y2=0
cc_413 N_Y_M1016_s N_VGND_c_752_n 0.00304497f $X=4.065 $Y=0.235 $X2=0 $Y2=0
cc_414 N_Y_M1019_s N_VGND_c_752_n 0.00304497f $X=4.925 $Y=0.235 $X2=0 $Y2=0
cc_415 N_Y_M1023_s N_VGND_c_752_n 0.00304497f $X=5.785 $Y=0.235 $X2=0 $Y2=0
cc_416 N_Y_M1026_s N_VGND_c_752_n 0.00304497f $X=6.645 $Y=0.235 $X2=0 $Y2=0
cc_417 N_Y_c_548_n N_VGND_c_752_n 0.00977851f $X=0.765 $Y=0.47 $X2=0 $Y2=0
cc_418 N_Y_c_549_n N_VGND_c_752_n 0.00977851f $X=1.625 $Y=0.47 $X2=0 $Y2=0
cc_419 N_Y_c_550_n N_VGND_c_752_n 0.00977851f $X=2.485 $Y=0.47 $X2=0 $Y2=0
cc_420 N_Y_c_551_n N_VGND_c_752_n 0.00977851f $X=3.345 $Y=0.47 $X2=0 $Y2=0
cc_421 N_Y_c_552_n N_VGND_c_752_n 0.00977851f $X=4.205 $Y=0.47 $X2=0 $Y2=0
cc_422 N_Y_c_553_n N_VGND_c_752_n 0.00977851f $X=5.065 $Y=0.47 $X2=0 $Y2=0
cc_423 N_Y_c_554_n N_VGND_c_752_n 0.00977851f $X=5.925 $Y=0.47 $X2=0 $Y2=0
cc_424 N_Y_c_555_n N_VGND_c_752_n 0.00977851f $X=6.785 $Y=0.47 $X2=0 $Y2=0
