* File: sky130_fd_sc_lp__mux4_lp.pex.spice
* Created: Wed Sep  2 10:02:14 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__MUX4_LP%A_84_21# 1 2 9 13 15 17 19 20 21 24 28 32 34
c80 32 0 2.63772e-19 $X=2.07 $Y=2.2
r81 30 34 7.34436 $w=1.7e-07 $l=1.35477e-07 $layer=LI1_cond $X=2.07 $Y=1.26
+ $X2=2.065 $Y2=1.127
r82 30 32 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=2.07 $Y=1.26
+ $X2=2.07 $Y2=2.2
r83 26 34 7.34436 $w=1.7e-07 $l=1.34477e-07 $layer=LI1_cond $X=2.06 $Y=0.995
+ $X2=2.065 $Y2=1.127
r84 26 28 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=2.06 $Y=0.995 $X2=2.06
+ $Y2=0.495
r85 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.14
+ $Y=1.095 $X2=1.14 $Y2=1.095
r86 21 34 0.195364 $w=2.65e-07 $l=9e-08 $layer=LI1_cond $X=1.975 $Y=1.127
+ $X2=2.065 $Y2=1.127
r87 21 23 36.3128 $w=2.63e-07 $l=8.35e-07 $layer=LI1_cond $X=1.975 $Y=1.127
+ $X2=1.14 $Y2=1.127
r88 17 24 68.9507 $w=3.17e-07 $l=4.48865e-07 $layer=POLY_cond $X=0.855 $Y=0.73
+ $X2=1.042 $Y2=1.095
r89 17 19 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.855 $Y=0.73
+ $X2=0.855 $Y2=0.445
r90 16 20 9.46703 $w=1.5e-07 $l=1.25e-07 $layer=POLY_cond $X=0.67 $Y=1.185
+ $X2=0.545 $Y2=1.185
r91 15 24 13.6845 $w=3.17e-07 $l=9e-08 $layer=POLY_cond $X=1.042 $Y=1.185
+ $X2=1.042 $Y2=1.095
r92 15 16 156.394 $w=1.5e-07 $l=3.05e-07 $layer=POLY_cond $X=0.975 $Y=1.185
+ $X2=0.67 $Y2=1.185
r93 11 20 15.9654 $w=2e-07 $l=7.5e-08 $layer=POLY_cond $X=0.545 $Y=1.26
+ $X2=0.545 $Y2=1.185
r94 11 13 319.263 $w=2.5e-07 $l=1.285e-06 $layer=POLY_cond $X=0.545 $Y=1.26
+ $X2=0.545 $Y2=2.545
r95 7 20 15.9654 $w=2e-07 $l=9.68246e-08 $layer=POLY_cond $X=0.495 $Y=1.11
+ $X2=0.545 $Y2=1.185
r96 7 9 340.989 $w=1.5e-07 $l=6.65e-07 $layer=POLY_cond $X=0.495 $Y=1.11
+ $X2=0.495 $Y2=0.445
r97 2 32 600 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_PDIFF $count=1 $X=1.85
+ $Y=2.055 $X2=2.07 $Y2=2.2
r98 1 28 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.92
+ $Y=0.285 $X2=2.06 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__MUX4_LP%S1 1 4 5 7 8 10 11 12 13 15 17 18 20 22 24
+ 26 29 31 35 41 42 43 45 46 48
c150 48 0 1.2079e-19 $X=1.195 $Y=1.545
c151 45 0 9.8611e-20 $X=2.42 $Y=2.545
c152 24 0 1.80147e-19 $X=3.705 $Y=1
c153 18 0 1.91813e-19 $X=3.63 $Y=1.075
c154 12 0 3.83947e-20 $X=3.025 $Y=1.525
c155 4 0 1.60848e-19 $X=1.62 $Y=1.47
c156 1 0 1.42982e-19 $X=1.545 $Y=1.545
r157 52 54 24.0142 $w=2.81e-07 $l=1.4e-07 $layer=POLY_cond $X=2.45 $Y=1.732
+ $X2=2.59 $Y2=1.732
r158 46 56 5.76222 $w=3.38e-07 $l=1.7e-07 $layer=LI1_cond $X=2.59 $Y=1.72
+ $X2=2.42 $Y2=1.72
r159 46 54 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.59
+ $Y=1.725 $X2=2.59 $Y2=1.725
r160 44 56 4.80115 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=2.42 $Y=1.89
+ $X2=2.42 $Y2=1.72
r161 44 45 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=2.42 $Y=1.89
+ $X2=2.42 $Y2=2.545
r162 42 45 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.335 $Y=2.63
+ $X2=2.42 $Y2=2.545
r163 42 43 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=2.335 $Y=2.63
+ $X2=1.805 $Y2=2.63
r164 41 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.72 $Y=2.545
+ $X2=1.805 $Y2=2.63
r165 40 41 48.6043 $w=1.68e-07 $l=7.45e-07 $layer=LI1_cond $X=1.72 $Y=1.8
+ $X2=1.72 $Y2=2.545
r166 38 48 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=1.195 $Y=1.635
+ $X2=1.195 $Y2=1.545
r167 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.195
+ $Y=1.635 $X2=1.195 $Y2=1.635
r168 35 40 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.635 $Y=1.635
+ $X2=1.72 $Y2=1.8
r169 35 37 15.3659 $w=3.28e-07 $l=4.4e-07 $layer=LI1_cond $X=1.635 $Y=1.635
+ $X2=1.195 $Y2=1.635
r170 27 29 115.372 $w=1.5e-07 $l=2.25e-07 $layer=POLY_cond $X=1.62 $Y=0.855
+ $X2=1.845 $Y2=0.855
r171 24 26 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.705 $Y=1 $X2=3.705
+ $Y2=0.715
r172 20 32 169.213 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=3.675 $Y=1.525
+ $X2=3.345 $Y2=1.525
r173 20 22 247.211 $w=2.5e-07 $l=9.95e-07 $layer=POLY_cond $X=3.675 $Y=1.6
+ $X2=3.675 $Y2=2.595
r174 19 31 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.42 $Y=1.075
+ $X2=3.345 $Y2=1.075
r175 18 24 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.63 $Y=1.075
+ $X2=3.705 $Y2=1
r176 18 19 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=3.63 $Y=1.075
+ $X2=3.42 $Y2=1.075
r177 17 32 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.345 $Y=1.45
+ $X2=3.345 $Y2=1.525
r178 16 31 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.345 $Y=1.15
+ $X2=3.345 $Y2=1.075
r179 16 17 153.83 $w=1.5e-07 $l=3e-07 $layer=POLY_cond $X=3.345 $Y=1.15
+ $X2=3.345 $Y2=1.45
r180 13 31 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.345 $Y=1
+ $X2=3.345 $Y2=1.075
r181 13 15 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.345 $Y=1 $X2=3.345
+ $Y2=0.715
r182 12 54 85.0291 $w=2.81e-07 $l=5.2846e-07 $layer=POLY_cond $X=3.025 $Y=1.525
+ $X2=2.59 $Y2=1.732
r183 11 32 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.27 $Y=1.525
+ $X2=3.345 $Y2=1.525
r184 11 12 125.628 $w=1.5e-07 $l=2.45e-07 $layer=POLY_cond $X=3.27 $Y=1.525
+ $X2=3.025 $Y2=1.525
r185 8 52 5.60901 $w=2.5e-07 $l=2.83e-07 $layer=POLY_cond $X=2.45 $Y=2.015
+ $X2=2.45 $Y2=1.732
r186 8 10 104.112 $w=2.5e-07 $l=5.4e-07 $layer=POLY_cond $X=2.45 $Y=2.015
+ $X2=2.45 $Y2=2.555
r187 5 29 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.845 $Y=0.78
+ $X2=1.845 $Y2=0.855
r188 5 7 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=1.845 $Y=0.78
+ $X2=1.845 $Y2=0.495
r189 3 27 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.62 $Y=0.93
+ $X2=1.62 $Y2=0.855
r190 3 4 276.894 $w=1.5e-07 $l=5.4e-07 $layer=POLY_cond $X=1.62 $Y=0.93 $X2=1.62
+ $Y2=1.47
r191 2 48 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.36 $Y=1.545
+ $X2=1.195 $Y2=1.545
r192 1 4 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.545 $Y=1.545
+ $X2=1.62 $Y2=1.47
r193 1 2 94.8617 $w=1.5e-07 $l=1.85e-07 $layer=POLY_cond $X=1.545 $Y=1.545
+ $X2=1.36 $Y2=1.545
.ends

.subckt PM_SKY130_FD_SC_LP__MUX4_LP%A_320_366# 1 2 7 9 11 14 18 20 27 30 31 35
+ 38
c87 38 0 1.67023e-19 $X=2.275 $Y=1.155
c88 20 0 1.60848e-19 $X=2.885 $Y=1.155
c89 18 0 9.8611e-20 $X=2.01 $Y=1.905
c90 14 0 1.1902e-19 $X=2.275 $Y=0.495
r91 32 35 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=3.13 $Y=1.82 $X2=3.33
+ $Y2=1.82
r92 30 32 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.13 $Y=1.655
+ $X2=3.13 $Y2=1.82
r93 29 31 6.46576 $w=2.5e-07 $l=2.0106e-07 $layer=LI1_cond $X=3.13 $Y=1.32
+ $X2=3.05 $Y2=1.155
r94 29 30 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=3.13 $Y=1.32
+ $X2=3.13 $Y2=1.655
r95 25 31 6.46576 $w=2.5e-07 $l=1.65e-07 $layer=LI1_cond $X=3.05 $Y=0.99
+ $X2=3.05 $Y2=1.155
r96 25 27 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=3.05 $Y=0.99
+ $X2=3.05 $Y2=0.78
r97 23 38 41.0795 $w=2.64e-07 $l=2.25e-07 $layer=POLY_cond $X=2.5 $Y=1.155
+ $X2=2.275 $Y2=1.155
r98 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.5
+ $Y=1.155 $X2=2.5 $Y2=1.155
r99 20 31 0.364692 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=2.885 $Y=1.155
+ $X2=3.05 $Y2=1.155
r100 20 22 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=2.885 $Y=1.155
+ $X2=2.5 $Y2=1.155
r101 12 38 15.9823 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.275 $Y=0.99
+ $X2=2.275 $Y2=1.155
r102 12 14 253.819 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=2.275 $Y=0.99
+ $X2=2.275 $Y2=0.495
r103 11 18 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.01 $Y=1.83
+ $X2=2.01 $Y2=1.905
r104 10 38 48.3826 $w=2.64e-07 $l=3.37565e-07 $layer=POLY_cond $X=2.01 $Y=1.32
+ $X2=2.275 $Y2=1.155
r105 10 11 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=2.01 $Y=1.32
+ $X2=2.01 $Y2=1.83
r106 7 18 146.138 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=1.725 $Y=1.905
+ $X2=2.01 $Y2=1.905
r107 7 9 110.86 $w=2.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.725 $Y=1.98
+ $X2=1.725 $Y2=2.555
r108 2 35 600 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=3.185
+ $Y=1.675 $X2=3.33 $Y2=1.82
r109 1 27 182 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=1 $X=2.905
+ $Y=0.505 $X2=3.05 $Y2=0.78
.ends

.subckt PM_SKY130_FD_SC_LP__MUX4_LP%A3 3 6 7 9 12 14 15 23
c47 12 0 1.04379e-19 $X=4.5 $Y=1.075
r48 22 23 8.74306 $w=3.3e-07 $l=5e-08 $layer=POLY_cond $X=4.365 $Y=1.715
+ $X2=4.415 $Y2=1.715
r49 19 22 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=4.185 $Y=1.715
+ $X2=4.365 $Y2=1.715
r50 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.185
+ $Y=1.715 $X2=4.185 $Y2=1.715
r51 15 20 9.57875 $w=3.83e-07 $l=3.2e-07 $layer=LI1_cond $X=4.157 $Y=2.035
+ $X2=4.157 $Y2=1.715
r52 14 20 1.49668 $w=3.83e-07 $l=5e-08 $layer=LI1_cond $X=4.157 $Y=1.665
+ $X2=4.157 $Y2=1.715
r53 10 12 43.5851 $w=1.5e-07 $l=8.5e-08 $layer=POLY_cond $X=4.415 $Y=1.075
+ $X2=4.5 $Y2=1.075
r54 7 12 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.5 $Y=1 $X2=4.5
+ $Y2=1.075
r55 7 9 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=4.5 $Y=1 $X2=4.5
+ $Y2=0.715
r56 6 23 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.415 $Y=1.55
+ $X2=4.415 $Y2=1.715
r57 5 10 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.415 $Y=1.15
+ $X2=4.415 $Y2=1.075
r58 5 6 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=4.415 $Y=1.15 $X2=4.415
+ $Y2=1.55
r59 1 22 9.34494 $w=2.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.365 $Y=1.88
+ $X2=4.365 $Y2=1.715
r60 1 3 177.644 $w=2.5e-07 $l=7.15e-07 $layer=POLY_cond $X=4.365 $Y=1.88
+ $X2=4.365 $Y2=2.595
.ends

.subckt PM_SKY130_FD_SC_LP__MUX4_LP%S0 3 6 10 14 16 18 23 25 27 31 36 38 40 43
+ 44 45 48 49 52 53 54 55 56 57 58 59 63 65 66 67 68 74 83 88 89 90 94
c210 59 0 4.86698e-20 $X=5.98 $Y=1.36
c211 58 0 1.89825e-19 $X=5.565 $Y=1.245
c212 57 0 1.04379e-19 $X=5.395 $Y=1.245
c213 55 0 1.01928e-19 $X=8.265 $Y=2.15
c214 54 0 1.70305e-19 $X=7.61 $Y=2.63
c215 53 0 1.56872e-19 $X=8.18 $Y=2.63
c216 40 0 3.61697e-19 $X=6.325 $Y=1.36
c217 10 0 8.47076e-20 $X=7.385 $Y=0.445
r218 92 94 1.17263 $w=5.08e-07 $l=5e-08 $layer=LI1_cond $X=8.35 $Y=1.895 $X2=8.4
+ $Y2=1.895
r219 88 91 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=9.455 $Y=1.77
+ $X2=9.455 $Y2=1.935
r220 88 90 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=9.455 $Y=1.77
+ $X2=9.455 $Y2=1.605
r221 88 89 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.455
+ $Y=1.77 $X2=9.455 $Y2=1.77
r222 83 86 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.345 $Y=1.77
+ $X2=8.345 $Y2=1.935
r223 68 89 2.22799 $w=5.08e-07 $l=9.5e-08 $layer=LI1_cond $X=9.36 $Y=1.895
+ $X2=9.455 $Y2=1.895
r224 67 68 11.2572 $w=5.08e-07 $l=4.8e-07 $layer=LI1_cond $X=8.88 $Y=1.895
+ $X2=9.36 $Y2=1.895
r225 66 92 2.32863 $w=5.1e-07 $l=8.5e-08 $layer=LI1_cond $X=8.265 $Y=1.895
+ $X2=8.35 $Y2=1.895
r226 66 67 10.8585 $w=5.08e-07 $l=4.63e-07 $layer=LI1_cond $X=8.417 $Y=1.895
+ $X2=8.88 $Y2=1.895
r227 66 94 0.398693 $w=5.08e-07 $l=1.7e-08 $layer=LI1_cond $X=8.417 $Y=1.895
+ $X2=8.4 $Y2=1.895
r228 66 83 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.345
+ $Y=1.77 $X2=8.345 $Y2=1.77
r229 63 78 32.0725 $w=3.45e-07 $l=1.65e-07 $layer=POLY_cond $X=5.972 $Y=1.595
+ $X2=5.972 $Y2=1.76
r230 62 63 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.98
+ $Y=1.595 $X2=5.98 $Y2=1.595
r231 59 62 8.20679 $w=3.28e-07 $l=2.35e-07 $layer=LI1_cond $X=5.98 $Y=1.36
+ $X2=5.98 $Y2=1.595
r232 57 58 8.63679 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=5.395 $Y=1.245
+ $X2=5.565 $Y2=1.245
r233 55 66 6.98588 $w=1.7e-07 $l=2.55e-07 $layer=LI1_cond $X=8.265 $Y=2.15
+ $X2=8.265 $Y2=1.895
r234 55 56 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=8.265 $Y=2.15
+ $X2=8.265 $Y2=2.545
r235 53 56 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.18 $Y=2.63
+ $X2=8.265 $Y2=2.545
r236 53 54 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=8.18 $Y=2.63
+ $X2=7.61 $Y2=2.63
r237 52 54 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.525 $Y=2.545
+ $X2=7.61 $Y2=2.63
r238 51 65 3.70735 $w=2.5e-07 $l=1.18427e-07 $layer=LI1_cond $X=7.525 $Y=1.76
+ $X2=7.445 $Y2=1.675
r239 51 52 51.2139 $w=1.68e-07 $l=7.85e-07 $layer=LI1_cond $X=7.525 $Y=1.76
+ $X2=7.525 $Y2=2.545
r240 49 80 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.445 $Y=1.245
+ $X2=7.445 $Y2=1.08
r241 48 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.445
+ $Y=1.245 $X2=7.445 $Y2=1.245
r242 46 65 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.445 $Y=1.59
+ $X2=7.445 $Y2=1.675
r243 46 48 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=7.445 $Y=1.59
+ $X2=7.445 $Y2=1.245
r244 44 65 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.28 $Y=1.675
+ $X2=7.445 $Y2=1.675
r245 44 45 51.2139 $w=1.68e-07 $l=7.85e-07 $layer=LI1_cond $X=7.28 $Y=1.675
+ $X2=6.495 $Y2=1.675
r246 43 45 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.41 $Y=1.59
+ $X2=6.495 $Y2=1.675
r247 42 43 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=6.41 $Y=1.445
+ $X2=6.41 $Y2=1.59
r248 41 59 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.145 $Y=1.36
+ $X2=5.98 $Y2=1.36
r249 40 42 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.325 $Y=1.36
+ $X2=6.41 $Y2=1.445
r250 40 41 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=6.325 $Y=1.36
+ $X2=6.145 $Y2=1.36
r251 38 59 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.815 $Y=1.36
+ $X2=5.98 $Y2=1.36
r252 38 58 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=5.815 $Y=1.36
+ $X2=5.565 $Y2=1.36
r253 36 74 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.035 $Y=1.21
+ $X2=5.035 $Y2=1.045
r254 35 57 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=5.035 $Y=1.21
+ $X2=5.395 $Y2=1.21
r255 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.035
+ $Y=1.21 $X2=5.035 $Y2=1.21
r256 30 31 112.809 $w=1.5e-07 $l=2.2e-07 $layer=POLY_cond $X=9.365 $Y=0.805
+ $X2=9.585 $Y2=0.805
r257 28 30 71.7872 $w=1.5e-07 $l=1.4e-07 $layer=POLY_cond $X=9.225 $Y=0.805
+ $X2=9.365 $Y2=0.805
r258 25 31 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.585 $Y=0.73
+ $X2=9.585 $Y2=0.805
r259 25 27 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=9.585 $Y=0.73
+ $X2=9.585 $Y2=0.445
r260 23 91 163.979 $w=2.5e-07 $l=6.6e-07 $layer=POLY_cond $X=9.415 $Y=2.595
+ $X2=9.415 $Y2=1.935
r261 19 30 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.365 $Y=0.88
+ $X2=9.365 $Y2=0.805
r262 19 90 371.755 $w=1.5e-07 $l=7.25e-07 $layer=POLY_cond $X=9.365 $Y=0.88
+ $X2=9.365 $Y2=1.605
r263 16 28 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.225 $Y=0.73
+ $X2=9.225 $Y2=0.805
r264 16 18 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=9.225 $Y=0.73
+ $X2=9.225 $Y2=0.445
r265 14 86 163.979 $w=2.5e-07 $l=6.6e-07 $layer=POLY_cond $X=8.335 $Y=2.595
+ $X2=8.335 $Y2=1.935
r266 10 80 325.606 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=7.385 $Y=0.445
+ $X2=7.385 $Y2=1.08
r267 6 78 207.459 $w=2.5e-07 $l=8.35e-07 $layer=POLY_cond $X=5.925 $Y=2.595
+ $X2=5.925 $Y2=1.76
r268 3 74 106.04 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=4.975 $Y=0.715
+ $X2=4.975 $Y2=1.045
.ends

.subckt PM_SKY130_FD_SC_LP__MUX4_LP%A_946_317# 1 2 9 11 15 19 21 22 24 25 27 29
+ 30 32 35 36 37 38 41 42 43 48 51 53 58 64 66 68 69 75
c193 75 0 4.86698e-20 $X=5.215 $Y=1.75
c194 66 0 8.47076e-20 $X=8.47 $Y=0.897
c195 32 0 1.3249e-19 $X=7.09 $Y=2.025
r196 63 66 8.65224 $w=2.63e-07 $l=1.65e-07 $layer=LI1_cond $X=8.305 $Y=0.897
+ $X2=8.47 $Y2=0.897
r197 63 64 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.305
+ $Y=0.93 $X2=8.305 $Y2=0.93
r198 58 60 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=5.55 $Y=1.83
+ $X2=5.55 $Y2=2.025
r199 54 75 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.05 $Y=1.75
+ $X2=5.215 $Y2=1.75
r200 54 72 34.0979 $w=3.3e-07 $l=1.95e-07 $layer=POLY_cond $X=5.05 $Y=1.75
+ $X2=4.855 $Y2=1.75
r201 53 56 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=5.05 $Y=1.75 $X2=5.05
+ $Y2=1.83
r202 53 54 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.05
+ $Y=1.75 $X2=5.05 $Y2=1.75
r203 51 68 3.03453 $w=3.12e-07 $l=1.80566e-07 $layer=LI1_cond $X=9.885 $Y=2.33
+ $X2=9.742 $Y2=2.415
r204 50 69 3.67481 $w=2.52e-07 $l=1.19499e-07 $layer=LI1_cond $X=9.885 $Y=1.03
+ $X2=9.802 $Y2=0.945
r205 50 51 84.8128 $w=1.68e-07 $l=1.3e-06 $layer=LI1_cond $X=9.885 $Y=1.03
+ $X2=9.885 $Y2=2.33
r206 46 69 3.67481 $w=2.52e-07 $l=8.5e-08 $layer=LI1_cond $X=9.802 $Y=0.86
+ $X2=9.802 $Y2=0.945
r207 46 48 13.4165 $w=3.33e-07 $l=3.9e-07 $layer=LI1_cond $X=9.802 $Y=0.86
+ $X2=9.802 $Y2=0.47
r208 42 68 3.60271 $w=1.7e-07 $l=2.27e-07 $layer=LI1_cond $X=9.515 $Y=2.415
+ $X2=9.742 $Y2=2.415
r209 42 43 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=9.515 $Y=2.415
+ $X2=8.805 $Y2=2.415
r210 40 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.72 $Y=2.5
+ $X2=8.805 $Y2=2.415
r211 40 41 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=8.72 $Y=2.5
+ $X2=8.72 $Y2=2.895
r212 38 69 2.79892 $w=1.7e-07 $l=1.67e-07 $layer=LI1_cond $X=9.635 $Y=0.945
+ $X2=9.802 $Y2=0.945
r213 38 66 76.0053 $w=1.68e-07 $l=1.165e-06 $layer=LI1_cond $X=9.635 $Y=0.945
+ $X2=8.47 $Y2=0.945
r214 36 41 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.635 $Y=2.98
+ $X2=8.72 $Y2=2.895
r215 36 37 89.7059 $w=1.68e-07 $l=1.375e-06 $layer=LI1_cond $X=8.635 $Y=2.98
+ $X2=7.26 $Y2=2.98
r216 35 37 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.175 $Y=2.895
+ $X2=7.26 $Y2=2.98
r217 34 35 51.2139 $w=1.68e-07 $l=7.85e-07 $layer=LI1_cond $X=7.175 $Y=2.11
+ $X2=7.175 $Y2=2.895
r218 33 60 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.635 $Y=2.025
+ $X2=5.55 $Y2=2.025
r219 32 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.09 $Y=2.025
+ $X2=7.175 $Y2=2.11
r220 32 33 94.9251 $w=1.68e-07 $l=1.455e-06 $layer=LI1_cond $X=7.09 $Y=2.025
+ $X2=5.635 $Y2=2.025
r221 31 56 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.215 $Y=1.83
+ $X2=5.05 $Y2=1.83
r222 30 58 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.465 $Y=1.83
+ $X2=5.55 $Y2=1.83
r223 30 31 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=5.465 $Y=1.83
+ $X2=5.215 $Y2=1.83
r224 28 64 53.3327 $w=3.3e-07 $l=3.05e-07 $layer=POLY_cond $X=8 $Y=0.93
+ $X2=8.305 $Y2=0.93
r225 28 29 5.03009 $w=3.3e-07 $l=1.8735e-07 $layer=POLY_cond $X=8 $Y=0.93
+ $X2=7.82 $Y2=0.945
r226 25 29 37.0704 $w=1.5e-07 $l=2.26495e-07 $layer=POLY_cond $X=7.925 $Y=0.765
+ $X2=7.82 $Y2=0.945
r227 25 27 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=7.925 $Y=0.765
+ $X2=7.925 $Y2=0.445
r228 23 29 37.0704 $w=1.5e-07 $l=1.83712e-07 $layer=POLY_cond $X=7.895 $Y=1.095
+ $X2=7.82 $Y2=0.945
r229 23 24 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=7.895 $Y=1.095
+ $X2=7.895 $Y2=1.65
r230 21 24 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.82 $Y=1.725
+ $X2=7.895 $Y2=1.65
r231 21 22 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.82 $Y=1.725
+ $X2=7.655 $Y2=1.725
r232 17 22 29.1797 $w=1.5e-07 $l=1.58114e-07 $layer=POLY_cond $X=7.53 $Y=1.8
+ $X2=7.655 $Y2=1.725
r233 17 19 197.521 $w=2.5e-07 $l=7.95e-07 $layer=POLY_cond $X=7.53 $Y=1.8
+ $X2=7.53 $Y2=2.595
r234 13 15 584.553 $w=1.5e-07 $l=1.14e-06 $layer=POLY_cond $X=5.485 $Y=1.585
+ $X2=5.485 $Y2=0.445
r235 11 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.41 $Y=1.66
+ $X2=5.485 $Y2=1.585
r236 11 75 99.9894 $w=1.5e-07 $l=1.95e-07 $layer=POLY_cond $X=5.41 $Y=1.66
+ $X2=5.215 $Y2=1.66
r237 7 72 9.34494 $w=2.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.855 $Y=1.915
+ $X2=4.855 $Y2=1.75
r238 7 9 168.948 $w=2.5e-07 $l=6.8e-07 $layer=POLY_cond $X=4.855 $Y=1.915
+ $X2=4.855 $Y2=2.595
r239 2 68 300 $w=1.7e-07 $l=4.64758e-07 $layer=licon1_PDIFF $count=2 $X=9.54
+ $Y=2.095 $X2=9.68 $Y2=2.495
r240 1 48 182 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=1 $X=9.66
+ $Y=0.235 $X2=9.8 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_LP__MUX4_LP%A2 3 4 8 10 12 13 16 18
c54 16 0 1.89825e-19 $X=5.935 $Y=0.93
c55 13 0 9.51642e-21 $X=6 $Y=0.925
r56 16 19 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=5.935 $Y=0.93
+ $X2=5.935 $Y2=1.02
r57 16 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.935 $Y=0.93
+ $X2=5.935 $Y2=0.765
r58 13 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.935
+ $Y=0.93 $X2=5.935 $Y2=0.93
r59 8 12 40.9178 $w=2.5e-07 $l=1.25e-07 $layer=POLY_cond $X=6.48 $Y=1.775
+ $X2=6.48 $Y2=1.65
r60 8 10 203.732 $w=2.5e-07 $l=8.2e-07 $layer=POLY_cond $X=6.48 $Y=1.775
+ $X2=6.48 $Y2=2.595
r61 6 12 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=6.43 $Y=1.095
+ $X2=6.43 $Y2=1.65
r62 5 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.1 $Y=1.02
+ $X2=5.935 $Y2=1.02
r63 4 6 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.355 $Y=1.02
+ $X2=6.43 $Y2=1.095
r64 4 5 130.755 $w=1.5e-07 $l=2.55e-07 $layer=POLY_cond $X=6.355 $Y=1.02 $X2=6.1
+ $Y2=1.02
r65 3 18 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=5.875 $Y=0.445
+ $X2=5.875 $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_LP__MUX4_LP%A1 3 5 9 11 12 15
c43 15 0 1.78025e-19 $X=6.905 $Y=1.245
c44 11 0 1.93189e-19 $X=7.04 $Y=1.65
c45 5 0 1.70305e-19 $X=7.04 $Y=2.595
c46 3 0 5.29209e-20 $X=7.04 $Y=1.775
r47 15 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.905 $Y=1.245
+ $X2=6.905 $Y2=1.41
r48 15 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.905 $Y=1.245
+ $X2=6.905 $Y2=1.08
r49 12 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.905
+ $Y=1.245 $X2=6.905 $Y2=1.245
r50 11 18 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=6.99 $Y=1.65
+ $X2=6.99 $Y2=1.41
r51 9 17 325.606 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=6.995 $Y=0.445
+ $X2=6.995 $Y2=1.08
r52 3 11 40.9178 $w=2.5e-07 $l=1.25e-07 $layer=POLY_cond $X=7.04 $Y=1.775
+ $X2=7.04 $Y2=1.65
r53 3 5 203.732 $w=2.5e-07 $l=8.2e-07 $layer=POLY_cond $X=7.04 $Y=1.775 $X2=7.04
+ $Y2=2.595
.ends

.subckt PM_SKY130_FD_SC_LP__MUX4_LP%A0 3 7 9 10 11 16
c41 7 0 1.56872e-19 $X=8.875 $Y=2.595
r42 16 19 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.885 $Y=1.335
+ $X2=8.885 $Y2=1.5
r43 16 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.885 $Y=1.335
+ $X2=8.885 $Y2=1.17
r44 10 11 22.1269 $w=2.48e-07 $l=4.8e-07 $layer=LI1_cond $X=8.88 $Y=1.335
+ $X2=9.36 $Y2=1.335
r45 10 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.885
+ $Y=1.335 $X2=8.885 $Y2=1.335
r46 9 10 22.1269 $w=2.48e-07 $l=4.8e-07 $layer=LI1_cond $X=8.4 $Y=1.335 $X2=8.88
+ $Y2=1.335
r47 7 19 272.057 $w=2.5e-07 $l=1.095e-06 $layer=POLY_cond $X=8.875 $Y=2.595
+ $X2=8.875 $Y2=1.5
r48 3 18 371.755 $w=1.5e-07 $l=7.25e-07 $layer=POLY_cond $X=8.795 $Y=0.445
+ $X2=8.795 $Y2=1.17
.ends

.subckt PM_SKY130_FD_SC_LP__MUX4_LP%X 1 2 7 8 9 10 11 12 13
r16 13 40 4.36531 $w=3.28e-07 $l=1.25e-07 $layer=LI1_cond $X=0.28 $Y=2.775
+ $X2=0.28 $Y2=2.9
r17 12 13 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.28 $Y=2.405
+ $X2=0.28 $Y2=2.775
r18 12 34 7.50834 $w=3.28e-07 $l=2.15e-07 $layer=LI1_cond $X=0.28 $Y=2.405
+ $X2=0.28 $Y2=2.19
r19 11 34 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=0.28 $Y=2.035
+ $X2=0.28 $Y2=2.19
r20 10 11 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.28 $Y=1.665
+ $X2=0.28 $Y2=2.035
r21 9 10 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.28 $Y=1.295
+ $X2=0.28 $Y2=1.665
r22 8 9 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.28 $Y=0.925 $X2=0.28
+ $Y2=1.295
r23 7 8 15.8897 $w=3.28e-07 $l=4.55e-07 $layer=LI1_cond $X=0.28 $Y=0.47 $X2=0.28
+ $Y2=0.925
r24 2 40 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.045 $X2=0.28 $Y2=2.9
r25 2 34 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.045 $X2=0.28 $Y2=2.19
r26 1 7 182 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.28 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_LP__MUX4_LP%VPWR 1 2 3 4 17 21 25 29 32 33 35 36 37 39
+ 61 62 65 68
r98 68 69 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r99 65 66 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r100 61 62 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r101 59 62 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=9.84 $Y2=3.33
r102 58 59 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r103 56 59 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=8.88 $Y2=3.33
r104 55 58 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=6.96 $Y=3.33
+ $X2=8.88 $Y2=3.33
r105 55 56 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r106 53 56 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=6.96 $Y2=3.33
r107 52 53 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r108 50 69 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=4.08 $Y2=3.33
r109 49 52 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=4.56 $Y=3.33
+ $X2=6.48 $Y2=3.33
r110 49 50 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r111 47 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.185 $Y=3.33
+ $X2=4.02 $Y2=3.33
r112 47 49 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=4.185 $Y=3.33
+ $X2=4.56 $Y2=3.33
r113 46 69 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r114 45 46 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r115 43 46 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=3.6 $Y2=3.33
r116 43 66 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r117 42 45 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=1.2 $Y=3.33 $X2=3.6
+ $Y2=3.33
r118 42 43 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r119 40 65 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.975 $Y=3.33
+ $X2=0.81 $Y2=3.33
r120 40 42 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=0.975 $Y=3.33
+ $X2=1.2 $Y2=3.33
r121 39 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.855 $Y=3.33
+ $X2=4.02 $Y2=3.33
r122 39 45 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=3.855 $Y=3.33
+ $X2=3.6 $Y2=3.33
r123 37 53 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=6.48 $Y2=3.33
r124 37 50 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=4.56 $Y2=3.33
r125 35 58 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=8.985 $Y=3.33
+ $X2=8.88 $Y2=3.33
r126 35 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.985 $Y=3.33
+ $X2=9.15 $Y2=3.33
r127 34 61 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=9.315 $Y=3.33
+ $X2=9.84 $Y2=3.33
r128 34 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.315 $Y=3.33
+ $X2=9.15 $Y2=3.33
r129 32 52 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=6.58 $Y=3.33 $X2=6.48
+ $Y2=3.33
r130 32 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.58 $Y=3.33
+ $X2=6.745 $Y2=3.33
r131 31 55 3.26203 $w=1.68e-07 $l=5e-08 $layer=LI1_cond $X=6.91 $Y=3.33 $X2=6.96
+ $Y2=3.33
r132 31 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.91 $Y=3.33
+ $X2=6.745 $Y2=3.33
r133 27 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.15 $Y=3.245
+ $X2=9.15 $Y2=3.33
r134 27 29 12.2229 $w=3.28e-07 $l=3.5e-07 $layer=LI1_cond $X=9.15 $Y=3.245
+ $X2=9.15 $Y2=2.895
r135 23 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.745 $Y=3.245
+ $X2=6.745 $Y2=3.33
r136 23 25 27.5888 $w=3.28e-07 $l=7.9e-07 $layer=LI1_cond $X=6.745 $Y=3.245
+ $X2=6.745 $Y2=2.455
r137 19 68 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.02 $Y=3.245
+ $X2=4.02 $Y2=3.33
r138 19 21 7.50834 $w=3.28e-07 $l=2.15e-07 $layer=LI1_cond $X=4.02 $Y=3.245
+ $X2=4.02 $Y2=3.03
r139 15 65 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.81 $Y=3.245
+ $X2=0.81 $Y2=3.33
r140 15 17 26.1919 $w=3.28e-07 $l=7.5e-07 $layer=LI1_cond $X=0.81 $Y=3.245
+ $X2=0.81 $Y2=2.495
r141 4 29 600 $w=1.7e-07 $l=8.7178e-07 $layer=licon1_PDIFF $count=1 $X=9
+ $Y=2.095 $X2=9.15 $Y2=2.895
r142 3 25 300 $w=1.7e-07 $l=4.24264e-07 $layer=licon1_PDIFF $count=2 $X=6.605
+ $Y=2.095 $X2=6.745 $Y2=2.455
r143 2 21 600 $w=1.7e-07 $l=1.03919e-06 $layer=licon1_PDIFF $count=1 $X=3.8
+ $Y=2.095 $X2=4.02 $Y2=3.03
r144 1 17 300 $w=1.7e-07 $l=5.15267e-07 $layer=licon1_PDIFF $count=2 $X=0.67
+ $Y=2.045 $X2=0.81 $Y2=2.495
.ends

.subckt PM_SKY130_FD_SC_LP__MUX4_LP%A_245_411# 1 2 3 4 14 15 16 17 18 20 22 23
+ 27 30 31 32 34 35 37 39 43 49 50
r146 41 50 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.12 $Y=2.515
+ $X2=5.12 $Y2=2.6
r147 41 43 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=5.12 $Y=2.515
+ $X2=5.12 $Y2=2.26
r148 40 49 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.705 $Y=2.6
+ $X2=4.62 $Y2=2.6
r149 39 50 3.80956 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.955 $Y=2.6
+ $X2=5.12 $Y2=2.6
r150 39 40 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=4.955 $Y=2.6
+ $X2=4.705 $Y2=2.6
r151 35 37 22.3574 $w=2.48e-07 $l=4.85e-07 $layer=LI1_cond $X=4.705 $Y=0.74
+ $X2=5.19 $Y2=0.74
r152 34 49 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.62 $Y=2.515
+ $X2=4.62 $Y2=2.6
r153 33 35 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=4.62 $Y=0.865
+ $X2=4.705 $Y2=0.74
r154 33 34 107.647 $w=1.68e-07 $l=1.65e-06 $layer=LI1_cond $X=4.62 $Y=0.865
+ $X2=4.62 $Y2=2.515
r155 31 49 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.535 $Y=2.6
+ $X2=4.62 $Y2=2.6
r156 31 32 81.5508 $w=1.68e-07 $l=1.25e-06 $layer=LI1_cond $X=4.535 $Y=2.6
+ $X2=3.285 $Y2=2.6
r157 29 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.2 $Y=2.685
+ $X2=3.285 $Y2=2.6
r158 29 30 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=3.2 $Y=2.685
+ $X2=3.2 $Y2=2.895
r159 25 27 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=1.63 $Y=0.645
+ $X2=1.63 $Y2=0.495
r160 24 48 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.455 $Y=2.98
+ $X2=1.33 $Y2=2.98
r161 23 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.115 $Y=2.98
+ $X2=3.2 $Y2=2.895
r162 23 24 108.299 $w=1.68e-07 $l=1.66e-06 $layer=LI1_cond $X=3.115 $Y=2.98
+ $X2=1.455 $Y2=2.98
r163 20 48 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.33 $Y=2.895
+ $X2=1.33 $Y2=2.98
r164 20 22 32.0379 $w=2.48e-07 $l=6.95e-07 $layer=LI1_cond $X=1.33 $Y=2.895
+ $X2=1.33 $Y2=2.2
r165 19 22 2.30489 $w=2.48e-07 $l=5e-08 $layer=LI1_cond $X=1.33 $Y=2.15 $X2=1.33
+ $Y2=2.2
r166 17 19 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.205 $Y=2.065
+ $X2=1.33 $Y2=2.15
r167 17 18 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=1.205 $Y=2.065
+ $X2=0.795 $Y2=2.065
r168 15 25 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.465 $Y=0.73
+ $X2=1.63 $Y2=0.645
r169 15 16 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.465 $Y=0.73
+ $X2=0.795 $Y2=0.73
r170 14 18 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.71 $Y=1.98
+ $X2=0.795 $Y2=2.065
r171 13 16 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.71 $Y=0.815
+ $X2=0.795 $Y2=0.73
r172 13 14 76.0053 $w=1.68e-07 $l=1.165e-06 $layer=LI1_cond $X=0.71 $Y=0.815
+ $X2=0.71 $Y2=1.98
r173 4 43 300 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_PDIFF $count=2 $X=4.98
+ $Y=2.095 $X2=5.12 $Y2=2.26
r174 3 48 400 $w=1.7e-07 $l=9.14631e-07 $layer=licon1_PDIFF $count=1 $X=1.225
+ $Y=2.055 $X2=1.37 $Y2=2.9
r175 3 22 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=1.225
+ $Y=2.055 $X2=1.37 $Y2=2.2
r176 2 37 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=5.05
+ $Y=0.505 $X2=5.19 $Y2=0.78
r177 1 27 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=1.485
+ $Y=0.285 $X2=1.63 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__MUX4_LP%A_470_57# 1 2 3 4 13 17 19 20 22 24 25 26 28
+ 29 30 32 33 34 37 41 43 51
c163 41 0 5.29209e-20 $X=7.875 $Y=2.2
c164 30 0 1.80147e-19 $X=4.355 $Y=0.35
c165 24 0 2.30208e-19 $X=3.68 $Y=2.165
c166 13 0 2.86043e-19 $X=3.395 $Y=0.35
r167 48 50 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=3.48 $Y=1.21 $X2=3.68
+ $Y2=1.21
r168 43 46 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=2.49 $Y=0.35
+ $X2=2.49 $Y2=0.495
r169 39 51 3.22182 $w=2.92e-07 $l=1.5995e-07 $layer=LI1_cond $X=7.875 $Y=0.9
+ $X2=7.752 $Y2=0.815
r170 39 41 84.8128 $w=1.68e-07 $l=1.3e-06 $layer=LI1_cond $X=7.875 $Y=0.9
+ $X2=7.875 $Y2=2.2
r171 35 51 3.22182 $w=2.92e-07 $l=8.5e-08 $layer=LI1_cond $X=7.752 $Y=0.73
+ $X2=7.752 $Y2=0.815
r172 35 37 7.22012 $w=4.13e-07 $l=2.6e-07 $layer=LI1_cond $X=7.752 $Y=0.73
+ $X2=7.752 $Y2=0.47
r173 33 51 3.35233 $w=1.7e-07 $l=2.07e-07 $layer=LI1_cond $X=7.545 $Y=0.815
+ $X2=7.752 $Y2=0.815
r174 33 34 72.4171 $w=1.68e-07 $l=1.11e-06 $layer=LI1_cond $X=7.545 $Y=0.815
+ $X2=6.435 $Y2=0.815
r175 32 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.35 $Y=0.73
+ $X2=6.435 $Y2=0.815
r176 31 32 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=6.35 $Y=0.435
+ $X2=6.35 $Y2=0.73
r177 29 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.265 $Y=0.35
+ $X2=6.35 $Y2=0.435
r178 29 30 124.61 $w=1.68e-07 $l=1.91e-06 $layer=LI1_cond $X=6.265 $Y=0.35
+ $X2=4.355 $Y2=0.35
r179 27 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.27 $Y=0.435
+ $X2=4.355 $Y2=0.35
r180 27 28 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=4.27 $Y=0.435
+ $X2=4.27 $Y2=1.125
r181 26 50 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=3.765 $Y=1.21
+ $X2=3.68 $Y2=1.21
r182 25 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.185 $Y=1.21
+ $X2=4.27 $Y2=1.125
r183 25 26 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=4.185 $Y=1.21
+ $X2=3.765 $Y2=1.21
r184 23 50 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.68 $Y=1.295
+ $X2=3.68 $Y2=1.21
r185 23 24 56.7594 $w=1.68e-07 $l=8.7e-07 $layer=LI1_cond $X=3.68 $Y=1.295
+ $X2=3.68 $Y2=2.165
r186 22 48 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.48 $Y=1.125
+ $X2=3.48 $Y2=1.21
r187 21 22 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.48 $Y=0.435
+ $X2=3.48 $Y2=1.125
r188 19 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.595 $Y=2.25
+ $X2=3.68 $Y2=2.165
r189 19 20 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=3.595 $Y=2.25
+ $X2=2.935 $Y2=2.25
r190 15 20 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.81 $Y=2.335
+ $X2=2.935 $Y2=2.25
r191 15 17 4.84026 $w=2.48e-07 $l=1.05e-07 $layer=LI1_cond $X=2.81 $Y=2.335
+ $X2=2.81 $Y2=2.44
r192 14 43 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.655 $Y=0.35
+ $X2=2.49 $Y2=0.35
r193 13 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.395 $Y=0.35
+ $X2=3.48 $Y2=0.435
r194 13 14 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=3.395 $Y=0.35
+ $X2=2.655 $Y2=0.35
r195 4 41 600 $w=1.7e-07 $l=2.67395e-07 $layer=licon1_PDIFF $count=1 $X=7.655
+ $Y=2.095 $X2=7.875 $Y2=2.2
r196 3 17 600 $w=1.7e-07 $l=4.72546e-07 $layer=licon1_PDIFF $count=1 $X=2.575
+ $Y=2.055 $X2=2.77 $Y2=2.44
r197 2 37 182 $w=1.7e-07 $l=3.4821e-07 $layer=licon1_NDIFF $count=1 $X=7.46
+ $Y=0.235 $X2=7.71 $Y2=0.47
r198 1 46 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.35
+ $Y=0.285 $X2=2.49 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__MUX4_LP%VGND 1 2 3 4 15 19 23 27 30 31 33 34 35 37
+ 52 58 59 62 65
r114 65 66 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=8.88 $Y=0
+ $X2=8.88 $Y2=0
r115 62 63 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r116 59 66 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=9.84 $Y=0 $X2=8.88
+ $Y2=0
r117 58 59 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.84 $Y=0 $X2=9.84
+ $Y2=0
r118 56 65 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.175 $Y=0 $X2=9.01
+ $Y2=0
r119 56 58 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=9.175 $Y=0 $X2=9.84
+ $Y2=0
r120 55 66 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=6.96 $Y=0
+ $X2=8.88 $Y2=0
r121 54 55 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.96 $Y=0
+ $X2=6.96 $Y2=0
r122 52 65 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.845 $Y=0 $X2=9.01
+ $Y2=0
r123 52 54 122.979 $w=1.68e-07 $l=1.885e-06 $layer=LI1_cond $X=8.845 $Y=0
+ $X2=6.96 $Y2=0
r124 51 55 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6.96
+ $Y2=0
r125 50 51 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r126 47 50 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=4.08 $Y=0 $X2=6.48
+ $Y2=0
r127 47 48 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r128 45 48 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r129 45 63 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=3.6 $Y=0 $X2=1.2
+ $Y2=0
r130 44 45 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r131 42 62 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.235 $Y=0 $X2=1.07
+ $Y2=0
r132 42 44 154.294 $w=1.68e-07 $l=2.365e-06 $layer=LI1_cond $X=1.235 $Y=0
+ $X2=3.6 $Y2=0
r133 40 63 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r134 39 40 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r135 37 62 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.905 $Y=0 $X2=1.07
+ $Y2=0
r136 37 39 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=0.905 $Y=0
+ $X2=0.72 $Y2=0
r137 35 51 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=5.04 $Y=0
+ $X2=6.48 $Y2=0
r138 35 48 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=4.08
+ $Y2=0
r139 33 50 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=6.615 $Y=0
+ $X2=6.48 $Y2=0
r140 33 34 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.615 $Y=0 $X2=6.74
+ $Y2=0
r141 32 54 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=6.865 $Y=0 $X2=6.96
+ $Y2=0
r142 32 34 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.865 $Y=0 $X2=6.74
+ $Y2=0
r143 30 44 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=3.755 $Y=0 $X2=3.6
+ $Y2=0
r144 30 31 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.755 $Y=0 $X2=3.88
+ $Y2=0
r145 29 47 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=4.005 $Y=0 $X2=4.08
+ $Y2=0
r146 29 31 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.005 $Y=0 $X2=3.88
+ $Y2=0
r147 25 65 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.01 $Y=0.085
+ $X2=9.01 $Y2=0
r148 25 27 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=9.01 $Y=0.085
+ $X2=9.01 $Y2=0.445
r149 21 34 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.74 $Y=0.085
+ $X2=6.74 $Y2=0
r150 21 23 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=6.74 $Y=0.085
+ $X2=6.74 $Y2=0.38
r151 17 31 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.88 $Y=0.085
+ $X2=3.88 $Y2=0
r152 17 19 29.0416 $w=2.48e-07 $l=6.3e-07 $layer=LI1_cond $X=3.88 $Y=0.085
+ $X2=3.88 $Y2=0.715
r153 13 62 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.07 $Y=0.085
+ $X2=1.07 $Y2=0
r154 13 15 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.07 $Y=0.085
+ $X2=1.07 $Y2=0.38
r155 4 27 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=8.87
+ $Y=0.235 $X2=9.01 $Y2=0.445
r156 3 23 182 $w=1.7e-07 $l=8.19298e-07 $layer=licon1_NDIFF $count=1 $X=5.95
+ $Y=0.235 $X2=6.7 $Y2=0.38
r157 2 19 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=3.78
+ $Y=0.505 $X2=3.92 $Y2=0.715
r158 1 15 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=0.93
+ $Y=0.235 $X2=1.07 $Y2=0.38
.ends

