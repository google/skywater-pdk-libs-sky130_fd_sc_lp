* File: sky130_fd_sc_lp__o211a_lp.pxi.spice
* Created: Wed Sep  2 10:14:07 2020
* 
x_PM_SKY130_FD_SC_LP__O211A_LP%A1 N_A1_M1010_g N_A1_c_68_n N_A1_M1009_g
+ N_A1_c_69_n A1 A1 N_A1_c_66_n N_A1_c_67_n PM_SKY130_FD_SC_LP__O211A_LP%A1
x_PM_SKY130_FD_SC_LP__O211A_LP%A2 N_A2_M1003_g N_A2_M1002_g A2 A2 N_A2_c_101_n
+ N_A2_c_102_n PM_SKY130_FD_SC_LP__O211A_LP%A2
x_PM_SKY130_FD_SC_LP__O211A_LP%B1 N_B1_M1008_g N_B1_M1007_g B1 B1 N_B1_c_139_n
+ PM_SKY130_FD_SC_LP__O211A_LP%B1
x_PM_SKY130_FD_SC_LP__O211A_LP%C1 N_C1_c_172_n N_C1_M1006_g N_C1_M1005_g
+ N_C1_c_173_n C1 C1 N_C1_c_175_n PM_SKY130_FD_SC_LP__O211A_LP%C1
x_PM_SKY130_FD_SC_LP__O211A_LP%A_232_419# N_A_232_419#_M1006_d
+ N_A_232_419#_M1003_d N_A_232_419#_M1005_d N_A_232_419#_M1000_g
+ N_A_232_419#_c_222_n N_A_232_419#_M1004_g N_A_232_419#_M1001_g
+ N_A_232_419#_c_217_n N_A_232_419#_c_231_n N_A_232_419#_c_218_n
+ N_A_232_419#_c_219_n N_A_232_419#_c_227_n N_A_232_419#_c_224_n
+ N_A_232_419#_c_220_n N_A_232_419#_c_226_n N_A_232_419#_c_221_n
+ PM_SKY130_FD_SC_LP__O211A_LP%A_232_419#
x_PM_SKY130_FD_SC_LP__O211A_LP%VPWR N_VPWR_M1009_s N_VPWR_M1007_d N_VPWR_M1004_s
+ N_VPWR_c_293_n N_VPWR_c_294_n N_VPWR_c_295_n N_VPWR_c_296_n N_VPWR_c_297_n
+ N_VPWR_c_298_n VPWR N_VPWR_c_299_n N_VPWR_c_300_n N_VPWR_c_292_n
+ N_VPWR_c_302_n PM_SKY130_FD_SC_LP__O211A_LP%VPWR
x_PM_SKY130_FD_SC_LP__O211A_LP%X N_X_M1001_d N_X_M1004_d X X X X X X X
+ PM_SKY130_FD_SC_LP__O211A_LP%X
x_PM_SKY130_FD_SC_LP__O211A_LP%A_27_144# N_A_27_144#_M1010_s N_A_27_144#_M1002_d
+ N_A_27_144#_c_359_n N_A_27_144#_c_360_n N_A_27_144#_c_361_n
+ PM_SKY130_FD_SC_LP__O211A_LP%A_27_144#
x_PM_SKY130_FD_SC_LP__O211A_LP%VGND N_VGND_M1010_d N_VGND_M1000_s N_VGND_c_385_n
+ N_VGND_c_386_n VGND N_VGND_c_387_n N_VGND_c_388_n N_VGND_c_389_n
+ N_VGND_c_390_n N_VGND_c_391_n N_VGND_c_392_n PM_SKY130_FD_SC_LP__O211A_LP%VGND
cc_1 VNB N_A1_M1010_g 0.035342f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.93
cc_2 VNB N_A1_c_66_n 0.0260969f $X=-0.19 $Y=-0.245 $X2=0.405 $Y2=1.56
cc_3 VNB N_A1_c_67_n 0.00949665f $X=-0.19 $Y=-0.245 $X2=0.405 $Y2=1.56
cc_4 VNB N_A2_M1002_g 0.0261292f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=2.09
cc_5 VNB N_A2_c_101_n 0.024203f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_6 VNB N_A2_c_102_n 0.00479805f $X=-0.19 $Y=-0.245 $X2=0.405 $Y2=1.56
cc_7 VNB N_B1_M1008_g 0.0378848f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.93
cc_8 VNB B1 0.0107409f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=2.595
cc_9 VNB N_B1_c_139_n 0.0113702f $X=-0.19 $Y=-0.245 $X2=0.405 $Y2=1.56
cc_10 VNB N_C1_c_172_n 0.0188803f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.395
cc_11 VNB N_C1_c_173_n 0.0498817f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=2.595
cc_12 VNB C1 0.0071012f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.95
cc_13 VNB N_C1_c_175_n 0.0358748f $X=-0.19 $Y=-0.245 $X2=0.405 $Y2=1.56
cc_14 VNB N_A_232_419#_M1000_g 0.0215622f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.95
cc_15 VNB N_A_232_419#_M1001_g 0.0205619f $X=-0.19 $Y=-0.245 $X2=0.405 $Y2=1.725
cc_16 VNB N_A_232_419#_c_217_n 0.0371358f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_232_419#_c_218_n 0.0111465f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_232_419#_c_219_n 0.0150063f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_232_419#_c_220_n 0.00684859f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_232_419#_c_221_n 0.0500026f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_VPWR_c_292_n 0.163682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB X 0.0178929f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=2.09
cc_23 VNB X 0.0508844f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=2.595
cc_24 VNB N_A_27_144#_c_359_n 0.0121136f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=2.09
cc_25 VNB N_A_27_144#_c_360_n 0.00399101f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_26 VNB N_A_27_144#_c_361_n 0.0183843f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_385_n 0.039968f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=2.595
cc_28 VNB N_VGND_c_386_n 0.0166594f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_387_n 0.022032f $X=-0.19 $Y=-0.245 $X2=0.405 $Y2=1.56
cc_30 VNB N_VGND_c_388_n 0.0489145f $X=-0.19 $Y=-0.245 $X2=0.342 $Y2=1.665
cc_31 VNB N_VGND_c_389_n 0.027824f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_390_n 0.251397f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_391_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_392_n 0.00510939f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VPB N_A1_c_68_n 0.0299907f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=2.09
cc_36 VPB N_A1_c_69_n 0.0156111f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=1.965
cc_37 VPB N_A1_c_66_n 0.0107608f $X=-0.19 $Y=1.655 $X2=0.405 $Y2=1.56
cc_38 VPB N_A1_c_67_n 0.019881f $X=-0.19 $Y=1.655 $X2=0.405 $Y2=1.56
cc_39 VPB N_A2_M1003_g 0.0352355f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=0.93
cc_40 VPB N_A2_c_101_n 0.00861043f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_41 VPB N_A2_c_102_n 0.00618433f $X=-0.19 $Y=1.655 $X2=0.405 $Y2=1.56
cc_42 VPB N_B1_M1007_g 0.0257803f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=2.09
cc_43 VPB B1 0.00120407f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=2.595
cc_44 VPB N_B1_c_139_n 0.0280218f $X=-0.19 $Y=1.655 $X2=0.405 $Y2=1.56
cc_45 VPB N_C1_M1005_g 0.0496376f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=1.965
cc_46 VPB N_C1_c_173_n 8.70029e-19 $X=-0.19 $Y=1.655 $X2=0.545 $Y2=2.595
cc_47 VPB C1 0.0164292f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.95
cc_48 VPB N_C1_c_175_n 0.0163946f $X=-0.19 $Y=1.655 $X2=0.405 $Y2=1.56
cc_49 VPB N_A_232_419#_c_222_n 0.0356764f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_50 VPB N_A_232_419#_c_217_n 0.0186568f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_51 VPB N_A_232_419#_c_224_n 0.00709126f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_52 VPB N_A_232_419#_c_220_n 0.0101473f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_53 VPB N_A_232_419#_c_226_n 0.00533603f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_54 VPB N_VPWR_c_293_n 0.0109777f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=1.965
cc_55 VPB N_VPWR_c_294_n 0.0325875f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.95
cc_56 VPB N_VPWR_c_295_n 0.00284591f $X=-0.19 $Y=1.655 $X2=0.405 $Y2=1.56
cc_57 VPB N_VPWR_c_296_n 0.0168232f $X=-0.19 $Y=1.655 $X2=0.342 $Y2=1.56
cc_58 VPB N_VPWR_c_297_n 0.0233961f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_59 VPB N_VPWR_c_298_n 0.00548753f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_60 VPB N_VPWR_c_299_n 0.0336396f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_61 VPB N_VPWR_c_300_n 0.0196629f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_62 VPB N_VPWR_c_292_n 0.0593177f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_63 VPB N_VPWR_c_302_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_64 VPB X 0.0605003f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=2.595
cc_65 N_A1_c_68_n N_A2_M1003_g 0.070416f $X=0.545 $Y=2.09 $X2=0 $Y2=0
cc_66 N_A1_c_69_n N_A2_M1003_g 0.00750739f $X=0.545 $Y=1.965 $X2=0 $Y2=0
cc_67 N_A1_c_67_n N_A2_M1003_g 4.03625e-19 $X=0.405 $Y=1.56 $X2=0 $Y2=0
cc_68 N_A1_M1010_g N_A2_M1002_g 0.0183692f $X=0.495 $Y=0.93 $X2=0 $Y2=0
cc_69 N_A1_c_66_n N_A2_c_101_n 0.0209351f $X=0.405 $Y=1.56 $X2=0 $Y2=0
cc_70 N_A1_c_67_n N_A2_c_101_n 0.00101771f $X=0.405 $Y=1.56 $X2=0 $Y2=0
cc_71 N_A1_c_68_n N_A2_c_102_n 0.00135336f $X=0.545 $Y=2.09 $X2=0 $Y2=0
cc_72 N_A1_c_69_n N_A2_c_102_n 0.00167518f $X=0.545 $Y=1.965 $X2=0 $Y2=0
cc_73 N_A1_c_66_n N_A2_c_102_n 9.89635e-19 $X=0.405 $Y=1.56 $X2=0 $Y2=0
cc_74 N_A1_c_67_n N_A2_c_102_n 0.0495665f $X=0.405 $Y=1.56 $X2=0 $Y2=0
cc_75 N_A1_c_68_n N_A_232_419#_c_227_n 0.00325465f $X=0.545 $Y=2.09 $X2=0 $Y2=0
cc_76 N_A1_c_67_n N_VPWR_M1009_s 0.00278687f $X=0.405 $Y=1.56 $X2=-0.19
+ $Y2=-0.245
cc_77 N_A1_c_68_n N_VPWR_c_294_n 0.0235505f $X=0.545 $Y=2.09 $X2=0 $Y2=0
cc_78 N_A1_c_66_n N_VPWR_c_294_n 5.31596e-19 $X=0.405 $Y=1.56 $X2=0 $Y2=0
cc_79 N_A1_c_67_n N_VPWR_c_294_n 0.0243791f $X=0.405 $Y=1.56 $X2=0 $Y2=0
cc_80 N_A1_c_68_n N_VPWR_c_299_n 0.008763f $X=0.545 $Y=2.09 $X2=0 $Y2=0
cc_81 N_A1_c_68_n N_VPWR_c_292_n 0.0144563f $X=0.545 $Y=2.09 $X2=0 $Y2=0
cc_82 N_A1_M1010_g N_A_27_144#_c_359_n 0.0153124f $X=0.495 $Y=0.93 $X2=0 $Y2=0
cc_83 N_A1_c_68_n N_A_27_144#_c_359_n 0.00241987f $X=0.545 $Y=2.09 $X2=0 $Y2=0
cc_84 N_A1_c_66_n N_A_27_144#_c_359_n 0.00129952f $X=0.405 $Y=1.56 $X2=0 $Y2=0
cc_85 N_A1_c_67_n N_A_27_144#_c_359_n 0.0157832f $X=0.405 $Y=1.56 $X2=0 $Y2=0
cc_86 N_A1_M1010_g N_A_27_144#_c_360_n 8.11586e-19 $X=0.495 $Y=0.93 $X2=0 $Y2=0
cc_87 N_A1_M1010_g N_A_27_144#_c_361_n 0.00115543f $X=0.495 $Y=0.93 $X2=0 $Y2=0
cc_88 N_A1_c_66_n N_A_27_144#_c_361_n 0.00300031f $X=0.405 $Y=1.56 $X2=0 $Y2=0
cc_89 N_A1_c_67_n N_A_27_144#_c_361_n 0.0219098f $X=0.405 $Y=1.56 $X2=0 $Y2=0
cc_90 N_A1_M1010_g N_VGND_c_385_n 0.00505645f $X=0.495 $Y=0.93 $X2=0 $Y2=0
cc_91 N_A1_M1010_g N_VGND_c_387_n 0.00368595f $X=0.495 $Y=0.93 $X2=0 $Y2=0
cc_92 N_A1_M1010_g N_VGND_c_390_n 0.00443953f $X=0.495 $Y=0.93 $X2=0 $Y2=0
cc_93 N_A2_M1002_g N_B1_M1008_g 0.0222041f $X=1.085 $Y=0.93 $X2=0 $Y2=0
cc_94 N_A2_c_102_n N_B1_M1008_g 0.0089364f $X=0.945 $Y=1.56 $X2=0 $Y2=0
cc_95 N_A2_M1003_g N_B1_M1007_g 0.0222041f $X=1.035 $Y=2.595 $X2=0 $Y2=0
cc_96 N_A2_c_101_n B1 3.65501e-19 $X=0.945 $Y=1.56 $X2=0 $Y2=0
cc_97 N_A2_c_102_n B1 0.0467848f $X=0.945 $Y=1.56 $X2=0 $Y2=0
cc_98 N_A2_c_101_n N_B1_c_139_n 0.0222041f $X=0.945 $Y=1.56 $X2=0 $Y2=0
cc_99 N_A2_c_102_n N_A_232_419#_M1003_d 0.00192192f $X=0.945 $Y=1.56 $X2=0 $Y2=0
cc_100 N_A2_M1003_g N_A_232_419#_c_227_n 0.0160617f $X=1.035 $Y=2.595 $X2=0
+ $Y2=0
cc_101 N_A2_c_102_n N_A_232_419#_c_227_n 0.0170777f $X=0.945 $Y=1.56 $X2=0 $Y2=0
cc_102 N_A2_M1003_g N_VPWR_c_294_n 0.00429931f $X=1.035 $Y=2.595 $X2=0 $Y2=0
cc_103 N_A2_M1003_g N_VPWR_c_295_n 0.00105123f $X=1.035 $Y=2.595 $X2=0 $Y2=0
cc_104 N_A2_M1003_g N_VPWR_c_299_n 0.00939541f $X=1.035 $Y=2.595 $X2=0 $Y2=0
cc_105 N_A2_M1003_g N_VPWR_c_292_n 0.0161521f $X=1.035 $Y=2.595 $X2=0 $Y2=0
cc_106 N_A2_c_102_n A_134_419# 0.00367761f $X=0.945 $Y=1.56 $X2=-0.19 $Y2=-0.245
cc_107 N_A2_M1002_g N_A_27_144#_c_359_n 0.0137785f $X=1.085 $Y=0.93 $X2=0 $Y2=0
cc_108 N_A2_c_101_n N_A_27_144#_c_359_n 0.00586385f $X=0.945 $Y=1.56 $X2=0 $Y2=0
cc_109 N_A2_c_102_n N_A_27_144#_c_359_n 0.053695f $X=0.945 $Y=1.56 $X2=0 $Y2=0
cc_110 N_A2_M1002_g N_A_27_144#_c_360_n 0.00676736f $X=1.085 $Y=0.93 $X2=0 $Y2=0
cc_111 N_A2_M1002_g N_VGND_c_385_n 0.00468619f $X=1.085 $Y=0.93 $X2=0 $Y2=0
cc_112 N_A2_M1002_g N_VGND_c_388_n 0.00355997f $X=1.085 $Y=0.93 $X2=0 $Y2=0
cc_113 N_A2_M1002_g N_VGND_c_390_n 0.00443953f $X=1.085 $Y=0.93 $X2=0 $Y2=0
cc_114 N_B1_M1008_g N_C1_c_172_n 0.040424f $X=1.515 $Y=0.93 $X2=-0.19 $Y2=-0.245
cc_115 N_B1_M1007_g N_C1_M1005_g 0.0316281f $X=1.565 $Y=2.595 $X2=0 $Y2=0
cc_116 B1 N_C1_M1005_g 0.00174479f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_117 N_B1_M1008_g N_C1_c_173_n 0.00579465f $X=1.515 $Y=0.93 $X2=0 $Y2=0
cc_118 B1 N_C1_c_173_n 0.00287676f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_119 N_B1_c_139_n N_C1_c_173_n 0.0230547f $X=1.705 $Y=1.77 $X2=0 $Y2=0
cc_120 N_B1_M1007_g N_A_232_419#_c_231_n 0.018159f $X=1.565 $Y=2.595 $X2=0 $Y2=0
cc_121 B1 N_A_232_419#_c_231_n 0.0172639f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_122 N_B1_c_139_n N_A_232_419#_c_231_n 6.96397e-19 $X=1.705 $Y=1.77 $X2=0
+ $Y2=0
cc_123 N_B1_M1008_g N_A_232_419#_c_218_n 0.00129863f $X=1.515 $Y=0.93 $X2=0
+ $Y2=0
cc_124 N_B1_M1007_g N_A_232_419#_c_227_n 0.0130701f $X=1.565 $Y=2.595 $X2=0
+ $Y2=0
cc_125 N_B1_M1007_g N_A_232_419#_c_224_n 0.00190124f $X=1.565 $Y=2.595 $X2=0
+ $Y2=0
cc_126 N_B1_M1008_g N_A_232_419#_c_220_n 0.00138421f $X=1.515 $Y=0.93 $X2=0
+ $Y2=0
cc_127 B1 N_A_232_419#_c_220_n 0.027237f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_128 N_B1_c_139_n N_A_232_419#_c_220_n 0.00104894f $X=1.705 $Y=1.77 $X2=0
+ $Y2=0
cc_129 B1 N_VPWR_M1007_d 0.00184052f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_130 N_B1_M1007_g N_VPWR_c_295_n 0.0134447f $X=1.565 $Y=2.595 $X2=0 $Y2=0
cc_131 N_B1_M1007_g N_VPWR_c_299_n 0.00840199f $X=1.565 $Y=2.595 $X2=0 $Y2=0
cc_132 N_B1_M1007_g N_VPWR_c_292_n 0.00763111f $X=1.565 $Y=2.595 $X2=0 $Y2=0
cc_133 N_B1_M1008_g N_A_27_144#_c_359_n 0.00618973f $X=1.515 $Y=0.93 $X2=0 $Y2=0
cc_134 N_B1_M1008_g N_A_27_144#_c_360_n 0.00745101f $X=1.515 $Y=0.93 $X2=0 $Y2=0
cc_135 N_B1_M1008_g N_VGND_c_388_n 0.00355997f $X=1.515 $Y=0.93 $X2=0 $Y2=0
cc_136 N_B1_M1008_g N_VGND_c_390_n 0.00443953f $X=1.515 $Y=0.93 $X2=0 $Y2=0
cc_137 C1 N_A_232_419#_c_222_n 0.00264535f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_138 C1 N_A_232_419#_c_217_n 0.00643806f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_139 N_C1_c_175_n N_A_232_419#_c_217_n 0.00758545f $X=2.69 $Y=1.51 $X2=0 $Y2=0
cc_140 N_C1_M1005_g N_A_232_419#_c_231_n 0.0110863f $X=2.205 $Y=2.595 $X2=0
+ $Y2=0
cc_141 N_C1_c_172_n N_A_232_419#_c_218_n 0.0106441f $X=1.905 $Y=1.215 $X2=0
+ $Y2=0
cc_142 N_C1_c_173_n N_A_232_419#_c_218_n 0.00935161f $X=2.33 $Y=1.51 $X2=0 $Y2=0
cc_143 C1 N_A_232_419#_c_219_n 0.0457814f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_144 N_C1_c_175_n N_A_232_419#_c_219_n 0.0141701f $X=2.69 $Y=1.51 $X2=0 $Y2=0
cc_145 N_C1_M1005_g N_A_232_419#_c_227_n 8.31599e-19 $X=2.205 $Y=2.595 $X2=0
+ $Y2=0
cc_146 N_C1_M1005_g N_A_232_419#_c_224_n 0.0113701f $X=2.205 $Y=2.595 $X2=0
+ $Y2=0
cc_147 C1 N_A_232_419#_c_224_n 0.0066981f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_148 N_C1_c_175_n N_A_232_419#_c_224_n 0.00692787f $X=2.69 $Y=1.51 $X2=0 $Y2=0
cc_149 N_C1_c_172_n N_A_232_419#_c_220_n 0.00179961f $X=1.905 $Y=1.215 $X2=0
+ $Y2=0
cc_150 N_C1_M1005_g N_A_232_419#_c_220_n 0.0154208f $X=2.205 $Y=2.595 $X2=0
+ $Y2=0
cc_151 N_C1_c_173_n N_A_232_419#_c_220_n 0.0191927f $X=2.33 $Y=1.51 $X2=0 $Y2=0
cc_152 C1 N_A_232_419#_c_220_n 0.0324829f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_153 N_C1_c_175_n N_A_232_419#_c_220_n 0.00564651f $X=2.69 $Y=1.51 $X2=0 $Y2=0
cc_154 N_C1_M1005_g N_A_232_419#_c_226_n 0.0205801f $X=2.205 $Y=2.595 $X2=0
+ $Y2=0
cc_155 C1 N_A_232_419#_c_221_n 0.00944757f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_156 N_C1_M1005_g N_VPWR_c_295_n 0.00732786f $X=2.205 $Y=2.595 $X2=0 $Y2=0
cc_157 N_C1_M1005_g N_VPWR_c_296_n 0.00499994f $X=2.205 $Y=2.595 $X2=0 $Y2=0
cc_158 C1 N_VPWR_c_296_n 0.0227986f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_159 N_C1_M1005_g N_VPWR_c_297_n 0.00743996f $X=2.205 $Y=2.595 $X2=0 $Y2=0
cc_160 N_C1_M1005_g N_VPWR_c_292_n 0.0101159f $X=2.205 $Y=2.595 $X2=0 $Y2=0
cc_161 C1 X 0.0295474f $X=3.035 $Y=1.58 $X2=0 $Y2=0
cc_162 N_C1_c_172_n N_A_27_144#_c_360_n 0.00113083f $X=1.905 $Y=1.215 $X2=0
+ $Y2=0
cc_163 N_C1_c_172_n N_VGND_c_386_n 5.96445e-19 $X=1.905 $Y=1.215 $X2=0 $Y2=0
cc_164 N_C1_c_172_n N_VGND_c_388_n 0.00355472f $X=1.905 $Y=1.215 $X2=0 $Y2=0
cc_165 N_C1_c_172_n N_VGND_c_390_n 0.00443953f $X=1.905 $Y=1.215 $X2=0 $Y2=0
cc_166 N_A_232_419#_c_231_n N_VPWR_M1007_d 0.0104996f $X=2.175 $Y=2.395 $X2=0
+ $Y2=0
cc_167 N_A_232_419#_c_231_n N_VPWR_c_295_n 0.0204762f $X=2.175 $Y=2.395 $X2=0
+ $Y2=0
cc_168 N_A_232_419#_c_227_n N_VPWR_c_295_n 0.0266857f $X=1.3 $Y=2.475 $X2=0
+ $Y2=0
cc_169 N_A_232_419#_c_226_n N_VPWR_c_295_n 0.0308377f $X=2.405 $Y=2.395 $X2=0
+ $Y2=0
cc_170 N_A_232_419#_c_222_n N_VPWR_c_296_n 0.0229639f $X=3.295 $Y=2.04 $X2=0
+ $Y2=0
cc_171 N_A_232_419#_c_224_n N_VPWR_c_296_n 0.0684268f $X=2.47 $Y=2.24 $X2=0
+ $Y2=0
cc_172 N_A_232_419#_c_220_n N_VPWR_c_296_n 0.00180986f $X=2.405 $Y=2.075 $X2=0
+ $Y2=0
cc_173 N_A_232_419#_c_226_n N_VPWR_c_297_n 0.028073f $X=2.405 $Y=2.395 $X2=0
+ $Y2=0
cc_174 N_A_232_419#_c_227_n N_VPWR_c_299_n 0.0177952f $X=1.3 $Y=2.475 $X2=0
+ $Y2=0
cc_175 N_A_232_419#_c_222_n N_VPWR_c_300_n 0.00802402f $X=3.295 $Y=2.04 $X2=0
+ $Y2=0
cc_176 N_A_232_419#_M1003_d N_VPWR_c_292_n 0.00223819f $X=1.16 $Y=2.095 $X2=0
+ $Y2=0
cc_177 N_A_232_419#_M1005_d N_VPWR_c_292_n 0.0023218f $X=2.33 $Y=2.095 $X2=0
+ $Y2=0
cc_178 N_A_232_419#_c_222_n N_VPWR_c_292_n 0.0149742f $X=3.295 $Y=2.04 $X2=0
+ $Y2=0
cc_179 N_A_232_419#_c_231_n N_VPWR_c_292_n 0.0120118f $X=2.175 $Y=2.395 $X2=0
+ $Y2=0
cc_180 N_A_232_419#_c_227_n N_VPWR_c_292_n 0.0123247f $X=1.3 $Y=2.475 $X2=0
+ $Y2=0
cc_181 N_A_232_419#_c_226_n N_VPWR_c_292_n 0.0169393f $X=2.405 $Y=2.395 $X2=0
+ $Y2=0
cc_182 N_A_232_419#_M1000_g X 0.0012881f $X=2.955 $Y=0.445 $X2=0 $Y2=0
cc_183 N_A_232_419#_M1001_g X 0.00884521f $X=3.345 $Y=0.445 $X2=0 $Y2=0
cc_184 N_A_232_419#_M1001_g X 0.0451276f $X=3.345 $Y=0.445 $X2=0 $Y2=0
cc_185 N_A_232_419#_c_219_n X 0.0192963f $X=3.045 $Y=0.96 $X2=0 $Y2=0
cc_186 N_A_232_419#_c_218_n N_A_27_144#_c_359_n 0.00208102f $X=2.345 $Y=0.96
+ $X2=0 $Y2=0
cc_187 N_A_232_419#_c_218_n N_A_27_144#_c_360_n 0.0132482f $X=2.345 $Y=0.96
+ $X2=0 $Y2=0
cc_188 N_A_232_419#_M1000_g N_VGND_c_386_n 0.0126731f $X=2.955 $Y=0.445 $X2=0
+ $Y2=0
cc_189 N_A_232_419#_M1001_g N_VGND_c_386_n 0.00222718f $X=3.345 $Y=0.445 $X2=0
+ $Y2=0
cc_190 N_A_232_419#_c_219_n N_VGND_c_386_n 0.0238544f $X=3.045 $Y=0.96 $X2=0
+ $Y2=0
cc_191 N_A_232_419#_c_218_n N_VGND_c_388_n 0.0057001f $X=2.345 $Y=0.96 $X2=0
+ $Y2=0
cc_192 N_A_232_419#_M1000_g N_VGND_c_389_n 0.00486043f $X=2.955 $Y=0.445 $X2=0
+ $Y2=0
cc_193 N_A_232_419#_M1001_g N_VGND_c_389_n 0.00549284f $X=3.345 $Y=0.445 $X2=0
+ $Y2=0
cc_194 N_A_232_419#_M1000_g N_VGND_c_390_n 0.00440794f $X=2.955 $Y=0.445 $X2=0
+ $Y2=0
cc_195 N_A_232_419#_M1001_g N_VGND_c_390_n 0.0109988f $X=3.345 $Y=0.445 $X2=0
+ $Y2=0
cc_196 N_A_232_419#_c_218_n N_VGND_c_390_n 0.011858f $X=2.345 $Y=0.96 $X2=0
+ $Y2=0
cc_197 N_A_232_419#_c_219_n N_VGND_c_390_n 0.0201024f $X=3.045 $Y=0.96 $X2=0
+ $Y2=0
cc_198 N_A_232_419#_c_221_n N_VGND_c_390_n 0.00139702f $X=3.345 $Y=0.96 $X2=0
+ $Y2=0
cc_199 N_VPWR_c_292_n A_134_419# 0.010279f $X=3.6 $Y=3.33 $X2=-0.19 $Y2=-0.245
cc_200 N_VPWR_c_296_n X 0.0272354f $X=3.03 $Y=2.19 $X2=0 $Y2=0
cc_201 N_VPWR_c_300_n X 0.0167213f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_202 N_VPWR_c_292_n X 0.0095959f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_203 X N_VGND_c_386_n 0.0110882f $X=3.515 $Y=0.47 $X2=0 $Y2=0
cc_204 X N_VGND_c_389_n 0.0197343f $X=3.515 $Y=0.47 $X2=0 $Y2=0
cc_205 N_X_M1001_d N_VGND_c_390_n 0.00232985f $X=3.42 $Y=0.235 $X2=0 $Y2=0
cc_206 X N_VGND_c_390_n 0.0125406f $X=3.515 $Y=0.47 $X2=0 $Y2=0
cc_207 N_A_27_144#_c_359_n N_VGND_M1010_d 0.00363814f $X=1.135 $Y=1.185
+ $X2=-0.19 $Y2=-0.245
cc_208 N_A_27_144#_c_359_n N_VGND_c_385_n 0.0265229f $X=1.135 $Y=1.185 $X2=0
+ $Y2=0
cc_209 N_A_27_144#_c_360_n N_VGND_c_385_n 0.00900273f $X=1.3 $Y=0.93 $X2=0 $Y2=0
cc_210 N_A_27_144#_c_360_n N_VGND_c_388_n 0.00563531f $X=1.3 $Y=0.93 $X2=0 $Y2=0
cc_211 N_A_27_144#_c_360_n N_VGND_c_390_n 0.00933109f $X=1.3 $Y=0.93 $X2=0 $Y2=0
cc_212 N_A_27_144#_c_361_n N_VGND_c_390_n 0.00922788f $X=0.28 $Y=1.015 $X2=0
+ $Y2=0
cc_213 N_VGND_c_390_n A_606_47# 0.00508983f $X=3.6 $Y=0 $X2=-0.19 $Y2=-0.245
