# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__dlrtp_2
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__dlrtp_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.200000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.580000 0.315000 0.805000 0.815000 ;
        RECT 0.580000 0.815000 0.880000 2.120000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.684600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.160000 0.345000 6.565000 1.175000 ;
        RECT 6.385000 1.175000 6.565000 3.075000 ;
    END
  END Q
  PIN RESET_B
    ANTENNAGATEAREA  0.315000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.355000 1.210000 5.675000 1.755000 ;
    END
  END RESET_B
  PIN GATE
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 1.050000 0.815000 1.300000 2.120000 ;
    END
  END GATE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 7.200000 0.085000 ;
        RECT 0.975000  0.085000 1.175000 0.645000 ;
        RECT 2.465000  0.085000 2.745000 0.535000 ;
        RECT 4.280000  0.085000 4.480000 0.555000 ;
        RECT 5.605000  0.085000 5.935000 1.040000 ;
        RECT 6.735000  0.085000 6.985000 1.225000 ;
      LAYER mcon ;
        RECT 0.155000 -0.085000 0.325000 0.085000 ;
        RECT 0.635000 -0.085000 0.805000 0.085000 ;
        RECT 1.115000 -0.085000 1.285000 0.085000 ;
        RECT 1.595000 -0.085000 1.765000 0.085000 ;
        RECT 2.075000 -0.085000 2.245000 0.085000 ;
        RECT 2.555000 -0.085000 2.725000 0.085000 ;
        RECT 3.035000 -0.085000 3.205000 0.085000 ;
        RECT 3.515000 -0.085000 3.685000 0.085000 ;
        RECT 3.995000 -0.085000 4.165000 0.085000 ;
        RECT 4.475000 -0.085000 4.645000 0.085000 ;
        RECT 4.955000 -0.085000 5.125000 0.085000 ;
        RECT 5.435000 -0.085000 5.605000 0.085000 ;
        RECT 5.915000 -0.085000 6.085000 0.085000 ;
        RECT 6.395000 -0.085000 6.565000 0.085000 ;
        RECT 6.875000 -0.085000 7.045000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 7.200000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.245000 7.200000 3.415000 ;
        RECT 0.600000 2.695000 0.850000 3.245000 ;
        RECT 2.645000 2.395000 2.835000 3.245000 ;
        RECT 4.290000 2.440000 4.785000 2.630000 ;
        RECT 4.290000 2.630000 5.050000 3.245000 ;
        RECT 5.750000 2.265000 6.080000 3.245000 ;
        RECT 6.735000 1.815000 7.075000 3.245000 ;
      LAYER mcon ;
        RECT 0.155000 3.245000 0.325000 3.415000 ;
        RECT 0.635000 3.245000 0.805000 3.415000 ;
        RECT 1.115000 3.245000 1.285000 3.415000 ;
        RECT 1.595000 3.245000 1.765000 3.415000 ;
        RECT 2.075000 3.245000 2.245000 3.415000 ;
        RECT 2.555000 3.245000 2.725000 3.415000 ;
        RECT 3.035000 3.245000 3.205000 3.415000 ;
        RECT 3.515000 3.245000 3.685000 3.415000 ;
        RECT 3.995000 3.245000 4.165000 3.415000 ;
        RECT 4.475000 3.245000 4.645000 3.415000 ;
        RECT 4.955000 3.245000 5.125000 3.415000 ;
        RECT 5.435000 3.245000 5.605000 3.415000 ;
        RECT 5.915000 3.245000 6.085000 3.415000 ;
        RECT 6.395000 3.245000 6.565000 3.415000 ;
        RECT 6.875000 3.245000 7.045000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 7.200000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.160000 0.315000 0.410000 2.355000 ;
      RECT 0.160000 2.355000 1.190000 2.525000 ;
      RECT 0.160000 2.525000 0.430000 3.025000 ;
      RECT 1.020000 2.525000 1.190000 2.885000 ;
      RECT 1.020000 2.885000 2.475000 3.055000 ;
      RECT 1.360000 2.355000 1.715000 2.715000 ;
      RECT 1.425000 0.330000 1.650000 0.660000 ;
      RECT 1.480000 0.660000 1.650000 1.885000 ;
      RECT 1.480000 1.885000 1.715000 2.355000 ;
      RECT 1.820000 0.255000 2.295000 0.535000 ;
      RECT 1.820000 0.535000 2.010000 1.535000 ;
      RECT 1.820000 1.535000 3.175000 1.705000 ;
      RECT 1.885000 1.705000 2.135000 2.715000 ;
      RECT 2.180000 0.705000 3.760000 0.875000 ;
      RECT 2.180000 0.875000 2.510000 1.365000 ;
      RECT 2.305000 1.895000 2.835000 2.225000 ;
      RECT 2.305000 2.225000 2.475000 2.885000 ;
      RECT 3.005000 1.045000 3.410000 1.305000 ;
      RECT 3.005000 1.305000 3.175000 1.535000 ;
      RECT 3.005000 1.705000 3.175000 2.825000 ;
      RECT 3.005000 2.825000 4.070000 2.995000 ;
      RECT 3.315000 0.255000 4.110000 0.535000 ;
      RECT 3.355000 1.555000 4.775000 1.725000 ;
      RECT 3.355000 1.725000 3.525000 2.405000 ;
      RECT 3.355000 2.405000 3.720000 2.655000 ;
      RECT 3.590000 0.875000 3.760000 1.125000 ;
      RECT 3.590000 1.125000 3.950000 1.385000 ;
      RECT 3.705000 1.905000 4.070000 2.235000 ;
      RECT 3.900000 2.235000 4.070000 2.825000 ;
      RECT 3.940000 0.535000 4.110000 0.725000 ;
      RECT 3.940000 0.725000 4.640000 0.895000 ;
      RECT 4.240000 1.905000 5.125000 1.925000 ;
      RECT 4.240000 1.925000 6.215000 2.095000 ;
      RECT 4.240000 2.095000 5.470000 2.235000 ;
      RECT 4.470000 0.895000 4.640000 1.335000 ;
      RECT 4.470000 1.335000 4.775000 1.555000 ;
      RECT 4.810000 0.345000 5.125000 1.165000 ;
      RECT 4.955000 1.165000 5.125000 1.905000 ;
      RECT 4.955000 2.235000 5.470000 2.460000 ;
      RECT 5.220000 2.460000 5.470000 3.075000 ;
      RECT 5.965000 1.345000 6.215000 1.925000 ;
  END
END sky130_fd_sc_lp__dlrtp_2
