# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__mux2i_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_lp__mux2i_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.840000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A0
    ANTENNAGATEAREA  0.315000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.345000 0.470000 1.760000 ;
    END
  END A0
  PIN A1
    ANTENNAGATEAREA  0.315000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.980000 1.425000 1.310000 1.750000 ;
    END
  END A1
  PIN S
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.375000 1.210000 3.755000 1.750000 ;
    END
  END S
  PIN Y
    ANTENNADIFFAREA  0.693000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.555000 0.595000 0.885000 1.165000 ;
        RECT 0.555000 1.165000 0.810000 1.175000 ;
        RECT 0.640000 1.175000 0.810000 1.930000 ;
        RECT 0.640000 1.930000 1.285000 2.140000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.840000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.840000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.840000 0.085000 ;
      RECT 0.000000  3.245000 3.840000 3.415000 ;
      RECT 0.105000  0.255000 1.915000 0.425000 ;
      RECT 0.105000  0.425000 0.385000 1.175000 ;
      RECT 0.200000  1.930000 0.470000 2.310000 ;
      RECT 0.200000  2.310000 1.625000 2.550000 ;
      RECT 0.200000  2.550000 0.530000 3.075000 ;
      RECT 1.055000  0.595000 1.385000 1.075000 ;
      RECT 1.055000  1.075000 2.775000 1.245000 ;
      RECT 1.455000  1.840000 2.595000 1.985000 ;
      RECT 1.455000  1.985000 1.625000 2.310000 ;
      RECT 1.470000  1.815000 2.595000 1.840000 ;
      RECT 1.520000  1.415000 3.205000 1.585000 ;
      RECT 1.585000  0.425000 1.915000 0.905000 ;
      RECT 1.795000  2.155000 2.125000 3.245000 ;
      RECT 2.085000  0.085000 2.305000 0.905000 ;
      RECT 2.295000  1.985000 2.595000 3.075000 ;
      RECT 2.490000  0.255000 2.775000 1.075000 ;
      RECT 2.945000  1.585000 3.205000 3.075000 ;
      RECT 2.985000  0.360000 3.245000 1.095000 ;
      RECT 2.985000  1.095000 3.205000 1.415000 ;
      RECT 3.375000  1.920000 3.705000 3.245000 ;
      RECT 3.415000  0.085000 3.745000 1.040000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
  END
END sky130_fd_sc_lp__mux2i_1
END LIBRARY
