* File: sky130_fd_sc_lp__buflp_0.spice
* Created: Wed Sep  2 09:36:21 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__buflp_0.pex.spice"
.subckt sky130_fd_sc_lp__buflp_0  VNB VPB A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* VPB	VPB
* VNB	VNB
MM1007 A_123_120# N_A_M1007_g N_A_36_120#_M1007_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.1197 PD=0.66 PS=1.41 NRD=18.564 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1003 N_VGND_M1003_d N_A_M1003_g A_123_120# VNB NSHORT L=0.15 W=0.42 AD=0.0588
+ AS=0.0504 PD=0.7 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75000.6 SB=75001
+ A=0.063 P=1.14 MULT=1
MM1002 A_287_120# N_A_36_120#_M1002_g N_VGND_M1003_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.0588 PD=0.66 PS=0.7 NRD=18.564 NRS=0 M=1 R=2.8 SA=75001
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1005 N_X_M1005_d N_A_36_120#_M1005_g A_287_120# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0504 PD=1.41 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75001.4
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1006 A_128_490# N_A_M1006_g N_A_36_120#_M1006_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0504 AS=0.1197 PD=0.66 PS=1.41 NRD=30.4759 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.5 A=0.063 P=1.14 MULT=1
MM1000 N_VPWR_M1000_d N_A_M1000_g A_128_490# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0905774 AS=0.0504 PD=0.820189 PS=0.66 NRD=55.1009 NRS=30.4759 M=1 R=2.8
+ SA=75000.6 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1004 A_315_446# N_A_36_120#_M1004_g N_VPWR_M1000_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0768 AS=0.138023 PD=0.88 PS=1.24981 NRD=19.9955 NRS=0 M=1 R=4.26667
+ SA=75000.8 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1001 N_X_M1001_d N_A_36_120#_M1001_g A_315_446# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1824 AS=0.0768 PD=1.85 PS=0.88 NRD=0 NRS=19.9955 M=1 R=4.26667 SA=75001.2
+ SB=75000.2 A=0.096 P=1.58 MULT=1
DX8_noxref VNB VPB NWDIODE A=5.1847 P=9.29
*
.include "sky130_fd_sc_lp__buflp_0.pxi.spice"
*
.ends
*
*
