# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__sdfxbp_1
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__sdfxbp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  14.40000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.020000 1.345000 1.520000 2.120000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.556500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.990000 0.375000 13.285000 1.345000 ;
        RECT 12.990000 1.345000 13.405000 2.145000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.615300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 13.845000 0.375000 14.315000 1.175000 ;
        RECT 14.045000 1.175000 14.315000 3.075000 ;
    END
  END Q_N
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.140000 0.550000 2.120000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.975000 0.265000 3.215000 1.390000 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 7.825000 1.120000 8.520000 1.455000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 14.400000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 14.400000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 14.400000 0.085000 ;
      RECT  0.000000  3.245000 14.400000 3.415000 ;
      RECT  0.095000  2.290000  2.075000 2.460000 ;
      RECT  0.095000  2.460000  0.355000 3.065000 ;
      RECT  0.165000  0.085000  0.495000 0.970000 ;
      RECT  0.525000  2.630000  0.855000 3.245000 ;
      RECT  1.010000  0.640000  1.340000 1.005000 ;
      RECT  1.010000  1.005000  1.870000 1.175000 ;
      RECT  1.315000  2.835000  2.425000 2.895000 ;
      RECT  1.315000  2.895000  3.145000 3.065000 ;
      RECT  1.700000  1.175000  1.870000 1.205000 ;
      RECT  1.700000  1.205000  2.425000 1.415000 ;
      RECT  1.745000  2.460000  2.075000 2.665000 ;
      RECT  1.855000  0.085000  2.185000 0.835000 ;
      RECT  2.255000  1.415000  2.425000 2.835000 ;
      RECT  2.355000  0.640000  2.805000 0.970000 ;
      RECT  2.595000  0.970000  2.805000 2.725000 ;
      RECT  2.975000  1.560000  3.555000 1.730000 ;
      RECT  2.975000  1.730000  3.145000 2.385000 ;
      RECT  2.975000  2.385000  5.875000 2.555000 ;
      RECT  2.975000  2.555000  3.145000 2.895000 ;
      RECT  3.315000  2.725000  3.575000 3.245000 ;
      RECT  3.385000  0.265000  4.405000 0.435000 ;
      RECT  3.385000  0.435000  3.555000 1.560000 ;
      RECT  3.795000  0.615000  4.065000 1.685000 ;
      RECT  3.795000  1.685000  6.735000 1.855000 ;
      RECT  3.795000  1.855000  5.050000 2.215000 ;
      RECT  4.235000  0.435000  4.405000 1.335000 ;
      RECT  4.235000  1.335000  6.200000 1.505000 ;
      RECT  4.320000  2.725000  4.650000 3.245000 ;
      RECT  4.575000  0.085000  4.905000 1.165000 ;
      RECT  4.940000  2.725000  5.270000 2.895000 ;
      RECT  4.940000  2.895000  6.895000 3.065000 ;
      RECT  5.390000  2.025000  6.385000 2.215000 ;
      RECT  5.500000  0.255000  6.710000 0.435000 ;
      RECT  5.500000  0.435000  5.795000 0.980000 ;
      RECT  5.545000  2.555000  5.875000 2.725000 ;
      RECT  5.965000  0.650000  6.200000 1.335000 ;
      RECT  6.055000  2.215000  6.385000 2.725000 ;
      RECT  6.380000  0.435000  6.710000 0.855000 ;
      RECT  6.565000  1.855000  6.735000 2.345000 ;
      RECT  6.565000  2.345000 10.240000 2.515000 ;
      RECT  6.565000  2.685000  6.895000 2.895000 ;
      RECT  6.905000  0.615000  7.635000 0.945000 ;
      RECT  6.905000  0.945000  7.165000 1.975000 ;
      RECT  6.905000  1.975000  7.635000 2.165000 ;
      RECT  6.950000  0.255000  7.280000 0.615000 ;
      RECT  7.405000  1.125000  7.655000 1.625000 ;
      RECT  7.405000  1.625000  8.915000 1.795000 ;
      RECT  7.805000  0.085000  8.080000 0.950000 ;
      RECT  7.830000  2.685000  8.160000 3.245000 ;
      RECT  8.250000  0.615000  8.915000 0.945000 ;
      RECT  8.320000  1.795000  8.915000 2.175000 ;
      RECT  8.690000  0.945000  8.915000 1.625000 ;
      RECT  8.910000  2.685000  9.240000 2.725000 ;
      RECT  8.910000  2.725000 10.810000 2.945000 ;
      RECT  9.085000  0.670000  9.575000 1.000000 ;
      RECT  9.085000  1.000000  9.255000 2.345000 ;
      RECT  9.530000  1.445000 11.335000 1.615000 ;
      RECT  9.530000  1.615000  9.860000 2.175000 ;
      RECT  9.745000  0.795000 10.075000 1.445000 ;
      RECT 10.020000  2.515000 10.240000 2.555000 ;
      RECT 10.030000  1.875000 10.240000 2.345000 ;
      RECT 10.410000  1.785000 10.740000 1.805000 ;
      RECT 10.410000  1.805000 11.785000 1.975000 ;
      RECT 10.480000  2.245000 10.810000 2.725000 ;
      RECT 10.680000  0.085000 11.010000 1.215000 ;
      RECT 10.980000  2.145000 11.335000 3.245000 ;
      RECT 11.005000  1.615000 11.335000 1.635000 ;
      RECT 11.180000  0.595000 11.685000 0.975000 ;
      RECT 11.180000  0.975000 12.460000 1.265000 ;
      RECT 11.505000  1.265000 12.460000 1.645000 ;
      RECT 11.505000  1.645000 11.785000 1.805000 ;
      RECT 11.505000  1.975000 11.785000 2.755000 ;
      RECT 11.980000  0.085000 12.270000 0.805000 ;
      RECT 12.005000  1.815000 12.810000 2.325000 ;
      RECT 12.005000  2.325000 13.875000 2.495000 ;
      RECT 12.440000  0.475000 12.810000 0.805000 ;
      RECT 12.530000  2.665000 12.860000 3.245000 ;
      RECT 12.640000  0.805000 12.810000 1.815000 ;
      RECT 13.455000  0.085000 13.675000 1.175000 ;
      RECT 13.545000  2.665000 13.875000 3.245000 ;
      RECT 13.625000  1.345000 13.875000 2.325000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.245000 10.885000 3.415000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  3.245000 11.365000 3.415000 ;
      RECT 11.675000 -0.085000 11.845000 0.085000 ;
      RECT 11.675000  3.245000 11.845000 3.415000 ;
      RECT 12.155000 -0.085000 12.325000 0.085000 ;
      RECT 12.155000  3.245000 12.325000 3.415000 ;
      RECT 12.635000 -0.085000 12.805000 0.085000 ;
      RECT 12.635000  3.245000 12.805000 3.415000 ;
      RECT 13.115000 -0.085000 13.285000 0.085000 ;
      RECT 13.115000  3.245000 13.285000 3.415000 ;
      RECT 13.595000 -0.085000 13.765000 0.085000 ;
      RECT 13.595000  3.245000 13.765000 3.415000 ;
      RECT 14.075000 -0.085000 14.245000 0.085000 ;
      RECT 14.075000  3.245000 14.245000 3.415000 ;
  END
END sky130_fd_sc_lp__sdfxbp_1
END LIBRARY
