* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__o2bb2a_0 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
X0 VPWR A1_N a_229_483# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X1 a_229_483# A2_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X2 X a_80_176# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 a_224_70# A2_N a_229_483# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 a_80_176# B2 a_598_483# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X5 VPWR a_229_483# a_80_176# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X6 a_80_176# a_229_483# a_512_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 X a_80_176# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X8 VGND A1_N a_224_70# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 a_598_483# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X10 a_512_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X11 VGND B1 a_512_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
