* File: sky130_fd_sc_lp__a31o_lp.pex.spice
* Created: Wed Sep  2 09:26:37 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A31O_LP%B1 1 3 5 8 12 14 15 18
r39 18 20 32.0725 $w=3.45e-07 $l=1.65e-07 $layer=POLY_cond $X=0.602 $Y=1.33
+ $X2=0.602 $Y2=1.495
r40 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.61
+ $Y=1.33 $X2=0.61 $Y2=1.33
r41 15 19 3.84148 $w=3.28e-07 $l=1.1e-07 $layer=LI1_cond $X=0.72 $Y=1.33
+ $X2=0.61 $Y2=1.33
r42 8 20 260.876 $w=2.5e-07 $l=1.05e-06 $layer=POLY_cond $X=0.65 $Y=2.545
+ $X2=0.65 $Y2=1.495
r43 5 18 1.17081 $w=3.45e-07 $l=7e-09 $layer=POLY_cond $X=0.602 $Y=1.323
+ $X2=0.602 $Y2=1.33
r44 5 14 66.5689 $w=3.45e-07 $l=3.98e-07 $layer=POLY_cond $X=0.602 $Y=1.323
+ $X2=0.602 $Y2=0.925
r45 1 14 26.2249 $w=3.45e-07 $l=1.5e-07 $layer=POLY_cond $X=0.685 $Y=0.775
+ $X2=0.685 $Y2=0.925
r46 1 12 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.865 $Y=0.775
+ $X2=0.865 $Y2=0.49
r47 1 3 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.505 $Y=0.775
+ $X2=0.505 $Y2=0.49
.ends

.subckt PM_SKY130_FD_SC_LP__A31O_LP%A1 3 9 10 11 12 15 17
c43 11 0 1.17441e-19 $X=1.267 $Y=0.925
r44 15 18 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.15 $Y=1.33
+ $X2=1.15 $Y2=1.495
r45 15 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.15 $Y=1.33
+ $X2=1.15 $Y2=1.165
r46 12 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.15
+ $Y=1.33 $X2=1.15 $Y2=1.33
r47 11 17 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=1.24 $Y=0.925
+ $X2=1.24 $Y2=1.165
r48 10 11 48.5235 $w=2.05e-07 $l=1.5e-07 $layer=POLY_cond $X=1.267 $Y=0.775
+ $X2=1.267 $Y2=0.925
r49 9 10 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=1.295 $Y=0.49
+ $X2=1.295 $Y2=0.775
r50 3 18 260.876 $w=2.5e-07 $l=1.05e-06 $layer=POLY_cond $X=1.18 $Y=2.545
+ $X2=1.18 $Y2=1.495
.ends

.subckt PM_SKY130_FD_SC_LP__A31O_LP%A2 3 7 9 10 11 16
c45 7 0 1.63368e-19 $X=1.685 $Y=0.49
r46 16 19 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.69 $Y=1.33
+ $X2=1.69 $Y2=1.495
r47 16 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.69 $Y=1.33
+ $X2=1.69 $Y2=1.165
r48 11 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.69
+ $Y=1.33 $X2=1.69 $Y2=1.33
r49 10 11 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.69 $Y=0.925
+ $X2=1.69 $Y2=1.295
r50 9 10 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.69 $Y=0.555
+ $X2=1.69 $Y2=0.925
r51 7 18 346.117 $w=1.5e-07 $l=6.75e-07 $layer=POLY_cond $X=1.685 $Y=0.49
+ $X2=1.685 $Y2=1.165
r52 3 19 260.876 $w=2.5e-07 $l=1.05e-06 $layer=POLY_cond $X=1.71 $Y=2.545
+ $X2=1.71 $Y2=1.495
.ends

.subckt PM_SKY130_FD_SC_LP__A31O_LP%A3 3 8 10 11 12 15 17
c43 12 0 4.91139e-20 $X=2.16 $Y=1.295
r44 15 18 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.23 $Y=1.33
+ $X2=2.23 $Y2=1.495
r45 15 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.23 $Y=1.33
+ $X2=2.23 $Y2=1.165
r46 12 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.23
+ $Y=1.33 $X2=2.23 $Y2=1.33
r47 11 17 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=2.14 $Y=0.925
+ $X2=2.14 $Y2=1.165
r48 10 11 44.7709 $w=2.15e-07 $l=1.5e-07 $layer=POLY_cond $X=2.107 $Y=0.775
+ $X2=2.107 $Y2=0.925
r49 8 18 260.876 $w=2.5e-07 $l=1.05e-06 $layer=POLY_cond $X=2.24 $Y=2.545
+ $X2=2.24 $Y2=1.495
r50 3 10 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.075 $Y=0.49
+ $X2=2.075 $Y2=0.775
.ends

.subckt PM_SKY130_FD_SC_LP__A31O_LP%A_48_409# 1 2 7 9 10 11 12 14 18 20 22 23 24
+ 26 29 33 34 35 39 43 44 46
c103 33 0 1.63368e-19 $X=0.915 $Y=0.9
c104 22 0 4.91139e-20 $X=2.77 $Y=1.175
c105 14 0 4.93603e-20 $X=2.77 $Y=2.545
r106 43 44 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.77
+ $Y=1.34 $X2=2.77 $Y2=1.34
r107 41 43 12.2561 $w=3.13e-07 $l=3.35e-07 $layer=LI1_cond $X=2.762 $Y=1.675
+ $X2=2.762 $Y2=1.34
r108 37 39 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=1.08 $Y=0.815
+ $X2=1.08 $Y2=0.49
r109 36 46 3.60271 $w=1.7e-07 $l=2.28e-07 $layer=LI1_cond $X=0.55 $Y=1.76
+ $X2=0.322 $Y2=1.76
r110 35 41 7.64049 $w=1.7e-07 $l=1.94921e-07 $layer=LI1_cond $X=2.605 $Y=1.76
+ $X2=2.762 $Y2=1.675
r111 35 36 134.07 $w=1.68e-07 $l=2.055e-06 $layer=LI1_cond $X=2.605 $Y=1.76
+ $X2=0.55 $Y2=1.76
r112 33 37 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.915 $Y=0.9
+ $X2=1.08 $Y2=0.815
r113 33 34 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=0.915 $Y=0.9
+ $X2=0.265 $Y2=0.9
r114 29 31 18.6641 $w=4.53e-07 $l=7.1e-07 $layer=LI1_cond $X=0.322 $Y=2.19
+ $X2=0.322 $Y2=2.9
r115 27 46 3.03453 $w=3.12e-07 $l=8.5e-08 $layer=LI1_cond $X=0.322 $Y=1.845
+ $X2=0.322 $Y2=1.76
r116 27 29 9.06917 $w=4.53e-07 $l=3.45e-07 $layer=LI1_cond $X=0.322 $Y=1.845
+ $X2=0.322 $Y2=2.19
r117 26 46 3.03453 $w=3.12e-07 $l=1.79538e-07 $layer=LI1_cond $X=0.18 $Y=1.675
+ $X2=0.322 $Y2=1.76
r118 25 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.18 $Y=0.985
+ $X2=0.265 $Y2=0.9
r119 25 26 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=0.18 $Y=0.985
+ $X2=0.18 $Y2=1.675
r120 23 44 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.77 $Y=1.68
+ $X2=2.77 $Y2=1.34
r121 22 44 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.77 $Y=1.175
+ $X2=2.77 $Y2=1.34
r122 18 24 20.4101 $w=1.5e-07 $l=7.64853e-08 $layer=POLY_cond $X=2.865 $Y=0.775
+ $X2=2.862 $Y2=0.85
r123 18 20 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.865 $Y=0.775
+ $X2=2.865 $Y2=0.49
r124 16 24 20.4101 $w=1.5e-07 $l=7.59934e-08 $layer=POLY_cond $X=2.86 $Y=0.925
+ $X2=2.862 $Y2=0.85
r125 16 22 128.191 $w=1.5e-07 $l=2.5e-07 $layer=POLY_cond $X=2.86 $Y=0.925
+ $X2=2.86 $Y2=1.175
r126 12 23 30.6163 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.77 $Y=1.845
+ $X2=2.77 $Y2=1.68
r127 12 14 173.918 $w=2.5e-07 $l=7e-07 $layer=POLY_cond $X=2.77 $Y=1.845
+ $X2=2.77 $Y2=2.545
r128 10 24 5.30422 $w=1.5e-07 $l=7.7e-08 $layer=POLY_cond $X=2.785 $Y=0.85
+ $X2=2.862 $Y2=0.85
r129 10 11 105.117 $w=1.5e-07 $l=2.05e-07 $layer=POLY_cond $X=2.785 $Y=0.85
+ $X2=2.58 $Y2=0.85
r130 7 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.505 $Y=0.775
+ $X2=2.58 $Y2=0.85
r131 7 9 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.505 $Y=0.775
+ $X2=2.505 $Y2=0.49
r132 2 31 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.24
+ $Y=2.045 $X2=0.385 $Y2=2.9
r133 2 29 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.24
+ $Y=2.045 $X2=0.385 $Y2=2.19
r134 1 39 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.94
+ $Y=0.28 $X2=1.08 $Y2=0.49
.ends

.subckt PM_SKY130_FD_SC_LP__A31O_LP%A_155_409# 1 2 7 9 11 13 15
c33 13 0 4.93603e-20 $X=1.975 $Y=2.195
r34 13 20 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.975 $Y=2.195
+ $X2=1.975 $Y2=2.11
r35 13 15 24.6204 $w=3.28e-07 $l=7.05e-07 $layer=LI1_cond $X=1.975 $Y=2.195
+ $X2=1.975 $Y2=2.9
r36 12 18 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.08 $Y=2.11
+ $X2=0.915 $Y2=2.11
r37 11 20 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.81 $Y=2.11
+ $X2=1.975 $Y2=2.11
r38 11 12 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=1.81 $Y=2.11
+ $X2=1.08 $Y2=2.11
r39 7 18 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.915 $Y=2.195
+ $X2=0.915 $Y2=2.11
r40 7 9 24.6204 $w=3.28e-07 $l=7.05e-07 $layer=LI1_cond $X=0.915 $Y=2.195
+ $X2=0.915 $Y2=2.9
r41 2 20 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.835
+ $Y=2.045 $X2=1.975 $Y2=2.19
r42 2 15 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=1.835
+ $Y=2.045 $X2=1.975 $Y2=2.9
r43 1 18 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.775
+ $Y=2.045 $X2=0.915 $Y2=2.19
r44 1 9 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=0.775
+ $Y=2.045 $X2=0.915 $Y2=2.9
.ends

.subckt PM_SKY130_FD_SC_LP__A31O_LP%VPWR 1 2 9 13 18 19 21 22 23 36 37
r43 36 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r44 34 37 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r45 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r46 30 31 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r47 27 31 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.2 $Y2=3.33
r48 26 30 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.24 $Y=3.33 $X2=1.2
+ $Y2=3.33
r49 26 27 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r50 23 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r51 23 31 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r52 21 33 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=2.34 $Y=3.33
+ $X2=2.16 $Y2=3.33
r53 21 22 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.34 $Y=3.33
+ $X2=2.505 $Y2=3.33
r54 20 36 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=2.67 $Y=3.33
+ $X2=3.12 $Y2=3.33
r55 20 22 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.67 $Y=3.33
+ $X2=2.505 $Y2=3.33
r56 18 30 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=1.28 $Y=3.33 $X2=1.2
+ $Y2=3.33
r57 18 19 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.28 $Y=3.33
+ $X2=1.445 $Y2=3.33
r58 17 33 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=1.61 $Y=3.33
+ $X2=2.16 $Y2=3.33
r59 17 19 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.61 $Y=3.33
+ $X2=1.445 $Y2=3.33
r60 13 16 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=2.505 $Y=2.19
+ $X2=2.505 $Y2=2.9
r61 11 22 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.505 $Y=3.245
+ $X2=2.505 $Y2=3.33
r62 11 16 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=2.505 $Y=3.245
+ $X2=2.505 $Y2=2.9
r63 7 19 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.445 $Y=3.245
+ $X2=1.445 $Y2=3.33
r64 7 9 24.6204 $w=3.28e-07 $l=7.05e-07 $layer=LI1_cond $X=1.445 $Y=3.245
+ $X2=1.445 $Y2=2.54
r65 2 16 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=2.365
+ $Y=2.045 $X2=2.505 $Y2=2.9
r66 2 13 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.365
+ $Y=2.045 $X2=2.505 $Y2=2.19
r67 1 9 300 $w=1.7e-07 $l=5.60647e-07 $layer=licon1_PDIFF $count=2 $X=1.305
+ $Y=2.045 $X2=1.445 $Y2=2.54
.ends

.subckt PM_SKY130_FD_SC_LP__A31O_LP%X 1 2 11 12 14 17 18
r23 18 26 3.60138 $w=3.98e-07 $l=1.25e-07 $layer=LI1_cond $X=3.07 $Y=2.775
+ $X2=3.07 $Y2=2.9
r24 17 18 10.6601 $w=3.98e-07 $l=3.7e-07 $layer=LI1_cond $X=3.07 $Y=2.405
+ $X2=3.07 $Y2=2.775
r25 14 16 10.6092 $w=3.53e-07 $l=2.3e-07 $layer=LI1_cond $X=3.092 $Y=0.49
+ $X2=3.092 $Y2=0.72
r26 12 16 85.139 $w=1.68e-07 $l=1.305e-06 $layer=LI1_cond $X=3.185 $Y=2.025
+ $X2=3.185 $Y2=0.72
r27 11 12 8.64761 $w=3.98e-07 $l=1.65e-07 $layer=LI1_cond $X=3.07 $Y=2.19
+ $X2=3.07 $Y2=2.025
r28 9 17 5.18599 $w=3.98e-07 $l=1.8e-07 $layer=LI1_cond $X=3.07 $Y=2.225
+ $X2=3.07 $Y2=2.405
r29 9 11 1.00839 $w=3.98e-07 $l=3.5e-08 $layer=LI1_cond $X=3.07 $Y=2.225
+ $X2=3.07 $Y2=2.19
r30 2 26 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=2.895
+ $Y=2.045 $X2=3.035 $Y2=2.9
r31 2 11 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.895
+ $Y=2.045 $X2=3.035 $Y2=2.19
r32 1 14 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.94
+ $Y=0.28 $X2=3.08 $Y2=0.49
.ends

.subckt PM_SKY130_FD_SC_LP__A31O_LP%VGND 1 2 7 9 13 15 17 24 25 31
c44 17 0 1.17441e-19 $X=2.125 $Y=0
r45 31 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r46 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r47 25 32 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.16
+ $Y2=0
r48 24 25 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r49 22 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.455 $Y=0 $X2=2.29
+ $Y2=0
r50 22 24 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=2.455 $Y=0 $X2=3.12
+ $Y2=0
r51 21 29 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r52 20 21 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r53 18 28 4.70928 $w=1.7e-07 $l=2.28e-07 $layer=LI1_cond $X=0.455 $Y=0 $X2=0.227
+ $Y2=0
r54 18 20 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.455 $Y=0 $X2=0.72
+ $Y2=0
r55 17 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.125 $Y=0 $X2=2.29
+ $Y2=0
r56 17 20 91.6631 $w=1.68e-07 $l=1.405e-06 $layer=LI1_cond $X=2.125 $Y=0
+ $X2=0.72 $Y2=0
r57 15 32 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r58 15 21 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=0.72
+ $Y2=0
r59 11 31 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.29 $Y=0.085
+ $X2=2.29 $Y2=0
r60 11 13 14.1436 $w=3.28e-07 $l=4.05e-07 $layer=LI1_cond $X=2.29 $Y=0.085
+ $X2=2.29 $Y2=0.49
r61 7 28 3.0569 $w=3.3e-07 $l=1.12161e-07 $layer=LI1_cond $X=0.29 $Y=0.085
+ $X2=0.227 $Y2=0
r62 7 9 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=0.29 $Y=0.085 $X2=0.29
+ $Y2=0.445
r63 2 13 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.15
+ $Y=0.28 $X2=2.29 $Y2=0.49
r64 1 9 182 $w=1.7e-07 $l=2.26164e-07 $layer=licon1_NDIFF $count=1 $X=0.145
+ $Y=0.28 $X2=0.29 $Y2=0.445
.ends

