* File: sky130_fd_sc_lp__buf_2.pex.spice
* Created: Fri Aug 28 10:10:18 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__BUF_2%A_90_21# 1 2 9 11 13 14 18 21 22 25 26 28 29
+ 32 36 38 40 42
r64 34 38 3.58051 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=2.085 $Y=1.855
+ $X2=2.085 $Y2=1.77
r65 34 36 5.54059 $w=2.58e-07 $l=1.25e-07 $layer=LI1_cond $X=2.085 $Y=1.855
+ $X2=2.085 $Y2=1.98
r66 30 38 3.58051 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=2.085 $Y=1.685
+ $X2=2.085 $Y2=1.77
r67 30 32 36.3463 $w=2.58e-07 $l=8.2e-07 $layer=LI1_cond $X=2.085 $Y=1.685
+ $X2=2.085 $Y2=0.865
r68 28 38 2.90867 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.955 $Y=1.77
+ $X2=2.085 $Y2=1.77
r69 28 29 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.955 $Y=1.77
+ $X2=1.275 $Y2=1.77
r70 26 40 68.0917 $w=3.95e-07 $l=3.25e-07 $layer=POLY_cond $X=1.077 $Y=1.51
+ $X2=1.077 $Y2=1.185
r71 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.11
+ $Y=1.51 $X2=1.11 $Y2=1.51
r72 23 29 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=1.14 $Y=1.685
+ $X2=1.275 $Y2=1.77
r73 23 25 7.46954 $w=2.68e-07 $l=1.75e-07 $layer=LI1_cond $X=1.14 $Y=1.685
+ $X2=1.14 $Y2=1.51
r74 21 42 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=0.995 $Y=2.465
+ $X2=0.995 $Y2=1.725
r75 18 40 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.955 $Y=0.655
+ $X2=0.955 $Y2=1.185
r76 15 22 5.30422 $w=1.5e-07 $l=9.5e-08 $layer=POLY_cond $X=0.64 $Y=1.65
+ $X2=0.545 $Y2=1.65
r77 14 42 32.8921 $w=3.95e-07 $l=7.5e-08 $layer=POLY_cond $X=1.077 $Y=1.65
+ $X2=1.077 $Y2=1.725
r78 14 26 19.7118 $w=3.95e-07 $l=1.4e-07 $layer=POLY_cond $X=1.077 $Y=1.65
+ $X2=1.077 $Y2=1.51
r79 14 15 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=0.88 $Y=1.65
+ $X2=0.64 $Y2=1.65
r80 11 22 20.4101 $w=1.5e-07 $l=8.44097e-08 $layer=POLY_cond $X=0.565 $Y=1.725
+ $X2=0.545 $Y2=1.65
r81 11 13 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=0.565 $Y=1.725
+ $X2=0.565 $Y2=2.465
r82 7 22 20.4101 $w=1.5e-07 $l=8.44097e-08 $layer=POLY_cond $X=0.525 $Y=1.575
+ $X2=0.545 $Y2=1.65
r83 7 9 471.745 $w=1.5e-07 $l=9.2e-07 $layer=POLY_cond $X=0.525 $Y=1.575
+ $X2=0.525 $Y2=0.655
r84 2 36 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=1.91
+ $Y=1.835 $X2=2.05 $Y2=1.98
r85 1 32 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.91
+ $Y=0.655 $X2=2.05 $Y2=0.865
.ends

.subckt PM_SKY130_FD_SC_LP__BUF_2%A 3 6 8 11 13
r26 11 14 56.1238 $w=3.95e-07 $l=2.4e-07 $layer=POLY_cond $X=1.712 $Y=1.35
+ $X2=1.712 $Y2=1.59
r27 11 13 45.5639 $w=3.95e-07 $l=1.65e-07 $layer=POLY_cond $X=1.712 $Y=1.35
+ $X2=1.712 $Y2=1.185
r28 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.68
+ $Y=1.35 $X2=1.68 $Y2=1.35
r29 6 14 289.713 $w=1.5e-07 $l=5.65e-07 $layer=POLY_cond $X=1.835 $Y=2.155
+ $X2=1.835 $Y2=1.59
r30 3 13 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.835 $Y=0.865
+ $X2=1.835 $Y2=1.185
.ends

.subckt PM_SKY130_FD_SC_LP__BUF_2%VPWR 1 2 7 9 15 19 21 28 29 35
r29 35 36 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r30 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r31 29 36 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r32 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r33 26 35 14.0645 $w=1.7e-07 $l=3.7e-07 $layer=LI1_cond $X=1.785 $Y=3.33
+ $X2=1.415 $Y2=3.33
r34 26 28 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.785 $Y=3.33
+ $X2=2.16 $Y2=3.33
r35 25 33 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r36 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r37 22 32 3.53348 $w=1.7e-07 $l=2.2e-07 $layer=LI1_cond $X=0.44 $Y=3.33 $X2=0.22
+ $Y2=3.33
r38 22 24 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=0.44 $Y=3.33
+ $X2=0.72 $Y2=3.33
r39 21 35 14.0645 $w=1.7e-07 $l=3.7e-07 $layer=LI1_cond $X=1.045 $Y=3.33
+ $X2=1.415 $Y2=3.33
r40 21 24 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=1.045 $Y=3.33
+ $X2=0.72 $Y2=3.33
r41 19 36 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r42 19 25 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r43 15 18 6.95019 $w=7.38e-07 $l=4.3e-07 $layer=LI1_cond $X=1.415 $Y=2.11
+ $X2=1.415 $Y2=2.54
r44 13 35 2.97738 $w=7.4e-07 $l=8.5e-08 $layer=LI1_cond $X=1.415 $Y=3.245
+ $X2=1.415 $Y2=3.33
r45 13 18 11.3951 $w=7.38e-07 $l=7.05e-07 $layer=LI1_cond $X=1.415 $Y=3.245
+ $X2=1.415 $Y2=2.54
r46 9 12 38.676 $w=1.93e-07 $l=6.8e-07 $layer=LI1_cond $X=0.342 $Y=2.27
+ $X2=0.342 $Y2=2.95
r47 7 32 3.32469 $w=1.95e-07 $l=1.58915e-07 $layer=LI1_cond $X=0.342 $Y=3.245
+ $X2=0.22 $Y2=3.33
r48 7 12 16.7786 $w=1.93e-07 $l=2.95e-07 $layer=LI1_cond $X=0.342 $Y=3.245
+ $X2=0.342 $Y2=2.95
r49 2 18 300 $w=1.7e-07 $l=7.71832e-07 $layer=licon1_PDIFF $count=2 $X=1.07
+ $Y=1.835 $X2=1.21 $Y2=2.54
r50 2 15 300 $w=1.7e-07 $l=6.7361e-07 $layer=licon1_PDIFF $count=2 $X=1.07
+ $Y=1.835 $X2=1.62 $Y2=2.11
r51 1 12 400 $w=1.7e-07 $l=1.17584e-06 $layer=licon1_PDIFF $count=1 $X=0.225
+ $Y=1.835 $X2=0.35 $Y2=2.95
r52 1 9 400 $w=1.7e-07 $l=4.93559e-07 $layer=licon1_PDIFF $count=1 $X=0.225
+ $Y=1.835 $X2=0.35 $Y2=2.27
.ends

.subckt PM_SKY130_FD_SC_LP__BUF_2%X 1 2 7 8 9 10 11 12 13 24 36 39
r20 37 39 1.43512 $w=2.63e-07 $l=3.3e-08 $layer=LI1_cond $X=0.742 $Y=2.177
+ $X2=0.742 $Y2=2.21
r21 36 48 0.512197 $w=2.23e-07 $l=1e-08 $layer=LI1_cond $X=0.722 $Y=2.035
+ $X2=0.722 $Y2=2.045
r22 13 45 5.00117 $w=2.63e-07 $l=1.15e-07 $layer=LI1_cond $X=0.742 $Y=2.775
+ $X2=0.742 $Y2=2.89
r23 12 13 16.0907 $w=2.63e-07 $l=3.7e-07 $layer=LI1_cond $X=0.742 $Y=2.405
+ $X2=0.742 $Y2=2.775
r24 12 39 8.48024 $w=2.63e-07 $l=1.95e-07 $layer=LI1_cond $X=0.742 $Y=2.405
+ $X2=0.742 $Y2=2.21
r25 11 37 4.1314 $w=2.63e-07 $l=9.5e-08 $layer=LI1_cond $X=0.742 $Y=2.082
+ $X2=0.742 $Y2=2.177
r26 11 48 1.90476 $w=2.63e-07 $l=3.7e-08 $layer=LI1_cond $X=0.742 $Y=2.082
+ $X2=0.742 $Y2=2.045
r27 11 36 1.94635 $w=2.23e-07 $l=3.8e-08 $layer=LI1_cond $X=0.722 $Y=1.997
+ $X2=0.722 $Y2=2.035
r28 10 11 17.0049 $w=2.23e-07 $l=3.32e-07 $layer=LI1_cond $X=0.722 $Y=1.665
+ $X2=0.722 $Y2=1.997
r29 9 10 18.9513 $w=2.23e-07 $l=3.7e-07 $layer=LI1_cond $X=0.722 $Y=1.295
+ $X2=0.722 $Y2=1.665
r30 8 9 18.9513 $w=2.23e-07 $l=3.7e-07 $layer=LI1_cond $X=0.722 $Y=0.925
+ $X2=0.722 $Y2=1.295
r31 7 8 18.9513 $w=2.23e-07 $l=3.7e-07 $layer=LI1_cond $X=0.722 $Y=0.555
+ $X2=0.722 $Y2=0.925
r32 7 24 6.91466 $w=2.23e-07 $l=1.35e-07 $layer=LI1_cond $X=0.722 $Y=0.555
+ $X2=0.722 $Y2=0.42
r33 2 45 400 $w=1.7e-07 $l=1.12282e-06 $layer=licon1_PDIFF $count=1 $X=0.64
+ $Y=1.835 $X2=0.78 $Y2=2.89
r34 2 39 400 $w=1.7e-07 $l=4.3946e-07 $layer=licon1_PDIFF $count=1 $X=0.64
+ $Y=1.835 $X2=0.78 $Y2=2.21
r35 1 24 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=0.6
+ $Y=0.235 $X2=0.74 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__BUF_2%VGND 1 2 7 9 13 18 20 27 28 34
r28 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r29 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r30 28 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.68
+ $Y2=0
r31 27 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r32 25 34 14.449 $w=1.7e-07 $l=3.9e-07 $layer=LI1_cond $X=1.785 $Y=0 $X2=1.395
+ $Y2=0
r33 25 27 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.785 $Y=0 $X2=2.16
+ $Y2=0
r34 24 32 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r35 23 24 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r36 21 31 4.36354 $w=1.7e-07 $l=2.2e-07 $layer=LI1_cond $X=0.44 $Y=0 $X2=0.22
+ $Y2=0
r37 21 23 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=0.44 $Y=0 $X2=0.72
+ $Y2=0
r38 20 34 14.449 $w=1.7e-07 $l=3.9e-07 $layer=LI1_cond $X=1.005 $Y=0 $X2=1.395
+ $Y2=0
r39 20 23 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.005 $Y=0 $X2=0.72
+ $Y2=0
r40 18 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r41 18 24 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r42 18 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r43 13 15 8.43389 $w=7.78e-07 $l=5.5e-07 $layer=LI1_cond $X=1.395 $Y=0.38
+ $X2=1.395 $Y2=0.93
r44 11 34 3.08259 $w=7.8e-07 $l=8.5e-08 $layer=LI1_cond $X=1.395 $Y=0.085
+ $X2=1.395 $Y2=0
r45 11 13 4.52363 $w=7.78e-07 $l=2.95e-07 $layer=LI1_cond $X=1.395 $Y=0.085
+ $X2=1.395 $Y2=0.38
r46 7 31 3.11398 $w=2.95e-07 $l=1.15521e-07 $layer=LI1_cond $X=0.292 $Y=0.085
+ $X2=0.22 $Y2=0
r47 7 9 11.5244 $w=2.93e-07 $l=2.95e-07 $layer=LI1_cond $X=0.292 $Y=0.085
+ $X2=0.292 $Y2=0.38
r48 2 15 182 $w=1.7e-07 $l=9.45026e-07 $layer=licon1_NDIFF $count=1 $X=1.03
+ $Y=0.235 $X2=1.62 $Y2=0.93
r49 2 15 182 $w=1.7e-07 $l=7.61791e-07 $layer=licon1_NDIFF $count=1 $X=1.03
+ $Y=0.235 $X2=1.17 $Y2=0.93
r50 2 13 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=1.03
+ $Y=0.235 $X2=1.17 $Y2=0.38
r51 1 9 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.185
+ $Y=0.235 $X2=0.31 $Y2=0.38
.ends

