* NGSPICE file created from sky130_fd_sc_lp__mux2i_0.ext - technology: sky130A

.subckt sky130_fd_sc_lp__mux2i_0 A0 A1 S VGND VNB VPB VPWR Y
M1000 a_465_491# A0 Y VPB phighvt w=640000u l=150000u
+  ad=1.76e+11p pd=1.83e+06u as=2.272e+11p ps=1.99e+06u
M1001 a_244_48# a_47_48# VGND VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=3.969e+11p ps=3.57e+06u
M1002 VPWR S a_47_48# VPB phighvt w=640000u l=150000u
+  ad=4.896e+11p pd=4.09e+06u as=1.696e+11p ps=1.81e+06u
M1003 VGND S a_436_48# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1004 VPWR S a_465_491# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_436_48# A1 Y VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.764e+11p ps=1.68e+06u
M1006 VGND S a_47_48# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1007 a_292_491# a_47_48# VPWR VPB phighvt w=640000u l=150000u
+  ad=1.344e+11p pd=1.7e+06u as=0p ps=0u
M1008 Y A0 a_244_48# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 Y A1 a_292_491# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

