* File: sky130_fd_sc_lp__clkinvlp_2.pxi.spice
* Created: Fri Aug 28 10:18:48 2020
* 
x_PM_SKY130_FD_SC_LP__CLKINVLP_2%A N_A_M1000_g N_A_c_27_n N_A_M1001_g N_A_c_28_n
+ N_A_M1002_g N_A_M1003_g A A N_A_c_30_n PM_SKY130_FD_SC_LP__CLKINVLP_2%A
x_PM_SKY130_FD_SC_LP__CLKINVLP_2%VPWR N_VPWR_M1000_s N_VPWR_M1003_s
+ N_VPWR_c_66_n N_VPWR_c_67_n N_VPWR_c_68_n N_VPWR_c_69_n N_VPWR_c_70_n VPWR
+ N_VPWR_c_71_n N_VPWR_c_65_n PM_SKY130_FD_SC_LP__CLKINVLP_2%VPWR
x_PM_SKY130_FD_SC_LP__CLKINVLP_2%Y N_Y_M1002_d N_Y_M1000_d N_Y_c_86_n Y Y Y Y Y
+ Y Y PM_SKY130_FD_SC_LP__CLKINVLP_2%Y
x_PM_SKY130_FD_SC_LP__CLKINVLP_2%VGND N_VGND_M1001_s N_VGND_c_113_n VGND
+ N_VGND_c_114_n N_VGND_c_115_n N_VGND_c_116_n N_VGND_c_117_n
+ PM_SKY130_FD_SC_LP__CLKINVLP_2%VGND
cc_1 VNB N_A_c_27_n 0.0211447f $X=-0.19 $Y=-0.245 $X2=0.85 $Y2=0.995
cc_2 VNB N_A_c_28_n 0.0202123f $X=-0.19 $Y=-0.245 $X2=1.24 $Y2=0.995
cc_3 VNB A 0.040355f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_4 VNB N_A_c_30_n 0.138812f $X=-0.19 $Y=-0.245 $X2=1.24 $Y2=1.33
cc_5 VNB N_VPWR_c_65_n 0.0840719f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=1.387
cc_6 VNB N_Y_c_86_n 0.023331f $X=-0.19 $Y=-0.245 $X2=1.36 $Y2=1.665
cc_7 VNB Y 0.0178881f $X=-0.19 $Y=-0.245 $X2=1.36 $Y2=2.48
cc_8 VNB N_VGND_c_113_n 0.0249118f $X=-0.19 $Y=-0.245 $X2=0.85 $Y2=0.61
cc_9 VNB N_VGND_c_114_n 0.0170996f $X=-0.19 $Y=-0.245 $X2=1.24 $Y2=0.61
cc_10 VNB N_VGND_c_115_n 0.0325108f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_11 VNB N_VGND_c_116_n 0.159247f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_VGND_c_117_n 0.00589254f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VPB N_A_M1000_g 0.0439229f $X=-0.19 $Y=1.655 $X2=0.83 $Y2=2.48
cc_14 VPB N_A_M1003_g 0.0446986f $X=-0.19 $Y=1.655 $X2=1.36 $Y2=2.48
cc_15 VPB A 0.0206558f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_16 VPB N_A_c_30_n 0.0142895f $X=-0.19 $Y=1.655 $X2=1.24 $Y2=1.33
cc_17 VPB N_VPWR_c_66_n 0.0504708f $X=-0.19 $Y=1.655 $X2=1.24 $Y2=0.61
cc_18 VPB N_VPWR_c_67_n 0.0120923f $X=-0.19 $Y=1.655 $X2=1.36 $Y2=2.48
cc_19 VPB N_VPWR_c_68_n 0.0632149f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_20 VPB N_VPWR_c_69_n 0.0148721f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_21 VPB N_VPWR_c_70_n 0.00598038f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_22 VPB N_VPWR_c_71_n 0.020628f $X=-0.19 $Y=1.655 $X2=1.24 $Y2=1.33
cc_23 VPB N_VPWR_c_65_n 0.0596418f $X=-0.19 $Y=1.655 $X2=0.69 $Y2=1.387
cc_24 VPB Y 0.00243503f $X=-0.19 $Y=1.655 $X2=1.36 $Y2=2.48
cc_25 VPB Y 0.00232136f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_26 VPB Y 0.0032582f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_27 N_A_M1000_g N_VPWR_c_66_n 0.0235567f $X=0.83 $Y=2.48 $X2=0 $Y2=0
cc_28 N_A_M1003_g N_VPWR_c_66_n 8.05893e-19 $X=1.36 $Y=2.48 $X2=0 $Y2=0
cc_29 A N_VPWR_c_66_n 0.0291664f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_30 N_A_c_30_n N_VPWR_c_66_n 0.00179491f $X=1.24 $Y=1.33 $X2=0 $Y2=0
cc_31 N_A_M1003_g N_VPWR_c_68_n 0.00595795f $X=1.36 $Y=2.48 $X2=0 $Y2=0
cc_32 N_A_M1000_g N_VPWR_c_71_n 0.00687065f $X=0.83 $Y=2.48 $X2=0 $Y2=0
cc_33 N_A_M1003_g N_VPWR_c_71_n 0.00696917f $X=1.36 $Y=2.48 $X2=0 $Y2=0
cc_34 N_A_M1000_g N_VPWR_c_65_n 0.0129282f $X=0.83 $Y=2.48 $X2=0 $Y2=0
cc_35 N_A_M1003_g N_VPWR_c_65_n 0.012542f $X=1.36 $Y=2.48 $X2=0 $Y2=0
cc_36 N_A_c_27_n N_Y_c_86_n 0.0036434f $X=0.85 $Y=0.995 $X2=0 $Y2=0
cc_37 N_A_c_28_n N_Y_c_86_n 0.012538f $X=1.24 $Y=0.995 $X2=0 $Y2=0
cc_38 N_A_c_30_n N_Y_c_86_n 0.00445703f $X=1.24 $Y=1.33 $X2=0 $Y2=0
cc_39 N_A_M1000_g Y 0.00555265f $X=0.83 $Y=2.48 $X2=0 $Y2=0
cc_40 N_A_c_27_n Y 0.00518284f $X=0.85 $Y=0.995 $X2=0 $Y2=0
cc_41 N_A_c_28_n Y 0.00817338f $X=1.24 $Y=0.995 $X2=0 $Y2=0
cc_42 N_A_M1003_g Y 0.0168263f $X=1.36 $Y=2.48 $X2=0 $Y2=0
cc_43 A Y 0.0594801f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_44 N_A_c_30_n Y 0.0485337f $X=1.24 $Y=1.33 $X2=0 $Y2=0
cc_45 N_A_M1000_g Y 0.0153217f $X=0.83 $Y=2.48 $X2=0 $Y2=0
cc_46 N_A_M1003_g Y 0.0155972f $X=1.36 $Y=2.48 $X2=0 $Y2=0
cc_47 N_A_M1000_g Y 0.00490991f $X=0.83 $Y=2.48 $X2=0 $Y2=0
cc_48 N_A_M1003_g Y 0.00359763f $X=1.36 $Y=2.48 $X2=0 $Y2=0
cc_49 N_A_c_27_n N_VGND_c_113_n 0.0125054f $X=0.85 $Y=0.995 $X2=0 $Y2=0
cc_50 N_A_c_28_n N_VGND_c_113_n 0.00107387f $X=1.24 $Y=0.995 $X2=0 $Y2=0
cc_51 A N_VGND_c_113_n 0.0212051f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_52 N_A_c_30_n N_VGND_c_113_n 0.00774745f $X=1.24 $Y=1.33 $X2=0 $Y2=0
cc_53 N_A_c_27_n N_VGND_c_115_n 0.00407525f $X=0.85 $Y=0.995 $X2=0 $Y2=0
cc_54 N_A_c_28_n N_VGND_c_115_n 0.00306316f $X=1.24 $Y=0.995 $X2=0 $Y2=0
cc_55 N_A_c_27_n N_VGND_c_116_n 0.00777674f $X=0.85 $Y=0.995 $X2=0 $Y2=0
cc_56 N_A_c_28_n N_VGND_c_116_n 0.00449031f $X=1.24 $Y=0.995 $X2=0 $Y2=0
cc_57 N_VPWR_c_71_n Y 0.0184863f $X=1.49 $Y=3.33 $X2=0 $Y2=0
cc_58 N_VPWR_c_65_n Y 0.0139841f $X=1.68 $Y=3.33 $X2=0 $Y2=0
cc_59 N_VPWR_c_66_n Y 0.0693797f $X=0.565 $Y=2.125 $X2=0 $Y2=0
cc_60 N_VPWR_c_68_n Y 0.0415535f $X=1.625 $Y=2.125 $X2=0 $Y2=0
cc_61 N_Y_c_86_n N_VGND_c_113_n 0.0292162f $X=1.455 $Y=0.545 $X2=0 $Y2=0
cc_62 N_Y_c_86_n N_VGND_c_115_n 0.0289255f $X=1.455 $Y=0.545 $X2=0 $Y2=0
cc_63 N_Y_c_86_n N_VGND_c_116_n 0.0210679f $X=1.455 $Y=0.545 $X2=0 $Y2=0
cc_64 N_Y_c_86_n A_185_67# 0.00445571f $X=1.455 $Y=0.545 $X2=-0.19 $Y2=-0.245
cc_65 Y A_185_67# 0.00146339f $X=1.115 $Y=0.84 $X2=-0.19 $Y2=-0.245
