* File: sky130_fd_sc_lp__nand2_lp.pex.spice
* Created: Wed Sep  2 10:03:12 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__NAND2_LP%B 3 7 9 11 12 13 14 15 22 23
r29 22 25 82.9202 $w=5e-07 $l=5.05e-07 $layer=POLY_cond $X=0.355 $Y=1.12
+ $X2=0.355 $Y2=1.625
r30 22 24 46.5382 $w=5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.355 $Y=1.12
+ $X2=0.355 $Y2=0.955
r31 22 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.27
+ $Y=1.12 $X2=0.27 $Y2=1.12
r32 14 15 14.4544 $w=2.93e-07 $l=3.7e-07 $layer=LI1_cond $X=0.252 $Y=2.405
+ $X2=0.252 $Y2=2.775
r33 13 14 14.4544 $w=2.93e-07 $l=3.7e-07 $layer=LI1_cond $X=0.252 $Y=2.035
+ $X2=0.252 $Y2=2.405
r34 12 13 14.4544 $w=2.93e-07 $l=3.7e-07 $layer=LI1_cond $X=0.252 $Y=1.665
+ $X2=0.252 $Y2=2.035
r35 11 12 14.4544 $w=2.93e-07 $l=3.7e-07 $layer=LI1_cond $X=0.252 $Y=1.295
+ $X2=0.252 $Y2=1.665
r36 11 23 6.83653 $w=2.93e-07 $l=1.75e-07 $layer=LI1_cond $X=0.252 $Y=1.295
+ $X2=0.252 $Y2=1.12
r37 7 9 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=0.53 $Y=2.045 $X2=0.53
+ $Y2=2.735
r38 7 25 215.362 $w=1.5e-07 $l=4.2e-07 $layer=POLY_cond $X=0.53 $Y=2.045
+ $X2=0.53 $Y2=1.625
r39 3 24 235.872 $w=1.5e-07 $l=4.6e-07 $layer=POLY_cond $X=0.53 $Y=0.495
+ $X2=0.53 $Y2=0.955
.ends

.subckt PM_SKY130_FD_SC_LP__NAND2_LP%A 3 7 9 13 15 16 19
r28 19 20 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.055
+ $Y=1.07 $X2=1.055 $Y2=1.07
r29 16 20 2.93854 $w=6.02e-07 $l=1.45e-07 $layer=LI1_cond $X=1.2 $Y=1.24
+ $X2=1.055 $Y2=1.24
r30 14 19 58.221 $w=3.35e-07 $l=3.38e-07 $layer=POLY_cond $X=1.052 $Y=1.408
+ $X2=1.052 $Y2=1.07
r31 14 15 46.5995 $w=3.35e-07 $l=1.67e-07 $layer=POLY_cond $X=1.052 $Y=1.408
+ $X2=1.052 $Y2=1.575
r32 13 19 2.58377 $w=3.35e-07 $l=1.5e-08 $layer=POLY_cond $X=1.052 $Y=1.055
+ $X2=1.052 $Y2=1.07
r33 12 13 43.6712 $w=3.35e-07 $l=1.5e-07 $layer=POLY_cond $X=1.032 $Y=0.905
+ $X2=1.032 $Y2=1.055
r34 7 9 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=0.96 $Y=2.045 $X2=0.96
+ $Y2=2.735
r35 7 15 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=0.96 $Y=2.045 $X2=0.96
+ $Y2=1.575
r36 3 12 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=0.92 $Y=0.495
+ $X2=0.92 $Y2=0.905
.ends

.subckt PM_SKY130_FD_SC_LP__NAND2_LP%Y 1 2 8 9 10 12 16 17
r35 16 21 2.39909 $w=4.6e-07 $l=8.5e-08 $layer=LI1_cond $X=0.665 $Y=2.045
+ $X2=0.75 $Y2=2.045
r36 16 17 10.9987 $w=4.58e-07 $l=4.23e-07 $layer=LI1_cond $X=0.777 $Y=2.045
+ $X2=1.2 $Y2=2.045
r37 16 21 0.702046 $w=4.58e-07 $l=2.7e-08 $layer=LI1_cond $X=0.777 $Y=2.045
+ $X2=0.75 $Y2=2.045
r38 12 14 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=1.135 $Y=0.495
+ $X2=1.135 $Y2=0.64
r39 9 14 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.97 $Y=0.64
+ $X2=1.135 $Y2=0.64
r40 9 10 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=0.97 $Y=0.64 $X2=0.75
+ $Y2=0.64
r41 8 16 6.49166 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=0.665 $Y=1.815
+ $X2=0.665 $Y2=2.045
r42 7 10 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.665 $Y=0.725
+ $X2=0.75 $Y2=0.64
r43 7 8 71.1123 $w=1.68e-07 $l=1.09e-06 $layer=LI1_cond $X=0.665 $Y=0.725
+ $X2=0.665 $Y2=1.815
r44 2 16 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=0.605
+ $Y=1.835 $X2=0.745 $Y2=2.045
r45 1 12 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.995
+ $Y=0.285 $X2=1.135 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__NAND2_LP%VPWR 1 6 8 10 17 18 21
r17 17 18 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r18 15 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.91 $Y=3.33
+ $X2=0.745 $Y2=3.33
r19 15 17 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=0.91 $Y=3.33 $X2=1.2
+ $Y2=3.33
r20 12 13 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r21 10 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.58 $Y=3.33
+ $X2=0.745 $Y2=3.33
r22 10 12 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=0.58 $Y=3.33
+ $X2=0.24 $Y2=3.33
r23 8 18 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33 $X2=1.2
+ $Y2=3.33
r24 8 13 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r25 8 21 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33 $X2=0.72
+ $Y2=3.33
r26 4 21 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.745 $Y=3.245
+ $X2=0.745 $Y2=3.33
r27 4 6 17.8105 $w=3.28e-07 $l=5.1e-07 $layer=LI1_cond $X=0.745 $Y=3.245
+ $X2=0.745 $Y2=2.735
r28 1 6 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=0.605
+ $Y=2.525 $X2=0.745 $Y2=2.735
.ends

.subckt PM_SKY130_FD_SC_LP__NAND2_LP%VGND 1 4 6 8 12 13
r19 16 17 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r20 12 13 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r21 10 16 3.96842 $w=1.7e-07 $l=2e-07 $layer=LI1_cond $X=0.4 $Y=0 $X2=0.2 $Y2=0
r22 10 12 52.1925 $w=1.68e-07 $l=8e-07 $layer=LI1_cond $X=0.4 $Y=0 $X2=1.2 $Y2=0
r23 8 13 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r24 8 17 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r25 4 16 3.17474 $w=2.5e-07 $l=1.16619e-07 $layer=LI1_cond $X=0.275 $Y=0.085
+ $X2=0.2 $Y2=0
r26 4 6 18.9001 $w=2.48e-07 $l=4.1e-07 $layer=LI1_cond $X=0.275 $Y=0.085
+ $X2=0.275 $Y2=0.495
r27 1 6 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.17
+ $Y=0.285 $X2=0.315 $Y2=0.495
.ends

