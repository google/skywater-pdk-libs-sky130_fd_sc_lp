* File: sky130_fd_sc_lp__nor4b_2.spice
* Created: Fri Aug 28 10:58:15 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__nor4b_2.pex.spice"
.subckt sky130_fd_sc_lp__nor4b_2  VNB VPB D_N C B A VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A	A
* B	B
* C	C
* D_N	D_N
* VPB	VPB
* VNB	VNB
MM1008 N_VGND_M1008_d N_D_N_M1008_g N_A_27_535#_M1008_s VNB NSHORT L=0.15 W=0.42
+ AD=0.161 AS=0.1113 PD=1.09667 PS=1.37 NRD=81.42 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75004.5 A=0.063 P=1.14 MULT=1
MM1003 N_Y_M1003_d N_C_M1003_g N_VGND_M1008_d VNB NSHORT L=0.15 W=0.84 AD=0.1176
+ AS=0.322 PD=1.12 PS=2.19333 NRD=0 NRS=22.848 M=1 R=5.6 SA=75000.7 SB=75003.5
+ A=0.126 P=1.98 MULT=1
MM1002 N_Y_M1003_d N_A_27_535#_M1002_g N_VGND_M1002_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.1
+ SB=75003.1 A=0.126 P=1.98 MULT=1
MM1014 N_Y_M1014_d N_A_27_535#_M1014_g N_VGND_M1002_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.6
+ SB=75002.6 A=0.126 P=1.98 MULT=1
MM1009 N_Y_M1014_d N_C_M1009_g N_VGND_M1009_s VNB NSHORT L=0.15 W=0.84 AD=0.1176
+ AS=0.2478 PD=1.12 PS=1.43 NRD=0 NRS=22.848 M=1 R=5.6 SA=75002 SB=75002.2
+ A=0.126 P=1.98 MULT=1
MM1000 N_Y_M1000_d N_B_M1000_g N_VGND_M1009_s VNB NSHORT L=0.15 W=0.84 AD=0.1176
+ AS=0.2478 PD=1.12 PS=1.43 NRD=0 NRS=21.42 M=1 R=5.6 SA=75002.7 SB=75001.5
+ A=0.126 P=1.98 MULT=1
MM1007 N_VGND_M1007_d N_A_M1007_g N_Y_M1000_d VNB NSHORT L=0.15 W=0.84 AD=0.1176
+ AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75003.2 SB=75001.1 A=0.126
+ P=1.98 MULT=1
MM1011 N_VGND_M1007_d N_A_M1011_g N_Y_M1011_s VNB NSHORT L=0.15 W=0.84 AD=0.1176
+ AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75003.6 SB=75000.6 A=0.126
+ P=1.98 MULT=1
MM1005 N_Y_M1011_s N_B_M1005_g N_VGND_M1005_s VNB NSHORT L=0.15 W=0.84 AD=0.1176
+ AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75004 SB=75000.2 A=0.126
+ P=1.98 MULT=1
MM1012 N_VPWR_M1012_d N_D_N_M1012_g N_A_27_535#_M1012_s VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1113 AS=0.1113 PD=1.37 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1015 N_A_229_367#_M1015_d N_C_M1015_g N_A_312_367#_M1015_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75003.5 A=0.189 P=2.82 MULT=1
MM1004 N_A_312_367#_M1015_s N_A_27_535#_M1004_g N_Y_M1004_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75003.1 A=0.189 P=2.82 MULT=1
MM1010 N_A_312_367#_M1010_d N_A_27_535#_M1010_g N_Y_M1004_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75002.6 A=0.189 P=2.82 MULT=1
MM1017 N_A_229_367#_M1017_d N_C_M1017_g N_A_312_367#_M1010_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.2268 AS=0.1764 PD=1.62 PS=1.54 NRD=12.4898 NRS=0 M=1 R=8.4
+ SA=75001.5 SB=75002.2 A=0.189 P=2.82 MULT=1
MM1001 N_A_229_367#_M1017_d N_B_M1001_g N_A_672_367#_M1001_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.2268 AS=0.3213 PD=1.62 PS=1.77 NRD=0 NRS=16.4101 M=1 R=8.4
+ SA=75002 SB=75001.7 A=0.189 P=2.82 MULT=1
MM1006 N_A_672_367#_M1001_s N_A_M1006_g N_VPWR_M1006_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3213 AS=0.1764 PD=1.77 PS=1.54 NRD=19.5424 NRS=0 M=1 R=8.4 SA=75002.6
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1013 N_A_672_367#_M1013_d N_A_M1013_g N_VPWR_M1006_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75003.1
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1016 N_A_229_367#_M1016_d N_B_M1016_g N_A_672_367#_M1013_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75003.5
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX18_noxref VNB VPB NWDIODE A=10.5559 P=15.05
*
.include "sky130_fd_sc_lp__nor4b_2.pxi.spice"
*
.ends
*
*
