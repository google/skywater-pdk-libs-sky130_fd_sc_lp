* File: sky130_fd_sc_lp__o2bb2a_1.pex.spice
* Created: Fri Aug 28 11:11:41 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O2BB2A_1%A_80_21# 1 2 9 12 16 17 19 20 22 24 26 27
+ 28 30 33 34 39 42
c102 28 0 1.7714e-19 $X=2.37 $Y=1.14
c103 27 0 7.16669e-20 $X=2.67 $Y=1.14
r104 37 39 3.62806 $w=2.68e-07 $l=8.5e-08 $layer=LI1_cond $X=2.67 $Y=2.785
+ $X2=2.755 $Y2=2.785
r105 32 34 1.08465 $w=3.38e-07 $l=3.2e-08 $layer=LI1_cond $X=2.24 $Y=0.45
+ $X2=2.272 $Y2=0.45
r106 32 33 6.42278 $w=3.38e-07 $l=1.65e-07 $layer=LI1_cond $X=2.24 $Y=0.45
+ $X2=2.075 $Y2=0.45
r107 30 39 3.44395 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=2.755 $Y=2.65
+ $X2=2.755 $Y2=2.785
r108 29 30 92.9679 $w=1.68e-07 $l=1.425e-06 $layer=LI1_cond $X=2.755 $Y=1.225
+ $X2=2.755 $Y2=2.65
r109 27 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.67 $Y=1.14
+ $X2=2.755 $Y2=1.225
r110 27 28 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=2.67 $Y=1.14 $X2=2.37
+ $Y2=1.14
r111 26 28 6.85817 $w=1.7e-07 $l=1.33918e-07 $layer=LI1_cond $X=2.272 $Y=1.055
+ $X2=2.37 $Y2=1.14
r112 25 34 4.00821 $w=1.95e-07 $l=1.7e-07 $layer=LI1_cond $X=2.272 $Y=0.62
+ $X2=2.272 $Y2=0.45
r113 25 26 24.7413 $w=1.93e-07 $l=4.35e-07 $layer=LI1_cond $X=2.272 $Y=0.62
+ $X2=2.272 $Y2=1.055
r114 24 33 34.8038 $w=2.48e-07 $l=7.55e-07 $layer=LI1_cond $X=1.32 $Y=0.405
+ $X2=2.075 $Y2=0.405
r115 21 24 6.83662 $w=2.5e-07 $l=1.9051e-07 $layer=LI1_cond $X=1.182 $Y=0.53
+ $X2=1.32 $Y2=0.405
r116 21 22 13.8293 $w=2.73e-07 $l=3.3e-07 $layer=LI1_cond $X=1.182 $Y=0.53
+ $X2=1.182 $Y2=0.86
r117 19 22 7.32204 $w=1.7e-07 $l=1.74396e-07 $layer=LI1_cond $X=1.045 $Y=0.945
+ $X2=1.182 $Y2=0.86
r118 19 20 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=1.045 $Y=0.945
+ $X2=0.865 $Y2=0.945
r119 17 43 45.5639 $w=3.95e-07 $l=1.65e-07 $layer=POLY_cond $X=0.597 $Y=1.35
+ $X2=0.597 $Y2=1.515
r120 17 42 45.5639 $w=3.95e-07 $l=1.65e-07 $layer=POLY_cond $X=0.597 $Y=1.35
+ $X2=0.597 $Y2=1.185
r121 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.63
+ $Y=1.35 $X2=0.63 $Y2=1.35
r122 14 20 7.85115 $w=1.7e-07 $l=2.08207e-07 $layer=LI1_cond $X=0.695 $Y=1.03
+ $X2=0.865 $Y2=0.945
r123 14 16 10.8465 $w=3.38e-07 $l=3.2e-07 $layer=LI1_cond $X=0.695 $Y=1.03
+ $X2=0.695 $Y2=1.35
r124 12 43 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=0.475 $Y=2.465
+ $X2=0.475 $Y2=1.515
r125 9 42 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.475 $Y=0.655
+ $X2=0.475 $Y2=1.185
r126 2 37 600 $w=1.7e-07 $l=3.58225e-07 $layer=licon1_PDIFF $count=1 $X=2.53
+ $Y=2.46 $X2=2.67 $Y2=2.755
r127 1 32 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=2.115
+ $Y=0.235 $X2=2.24 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__O2BB2A_1%A1_N 3 6 9 11 12 13 14 19
c45 12 0 1.62131e-19 $X=1.2 $Y=1.295
r46 19 21 45.5639 $w=3.95e-07 $l=1.65e-07 $layer=POLY_cond $X=1.232 $Y=1.74
+ $X2=1.232 $Y2=1.575
r47 13 14 12.3595 $w=3.43e-07 $l=3.7e-07 $layer=LI1_cond $X=1.207 $Y=1.665
+ $X2=1.207 $Y2=2.035
r48 13 19 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.2 $Y=1.74
+ $X2=1.2 $Y2=1.74
r49 12 13 12.3595 $w=3.43e-07 $l=3.7e-07 $layer=LI1_cond $X=1.207 $Y=1.295
+ $X2=1.207 $Y2=1.665
r50 9 11 217.926 $w=1.5e-07 $l=4.25e-07 $layer=POLY_cond $X=1.355 $Y=2.67
+ $X2=1.355 $Y2=2.245
r51 6 11 50.0695 $w=3.95e-07 $l=1.97e-07 $layer=POLY_cond $X=1.232 $Y=2.048
+ $X2=1.232 $Y2=2.245
r52 5 19 4.50555 $w=3.95e-07 $l=3.2e-08 $layer=POLY_cond $X=1.232 $Y=1.772
+ $X2=1.232 $Y2=1.74
r53 5 6 38.8604 $w=3.95e-07 $l=2.76e-07 $layer=POLY_cond $X=1.232 $Y=1.772
+ $X2=1.232 $Y2=2.048
r54 3 21 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=1.11 $Y=0.865
+ $X2=1.11 $Y2=1.575
.ends

.subckt PM_SKY130_FD_SC_LP__O2BB2A_1%A2_N 1 3 8 12 14 17 18 19
c50 18 0 6.68251e-20 $X=1.835 $Y=2.035
c51 17 0 3.07487e-19 $X=1.835 $Y=2.035
c52 12 0 1.7714e-19 $X=1.745 $Y=1.26
r53 17 20 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.835 $Y=2.035
+ $X2=1.835 $Y2=2.2
r54 17 19 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.835 $Y=2.035
+ $X2=1.835 $Y2=1.87
r55 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.835
+ $Y=2.035 $X2=1.835 $Y2=2.035
r56 14 18 4.63971 $w=3.83e-07 $l=1.55e-07 $layer=LI1_cond $X=1.68 $Y=1.947
+ $X2=1.835 $Y2=1.947
r57 10 12 125.628 $w=1.5e-07 $l=2.45e-07 $layer=POLY_cond $X=1.5 $Y=1.26
+ $X2=1.745 $Y2=1.26
r58 8 20 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=1.785 $Y=2.67 $X2=1.785
+ $Y2=2.2
r59 4 12 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.745 $Y=1.335
+ $X2=1.745 $Y2=1.26
r60 4 19 274.33 $w=1.5e-07 $l=5.35e-07 $layer=POLY_cond $X=1.745 $Y=1.335
+ $X2=1.745 $Y2=1.87
r61 1 10 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.5 $Y=1.185 $X2=1.5
+ $Y2=1.26
r62 1 3 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.5 $Y=1.185 $X2=1.5
+ $Y2=0.865
.ends

.subckt PM_SKY130_FD_SC_LP__O2BB2A_1%A_286_492# 1 2 9 13 17 18 21 25 27 28 29 30
+ 31 32 35
c78 31 0 1.47281e-19 $X=2.37 $Y=1.575
c79 28 0 1.45356e-19 $X=1.675 $Y=2.395
c80 27 0 1.63416e-19 $X=2.24 $Y=2.395
c81 18 0 1.98721e-19 $X=2.405 $Y=2.075
c82 13 0 6.68251e-20 $X=2.455 $Y=2.67
r83 34 35 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.405
+ $Y=1.57 $X2=2.405 $Y2=1.57
r84 31 34 2.85134 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=2.37 $Y=1.575
+ $X2=2.37 $Y2=1.49
r85 31 32 32.5787 $w=2.58e-07 $l=7.35e-07 $layer=LI1_cond $X=2.37 $Y=1.575
+ $X2=2.37 $Y2=2.31
r86 29 34 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.24 $Y=1.49 $X2=2.37
+ $Y2=1.49
r87 29 30 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=2.24 $Y=1.49
+ $X2=1.88 $Y2=1.49
r88 27 32 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=2.24 $Y=2.395
+ $X2=2.37 $Y2=2.31
r89 27 28 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=2.24 $Y=2.395
+ $X2=1.675 $Y2=2.395
r90 23 30 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.715 $Y=1.405
+ $X2=1.88 $Y2=1.49
r91 23 25 18.8582 $w=3.28e-07 $l=5.4e-07 $layer=LI1_cond $X=1.715 $Y=1.405
+ $X2=1.715 $Y2=0.865
r92 19 28 10.5078 $w=1.38e-07 $l=1.56844e-07 $layer=LI1_cond $X=1.555 $Y=2.48
+ $X2=1.675 $Y2=2.395
r93 19 21 9.12351 $w=2.38e-07 $l=1.9e-07 $layer=LI1_cond $X=1.555 $Y=2.48
+ $X2=1.555 $Y2=2.67
r94 17 35 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.405 $Y=1.91
+ $X2=2.405 $Y2=1.57
r95 17 18 40.8701 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.405 $Y=1.91
+ $X2=2.405 $Y2=2.075
r96 16 35 40.8701 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.405 $Y=1.405
+ $X2=2.405 $Y2=1.57
r97 13 18 305.096 $w=1.5e-07 $l=5.95e-07 $layer=POLY_cond $X=2.455 $Y=2.67
+ $X2=2.455 $Y2=2.075
r98 9 16 492.255 $w=1.5e-07 $l=9.6e-07 $layer=POLY_cond $X=2.455 $Y=0.445
+ $X2=2.455 $Y2=1.405
r99 2 21 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=1.43
+ $Y=2.46 $X2=1.57 $Y2=2.67
r100 1 25 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.575
+ $Y=0.655 $X2=1.715 $Y2=0.865
.ends

.subckt PM_SKY130_FD_SC_LP__O2BB2A_1%B2 3 7 9 11 20
c41 20 0 1.47281e-19 $X=3.105 $Y=1.465
c42 7 0 1.63416e-19 $X=2.885 $Y=2.67
r43 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.105
+ $Y=1.465 $X2=3.105 $Y2=1.465
r44 17 20 38.4695 $w=3.3e-07 $l=2.2e-07 $layer=POLY_cond $X=2.885 $Y=1.465
+ $X2=3.105 $Y2=1.465
r45 9 11 8.97059 $w=6.38e-07 $l=4.8e-07 $layer=LI1_cond $X=3.12 $Y=1.43 $X2=3.6
+ $Y2=1.43
r46 9 21 0.280331 $w=6.38e-07 $l=1.5e-08 $layer=LI1_cond $X=3.12 $Y=1.43
+ $X2=3.105 $Y2=1.43
r47 5 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.885 $Y=1.63
+ $X2=2.885 $Y2=1.465
r48 5 7 533.277 $w=1.5e-07 $l=1.04e-06 $layer=POLY_cond $X=2.885 $Y=1.63
+ $X2=2.885 $Y2=2.67
r49 1 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.885 $Y=1.3
+ $X2=2.885 $Y2=1.465
r50 1 3 438.415 $w=1.5e-07 $l=8.55e-07 $layer=POLY_cond $X=2.885 $Y=1.3
+ $X2=2.885 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__O2BB2A_1%B1 3 7 10 13 15 16 24
c36 13 0 2.73064e-20 $X=3.585 $Y=0.985
c37 10 0 4.43605e-20 $X=3.585 $Y=1.87
r38 22 24 38.4695 $w=3.3e-07 $l=2.2e-07 $layer=POLY_cond $X=3.365 $Y=2.035
+ $X2=3.585 $Y2=2.035
r39 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.365
+ $Y=2.035 $X2=3.365 $Y2=2.035
r40 19 22 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=3.275 $Y=2.035
+ $X2=3.365 $Y2=2.035
r41 16 23 9.33876 $w=2.88e-07 $l=2.35e-07 $layer=LI1_cond $X=3.6 $Y=2.065
+ $X2=3.365 $Y2=2.065
r42 15 23 9.73616 $w=2.88e-07 $l=2.45e-07 $layer=LI1_cond $X=3.12 $Y=2.065
+ $X2=3.365 $Y2=2.065
r43 11 13 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=3.315 $Y=0.985
+ $X2=3.585 $Y2=0.985
r44 10 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.585 $Y=1.87
+ $X2=3.585 $Y2=2.035
r45 9 13 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.585 $Y=1.06
+ $X2=3.585 $Y2=0.985
r46 9 10 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=3.585 $Y=1.06
+ $X2=3.585 $Y2=1.87
r47 5 11 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.315 $Y=0.91
+ $X2=3.315 $Y2=0.985
r48 5 7 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.315 $Y=0.91
+ $X2=3.315 $Y2=0.445
r49 1 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.275 $Y=2.2
+ $X2=3.275 $Y2=2.035
r50 1 3 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=3.275 $Y=2.2 $X2=3.275
+ $Y2=2.67
.ends

.subckt PM_SKY130_FD_SC_LP__O2BB2A_1%X 1 2 7 8 9 10 11 12 13 22
r11 13 40 5.98384 $w=2.58e-07 $l=1.35e-07 $layer=LI1_cond $X=0.225 $Y=2.775
+ $X2=0.225 $Y2=2.91
r12 12 13 16.4002 $w=2.58e-07 $l=3.7e-07 $layer=LI1_cond $X=0.225 $Y=2.405
+ $X2=0.225 $Y2=2.775
r13 11 12 18.838 $w=2.58e-07 $l=4.25e-07 $layer=LI1_cond $X=0.225 $Y=1.98
+ $X2=0.225 $Y2=2.405
r14 10 11 13.9623 $w=2.58e-07 $l=3.15e-07 $layer=LI1_cond $X=0.225 $Y=1.665
+ $X2=0.225 $Y2=1.98
r15 9 10 16.4002 $w=2.58e-07 $l=3.7e-07 $layer=LI1_cond $X=0.225 $Y=1.295
+ $X2=0.225 $Y2=1.665
r16 8 9 16.4002 $w=2.58e-07 $l=3.7e-07 $layer=LI1_cond $X=0.225 $Y=0.925
+ $X2=0.225 $Y2=1.295
r17 7 8 16.4002 $w=2.58e-07 $l=3.7e-07 $layer=LI1_cond $X=0.225 $Y=0.555
+ $X2=0.225 $Y2=0.925
r18 7 22 5.98384 $w=2.58e-07 $l=1.35e-07 $layer=LI1_cond $X=0.225 $Y=0.555
+ $X2=0.225 $Y2=0.42
r19 2 40 400 $w=1.7e-07 $l=1.13578e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.835 $X2=0.26 $Y2=2.91
r20 2 11 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.835 $X2=0.26 $Y2=1.98
r21 1 22 91 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__O2BB2A_1%VPWR 1 2 3 12 16 18 20 22 24 29 34 40 47 51
c54 16 0 1.98721e-19 $X=2.135 $Y=2.755
r55 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r56 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r57 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r58 40 43 10.6677 $w=7.38e-07 $l=6.6e-07 $layer=LI1_cond $X=0.895 $Y=2.67
+ $X2=0.895 $Y2=3.33
r59 40 41 6.39005 $w=7.38e-07 $l=1.65e-07 $layer=LI1_cond $X=0.895 $Y=2.67
+ $X2=0.895 $Y2=2.505
r60 38 51 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r61 38 48 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.16 $Y2=3.33
r62 37 38 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r63 35 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.3 $Y=3.33
+ $X2=2.135 $Y2=3.33
r64 35 37 53.4973 $w=1.68e-07 $l=8.2e-07 $layer=LI1_cond $X=2.3 $Y=3.33 $X2=3.12
+ $Y2=3.33
r65 34 50 4.59886 $w=1.7e-07 $l=2.57e-07 $layer=LI1_cond $X=3.325 $Y=3.33
+ $X2=3.582 $Y2=3.33
r66 34 37 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=3.325 $Y=3.33
+ $X2=3.12 $Y2=3.33
r67 33 44 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.72 $Y2=3.33
r68 32 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r69 30 43 9.68893 $w=1.7e-07 $l=3.7e-07 $layer=LI1_cond $X=1.265 $Y=3.33
+ $X2=0.895 $Y2=3.33
r70 30 32 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=1.265 $Y=3.33
+ $X2=1.68 $Y2=3.33
r71 29 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.97 $Y=3.33
+ $X2=2.135 $Y2=3.33
r72 29 32 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=1.97 $Y=3.33
+ $X2=1.68 $Y2=3.33
r73 27 44 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r74 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r75 24 43 9.68893 $w=1.7e-07 $l=3.7e-07 $layer=LI1_cond $X=0.525 $Y=3.33
+ $X2=0.895 $Y2=3.33
r76 24 26 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.525 $Y=3.33
+ $X2=0.24 $Y2=3.33
r77 22 48 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=2.16 $Y2=3.33
r78 22 33 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=1.68 $Y2=3.33
r79 18 50 3.16731 $w=3.3e-07 $l=1.27609e-07 $layer=LI1_cond $X=3.49 $Y=3.245
+ $X2=3.582 $Y2=3.33
r80 18 20 19.9058 $w=3.28e-07 $l=5.7e-07 $layer=LI1_cond $X=3.49 $Y=3.245
+ $X2=3.49 $Y2=2.675
r81 14 47 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.135 $Y=3.245
+ $X2=2.135 $Y2=3.33
r82 14 16 17.112 $w=3.28e-07 $l=4.9e-07 $layer=LI1_cond $X=2.135 $Y=3.245
+ $X2=2.135 $Y2=2.755
r83 12 41 18.3343 $w=3.28e-07 $l=5.25e-07 $layer=LI1_cond $X=0.69 $Y=1.98
+ $X2=0.69 $Y2=2.505
r84 3 20 600 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_PDIFF $count=1 $X=3.35
+ $Y=2.46 $X2=3.49 $Y2=2.675
r85 2 16 600 $w=1.7e-07 $l=4.10061e-07 $layer=licon1_PDIFF $count=1 $X=1.86
+ $Y=2.46 $X2=2.135 $Y2=2.755
r86 1 40 300 $w=1.7e-07 $l=1.08698e-06 $layer=licon1_PDIFF $count=2 $X=0.55
+ $Y=1.835 $X2=1.13 $Y2=2.67
r87 1 12 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=0.55
+ $Y=1.835 $X2=0.69 $Y2=1.98
.ends

.subckt PM_SKY130_FD_SC_LP__O2BB2A_1%VGND 1 2 9 13 15 17 22 32 33 36 39
r52 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r53 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r54 33 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=3.12
+ $Y2=0
r55 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r56 30 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.265 $Y=0 $X2=3.1
+ $Y2=0
r57 30 32 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=3.265 $Y=0 $X2=3.6
+ $Y2=0
r58 29 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r59 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r60 26 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r61 25 28 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.64
+ $Y2=0
r62 25 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r63 23 36 8.9695 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=0.875 $Y=0 $X2=0.7
+ $Y2=0
r64 23 25 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.875 $Y=0 $X2=1.2
+ $Y2=0
r65 22 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.935 $Y=0 $X2=3.1
+ $Y2=0
r66 22 28 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=2.935 $Y=0 $X2=2.64
+ $Y2=0
r67 20 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r68 19 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r69 17 36 8.9695 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=0.525 $Y=0 $X2=0.7
+ $Y2=0
r70 17 19 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.525 $Y=0 $X2=0.24
+ $Y2=0
r71 15 29 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=2.64
+ $Y2=0
r72 15 26 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=1.2
+ $Y2=0
r73 11 39 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.1 $Y=0.085 $X2=3.1
+ $Y2=0
r74 11 13 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=3.1 $Y=0.085 $X2=3.1
+ $Y2=0.445
r75 7 36 1.07557 $w=3.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.7 $Y=0.085 $X2=0.7
+ $Y2=0
r76 7 9 15.6403 $w=3.48e-07 $l=4.75e-07 $layer=LI1_cond $X=0.7 $Y=0.085 $X2=0.7
+ $Y2=0.56
r77 2 13 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.96
+ $Y=0.235 $X2=3.1 $Y2=0.445
r78 1 9 182 $w=1.7e-07 $l=3.88748e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.235 $X2=0.69 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_LP__O2BB2A_1%A_506_47# 1 2 9 11 12 15
r27 13 15 11.9677 $w=2.58e-07 $l=2.7e-07 $layer=LI1_cond $X=3.565 $Y=0.715
+ $X2=3.565 $Y2=0.445
r28 11 13 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=3.435 $Y=0.8
+ $X2=3.565 $Y2=0.715
r29 11 12 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.435 $Y=0.8
+ $X2=2.765 $Y2=0.8
r30 7 12 6.9898 $w=1.7e-07 $l=1.49579e-07 $layer=LI1_cond $X=2.652 $Y=0.715
+ $X2=2.765 $Y2=0.8
r31 7 9 13.8293 $w=2.23e-07 $l=2.7e-07 $layer=LI1_cond $X=2.652 $Y=0.715
+ $X2=2.652 $Y2=0.445
r32 2 15 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=3.39
+ $Y=0.235 $X2=3.53 $Y2=0.445
r33 1 9 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.53
+ $Y=0.235 $X2=2.67 $Y2=0.445
.ends

