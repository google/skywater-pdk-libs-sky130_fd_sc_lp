* NGSPICE file created from sky130_fd_sc_lp__o41ai_2.ext - technology: sky130A

.subckt sky130_fd_sc_lp__o41ai_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
M1000 a_808_367# A2 a_615_365# VPB phighvt w=1.26e+06u l=150000u
+  ad=1.0206e+12p pd=9.18e+06u as=7.056e+11p ps=6.16e+06u
M1001 VGND A3 a_155_47# VNB nshort w=840000u l=150000u
+  ad=1.1298e+12p pd=9.41e+06u as=1.4028e+12p ps=1.342e+07u
M1002 a_313_365# A4 Y VPB phighvt w=1.26e+06u l=150000u
+  ad=1.3167e+12p pd=9.65e+06u as=7.056e+11p ps=6.16e+06u
M1003 VGND A2 a_155_47# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_808_367# A1 VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=1.0206e+12p ps=9.18e+06u
M1005 a_155_47# A1 VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_615_365# A2 a_808_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 Y B1 a_155_47# VNB nshort w=840000u l=150000u
+  ad=2.352e+11p pd=2.24e+06u as=0p ps=0u
M1008 a_155_47# B1 Y VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR B1 Y VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR A1 a_808_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 Y A4 a_313_365# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_155_47# A2 VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_313_365# A3 a_615_365# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_155_47# A3 VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VGND A4 a_155_47# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_155_47# A4 VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VGND A1 a_155_47# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 Y B1 VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_615_365# A3 a_313_365# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

