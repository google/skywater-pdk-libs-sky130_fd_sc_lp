* File: sky130_fd_sc_lp__bushold0_1.spice
* Created: Wed Sep  2 09:37:40 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__bushold0_1.pex.spice"
.subckt sky130_fd_sc_lp__bushold0_1  VNB VPB X RESET VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* RESET	RESET
* X	X
* VPB	VPB
* VNB	VNB
MM1005 N_VGND_M1005_d N_X_M1005_g N_A_27_535#_M1005_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75001.4
+ A=0.063 P=1.14 MULT=1
MM1000 N_X_M1000_d N_RESET_M1000_g N_VGND_M1005_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6 SB=75001
+ A=0.063 P=1.14 MULT=1
MM1004 N_VGND_M1004_d N_A_27_535#_M1004_g N_X_M1000_d VNB NSHORT L=0.5 W=0.42
+ AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=0.84 SA=250001 SB=250000
+ A=0.21 P=1.84 MULT=1
MM1003 N_VPWR_M1003_d N_X_M1003_g N_A_27_535#_M1003_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.06825 AS=0.2226 PD=0.745 PS=1.9 NRD=21.0987 NRS=124.287 M=1 R=2.8
+ SA=75000.5 SB=75001.4 A=0.063 P=1.14 MULT=1
MM1002 A_258_535# N_RESET_M1002_g N_VPWR_M1003_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0441 AS=0.06825 PD=0.63 PS=0.745 NRD=23.443 NRS=0 M=1 R=2.8 SA=75000.9
+ SB=75000.9 A=0.063 P=1.14 MULT=1
MM1001 N_X_M1001_d N_A_27_535#_M1001_g A_258_535# VPB PHIGHVT L=0.5 W=0.42
+ AD=0.1113 AS=0.0441 PD=1.37 PS=0.63 NRD=0 NRS=23.443 M=1 R=0.84 SA=250001
+ SB=250000 A=0.21 P=1.84 MULT=1
DX6_noxref VNB VPB NWDIODE A=5.1847 P=9.29
*
.include "sky130_fd_sc_lp__bushold0_1.pxi.spice"
*
.ends
*
*
