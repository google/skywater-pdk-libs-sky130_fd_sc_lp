* File: sky130_fd_sc_lp__o22a_m.pex.spice
* Created: Wed Sep  2 10:20:19 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O22A_M%A_88_187# 1 2 8 11 15 16 20 21 22 23 24 25 28
+ 31 36
c80 22 0 9.68398e-20 $X=1.67 $Y=0.9
c81 11 0 7.49253e-20 $X=0.515 $Y=2.885
r82 31 33 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=1.835 $Y=0.7 $X2=1.835
+ $Y2=0.9
r83 26 28 6.07359 $w=2.08e-07 $l=1.15e-07 $layer=LI1_cond $X=2.195 $Y=2.705
+ $X2=2.195 $Y2=2.82
r84 24 26 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=2.09 $Y=2.62
+ $X2=2.195 $Y2=2.705
r85 24 25 89.7059 $w=1.68e-07 $l=1.375e-06 $layer=LI1_cond $X=2.09 $Y=2.62
+ $X2=0.715 $Y2=2.62
r86 22 33 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.67 $Y=0.9
+ $X2=1.835 $Y2=0.9
r87 22 23 62.3048 $w=1.68e-07 $l=9.55e-07 $layer=LI1_cond $X=1.67 $Y=0.9
+ $X2=0.715 $Y2=0.9
r88 21 36 46.504 $w=3.55e-07 $l=1.65e-07 $layer=POLY_cond $X=0.617 $Y=1.1
+ $X2=0.617 $Y2=0.935
r89 20 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.63 $Y=1.1
+ $X2=0.63 $Y2=1.1
r90 18 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.63 $Y=2.535
+ $X2=0.715 $Y2=2.62
r91 18 20 93.6203 $w=1.68e-07 $l=1.435e-06 $layer=LI1_cond $X=0.63 $Y=2.535
+ $X2=0.63 $Y2=1.1
r92 17 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.63 $Y=0.985
+ $X2=0.715 $Y2=0.9
r93 17 20 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=0.63 $Y=0.985
+ $X2=0.63 $Y2=1.1
r94 15 36 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.54 $Y=0.615
+ $X2=0.54 $Y2=0.935
r95 11 16 656.34 $w=1.5e-07 $l=1.28e-06 $layer=POLY_cond $X=0.515 $Y=2.885
+ $X2=0.515 $Y2=1.605
r96 8 16 48.4546 $w=3.55e-07 $l=1.77e-07 $layer=POLY_cond $X=0.617 $Y=1.428
+ $X2=0.617 $Y2=1.605
r97 7 21 1.95057 $w=3.55e-07 $l=1.2e-08 $layer=POLY_cond $X=0.617 $Y=1.112
+ $X2=0.617 $Y2=1.1
r98 7 8 51.3649 $w=3.55e-07 $l=3.16e-07 $layer=POLY_cond $X=0.617 $Y=1.112
+ $X2=0.617 $Y2=1.428
r99 2 28 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.055
+ $Y=2.675 $X2=2.195 $Y2=2.82
r100 1 31 182 $w=1.7e-07 $l=3.58225e-07 $layer=licon1_NDIFF $count=1 $X=1.695
+ $Y=0.405 $X2=1.835 $Y2=0.7
.ends

.subckt PM_SKY130_FD_SC_LP__O22A_M%A1 3 7 12 13 16 17 21 22 23 31
c57 16 0 7.49253e-20 $X=1.17 $Y=1.25
c58 3 0 1.00575e-19 $X=1.11 $Y=0.615
r59 31 32 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.97
+ $Y=1.82 $X2=2.97 $Y2=1.82
r60 22 23 13.3251 $w=3.18e-07 $l=3.7e-07 $layer=LI1_cond $X=3.045 $Y=2.035
+ $X2=3.045 $Y2=2.405
r61 22 32 7.74298 $w=3.18e-07 $l=2.15e-07 $layer=LI1_cond $X=3.045 $Y=2.035
+ $X2=3.045 $Y2=1.82
r62 21 32 4.06956 $w=3.18e-07 $l=1.13e-07 $layer=LI1_cond $X=3.045 $Y=1.707
+ $X2=3.045 $Y2=1.82
r63 16 19 11.5244 $w=3.28e-07 $l=3.3e-07 $layer=LI1_cond $X=1.17 $Y=1.25
+ $X2=1.17 $Y2=1.58
r64 16 17 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.17
+ $Y=1.25 $X2=1.17 $Y2=1.25
r65 14 19 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.335 $Y=1.58
+ $X2=1.17 $Y2=1.58
r66 13 21 5.01689 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=2.885 $Y=1.58
+ $X2=3.045 $Y2=1.58
r67 13 14 101.123 $w=1.68e-07 $l=1.55e-06 $layer=LI1_cond $X=2.885 $Y=1.58
+ $X2=1.335 $Y2=1.58
r68 11 31 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.97 $Y=2.16
+ $X2=2.97 $Y2=1.82
r69 11 12 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.97 $Y=2.16
+ $X2=2.97 $Y2=2.325
r70 10 17 41.8716 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.17 $Y=1.085
+ $X2=1.17 $Y2=1.25
r71 7 12 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=2.88 $Y=2.885
+ $X2=2.88 $Y2=2.325
r72 3 10 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=1.11 $Y=0.615 $X2=1.11
+ $Y2=1.085
.ends

.subckt PM_SKY130_FD_SC_LP__O22A_M%B1 3 7 9 10 11
c38 11 0 1.64512e-19 $X=1.2 $Y=2.035
r39 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.2
+ $Y=2.16 $X2=1.2 $Y2=2.16
r40 11 15 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=1.2 $Y=2.035
+ $X2=1.2 $Y2=2.16
r41 9 14 60.3271 $w=3.3e-07 $l=3.45e-07 $layer=POLY_cond $X=1.545 $Y=2.16
+ $X2=1.2 $Y2=2.16
r42 9 10 5.03009 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=1.545 $Y=2.16
+ $X2=1.62 $Y2=2.16
r43 5 10 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.62 $Y=2.325
+ $X2=1.62 $Y2=2.16
r44 5 7 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=1.62 $Y=2.325 $X2=1.62
+ $Y2=2.885
r45 1 10 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.62 $Y=1.995
+ $X2=1.62 $Y2=2.16
r46 1 3 707.617 $w=1.5e-07 $l=1.38e-06 $layer=POLY_cond $X=1.62 $Y=1.995
+ $X2=1.62 $Y2=0.615
.ends

.subckt PM_SKY130_FD_SC_LP__O22A_M%B2 3 7 11 12 13 14 18
c34 11 0 1.64512e-19 $X=2.07 $Y=2.27
c35 7 0 9.68398e-20 $X=2.05 $Y=0.615
r36 18 19 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.07
+ $Y=1.93 $X2=2.07 $Y2=1.93
r37 14 19 2.11073 $w=5.08e-07 $l=9e-08 $layer=LI1_cond $X=2.16 $Y=2.1 $X2=2.07
+ $Y2=2.1
r38 13 19 9.14648 $w=5.08e-07 $l=3.9e-07 $layer=LI1_cond $X=1.68 $Y=2.1 $X2=2.07
+ $Y2=2.1
r39 11 18 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.07 $Y=2.27
+ $X2=2.07 $Y2=1.93
r40 11 12 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.07 $Y=2.27
+ $X2=2.07 $Y2=2.435
r41 10 18 38.6168 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.07 $Y=1.765
+ $X2=2.07 $Y2=1.93
r42 7 10 589.681 $w=1.5e-07 $l=1.15e-06 $layer=POLY_cond $X=2.05 $Y=0.615
+ $X2=2.05 $Y2=1.765
r43 3 12 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=1.98 $Y=2.885
+ $X2=1.98 $Y2=2.435
.ends

.subckt PM_SKY130_FD_SC_LP__O22A_M%A2 1 3 5 7 8 9
c34 5 0 1.00575e-19 $X=2.56 $Y=0.935
r35 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.65
+ $Y=1.1 $X2=2.65 $Y2=1.1
r36 9 14 15.6999 $w=3.43e-07 $l=4.7e-07 $layer=LI1_cond $X=3.12 $Y=1.012
+ $X2=2.65 $Y2=1.012
r37 8 14 0.334041 $w=3.43e-07 $l=1e-08 $layer=LI1_cond $X=2.64 $Y=1.012 $X2=2.65
+ $Y2=1.012
r38 5 13 38.7595 $w=2.78e-07 $l=1.96914e-07 $layer=POLY_cond $X=2.56 $Y=0.935
+ $X2=2.63 $Y2=1.1
r39 5 7 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.56 $Y=0.935 $X2=2.56
+ $Y2=0.615
r40 1 13 69.9681 $w=2.78e-07 $l=3.96201e-07 $layer=POLY_cond $X=2.52 $Y=1.445
+ $X2=2.63 $Y2=1.1
r41 1 3 738.383 $w=1.5e-07 $l=1.44e-06 $layer=POLY_cond $X=2.52 $Y=1.445
+ $X2=2.52 $Y2=2.885
.ends

.subckt PM_SKY130_FD_SC_LP__O22A_M%X 1 2 9 12 13 14 15 16 17
r15 16 17 18.9513 $w=2.23e-07 $l=3.7e-07 $layer=LI1_cond $X=0.252 $Y=2.405
+ $X2=0.252 $Y2=2.775
r16 15 16 18.9513 $w=2.23e-07 $l=3.7e-07 $layer=LI1_cond $X=0.252 $Y=2.035
+ $X2=0.252 $Y2=2.405
r17 14 15 18.9513 $w=2.23e-07 $l=3.7e-07 $layer=LI1_cond $X=0.252 $Y=1.665
+ $X2=0.252 $Y2=2.035
r18 13 14 18.9513 $w=2.23e-07 $l=3.7e-07 $layer=LI1_cond $X=0.252 $Y=1.295
+ $X2=0.252 $Y2=1.665
r19 12 13 18.9513 $w=2.23e-07 $l=3.7e-07 $layer=LI1_cond $X=0.252 $Y=0.925
+ $X2=0.252 $Y2=1.295
r20 11 12 14.8537 $w=2.23e-07 $l=2.9e-07 $layer=LI1_cond $X=0.252 $Y=0.635
+ $X2=0.252 $Y2=0.925
r21 9 11 4.14275 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=0.305 $Y=0.55
+ $X2=0.305 $Y2=0.635
r22 2 17 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.155
+ $Y=2.675 $X2=0.28 $Y2=2.82
r23 1 9 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.18
+ $Y=0.405 $X2=0.305 $Y2=0.55
.ends

.subckt PM_SKY130_FD_SC_LP__O22A_M%VPWR 1 2 9 11 13 15 17 22 31 35
r43 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r44 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r45 29 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r46 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r47 26 32 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r48 25 28 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r49 25 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r50 23 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.895 $Y=3.33
+ $X2=0.73 $Y2=3.33
r51 23 25 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.895 $Y=3.33
+ $X2=1.2 $Y2=3.33
r52 22 34 4.77065 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=2.93 $Y=3.33
+ $X2=3.145 $Y2=3.33
r53 22 28 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=2.93 $Y=3.33
+ $X2=2.64 $Y2=3.33
r54 20 32 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r55 19 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r56 17 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.565 $Y=3.33
+ $X2=0.73 $Y2=3.33
r57 17 19 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.565 $Y=3.33
+ $X2=0.24 $Y2=3.33
r58 15 29 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r59 15 26 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r60 11 34 2.99552 $w=3.3e-07 $l=1.07121e-07 $layer=LI1_cond $X=3.095 $Y=3.245
+ $X2=3.145 $Y2=3.33
r61 11 13 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=3.095 $Y=3.245
+ $X2=3.095 $Y2=2.95
r62 7 31 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=3.245 $X2=0.73
+ $Y2=3.33
r63 7 9 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=0.73 $Y=3.245
+ $X2=0.73 $Y2=2.97
r64 2 13 600 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=1 $X=2.955
+ $Y=2.675 $X2=3.095 $Y2=2.95
r65 1 9 600 $w=1.7e-07 $l=3.58225e-07 $layer=licon1_PDIFF $count=1 $X=0.59
+ $Y=2.675 $X2=0.73 $Y2=2.97
.ends

.subckt PM_SKY130_FD_SC_LP__O22A_M%VGND 1 2 11 15 18 19 20 30 31 34
r38 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r39 30 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r40 28 31 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r41 27 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r42 25 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r43 24 27 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.64
+ $Y2=0
r44 24 25 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r45 22 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.98 $Y=0 $X2=0.815
+ $Y2=0
r46 22 24 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=0.98 $Y=0 $X2=1.2
+ $Y2=0
r47 20 28 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r48 20 25 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r49 18 27 3.26203 $w=1.68e-07 $l=5e-08 $layer=LI1_cond $X=2.69 $Y=0 $X2=2.64
+ $Y2=0
r50 18 19 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.69 $Y=0 $X2=2.855
+ $Y2=0
r51 17 30 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=3.02 $Y=0 $X2=3.12
+ $Y2=0
r52 17 19 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.02 $Y=0 $X2=2.855
+ $Y2=0
r53 13 19 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.855 $Y=0.085
+ $X2=2.855 $Y2=0
r54 13 15 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=2.855 $Y=0.085
+ $X2=2.855 $Y2=0.55
r55 9 34 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.815 $Y=0.085
+ $X2=0.815 $Y2=0
r56 9 11 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=0.815 $Y=0.085
+ $X2=0.815 $Y2=0.53
r57 2 15 182 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_NDIFF $count=1 $X=2.635
+ $Y=0.405 $X2=2.855 $Y2=0.55
r58 1 11 182 $w=1.7e-07 $l=2.54951e-07 $layer=licon1_NDIFF $count=1 $X=0.615
+ $Y=0.405 $X2=0.815 $Y2=0.53
.ends

.subckt PM_SKY130_FD_SC_LP__O22A_M%A_237_81# 1 2 7 9 14
c23 7 0 2.01149e-19 $X=2.18 $Y=0.35
r24 14 17 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=2.345 $Y=0.35 $X2=2.345
+ $Y2=0.55
r25 9 12 6.28605 $w=3.28e-07 $l=1.8e-07 $layer=LI1_cond $X=1.325 $Y=0.35
+ $X2=1.325 $Y2=0.53
r26 8 9 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.49 $Y=0.35 $X2=1.325
+ $Y2=0.35
r27 7 14 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.18 $Y=0.35
+ $X2=2.345 $Y2=0.35
r28 7 8 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.18 $Y=0.35 $X2=1.49
+ $Y2=0.35
r29 2 17 182 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_NDIFF $count=1 $X=2.125
+ $Y=0.405 $X2=2.345 $Y2=0.55
r30 1 12 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=1.185
+ $Y=0.405 $X2=1.325 $Y2=0.53
.ends

