* File: sky130_fd_sc_lp__o22ai_0.spice
* Created: Fri Aug 28 11:10:22 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__o22ai_0.pex.spice"
.subckt sky130_fd_sc_lp__o22ai_0  VNB VPB B1 B2 A2 A1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A1	A1
* A2	A2
* B2	B2
* B1	B1
* VPB	VPB
* VNB	VNB
MM1004 N_Y_M1004_d N_B1_M1004_g N_A_27_85#_M1004_s VNB NSHORT L=0.15 W=0.42
+ AD=0.07455 AS=0.1218 PD=0.775 PS=1.42 NRD=21.42 NRS=1.428 M=1 R=2.8 SA=75000.2
+ SB=75001.6 A=0.063 P=1.14 MULT=1
MM1007 N_A_27_85#_M1007_d N_B2_M1007_g N_Y_M1004_d VNB NSHORT L=0.15 W=0.42
+ AD=0.06405 AS=0.07455 PD=0.725 PS=0.775 NRD=5.712 NRS=0 M=1 R=2.8 SA=75000.7
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1005 N_VGND_M1005_d N_A2_M1005_g N_A_27_85#_M1007_d VNB NSHORT L=0.15 W=0.42
+ AD=0.06615 AS=0.06405 PD=0.735 PS=0.725 NRD=4.284 NRS=1.428 M=1 R=2.8
+ SA=75001.2 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1006 N_A_27_85#_M1006_d N_A1_M1006_g N_VGND_M1005_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.06615 PD=1.37 PS=0.735 NRD=0 NRS=5.712 M=1 R=2.8 SA=75001.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1001 A_143_483# N_B1_M1001_g N_VPWR_M1001_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0768 AS=0.256 PD=0.88 PS=2.08 NRD=19.9955 NRS=20.7638 M=1 R=4.26667
+ SA=75000.3 SB=75001.4 A=0.096 P=1.58 MULT=1
MM1002 N_Y_M1002_d N_B2_M1002_g A_143_483# VPB PHIGHVT L=0.15 W=0.64 AD=0.0896
+ AS=0.0768 PD=0.92 PS=0.88 NRD=0 NRS=19.9955 M=1 R=4.26667 SA=75000.7 SB=75001
+ A=0.096 P=1.58 MULT=1
MM1000 A_307_483# N_A2_M1000_g N_Y_M1002_d VPB PHIGHVT L=0.15 W=0.64 AD=0.0768
+ AS=0.0896 PD=0.88 PS=0.92 NRD=19.9955 NRS=0 M=1 R=4.26667 SA=75001.1
+ SB=75000.6 A=0.096 P=1.58 MULT=1
MM1003 N_VPWR_M1003_d N_A1_M1003_g A_307_483# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1696 AS=0.0768 PD=1.81 PS=0.88 NRD=0 NRS=19.9955 M=1 R=4.26667 SA=75001.5
+ SB=75000.2 A=0.096 P=1.58 MULT=1
DX8_noxref VNB VPB NWDIODE A=5.1847 P=9.29
c_276 A_307_483# 0 1.06273e-19 $X=1.535 $Y=2.415
*
.include "sky130_fd_sc_lp__o22ai_0.pxi.spice"
*
.ends
*
*
