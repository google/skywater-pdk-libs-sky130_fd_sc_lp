* File: sky130_fd_sc_lp__o21bai_lp.pxi.spice
* Created: Wed Sep  2 10:17:51 2020
* 
x_PM_SKY130_FD_SC_LP__O21BAI_LP%A1 N_A1_c_61_n N_A1_M1003_g N_A1_M1002_g
+ N_A1_c_62_n N_A1_c_66_n A1 A1 N_A1_c_63_n N_A1_c_64_n
+ PM_SKY130_FD_SC_LP__O21BAI_LP%A1
x_PM_SKY130_FD_SC_LP__O21BAI_LP%A2 N_A2_M1000_g N_A2_M1006_g A2 A2 N_A2_c_92_n
+ N_A2_c_93_n N_A2_c_94_n PM_SKY130_FD_SC_LP__O21BAI_LP%A2
x_PM_SKY130_FD_SC_LP__O21BAI_LP%A_288_21# N_A_288_21#_M1008_d
+ N_A_288_21#_M1001_d N_A_288_21#_c_131_n N_A_288_21#_M1004_g
+ N_A_288_21#_M1005_g N_A_288_21#_c_133_n N_A_288_21#_c_140_n
+ N_A_288_21#_c_134_n N_A_288_21#_c_135_n N_A_288_21#_c_136_n
+ N_A_288_21#_c_137_n N_A_288_21#_c_138_n
+ PM_SKY130_FD_SC_LP__O21BAI_LP%A_288_21#
x_PM_SKY130_FD_SC_LP__O21BAI_LP%B1_N N_B1_N_c_207_n N_B1_N_M1001_g
+ N_B1_N_M1007_g N_B1_N_c_208_n N_B1_N_c_209_n N_B1_N_c_201_n N_B1_N_M1008_g
+ N_B1_N_c_203_n N_B1_N_c_204_n B1_N N_B1_N_c_206_n
+ PM_SKY130_FD_SC_LP__O21BAI_LP%B1_N
x_PM_SKY130_FD_SC_LP__O21BAI_LP%VPWR N_VPWR_M1002_s N_VPWR_M1005_d
+ N_VPWR_c_255_n N_VPWR_c_256_n N_VPWR_c_257_n VPWR N_VPWR_c_258_n
+ N_VPWR_c_259_n N_VPWR_c_254_n N_VPWR_c_261_n
+ PM_SKY130_FD_SC_LP__O21BAI_LP%VPWR
x_PM_SKY130_FD_SC_LP__O21BAI_LP%Y N_Y_M1004_d N_Y_M1000_d N_Y_c_303_n
+ N_Y_c_290_n N_Y_c_292_n Y Y PM_SKY130_FD_SC_LP__O21BAI_LP%Y
x_PM_SKY130_FD_SC_LP__O21BAI_LP%A_28_110# N_A_28_110#_M1003_s
+ N_A_28_110#_M1006_d N_A_28_110#_c_336_n N_A_28_110#_c_337_n
+ N_A_28_110#_c_338_n PM_SKY130_FD_SC_LP__O21BAI_LP%A_28_110#
x_PM_SKY130_FD_SC_LP__O21BAI_LP%VGND N_VGND_M1003_d N_VGND_M1007_s
+ N_VGND_c_359_n N_VGND_c_360_n VGND N_VGND_c_361_n N_VGND_c_362_n
+ N_VGND_c_363_n N_VGND_c_364_n N_VGND_c_365_n N_VGND_c_366_n
+ PM_SKY130_FD_SC_LP__O21BAI_LP%VGND
cc_1 VNB N_A1_c_61_n 0.0641406f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=1.27
cc_2 VNB N_A1_c_62_n 0.00370103f $X=-0.19 $Y=-0.245 $X2=0.547 $Y2=1.84
cc_3 VNB N_A1_c_63_n 0.00483634f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.435
cc_4 VNB N_A1_c_64_n 0.0548803f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=1.435
cc_5 VNB N_A2_M1000_g 0.00298717f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=1.27
cc_6 VNB N_A2_c_92_n 0.0308885f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.435
cc_7 VNB N_A2_c_93_n 0.0104363f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A2_c_94_n 0.0461308f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=1.435
cc_9 VNB N_A_288_21#_c_131_n 0.0557027f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=2.565
cc_10 VNB N_A_288_21#_M1005_g 0.0106682f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.95
cc_11 VNB N_A_288_21#_c_133_n 0.0112909f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.435
cc_12 VNB N_A_288_21#_c_134_n 0.0277776f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=1.665
cc_13 VNB N_A_288_21#_c_135_n 0.0258453f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_288_21#_c_136_n 0.0181241f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_288_21#_c_137_n 0.0121093f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_288_21#_c_138_n 0.0561221f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_B1_N_M1007_g 0.0199771f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=1.99
cc_18 VNB N_B1_N_c_201_n 0.00671477f $X=-0.19 $Y=-0.245 $X2=0.547 $Y2=1.99
cc_19 VNB N_B1_N_M1008_g 0.0277118f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_B1_N_c_203_n 0.035923f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.435
cc_21 VNB N_B1_N_c_204_n 0.0228961f $X=-0.19 $Y=-0.245 $X2=0.485 $Y2=1.435
cc_22 VNB B1_N 0.00907485f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_B1_N_c_206_n 0.0316621f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=1.665
cc_24 VNB N_VPWR_c_254_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_Y_c_290_n 0.0193472f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB Y 0.00544117f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_28_110#_c_336_n 0.00438843f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=2.565
cc_28 VNB N_A_28_110#_c_337_n 0.0215136f $X=-0.19 $Y=-0.245 $X2=0.547 $Y2=1.99
cc_29 VNB N_A_28_110#_c_338_n 0.00637255f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.435
cc_30 VNB N_VGND_c_359_n 0.0156825f $X=-0.19 $Y=-0.245 $X2=0.547 $Y2=1.84
cc_31 VNB N_VGND_c_360_n 0.00916183f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_361_n 0.0208004f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.435
cc_33 VNB N_VGND_c_362_n 0.0341047f $X=-0.19 $Y=-0.245 $X2=0.28 $Y2=1.435
cc_34 VNB N_VGND_c_363_n 0.0270417f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_364_n 0.214242f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_365_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_366_n 0.00510915f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VPB N_A1_c_62_n 0.0126109f $X=-0.19 $Y=1.655 $X2=0.547 $Y2=1.84
cc_39 VPB N_A1_c_66_n 0.0379886f $X=-0.19 $Y=1.655 $X2=0.547 $Y2=1.99
cc_40 VPB N_A1_c_63_n 0.0204072f $X=-0.19 $Y=1.655 $X2=0.29 $Y2=1.435
cc_41 VPB N_A2_M1000_g 0.0368089f $X=-0.19 $Y=1.655 $X2=0.5 $Y2=1.27
cc_42 VPB N_A2_c_93_n 0.00420665f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_43 VPB N_A_288_21#_M1005_g 0.0452096f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.95
cc_44 VPB N_A_288_21#_c_140_n 0.0211635f $X=-0.19 $Y=1.655 $X2=0.485 $Y2=1.435
cc_45 VPB N_A_288_21#_c_135_n 0.0091103f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_46 VPB N_A_288_21#_c_136_n 0.0115533f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_47 VPB N_B1_N_c_207_n 0.0212316f $X=-0.19 $Y=1.655 $X2=0.485 $Y2=1.6
cc_48 VPB N_B1_N_c_208_n 0.0514531f $X=-0.19 $Y=1.655 $X2=0.575 $Y2=2.565
cc_49 VPB N_B1_N_c_209_n 0.0162002f $X=-0.19 $Y=1.655 $X2=0.547 $Y2=1.84
cc_50 VPB N_B1_N_c_203_n 0.123685f $X=-0.19 $Y=1.655 $X2=0.29 $Y2=1.435
cc_51 VPB N_VPWR_c_255_n 0.0121621f $X=-0.19 $Y=1.655 $X2=0.575 $Y2=2.565
cc_52 VPB N_VPWR_c_256_n 0.0330902f $X=-0.19 $Y=1.655 $X2=0.547 $Y2=1.84
cc_53 VPB N_VPWR_c_257_n 0.00443446f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_54 VPB N_VPWR_c_258_n 0.03308f $X=-0.19 $Y=1.655 $X2=0.29 $Y2=1.435
cc_55 VPB N_VPWR_c_259_n 0.0428092f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_56 VPB N_VPWR_c_254_n 0.0625539f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_57 VPB N_VPWR_c_261_n 0.00533588f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_58 VPB N_Y_c_292_n 0.0012299f $X=-0.19 $Y=1.655 $X2=0.29 $Y2=1.435
cc_59 VPB Y 0.00338806f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_60 VPB Y 0.00114455f $X=-0.19 $Y=1.655 $X2=0.485 $Y2=1.435
cc_61 N_A1_c_62_n N_A2_M1000_g 0.00755557f $X=0.547 $Y=1.84 $X2=0 $Y2=0
cc_62 N_A1_c_66_n N_A2_M1000_g 0.0883737f $X=0.547 $Y=1.99 $X2=0 $Y2=0
cc_63 N_A1_c_63_n N_A2_M1000_g 2.39932e-19 $X=0.29 $Y=1.435 $X2=0 $Y2=0
cc_64 N_A1_c_63_n N_A2_c_92_n 2.39968e-19 $X=0.29 $Y=1.435 $X2=0 $Y2=0
cc_65 N_A1_c_64_n N_A2_c_92_n 0.020826f $X=0.5 $Y=1.435 $X2=0 $Y2=0
cc_66 N_A1_c_66_n N_A2_c_93_n 0.0159586f $X=0.547 $Y=1.99 $X2=0 $Y2=0
cc_67 N_A1_c_63_n N_A2_c_93_n 0.06897f $X=0.29 $Y=1.435 $X2=0 $Y2=0
cc_68 N_A1_c_64_n N_A2_c_93_n 0.00505842f $X=0.5 $Y=1.435 $X2=0 $Y2=0
cc_69 N_A1_c_61_n N_A2_c_94_n 0.0274576f $X=0.5 $Y=1.27 $X2=0 $Y2=0
cc_70 N_A1_c_63_n N_VPWR_M1002_s 0.00273067f $X=0.29 $Y=1.435 $X2=-0.19
+ $Y2=-0.245
cc_71 N_A1_c_66_n N_VPWR_c_256_n 0.0244465f $X=0.547 $Y=1.99 $X2=0 $Y2=0
cc_72 N_A1_c_63_n N_VPWR_c_256_n 0.0223371f $X=0.29 $Y=1.435 $X2=0 $Y2=0
cc_73 N_A1_c_66_n N_VPWR_c_258_n 0.00831182f $X=0.547 $Y=1.99 $X2=0 $Y2=0
cc_74 N_A1_c_66_n N_VPWR_c_254_n 0.0142754f $X=0.547 $Y=1.99 $X2=0 $Y2=0
cc_75 N_A1_c_66_n N_Y_c_292_n 0.00198508f $X=0.547 $Y=1.99 $X2=0 $Y2=0
cc_76 N_A1_c_61_n N_A_28_110#_c_336_n 0.0162799f $X=0.5 $Y=1.27 $X2=0 $Y2=0
cc_77 N_A1_c_61_n N_A_28_110#_c_337_n 0.0101824f $X=0.5 $Y=1.27 $X2=0 $Y2=0
cc_78 N_A1_c_63_n N_A_28_110#_c_337_n 0.0267483f $X=0.29 $Y=1.435 $X2=0 $Y2=0
cc_79 N_A1_c_64_n N_A_28_110#_c_337_n 0.00228944f $X=0.5 $Y=1.435 $X2=0 $Y2=0
cc_80 N_A1_c_61_n N_A_28_110#_c_338_n 8.81474e-19 $X=0.5 $Y=1.27 $X2=0 $Y2=0
cc_81 N_A1_c_61_n N_VGND_c_359_n 0.0151037f $X=0.5 $Y=1.27 $X2=0 $Y2=0
cc_82 N_A1_c_61_n N_VGND_c_361_n 0.00558995f $X=0.5 $Y=1.27 $X2=0 $Y2=0
cc_83 N_A1_c_61_n N_VGND_c_364_n 0.0114789f $X=0.5 $Y=1.27 $X2=0 $Y2=0
cc_84 N_A2_c_93_n N_A_288_21#_c_131_n 0.00894383f $X=0.95 $Y=1.435 $X2=0 $Y2=0
cc_85 N_A2_c_94_n N_A_288_21#_c_131_n 0.0293873f $X=0.972 $Y=1.27 $X2=0 $Y2=0
cc_86 N_A2_M1000_g N_A_288_21#_M1005_g 0.0293873f $X=1.035 $Y=2.565 $X2=0 $Y2=0
cc_87 N_A2_c_92_n N_A_288_21#_c_133_n 0.0293873f $X=0.95 $Y=1.435 $X2=0 $Y2=0
cc_88 N_A2_M1000_g N_VPWR_c_256_n 0.00284782f $X=1.035 $Y=2.565 $X2=0 $Y2=0
cc_89 N_A2_M1000_g N_VPWR_c_257_n 9.08728e-19 $X=1.035 $Y=2.565 $X2=0 $Y2=0
cc_90 N_A2_M1000_g N_VPWR_c_258_n 0.00890977f $X=1.035 $Y=2.565 $X2=0 $Y2=0
cc_91 N_A2_M1000_g N_VPWR_c_254_n 0.0158598f $X=1.035 $Y=2.565 $X2=0 $Y2=0
cc_92 N_A2_c_93_n A_140_413# 0.00433061f $X=0.95 $Y=1.435 $X2=-0.19 $Y2=-0.245
cc_93 N_A2_c_93_n N_Y_M1000_d 0.00192361f $X=0.95 $Y=1.435 $X2=0 $Y2=0
cc_94 N_A2_c_92_n N_Y_c_290_n 3.04604e-19 $X=0.95 $Y=1.435 $X2=0 $Y2=0
cc_95 N_A2_c_93_n N_Y_c_290_n 0.0460593f $X=0.95 $Y=1.435 $X2=0 $Y2=0
cc_96 N_A2_M1000_g N_Y_c_292_n 0.0171087f $X=1.035 $Y=2.565 $X2=0 $Y2=0
cc_97 N_A2_c_93_n N_Y_c_292_n 0.0108196f $X=0.95 $Y=1.435 $X2=0 $Y2=0
cc_98 N_A2_M1000_g Y 3.04604e-19 $X=1.035 $Y=2.565 $X2=0 $Y2=0
cc_99 N_A2_M1000_g Y 6.85028e-19 $X=1.035 $Y=2.565 $X2=0 $Y2=0
cc_100 N_A2_c_92_n N_A_28_110#_c_336_n 0.00157672f $X=0.95 $Y=1.435 $X2=0 $Y2=0
cc_101 N_A2_c_93_n N_A_28_110#_c_336_n 0.0426214f $X=0.95 $Y=1.435 $X2=0 $Y2=0
cc_102 N_A2_c_94_n N_A_28_110#_c_336_n 0.0124254f $X=0.972 $Y=1.27 $X2=0 $Y2=0
cc_103 N_A2_c_94_n N_A_28_110#_c_337_n 8.83935e-19 $X=0.972 $Y=1.27 $X2=0 $Y2=0
cc_104 N_A2_c_93_n N_A_28_110#_c_338_n 0.0160768f $X=0.95 $Y=1.435 $X2=0 $Y2=0
cc_105 N_A2_c_94_n N_A_28_110#_c_338_n 0.00843905f $X=0.972 $Y=1.27 $X2=0 $Y2=0
cc_106 N_A2_c_94_n N_VGND_c_359_n 0.0136f $X=0.972 $Y=1.27 $X2=0 $Y2=0
cc_107 N_A2_c_94_n N_VGND_c_362_n 0.00558995f $X=0.972 $Y=1.27 $X2=0 $Y2=0
cc_108 N_A2_c_94_n N_VGND_c_364_n 0.0104363f $X=0.972 $Y=1.27 $X2=0 $Y2=0
cc_109 N_A_288_21#_M1005_g N_B1_N_c_207_n 0.0213578f $X=1.565 $Y=2.565 $X2=-0.19
+ $Y2=-0.245
cc_110 N_A_288_21#_c_140_n N_B1_N_c_207_n 0.0282709f $X=2.62 $Y=2.145 $X2=-0.19
+ $Y2=-0.245
cc_111 N_A_288_21#_c_135_n N_B1_N_c_207_n 0.0016425f $X=2.62 $Y=1.495 $X2=-0.19
+ $Y2=-0.245
cc_112 N_A_288_21#_c_138_n N_B1_N_c_207_n 0.0095366f $X=2.455 $Y=1.495 $X2=-0.19
+ $Y2=-0.245
cc_113 N_A_288_21#_c_137_n N_B1_N_M1007_g 8.57376e-19 $X=3.08 $Y=0.41 $X2=0
+ $Y2=0
cc_114 N_A_288_21#_c_140_n N_B1_N_c_208_n 0.00516985f $X=2.62 $Y=2.145 $X2=0
+ $Y2=0
cc_115 N_A_288_21#_c_135_n N_B1_N_c_201_n 0.011146f $X=2.62 $Y=1.495 $X2=0 $Y2=0
cc_116 N_A_288_21#_c_136_n N_B1_N_c_201_n 0.00971735f $X=3.16 $Y=1.495 $X2=0
+ $Y2=0
cc_117 N_A_288_21#_c_134_n N_B1_N_M1008_g 0.00963308f $X=3.16 $Y=1.33 $X2=0
+ $Y2=0
cc_118 N_A_288_21#_c_137_n N_B1_N_M1008_g 0.0064251f $X=3.08 $Y=0.41 $X2=0 $Y2=0
cc_119 N_A_288_21#_c_140_n N_B1_N_c_203_n 0.0338914f $X=2.62 $Y=2.145 $X2=0
+ $Y2=0
cc_120 N_A_288_21#_c_134_n N_B1_N_c_203_n 0.0150165f $X=3.16 $Y=1.33 $X2=0 $Y2=0
cc_121 N_A_288_21#_c_135_n N_B1_N_c_203_n 0.0181258f $X=2.62 $Y=1.495 $X2=0
+ $Y2=0
cc_122 N_A_288_21#_c_136_n N_B1_N_c_203_n 0.0226838f $X=3.16 $Y=1.495 $X2=0
+ $Y2=0
cc_123 N_A_288_21#_c_134_n N_B1_N_c_204_n 0.00894354f $X=3.16 $Y=1.33 $X2=0
+ $Y2=0
cc_124 N_A_288_21#_c_137_n N_B1_N_c_204_n 0.00355012f $X=3.08 $Y=0.41 $X2=0
+ $Y2=0
cc_125 N_A_288_21#_c_134_n B1_N 0.0159955f $X=3.16 $Y=1.33 $X2=0 $Y2=0
cc_126 N_A_288_21#_c_135_n B1_N 0.00150048f $X=2.62 $Y=1.495 $X2=0 $Y2=0
cc_127 N_A_288_21#_c_136_n B1_N 0.0197467f $X=3.16 $Y=1.495 $X2=0 $Y2=0
cc_128 N_A_288_21#_c_138_n B1_N 0.00125691f $X=2.455 $Y=1.495 $X2=0 $Y2=0
cc_129 N_A_288_21#_c_131_n N_B1_N_c_206_n 0.00259672f $X=1.515 $Y=1.36 $X2=0
+ $Y2=0
cc_130 N_A_288_21#_c_135_n N_B1_N_c_206_n 0.00809447f $X=2.62 $Y=1.495 $X2=0
+ $Y2=0
cc_131 N_A_288_21#_c_136_n N_B1_N_c_206_n 5.04688e-19 $X=3.16 $Y=1.495 $X2=0
+ $Y2=0
cc_132 N_A_288_21#_c_138_n N_B1_N_c_206_n 0.0114175f $X=2.455 $Y=1.495 $X2=0
+ $Y2=0
cc_133 N_A_288_21#_M1005_g N_VPWR_c_257_n 0.0127118f $X=1.565 $Y=2.565 $X2=0
+ $Y2=0
cc_134 N_A_288_21#_c_140_n N_VPWR_c_257_n 0.0129681f $X=2.62 $Y=2.145 $X2=0
+ $Y2=0
cc_135 N_A_288_21#_M1005_g N_VPWR_c_258_n 0.0079675f $X=1.565 $Y=2.565 $X2=0
+ $Y2=0
cc_136 N_A_288_21#_c_140_n N_VPWR_c_259_n 0.0173367f $X=2.62 $Y=2.145 $X2=0
+ $Y2=0
cc_137 N_A_288_21#_M1005_g N_VPWR_c_254_n 0.00756802f $X=1.565 $Y=2.565 $X2=0
+ $Y2=0
cc_138 N_A_288_21#_c_140_n N_VPWR_c_254_n 0.0110393f $X=2.62 $Y=2.145 $X2=0
+ $Y2=0
cc_139 N_A_288_21#_M1005_g N_Y_c_303_n 0.0197938f $X=1.565 $Y=2.565 $X2=0 $Y2=0
cc_140 N_A_288_21#_c_140_n N_Y_c_303_n 0.0129587f $X=2.62 $Y=2.145 $X2=0 $Y2=0
cc_141 N_A_288_21#_c_131_n N_Y_c_290_n 0.0105351f $X=1.515 $Y=1.36 $X2=0 $Y2=0
cc_142 N_A_288_21#_M1005_g N_Y_c_290_n 0.00137061f $X=1.565 $Y=2.565 $X2=0 $Y2=0
cc_143 N_A_288_21#_c_133_n N_Y_c_290_n 0.00374726f $X=1.565 $Y=1.435 $X2=0 $Y2=0
cc_144 N_A_288_21#_c_135_n N_Y_c_290_n 3.76673e-19 $X=2.62 $Y=1.495 $X2=0 $Y2=0
cc_145 N_A_288_21#_c_136_n N_Y_c_290_n 0.00666596f $X=3.16 $Y=1.495 $X2=0 $Y2=0
cc_146 N_A_288_21#_c_138_n N_Y_c_290_n 0.016663f $X=2.455 $Y=1.495 $X2=0 $Y2=0
cc_147 N_A_288_21#_M1005_g N_Y_c_292_n 0.0173016f $X=1.565 $Y=2.565 $X2=0 $Y2=0
cc_148 N_A_288_21#_M1005_g Y 0.012844f $X=1.565 $Y=2.565 $X2=0 $Y2=0
cc_149 N_A_288_21#_c_140_n Y 0.0507529f $X=2.62 $Y=2.145 $X2=0 $Y2=0
cc_150 N_A_288_21#_c_135_n Y 8.45163e-19 $X=2.62 $Y=1.495 $X2=0 $Y2=0
cc_151 N_A_288_21#_c_136_n Y 0.00920749f $X=3.16 $Y=1.495 $X2=0 $Y2=0
cc_152 N_A_288_21#_c_138_n Y 0.016883f $X=2.455 $Y=1.495 $X2=0 $Y2=0
cc_153 N_A_288_21#_M1005_g Y 0.0168606f $X=1.565 $Y=2.565 $X2=0 $Y2=0
cc_154 N_A_288_21#_c_131_n N_A_28_110#_c_338_n 0.00868289f $X=1.515 $Y=1.36
+ $X2=0 $Y2=0
cc_155 N_A_288_21#_c_131_n N_VGND_c_360_n 0.0106269f $X=1.515 $Y=1.36 $X2=0
+ $Y2=0
cc_156 N_A_288_21#_c_137_n N_VGND_c_360_n 0.0105391f $X=3.08 $Y=0.41 $X2=0 $Y2=0
cc_157 N_A_288_21#_c_131_n N_VGND_c_362_n 0.00558995f $X=1.515 $Y=1.36 $X2=0
+ $Y2=0
cc_158 N_A_288_21#_c_137_n N_VGND_c_363_n 0.0164408f $X=3.08 $Y=0.41 $X2=0 $Y2=0
cc_159 N_A_288_21#_M1008_d N_VGND_c_364_n 0.00234032f $X=2.94 $Y=0.235 $X2=0
+ $Y2=0
cc_160 N_A_288_21#_c_131_n N_VGND_c_364_n 0.011603f $X=1.515 $Y=1.36 $X2=0 $Y2=0
cc_161 N_A_288_21#_c_137_n N_VGND_c_364_n 0.0121866f $X=3.08 $Y=0.41 $X2=0 $Y2=0
cc_162 N_B1_N_c_207_n N_VPWR_c_257_n 0.00848723f $X=2.355 $Y=3.075 $X2=0 $Y2=0
cc_163 N_B1_N_c_209_n N_VPWR_c_259_n 0.0307431f $X=2.48 $Y=3.15 $X2=0 $Y2=0
cc_164 N_B1_N_c_208_n N_VPWR_c_254_n 0.0317841f $X=3.025 $Y=3.15 $X2=0 $Y2=0
cc_165 N_B1_N_c_209_n N_VPWR_c_254_n 0.0148748f $X=2.48 $Y=3.15 $X2=0 $Y2=0
cc_166 N_B1_N_c_207_n N_Y_c_303_n 0.00765179f $X=2.355 $Y=3.075 $X2=0 $Y2=0
cc_167 N_B1_N_M1007_g N_Y_c_290_n 0.00443037f $X=2.505 $Y=0.445 $X2=0 $Y2=0
cc_168 B1_N N_Y_c_290_n 0.0151748f $X=2.555 $Y=0.84 $X2=0 $Y2=0
cc_169 N_B1_N_c_206_n N_Y_c_290_n 0.00142535f $X=2.415 $Y=0.955 $X2=0 $Y2=0
cc_170 B1_N Y 0.00101005f $X=2.555 $Y=0.84 $X2=0 $Y2=0
cc_171 N_B1_N_c_207_n Y 0.0170298f $X=2.355 $Y=3.075 $X2=0 $Y2=0
cc_172 N_B1_N_M1007_g N_VGND_c_360_n 0.0123954f $X=2.505 $Y=0.445 $X2=0 $Y2=0
cc_173 N_B1_N_M1008_g N_VGND_c_360_n 0.00228984f $X=2.865 $Y=0.445 $X2=0 $Y2=0
cc_174 B1_N N_VGND_c_360_n 0.0131124f $X=2.555 $Y=0.84 $X2=0 $Y2=0
cc_175 N_B1_N_c_206_n N_VGND_c_360_n 0.0039899f $X=2.415 $Y=0.955 $X2=0 $Y2=0
cc_176 N_B1_N_M1007_g N_VGND_c_363_n 0.00486043f $X=2.505 $Y=0.445 $X2=0 $Y2=0
cc_177 N_B1_N_M1008_g N_VGND_c_363_n 0.00550269f $X=2.865 $Y=0.445 $X2=0 $Y2=0
cc_178 N_B1_N_M1007_g N_VGND_c_364_n 0.00430361f $X=2.505 $Y=0.445 $X2=0 $Y2=0
cc_179 N_B1_N_M1008_g N_VGND_c_364_n 0.0107628f $X=2.865 $Y=0.445 $X2=0 $Y2=0
cc_180 B1_N N_VGND_c_364_n 0.0112956f $X=2.555 $Y=0.84 $X2=0 $Y2=0
cc_181 N_VPWR_M1005_d N_Y_c_303_n 0.00874403f $X=1.69 $Y=2.065 $X2=0 $Y2=0
cc_182 N_VPWR_c_257_n N_Y_c_303_n 0.0226318f $X=1.83 $Y=2.87 $X2=0 $Y2=0
cc_183 N_VPWR_c_254_n N_Y_c_303_n 0.0173205f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_184 N_VPWR_c_256_n N_Y_c_292_n 0.0184795f $X=0.31 $Y=2.475 $X2=0 $Y2=0
cc_185 N_VPWR_c_257_n N_Y_c_292_n 0.0266857f $X=1.83 $Y=2.87 $X2=0 $Y2=0
cc_186 N_VPWR_c_258_n N_Y_c_292_n 0.0177952f $X=1.665 $Y=3.33 $X2=0 $Y2=0
cc_187 N_VPWR_c_254_n N_Y_c_292_n 0.0124497f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_188 N_VPWR_M1005_d Y 0.00270082f $X=1.69 $Y=2.065 $X2=0 $Y2=0
cc_189 N_Y_c_290_n N_A_28_110#_c_338_n 0.022684f $X=1.73 $Y=0.76 $X2=0 $Y2=0
cc_190 N_Y_c_290_n N_VGND_c_360_n 9.90462e-19 $X=1.73 $Y=0.76 $X2=0 $Y2=0
cc_191 N_Y_c_290_n N_VGND_c_362_n 0.00523326f $X=1.73 $Y=0.76 $X2=0 $Y2=0
cc_192 N_Y_c_290_n N_VGND_c_364_n 0.00774263f $X=1.73 $Y=0.76 $X2=0 $Y2=0
cc_193 N_A_28_110#_c_336_n N_VGND_M1003_d 0.00353167f $X=1.135 $Y=1.015
+ $X2=-0.19 $Y2=-0.245
cc_194 N_A_28_110#_c_336_n N_VGND_c_359_n 0.0257907f $X=1.135 $Y=1.015 $X2=0
+ $Y2=0
cc_195 N_A_28_110#_c_337_n N_VGND_c_359_n 0.0112721f $X=0.285 $Y=0.77 $X2=0
+ $Y2=0
cc_196 N_A_28_110#_c_337_n N_VGND_c_361_n 0.00604016f $X=0.285 $Y=0.77 $X2=0
+ $Y2=0
cc_197 N_A_28_110#_c_338_n N_VGND_c_362_n 0.00544019f $X=1.3 $Y=0.77 $X2=0 $Y2=0
cc_198 N_A_28_110#_c_337_n N_VGND_c_364_n 0.00989534f $X=0.285 $Y=0.77 $X2=0
+ $Y2=0
cc_199 N_A_28_110#_c_338_n N_VGND_c_364_n 0.00976012f $X=1.3 $Y=0.77 $X2=0 $Y2=0
cc_200 N_VGND_c_364_n A_516_47# 0.00393598f $X=3.12 $Y=0 $X2=-0.19 $Y2=-0.245
