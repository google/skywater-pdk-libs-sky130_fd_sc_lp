* File: sky130_fd_sc_lp__nand2b_4.pex.spice
* Created: Wed Sep  2 10:03:40 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__NAND2B_4%A_N 3 7 9 12 13
r33 12 15 45.3519 $w=3.85e-07 $l=1.65e-07 $layer=POLY_cond $X=0.357 $Y=1.46
+ $X2=0.357 $Y2=1.625
r34 12 14 45.3519 $w=3.85e-07 $l=1.65e-07 $layer=POLY_cond $X=0.357 $Y=1.46
+ $X2=0.357 $Y2=1.295
r35 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.33
+ $Y=1.46 $X2=0.33 $Y2=1.46
r36 9 13 6.94855 $w=3.38e-07 $l=2.05e-07 $layer=LI1_cond $X=0.325 $Y=1.665
+ $X2=0.325 $Y2=1.46
r37 7 15 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=0.475 $Y=2.465
+ $X2=0.475 $Y2=1.625
r38 3 14 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=0.475 $Y=0.675
+ $X2=0.475 $Y2=1.295
.ends

.subckt PM_SKY130_FD_SC_LP__NAND2B_4%A_27_51# 1 2 9 13 17 21 25 29 33 37 41 43
+ 45 47 48 49 52 54 60 65 66 76
c129 33 0 6.6899e-20 $X=2.715 $Y=2.465
r130 75 76 24.4806 $w=3.3e-07 $l=1.4e-07 $layer=POLY_cond $X=2.715 $Y=1.51
+ $X2=2.855 $Y2=1.51
r131 74 75 62.9501 $w=3.3e-07 $l=3.6e-07 $layer=POLY_cond $X=2.355 $Y=1.51
+ $X2=2.715 $Y2=1.51
r132 71 72 13.9889 $w=3.3e-07 $l=8e-08 $layer=POLY_cond $X=1.775 $Y=1.51
+ $X2=1.855 $Y2=1.51
r133 70 71 61.2015 $w=3.3e-07 $l=3.5e-07 $layer=POLY_cond $X=1.425 $Y=1.51
+ $X2=1.775 $Y2=1.51
r134 69 70 13.9889 $w=3.3e-07 $l=8e-08 $layer=POLY_cond $X=1.345 $Y=1.51
+ $X2=1.425 $Y2=1.51
r135 66 69 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=1.27 $Y=1.51
+ $X2=1.345 $Y2=1.51
r136 61 74 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=2.285 $Y=1.51
+ $X2=2.355 $Y2=1.51
r137 61 72 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=2.285 $Y=1.51
+ $X2=1.855 $Y2=1.51
r138 60 61 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=2.285
+ $Y=1.51 $X2=2.285 $Y2=1.51
r139 58 66 60.3271 $w=3.3e-07 $l=3.45e-07 $layer=POLY_cond $X=0.925 $Y=1.51
+ $X2=1.27 $Y2=1.51
r140 57 60 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=0.925 $Y=1.51
+ $X2=2.285 $Y2=1.51
r141 57 58 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=0.925
+ $Y=1.51 $X2=0.925 $Y2=1.51
r142 55 65 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.835 $Y=1.51
+ $X2=0.75 $Y2=1.51
r143 55 57 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=0.835 $Y=1.51
+ $X2=0.925 $Y2=1.51
r144 53 65 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.75 $Y=1.595
+ $X2=0.75 $Y2=1.51
r145 53 54 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=0.75 $Y=1.595
+ $X2=0.75 $Y2=1.93
r146 52 65 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.75 $Y=1.425
+ $X2=0.75 $Y2=1.51
r147 51 52 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=0.75 $Y=1.195
+ $X2=0.75 $Y2=1.425
r148 50 64 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.355 $Y=2.015
+ $X2=0.225 $Y2=2.015
r149 49 54 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.665 $Y=2.015
+ $X2=0.75 $Y2=1.93
r150 49 50 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=0.665 $Y=2.015
+ $X2=0.355 $Y2=2.015
r151 47 51 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.665 $Y=1.11
+ $X2=0.75 $Y2=1.195
r152 47 48 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=0.665 $Y=1.11
+ $X2=0.345 $Y2=1.11
r153 43 64 2.85134 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=0.225 $Y=2.1
+ $X2=0.225 $Y2=2.015
r154 43 45 35.903 $w=2.58e-07 $l=8.1e-07 $layer=LI1_cond $X=0.225 $Y=2.1
+ $X2=0.225 $Y2=2.91
r155 39 48 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.22 $Y=1.025
+ $X2=0.345 $Y2=1.11
r156 39 41 27.8891 $w=2.48e-07 $l=6.05e-07 $layer=LI1_cond $X=0.22 $Y=1.025
+ $X2=0.22 $Y2=0.42
r157 35 76 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.855 $Y=1.345
+ $X2=2.855 $Y2=1.51
r158 35 37 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=2.855 $Y=1.345
+ $X2=2.855 $Y2=0.745
r159 31 75 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.715 $Y=1.675
+ $X2=2.715 $Y2=1.51
r160 31 33 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.715 $Y=1.675
+ $X2=2.715 $Y2=2.465
r161 27 74 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.355 $Y=1.345
+ $X2=2.355 $Y2=1.51
r162 27 29 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=2.355 $Y=1.345
+ $X2=2.355 $Y2=0.745
r163 23 61 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.285 $Y=1.675
+ $X2=2.285 $Y2=1.51
r164 23 25 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.285 $Y=1.675
+ $X2=2.285 $Y2=2.465
r165 19 72 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.855 $Y=1.345
+ $X2=1.855 $Y2=1.51
r166 19 21 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=1.855 $Y=1.345
+ $X2=1.855 $Y2=0.745
r167 15 71 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.775 $Y=1.675
+ $X2=1.775 $Y2=1.51
r168 15 17 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.775 $Y=1.675
+ $X2=1.775 $Y2=2.465
r169 11 70 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.425 $Y=1.345
+ $X2=1.425 $Y2=1.51
r170 11 13 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=1.425 $Y=1.345
+ $X2=1.425 $Y2=0.745
r171 7 69 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.345 $Y=1.675
+ $X2=1.345 $Y2=1.51
r172 7 9 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.345 $Y=1.675
+ $X2=1.345 $Y2=2.465
r173 2 64 400 $w=1.7e-07 $l=3.16386e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.835 $X2=0.26 $Y2=2.095
r174 2 45 400 $w=1.7e-07 $l=1.13578e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.835 $X2=0.26 $Y2=2.91
r175 1 41 91 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.255 $X2=0.26 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__NAND2B_4%B 3 7 11 15 19 23 27 31 33 34 35 57
c74 35 0 6.6899e-20 $X=5.04 $Y=1.665
c75 3 0 8.67364e-20 $X=3.285 $Y=0.745
r76 57 58 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.775
+ $Y=1.51 $X2=4.775 $Y2=1.51
r77 55 57 24.4806 $w=3.3e-07 $l=1.4e-07 $layer=POLY_cond $X=4.635 $Y=1.51
+ $X2=4.775 $Y2=1.51
r78 54 55 10.4917 $w=3.3e-07 $l=6e-08 $layer=POLY_cond $X=4.575 $Y=1.51
+ $X2=4.635 $Y2=1.51
r79 52 54 24.4806 $w=3.3e-07 $l=1.4e-07 $layer=POLY_cond $X=4.435 $Y=1.51
+ $X2=4.575 $Y2=1.51
r80 52 53 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.435
+ $Y=1.51 $X2=4.435 $Y2=1.51
r81 50 52 40.2181 $w=3.3e-07 $l=2.3e-07 $layer=POLY_cond $X=4.205 $Y=1.51
+ $X2=4.435 $Y2=1.51
r82 49 50 10.4917 $w=3.3e-07 $l=6e-08 $layer=POLY_cond $X=4.145 $Y=1.51
+ $X2=4.205 $Y2=1.51
r83 48 53 11.6964 $w=3.33e-07 $l=3.4e-07 $layer=LI1_cond $X=4.095 $Y=1.592
+ $X2=4.435 $Y2=1.592
r84 47 49 8.74306 $w=3.3e-07 $l=5e-08 $layer=POLY_cond $X=4.095 $Y=1.51
+ $X2=4.145 $Y2=1.51
r85 47 48 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.095
+ $Y=1.51 $X2=4.095 $Y2=1.51
r86 45 47 55.9556 $w=3.3e-07 $l=3.2e-07 $layer=POLY_cond $X=3.775 $Y=1.51
+ $X2=4.095 $Y2=1.51
r87 43 45 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=3.755 $Y=1.51
+ $X2=3.775 $Y2=1.51
r88 43 44 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.755
+ $Y=1.51 $X2=3.755 $Y2=1.51
r89 41 43 6.99445 $w=3.3e-07 $l=4e-08 $layer=POLY_cond $X=3.715 $Y=1.51
+ $X2=3.755 $Y2=1.51
r90 39 41 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=3.285 $Y=1.51
+ $X2=3.715 $Y2=1.51
r91 35 58 9.11634 $w=3.33e-07 $l=2.65e-07 $layer=LI1_cond $X=5.04 $Y=1.592
+ $X2=4.775 $Y2=1.592
r92 34 58 7.39628 $w=3.33e-07 $l=2.15e-07 $layer=LI1_cond $X=4.56 $Y=1.592
+ $X2=4.775 $Y2=1.592
r93 34 53 4.30016 $w=3.33e-07 $l=1.25e-07 $layer=LI1_cond $X=4.56 $Y=1.592
+ $X2=4.435 $Y2=1.592
r94 33 48 0.516019 $w=3.33e-07 $l=1.5e-08 $layer=LI1_cond $X=4.08 $Y=1.592
+ $X2=4.095 $Y2=1.592
r95 33 44 11.1804 $w=3.33e-07 $l=3.25e-07 $layer=LI1_cond $X=4.08 $Y=1.592
+ $X2=3.755 $Y2=1.592
r96 29 55 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.635 $Y=1.675
+ $X2=4.635 $Y2=1.51
r97 29 31 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=4.635 $Y=1.675
+ $X2=4.635 $Y2=2.465
r98 25 54 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.575 $Y=1.345
+ $X2=4.575 $Y2=1.51
r99 25 27 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=4.575 $Y=1.345
+ $X2=4.575 $Y2=0.745
r100 21 50 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.205 $Y=1.675
+ $X2=4.205 $Y2=1.51
r101 21 23 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=4.205 $Y=1.675
+ $X2=4.205 $Y2=2.465
r102 17 49 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.145 $Y=1.345
+ $X2=4.145 $Y2=1.51
r103 17 19 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=4.145 $Y=1.345
+ $X2=4.145 $Y2=0.745
r104 13 45 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.775 $Y=1.675
+ $X2=3.775 $Y2=1.51
r105 13 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.775 $Y=1.675
+ $X2=3.775 $Y2=2.465
r106 9 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.715 $Y=1.345
+ $X2=3.715 $Y2=1.51
r107 9 11 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=3.715 $Y=1.345
+ $X2=3.715 $Y2=0.745
r108 5 39 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.285 $Y=1.675
+ $X2=3.285 $Y2=1.51
r109 5 7 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.285 $Y=1.675
+ $X2=3.285 $Y2=2.465
r110 1 39 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.285 $Y=1.345
+ $X2=3.285 $Y2=1.51
r111 1 3 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=3.285 $Y=1.345 $X2=3.285
+ $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_LP__NAND2B_4%VPWR 1 2 3 4 5 19 22 26 32 36 38 40 45 48
+ 49 51 52 54 55 56 58 73 78 82
r84 81 82 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r85 78 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r86 76 82 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.04 $Y2=3.33
r87 75 76 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r88 73 81 4.48746 $w=1.7e-07 $l=2.97e-07 $layer=LI1_cond $X=4.685 $Y=3.33
+ $X2=4.982 $Y2=3.33
r89 73 75 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=4.685 $Y=3.33
+ $X2=4.56 $Y2=3.33
r90 72 76 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.56 $Y2=3.33
r91 71 72 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r92 66 79 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.72 $Y2=3.33
r93 65 66 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r94 63 78 14.0645 $w=1.7e-07 $l=3.7e-07 $layer=LI1_cond $X=1.265 $Y=3.33
+ $X2=0.895 $Y2=3.33
r95 63 65 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=1.265 $Y=3.33
+ $X2=1.68 $Y2=3.33
r96 61 79 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r97 60 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r98 58 78 14.0645 $w=1.7e-07 $l=3.7e-07 $layer=LI1_cond $X=0.525 $Y=3.33
+ $X2=0.895 $Y2=3.33
r99 58 60 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.525 $Y=3.33
+ $X2=0.24 $Y2=3.33
r100 56 72 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r101 56 66 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=1.68 $Y2=3.33
r102 56 68 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r103 54 71 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=3.86 $Y=3.33
+ $X2=3.6 $Y2=3.33
r104 54 55 7.34436 $w=1.7e-07 $l=1.32e-07 $layer=LI1_cond $X=3.86 $Y=3.33
+ $X2=3.992 $Y2=3.33
r105 53 75 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=4.125 $Y=3.33
+ $X2=4.56 $Y2=3.33
r106 53 55 7.34436 $w=1.7e-07 $l=1.33e-07 $layer=LI1_cond $X=4.125 $Y=3.33
+ $X2=3.992 $Y2=3.33
r107 51 68 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=2.835 $Y=3.33
+ $X2=2.64 $Y2=3.33
r108 51 52 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.835 $Y=3.33 $X2=3
+ $Y2=3.33
r109 50 71 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=3.165 $Y=3.33
+ $X2=3.6 $Y2=3.33
r110 50 52 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.165 $Y=3.33 $X2=3
+ $Y2=3.33
r111 48 65 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=1.865 $Y=3.33
+ $X2=1.68 $Y2=3.33
r112 48 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.865 $Y=3.33
+ $X2=2.03 $Y2=3.33
r113 47 68 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=2.195 $Y=3.33
+ $X2=2.64 $Y2=3.33
r114 47 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.195 $Y=3.33
+ $X2=2.03 $Y2=3.33
r115 45 46 6.71429 $w=7.38e-07 $l=8.5e-08 $layer=LI1_cond $X=0.895 $Y=2.355
+ $X2=0.895 $Y2=2.27
r116 40 43 32.6526 $w=3.28e-07 $l=9.35e-07 $layer=LI1_cond $X=4.85 $Y=2.015
+ $X2=4.85 $Y2=2.95
r117 38 81 3.27872 $w=3.3e-07 $l=1.69245e-07 $layer=LI1_cond $X=4.85 $Y=3.245
+ $X2=4.982 $Y2=3.33
r118 38 43 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=4.85 $Y=3.245
+ $X2=4.85 $Y2=2.95
r119 34 55 0.195364 $w=2.65e-07 $l=8.5e-08 $layer=LI1_cond $X=3.992 $Y=3.245
+ $X2=3.992 $Y2=3.33
r120 34 36 35.2256 $w=2.63e-07 $l=8.1e-07 $layer=LI1_cond $X=3.992 $Y=3.245
+ $X2=3.992 $Y2=2.435
r121 30 52 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3 $Y=3.245 $X2=3
+ $Y2=3.33
r122 30 32 30.3826 $w=3.28e-07 $l=8.7e-07 $layer=LI1_cond $X=3 $Y=3.245 $X2=3
+ $Y2=2.375
r123 26 29 27.2396 $w=3.28e-07 $l=7.8e-07 $layer=LI1_cond $X=2.03 $Y=2.19
+ $X2=2.03 $Y2=2.97
r124 24 49 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.03 $Y=3.245
+ $X2=2.03 $Y2=3.33
r125 24 29 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.03 $Y=3.245
+ $X2=2.03 $Y2=2.97
r126 22 46 13.519 $w=2.58e-07 $l=3.05e-07 $layer=LI1_cond $X=1.135 $Y=1.965
+ $X2=1.135 $Y2=2.27
r127 17 78 2.97738 $w=7.4e-07 $l=8.5e-08 $layer=LI1_cond $X=0.895 $Y=3.245
+ $X2=0.895 $Y2=3.33
r128 17 19 4.76815 $w=7.38e-07 $l=2.95e-07 $layer=LI1_cond $X=0.895 $Y=3.245
+ $X2=0.895 $Y2=2.95
r129 16 45 4.60652 $w=7.38e-07 $l=2.85e-07 $layer=LI1_cond $X=0.895 $Y=2.64
+ $X2=0.895 $Y2=2.355
r130 16 19 5.0106 $w=7.38e-07 $l=3.1e-07 $layer=LI1_cond $X=0.895 $Y=2.64
+ $X2=0.895 $Y2=2.95
r131 5 43 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=4.71
+ $Y=1.835 $X2=4.85 $Y2=2.95
r132 5 40 400 $w=1.7e-07 $l=2.4e-07 $layer=licon1_PDIFF $count=1 $X=4.71
+ $Y=1.835 $X2=4.85 $Y2=2.015
r133 4 36 300 $w=1.7e-07 $l=6.66333e-07 $layer=licon1_PDIFF $count=2 $X=3.85
+ $Y=1.835 $X2=3.99 $Y2=2.435
r134 3 32 300 $w=1.7e-07 $l=6.36396e-07 $layer=licon1_PDIFF $count=2 $X=2.79
+ $Y=1.835 $X2=3 $Y2=2.375
r135 2 29 400 $w=1.7e-07 $l=1.22169e-06 $layer=licon1_PDIFF $count=1 $X=1.85
+ $Y=1.835 $X2=2.03 $Y2=2.97
r136 2 26 400 $w=1.7e-07 $l=4.35804e-07 $layer=licon1_PDIFF $count=1 $X=1.85
+ $Y=1.835 $X2=2.03 $Y2=2.19
r137 1 45 300 $w=1.7e-07 $l=5.85833e-07 $layer=licon1_PDIFF $count=2 $X=0.55
+ $Y=1.835 $X2=0.69 $Y2=2.355
r138 1 22 600 $w=1.7e-07 $l=6.41716e-07 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=1.835 $X2=1.13 $Y2=1.965
r139 1 19 300 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=2 $X=0.55
+ $Y=1.835 $X2=0.69 $Y2=2.95
.ends

.subckt PM_SKY130_FD_SC_LP__NAND2B_4%Y 1 2 3 4 5 6 21 27 29 30 31 32 35 38 39 41
+ 43 45 48 49 50 57 58 60 64 69
c90 45 0 8.67364e-20 $X=2.64 $Y=1.17
r91 73 74 0.324468 $w=5.64e-07 $l=1.5e-08 $layer=LI1_cond $X=2.5 $Y=1.78
+ $X2=2.515 $Y2=1.78
r92 58 60 2.33493 $w=1.88e-07 $l=4e-08 $layer=LI1_cond $X=3.08 $Y=2.025 $X2=3.12
+ $Y2=2.025
r93 50 57 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=3.525 $Y=2.025
+ $X2=3.36 $Y2=2.025
r94 50 69 20.2817 $w=4.98e-07 $l=7.9e-07 $layer=LI1_cond $X=3.525 $Y=2.12
+ $X2=3.525 $Y2=2.91
r95 49 58 6.24499 $w=5.64e-07 $l=2.56242e-07 $layer=LI1_cond $X=3.057 $Y=1.78
+ $X2=3.08 $Y2=2.025
r96 49 77 7.46277 $w=5.64e-07 $l=3.45e-07 $layer=LI1_cond $X=3.057 $Y=1.78
+ $X2=2.712 $Y2=1.78
r97 49 57 12.7254 $w=1.88e-07 $l=2.18e-07 $layer=LI1_cond $X=3.142 $Y=2.025
+ $X2=3.36 $Y2=2.025
r98 49 60 1.28421 $w=1.88e-07 $l=2.2e-08 $layer=LI1_cond $X=3.142 $Y=2.025
+ $X2=3.12 $Y2=2.025
r99 48 77 1.55745 $w=5.64e-07 $l=7.2e-08 $layer=LI1_cond $X=2.64 $Y=1.78
+ $X2=2.712 $Y2=1.78
r100 48 74 2.7039 $w=5.64e-07 $l=1.25e-07 $layer=LI1_cond $X=2.64 $Y=1.78
+ $X2=2.515 $Y2=1.78
r101 48 74 4.43409 $w=3e-07 $l=3.4e-07 $layer=LI1_cond $X=2.515 $Y=2.12
+ $X2=2.515 $Y2=1.78
r102 48 64 23.0568 $w=4.08e-07 $l=7.9e-07 $layer=LI1_cond $X=2.515 $Y=2.12
+ $X2=2.515 $Y2=2.91
r103 41 47 3.03526 $w=2.2e-07 $l=8.5e-08 $layer=LI1_cond $X=4.405 $Y=2.1
+ $X2=4.405 $Y2=2.015
r104 41 43 42.4309 $w=2.18e-07 $l=8.1e-07 $layer=LI1_cond $X=4.405 $Y=2.1
+ $X2=4.405 $Y2=2.91
r105 40 50 8.26956 $w=1.8e-07 $l=1.69926e-07 $layer=LI1_cond $X=3.69 $Y=2.015
+ $X2=3.525 $Y2=2.025
r106 39 47 3.92798 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=4.295 $Y=2.015
+ $X2=4.405 $Y2=2.015
r107 39 40 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=4.295 $Y=2.015
+ $X2=3.69 $Y2=2.015
r108 38 77 7.3934 $w=1.85e-07 $l=3.4e-07 $layer=LI1_cond $X=2.712 $Y=1.44
+ $X2=2.712 $Y2=1.78
r109 37 45 3.6114 $w=2.57e-07 $l=1.15521e-07 $layer=LI1_cond $X=2.712 $Y=1.255
+ $X2=2.64 $Y2=1.17
r110 37 38 11.0909 $w=1.83e-07 $l=1.85e-07 $layer=LI1_cond $X=2.712 $Y=1.255
+ $X2=2.712 $Y2=1.44
r111 33 45 3.6114 $w=2.57e-07 $l=8.5e-08 $layer=LI1_cond $X=2.64 $Y=1.085
+ $X2=2.64 $Y2=1.17
r112 33 35 13.7944 $w=3.28e-07 $l=3.95e-07 $layer=LI1_cond $X=2.64 $Y=1.085
+ $X2=2.64 $Y2=0.69
r113 31 45 2.87242 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.475 $Y=1.17
+ $X2=2.64 $Y2=1.17
r114 31 32 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.475 $Y=1.17
+ $X2=1.805 $Y2=1.17
r115 29 73 9.4717 $w=5.64e-07 $l=1.66358e-07 $layer=LI1_cond $X=2.365 $Y=1.85
+ $X2=2.5 $Y2=1.78
r116 29 30 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.365 $Y=1.85
+ $X2=1.695 $Y2=1.85
r117 25 32 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.64 $Y=1.085
+ $X2=1.805 $Y2=1.17
r118 25 27 13.7944 $w=3.28e-07 $l=3.95e-07 $layer=LI1_cond $X=1.64 $Y=1.085
+ $X2=1.64 $Y2=0.69
r119 21 23 41.8869 $w=2.58e-07 $l=9.45e-07 $layer=LI1_cond $X=1.565 $Y=1.965
+ $X2=1.565 $Y2=2.91
r120 19 30 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=1.565 $Y=1.935
+ $X2=1.695 $Y2=1.85
r121 19 21 1.32974 $w=2.58e-07 $l=3e-08 $layer=LI1_cond $X=1.565 $Y=1.935
+ $X2=1.565 $Y2=1.965
r122 6 47 400 $w=1.7e-07 $l=3.2249e-07 $layer=licon1_PDIFF $count=1 $X=4.28
+ $Y=1.835 $X2=4.42 $Y2=2.095
r123 6 43 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=4.28
+ $Y=1.835 $X2=4.42 $Y2=2.91
r124 5 50 400 $w=1.7e-07 $l=3.32415e-07 $layer=licon1_PDIFF $count=1 $X=3.36
+ $Y=1.835 $X2=3.525 $Y2=2.095
r125 5 69 400 $w=1.7e-07 $l=1.15456e-06 $layer=licon1_PDIFF $count=1 $X=3.36
+ $Y=1.835 $X2=3.525 $Y2=2.91
r126 4 73 400 $w=1.7e-07 $l=1.94422e-07 $layer=licon1_PDIFF $count=1 $X=2.36
+ $Y=1.835 $X2=2.5 $Y2=1.965
r127 4 64 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=2.36
+ $Y=1.835 $X2=2.5 $Y2=2.91
r128 3 23 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=1.42
+ $Y=1.835 $X2=1.56 $Y2=2.91
r129 3 21 400 $w=1.7e-07 $l=1.94422e-07 $layer=licon1_PDIFF $count=1 $X=1.42
+ $Y=1.835 $X2=1.56 $Y2=1.965
r130 2 35 91 $w=1.7e-07 $l=4.58121e-07 $layer=licon1_NDIFF $count=2 $X=2.43
+ $Y=0.325 $X2=2.64 $Y2=0.69
r131 1 27 91 $w=1.7e-07 $l=4.29331e-07 $layer=licon1_NDIFF $count=2 $X=1.5
+ $Y=0.325 $X2=1.64 $Y2=0.69
.ends

.subckt PM_SKY130_FD_SC_LP__NAND2B_4%VGND 1 2 3 12 16 20 23 24 26 27 28 30 46 47
+ 50
r66 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r67 46 47 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r68 44 47 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=5.04
+ $Y2=0
r69 43 44 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r70 41 44 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=4.08
+ $Y2=0
r71 40 41 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r72 38 51 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r73 37 40 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=3.12
+ $Y2=0
r74 37 38 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r75 35 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.855 $Y=0 $X2=0.69
+ $Y2=0
r76 35 37 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.855 $Y=0 $X2=1.2
+ $Y2=0
r77 33 51 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r78 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r79 30 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.525 $Y=0 $X2=0.69
+ $Y2=0
r80 30 32 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.525 $Y=0 $X2=0.24
+ $Y2=0
r81 28 41 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r82 28 38 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=2.64 $Y=0 $X2=1.2
+ $Y2=0
r83 26 43 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=4.195 $Y=0 $X2=4.08
+ $Y2=0
r84 26 27 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.195 $Y=0 $X2=4.36
+ $Y2=0
r85 25 46 33.5989 $w=1.68e-07 $l=5.15e-07 $layer=LI1_cond $X=4.525 $Y=0 $X2=5.04
+ $Y2=0
r86 25 27 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.525 $Y=0 $X2=4.36
+ $Y2=0
r87 23 40 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=3.335 $Y=0 $X2=3.12
+ $Y2=0
r88 23 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.335 $Y=0 $X2=3.5
+ $Y2=0
r89 22 43 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=3.665 $Y=0 $X2=4.08
+ $Y2=0
r90 22 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.665 $Y=0 $X2=3.5
+ $Y2=0
r91 18 27 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.36 $Y=0.085
+ $X2=4.36 $Y2=0
r92 18 20 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=4.36 $Y=0.085
+ $X2=4.36 $Y2=0.45
r93 14 24 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.5 $Y=0.085 $X2=3.5
+ $Y2=0
r94 14 16 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=3.5 $Y=0.085
+ $X2=3.5 $Y2=0.45
r95 10 50 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=0.085
+ $X2=0.69 $Y2=0
r96 10 12 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=0.69 $Y=0.085
+ $X2=0.69 $Y2=0.4
r97 3 20 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=4.22
+ $Y=0.325 $X2=4.36 $Y2=0.45
r98 2 16 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=3.36
+ $Y=0.325 $X2=3.5 $Y2=0.45
r99 1 12 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=0.55
+ $Y=0.255 $X2=0.69 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_LP__NAND2B_4%A_217_65# 1 2 3 4 5 18 20 21 24 26 32 33 36
+ 38 42 44 45
r73 40 42 26.8165 $w=2.58e-07 $l=6.05e-07 $layer=LI1_cond $X=4.825 $Y=1.075
+ $X2=4.825 $Y2=0.47
r74 39 45 5.52892 $w=1.75e-07 $l=9.5e-08 $layer=LI1_cond $X=4.025 $Y=1.165
+ $X2=3.93 $Y2=1.165
r75 38 40 7.11373 $w=1.8e-07 $l=1.69115e-07 $layer=LI1_cond $X=4.695 $Y=1.165
+ $X2=4.825 $Y2=1.075
r76 38 39 41.2828 $w=1.78e-07 $l=6.7e-07 $layer=LI1_cond $X=4.695 $Y=1.165
+ $X2=4.025 $Y2=1.165
r77 34 45 1.04816 $w=1.9e-07 $l=9e-08 $layer=LI1_cond $X=3.93 $Y=1.075 $X2=3.93
+ $Y2=1.165
r78 34 36 36.4833 $w=1.88e-07 $l=6.25e-07 $layer=LI1_cond $X=3.93 $Y=1.075
+ $X2=3.93 $Y2=0.45
r79 32 45 5.52892 $w=1.75e-07 $l=9.74679e-08 $layer=LI1_cond $X=3.835 $Y=1.17
+ $X2=3.93 $Y2=1.165
r80 32 33 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.835 $Y=1.17
+ $X2=3.165 $Y2=1.17
r81 29 33 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=3.07 $Y=1.085
+ $X2=3.165 $Y2=1.17
r82 29 31 37.067 $w=1.88e-07 $l=6.35e-07 $layer=LI1_cond $X=3.07 $Y=1.085
+ $X2=3.07 $Y2=0.45
r83 28 31 1.45933 $w=1.88e-07 $l=2.5e-08 $layer=LI1_cond $X=3.07 $Y=0.425
+ $X2=3.07 $Y2=0.45
r84 27 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.305 $Y=0.34
+ $X2=2.14 $Y2=0.34
r85 26 28 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=2.975 $Y=0.34
+ $X2=3.07 $Y2=0.425
r86 26 27 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.975 $Y=0.34
+ $X2=2.305 $Y2=0.34
r87 22 44 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.14 $Y=0.425
+ $X2=2.14 $Y2=0.34
r88 22 24 0.873063 $w=3.28e-07 $l=2.5e-08 $layer=LI1_cond $X=2.14 $Y=0.425
+ $X2=2.14 $Y2=0.45
r89 20 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.975 $Y=0.34
+ $X2=2.14 $Y2=0.34
r90 20 21 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.975 $Y=0.34
+ $X2=1.305 $Y2=0.34
r91 16 21 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=1.175 $Y=0.425
+ $X2=1.305 $Y2=0.34
r92 16 18 1.99461 $w=2.58e-07 $l=4.5e-08 $layer=LI1_cond $X=1.175 $Y=0.425
+ $X2=1.175 $Y2=0.47
r93 5 42 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.65
+ $Y=0.325 $X2=4.79 $Y2=0.47
r94 4 36 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=3.79
+ $Y=0.325 $X2=3.93 $Y2=0.45
r95 3 31 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=2.93
+ $Y=0.325 $X2=3.07 $Y2=0.45
r96 2 24 91 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=2 $X=1.93
+ $Y=0.325 $X2=2.14 $Y2=0.45
r97 1 18 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=1.085
+ $Y=0.325 $X2=1.21 $Y2=0.47
.ends

