* File: sky130_fd_sc_lp__srsdfxtp_1.spice
* Created: Wed Sep  2 10:39:30 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__srsdfxtp_1.pex.spice"
.subckt sky130_fd_sc_lp__srsdfxtp_1  VNB VPB SCE D SCD SLEEP_B CLK VPWR KAPWR Q
+ VGND
* 
* VGND	VGND
* Q	Q
* KAPWR	KAPWR
* VPWR	VPWR
* CLK	CLK
* SLEEP_B	SLEEP_B
* SCD	SCD
* D	D
* SCE	SCE
* VPB	VPB
* VNB	VNB
MM1040 N_VGND_M1040_d N_SCE_M1040_g N_A_31_477#_M1040_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.1197 PD=0.7 PS=1.41 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75002.4
+ A=0.063 P=1.14 MULT=1
MM1037 A_210_47# N_A_31_477#_M1037_g N_VGND_M1040_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.0588 PD=0.66 PS=0.7 NRD=18.564 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75002 A=0.063 P=1.14 MULT=1
MM1003 N_A_282_477#_M1003_d N_D_M1003_g A_210_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.0819 AS=0.0504 PD=0.81 PS=0.66 NRD=31.428 NRS=18.564 M=1 R=2.8 SA=75001
+ SB=75001.6 A=0.063 P=1.14 MULT=1
MM1018 A_396_47# N_SCE_M1018_g N_A_282_477#_M1003_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.0819 PD=0.66 PS=0.81 NRD=18.564 NRS=0 M=1 R=2.8 SA=75001.6
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1016 N_VGND_M1016_d N_SCD_M1016_g A_396_47# VNB NSHORT L=0.15 W=0.42 AD=0.0693
+ AS=0.0504 PD=0.75 PS=0.66 NRD=14.28 NRS=18.564 M=1 R=2.8 SA=75002 SB=75000.7
+ A=0.063 P=1.14 MULT=1
MM1025 N_A_570_47#_M1025_d N_A_540_21#_M1025_g N_VGND_M1016_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1176 AS=0.0693 PD=1.4 PS=0.75 NRD=0 NRS=0 M=1 R=2.8 SA=75002.4
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1005 N_A_786_139#_M1005_d N_A_540_21#_M1005_g N_A_282_477#_M1005_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.0588 AS=0.1197 PD=0.7 PS=1.41 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75004 A=0.063 P=1.14 MULT=1
MM1008 A_872_139# N_A_570_47#_M1008_g N_A_786_139#_M1005_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0504 AS=0.0588 PD=0.66 PS=0.7 NRD=18.564 NRS=0 M=1 R=2.8
+ SA=75000.6 SB=75003.6 A=0.063 P=1.14 MULT=1
MM1034 N_VGND_M1034_d N_A_914_245#_M1034_g A_872_139# VNB NSHORT L=0.15 W=0.42
+ AD=0.198628 AS=0.0504 PD=1.29566 PS=0.66 NRD=119.4 NRS=18.564 M=1 R=2.8
+ SA=75001 SB=75003.2 A=0.063 P=1.14 MULT=1
MM1038 N_A_914_245#_M1038_d N_A_786_139#_M1038_g N_VGND_M1034_d VNB NSHORT
+ L=0.15 W=0.64 AD=0.1696 AS=0.302672 PD=1.17 PS=1.97434 NRD=0 NRS=78.36 M=1
+ R=4.26667 SA=75001.1 SB=75002.8 A=0.096 P=1.58 MULT=1
MM1028 A_1247_69# N_A_570_47#_M1028_g N_A_914_245#_M1038_d VNB NSHORT L=0.15
+ W=0.64 AD=0.0672 AS=0.1696 PD=0.85 PS=1.17 NRD=9.372 NRS=46.872 M=1 R=4.26667
+ SA=75001.8 SB=75002.1 A=0.096 P=1.58 MULT=1
MM1012 N_A_1319_69#_M1012_d N_A_570_47#_M1012_g A_1247_69# VNB NSHORT L=0.15
+ W=0.64 AD=0.187109 AS=0.0672 PD=1.38868 PS=0.85 NRD=43.116 NRS=9.372 M=1
+ R=4.26667 SA=75002.1 SB=75001.7 A=0.096 P=1.58 MULT=1
MM1026 A_1451_113# N_A_540_21#_M1026_g N_A_1319_69#_M1012_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.122791 PD=0.63 PS=0.911321 NRD=14.28 NRS=0 M=1 R=2.8
+ SA=75003.1 SB=75001.8 A=0.063 P=1.14 MULT=1
MM1019 A_1523_113# N_A_1493_21#_M1019_g A_1451_113# VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0441 PD=0.63 PS=0.63 NRD=14.28 NRS=14.28 M=1 R=2.8 SA=75003.5
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1006 N_VGND_M1006_d N_A_1493_21#_M1006_g A_1523_113# VNB NSHORT L=0.15 W=0.42
+ AD=0.08715 AS=0.0441 PD=0.875 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75003.8
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1020 A_1704_125# N_A_1319_69#_M1020_g N_VGND_M1006_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.08715 PD=0.63 PS=0.875 NRD=14.28 NRS=32.856 M=1 R=2.8
+ SA=75003.9 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1007 N_A_1493_21#_M1007_d N_A_1319_69#_M1007_g A_1704_125# VNB NSHORT L=0.15
+ W=0.42 AD=0.1738 AS=0.0441 PD=1.68 PS=0.63 NRD=32.856 NRS=14.28 M=1 R=2.8
+ SA=75004.3 SB=75000.3 A=0.063 P=1.14 MULT=1
MM1013 A_2243_178# N_CLK_M1013_g N_A_540_21#_M1013_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.168 PD=0.66 PS=1.64 NRD=18.564 NRS=32.856 M=1 R=2.8 SA=75000.3
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1002 A_2321_178# N_SLEEP_B_M1002_g A_2243_178# VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0504 PD=0.63 PS=0.66 NRD=14.28 NRS=18.564 M=1 R=2.8 SA=75000.7
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1033 N_VGND_M1033_d N_SLEEP_B_M1033_g A_2321_178# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.1
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1032 N_VGND_M1032_d N_A_1319_69#_M1032_g N_A_2504_57#_M1032_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.0952 AS=0.1197 PD=0.823333 PS=1.41 NRD=32.856 NRS=0 M=1
+ R=2.8 SA=75000.2 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1031 N_Q_M1031_d N_A_2504_57#_M1031_g N_VGND_M1032_d VNB NSHORT L=0.15 W=0.84
+ AD=0.2394 AS=0.1904 PD=2.25 PS=1.64667 NRD=0 NRS=0 M=1 R=5.6 SA=75000.5
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1030 N_VPWR_M1030_d N_SCE_M1030_g N_A_31_477#_M1030_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.0896 AS=0.1824 PD=0.92 PS=1.85 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75002.8 A=0.096 P=1.58 MULT=1
MM1000 A_204_477# N_SCE_M1000_g N_VPWR_M1030_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0768 AS=0.0896 PD=0.88 PS=0.92 NRD=19.9955 NRS=0 M=1 R=4.26667 SA=75000.6
+ SB=75002.3 A=0.096 P=1.58 MULT=1
MM1021 N_A_282_477#_M1021_d N_D_M1021_g A_204_477# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0896 AS=0.0768 PD=0.92 PS=0.88 NRD=0 NRS=19.9955 M=1 R=4.26667 SA=75001
+ SB=75001.9 A=0.096 P=1.58 MULT=1
MM1004 A_368_477# N_A_31_477#_M1004_g N_A_282_477#_M1021_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1024 AS=0.0896 PD=0.96 PS=0.92 NRD=32.308 NRS=0 M=1 R=4.26667
+ SA=75001.5 SB=75001.5 A=0.096 P=1.58 MULT=1
MM1039 N_VPWR_M1039_d N_SCD_M1039_g A_368_477# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.2208 AS=0.1024 PD=1.33 PS=0.96 NRD=35.3812 NRS=32.308 M=1 R=4.26667
+ SA=75001.9 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1027 N_A_570_47#_M1027_d N_A_540_21#_M1027_g N_VPWR_M1039_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1824 AS=0.2208 PD=1.85 PS=1.33 NRD=0 NRS=90.7973 M=1 R=4.26667
+ SA=75002.8 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1035 N_A_786_139#_M1035_d N_A_570_47#_M1035_g N_A_282_477#_M1035_s VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.0588 AS=0.1491 PD=0.7 PS=1.55 NRD=0 NRS=32.8202 M=1 R=2.8
+ SA=75000.3 SB=75001.9 A=0.063 P=1.14 MULT=1
MM1022 A_1010_530# N_A_540_21#_M1022_g N_A_786_139#_M1035_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0504 AS=0.0588 PD=0.66 PS=0.7 NRD=30.4759 NRS=0 M=1 R=2.8
+ SA=75000.7 SB=75001.5 A=0.063 P=1.14 MULT=1
MM1036 N_VPWR_M1036_d N_A_914_245#_M1036_g A_1010_530# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.159525 AS=0.0504 PD=1.22 PS=0.66 NRD=39.8531 NRS=30.4759 M=1 R=2.8
+ SA=75001.1 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1023 N_A_914_245#_M1023_d N_A_786_139#_M1023_g N_VPWR_M1036_d VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.1673 AS=0.31905 PD=1.43 PS=2.44 NRD=2.3443 NRS=76.1602 M=1
+ R=5.6 SA=75000.9 SB=75000.8 A=0.126 P=1.98 MULT=1
MM1009 A_1372_379# N_A_540_21#_M1009_g N_A_914_245#_M1023_d VPB PHIGHVT L=0.15
+ W=0.84 AD=0.0882 AS=0.1673 PD=1.05 PS=1.43 NRD=11.7215 NRS=16.4101 M=1 R=5.6
+ SA=75000.7 SB=75000.6 A=0.126 P=1.98 MULT=1
MM1014 N_A_1319_69#_M1014_d N_A_540_21#_M1014_g A_1372_379# VPB PHIGHVT L=0.15
+ W=0.84 AD=0.2394 AS=0.0882 PD=2.25 PS=1.05 NRD=0 NRS=11.7215 M=1 R=5.6
+ SA=75001.1 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1001 A_1858_419# N_A_570_47#_M1001_g N_A_1319_69#_M1001_s VPB PHIGHVT L=0.25
+ W=1 AD=0.12 AS=0.285 PD=1.24 PS=2.57 NRD=12.7853 NRS=0 M=1 R=4 SA=125000
+ SB=125002 A=0.25 P=2.5 MULT=1
MM1017 N_KAPWR_M1017_d N_A_1493_21#_M1017_g A_1858_419# VPB PHIGHVT L=0.25 W=1
+ AD=0.216707 AS=0.12 PD=1.70122 PS=1.24 NRD=0 NRS=12.7853 M=1 R=4 SA=125001
+ SB=125001 A=0.25 P=2.5 MULT=1
MM1010 N_A_540_21#_M1010_d N_SLEEP_B_M1010_g N_KAPWR_M1017_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.176 AS=0.138693 PD=1.19 PS=1.08878 NRD=41.5473 NRS=49.7622 M=1
+ R=4.26667 SA=75001.3 SB=75001.7 A=0.096 P=1.58 MULT=1
MM1015 N_KAPWR_M1015_d N_CLK_M1015_g N_A_540_21#_M1010_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.138693 AS=0.176 PD=1.08878 PS=1.19 NRD=49.7622 NRS=41.5473 M=1
+ R=4.26667 SA=75002 SB=75001 A=0.096 P=1.58 MULT=1
MM1029 N_A_1493_21#_M1029_d N_A_1319_69#_M1029_g N_KAPWR_M1015_d VPB PHIGHVT
+ L=0.25 W=1 AD=0.435 AS=0.216707 PD=2.87 PS=1.70122 NRD=29.55 NRS=0 M=1 R=4
+ SA=125002 SB=125000 A=0.25 P=2.5 MULT=1
MM1011 N_VPWR_M1011_d N_A_1319_69#_M1011_g N_A_2504_57#_M1011_s VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.144674 AS=0.1824 PD=1.11495 PS=1.85 NRD=36.1495 NRS=0 M=1
+ R=4.26667 SA=75000.2 SB=75000.8 A=0.096 P=1.58 MULT=1
MM1024 N_Q_M1024_d N_A_2504_57#_M1024_g N_VPWR_M1011_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3591 AS=0.284826 PD=3.09 PS=2.19505 NRD=0 NRS=0 M=1 R=8.4 SA=75000.5
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX41_noxref VNB VPB NWDIODE A=26.6695 P=32.33
c_153 VNB 0 7.12721e-20 $X=0 $Y=0
*
.include "sky130_fd_sc_lp__srsdfxtp_1.pxi.spice"
*
.ends
*
*
