* File: sky130_fd_sc_lp__o32ai_m.pxi.spice
* Created: Wed Sep  2 10:27:11 2020
* 
x_PM_SKY130_FD_SC_LP__O32AI_M%B1 N_B1_c_72_n N_B1_c_73_n N_B1_c_74_n N_B1_c_80_n
+ N_B1_c_81_n N_B1_c_75_n N_B1_M1007_g N_B1_M1001_g N_B1_c_76_n B1 B1 B1 B1 B1
+ N_B1_c_78_n PM_SKY130_FD_SC_LP__O32AI_M%B1
x_PM_SKY130_FD_SC_LP__O32AI_M%B2 N_B2_M1009_g N_B2_M1000_g N_B2_c_114_n
+ N_B2_c_119_n B2 B2 B2 B2 N_B2_c_116_n PM_SKY130_FD_SC_LP__O32AI_M%B2
x_PM_SKY130_FD_SC_LP__O32AI_M%A3 N_A3_M1006_g N_A3_M1008_g N_A3_c_154_n
+ N_A3_c_159_n A3 A3 A3 A3 N_A3_c_156_n PM_SKY130_FD_SC_LP__O32AI_M%A3
x_PM_SKY130_FD_SC_LP__O32AI_M%A2 N_A2_M1003_g N_A2_M1005_g N_A2_c_194_n
+ N_A2_c_199_n A2 A2 A2 A2 N_A2_c_196_n PM_SKY130_FD_SC_LP__O32AI_M%A2
x_PM_SKY130_FD_SC_LP__O32AI_M%A1 N_A1_M1002_g N_A1_c_235_n N_A1_M1004_g
+ N_A1_c_243_n N_A1_c_244_n N_A1_c_236_n N_A1_c_237_n N_A1_c_238_n N_A1_c_239_n
+ A1 A1 A1 A1 A1 N_A1_c_241_n PM_SKY130_FD_SC_LP__O32AI_M%A1
x_PM_SKY130_FD_SC_LP__O32AI_M%VPWR N_VPWR_M1001_s N_VPWR_M1002_d N_VPWR_c_276_n
+ N_VPWR_c_277_n N_VPWR_c_278_n N_VPWR_c_279_n VPWR N_VPWR_c_280_n
+ N_VPWR_c_275_n PM_SKY130_FD_SC_LP__O32AI_M%VPWR
x_PM_SKY130_FD_SC_LP__O32AI_M%Y N_Y_M1007_d N_Y_M1000_d N_Y_c_314_n N_Y_c_315_n
+ Y Y Y Y Y PM_SKY130_FD_SC_LP__O32AI_M%Y
x_PM_SKY130_FD_SC_LP__O32AI_M%A_66_82# N_A_66_82#_M1007_s N_A_66_82#_M1009_d
+ N_A_66_82#_M1003_d N_A_66_82#_c_364_n N_A_66_82#_c_365_n N_A_66_82#_c_366_n
+ N_A_66_82#_c_390_p N_A_66_82#_c_367_n PM_SKY130_FD_SC_LP__O32AI_M%A_66_82#
x_PM_SKY130_FD_SC_LP__O32AI_M%VGND N_VGND_M1006_d N_VGND_M1004_d N_VGND_c_397_n
+ N_VGND_c_398_n N_VGND_c_399_n VGND N_VGND_c_400_n N_VGND_c_401_n
+ N_VGND_c_402_n N_VGND_c_403_n N_VGND_c_404_n PM_SKY130_FD_SC_LP__O32AI_M%VGND
cc_1 VNB N_B1_c_72_n 0.00308084f $X=-0.19 $Y=-0.245 $X2=0.36 $Y2=2.24
cc_2 VNB N_B1_c_73_n 0.0297575f $X=-0.19 $Y=-0.245 $X2=0.675 $Y2=1.015
cc_3 VNB N_B1_c_74_n 0.0242726f $X=-0.19 $Y=-0.245 $X2=0.435 $Y2=1.015
cc_4 VNB N_B1_c_75_n 0.0182338f $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=0.94
cc_5 VNB N_B1_c_76_n 0.024983f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.61
cc_6 VNB B1 0.00919959f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_7 VNB N_B1_c_78_n 0.0382498f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.105
cc_8 VNB N_B2_M1009_g 0.0359061f $X=-0.19 $Y=-0.245 $X2=0.675 $Y2=1.015
cc_9 VNB N_B2_c_114_n 0.0112894f $X=-0.19 $Y=-0.245 $X2=0.82 $Y2=2.885
cc_10 VNB B2 0.00618848f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_B2_c_116_n 0.0168717f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A3_M1006_g 0.0295382f $X=-0.19 $Y=-0.245 $X2=0.675 $Y2=1.015
cc_13 VNB N_A3_c_154_n 0.0190404f $X=-0.19 $Y=-0.245 $X2=0.82 $Y2=2.885
cc_14 VNB A3 8.14036e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A3_c_156_n 0.0162214f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A2_M1003_g 0.0390674f $X=-0.19 $Y=-0.245 $X2=0.675 $Y2=1.015
cc_17 VNB N_A2_c_194_n 0.0123834f $X=-0.19 $Y=-0.245 $X2=0.82 $Y2=2.885
cc_18 VNB A2 0.0024827f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A2_c_196_n 0.0180423f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A1_c_235_n 0.0189261f $X=-0.19 $Y=-0.245 $X2=0.745 $Y2=2.315
cc_21 VNB N_A1_c_236_n 0.0382595f $X=-0.19 $Y=-0.245 $X2=0.82 $Y2=2.39
cc_22 VNB N_A1_c_237_n 0.0136665f $X=-0.19 $Y=-0.245 $X2=0.82 $Y2=2.885
cc_23 VNB N_A1_c_238_n 0.00308801f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A1_c_239_n 0.0199637f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.61
cc_25 VNB A1 0.0375654f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_26 VNB N_A1_c_241_n 0.0300924f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.105
cc_27 VNB N_VPWR_c_275_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0.255 $Y2=0.925
cc_28 VNB N_Y_c_314_n 0.006876f $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=0.94
cc_29 VNB N_Y_c_315_n 0.0109252f $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=0.62
cc_30 VNB N_A_66_82#_c_364_n 0.00805683f $X=-0.19 $Y=-0.245 $X2=0.82 $Y2=2.39
cc_31 VNB N_A_66_82#_c_365_n 0.0135005f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.61
cc_32 VNB N_A_66_82#_c_366_n 0.0079944f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_33 VNB N_A_66_82#_c_367_n 0.0189017f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_397_n 0.00503474f $X=-0.19 $Y=-0.245 $X2=0.75 $Y2=0.62
cc_35 VNB N_VGND_c_398_n 0.0163873f $X=-0.19 $Y=-0.245 $X2=0.82 $Y2=2.885
cc_36 VNB N_VGND_c_399_n 0.0217412f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.445
cc_37 VNB N_VGND_c_400_n 0.0445675f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_38 VNB N_VGND_c_401_n 0.0170996f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_402_n 0.22032f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.105
cc_40 VNB N_VGND_c_403_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0.255 $Y2=0.925
cc_41 VNB N_VGND_c_404_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0.255 $Y2=1.105
cc_42 VPB N_B1_c_72_n 0.0392062f $X=-0.19 $Y=1.655 $X2=0.36 $Y2=2.24
cc_43 VPB N_B1_c_80_n 0.0408668f $X=-0.19 $Y=1.655 $X2=0.745 $Y2=2.315
cc_44 VPB N_B1_c_81_n 0.011124f $X=-0.19 $Y=1.655 $X2=0.435 $Y2=2.315
cc_45 VPB N_B1_M1001_g 0.0300046f $X=-0.19 $Y=1.655 $X2=0.82 $Y2=2.885
cc_46 VPB B1 0.0332937f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_47 VPB N_B2_M1000_g 0.0426347f $X=-0.19 $Y=1.655 $X2=0.75 $Y2=0.94
cc_48 VPB N_B2_c_114_n 0.0127095f $X=-0.19 $Y=1.655 $X2=0.82 $Y2=2.885
cc_49 VPB N_B2_c_119_n 0.0178922f $X=-0.19 $Y=1.655 $X2=0.82 $Y2=2.885
cc_50 VPB B2 0.0106588f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_51 VPB N_A3_M1008_g 0.0514452f $X=-0.19 $Y=1.655 $X2=0.75 $Y2=0.94
cc_52 VPB N_A3_c_154_n 0.00402647f $X=-0.19 $Y=1.655 $X2=0.82 $Y2=2.885
cc_53 VPB N_A3_c_159_n 0.0190569f $X=-0.19 $Y=1.655 $X2=0.82 $Y2=2.885
cc_54 VPB A3 0.0053906f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_55 VPB N_A2_M1005_g 0.046543f $X=-0.19 $Y=1.655 $X2=0.75 $Y2=0.94
cc_56 VPB N_A2_c_194_n 0.013941f $X=-0.19 $Y=1.655 $X2=0.82 $Y2=2.885
cc_57 VPB N_A2_c_199_n 0.0191585f $X=-0.19 $Y=1.655 $X2=0.82 $Y2=2.885
cc_58 VPB A2 0.00657003f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_59 VPB N_A1_M1002_g 0.0331156f $X=-0.19 $Y=1.655 $X2=0.675 $Y2=1.015
cc_60 VPB N_A1_c_243_n 0.0405459f $X=-0.19 $Y=1.655 $X2=0.75 $Y2=0.62
cc_61 VPB N_A1_c_244_n 0.0132019f $X=-0.19 $Y=1.655 $X2=0.75 $Y2=0.62
cc_62 VPB N_A1_c_238_n 0.0393786f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_63 VPB A1 0.038314f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_64 VPB N_VPWR_c_276_n 0.0142813f $X=-0.19 $Y=1.655 $X2=0.75 $Y2=0.94
cc_65 VPB N_VPWR_c_277_n 0.00485511f $X=-0.19 $Y=1.655 $X2=0.75 $Y2=0.62
cc_66 VPB N_VPWR_c_278_n 0.0142813f $X=-0.19 $Y=1.655 $X2=0.82 $Y2=2.885
cc_67 VPB N_VPWR_c_279_n 0.00485511f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_280_n 0.0609464f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_69 VPB N_VPWR_c_275_n 0.0512397f $X=-0.19 $Y=1.655 $X2=0.255 $Y2=0.925
cc_70 VPB N_Y_c_315_n 0.018559f $X=-0.19 $Y=1.655 $X2=0.75 $Y2=0.62
cc_71 VPB Y 0.0281531f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.61
cc_72 N_B1_c_75_n N_B2_M1009_g 0.0223414f $X=0.75 $Y=0.94 $X2=0 $Y2=0
cc_73 N_B1_c_78_n N_B2_M1009_g 0.00158523f $X=0.27 $Y=1.105 $X2=0 $Y2=0
cc_74 N_B1_c_72_n N_B2_M1000_g 0.00150624f $X=0.36 $Y=2.24 $X2=0 $Y2=0
cc_75 N_B1_c_80_n N_B2_M1000_g 0.0628087f $X=0.745 $Y=2.315 $X2=0 $Y2=0
cc_76 N_B1_c_76_n N_B2_c_114_n 0.00375903f $X=0.27 $Y=1.61 $X2=0 $Y2=0
cc_77 N_B1_c_72_n N_B2_c_119_n 0.00375903f $X=0.36 $Y=2.24 $X2=0 $Y2=0
cc_78 N_B1_c_80_n B2 0.0016189f $X=0.745 $Y=2.315 $X2=0 $Y2=0
cc_79 N_B1_c_78_n N_B2_c_116_n 0.00375903f $X=0.27 $Y=1.105 $X2=0 $Y2=0
cc_80 N_B1_c_81_n N_VPWR_c_277_n 0.00404181f $X=0.435 $Y=2.315 $X2=0 $Y2=0
cc_81 N_B1_M1001_g N_VPWR_c_277_n 0.00685007f $X=0.82 $Y=2.885 $X2=0 $Y2=0
cc_82 B1 N_VPWR_c_277_n 0.00491962f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_83 N_B1_M1001_g N_VPWR_c_280_n 0.00372967f $X=0.82 $Y=2.885 $X2=0 $Y2=0
cc_84 N_B1_M1001_g N_VPWR_c_275_n 0.00669081f $X=0.82 $Y=2.885 $X2=0 $Y2=0
cc_85 B1 N_VPWR_c_275_n 0.00476695f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_86 N_B1_c_73_n N_Y_c_314_n 0.0036213f $X=0.675 $Y=1.015 $X2=0 $Y2=0
cc_87 N_B1_c_75_n N_Y_c_314_n 0.0155643f $X=0.75 $Y=0.94 $X2=0 $Y2=0
cc_88 B1 N_Y_c_314_n 0.00890083f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_89 N_B1_c_73_n N_Y_c_315_n 0.00789973f $X=0.675 $Y=1.015 $X2=0 $Y2=0
cc_90 N_B1_c_80_n N_Y_c_315_n 0.0129551f $X=0.745 $Y=2.315 $X2=0 $Y2=0
cc_91 N_B1_M1001_g N_Y_c_315_n 0.0182989f $X=0.82 $Y=2.885 $X2=0 $Y2=0
cc_92 B1 N_Y_c_315_n 0.0695984f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_93 N_B1_c_78_n N_Y_c_315_n 0.00887328f $X=0.27 $Y=1.105 $X2=0 $Y2=0
cc_94 N_B1_M1001_g Y 0.00892919f $X=0.82 $Y=2.885 $X2=0 $Y2=0
cc_95 N_B1_c_75_n N_A_66_82#_c_364_n 0.0116881f $X=0.75 $Y=0.94 $X2=0 $Y2=0
cc_96 N_B1_c_74_n N_A_66_82#_c_367_n 0.00979176f $X=0.435 $Y=1.015 $X2=0 $Y2=0
cc_97 N_B1_c_75_n N_A_66_82#_c_367_n 0.00142375f $X=0.75 $Y=0.94 $X2=0 $Y2=0
cc_98 B1 N_A_66_82#_c_367_n 0.00523932f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_99 N_B1_c_75_n N_VGND_c_400_n 9.21892e-19 $X=0.75 $Y=0.94 $X2=0 $Y2=0
cc_100 B1 N_VGND_c_402_n 0.00544513f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_101 N_B2_M1009_g N_A3_M1006_g 0.025475f $X=1.18 $Y=0.62 $X2=0 $Y2=0
cc_102 N_B2_c_119_n N_A3_M1008_g 0.0443528f $X=1.09 $Y=2 $X2=0 $Y2=0
cc_103 B2 N_A3_M1008_g 0.00363888f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_104 N_B2_c_116_n N_A3_c_154_n 0.0139197f $X=1.09 $Y=1.495 $X2=0 $Y2=0
cc_105 N_B2_c_114_n N_A3_c_159_n 0.0139197f $X=1.09 $Y=1.835 $X2=0 $Y2=0
cc_106 N_B2_M1009_g A3 0.00145893f $X=1.18 $Y=0.62 $X2=0 $Y2=0
cc_107 B2 A3 0.0707075f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_108 N_B2_M1009_g N_A3_c_156_n 0.0139197f $X=1.18 $Y=0.62 $X2=0 $Y2=0
cc_109 B2 N_A3_c_156_n 0.00439653f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_110 N_B2_M1000_g N_VPWR_c_280_n 0.00373071f $X=1.18 $Y=2.885 $X2=0 $Y2=0
cc_111 N_B2_M1000_g N_VPWR_c_275_n 0.00531889f $X=1.18 $Y=2.885 $X2=0 $Y2=0
cc_112 N_B2_M1009_g N_Y_c_314_n 0.00703622f $X=1.18 $Y=0.62 $X2=0 $Y2=0
cc_113 B2 N_Y_c_314_n 0.00971283f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_114 N_B2_c_116_n N_Y_c_314_n 0.00363823f $X=1.09 $Y=1.495 $X2=0 $Y2=0
cc_115 N_B2_M1009_g N_Y_c_315_n 0.00426241f $X=1.18 $Y=0.62 $X2=0 $Y2=0
cc_116 N_B2_M1000_g N_Y_c_315_n 0.00223717f $X=1.18 $Y=2.885 $X2=0 $Y2=0
cc_117 B2 N_Y_c_315_n 0.0924254f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_118 N_B2_c_116_n N_Y_c_315_n 0.00672467f $X=1.09 $Y=1.495 $X2=0 $Y2=0
cc_119 N_B2_M1000_g Y 0.0114587f $X=1.18 $Y=2.885 $X2=0 $Y2=0
cc_120 N_B2_c_119_n Y 0.00240463f $X=1.09 $Y=2 $X2=0 $Y2=0
cc_121 B2 Y 0.0216255f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_122 N_B2_M1009_g N_A_66_82#_c_364_n 0.0132483f $X=1.18 $Y=0.62 $X2=0 $Y2=0
cc_123 N_B2_M1009_g N_A_66_82#_c_366_n 0.00136047f $X=1.18 $Y=0.62 $X2=0 $Y2=0
cc_124 N_B2_M1009_g N_VGND_c_400_n 9.21892e-19 $X=1.18 $Y=0.62 $X2=0 $Y2=0
cc_125 N_A3_M1006_g N_A2_M1003_g 0.0237503f $X=1.61 $Y=0.62 $X2=0 $Y2=0
cc_126 A3 N_A2_M1003_g 0.00228558f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_127 N_A3_c_156_n N_A2_M1003_g 0.0136684f $X=1.63 $Y=1.375 $X2=0 $Y2=0
cc_128 N_A3_c_159_n N_A2_c_194_n 0.0136684f $X=1.63 $Y=1.88 $X2=0 $Y2=0
cc_129 N_A3_M1008_g N_A2_c_199_n 0.0516938f $X=1.61 $Y=2.885 $X2=0 $Y2=0
cc_130 A3 N_A2_c_199_n 0.00421755f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_131 N_A3_M1008_g A2 6.41364e-19 $X=1.61 $Y=2.885 $X2=0 $Y2=0
cc_132 A3 A2 0.0572718f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_133 N_A3_c_156_n A2 0.00214301f $X=1.63 $Y=1.375 $X2=0 $Y2=0
cc_134 N_A3_c_154_n N_A2_c_196_n 0.0136684f $X=1.63 $Y=1.715 $X2=0 $Y2=0
cc_135 N_A3_M1008_g N_VPWR_c_280_n 0.00373071f $X=1.61 $Y=2.885 $X2=0 $Y2=0
cc_136 N_A3_M1008_g N_VPWR_c_275_n 0.00561503f $X=1.61 $Y=2.885 $X2=0 $Y2=0
cc_137 N_A3_M1006_g N_Y_c_314_n 2.87482e-19 $X=1.61 $Y=0.62 $X2=0 $Y2=0
cc_138 N_A3_M1008_g Y 0.0131409f $X=1.61 $Y=2.885 $X2=0 $Y2=0
cc_139 A3 Y 0.0167774f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_140 N_A3_M1006_g N_A_66_82#_c_364_n 0.00111918f $X=1.61 $Y=0.62 $X2=0 $Y2=0
cc_141 N_A3_M1006_g N_A_66_82#_c_365_n 0.0119653f $X=1.61 $Y=0.62 $X2=0 $Y2=0
cc_142 A3 N_A_66_82#_c_365_n 0.0138013f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_143 N_A3_c_156_n N_A_66_82#_c_365_n 0.00307639f $X=1.63 $Y=1.375 $X2=0 $Y2=0
cc_144 N_A3_c_156_n N_A_66_82#_c_366_n 0.00159171f $X=1.63 $Y=1.375 $X2=0 $Y2=0
cc_145 N_A3_M1006_g N_VGND_c_397_n 0.00490157f $X=1.61 $Y=0.62 $X2=0 $Y2=0
cc_146 N_A3_M1006_g N_VGND_c_400_n 0.00529112f $X=1.61 $Y=0.62 $X2=0 $Y2=0
cc_147 N_A3_M1006_g N_VGND_c_402_n 0.00518865f $X=1.61 $Y=0.62 $X2=0 $Y2=0
cc_148 N_A2_M1003_g N_A1_c_235_n 0.0208929f $X=2.08 $Y=0.62 $X2=0 $Y2=0
cc_149 N_A2_M1005_g N_A1_c_244_n 0.0639066f $X=2.08 $Y=2.885 $X2=0 $Y2=0
cc_150 A2 N_A1_c_244_n 0.00281813f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_151 N_A2_M1005_g N_A1_c_238_n 0.00179839f $X=2.08 $Y=2.885 $X2=0 $Y2=0
cc_152 N_A2_c_199_n N_A1_c_238_n 0.00511802f $X=2.17 $Y=2 $X2=0 $Y2=0
cc_153 A2 N_A1_c_238_n 0.00106794f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_154 N_A2_c_194_n N_A1_c_239_n 0.00511802f $X=2.17 $Y=1.835 $X2=0 $Y2=0
cc_155 A2 A1 0.0331087f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_156 N_A2_c_196_n A1 0.00257337f $X=2.17 $Y=1.495 $X2=0 $Y2=0
cc_157 N_A2_M1003_g N_A1_c_241_n 0.00227382f $X=2.08 $Y=0.62 $X2=0 $Y2=0
cc_158 A2 N_A1_c_241_n 0.00331116f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_159 N_A2_c_196_n N_A1_c_241_n 0.00511802f $X=2.17 $Y=1.495 $X2=0 $Y2=0
cc_160 N_A2_M1005_g N_VPWR_c_280_n 0.00373071f $X=2.08 $Y=2.885 $X2=0 $Y2=0
cc_161 N_A2_M1005_g N_VPWR_c_275_n 0.0054198f $X=2.08 $Y=2.885 $X2=0 $Y2=0
cc_162 N_A2_M1005_g Y 0.0180916f $X=2.08 $Y=2.885 $X2=0 $Y2=0
cc_163 N_A2_c_199_n Y 0.00240463f $X=2.17 $Y=2 $X2=0 $Y2=0
cc_164 A2 Y 0.0139906f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_165 N_A2_M1003_g N_A_66_82#_c_365_n 0.0134521f $X=2.08 $Y=0.62 $X2=0 $Y2=0
cc_166 A2 N_A_66_82#_c_365_n 0.0121889f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_167 N_A2_c_196_n N_A_66_82#_c_365_n 0.00362437f $X=2.17 $Y=1.495 $X2=0 $Y2=0
cc_168 N_A2_M1003_g N_VGND_c_397_n 0.00670336f $X=2.08 $Y=0.62 $X2=0 $Y2=0
cc_169 N_A2_M1003_g N_VGND_c_398_n 0.00529112f $X=2.08 $Y=0.62 $X2=0 $Y2=0
cc_170 N_A2_M1003_g N_VGND_c_399_n 6.89375e-19 $X=2.08 $Y=0.62 $X2=0 $Y2=0
cc_171 N_A2_M1003_g N_VGND_c_402_n 0.00518865f $X=2.08 $Y=0.62 $X2=0 $Y2=0
cc_172 N_A1_M1002_g N_VPWR_c_279_n 0.00589957f $X=2.44 $Y=2.885 $X2=0 $Y2=0
cc_173 N_A1_c_243_n N_VPWR_c_279_n 3.19995e-19 $X=2.81 $Y=2.315 $X2=0 $Y2=0
cc_174 A1 N_VPWR_c_279_n 0.0105102f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_175 N_A1_M1002_g N_VPWR_c_280_n 0.00373071f $X=2.44 $Y=2.885 $X2=0 $Y2=0
cc_176 N_A1_M1002_g N_VPWR_c_275_n 0.00669127f $X=2.44 $Y=2.885 $X2=0 $Y2=0
cc_177 A1 N_VPWR_c_275_n 0.00584664f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_178 N_A1_M1002_g Y 0.0220309f $X=2.44 $Y=2.885 $X2=0 $Y2=0
cc_179 N_A1_c_243_n Y 0.00690984f $X=2.81 $Y=2.315 $X2=0 $Y2=0
cc_180 N_A1_c_235_n N_A_66_82#_c_365_n 0.00250601f $X=2.51 $Y=0.94 $X2=0 $Y2=0
cc_181 A1 N_A_66_82#_c_365_n 0.00591572f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_182 N_A1_c_235_n N_VGND_c_397_n 6.56138e-19 $X=2.51 $Y=0.94 $X2=0 $Y2=0
cc_183 N_A1_c_235_n N_VGND_c_398_n 0.00455951f $X=2.51 $Y=0.94 $X2=0 $Y2=0
cc_184 N_A1_c_235_n N_VGND_c_399_n 0.00994346f $X=2.51 $Y=0.94 $X2=0 $Y2=0
cc_185 N_A1_c_236_n N_VGND_c_399_n 0.0103638f $X=2.81 $Y=1.015 $X2=0 $Y2=0
cc_186 N_A1_c_235_n N_VGND_c_402_n 0.00447788f $X=2.51 $Y=0.94 $X2=0 $Y2=0
cc_187 A1 N_VGND_c_402_n 0.0123416f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_188 N_VPWR_c_275_n A_179_535# 0.00173577f $X=3.12 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_189 N_VPWR_c_275_n N_Y_M1000_d 0.00231436f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_190 N_VPWR_M1001_s N_Y_c_315_n 0.00800578f $X=0.245 $Y=2.675 $X2=0 $Y2=0
cc_191 N_VPWR_c_277_n N_Y_c_315_n 0.0168863f $X=0.37 $Y=2.95 $X2=0 $Y2=0
cc_192 N_VPWR_c_280_n N_Y_c_315_n 0.00748325f $X=2.905 $Y=3.33 $X2=0 $Y2=0
cc_193 N_VPWR_c_275_n N_Y_c_315_n 0.00669622f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_194 N_VPWR_M1002_d Y 0.0096436f $X=2.515 $Y=2.675 $X2=0 $Y2=0
cc_195 N_VPWR_c_279_n Y 0.0168078f $X=2.99 $Y=2.95 $X2=0 $Y2=0
cc_196 N_VPWR_c_280_n Y 0.0735372f $X=2.905 $Y=3.33 $X2=0 $Y2=0
cc_197 N_VPWR_c_275_n Y 0.0661651f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_198 N_VPWR_c_275_n A_337_535# 0.00264498f $X=3.12 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_199 N_VPWR_c_275_n A_431_535# 0.00173577f $X=3.12 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_200 A_179_535# Y 0.00107385f $X=0.895 $Y=2.675 $X2=0 $Y2=0
cc_201 Y A_337_535# 0.00230429f $X=2.555 $Y=2.69 $X2=-0.19 $Y2=-0.245
cc_202 Y A_431_535# 0.00107385f $X=2.555 $Y=2.69 $X2=-0.19 $Y2=-0.245
cc_203 N_Y_M1007_d N_A_66_82#_c_364_n 0.00180746f $X=0.825 $Y=0.41 $X2=0 $Y2=0
cc_204 N_Y_c_314_n N_A_66_82#_c_364_n 0.0192361f $X=0.74 $Y=1.01 $X2=0 $Y2=0
cc_205 N_Y_c_314_n N_A_66_82#_c_366_n 0.0136086f $X=0.74 $Y=1.01 $X2=0 $Y2=0
cc_206 N_A_66_82#_c_365_n N_VGND_M1006_d 0.00220794f $X=2.19 $Y=0.905 $X2=-0.19
+ $Y2=-0.245
cc_207 N_A_66_82#_c_364_n N_VGND_c_397_n 0.0123841f $X=1.31 $Y=0.355 $X2=0 $Y2=0
cc_208 N_A_66_82#_c_365_n N_VGND_c_397_n 0.0160971f $X=2.19 $Y=0.905 $X2=0 $Y2=0
cc_209 N_A_66_82#_c_390_p N_VGND_c_398_n 0.00438316f $X=2.295 $Y=0.685 $X2=0
+ $Y2=0
cc_210 N_A_66_82#_c_364_n N_VGND_c_400_n 0.0531105f $X=1.31 $Y=0.355 $X2=0 $Y2=0
cc_211 N_A_66_82#_c_367_n N_VGND_c_400_n 0.0206108f $X=0.455 $Y=0.355 $X2=0
+ $Y2=0
cc_212 N_A_66_82#_c_364_n N_VGND_c_402_n 0.0330503f $X=1.31 $Y=0.355 $X2=0 $Y2=0
cc_213 N_A_66_82#_c_365_n N_VGND_c_402_n 0.0127863f $X=2.19 $Y=0.905 $X2=0 $Y2=0
cc_214 N_A_66_82#_c_390_p N_VGND_c_402_n 0.00609927f $X=2.295 $Y=0.685 $X2=0
+ $Y2=0
cc_215 N_A_66_82#_c_367_n N_VGND_c_402_n 0.0124745f $X=0.455 $Y=0.355 $X2=0
+ $Y2=0
