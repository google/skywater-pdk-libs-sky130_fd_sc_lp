* File: sky130_fd_sc_lp__sdfstp_4.pex.spice
* Created: Fri Aug 28 11:29:51 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__SDFSTP_4%SCD 3 5 7 11 14 15 16 20 21
r36 20 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.385
+ $Y=1.29 $X2=0.385 $Y2=1.29
r37 15 16 9.51718 $w=4.63e-07 $l=3.7e-07 $layer=LI1_cond $X=0.317 $Y=1.295
+ $X2=0.317 $Y2=1.665
r38 15 21 0.128611 $w=4.63e-07 $l=5e-09 $layer=LI1_cond $X=0.317 $Y=1.295
+ $X2=0.317 $Y2=1.29
r39 13 20 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.385 $Y=1.63
+ $X2=0.385 $Y2=1.29
r40 13 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.385 $Y=1.63
+ $X2=0.385 $Y2=1.795
r41 9 20 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=0.385 $Y=1.275
+ $X2=0.385 $Y2=1.29
r42 9 11 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=0.385 $Y=1.2
+ $X2=0.655 $Y2=1.2
r43 5 11 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.655 $Y=1.125
+ $X2=0.655 $Y2=1.2
r44 5 7 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.655 $Y=1.125
+ $X2=0.655 $Y2=0.805
r45 3 14 471.745 $w=1.5e-07 $l=9.2e-07 $layer=POLY_cond $X=0.475 $Y=2.715
+ $X2=0.475 $Y2=1.795
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSTP_4%D 3 9 12 13 14 15 16 17 25 27 35 36
c54 25 0 1.1672e-19 $X=1.355 $Y=2.07
r55 25 28 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.355 $Y=2.07
+ $X2=1.355 $Y2=2.235
r56 25 27 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.355 $Y=2.07
+ $X2=1.355 $Y2=1.905
r57 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.355
+ $Y=2.07 $X2=1.355 $Y2=2.07
r58 16 17 19.4096 $w=2.83e-07 $l=4.8e-07 $layer=LI1_cond $X=1.68 $Y=2.012
+ $X2=2.16 $Y2=2.012
r59 16 26 13.1419 $w=2.83e-07 $l=3.25e-07 $layer=LI1_cond $X=1.68 $Y=2.012
+ $X2=1.355 $Y2=2.012
r60 15 26 6.26767 $w=2.83e-07 $l=1.55e-07 $layer=LI1_cond $X=1.2 $Y=2.012
+ $X2=1.355 $Y2=2.012
r61 15 36 13.6676 $w=2.83e-07 $l=3.38e-07 $layer=LI1_cond $X=1.2 $Y=2.012
+ $X2=0.862 $Y2=2.012
r62 14 36 4.04366 $w=2.83e-07 $l=1e-07 $layer=LI1_cond $X=0.762 $Y=2.012
+ $X2=0.862 $Y2=2.012
r63 14 35 1.69834 $w=2.83e-07 $l=4.2e-08 $layer=LI1_cond $X=0.762 $Y=2.012
+ $X2=0.72 $Y2=2.012
r64 14 35 2.2525 $w=2.18e-07 $l=4.3e-08 $layer=LI1_cond $X=0.677 $Y=2.045
+ $X2=0.72 $Y2=2.045
r65 13 14 22.8917 $w=2.18e-07 $l=4.37e-07 $layer=LI1_cond $X=0.24 $Y=2.045
+ $X2=0.677 $Y2=2.045
r66 12 27 199.979 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=1.415 $Y=1.515
+ $X2=1.415 $Y2=1.905
r67 11 12 58.3064 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=1.43 $Y=1.365
+ $X2=1.43 $Y2=1.515
r68 9 11 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=1.445 $Y=0.805
+ $X2=1.445 $Y2=1.365
r69 3 28 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.265 $Y=2.715
+ $X2=1.265 $Y2=2.235
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSTP_4%A_346_93# 1 2 9 13 15 17 19 26 27 28 29 32
r75 30 32 20.8326 $w=2.58e-07 $l=4.7e-07 $layer=LI1_cond $X=3.495 $Y=2.1
+ $X2=3.495 $Y2=2.57
r76 28 30 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=3.365 $Y=2.015
+ $X2=3.495 $Y2=2.1
r77 28 29 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=3.365 $Y=2.015
+ $X2=3.025 $Y2=2.015
r78 26 27 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.86 $Y=1.4
+ $X2=2.86 $Y2=1.4
r79 24 29 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=2.895 $Y=1.93
+ $X2=3.025 $Y2=2.015
r80 24 26 23.4921 $w=2.58e-07 $l=5.3e-07 $layer=LI1_cond $X=2.895 $Y=1.93
+ $X2=2.895 $Y2=1.4
r81 23 26 19.0596 $w=2.58e-07 $l=4.3e-07 $layer=LI1_cond $X=2.895 $Y=0.97
+ $X2=2.895 $Y2=1.4
r82 19 23 6.94204 $w=3.3e-07 $l=2.20624e-07 $layer=LI1_cond $X=2.765 $Y=0.805
+ $X2=2.895 $Y2=0.97
r83 19 21 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=2.765 $Y=0.805
+ $X2=2.45 $Y2=0.805
r84 18 27 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=2.86 $Y=1.755
+ $X2=2.86 $Y2=1.4
r85 16 17 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.88 $Y=1.83
+ $X2=1.805 $Y2=1.83
r86 15 18 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=2.695 $Y=1.83
+ $X2=2.86 $Y2=1.755
r87 15 16 417.904 $w=1.5e-07 $l=8.15e-07 $layer=POLY_cond $X=2.695 $Y=1.83
+ $X2=1.88 $Y2=1.83
r88 11 17 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.805 $Y=1.905
+ $X2=1.805 $Y2=1.83
r89 11 13 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=1.805 $Y=1.905
+ $X2=1.805 $Y2=2.715
r90 7 17 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.805 $Y=1.755
+ $X2=1.805 $Y2=1.83
r91 7 9 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=1.805 $Y=1.755
+ $X2=1.805 $Y2=0.805
r92 2 32 600 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_PDIFF $count=1 $X=3.32
+ $Y=2.405 $X2=3.46 $Y2=2.57
r93 1 21 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.31
+ $Y=0.595 $X2=2.45 $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSTP_4%SCE 3 8 9 10 13 15 17 19 23 26 28 31 34 35
+ 36 37 38 39 40 46
r101 39 40 16.4002 $w=2.58e-07 $l=3.7e-07 $layer=LI1_cond $X=3.565 $Y=1.295
+ $X2=3.565 $Y2=1.665
r102 38 39 16.4002 $w=2.58e-07 $l=3.7e-07 $layer=LI1_cond $X=3.565 $Y=0.925
+ $X2=3.565 $Y2=1.295
r103 37 38 16.4002 $w=2.58e-07 $l=3.7e-07 $layer=LI1_cond $X=3.565 $Y=0.555
+ $X2=3.565 $Y2=0.925
r104 37 46 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.6
+ $Y=0.635 $X2=3.6 $Y2=0.635
r105 35 46 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=3.6 $Y=0.975
+ $X2=3.6 $Y2=0.635
r106 35 36 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.6 $Y=0.975
+ $X2=3.6 $Y2=1.14
r107 34 46 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.6 $Y=0.47
+ $X2=3.6 $Y2=0.635
r108 29 31 135.883 $w=1.5e-07 $l=2.65e-07 $layer=POLY_cond $X=3.245 $Y=2.22
+ $X2=3.51 $Y2=2.22
r109 24 26 56.4043 $w=1.5e-07 $l=1.1e-07 $layer=POLY_cond $X=0.905 $Y=1.59
+ $X2=1.015 $Y2=1.59
r110 23 31 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.51 $Y=2.145
+ $X2=3.51 $Y2=2.22
r111 23 36 515.33 $w=1.5e-07 $l=1.005e-06 $layer=POLY_cond $X=3.51 $Y=2.145
+ $X2=3.51 $Y2=1.14
r112 20 34 110.245 $w=1.5e-07 $l=2.15e-07 $layer=POLY_cond $X=3.51 $Y=0.255
+ $X2=3.51 $Y2=0.47
r113 17 29 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.245 $Y=2.295
+ $X2=3.245 $Y2=2.22
r114 17 19 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=3.245 $Y=2.295
+ $X2=3.245 $Y2=2.725
r115 16 28 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.31 $Y=0.18
+ $X2=2.235 $Y2=0.18
r116 15 20 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.435 $Y=0.18
+ $X2=3.51 $Y2=0.255
r117 15 16 576.862 $w=1.5e-07 $l=1.125e-06 $layer=POLY_cond $X=3.435 $Y=0.18
+ $X2=2.31 $Y2=0.18
r118 11 28 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.235 $Y=0.255
+ $X2=2.235 $Y2=0.18
r119 11 13 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=2.235 $Y=0.255
+ $X2=2.235 $Y2=0.805
r120 9 28 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.16 $Y=0.18
+ $X2=2.235 $Y2=0.18
r121 9 10 548.66 $w=1.5e-07 $l=1.07e-06 $layer=POLY_cond $X=2.16 $Y=0.18
+ $X2=1.09 $Y2=0.18
r122 6 26 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.015 $Y=1.515
+ $X2=1.015 $Y2=1.59
r123 6 8 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=1.015 $Y=1.515
+ $X2=1.015 $Y2=0.805
r124 5 10 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.015 $Y=0.255
+ $X2=1.09 $Y2=0.18
r125 5 8 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=1.015 $Y=0.255
+ $X2=1.015 $Y2=0.805
r126 1 24 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.905 $Y=1.665
+ $X2=0.905 $Y2=1.59
r127 1 3 538.404 $w=1.5e-07 $l=1.05e-06 $layer=POLY_cond $X=0.905 $Y=1.665
+ $X2=0.905 $Y2=2.715
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSTP_4%CLK 1 3 7 11 12 13 14 19
r45 19 20 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.3
+ $Y=1.005 $X2=4.3 $Y2=1.005
r46 13 14 7.6965 $w=5.73e-07 $l=3.7e-07 $layer=LI1_cond $X=4.492 $Y=1.295
+ $X2=4.492 $Y2=1.665
r47 13 20 6.0324 $w=5.73e-07 $l=2.9e-07 $layer=LI1_cond $X=4.492 $Y=1.295
+ $X2=4.492 $Y2=1.005
r48 12 20 1.66411 $w=5.73e-07 $l=8e-08 $layer=LI1_cond $X=4.492 $Y=0.925
+ $X2=4.492 $Y2=1.005
r49 11 19 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=4.3 $Y=1.345 $X2=4.3
+ $Y2=1.005
r50 10 19 38.6168 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.3 $Y=0.84 $X2=4.3
+ $Y2=1.005
r51 7 10 176.904 $w=1.5e-07 $l=3.45e-07 $layer=POLY_cond $X=4.32 $Y=0.495
+ $X2=4.32 $Y2=0.84
r52 1 11 37.5318 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.3 $Y=1.51 $X2=4.3
+ $Y2=1.345
r53 1 3 648.649 $w=1.5e-07 $l=1.265e-06 $layer=POLY_cond $X=4.3 $Y=1.51 $X2=4.3
+ $Y2=2.775
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSTP_4%A_961_491# 1 2 9 13 17 21 23 27 29 32 35 38
+ 41 42 43 45 46 47 49 51 52 57 59 61 63 66 70
c183 61 0 9.96682e-20 $X=9.525 $Y=1.93
c184 59 0 2.18911e-19 $X=5.845 $Y=2.935
c185 51 0 1.49949e-19 $X=8.12 $Y=1.88
c186 9 0 7.13856e-20 $X=5.98 $Y=2.525
r187 62 70 34.9723 $w=3.3e-07 $l=2e-07 $layer=POLY_cond $X=9.525 $Y=1.93
+ $X2=9.725 $Y2=1.93
r188 61 63 9.26861 $w=2.18e-07 $l=1.65e-07 $layer=LI1_cond $X=9.525 $Y=1.905
+ $X2=9.36 $Y2=1.905
r189 61 62 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.525
+ $Y=1.93 $X2=9.525 $Y2=1.93
r190 52 55 7.44286 $w=2.38e-07 $l=1.55e-07 $layer=LI1_cond $X=4.95 $Y=0.34
+ $X2=4.95 $Y2=0.495
r191 51 63 80.8984 $w=1.68e-07 $l=1.24e-06 $layer=LI1_cond $X=8.12 $Y=1.88
+ $X2=9.36 $Y2=1.88
r192 48 51 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.035 $Y=1.965
+ $X2=8.12 $Y2=1.88
r193 48 49 53.4973 $w=1.68e-07 $l=8.2e-07 $layer=LI1_cond $X=8.035 $Y=1.965
+ $X2=8.035 $Y2=2.785
r194 46 49 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.95 $Y=2.87
+ $X2=8.035 $Y2=2.785
r195 46 47 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=7.95 $Y=2.87
+ $X2=7.42 $Y2=2.87
r196 45 47 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.335 $Y=2.785
+ $X2=7.42 $Y2=2.87
r197 44 45 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=7.335 $Y=2.265
+ $X2=7.335 $Y2=2.785
r198 42 44 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.25 $Y=2.18
+ $X2=7.335 $Y2=2.265
r199 42 43 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=7.25 $Y=2.18
+ $X2=6.72 $Y2=2.18
r200 40 43 6.82373 $w=1.7e-07 $l=1.25499e-07 $layer=LI1_cond $X=6.63 $Y=2.265
+ $X2=6.72 $Y2=2.18
r201 40 41 33.2727 $w=1.78e-07 $l=5.4e-07 $layer=LI1_cond $X=6.63 $Y=2.265
+ $X2=6.63 $Y2=2.805
r202 39 59 3.40559 $w=2.75e-07 $l=8.74643e-08 $layer=LI1_cond $X=5.93 $Y=2.94
+ $X2=5.845 $Y2=2.935
r203 38 41 7.17723 $w=2.7e-07 $l=1.74284e-07 $layer=LI1_cond $X=6.54 $Y=2.94
+ $X2=6.63 $Y2=2.805
r204 38 39 26.0367 $w=2.68e-07 $l=6.1e-07 $layer=LI1_cond $X=6.54 $Y=2.94
+ $X2=5.93 $Y2=2.94
r205 36 57 56.7594 $w=1.68e-07 $l=8.7e-07 $layer=LI1_cond $X=5.935 $Y=0.425
+ $X2=5.935 $Y2=1.295
r206 35 59 3.11956 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=5.845 $Y=2.795
+ $X2=5.845 $Y2=2.935
r207 35 58 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=5.845 $Y=2.795
+ $X2=5.845 $Y2=1.965
r208 33 66 11.1804 $w=5.82e-07 $l=1.35e-07 $layer=POLY_cond $X=5.845 $Y=1.63
+ $X2=5.98 $Y2=1.63
r209 32 33 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.845
+ $Y=1.46 $X2=5.845 $Y2=1.46
r210 30 58 7.14225 $w=2.58e-07 $l=1.3e-07 $layer=LI1_cond $X=5.89 $Y=1.835
+ $X2=5.89 $Y2=1.965
r211 30 32 16.6218 $w=2.58e-07 $l=3.75e-07 $layer=LI1_cond $X=5.89 $Y=1.835
+ $X2=5.89 $Y2=1.46
r212 29 57 7.14225 $w=2.58e-07 $l=1.3e-07 $layer=LI1_cond $X=5.89 $Y=1.425
+ $X2=5.89 $Y2=1.295
r213 29 32 1.55137 $w=2.58e-07 $l=3.5e-08 $layer=LI1_cond $X=5.89 $Y=1.425
+ $X2=5.89 $Y2=1.46
r214 28 52 2.75731 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=5.07 $Y=0.34
+ $X2=4.95 $Y2=0.34
r215 27 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.85 $Y=0.34
+ $X2=5.935 $Y2=0.425
r216 27 28 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=5.85 $Y=0.34
+ $X2=5.07 $Y2=0.34
r217 23 59 3.40559 $w=2.75e-07 $l=8.5e-08 $layer=LI1_cond $X=5.76 $Y=2.935
+ $X2=5.845 $Y2=2.935
r218 23 25 33.5443 $w=2.78e-07 $l=8.15e-07 $layer=LI1_cond $X=5.76 $Y=2.935
+ $X2=4.945 $Y2=2.935
r219 19 70 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.725 $Y=2.095
+ $X2=9.725 $Y2=1.93
r220 19 21 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=9.725 $Y=2.095
+ $X2=9.725 $Y2=2.525
r221 15 70 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.725 $Y=1.765
+ $X2=9.725 $Y2=1.93
r222 15 17 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=9.725 $Y=1.765
+ $X2=9.725 $Y2=0.945
r223 11 66 43.0653 $w=5.82e-07 $l=6.66783e-07 $layer=POLY_cond $X=6.5 $Y=1.295
+ $X2=5.98 $Y2=1.63
r224 11 13 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=6.5 $Y=1.295
+ $X2=6.5 $Y2=0.615
r225 7 66 35.2868 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=5.98 $Y=1.965
+ $X2=5.98 $Y2=1.63
r226 7 9 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=5.98 $Y=1.965
+ $X2=5.98 $Y2=2.525
r227 2 25 600 $w=1.7e-07 $l=5.20312e-07 $layer=licon1_PDIFF $count=1 $X=4.805
+ $Y=2.455 $X2=4.945 $Y2=2.91
r228 1 55 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=4.825
+ $Y=0.285 $X2=4.965 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSTP_4%A_1339_331# 1 2 9 13 16 19 21 24 28 31 36
+ 39
r69 26 28 30.6459 $w=1.88e-07 $l=5.25e-07 $layer=LI1_cond $X=7.685 $Y=1.925
+ $X2=7.685 $Y2=2.45
r70 24 39 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.95 $Y=1.1
+ $X2=6.95 $Y2=0.935
r71 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.95
+ $Y=1.1 $X2=6.95 $Y2=1.1
r72 21 31 9.74833 $w=1.88e-07 $l=1.67e-07 $layer=LI1_cond $X=7.69 $Y=1.067
+ $X2=7.69 $Y2=0.9
r73 21 23 31.6309 $w=2.33e-07 $l=6.45e-07 $layer=LI1_cond $X=7.595 $Y=1.067
+ $X2=6.95 $Y2=1.067
r74 19 37 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.86 $Y=1.82
+ $X2=6.86 $Y2=1.985
r75 19 36 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.86 $Y=1.82
+ $X2=6.86 $Y2=1.655
r76 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.86
+ $Y=1.82 $X2=6.86 $Y2=1.82
r77 16 26 6.83868 $w=2.1e-07 $l=1.44914e-07 $layer=LI1_cond $X=7.59 $Y=1.82
+ $X2=7.685 $Y2=1.925
r78 16 18 38.5541 $w=2.08e-07 $l=7.3e-07 $layer=LI1_cond $X=7.59 $Y=1.82
+ $X2=6.86 $Y2=1.82
r79 14 24 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.95 $Y=1.265
+ $X2=6.95 $Y2=1.1
r80 14 36 199.979 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=6.95 $Y=1.265
+ $X2=6.95 $Y2=1.655
r81 13 39 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=6.86 $Y=0.615
+ $X2=6.86 $Y2=0.935
r82 9 37 276.894 $w=1.5e-07 $l=5.4e-07 $layer=POLY_cond $X=6.77 $Y=2.525
+ $X2=6.77 $Y2=1.985
r83 2 28 600 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_PDIFF $count=1 $X=7.545
+ $Y=2.315 $X2=7.685 $Y2=2.45
r84 1 31 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=7.575
+ $Y=0.625 $X2=7.7 $Y2=0.9
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSTP_4%A_1211_463# 1 2 9 11 15 19 21 23 25 27 36
+ 37 40 43 45 47 49 53
c117 36 0 7.13856e-20 $X=6.195 $Y=2.47
c118 15 0 1.36539e-19 $X=7.915 $Y=0.835
c119 11 0 3.46573e-20 $X=7.84 $Y=1.355
c120 9 0 1.15292e-19 $X=7.47 $Y=2.525
r121 46 56 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.77 $Y=1.54
+ $X2=8.77 $Y2=1.705
r122 46 53 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=8.77 $Y=1.54 $X2=8.77
+ $Y2=1.45
r123 45 47 8.06855 $w=2.68e-07 $l=1.65e-07 $layer=LI1_cond $X=8.77 $Y=1.49
+ $X2=8.605 $Y2=1.49
r124 45 46 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.77
+ $Y=1.54 $X2=8.77 $Y2=1.54
r125 40 42 8.41541 $w=2.58e-07 $l=1.65e-07 $layer=LI1_cond $X=6.32 $Y=0.7
+ $X2=6.32 $Y2=0.865
r126 36 37 8.3262 $w=2.68e-07 $l=1.65e-07 $layer=LI1_cond $X=6.235 $Y=2.47
+ $X2=6.235 $Y2=2.305
r127 34 52 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.49 $Y=1.45
+ $X2=7.49 $Y2=1.615
r128 34 49 16.6118 $w=3.3e-07 $l=9.5e-08 $layer=POLY_cond $X=7.49 $Y=1.45
+ $X2=7.49 $Y2=1.355
r129 33 47 65.0861 $w=1.88e-07 $l=1.115e-06 $layer=LI1_cond $X=7.49 $Y=1.45
+ $X2=8.605 $Y2=1.45
r130 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.49
+ $Y=1.45 $X2=7.49 $Y2=1.45
r131 31 43 1.14861 $w=1.9e-07 $l=9e-08 $layer=LI1_cond $X=6.37 $Y=1.45 $X2=6.28
+ $Y2=1.45
r132 31 33 65.378 $w=1.88e-07 $l=1.12e-06 $layer=LI1_cond $X=6.37 $Y=1.45
+ $X2=7.49 $Y2=1.45
r133 28 43 5.40251 $w=1.8e-07 $l=9.5e-08 $layer=LI1_cond $X=6.28 $Y=1.545
+ $X2=6.28 $Y2=1.45
r134 28 37 46.8283 $w=1.78e-07 $l=7.6e-07 $layer=LI1_cond $X=6.28 $Y=1.545
+ $X2=6.28 $Y2=2.305
r135 27 43 5.40251 $w=1.8e-07 $l=9.5e-08 $layer=LI1_cond $X=6.28 $Y=1.355
+ $X2=6.28 $Y2=1.45
r136 27 42 30.1919 $w=1.78e-07 $l=4.9e-07 $layer=LI1_cond $X=6.28 $Y=1.355
+ $X2=6.28 $Y2=0.865
r137 23 25 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=9.365 $Y=1.375
+ $X2=9.365 $Y2=0.945
r138 22 53 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.935 $Y=1.45
+ $X2=8.77 $Y2=1.45
r139 21 23 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.29 $Y=1.45
+ $X2=9.365 $Y2=1.375
r140 21 22 182.032 $w=1.5e-07 $l=3.55e-07 $layer=POLY_cond $X=9.29 $Y=1.45
+ $X2=8.935 $Y2=1.45
r141 19 56 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=8.68 $Y=2.315
+ $X2=8.68 $Y2=1.705
r142 13 15 228.181 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=7.915 $Y=1.28
+ $X2=7.915 $Y2=0.835
r143 12 49 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.655 $Y=1.355
+ $X2=7.49 $Y2=1.355
r144 11 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.84 $Y=1.355
+ $X2=7.915 $Y2=1.28
r145 11 12 94.8617 $w=1.5e-07 $l=1.85e-07 $layer=POLY_cond $X=7.84 $Y=1.355
+ $X2=7.655 $Y2=1.355
r146 9 52 466.617 $w=1.5e-07 $l=9.1e-07 $layer=POLY_cond $X=7.47 $Y=2.525
+ $X2=7.47 $Y2=1.615
r147 2 36 600 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_PDIFF $count=1 $X=6.055
+ $Y=2.315 $X2=6.195 $Y2=2.47
r148 1 40 182 $w=1.7e-07 $l=3.58225e-07 $layer=licon1_NDIFF $count=1 $X=6.145
+ $Y=0.405 $X2=6.285 $Y2=0.7
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSTP_4%SET_B 3 5 6 7 10 13 17 20 21 23 24 26 27 28
+ 29 30 31
c97 26 0 1.36539e-19 $X=10.685 $Y=0.46
r98 39 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.48
+ $Y=0.35 $X2=8.48 $Y2=0.35
r99 30 31 13.492 $w=4.08e-07 $l=4.8e-07 $layer=LI1_cond $X=9.84 $Y=0.46
+ $X2=10.32 $Y2=0.46
r100 29 30 13.492 $w=4.08e-07 $l=4.8e-07 $layer=LI1_cond $X=9.36 $Y=0.46
+ $X2=9.84 $Y2=0.46
r101 28 29 13.492 $w=4.08e-07 $l=4.8e-07 $layer=LI1_cond $X=8.88 $Y=0.46
+ $X2=9.36 $Y2=0.46
r102 28 40 11.2433 $w=4.08e-07 $l=4e-07 $layer=LI1_cond $X=8.88 $Y=0.46 $X2=8.48
+ $Y2=0.46
r103 27 40 2.24867 $w=4.08e-07 $l=8e-08 $layer=LI1_cond $X=8.4 $Y=0.46 $X2=8.48
+ $Y2=0.46
r104 26 31 10.2596 $w=4.08e-07 $l=3.65e-07 $layer=LI1_cond $X=10.685 $Y=0.46
+ $X2=10.32 $Y2=0.46
r105 24 43 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=11.73 $Y=1.67
+ $X2=11.73 $Y2=1.835
r106 24 42 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=11.73 $Y=1.67
+ $X2=11.73 $Y2=1.505
r107 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.73
+ $Y=1.67 $X2=11.73 $Y2=1.67
r108 21 23 53.9141 $w=1.78e-07 $l=8.75e-07 $layer=LI1_cond $X=10.855 $Y=1.675
+ $X2=11.73 $Y2=1.675
r109 20 21 6.82373 $w=1.8e-07 $l=1.25499e-07 $layer=LI1_cond $X=10.77 $Y=1.585
+ $X2=10.855 $Y2=1.675
r110 19 26 8.45803 $w=4.1e-07 $l=2.43824e-07 $layer=LI1_cond $X=10.77 $Y=0.665
+ $X2=10.685 $Y2=0.46
r111 19 20 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=10.77 $Y=0.665
+ $X2=10.77 $Y2=1.585
r112 17 43 492.255 $w=1.5e-07 $l=9.6e-07 $layer=POLY_cond $X=11.66 $Y=2.795
+ $X2=11.66 $Y2=1.835
r113 13 42 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=11.64 $Y=0.835
+ $X2=11.64 $Y2=1.505
r114 8 10 428.16 $w=1.5e-07 $l=8.35e-07 $layer=POLY_cond $X=8.275 $Y=1.67
+ $X2=8.275 $Y2=0.835
r115 7 39 34.9152 $w=2.83e-07 $l=2.75409e-07 $layer=POLY_cond $X=8.275 $Y=0.515
+ $X2=8.48 $Y2=0.35
r116 7 10 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=8.275 $Y=0.515
+ $X2=8.275 $Y2=0.835
r117 5 8 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.2 $Y=1.745
+ $X2=8.275 $Y2=1.67
r118 5 6 94.8617 $w=1.5e-07 $l=1.85e-07 $layer=POLY_cond $X=8.2 $Y=1.745
+ $X2=8.015 $Y2=1.745
r119 1 6 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.94 $Y=1.82
+ $X2=8.015 $Y2=1.745
r120 1 3 361.5 $w=1.5e-07 $l=7.05e-07 $layer=POLY_cond $X=7.94 $Y=1.82 $X2=7.94
+ $Y2=2.525
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSTP_4%A_773_409# 1 2 9 13 17 18 19 22 23 24 25 27
+ 30 32 36 38 39 42 45 49 50 52 55 56 63 66
c164 36 0 9.96682e-20 $X=10.25 $Y=2.315
c165 30 0 3.02798e-20 $X=6.41 $Y=2.525
r166 67 68 30.474 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=4.82 $Y=2.2 $X2=4.82
+ $Y2=2.275
r167 60 63 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=3.95 $Y=0.495
+ $X2=4.105 $Y2=0.495
r168 56 67 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=4.82 $Y=2.11 $X2=4.82
+ $Y2=2.2
r169 56 66 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.82 $Y=2.11
+ $X2=4.82 $Y2=1.945
r170 55 56 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.82
+ $Y=2.11 $X2=4.82 $Y2=2.11
r171 53 59 2.79448 $w=3.4e-07 $l=1.05e-07 $layer=LI1_cond $X=4.035 $Y=2.115
+ $X2=3.93 $Y2=2.115
r172 53 55 26.6079 $w=3.38e-07 $l=7.85e-07 $layer=LI1_cond $X=4.035 $Y=2.115
+ $X2=4.82 $Y2=2.115
r173 52 59 5.05668 $w=1.7e-07 $l=1.79722e-07 $layer=LI1_cond $X=3.95 $Y=1.945
+ $X2=3.93 $Y2=2.115
r174 51 60 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.95 $Y=0.66
+ $X2=3.95 $Y2=0.495
r175 51 52 83.8342 $w=1.68e-07 $l=1.285e-06 $layer=LI1_cond $X=3.95 $Y=0.66
+ $X2=3.95 $Y2=1.945
r176 46 48 82.0426 $w=1.5e-07 $l=1.6e-07 $layer=POLY_cond $X=4.75 $Y=1.01
+ $X2=4.91 $Y2=1.01
r177 44 50 26.7401 $w=1.5e-07 $l=1.05e-07 $layer=POLY_cond $X=10.74 $Y=1.695
+ $X2=10.74 $Y2=1.59
r178 44 45 707.617 $w=1.5e-07 $l=1.38e-06 $layer=POLY_cond $X=10.74 $Y=1.695
+ $X2=10.74 $Y2=3.075
r179 40 50 26.7401 $w=1.5e-07 $l=1.05e-07 $layer=POLY_cond $X=10.74 $Y=1.485
+ $X2=10.74 $Y2=1.59
r180 40 42 333.298 $w=1.5e-07 $l=6.5e-07 $layer=POLY_cond $X=10.74 $Y=1.485
+ $X2=10.74 $Y2=0.835
r181 38 50 0.647981 $w=2.1e-07 $l=7.5e-08 $layer=POLY_cond $X=10.665 $Y=1.59
+ $X2=10.74 $Y2=1.59
r182 38 39 107.368 $w=2.1e-07 $l=3.4e-07 $layer=POLY_cond $X=10.665 $Y=1.59
+ $X2=10.325 $Y2=1.59
r183 34 39 27.9153 $w=2.1e-07 $l=1.37477e-07 $layer=POLY_cond $X=10.25 $Y=1.695
+ $X2=10.325 $Y2=1.59
r184 34 36 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=10.25 $Y=1.695
+ $X2=10.25 $Y2=2.315
r185 33 49 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.485 $Y=3.15
+ $X2=6.41 $Y2=3.15
r186 32 45 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=10.665 $Y=3.15
+ $X2=10.74 $Y2=3.075
r187 32 33 2143.36 $w=1.5e-07 $l=4.18e-06 $layer=POLY_cond $X=10.665 $Y=3.15
+ $X2=6.485 $Y2=3.15
r188 28 49 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.41 $Y=3.075
+ $X2=6.41 $Y2=3.15
r189 28 30 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=6.41 $Y=3.075
+ $X2=6.41 $Y2=2.525
r190 25 27 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=6.07 $Y=0.935
+ $X2=6.07 $Y2=0.615
r191 23 49 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.335 $Y=3.15
+ $X2=6.41 $Y2=3.15
r192 23 24 533.277 $w=1.5e-07 $l=1.04e-06 $layer=POLY_cond $X=6.335 $Y=3.15
+ $X2=5.295 $Y2=3.15
r193 22 24 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.22 $Y=3.075
+ $X2=5.295 $Y2=3.15
r194 21 22 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=5.22 $Y=2.275
+ $X2=5.22 $Y2=3.075
r195 20 67 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.985 $Y=2.2
+ $X2=4.82 $Y2=2.2
r196 19 21 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.145 $Y=2.2
+ $X2=5.22 $Y2=2.275
r197 19 20 82.0426 $w=1.5e-07 $l=1.6e-07 $layer=POLY_cond $X=5.145 $Y=2.2
+ $X2=4.985 $Y2=2.2
r198 18 48 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.985 $Y=1.01
+ $X2=4.91 $Y2=1.01
r199 17 25 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.995 $Y=1.01
+ $X2=6.07 $Y2=0.935
r200 17 18 517.894 $w=1.5e-07 $l=1.01e-06 $layer=POLY_cond $X=5.995 $Y=1.01
+ $X2=4.985 $Y2=1.01
r201 15 48 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.91 $Y=1.085
+ $X2=4.91 $Y2=1.01
r202 15 66 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=4.91 $Y=1.085
+ $X2=4.91 $Y2=1.945
r203 11 46 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.75 $Y=0.935
+ $X2=4.75 $Y2=1.01
r204 11 13 225.617 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=4.75 $Y=0.935
+ $X2=4.75 $Y2=0.495
r205 9 68 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=4.73 $Y=2.775 $X2=4.73
+ $Y2=2.275
r206 2 59 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=3.865
+ $Y=2.045 $X2=3.99 $Y2=2.19
r207 1 63 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=3.98
+ $Y=0.285 $X2=4.105 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSTP_4%A_2205_231# 1 2 9 12 14 17 19 21 25 30
c55 12 0 1.90511e-19 $X=11.23 $Y=2.795
r56 23 25 47.2697 $w=2.93e-07 $l=1.21e-06 $layer=LI1_cond $X=12.842 $Y=1.415
+ $X2=12.842 $Y2=2.625
r57 19 23 25.7157 $w=2.04e-07 $l=4.3e-07 $layer=LI1_cond $X=12.412 $Y=1.295
+ $X2=12.842 $Y2=1.295
r58 19 21 13.0871 $w=2.93e-07 $l=3.35e-07 $layer=LI1_cond $X=12.412 $Y=1.175
+ $X2=12.412 $Y2=0.84
r59 17 31 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=11.19 $Y=1.32
+ $X2=11.19 $Y2=1.485
r60 17 30 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=11.19 $Y=1.32
+ $X2=11.19 $Y2=1.155
r61 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.19
+ $Y=1.32 $X2=11.19 $Y2=1.32
r62 14 19 7.78198 $w=2.4e-07 $l=1.47e-07 $layer=LI1_cond $X=12.265 $Y=1.295
+ $X2=12.412 $Y2=1.295
r63 14 16 51.6198 $w=2.38e-07 $l=1.075e-06 $layer=LI1_cond $X=12.265 $Y=1.295
+ $X2=11.19 $Y2=1.295
r64 12 31 671.723 $w=1.5e-07 $l=1.31e-06 $layer=POLY_cond $X=11.23 $Y=2.795
+ $X2=11.23 $Y2=1.485
r65 9 30 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=11.165 $Y=0.835
+ $X2=11.165 $Y2=1.155
r66 2 25 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=12.685
+ $Y=2.415 $X2=12.825 $Y2=2.625
r67 1 21 182 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_NDIFF $count=1 $X=12.255
+ $Y=0.625 $X2=12.395 $Y2=0.84
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSTP_4%A_1960_125# 1 2 3 12 14 16 18 22 24 26 27
+ 28 30 32 34 36
c98 27 0 2.12354e-19 $X=13.545 $Y=1.65
r99 43 44 8.66906 $w=5.56e-07 $l=1e-07 $layer=POLY_cond $X=12.395 $Y=1.75
+ $X2=12.395 $Y2=1.65
r100 42 43 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=12.3
+ $Y=1.75 $X2=12.3 $Y2=1.75
r101 34 42 9.43173 $w=4.98e-07 $l=5.26498e-07 $layer=LI1_cond $X=11.915 $Y=2.255
+ $X2=12.3 $Y2=1.92
r102 34 36 21.4593 $w=2.88e-07 $l=5.4e-07 $layer=LI1_cond $X=11.915 $Y=2.255
+ $X2=11.915 $Y2=2.795
r103 33 39 7.62182 $w=1.9e-07 $l=3.23e-07 $layer=LI1_cond $X=10.515 $Y=2.03
+ $X2=10.192 $Y2=2.03
r104 32 34 8.4184 $w=4.98e-07 $l=2.88531e-07 $layer=LI1_cond $X=11.77 $Y=2.03
+ $X2=11.915 $Y2=2.255
r105 32 33 73.2584 $w=1.88e-07 $l=1.255e-06 $layer=LI1_cond $X=11.77 $Y=2.03
+ $X2=10.515 $Y2=2.03
r106 28 39 2.24171 $w=6.45e-07 $l=9.5e-08 $layer=LI1_cond $X=10.192 $Y=1.935
+ $X2=10.192 $Y2=2.03
r107 28 30 17.3385 $w=6.43e-07 $l=9.35e-07 $layer=LI1_cond $X=10.192 $Y=1.935
+ $X2=10.192 $Y2=1
r108 24 27 20.4101 $w=1.5e-07 $l=8.21584e-08 $layer=POLY_cond $X=13.56 $Y=1.725
+ $X2=13.545 $Y2=1.65
r109 24 26 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=13.56 $Y=1.725
+ $X2=13.56 $Y2=2.465
r110 20 27 20.4101 $w=1.5e-07 $l=8.21584e-08 $layer=POLY_cond $X=13.53 $Y=1.575
+ $X2=13.545 $Y2=1.65
r111 20 22 456.362 $w=1.5e-07 $l=8.9e-07 $layer=POLY_cond $X=13.53 $Y=1.575
+ $X2=13.53 $Y2=0.685
r112 19 44 34.1107 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=12.685 $Y=1.65
+ $X2=12.395 $Y2=1.65
r113 18 27 5.30422 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=13.455 $Y=1.65
+ $X2=13.545 $Y2=1.65
r114 18 19 394.83 $w=1.5e-07 $l=7.7e-07 $layer=POLY_cond $X=13.455 $Y=1.65
+ $X2=12.685 $Y2=1.65
r115 14 43 72.8768 $w=5.56e-07 $l=6.02993e-07 $layer=POLY_cond $X=12.61 $Y=2.255
+ $X2=12.395 $Y2=1.75
r116 14 16 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=12.61 $Y=2.255
+ $X2=12.61 $Y2=2.625
r117 10 44 35.5998 $w=5.56e-07 $l=2.497e-07 $layer=POLY_cond $X=12.18 $Y=1.575
+ $X2=12.395 $Y2=1.65
r118 10 12 379.447 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=12.18 $Y=1.575
+ $X2=12.18 $Y2=0.835
r119 3 36 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=11.735
+ $Y=2.585 $X2=11.875 $Y2=2.795
r120 2 39 600 $w=1.7e-07 $l=3.745e-07 $layer=licon1_PDIFF $count=1 $X=9.8
+ $Y=2.315 $X2=10.035 $Y2=2.04
r121 1 30 91 $w=1.7e-07 $l=7.95707e-07 $layer=licon1_NDIFF $count=2 $X=9.8
+ $Y=0.625 $X2=10.43 $Y2=1
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSTP_4%A_2638_53# 1 2 9 13 17 21 25 29 33 37 41 45
+ 54 57 68
c105 57 0 4.70822e-20 $X=13.32 $Y=1.51
r106 67 68 5.24584 $w=3.3e-07 $l=3e-08 $layer=POLY_cond $X=15.25 $Y=1.51
+ $X2=15.28 $Y2=1.51
r107 66 67 69.9445 $w=3.3e-07 $l=4e-07 $layer=POLY_cond $X=14.85 $Y=1.51
+ $X2=15.25 $Y2=1.51
r108 65 66 5.24584 $w=3.3e-07 $l=3e-08 $layer=POLY_cond $X=14.82 $Y=1.51
+ $X2=14.85 $Y2=1.51
r109 62 63 5.24584 $w=3.3e-07 $l=3e-08 $layer=POLY_cond $X=14.39 $Y=1.51
+ $X2=14.42 $Y2=1.51
r110 58 60 5.24584 $w=3.3e-07 $l=3e-08 $layer=POLY_cond $X=13.96 $Y=1.51
+ $X2=13.99 $Y2=1.51
r111 55 65 22.732 $w=3.3e-07 $l=1.3e-07 $layer=POLY_cond $X=14.69 $Y=1.51
+ $X2=14.82 $Y2=1.51
r112 55 63 47.2125 $w=3.3e-07 $l=2.7e-07 $layer=POLY_cond $X=14.69 $Y=1.51
+ $X2=14.42 $Y2=1.51
r113 54 55 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=14.69
+ $Y=1.51 $X2=14.69 $Y2=1.51
r114 52 62 66.4473 $w=3.3e-07 $l=3.8e-07 $layer=POLY_cond $X=14.01 $Y=1.51
+ $X2=14.39 $Y2=1.51
r115 52 60 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=14.01 $Y=1.51
+ $X2=13.99 $Y2=1.51
r116 51 54 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=14.01 $Y=1.51
+ $X2=14.69 $Y2=1.51
r117 51 52 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=14.01
+ $Y=1.51 $X2=14.01 $Y2=1.51
r118 49 57 3.25423 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=13.48 $Y=1.51
+ $X2=13.32 $Y2=1.51
r119 49 51 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=13.48 $Y=1.51
+ $X2=14.01 $Y2=1.51
r120 45 47 33.4929 $w=3.18e-07 $l=9.3e-07 $layer=LI1_cond $X=13.32 $Y=1.98
+ $X2=13.32 $Y2=2.91
r121 43 57 3.29812 $w=2.85e-07 $l=8.5e-08 $layer=LI1_cond $X=13.32 $Y=1.595
+ $X2=13.32 $Y2=1.51
r122 43 45 13.8653 $w=3.18e-07 $l=3.85e-07 $layer=LI1_cond $X=13.32 $Y=1.595
+ $X2=13.32 $Y2=1.98
r123 39 57 3.29812 $w=2.85e-07 $l=1.00995e-07 $layer=LI1_cond $X=13.285 $Y=1.425
+ $X2=13.32 $Y2=1.51
r124 39 41 46.3282 $w=2.48e-07 $l=1.005e-06 $layer=LI1_cond $X=13.285 $Y=1.425
+ $X2=13.285 $Y2=0.42
r125 35 68 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=15.28 $Y=1.675
+ $X2=15.28 $Y2=1.51
r126 35 37 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=15.28 $Y=1.675
+ $X2=15.28 $Y2=2.465
r127 31 67 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=15.25 $Y=1.345
+ $X2=15.25 $Y2=1.51
r128 31 33 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=15.25 $Y=1.345
+ $X2=15.25 $Y2=0.685
r129 27 66 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=14.85 $Y=1.675
+ $X2=14.85 $Y2=1.51
r130 27 29 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=14.85 $Y=1.675
+ $X2=14.85 $Y2=2.465
r131 23 65 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=14.82 $Y=1.345
+ $X2=14.82 $Y2=1.51
r132 23 25 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=14.82 $Y=1.345
+ $X2=14.82 $Y2=0.685
r133 19 63 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=14.42 $Y=1.675
+ $X2=14.42 $Y2=1.51
r134 19 21 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=14.42 $Y=1.675
+ $X2=14.42 $Y2=2.465
r135 15 62 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=14.39 $Y=1.345
+ $X2=14.39 $Y2=1.51
r136 15 17 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=14.39 $Y=1.345
+ $X2=14.39 $Y2=0.685
r137 11 60 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=13.99 $Y=1.675
+ $X2=13.99 $Y2=1.51
r138 11 13 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=13.99 $Y=1.675
+ $X2=13.99 $Y2=2.465
r139 7 58 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=13.96 $Y=1.345
+ $X2=13.96 $Y2=1.51
r140 7 9 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=13.96 $Y=1.345
+ $X2=13.96 $Y2=0.685
r141 2 47 400 $w=1.7e-07 $l=1.13578e-06 $layer=licon1_PDIFF $count=1 $X=13.22
+ $Y=1.835 $X2=13.345 $Y2=2.91
r142 2 45 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=13.22
+ $Y=1.835 $X2=13.345 $Y2=1.98
r143 1 41 91 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=2 $X=13.19
+ $Y=0.265 $X2=13.315 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSTP_4%A_27_479# 1 2 9 11 12
r27 11 16 6.95815 $w=2.63e-07 $l=1.6e-07 $layer=LI1_cond $X=2.002 $Y=2.41
+ $X2=2.002 $Y2=2.57
r28 11 12 98.8396 $w=1.68e-07 $l=1.515e-06 $layer=LI1_cond $X=1.87 $Y=2.41
+ $X2=0.355 $Y2=2.41
r29 7 12 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=0.225 $Y=2.495
+ $X2=0.355 $Y2=2.41
r30 7 9 1.99461 $w=2.58e-07 $l=4.5e-08 $layer=LI1_cond $X=0.225 $Y=2.495
+ $X2=0.225 $Y2=2.54
r31 2 16 600 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_PDIFF $count=1 $X=1.88
+ $Y=2.395 $X2=2.02 $Y2=2.57
r32 1 9 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.395 $X2=0.26 $Y2=2.54
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSTP_4%VPWR 1 2 3 4 5 6 7 8 9 10 33 37 41 43 47 51
+ 55 57 61 65 71 75 77 82 83 84 85 86 88 100 107 119 124 129 135 138 141 144 147
+ 150 153 157
r184 156 157 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=15.6 $Y=3.33
+ $X2=15.6 $Y2=3.33
r185 153 154 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.64 $Y=3.33
+ $X2=14.64 $Y2=3.33
r186 150 151 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=13.68 $Y=3.33
+ $X2=13.68 $Y2=3.33
r187 147 148 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=12.24 $Y=3.33
+ $X2=12.24 $Y2=3.33
r188 144 145 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r189 141 142 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r190 139 142 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=6.96 $Y2=3.33
r191 138 139 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r192 135 136 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r193 133 157 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=15.12 $Y=3.33
+ $X2=15.6 $Y2=3.33
r194 133 154 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=15.12 $Y=3.33
+ $X2=14.64 $Y2=3.33
r195 132 133 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=15.12 $Y=3.33
+ $X2=15.12 $Y2=3.33
r196 130 153 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=14.8 $Y=3.33
+ $X2=14.635 $Y2=3.33
r197 130 132 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=14.8 $Y=3.33
+ $X2=15.12 $Y2=3.33
r198 129 156 4.60552 $w=1.7e-07 $l=2.55e-07 $layer=LI1_cond $X=15.33 $Y=3.33
+ $X2=15.585 $Y2=3.33
r199 129 132 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=15.33 $Y=3.33
+ $X2=15.12 $Y2=3.33
r200 128 154 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=14.16 $Y=3.33
+ $X2=14.64 $Y2=3.33
r201 128 151 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=14.16 $Y=3.33
+ $X2=13.68 $Y2=3.33
r202 127 128 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.16 $Y=3.33
+ $X2=14.16 $Y2=3.33
r203 125 150 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=13.9 $Y=3.33
+ $X2=13.775 $Y2=3.33
r204 125 127 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=13.9 $Y=3.33
+ $X2=14.16 $Y2=3.33
r205 124 153 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=14.47 $Y=3.33
+ $X2=14.635 $Y2=3.33
r206 124 127 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=14.47 $Y=3.33
+ $X2=14.16 $Y2=3.33
r207 123 151 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=12.72 $Y=3.33
+ $X2=13.68 $Y2=3.33
r208 123 148 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.72 $Y=3.33
+ $X2=12.24 $Y2=3.33
r209 122 123 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=12.72 $Y=3.33
+ $X2=12.72 $Y2=3.33
r210 120 147 7.94884 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=12.525 $Y=3.33
+ $X2=12.377 $Y2=3.33
r211 120 122 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=12.525 $Y=3.33
+ $X2=12.72 $Y2=3.33
r212 119 150 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=13.65 $Y=3.33
+ $X2=13.775 $Y2=3.33
r213 119 122 60.6738 $w=1.68e-07 $l=9.3e-07 $layer=LI1_cond $X=13.65 $Y=3.33
+ $X2=12.72 $Y2=3.33
r214 118 148 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=11.28 $Y=3.33
+ $X2=12.24 $Y2=3.33
r215 117 118 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=11.28 $Y=3.33
+ $X2=11.28 $Y2=3.33
r216 115 118 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=11.28 $Y2=3.33
r217 115 145 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=8.4 $Y2=3.33
r218 114 117 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=8.88 $Y=3.33
+ $X2=11.28 $Y2=3.33
r219 114 115 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r220 112 144 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.63 $Y=3.33
+ $X2=8.465 $Y2=3.33
r221 112 114 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=8.63 $Y=3.33
+ $X2=8.88 $Y2=3.33
r222 108 141 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=7.08 $Y=3.33
+ $X2=6.985 $Y2=3.33
r223 108 110 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=7.08 $Y=3.33
+ $X2=7.92 $Y2=3.33
r224 107 144 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.3 $Y=3.33
+ $X2=8.465 $Y2=3.33
r225 107 110 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=8.3 $Y=3.33
+ $X2=7.92 $Y2=3.33
r226 106 139 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r227 105 106 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r228 103 106 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=4.08 $Y2=3.33
r229 102 105 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=3.12 $Y=3.33
+ $X2=4.08 $Y2=3.33
r230 102 103 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r231 100 138 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=4.35 $Y=3.33
+ $X2=4.48 $Y2=3.33
r232 100 105 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=4.35 $Y=3.33
+ $X2=4.08 $Y2=3.33
r233 99 103 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r234 98 99 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r235 96 99 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r236 96 136 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r237 95 98 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r238 95 96 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r239 93 135 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.855 $Y=3.33
+ $X2=0.69 $Y2=3.33
r240 93 95 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.855 $Y=3.33
+ $X2=1.2 $Y2=3.33
r241 91 136 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r242 90 91 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r243 88 135 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.525 $Y=3.33
+ $X2=0.69 $Y2=3.33
r244 88 90 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.525 $Y=3.33
+ $X2=0.24 $Y2=3.33
r245 86 145 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=8.4 $Y2=3.33
r246 86 142 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=6.96 $Y2=3.33
r247 86 110 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r248 84 117 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=11.34 $Y=3.33
+ $X2=11.28 $Y2=3.33
r249 84 85 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=11.34 $Y=3.33
+ $X2=11.445 $Y2=3.33
r250 82 98 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=2.645 $Y=3.33
+ $X2=2.64 $Y2=3.33
r251 82 83 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=2.645 $Y=3.33
+ $X2=2.75 $Y2=3.33
r252 81 102 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=2.855 $Y=3.33
+ $X2=3.12 $Y2=3.33
r253 81 83 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=2.855 $Y=3.33
+ $X2=2.75 $Y2=3.33
r254 77 80 26.5411 $w=3.28e-07 $l=7.6e-07 $layer=LI1_cond $X=15.495 $Y=2.19
+ $X2=15.495 $Y2=2.95
r255 75 156 3.16065 $w=3.3e-07 $l=1.25499e-07 $layer=LI1_cond $X=15.495 $Y=3.245
+ $X2=15.585 $Y2=3.33
r256 75 80 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=15.495 $Y=3.245
+ $X2=15.495 $Y2=2.95
r257 71 74 27.2396 $w=3.28e-07 $l=7.8e-07 $layer=LI1_cond $X=14.635 $Y=2.19
+ $X2=14.635 $Y2=2.97
r258 69 153 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=14.635 $Y=3.245
+ $X2=14.635 $Y2=3.33
r259 69 74 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=14.635 $Y=3.245
+ $X2=14.635 $Y2=2.97
r260 65 68 45.6367 $w=2.48e-07 $l=9.9e-07 $layer=LI1_cond $X=13.775 $Y=1.98
+ $X2=13.775 $Y2=2.97
r261 63 150 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=13.775 $Y=3.245
+ $X2=13.775 $Y2=3.33
r262 63 68 12.6769 $w=2.48e-07 $l=2.75e-07 $layer=LI1_cond $X=13.775 $Y=3.245
+ $X2=13.775 $Y2=2.97
r263 59 147 0.543863 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=12.377 $Y=3.245
+ $X2=12.377 $Y2=3.33
r264 59 61 24.2208 $w=2.93e-07 $l=6.2e-07 $layer=LI1_cond $X=12.377 $Y=3.245
+ $X2=12.377 $Y2=2.625
r265 58 85 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=11.55 $Y=3.33
+ $X2=11.445 $Y2=3.33
r266 57 147 7.94884 $w=1.7e-07 $l=1.47e-07 $layer=LI1_cond $X=12.23 $Y=3.33
+ $X2=12.377 $Y2=3.33
r267 57 58 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=12.23 $Y=3.33
+ $X2=11.55 $Y2=3.33
r268 53 85 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=11.445 $Y=3.245
+ $X2=11.445 $Y2=3.33
r269 53 55 23.7662 $w=2.08e-07 $l=4.5e-07 $layer=LI1_cond $X=11.445 $Y=3.245
+ $X2=11.445 $Y2=2.795
r270 49 144 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.465 $Y=3.245
+ $X2=8.465 $Y2=3.33
r271 49 51 35.7956 $w=3.28e-07 $l=1.025e-06 $layer=LI1_cond $X=8.465 $Y=3.245
+ $X2=8.465 $Y2=2.22
r272 45 141 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=6.985 $Y=3.245
+ $X2=6.985 $Y2=3.33
r273 45 47 37.6507 $w=1.88e-07 $l=6.45e-07 $layer=LI1_cond $X=6.985 $Y=3.245
+ $X2=6.985 $Y2=2.6
r274 44 138 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=4.61 $Y=3.33
+ $X2=4.48 $Y2=3.33
r275 43 141 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=6.89 $Y=3.33
+ $X2=6.985 $Y2=3.33
r276 43 44 148.749 $w=1.68e-07 $l=2.28e-06 $layer=LI1_cond $X=6.89 $Y=3.33
+ $X2=4.61 $Y2=3.33
r277 39 138 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=4.48 $Y=3.245
+ $X2=4.48 $Y2=3.33
r278 39 41 12.6325 $w=2.58e-07 $l=2.85e-07 $layer=LI1_cond $X=4.48 $Y=3.245
+ $X2=4.48 $Y2=2.96
r279 35 83 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=2.75 $Y=3.245
+ $X2=2.75 $Y2=3.33
r280 35 37 18.7489 $w=2.08e-07 $l=3.55e-07 $layer=LI1_cond $X=2.75 $Y=3.245
+ $X2=2.75 $Y2=2.89
r281 31 135 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=3.245
+ $X2=0.69 $Y2=3.33
r282 31 33 15.8897 $w=3.28e-07 $l=4.55e-07 $layer=LI1_cond $X=0.69 $Y=3.245
+ $X2=0.69 $Y2=2.79
r283 10 80 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=15.355
+ $Y=1.835 $X2=15.495 $Y2=2.95
r284 10 77 400 $w=1.7e-07 $l=4.19196e-07 $layer=licon1_PDIFF $count=1 $X=15.355
+ $Y=1.835 $X2=15.495 $Y2=2.19
r285 9 74 400 $w=1.7e-07 $l=1.20297e-06 $layer=licon1_PDIFF $count=1 $X=14.495
+ $Y=1.835 $X2=14.635 $Y2=2.97
r286 9 71 400 $w=1.7e-07 $l=4.19196e-07 $layer=licon1_PDIFF $count=1 $X=14.495
+ $Y=1.835 $X2=14.635 $Y2=2.19
r287 8 68 400 $w=1.7e-07 $l=1.20297e-06 $layer=licon1_PDIFF $count=1 $X=13.635
+ $Y=1.835 $X2=13.775 $Y2=2.97
r288 8 65 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=13.635
+ $Y=1.835 $X2=13.775 $Y2=1.98
r289 7 61 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=12.27
+ $Y=2.415 $X2=12.395 $Y2=2.625
r290 6 55 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=11.305
+ $Y=2.585 $X2=11.445 $Y2=2.795
r291 5 51 300 $w=1.7e-07 $l=4.95227e-07 $layer=licon1_PDIFF $count=2 $X=8.015
+ $Y=2.315 $X2=8.465 $Y2=2.22
r292 4 47 600 $w=1.7e-07 $l=3.4803e-07 $layer=licon1_PDIFF $count=1 $X=6.845
+ $Y=2.315 $X2=6.985 $Y2=2.6
r293 3 41 600 $w=1.7e-07 $l=5.70723e-07 $layer=licon1_PDIFF $count=1 $X=4.375
+ $Y=2.455 $X2=4.515 $Y2=2.96
r294 2 37 600 $w=1.7e-07 $l=5.43921e-07 $layer=licon1_PDIFF $count=1 $X=2.635
+ $Y=2.405 $X2=2.76 $Y2=2.89
r295 1 33 600 $w=1.7e-07 $l=4.59701e-07 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=2.395 $X2=0.69 $Y2=2.79
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSTP_4%A_218_119# 1 2 3 4 15 17 18 19 22 24 25 26
+ 28 29 30 32 33 34 36 38 46
c143 17 0 1.1672e-19 $X=2.425 $Y=1.377
r144 46 48 4.38905 $w=3.38e-07 $l=1.05e-07 $layer=LI1_cond $X=5.51 $Y=0.7
+ $X2=5.51 $Y2=0.805
r145 42 44 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=2.39 $Y=2.47
+ $X2=2.51 $Y2=2.47
r146 38 40 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=1.535 $Y=2.79
+ $X2=1.535 $Y2=2.99
r147 36 50 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.465 $Y=2.455
+ $X2=5.465 $Y2=2.54
r148 36 48 76.0612 $w=2.48e-07 $l=1.65e-06 $layer=LI1_cond $X=5.465 $Y=2.455
+ $X2=5.465 $Y2=0.805
r149 33 50 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.34 $Y=2.54
+ $X2=5.465 $Y2=2.54
r150 33 34 75.6791 $w=1.68e-07 $l=1.16e-06 $layer=LI1_cond $X=5.34 $Y=2.54
+ $X2=4.18 $Y2=2.54
r151 31 34 6.9898 $w=1.7e-07 $l=1.49579e-07 $layer=LI1_cond $X=4.067 $Y=2.625
+ $X2=4.18 $Y2=2.54
r152 31 32 14.3415 $w=2.23e-07 $l=2.8e-07 $layer=LI1_cond $X=4.067 $Y=2.625
+ $X2=4.067 $Y2=2.905
r153 29 32 6.9898 $w=1.7e-07 $l=1.4854e-07 $layer=LI1_cond $X=3.955 $Y=2.99
+ $X2=4.067 $Y2=2.905
r154 29 30 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=3.955 $Y=2.99
+ $X2=3.195 $Y2=2.99
r155 28 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.11 $Y=2.905
+ $X2=3.195 $Y2=2.99
r156 27 28 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=3.11 $Y=2.555
+ $X2=3.11 $Y2=2.905
r157 26 44 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=2.595 $Y=2.47
+ $X2=2.51 $Y2=2.47
r158 25 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.025 $Y=2.47
+ $X2=3.11 $Y2=2.555
r159 25 26 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=3.025 $Y=2.47
+ $X2=2.595 $Y2=2.47
r160 24 44 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.51 $Y=2.385
+ $X2=2.51 $Y2=2.47
r161 23 24 55.1283 $w=1.68e-07 $l=8.45e-07 $layer=LI1_cond $X=2.51 $Y=1.54
+ $X2=2.51 $Y2=2.385
r162 21 42 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.39 $Y=2.555
+ $X2=2.39 $Y2=2.47
r163 21 22 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=2.39 $Y=2.555
+ $X2=2.39 $Y2=2.905
r164 20 40 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.7 $Y=2.99
+ $X2=1.535 $Y2=2.99
r165 19 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.305 $Y=2.99
+ $X2=2.39 $Y2=2.905
r166 19 20 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=2.305 $Y=2.99
+ $X2=1.7 $Y2=2.99
r167 17 23 7.72402 $w=3.25e-07 $l=2.01057e-07 $layer=LI1_cond $X=2.425 $Y=1.377
+ $X2=2.51 $Y2=1.54
r168 17 18 36.5236 $w=3.23e-07 $l=1.03e-06 $layer=LI1_cond $X=2.425 $Y=1.377
+ $X2=1.395 $Y2=1.377
r169 13 18 6.81701 $w=3.25e-07 $l=2.32282e-07 $layer=LI1_cond $X=1.23 $Y=1.215
+ $X2=1.395 $Y2=1.377
r170 13 15 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=1.23 $Y=1.215
+ $X2=1.23 $Y2=0.805
r171 4 50 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=5.37
+ $Y=2.315 $X2=5.495 $Y2=2.46
r172 3 38 600 $w=1.7e-07 $l=4.82753e-07 $layer=licon1_PDIFF $count=1 $X=1.34
+ $Y=2.395 $X2=1.535 $Y2=2.79
r173 2 46 182 $w=1.7e-07 $l=3.64349e-07 $layer=licon1_NDIFF $count=1 $X=5.36
+ $Y=0.405 $X2=5.515 $Y2=0.7
r174 1 15 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.09
+ $Y=0.595 $X2=1.23 $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSTP_4%A_1751_379# 1 2 9 15 16
r30 15 16 8.84356 $w=2.28e-07 $l=1.65e-07 $layer=LI1_cond $X=10.465 $Y=2.41
+ $X2=10.3 $Y2=2.41
r31 9 12 4.15909 $w=1.98e-07 $l=7.5e-08 $layer=LI1_cond $X=8.9 $Y=2.385 $X2=8.9
+ $Y2=2.46
r32 8 9 1.35108 $w=1.8e-07 $l=1e-07 $layer=LI1_cond $X=9 $Y=2.385 $X2=8.9
+ $Y2=2.385
r33 8 16 80.101 $w=1.78e-07 $l=1.3e-06 $layer=LI1_cond $X=9 $Y=2.385 $X2=10.3
+ $Y2=2.385
r34 2 15 600 $w=1.7e-07 $l=5.80797e-07 $layer=licon1_PDIFF $count=1 $X=10.325
+ $Y=1.895 $X2=10.465 $Y2=2.41
r35 1 12 600 $w=1.7e-07 $l=6.3113e-07 $layer=licon1_PDIFF $count=1 $X=8.755
+ $Y=1.895 $X2=8.895 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSTP_4%A_1858_463# 1 2 9 14
c19 9 0 1.90511e-19 $X=11.015 $Y=2.86
r20 12 14 5.23454 $w=3.78e-07 $l=1.65e-07 $layer=LI1_cond $X=9.415 $Y=2.835
+ $X2=9.58 $Y2=2.835
r21 9 14 50.1138 $w=3.28e-07 $l=1.435e-06 $layer=LI1_cond $X=11.015 $Y=2.86
+ $X2=9.58 $Y2=2.86
r22 2 9 600 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_PDIFF $count=1 $X=10.89
+ $Y=2.585 $X2=11.015 $Y2=2.86
r23 1 12 600 $w=1.7e-07 $l=4.83477e-07 $layer=licon1_PDIFF $count=1 $X=9.29
+ $Y=2.315 $X2=9.415 $Y2=2.74
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSTP_4%Q 1 2 3 4 15 21 23 24 25 26 29 33 38 39 47
r64 45 47 0.736048 $w=6.48e-07 $l=4e-08 $layer=LI1_cond $X=15.36 $Y=1.255
+ $X2=15.36 $Y2=1.295
r65 39 45 2.43731 $w=4.2e-07 $l=1.11445e-07 $layer=LI1_cond $X=15.312 $Y=1.165
+ $X2=15.36 $Y2=1.255
r66 39 47 0.404827 $w=6.48e-07 $l=2.2e-08 $layer=LI1_cond $X=15.36 $Y=1.317
+ $X2=15.36 $Y2=1.295
r67 37 39 8.24374 $w=6.48e-07 $l=4.48e-07 $layer=LI1_cond $X=15.36 $Y=1.765
+ $X2=15.36 $Y2=1.317
r68 37 38 2.31106 $w=4.2e-07 $l=1.0015e-07 $layer=LI1_cond $X=15.36 $Y=1.765
+ $X2=15.327 $Y2=1.85
r69 33 35 55.4545 $w=1.88e-07 $l=9.5e-07 $layer=LI1_cond $X=15.065 $Y=1.96
+ $X2=15.065 $Y2=2.91
r70 31 38 2.31106 $w=4.2e-07 $l=3.01519e-07 $layer=LI1_cond $X=15.065 $Y=1.935
+ $X2=15.327 $Y2=1.85
r71 31 33 1.45933 $w=1.88e-07 $l=2.5e-08 $layer=LI1_cond $X=15.065 $Y=1.935
+ $X2=15.065 $Y2=1.96
r72 27 39 2.43731 $w=4.2e-07 $l=3.1884e-07 $layer=LI1_cond $X=15.035 $Y=1.075
+ $X2=15.312 $Y2=1.165
r73 27 29 38.2345 $w=1.88e-07 $l=6.55e-07 $layer=LI1_cond $X=15.035 $Y=1.075
+ $X2=15.035 $Y2=0.42
r74 25 38 4.73016 $w=1.7e-07 $l=3.57e-07 $layer=LI1_cond $X=14.97 $Y=1.85
+ $X2=15.327 $Y2=1.85
r75 25 26 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=14.97 $Y=1.85
+ $X2=14.3 $Y2=1.85
r76 23 39 4.51133 $w=1.8e-07 $l=3.72e-07 $layer=LI1_cond $X=14.94 $Y=1.165
+ $X2=15.312 $Y2=1.165
r77 23 24 41.2828 $w=1.78e-07 $l=6.7e-07 $layer=LI1_cond $X=14.94 $Y=1.165
+ $X2=14.27 $Y2=1.165
r78 19 24 6.82297 $w=1.8e-07 $l=1.32571e-07 $layer=LI1_cond $X=14.175 $Y=1.075
+ $X2=14.27 $Y2=1.165
r79 19 21 38.2345 $w=1.88e-07 $l=6.55e-07 $layer=LI1_cond $X=14.175 $Y=1.075
+ $X2=14.175 $Y2=0.42
r80 15 17 47.6009 $w=2.28e-07 $l=9.5e-07 $layer=LI1_cond $X=14.185 $Y=1.96
+ $X2=14.185 $Y2=2.91
r81 13 26 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=14.185 $Y=1.935
+ $X2=14.3 $Y2=1.85
r82 13 15 1.25266 $w=2.28e-07 $l=2.5e-08 $layer=LI1_cond $X=14.185 $Y=1.935
+ $X2=14.185 $Y2=1.96
r83 4 35 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=14.925
+ $Y=1.835 $X2=15.065 $Y2=2.91
r84 4 33 400 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=14.925
+ $Y=1.835 $X2=15.065 $Y2=1.96
r85 3 17 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=14.065
+ $Y=1.835 $X2=14.205 $Y2=2.91
r86 3 15 400 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=14.065
+ $Y=1.835 $X2=14.205 $Y2=1.96
r87 2 29 91 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=2 $X=14.895
+ $Y=0.265 $X2=15.035 $Y2=0.42
r88 1 21 91 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=2 $X=14.035
+ $Y=0.265 $X2=14.175 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSTP_4%VGND 1 2 3 4 5 6 7 8 9 30 34 38 42 45 46 50
+ 54 58 62 64 66 69 70 72 73 74 79 86 91 100 104 112 117 123 126 129 132 135 138
+ 142
c169 58 0 1.65272e-19 $X=13.745 $Y=0.39
c170 50 0 1.52906e-19 $X=9.15 $Y=1.015
r171 141 142 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=15.6 $Y=0
+ $X2=15.6 $Y2=0
r172 138 139 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.64 $Y=0
+ $X2=14.64 $Y2=0
r173 135 136 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.68 $Y=0
+ $X2=13.68 $Y2=0
r174 132 133 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=11.76 $Y=0
+ $X2=11.76 $Y2=0
r175 129 130 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.96 $Y=0
+ $X2=6.96 $Y2=0
r176 126 127 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=0
+ $X2=4.56 $Y2=0
r177 123 124 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.16 $Y=0
+ $X2=2.16 $Y2=0
r178 121 142 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=15.12 $Y=0
+ $X2=15.6 $Y2=0
r179 121 139 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=15.12 $Y=0
+ $X2=14.64 $Y2=0
r180 120 121 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=15.12 $Y=0
+ $X2=15.12 $Y2=0
r181 118 138 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=14.77 $Y=0
+ $X2=14.605 $Y2=0
r182 118 120 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=14.77 $Y=0
+ $X2=15.12 $Y2=0
r183 117 141 4.55841 $w=1.7e-07 $l=2.7e-07 $layer=LI1_cond $X=15.3 $Y=0
+ $X2=15.57 $Y2=0
r184 117 120 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=15.3 $Y=0
+ $X2=15.12 $Y2=0
r185 116 139 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=14.16 $Y=0
+ $X2=14.64 $Y2=0
r186 116 136 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=14.16 $Y=0
+ $X2=13.68 $Y2=0
r187 115 116 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.16 $Y=0
+ $X2=14.16 $Y2=0
r188 113 135 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.91 $Y=0
+ $X2=13.745 $Y2=0
r189 113 115 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=13.91 $Y=0
+ $X2=14.16 $Y2=0
r190 112 138 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=14.44 $Y=0
+ $X2=14.605 $Y2=0
r191 112 115 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=14.44 $Y=0
+ $X2=14.16 $Y2=0
r192 111 136 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.2 $Y=0
+ $X2=13.68 $Y2=0
r193 110 111 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=13.2 $Y=0
+ $X2=13.2 $Y2=0
r194 108 111 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=12.24 $Y=0
+ $X2=13.2 $Y2=0
r195 108 133 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.24 $Y=0
+ $X2=11.76 $Y2=0
r196 107 110 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=12.24 $Y=0
+ $X2=13.2 $Y2=0
r197 107 108 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=12.24 $Y=0
+ $X2=12.24 $Y2=0
r198 105 132 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.075 $Y=0
+ $X2=11.91 $Y2=0
r199 105 107 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=12.075 $Y=0
+ $X2=12.24 $Y2=0
r200 104 135 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.58 $Y=0
+ $X2=13.745 $Y2=0
r201 104 110 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=13.58 $Y=0
+ $X2=13.2 $Y2=0
r202 103 133 0.936549 $w=4.9e-07 $l=3.36e-06 $layer=MET1_cond $X=8.4 $Y=0
+ $X2=11.76 $Y2=0
r203 102 103 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=8.4 $Y=0
+ $X2=8.4 $Y2=0
r204 100 132 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.745 $Y=0
+ $X2=11.91 $Y2=0
r205 100 102 218.23 $w=1.68e-07 $l=3.345e-06 $layer=LI1_cond $X=11.745 $Y=0
+ $X2=8.4 $Y2=0
r206 96 129 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.24 $Y=0
+ $X2=7.075 $Y2=0
r207 96 98 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=7.24 $Y=0 $X2=7.92
+ $Y2=0
r208 95 130 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=5.04 $Y=0
+ $X2=6.96 $Y2=0
r209 95 127 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0
+ $X2=4.56 $Y2=0
r210 94 95 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.04 $Y=0
+ $X2=5.04 $Y2=0
r211 92 126 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.66 $Y=0
+ $X2=4.535 $Y2=0
r212 92 94 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=4.66 $Y=0 $X2=5.04
+ $Y2=0
r213 91 129 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.91 $Y=0
+ $X2=7.075 $Y2=0
r214 91 94 122 $w=1.68e-07 $l=1.87e-06 $layer=LI1_cond $X=6.91 $Y=0 $X2=5.04
+ $Y2=0
r215 90 127 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0
+ $X2=4.56 $Y2=0
r216 90 124 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=4.08 $Y=0
+ $X2=2.16 $Y2=0
r217 89 90 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.08 $Y=0
+ $X2=4.08 $Y2=0
r218 87 123 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.185 $Y=0
+ $X2=2.02 $Y2=0
r219 87 89 123.631 $w=1.68e-07 $l=1.895e-06 $layer=LI1_cond $X=2.185 $Y=0
+ $X2=4.08 $Y2=0
r220 86 126 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.41 $Y=0
+ $X2=4.535 $Y2=0
r221 86 89 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=4.41 $Y=0 $X2=4.08
+ $Y2=0
r222 85 124 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0
+ $X2=2.16 $Y2=0
r223 84 85 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r224 82 85 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r225 81 84 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r226 81 82 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r227 79 123 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.855 $Y=0
+ $X2=2.02 $Y2=0
r228 79 84 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=1.855 $Y=0
+ $X2=1.68 $Y2=0
r229 78 82 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r230 77 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r231 74 103 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=8.4
+ $Y2=0
r232 74 130 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.92 $Y=0
+ $X2=6.96 $Y2=0
r233 74 98 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r234 72 98 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=7.965 $Y=0 $X2=7.92
+ $Y2=0
r235 72 73 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.965 $Y=0 $X2=8.05
+ $Y2=0
r236 71 102 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=8.135 $Y=0
+ $X2=8.4 $Y2=0
r237 71 73 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.135 $Y=0 $X2=8.05
+ $Y2=0
r238 69 77 2.51176 $w=1.7e-07 $l=3.5e-08 $layer=LI1_cond $X=0.275 $Y=0 $X2=0.24
+ $Y2=0
r239 69 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.275 $Y=0 $X2=0.44
+ $Y2=0
r240 68 81 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=0.605 $Y=0
+ $X2=0.72 $Y2=0
r241 68 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.605 $Y=0 $X2=0.44
+ $Y2=0
r242 64 141 3.20777 $w=3.3e-07 $l=1.41244e-07 $layer=LI1_cond $X=15.465 $Y=0.085
+ $X2=15.57 $Y2=0
r243 64 66 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=15.465 $Y=0.085
+ $X2=15.465 $Y2=0.41
r244 60 138 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=14.605 $Y=0.085
+ $X2=14.605 $Y2=0
r245 60 62 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=14.605 $Y=0.085
+ $X2=14.605 $Y2=0.39
r246 56 135 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=13.745 $Y=0.085
+ $X2=13.745 $Y2=0
r247 56 58 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=13.745 $Y=0.085
+ $X2=13.745 $Y2=0.39
r248 52 132 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=11.91 $Y=0.085
+ $X2=11.91 $Y2=0
r249 52 54 26.3665 $w=3.28e-07 $l=7.55e-07 $layer=LI1_cond $X=11.91 $Y=0.085
+ $X2=11.91 $Y2=0.84
r250 48 50 21.7318 $w=3.48e-07 $l=6.6e-07 $layer=LI1_cond $X=8.49 $Y=1.01
+ $X2=9.15 $Y2=1.01
r251 46 48 11.6891 $w=3.48e-07 $l=3.55e-07 $layer=LI1_cond $X=8.135 $Y=1.01
+ $X2=8.49 $Y2=1.01
r252 45 46 7.93686 $w=3.5e-07 $l=2.13307e-07 $layer=LI1_cond $X=8.05 $Y=0.835
+ $X2=8.135 $Y2=1.01
r253 44 73 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.05 $Y=0.085
+ $X2=8.05 $Y2=0
r254 44 45 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=8.05 $Y=0.085
+ $X2=8.05 $Y2=0.835
r255 40 129 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.075 $Y=0.085
+ $X2=7.075 $Y2=0
r256 40 42 18.5089 $w=3.28e-07 $l=5.3e-07 $layer=LI1_cond $X=7.075 $Y=0.085
+ $X2=7.075 $Y2=0.615
r257 36 126 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.535 $Y=0.085
+ $X2=4.535 $Y2=0
r258 36 38 18.9001 $w=2.48e-07 $l=4.1e-07 $layer=LI1_cond $X=4.535 $Y=0.085
+ $X2=4.535 $Y2=0.495
r259 32 123 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.02 $Y=0.085
+ $X2=2.02 $Y2=0
r260 32 34 25.1442 $w=3.28e-07 $l=7.2e-07 $layer=LI1_cond $X=2.02 $Y=0.085
+ $X2=2.02 $Y2=0.805
r261 28 70 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.44 $Y=0.085
+ $X2=0.44 $Y2=0
r262 28 30 25.1442 $w=3.28e-07 $l=7.2e-07 $layer=LI1_cond $X=0.44 $Y=0.085
+ $X2=0.44 $Y2=0.805
r263 9 66 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=15.325
+ $Y=0.265 $X2=15.465 $Y2=0.41
r264 8 62 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=14.465
+ $Y=0.265 $X2=14.605 $Y2=0.39
r265 7 58 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=13.605
+ $Y=0.265 $X2=13.745 $Y2=0.39
r266 6 54 182 $w=1.7e-07 $l=2.96901e-07 $layer=licon1_NDIFF $count=1 $X=11.715
+ $Y=0.625 $X2=11.91 $Y2=0.84
r267 5 50 182 $w=1.7e-07 $l=9.75705e-07 $layer=licon1_NDIFF $count=1 $X=8.35
+ $Y=0.625 $X2=9.15 $Y2=1.015
r268 5 48 182 $w=1.7e-07 $l=3.58225e-07 $layer=licon1_NDIFF $count=1 $X=8.35
+ $Y=0.625 $X2=8.49 $Y2=0.92
r269 4 42 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=6.935
+ $Y=0.405 $X2=7.075 $Y2=0.615
r270 3 38 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=4.395
+ $Y=0.285 $X2=4.535 $Y2=0.495
r271 2 34 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.88
+ $Y=0.595 $X2=2.02 $Y2=0.805
r272 1 30 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.315
+ $Y=0.595 $X2=0.44 $Y2=0.805
.ends

