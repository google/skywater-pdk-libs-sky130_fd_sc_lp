* File: sky130_fd_sc_lp__dlxtp_1.pex.spice
* Created: Fri Aug 28 10:28:56 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__DLXTP_1%D 3 7 9 10 11 12 13 17
c34 17 0 1.68254e-19 $X=0.565 $Y=0.94
c35 11 0 8.46584e-20 $X=0.565 $Y=1.445
r36 17 18 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.565
+ $Y=0.94 $X2=0.565 $Y2=0.94
r37 13 18 11.8585 $w=3.43e-07 $l=3.55e-07 $layer=LI1_cond $X=0.642 $Y=1.295
+ $X2=0.642 $Y2=0.94
r38 12 18 0.501062 $w=3.43e-07 $l=1.5e-08 $layer=LI1_cond $X=0.642 $Y=0.925
+ $X2=0.642 $Y2=0.94
r39 10 17 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.565 $Y=1.28
+ $X2=0.565 $Y2=0.94
r40 10 11 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.565 $Y=1.28
+ $X2=0.565 $Y2=1.445
r41 9 17 40.8701 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.565 $Y=0.775
+ $X2=0.565 $Y2=0.94
r42 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.615 $Y=0.455
+ $X2=0.615 $Y2=0.775
r43 3 11 512.766 $w=1.5e-07 $l=1e-06 $layer=POLY_cond $X=0.475 $Y=2.445
+ $X2=0.475 $Y2=1.445
.ends

.subckt PM_SKY130_FD_SC_LP__DLXTP_1%GATE 3 7 9 12 14 17 19
c42 17 0 1.00661e-19 $X=1.135 $Y=0.94
c43 3 0 9.51503e-20 $X=0.905 $Y=2.445
r44 17 20 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.135 $Y=0.94
+ $X2=1.135 $Y2=1.105
r45 17 19 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.135 $Y=0.94
+ $X2=1.135 $Y2=0.775
r46 14 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.135
+ $Y=0.94 $X2=1.135 $Y2=0.94
r47 10 12 71.7872 $w=1.5e-07 $l=1.4e-07 $layer=POLY_cond $X=0.905 $Y=1.76
+ $X2=1.045 $Y2=1.76
r48 9 12 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.045 $Y=1.685
+ $X2=1.045 $Y2=1.76
r49 9 20 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=1.045 $Y=1.685
+ $X2=1.045 $Y2=1.105
r50 7 19 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.045 $Y=0.455
+ $X2=1.045 $Y2=0.775
r51 1 10 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.905 $Y=1.835
+ $X2=0.905 $Y2=1.76
r52 1 3 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=0.905 $Y=1.835
+ $X2=0.905 $Y2=2.445
.ends

.subckt PM_SKY130_FD_SC_LP__DLXTP_1%A_27_425# 1 2 9 13 16 19 21 23 28 30 31 35
+ 42
c85 42 0 2.72916e-19 $X=2.545 $Y=1.58
c86 35 0 4.61158e-20 $X=2.35 $Y=1.45
c87 31 0 8.46584e-20 $X=1.07 $Y=1.45
r88 42 43 4.56151 $w=3.17e-07 $l=3e-08 $layer=POLY_cond $X=2.545 $Y=1.58
+ $X2=2.575 $Y2=1.58
r89 39 42 24.3281 $w=3.17e-07 $l=1.6e-07 $layer=POLY_cond $X=2.385 $Y=1.58
+ $X2=2.545 $Y2=1.58
r90 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.385
+ $Y=1.58 $X2=2.385 $Y2=1.58
r91 35 38 5.76222 $w=2.58e-07 $l=1.3e-07 $layer=LI1_cond $X=2.35 $Y=1.45
+ $X2=2.35 $Y2=1.58
r92 31 33 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=1.07 $Y=1.45
+ $X2=1.07 $Y2=1.71
r93 25 28 7.05024 $w=3.38e-07 $l=2.08e-07 $layer=LI1_cond $X=0.192 $Y=0.435
+ $X2=0.4 $Y2=0.435
r94 24 31 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.155 $Y=1.45
+ $X2=1.07 $Y2=1.45
r95 23 35 3.22376 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.22 $Y=1.45 $X2=2.35
+ $Y2=1.45
r96 23 24 69.4813 $w=1.68e-07 $l=1.065e-06 $layer=LI1_cond $X=2.22 $Y=1.45
+ $X2=1.155 $Y2=1.45
r97 22 30 2.72405 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=0.365 $Y=1.71
+ $X2=0.225 $Y2=1.71
r98 21 33 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.985 $Y=1.71
+ $X2=1.07 $Y2=1.71
r99 21 22 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=0.985 $Y=1.71
+ $X2=0.365 $Y2=1.71
r100 17 30 3.74047 $w=2.47e-07 $l=8.5e-08 $layer=LI1_cond $X=0.225 $Y=1.795
+ $X2=0.225 $Y2=1.71
r101 17 19 19.5504 $w=2.78e-07 $l=4.75e-07 $layer=LI1_cond $X=0.225 $Y=1.795
+ $X2=0.225 $Y2=2.27
r102 16 30 3.74047 $w=2.47e-07 $l=1.0015e-07 $layer=LI1_cond $X=0.192 $Y=1.625
+ $X2=0.225 $Y2=1.71
r103 15 25 3.4367 $w=2.15e-07 $l=1.7e-07 $layer=LI1_cond $X=0.192 $Y=0.605
+ $X2=0.192 $Y2=0.435
r104 15 16 54.674 $w=2.13e-07 $l=1.02e-06 $layer=LI1_cond $X=0.192 $Y=0.605
+ $X2=0.192 $Y2=1.625
r105 11 43 20.269 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.575 $Y=1.415
+ $X2=2.575 $Y2=1.58
r106 11 13 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=2.575 $Y=1.415
+ $X2=2.575 $Y2=0.835
r107 7 42 20.269 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.545 $Y=1.745
+ $X2=2.545 $Y2=1.58
r108 7 9 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=2.545 $Y=1.745
+ $X2=2.545 $Y2=2.415
r109 2 19 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.125 $X2=0.26 $Y2=2.27
r110 1 28 182 $w=1.7e-07 $l=2.498e-07 $layer=licon1_NDIFF $count=1 $X=0.275
+ $Y=0.245 $X2=0.4 $Y2=0.44
.ends

.subckt PM_SKY130_FD_SC_LP__DLXTP_1%A_196_425# 1 2 8 9 10 13 14 17 19 23 24 28
+ 32 34 35 37 41 47 48 54 56 60
c105 47 0 4.61158e-20 $X=1.525 $Y=1.8
c106 37 0 9.51503e-20 $X=1.12 $Y=2.27
c107 35 0 1.77226e-19 $X=1.175 $Y=2.135
r108 59 60 30.474 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=2.055 $Y=0.44
+ $X2=2.055 $Y2=0.515
r109 48 51 3.58958 $w=3.03e-07 $l=9.5e-08 $layer=LI1_cond $X=1.272 $Y=0.345
+ $X2=1.272 $Y2=0.44
r110 47 55 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.525 $Y=1.8
+ $X2=1.525 $Y2=1.965
r111 47 54 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.525 $Y=1.8
+ $X2=1.525 $Y2=1.635
r112 46 47 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.525
+ $Y=1.8 $X2=1.525 $Y2=1.8
r113 42 59 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=2.055 $Y=0.35
+ $X2=2.055 $Y2=0.44
r114 42 56 29.7264 $w=3.3e-07 $l=1.7e-07 $layer=POLY_cond $X=2.055 $Y=0.35
+ $X2=2.055 $Y2=0.18
r115 41 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.055
+ $Y=0.35 $X2=2.055 $Y2=0.35
r116 39 48 3.82255 $w=1.8e-07 $l=1.53e-07 $layer=LI1_cond $X=1.425 $Y=0.345
+ $X2=1.272 $Y2=0.345
r117 39 41 38.8182 $w=1.78e-07 $l=6.3e-07 $layer=LI1_cond $X=1.425 $Y=0.345
+ $X2=2.055 $Y2=0.345
r118 35 46 13.9542 $w=3.06e-07 $l=4.44691e-07 $layer=LI1_cond $X=1.175 $Y=2.135
+ $X2=1.525 $Y2=1.92
r119 35 37 4.86187 $w=3.18e-07 $l=1.35e-07 $layer=LI1_cond $X=1.175 $Y=2.135
+ $X2=1.175 $Y2=2.27
r120 30 32 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=3.38 $Y=0.255
+ $X2=3.38 $Y2=0.835
r121 26 28 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.905 $Y=3.075
+ $X2=2.905 $Y2=2.415
r122 25 56 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.22 $Y=0.18
+ $X2=2.055 $Y2=0.18
r123 24 30 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.305 $Y=0.18
+ $X2=3.38 $Y2=0.255
r124 24 25 556.351 $w=1.5e-07 $l=1.085e-06 $layer=POLY_cond $X=3.305 $Y=0.18
+ $X2=2.22 $Y2=0.18
r125 23 60 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.145 $Y=0.835
+ $X2=2.145 $Y2=0.515
r126 20 34 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2 $Y=3.15 $X2=1.925
+ $Y2=3.15
r127 19 26 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.83 $Y=3.15
+ $X2=2.905 $Y2=3.075
r128 19 20 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=2.83 $Y=3.15 $X2=2
+ $Y2=3.15
r129 15 34 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.925 $Y=3.075
+ $X2=1.925 $Y2=3.15
r130 15 17 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=1.925 $Y=3.075
+ $X2=1.925 $Y2=2.625
r131 13 59 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.89 $Y=0.44
+ $X2=2.055 $Y2=0.44
r132 13 14 102.553 $w=1.5e-07 $l=2e-07 $layer=POLY_cond $X=1.89 $Y=0.44 $X2=1.69
+ $Y2=0.44
r133 11 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.615 $Y=0.515
+ $X2=1.69 $Y2=0.44
r134 11 54 574.298 $w=1.5e-07 $l=1.12e-06 $layer=POLY_cond $X=1.615 $Y=0.515
+ $X2=1.615 $Y2=1.635
r135 9 34 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.85 $Y=3.15
+ $X2=1.925 $Y2=3.15
r136 9 10 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=1.85 $Y=3.15 $X2=1.51
+ $Y2=3.15
r137 8 10 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.435 $Y=3.075
+ $X2=1.51 $Y2=3.15
r138 8 55 569.17 $w=1.5e-07 $l=1.11e-06 $layer=POLY_cond $X=1.435 $Y=3.075
+ $X2=1.435 $Y2=1.965
r139 2 37 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=0.98
+ $Y=2.125 $X2=1.12 $Y2=2.27
r140 1 51 182 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_NDIFF $count=1 $X=1.12
+ $Y=0.245 $X2=1.26 $Y2=0.44
.ends

.subckt PM_SKY130_FD_SC_LP__DLXTP_1%A_317_461# 1 2 9 13 19 21 23 24 26 28 30 34
+ 35
c88 28 0 1.64722e-19 $X=2.735 $Y=2.305
r89 35 37 15.3286 $w=2.83e-07 $l=9e-08 $layer=POLY_cond $X=3.025 $Y=1.65
+ $X2=2.935 $Y2=1.65
r90 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.025
+ $Y=1.56 $X2=3.025 $Y2=1.56
r91 31 34 10.1275 $w=3.28e-07 $l=2.9e-07 $layer=LI1_cond $X=2.735 $Y=1.56
+ $X2=3.025 $Y2=1.56
r92 27 31 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.735 $Y=1.725
+ $X2=2.735 $Y2=1.56
r93 27 28 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=2.735 $Y=1.725
+ $X2=2.735 $Y2=2.305
r94 26 31 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.735 $Y=1.395
+ $X2=2.735 $Y2=1.56
r95 25 26 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=2.735 $Y=1.185
+ $X2=2.735 $Y2=1.395
r96 23 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.65 $Y=1.1
+ $X2=2.735 $Y2=1.185
r97 23 24 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=2.65 $Y=1.1
+ $X2=2.025 $Y2=1.1
r98 22 30 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.875 $Y=2.39
+ $X2=1.71 $Y2=2.39
r99 21 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.65 $Y=2.39
+ $X2=2.735 $Y2=2.305
r100 21 22 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=2.65 $Y=2.39
+ $X2=1.875 $Y2=2.39
r101 17 24 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=1.895 $Y=1.015
+ $X2=2.025 $Y2=1.1
r102 17 19 7.75683 $w=2.58e-07 $l=1.75e-07 $layer=LI1_cond $X=1.895 $Y=1.015
+ $X2=1.895 $Y2=0.84
r103 11 35 68.9788 $w=2.83e-07 $l=5.17011e-07 $layer=POLY_cond $X=3.43 $Y=1.905
+ $X2=3.025 $Y2=1.65
r104 11 13 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=3.43 $Y=1.905
+ $X2=3.43 $Y2=2.305
r105 7 37 17.601 $w=1.5e-07 $l=2.55e-07 $layer=POLY_cond $X=2.935 $Y=1.395
+ $X2=2.935 $Y2=1.65
r106 7 9 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=2.935 $Y=1.395
+ $X2=2.935 $Y2=0.835
r107 2 30 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=1.585
+ $Y=2.305 $X2=1.71 $Y2=2.45
r108 1 19 182 $w=1.7e-07 $l=2.7037e-07 $layer=licon1_NDIFF $count=1 $X=1.805
+ $Y=0.625 $X2=1.93 $Y2=0.84
.ends

.subckt PM_SKY130_FD_SC_LP__DLXTP_1%A_733_99# 1 2 9 13 17 20 24 25 27 28 31 34
+ 38 42 45 50
c89 45 0 1.83405e-19 $X=5.13 $Y=1.43
c90 25 0 1.4427e-19 $X=3.83 $Y=1.35
r91 45 51 45.5639 $w=3.95e-07 $l=1.65e-07 $layer=POLY_cond $X=5.162 $Y=1.43
+ $X2=5.162 $Y2=1.595
r92 45 50 45.5639 $w=3.95e-07 $l=1.65e-07 $layer=POLY_cond $X=5.162 $Y=1.43
+ $X2=5.162 $Y2=1.265
r93 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.13
+ $Y=1.43 $X2=5.13 $Y2=1.43
r94 42 44 14.2102 $w=3.52e-07 $l=4.1e-07 $layer=LI1_cond $X=4.72 $Y=1.565
+ $X2=5.13 $Y2=1.565
r95 41 42 5.89205 $w=3.52e-07 $l=3.70371e-07 $layer=LI1_cond $X=4.55 $Y=1.86
+ $X2=4.72 $Y2=1.565
r96 36 38 7.62646 $w=3.38e-07 $l=2.25e-07 $layer=LI1_cond $X=4.495 $Y=0.455
+ $X2=4.72 $Y2=0.455
r97 34 42 5.00804 $w=1.7e-07 $l=3e-07 $layer=LI1_cond $X=4.72 $Y=1.265 $X2=4.72
+ $Y2=1.565
r98 33 38 4.80115 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=4.72 $Y=0.625
+ $X2=4.72 $Y2=0.455
r99 33 34 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=4.72 $Y=0.625
+ $X2=4.72 $Y2=1.265
r100 29 41 2.51309 $w=2.6e-07 $l=3.74166e-08 $layer=LI1_cond $X=4.585 $Y=1.865
+ $X2=4.55 $Y2=1.86
r101 29 31 40.7788 $w=2.58e-07 $l=9.2e-07 $layer=LI1_cond $X=4.585 $Y=1.865
+ $X2=4.585 $Y2=2.785
r102 27 41 6.56424 $w=3.52e-07 $l=1.28938e-07 $layer=LI1_cond $X=4.455 $Y=1.78
+ $X2=4.55 $Y2=1.86
r103 27 28 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=4.455 $Y=1.78
+ $X2=3.995 $Y2=1.78
r104 25 48 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.83 $Y=1.35
+ $X2=3.83 $Y2=1.515
r105 25 47 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.83 $Y=1.35
+ $X2=3.83 $Y2=1.185
r106 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.83
+ $Y=1.35 $X2=3.83 $Y2=1.35
r107 22 28 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.83 $Y=1.695
+ $X2=3.995 $Y2=1.78
r108 22 24 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=3.83 $Y=1.695
+ $X2=3.83 $Y2=1.35
r109 20 51 446.106 $w=1.5e-07 $l=8.7e-07 $layer=POLY_cond $X=5.285 $Y=2.465
+ $X2=5.285 $Y2=1.595
r110 17 50 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=5.285 $Y=0.735
+ $X2=5.285 $Y2=1.265
r111 13 48 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.79 $Y=2.305
+ $X2=3.79 $Y2=1.515
r112 9 47 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=3.74 $Y=0.835
+ $X2=3.74 $Y2=1.185
r113 2 41 400 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_PDIFF $count=1 $X=4.41
+ $Y=1.675 $X2=4.55 $Y2=1.86
r114 2 31 400 $w=1.7e-07 $l=1.17792e-06 $layer=licon1_PDIFF $count=1 $X=4.41
+ $Y=1.675 $X2=4.55 $Y2=2.785
r115 1 36 182 $w=1.7e-07 $l=2.86575e-07 $layer=licon1_NDIFF $count=1 $X=4.355
+ $Y=0.235 $X2=4.495 $Y2=0.46
.ends

.subckt PM_SKY130_FD_SC_LP__DLXTP_1%A_596_419# 1 2 9 12 14 22 26 27 30 31 32 34
c80 31 0 9.56904e-20 $X=3.237 $Y=2.075
c81 26 0 1.83405e-19 $X=4.37 $Y=1.35
r82 30 31 8.86124 $w=4.43e-07 $l=1.65e-07 $layer=LI1_cond $X=3.237 $Y=2.24
+ $X2=3.237 $Y2=2.075
r83 27 35 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.37 $Y=1.35
+ $X2=4.37 $Y2=1.515
r84 27 34 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.37 $Y=1.35
+ $X2=4.37 $Y2=1.185
r85 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.37
+ $Y=1.35 $X2=4.37 $Y2=1.35
r86 24 26 15.292 $w=2.58e-07 $l=3.45e-07 $layer=LI1_cond $X=4.335 $Y=1.005
+ $X2=4.335 $Y2=1.35
r87 23 32 4.3182 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=3.46 $Y=0.9 $X2=3.375
+ $Y2=0.9
r88 22 24 6.91731 $w=2.1e-07 $l=1.74786e-07 $layer=LI1_cond $X=4.205 $Y=0.9
+ $X2=4.335 $Y2=1.005
r89 22 23 39.3463 $w=2.08e-07 $l=7.45e-07 $layer=LI1_cond $X=4.205 $Y=0.9
+ $X2=3.46 $Y2=0.9
r90 20 32 2.11342 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=3.375 $Y=1.005
+ $X2=3.375 $Y2=0.9
r91 20 31 69.8075 $w=1.68e-07 $l=1.07e-06 $layer=LI1_cond $X=3.375 $Y=1.005
+ $X2=3.375 $Y2=2.075
r92 14 32 4.3182 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=3.29 $Y=0.9 $X2=3.375
+ $Y2=0.9
r93 14 16 6.60173 $w=2.08e-07 $l=1.25e-07 $layer=LI1_cond $X=3.29 $Y=0.9
+ $X2=3.165 $Y2=0.9
r94 12 35 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=4.335 $Y=2.305
+ $X2=4.335 $Y2=1.515
r95 9 34 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=4.28 $Y=0.655
+ $X2=4.28 $Y2=1.185
r96 2 30 300 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_PDIFF $count=2 $X=2.98
+ $Y=2.095 $X2=3.18 $Y2=2.24
r97 1 16 182 $w=1.7e-07 $l=3.43875e-07 $layer=licon1_NDIFF $count=1 $X=3.01
+ $Y=0.625 $X2=3.165 $Y2=0.9
.ends

.subckt PM_SKY130_FD_SC_LP__DLXTP_1%VPWR 1 2 3 4 15 19 23 27 30 33 35 40 45 53
+ 60 61 64 67 70 73
c80 23 0 1.4427e-19 $X=4.12 $Y=2.12
r81 73 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r82 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r83 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r84 64 65 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r85 61 74 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=5.04 $Y2=3.33
r86 60 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r87 58 73 8.23795 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=5.215 $Y=3.33
+ $X2=5.06 $Y2=3.33
r88 58 60 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=5.215 $Y=3.33
+ $X2=5.52 $Y2=3.33
r89 57 74 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.04 $Y2=3.33
r90 57 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=4.08 $Y2=3.33
r91 56 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r92 54 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.285 $Y=3.33
+ $X2=4.12 $Y2=3.33
r93 54 56 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=4.285 $Y=3.33
+ $X2=4.56 $Y2=3.33
r94 53 73 8.23795 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=4.905 $Y=3.33
+ $X2=5.06 $Y2=3.33
r95 53 56 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=4.905 $Y=3.33
+ $X2=4.56 $Y2=3.33
r96 52 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r97 51 52 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r98 49 68 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r99 48 51 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.64 $Y=3.33 $X2=3.6
+ $Y2=3.33
r100 48 49 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r101 46 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.4 $Y=3.33
+ $X2=2.235 $Y2=3.33
r102 46 48 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=2.4 $Y=3.33
+ $X2=2.64 $Y2=3.33
r103 45 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.955 $Y=3.33
+ $X2=4.12 $Y2=3.33
r104 45 51 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=3.955 $Y=3.33
+ $X2=3.6 $Y2=3.33
r105 44 68 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r106 44 65 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.72 $Y2=3.33
r107 43 44 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r108 41 64 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=0.795 $Y=3.33
+ $X2=0.69 $Y2=3.33
r109 41 43 57.738 $w=1.68e-07 $l=8.85e-07 $layer=LI1_cond $X=0.795 $Y=3.33
+ $X2=1.68 $Y2=3.33
r110 40 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.07 $Y=3.33
+ $X2=2.235 $Y2=3.33
r111 40 43 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=2.07 $Y=3.33
+ $X2=1.68 $Y2=3.33
r112 38 65 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r113 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r114 35 64 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=0.585 $Y=3.33
+ $X2=0.69 $Y2=3.33
r115 35 37 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.585 $Y=3.33
+ $X2=0.24 $Y2=3.33
r116 33 52 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.88 $Y=3.33
+ $X2=3.6 $Y2=3.33
r117 33 49 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.88 $Y=3.33
+ $X2=2.64 $Y2=3.33
r118 28 73 0.701276 $w=3.1e-07 $l=8.5e-08 $layer=LI1_cond $X=5.06 $Y=3.245
+ $X2=5.06 $Y2=3.33
r119 28 30 29.5546 $w=3.08e-07 $l=7.95e-07 $layer=LI1_cond $X=5.06 $Y=3.245
+ $X2=5.06 $Y2=2.45
r120 27 32 8.52182 $w=3.1e-07 $l=2.1e-07 $layer=LI1_cond $X=5.06 $Y=2.19
+ $X2=5.06 $Y2=1.98
r121 27 30 9.66565 $w=3.08e-07 $l=2.6e-07 $layer=LI1_cond $X=5.06 $Y=2.19
+ $X2=5.06 $Y2=2.45
r122 23 26 12.2229 $w=3.28e-07 $l=3.5e-07 $layer=LI1_cond $X=4.12 $Y=2.12
+ $X2=4.12 $Y2=2.47
r123 21 70 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.12 $Y=3.245
+ $X2=4.12 $Y2=3.33
r124 21 26 27.0649 $w=3.28e-07 $l=7.75e-07 $layer=LI1_cond $X=4.12 $Y=3.245
+ $X2=4.12 $Y2=2.47
r125 17 67 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.235 $Y=3.245
+ $X2=2.235 $Y2=3.33
r126 17 19 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=2.235 $Y=3.245
+ $X2=2.235 $Y2=2.75
r127 13 64 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=3.245
+ $X2=0.69 $Y2=3.33
r128 13 15 49.9091 $w=2.08e-07 $l=9.45e-07 $layer=LI1_cond $X=0.69 $Y=3.245
+ $X2=0.69 $Y2=2.3
r129 4 32 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=4.945
+ $Y=1.835 $X2=5.07 $Y2=1.98
r130 4 30 300 $w=1.7e-07 $l=6.74611e-07 $layer=licon1_PDIFF $count=2 $X=4.945
+ $Y=1.835 $X2=5.07 $Y2=2.45
r131 3 26 300 $w=1.7e-07 $l=4.86056e-07 $layer=licon1_PDIFF $count=2 $X=3.865
+ $Y=2.095 $X2=4.12 $Y2=2.47
r132 3 23 600 $w=1.7e-07 $l=2.67208e-07 $layer=licon1_PDIFF $count=1 $X=3.865
+ $Y=2.095 $X2=4.12 $Y2=2.12
r133 2 19 600 $w=1.7e-07 $l=5.50091e-07 $layer=licon1_PDIFF $count=1 $X=2
+ $Y=2.305 $X2=2.235 $Y2=2.75
r134 1 15 300 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_PDIFF $count=2 $X=0.55
+ $Y=2.125 $X2=0.69 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_LP__DLXTP_1%Q 1 2 7 8 9 10 11 12 13 22
r12 13 40 5.36482 $w=2.88e-07 $l=1.35e-07 $layer=LI1_cond $X=5.53 $Y=2.775
+ $X2=5.53 $Y2=2.91
r13 12 13 14.7036 $w=2.88e-07 $l=3.7e-07 $layer=LI1_cond $X=5.53 $Y=2.405
+ $X2=5.53 $Y2=2.775
r14 11 12 16.8893 $w=2.88e-07 $l=4.25e-07 $layer=LI1_cond $X=5.53 $Y=1.98
+ $X2=5.53 $Y2=2.405
r15 10 11 12.5179 $w=2.88e-07 $l=3.15e-07 $layer=LI1_cond $X=5.53 $Y=1.665
+ $X2=5.53 $Y2=1.98
r16 9 10 14.7036 $w=2.88e-07 $l=3.7e-07 $layer=LI1_cond $X=5.53 $Y=1.295
+ $X2=5.53 $Y2=1.665
r17 8 9 14.7036 $w=2.88e-07 $l=3.7e-07 $layer=LI1_cond $X=5.53 $Y=0.925 $X2=5.53
+ $Y2=1.295
r18 7 8 14.7036 $w=2.88e-07 $l=3.7e-07 $layer=LI1_cond $X=5.53 $Y=0.555 $X2=5.53
+ $Y2=0.925
r19 7 22 3.77524 $w=2.88e-07 $l=9.5e-08 $layer=LI1_cond $X=5.53 $Y=0.555
+ $X2=5.53 $Y2=0.46
r20 2 40 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=5.36
+ $Y=1.835 $X2=5.5 $Y2=2.91
r21 2 11 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=5.36
+ $Y=1.835 $X2=5.5 $Y2=1.98
r22 1 22 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.36
+ $Y=0.315 $X2=5.5 $Y2=0.46
.ends

.subckt PM_SKY130_FD_SC_LP__DLXTP_1%VGND 1 2 3 4 17 20 23 25 29 34 37 38 39 48
+ 57 58 61 64 67
c78 61 0 1.68254e-19 $X=0.72 $Y=0
c79 37 0 1.00661e-19 $X=2.4 $Y=0
r80 67 68 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r81 65 68 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=5.04
+ $Y2=0
r82 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r83 61 62 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r84 58 68 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=5.04
+ $Y2=0
r85 57 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r86 55 67 6.81202 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=5.215 $Y=0 $X2=5.095
+ $Y2=0
r87 55 57 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=5.215 $Y=0 $X2=5.52
+ $Y2=0
r88 54 65 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r89 53 54 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r90 50 53 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r91 50 51 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r92 48 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.9 $Y=0 $X2=4.065
+ $Y2=0
r93 48 53 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=3.9 $Y=0 $X2=3.6 $Y2=0
r94 47 51 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r95 46 47 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r96 44 47 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r97 44 62 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r98 43 46 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r99 43 44 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r100 41 61 6.92067 $w=1.7e-07 $l=1.23e-07 $layer=LI1_cond $X=0.95 $Y=0 $X2=0.827
+ $Y2=0
r101 41 43 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=0.95 $Y=0 $X2=1.2
+ $Y2=0
r102 39 54 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.88 $Y=0 $X2=3.6
+ $Y2=0
r103 39 51 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.88 $Y=0
+ $X2=2.64 $Y2=0
r104 37 46 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=2.4 $Y=0 $X2=2.16
+ $Y2=0
r105 37 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.4 $Y=0 $X2=2.485
+ $Y2=0
r106 36 50 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=2.57 $Y=0 $X2=2.64
+ $Y2=0
r107 36 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.57 $Y=0 $X2=2.485
+ $Y2=0
r108 32 34 6.00231 $w=2.38e-07 $l=1.25e-07 $layer=LI1_cond $X=2.36 $Y=0.725
+ $X2=2.485 $Y2=0.725
r109 27 67 0.135687 $w=2.4e-07 $l=8.5e-08 $layer=LI1_cond $X=5.095 $Y=0.085
+ $X2=5.095 $Y2=0
r110 27 29 18.0069 $w=2.38e-07 $l=3.75e-07 $layer=LI1_cond $X=5.095 $Y=0.085
+ $X2=5.095 $Y2=0.46
r111 26 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.23 $Y=0 $X2=4.065
+ $Y2=0
r112 25 67 6.81202 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=4.975 $Y=0 $X2=5.095
+ $Y2=0
r113 25 26 48.6043 $w=1.68e-07 $l=7.45e-07 $layer=LI1_cond $X=4.975 $Y=0
+ $X2=4.23 $Y2=0
r114 21 64 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.065 $Y=0.085
+ $X2=4.065 $Y2=0
r115 21 23 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=4.065 $Y=0.085
+ $X2=4.065 $Y2=0.5
r116 20 34 2.75731 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=2.485 $Y=0.605
+ $X2=2.485 $Y2=0.725
r117 19 38 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.485 $Y=0.085
+ $X2=2.485 $Y2=0
r118 19 20 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=2.485 $Y=0.085
+ $X2=2.485 $Y2=0.605
r119 15 61 0.066131 $w=2.45e-07 $l=8.5e-08 $layer=LI1_cond $X=0.827 $Y=0.085
+ $X2=0.827 $Y2=0
r120 15 17 16.6987 $w=2.43e-07 $l=3.55e-07 $layer=LI1_cond $X=0.827 $Y=0.085
+ $X2=0.827 $Y2=0.44
r121 4 29 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=4.945
+ $Y=0.315 $X2=5.07 $Y2=0.46
r122 3 23 182 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_NDIFF $count=1 $X=3.815
+ $Y=0.625 $X2=4.065 $Y2=0.5
r123 2 32 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=2.22
+ $Y=0.625 $X2=2.36 $Y2=0.75
r124 1 17 182 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_NDIFF $count=1 $X=0.69
+ $Y=0.245 $X2=0.83 $Y2=0.44
.ends

