* File: sky130_fd_sc_lp__o41a_2.pxi.spice
* Created: Wed Sep  2 10:27:33 2020
* 
x_PM_SKY130_FD_SC_LP__O41A_2%A_102_53# N_A_102_53#_M1004_s N_A_102_53#_M1007_d
+ N_A_102_53#_c_74_n N_A_102_53#_M1000_g N_A_102_53#_M1003_g N_A_102_53#_c_75_n
+ N_A_102_53#_M1011_g N_A_102_53#_M1013_g N_A_102_53#_c_76_n N_A_102_53#_c_121_p
+ N_A_102_53#_c_77_n N_A_102_53#_c_78_n N_A_102_53#_c_85_n N_A_102_53#_c_87_p
+ N_A_102_53#_c_79_n N_A_102_53#_c_80_n N_A_102_53#_c_88_p N_A_102_53#_c_89_p
+ PM_SKY130_FD_SC_LP__O41A_2%A_102_53#
x_PM_SKY130_FD_SC_LP__O41A_2%B1 N_B1_M1007_g N_B1_c_162_n N_B1_M1004_g B1 B1
+ N_B1_c_164_n PM_SKY130_FD_SC_LP__O41A_2%B1
x_PM_SKY130_FD_SC_LP__O41A_2%A4 N_A4_M1010_g N_A4_M1008_g A4 A4 N_A4_c_202_n
+ N_A4_c_203_n PM_SKY130_FD_SC_LP__O41A_2%A4
x_PM_SKY130_FD_SC_LP__O41A_2%A3 N_A3_M1009_g N_A3_M1006_g A3 A3 A3 A3
+ N_A3_c_246_n N_A3_c_247_n PM_SKY130_FD_SC_LP__O41A_2%A3
x_PM_SKY130_FD_SC_LP__O41A_2%A2 N_A2_M1012_g N_A2_M1001_g A2 A2 A2 A2
+ N_A2_c_285_n N_A2_c_286_n PM_SKY130_FD_SC_LP__O41A_2%A2
x_PM_SKY130_FD_SC_LP__O41A_2%A1 N_A1_M1002_g N_A1_M1005_g A1 N_A1_c_322_n
+ N_A1_c_323_n PM_SKY130_FD_SC_LP__O41A_2%A1
x_PM_SKY130_FD_SC_LP__O41A_2%VPWR N_VPWR_M1003_d N_VPWR_M1013_d N_VPWR_M1005_d
+ N_VPWR_c_346_n N_VPWR_c_347_n N_VPWR_c_358_n N_VPWR_c_348_n N_VPWR_c_349_n
+ N_VPWR_c_350_n N_VPWR_c_367_n VPWR N_VPWR_c_351_n N_VPWR_c_352_n
+ N_VPWR_c_353_n N_VPWR_c_345_n PM_SKY130_FD_SC_LP__O41A_2%VPWR
x_PM_SKY130_FD_SC_LP__O41A_2%X N_X_M1000_s N_X_M1003_s X X X X X X X
+ PM_SKY130_FD_SC_LP__O41A_2%X
x_PM_SKY130_FD_SC_LP__O41A_2%VGND N_VGND_M1000_d N_VGND_M1011_d N_VGND_M1010_d
+ N_VGND_M1012_d N_VGND_c_428_n N_VGND_c_429_n N_VGND_c_430_n N_VGND_c_431_n
+ N_VGND_c_432_n N_VGND_c_433_n N_VGND_c_434_n N_VGND_c_435_n N_VGND_c_436_n
+ VGND N_VGND_c_437_n N_VGND_c_438_n N_VGND_c_439_n N_VGND_c_440_n
+ PM_SKY130_FD_SC_LP__O41A_2%VGND
x_PM_SKY130_FD_SC_LP__O41A_2%A_465_49# N_A_465_49#_M1004_d N_A_465_49#_M1006_d
+ N_A_465_49#_M1002_d N_A_465_49#_c_491_n N_A_465_49#_c_486_n
+ N_A_465_49#_c_487_n N_A_465_49#_c_503_n N_A_465_49#_c_488_n
+ N_A_465_49#_c_489_n N_A_465_49#_c_490_n PM_SKY130_FD_SC_LP__O41A_2%A_465_49#
cc_1 VNB N_A_102_53#_c_74_n 0.0187244f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.345
cc_2 VNB N_A_102_53#_c_75_n 0.0187429f $X=-0.19 $Y=-0.245 $X2=1.015 $Y2=1.345
cc_3 VNB N_A_102_53#_c_76_n 0.0390751f $X=-0.19 $Y=-0.245 $X2=1.09 $Y2=1.51
cc_4 VNB N_A_102_53#_c_77_n 0.042903f $X=-0.19 $Y=-0.245 $X2=1.495 $Y2=1.51
cc_5 VNB N_A_102_53#_c_78_n 0.00743151f $X=-0.19 $Y=-0.245 $X2=1.757 $Y2=1.345
cc_6 VNB N_A_102_53#_c_79_n 0.0175126f $X=-0.19 $Y=-0.245 $X2=2.035 $Y2=0.39
cc_7 VNB N_A_102_53#_c_80_n 0.0023602f $X=-0.19 $Y=-0.245 $X2=1.757 $Y2=1.51
cc_8 VNB N_B1_M1007_g 0.0061156f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_B1_c_162_n 0.02108f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB B1 0.0018365f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=0.815
cc_11 VNB N_B1_c_164_n 0.0394151f $X=-0.19 $Y=-0.245 $X2=1.015 $Y2=1.675
cc_12 VNB N_A4_M1010_g 0.0258459f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A4_c_202_n 0.0251432f $X=-0.19 $Y=-0.245 $X2=1.015 $Y2=1.345
cc_14 VNB N_A4_c_203_n 0.00378369f $X=-0.19 $Y=-0.245 $X2=1.015 $Y2=0.815
cc_15 VNB N_A3_M1006_g 0.025201f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.345
cc_16 VNB N_A3_c_246_n 0.0239673f $X=-0.19 $Y=-0.245 $X2=1.015 $Y2=2.465
cc_17 VNB N_A3_c_247_n 0.00371614f $X=-0.19 $Y=-0.245 $X2=1.015 $Y2=2.465
cc_18 VNB N_A2_M1012_g 0.025264f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A2_c_285_n 0.0223114f $X=-0.19 $Y=-0.245 $X2=1.495 $Y2=1.51
cc_20 VNB N_A2_c_286_n 0.00662975f $X=-0.19 $Y=-0.245 $X2=1.495 $Y2=1.51
cc_21 VNB N_A1_M1002_g 0.0296317f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A1_M1005_g 0.00137264f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.345
cc_23 VNB N_A1_c_322_n 0.0618679f $X=-0.19 $Y=-0.245 $X2=1.015 $Y2=1.345
cc_24 VNB N_A1_c_323_n 0.0012933f $X=-0.19 $Y=-0.245 $X2=1.015 $Y2=0.815
cc_25 VNB N_VPWR_c_345_n 0.203486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB X 0.0032792f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.345
cc_27 VNB N_VGND_c_428_n 0.0137412f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_429_n 0.0497502f $X=-0.19 $Y=-0.245 $X2=1.015 $Y2=0.815
cc_29 VNB N_VGND_c_430_n 0.0163188f $X=-0.19 $Y=-0.245 $X2=1.015 $Y2=2.465
cc_30 VNB N_VGND_c_431_n 0.00530065f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_432_n 0.00530084f $X=-0.19 $Y=-0.245 $X2=1.495 $Y2=1.51
cc_32 VNB N_VGND_c_433_n 0.0377247f $X=-0.19 $Y=-0.245 $X2=1.757 $Y2=1.04
cc_33 VNB N_VGND_c_434_n 0.00634081f $X=-0.19 $Y=-0.245 $X2=1.757 $Y2=1.345
cc_34 VNB N_VGND_c_435_n 0.017273f $X=-0.19 $Y=-0.245 $X2=1.757 $Y2=1.96
cc_35 VNB N_VGND_c_436_n 0.00634081f $X=-0.19 $Y=-0.245 $X2=2.197 $Y2=2.14
cc_36 VNB N_VGND_c_437_n 0.0171105f $X=-0.19 $Y=-0.245 $X2=2.035 $Y2=0.39
cc_37 VNB N_VGND_c_438_n 0.0204354f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_439_n 0.278351f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_440_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_465_49#_c_486_n 0.00627992f $X=-0.19 $Y=-0.245 $X2=1.015 $Y2=1.345
cc_41 VNB N_A_465_49#_c_487_n 0.00488348f $X=-0.19 $Y=-0.245 $X2=1.015 $Y2=0.815
cc_42 VNB N_A_465_49#_c_488_n 0.0125442f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_465_49#_c_489_n 0.0290655f $X=-0.19 $Y=-0.245 $X2=1.015 $Y2=1.51
cc_44 VNB N_A_465_49#_c_490_n 0.00561742f $X=-0.19 $Y=-0.245 $X2=1.495 $Y2=1.51
cc_45 VPB N_A_102_53#_M1003_g 0.0249072f $X=-0.19 $Y=1.655 $X2=0.585 $Y2=2.465
cc_46 VPB N_A_102_53#_M1013_g 0.0222849f $X=-0.19 $Y=1.655 $X2=1.015 $Y2=2.465
cc_47 VPB N_A_102_53#_c_76_n 0.00519541f $X=-0.19 $Y=1.655 $X2=1.09 $Y2=1.51
cc_48 VPB N_A_102_53#_c_77_n 0.0169199f $X=-0.19 $Y=1.655 $X2=1.495 $Y2=1.51
cc_49 VPB N_A_102_53#_c_85_n 0.00360655f $X=-0.19 $Y=1.655 $X2=1.757 $Y2=1.96
cc_50 VPB N_B1_M1007_g 0.0258354f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_51 VPB B1 0.00233675f $X=-0.19 $Y=1.655 $X2=0.585 $Y2=0.815
cc_52 VPB N_A4_M1008_g 0.0203311f $X=-0.19 $Y=1.655 $X2=0.585 $Y2=1.345
cc_53 VPB N_A4_c_202_n 0.00654804f $X=-0.19 $Y=1.655 $X2=1.015 $Y2=1.345
cc_54 VPB N_A4_c_203_n 0.00167067f $X=-0.19 $Y=1.655 $X2=1.015 $Y2=0.815
cc_55 VPB N_A3_M1009_g 0.0177506f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_56 VPB N_A3_c_246_n 0.00824058f $X=-0.19 $Y=1.655 $X2=1.015 $Y2=2.465
cc_57 VPB N_A3_c_247_n 0.00210806f $X=-0.19 $Y=1.655 $X2=1.015 $Y2=2.465
cc_58 VPB N_A2_M1001_g 0.0197733f $X=-0.19 $Y=1.655 $X2=0.585 $Y2=1.345
cc_59 VPB N_A2_c_285_n 0.00625343f $X=-0.19 $Y=1.655 $X2=1.495 $Y2=1.51
cc_60 VPB N_A2_c_286_n 0.00115564f $X=-0.19 $Y=1.655 $X2=1.495 $Y2=1.51
cc_61 VPB N_A1_M1005_g 0.0257099f $X=-0.19 $Y=1.655 $X2=0.585 $Y2=1.345
cc_62 VPB N_A1_c_323_n 0.0089038f $X=-0.19 $Y=1.655 $X2=1.015 $Y2=0.815
cc_63 VPB N_VPWR_c_346_n 0.013712f $X=-0.19 $Y=1.655 $X2=0.585 $Y2=1.675
cc_64 VPB N_VPWR_c_347_n 0.0568716f $X=-0.19 $Y=1.655 $X2=0.585 $Y2=2.465
cc_65 VPB N_VPWR_c_348_n 0.00550473f $X=-0.19 $Y=1.655 $X2=1.09 $Y2=1.51
cc_66 VPB N_VPWR_c_349_n 0.0132697f $X=-0.19 $Y=1.655 $X2=0.585 $Y2=1.51
cc_67 VPB N_VPWR_c_350_n 0.0495344f $X=-0.19 $Y=1.655 $X2=1.015 $Y2=1.51
cc_68 VPB N_VPWR_c_351_n 0.0154314f $X=-0.19 $Y=1.655 $X2=1.757 $Y2=1.96
cc_69 VPB N_VPWR_c_352_n 0.0634983f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_70 VPB N_VPWR_c_353_n 0.0147669f $X=-0.19 $Y=1.655 $X2=1.495 $Y2=1.51
cc_71 VPB N_VPWR_c_345_n 0.0523956f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_72 VPB X 0.00151789f $X=-0.19 $Y=1.655 $X2=0.585 $Y2=1.345
cc_73 N_A_102_53#_c_85_n N_B1_M1007_g 0.00649141f $X=1.757 $Y=1.96 $X2=0 $Y2=0
cc_74 N_A_102_53#_c_87_p N_B1_M1007_g 0.0176448f $X=2.197 $Y=2.14 $X2=0 $Y2=0
cc_75 N_A_102_53#_c_88_p N_B1_M1007_g 0.00941422f $X=2.575 $Y=2.495 $X2=0 $Y2=0
cc_76 N_A_102_53#_c_89_p N_B1_M1007_g 0.00390647f $X=2.405 $Y=2.33 $X2=0 $Y2=0
cc_77 N_A_102_53#_c_78_n N_B1_c_162_n 0.00319002f $X=1.757 $Y=1.345 $X2=0 $Y2=0
cc_78 N_A_102_53#_c_79_n N_B1_c_162_n 0.0132101f $X=2.035 $Y=0.39 $X2=0 $Y2=0
cc_79 N_A_102_53#_c_77_n B1 2.40288e-19 $X=1.495 $Y=1.51 $X2=0 $Y2=0
cc_80 N_A_102_53#_c_78_n B1 0.0100775f $X=1.757 $Y=1.345 $X2=0 $Y2=0
cc_81 N_A_102_53#_c_85_n B1 0.00558065f $X=1.757 $Y=1.96 $X2=0 $Y2=0
cc_82 N_A_102_53#_c_87_p B1 0.011187f $X=2.197 $Y=2.14 $X2=0 $Y2=0
cc_83 N_A_102_53#_c_79_n B1 0.00875283f $X=2.035 $Y=0.39 $X2=0 $Y2=0
cc_84 N_A_102_53#_c_80_n B1 0.0267808f $X=1.757 $Y=1.51 $X2=0 $Y2=0
cc_85 N_A_102_53#_c_77_n N_B1_c_164_n 0.0134824f $X=1.495 $Y=1.51 $X2=0 $Y2=0
cc_86 N_A_102_53#_c_78_n N_B1_c_164_n 0.00363476f $X=1.757 $Y=1.345 $X2=0 $Y2=0
cc_87 N_A_102_53#_c_87_p N_B1_c_164_n 0.0028625f $X=2.197 $Y=2.14 $X2=0 $Y2=0
cc_88 N_A_102_53#_c_79_n N_B1_c_164_n 0.00654187f $X=2.035 $Y=0.39 $X2=0 $Y2=0
cc_89 N_A_102_53#_c_80_n N_B1_c_164_n 0.0029107f $X=1.757 $Y=1.51 $X2=0 $Y2=0
cc_90 N_A_102_53#_c_79_n N_A4_M1010_g 3.1246e-19 $X=2.035 $Y=0.39 $X2=0 $Y2=0
cc_91 N_A_102_53#_c_87_p N_A4_M1008_g 5.24242e-19 $X=2.197 $Y=2.14 $X2=0 $Y2=0
cc_92 N_A_102_53#_c_88_p N_A4_M1008_g 0.0112541f $X=2.575 $Y=2.495 $X2=0 $Y2=0
cc_93 N_A_102_53#_c_89_p N_A4_M1008_g 0.00155815f $X=2.405 $Y=2.33 $X2=0 $Y2=0
cc_94 N_A_102_53#_c_88_p N_A4_c_202_n 4.73027e-19 $X=2.575 $Y=2.495 $X2=0 $Y2=0
cc_95 N_A_102_53#_M1007_d N_A4_c_203_n 0.00631361f $X=2.095 $Y=1.835 $X2=0 $Y2=0
cc_96 N_A_102_53#_c_85_n N_A4_c_203_n 0.00479347f $X=1.757 $Y=1.96 $X2=0 $Y2=0
cc_97 N_A_102_53#_c_87_p N_A4_c_203_n 0.0151692f $X=2.197 $Y=2.14 $X2=0 $Y2=0
cc_98 N_A_102_53#_c_88_p N_A4_c_203_n 0.0165955f $X=2.575 $Y=2.495 $X2=0 $Y2=0
cc_99 N_A_102_53#_c_89_p N_A4_c_203_n 0.00157023f $X=2.405 $Y=2.33 $X2=0 $Y2=0
cc_100 N_A_102_53#_c_88_p N_A3_M1009_g 0.00111629f $X=2.575 $Y=2.495 $X2=0 $Y2=0
cc_101 N_A_102_53#_c_88_p N_A3_c_247_n 0.0393605f $X=2.575 $Y=2.495 $X2=0 $Y2=0
cc_102 N_A_102_53#_c_89_p N_A3_c_247_n 0.00478617f $X=2.405 $Y=2.33 $X2=0 $Y2=0
cc_103 N_A_102_53#_c_85_n N_VPWR_M1013_d 0.00290954f $X=1.757 $Y=1.96 $X2=0
+ $Y2=0
cc_104 N_A_102_53#_c_87_p N_VPWR_M1013_d 0.0068169f $X=2.197 $Y=2.14 $X2=0 $Y2=0
cc_105 N_A_102_53#_M1003_g N_VPWR_c_347_n 0.00731199f $X=0.585 $Y=2.465 $X2=0
+ $Y2=0
cc_106 N_A_102_53#_M1003_g N_VPWR_c_358_n 4.10802e-19 $X=0.585 $Y=2.465 $X2=0
+ $Y2=0
cc_107 N_A_102_53#_M1013_g N_VPWR_c_358_n 0.00723432f $X=1.015 $Y=2.465 $X2=0
+ $Y2=0
cc_108 N_A_102_53#_c_121_p N_VPWR_c_358_n 0.0289242f $X=1.62 $Y=1.51 $X2=0 $Y2=0
cc_109 N_A_102_53#_c_77_n N_VPWR_c_358_n 0.00816921f $X=1.495 $Y=1.51 $X2=0
+ $Y2=0
cc_110 N_A_102_53#_c_85_n N_VPWR_c_358_n 0.00920761f $X=1.757 $Y=1.96 $X2=0
+ $Y2=0
cc_111 N_A_102_53#_c_87_p N_VPWR_c_358_n 0.0153688f $X=2.197 $Y=2.14 $X2=0 $Y2=0
cc_112 N_A_102_53#_c_89_p N_VPWR_c_358_n 0.00472484f $X=2.405 $Y=2.33 $X2=0
+ $Y2=0
cc_113 N_A_102_53#_M1003_g N_VPWR_c_348_n 4.98916e-19 $X=0.585 $Y=2.465 $X2=0
+ $Y2=0
cc_114 N_A_102_53#_M1013_g N_VPWR_c_348_n 0.00986717f $X=1.015 $Y=2.465 $X2=0
+ $Y2=0
cc_115 N_A_102_53#_M1013_g N_VPWR_c_367_n 0.0055922f $X=1.015 $Y=2.465 $X2=0
+ $Y2=0
cc_116 N_A_102_53#_c_121_p N_VPWR_c_367_n 0.00495202f $X=1.62 $Y=1.51 $X2=0
+ $Y2=0
cc_117 N_A_102_53#_c_77_n N_VPWR_c_367_n 0.00286807f $X=1.495 $Y=1.51 $X2=0
+ $Y2=0
cc_118 N_A_102_53#_c_87_p N_VPWR_c_367_n 0.0218515f $X=2.197 $Y=2.14 $X2=0 $Y2=0
cc_119 N_A_102_53#_M1003_g N_VPWR_c_351_n 0.0054895f $X=0.585 $Y=2.465 $X2=0
+ $Y2=0
cc_120 N_A_102_53#_M1013_g N_VPWR_c_351_n 0.00486043f $X=1.015 $Y=2.465 $X2=0
+ $Y2=0
cc_121 N_A_102_53#_c_88_p N_VPWR_c_352_n 0.0428299f $X=2.575 $Y=2.495 $X2=0
+ $Y2=0
cc_122 N_A_102_53#_M1007_d N_VPWR_c_345_n 0.00505717f $X=2.095 $Y=1.835 $X2=0
+ $Y2=0
cc_123 N_A_102_53#_M1003_g N_VPWR_c_345_n 0.010787f $X=0.585 $Y=2.465 $X2=0
+ $Y2=0
cc_124 N_A_102_53#_M1013_g N_VPWR_c_345_n 0.00824727f $X=1.015 $Y=2.465 $X2=0
+ $Y2=0
cc_125 N_A_102_53#_c_88_p N_VPWR_c_345_n 0.0256043f $X=2.575 $Y=2.495 $X2=0
+ $Y2=0
cc_126 N_A_102_53#_c_74_n X 0.0160634f $X=0.585 $Y=1.345 $X2=0 $Y2=0
cc_127 N_A_102_53#_M1003_g X 0.0223641f $X=0.585 $Y=2.465 $X2=0 $Y2=0
cc_128 N_A_102_53#_c_75_n X 0.00369031f $X=1.015 $Y=1.345 $X2=0 $Y2=0
cc_129 N_A_102_53#_M1013_g X 0.00481266f $X=1.015 $Y=2.465 $X2=0 $Y2=0
cc_130 N_A_102_53#_c_76_n X 0.0307133f $X=1.09 $Y=1.51 $X2=0 $Y2=0
cc_131 N_A_102_53#_c_121_p X 0.0257389f $X=1.62 $Y=1.51 $X2=0 $Y2=0
cc_132 N_A_102_53#_c_74_n N_VGND_c_429_n 0.00712782f $X=0.585 $Y=1.345 $X2=0
+ $Y2=0
cc_133 N_A_102_53#_c_74_n N_VGND_c_430_n 6.4119e-19 $X=0.585 $Y=1.345 $X2=0
+ $Y2=0
cc_134 N_A_102_53#_c_75_n N_VGND_c_430_n 0.0168197f $X=1.015 $Y=1.345 $X2=0
+ $Y2=0
cc_135 N_A_102_53#_c_121_p N_VGND_c_430_n 0.0244507f $X=1.62 $Y=1.51 $X2=0 $Y2=0
cc_136 N_A_102_53#_c_77_n N_VGND_c_430_n 0.00688795f $X=1.495 $Y=1.51 $X2=0
+ $Y2=0
cc_137 N_A_102_53#_c_79_n N_VGND_c_430_n 0.0652063f $X=2.035 $Y=0.39 $X2=0 $Y2=0
cc_138 N_A_102_53#_c_79_n N_VGND_c_433_n 0.0389683f $X=2.035 $Y=0.39 $X2=0 $Y2=0
cc_139 N_A_102_53#_c_74_n N_VGND_c_437_n 0.00534051f $X=0.585 $Y=1.345 $X2=0
+ $Y2=0
cc_140 N_A_102_53#_c_75_n N_VGND_c_437_n 0.00465077f $X=1.015 $Y=1.345 $X2=0
+ $Y2=0
cc_141 N_A_102_53#_M1004_s N_VGND_c_439_n 0.00212301f $X=1.91 $Y=0.245 $X2=0
+ $Y2=0
cc_142 N_A_102_53#_c_74_n N_VGND_c_439_n 0.00537853f $X=0.585 $Y=1.345 $X2=0
+ $Y2=0
cc_143 N_A_102_53#_c_75_n N_VGND_c_439_n 0.00451796f $X=1.015 $Y=1.345 $X2=0
+ $Y2=0
cc_144 N_A_102_53#_c_79_n N_VGND_c_439_n 0.0222883f $X=2.035 $Y=0.39 $X2=0 $Y2=0
cc_145 N_A_102_53#_c_79_n N_A_465_49#_c_491_n 0.0477265f $X=2.035 $Y=0.39 $X2=0
+ $Y2=0
cc_146 N_A_102_53#_c_78_n N_A_465_49#_c_487_n 0.00520417f $X=1.757 $Y=1.345
+ $X2=0 $Y2=0
cc_147 N_A_102_53#_c_79_n N_A_465_49#_c_487_n 0.00242364f $X=2.035 $Y=0.39 $X2=0
+ $Y2=0
cc_148 N_B1_c_162_n N_A4_M1010_g 0.0199379f $X=2.25 $Y=1.21 $X2=0 $Y2=0
cc_149 B1 N_A4_M1010_g 7.16407e-19 $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_150 N_B1_M1007_g N_A4_M1008_g 0.00872161f $X=2.02 $Y=2.465 $X2=0 $Y2=0
cc_151 N_B1_M1007_g N_A4_c_202_n 0.00322065f $X=2.02 $Y=2.465 $X2=0 $Y2=0
cc_152 B1 N_A4_c_202_n 6.7325e-19 $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_153 N_B1_c_164_n N_A4_c_202_n 0.0123166f $X=2.25 $Y=1.375 $X2=0 $Y2=0
cc_154 N_B1_M1007_g N_A4_c_203_n 0.00249362f $X=2.02 $Y=2.465 $X2=0 $Y2=0
cc_155 B1 N_A4_c_203_n 0.0246118f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_156 N_B1_c_164_n N_A4_c_203_n 0.00129794f $X=2.25 $Y=1.375 $X2=0 $Y2=0
cc_157 N_B1_M1007_g N_VPWR_c_358_n 0.00335725f $X=2.02 $Y=2.465 $X2=0 $Y2=0
cc_158 N_B1_M1007_g N_VPWR_c_348_n 0.00656185f $X=2.02 $Y=2.465 $X2=0 $Y2=0
cc_159 N_B1_M1007_g N_VPWR_c_352_n 0.0054895f $X=2.02 $Y=2.465 $X2=0 $Y2=0
cc_160 N_B1_M1007_g N_VPWR_c_345_n 0.0117066f $X=2.02 $Y=2.465 $X2=0 $Y2=0
cc_161 N_B1_c_162_n N_VGND_c_433_n 0.00539298f $X=2.25 $Y=1.21 $X2=0 $Y2=0
cc_162 N_B1_c_162_n N_VGND_c_439_n 0.0113563f $X=2.25 $Y=1.21 $X2=0 $Y2=0
cc_163 N_B1_c_162_n N_A_465_49#_c_491_n 0.00320203f $X=2.25 $Y=1.21 $X2=0 $Y2=0
cc_164 N_B1_c_162_n N_A_465_49#_c_487_n 0.00182767f $X=2.25 $Y=1.21 $X2=0 $Y2=0
cc_165 N_A4_M1008_g N_A3_M1009_g 0.0564942f $X=2.79 $Y=2.465 $X2=0 $Y2=0
cc_166 N_A4_M1010_g N_A3_M1006_g 0.0176694f $X=2.725 $Y=0.665 $X2=0 $Y2=0
cc_167 N_A4_c_202_n N_A3_c_246_n 0.0564942f $X=2.7 $Y=1.51 $X2=0 $Y2=0
cc_168 N_A4_c_203_n N_A3_c_246_n 7.90116e-19 $X=2.7 $Y=1.51 $X2=0 $Y2=0
cc_169 N_A4_c_202_n N_A3_c_247_n 0.011166f $X=2.7 $Y=1.51 $X2=0 $Y2=0
cc_170 N_A4_c_203_n N_A3_c_247_n 0.0639731f $X=2.7 $Y=1.51 $X2=0 $Y2=0
cc_171 N_A4_M1008_g N_VPWR_c_352_n 0.0054895f $X=2.79 $Y=2.465 $X2=0 $Y2=0
cc_172 N_A4_M1008_g N_VPWR_c_345_n 0.0104939f $X=2.79 $Y=2.465 $X2=0 $Y2=0
cc_173 N_A4_M1010_g N_VGND_c_431_n 0.00311747f $X=2.725 $Y=0.665 $X2=0 $Y2=0
cc_174 N_A4_M1010_g N_VGND_c_433_n 0.00561712f $X=2.725 $Y=0.665 $X2=0 $Y2=0
cc_175 N_A4_M1010_g N_VGND_c_439_n 0.0106814f $X=2.725 $Y=0.665 $X2=0 $Y2=0
cc_176 N_A4_M1010_g N_A_465_49#_c_491_n 0.00998098f $X=2.725 $Y=0.665 $X2=0
+ $Y2=0
cc_177 N_A4_M1010_g N_A_465_49#_c_486_n 0.012748f $X=2.725 $Y=0.665 $X2=0 $Y2=0
cc_178 N_A4_c_202_n N_A_465_49#_c_486_n 0.00221419f $X=2.7 $Y=1.51 $X2=0 $Y2=0
cc_179 N_A4_c_203_n N_A_465_49#_c_486_n 0.0117493f $X=2.7 $Y=1.51 $X2=0 $Y2=0
cc_180 N_A4_M1010_g N_A_465_49#_c_487_n 0.0011945f $X=2.725 $Y=0.665 $X2=0 $Y2=0
cc_181 N_A4_c_202_n N_A_465_49#_c_487_n 9.10195e-19 $X=2.7 $Y=1.51 $X2=0 $Y2=0
cc_182 N_A4_c_203_n N_A_465_49#_c_487_n 0.0147535f $X=2.7 $Y=1.51 $X2=0 $Y2=0
cc_183 N_A4_M1010_g N_A_465_49#_c_503_n 3.78115e-19 $X=2.725 $Y=0.665 $X2=0
+ $Y2=0
cc_184 N_A3_M1006_g N_A2_M1012_g 0.0250312f $X=3.26 $Y=0.665 $X2=0 $Y2=0
cc_185 N_A3_M1009_g N_A2_M1001_g 0.0463739f $X=3.15 $Y=2.465 $X2=0 $Y2=0
cc_186 N_A3_c_247_n N_A2_M1001_g 0.00372779f $X=3.24 $Y=1.51 $X2=0 $Y2=0
cc_187 N_A3_c_246_n N_A2_c_285_n 0.0204266f $X=3.24 $Y=1.51 $X2=0 $Y2=0
cc_188 N_A3_c_247_n N_A2_c_285_n 2.88166e-19 $X=3.24 $Y=1.51 $X2=0 $Y2=0
cc_189 N_A3_M1009_g N_A2_c_286_n 0.00437184f $X=3.15 $Y=2.465 $X2=0 $Y2=0
cc_190 N_A3_c_246_n N_A2_c_286_n 0.00236569f $X=3.24 $Y=1.51 $X2=0 $Y2=0
cc_191 N_A3_c_247_n N_A2_c_286_n 0.137865f $X=3.24 $Y=1.51 $X2=0 $Y2=0
cc_192 N_A3_M1009_g N_VPWR_c_352_n 0.0037962f $X=3.15 $Y=2.465 $X2=0 $Y2=0
cc_193 N_A3_c_247_n N_VPWR_c_352_n 0.0113755f $X=3.24 $Y=1.51 $X2=0 $Y2=0
cc_194 N_A3_M1009_g N_VPWR_c_345_n 0.00561463f $X=3.15 $Y=2.465 $X2=0 $Y2=0
cc_195 N_A3_c_247_n N_VPWR_c_345_n 0.0116419f $X=3.24 $Y=1.51 $X2=0 $Y2=0
cc_196 N_A3_c_247_n A_573_367# 0.0118132f $X=3.24 $Y=1.51 $X2=-0.19 $Y2=-0.245
cc_197 N_A3_c_247_n A_645_367# 0.0106255f $X=3.24 $Y=1.51 $X2=-0.19 $Y2=-0.245
cc_198 N_A3_M1006_g N_VGND_c_431_n 0.00177287f $X=3.26 $Y=0.665 $X2=0 $Y2=0
cc_199 N_A3_M1006_g N_VGND_c_435_n 0.00569184f $X=3.26 $Y=0.665 $X2=0 $Y2=0
cc_200 N_A3_M1006_g N_VGND_c_439_n 0.0107208f $X=3.26 $Y=0.665 $X2=0 $Y2=0
cc_201 N_A3_M1006_g N_A_465_49#_c_491_n 3.83578e-19 $X=3.26 $Y=0.665 $X2=0 $Y2=0
cc_202 N_A3_M1006_g N_A_465_49#_c_486_n 0.0132571f $X=3.26 $Y=0.665 $X2=0 $Y2=0
cc_203 N_A3_c_246_n N_A_465_49#_c_486_n 7.65086e-19 $X=3.24 $Y=1.51 $X2=0 $Y2=0
cc_204 N_A3_c_247_n N_A_465_49#_c_486_n 0.0268961f $X=3.24 $Y=1.51 $X2=0 $Y2=0
cc_205 N_A3_M1006_g N_A_465_49#_c_503_n 0.00986364f $X=3.26 $Y=0.665 $X2=0 $Y2=0
cc_206 N_A3_M1006_g N_A_465_49#_c_490_n 0.0013549f $X=3.26 $Y=0.665 $X2=0 $Y2=0
cc_207 N_A3_c_246_n N_A_465_49#_c_490_n 0.00311089f $X=3.24 $Y=1.51 $X2=0 $Y2=0
cc_208 N_A2_M1012_g N_A1_M1002_g 0.0253902f $X=3.69 $Y=0.665 $X2=0 $Y2=0
cc_209 N_A2_M1001_g N_A1_M1005_g 0.0458281f $X=3.69 $Y=2.465 $X2=0 $Y2=0
cc_210 N_A2_c_286_n N_A1_M1005_g 0.0403697f $X=3.78 $Y=1.51 $X2=0 $Y2=0
cc_211 N_A2_c_285_n N_A1_c_322_n 0.0214098f $X=3.78 $Y=1.51 $X2=0 $Y2=0
cc_212 N_A2_c_286_n N_A1_c_322_n 0.00740406f $X=3.78 $Y=1.51 $X2=0 $Y2=0
cc_213 N_A2_c_286_n N_A1_c_323_n 0.032637f $X=3.78 $Y=1.51 $X2=0 $Y2=0
cc_214 N_A2_M1001_g N_VPWR_c_352_n 0.0037962f $X=3.69 $Y=2.465 $X2=0 $Y2=0
cc_215 N_A2_c_286_n N_VPWR_c_352_n 0.0241565f $X=3.78 $Y=1.51 $X2=0 $Y2=0
cc_216 N_A2_M1001_g N_VPWR_c_345_n 0.00607065f $X=3.69 $Y=2.465 $X2=0 $Y2=0
cc_217 N_A2_c_286_n N_VPWR_c_345_n 0.023993f $X=3.78 $Y=1.51 $X2=0 $Y2=0
cc_218 N_A2_c_286_n A_645_367# 0.0110038f $X=3.78 $Y=1.51 $X2=-0.19 $Y2=-0.245
cc_219 N_A2_c_286_n A_753_367# 0.00520986f $X=3.78 $Y=1.51 $X2=-0.19 $Y2=-0.245
cc_220 N_A2_M1012_g N_VGND_c_432_n 0.00517281f $X=3.69 $Y=0.665 $X2=0 $Y2=0
cc_221 N_A2_M1012_g N_VGND_c_435_n 0.00554241f $X=3.69 $Y=0.665 $X2=0 $Y2=0
cc_222 N_A2_M1012_g N_VGND_c_439_n 0.0104609f $X=3.69 $Y=0.665 $X2=0 $Y2=0
cc_223 N_A2_M1012_g N_A_465_49#_c_503_n 0.0104977f $X=3.69 $Y=0.665 $X2=0 $Y2=0
cc_224 N_A2_M1012_g N_A_465_49#_c_488_n 0.0124019f $X=3.69 $Y=0.665 $X2=0 $Y2=0
cc_225 N_A2_c_285_n N_A_465_49#_c_488_n 0.00126891f $X=3.78 $Y=1.51 $X2=0 $Y2=0
cc_226 N_A2_c_286_n N_A_465_49#_c_488_n 0.0438185f $X=3.78 $Y=1.51 $X2=0 $Y2=0
cc_227 N_A2_M1012_g N_A_465_49#_c_489_n 6.32452e-19 $X=3.69 $Y=0.665 $X2=0 $Y2=0
cc_228 N_A2_M1012_g N_A_465_49#_c_490_n 0.00148772f $X=3.69 $Y=0.665 $X2=0 $Y2=0
cc_229 N_A2_c_286_n N_A_465_49#_c_490_n 0.0124198f $X=3.78 $Y=1.51 $X2=0 $Y2=0
cc_230 N_A1_M1005_g N_VPWR_c_350_n 0.00620143f $X=4.23 $Y=2.465 $X2=0 $Y2=0
cc_231 N_A1_c_322_n N_VPWR_c_350_n 0.00152187f $X=4.51 $Y=1.46 $X2=0 $Y2=0
cc_232 N_A1_c_323_n N_VPWR_c_350_n 0.0225603f $X=4.51 $Y=1.46 $X2=0 $Y2=0
cc_233 N_A1_M1005_g N_VPWR_c_352_n 0.00559321f $X=4.23 $Y=2.465 $X2=0 $Y2=0
cc_234 N_A1_M1005_g N_VPWR_c_345_n 0.0113162f $X=4.23 $Y=2.465 $X2=0 $Y2=0
cc_235 N_A1_M1002_g N_VGND_c_432_n 0.00315548f $X=4.23 $Y=0.665 $X2=0 $Y2=0
cc_236 N_A1_M1002_g N_VGND_c_438_n 0.00569184f $X=4.23 $Y=0.665 $X2=0 $Y2=0
cc_237 N_A1_M1002_g N_VGND_c_439_n 0.0117163f $X=4.23 $Y=0.665 $X2=0 $Y2=0
cc_238 N_A1_M1002_g N_A_465_49#_c_503_n 3.83715e-19 $X=4.23 $Y=0.665 $X2=0 $Y2=0
cc_239 N_A1_M1002_g N_A_465_49#_c_488_n 0.0190919f $X=4.23 $Y=0.665 $X2=0 $Y2=0
cc_240 N_A1_c_322_n N_A_465_49#_c_488_n 0.00845246f $X=4.51 $Y=1.46 $X2=0 $Y2=0
cc_241 N_A1_c_323_n N_A_465_49#_c_488_n 0.0226879f $X=4.51 $Y=1.46 $X2=0 $Y2=0
cc_242 N_A1_M1002_g N_A_465_49#_c_489_n 0.0109799f $X=4.23 $Y=0.665 $X2=0 $Y2=0
cc_243 N_VPWR_c_345_n N_X_M1003_s 0.00380103f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_244 N_VPWR_c_347_n X 0.0463448f $X=0.37 $Y=1.98 $X2=0 $Y2=0
cc_245 N_VPWR_c_351_n X 0.015688f $X=1.065 $Y=3.33 $X2=0 $Y2=0
cc_246 N_VPWR_c_345_n X 0.00984745f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_247 N_VPWR_c_345_n A_573_367# 0.00593643f $X=4.56 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_248 N_VPWR_c_345_n A_645_367# 0.00922383f $X=4.56 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_249 N_VPWR_c_345_n A_753_367# 0.00331457f $X=4.56 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_250 N_VPWR_c_347_n N_VGND_c_429_n 0.0105123f $X=0.37 $Y=1.98 $X2=0 $Y2=0
cc_251 X N_VGND_c_429_n 0.0333602f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_252 X N_VGND_c_430_n 0.0307804f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_253 X N_VGND_c_437_n 0.0103916f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_254 X N_VGND_c_439_n 0.0093632f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_255 N_VGND_c_439_n N_A_465_49#_M1004_d 0.00607622f $X=4.56 $Y=0 $X2=-0.19
+ $Y2=-0.245
cc_256 N_VGND_c_439_n N_A_465_49#_M1006_d 0.00223559f $X=4.56 $Y=0 $X2=0 $Y2=0
cc_257 N_VGND_c_439_n N_A_465_49#_M1002_d 0.00212301f $X=4.56 $Y=0 $X2=0 $Y2=0
cc_258 N_VGND_c_433_n N_A_465_49#_c_491_n 0.0143455f $X=2.83 $Y=0 $X2=0 $Y2=0
cc_259 N_VGND_c_439_n N_A_465_49#_c_491_n 0.00894414f $X=4.56 $Y=0 $X2=0 $Y2=0
cc_260 N_VGND_M1010_d N_A_465_49#_c_486_n 0.0029901f $X=2.8 $Y=0.245 $X2=0 $Y2=0
cc_261 N_VGND_c_431_n N_A_465_49#_c_486_n 0.0220482f $X=2.995 $Y=0.37 $X2=0
+ $Y2=0
cc_262 N_VGND_c_435_n N_A_465_49#_c_503_n 0.0168785f $X=3.8 $Y=0 $X2=0 $Y2=0
cc_263 N_VGND_c_439_n N_A_465_49#_c_503_n 0.0113568f $X=4.56 $Y=0 $X2=0 $Y2=0
cc_264 N_VGND_M1012_d N_A_465_49#_c_488_n 0.00306511f $X=3.765 $Y=0.245 $X2=0
+ $Y2=0
cc_265 N_VGND_c_432_n N_A_465_49#_c_488_n 0.022455f $X=3.965 $Y=0.37 $X2=0 $Y2=0
cc_266 N_VGND_c_438_n N_A_465_49#_c_489_n 0.0196832f $X=4.56 $Y=0 $X2=0 $Y2=0
cc_267 N_VGND_c_439_n N_A_465_49#_c_489_n 0.0118828f $X=4.56 $Y=0 $X2=0 $Y2=0
