# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__bufbuf_8
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__bufbuf_8 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.200000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.650000 1.405000 7.115000 1.755000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  2.352000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.055000 3.665000 1.225000 ;
        RECT 0.085000 1.225000 0.405000 1.755000 ;
        RECT 0.085000 1.755000 3.665000 1.925000 ;
        RECT 0.860000 1.925000 1.120000 3.075000 ;
        RECT 0.895000 0.290000 1.085000 1.055000 ;
        RECT 1.720000 1.925000 1.980000 3.075000 ;
        RECT 1.755000 0.290000 1.945000 1.055000 ;
        RECT 2.580000 1.925000 2.840000 3.075000 ;
        RECT 2.615000 0.290000 2.805000 1.055000 ;
        RECT 3.440000 1.925000 3.665000 3.075000 ;
        RECT 3.475000 0.290000 3.665000 1.055000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 7.200000 0.085000 ;
        RECT 0.395000  0.085000 0.725000 0.885000 ;
        RECT 1.255000  0.085000 1.585000 0.885000 ;
        RECT 2.115000  0.085000 2.445000 0.885000 ;
        RECT 2.975000  0.085000 3.305000 0.885000 ;
        RECT 3.835000  0.085000 4.190000 0.885000 ;
        RECT 4.740000  0.085000 5.070000 0.885000 ;
        RECT 6.210000  0.085000 6.540000 0.895000 ;
      LAYER mcon ;
        RECT 0.155000 -0.085000 0.325000 0.085000 ;
        RECT 0.635000 -0.085000 0.805000 0.085000 ;
        RECT 1.115000 -0.085000 1.285000 0.085000 ;
        RECT 1.595000 -0.085000 1.765000 0.085000 ;
        RECT 2.075000 -0.085000 2.245000 0.085000 ;
        RECT 2.555000 -0.085000 2.725000 0.085000 ;
        RECT 3.035000 -0.085000 3.205000 0.085000 ;
        RECT 3.515000 -0.085000 3.685000 0.085000 ;
        RECT 3.995000 -0.085000 4.165000 0.085000 ;
        RECT 4.475000 -0.085000 4.645000 0.085000 ;
        RECT 4.955000 -0.085000 5.125000 0.085000 ;
        RECT 5.435000 -0.085000 5.605000 0.085000 ;
        RECT 5.915000 -0.085000 6.085000 0.085000 ;
        RECT 6.395000 -0.085000 6.565000 0.085000 ;
        RECT 6.875000 -0.085000 7.045000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 7.200000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.245000 7.200000 3.415000 ;
        RECT 0.395000 2.105000 0.690000 3.245000 ;
        RECT 1.290000 2.105000 1.550000 3.245000 ;
        RECT 2.150000 2.105000 2.410000 3.245000 ;
        RECT 3.010000 2.105000 3.270000 3.245000 ;
        RECT 3.835000 2.095000 4.165000 3.245000 ;
        RECT 4.780000 2.095000 5.040000 3.245000 ;
        RECT 6.250000 2.370000 6.580000 3.245000 ;
      LAYER mcon ;
        RECT 0.155000 3.245000 0.325000 3.415000 ;
        RECT 0.635000 3.245000 0.805000 3.415000 ;
        RECT 1.115000 3.245000 1.285000 3.415000 ;
        RECT 1.595000 3.245000 1.765000 3.415000 ;
        RECT 2.075000 3.245000 2.245000 3.415000 ;
        RECT 2.555000 3.245000 2.725000 3.415000 ;
        RECT 3.035000 3.245000 3.205000 3.415000 ;
        RECT 3.515000 3.245000 3.685000 3.415000 ;
        RECT 3.995000 3.245000 4.165000 3.415000 ;
        RECT 4.475000 3.245000 4.645000 3.415000 ;
        RECT 4.955000 3.245000 5.125000 3.415000 ;
        RECT 5.435000 3.245000 5.605000 3.415000 ;
        RECT 5.915000 3.245000 6.085000 3.415000 ;
        RECT 6.395000 3.245000 6.565000 3.415000 ;
        RECT 6.875000 3.245000 7.045000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 7.200000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.585000 1.395000 4.005000 1.585000 ;
      RECT 3.835000 1.055000 5.500000 1.225000 ;
      RECT 3.835000 1.225000 4.005000 1.395000 ;
      RECT 3.835000 1.585000 4.005000 1.755000 ;
      RECT 3.835000 1.755000 5.500000 1.925000 ;
      RECT 4.185000 1.395000 6.020000 1.585000 ;
      RECT 4.335000 1.925000 4.610000 3.075000 ;
      RECT 4.360000 0.290000 4.570000 1.055000 ;
      RECT 5.210000 1.925000 5.500000 3.075000 ;
      RECT 5.240000 0.290000 5.500000 1.055000 ;
      RECT 5.760000 0.435000 6.020000 1.395000 ;
      RECT 5.840000 1.585000 6.020000 1.815000 ;
      RECT 5.840000 1.815000 6.070000 2.825000 ;
      RECT 6.190000 1.065000 7.105000 1.235000 ;
      RECT 6.190000 1.235000 6.440000 1.525000 ;
      RECT 6.240000 1.525000 6.440000 1.925000 ;
      RECT 6.240000 1.925000 7.105000 2.200000 ;
      RECT 6.775000 0.665000 7.105000 1.065000 ;
  END
END sky130_fd_sc_lp__bufbuf_8
