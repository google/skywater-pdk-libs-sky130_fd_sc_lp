* File: sky130_fd_sc_lp__o2bb2ai_lp.pxi.spice
* Created: Fri Aug 28 11:13:06 2020
* 
x_PM_SKY130_FD_SC_LP__O2BB2AI_LP%A1_N N_A1_N_M1001_g N_A1_N_M1006_g A1_N A1_N
+ N_A1_N_c_67_n PM_SKY130_FD_SC_LP__O2BB2AI_LP%A1_N
x_PM_SKY130_FD_SC_LP__O2BB2AI_LP%A2_N N_A2_N_M1009_g N_A2_N_c_97_n
+ N_A2_N_M1005_g N_A2_N_c_99_n A2_N N_A2_N_c_101_n
+ PM_SKY130_FD_SC_LP__O2BB2AI_LP%A2_N
x_PM_SKY130_FD_SC_LP__O2BB2AI_LP%A_145_419# N_A_145_419#_M1009_d
+ N_A_145_419#_M1006_d N_A_145_419#_M1002_g N_A_145_419#_c_148_n
+ N_A_145_419#_c_149_n N_A_145_419#_M1007_g N_A_145_419#_c_150_n
+ N_A_145_419#_c_151_n N_A_145_419#_c_152_n N_A_145_419#_c_165_n
+ N_A_145_419#_c_157_n N_A_145_419#_c_158_n N_A_145_419#_c_153_n
+ N_A_145_419#_c_154_n PM_SKY130_FD_SC_LP__O2BB2AI_LP%A_145_419#
x_PM_SKY130_FD_SC_LP__O2BB2AI_LP%B2 N_B2_M1008_g N_B2_M1003_g B2 B2 N_B2_c_230_n
+ PM_SKY130_FD_SC_LP__O2BB2AI_LP%B2
x_PM_SKY130_FD_SC_LP__O2BB2AI_LP%B1 N_B1_c_269_n N_B1_M1004_g N_B1_M1000_g
+ N_B1_c_270_n B1 B1 N_B1_c_268_n PM_SKY130_FD_SC_LP__O2BB2AI_LP%B1
x_PM_SKY130_FD_SC_LP__O2BB2AI_LP%VPWR N_VPWR_M1006_s N_VPWR_M1005_d
+ N_VPWR_M1004_d N_VPWR_c_295_n N_VPWR_c_296_n N_VPWR_c_297_n N_VPWR_c_298_n
+ N_VPWR_c_299_n N_VPWR_c_300_n N_VPWR_c_301_n VPWR N_VPWR_c_302_n
+ N_VPWR_c_294_n PM_SKY130_FD_SC_LP__O2BB2AI_LP%VPWR
x_PM_SKY130_FD_SC_LP__O2BB2AI_LP%Y N_Y_M1007_s N_Y_M1002_d N_Y_c_342_n
+ N_Y_c_338_n N_Y_c_339_n Y Y PM_SKY130_FD_SC_LP__O2BB2AI_LP%Y
x_PM_SKY130_FD_SC_LP__O2BB2AI_LP%VGND N_VGND_M1001_s N_VGND_M1003_d
+ N_VGND_c_380_n N_VGND_c_381_n N_VGND_c_382_n VGND N_VGND_c_383_n
+ N_VGND_c_384_n N_VGND_c_385_n N_VGND_c_386_n
+ PM_SKY130_FD_SC_LP__O2BB2AI_LP%VGND
x_PM_SKY130_FD_SC_LP__O2BB2AI_LP%A_400_83# N_A_400_83#_M1007_d
+ N_A_400_83#_M1000_d N_A_400_83#_c_422_n N_A_400_83#_c_418_n
+ N_A_400_83#_c_419_n N_A_400_83#_c_420_n
+ PM_SKY130_FD_SC_LP__O2BB2AI_LP%A_400_83#
cc_1 VNB N_A1_N_M1001_g 0.054249f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.495
cc_2 VNB A1_N 0.0221065f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_3 VNB N_A1_N_c_67_n 0.0532678f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.39
cc_4 VNB N_A2_N_M1009_g 0.0208099f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.495
cc_5 VNB N_A2_N_c_97_n 0.0140219f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=1.895
cc_6 VNB N_A2_N_M1005_g 0.00530684f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=2.595
cc_7 VNB N_A2_N_c_99_n 0.0296754f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB A2_N 0.00671148f $X=-0.19 $Y=-0.245 $X2=0.472 $Y2=1.39
cc_9 VNB N_A2_N_c_101_n 0.0318923f $X=-0.19 $Y=-0.245 $X2=0.472 $Y2=1.225
cc_10 VNB N_A_145_419#_c_148_n 0.0306721f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_145_419#_c_149_n 0.0165068f $X=-0.19 $Y=-0.245 $X2=0.472 $Y2=1.39
cc_12 VNB N_A_145_419#_c_150_n 0.0138852f $X=-0.19 $Y=-0.245 $X2=0.307 $Y2=1.295
cc_13 VNB N_A_145_419#_c_151_n 0.0103477f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_145_419#_c_152_n 0.00880095f $X=-0.19 $Y=-0.245 $X2=0.307 $Y2=1.39
cc_15 VNB N_A_145_419#_c_153_n 0.0034216f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_145_419#_c_154_n 0.0115749f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_B2_M1003_g 0.0379523f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=2.595
cc_18 VNB B2 0.00739033f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_19 VNB N_B2_c_230_n 0.0220053f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.39
cc_20 VNB N_B1_M1000_g 0.05143f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=2.595
cc_21 VNB B1 0.0246527f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_B1_c_268_n 0.0302061f $X=-0.19 $Y=-0.245 $X2=0.472 $Y2=1.225
cc_23 VNB N_VPWR_c_294_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_Y_c_338_n 0.00833442f $X=-0.19 $Y=-0.245 $X2=0.472 $Y2=1.225
cc_25 VNB N_Y_c_339_n 0.00397852f $X=-0.19 $Y=-0.245 $X2=0.307 $Y2=1.295
cc_26 VNB Y 0.0121765f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_380_n 0.0113827f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=2.595
cc_28 VNB N_VGND_c_381_n 0.0259837f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_29 VNB N_VGND_c_382_n 0.00998722f $X=-0.19 $Y=-0.245 $X2=0.472 $Y2=1.39
cc_30 VNB N_VGND_c_383_n 0.0537597f $X=-0.19 $Y=-0.245 $X2=0.472 $Y2=1.895
cc_31 VNB N_VGND_c_384_n 0.0202312f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_385_n 0.226555f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_386_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_400_83#_c_418_n 0.0175826f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_400_83#_c_419_n 0.00620038f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_400_83#_c_420_n 0.0150847f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.39
cc_37 VPB N_A1_N_M1006_g 0.0346523f $X=-0.19 $Y=1.655 $X2=0.6 $Y2=2.595
cc_38 VPB A1_N 0.0134933f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_39 VPB N_A1_N_c_67_n 0.0301782f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.39
cc_40 VPB N_A2_N_M1005_g 0.0419864f $X=-0.19 $Y=1.655 $X2=0.6 $Y2=2.595
cc_41 VPB N_A_145_419#_M1002_g 0.0272675f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_42 VPB N_A_145_419#_c_152_n 5.3438e-19 $X=-0.19 $Y=1.655 $X2=0.307 $Y2=1.39
cc_43 VPB N_A_145_419#_c_157_n 0.00930583f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_44 VPB N_A_145_419#_c_158_n 0.00555217f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_45 VPB N_A_145_419#_c_153_n 0.00464013f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_46 VPB N_A_145_419#_c_154_n 0.0265227f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_47 VPB N_B2_M1008_g 0.038894f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=0.495
cc_48 VPB B2 0.0108484f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_49 VPB N_B2_c_230_n 0.00680067f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.39
cc_50 VPB N_B1_c_269_n 0.0303743f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=1.225
cc_51 VPB N_B1_c_270_n 0.0205845f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_52 VPB B1 0.00818035f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_53 VPB N_B1_c_268_n 0.0120326f $X=-0.19 $Y=1.655 $X2=0.472 $Y2=1.225
cc_54 VPB N_VPWR_c_295_n 0.0124723f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_55 VPB N_VPWR_c_296_n 0.0436343f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_56 VPB N_VPWR_c_297_n 0.00284591f $X=-0.19 $Y=1.655 $X2=0.307 $Y2=1.295
cc_57 VPB N_VPWR_c_298_n 0.0109777f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_58 VPB N_VPWR_c_299_n 0.045048f $X=-0.19 $Y=1.655 $X2=0.307 $Y2=1.665
cc_59 VPB N_VPWR_c_300_n 0.0180883f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_60 VPB N_VPWR_c_301_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_61 VPB N_VPWR_c_302_n 0.0389824f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_62 VPB N_VPWR_c_294_n 0.0469817f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_63 VPB N_Y_c_339_n 0.00826014f $X=-0.19 $Y=1.655 $X2=0.307 $Y2=1.295
cc_64 N_A1_N_M1001_g N_A2_N_M1009_g 0.041651f $X=0.495 $Y=0.495 $X2=0 $Y2=0
cc_65 A1_N N_A2_N_M1005_g 2.16378e-19 $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_66 N_A1_N_c_67_n N_A2_N_M1005_g 0.0419994f $X=0.385 $Y=1.39 $X2=0 $Y2=0
cc_67 N_A1_N_c_67_n A2_N 3.27285e-19 $X=0.385 $Y=1.39 $X2=0 $Y2=0
cc_68 N_A1_N_M1001_g N_A2_N_c_101_n 0.00540337f $X=0.495 $Y=0.495 $X2=0 $Y2=0
cc_69 N_A1_N_c_67_n N_A2_N_c_101_n 0.0183313f $X=0.385 $Y=1.39 $X2=0 $Y2=0
cc_70 N_A1_N_M1001_g N_A_145_419#_c_151_n 0.0021305f $X=0.495 $Y=0.495 $X2=0
+ $Y2=0
cc_71 N_A1_N_M1001_g N_A_145_419#_c_152_n 0.0110804f $X=0.495 $Y=0.495 $X2=0
+ $Y2=0
cc_72 A1_N N_A_145_419#_c_152_n 0.0407075f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_73 N_A1_N_c_67_n N_A_145_419#_c_152_n 0.0150765f $X=0.385 $Y=1.39 $X2=0 $Y2=0
cc_74 N_A1_N_M1006_g N_A_145_419#_c_165_n 0.0315103f $X=0.6 $Y=2.595 $X2=0 $Y2=0
cc_75 N_A1_N_M1006_g N_A_145_419#_c_158_n 0.00244432f $X=0.6 $Y=2.595 $X2=0
+ $Y2=0
cc_76 A1_N N_A_145_419#_c_158_n 0.00998235f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_77 N_A1_N_c_67_n N_A_145_419#_c_158_n 0.00416038f $X=0.385 $Y=1.39 $X2=0
+ $Y2=0
cc_78 N_A1_N_M1006_g N_VPWR_c_296_n 0.0218955f $X=0.6 $Y=2.595 $X2=0 $Y2=0
cc_79 A1_N N_VPWR_c_296_n 0.0283096f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_80 N_A1_N_c_67_n N_VPWR_c_296_n 0.00198162f $X=0.385 $Y=1.39 $X2=0 $Y2=0
cc_81 N_A1_N_M1006_g N_VPWR_c_297_n 0.00127185f $X=0.6 $Y=2.595 $X2=0 $Y2=0
cc_82 N_A1_N_M1006_g N_VPWR_c_300_n 0.00834099f $X=0.6 $Y=2.595 $X2=0 $Y2=0
cc_83 N_A1_N_M1006_g N_VPWR_c_294_n 0.0131096f $X=0.6 $Y=2.595 $X2=0 $Y2=0
cc_84 N_A1_N_M1001_g N_VGND_c_381_n 0.0137106f $X=0.495 $Y=0.495 $X2=0 $Y2=0
cc_85 A1_N N_VGND_c_381_n 0.0148402f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_86 N_A1_N_c_67_n N_VGND_c_381_n 0.00126057f $X=0.385 $Y=1.39 $X2=0 $Y2=0
cc_87 N_A1_N_M1001_g N_VGND_c_383_n 0.00445056f $X=0.495 $Y=0.495 $X2=0 $Y2=0
cc_88 N_A1_N_M1001_g N_VGND_c_385_n 0.00804604f $X=0.495 $Y=0.495 $X2=0 $Y2=0
cc_89 N_A2_N_M1005_g N_A_145_419#_M1002_g 0.0229058f $X=1.13 $Y=2.595 $X2=0
+ $Y2=0
cc_90 N_A2_N_M1005_g N_A_145_419#_c_148_n 7.36371e-19 $X=1.13 $Y=2.595 $X2=0
+ $Y2=0
cc_91 A2_N N_A_145_419#_c_148_n 0.00160572f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_92 N_A2_N_c_101_n N_A_145_419#_c_148_n 0.00696522f $X=1.13 $Y=1.07 $X2=0
+ $Y2=0
cc_93 N_A2_N_c_99_n N_A_145_419#_c_149_n 0.00118305f $X=1.052 $Y=0.985 $X2=0
+ $Y2=0
cc_94 N_A2_N_c_99_n N_A_145_419#_c_150_n 0.00696522f $X=1.052 $Y=0.985 $X2=0
+ $Y2=0
cc_95 A2_N N_A_145_419#_c_150_n 8.87685e-19 $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_96 N_A2_N_M1009_g N_A_145_419#_c_151_n 0.0172334f $X=0.885 $Y=0.495 $X2=0
+ $Y2=0
cc_97 N_A2_N_c_99_n N_A_145_419#_c_151_n 0.0100379f $X=1.052 $Y=0.985 $X2=0
+ $Y2=0
cc_98 A2_N N_A_145_419#_c_151_n 0.0201712f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_99 N_A2_N_M1009_g N_A_145_419#_c_152_n 0.00320595f $X=0.885 $Y=0.495 $X2=0
+ $Y2=0
cc_100 N_A2_N_M1005_g N_A_145_419#_c_152_n 0.00183545f $X=1.13 $Y=2.595 $X2=0
+ $Y2=0
cc_101 N_A2_N_c_99_n N_A_145_419#_c_152_n 0.00611612f $X=1.052 $Y=0.985 $X2=0
+ $Y2=0
cc_102 A2_N N_A_145_419#_c_152_n 0.047533f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_103 N_A2_N_c_101_n N_A_145_419#_c_152_n 0.00423807f $X=1.13 $Y=1.07 $X2=0
+ $Y2=0
cc_104 N_A2_N_M1005_g N_A_145_419#_c_165_n 0.0255632f $X=1.13 $Y=2.595 $X2=0
+ $Y2=0
cc_105 N_A2_N_c_97_n N_A_145_419#_c_157_n 0.00103948f $X=1.13 $Y=1.575 $X2=0
+ $Y2=0
cc_106 N_A2_N_M1005_g N_A_145_419#_c_157_n 0.0177643f $X=1.13 $Y=2.595 $X2=0
+ $Y2=0
cc_107 A2_N N_A_145_419#_c_157_n 0.0200251f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_108 N_A2_N_c_97_n N_A_145_419#_c_158_n 0.0018941f $X=1.13 $Y=1.575 $X2=0
+ $Y2=0
cc_109 N_A2_N_M1005_g N_A_145_419#_c_158_n 0.00333192f $X=1.13 $Y=2.595 $X2=0
+ $Y2=0
cc_110 A2_N N_A_145_419#_c_158_n 7.69221e-19 $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_111 N_A2_N_M1005_g N_A_145_419#_c_153_n 9.37255e-19 $X=1.13 $Y=2.595 $X2=0
+ $Y2=0
cc_112 N_A2_N_M1005_g N_A_145_419#_c_154_n 0.017597f $X=1.13 $Y=2.595 $X2=0
+ $Y2=0
cc_113 N_A2_N_M1005_g N_VPWR_c_296_n 0.00124014f $X=1.13 $Y=2.595 $X2=0 $Y2=0
cc_114 N_A2_N_M1005_g N_VPWR_c_297_n 0.0257535f $X=1.13 $Y=2.595 $X2=0 $Y2=0
cc_115 N_A2_N_M1005_g N_VPWR_c_300_n 0.00840199f $X=1.13 $Y=2.595 $X2=0 $Y2=0
cc_116 N_A2_N_M1005_g N_VPWR_c_294_n 0.0136033f $X=1.13 $Y=2.595 $X2=0 $Y2=0
cc_117 N_A2_N_M1005_g N_Y_c_342_n 3.87543e-19 $X=1.13 $Y=2.595 $X2=0 $Y2=0
cc_118 A2_N N_Y_c_338_n 0.011762f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_119 N_A2_N_c_101_n N_Y_c_338_n 7.3054e-19 $X=1.13 $Y=1.07 $X2=0 $Y2=0
cc_120 A2_N N_Y_c_339_n 0.00477482f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_121 N_A2_N_M1009_g Y 0.00334007f $X=0.885 $Y=0.495 $X2=0 $Y2=0
cc_122 N_A2_N_c_99_n Y 0.00318923f $X=1.052 $Y=0.985 $X2=0 $Y2=0
cc_123 A2_N Y 0.023407f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_124 N_A2_N_M1009_g N_VGND_c_381_n 0.00179493f $X=0.885 $Y=0.495 $X2=0 $Y2=0
cc_125 N_A2_N_M1009_g N_VGND_c_383_n 0.00366349f $X=0.885 $Y=0.495 $X2=0 $Y2=0
cc_126 N_A2_N_M1009_g N_VGND_c_385_n 0.00606156f $X=0.885 $Y=0.495 $X2=0 $Y2=0
cc_127 N_A2_N_c_99_n N_VGND_c_385_n 7.69802e-19 $X=1.052 $Y=0.985 $X2=0 $Y2=0
cc_128 N_A_145_419#_c_154_n N_B2_M1008_g 0.0220743f $X=1.845 $Y=1.77 $X2=0 $Y2=0
cc_129 N_A_145_419#_c_148_n N_B2_M1003_g 0.0108975f $X=1.845 $Y=1.605 $X2=0
+ $Y2=0
cc_130 N_A_145_419#_c_149_n N_B2_M1003_g 0.016333f $X=1.925 $Y=0.91 $X2=0 $Y2=0
cc_131 N_A_145_419#_c_148_n B2 0.00103962f $X=1.845 $Y=1.605 $X2=0 $Y2=0
cc_132 N_A_145_419#_c_148_n N_B2_c_230_n 0.0220743f $X=1.845 $Y=1.605 $X2=0
+ $Y2=0
cc_133 N_A_145_419#_c_165_n N_VPWR_c_296_n 0.0714415f $X=0.865 $Y=2.24 $X2=0
+ $Y2=0
cc_134 N_A_145_419#_M1002_g N_VPWR_c_297_n 0.0141743f $X=1.795 $Y=2.595 $X2=0
+ $Y2=0
cc_135 N_A_145_419#_c_165_n N_VPWR_c_297_n 0.0630158f $X=0.865 $Y=2.24 $X2=0
+ $Y2=0
cc_136 N_A_145_419#_c_157_n N_VPWR_c_297_n 0.0190817f $X=1.505 $Y=1.85 $X2=0
+ $Y2=0
cc_137 N_A_145_419#_c_153_n N_VPWR_c_297_n 0.00420702f $X=1.67 $Y=1.77 $X2=0
+ $Y2=0
cc_138 N_A_145_419#_c_154_n N_VPWR_c_297_n 4.16361e-19 $X=1.845 $Y=1.77 $X2=0
+ $Y2=0
cc_139 N_A_145_419#_c_165_n N_VPWR_c_300_n 0.019714f $X=0.865 $Y=2.24 $X2=0
+ $Y2=0
cc_140 N_A_145_419#_M1002_g N_VPWR_c_302_n 0.00939541f $X=1.795 $Y=2.595 $X2=0
+ $Y2=0
cc_141 N_A_145_419#_M1006_d N_VPWR_c_294_n 0.00223819f $X=0.725 $Y=2.095 $X2=0
+ $Y2=0
cc_142 N_A_145_419#_M1002_g N_VPWR_c_294_n 0.0165766f $X=1.795 $Y=2.595 $X2=0
+ $Y2=0
cc_143 N_A_145_419#_c_165_n N_VPWR_c_294_n 0.0133473f $X=0.865 $Y=2.24 $X2=0
+ $Y2=0
cc_144 N_A_145_419#_M1002_g N_Y_c_342_n 0.0198138f $X=1.795 $Y=2.595 $X2=0 $Y2=0
cc_145 N_A_145_419#_c_148_n N_Y_c_338_n 0.0151096f $X=1.845 $Y=1.605 $X2=0 $Y2=0
cc_146 N_A_145_419#_c_150_n N_Y_c_338_n 0.00323218f $X=1.925 $Y=0.985 $X2=0
+ $Y2=0
cc_147 N_A_145_419#_c_153_n N_Y_c_338_n 0.0151158f $X=1.67 $Y=1.77 $X2=0 $Y2=0
cc_148 N_A_145_419#_c_154_n N_Y_c_338_n 0.00210444f $X=1.845 $Y=1.77 $X2=0 $Y2=0
cc_149 N_A_145_419#_c_148_n N_Y_c_339_n 0.0099351f $X=1.845 $Y=1.605 $X2=0 $Y2=0
cc_150 N_A_145_419#_c_153_n N_Y_c_339_n 0.024282f $X=1.67 $Y=1.77 $X2=0 $Y2=0
cc_151 N_A_145_419#_c_148_n Y 0.00740804f $X=1.845 $Y=1.605 $X2=0 $Y2=0
cc_152 N_A_145_419#_c_149_n Y 0.00816863f $X=1.925 $Y=0.91 $X2=0 $Y2=0
cc_153 N_A_145_419#_c_150_n Y 0.00677295f $X=1.925 $Y=0.985 $X2=0 $Y2=0
cc_154 N_A_145_419#_c_151_n Y 0.019953f $X=0.755 $Y=0.725 $X2=0 $Y2=0
cc_155 N_A_145_419#_c_151_n N_VGND_c_381_n 0.0204334f $X=0.755 $Y=0.725 $X2=0
+ $Y2=0
cc_156 N_A_145_419#_c_149_n N_VGND_c_382_n 7.2708e-19 $X=1.925 $Y=0.91 $X2=0
+ $Y2=0
cc_157 N_A_145_419#_c_149_n N_VGND_c_383_n 0.00520606f $X=1.925 $Y=0.91 $X2=0
+ $Y2=0
cc_158 N_A_145_419#_c_151_n N_VGND_c_383_n 0.0266861f $X=0.755 $Y=0.725 $X2=0
+ $Y2=0
cc_159 N_A_145_419#_c_149_n N_VGND_c_385_n 0.005315f $X=1.925 $Y=0.91 $X2=0
+ $Y2=0
cc_160 N_A_145_419#_c_151_n N_VGND_c_385_n 0.0202553f $X=0.755 $Y=0.725 $X2=0
+ $Y2=0
cc_161 N_A_145_419#_c_151_n A_114_57# 0.00279363f $X=0.755 $Y=0.725 $X2=-0.19
+ $Y2=-0.245
cc_162 N_A_145_419#_c_149_n N_A_400_83#_c_419_n 0.00144965f $X=1.925 $Y=0.91
+ $X2=0 $Y2=0
cc_163 N_B2_M1008_g N_B1_c_269_n 0.0701758f $X=2.325 $Y=2.595 $X2=-0.19
+ $Y2=-0.245
cc_164 B2 N_B1_c_269_n 0.00158423f $X=2.555 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_165 N_B2_M1003_g N_B1_M1000_g 0.0297177f $X=2.355 $Y=0.625 $X2=0 $Y2=0
cc_166 B2 N_B1_M1000_g 0.00548747f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_167 N_B2_M1008_g N_B1_c_270_n 0.0111173f $X=2.325 $Y=2.595 $X2=0 $Y2=0
cc_168 B2 B1 0.0478954f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_169 N_B2_c_230_n B1 2.2983e-19 $X=2.365 $Y=1.56 $X2=0 $Y2=0
cc_170 N_B2_c_230_n N_B1_c_268_n 0.0206442f $X=2.365 $Y=1.56 $X2=0 $Y2=0
cc_171 N_B2_M1008_g N_VPWR_c_299_n 0.00531277f $X=2.325 $Y=2.595 $X2=0 $Y2=0
cc_172 N_B2_M1008_g N_VPWR_c_302_n 0.00939541f $X=2.325 $Y=2.595 $X2=0 $Y2=0
cc_173 N_B2_M1008_g N_VPWR_c_294_n 0.0161521f $X=2.325 $Y=2.595 $X2=0 $Y2=0
cc_174 N_B2_M1008_g N_Y_c_342_n 0.0227798f $X=2.325 $Y=2.595 $X2=0 $Y2=0
cc_175 N_B2_M1003_g N_Y_c_338_n 5.45964e-19 $X=2.355 $Y=0.625 $X2=0 $Y2=0
cc_176 B2 N_Y_c_338_n 0.0148487f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_177 N_B2_c_230_n N_Y_c_338_n 2.26987e-19 $X=2.365 $Y=1.56 $X2=0 $Y2=0
cc_178 B2 N_Y_c_339_n 0.0273331f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_179 N_B2_c_230_n N_Y_c_339_n 0.0100436f $X=2.365 $Y=1.56 $X2=0 $Y2=0
cc_180 N_B2_M1003_g Y 0.00134917f $X=2.355 $Y=0.625 $X2=0 $Y2=0
cc_181 B2 Y 0.00307067f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_182 N_B2_M1003_g N_VGND_c_382_n 0.00765684f $X=2.355 $Y=0.625 $X2=0 $Y2=0
cc_183 N_B2_M1003_g N_VGND_c_383_n 0.00452954f $X=2.355 $Y=0.625 $X2=0 $Y2=0
cc_184 N_B2_M1003_g N_VGND_c_385_n 0.0044646f $X=2.355 $Y=0.625 $X2=0 $Y2=0
cc_185 N_B2_M1003_g N_A_400_83#_c_422_n 2.62469e-19 $X=2.355 $Y=0.625 $X2=0
+ $Y2=0
cc_186 N_B2_M1003_g N_A_400_83#_c_418_n 0.0113065f $X=2.355 $Y=0.625 $X2=0 $Y2=0
cc_187 B2 N_A_400_83#_c_418_n 0.0370271f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_188 N_B2_c_230_n N_A_400_83#_c_418_n 0.00183855f $X=2.365 $Y=1.56 $X2=0 $Y2=0
cc_189 N_B2_c_230_n N_A_400_83#_c_419_n 9.41275e-19 $X=2.365 $Y=1.56 $X2=0 $Y2=0
cc_190 N_B1_c_269_n N_VPWR_c_299_n 0.0268844f $X=2.815 $Y=2.09 $X2=0 $Y2=0
cc_191 B1 N_VPWR_c_299_n 0.0194919f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_192 N_B1_c_268_n N_VPWR_c_299_n 0.00140236f $X=2.98 $Y=1.56 $X2=0 $Y2=0
cc_193 N_B1_c_269_n N_VPWR_c_302_n 0.008763f $X=2.815 $Y=2.09 $X2=0 $Y2=0
cc_194 N_B1_c_269_n N_VPWR_c_294_n 0.0144563f $X=2.815 $Y=2.09 $X2=0 $Y2=0
cc_195 N_B1_c_269_n N_Y_c_342_n 0.00410437f $X=2.815 $Y=2.09 $X2=0 $Y2=0
cc_196 N_B1_M1000_g N_VGND_c_382_n 0.00378536f $X=2.815 $Y=0.625 $X2=0 $Y2=0
cc_197 N_B1_M1000_g N_VGND_c_384_n 0.00545098f $X=2.815 $Y=0.625 $X2=0 $Y2=0
cc_198 N_B1_M1000_g N_VGND_c_385_n 0.005315f $X=2.815 $Y=0.625 $X2=0 $Y2=0
cc_199 N_B1_M1000_g N_A_400_83#_c_418_n 0.0179903f $X=2.815 $Y=0.625 $X2=0 $Y2=0
cc_200 B1 N_A_400_83#_c_418_n 0.0270611f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_201 N_B1_c_268_n N_A_400_83#_c_418_n 0.00137622f $X=2.98 $Y=1.56 $X2=0 $Y2=0
cc_202 N_B1_M1000_g N_A_400_83#_c_420_n 6.77323e-19 $X=2.815 $Y=0.625 $X2=0
+ $Y2=0
cc_203 N_VPWR_c_294_n N_Y_M1002_d 0.00223819f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_204 N_VPWR_c_297_n N_Y_c_342_n 0.0438f $X=1.395 $Y=2.28 $X2=0 $Y2=0
cc_205 N_VPWR_c_302_n N_Y_c_342_n 0.0177952f $X=2.915 $Y=3.33 $X2=0 $Y2=0
cc_206 N_VPWR_c_294_n N_Y_c_342_n 0.0123247f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_207 N_VPWR_c_294_n A_490_419# 0.010279f $X=3.12 $Y=3.33 $X2=-0.19 $Y2=-0.245
cc_208 Y N_VGND_c_382_n 0.00192202f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_209 Y N_VGND_c_383_n 0.0123222f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_210 Y N_VGND_c_385_n 0.0117582f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_211 Y N_A_400_83#_c_422_n 0.014088f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_212 N_Y_c_338_n N_A_400_83#_c_419_n 0.00260975f $X=2.01 $Y=1.34 $X2=0 $Y2=0
cc_213 Y N_A_400_83#_c_419_n 0.0136942f $X=1.595 $Y=0.47 $X2=0 $Y2=0
cc_214 N_VGND_c_383_n N_A_400_83#_c_422_n 0.00490703f $X=2.405 $Y=0 $X2=0 $Y2=0
cc_215 N_VGND_c_385_n N_A_400_83#_c_422_n 0.00571825f $X=3.12 $Y=0 $X2=0 $Y2=0
cc_216 N_VGND_c_382_n N_A_400_83#_c_418_n 0.0214863f $X=2.57 $Y=0.56 $X2=0 $Y2=0
cc_217 N_VGND_c_385_n N_A_400_83#_c_418_n 0.0125297f $X=3.12 $Y=0 $X2=0 $Y2=0
cc_218 N_VGND_c_384_n N_A_400_83#_c_420_n 0.00778817f $X=3.12 $Y=0 $X2=0 $Y2=0
cc_219 N_VGND_c_385_n N_A_400_83#_c_420_n 0.00948514f $X=3.12 $Y=0 $X2=0 $Y2=0
