* File: sky130_fd_sc_lp__o32a_2.pex.spice
* Created: Fri Aug 28 11:17:25 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O32A_2%A_85_21# 1 2 9 13 17 21 23 27 31 34 36 37 39
+ 43
c90 37 0 1.54109e-19 $X=1.07 $Y=1.505
c91 36 0 2.89487e-20 $X=1.07 $Y=1.505
c92 34 0 2.77137e-20 $X=3.57 $Y=1.71
c93 23 0 1.74055e-19 $X=2.7 $Y=1.77
r94 45 47 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=0.5 $Y=1.505
+ $X2=0.93 $Y2=1.505
r95 41 43 3.55902 $w=3.38e-07 $l=1.05e-07 $layer=LI1_cond $X=3.465 $Y=0.765
+ $X2=3.57 $Y2=0.765
r96 37 47 24.4806 $w=3.3e-07 $l=1.4e-07 $layer=POLY_cond $X=1.07 $Y=1.505
+ $X2=0.93 $Y2=1.505
r97 36 37 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.07
+ $Y=1.505 $X2=1.07 $Y2=1.505
r98 33 43 4.80115 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=3.57 $Y=0.935
+ $X2=3.57 $Y2=0.765
r99 33 34 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=3.57 $Y=0.935
+ $X2=3.57 $Y2=1.71
r100 32 39 7.87875 $w=1.92e-07 $l=3.90461e-07 $layer=LI1_cond $X=3.03 $Y=1.817
+ $X2=2.7 $Y2=1.685
r101 31 34 6.93832 $w=2.15e-07 $l=1.43332e-07 $layer=LI1_cond $X=3.485 $Y=1.817
+ $X2=3.57 $Y2=1.71
r102 31 32 24.3889 $w=2.13e-07 $l=4.55e-07 $layer=LI1_cond $X=3.485 $Y=1.817
+ $X2=3.03 $Y2=1.817
r103 27 29 32.4779 $w=3.28e-07 $l=9.3e-07 $layer=LI1_cond $X=2.865 $Y=1.98
+ $X2=2.865 $Y2=2.91
r104 25 39 0.50483 $w=3.3e-07 $l=3.11769e-07 $layer=LI1_cond $X=2.865 $Y=1.925
+ $X2=2.7 $Y2=1.685
r105 25 27 1.92074 $w=3.28e-07 $l=5.5e-08 $layer=LI1_cond $X=2.865 $Y=1.925
+ $X2=2.865 $Y2=1.98
r106 24 36 11.11 $w=2.91e-07 $l=3.43402e-07 $layer=LI1_cond $X=1.345 $Y=1.77
+ $X2=1.165 $Y2=1.505
r107 23 39 7.87875 $w=1.92e-07 $l=8.5e-08 $layer=LI1_cond $X=2.7 $Y=1.77 $X2=2.7
+ $Y2=1.685
r108 23 24 88.4011 $w=1.68e-07 $l=1.355e-06 $layer=LI1_cond $X=2.7 $Y=1.77
+ $X2=1.345 $Y2=1.77
r109 19 47 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.93 $Y=1.67
+ $X2=0.93 $Y2=1.505
r110 19 21 407.649 $w=1.5e-07 $l=7.95e-07 $layer=POLY_cond $X=0.93 $Y=1.67
+ $X2=0.93 $Y2=2.465
r111 15 47 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.93 $Y=1.34
+ $X2=0.93 $Y2=1.505
r112 15 17 351.245 $w=1.5e-07 $l=6.85e-07 $layer=POLY_cond $X=0.93 $Y=1.34
+ $X2=0.93 $Y2=0.655
r113 11 45 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.5 $Y=1.67
+ $X2=0.5 $Y2=1.505
r114 11 13 407.649 $w=1.5e-07 $l=7.95e-07 $layer=POLY_cond $X=0.5 $Y=1.67
+ $X2=0.5 $Y2=2.465
r115 7 45 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.5 $Y=1.34 $X2=0.5
+ $Y2=1.505
r116 7 9 351.245 $w=1.5e-07 $l=6.85e-07 $layer=POLY_cond $X=0.5 $Y=1.34 $X2=0.5
+ $Y2=0.655
r117 2 29 400 $w=1.7e-07 $l=1.16614e-06 $layer=licon1_PDIFF $count=1 $X=2.675
+ $Y=1.835 $X2=2.865 $Y2=2.91
r118 2 27 400 $w=1.7e-07 $l=2.5229e-07 $layer=licon1_PDIFF $count=1 $X=2.675
+ $Y=1.835 $X2=2.865 $Y2=1.98
r119 1 41 182 $w=1.7e-07 $l=6.08379e-07 $layer=licon1_NDIFF $count=1 $X=3.285
+ $Y=0.235 $X2=3.465 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_LP__O32A_2%A1 3 6 8 11 13
c33 8 0 1.54109e-19 $X=1.68 $Y=1.295
r34 11 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.61 $Y=1.35
+ $X2=1.61 $Y2=1.515
r35 11 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.61 $Y=1.35
+ $X2=1.61 $Y2=1.185
r36 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.61
+ $Y=1.35 $X2=1.61 $Y2=1.35
r37 6 14 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=1.7 $Y=2.465 $X2=1.7
+ $Y2=1.515
r38 3 13 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.63 $Y=0.655
+ $X2=1.63 $Y2=1.185
.ends

.subckt PM_SKY130_FD_SC_LP__O32A_2%A2 3 6 8 11 13
c33 8 0 2.89487e-20 $X=2.16 $Y=1.295
r34 11 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.15 $Y=1.35
+ $X2=2.15 $Y2=1.515
r35 11 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.15 $Y=1.35
+ $X2=2.15 $Y2=1.185
r36 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.15
+ $Y=1.35 $X2=2.15 $Y2=1.35
r37 6 14 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=2.06 $Y=2.465
+ $X2=2.06 $Y2=1.515
r38 3 13 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.06 $Y=0.655
+ $X2=2.06 $Y2=1.185
.ends

.subckt PM_SKY130_FD_SC_LP__O32A_2%A3 3 7 8 11 13
c33 11 0 1.74055e-19 $X=2.69 $Y=1.35
c34 8 0 2.77137e-20 $X=2.64 $Y=1.295
r35 11 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.69 $Y=1.35
+ $X2=2.69 $Y2=1.515
r36 11 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.69 $Y=1.35
+ $X2=2.69 $Y2=1.185
r37 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.69
+ $Y=1.35 $X2=2.69 $Y2=1.35
r38 7 13 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.78 $Y=0.655
+ $X2=2.78 $Y2=1.185
r39 3 14 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=2.6 $Y=2.465 $X2=2.6
+ $Y2=1.515
.ends

.subckt PM_SKY130_FD_SC_LP__O32A_2%B2 3 7 9 12 13
r33 12 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.23 $Y=1.375
+ $X2=3.23 $Y2=1.54
r34 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.23 $Y=1.375
+ $X2=3.23 $Y2=1.21
r35 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.23
+ $Y=1.375 $X2=3.23 $Y2=1.375
r36 9 13 3.84148 $w=3.28e-07 $l=1.1e-07 $layer=LI1_cond $X=3.12 $Y=1.375
+ $X2=3.23 $Y2=1.375
r37 7 14 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=3.21 $Y=0.655
+ $X2=3.21 $Y2=1.21
r38 3 15 474.309 $w=1.5e-07 $l=9.25e-07 $layer=POLY_cond $X=3.14 $Y=2.465
+ $X2=3.14 $Y2=1.54
.ends

.subckt PM_SKY130_FD_SC_LP__O32A_2%B1 3 7 9 10 16
r28 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.93
+ $Y=1.375 $X2=3.93 $Y2=1.375
r29 13 16 43.7153 $w=3.3e-07 $l=2.5e-07 $layer=POLY_cond $X=3.68 $Y=1.375
+ $X2=3.93 $Y2=1.375
r30 10 17 8.56945 $w=3.88e-07 $l=2.9e-07 $layer=LI1_cond $X=4.04 $Y=1.665
+ $X2=4.04 $Y2=1.375
r31 9 17 2.36399 $w=3.88e-07 $l=8e-08 $layer=LI1_cond $X=4.04 $Y=1.295 $X2=4.04
+ $Y2=1.375
r32 5 13 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.68 $Y=1.54
+ $X2=3.68 $Y2=1.375
r33 5 7 474.309 $w=1.5e-07 $l=9.25e-07 $layer=POLY_cond $X=3.68 $Y=1.54 $X2=3.68
+ $Y2=2.465
r34 1 13 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.68 $Y=1.21
+ $X2=3.68 $Y2=1.375
r35 1 3 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=3.68 $Y=1.21 $X2=3.68
+ $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__O32A_2%VPWR 1 2 3 10 12 18 22 24 28 30 35 47 51
r47 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r48 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r49 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r50 42 51 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r51 41 42 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r52 39 48 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r53 38 41 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=1.68 $Y=3.33
+ $X2=3.6 $Y2=3.33
r54 38 39 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r55 36 47 13.3456 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=1.65 $Y=3.33
+ $X2=1.315 $Y2=3.33
r56 36 38 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=1.65 $Y=3.33 $X2=1.68
+ $Y2=3.33
r57 35 50 3.87555 $w=1.7e-07 $l=2.55e-07 $layer=LI1_cond $X=3.81 $Y=3.33
+ $X2=4.065 $Y2=3.33
r58 35 41 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=3.81 $Y=3.33 $X2=3.6
+ $Y2=3.33
r59 34 48 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r60 34 45 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r61 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r62 31 44 4.40602 $w=1.7e-07 $l=2.08e-07 $layer=LI1_cond $X=0.415 $Y=3.33
+ $X2=0.207 $Y2=3.33
r63 31 33 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.415 $Y=3.33
+ $X2=0.72 $Y2=3.33
r64 30 47 13.3456 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=0.98 $Y=3.33
+ $X2=1.315 $Y2=3.33
r65 30 33 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=0.98 $Y=3.33
+ $X2=0.72 $Y2=3.33
r66 28 42 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.6 $Y2=3.33
r67 28 39 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r68 24 27 36.1867 $w=2.48e-07 $l=7.85e-07 $layer=LI1_cond $X=3.935 $Y=2.165
+ $X2=3.935 $Y2=2.95
r69 22 50 3.26762 $w=2.5e-07 $l=1.67183e-07 $layer=LI1_cond $X=3.935 $Y=3.245
+ $X2=4.065 $Y2=3.33
r70 22 27 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=3.935 $Y=3.245
+ $X2=3.935 $Y2=2.95
r71 18 21 14.9956 $w=6.68e-07 $l=8.4e-07 $layer=LI1_cond $X=1.315 $Y=2.11
+ $X2=1.315 $Y2=2.95
r72 16 47 2.76849 $w=6.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.315 $Y=3.245
+ $X2=1.315 $Y2=3.33
r73 16 21 5.26632 $w=6.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.315 $Y=3.245
+ $X2=1.315 $Y2=2.95
r74 12 15 37.8939 $w=2.93e-07 $l=9.7e-07 $layer=LI1_cond $X=0.267 $Y=1.98
+ $X2=0.267 $Y2=2.95
r75 10 44 3.0715 $w=2.95e-07 $l=1.11018e-07 $layer=LI1_cond $X=0.267 $Y=3.245
+ $X2=0.207 $Y2=3.33
r76 10 15 11.5244 $w=2.93e-07 $l=2.95e-07 $layer=LI1_cond $X=0.267 $Y=3.245
+ $X2=0.267 $Y2=2.95
r77 3 27 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=3.755
+ $Y=1.835 $X2=3.895 $Y2=2.95
r78 3 24 400 $w=1.7e-07 $l=3.93827e-07 $layer=licon1_PDIFF $count=1 $X=3.755
+ $Y=1.835 $X2=3.895 $Y2=2.165
r79 2 21 200 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=3 $X=1.005
+ $Y=1.835 $X2=1.145 $Y2=2.95
r80 2 18 200 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=3 $X=1.005
+ $Y=1.835 $X2=1.145 $Y2=2.11
r81 1 15 400 $w=1.7e-07 $l=1.17584e-06 $layer=licon1_PDIFF $count=1 $X=0.16
+ $Y=1.835 $X2=0.285 $Y2=2.95
r82 1 12 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.16
+ $Y=1.835 $X2=0.285 $Y2=1.98
.ends

.subckt PM_SKY130_FD_SC_LP__O32A_2%X 1 2 7 8 9 10 11 12 13 22
r16 13 40 6.91466 $w=2.23e-07 $l=1.35e-07 $layer=LI1_cond $X=0.697 $Y=2.775
+ $X2=0.697 $Y2=2.91
r17 12 13 18.9513 $w=2.23e-07 $l=3.7e-07 $layer=LI1_cond $X=0.697 $Y=2.405
+ $X2=0.697 $Y2=2.775
r18 11 12 19.9757 $w=2.23e-07 $l=3.9e-07 $layer=LI1_cond $X=0.697 $Y=2.015
+ $X2=0.697 $Y2=2.405
r19 10 11 17.9269 $w=2.23e-07 $l=3.5e-07 $layer=LI1_cond $X=0.697 $Y=1.665
+ $X2=0.697 $Y2=2.015
r20 9 10 18.9513 $w=2.23e-07 $l=3.7e-07 $layer=LI1_cond $X=0.697 $Y=1.295
+ $X2=0.697 $Y2=1.665
r21 8 9 18.9513 $w=2.23e-07 $l=3.7e-07 $layer=LI1_cond $X=0.697 $Y=0.925
+ $X2=0.697 $Y2=1.295
r22 7 8 18.9513 $w=2.23e-07 $l=3.7e-07 $layer=LI1_cond $X=0.697 $Y=0.555
+ $X2=0.697 $Y2=0.925
r23 7 22 6.91466 $w=2.23e-07 $l=1.35e-07 $layer=LI1_cond $X=0.697 $Y=0.555
+ $X2=0.697 $Y2=0.42
r24 2 40 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=0.575
+ $Y=1.835 $X2=0.715 $Y2=2.91
r25 2 11 400 $w=1.7e-07 $l=2.4e-07 $layer=licon1_PDIFF $count=1 $X=0.575
+ $Y=1.835 $X2=0.715 $Y2=2.015
r26 1 22 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=0.575
+ $Y=0.235 $X2=0.715 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__O32A_2%VGND 1 2 3 10 12 16 20 23 24 25 27 40 41 47
r55 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r56 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r57 40 41 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r58 38 41 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=2.64 $Y=0 $X2=4.08
+ $Y2=0
r59 37 40 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=2.64 $Y=0 $X2=4.08
+ $Y2=0
r60 37 38 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r61 32 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.44 $Y=0 $X2=1.275
+ $Y2=0
r62 32 34 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=1.44 $Y=0 $X2=2.16
+ $Y2=0
r63 31 48 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r64 31 45 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r65 30 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r66 28 44 4.40602 $w=1.7e-07 $l=2.08e-07 $layer=LI1_cond $X=0.415 $Y=0 $X2=0.207
+ $Y2=0
r67 28 30 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.415 $Y=0 $X2=0.72
+ $Y2=0
r68 27 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.11 $Y=0 $X2=1.275
+ $Y2=0
r69 27 30 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=1.11 $Y=0 $X2=0.72
+ $Y2=0
r70 25 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r71 25 48 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.2
+ $Y2=0
r72 25 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r73 23 34 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=2.25 $Y=0 $X2=2.16
+ $Y2=0
r74 23 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.25 $Y=0 $X2=2.415
+ $Y2=0
r75 22 37 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=2.58 $Y=0 $X2=2.64
+ $Y2=0
r76 22 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.58 $Y=0 $X2=2.415
+ $Y2=0
r77 18 24 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.415 $Y=0.085
+ $X2=2.415 $Y2=0
r78 18 20 17.112 $w=3.28e-07 $l=4.9e-07 $layer=LI1_cond $X=2.415 $Y=0.085
+ $X2=2.415 $Y2=0.575
r79 14 47 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.275 $Y=0.085
+ $X2=1.275 $Y2=0
r80 14 16 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.275 $Y=0.085
+ $X2=1.275 $Y2=0.38
r81 10 44 3.0715 $w=2.95e-07 $l=1.11018e-07 $layer=LI1_cond $X=0.267 $Y=0.085
+ $X2=0.207 $Y2=0
r82 10 12 11.5244 $w=2.93e-07 $l=2.95e-07 $layer=LI1_cond $X=0.267 $Y=0.085
+ $X2=0.267 $Y2=0.38
r83 3 20 182 $w=1.7e-07 $l=4.5913e-07 $layer=licon1_NDIFF $count=1 $X=2.135
+ $Y=0.235 $X2=2.415 $Y2=0.575
r84 2 16 91 $w=1.7e-07 $l=3.34739e-07 $layer=licon1_NDIFF $count=2 $X=1.005
+ $Y=0.235 $X2=1.275 $Y2=0.38
r85 1 12 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.16
+ $Y=0.235 $X2=0.285 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_LP__O32A_2%A_341_47# 1 2 3 12 14 15 16 17 18 25
r50 19 23 4.79851 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=3.13 $Y=0.34 $X2=2.98
+ $Y2=0.34
r51 18 25 4.47015 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=3.825 $Y=0.34
+ $X2=3.96 $Y2=0.34
r52 18 19 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=3.825 $Y=0.34
+ $X2=3.13 $Y2=0.34
r53 16 23 2.71916 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.98 $Y=0.425 $X2=2.98
+ $Y2=0.34
r54 16 17 17.0946 $w=2.98e-07 $l=4.45e-07 $layer=LI1_cond $X=2.98 $Y=0.425
+ $X2=2.98 $Y2=0.87
r55 14 17 7.51767 $w=1.7e-07 $l=1.8775e-07 $layer=LI1_cond $X=2.83 $Y=0.955
+ $X2=2.98 $Y2=0.87
r56 14 15 53.4973 $w=1.68e-07 $l=8.2e-07 $layer=LI1_cond $X=2.83 $Y=0.955
+ $X2=2.01 $Y2=0.955
r57 10 15 16.7971 $w=1.15e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.845 $Y=0.87
+ $X2=2.01 $Y2=0.955
r58 10 12 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=1.845 $Y=0.87
+ $X2=1.845 $Y2=0.42
r59 3 25 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=3.755
+ $Y=0.235 $X2=3.91 $Y2=0.42
r60 2 23 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=2.855
+ $Y=0.235 $X2=2.995 $Y2=0.42
r61 1 12 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=1.705
+ $Y=0.235 $X2=1.845 $Y2=0.42
.ends

