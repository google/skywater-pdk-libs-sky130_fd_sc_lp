* File: sky130_fd_sc_lp__a211oi_1.pex.spice
* Created: Fri Aug 28 09:48:16 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A211OI_1%A2 1 3 6 8 9 16
r27 13 16 30.6007 $w=3.3e-07 $l=1.75e-07 $layer=POLY_cond $X=0.3 $Y=1.375
+ $X2=0.475 $Y2=1.375
r28 8 9 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.26 $Y=1.295 $X2=0.26
+ $Y2=1.665
r29 8 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.3
+ $Y=1.375 $X2=0.3 $Y2=1.375
r30 4 16 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=1.54
+ $X2=0.475 $Y2=1.375
r31 4 6 474.309 $w=1.5e-07 $l=9.25e-07 $layer=POLY_cond $X=0.475 $Y=1.54
+ $X2=0.475 $Y2=2.465
r32 1 16 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=1.21
+ $X2=0.475 $Y2=1.375
r33 1 3 175.127 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=0.475 $Y=1.21
+ $X2=0.475 $Y2=0.665
.ends

.subckt PM_SKY130_FD_SC_LP__A211OI_1%A1 3 6 8 9 10 11 17 19
c40 11 0 1.87627e-19 $X=0.72 $Y=1.665
r41 17 20 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.925 $Y=1.36
+ $X2=0.925 $Y2=1.525
r42 17 19 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.925 $Y=1.36
+ $X2=0.925 $Y2=1.195
r43 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.925
+ $Y=1.36 $X2=0.925 $Y2=1.36
r44 11 18 10.3939 $w=3.58e-07 $l=3.05e-07 $layer=LI1_cond $X=0.802 $Y=1.665
+ $X2=0.802 $Y2=1.36
r45 10 18 2.21508 $w=3.58e-07 $l=6.5e-08 $layer=LI1_cond $X=0.802 $Y=1.295
+ $X2=0.802 $Y2=1.36
r46 10 21 4.53139 $w=3.58e-07 $l=1.34907e-07 $layer=LI1_cond $X=0.802 $Y=1.295
+ $X2=0.72 $Y2=1.195
r47 9 21 12.4464 $w=2.48e-07 $l=2.7e-07 $layer=LI1_cond $X=0.72 $Y=0.925
+ $X2=0.72 $Y2=1.195
r48 8 9 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=0.72 $Y=0.555 $X2=0.72
+ $Y2=0.925
r49 6 20 482 $w=1.5e-07 $l=9.4e-07 $layer=POLY_cond $X=1.015 $Y=2.465 $X2=1.015
+ $Y2=1.525
r50 3 19 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.835 $Y=0.665
+ $X2=0.835 $Y2=1.195
.ends

.subckt PM_SKY130_FD_SC_LP__A211OI_1%B1 3 7 9 12
c34 12 0 1.87627e-19 $X=1.465 $Y=1.51
r35 12 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.465 $Y=1.51
+ $X2=1.465 $Y2=1.675
r36 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.465 $Y=1.51
+ $X2=1.465 $Y2=1.345
r37 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.465
+ $Y=1.51 $X2=1.465 $Y2=1.51
r38 9 13 5.97049 $w=4.13e-07 $l=2.15e-07 $layer=LI1_cond $X=1.68 $Y=1.552
+ $X2=1.465 $Y2=1.552
r39 7 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.555 $Y=2.465
+ $X2=1.555 $Y2=1.675
r40 3 14 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=1.375 $Y=0.665
+ $X2=1.375 $Y2=1.345
.ends

.subckt PM_SKY130_FD_SC_LP__A211OI_1%C1 3 7 9 14 15
r28 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.135
+ $Y=1.46 $X2=2.135 $Y2=1.46
r29 11 14 38.4695 $w=3.3e-07 $l=2.2e-07 $layer=POLY_cond $X=1.915 $Y=1.46
+ $X2=2.135 $Y2=1.46
r30 9 15 7.05226 $w=3.33e-07 $l=2.05e-07 $layer=LI1_cond $X=2.137 $Y=1.665
+ $X2=2.137 $Y2=1.46
r31 5 11 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.915 $Y=1.625
+ $X2=1.915 $Y2=1.46
r32 5 7 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=1.915 $Y=1.625
+ $X2=1.915 $Y2=2.465
r33 1 11 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.915 $Y=1.295
+ $X2=1.915 $Y2=1.46
r34 1 3 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=1.915 $Y=1.295
+ $X2=1.915 $Y2=0.665
.ends

.subckt PM_SKY130_FD_SC_LP__A211OI_1%A_27_367# 1 2 7 9 11 13 15
r22 13 20 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.29 $Y=2.1 $X2=1.29
+ $Y2=2.015
r23 13 15 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=1.29 $Y=2.1
+ $X2=1.29 $Y2=2.455
r24 12 18 4.96789 $w=1.7e-07 $l=1.58e-07 $layer=LI1_cond $X=0.41 $Y=2.015
+ $X2=0.252 $Y2=2.015
r25 11 20 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.125 $Y=2.015
+ $X2=1.29 $Y2=2.015
r26 11 12 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=1.125 $Y=2.015
+ $X2=0.41 $Y2=2.015
r27 7 18 2.6726 $w=3.15e-07 $l=8.5e-08 $layer=LI1_cond $X=0.252 $Y=2.1 $X2=0.252
+ $Y2=2.015
r28 7 9 29.6342 $w=3.13e-07 $l=8.1e-07 $layer=LI1_cond $X=0.252 $Y=2.1 $X2=0.252
+ $Y2=2.91
r29 2 20 600 $w=1.7e-07 $l=2.75681e-07 $layer=licon1_PDIFF $count=1 $X=1.09
+ $Y=1.835 $X2=1.29 $Y2=2.015
r30 2 15 300 $w=1.7e-07 $l=7.13022e-07 $layer=licon1_PDIFF $count=2 $X=1.09
+ $Y=1.835 $X2=1.29 $Y2=2.455
r31 1 18 400 $w=1.7e-07 $l=2.34307e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.835 $X2=0.26 $Y2=2.015
r32 1 9 400 $w=1.7e-07 $l=1.13578e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.835 $X2=0.26 $Y2=2.91
.ends

.subckt PM_SKY130_FD_SC_LP__A211OI_1%VPWR 1 6 8 10 20 21 24
r28 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r29 20 21 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r30 18 25 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r31 17 20 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r32 17 18 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r33 15 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.91 $Y=3.33
+ $X2=0.745 $Y2=3.33
r34 15 17 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=0.91 $Y=3.33 $X2=1.2
+ $Y2=3.33
r35 13 25 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r36 12 13 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r37 10 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.58 $Y=3.33
+ $X2=0.745 $Y2=3.33
r38 10 12 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=0.58 $Y=3.33
+ $X2=0.24 $Y2=3.33
r39 8 21 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=2.64 $Y2=3.33
r40 8 18 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=1.2 $Y2=3.33
r41 4 24 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.745 $Y=3.245
+ $X2=0.745 $Y2=3.33
r42 4 6 29.6841 $w=3.28e-07 $l=8.5e-07 $layer=LI1_cond $X=0.745 $Y=3.245
+ $X2=0.745 $Y2=2.395
r43 1 6 300 $w=1.7e-07 $l=6.50231e-07 $layer=licon1_PDIFF $count=2 $X=0.55
+ $Y=1.835 $X2=0.745 $Y2=2.395
.ends

.subckt PM_SKY130_FD_SC_LP__A211OI_1%Y 1 2 3 10 12 18 24 25 27 28 29 34 35
r44 34 35 6.65594 $w=8.18e-07 $l=8.5e-08 $layer=LI1_cond $X=2.375 $Y=2.01
+ $X2=2.375 $Y2=1.925
r45 29 43 2.55261 $w=8.18e-07 $l=1.75e-07 $layer=LI1_cond $X=2.375 $Y=2.775
+ $X2=2.375 $Y2=2.95
r46 28 29 5.39694 $w=8.18e-07 $l=3.7e-07 $layer=LI1_cond $X=2.375 $Y=2.405
+ $X2=2.375 $Y2=2.775
r47 27 28 5.39694 $w=8.18e-07 $l=3.7e-07 $layer=LI1_cond $X=2.375 $Y=2.035
+ $X2=2.375 $Y2=2.405
r48 27 34 0.364658 $w=8.18e-07 $l=2.5e-08 $layer=LI1_cond $X=2.375 $Y=2.035
+ $X2=2.375 $Y2=2.01
r49 23 25 19.2736 $w=2.88e-07 $l=4.85e-07 $layer=LI1_cond $X=2.157 $Y=1.03
+ $X2=2.642 $Y2=1.03
r50 23 24 7.09248 $w=2.88e-07 $l=1.37e-07 $layer=LI1_cond $X=2.157 $Y=1.03
+ $X2=2.02 $Y2=1.03
r51 20 25 0.843369 $w=2.85e-07 $l=1.45e-07 $layer=LI1_cond $X=2.642 $Y=1.175
+ $X2=2.642 $Y2=1.03
r52 20 35 30.3274 $w=2.83e-07 $l=7.5e-07 $layer=LI1_cond $X=2.642 $Y=1.175
+ $X2=2.642 $Y2=1.925
r53 16 23 1.05929 $w=2.75e-07 $l=1.45e-07 $layer=LI1_cond $X=2.157 $Y=0.885
+ $X2=2.157 $Y2=1.03
r54 16 18 19.4868 $w=2.73e-07 $l=4.65e-07 $layer=LI1_cond $X=2.157 $Y=0.885
+ $X2=2.157 $Y2=0.42
r55 15 22 2.49649 $w=1.8e-07 $l=1.68e-07 $layer=LI1_cond $X=1.35 $Y=1.085
+ $X2=1.182 $Y2=1.085
r56 15 24 41.2828 $w=1.78e-07 $l=6.7e-07 $layer=LI1_cond $X=1.35 $Y=1.085
+ $X2=2.02 $Y2=1.085
r57 10 22 11.3933 $w=3.35e-07 $l=2.87e-07 $layer=LI1_cond $X=1.182 $Y=0.798
+ $X2=1.182 $Y2=1.085
r58 10 12 13.0037 $w=3.33e-07 $l=3.78e-07 $layer=LI1_cond $X=1.182 $Y=0.798
+ $X2=1.182 $Y2=0.42
r59 3 43 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=1.99
+ $Y=1.835 $X2=2.13 $Y2=2.95
r60 3 34 400 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_PDIFF $count=1 $X=1.99
+ $Y=1.835 $X2=2.13 $Y2=2.01
r61 2 18 91 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=2 $X=1.99
+ $Y=0.245 $X2=2.13 $Y2=0.42
r62 1 12 91 $w=1.7e-07 $l=2.94788e-07 $layer=licon1_NDIFF $count=2 $X=0.91
+ $Y=0.245 $X2=1.13 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__A211OI_1%VGND 1 2 7 9 13 15 17 24 25 31
r35 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r36 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r37 25 32 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=1.68
+ $Y2=0
r38 24 25 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r39 22 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.85 $Y=0 $X2=1.685
+ $Y2=0
r40 22 24 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=1.85 $Y=0 $X2=2.64
+ $Y2=0
r41 21 29 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.24
+ $Y2=0
r42 20 21 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r43 18 28 4.78091 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=0 $X2=0.212
+ $Y2=0
r44 18 20 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=0.425 $Y=0 $X2=1.2
+ $Y2=0
r45 17 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.52 $Y=0 $X2=1.685
+ $Y2=0
r46 17 20 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=1.52 $Y=0 $X2=1.2
+ $Y2=0
r47 15 32 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=1.68
+ $Y2=0
r48 15 21 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=1.2
+ $Y2=0
r49 11 31 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.685 $Y=0.085
+ $X2=1.685 $Y2=0
r50 11 13 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=1.685 $Y=0.085
+ $X2=1.685 $Y2=0.37
r51 7 28 2.98526 $w=3.3e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.212 $Y2=0
r52 7 9 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.26 $Y2=0.39
r53 2 13 91 $w=1.7e-07 $l=2.90861e-07 $layer=licon1_NDIFF $count=2 $X=1.45
+ $Y=0.245 $X2=1.685 $Y2=0.37
r54 1 9 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.245 $X2=0.26 $Y2=0.39
.ends

