* File: sky130_fd_sc_lp__invkapwr_1.pex.spice
* Created: Wed Sep  2 09:56:26 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__INVKAPWR_1%A 3 7 9 11 13 14 15
r32 20 22 12.5087 $w=5.78e-07 $l=1.5e-07 $layer=POLY_cond $X=0.385 $Y=1.44
+ $X2=0.535 $Y2=1.44
r33 20 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.385
+ $Y=1.27 $X2=0.385 $Y2=1.27
r34 14 15 11.5244 $w=3.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.29 $Y=1.295
+ $X2=0.29 $Y2=1.665
r35 14 21 0.778678 $w=3.68e-07 $l=2.5e-08 $layer=LI1_cond $X=0.29 $Y=1.295
+ $X2=0.29 $Y2=1.27
r36 13 21 10.7458 $w=3.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.29 $Y=0.925
+ $X2=0.29 $Y2=1.27
r37 9 22 35.8581 $w=5.78e-07 $l=4.3e-07 $layer=POLY_cond $X=0.965 $Y=1.44
+ $X2=0.535 $Y2=1.44
r38 9 11 476.872 $w=1.5e-07 $l=9.3e-07 $layer=POLY_cond $X=0.965 $Y=1.6
+ $X2=0.965 $Y2=2.53
r39 5 9 35.1088 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=0.965 $Y=1.105
+ $X2=0.965 $Y2=1.44
r40 5 7 279.457 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=0.965 $Y=1.105
+ $X2=0.965 $Y2=0.56
r41 1 22 35.1088 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=0.535 $Y=1.775
+ $X2=0.535 $Y2=1.44
r42 1 3 387.138 $w=1.5e-07 $l=7.55e-07 $layer=POLY_cond $X=0.535 $Y=1.775
+ $X2=0.535 $Y2=2.53
.ends

.subckt PM_SKY130_FD_SC_LP__INVKAPWR_1%KAPWR 1 2 7 10 17 21 27
r21 21 27 0.245948 $w=2.55e-07 $l=4.25e-07 $layer=MET1_cond $X=1.175 $Y=2.817
+ $X2=0.75 $Y2=2.817
r22 20 21 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.175 $Y=2.81
+ $X2=1.175 $Y2=2.81
r23 17 20 17.8629 $w=2.98e-07 $l=4.65e-07 $layer=LI1_cond $X=1.195 $Y=2.345
+ $X2=1.195 $Y2=2.81
r24 13 14 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.305 $Y=2.81
+ $X2=0.305 $Y2=2.81
r25 10 13 16.7464 $w=3.18e-07 $l=4.65e-07 $layer=LI1_cond $X=0.315 $Y=2.345
+ $X2=0.315 $Y2=2.81
r26 7 27 0.0173611 $w=2.55e-07 $l=3e-08 $layer=MET1_cond $X=0.72 $Y=2.817
+ $X2=0.75 $Y2=2.817
r27 7 14 0.240161 $w=2.55e-07 $l=4.15e-07 $layer=MET1_cond $X=0.72 $Y=2.817
+ $X2=0.305 $Y2=2.817
r28 2 17 300 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_PDIFF $count=2 $X=1.04
+ $Y=2.11 $X2=1.18 $Y2=2.345
r29 1 10 300 $w=1.7e-07 $l=2.90861e-07 $layer=licon1_PDIFF $count=2 $X=0.195
+ $Y=2.11 $X2=0.32 $Y2=2.345
.ends

.subckt PM_SKY130_FD_SC_LP__INVKAPWR_1%Y 1 2 9 13 15 16 17
r26 17 32 9.57519 $w=6.38e-07 $l=2.35e-07 $layer=LI1_cond $X=0.965 $Y=1.665
+ $X2=0.965 $Y2=1.9
r27 16 17 4.76877 $w=8.08e-07 $l=2.85e-07 $layer=LI1_cond $X=0.965 $Y=1.295
+ $X2=0.965 $Y2=1.58
r28 16 22 2.52298 $w=6.38e-07 $l=1.35e-07 $layer=LI1_cond $X=0.965 $Y=1.295
+ $X2=0.965 $Y2=1.16
r29 15 22 4.39185 $w=6.38e-07 $l=2.35e-07 $layer=LI1_cond $X=0.965 $Y=0.925
+ $X2=0.965 $Y2=1.16
r30 15 28 7.75425 $w=6.38e-07 $l=8.5e-08 $layer=LI1_cond $X=0.965 $Y=0.925
+ $X2=0.965 $Y2=0.84
r31 13 32 22.2973 $w=2.28e-07 $l=4.45e-07 $layer=LI1_cond $X=0.76 $Y=2.345
+ $X2=0.76 $Y2=1.9
r32 9 28 15.5273 $w=1.98e-07 $l=2.8e-07 $layer=LI1_cond $X=0.745 $Y=0.56
+ $X2=0.745 $Y2=0.84
r33 2 13 300 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_PDIFF $count=2 $X=0.61
+ $Y=2.11 $X2=0.75 $Y2=2.345
r34 1 9 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.625
+ $Y=0.35 $X2=0.75 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_LP__INVKAPWR_1%VGND 1 4 6 8 10 17
r12 16 17 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r13 10 16 4.78613 $w=1.7e-07 $l=2.12e-07 $layer=LI1_cond $X=1.015 $Y=0 $X2=1.227
+ $Y2=0
r14 10 12 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.015 $Y=0 $X2=0.72
+ $Y2=0
r15 8 17 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r16 8 12 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r17 4 16 2.98004 $w=3.3e-07 $l=1.05924e-07 $layer=LI1_cond $X=1.18 $Y=0.085
+ $X2=1.227 $Y2=0
r18 4 6 16.5882 $w=3.28e-07 $l=4.75e-07 $layer=LI1_cond $X=1.18 $Y=0.085
+ $X2=1.18 $Y2=0.56
r19 1 6 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.04
+ $Y=0.35 $X2=1.18 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_LP__INVKAPWR_1%VPWR 1 8 14
r15 5 14 0.0108064 $w=1.44e-06 $l=1.22e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.208
r16 5 8 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r17 4 8 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.24 $Y=3.33 $X2=1.2
+ $Y2=3.33
r18 4 5 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33 $X2=0.24
+ $Y2=3.33
r19 1 14 8.85771e-05 $w=1.44e-06 $l=1e-09 $layer=MET1_cond $X=0.72 $Y=3.207
+ $X2=0.72 $Y2=3.208
.ends

