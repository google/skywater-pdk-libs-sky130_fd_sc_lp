* File: sky130_fd_sc_lp__a21bo_lp.pex.spice
* Created: Wed Sep  2 09:18:59 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A21BO_LP%A_84_29# 1 2 9 11 13 17 21 23 24 26 27 29
+ 30 33 37 41 42
c94 13 0 2.1464e-19 $X=0.595 $Y=2.545
r95 40 41 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.605
+ $Y=1.06 $X2=0.605 $Y2=1.06
r96 35 37 2.09535 $w=3.28e-07 $l=6e-08 $layer=LI1_cond $X=1.93 $Y=2.13 $X2=1.93
+ $Y2=2.19
r97 31 33 14.1436 $w=3.28e-07 $l=4.05e-07 $layer=LI1_cond $X=1.89 $Y=0.895
+ $X2=1.89 $Y2=0.49
r98 29 35 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.765 $Y=2.045
+ $X2=1.93 $Y2=2.13
r99 29 30 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=1.765 $Y=2.045
+ $X2=0.845 $Y2=2.045
r100 28 40 5.93104 $w=1.7e-07 $l=2.03e-07 $layer=LI1_cond $X=0.845 $Y=0.98
+ $X2=0.642 $Y2=0.98
r101 27 31 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.725 $Y=0.98
+ $X2=1.89 $Y2=0.895
r102 27 28 57.4118 $w=1.68e-07 $l=8.8e-07 $layer=LI1_cond $X=1.725 $Y=0.98
+ $X2=0.845 $Y2=0.98
r103 26 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.76 $Y=1.96
+ $X2=0.845 $Y2=2.045
r104 26 42 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=0.76 $Y=1.96
+ $X2=0.76 $Y2=1.565
r105 24 42 9.72165 $w=4.03e-07 $l=2.02e-07 $layer=LI1_cond $X=0.642 $Y=1.363
+ $X2=0.642 $Y2=1.565
r106 23 40 2.48344 $w=4.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.642 $Y=1.065
+ $X2=0.642 $Y2=0.98
r107 23 24 8.4797 $w=4.03e-07 $l=2.98e-07 $layer=LI1_cond $X=0.642 $Y=1.065
+ $X2=0.642 $Y2=1.363
r108 22 41 54.4068 $w=3.5e-07 $l=3.3e-07 $layer=POLY_cond $X=0.595 $Y=1.39
+ $X2=0.595 $Y2=1.06
r109 21 41 3.29738 $w=3.5e-07 $l=2e-08 $layer=POLY_cond $X=0.595 $Y=1.04
+ $X2=0.595 $Y2=1.06
r110 11 22 31.2502 $w=3.5e-07 $l=1.75e-07 $layer=POLY_cond $X=0.595 $Y=1.565
+ $X2=0.595 $Y2=1.39
r111 11 13 243.485 $w=2.5e-07 $l=9.8e-07 $layer=POLY_cond $X=0.595 $Y=1.565
+ $X2=0.595 $Y2=2.545
r112 7 21 26.0701 $w=3.5e-07 $l=1.5e-07 $layer=POLY_cond $X=0.675 $Y=0.89
+ $X2=0.675 $Y2=1.04
r113 7 17 207.67 $w=1.5e-07 $l=4.05e-07 $layer=POLY_cond $X=0.855 $Y=0.89
+ $X2=0.855 $Y2=0.485
r114 7 9 207.67 $w=1.5e-07 $l=4.05e-07 $layer=POLY_cond $X=0.495 $Y=0.89
+ $X2=0.495 $Y2=0.485
r115 2 37 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=1.79
+ $Y=2.045 $X2=1.93 $Y2=2.19
r116 1 33 182 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_NDIFF $count=1 $X=1.75
+ $Y=0.275 $X2=1.89 $Y2=0.49
.ends

.subckt PM_SKY130_FD_SC_LP__A21BO_LP%A2 3 9 10 11 12 15 16 17
c48 11 0 1.57471e-19 $X=1.282 $Y=0.92
r49 15 18 32.0725 $w=3.45e-07 $l=1.65e-07 $layer=POLY_cond $X=1.182 $Y=1.445
+ $X2=1.182 $Y2=1.61
r50 15 17 46.3655 $w=3.45e-07 $l=1.65e-07 $layer=POLY_cond $X=1.182 $Y=1.445
+ $X2=1.182 $Y2=1.28
r51 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.19
+ $Y=1.445 $X2=1.19 $Y2=1.445
r52 12 16 7.68295 $w=3.28e-07 $l=2.2e-07 $layer=LI1_cond $X=1.19 $Y=1.665
+ $X2=1.19 $Y2=1.445
r53 11 17 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=1.28 $Y=0.92
+ $X2=1.28 $Y2=1.28
r54 10 11 71.7618 $w=1.55e-07 $l=1.5e-07 $layer=POLY_cond $X=1.282 $Y=0.77
+ $X2=1.282 $Y2=0.92
r55 9 10 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=1.285 $Y=0.485
+ $X2=1.285 $Y2=0.77
r56 3 18 232.304 $w=2.5e-07 $l=9.35e-07 $layer=POLY_cond $X=1.135 $Y=2.545
+ $X2=1.135 $Y2=1.61
.ends

.subckt PM_SKY130_FD_SC_LP__A21BO_LP%A1 3 7 12 13 17 24 26 29
c61 26 0 9.52166e-20 $X=2.755 $Y=1.77
c62 24 0 1.08855e-19 $X=2.66 $Y=1.77
r63 23 26 16.6118 $w=3.3e-07 $l=9.5e-08 $layer=POLY_cond $X=2.66 $Y=1.77
+ $X2=2.755 $Y2=1.77
r64 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.66
+ $Y=1.77 $X2=2.66 $Y2=1.77
r65 17 24 0.598672 $w=3.83e-07 $l=2e-08 $layer=LI1_cond $X=2.64 $Y=1.742
+ $X2=2.66 $Y2=1.742
r66 17 29 7.99026 $w=3.83e-07 $l=1.45e-07 $layer=LI1_cond $X=2.64 $Y=1.742
+ $X2=2.495 $Y2=1.742
r67 13 20 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.76 $Y=1.415
+ $X2=1.76 $Y2=1.25
r68 12 15 7.68295 $w=3.28e-07 $l=2.2e-07 $layer=LI1_cond $X=1.76 $Y=1.415
+ $X2=1.76 $Y2=1.635
r69 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.76
+ $Y=1.415 $X2=1.76 $Y2=1.415
r70 10 15 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.925 $Y=1.635
+ $X2=1.76 $Y2=1.635
r71 10 29 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=1.925 $Y=1.635
+ $X2=2.495 $Y2=1.635
r72 5 26 9.34494 $w=2.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.755 $Y=1.935
+ $X2=2.755 $Y2=1.77
r73 5 7 163.979 $w=2.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.755 $Y=1.935
+ $X2=2.755 $Y2=2.595
r74 3 20 392.266 $w=1.5e-07 $l=7.65e-07 $layer=POLY_cond $X=1.675 $Y=0.485
+ $X2=1.675 $Y2=1.25
.ends

.subckt PM_SKY130_FD_SC_LP__A21BO_LP%A_308_364# 1 2 7 9 10 11 12 14 16 17 19 20
+ 24 28 32 36 38 39
c92 32 0 9.52166e-20 $X=2.415 $Y=0.77
r93 36 43 8.16949 $w=2.95e-07 $l=5e-08 $layer=POLY_cond $X=2.415 $Y=0.97
+ $X2=2.465 $Y2=0.97
r94 36 41 33.4949 $w=2.95e-07 $l=2.05e-07 $layer=POLY_cond $X=2.415 $Y=0.97
+ $X2=2.21 $Y2=0.97
r95 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.415
+ $Y=0.97 $X2=2.415 $Y2=0.97
r96 32 35 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=2.415 $Y=0.77 $X2=2.415
+ $Y2=0.97
r97 30 38 3.70735 $w=2.5e-07 $l=1.56844e-07 $layer=LI1_cond $X=3.63 $Y=0.855
+ $X2=3.51 $Y2=0.77
r98 30 39 79.5936 $w=1.68e-07 $l=1.22e-06 $layer=LI1_cond $X=3.63 $Y=0.855
+ $X2=3.63 $Y2=2.075
r99 28 39 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=3.55 $Y=2.24
+ $X2=3.55 $Y2=2.075
r100 22 38 3.70735 $w=2.5e-07 $l=1.03078e-07 $layer=LI1_cond $X=3.47 $Y=0.685
+ $X2=3.51 $Y2=0.77
r101 22 24 6.80989 $w=3.28e-07 $l=1.95e-07 $layer=LI1_cond $X=3.47 $Y=0.685
+ $X2=3.47 $Y2=0.49
r102 21 32 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.58 $Y=0.77
+ $X2=2.415 $Y2=0.77
r103 20 38 2.76166 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=3.305 $Y=0.77
+ $X2=3.51 $Y2=0.77
r104 20 21 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=3.305 $Y=0.77
+ $X2=2.58 $Y2=0.77
r105 17 43 18.5736 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.465 $Y=0.805
+ $X2=2.465 $Y2=0.97
r106 17 19 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.465 $Y=0.805
+ $X2=2.465 $Y2=0.485
r107 15 41 18.5736 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.21 $Y=1.135
+ $X2=2.21 $Y2=0.97
r108 15 16 351.245 $w=1.5e-07 $l=6.85e-07 $layer=POLY_cond $X=2.21 $Y=1.135
+ $X2=2.21 $Y2=1.82
r109 12 41 17.1559 $w=2.95e-07 $l=2.11069e-07 $layer=POLY_cond $X=2.105 $Y=0.805
+ $X2=2.21 $Y2=0.97
r110 12 14 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.105 $Y=0.805
+ $X2=2.105 $Y2=0.485
r111 10 16 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.135 $Y=1.895
+ $X2=2.21 $Y2=1.82
r112 10 11 176.904 $w=1.5e-07 $l=3.45e-07 $layer=POLY_cond $X=2.135 $Y=1.895
+ $X2=1.79 $Y2=1.895
r113 7 11 29.1797 $w=1.5e-07 $l=1.58114e-07 $layer=POLY_cond $X=1.665 $Y=1.97
+ $X2=1.79 $Y2=1.895
r114 7 9 110.86 $w=2.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.665 $Y=1.97
+ $X2=1.665 $Y2=2.545
r115 2 28 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=3.41
+ $Y=2.095 $X2=3.55 $Y2=2.24
r116 1 24 182 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_NDIFF $count=1 $X=3.33
+ $Y=0.275 $X2=3.47 $Y2=0.49
.ends

.subckt PM_SKY130_FD_SC_LP__A21BO_LP%B1_N 3 7 11 13 14 20 21
c42 21 0 1.08855e-19 $X=3.255 $Y=1.292
r43 21 22 4.78808 $w=3.02e-07 $l=3e-08 $layer=POLY_cond $X=3.255 $Y=1.292
+ $X2=3.285 $Y2=1.292
r44 19 21 13.5662 $w=3.02e-07 $l=8.5e-08 $layer=POLY_cond $X=3.17 $Y=1.292
+ $X2=3.255 $Y2=1.292
r45 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.17
+ $Y=1.2 $X2=3.17 $Y2=1.2
r46 13 14 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=3.17 $Y=1.295
+ $X2=3.17 $Y2=1.665
r47 13 20 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=3.17 $Y=1.295
+ $X2=3.17 $Y2=1.2
r48 9 21 19.1248 $w=1.5e-07 $l=2.57e-07 $layer=POLY_cond $X=3.255 $Y=1.035
+ $X2=3.255 $Y2=1.292
r49 9 11 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=3.255 $Y=1.035
+ $X2=3.255 $Y2=0.485
r50 5 22 7.29241 $w=2.5e-07 $l=2.58e-07 $layer=POLY_cond $X=3.285 $Y=1.55
+ $X2=3.285 $Y2=1.292
r51 5 7 259.634 $w=2.5e-07 $l=1.045e-06 $layer=POLY_cond $X=3.285 $Y=1.55
+ $X2=3.285 $Y2=2.595
r52 1 19 43.8907 $w=3.02e-07 $l=3.82492e-07 $layer=POLY_cond $X=2.895 $Y=1.035
+ $X2=3.17 $Y2=1.292
r53 1 3 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=2.895 $Y=1.035
+ $X2=2.895 $Y2=0.485
.ends

.subckt PM_SKY130_FD_SC_LP__A21BO_LP%X 1 2 11 14 15 16
r26 16 22 10.4468 $w=3.53e-07 $l=2.25e-07 $layer=LI1_cond $X=0.267 $Y=0.49
+ $X2=0.267 $Y2=0.715
r27 15 22 85.4652 $w=1.68e-07 $l=1.31e-06 $layer=LI1_cond $X=0.175 $Y=2.025
+ $X2=0.175 $Y2=0.715
r28 14 15 8.6688 $w=4.03e-07 $l=1.65e-07 $layer=LI1_cond $X=0.292 $Y=2.19
+ $X2=0.292 $Y2=2.025
r29 9 14 1.05285 $w=4.03e-07 $l=3.7e-08 $layer=LI1_cond $X=0.292 $Y=2.227
+ $X2=0.292 $Y2=2.19
r30 9 11 19.1505 $w=4.03e-07 $l=6.73e-07 $layer=LI1_cond $X=0.292 $Y=2.227
+ $X2=0.292 $Y2=2.9
r31 2 14 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.185
+ $Y=2.045 $X2=0.33 $Y2=2.19
r32 2 11 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.185
+ $Y=2.045 $X2=0.33 $Y2=2.9
r33 1 16 182 $w=1.7e-07 $l=2.78209e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.275 $X2=0.28 $Y2=0.49
.ends

.subckt PM_SKY130_FD_SC_LP__A21BO_LP%VPWR 1 2 11 15 18 19 20 30 31 34
r44 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r45 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r46 28 31 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r47 27 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r48 25 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r49 24 27 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r50 24 25 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r51 22 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.025 $Y=3.33
+ $X2=0.86 $Y2=3.33
r52 22 24 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=1.025 $Y=3.33
+ $X2=1.2 $Y2=3.33
r53 20 28 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=2.64 $Y2=3.33
r54 20 25 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=1.2 $Y2=3.33
r55 18 27 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=2.855 $Y=3.33
+ $X2=2.64 $Y2=3.33
r56 18 19 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.855 $Y=3.33
+ $X2=3.02 $Y2=3.33
r57 17 30 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=3.185 $Y=3.33
+ $X2=3.6 $Y2=3.33
r58 17 19 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.185 $Y=3.33
+ $X2=3.02 $Y2=3.33
r59 13 19 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.02 $Y=3.245
+ $X2=3.02 $Y2=3.33
r60 13 15 33.7002 $w=3.28e-07 $l=9.65e-07 $layer=LI1_cond $X=3.02 $Y=3.245
+ $X2=3.02 $Y2=2.28
r61 9 34 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.86 $Y=3.245 $X2=0.86
+ $Y2=3.33
r62 9 11 26.8903 $w=3.28e-07 $l=7.7e-07 $layer=LI1_cond $X=0.86 $Y=3.245
+ $X2=0.86 $Y2=2.475
r63 2 15 300 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_PDIFF $count=2 $X=2.88
+ $Y=2.095 $X2=3.02 $Y2=2.28
r64 1 11 300 $w=1.7e-07 $l=4.95076e-07 $layer=licon1_PDIFF $count=2 $X=0.72
+ $Y=2.045 $X2=0.86 $Y2=2.475
.ends

.subckt PM_SKY130_FD_SC_LP__A21BO_LP%A_252_409# 1 2 9 11 12 15
c31 12 0 5.03348e-20 $X=1.565 $Y=2.98
c32 9 0 1.64305e-19 $X=1.4 $Y=2.475
r33 13 15 21.4773 $w=3.28e-07 $l=6.15e-07 $layer=LI1_cond $X=2.49 $Y=2.895
+ $X2=2.49 $Y2=2.28
r34 11 13 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.325 $Y=2.98
+ $X2=2.49 $Y2=2.895
r35 11 12 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=2.325 $Y=2.98
+ $X2=1.565 $Y2=2.98
r36 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.4 $Y=2.895
+ $X2=1.565 $Y2=2.98
r37 7 9 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=1.4 $Y=2.895 $X2=1.4
+ $Y2=2.475
r38 2 15 300 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_PDIFF $count=2 $X=2.345
+ $Y=2.095 $X2=2.49 $Y2=2.28
r39 1 9 300 $w=1.7e-07 $l=4.95076e-07 $layer=licon1_PDIFF $count=2 $X=1.26
+ $Y=2.045 $X2=1.4 $Y2=2.475
.ends

.subckt PM_SKY130_FD_SC_LP__A21BO_LP%VGND 1 2 9 13 15 17 22 29 30 33 36
c52 9 0 1.57471e-19 $X=1.07 $Y=0.485
r53 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r54 33 34 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r55 30 37 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=2.64
+ $Y2=0
r56 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r57 27 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.845 $Y=0 $X2=2.68
+ $Y2=0
r58 27 29 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=2.845 $Y=0 $X2=3.6
+ $Y2=0
r59 26 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r60 25 26 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r61 23 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.235 $Y=0 $X2=1.07
+ $Y2=0
r62 23 25 60.3476 $w=1.68e-07 $l=9.25e-07 $layer=LI1_cond $X=1.235 $Y=0 $X2=2.16
+ $Y2=0
r63 22 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.515 $Y=0 $X2=2.68
+ $Y2=0
r64 22 25 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=2.515 $Y=0 $X2=2.16
+ $Y2=0
r65 20 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r66 19 20 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r67 17 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.905 $Y=0 $X2=1.07
+ $Y2=0
r68 17 19 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=0.905 $Y=0 $X2=0.72
+ $Y2=0
r69 15 26 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=2.16
+ $Y2=0
r70 15 34 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=1.2
+ $Y2=0
r71 11 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.68 $Y=0.085
+ $X2=2.68 $Y2=0
r72 11 13 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=2.68 $Y=0.085
+ $X2=2.68 $Y2=0.42
r73 7 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.07 $Y=0.085 $X2=1.07
+ $Y2=0
r74 7 9 13.969 $w=3.28e-07 $l=4e-07 $layer=LI1_cond $X=1.07 $Y=0.085 $X2=1.07
+ $Y2=0.485
r75 2 13 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=2.54
+ $Y=0.275 $X2=2.68 $Y2=0.42
r76 1 9 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.93
+ $Y=0.275 $X2=1.07 $Y2=0.485
.ends

