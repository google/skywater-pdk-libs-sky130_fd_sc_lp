* NGSPICE file created from sky130_fd_sc_lp__and3b_4.ext - technology: sky130A

.subckt sky130_fd_sc_lp__and3b_4 A_N B C VGND VNB VPB VPWR X
M1000 X a_242_23# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=7.056e+11p pd=6.16e+06u as=1.7808e+12p ps=1.326e+07u
M1001 a_242_23# C VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=6.867e+11p pd=6.13e+06u as=0p ps=0u
M1002 X a_242_23# VGND VNB nshort w=840000u l=150000u
+  ad=4.704e+11p pd=4.48e+06u as=9.261e+11p ps=7.51e+06u
M1003 X a_242_23# VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_717_49# B a_645_49# VNB nshort w=840000u l=150000u
+  ad=3.276e+11p pd=2.46e+06u as=1.764e+11p ps=2.1e+06u
M1005 VPWR B a_242_23# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 X a_242_23# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_242_23# a_49_133# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND a_242_23# X VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR A_N a_49_133# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1010 a_242_23# a_49_133# a_717_49# VNB nshort w=840000u l=150000u
+  ad=2.226e+11p pd=2.21e+06u as=0p ps=0u
M1011 a_645_49# C VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VGND a_242_23# X VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VPWR a_242_23# X VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VPWR a_242_23# X VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VGND A_N a_49_133# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
.ends

