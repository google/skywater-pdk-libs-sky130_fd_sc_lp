* File: sky130_fd_sc_lp__einvn_1.spice
* Created: Wed Sep  2 09:51:32 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__einvn_1.pex.spice"
.subckt sky130_fd_sc_lp__einvn_1  VNB VPB A TE_B Z VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Z	Z
* TE_B	TE_B
* A	A
* VPB	VPB
* VNB	VNB
MM1000 A_166_73# N_A_M1000_g N_Z_M1000_s VNB NSHORT L=0.15 W=0.84 AD=0.1008
+ AS=0.2226 PD=1.08 PS=2.21 NRD=9.276 NRS=0 M=1 R=5.6 SA=75000.2 SB=75000.9
+ A=0.126 P=1.98 MULT=1
MM1001 N_VGND_M1001_d N_A_214_21#_M1001_g A_166_73# VNB NSHORT L=0.15 W=0.84
+ AD=0.2604 AS=0.1008 PD=1.96667 PS=1.08 NRD=12.372 NRS=9.276 M=1 R=5.6
+ SA=75000.6 SB=75000.5 A=0.126 P=1.98 MULT=1
MM1002 N_A_214_21#_M1002_d N_TE_B_M1002_g N_VGND_M1001_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1113 AS=0.1302 PD=1.37 PS=0.983333 NRD=0 NRS=37.14 M=1 R=2.8
+ SA=75001 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1004 A_166_367# N_A_M1004_g N_Z_M1004_s VPB PHIGHVT L=0.15 W=1.26 AD=0.1512
+ AS=0.3339 PD=1.5 PS=3.05 NRD=10.1455 NRS=0 M=1 R=8.4 SA=75000.2 SB=75000.9
+ A=0.189 P=2.82 MULT=1
MM1005 N_VPWR_M1005_d N_TE_B_M1005_g A_166_367# VPB PHIGHVT L=0.15 W=1.26
+ AD=0.330551 AS=0.1512 PD=2.27463 PS=1.5 NRD=13.2778 NRS=10.1455 M=1 R=8.4
+ SA=75000.6 SB=75000.5 A=0.189 P=2.82 MULT=1
MM1003 N_A_214_21#_M1003_d N_TE_B_M1003_g N_VPWR_M1005_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1696 AS=0.167899 PD=1.81 PS=1.15537 NRD=0 NRS=15.3857 M=1
+ R=4.26667 SA=75001.2 SB=75000.2 A=0.096 P=1.58 MULT=1
DX6_noxref VNB VPB NWDIODE A=5.1847 P=9.29
*
.include "sky130_fd_sc_lp__einvn_1.pxi.spice"
*
.ends
*
*
