* File: sky130_fd_sc_lp__o21ba_2.pex.spice
* Created: Wed Sep  2 10:16:50 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O21BA_2%B1_N 3 7 9 10 14
c29 9 0 7.43928e-20 $X=0.72 $Y=1.295
r30 14 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.555 $Y=1.375
+ $X2=0.555 $Y2=1.54
r31 14 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.555 $Y=1.375
+ $X2=0.555 $Y2=1.21
r32 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.555
+ $Y=1.375 $X2=0.555 $Y2=1.375
r33 10 15 7.62336 $w=4.53e-07 $l=2.9e-07 $layer=LI1_cond $X=0.667 $Y=1.665
+ $X2=0.667 $Y2=1.375
r34 9 15 2.10299 $w=4.53e-07 $l=8e-08 $layer=LI1_cond $X=0.667 $Y=1.295
+ $X2=0.667 $Y2=1.375
r35 7 17 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=0.645 $Y=2.045
+ $X2=0.645 $Y2=1.54
r36 3 16 176.904 $w=1.5e-07 $l=3.45e-07 $layer=POLY_cond $X=0.48 $Y=0.865
+ $X2=0.48 $Y2=1.21
.ends

.subckt PM_SKY130_FD_SC_LP__O21BA_2%A_186_21# 1 2 7 9 10 12 13 15 16 18 21 24 25
+ 28 32 39 41 47
c77 25 0 1.77193e-19 $X=1.795 $Y=1.09
c78 21 0 9.68575e-20 $X=1.63 $Y=1.35
c79 10 0 7.43928e-20 $X=1.29 $Y=1.725
r80 44 45 14.3665 $w=5.4e-07 $l=1.45e-07 $layer=POLY_cond $X=1.29 $Y=1.455
+ $X2=1.435 $Y2=1.455
r81 42 44 28.2377 $w=5.4e-07 $l=2.85e-07 $layer=POLY_cond $X=1.005 $Y=1.455
+ $X2=1.29 $Y2=1.455
r82 36 39 0.364908 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.525 $Y=1.175
+ $X2=2.525 $Y2=1.09
r83 36 41 41.899 $w=1.78e-07 $l=6.8e-07 $layer=LI1_cond $X=2.525 $Y=1.175
+ $X2=2.525 $Y2=1.855
r84 32 34 47.0043 $w=2.08e-07 $l=8.9e-07 $layer=LI1_cond $X=2.51 $Y=2.02
+ $X2=2.51 $Y2=2.91
r85 30 41 5.80296 $w=2.08e-07 $l=1.05e-07 $layer=LI1_cond $X=2.51 $Y=1.96
+ $X2=2.51 $Y2=1.855
r86 30 32 3.16883 $w=2.08e-07 $l=6e-08 $layer=LI1_cond $X=2.51 $Y=1.96 $X2=2.51
+ $Y2=2.02
r87 26 39 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=2.135 $Y=1.09
+ $X2=2.525 $Y2=1.09
r88 26 28 25.93 $w=2.58e-07 $l=5.85e-07 $layer=LI1_cond $X=2.135 $Y=1.005
+ $X2=2.135 $Y2=0.42
r89 24 26 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=2.005 $Y=1.09
+ $X2=2.135 $Y2=1.09
r90 24 25 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=2.005 $Y=1.09
+ $X2=1.795 $Y2=1.09
r91 22 47 8.91716 $w=5.4e-07 $l=9e-08 $layer=POLY_cond $X=1.63 $Y=1.455 $X2=1.72
+ $Y2=1.455
r92 22 45 19.3205 $w=5.4e-07 $l=1.95e-07 $layer=POLY_cond $X=1.63 $Y=1.455
+ $X2=1.435 $Y2=1.455
r93 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.63
+ $Y=1.35 $X2=1.63 $Y2=1.35
r94 19 25 7.59919 $w=1.7e-07 $l=1.92873e-07 $layer=LI1_cond $X=1.64 $Y=1.175
+ $X2=1.795 $Y2=1.09
r95 19 21 6.50573 $w=3.08e-07 $l=1.75e-07 $layer=LI1_cond $X=1.64 $Y=1.175
+ $X2=1.64 $Y2=1.35
r96 16 47 33.3633 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=1.72 $Y=1.725
+ $X2=1.72 $Y2=1.455
r97 16 18 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=1.72 $Y=1.725
+ $X2=1.72 $Y2=2.465
r98 13 45 33.3633 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=1.435 $Y=1.185
+ $X2=1.435 $Y2=1.455
r99 13 15 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.435 $Y=1.185
+ $X2=1.435 $Y2=0.655
r100 10 44 33.3633 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=1.29 $Y=1.725
+ $X2=1.29 $Y2=1.455
r101 10 12 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=1.29 $Y=1.725
+ $X2=1.29 $Y2=2.465
r102 7 42 33.3633 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=1.005 $Y=1.185
+ $X2=1.005 $Y2=1.455
r103 7 9 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.005 $Y=1.185
+ $X2=1.005 $Y2=0.655
r104 2 34 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=2.38
+ $Y=1.835 $X2=2.52 $Y2=2.91
r105 2 32 400 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_PDIFF $count=1 $X=2.38
+ $Y=1.835 $X2=2.52 $Y2=2.02
r106 1 28 91 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=2 $X=2.045
+ $Y=0.235 $X2=2.17 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__O21BA_2%A_28_131# 1 2 9 13 17 20 22 26 27 31 36
r67 32 36 21.8356 $w=2.98e-07 $l=1.35e-07 $layer=POLY_cond $X=2.17 $Y=1.51
+ $X2=2.305 $Y2=1.51
r68 31 34 7.49534 $w=2.58e-07 $l=1.65e-07 $layer=LI1_cond $X=2.135 $Y=1.51
+ $X2=2.135 $Y2=1.675
r69 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.17
+ $Y=1.51 $X2=2.17 $Y2=1.51
r70 26 28 6.80123 $w=5.08e-07 $l=2.9e-07 $layer=LI1_cond $X=0.34 $Y=2.085
+ $X2=0.34 $Y2=2.375
r71 26 27 8.98828 $w=5.08e-07 $l=1.65e-07 $layer=LI1_cond $X=0.34 $Y=2.085
+ $X2=0.34 $Y2=1.92
r72 24 27 53.3563 $w=1.83e-07 $l=8.9e-07 $layer=LI1_cond $X=0.177 $Y=1.03
+ $X2=0.177 $Y2=1.92
r73 22 24 8.15385 $w=2.73e-07 $l=1.65e-07 $layer=LI1_cond $X=0.222 $Y=0.865
+ $X2=0.222 $Y2=1.03
r74 20 34 30.8153 $w=2.28e-07 $l=6.15e-07 $layer=LI1_cond $X=2.12 $Y=2.29
+ $X2=2.12 $Y2=1.675
r75 18 28 7.28118 $w=1.7e-07 $l=2.55e-07 $layer=LI1_cond $X=0.595 $Y=2.375
+ $X2=0.34 $Y2=2.375
r76 17 20 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=2.005 $Y=2.375
+ $X2=2.12 $Y2=2.29
r77 17 18 91.9893 $w=1.68e-07 $l=1.41e-06 $layer=LI1_cond $X=2.005 $Y=2.375
+ $X2=0.595 $Y2=2.375
r78 11 36 12.9396 $w=2.98e-07 $l=2.0106e-07 $layer=POLY_cond $X=2.385 $Y=1.345
+ $X2=2.305 $Y2=1.51
r79 11 13 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.385 $Y=1.345
+ $X2=2.385 $Y2=0.655
r80 7 36 18.8112 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.305 $Y=1.675
+ $X2=2.305 $Y2=1.51
r81 7 9 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.305 $Y=1.675
+ $X2=2.305 $Y2=2.465
r82 2 26 600 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_PDIFF $count=1 $X=0.305
+ $Y=1.835 $X2=0.43 $Y2=2.085
r83 1 22 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.14
+ $Y=0.655 $X2=0.265 $Y2=0.865
.ends

.subckt PM_SKY130_FD_SC_LP__O21BA_2%A2 3 7 9 10 11 12 18
c37 3 0 1.32777e-19 $X=2.745 $Y=2.465
r38 18 21 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=2.852 $Y=1.375
+ $X2=2.852 $Y2=1.54
r39 18 20 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=2.852 $Y=1.375
+ $X2=2.852 $Y2=1.21
r40 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.87
+ $Y=1.375 $X2=2.87 $Y2=1.375
r41 11 12 9.91637 $w=4.28e-07 $l=3.7e-07 $layer=LI1_cond $X=3 $Y=2.035 $X2=3
+ $Y2=2.405
r42 10 11 9.91637 $w=4.28e-07 $l=3.7e-07 $layer=LI1_cond $X=3 $Y=1.665 $X2=3
+ $Y2=2.035
r43 10 19 7.77229 $w=4.28e-07 $l=2.9e-07 $layer=LI1_cond $X=3 $Y=1.665 $X2=3
+ $Y2=1.375
r44 9 19 2.14408 $w=4.28e-07 $l=8e-08 $layer=LI1_cond $X=3 $Y=1.295 $X2=3
+ $Y2=1.375
r45 7 20 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=2.815 $Y=0.655
+ $X2=2.815 $Y2=1.21
r46 3 21 474.309 $w=1.5e-07 $l=9.25e-07 $layer=POLY_cond $X=2.745 $Y=2.465
+ $X2=2.745 $Y2=1.54
.ends

.subckt PM_SKY130_FD_SC_LP__O21BA_2%A1 3 7 9 10 14
c25 9 0 1.32777e-19 $X=3.6 $Y=1.295
r26 14 17 45.456 $w=3.9e-07 $l=1.65e-07 $layer=POLY_cond $X=3.44 $Y=1.375
+ $X2=3.44 $Y2=1.54
r27 14 16 45.456 $w=3.9e-07 $l=1.65e-07 $layer=POLY_cond $X=3.44 $Y=1.375
+ $X2=3.44 $Y2=1.21
r28 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.47
+ $Y=1.375 $X2=3.47 $Y2=1.375
r29 10 15 9.03266 $w=3.68e-07 $l=2.9e-07 $layer=LI1_cond $X=3.57 $Y=1.665
+ $X2=3.57 $Y2=1.375
r30 9 15 2.49177 $w=3.68e-07 $l=8e-08 $layer=LI1_cond $X=3.57 $Y=1.295 $X2=3.57
+ $Y2=1.375
r31 7 16 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=3.325 $Y=0.655
+ $X2=3.325 $Y2=1.21
r32 3 17 474.309 $w=1.5e-07 $l=9.25e-07 $layer=POLY_cond $X=3.32 $Y=2.465
+ $X2=3.32 $Y2=1.54
.ends

.subckt PM_SKY130_FD_SC_LP__O21BA_2%VPWR 1 2 3 12 16 18 20 25 26 27 33 37 43 47
c42 1 0 1.96412e-19 $X=0.72 $Y=1.835
r43 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r44 43 44 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r45 41 47 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r46 41 44 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.16 $Y2=3.33
r47 40 41 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r48 38 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.17 $Y=3.33
+ $X2=2.005 $Y2=3.33
r49 38 40 61.9786 $w=1.68e-07 $l=9.5e-07 $layer=LI1_cond $X=2.17 $Y=3.33
+ $X2=3.12 $Y2=3.33
r50 37 46 4.54029 $w=1.7e-07 $l=2.27e-07 $layer=LI1_cond $X=3.385 $Y=3.33
+ $X2=3.612 $Y2=3.33
r51 37 40 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=3.385 $Y=3.33
+ $X2=3.12 $Y2=3.33
r52 35 36 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r53 33 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.84 $Y=3.33
+ $X2=2.005 $Y2=3.33
r54 33 35 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=1.84 $Y=3.33
+ $X2=1.68 $Y2=3.33
r55 31 36 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r56 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r57 27 44 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=2.16 $Y2=3.33
r58 27 36 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=1.68 $Y2=3.33
r59 25 30 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=0.91 $Y=3.33
+ $X2=0.72 $Y2=3.33
r60 25 26 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.91 $Y=3.33
+ $X2=1.075 $Y2=3.33
r61 24 35 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=1.24 $Y=3.33
+ $X2=1.68 $Y2=3.33
r62 24 26 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.24 $Y=3.33
+ $X2=1.075 $Y2=3.33
r63 20 23 31.6465 $w=3.13e-07 $l=8.65e-07 $layer=LI1_cond $X=3.542 $Y=2.085
+ $X2=3.542 $Y2=2.95
r64 18 46 3.1002 $w=3.15e-07 $l=1.14782e-07 $layer=LI1_cond $X=3.542 $Y=3.245
+ $X2=3.612 $Y2=3.33
r65 18 23 10.7927 $w=3.13e-07 $l=2.95e-07 $layer=LI1_cond $X=3.542 $Y=3.245
+ $X2=3.542 $Y2=2.95
r66 14 43 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.005 $Y=3.245
+ $X2=2.005 $Y2=3.33
r67 14 16 17.112 $w=3.28e-07 $l=4.9e-07 $layer=LI1_cond $X=2.005 $Y=3.245
+ $X2=2.005 $Y2=2.755
r68 10 26 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.075 $Y=3.245
+ $X2=1.075 $Y2=3.33
r69 10 12 17.112 $w=3.28e-07 $l=4.9e-07 $layer=LI1_cond $X=1.075 $Y=3.245
+ $X2=1.075 $Y2=2.755
r70 3 23 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=3.395
+ $Y=1.835 $X2=3.535 $Y2=2.95
r71 3 20 400 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_PDIFF $count=1 $X=3.395
+ $Y=1.835 $X2=3.535 $Y2=2.085
r72 2 16 600 $w=1.7e-07 $l=1.01961e-06 $layer=licon1_PDIFF $count=1 $X=1.795
+ $Y=1.835 $X2=2.005 $Y2=2.755
r73 1 12 600 $w=1.7e-07 $l=1.08305e-06 $layer=licon1_PDIFF $count=1 $X=0.72
+ $Y=1.835 $X2=1.075 $Y2=2.755
.ends

.subckt PM_SKY130_FD_SC_LP__O21BA_2%X 1 2 9 11 12 13 14 15 21 23
c31 23 0 1.96412e-19 $X=1.22 $Y=0.42
r32 15 21 3.54615 $w=2.5e-07 $l=1.35e-07 $layer=LI1_cond $X=1.19 $Y=1.985
+ $X2=1.19 $Y2=1.85
r33 14 21 8.52808 $w=2.48e-07 $l=1.85e-07 $layer=LI1_cond $X=1.19 $Y=1.665
+ $X2=1.19 $Y2=1.85
r34 13 14 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=1.19 $Y=1.295
+ $X2=1.19 $Y2=1.665
r35 12 13 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=1.19 $Y=0.925
+ $X2=1.19 $Y2=1.295
r36 11 12 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=1.19 $Y=0.555
+ $X2=1.19 $Y2=0.925
r37 11 23 6.22319 $w=2.48e-07 $l=1.35e-07 $layer=LI1_cond $X=1.19 $Y=0.555
+ $X2=1.19 $Y2=0.42
r38 7 15 3.28347 $w=2.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.315 $Y=1.985
+ $X2=1.19 $Y2=1.985
r39 7 9 8.10978 $w=2.68e-07 $l=1.9e-07 $layer=LI1_cond $X=1.315 $Y=1.985
+ $X2=1.505 $Y2=1.985
r40 2 9 600 $w=1.7e-07 $l=2.4e-07 $layer=licon1_PDIFF $count=1 $X=1.365 $Y=1.835
+ $X2=1.505 $Y2=2.015
r41 1 23 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=1.08
+ $Y=0.235 $X2=1.22 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__O21BA_2%VGND 1 2 3 12 18 22 24 26 31 36 43 44 47 50
+ 53
r59 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r60 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r61 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r62 44 54 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=3.12
+ $Y2=0
r63 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r64 41 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.265 $Y=0 $X2=3.1
+ $Y2=0
r65 41 43 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=3.265 $Y=0 $X2=3.6
+ $Y2=0
r66 40 54 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r67 39 40 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r68 37 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.815 $Y=0 $X2=1.65
+ $Y2=0
r69 37 39 53.8235 $w=1.68e-07 $l=8.25e-07 $layer=LI1_cond $X=1.815 $Y=0 $X2=2.64
+ $Y2=0
r70 36 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.935 $Y=0 $X2=3.1
+ $Y2=0
r71 36 39 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=2.935 $Y=0 $X2=2.64
+ $Y2=0
r72 35 51 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r73 35 48 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r74 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r75 32 47 9.23004 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=0.895 $Y=0 $X2=0.712
+ $Y2=0
r76 32 34 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.895 $Y=0 $X2=1.2
+ $Y2=0
r77 31 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.485 $Y=0 $X2=1.65
+ $Y2=0
r78 31 34 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.485 $Y=0 $X2=1.2
+ $Y2=0
r79 29 48 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r80 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r81 26 47 9.23004 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=0.53 $Y=0 $X2=0.712
+ $Y2=0
r82 26 28 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=0.53 $Y=0 $X2=0.24
+ $Y2=0
r83 24 40 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=2.64
+ $Y2=0
r84 24 51 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=1.68
+ $Y2=0
r85 20 53 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.1 $Y=0.085 $X2=3.1
+ $Y2=0
r86 20 22 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=3.1 $Y=0.085
+ $X2=3.1 $Y2=0.38
r87 16 50 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.65 $Y=0.085
+ $X2=1.65 $Y2=0
r88 16 18 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.65 $Y=0.085
+ $X2=1.65 $Y2=0.38
r89 12 14 15.629 $w=3.63e-07 $l=4.95e-07 $layer=LI1_cond $X=0.712 $Y=0.38
+ $X2=0.712 $Y2=0.875
r90 10 47 1.2012 $w=3.65e-07 $l=8.5e-08 $layer=LI1_cond $X=0.712 $Y=0.085
+ $X2=0.712 $Y2=0
r91 10 12 9.31427 $w=3.63e-07 $l=2.95e-07 $layer=LI1_cond $X=0.712 $Y=0.085
+ $X2=0.712 $Y2=0.38
r92 3 22 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=2.89
+ $Y=0.235 $X2=3.1 $Y2=0.38
r93 2 18 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.51
+ $Y=0.235 $X2=1.65 $Y2=0.38
r94 1 14 182 $w=1.7e-07 $l=2.81425e-07 $layer=licon1_NDIFF $count=1 $X=0.555
+ $Y=0.655 $X2=0.695 $Y2=0.875
r95 1 12 182 $w=1.7e-07 $l=3.745e-07 $layer=licon1_NDIFF $count=1 $X=0.555
+ $Y=0.655 $X2=0.79 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_LP__O21BA_2%A_492_47# 1 2 9 11 12 15 17
r31 17 20 6.46067 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=3.54 $Y=0.745
+ $X2=3.54 $Y2=0.93
r32 17 18 3.55804 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=3.54 $Y=0.745 $X2=3.54
+ $Y2=0.655
r33 15 18 10.0305 $w=2.68e-07 $l=2.35e-07 $layer=LI1_cond $X=3.57 $Y=0.42
+ $X2=3.57 $Y2=0.655
r34 11 17 4.28565 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=3.375 $Y=0.745
+ $X2=3.54 $Y2=0.745
r35 11 12 37.5859 $w=1.78e-07 $l=6.1e-07 $layer=LI1_cond $X=3.375 $Y=0.745
+ $X2=2.765 $Y2=0.745
r36 7 12 7.61292 $w=1.8e-07 $l=2.05122e-07 $layer=LI1_cond $X=2.6 $Y=0.655
+ $X2=2.765 $Y2=0.745
r37 7 9 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=2.6 $Y=0.655 $X2=2.6
+ $Y2=0.37
r38 2 20 182 $w=1.7e-07 $l=7.61791e-07 $layer=licon1_NDIFF $count=1 $X=3.4
+ $Y=0.235 $X2=3.54 $Y2=0.93
r39 2 15 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=3.4
+ $Y=0.235 $X2=3.54 $Y2=0.42
r40 1 9 91 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_NDIFF $count=2 $X=2.46
+ $Y=0.235 $X2=2.6 $Y2=0.37
.ends

