* File: sky130_fd_sc_lp__nand2_m.spice
* Created: Wed Sep  2 10:03:19 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__nand2_m.pex.spice"
.subckt sky130_fd_sc_lp__nand2_m  VNB VPB B A VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A	A
* B	B
* VPB	VPB
* VNB	VNB
MM1003 A_124_47# N_B_M1003_g N_VGND_M1003_s VNB NSHORT L=0.15 W=0.42 AD=0.0504
+ AS=0.1113 PD=0.66 PS=1.37 NRD=18.564 NRS=0 M=1 R=2.8 SA=75000.2 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1001 N_Y_M1001_d N_A_M1001_g A_124_47# VNB NSHORT L=0.15 W=0.42 AD=0.1113
+ AS=0.0504 PD=1.37 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75000.6 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1000 N_Y_M1000_d N_B_M1000_g N_VPWR_M1000_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1002 N_VPWR_M1002_d N_A_M1002_g N_Y_M1000_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6 SB=75000.2
+ A=0.063 P=1.14 MULT=1
DX4_noxref VNB VPB NWDIODE A=3.3943 P=7.37
*
.include "sky130_fd_sc_lp__nand2_m.pxi.spice"
*
.ends
*
*
