# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__busdrivernovlp_20
  CLASS CORE ;
  FOREIGN sky130_fd_sc_lp__busdrivernovlp_20 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  17.76000 BY  3.330000 ;
  SYMMETRY X Y ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.925000 1.345000 5.255000 1.675000 ;
        RECT 4.925000 1.675000 5.155000 2.150000 ;
    END
  END A
  PIN TE_B
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.505000 0.995000 1.740000 1.165000 ;
        RECT 0.505000 1.165000 0.835000 1.410000 ;
        RECT 1.570000 0.265000 2.805000 0.435000 ;
        RECT 1.570000 0.435000 1.740000 0.995000 ;
        RECT 2.475000 0.435000 2.805000 0.850000 ;
        RECT 2.475000 0.850000 3.505000 1.020000 ;
        RECT 3.335000 0.265000 4.205000 0.435000 ;
        RECT 3.335000 0.435000 3.505000 0.850000 ;
        RECT 4.035000 0.435000 4.205000 0.645000 ;
        RECT 4.035000 0.645000 5.985000 0.815000 ;
        RECT 5.815000 0.815000 5.985000 0.995000 ;
        RECT 5.815000 0.995000 6.215000 1.325000 ;
    END
  END TE_B
  PIN Z
    ANTENNADIFFAREA  4.968000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 9.160000 1.920000 17.190000 2.150000 ;
    END
  END Z
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 17.760000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 17.760000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 17.760000 0.085000 ;
      RECT  0.000000  3.245000 17.760000 3.415000 ;
      RECT  0.100000  0.645000  0.880000 0.815000 ;
      RECT  0.100000  0.815000  0.270000 1.590000 ;
      RECT  0.100000  1.590000  1.415000 1.760000 ;
      RECT  0.100000  1.760000  0.430000 2.695000 ;
      RECT  0.550000  0.405000  0.880000 0.645000 ;
      RECT  0.630000  1.940000  0.880000 3.245000 ;
      RECT  1.060000  0.085000  1.390000 0.815000 ;
      RECT  1.060000  1.940000  1.765000 2.110000 ;
      RECT  1.060000  2.110000  1.390000 3.065000 ;
      RECT  1.085000  1.345000  1.415000 1.590000 ;
      RECT  1.570000  2.290000  1.820000 3.245000 ;
      RECT  1.595000  1.550000  2.565000 1.720000 ;
      RECT  1.595000  1.720000  1.765000 1.940000 ;
      RECT  1.995000  0.615000  2.245000 1.200000 ;
      RECT  1.995000  1.200000  2.970000 1.370000 ;
      RECT  2.000000  2.085000  3.130000 2.255000 ;
      RECT  2.000000  2.255000  2.330000 3.065000 ;
      RECT  2.045000  1.720000  2.565000 1.905000 ;
      RECT  2.510000  2.435000  2.760000 3.245000 ;
      RECT  2.800000  1.370000  2.970000 1.575000 ;
      RECT  2.800000  1.575000  3.130000 2.085000 ;
      RECT  2.985000  0.085000  3.155000 0.670000 ;
      RECT  3.335000  1.815000  3.505000 2.895000 ;
      RECT  3.335000  2.895000  4.485000 3.065000 ;
      RECT  3.685000  0.615000  3.855000 0.995000 ;
      RECT  3.685000  0.995000  5.635000 1.165000 ;
      RECT  3.685000  1.165000  3.855000 1.815000 ;
      RECT  3.685000  1.815000  3.975000 2.715000 ;
      RECT  4.155000  1.815000  4.485000 2.330000 ;
      RECT  4.155000  2.330000  5.585000 2.500000 ;
      RECT  4.155000  2.500000  4.485000 2.895000 ;
      RECT  4.385000  0.085000  4.715000 0.465000 ;
      RECT  4.665000  2.680000  4.995000 3.245000 ;
      RECT  5.335000  1.855000  5.585000 2.330000 ;
      RECT  5.335000  2.500000  5.585000 3.065000 ;
      RECT  5.435000  1.165000  5.635000 1.410000 ;
      RECT  5.545000  0.085000  5.875000 0.465000 ;
      RECT  5.845000  1.845000  6.175000 3.245000 ;
      RECT  6.165000  0.265000  6.495000 0.645000 ;
      RECT  6.165000  0.645000  7.190000 0.815000 ;
      RECT  6.395000  0.995000  6.840000 1.665000 ;
      RECT  6.665000  1.845000  7.190000 2.015000 ;
      RECT  6.665000  2.015000  6.995000 2.725000 ;
      RECT  6.675000  0.085000  7.005000 0.465000 ;
      RECT  7.020000  0.815000  7.190000 1.275000 ;
      RECT  7.020000  1.275000  8.690000 1.605000 ;
      RECT  7.020000  1.605000  7.190000 1.845000 ;
      RECT  7.235000  0.295000  7.565000 0.465000 ;
      RECT  7.265000  2.185000  7.515000 3.245000 ;
      RECT  7.360000  0.465000  7.565000 0.925000 ;
      RECT  7.360000  0.925000  8.505000 1.095000 ;
      RECT  7.695000  1.785000  9.040000 1.955000 ;
      RECT  7.695000  1.955000  8.025000 3.065000 ;
      RECT  7.745000  0.085000  7.995000 0.745000 ;
      RECT  8.175000  0.265000  9.470000 0.435000 ;
      RECT  8.175000  0.435000  8.505000 0.925000 ;
      RECT  8.205000  2.135000  8.875000 3.245000 ;
      RECT  8.685000  0.615000  9.040000 1.095000 ;
      RECT  8.870000  1.095000  9.040000 1.550000 ;
      RECT  8.870000  1.550000  9.475000 1.780000 ;
      RECT  8.870000  1.780000  9.040000 1.785000 ;
      RECT  9.220000  0.435000  9.470000 1.095000 ;
      RECT  9.220000  1.950000 10.330000 2.130000 ;
      RECT  9.220000  2.130000  9.390000 3.065000 ;
      RECT  9.570000  2.310000  9.820000 3.245000 ;
      RECT  9.640000  1.035000  9.830000 1.410000 ;
      RECT 10.000000  0.255000 10.330000 1.950000 ;
      RECT 10.000000  2.130000 10.330000 3.065000 ;
      RECT 10.500000  1.035000 10.690000 1.410000 ;
      RECT 10.510000  0.085000 10.680000 0.865000 ;
      RECT 10.510000  2.290000 10.680000 3.245000 ;
      RECT 10.860000  0.255000 11.190000 3.065000 ;
      RECT 11.360000  1.035000 11.550000 1.410000 ;
      RECT 11.370000  0.085000 11.540000 0.865000 ;
      RECT 11.370000  2.290000 11.540000 3.245000 ;
      RECT 11.720000  0.255000 12.050000 3.065000 ;
      RECT 12.220000  1.035000 12.410000 1.410000 ;
      RECT 12.230000  0.085000 12.400000 0.865000 ;
      RECT 12.230000  2.290000 12.400000 3.245000 ;
      RECT 12.580000  0.255000 12.910000 3.065000 ;
      RECT 13.080000  1.035000 13.270000 1.410000 ;
      RECT 13.090000  0.085000 13.260000 0.865000 ;
      RECT 13.090000  2.290000 13.260000 3.245000 ;
      RECT 13.440000  0.255000 13.770000 3.065000 ;
      RECT 13.940000  1.345000 14.130000 1.760000 ;
      RECT 13.950000  0.085000 14.120000 0.865000 ;
      RECT 13.950000  2.290000 14.120000 3.245000 ;
      RECT 14.300000  0.255000 14.630000 3.065000 ;
      RECT 14.800000  1.345000 14.990000 1.760000 ;
      RECT 14.810000  0.085000 14.980000 0.865000 ;
      RECT 14.810000  2.290000 14.980000 3.245000 ;
      RECT 15.160000  0.260000 15.490000 3.065000 ;
      RECT 15.660000  1.345000 15.850000 1.760000 ;
      RECT 15.670000  0.085000 15.840000 0.865000 ;
      RECT 15.670000  2.290000 15.840000 3.245000 ;
      RECT 16.020000  0.255000 16.350000 3.065000 ;
      RECT 16.520000  1.345000 17.110000 1.760000 ;
      RECT 16.530000  2.290000 16.700000 3.245000 ;
      RECT 16.880000  1.940000 17.210000 3.065000 ;
      RECT 17.390000  2.290000 17.640000 3.245000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  1.580000  2.245000 1.750000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  1.210000  5.605000 1.380000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  1.210000  6.565000 1.380000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  1.580000  9.445000 1.750000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.660000  1.210000  9.830000 1.380000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.080000  1.950000 10.250000 2.120000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
      RECT 10.520000  1.210000 10.690000 1.380000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  3.245000 10.885000 3.415000 ;
      RECT 10.940000  1.950000 11.110000 2.120000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  3.245000 11.365000 3.415000 ;
      RECT 11.380000  1.210000 11.550000 1.380000 ;
      RECT 11.675000 -0.085000 11.845000 0.085000 ;
      RECT 11.675000  3.245000 11.845000 3.415000 ;
      RECT 11.800000  1.950000 11.970000 2.120000 ;
      RECT 12.155000 -0.085000 12.325000 0.085000 ;
      RECT 12.155000  3.245000 12.325000 3.415000 ;
      RECT 12.240000  1.210000 12.410000 1.380000 ;
      RECT 12.635000 -0.085000 12.805000 0.085000 ;
      RECT 12.635000  3.245000 12.805000 3.415000 ;
      RECT 12.660000  1.950000 12.830000 2.120000 ;
      RECT 13.100000  1.210000 13.270000 1.380000 ;
      RECT 13.115000 -0.085000 13.285000 0.085000 ;
      RECT 13.115000  3.245000 13.285000 3.415000 ;
      RECT 13.520000  1.950000 13.690000 2.120000 ;
      RECT 13.595000 -0.085000 13.765000 0.085000 ;
      RECT 13.595000  3.245000 13.765000 3.415000 ;
      RECT 13.940000  1.580000 14.110000 1.750000 ;
      RECT 14.075000 -0.085000 14.245000 0.085000 ;
      RECT 14.075000  3.245000 14.245000 3.415000 ;
      RECT 14.380000  1.950000 14.550000 2.120000 ;
      RECT 14.555000 -0.085000 14.725000 0.085000 ;
      RECT 14.555000  3.245000 14.725000 3.415000 ;
      RECT 14.800000  1.580000 14.970000 1.750000 ;
      RECT 15.035000 -0.085000 15.205000 0.085000 ;
      RECT 15.035000  3.245000 15.205000 3.415000 ;
      RECT 15.240000  1.950000 15.410000 2.120000 ;
      RECT 15.515000 -0.085000 15.685000 0.085000 ;
      RECT 15.515000  3.245000 15.685000 3.415000 ;
      RECT 15.660000  1.580000 15.830000 1.750000 ;
      RECT 15.995000 -0.085000 16.165000 0.085000 ;
      RECT 15.995000  3.245000 16.165000 3.415000 ;
      RECT 16.100000  1.950000 16.270000 2.120000 ;
      RECT 16.475000 -0.085000 16.645000 0.085000 ;
      RECT 16.475000  3.245000 16.645000 3.415000 ;
      RECT 16.520000  1.580000 16.690000 1.750000 ;
      RECT 16.880000  1.580000 17.050000 1.750000 ;
      RECT 16.955000 -0.085000 17.125000 0.085000 ;
      RECT 16.955000  3.245000 17.125000 3.415000 ;
      RECT 16.960000  1.950000 17.130000 2.120000 ;
      RECT 17.435000 -0.085000 17.605000 0.085000 ;
      RECT 17.435000  3.245000 17.605000 3.415000 ;
    LAYER met1 ;
      RECT 2.015000 1.550000  2.305000 1.595000 ;
      RECT 2.015000 1.595000 17.110000 1.735000 ;
      RECT 2.015000 1.735000  2.305000 1.780000 ;
      RECT 5.375000 1.180000  5.665000 1.225000 ;
      RECT 5.375000 1.225000 13.330000 1.365000 ;
      RECT 5.375000 1.365000  5.665000 1.410000 ;
      RECT 6.335000 1.180000  6.625000 1.225000 ;
      RECT 6.335000 1.365000  6.625000 1.410000 ;
      RECT 9.215000 1.550000 17.110000 1.595000 ;
      RECT 9.215000 1.735000 17.110000 1.780000 ;
      RECT 9.600000 1.180000 13.330000 1.225000 ;
      RECT 9.600000 1.365000 13.330000 1.410000 ;
  END
END sky130_fd_sc_lp__busdrivernovlp_20
END LIBRARY
