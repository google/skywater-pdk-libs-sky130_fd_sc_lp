* File: sky130_fd_sc_lp__or2_4.spice
* Created: Wed Sep  2 10:29:12 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__or2_4.pex.spice"
.subckt sky130_fd_sc_lp__or2_4  VNB VPB B A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* B	B
* VPB	VPB
* VNB	VNB
MM1003 N_A_27_367#_M1003_d N_B_M1003_g N_VGND_M1003_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1239 AS=0.2226 PD=1.135 PS=2.21 NRD=2.136 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75002.4 A=0.126 P=1.98 MULT=1
MM1008 N_VGND_M1008_d N_A_M1008_g N_A_27_367#_M1003_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1428 AS=0.1239 PD=1.18 PS=1.135 NRD=4.284 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75002 A=0.126 P=1.98 MULT=1
MM1001 N_X_M1001_d N_A_27_367#_M1001_g N_VGND_M1008_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1428 PD=1.12 PS=1.18 NRD=0 NRS=4.284 M=1 R=5.6 SA=75001.1
+ SB=75001.5 A=0.126 P=1.98 MULT=1
MM1002 N_X_M1001_d N_A_27_367#_M1002_g N_VGND_M1002_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.6
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1005 N_X_M1005_d N_A_27_367#_M1005_g N_VGND_M1002_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002 SB=75000.6
+ A=0.126 P=1.98 MULT=1
MM1007 N_X_M1005_d N_A_27_367#_M1007_g N_VGND_M1007_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75002.4
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1011 A_110_367# N_B_M1011_g N_A_27_367#_M1011_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1323 AS=0.3339 PD=1.47 PS=3.05 NRD=7.8012 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75002.4 A=0.189 P=2.82 MULT=1
MM1009 N_VPWR_M1009_d N_A_M1009_g A_110_367# VPB PHIGHVT L=0.15 W=1.26
+ AD=0.26775 AS=0.1323 PD=1.685 PS=1.47 NRD=11.7215 NRS=7.8012 M=1 R=8.4
+ SA=75000.6 SB=75002.1 A=0.189 P=2.82 MULT=1
MM1000 N_VPWR_M1009_d N_A_27_367#_M1000_g N_X_M1000_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.26775 AS=0.1764 PD=1.685 PS=1.54 NRD=10.9335 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75001.5 A=0.189 P=2.82 MULT=1
MM1004 N_VPWR_M1004_d N_A_27_367#_M1004_g N_X_M1000_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.6
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1006 N_VPWR_M1004_d N_A_27_367#_M1006_g N_X_M1006_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002 SB=75000.6
+ A=0.189 P=2.82 MULT=1
MM1010 N_VPWR_M1010_d N_A_27_367#_M1010_g N_X_M1006_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.4
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX12_noxref VNB VPB NWDIODE A=6.9751 P=11.21
*
.include "sky130_fd_sc_lp__or2_4.pxi.spice"
*
.ends
*
*
