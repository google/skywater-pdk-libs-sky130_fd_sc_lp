* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__dfstp_4 CLK D SET_B VGND VNB VPB VPWR Q
X0 VPWR a_562_119# a_690_93# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X1 a_562_119# a_30_99# a_690_463# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X2 a_690_463# a_690_93# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X3 a_30_99# CLK VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 a_648_119# a_690_93# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 a_1247_47# a_30_99# a_1356_91# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 VPWR a_30_99# a_230_465# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X7 VGND D a_476_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 a_1356_91# a_1398_65# a_1428_91# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 VPWR a_562_119# a_1094_379# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X10 a_562_119# a_230_465# a_648_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X11 a_1247_47# a_30_99# a_1094_379# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X12 VPWR a_1247_47# a_1398_65# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X13 a_1989_49# a_1247_47# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X14 Q a_1989_49# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X15 Q a_1989_49# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X16 a_1201_407# a_1398_65# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X17 VPWR a_1989_49# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X18 a_1989_49# a_1247_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X19 a_476_119# a_30_99# a_562_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X20 a_914_47# SET_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X21 a_1175_47# a_230_465# a_1247_47# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X22 VGND a_1989_49# Q VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X23 VPWR D a_476_119# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X24 Q a_1989_49# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X25 a_1428_91# SET_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X26 VGND a_1989_49# Q VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X27 VPWR SET_B a_1247_47# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X28 Q a_1989_49# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X29 VGND a_1247_47# a_1398_65# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X30 a_1201_407# a_230_465# a_1247_47# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X31 VGND a_30_99# a_230_465# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X32 a_476_119# a_230_465# a_562_119# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X33 a_690_93# a_562_119# a_914_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X34 VGND a_562_119# a_1175_47# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X35 a_30_99# CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X36 VPWR a_1989_49# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X37 a_690_93# SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
.ends
