* File: sky130_fd_sc_lp__nand2b_lp.pxi.spice
* Created: Fri Aug 28 10:48:31 2020
* 
x_PM_SKY130_FD_SC_LP__NAND2B_LP%A_N N_A_N_c_52_n N_A_N_M1000_g N_A_N_c_53_n
+ N_A_N_M1003_g N_A_N_c_54_n N_A_N_c_55_n N_A_N_M1005_g N_A_N_c_56_n
+ N_A_N_c_62_n A_N N_A_N_c_57_n N_A_N_c_58_n N_A_N_c_59_n
+ PM_SKY130_FD_SC_LP__NAND2B_LP%A_N
x_PM_SKY130_FD_SC_LP__NAND2B_LP%B N_B_c_105_n N_B_M1006_g N_B_M1001_g
+ N_B_c_102_n B N_B_c_103_n N_B_c_104_n PM_SKY130_FD_SC_LP__NAND2B_LP%B
x_PM_SKY130_FD_SC_LP__NAND2B_LP%A_32_51# N_A_32_51#_M1000_s N_A_32_51#_M1003_s
+ N_A_32_51#_M1002_g N_A_32_51#_M1004_g N_A_32_51#_c_145_n N_A_32_51#_c_146_n
+ N_A_32_51#_c_147_n N_A_32_51#_c_148_n N_A_32_51#_c_149_n N_A_32_51#_c_154_n
+ N_A_32_51#_c_150_n N_A_32_51#_c_151_n N_A_32_51#_c_152_n
+ PM_SKY130_FD_SC_LP__NAND2B_LP%A_32_51#
x_PM_SKY130_FD_SC_LP__NAND2B_LP%VPWR N_VPWR_M1003_d N_VPWR_M1004_d
+ N_VPWR_c_214_n N_VPWR_c_215_n N_VPWR_c_216_n N_VPWR_c_217_n N_VPWR_c_218_n
+ VPWR N_VPWR_c_219_n N_VPWR_c_213_n PM_SKY130_FD_SC_LP__NAND2B_LP%VPWR
x_PM_SKY130_FD_SC_LP__NAND2B_LP%Y N_Y_M1002_d N_Y_M1006_d N_Y_c_249_n
+ N_Y_c_255_n N_Y_c_247_n N_Y_c_248_n Y Y N_Y_c_251_n
+ PM_SKY130_FD_SC_LP__NAND2B_LP%Y
x_PM_SKY130_FD_SC_LP__NAND2B_LP%VGND N_VGND_M1005_d N_VGND_c_283_n VGND
+ N_VGND_c_284_n N_VGND_c_285_n N_VGND_c_286_n N_VGND_c_287_n
+ PM_SKY130_FD_SC_LP__NAND2B_LP%VGND
cc_1 VNB N_A_N_c_52_n 0.0174092f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=0.75
cc_2 VNB N_A_N_c_53_n 0.0182818f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.71
cc_3 VNB N_A_N_c_54_n 0.0167417f $X=-0.19 $Y=-0.245 $X2=0.805 $Y2=0.825
cc_4 VNB N_A_N_c_55_n 0.0136346f $X=-0.19 $Y=-0.245 $X2=0.88 $Y2=0.75
cc_5 VNB N_A_N_c_56_n 0.00664349f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=0.825
cc_6 VNB N_A_N_c_57_n 0.0171752f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=1.39
cc_7 VNB N_A_N_c_58_n 0.00452877f $X=-0.19 $Y=-0.245 $X2=0.65 $Y2=1.39
cc_8 VNB N_A_N_c_59_n 0.0187633f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.225
cc_9 VNB N_B_M1001_g 0.0425078f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.71
cc_10 VNB N_B_c_102_n 0.018682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_B_c_103_n 0.0167746f $X=-0.19 $Y=-0.245 $X2=0.88 $Y2=0.465
cc_12 VNB N_B_c_104_n 0.00171359f $X=-0.19 $Y=-0.245 $X2=0.88 $Y2=0.465
cc_13 VNB N_A_32_51#_M1002_g 0.0250734f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=2.595
cc_14 VNB N_A_32_51#_M1004_g 0.00753721f $X=-0.19 $Y=-0.245 $X2=0.595 $Y2=0.825
cc_15 VNB N_A_32_51#_c_145_n 0.0259442f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=0.825
cc_16 VNB N_A_32_51#_c_146_n 0.0149892f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.895
cc_17 VNB N_A_32_51#_c_147_n 0.0242296f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.39
cc_18 VNB N_A_32_51#_c_148_n 0.029288f $X=-0.19 $Y=-0.245 $X2=0.66 $Y2=1.665
cc_19 VNB N_A_32_51#_c_149_n 0.0134429f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_32_51#_c_150_n 0.0285788f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_32_51#_c_151_n 0.0043171f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_32_51#_c_152_n 0.017547f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_VPWR_c_213_n 0.103974f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_Y_c_247_n 0.0466659f $X=-0.19 $Y=-0.245 $X2=0.805 $Y2=0.825
cc_25 VNB N_Y_c_248_n 0.0313303f $X=-0.19 $Y=-0.245 $X2=0.88 $Y2=0.465
cc_26 VNB N_VGND_c_283_n 0.00332502f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.41
cc_27 VNB N_VGND_c_284_n 0.0277505f $X=-0.19 $Y=-0.245 $X2=0.69 $Y2=2.595
cc_28 VNB N_VGND_c_285_n 0.0323914f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=0.825
cc_29 VNB N_VGND_c_286_n 0.173204f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.895
cc_30 VNB N_VGND_c_287_n 0.00463869f $X=-0.19 $Y=-0.245 $X2=0.63 $Y2=1.39
cc_31 VPB N_A_N_c_53_n 0.00404596f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=1.71
cc_32 VPB N_A_N_M1003_g 0.0331558f $X=-0.19 $Y=1.655 $X2=0.69 $Y2=2.595
cc_33 VPB N_A_N_c_62_n 0.0171944f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=1.895
cc_34 VPB N_A_N_c_58_n 0.00255957f $X=-0.19 $Y=1.655 $X2=0.65 $Y2=1.39
cc_35 VPB N_B_c_105_n 0.0139168f $X=-0.19 $Y=1.655 $X2=0.52 $Y2=0.75
cc_36 VPB N_B_M1006_g 0.0280138f $X=-0.19 $Y=1.655 $X2=0.52 $Y2=0.465
cc_37 VPB N_B_c_102_n 0.00524306f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_38 VPB N_B_c_104_n 7.45264e-19 $X=-0.19 $Y=1.655 $X2=0.88 $Y2=0.465
cc_39 VPB N_A_32_51#_M1004_g 0.0484076f $X=-0.19 $Y=1.655 $X2=0.595 $Y2=0.825
cc_40 VPB N_A_32_51#_c_154_n 0.0514144f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_41 VPB N_A_32_51#_c_150_n 0.0200965f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_42 VPB N_VPWR_c_214_n 0.00995657f $X=-0.19 $Y=1.655 $X2=0.69 $Y2=2.595
cc_43 VPB N_VPWR_c_215_n 0.0134668f $X=-0.19 $Y=1.655 $X2=0.595 $Y2=0.825
cc_44 VPB N_VPWR_c_216_n 0.0346158f $X=-0.19 $Y=1.655 $X2=0.88 $Y2=0.465
cc_45 VPB N_VPWR_c_217_n 0.0220566f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=1.895
cc_46 VPB N_VPWR_c_218_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_47 VPB N_VPWR_c_219_n 0.0203779f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_48 VPB N_VPWR_c_213_n 0.0490028f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_49 VPB N_Y_c_249_n 0.0118881f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=1.71
cc_50 VPB N_Y_c_247_n 0.026683f $X=-0.19 $Y=1.655 $X2=0.805 $Y2=0.825
cc_51 VPB N_Y_c_251_n 0.00763087f $X=-0.19 $Y=1.655 $X2=0.63 $Y2=1.225
cc_52 N_A_N_c_62_n N_B_c_105_n 0.0118472f $X=0.63 $Y=1.895 $X2=-0.19 $Y2=-0.245
cc_53 N_A_N_M1003_g N_B_M1006_g 0.0166121f $X=0.69 $Y=2.595 $X2=0 $Y2=0
cc_54 N_A_N_c_55_n N_B_M1001_g 0.0190109f $X=0.88 $Y=0.75 $X2=0 $Y2=0
cc_55 N_A_N_c_59_n N_B_M1001_g 0.00279366f $X=0.63 $Y=1.225 $X2=0 $Y2=0
cc_56 N_A_N_c_53_n N_B_c_102_n 0.0118472f $X=0.63 $Y=1.71 $X2=0 $Y2=0
cc_57 N_A_N_c_57_n N_B_c_103_n 0.0118472f $X=0.65 $Y=1.39 $X2=0 $Y2=0
cc_58 N_A_N_c_58_n N_B_c_103_n 0.00410205f $X=0.65 $Y=1.39 $X2=0 $Y2=0
cc_59 N_A_N_c_57_n N_B_c_104_n 8.22042e-19 $X=0.65 $Y=1.39 $X2=0 $Y2=0
cc_60 N_A_N_c_58_n N_B_c_104_n 0.0438819f $X=0.65 $Y=1.39 $X2=0 $Y2=0
cc_61 N_A_N_c_52_n N_A_32_51#_c_147_n 0.00987934f $X=0.52 $Y=0.75 $X2=0 $Y2=0
cc_62 N_A_N_c_55_n N_A_32_51#_c_147_n 0.00144103f $X=0.88 $Y=0.75 $X2=0 $Y2=0
cc_63 N_A_N_c_56_n N_A_32_51#_c_147_n 0.00836616f $X=0.52 $Y=0.825 $X2=0 $Y2=0
cc_64 N_A_N_c_54_n N_A_32_51#_c_148_n 0.0202378f $X=0.805 $Y=0.825 $X2=0 $Y2=0
cc_65 N_A_N_c_56_n N_A_32_51#_c_148_n 0.00576469f $X=0.52 $Y=0.825 $X2=0 $Y2=0
cc_66 N_A_N_c_57_n N_A_32_51#_c_148_n 7.23299e-19 $X=0.65 $Y=1.39 $X2=0 $Y2=0
cc_67 N_A_N_c_58_n N_A_32_51#_c_148_n 0.0262715f $X=0.65 $Y=1.39 $X2=0 $Y2=0
cc_68 N_A_N_c_59_n N_A_32_51#_c_148_n 0.00493967f $X=0.63 $Y=1.225 $X2=0 $Y2=0
cc_69 N_A_N_c_56_n N_A_32_51#_c_149_n 5.65839e-19 $X=0.52 $Y=0.825 $X2=0 $Y2=0
cc_70 N_A_N_c_59_n N_A_32_51#_c_149_n 0.00455711f $X=0.63 $Y=1.225 $X2=0 $Y2=0
cc_71 N_A_N_M1003_g N_A_32_51#_c_154_n 0.0236634f $X=0.69 $Y=2.595 $X2=0 $Y2=0
cc_72 N_A_N_c_62_n N_A_32_51#_c_154_n 0.0025759f $X=0.63 $Y=1.895 $X2=0 $Y2=0
cc_73 N_A_N_c_58_n N_A_32_51#_c_154_n 0.00867382f $X=0.65 $Y=1.39 $X2=0 $Y2=0
cc_74 N_A_N_M1003_g N_A_32_51#_c_150_n 0.00427061f $X=0.69 $Y=2.595 $X2=0 $Y2=0
cc_75 N_A_N_c_58_n N_A_32_51#_c_150_n 0.0483743f $X=0.65 $Y=1.39 $X2=0 $Y2=0
cc_76 N_A_N_c_59_n N_A_32_51#_c_150_n 0.0212209f $X=0.63 $Y=1.225 $X2=0 $Y2=0
cc_77 N_A_N_M1003_g N_VPWR_c_214_n 0.0239778f $X=0.69 $Y=2.595 $X2=0 $Y2=0
cc_78 N_A_N_c_58_n N_VPWR_c_214_n 0.00364455f $X=0.65 $Y=1.39 $X2=0 $Y2=0
cc_79 N_A_N_M1003_g N_VPWR_c_217_n 0.00840199f $X=0.69 $Y=2.595 $X2=0 $Y2=0
cc_80 N_A_N_M1003_g N_VPWR_c_213_n 0.014629f $X=0.69 $Y=2.595 $X2=0 $Y2=0
cc_81 N_A_N_c_52_n N_VGND_c_283_n 0.00228357f $X=0.52 $Y=0.75 $X2=0 $Y2=0
cc_82 N_A_N_c_55_n N_VGND_c_283_n 0.0126864f $X=0.88 $Y=0.75 $X2=0 $Y2=0
cc_83 N_A_N_c_52_n N_VGND_c_284_n 0.00530134f $X=0.52 $Y=0.75 $X2=0 $Y2=0
cc_84 N_A_N_c_54_n N_VGND_c_284_n 4.75415e-19 $X=0.805 $Y=0.825 $X2=0 $Y2=0
cc_85 N_A_N_c_55_n N_VGND_c_284_n 0.00469214f $X=0.88 $Y=0.75 $X2=0 $Y2=0
cc_86 N_A_N_c_52_n N_VGND_c_286_n 0.0105885f $X=0.52 $Y=0.75 $X2=0 $Y2=0
cc_87 N_A_N_c_54_n N_VGND_c_286_n 6.44251e-19 $X=0.805 $Y=0.825 $X2=0 $Y2=0
cc_88 N_A_N_c_55_n N_VGND_c_286_n 0.00807254f $X=0.88 $Y=0.75 $X2=0 $Y2=0
cc_89 N_B_M1001_g N_A_32_51#_M1002_g 0.0238835f $X=1.31 $Y=0.465 $X2=0 $Y2=0
cc_90 N_B_M1006_g N_A_32_51#_M1004_g 0.0277122f $X=1.22 $Y=2.595 $X2=0 $Y2=0
cc_91 N_B_c_102_n N_A_32_51#_c_145_n 0.0238835f $X=1.22 $Y=1.73 $X2=0 $Y2=0
cc_92 N_B_c_104_n N_A_32_51#_c_145_n 0.00354526f $X=1.22 $Y=1.39 $X2=0 $Y2=0
cc_93 N_B_c_105_n N_A_32_51#_c_146_n 0.0238835f $X=1.22 $Y=1.895 $X2=0 $Y2=0
cc_94 N_B_M1001_g N_A_32_51#_c_148_n 0.0156102f $X=1.31 $Y=0.465 $X2=0 $Y2=0
cc_95 N_B_c_103_n N_A_32_51#_c_148_n 0.00123028f $X=1.22 $Y=1.39 $X2=0 $Y2=0
cc_96 N_B_c_104_n N_A_32_51#_c_148_n 0.0245051f $X=1.22 $Y=1.39 $X2=0 $Y2=0
cc_97 N_B_M1006_g N_A_32_51#_c_154_n 2.56991e-19 $X=1.22 $Y=2.595 $X2=0 $Y2=0
cc_98 N_B_M1001_g N_A_32_51#_c_151_n 0.00233424f $X=1.31 $Y=0.465 $X2=0 $Y2=0
cc_99 N_B_c_104_n N_A_32_51#_c_151_n 0.0181736f $X=1.22 $Y=1.39 $X2=0 $Y2=0
cc_100 N_B_c_103_n N_A_32_51#_c_152_n 0.0238835f $X=1.22 $Y=1.39 $X2=0 $Y2=0
cc_101 N_B_c_105_n N_VPWR_c_214_n 3.03142e-19 $X=1.22 $Y=1.895 $X2=0 $Y2=0
cc_102 N_B_M1006_g N_VPWR_c_214_n 0.0227385f $X=1.22 $Y=2.595 $X2=0 $Y2=0
cc_103 N_B_c_104_n N_VPWR_c_214_n 0.00526295f $X=1.22 $Y=1.39 $X2=0 $Y2=0
cc_104 N_B_M1006_g N_VPWR_c_219_n 0.00840199f $X=1.22 $Y=2.595 $X2=0 $Y2=0
cc_105 N_B_M1006_g N_VPWR_c_213_n 0.0136033f $X=1.22 $Y=2.595 $X2=0 $Y2=0
cc_106 N_B_c_105_n N_Y_c_249_n 3.02817e-19 $X=1.22 $Y=1.895 $X2=0 $Y2=0
cc_107 N_B_M1006_g N_Y_c_249_n 0.00597514f $X=1.22 $Y=2.595 $X2=0 $Y2=0
cc_108 N_B_c_104_n N_Y_c_249_n 0.00534367f $X=1.22 $Y=1.39 $X2=0 $Y2=0
cc_109 N_B_M1006_g N_Y_c_255_n 0.0188476f $X=1.22 $Y=2.595 $X2=0 $Y2=0
cc_110 N_B_M1001_g N_Y_c_248_n 0.00120881f $X=1.31 $Y=0.465 $X2=0 $Y2=0
cc_111 N_B_M1001_g N_VGND_c_283_n 0.0129577f $X=1.31 $Y=0.465 $X2=0 $Y2=0
cc_112 N_B_M1001_g N_VGND_c_285_n 0.00469214f $X=1.31 $Y=0.465 $X2=0 $Y2=0
cc_113 N_B_M1001_g N_VGND_c_286_n 0.00818361f $X=1.31 $Y=0.465 $X2=0 $Y2=0
cc_114 N_A_32_51#_M1004_g N_VPWR_c_214_n 0.00128891f $X=1.75 $Y=2.595 $X2=0
+ $Y2=0
cc_115 N_A_32_51#_c_154_n N_VPWR_c_214_n 0.0668397f $X=0.425 $Y=2.24 $X2=0 $Y2=0
cc_116 N_A_32_51#_M1004_g N_VPWR_c_216_n 0.0215478f $X=1.75 $Y=2.595 $X2=0 $Y2=0
cc_117 N_A_32_51#_c_154_n N_VPWR_c_217_n 0.0281861f $X=0.425 $Y=2.24 $X2=0 $Y2=0
cc_118 N_A_32_51#_M1004_g N_VPWR_c_219_n 0.00811685f $X=1.75 $Y=2.595 $X2=0
+ $Y2=0
cc_119 N_A_32_51#_M1003_s N_VPWR_c_213_n 0.0023218f $X=0.28 $Y=2.095 $X2=0 $Y2=0
cc_120 N_A_32_51#_M1004_g N_VPWR_c_213_n 0.0140291f $X=1.75 $Y=2.595 $X2=0 $Y2=0
cc_121 N_A_32_51#_c_154_n N_VPWR_c_213_n 0.0173447f $X=0.425 $Y=2.24 $X2=0 $Y2=0
cc_122 N_A_32_51#_M1004_g N_Y_c_249_n 0.0058008f $X=1.75 $Y=2.595 $X2=0 $Y2=0
cc_123 N_A_32_51#_c_151_n N_Y_c_249_n 0.00485508f $X=1.79 $Y=1.04 $X2=0 $Y2=0
cc_124 N_A_32_51#_M1004_g N_Y_c_255_n 0.0277805f $X=1.75 $Y=2.595 $X2=0 $Y2=0
cc_125 N_A_32_51#_M1002_g N_Y_c_247_n 0.00502213f $X=1.7 $Y=0.465 $X2=0 $Y2=0
cc_126 N_A_32_51#_M1004_g N_Y_c_247_n 0.0123358f $X=1.75 $Y=2.595 $X2=0 $Y2=0
cc_127 N_A_32_51#_c_145_n N_Y_c_247_n 0.0111183f $X=1.79 $Y=1.38 $X2=0 $Y2=0
cc_128 N_A_32_51#_c_151_n N_Y_c_247_n 0.0488899f $X=1.79 $Y=1.04 $X2=0 $Y2=0
cc_129 N_A_32_51#_c_152_n N_Y_c_247_n 0.00117888f $X=1.79 $Y=1.04 $X2=0 $Y2=0
cc_130 N_A_32_51#_M1002_g N_Y_c_248_n 0.00854485f $X=1.7 $Y=0.465 $X2=0 $Y2=0
cc_131 N_A_32_51#_c_151_n N_Y_c_248_n 0.0166833f $X=1.79 $Y=1.04 $X2=0 $Y2=0
cc_132 N_A_32_51#_c_152_n N_Y_c_248_n 0.00133403f $X=1.79 $Y=1.04 $X2=0 $Y2=0
cc_133 N_A_32_51#_M1004_g N_Y_c_251_n 0.0172989f $X=1.75 $Y=2.595 $X2=0 $Y2=0
cc_134 N_A_32_51#_c_146_n N_Y_c_251_n 4.81734e-19 $X=1.79 $Y=1.545 $X2=0 $Y2=0
cc_135 N_A_32_51#_c_151_n N_Y_c_251_n 0.00928407f $X=1.79 $Y=1.04 $X2=0 $Y2=0
cc_136 N_A_32_51#_M1002_g N_VGND_c_283_n 0.00229479f $X=1.7 $Y=0.465 $X2=0 $Y2=0
cc_137 N_A_32_51#_c_147_n N_VGND_c_283_n 0.0144032f $X=0.305 $Y=0.48 $X2=0 $Y2=0
cc_138 N_A_32_51#_c_148_n N_VGND_c_283_n 0.026201f $X=1.625 $Y=0.96 $X2=0 $Y2=0
cc_139 N_A_32_51#_c_147_n N_VGND_c_284_n 0.0201256f $X=0.305 $Y=0.48 $X2=0 $Y2=0
cc_140 N_A_32_51#_M1002_g N_VGND_c_285_n 0.0052871f $X=1.7 $Y=0.465 $X2=0 $Y2=0
cc_141 N_A_32_51#_M1002_g N_VGND_c_286_n 0.0107684f $X=1.7 $Y=0.465 $X2=0 $Y2=0
cc_142 N_A_32_51#_c_147_n N_VGND_c_286_n 0.0127743f $X=0.305 $Y=0.48 $X2=0 $Y2=0
cc_143 N_VPWR_c_213_n N_Y_M1006_d 0.00223819f $X=2.16 $Y=3.33 $X2=0 $Y2=0
cc_144 N_VPWR_c_214_n N_Y_c_249_n 0.00525271f $X=0.955 $Y=2.24 $X2=0 $Y2=0
cc_145 N_VPWR_c_214_n N_Y_c_255_n 0.0613317f $X=0.955 $Y=2.24 $X2=0 $Y2=0
cc_146 N_VPWR_c_219_n N_Y_c_255_n 0.0232319f $X=1.915 $Y=3.33 $X2=0 $Y2=0
cc_147 N_VPWR_c_213_n N_Y_c_255_n 0.0152221f $X=2.16 $Y=3.33 $X2=0 $Y2=0
cc_148 N_VPWR_M1004_d N_Y_c_247_n 0.00129436f $X=1.875 $Y=2.095 $X2=0 $Y2=0
cc_149 N_VPWR_c_216_n N_Y_c_247_n 0.00948199f $X=2.08 $Y=2.495 $X2=0 $Y2=0
cc_150 N_VPWR_M1004_d N_Y_c_251_n 0.00245622f $X=1.875 $Y=2.095 $X2=0 $Y2=0
cc_151 N_VPWR_c_216_n N_Y_c_251_n 0.0161167f $X=2.08 $Y=2.495 $X2=0 $Y2=0
cc_152 N_Y_c_248_n N_VGND_c_283_n 0.0141494f $X=2.22 $Y=0.48 $X2=0 $Y2=0
cc_153 N_Y_c_248_n N_VGND_c_285_n 0.0337853f $X=2.22 $Y=0.48 $X2=0 $Y2=0
cc_154 N_Y_c_248_n N_VGND_c_286_n 0.021088f $X=2.22 $Y=0.48 $X2=0 $Y2=0
