* NGSPICE file created from sky130_fd_sc_lp__sdfxtp_4.ext - technology: sky130A

.subckt sky130_fd_sc_lp__sdfxtp_4 CLK D SCD SCE VGND VNB VPB VPWR Q
M1000 a_483_123# SCE a_359_123# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=3.087e+11p ps=3.15e+06u
M1001 VPWR SCD a_454_491# VPB phighvt w=640000u l=150000u
+  ad=2.6409e+12p pd=2.195e+07u as=2.048e+11p ps=1.92e+06u
M1002 a_1203_99# a_1053_125# VPWR VPB phighvt w=840000u l=150000u
+  ad=2.352e+11p pd=2.24e+06u as=0p ps=0u
M1003 a_850_51# a_641_123# VPWR VPB phighvt w=640000u l=150000u
+  ad=1.696e+11p pd=1.81e+06u as=0p ps=0u
M1004 VPWR a_1673_409# Q VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=7.056e+11p ps=6.16e+06u
M1005 VGND a_1673_409# Q VNB nshort w=840000u l=150000u
+  ad=1.8691e+12p pd=1.667e+07u as=4.704e+11p ps=4.48e+06u
M1006 a_850_51# a_641_123# VGND VNB nshort w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1007 a_454_491# a_91_123# a_359_123# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=2.905e+11p ps=3.21e+06u
M1008 a_1053_125# a_850_51# a_359_123# VPB phighvt w=420000u l=150000u
+  ad=2.149e+11p pd=1.92e+06u as=0p ps=0u
M1009 a_1053_125# a_641_123# a_359_123# VNB nshort w=420000u l=150000u
+  ad=1.26e+11p pd=1.44e+06u as=0p ps=0u
M1010 a_1143_125# a_850_51# a_1053_125# VNB nshort w=420000u l=150000u
+  ad=1.26e+11p pd=1.44e+06u as=0p ps=0u
M1011 Q a_1673_409# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VGND a_1203_99# a_1143_125# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_1673_409# a_1475_449# VGND VNB nshort w=840000u l=150000u
+  ad=2.226e+11p pd=2.21e+06u as=0p ps=0u
M1014 Q a_1673_409# VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_1673_409# a_1475_449# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=3.339e+11p pd=3.05e+06u as=0p ps=0u
M1016 a_296_491# SCE VPWR VPB phighvt w=640000u l=150000u
+  ad=1.344e+11p pd=1.7e+06u as=0p ps=0u
M1017 Q a_1673_409# VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VPWR a_1673_409# a_1631_507# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1019 a_1203_99# a_1053_125# VGND VNB nshort w=640000u l=150000u
+  ad=2.286e+11p pd=2.07e+06u as=0p ps=0u
M1020 a_359_123# D a_296_491# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VPWR a_1203_99# a_1199_449# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1022 a_1199_449# a_641_123# a_1053_125# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_1475_449# a_641_123# a_1203_99# VPB phighvt w=840000u l=150000u
+  ad=3.696e+11p pd=2.94e+06u as=0p ps=0u
M1024 Q a_1673_409# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 VGND a_1673_409# Q VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 VGND SCD a_483_123# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 VPWR SCE a_91_123# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.696e+11p ps=1.81e+06u
M1028 a_641_123# CLK VGND VNB nshort w=420000u l=150000u
+  ad=1.512e+11p pd=1.56e+06u as=0p ps=0u
M1029 VGND a_1673_409# a_1670_61# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.155e+11p ps=1.39e+06u
M1030 a_359_123# D a_260_123# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.449e+11p ps=1.53e+06u
M1031 a_641_123# CLK VPWR VPB phighvt w=640000u l=150000u
+  ad=1.696e+11p pd=1.81e+06u as=0p ps=0u
M1032 a_1631_507# a_850_51# a_1475_449# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 a_1475_449# a_850_51# a_1203_99# VNB nshort w=420000u l=150000u
+  ad=2.163e+11p pd=1.87e+06u as=0p ps=0u
M1034 a_1670_61# a_641_123# a_1475_449# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1035 VGND SCE a_91_123# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1036 VPWR a_1673_409# Q VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1037 a_260_123# a_91_123# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

