* File: sky130_fd_sc_lp__a221o_2.spice
* Created: Fri Aug 28 09:52:34 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__a221o_2.pex.spice"
.subckt sky130_fd_sc_lp__a221o_2  VNB VPB A2 A1 C1 B1 B2 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* B2	B2
* B1	B1
* C1	C1
* A1	A1
* A2	A2
* VPB	VPB
* VNB	VNB
MM1011 N_VGND_M1011_d N_A_86_27#_M1011_g N_X_M1011_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75001.7 A=0.126 P=1.98 MULT=1
MM1012 N_VGND_M1012_d N_A_86_27#_M1012_g N_X_M1011_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2604 AS=0.1176 PD=1.46 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75001.3 A=0.126 P=1.98 MULT=1
MM1008 A_356_53# N_A2_M1008_g N_VGND_M1012_d VNB NSHORT L=0.15 W=0.84 AD=0.0882
+ AS=0.2604 PD=1.05 PS=1.46 NRD=7.14 NRS=0 M=1 R=5.6 SA=75001.4 SB=75000.6
+ A=0.126 P=1.98 MULT=1
MM1003 N_A_86_27#_M1003_d N_A1_M1003_g A_356_53# VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.0882 PD=2.21 PS=1.05 NRD=0 NRS=7.14 M=1 R=5.6 SA=75001.7
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1013 N_A_86_27#_M1013_d N_C1_M1013_g N_VGND_M1013_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1006 A_739_49# N_B1_M1006_g N_A_86_27#_M1013_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1344 AS=0.1176 PD=1.16 PS=1.12 NRD=15 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75000.7 A=0.126 P=1.98 MULT=1
MM1001 N_VGND_M1001_d N_B2_M1001_g A_739_49# VNB NSHORT L=0.15 W=0.84 AD=0.2226
+ AS=0.1344 PD=2.21 PS=1.16 NRD=0 NRS=15 M=1 R=5.6 SA=75001.1 SB=75000.2 A=0.126
+ P=1.98 MULT=1
MM1004 N_X_M1004_d N_A_86_27#_M1004_g N_VPWR_M1004_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75001.7 A=0.189 P=2.82 MULT=1
MM1009 N_X_M1004_d N_A_86_27#_M1009_g N_VPWR_M1009_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.3213 PD=1.54 PS=1.77 NRD=0 NRS=18.7544 M=1 R=8.4 SA=75000.6
+ SB=75001.3 A=0.189 P=2.82 MULT=1
MM1000 N_A_334_367#_M1000_d N_A2_M1000_g N_VPWR_M1009_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.19845 AS=0.3213 PD=1.575 PS=1.77 NRD=0 NRS=17.1981 M=1 R=8.4
+ SA=75001.3 SB=75000.7 A=0.189 P=2.82 MULT=1
MM1007 N_VPWR_M1007_d N_A1_M1007_g N_A_334_367#_M1000_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.19845 PD=3.05 PS=1.575 NRD=0 NRS=5.4569 M=1 R=8.4
+ SA=75001.7 SB=75000.2 A=0.189 P=2.82 MULT=1
MM1010 N_A_653_367#_M1010_d N_C1_M1010_g N_A_86_27#_M1010_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1005 N_A_334_367#_M1005_d N_B1_M1005_g N_A_653_367#_M1010_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.2016 AS=0.1764 PD=1.58 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75000.7 A=0.189 P=2.82 MULT=1
MM1002 N_A_653_367#_M1002_d N_B2_M1002_g N_A_334_367#_M1005_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.2016 PD=3.05 PS=1.58 NRD=0 NRS=6.2449 M=1 R=8.4
+ SA=75001.1 SB=75000.2 A=0.189 P=2.82 MULT=1
DX14_noxref VNB VPB NWDIODE A=9.6607 P=14.09
*
.include "sky130_fd_sc_lp__a221o_2.pxi.spice"
*
.ends
*
*
