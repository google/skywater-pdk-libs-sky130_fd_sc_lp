* File: sky130_fd_sc_lp__sdfstp_2.pxi.spice
* Created: Wed Sep  2 10:35:44 2020
* 
x_PM_SKY130_FD_SC_LP__SDFSTP_2%SCD N_SCD_M1037_g N_SCD_c_266_n N_SCD_M1022_g
+ N_SCD_c_267_n N_SCD_c_268_n SCD SCD N_SCD_c_270_n
+ PM_SKY130_FD_SC_LP__SDFSTP_2%SCD
x_PM_SKY130_FD_SC_LP__SDFSTP_2%D N_D_c_300_n N_D_M1018_g N_D_M1015_g D D D D D
+ PM_SKY130_FD_SC_LP__SDFSTP_2%D
x_PM_SKY130_FD_SC_LP__SDFSTP_2%A_358_429# N_A_358_429#_M1026_d
+ N_A_358_429#_M1014_d N_A_358_429#_M1033_g N_A_358_429#_M1009_g
+ N_A_358_429#_c_342_n N_A_358_429#_c_343_n N_A_358_429#_c_350_n
+ N_A_358_429#_c_344_n N_A_358_429#_c_345_n N_A_358_429#_c_346_n
+ N_A_358_429#_c_347_n N_A_358_429#_c_353_n N_A_358_429#_c_348_n
+ PM_SKY130_FD_SC_LP__SDFSTP_2%A_358_429#
x_PM_SKY130_FD_SC_LP__SDFSTP_2%SCE N_SCE_M1017_g N_SCE_M1011_g N_SCE_c_415_n
+ N_SCE_c_416_n N_SCE_M1026_g N_SCE_c_418_n N_SCE_c_426_n N_SCE_M1014_g
+ N_SCE_c_419_n N_SCE_c_420_n N_SCE_c_421_n N_SCE_c_429_n N_SCE_c_422_n SCE SCE
+ SCE N_SCE_c_423_n N_SCE_c_424_n PM_SKY130_FD_SC_LP__SDFSTP_2%SCE
x_PM_SKY130_FD_SC_LP__SDFSTP_2%CLK N_CLK_M1010_g N_CLK_M1020_g N_CLK_c_500_n
+ N_CLK_c_504_n CLK CLK CLK N_CLK_c_502_n PM_SKY130_FD_SC_LP__SDFSTP_2%CLK
x_PM_SKY130_FD_SC_LP__SDFSTP_2%A_963_47# N_A_963_47#_M1023_d N_A_963_47#_M1000_d
+ N_A_963_47#_M1029_g N_A_963_47#_M1035_g N_A_963_47#_M1032_g
+ N_A_963_47#_M1008_g N_A_963_47#_c_549_n N_A_963_47#_c_541_n
+ N_A_963_47#_c_550_n N_A_963_47#_c_551_n N_A_963_47#_c_552_n
+ N_A_963_47#_c_553_n N_A_963_47#_c_554_n N_A_963_47#_c_555_n
+ N_A_963_47#_c_556_n N_A_963_47#_c_557_n N_A_963_47#_c_558_n
+ N_A_963_47#_c_559_n N_A_963_47#_c_560_n N_A_963_47#_c_542_n
+ N_A_963_47#_c_543_n N_A_963_47#_c_544_n N_A_963_47#_c_562_n
+ N_A_963_47#_c_563_n N_A_963_47#_c_545_n N_A_963_47#_c_565_n
+ PM_SKY130_FD_SC_LP__SDFSTP_2%A_963_47#
x_PM_SKY130_FD_SC_LP__SDFSTP_2%A_1365_29# N_A_1365_29#_M1024_s
+ N_A_1365_29#_M1040_d N_A_1365_29#_M1038_g N_A_1365_29#_M1005_g
+ N_A_1365_29#_c_715_n N_A_1365_29#_c_716_n N_A_1365_29#_c_717_n
+ N_A_1365_29#_c_718_n N_A_1365_29#_c_724_n N_A_1365_29#_c_719_n
+ N_A_1365_29#_c_720_n PM_SKY130_FD_SC_LP__SDFSTP_2%A_1365_29#
x_PM_SKY130_FD_SC_LP__SDFSTP_2%A_1237_55# N_A_1237_55#_M1034_d
+ N_A_1237_55#_M1029_d N_A_1237_55#_M1040_g N_A_1237_55#_c_777_n
+ N_A_1237_55#_M1024_g N_A_1237_55#_M1007_g N_A_1237_55#_c_779_n
+ N_A_1237_55#_c_780_n N_A_1237_55#_M1013_g N_A_1237_55#_c_869_p
+ N_A_1237_55#_c_781_n N_A_1237_55#_c_789_n N_A_1237_55#_c_782_n
+ N_A_1237_55#_c_783_n N_A_1237_55#_c_784_n N_A_1237_55#_c_785_n
+ N_A_1237_55#_c_786_n PM_SKY130_FD_SC_LP__SDFSTP_2%A_1237_55#
x_PM_SKY130_FD_SC_LP__SDFSTP_2%SET_B N_SET_B_M1004_g N_SET_B_M1027_g
+ N_SET_B_M1019_g N_SET_B_c_874_n N_SET_B_M1012_g N_SET_B_c_875_n
+ N_SET_B_c_876_n N_SET_B_c_877_n N_SET_B_c_878_n N_SET_B_c_879_n SET_B SET_B
+ SET_B SET_B N_SET_B_c_881_n N_SET_B_c_882_n PM_SKY130_FD_SC_LP__SDFSTP_2%SET_B
x_PM_SKY130_FD_SC_LP__SDFSTP_2%A_794_47# N_A_794_47#_M1010_s N_A_794_47#_M1020_s
+ N_A_794_47#_c_968_n N_A_794_47#_M1023_g N_A_794_47#_M1000_g
+ N_A_794_47#_c_978_n N_A_794_47#_c_969_n N_A_794_47#_c_979_n
+ N_A_794_47#_c_980_n N_A_794_47#_M1034_g N_A_794_47#_M1001_g
+ N_A_794_47#_c_982_n N_A_794_47#_c_983_n N_A_794_47#_M1030_g
+ N_A_794_47#_M1002_g N_A_794_47#_c_984_n N_A_794_47#_c_972_n
+ N_A_794_47#_c_985_n N_A_794_47#_c_973_n N_A_794_47#_c_974_n
+ N_A_794_47#_c_988_n N_A_794_47#_c_1096_p N_A_794_47#_c_1009_n
+ N_A_794_47#_c_975_n N_A_794_47#_c_976_n N_A_794_47#_c_990_n
+ N_A_794_47#_c_991_n PM_SKY130_FD_SC_LP__SDFSTP_2%A_794_47#
x_PM_SKY130_FD_SC_LP__SDFSTP_2%A_2214_99# N_A_2214_99#_M1031_d
+ N_A_2214_99#_M1003_d N_A_2214_99#_c_1137_n N_A_2214_99#_M1016_g
+ N_A_2214_99#_M1025_g N_A_2214_99#_c_1139_n N_A_2214_99#_c_1140_n
+ N_A_2214_99#_c_1141_n N_A_2214_99#_c_1142_n N_A_2214_99#_c_1143_n
+ PM_SKY130_FD_SC_LP__SDFSTP_2%A_2214_99#
x_PM_SKY130_FD_SC_LP__SDFSTP_2%A_1998_463# N_A_1998_463#_M1008_d
+ N_A_1998_463#_M1032_d N_A_1998_463#_M1012_d N_A_1998_463#_M1031_g
+ N_A_1998_463#_M1003_g N_A_1998_463#_c_1200_n N_A_1998_463#_M1006_g
+ N_A_1998_463#_c_1207_n N_A_1998_463#_M1041_g N_A_1998_463#_c_1202_n
+ N_A_1998_463#_c_1209_n N_A_1998_463#_c_1203_n N_A_1998_463#_c_1211_n
+ N_A_1998_463#_c_1204_n N_A_1998_463#_c_1213_n N_A_1998_463#_c_1231_n
+ N_A_1998_463#_c_1214_n N_A_1998_463#_c_1215_n
+ PM_SKY130_FD_SC_LP__SDFSTP_2%A_1998_463#
x_PM_SKY130_FD_SC_LP__SDFSTP_2%A_2686_131# N_A_2686_131#_M1006_s
+ N_A_2686_131#_M1041_s N_A_2686_131#_M1021_g N_A_2686_131#_M1028_g
+ N_A_2686_131#_c_1300_n N_A_2686_131#_M1036_g N_A_2686_131#_M1039_g
+ N_A_2686_131#_c_1303_n N_A_2686_131#_c_1304_n N_A_2686_131#_c_1310_n
+ N_A_2686_131#_c_1305_n N_A_2686_131#_c_1306_n N_A_2686_131#_c_1307_n
+ PM_SKY130_FD_SC_LP__SDFSTP_2%A_2686_131#
x_PM_SKY130_FD_SC_LP__SDFSTP_2%A_39_481# N_A_39_481#_M1037_s N_A_39_481#_M1033_d
+ N_A_39_481#_c_1365_n N_A_39_481#_c_1366_n N_A_39_481#_c_1367_n
+ PM_SKY130_FD_SC_LP__SDFSTP_2%A_39_481#
x_PM_SKY130_FD_SC_LP__SDFSTP_2%VPWR N_VPWR_M1037_d N_VPWR_M1014_s N_VPWR_M1020_d
+ N_VPWR_M1005_d N_VPWR_M1004_d N_VPWR_M1025_d N_VPWR_M1003_s N_VPWR_M1041_d
+ N_VPWR_M1039_d N_VPWR_c_1390_n N_VPWR_c_1391_n N_VPWR_c_1392_n N_VPWR_c_1393_n
+ N_VPWR_c_1394_n N_VPWR_c_1395_n N_VPWR_c_1396_n N_VPWR_c_1397_n
+ N_VPWR_c_1398_n N_VPWR_c_1399_n N_VPWR_c_1400_n N_VPWR_c_1401_n
+ N_VPWR_c_1402_n N_VPWR_c_1403_n N_VPWR_c_1404_n N_VPWR_c_1405_n
+ N_VPWR_c_1406_n N_VPWR_c_1407_n N_VPWR_c_1408_n N_VPWR_c_1409_n VPWR
+ N_VPWR_c_1410_n N_VPWR_c_1411_n N_VPWR_c_1412_n N_VPWR_c_1413_n
+ N_VPWR_c_1414_n N_VPWR_c_1415_n N_VPWR_c_1416_n N_VPWR_c_1389_n
+ PM_SKY130_FD_SC_LP__SDFSTP_2%VPWR
x_PM_SKY130_FD_SC_LP__SDFSTP_2%A_244_121# N_A_244_121#_M1011_d
+ N_A_244_121#_M1034_s N_A_244_121#_M1018_d N_A_244_121#_M1029_s
+ N_A_244_121#_c_1575_n N_A_244_121#_c_1563_n N_A_244_121#_c_1559_n
+ N_A_244_121#_c_1560_n N_A_244_121#_c_1561_n N_A_244_121#_c_1565_n
+ N_A_244_121#_c_1566_n N_A_244_121#_c_1567_n N_A_244_121#_c_1568_n
+ N_A_244_121#_c_1569_n N_A_244_121#_c_1623_n N_A_244_121#_c_1570_n
+ N_A_244_121#_c_1562_n N_A_244_121#_c_1572_n N_A_244_121#_c_1611_n
+ N_A_244_121#_c_1573_n N_A_244_121#_c_1574_n
+ PM_SKY130_FD_SC_LP__SDFSTP_2%A_244_121#
x_PM_SKY130_FD_SC_LP__SDFSTP_2%A_1781_379# N_A_1781_379#_M1007_d
+ N_A_1781_379#_M1030_d N_A_1781_379#_c_1697_n N_A_1781_379#_c_1698_n
+ N_A_1781_379#_c_1699_n N_A_1781_379#_c_1700_n
+ PM_SKY130_FD_SC_LP__SDFSTP_2%A_1781_379#
x_PM_SKY130_FD_SC_LP__SDFSTP_2%A_1888_463# N_A_1888_463#_M1032_s
+ N_A_1888_463#_M1025_s N_A_1888_463#_c_1733_n N_A_1888_463#_c_1734_n
+ N_A_1888_463#_c_1735_n PM_SKY130_FD_SC_LP__SDFSTP_2%A_1888_463#
x_PM_SKY130_FD_SC_LP__SDFSTP_2%Q N_Q_M1021_s N_Q_M1028_s N_Q_c_1787_p
+ N_Q_c_1779_n N_Q_c_1759_n N_Q_c_1761_n Q PM_SKY130_FD_SC_LP__SDFSTP_2%Q
x_PM_SKY130_FD_SC_LP__SDFSTP_2%VGND N_VGND_M1022_s N_VGND_M1009_d N_VGND_M1010_d
+ N_VGND_M1038_d N_VGND_M1027_d N_VGND_M1019_d N_VGND_M1006_d N_VGND_M1036_d
+ N_VGND_c_1790_n N_VGND_c_1791_n N_VGND_c_1792_n N_VGND_c_1793_n
+ N_VGND_c_1794_n N_VGND_c_1859_n N_VGND_c_1846_n N_VGND_c_1795_n
+ N_VGND_c_1796_n N_VGND_c_1797_n N_VGND_c_1798_n N_VGND_c_1799_n
+ N_VGND_c_1800_n N_VGND_c_1801_n N_VGND_c_1802_n N_VGND_c_1803_n
+ N_VGND_c_1804_n VGND N_VGND_c_1805_n N_VGND_c_1806_n N_VGND_c_1807_n
+ N_VGND_c_1808_n N_VGND_c_1809_n N_VGND_c_1810_n N_VGND_c_1811_n
+ N_VGND_c_1812_n N_VGND_c_1813_n N_VGND_c_1814_n
+ PM_SKY130_FD_SC_LP__SDFSTP_2%VGND
cc_1 VNB N_SCD_c_266_n 0.0210405f $X=-0.19 $Y=-0.245 $X2=0.785 $Y2=1.135
cc_2 VNB N_SCD_c_267_n 0.0437741f $X=-0.19 $Y=-0.245 $X2=0.785 $Y2=1.21
cc_3 VNB N_SCD_c_268_n 0.00398085f $X=-0.19 $Y=-0.245 $X2=0.415 $Y2=1.805
cc_4 VNB SCD 0.0250342f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_5 VNB N_SCD_c_270_n 0.0303661f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.3
cc_6 VNB N_D_M1015_g 0.0378577f $X=-0.19 $Y=-0.245 $X2=0.785 $Y2=0.815
cc_7 VNB N_A_358_429#_M1009_g 0.035391f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_358_429#_c_342_n 0.0669849f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_9 VNB N_A_358_429#_c_343_n 0.0014119f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_358_429#_c_344_n 0.00495357f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.3
cc_11 VNB N_A_358_429#_c_345_n 0.0163549f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_358_429#_c_346_n 0.00814111f $X=-0.19 $Y=-0.245 $X2=0.317 $Y2=1.3
cc_13 VNB N_A_358_429#_c_347_n 2.46275e-19 $X=-0.19 $Y=-0.245 $X2=0.317
+ $Y2=1.665
cc_14 VNB N_A_358_429#_c_348_n 0.0240148f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_SCE_M1011_g 0.0506093f $X=-0.19 $Y=-0.245 $X2=0.415 $Y2=1.21
cc_16 VNB N_SCE_c_415_n 0.101431f $X=-0.19 $Y=-0.245 $X2=0.415 $Y2=1.285
cc_17 VNB N_SCE_c_416_n 0.0124998f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_SCE_M1026_g 0.0353814f $X=-0.19 $Y=-0.245 $X2=0.415 $Y2=1.61
cc_19 VNB N_SCE_c_418_n 0.069973f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_20 VNB N_SCE_c_419_n 0.0474166f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.3
cc_21 VNB N_SCE_c_420_n 0.0210223f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_SCE_c_421_n 0.00749069f $X=-0.19 $Y=-0.245 $X2=0.317 $Y2=1.665
cc_23 VNB N_SCE_c_422_n 0.0198493f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_SCE_c_423_n 0.0452768f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_SCE_c_424_n 0.00640764f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_CLK_M1010_g 0.0405345f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=2.725
cc_27 VNB N_CLK_c_500_n 0.0240162f $X=-0.19 $Y=-0.245 $X2=0.785 $Y2=1.21
cc_28 VNB CLK 0.00858713f $X=-0.19 $Y=-0.245 $X2=0.415 $Y2=1.61
cc_29 VNB N_CLK_c_502_n 0.0170015f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.3
cc_30 VNB N_A_963_47#_M1035_g 0.0320697f $X=-0.19 $Y=-0.245 $X2=0.415 $Y2=1.61
cc_31 VNB N_A_963_47#_M1008_g 0.0387383f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.3
cc_32 VNB N_A_963_47#_c_541_n 0.0126109f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_963_47#_c_542_n 0.00815578f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_963_47#_c_543_n 2.27796e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_963_47#_c_544_n 0.00617453f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_963_47#_c_545_n 0.0658183f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_1365_29#_c_715_n 0.0356155f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_1365_29#_c_716_n 0.018051f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.3
cc_39 VNB N_A_1365_29#_c_717_n 0.00713527f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_1365_29#_c_718_n 0.0148128f $X=-0.19 $Y=-0.245 $X2=0.317 $Y2=1.665
cc_41 VNB N_A_1365_29#_c_719_n 0.0190033f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_1365_29#_c_720_n 0.0210963f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_1237_55#_M1040_g 0.0102005f $X=-0.19 $Y=-0.245 $X2=0.415 $Y2=1.285
cc_44 VNB N_A_1237_55#_c_777_n 0.0213571f $X=-0.19 $Y=-0.245 $X2=0.785 $Y2=1.21
cc_45 VNB N_A_1237_55#_M1007_g 0.0109531f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_46 VNB N_A_1237_55#_c_779_n 0.0321704f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_1237_55#_c_780_n 0.0173557f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.3
cc_48 VNB N_A_1237_55#_c_781_n 0.00790391f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_1237_55#_c_782_n 0.0453387f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_1237_55#_c_783_n 0.0409411f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_1237_55#_c_784_n 7.2595e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_1237_55#_c_785_n 0.00146392f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_1237_55#_c_786_n 0.0372402f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_SET_B_M1027_g 0.0356565f $X=-0.19 $Y=-0.245 $X2=0.415 $Y2=1.21
cc_55 VNB N_SET_B_M1019_g 0.0284758f $X=-0.19 $Y=-0.245 $X2=0.785 $Y2=1.21
cc_56 VNB N_SET_B_c_874_n 0.0228474f $X=-0.19 $Y=-0.245 $X2=0.415 $Y2=1.61
cc_57 VNB N_SET_B_c_875_n 0.0104121f $X=-0.19 $Y=-0.245 $X2=0.415 $Y2=1.3
cc_58 VNB N_SET_B_c_876_n 0.0126503f $X=-0.19 $Y=-0.245 $X2=0.317 $Y2=1.295
cc_59 VNB N_SET_B_c_877_n 2.97037e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_SET_B_c_878_n 0.0061625f $X=-0.19 $Y=-0.245 $X2=0.317 $Y2=1.3
cc_61 VNB N_SET_B_c_879_n 0.0320343f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB SET_B 0.00171253f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_SET_B_c_881_n 0.0528459f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_SET_B_c_882_n 0.0155218f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_A_794_47#_c_968_n 0.0204004f $X=-0.19 $Y=-0.245 $X2=0.785 $Y2=0.815
cc_66 VNB N_A_794_47#_c_969_n 0.0474747f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_67 VNB N_A_794_47#_M1034_g 0.0318076f $X=-0.19 $Y=-0.245 $X2=0.317 $Y2=1.295
cc_68 VNB N_A_794_47#_M1002_g 0.0481647f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_794_47#_c_972_n 0.0535429f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_A_794_47#_c_973_n 0.0169555f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_A_794_47#_c_974_n 0.0194337f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_A_794_47#_c_975_n 0.0538325f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_A_794_47#_c_976_n 0.00217951f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_A_2214_99#_c_1137_n 0.0194987f $X=-0.19 $Y=-0.245 $X2=0.785
+ $Y2=0.815
cc_75 VNB N_A_2214_99#_M1025_g 0.00941713f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_A_2214_99#_c_1139_n 0.0200974f $X=-0.19 $Y=-0.245 $X2=0.415
+ $Y2=1.805
cc_77 VNB N_A_2214_99#_c_1140_n 0.0508197f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_A_2214_99#_c_1141_n 0.0128474f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.3
cc_79 VNB N_A_2214_99#_c_1142_n 0.0256076f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_A_2214_99#_c_1143_n 0.00409067f $X=-0.19 $Y=-0.245 $X2=0.317 $Y2=1.3
cc_81 VNB N_A_1998_463#_M1031_g 0.04967f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_A_1998_463#_c_1200_n 0.0305071f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_A_1998_463#_M1006_g 0.043447f $X=-0.19 $Y=-0.245 $X2=0.317 $Y2=1.295
cc_84 VNB N_A_1998_463#_c_1202_n 0.015619f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_A_1998_463#_c_1203_n 0.0023032f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_A_1998_463#_c_1204_n 0.00755538f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_A_2686_131#_M1021_g 0.026492f $X=-0.19 $Y=-0.245 $X2=0.415 $Y2=1.285
cc_88 VNB N_A_2686_131#_M1028_g 4.96559e-19 $X=-0.19 $Y=-0.245 $X2=0.415
+ $Y2=1.61
cc_89 VNB N_A_2686_131#_c_1300_n 0.0116475f $X=-0.19 $Y=-0.245 $X2=0.155
+ $Y2=1.21
cc_90 VNB N_A_2686_131#_M1036_g 0.0261688f $X=-0.19 $Y=-0.245 $X2=0.415 $Y2=1.3
cc_91 VNB N_A_2686_131#_M1039_g 0.0104331f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_A_2686_131#_c_1303_n 0.00666901f $X=-0.19 $Y=-0.245 $X2=0.317
+ $Y2=1.3
cc_93 VNB N_A_2686_131#_c_1304_n 0.0143336f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_94 VNB N_A_2686_131#_c_1305_n 0.005352f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_95 VNB N_A_2686_131#_c_1306_n 0.00350666f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_96 VNB N_A_2686_131#_c_1307_n 0.0274742f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_97 VNB N_VPWR_c_1389_n 0.641339f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_98 VNB N_A_244_121#_c_1559_n 0.0249508f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.3
cc_99 VNB N_A_244_121#_c_1560_n 0.00326949f $X=-0.19 $Y=-0.245 $X2=0.317
+ $Y2=1.295
cc_100 VNB N_A_244_121#_c_1561_n 0.00206099f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_101 VNB N_A_244_121#_c_1562_n 0.0114864f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_102 VNB N_Q_c_1759_n 0.0205955f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_103 VNB Q 0.0300142f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_104 VNB N_VGND_c_1790_n 0.0389543f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_105 VNB N_VGND_c_1791_n 0.0153594f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_106 VNB N_VGND_c_1792_n 0.00519343f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_107 VNB N_VGND_c_1793_n 0.0146786f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_108 VNB N_VGND_c_1794_n 0.0164213f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_109 VNB N_VGND_c_1795_n 0.0282207f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_110 VNB N_VGND_c_1796_n 0.0192477f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_111 VNB N_VGND_c_1797_n 0.0159479f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_112 VNB N_VGND_c_1798_n 0.0239641f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_113 VNB N_VGND_c_1799_n 0.0198259f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_114 VNB N_VGND_c_1800_n 0.00326991f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_115 VNB N_VGND_c_1801_n 0.0941749f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_116 VNB N_VGND_c_1802_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_117 VNB N_VGND_c_1803_n 0.0491843f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_118 VNB N_VGND_c_1804_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_119 VNB N_VGND_c_1805_n 0.0150312f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_120 VNB N_VGND_c_1806_n 0.0373156f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_121 VNB N_VGND_c_1807_n 0.0489375f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_122 VNB N_VGND_c_1808_n 0.0583576f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_123 VNB N_VGND_c_1809_n 0.0158018f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_124 VNB N_VGND_c_1810_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_125 VNB N_VGND_c_1811_n 0.0086911f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_126 VNB N_VGND_c_1812_n 0.00487954f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_127 VNB N_VGND_c_1813_n 0.00540966f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_128 VNB N_VGND_c_1814_n 0.851783f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_129 VPB N_SCD_M1037_g 0.0554593f $X=-0.19 $Y=1.655 $X2=0.535 $Y2=2.725
cc_130 VPB N_SCD_c_268_n 0.0201615f $X=-0.19 $Y=1.655 $X2=0.415 $Y2=1.805
cc_131 VPB SCD 0.0061149f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_132 VPB N_D_c_300_n 0.0440016f $X=-0.19 $Y=1.655 $X2=0.535 $Y2=1.805
cc_133 VPB N_D_M1018_g 0.0199571f $X=-0.19 $Y=1.655 $X2=0.535 $Y2=2.725
cc_134 VPB N_D_M1015_g 0.00557882f $X=-0.19 $Y=1.655 $X2=0.785 $Y2=0.815
cc_135 VPB D 0.0460346f $X=-0.19 $Y=1.655 $X2=0.415 $Y2=1.61
cc_136 VPB N_A_358_429#_c_343_n 0.0286942f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_137 VPB N_A_358_429#_c_350_n 0.0348568f $X=-0.19 $Y=1.655 $X2=0.415 $Y2=1.3
cc_138 VPB N_A_358_429#_c_346_n 0.00332035f $X=-0.19 $Y=1.655 $X2=0.317 $Y2=1.3
cc_139 VPB N_A_358_429#_c_347_n 0.00282776f $X=-0.19 $Y=1.655 $X2=0.317
+ $Y2=1.665
cc_140 VPB N_A_358_429#_c_353_n 0.0155467f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_141 VPB N_A_358_429#_c_348_n 0.0201812f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_142 VPB N_SCE_M1017_g 0.0462189f $X=-0.19 $Y=1.655 $X2=0.535 $Y2=2.725
cc_143 VPB N_SCE_c_426_n 0.0220856f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_144 VPB N_SCE_c_419_n 0.0237393f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.3
cc_145 VPB N_SCE_c_420_n 0.00716609f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_146 VPB N_SCE_c_429_n 0.0305575f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_147 VPB N_CLK_M1020_g 0.0478083f $X=-0.19 $Y=1.655 $X2=0.785 $Y2=0.815
cc_148 VPB N_CLK_c_504_n 0.0168049f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_149 VPB CLK 0.0031373f $X=-0.19 $Y=1.655 $X2=0.415 $Y2=1.61
cc_150 VPB N_A_963_47#_M1029_g 0.0343082f $X=-0.19 $Y=1.655 $X2=0.415 $Y2=1.285
cc_151 VPB N_A_963_47#_M1032_g 0.0244374f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_152 VPB N_A_963_47#_M1008_g 0.00864945f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.3
cc_153 VPB N_A_963_47#_c_549_n 0.0162198f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_154 VPB N_A_963_47#_c_550_n 0.0058973f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_155 VPB N_A_963_47#_c_551_n 0.0151349f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_156 VPB N_A_963_47#_c_552_n 0.00152609f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_157 VPB N_A_963_47#_c_553_n 0.00723901f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_158 VPB N_A_963_47#_c_554_n 0.00265738f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_159 VPB N_A_963_47#_c_555_n 4.9078e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_160 VPB N_A_963_47#_c_556_n 0.0170584f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_161 VPB N_A_963_47#_c_557_n 0.0029026f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_162 VPB N_A_963_47#_c_558_n 0.00277529f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_163 VPB N_A_963_47#_c_559_n 0.0191875f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_164 VPB N_A_963_47#_c_560_n 3.66301e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_165 VPB N_A_963_47#_c_543_n 0.0011811f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_166 VPB N_A_963_47#_c_562_n 0.00240678f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_167 VPB N_A_963_47#_c_563_n 0.0107523f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_168 VPB N_A_963_47#_c_545_n 0.0255343f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_169 VPB N_A_963_47#_c_565_n 0.0454838f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_170 VPB N_A_1365_29#_M1005_g 0.025286f $X=-0.19 $Y=1.655 $X2=0.415 $Y2=1.805
cc_171 VPB N_A_1365_29#_c_717_n 0.00834469f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_172 VPB N_A_1365_29#_c_718_n 0.0185056f $X=-0.19 $Y=1.655 $X2=0.317 $Y2=1.665
cc_173 VPB N_A_1365_29#_c_724_n 0.00367503f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_174 VPB N_A_1237_55#_M1040_g 0.0366587f $X=-0.19 $Y=1.655 $X2=0.415 $Y2=1.285
cc_175 VPB N_A_1237_55#_M1007_g 0.0273953f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_176 VPB N_A_1237_55#_c_789_n 0.00670709f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_177 VPB N_SET_B_M1004_g 0.0225759f $X=-0.19 $Y=1.655 $X2=0.535 $Y2=2.725
cc_178 VPB N_SET_B_c_874_n 0.0162783f $X=-0.19 $Y=1.655 $X2=0.415 $Y2=1.61
cc_179 VPB N_SET_B_M1012_g 0.0323425f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_180 VPB N_SET_B_c_875_n 0.00533633f $X=-0.19 $Y=1.655 $X2=0.415 $Y2=1.3
cc_181 VPB N_SET_B_c_878_n 0.00620862f $X=-0.19 $Y=1.655 $X2=0.317 $Y2=1.3
cc_182 VPB N_A_794_47#_M1000_g 0.0189789f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_183 VPB N_A_794_47#_c_978_n 0.0462455f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_184 VPB N_A_794_47#_c_979_n 0.0703139f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_185 VPB N_A_794_47#_c_980_n 0.0106266f $X=-0.19 $Y=1.655 $X2=0.415 $Y2=1.3
cc_186 VPB N_A_794_47#_M1001_g 0.0484463f $X=-0.19 $Y=1.655 $X2=0.317 $Y2=1.665
cc_187 VPB N_A_794_47#_c_982_n 0.32656f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_188 VPB N_A_794_47#_c_983_n 0.0135813f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_189 VPB N_A_794_47#_c_984_n 0.0718578f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_190 VPB N_A_794_47#_c_985_n 0.00749069f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_191 VPB N_A_794_47#_c_973_n 0.0275861f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_192 VPB N_A_794_47#_c_974_n 0.0073071f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_193 VPB N_A_794_47#_c_988_n 0.00964137f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_194 VPB N_A_794_47#_c_975_n 0.0301777f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_195 VPB N_A_794_47#_c_990_n 0.0108011f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_196 VPB N_A_794_47#_c_991_n 0.0380126f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_197 VPB N_A_2214_99#_M1025_g 0.038157f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_198 VPB N_A_2214_99#_c_1143_n 0.0207064f $X=-0.19 $Y=1.655 $X2=0.317 $Y2=1.3
cc_199 VPB N_A_1998_463#_M1003_g 0.0264563f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_200 VPB N_A_1998_463#_c_1200_n 0.0272266f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_201 VPB N_A_1998_463#_c_1207_n 0.0203394f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_202 VPB N_A_1998_463#_c_1202_n 0.0109685f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_203 VPB N_A_1998_463#_c_1209_n 0.0240693f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_204 VPB N_A_1998_463#_c_1203_n 0.00273241f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_205 VPB N_A_1998_463#_c_1211_n 0.00190829f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_206 VPB N_A_1998_463#_c_1204_n 0.00413407f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_207 VPB N_A_1998_463#_c_1213_n 0.0151524f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_208 VPB N_A_1998_463#_c_1214_n 0.0297696f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_209 VPB N_A_1998_463#_c_1215_n 0.0233827f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_210 VPB N_A_2686_131#_M1028_g 0.0223654f $X=-0.19 $Y=1.655 $X2=0.415 $Y2=1.61
cc_211 VPB N_A_2686_131#_M1039_g 0.0227559f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_212 VPB N_A_2686_131#_c_1310_n 0.013686f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_213 VPB N_A_39_481#_c_1365_n 0.0126642f $X=-0.19 $Y=1.655 $X2=0.785 $Y2=0.815
cc_214 VPB N_A_39_481#_c_1366_n 0.0179478f $X=-0.19 $Y=1.655 $X2=0.415 $Y2=1.285
cc_215 VPB N_A_39_481#_c_1367_n 0.0134114f $X=-0.19 $Y=1.655 $X2=0.415 $Y2=1.61
cc_216 VPB N_VPWR_c_1390_n 0.00177638f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_217 VPB N_VPWR_c_1391_n 0.0188507f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_218 VPB N_VPWR_c_1392_n 0.00151893f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_219 VPB N_VPWR_c_1393_n 0.0209706f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_220 VPB N_VPWR_c_1394_n 0.0206641f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_221 VPB N_VPWR_c_1395_n 0.0201529f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_222 VPB N_VPWR_c_1396_n 0.0194327f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_223 VPB N_VPWR_c_1397_n 0.0235737f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_224 VPB N_VPWR_c_1398_n 0.015922f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_225 VPB N_VPWR_c_1399_n 0.0388805f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_226 VPB N_VPWR_c_1400_n 0.0449228f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_227 VPB N_VPWR_c_1401_n 0.00497514f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_228 VPB N_VPWR_c_1402_n 0.0509705f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_229 VPB N_VPWR_c_1403_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_230 VPB N_VPWR_c_1404_n 0.0321592f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_231 VPB N_VPWR_c_1405_n 0.00297041f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_232 VPB N_VPWR_c_1406_n 0.0713504f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_233 VPB N_VPWR_c_1407_n 0.00487897f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_234 VPB N_VPWR_c_1408_n 0.0333411f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_235 VPB N_VPWR_c_1409_n 0.00584081f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_236 VPB N_VPWR_c_1410_n 0.0169688f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_237 VPB N_VPWR_c_1411_n 0.0367197f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_238 VPB N_VPWR_c_1412_n 0.0207798f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_239 VPB N_VPWR_c_1413_n 0.0131639f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_240 VPB N_VPWR_c_1414_n 0.00497475f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_241 VPB N_VPWR_c_1415_n 0.00485155f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_242 VPB N_VPWR_c_1416_n 0.00612923f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_243 VPB N_VPWR_c_1389_n 0.138812f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_244 VPB N_A_244_121#_c_1563_n 0.0206192f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_245 VPB N_A_244_121#_c_1561_n 0.0103352f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_246 VPB N_A_244_121#_c_1565_n 0.0183336f $X=-0.19 $Y=1.655 $X2=0.317
+ $Y2=1.665
cc_247 VPB N_A_244_121#_c_1566_n 0.0239213f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_248 VPB N_A_244_121#_c_1567_n 0.00262807f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_249 VPB N_A_244_121#_c_1568_n 0.013494f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_250 VPB N_A_244_121#_c_1569_n 0.0013657f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_251 VPB N_A_244_121#_c_1570_n 0.00575065f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_252 VPB N_A_244_121#_c_1562_n 0.00413225f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_253 VPB N_A_244_121#_c_1572_n 0.00225097f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_254 VPB N_A_244_121#_c_1573_n 0.00189763f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_255 VPB N_A_244_121#_c_1574_n 0.00259431f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_256 VPB N_A_1781_379#_c_1697_n 0.0140616f $X=-0.19 $Y=1.655 $X2=0.415
+ $Y2=1.285
cc_257 VPB N_A_1781_379#_c_1698_n 0.00419811f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_258 VPB N_A_1781_379#_c_1699_n 0.00687037f $X=-0.19 $Y=1.655 $X2=0.415
+ $Y2=1.805
cc_259 VPB N_A_1781_379#_c_1700_n 0.00325022f $X=-0.19 $Y=1.655 $X2=0.155
+ $Y2=1.21
cc_260 VPB N_A_1888_463#_c_1733_n 0.0236764f $X=-0.19 $Y=1.655 $X2=0.785
+ $Y2=0.815
cc_261 VPB N_A_1888_463#_c_1734_n 0.00732699f $X=-0.19 $Y=1.655 $X2=0.785
+ $Y2=1.21
cc_262 VPB N_A_1888_463#_c_1735_n 0.00837013f $X=-0.19 $Y=1.655 $X2=0.415
+ $Y2=1.805
cc_263 VPB N_Q_c_1761_n 0.0184805f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.3
cc_264 VPB Q 0.0102511f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_265 N_SCD_M1037_g D 0.0190136f $X=0.535 $Y=2.725 $X2=0 $Y2=0
cc_266 N_SCD_c_267_n D 0.00609731f $X=0.785 $Y=1.21 $X2=0 $Y2=0
cc_267 N_SCD_c_268_n D 0.00647718f $X=0.415 $Y=1.805 $X2=0 $Y2=0
cc_268 SCD D 0.0383479f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_269 N_SCD_c_268_n N_SCE_M1017_g 0.055676f $X=0.415 $Y=1.805 $X2=0 $Y2=0
cc_270 SCD N_SCE_M1017_g 5.75322e-19 $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_271 N_SCD_c_266_n N_SCE_M1011_g 0.0487148f $X=0.785 $Y=1.135 $X2=0 $Y2=0
cc_272 SCD N_SCE_M1011_g 0.0012814f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_273 N_SCD_c_270_n N_SCE_M1011_g 0.00637482f $X=0.385 $Y=1.3 $X2=0 $Y2=0
cc_274 SCD N_SCE_c_420_n 9.13167e-19 $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_275 N_SCD_c_270_n N_SCE_c_420_n 0.00868821f $X=0.385 $Y=1.3 $X2=0 $Y2=0
cc_276 N_SCD_M1037_g N_A_39_481#_c_1366_n 4.46816e-19 $X=0.535 $Y=2.725 $X2=0
+ $Y2=0
cc_277 N_SCD_M1037_g N_A_39_481#_c_1367_n 0.0119172f $X=0.535 $Y=2.725 $X2=0
+ $Y2=0
cc_278 N_SCD_M1037_g N_VPWR_c_1390_n 0.00776857f $X=0.535 $Y=2.725 $X2=0 $Y2=0
cc_279 N_SCD_M1037_g N_VPWR_c_1410_n 0.00325653f $X=0.535 $Y=2.725 $X2=0 $Y2=0
cc_280 N_SCD_M1037_g N_VPWR_c_1389_n 0.00471934f $X=0.535 $Y=2.725 $X2=0 $Y2=0
cc_281 N_SCD_c_266_n N_A_244_121#_c_1575_n 0.0017569f $X=0.785 $Y=1.135 $X2=0
+ $Y2=0
cc_282 N_SCD_c_267_n N_A_244_121#_c_1560_n 5.01393e-19 $X=0.785 $Y=1.21 $X2=0
+ $Y2=0
cc_283 SCD N_A_244_121#_c_1560_n 0.0068351f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_284 N_SCD_c_270_n N_A_244_121#_c_1560_n 4.3985e-19 $X=0.385 $Y=1.3 $X2=0
+ $Y2=0
cc_285 N_SCD_c_266_n N_VGND_c_1790_n 0.0128531f $X=0.785 $Y=1.135 $X2=0 $Y2=0
cc_286 N_SCD_c_267_n N_VGND_c_1790_n 0.00971745f $X=0.785 $Y=1.21 $X2=0 $Y2=0
cc_287 SCD N_VGND_c_1790_n 0.0124971f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_288 N_SCD_c_266_n N_VGND_c_1806_n 0.00354091f $X=0.785 $Y=1.135 $X2=0 $Y2=0
cc_289 N_SCD_c_266_n N_VGND_c_1814_n 0.00398995f $X=0.785 $Y=1.135 $X2=0 $Y2=0
cc_290 N_D_M1015_g N_A_358_429#_M1009_g 0.0453695f $X=1.575 $Y=0.815 $X2=0 $Y2=0
cc_291 D N_A_358_429#_c_342_n 0.0047786f $X=2.075 $Y=1.95 $X2=0 $Y2=0
cc_292 N_D_c_300_n N_A_358_429#_c_343_n 0.0111992f $X=1.325 $Y=2.245 $X2=0 $Y2=0
cc_293 D N_A_358_429#_c_343_n 0.0126651f $X=2.075 $Y=1.95 $X2=0 $Y2=0
cc_294 N_D_c_300_n N_A_358_429#_c_350_n 0.00662939f $X=1.325 $Y=2.245 $X2=0
+ $Y2=0
cc_295 N_D_M1018_g N_A_358_429#_c_350_n 0.0201196f $X=1.325 $Y=2.725 $X2=0 $Y2=0
cc_296 D N_A_358_429#_c_350_n 0.00773081f $X=2.075 $Y=1.95 $X2=0 $Y2=0
cc_297 N_D_c_300_n N_A_358_429#_c_344_n 0.0453695f $X=1.325 $Y=2.245 $X2=0 $Y2=0
cc_298 N_D_c_300_n N_SCE_M1017_g 0.0867094f $X=1.325 $Y=2.245 $X2=0 $Y2=0
cc_299 N_D_M1015_g N_SCE_M1017_g 0.00255628f $X=1.575 $Y=0.815 $X2=0 $Y2=0
cc_300 D N_SCE_M1017_g 0.0181042f $X=2.075 $Y=1.95 $X2=0 $Y2=0
cc_301 N_D_M1015_g N_SCE_M1011_g 0.0393847f $X=1.575 $Y=0.815 $X2=0 $Y2=0
cc_302 N_D_M1015_g N_SCE_c_415_n 0.0103352f $X=1.575 $Y=0.815 $X2=0 $Y2=0
cc_303 D N_SCE_c_420_n 0.00748754f $X=2.075 $Y=1.95 $X2=0 $Y2=0
cc_304 D N_A_39_481#_c_1365_n 0.0226773f $X=2.075 $Y=1.95 $X2=0 $Y2=0
cc_305 N_D_c_300_n N_A_39_481#_c_1367_n 0.00462833f $X=1.325 $Y=2.245 $X2=0
+ $Y2=0
cc_306 N_D_M1018_g N_A_39_481#_c_1367_n 0.0151271f $X=1.325 $Y=2.725 $X2=0 $Y2=0
cc_307 D N_A_39_481#_c_1367_n 0.141341f $X=2.075 $Y=1.95 $X2=0 $Y2=0
cc_308 N_D_M1018_g N_VPWR_c_1390_n 0.00154332f $X=1.325 $Y=2.725 $X2=0 $Y2=0
cc_309 N_D_M1018_g N_VPWR_c_1400_n 0.00391581f $X=1.325 $Y=2.725 $X2=0 $Y2=0
cc_310 N_D_M1018_g N_VPWR_c_1389_n 0.00567109f $X=1.325 $Y=2.725 $X2=0 $Y2=0
cc_311 N_D_M1015_g N_A_244_121#_c_1575_n 0.0101773f $X=1.575 $Y=0.815 $X2=0
+ $Y2=0
cc_312 N_D_M1018_g N_A_244_121#_c_1563_n 4.6748e-19 $X=1.325 $Y=2.725 $X2=0
+ $Y2=0
cc_313 D N_A_244_121#_c_1563_n 3.39772e-19 $X=2.075 $Y=1.95 $X2=0 $Y2=0
cc_314 N_D_M1015_g N_A_244_121#_c_1559_n 0.0138596f $X=1.575 $Y=0.815 $X2=0
+ $Y2=0
cc_315 D N_A_244_121#_c_1559_n 0.0241927f $X=2.075 $Y=1.95 $X2=0 $Y2=0
cc_316 N_D_c_300_n N_A_244_121#_c_1560_n 0.00551655f $X=1.325 $Y=2.245 $X2=0
+ $Y2=0
cc_317 N_D_M1015_g N_A_244_121#_c_1560_n 0.00426595f $X=1.575 $Y=0.815 $X2=0
+ $Y2=0
cc_318 D N_A_244_121#_c_1560_n 0.011463f $X=2.075 $Y=1.95 $X2=0 $Y2=0
cc_319 D N_A_244_121#_c_1565_n 0.00874591f $X=2.075 $Y=1.95 $X2=0 $Y2=0
cc_320 D N_A_244_121#_c_1572_n 0.0158346f $X=2.075 $Y=1.95 $X2=0 $Y2=0
cc_321 N_D_M1015_g N_VGND_c_1791_n 0.00176244f $X=1.575 $Y=0.815 $X2=0 $Y2=0
cc_322 N_D_M1015_g N_VGND_c_1814_n 9.27138e-19 $X=1.575 $Y=0.815 $X2=0 $Y2=0
cc_323 N_A_358_429#_M1009_g N_SCE_c_415_n 0.0103265f $X=1.935 $Y=0.815 $X2=0
+ $Y2=0
cc_324 N_A_358_429#_M1009_g N_SCE_M1026_g 0.0051197f $X=1.935 $Y=0.815 $X2=0
+ $Y2=0
cc_325 N_A_358_429#_c_342_n N_SCE_M1026_g 0.00755169f $X=2.96 $Y=1.555 $X2=0
+ $Y2=0
cc_326 N_A_358_429#_c_345_n N_SCE_M1026_g 0.00584673f $X=2.92 $Y=0.815 $X2=0
+ $Y2=0
cc_327 N_A_358_429#_c_345_n N_SCE_c_418_n 0.00415142f $X=2.92 $Y=0.815 $X2=0
+ $Y2=0
cc_328 N_A_358_429#_c_353_n N_SCE_c_426_n 0.00241891f $X=3.62 $Y=2.465 $X2=0
+ $Y2=0
cc_329 N_A_358_429#_c_345_n N_SCE_c_419_n 0.00489388f $X=2.92 $Y=0.815 $X2=0
+ $Y2=0
cc_330 N_A_358_429#_c_346_n N_SCE_c_419_n 0.010097f $X=3.535 $Y=1.665 $X2=0
+ $Y2=0
cc_331 N_A_358_429#_c_353_n N_SCE_c_419_n 0.010108f $X=3.62 $Y=2.465 $X2=0 $Y2=0
cc_332 N_A_358_429#_c_348_n N_SCE_c_419_n 0.012555f $X=3.125 $Y=1.555 $X2=0
+ $Y2=0
cc_333 N_A_358_429#_c_346_n N_SCE_c_429_n 0.00634697f $X=3.535 $Y=1.665 $X2=0
+ $Y2=0
cc_334 N_A_358_429#_c_353_n N_SCE_c_429_n 0.0134804f $X=3.62 $Y=2.465 $X2=0
+ $Y2=0
cc_335 N_A_358_429#_c_346_n N_SCE_c_422_n 5.42059e-19 $X=3.535 $Y=1.665 $X2=0
+ $Y2=0
cc_336 N_A_358_429#_c_345_n N_SCE_c_423_n 0.00265446f $X=2.92 $Y=0.815 $X2=0
+ $Y2=0
cc_337 N_A_358_429#_c_345_n N_SCE_c_424_n 0.0353441f $X=2.92 $Y=0.815 $X2=0
+ $Y2=0
cc_338 N_A_358_429#_c_346_n N_SCE_c_424_n 0.0286066f $X=3.535 $Y=1.665 $X2=0
+ $Y2=0
cc_339 N_A_358_429#_c_353_n N_CLK_M1020_g 0.00468876f $X=3.62 $Y=2.465 $X2=0
+ $Y2=0
cc_340 N_A_358_429#_c_346_n N_A_794_47#_c_974_n 0.0186505f $X=3.535 $Y=1.665
+ $X2=0 $Y2=0
cc_341 N_A_358_429#_c_353_n N_A_794_47#_c_974_n 0.0159778f $X=3.62 $Y=2.465
+ $X2=0 $Y2=0
cc_342 N_A_358_429#_c_353_n N_A_794_47#_c_990_n 0.0267005f $X=3.62 $Y=2.465
+ $X2=0 $Y2=0
cc_343 N_A_358_429#_c_350_n N_A_39_481#_c_1367_n 0.0135352f $X=1.9 $Y=2.295
+ $X2=0 $Y2=0
cc_344 N_A_358_429#_c_350_n N_VPWR_c_1400_n 0.00325902f $X=1.9 $Y=2.295 $X2=0
+ $Y2=0
cc_345 N_A_358_429#_c_350_n N_VPWR_c_1389_n 0.00595398f $X=1.9 $Y=2.295 $X2=0
+ $Y2=0
cc_346 N_A_358_429#_M1009_g N_A_244_121#_c_1575_n 0.00174772f $X=1.935 $Y=0.815
+ $X2=0 $Y2=0
cc_347 N_A_358_429#_c_350_n N_A_244_121#_c_1563_n 0.0132759f $X=1.9 $Y=2.295
+ $X2=0 $Y2=0
cc_348 N_A_358_429#_M1009_g N_A_244_121#_c_1559_n 0.0215609f $X=1.935 $Y=0.815
+ $X2=0 $Y2=0
cc_349 N_A_358_429#_c_342_n N_A_244_121#_c_1559_n 0.013279f $X=2.96 $Y=1.555
+ $X2=0 $Y2=0
cc_350 N_A_358_429#_c_345_n N_A_244_121#_c_1559_n 0.0203097f $X=2.92 $Y=0.815
+ $X2=0 $Y2=0
cc_351 N_A_358_429#_M1009_g N_A_244_121#_c_1561_n 0.00195541f $X=1.935 $Y=0.815
+ $X2=0 $Y2=0
cc_352 N_A_358_429#_c_342_n N_A_244_121#_c_1561_n 0.0184135f $X=2.96 $Y=1.555
+ $X2=0 $Y2=0
cc_353 N_A_358_429#_c_343_n N_A_244_121#_c_1561_n 0.00842938f $X=1.9 $Y=2.145
+ $X2=0 $Y2=0
cc_354 N_A_358_429#_c_345_n N_A_244_121#_c_1561_n 0.0097237f $X=2.92 $Y=0.815
+ $X2=0 $Y2=0
cc_355 N_A_358_429#_c_347_n N_A_244_121#_c_1561_n 0.0169541f $X=3.085 $Y=1.665
+ $X2=0 $Y2=0
cc_356 N_A_358_429#_c_348_n N_A_244_121#_c_1561_n 0.00161432f $X=3.125 $Y=1.555
+ $X2=0 $Y2=0
cc_357 N_A_358_429#_c_343_n N_A_244_121#_c_1565_n 4.19464e-19 $X=1.9 $Y=2.145
+ $X2=0 $Y2=0
cc_358 N_A_358_429#_c_350_n N_A_244_121#_c_1565_n 0.00773986f $X=1.9 $Y=2.295
+ $X2=0 $Y2=0
cc_359 N_A_358_429#_c_342_n N_A_244_121#_c_1566_n 0.00651116f $X=2.96 $Y=1.555
+ $X2=0 $Y2=0
cc_360 N_A_358_429#_c_346_n N_A_244_121#_c_1566_n 0.0222575f $X=3.535 $Y=1.665
+ $X2=0 $Y2=0
cc_361 N_A_358_429#_c_347_n N_A_244_121#_c_1566_n 0.0243045f $X=3.085 $Y=1.665
+ $X2=0 $Y2=0
cc_362 N_A_358_429#_c_353_n N_A_244_121#_c_1566_n 0.0141507f $X=3.62 $Y=2.465
+ $X2=0 $Y2=0
cc_363 N_A_358_429#_c_348_n N_A_244_121#_c_1566_n 0.00774857f $X=3.125 $Y=1.555
+ $X2=0 $Y2=0
cc_364 N_A_358_429#_c_353_n N_A_244_121#_c_1567_n 0.0244413f $X=3.62 $Y=2.465
+ $X2=0 $Y2=0
cc_365 N_A_358_429#_M1014_d N_A_244_121#_c_1568_n 0.00272304f $X=3.48 $Y=2.31
+ $X2=0 $Y2=0
cc_366 N_A_358_429#_c_353_n N_A_244_121#_c_1568_n 0.0192998f $X=3.62 $Y=2.465
+ $X2=0 $Y2=0
cc_367 N_A_358_429#_c_343_n N_A_244_121#_c_1572_n 7.8284e-19 $X=1.9 $Y=2.145
+ $X2=0 $Y2=0
cc_368 N_A_358_429#_c_353_n N_A_244_121#_c_1611_n 0.00597334f $X=3.62 $Y=2.465
+ $X2=0 $Y2=0
cc_369 N_A_358_429#_M1009_g N_VGND_c_1791_n 0.011862f $X=1.935 $Y=0.815 $X2=0
+ $Y2=0
cc_370 N_A_358_429#_c_342_n N_VGND_c_1791_n 0.00123976f $X=2.96 $Y=1.555 $X2=0
+ $Y2=0
cc_371 N_A_358_429#_c_345_n N_VGND_c_1807_n 0.00507875f $X=2.92 $Y=0.815 $X2=0
+ $Y2=0
cc_372 N_A_358_429#_M1009_g N_VGND_c_1814_n 7.78796e-19 $X=1.935 $Y=0.815 $X2=0
+ $Y2=0
cc_373 N_A_358_429#_c_345_n N_VGND_c_1814_n 0.00764386f $X=2.92 $Y=0.815 $X2=0
+ $Y2=0
cc_374 N_SCE_c_418_n N_CLK_M1010_g 0.00717511f $X=3.435 $Y=0.19 $X2=0 $Y2=0
cc_375 N_SCE_c_419_n N_CLK_M1020_g 0.00473751f $X=3.69 $Y=2.05 $X2=0 $Y2=0
cc_376 N_SCE_c_422_n N_CLK_c_500_n 0.00717511f $X=3.6 $Y=0.935 $X2=0 $Y2=0
cc_377 N_SCE_c_419_n N_CLK_c_504_n 0.00717511f $X=3.69 $Y=2.05 $X2=0 $Y2=0
cc_378 N_SCE_c_423_n N_CLK_c_502_n 0.00717511f $X=3.6 $Y=0.43 $X2=0 $Y2=0
cc_379 N_SCE_c_419_n N_A_794_47#_c_974_n 0.00163016f $X=3.69 $Y=2.05 $X2=0 $Y2=0
cc_380 N_SCE_c_422_n N_A_794_47#_c_974_n 0.00623631f $X=3.6 $Y=0.935 $X2=0 $Y2=0
cc_381 N_SCE_c_423_n N_A_794_47#_c_976_n 0.00623631f $X=3.6 $Y=0.43 $X2=0 $Y2=0
cc_382 N_SCE_c_424_n N_A_794_47#_c_976_n 0.0738436f $X=3.6 $Y=0.43 $X2=0 $Y2=0
cc_383 N_SCE_c_419_n N_A_794_47#_c_990_n 9.46006e-19 $X=3.69 $Y=2.05 $X2=0 $Y2=0
cc_384 N_SCE_M1017_g N_A_39_481#_c_1367_n 0.0140234f $X=0.965 $Y=2.725 $X2=0
+ $Y2=0
cc_385 N_SCE_M1017_g N_VPWR_c_1390_n 0.0087721f $X=0.965 $Y=2.725 $X2=0 $Y2=0
cc_386 N_SCE_c_426_n N_VPWR_c_1391_n 0.00698095f $X=3.405 $Y=2.2 $X2=0 $Y2=0
cc_387 N_SCE_M1017_g N_VPWR_c_1400_n 0.00325653f $X=0.965 $Y=2.725 $X2=0 $Y2=0
cc_388 N_SCE_c_426_n N_VPWR_c_1411_n 0.00405031f $X=3.405 $Y=2.2 $X2=0 $Y2=0
cc_389 N_SCE_M1017_g N_VPWR_c_1389_n 0.00392971f $X=0.965 $Y=2.725 $X2=0 $Y2=0
cc_390 N_SCE_c_426_n N_VPWR_c_1389_n 0.00542671f $X=3.405 $Y=2.2 $X2=0 $Y2=0
cc_391 N_SCE_M1011_g N_A_244_121#_c_1575_n 0.0103434f $X=1.145 $Y=0.815 $X2=0
+ $Y2=0
cc_392 N_SCE_c_415_n N_A_244_121#_c_1575_n 0.00340864f $X=2.63 $Y=0.19 $X2=0
+ $Y2=0
cc_393 N_SCE_M1011_g N_A_244_121#_c_1560_n 0.00847996f $X=1.145 $Y=0.815 $X2=0
+ $Y2=0
cc_394 N_SCE_c_419_n N_A_244_121#_c_1566_n 6.4911e-19 $X=3.69 $Y=2.05 $X2=0
+ $Y2=0
cc_395 N_SCE_c_429_n N_A_244_121#_c_1566_n 0.00354967f $X=3.69 $Y=2.125 $X2=0
+ $Y2=0
cc_396 N_SCE_c_426_n N_A_244_121#_c_1567_n 0.0220379f $X=3.405 $Y=2.2 $X2=0
+ $Y2=0
cc_397 N_SCE_c_429_n N_A_244_121#_c_1567_n 0.00267849f $X=3.69 $Y=2.125 $X2=0
+ $Y2=0
cc_398 N_SCE_c_426_n N_A_244_121#_c_1568_n 0.0119763f $X=3.405 $Y=2.2 $X2=0
+ $Y2=0
cc_399 N_SCE_c_429_n N_A_244_121#_c_1568_n 6.67519e-19 $X=3.69 $Y=2.125 $X2=0
+ $Y2=0
cc_400 N_SCE_c_426_n N_A_244_121#_c_1569_n 0.00379981f $X=3.405 $Y=2.2 $X2=0
+ $Y2=0
cc_401 N_SCE_c_426_n N_A_244_121#_c_1611_n 0.00373789f $X=3.405 $Y=2.2 $X2=0
+ $Y2=0
cc_402 N_SCE_M1011_g N_VGND_c_1790_n 0.00177594f $X=1.145 $Y=0.815 $X2=0 $Y2=0
cc_403 N_SCE_c_416_n N_VGND_c_1790_n 0.0102909f $X=1.22 $Y=0.19 $X2=0 $Y2=0
cc_404 N_SCE_c_415_n N_VGND_c_1791_n 0.0416955f $X=2.63 $Y=0.19 $X2=0 $Y2=0
cc_405 N_SCE_M1026_g N_VGND_c_1791_n 0.0149666f $X=2.705 $Y=0.815 $X2=0 $Y2=0
cc_406 N_SCE_c_416_n N_VGND_c_1806_n 0.029155f $X=1.22 $Y=0.19 $X2=0 $Y2=0
cc_407 N_SCE_c_415_n N_VGND_c_1807_n 0.0341729f $X=2.63 $Y=0.19 $X2=0 $Y2=0
cc_408 N_SCE_c_424_n N_VGND_c_1807_n 0.0209793f $X=3.6 $Y=0.43 $X2=0 $Y2=0
cc_409 N_SCE_c_415_n N_VGND_c_1814_n 0.028425f $X=2.63 $Y=0.19 $X2=0 $Y2=0
cc_410 N_SCE_c_416_n N_VGND_c_1814_n 0.0106621f $X=1.22 $Y=0.19 $X2=0 $Y2=0
cc_411 N_SCE_c_418_n N_VGND_c_1814_n 0.0378764f $X=3.435 $Y=0.19 $X2=0 $Y2=0
cc_412 N_SCE_c_421_n N_VGND_c_1814_n 0.00903659f $X=2.705 $Y=0.19 $X2=0 $Y2=0
cc_413 N_SCE_c_424_n N_VGND_c_1814_n 0.0111805f $X=3.6 $Y=0.43 $X2=0 $Y2=0
cc_414 N_CLK_M1010_g N_A_794_47#_c_968_n 0.0198743f $X=4.31 $Y=0.445 $X2=0 $Y2=0
cc_415 N_CLK_M1010_g N_A_794_47#_c_972_n 0.00582031f $X=4.31 $Y=0.445 $X2=0
+ $Y2=0
cc_416 CLK N_A_794_47#_c_972_n 0.0222832f $X=4.475 $Y=0.84 $X2=0 $Y2=0
cc_417 N_CLK_M1010_g N_A_794_47#_c_974_n 0.0136491f $X=4.31 $Y=0.445 $X2=0 $Y2=0
cc_418 N_CLK_M1020_g N_A_794_47#_c_974_n 0.00369244f $X=4.45 $Y=2.735 $X2=0
+ $Y2=0
cc_419 CLK N_A_794_47#_c_974_n 0.0792723f $X=4.475 $Y=0.84 $X2=0 $Y2=0
cc_420 N_CLK_M1020_g N_A_794_47#_c_988_n 0.0130439f $X=4.45 $Y=2.735 $X2=0 $Y2=0
cc_421 N_CLK_c_504_n N_A_794_47#_c_988_n 7.64656e-19 $X=4.4 $Y=1.825 $X2=0 $Y2=0
cc_422 CLK N_A_794_47#_c_988_n 0.0304231f $X=4.475 $Y=0.84 $X2=0 $Y2=0
cc_423 N_CLK_M1020_g N_A_794_47#_c_1009_n 9.5249e-19 $X=4.45 $Y=2.735 $X2=0
+ $Y2=0
cc_424 CLK N_A_794_47#_c_1009_n 0.0458771f $X=4.475 $Y=0.84 $X2=0 $Y2=0
cc_425 N_CLK_c_502_n N_A_794_47#_c_1009_n 5.42836e-19 $X=4.4 $Y=1.32 $X2=0 $Y2=0
cc_426 N_CLK_M1020_g N_A_794_47#_c_975_n 0.0472945f $X=4.45 $Y=2.735 $X2=0 $Y2=0
cc_427 N_CLK_c_502_n N_A_794_47#_c_975_n 0.0367636f $X=4.4 $Y=1.32 $X2=0 $Y2=0
cc_428 N_CLK_M1020_g N_A_794_47#_c_990_n 0.00561571f $X=4.45 $Y=2.735 $X2=0
+ $Y2=0
cc_429 N_CLK_c_504_n N_A_794_47#_c_990_n 0.00312973f $X=4.4 $Y=1.825 $X2=0 $Y2=0
cc_430 N_CLK_M1020_g N_VPWR_c_1392_n 0.0108967f $X=4.45 $Y=2.735 $X2=0 $Y2=0
cc_431 N_CLK_M1020_g N_VPWR_c_1411_n 0.0032999f $X=4.45 $Y=2.735 $X2=0 $Y2=0
cc_432 N_CLK_M1020_g N_VPWR_c_1389_n 0.00504806f $X=4.45 $Y=2.735 $X2=0 $Y2=0
cc_433 N_CLK_M1020_g N_A_244_121#_c_1623_n 0.012197f $X=4.45 $Y=2.735 $X2=0
+ $Y2=0
cc_434 N_CLK_M1020_g N_A_244_121#_c_1573_n 0.00322654f $X=4.45 $Y=2.735 $X2=0
+ $Y2=0
cc_435 N_CLK_M1010_g N_VGND_c_1792_n 0.0031247f $X=4.31 $Y=0.445 $X2=0 $Y2=0
cc_436 CLK N_VGND_c_1792_n 0.0186433f $X=4.475 $Y=0.84 $X2=0 $Y2=0
cc_437 N_CLK_c_502_n N_VGND_c_1792_n 5.26174e-19 $X=4.4 $Y=1.32 $X2=0 $Y2=0
cc_438 N_CLK_M1010_g N_VGND_c_1807_n 0.00585385f $X=4.31 $Y=0.445 $X2=0 $Y2=0
cc_439 N_CLK_M1010_g N_VGND_c_1814_n 0.0088715f $X=4.31 $Y=0.445 $X2=0 $Y2=0
cc_440 CLK N_VGND_c_1814_n 0.00536166f $X=4.475 $Y=0.84 $X2=0 $Y2=0
cc_441 N_A_963_47#_c_552_n N_A_1365_29#_M1005_g 0.00208785f $X=6.705 $Y=2.705
+ $X2=0 $Y2=0
cc_442 N_A_963_47#_c_553_n N_A_1365_29#_M1005_g 0.0151964f $X=7.48 $Y=2.02 $X2=0
+ $Y2=0
cc_443 N_A_963_47#_c_555_n N_A_1365_29#_M1005_g 0.00277946f $X=7.565 $Y=2.565
+ $X2=0 $Y2=0
cc_444 N_A_963_47#_c_545_n N_A_1365_29#_c_715_n 0.030163f $X=6.13 $Y=1.41 $X2=0
+ $Y2=0
cc_445 N_A_963_47#_M1035_g N_A_1365_29#_c_716_n 0.00113909f $X=6.54 $Y=0.485
+ $X2=0 $Y2=0
cc_446 N_A_963_47#_c_553_n N_A_1365_29#_c_717_n 0.0603749f $X=7.48 $Y=2.02 $X2=0
+ $Y2=0
cc_447 N_A_963_47#_c_560_n N_A_1365_29#_c_717_n 0.00267453f $X=8.35 $Y=1.82
+ $X2=0 $Y2=0
cc_448 N_A_963_47#_c_545_n N_A_1365_29#_c_717_n 5.6075e-19 $X=6.13 $Y=1.41 $X2=0
+ $Y2=0
cc_449 N_A_963_47#_M1029_g N_A_1365_29#_c_718_n 0.00259413f $X=6.13 $Y=2.285
+ $X2=0 $Y2=0
cc_450 N_A_963_47#_c_553_n N_A_1365_29#_c_718_n 0.00438376f $X=7.48 $Y=2.02
+ $X2=0 $Y2=0
cc_451 N_A_963_47#_c_553_n N_A_1365_29#_c_724_n 0.0125022f $X=7.48 $Y=2.02 $X2=0
+ $Y2=0
cc_452 N_A_963_47#_c_556_n N_A_1365_29#_c_724_n 0.0144371f $X=8.18 $Y=2.65 $X2=0
+ $Y2=0
cc_453 N_A_963_47#_c_558_n N_A_1365_29#_c_724_n 0.0339577f $X=8.265 $Y=2.565
+ $X2=0 $Y2=0
cc_454 N_A_963_47#_c_560_n N_A_1365_29#_c_724_n 0.0112262f $X=8.35 $Y=1.82 $X2=0
+ $Y2=0
cc_455 N_A_963_47#_M1035_g N_A_1365_29#_c_719_n 0.030163f $X=6.54 $Y=0.485 $X2=0
+ $Y2=0
cc_456 N_A_963_47#_c_545_n N_A_1365_29#_c_720_n 0.0298733f $X=6.13 $Y=1.41 $X2=0
+ $Y2=0
cc_457 N_A_963_47#_c_553_n N_A_1237_55#_M1040_g 0.00548785f $X=7.48 $Y=2.02
+ $X2=0 $Y2=0
cc_458 N_A_963_47#_c_555_n N_A_1237_55#_M1040_g 0.0123087f $X=7.565 $Y=2.565
+ $X2=0 $Y2=0
cc_459 N_A_963_47#_c_556_n N_A_1237_55#_M1040_g 0.00874058f $X=8.18 $Y=2.65
+ $X2=0 $Y2=0
cc_460 N_A_963_47#_c_557_n N_A_1237_55#_M1040_g 0.00117379f $X=7.65 $Y=2.65
+ $X2=0 $Y2=0
cc_461 N_A_963_47#_c_558_n N_A_1237_55#_M1040_g 0.00231522f $X=8.265 $Y=2.565
+ $X2=0 $Y2=0
cc_462 N_A_963_47#_c_558_n N_A_1237_55#_M1007_g 8.15145e-19 $X=8.265 $Y=2.565
+ $X2=0 $Y2=0
cc_463 N_A_963_47#_c_559_n N_A_1237_55#_M1007_g 0.0182659f $X=9.61 $Y=1.82 $X2=0
+ $Y2=0
cc_464 N_A_963_47#_c_565_n N_A_1237_55#_M1007_g 0.00510747f $X=9.95 $Y=1.93
+ $X2=0 $Y2=0
cc_465 N_A_963_47#_c_563_n N_A_1237_55#_c_779_n 0.00127635f $X=9.76 $Y=1.82
+ $X2=0 $Y2=0
cc_466 N_A_963_47#_c_565_n N_A_1237_55#_c_779_n 0.00310804f $X=9.95 $Y=1.93
+ $X2=0 $Y2=0
cc_467 N_A_963_47#_M1008_g N_A_1237_55#_c_780_n 0.0647377f $X=9.95 $Y=0.945
+ $X2=0 $Y2=0
cc_468 N_A_963_47#_c_544_n N_A_1237_55#_c_781_n 0.0340751f $X=5.985 $Y=1.375
+ $X2=0 $Y2=0
cc_469 N_A_963_47#_c_545_n N_A_1237_55#_c_781_n 0.00341259f $X=6.13 $Y=1.41
+ $X2=0 $Y2=0
cc_470 N_A_963_47#_M1029_g N_A_1237_55#_c_789_n 0.00358054f $X=6.13 $Y=2.285
+ $X2=0 $Y2=0
cc_471 N_A_963_47#_c_551_n N_A_1237_55#_c_789_n 0.00973275f $X=6.62 $Y=2.87
+ $X2=0 $Y2=0
cc_472 N_A_963_47#_c_554_n N_A_1237_55#_c_789_n 0.0125477f $X=6.79 $Y=2.02 $X2=0
+ $Y2=0
cc_473 N_A_963_47#_c_543_n N_A_1237_55#_c_789_n 0.057451f $X=5.995 $Y=1.54 $X2=0
+ $Y2=0
cc_474 N_A_963_47#_c_545_n N_A_1237_55#_c_789_n 0.017613f $X=6.13 $Y=1.41 $X2=0
+ $Y2=0
cc_475 N_A_963_47#_c_553_n N_A_1237_55#_c_783_n 0.0019087f $X=7.48 $Y=2.02 $X2=0
+ $Y2=0
cc_476 N_A_963_47#_c_554_n N_A_1237_55#_c_783_n 0.00665258f $X=6.79 $Y=2.02
+ $X2=0 $Y2=0
cc_477 N_A_963_47#_c_559_n N_A_1237_55#_c_783_n 0.0339104f $X=9.61 $Y=1.82 $X2=0
+ $Y2=0
cc_478 N_A_963_47#_c_560_n N_A_1237_55#_c_783_n 0.00834941f $X=8.35 $Y=1.82
+ $X2=0 $Y2=0
cc_479 N_A_963_47#_c_545_n N_A_1237_55#_c_783_n 0.0151956f $X=6.13 $Y=1.41 $X2=0
+ $Y2=0
cc_480 N_A_963_47#_M1035_g N_A_1237_55#_c_784_n 0.00568774f $X=6.54 $Y=0.485
+ $X2=0 $Y2=0
cc_481 N_A_963_47#_c_544_n N_A_1237_55#_c_784_n 0.0106904f $X=5.985 $Y=1.375
+ $X2=0 $Y2=0
cc_482 N_A_963_47#_c_545_n N_A_1237_55#_c_784_n 4.73118e-19 $X=6.13 $Y=1.41
+ $X2=0 $Y2=0
cc_483 N_A_963_47#_c_543_n N_A_1237_55#_c_785_n 0.00309201f $X=5.995 $Y=1.54
+ $X2=0 $Y2=0
cc_484 N_A_963_47#_c_544_n N_A_1237_55#_c_785_n 0.0117635f $X=5.985 $Y=1.375
+ $X2=0 $Y2=0
cc_485 N_A_963_47#_c_545_n N_A_1237_55#_c_785_n 0.00925348f $X=6.13 $Y=1.41
+ $X2=0 $Y2=0
cc_486 N_A_963_47#_c_559_n N_A_1237_55#_c_786_n 0.0233111f $X=9.61 $Y=1.82 $X2=0
+ $Y2=0
cc_487 N_A_963_47#_c_555_n N_SET_B_M1004_g 2.43971e-19 $X=7.565 $Y=2.565 $X2=0
+ $Y2=0
cc_488 N_A_963_47#_c_556_n N_SET_B_M1004_g 8.41666e-19 $X=8.18 $Y=2.65 $X2=0
+ $Y2=0
cc_489 N_A_963_47#_c_558_n N_SET_B_M1004_g 0.0156167f $X=8.265 $Y=2.565 $X2=0
+ $Y2=0
cc_490 N_A_963_47#_c_560_n N_SET_B_M1004_g 0.00764192f $X=8.35 $Y=1.82 $X2=0
+ $Y2=0
cc_491 N_A_963_47#_c_559_n N_SET_B_c_875_n 0.00163921f $X=9.61 $Y=1.82 $X2=0
+ $Y2=0
cc_492 N_A_963_47#_c_560_n N_SET_B_c_875_n 0.00174463f $X=8.35 $Y=1.82 $X2=0
+ $Y2=0
cc_493 N_A_963_47#_M1008_g N_SET_B_c_879_n 0.00645726f $X=9.95 $Y=0.945 $X2=0
+ $Y2=0
cc_494 N_A_963_47#_M1008_g SET_B 0.0115181f $X=9.95 $Y=0.945 $X2=0 $Y2=0
cc_495 N_A_963_47#_c_549_n N_A_794_47#_c_978_n 0.0188966f $X=5.91 $Y=2.87 $X2=0
+ $Y2=0
cc_496 N_A_963_47#_c_550_n N_A_794_47#_c_978_n 0.00368206f $X=6 $Y=2.705 $X2=0
+ $Y2=0
cc_497 N_A_963_47#_c_541_n N_A_794_47#_c_969_n 0.00388743f $X=5.88 $Y=0.34 $X2=0
+ $Y2=0
cc_498 N_A_963_47#_c_544_n N_A_794_47#_c_969_n 0.00940023f $X=5.985 $Y=1.375
+ $X2=0 $Y2=0
cc_499 N_A_963_47#_c_545_n N_A_794_47#_c_969_n 0.0228489f $X=6.13 $Y=1.41 $X2=0
+ $Y2=0
cc_500 N_A_963_47#_M1029_g N_A_794_47#_c_979_n 0.00293414f $X=6.13 $Y=2.285
+ $X2=0 $Y2=0
cc_501 N_A_963_47#_c_549_n N_A_794_47#_c_979_n 0.0088166f $X=5.91 $Y=2.87 $X2=0
+ $Y2=0
cc_502 N_A_963_47#_c_551_n N_A_794_47#_c_979_n 0.00567699f $X=6.62 $Y=2.87 $X2=0
+ $Y2=0
cc_503 N_A_963_47#_c_562_n N_A_794_47#_c_979_n 0.00392429f $X=6 $Y=2.87 $X2=0
+ $Y2=0
cc_504 N_A_963_47#_M1035_g N_A_794_47#_M1034_g 0.0229717f $X=6.54 $Y=0.485 $X2=0
+ $Y2=0
cc_505 N_A_963_47#_c_541_n N_A_794_47#_M1034_g 0.0068961f $X=5.88 $Y=0.34 $X2=0
+ $Y2=0
cc_506 N_A_963_47#_c_544_n N_A_794_47#_M1034_g 0.0159315f $X=5.985 $Y=1.375
+ $X2=0 $Y2=0
cc_507 N_A_963_47#_M1029_g N_A_794_47#_M1001_g 0.0130279f $X=6.13 $Y=2.285 $X2=0
+ $Y2=0
cc_508 N_A_963_47#_c_550_n N_A_794_47#_M1001_g 0.00217035f $X=6 $Y=2.705 $X2=0
+ $Y2=0
cc_509 N_A_963_47#_c_551_n N_A_794_47#_M1001_g 0.0262197f $X=6.62 $Y=2.87 $X2=0
+ $Y2=0
cc_510 N_A_963_47#_c_552_n N_A_794_47#_M1001_g 0.0125562f $X=6.705 $Y=2.705
+ $X2=0 $Y2=0
cc_511 N_A_963_47#_c_554_n N_A_794_47#_M1001_g 0.00317217f $X=6.79 $Y=2.02 $X2=0
+ $Y2=0
cc_512 N_A_963_47#_c_545_n N_A_794_47#_M1001_g 0.00678246f $X=6.13 $Y=1.41 $X2=0
+ $Y2=0
cc_513 N_A_963_47#_M1032_g N_A_794_47#_c_982_n 0.00884409f $X=9.915 $Y=2.525
+ $X2=0 $Y2=0
cc_514 N_A_963_47#_c_551_n N_A_794_47#_c_982_n 0.00158131f $X=6.62 $Y=2.87 $X2=0
+ $Y2=0
cc_515 N_A_963_47#_c_556_n N_A_794_47#_c_982_n 0.0104196f $X=8.18 $Y=2.65 $X2=0
+ $Y2=0
cc_516 N_A_963_47#_c_557_n N_A_794_47#_c_982_n 0.0031402f $X=7.65 $Y=2.65 $X2=0
+ $Y2=0
cc_517 N_A_963_47#_M1032_g N_A_794_47#_c_983_n 0.0225271f $X=9.915 $Y=2.525
+ $X2=0 $Y2=0
cc_518 N_A_963_47#_c_565_n N_A_794_47#_c_983_n 0.00520955f $X=9.95 $Y=1.93 $X2=0
+ $Y2=0
cc_519 N_A_963_47#_M1008_g N_A_794_47#_M1002_g 0.0109557f $X=9.95 $Y=0.945 $X2=0
+ $Y2=0
cc_520 N_A_963_47#_c_541_n N_A_794_47#_c_972_n 0.00824725f $X=5.88 $Y=0.34 $X2=0
+ $Y2=0
cc_521 N_A_963_47#_c_542_n N_A_794_47#_c_972_n 0.00572067f $X=4.972 $Y=0.34
+ $X2=0 $Y2=0
cc_522 N_A_963_47#_M1008_g N_A_794_47#_c_973_n 0.00520955f $X=9.95 $Y=0.945
+ $X2=0 $Y2=0
cc_523 N_A_963_47#_c_542_n N_A_794_47#_c_1009_n 0.00748769f $X=4.972 $Y=0.34
+ $X2=0 $Y2=0
cc_524 N_A_963_47#_M1029_g N_A_794_47#_c_975_n 0.0121016f $X=6.13 $Y=2.285 $X2=0
+ $Y2=0
cc_525 N_A_963_47#_c_550_n N_A_794_47#_c_975_n 0.00177117f $X=6 $Y=2.705 $X2=0
+ $Y2=0
cc_526 N_A_963_47#_c_543_n N_A_794_47#_c_975_n 2.65069e-19 $X=5.995 $Y=1.54
+ $X2=0 $Y2=0
cc_527 N_A_963_47#_c_544_n N_A_794_47#_c_975_n 5.82401e-19 $X=5.985 $Y=1.375
+ $X2=0 $Y2=0
cc_528 N_A_963_47#_c_545_n N_A_794_47#_c_975_n 0.0095402f $X=6.13 $Y=1.41 $X2=0
+ $Y2=0
cc_529 N_A_963_47#_M1032_g N_A_1998_463#_c_1211_n 3.11481e-19 $X=9.915 $Y=2.525
+ $X2=0 $Y2=0
cc_530 N_A_963_47#_c_563_n N_A_1998_463#_c_1211_n 0.0150666f $X=9.76 $Y=1.82
+ $X2=0 $Y2=0
cc_531 N_A_963_47#_c_565_n N_A_1998_463#_c_1211_n 0.00188233f $X=9.95 $Y=1.93
+ $X2=0 $Y2=0
cc_532 N_A_963_47#_M1008_g N_A_1998_463#_c_1204_n 0.0317911f $X=9.95 $Y=0.945
+ $X2=0 $Y2=0
cc_533 N_A_963_47#_c_563_n N_A_1998_463#_c_1204_n 0.0138743f $X=9.76 $Y=1.82
+ $X2=0 $Y2=0
cc_534 N_A_963_47#_c_553_n N_VPWR_M1005_d 0.0096518f $X=7.48 $Y=2.02 $X2=0 $Y2=0
cc_535 N_A_963_47#_c_555_n N_VPWR_M1005_d 0.00464265f $X=7.565 $Y=2.565 $X2=0
+ $Y2=0
cc_536 N_A_963_47#_c_559_n N_VPWR_M1004_d 0.00818638f $X=9.61 $Y=1.82 $X2=0
+ $Y2=0
cc_537 N_A_963_47#_c_551_n N_VPWR_c_1393_n 0.0269813f $X=6.62 $Y=2.87 $X2=0
+ $Y2=0
cc_538 N_A_963_47#_c_552_n N_VPWR_c_1393_n 0.022331f $X=6.705 $Y=2.705 $X2=0
+ $Y2=0
cc_539 N_A_963_47#_c_553_n N_VPWR_c_1393_n 0.0219335f $X=7.48 $Y=2.02 $X2=0
+ $Y2=0
cc_540 N_A_963_47#_c_555_n N_VPWR_c_1393_n 0.0223246f $X=7.565 $Y=2.565 $X2=0
+ $Y2=0
cc_541 N_A_963_47#_c_557_n N_VPWR_c_1393_n 0.0150381f $X=7.65 $Y=2.65 $X2=0
+ $Y2=0
cc_542 N_A_963_47#_c_556_n N_VPWR_c_1394_n 0.0143976f $X=8.18 $Y=2.65 $X2=0
+ $Y2=0
cc_543 N_A_963_47#_c_558_n N_VPWR_c_1394_n 0.027895f $X=8.265 $Y=2.565 $X2=0
+ $Y2=0
cc_544 N_A_963_47#_c_559_n N_VPWR_c_1394_n 0.0144005f $X=9.61 $Y=1.82 $X2=0
+ $Y2=0
cc_545 N_A_963_47#_c_549_n N_VPWR_c_1402_n 0.0480741f $X=5.91 $Y=2.87 $X2=0
+ $Y2=0
cc_546 N_A_963_47#_c_551_n N_VPWR_c_1402_n 0.0378038f $X=6.62 $Y=2.87 $X2=0
+ $Y2=0
cc_547 N_A_963_47#_c_562_n N_VPWR_c_1402_n 0.010285f $X=6 $Y=2.87 $X2=0 $Y2=0
cc_548 N_A_963_47#_c_556_n N_VPWR_c_1404_n 0.0142546f $X=8.18 $Y=2.65 $X2=0
+ $Y2=0
cc_549 N_A_963_47#_c_557_n N_VPWR_c_1404_n 0.00374304f $X=7.65 $Y=2.65 $X2=0
+ $Y2=0
cc_550 N_A_963_47#_c_549_n N_VPWR_c_1389_n 0.0313535f $X=5.91 $Y=2.87 $X2=0
+ $Y2=0
cc_551 N_A_963_47#_c_551_n N_VPWR_c_1389_n 0.0232827f $X=6.62 $Y=2.87 $X2=0
+ $Y2=0
cc_552 N_A_963_47#_c_556_n N_VPWR_c_1389_n 0.0181537f $X=8.18 $Y=2.65 $X2=0
+ $Y2=0
cc_553 N_A_963_47#_c_557_n N_VPWR_c_1389_n 0.00464028f $X=7.65 $Y=2.65 $X2=0
+ $Y2=0
cc_554 N_A_963_47#_c_562_n N_VPWR_c_1389_n 0.00613933f $X=6 $Y=2.87 $X2=0 $Y2=0
cc_555 N_A_963_47#_c_541_n N_A_244_121#_M1034_s 0.00948205f $X=5.88 $Y=0.34
+ $X2=0 $Y2=0
cc_556 N_A_963_47#_c_544_n N_A_244_121#_M1034_s 0.00760501f $X=5.985 $Y=1.375
+ $X2=0 $Y2=0
cc_557 N_A_963_47#_c_550_n N_A_244_121#_M1029_s 0.00400815f $X=6 $Y=2.705 $X2=0
+ $Y2=0
cc_558 N_A_963_47#_M1000_d N_A_244_121#_c_1570_n 0.00223155f $X=4.955 $Y=2.415
+ $X2=0 $Y2=0
cc_559 N_A_963_47#_c_549_n N_A_244_121#_c_1570_n 0.0259001f $X=5.91 $Y=2.87
+ $X2=0 $Y2=0
cc_560 N_A_963_47#_M1029_g N_A_244_121#_c_1562_n 0.00152292f $X=6.13 $Y=2.285
+ $X2=0 $Y2=0
cc_561 N_A_963_47#_c_541_n N_A_244_121#_c_1562_n 0.0250201f $X=5.88 $Y=0.34
+ $X2=0 $Y2=0
cc_562 N_A_963_47#_c_550_n N_A_244_121#_c_1562_n 0.0336923f $X=6 $Y=2.705 $X2=0
+ $Y2=0
cc_563 N_A_963_47#_c_542_n N_A_244_121#_c_1562_n 9.21522e-19 $X=4.972 $Y=0.34
+ $X2=0 $Y2=0
cc_564 N_A_963_47#_c_544_n N_A_244_121#_c_1562_n 0.0859113f $X=5.985 $Y=1.375
+ $X2=0 $Y2=0
cc_565 N_A_963_47#_c_545_n N_A_244_121#_c_1562_n 0.00322854f $X=6.13 $Y=1.41
+ $X2=0 $Y2=0
cc_566 N_A_963_47#_M1029_g N_A_244_121#_c_1574_n 0.00106064f $X=6.13 $Y=2.285
+ $X2=0 $Y2=0
cc_567 N_A_963_47#_c_549_n N_A_244_121#_c_1574_n 0.0286986f $X=5.91 $Y=2.87
+ $X2=0 $Y2=0
cc_568 N_A_963_47#_c_550_n N_A_244_121#_c_1574_n 0.0263548f $X=6 $Y=2.705 $X2=0
+ $Y2=0
cc_569 N_A_963_47#_c_559_n N_A_1781_379#_M1007_d 0.00225342f $X=9.61 $Y=1.82
+ $X2=-0.19 $Y2=-0.245
cc_570 N_A_963_47#_M1032_g N_A_1781_379#_c_1697_n 0.0163226f $X=9.915 $Y=2.525
+ $X2=0 $Y2=0
cc_571 N_A_963_47#_c_559_n N_A_1781_379#_c_1697_n 0.0175973f $X=9.61 $Y=1.82
+ $X2=0 $Y2=0
cc_572 N_A_963_47#_c_563_n N_A_1781_379#_c_1697_n 0.0214354f $X=9.76 $Y=1.82
+ $X2=0 $Y2=0
cc_573 N_A_963_47#_c_565_n N_A_1781_379#_c_1697_n 0.00303148f $X=9.95 $Y=1.93
+ $X2=0 $Y2=0
cc_574 N_A_963_47#_M1032_g N_A_1781_379#_c_1698_n 0.00847934f $X=9.915 $Y=2.525
+ $X2=0 $Y2=0
cc_575 N_A_963_47#_c_559_n N_A_1781_379#_c_1698_n 0.0202165f $X=9.61 $Y=1.82
+ $X2=0 $Y2=0
cc_576 N_A_963_47#_c_563_n N_A_1781_379#_c_1698_n 8.24085e-19 $X=9.76 $Y=1.82
+ $X2=0 $Y2=0
cc_577 N_A_963_47#_M1032_g N_A_1781_379#_c_1700_n 8.68604e-19 $X=9.915 $Y=2.525
+ $X2=0 $Y2=0
cc_578 N_A_963_47#_M1032_g N_A_1888_463#_c_1733_n 0.00681915f $X=9.915 $Y=2.525
+ $X2=0 $Y2=0
cc_579 N_A_963_47#_M1032_g N_A_1888_463#_c_1735_n 0.00780991f $X=9.915 $Y=2.525
+ $X2=0 $Y2=0
cc_580 N_A_963_47#_M1035_g N_VGND_c_1793_n 0.00189234f $X=6.54 $Y=0.485 $X2=0
+ $Y2=0
cc_581 N_A_963_47#_M1008_g N_VGND_c_1846_n 5.64369e-19 $X=9.95 $Y=0.945 $X2=0
+ $Y2=0
cc_582 N_A_963_47#_M1008_g N_VGND_c_1801_n 5.58455e-19 $X=9.95 $Y=0.945 $X2=0
+ $Y2=0
cc_583 N_A_963_47#_M1035_g N_VGND_c_1808_n 0.00545548f $X=6.54 $Y=0.485 $X2=0
+ $Y2=0
cc_584 N_A_963_47#_c_541_n N_VGND_c_1808_n 0.0624262f $X=5.88 $Y=0.34 $X2=0
+ $Y2=0
cc_585 N_A_963_47#_c_542_n N_VGND_c_1808_n 0.0182557f $X=4.972 $Y=0.34 $X2=0
+ $Y2=0
cc_586 N_A_963_47#_M1023_d N_VGND_c_1814_n 0.00228875f $X=4.815 $Y=0.235 $X2=0
+ $Y2=0
cc_587 N_A_963_47#_M1035_g N_VGND_c_1814_n 0.0104387f $X=6.54 $Y=0.485 $X2=0
+ $Y2=0
cc_588 N_A_963_47#_c_541_n N_VGND_c_1814_n 0.0357969f $X=5.88 $Y=0.34 $X2=0
+ $Y2=0
cc_589 N_A_963_47#_c_542_n N_VGND_c_1814_n 0.0112074f $X=4.972 $Y=0.34 $X2=0
+ $Y2=0
cc_590 N_A_1365_29#_M1005_g N_A_1237_55#_M1040_g 0.00891656f $X=6.92 $Y=2.285
+ $X2=0 $Y2=0
cc_591 N_A_1365_29#_c_717_n N_A_1237_55#_M1040_g 0.0154284f $X=7.82 $Y=1.675
+ $X2=0 $Y2=0
cc_592 N_A_1365_29#_c_718_n N_A_1237_55#_M1040_g 0.00909063f $X=7.01 $Y=1.67
+ $X2=0 $Y2=0
cc_593 N_A_1365_29#_c_724_n N_A_1237_55#_M1040_g 0.00556189f $X=7.915 $Y=2.22
+ $X2=0 $Y2=0
cc_594 N_A_1365_29#_c_720_n N_A_1237_55#_M1040_g 4.5701e-19 $X=7.01 $Y=1.505
+ $X2=0 $Y2=0
cc_595 N_A_1365_29#_c_716_n N_A_1237_55#_c_777_n 0.00232423f $X=7.71 $Y=0.89
+ $X2=0 $Y2=0
cc_596 N_A_1365_29#_c_716_n N_A_1237_55#_c_781_n 0.013835f $X=7.71 $Y=0.89 $X2=0
+ $Y2=0
cc_597 N_A_1365_29#_c_720_n N_A_1237_55#_c_781_n 3.98673e-19 $X=7.01 $Y=1.505
+ $X2=0 $Y2=0
cc_598 N_A_1365_29#_c_717_n N_A_1237_55#_c_789_n 0.00713994f $X=7.82 $Y=1.675
+ $X2=0 $Y2=0
cc_599 N_A_1365_29#_c_718_n N_A_1237_55#_c_789_n 0.00360078f $X=7.01 $Y=1.67
+ $X2=0 $Y2=0
cc_600 N_A_1365_29#_c_720_n N_A_1237_55#_c_789_n 8.73008e-19 $X=7.01 $Y=1.505
+ $X2=0 $Y2=0
cc_601 N_A_1365_29#_c_716_n N_A_1237_55#_c_782_n 0.0059635f $X=7.71 $Y=0.89
+ $X2=0 $Y2=0
cc_602 N_A_1365_29#_c_717_n N_A_1237_55#_c_782_n 0.00515594f $X=7.82 $Y=1.675
+ $X2=0 $Y2=0
cc_603 N_A_1365_29#_c_720_n N_A_1237_55#_c_782_n 0.00664958f $X=7.01 $Y=1.505
+ $X2=0 $Y2=0
cc_604 N_A_1365_29#_c_715_n N_A_1237_55#_c_783_n 0.00195978f $X=6.99 $Y=0.97
+ $X2=0 $Y2=0
cc_605 N_A_1365_29#_c_716_n N_A_1237_55#_c_783_n 0.0747694f $X=7.71 $Y=0.89
+ $X2=0 $Y2=0
cc_606 N_A_1365_29#_c_717_n N_A_1237_55#_c_783_n 0.0868362f $X=7.82 $Y=1.675
+ $X2=0 $Y2=0
cc_607 N_A_1365_29#_c_718_n N_A_1237_55#_c_783_n 0.00187382f $X=7.01 $Y=1.67
+ $X2=0 $Y2=0
cc_608 N_A_1365_29#_c_720_n N_A_1237_55#_c_783_n 0.0124359f $X=7.01 $Y=1.505
+ $X2=0 $Y2=0
cc_609 N_A_1365_29#_c_724_n N_SET_B_M1004_g 0.00431365f $X=7.915 $Y=2.22 $X2=0
+ $Y2=0
cc_610 N_A_1365_29#_c_717_n N_SET_B_c_875_n 0.00472792f $X=7.82 $Y=1.675 $X2=0
+ $Y2=0
cc_611 N_A_1365_29#_M1005_g N_A_794_47#_M1001_g 0.0405493f $X=6.92 $Y=2.285
+ $X2=0 $Y2=0
cc_612 N_A_1365_29#_M1005_g N_A_794_47#_c_982_n 0.00461292f $X=6.92 $Y=2.285
+ $X2=0 $Y2=0
cc_613 N_A_1365_29#_M1005_g N_VPWR_c_1393_n 0.00596035f $X=6.92 $Y=2.285 $X2=0
+ $Y2=0
cc_614 N_A_1365_29#_M1005_g N_VPWR_c_1389_n 8.80648e-19 $X=6.92 $Y=2.285 $X2=0
+ $Y2=0
cc_615 N_A_1365_29#_c_715_n N_VGND_c_1793_n 0.00100313f $X=6.99 $Y=0.97 $X2=0
+ $Y2=0
cc_616 N_A_1365_29#_c_716_n N_VGND_c_1793_n 0.0246094f $X=7.71 $Y=0.89 $X2=0
+ $Y2=0
cc_617 N_A_1365_29#_c_719_n N_VGND_c_1793_n 0.0108244f $X=6.99 $Y=0.805 $X2=0
+ $Y2=0
cc_618 N_A_1365_29#_c_716_n N_VGND_c_1794_n 0.00659607f $X=7.71 $Y=0.89 $X2=0
+ $Y2=0
cc_619 N_A_1365_29#_c_716_n N_VGND_c_1859_n 0.0174807f $X=7.71 $Y=0.89 $X2=0
+ $Y2=0
cc_620 N_A_1365_29#_c_716_n N_VGND_c_1799_n 0.00805088f $X=7.71 $Y=0.89 $X2=0
+ $Y2=0
cc_621 N_A_1365_29#_c_716_n N_VGND_c_1808_n 0.00173759f $X=7.71 $Y=0.89 $X2=0
+ $Y2=0
cc_622 N_A_1365_29#_c_719_n N_VGND_c_1808_n 0.00336323f $X=6.99 $Y=0.805 $X2=0
+ $Y2=0
cc_623 N_A_1365_29#_c_716_n N_VGND_c_1814_n 0.0183081f $X=7.71 $Y=0.89 $X2=0
+ $Y2=0
cc_624 N_A_1365_29#_c_719_n N_VGND_c_1814_n 0.00405306f $X=6.99 $Y=0.805 $X2=0
+ $Y2=0
cc_625 N_A_1237_55#_M1007_g N_SET_B_M1004_g 0.0126691f $X=8.83 $Y=2.315 $X2=0
+ $Y2=0
cc_626 N_A_1237_55#_M1040_g N_SET_B_M1027_g 0.00185333f $X=7.7 $Y=2.285 $X2=0
+ $Y2=0
cc_627 N_A_1237_55#_c_782_n N_SET_B_M1027_g 0.0325118f $X=7.745 $Y=1.32 $X2=0
+ $Y2=0
cc_628 N_A_1237_55#_c_783_n N_SET_B_M1027_g 0.012359f $X=8.92 $Y=1.32 $X2=0
+ $Y2=0
cc_629 N_A_1237_55#_c_786_n N_SET_B_M1027_g 0.0108203f $X=9.085 $Y=1.34 $X2=0
+ $Y2=0
cc_630 N_A_1237_55#_M1040_g N_SET_B_c_875_n 0.0185313f $X=7.7 $Y=2.285 $X2=0
+ $Y2=0
cc_631 N_A_1237_55#_M1007_g N_SET_B_c_875_n 0.0108203f $X=8.83 $Y=2.315 $X2=0
+ $Y2=0
cc_632 N_A_1237_55#_c_783_n N_SET_B_c_875_n 0.0033816f $X=8.92 $Y=1.32 $X2=0
+ $Y2=0
cc_633 N_A_1237_55#_c_777_n N_SET_B_c_881_n 0.0254737f $X=7.965 $Y=1.155 $X2=0
+ $Y2=0
cc_634 N_A_1237_55#_c_780_n N_SET_B_c_882_n 0.0160442f $X=9.59 $Y=1.375 $X2=0
+ $Y2=0
cc_635 N_A_1237_55#_c_781_n N_A_794_47#_M1034_g 0.00317354f $X=6.345 $Y=1.225
+ $X2=0 $Y2=0
cc_636 N_A_1237_55#_c_789_n N_A_794_47#_M1001_g 9.52094e-19 $X=6.345 $Y=2.22
+ $X2=0 $Y2=0
cc_637 N_A_1237_55#_c_783_n N_A_794_47#_M1001_g 0.00132099f $X=8.92 $Y=1.32
+ $X2=0 $Y2=0
cc_638 N_A_1237_55#_M1040_g N_A_794_47#_c_982_n 0.00324269f $X=7.7 $Y=2.285
+ $X2=0 $Y2=0
cc_639 N_A_1237_55#_M1007_g N_A_794_47#_c_982_n 0.0104164f $X=8.83 $Y=2.315
+ $X2=0 $Y2=0
cc_640 N_A_1237_55#_M1040_g N_VPWR_c_1393_n 0.00109199f $X=7.7 $Y=2.285 $X2=0
+ $Y2=0
cc_641 N_A_1237_55#_M1007_g N_VPWR_c_1394_n 0.00381353f $X=8.83 $Y=2.315 $X2=0
+ $Y2=0
cc_642 N_A_1237_55#_M1007_g N_VPWR_c_1389_n 9.39239e-19 $X=8.83 $Y=2.315 $X2=0
+ $Y2=0
cc_643 N_A_1237_55#_M1007_g N_A_1781_379#_c_1699_n 4.68635e-19 $X=8.83 $Y=2.315
+ $X2=0 $Y2=0
cc_644 N_A_1237_55#_M1007_g N_A_1888_463#_c_1735_n 0.00203475f $X=8.83 $Y=2.315
+ $X2=0 $Y2=0
cc_645 N_A_1237_55#_c_777_n N_VGND_c_1793_n 0.00141034f $X=7.965 $Y=1.155 $X2=0
+ $Y2=0
cc_646 N_A_1237_55#_c_777_n N_VGND_c_1794_n 0.014455f $X=7.965 $Y=1.155 $X2=0
+ $Y2=0
cc_647 N_A_1237_55#_c_777_n N_VGND_c_1859_n 0.00582867f $X=7.965 $Y=1.155 $X2=0
+ $Y2=0
cc_648 N_A_1237_55#_c_783_n N_VGND_c_1859_n 0.00922256f $X=8.92 $Y=1.32 $X2=0
+ $Y2=0
cc_649 N_A_1237_55#_c_779_n N_VGND_c_1846_n 0.00709255f $X=9.515 $Y=1.45 $X2=0
+ $Y2=0
cc_650 N_A_1237_55#_c_780_n N_VGND_c_1846_n 0.00482276f $X=9.59 $Y=1.375 $X2=0
+ $Y2=0
cc_651 N_A_1237_55#_c_783_n N_VGND_c_1846_n 0.0547f $X=8.92 $Y=1.32 $X2=0 $Y2=0
cc_652 N_A_1237_55#_c_786_n N_VGND_c_1846_n 0.00854365f $X=9.085 $Y=1.34 $X2=0
+ $Y2=0
cc_653 N_A_1237_55#_c_777_n N_VGND_c_1799_n 0.00206768f $X=7.965 $Y=1.155 $X2=0
+ $Y2=0
cc_654 N_A_1237_55#_c_780_n N_VGND_c_1801_n 5.42344e-19 $X=9.59 $Y=1.375 $X2=0
+ $Y2=0
cc_655 N_A_1237_55#_c_869_p N_VGND_c_1808_n 0.00854685f $X=6.325 $Y=0.49 $X2=0
+ $Y2=0
cc_656 N_A_1237_55#_c_777_n N_VGND_c_1814_n 0.00237845f $X=7.965 $Y=1.155 $X2=0
+ $Y2=0
cc_657 N_A_1237_55#_c_869_p N_VGND_c_1814_n 0.0070283f $X=6.325 $Y=0.49 $X2=0
+ $Y2=0
cc_658 N_SET_B_M1004_g N_A_794_47#_c_982_n 0.00180597f $X=8.225 $Y=2.105 $X2=0
+ $Y2=0
cc_659 N_SET_B_c_876_n N_A_794_47#_M1002_g 0.0106546f $X=10.955 $Y=1.585 $X2=0
+ $Y2=0
cc_660 N_SET_B_c_877_n N_A_794_47#_M1002_g 5.4374e-19 $X=11.04 $Y=1.675 $X2=0
+ $Y2=0
cc_661 N_SET_B_c_879_n N_A_794_47#_M1002_g 0.00805153f $X=10.87 $Y=0.382 $X2=0
+ $Y2=0
cc_662 N_SET_B_c_877_n N_A_794_47#_c_973_n 0.0116151f $X=11.04 $Y=1.675 $X2=0
+ $Y2=0
cc_663 N_SET_B_M1019_g N_A_2214_99#_c_1137_n 0.0160696f $X=11.835 $Y=0.835 $X2=0
+ $Y2=0
cc_664 N_SET_B_c_876_n N_A_2214_99#_c_1137_n 0.0102441f $X=10.955 $Y=1.585 $X2=0
+ $Y2=0
cc_665 N_SET_B_c_874_n N_A_2214_99#_M1025_g 0.0199052f $X=11.87 $Y=1.835 $X2=0
+ $Y2=0
cc_666 N_SET_B_M1012_g N_A_2214_99#_M1025_g 0.0236755f $X=11.87 $Y=2.385 $X2=0
+ $Y2=0
cc_667 N_SET_B_c_876_n N_A_2214_99#_M1025_g 0.00191246f $X=10.955 $Y=1.585 $X2=0
+ $Y2=0
cc_668 N_SET_B_c_878_n N_A_2214_99#_M1025_g 0.0111504f $X=11.925 $Y=1.67 $X2=0
+ $Y2=0
cc_669 N_SET_B_M1019_g N_A_2214_99#_c_1139_n 0.00974063f $X=11.835 $Y=0.835
+ $X2=0 $Y2=0
cc_670 N_SET_B_c_874_n N_A_2214_99#_c_1139_n 0.00985513f $X=11.87 $Y=1.835 $X2=0
+ $Y2=0
cc_671 N_SET_B_c_876_n N_A_2214_99#_c_1139_n 0.0136188f $X=10.955 $Y=1.585 $X2=0
+ $Y2=0
cc_672 N_SET_B_c_878_n N_A_2214_99#_c_1139_n 0.0623244f $X=11.925 $Y=1.67 $X2=0
+ $Y2=0
cc_673 N_SET_B_M1019_g N_A_2214_99#_c_1140_n 0.0223851f $X=11.835 $Y=0.835 $X2=0
+ $Y2=0
cc_674 N_SET_B_c_876_n N_A_2214_99#_c_1140_n 0.00200868f $X=10.955 $Y=1.585
+ $X2=0 $Y2=0
cc_675 N_SET_B_c_878_n N_A_2214_99#_c_1140_n 0.00995492f $X=11.925 $Y=1.67 $X2=0
+ $Y2=0
cc_676 N_SET_B_M1019_g N_A_2214_99#_c_1141_n 0.00103979f $X=11.835 $Y=0.835
+ $X2=0 $Y2=0
cc_677 N_SET_B_M1019_g N_A_1998_463#_M1031_g 0.0176345f $X=11.835 $Y=0.835 $X2=0
+ $Y2=0
cc_678 N_SET_B_c_874_n N_A_1998_463#_M1031_g 0.0213027f $X=11.87 $Y=1.835 $X2=0
+ $Y2=0
cc_679 N_SET_B_c_878_n N_A_1998_463#_c_1202_n 6.30604e-19 $X=11.925 $Y=1.67
+ $X2=0 $Y2=0
cc_680 N_SET_B_c_876_n N_A_1998_463#_c_1204_n 0.0715641f $X=10.955 $Y=1.585
+ $X2=0 $Y2=0
cc_681 N_SET_B_c_877_n N_A_1998_463#_c_1204_n 0.0152108f $X=11.04 $Y=1.675 $X2=0
+ $Y2=0
cc_682 N_SET_B_c_879_n N_A_1998_463#_c_1204_n 0.0458316f $X=10.87 $Y=0.382 $X2=0
+ $Y2=0
cc_683 N_SET_B_c_874_n N_A_1998_463#_c_1213_n 0.00124221f $X=11.87 $Y=1.835
+ $X2=0 $Y2=0
cc_684 N_SET_B_M1012_g N_A_1998_463#_c_1213_n 0.0158972f $X=11.87 $Y=2.385 $X2=0
+ $Y2=0
cc_685 N_SET_B_c_877_n N_A_1998_463#_c_1213_n 0.0130927f $X=11.04 $Y=1.675 $X2=0
+ $Y2=0
cc_686 N_SET_B_c_878_n N_A_1998_463#_c_1213_n 0.0666888f $X=11.925 $Y=1.67 $X2=0
+ $Y2=0
cc_687 N_SET_B_c_874_n N_A_1998_463#_c_1231_n 6.29432e-19 $X=11.87 $Y=1.835
+ $X2=0 $Y2=0
cc_688 N_SET_B_M1012_g N_A_1998_463#_c_1231_n 5.10999e-19 $X=11.87 $Y=2.385
+ $X2=0 $Y2=0
cc_689 N_SET_B_c_878_n N_A_1998_463#_c_1231_n 0.00682903f $X=11.925 $Y=1.67
+ $X2=0 $Y2=0
cc_690 N_SET_B_c_874_n N_A_1998_463#_c_1214_n 0.003482f $X=11.87 $Y=1.835 $X2=0
+ $Y2=0
cc_691 N_SET_B_M1012_g N_A_1998_463#_c_1214_n 0.00681672f $X=11.87 $Y=2.385
+ $X2=0 $Y2=0
cc_692 N_SET_B_c_874_n N_A_1998_463#_c_1215_n 0.00340711f $X=11.87 $Y=1.835
+ $X2=0 $Y2=0
cc_693 N_SET_B_M1012_g N_A_1998_463#_c_1215_n 0.00268139f $X=11.87 $Y=2.385
+ $X2=0 $Y2=0
cc_694 N_SET_B_c_878_n N_A_1998_463#_c_1215_n 0.0108374f $X=11.925 $Y=1.67 $X2=0
+ $Y2=0
cc_695 N_SET_B_M1004_g N_VPWR_c_1394_n 0.00123911f $X=8.225 $Y=2.105 $X2=0 $Y2=0
cc_696 N_SET_B_M1012_g N_VPWR_c_1395_n 0.00194124f $X=11.87 $Y=2.385 $X2=0 $Y2=0
cc_697 N_SET_B_M1012_g N_VPWR_c_1396_n 0.00269023f $X=11.87 $Y=2.385 $X2=0 $Y2=0
cc_698 N_SET_B_M1012_g N_VPWR_c_1412_n 0.00361794f $X=11.87 $Y=2.385 $X2=0 $Y2=0
cc_699 N_SET_B_M1012_g N_VPWR_c_1389_n 0.00440068f $X=11.87 $Y=2.385 $X2=0 $Y2=0
cc_700 N_SET_B_c_882_n N_VGND_M1027_d 0.0109389f $X=9.738 $Y=0.452 $X2=0 $Y2=0
cc_701 N_SET_B_c_881_n N_VGND_c_1794_n 0.0128871f $X=8.48 $Y=0.35 $X2=0 $Y2=0
cc_702 N_SET_B_c_882_n N_VGND_c_1794_n 0.0284786f $X=9.738 $Y=0.452 $X2=0 $Y2=0
cc_703 N_SET_B_M1027_g N_VGND_c_1846_n 0.00952524f $X=8.325 $Y=0.835 $X2=0 $Y2=0
cc_704 N_SET_B_c_881_n N_VGND_c_1846_n 0.00117733f $X=8.48 $Y=0.35 $X2=0 $Y2=0
cc_705 N_SET_B_c_882_n N_VGND_c_1846_n 0.0838459f $X=9.738 $Y=0.452 $X2=0 $Y2=0
cc_706 N_SET_B_M1019_g N_VGND_c_1795_n 0.0138423f $X=11.835 $Y=0.835 $X2=0 $Y2=0
cc_707 N_SET_B_M1019_g N_VGND_c_1801_n 0.00345209f $X=11.835 $Y=0.835 $X2=0
+ $Y2=0
cc_708 N_SET_B_c_879_n N_VGND_c_1801_n 0.0114622f $X=10.87 $Y=0.382 $X2=0 $Y2=0
cc_709 N_SET_B_c_881_n N_VGND_c_1801_n 0.00860664f $X=8.48 $Y=0.35 $X2=0 $Y2=0
cc_710 N_SET_B_c_882_n N_VGND_c_1801_n 0.160686f $X=9.738 $Y=0.452 $X2=0 $Y2=0
cc_711 N_SET_B_M1019_g N_VGND_c_1814_n 0.00394323f $X=11.835 $Y=0.835 $X2=0
+ $Y2=0
cc_712 N_SET_B_c_879_n N_VGND_c_1814_n 0.00657784f $X=10.87 $Y=0.382 $X2=0 $Y2=0
cc_713 N_SET_B_c_881_n N_VGND_c_1814_n 0.0121286f $X=8.48 $Y=0.35 $X2=0 $Y2=0
cc_714 N_SET_B_c_882_n N_VGND_c_1814_n 0.0953402f $X=9.738 $Y=0.452 $X2=0 $Y2=0
cc_715 SET_B A_1933_125# 0.00335841f $X=9.755 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_716 N_SET_B_c_882_n A_1933_125# 6.29702e-19 $X=9.738 $Y=0.452 $X2=-0.19
+ $Y2=-0.245
cc_717 N_SET_B_c_876_n A_2159_125# 0.00638609f $X=10.955 $Y=1.585 $X2=-0.19
+ $Y2=-0.245
cc_718 N_A_794_47#_M1002_g N_A_2214_99#_c_1137_n 0.0295842f $X=10.72 $Y=0.835
+ $X2=0 $Y2=0
cc_719 N_A_794_47#_M1002_g N_A_2214_99#_M1025_g 0.00190835f $X=10.72 $Y=0.835
+ $X2=0 $Y2=0
cc_720 N_A_794_47#_c_973_n N_A_2214_99#_M1025_g 0.0312735f $X=10.72 $Y=1.755
+ $X2=0 $Y2=0
cc_721 N_A_794_47#_M1002_g N_A_2214_99#_c_1140_n 0.00385253f $X=10.72 $Y=0.835
+ $X2=0 $Y2=0
cc_722 N_A_794_47#_c_983_n N_A_1998_463#_c_1211_n 0.00736821f $X=10.46 $Y=1.785
+ $X2=0 $Y2=0
cc_723 N_A_794_47#_c_984_n N_A_1998_463#_c_1211_n 5.43792e-19 $X=10.95 $Y=3.075
+ $X2=0 $Y2=0
cc_724 N_A_794_47#_c_983_n N_A_1998_463#_c_1204_n 0.00423205f $X=10.46 $Y=1.785
+ $X2=0 $Y2=0
cc_725 N_A_794_47#_M1002_g N_A_1998_463#_c_1204_n 0.0246745f $X=10.72 $Y=0.835
+ $X2=0 $Y2=0
cc_726 N_A_794_47#_c_984_n N_A_1998_463#_c_1204_n 0.00105339f $X=10.95 $Y=3.075
+ $X2=0 $Y2=0
cc_727 N_A_794_47#_c_973_n N_A_1998_463#_c_1204_n 0.020735f $X=10.72 $Y=1.755
+ $X2=0 $Y2=0
cc_728 N_A_794_47#_c_984_n N_A_1998_463#_c_1213_n 0.0156917f $X=10.95 $Y=3.075
+ $X2=0 $Y2=0
cc_729 N_A_794_47#_c_973_n N_A_1998_463#_c_1213_n 0.00681298f $X=10.72 $Y=1.755
+ $X2=0 $Y2=0
cc_730 N_A_794_47#_M1000_g N_VPWR_c_1392_n 0.00744981f $X=4.88 $Y=2.735 $X2=0
+ $Y2=0
cc_731 N_A_794_47#_c_978_n N_VPWR_c_1392_n 0.00117266f $X=5.37 $Y=3.075 $X2=0
+ $Y2=0
cc_732 N_A_794_47#_c_980_n N_VPWR_c_1392_n 7.40493e-19 $X=5.445 $Y=3.15 $X2=0
+ $Y2=0
cc_733 N_A_794_47#_M1001_g N_VPWR_c_1393_n 0.00361451f $X=6.56 $Y=2.285 $X2=0
+ $Y2=0
cc_734 N_A_794_47#_c_982_n N_VPWR_c_1393_n 0.026053f $X=10.875 $Y=3.15 $X2=0
+ $Y2=0
cc_735 N_A_794_47#_c_982_n N_VPWR_c_1394_n 0.0202126f $X=10.875 $Y=3.15 $X2=0
+ $Y2=0
cc_736 N_A_794_47#_c_984_n N_VPWR_c_1395_n 0.00617519f $X=10.95 $Y=3.075 $X2=0
+ $Y2=0
cc_737 N_A_794_47#_M1000_g N_VPWR_c_1402_n 0.00452967f $X=4.88 $Y=2.735 $X2=0
+ $Y2=0
cc_738 N_A_794_47#_c_980_n N_VPWR_c_1402_n 0.0396622f $X=5.445 $Y=3.15 $X2=0
+ $Y2=0
cc_739 N_A_794_47#_c_982_n N_VPWR_c_1404_n 0.0330265f $X=10.875 $Y=3.15 $X2=0
+ $Y2=0
cc_740 N_A_794_47#_c_982_n N_VPWR_c_1406_n 0.0560513f $X=10.875 $Y=3.15 $X2=0
+ $Y2=0
cc_741 N_A_794_47#_M1000_g N_VPWR_c_1389_n 0.00443906f $X=4.88 $Y=2.735 $X2=0
+ $Y2=0
cc_742 N_A_794_47#_c_979_n N_VPWR_c_1389_n 0.0245183f $X=6.485 $Y=3.15 $X2=0
+ $Y2=0
cc_743 N_A_794_47#_c_980_n N_VPWR_c_1389_n 0.00510574f $X=5.445 $Y=3.15 $X2=0
+ $Y2=0
cc_744 N_A_794_47#_c_982_n N_VPWR_c_1389_n 0.117579f $X=10.875 $Y=3.15 $X2=0
+ $Y2=0
cc_745 N_A_794_47#_c_985_n N_VPWR_c_1389_n 0.00372139f $X=6.56 $Y=3.15 $X2=0
+ $Y2=0
cc_746 N_A_794_47#_M1020_s N_A_244_121#_c_1568_n 0.00560524f $X=4.015 $Y=2.085
+ $X2=0 $Y2=0
cc_747 N_A_794_47#_c_990_n N_A_244_121#_c_1568_n 0.006755f $X=4.305 $Y=2.16
+ $X2=0 $Y2=0
cc_748 N_A_794_47#_c_988_n N_A_244_121#_c_1623_n 0.0129612f $X=4.855 $Y=2.09
+ $X2=0 $Y2=0
cc_749 N_A_794_47#_M1000_g N_A_244_121#_c_1570_n 0.00935405f $X=4.88 $Y=2.735
+ $X2=0 $Y2=0
cc_750 N_A_794_47#_c_978_n N_A_244_121#_c_1570_n 0.00916814f $X=5.37 $Y=3.075
+ $X2=0 $Y2=0
cc_751 N_A_794_47#_c_988_n N_A_244_121#_c_1570_n 0.00167466f $X=4.855 $Y=2.09
+ $X2=0 $Y2=0
cc_752 N_A_794_47#_c_1096_p N_A_244_121#_c_1570_n 0.021919f $X=4.995 $Y=1.995
+ $X2=0 $Y2=0
cc_753 N_A_794_47#_c_991_n N_A_244_121#_c_1570_n 0.00570835f $X=4.97 $Y=2.09
+ $X2=0 $Y2=0
cc_754 N_A_794_47#_c_968_n N_A_244_121#_c_1562_n 0.00349082f $X=4.74 $Y=0.765
+ $X2=0 $Y2=0
cc_755 N_A_794_47#_c_969_n N_A_244_121#_c_1562_n 0.0177845f $X=6.035 $Y=1.06
+ $X2=0 $Y2=0
cc_756 N_A_794_47#_M1034_g N_A_244_121#_c_1562_n 0.00201203f $X=6.11 $Y=0.485
+ $X2=0 $Y2=0
cc_757 N_A_794_47#_c_972_n N_A_244_121#_c_1562_n 0.0156491f $X=5.125 $Y=1.135
+ $X2=0 $Y2=0
cc_758 N_A_794_47#_c_1096_p N_A_244_121#_c_1562_n 0.0112814f $X=4.995 $Y=1.995
+ $X2=0 $Y2=0
cc_759 N_A_794_47#_c_1009_n N_A_244_121#_c_1562_n 0.0414264f $X=4.97 $Y=1.41
+ $X2=0 $Y2=0
cc_760 N_A_794_47#_c_975_n N_A_244_121#_c_1562_n 0.0319854f $X=4.97 $Y=1.41
+ $X2=0 $Y2=0
cc_761 N_A_794_47#_c_991_n N_A_244_121#_c_1562_n 0.00956563f $X=4.97 $Y=2.09
+ $X2=0 $Y2=0
cc_762 N_A_794_47#_M1020_s N_A_244_121#_c_1611_n 0.0111803f $X=4.015 $Y=2.085
+ $X2=0 $Y2=0
cc_763 N_A_794_47#_c_988_n N_A_244_121#_c_1611_n 6.84046e-19 $X=4.855 $Y=2.09
+ $X2=0 $Y2=0
cc_764 N_A_794_47#_c_990_n N_A_244_121#_c_1611_n 0.0128181f $X=4.305 $Y=2.16
+ $X2=0 $Y2=0
cc_765 N_A_794_47#_M1000_g N_A_244_121#_c_1573_n 0.00632142f $X=4.88 $Y=2.735
+ $X2=0 $Y2=0
cc_766 N_A_794_47#_c_978_n N_A_244_121#_c_1573_n 7.51633e-19 $X=5.37 $Y=3.075
+ $X2=0 $Y2=0
cc_767 N_A_794_47#_c_988_n N_A_244_121#_c_1573_n 0.0132352f $X=4.855 $Y=2.09
+ $X2=0 $Y2=0
cc_768 N_A_794_47#_M1000_g N_A_244_121#_c_1574_n 5.94155e-19 $X=4.88 $Y=2.735
+ $X2=0 $Y2=0
cc_769 N_A_794_47#_c_978_n N_A_244_121#_c_1574_n 0.00896705f $X=5.37 $Y=3.075
+ $X2=0 $Y2=0
cc_770 N_A_794_47#_c_991_n N_A_244_121#_c_1574_n 0.00475f $X=4.97 $Y=2.09 $X2=0
+ $Y2=0
cc_771 N_A_794_47#_c_982_n N_A_1781_379#_c_1697_n 0.00488407f $X=10.875 $Y=3.15
+ $X2=0 $Y2=0
cc_772 N_A_794_47#_c_983_n N_A_1781_379#_c_1697_n 0.00964289f $X=10.46 $Y=1.785
+ $X2=0 $Y2=0
cc_773 N_A_794_47#_c_982_n N_A_1781_379#_c_1699_n 0.00592942f $X=10.875 $Y=3.15
+ $X2=0 $Y2=0
cc_774 N_A_794_47#_c_983_n N_A_1781_379#_c_1700_n 0.00493282f $X=10.46 $Y=1.785
+ $X2=0 $Y2=0
cc_775 N_A_794_47#_c_984_n N_A_1781_379#_c_1700_n 0.00321516f $X=10.95 $Y=3.075
+ $X2=0 $Y2=0
cc_776 N_A_794_47#_c_973_n N_A_1781_379#_c_1700_n 7.50836e-19 $X=10.72 $Y=1.755
+ $X2=0 $Y2=0
cc_777 N_A_794_47#_c_982_n N_A_1888_463#_c_1733_n 0.0181467f $X=10.875 $Y=3.15
+ $X2=0 $Y2=0
cc_778 N_A_794_47#_c_983_n N_A_1888_463#_c_1733_n 0.00650876f $X=10.46 $Y=1.785
+ $X2=0 $Y2=0
cc_779 N_A_794_47#_c_984_n N_A_1888_463#_c_1733_n 0.0178301f $X=10.95 $Y=3.075
+ $X2=0 $Y2=0
cc_780 N_A_794_47#_c_984_n N_A_1888_463#_c_1734_n 0.00922496f $X=10.95 $Y=3.075
+ $X2=0 $Y2=0
cc_781 N_A_794_47#_c_982_n N_A_1888_463#_c_1735_n 0.00742651f $X=10.875 $Y=3.15
+ $X2=0 $Y2=0
cc_782 N_A_794_47#_c_968_n N_VGND_c_1792_n 0.00315529f $X=4.74 $Y=0.765 $X2=0
+ $Y2=0
cc_783 N_A_794_47#_M1002_g N_VGND_c_1801_n 5.42344e-19 $X=10.72 $Y=0.835 $X2=0
+ $Y2=0
cc_784 N_A_794_47#_c_976_n N_VGND_c_1807_n 0.0142913f $X=4.095 $Y=0.445 $X2=0
+ $Y2=0
cc_785 N_A_794_47#_c_968_n N_VGND_c_1808_n 0.00585385f $X=4.74 $Y=0.765 $X2=0
+ $Y2=0
cc_786 N_A_794_47#_M1034_g N_VGND_c_1808_n 0.00495687f $X=6.11 $Y=0.485 $X2=0
+ $Y2=0
cc_787 N_A_794_47#_c_972_n N_VGND_c_1808_n 2.79886e-19 $X=5.125 $Y=1.135 $X2=0
+ $Y2=0
cc_788 N_A_794_47#_M1010_s N_VGND_c_1814_n 0.00237743f $X=3.97 $Y=0.235 $X2=0
+ $Y2=0
cc_789 N_A_794_47#_c_968_n N_VGND_c_1814_n 0.0115819f $X=4.74 $Y=0.765 $X2=0
+ $Y2=0
cc_790 N_A_794_47#_M1034_g N_VGND_c_1814_n 0.0102613f $X=6.11 $Y=0.485 $X2=0
+ $Y2=0
cc_791 N_A_794_47#_c_972_n N_VGND_c_1814_n 2.93956e-19 $X=5.125 $Y=1.135 $X2=0
+ $Y2=0
cc_792 N_A_794_47#_c_976_n N_VGND_c_1814_n 0.0100306f $X=4.095 $Y=0.445 $X2=0
+ $Y2=0
cc_793 N_A_2214_99#_c_1139_n N_A_1998_463#_M1031_g 0.0127786f $X=12.425 $Y=1.325
+ $X2=0 $Y2=0
cc_794 N_A_2214_99#_c_1141_n N_A_1998_463#_M1031_g 0.0133149f $X=12.59 $Y=0.83
+ $X2=0 $Y2=0
cc_795 N_A_2214_99#_c_1142_n N_A_1998_463#_M1031_g 0.00530037f $X=13.065
+ $Y=1.415 $X2=0 $Y2=0
cc_796 N_A_2214_99#_c_1143_n N_A_1998_463#_M1031_g 0.00416818f $X=13.035
+ $Y=2.625 $X2=0 $Y2=0
cc_797 N_A_2214_99#_c_1142_n N_A_1998_463#_c_1200_n 0.00137108f $X=13.065
+ $Y=1.415 $X2=0 $Y2=0
cc_798 N_A_2214_99#_c_1143_n N_A_1998_463#_c_1200_n 0.0182569f $X=13.035
+ $Y=2.625 $X2=0 $Y2=0
cc_799 N_A_2214_99#_c_1142_n N_A_1998_463#_M1006_g 5.71476e-19 $X=13.065
+ $Y=1.415 $X2=0 $Y2=0
cc_800 N_A_2214_99#_c_1143_n N_A_1998_463#_M1006_g 6.09292e-19 $X=13.035
+ $Y=2.625 $X2=0 $Y2=0
cc_801 N_A_2214_99#_c_1143_n N_A_1998_463#_c_1207_n 0.00310459f $X=13.035
+ $Y=2.625 $X2=0 $Y2=0
cc_802 N_A_2214_99#_c_1142_n N_A_1998_463#_c_1202_n 0.0130114f $X=13.065
+ $Y=1.415 $X2=0 $Y2=0
cc_803 N_A_2214_99#_M1025_g N_A_1998_463#_c_1213_n 0.0150639f $X=11.44 $Y=2.385
+ $X2=0 $Y2=0
cc_804 N_A_2214_99#_c_1142_n N_A_1998_463#_c_1231_n 0.0206794f $X=13.065
+ $Y=1.415 $X2=0 $Y2=0
cc_805 N_A_2214_99#_c_1143_n N_A_1998_463#_c_1231_n 0.0261591f $X=13.035
+ $Y=2.625 $X2=0 $Y2=0
cc_806 N_A_2214_99#_c_1143_n N_A_1998_463#_c_1214_n 0.0215604f $X=13.035
+ $Y=2.625 $X2=0 $Y2=0
cc_807 N_A_2214_99#_c_1139_n N_A_1998_463#_c_1215_n 0.0147473f $X=12.425
+ $Y=1.325 $X2=0 $Y2=0
cc_808 N_A_2214_99#_c_1143_n N_A_1998_463#_c_1215_n 0.0264069f $X=13.035
+ $Y=2.625 $X2=0 $Y2=0
cc_809 N_A_2214_99#_c_1141_n N_A_2686_131#_c_1304_n 0.0175664f $X=12.59 $Y=0.83
+ $X2=0 $Y2=0
cc_810 N_A_2214_99#_c_1142_n N_A_2686_131#_c_1304_n 0.0063468f $X=13.065
+ $Y=1.415 $X2=0 $Y2=0
cc_811 N_A_2214_99#_c_1143_n N_A_2686_131#_c_1310_n 0.0624823f $X=13.035
+ $Y=2.625 $X2=0 $Y2=0
cc_812 N_A_2214_99#_c_1142_n N_A_2686_131#_c_1306_n 0.00856983f $X=13.065
+ $Y=1.415 $X2=0 $Y2=0
cc_813 N_A_2214_99#_c_1143_n N_A_2686_131#_c_1306_n 0.0179332f $X=13.035
+ $Y=2.625 $X2=0 $Y2=0
cc_814 N_A_2214_99#_M1025_g N_VPWR_c_1395_n 0.00102367f $X=11.44 $Y=2.385 $X2=0
+ $Y2=0
cc_815 N_A_2214_99#_c_1143_n N_VPWR_c_1397_n 0.00979029f $X=13.035 $Y=2.625
+ $X2=0 $Y2=0
cc_816 N_A_2214_99#_M1025_g N_VPWR_c_1406_n 0.00361794f $X=11.44 $Y=2.385 $X2=0
+ $Y2=0
cc_817 N_A_2214_99#_c_1143_n N_VPWR_c_1408_n 0.00623679f $X=13.035 $Y=2.625
+ $X2=0 $Y2=0
cc_818 N_A_2214_99#_M1025_g N_VPWR_c_1389_n 0.00440068f $X=11.44 $Y=2.385 $X2=0
+ $Y2=0
cc_819 N_A_2214_99#_c_1143_n N_VPWR_c_1389_n 0.00871514f $X=13.035 $Y=2.625
+ $X2=0 $Y2=0
cc_820 N_A_2214_99#_M1025_g N_A_1888_463#_c_1734_n 0.00117326f $X=11.44 $Y=2.385
+ $X2=0 $Y2=0
cc_821 N_A_2214_99#_c_1137_n N_VGND_c_1795_n 0.00213306f $X=11.145 $Y=1.155
+ $X2=0 $Y2=0
cc_822 N_A_2214_99#_c_1139_n N_VGND_c_1795_n 0.0190476f $X=12.425 $Y=1.325 $X2=0
+ $Y2=0
cc_823 N_A_2214_99#_c_1141_n N_VGND_c_1795_n 0.0217738f $X=12.59 $Y=0.83 $X2=0
+ $Y2=0
cc_824 N_A_2214_99#_c_1137_n N_VGND_c_1801_n 0.00415323f $X=11.145 $Y=1.155
+ $X2=0 $Y2=0
cc_825 N_A_2214_99#_c_1141_n N_VGND_c_1803_n 0.00535315f $X=12.59 $Y=0.83 $X2=0
+ $Y2=0
cc_826 N_A_2214_99#_c_1137_n N_VGND_c_1814_n 0.00469432f $X=11.145 $Y=1.155
+ $X2=0 $Y2=0
cc_827 N_A_2214_99#_c_1141_n N_VGND_c_1814_n 0.00961232f $X=12.59 $Y=0.83 $X2=0
+ $Y2=0
cc_828 N_A_1998_463#_M1006_g N_A_2686_131#_M1021_g 0.0172392f $X=13.77 $Y=0.865
+ $X2=0 $Y2=0
cc_829 N_A_1998_463#_c_1203_n N_A_2686_131#_M1028_g 0.0191288f $X=13.77 $Y=1.65
+ $X2=0 $Y2=0
cc_830 N_A_1998_463#_M1006_g N_A_2686_131#_c_1304_n 0.0101034f $X=13.77 $Y=0.865
+ $X2=0 $Y2=0
cc_831 N_A_1998_463#_c_1200_n N_A_2686_131#_c_1310_n 0.00991233f $X=13.695
+ $Y=1.65 $X2=0 $Y2=0
cc_832 N_A_1998_463#_c_1207_n N_A_2686_131#_c_1310_n 0.00480341f $X=13.77
+ $Y=1.725 $X2=0 $Y2=0
cc_833 N_A_1998_463#_c_1200_n N_A_2686_131#_c_1305_n 4.34011e-19 $X=13.695
+ $Y=1.65 $X2=0 $Y2=0
cc_834 N_A_1998_463#_M1006_g N_A_2686_131#_c_1305_n 0.0184348f $X=13.77 $Y=0.865
+ $X2=0 $Y2=0
cc_835 N_A_1998_463#_c_1203_n N_A_2686_131#_c_1305_n 0.00885751f $X=13.77
+ $Y=1.65 $X2=0 $Y2=0
cc_836 N_A_1998_463#_c_1200_n N_A_2686_131#_c_1306_n 0.00819928f $X=13.695
+ $Y=1.65 $X2=0 $Y2=0
cc_837 N_A_1998_463#_M1006_g N_A_2686_131#_c_1307_n 0.0181395f $X=13.77 $Y=0.865
+ $X2=0 $Y2=0
cc_838 N_A_1998_463#_c_1213_n N_VPWR_c_1395_n 0.0170158f $X=11.955 $Y=2.02 $X2=0
+ $Y2=0
cc_839 N_A_1998_463#_M1003_g N_VPWR_c_1396_n 0.0141614f $X=12.82 $Y=2.625 $X2=0
+ $Y2=0
cc_840 N_A_1998_463#_c_1209_n N_VPWR_c_1396_n 0.00168278f $X=12.697 $Y=2.255
+ $X2=0 $Y2=0
cc_841 N_A_1998_463#_c_1215_n N_VPWR_c_1396_n 0.0286682f $X=12.085 $Y=2.385
+ $X2=0 $Y2=0
cc_842 N_A_1998_463#_c_1207_n N_VPWR_c_1397_n 0.00388706f $X=13.77 $Y=1.725
+ $X2=0 $Y2=0
cc_843 N_A_1998_463#_M1003_g N_VPWR_c_1408_n 0.00440637f $X=12.82 $Y=2.625 $X2=0
+ $Y2=0
cc_844 N_A_1998_463#_c_1207_n N_VPWR_c_1408_n 0.00312414f $X=13.77 $Y=1.725
+ $X2=0 $Y2=0
cc_845 N_A_1998_463#_M1003_g N_VPWR_c_1389_n 0.00459568f $X=12.82 $Y=2.625 $X2=0
+ $Y2=0
cc_846 N_A_1998_463#_c_1207_n N_VPWR_c_1389_n 0.00410284f $X=13.77 $Y=1.725
+ $X2=0 $Y2=0
cc_847 N_A_1998_463#_c_1215_n N_VPWR_c_1389_n 0.0121434f $X=12.085 $Y=2.385
+ $X2=0 $Y2=0
cc_848 N_A_1998_463#_c_1211_n N_A_1781_379#_M1030_d 0.00145605f $X=10.397
+ $Y=1.915 $X2=0 $Y2=0
cc_849 N_A_1998_463#_c_1204_n N_A_1781_379#_M1030_d 2.57675e-19 $X=10.505 $Y=0.8
+ $X2=0 $Y2=0
cc_850 N_A_1998_463#_c_1213_n N_A_1781_379#_M1030_d 0.00201436f $X=11.955
+ $Y=2.02 $X2=0 $Y2=0
cc_851 N_A_1998_463#_M1032_d N_A_1781_379#_c_1697_n 0.00653602f $X=9.99 $Y=2.315
+ $X2=0 $Y2=0
cc_852 N_A_1998_463#_c_1211_n N_A_1781_379#_c_1697_n 0.0295967f $X=10.397
+ $Y=1.915 $X2=0 $Y2=0
cc_853 N_A_1998_463#_c_1211_n N_A_1781_379#_c_1700_n 0.0111086f $X=10.397
+ $Y=1.915 $X2=0 $Y2=0
cc_854 N_A_1998_463#_c_1213_n N_A_1781_379#_c_1700_n 0.0107747f $X=11.955
+ $Y=2.02 $X2=0 $Y2=0
cc_855 N_A_1998_463#_c_1213_n N_A_1888_463#_c_1734_n 0.0224458f $X=11.955
+ $Y=2.02 $X2=0 $Y2=0
cc_856 N_A_1998_463#_c_1204_n N_VGND_c_1846_n 0.00672688f $X=10.505 $Y=0.8 $X2=0
+ $Y2=0
cc_857 N_A_1998_463#_M1031_g N_VGND_c_1795_n 0.00761689f $X=12.375 $Y=0.835
+ $X2=0 $Y2=0
cc_858 N_A_1998_463#_M1006_g N_VGND_c_1796_n 0.0138477f $X=13.77 $Y=0.865 $X2=0
+ $Y2=0
cc_859 N_A_1998_463#_M1031_g N_VGND_c_1803_n 0.00400506f $X=12.375 $Y=0.835
+ $X2=0 $Y2=0
cc_860 N_A_1998_463#_M1006_g N_VGND_c_1803_n 0.00385681f $X=13.77 $Y=0.865 $X2=0
+ $Y2=0
cc_861 N_A_1998_463#_M1031_g N_VGND_c_1814_n 0.00469432f $X=12.375 $Y=0.835
+ $X2=0 $Y2=0
cc_862 N_A_1998_463#_M1006_g N_VGND_c_1814_n 0.0044892f $X=13.77 $Y=0.865 $X2=0
+ $Y2=0
cc_863 N_A_2686_131#_M1028_g N_VPWR_c_1397_n 0.0246053f $X=14.28 $Y=2.465 $X2=0
+ $Y2=0
cc_864 N_A_2686_131#_M1039_g N_VPWR_c_1397_n 7.93019e-19 $X=14.71 $Y=2.465 $X2=0
+ $Y2=0
cc_865 N_A_2686_131#_c_1310_n N_VPWR_c_1397_n 0.00149665f $X=13.555 $Y=1.98
+ $X2=0 $Y2=0
cc_866 N_A_2686_131#_c_1305_n N_VPWR_c_1397_n 0.0302138f $X=14.25 $Y=1.48 $X2=0
+ $Y2=0
cc_867 N_A_2686_131#_c_1307_n N_VPWR_c_1397_n 0.0027817f $X=14.25 $Y=1.39 $X2=0
+ $Y2=0
cc_868 N_A_2686_131#_M1028_g N_VPWR_c_1399_n 7.11463e-19 $X=14.28 $Y=2.465 $X2=0
+ $Y2=0
cc_869 N_A_2686_131#_M1039_g N_VPWR_c_1399_n 0.0145974f $X=14.71 $Y=2.465 $X2=0
+ $Y2=0
cc_870 N_A_2686_131#_M1028_g N_VPWR_c_1413_n 0.00525069f $X=14.28 $Y=2.465 $X2=0
+ $Y2=0
cc_871 N_A_2686_131#_M1039_g N_VPWR_c_1413_n 0.00486043f $X=14.71 $Y=2.465 $X2=0
+ $Y2=0
cc_872 N_A_2686_131#_M1028_g N_VPWR_c_1389_n 0.00886509f $X=14.28 $Y=2.465 $X2=0
+ $Y2=0
cc_873 N_A_2686_131#_M1039_g N_VPWR_c_1389_n 0.00824727f $X=14.71 $Y=2.465 $X2=0
+ $Y2=0
cc_874 N_A_2686_131#_c_1310_n N_VPWR_c_1389_n 0.0115026f $X=13.555 $Y=1.98 $X2=0
+ $Y2=0
cc_875 N_A_2686_131#_M1021_g N_Q_c_1759_n 0.00200698f $X=14.28 $Y=0.655 $X2=0
+ $Y2=0
cc_876 N_A_2686_131#_c_1300_n N_Q_c_1759_n 0.00406666f $X=14.635 $Y=1.39 $X2=0
+ $Y2=0
cc_877 N_A_2686_131#_M1036_g N_Q_c_1759_n 0.0135958f $X=14.71 $Y=0.655 $X2=0
+ $Y2=0
cc_878 N_A_2686_131#_M1028_g N_Q_c_1761_n 6.94505e-19 $X=14.28 $Y=2.465 $X2=0
+ $Y2=0
cc_879 N_A_2686_131#_c_1300_n N_Q_c_1761_n 0.00492089f $X=14.635 $Y=1.39 $X2=0
+ $Y2=0
cc_880 N_A_2686_131#_M1039_g N_Q_c_1761_n 0.0131192f $X=14.71 $Y=2.465 $X2=0
+ $Y2=0
cc_881 N_A_2686_131#_c_1307_n N_Q_c_1761_n 0.00114878f $X=14.25 $Y=1.39 $X2=0
+ $Y2=0
cc_882 N_A_2686_131#_M1021_g Q 0.00344624f $X=14.28 $Y=0.655 $X2=0 $Y2=0
cc_883 N_A_2686_131#_M1028_g Q 0.00344624f $X=14.28 $Y=2.465 $X2=0 $Y2=0
cc_884 N_A_2686_131#_c_1300_n Q 0.00544118f $X=14.635 $Y=1.39 $X2=0 $Y2=0
cc_885 N_A_2686_131#_M1036_g Q 0.00779839f $X=14.71 $Y=0.655 $X2=0 $Y2=0
cc_886 N_A_2686_131#_M1039_g Q 0.0150943f $X=14.71 $Y=2.465 $X2=0 $Y2=0
cc_887 N_A_2686_131#_c_1303_n Q 0.0054821f $X=14.71 $Y=1.39 $X2=0 $Y2=0
cc_888 N_A_2686_131#_c_1305_n Q 0.0233909f $X=14.25 $Y=1.48 $X2=0 $Y2=0
cc_889 N_A_2686_131#_c_1307_n Q 0.00137117f $X=14.25 $Y=1.39 $X2=0 $Y2=0
cc_890 N_A_2686_131#_M1021_g N_VGND_c_1796_n 0.00601974f $X=14.28 $Y=0.655 $X2=0
+ $Y2=0
cc_891 N_A_2686_131#_c_1304_n N_VGND_c_1796_n 0.0155924f $X=13.555 $Y=0.865
+ $X2=0 $Y2=0
cc_892 N_A_2686_131#_c_1305_n N_VGND_c_1796_n 0.0238096f $X=14.25 $Y=1.48 $X2=0
+ $Y2=0
cc_893 N_A_2686_131#_c_1307_n N_VGND_c_1796_n 0.00190611f $X=14.25 $Y=1.39 $X2=0
+ $Y2=0
cc_894 N_A_2686_131#_M1021_g N_VGND_c_1798_n 6.26874e-19 $X=14.28 $Y=0.655 $X2=0
+ $Y2=0
cc_895 N_A_2686_131#_M1036_g N_VGND_c_1798_n 0.0109716f $X=14.71 $Y=0.655 $X2=0
+ $Y2=0
cc_896 N_A_2686_131#_c_1304_n N_VGND_c_1803_n 0.00445281f $X=13.555 $Y=0.865
+ $X2=0 $Y2=0
cc_897 N_A_2686_131#_M1021_g N_VGND_c_1809_n 0.00585385f $X=14.28 $Y=0.655 $X2=0
+ $Y2=0
cc_898 N_A_2686_131#_M1036_g N_VGND_c_1809_n 0.00486043f $X=14.71 $Y=0.655 $X2=0
+ $Y2=0
cc_899 N_A_2686_131#_M1021_g N_VGND_c_1814_n 0.0118904f $X=14.28 $Y=0.655 $X2=0
+ $Y2=0
cc_900 N_A_2686_131#_M1036_g N_VGND_c_1814_n 0.00824727f $X=14.71 $Y=0.655 $X2=0
+ $Y2=0
cc_901 N_A_2686_131#_c_1304_n N_VGND_c_1814_n 0.00804028f $X=13.555 $Y=0.865
+ $X2=0 $Y2=0
cc_902 N_A_39_481#_c_1367_n N_VPWR_M1037_d 0.00173127f $X=2.08 $Y=2.55 $X2=-0.19
+ $Y2=1.655
cc_903 N_A_39_481#_c_1366_n N_VPWR_c_1390_n 0.0101431f $X=0.32 $Y=2.9 $X2=0
+ $Y2=0
cc_904 N_A_39_481#_c_1367_n N_VPWR_c_1390_n 0.0166605f $X=2.08 $Y=2.55 $X2=0
+ $Y2=0
cc_905 N_A_39_481#_c_1367_n N_VPWR_c_1400_n 0.00688458f $X=2.08 $Y=2.55 $X2=0
+ $Y2=0
cc_906 N_A_39_481#_c_1366_n N_VPWR_c_1410_n 0.017376f $X=0.32 $Y=2.9 $X2=0 $Y2=0
cc_907 N_A_39_481#_c_1367_n N_VPWR_c_1410_n 0.00223975f $X=2.08 $Y=2.55 $X2=0
+ $Y2=0
cc_908 N_A_39_481#_c_1366_n N_VPWR_c_1389_n 0.00997879f $X=0.32 $Y=2.9 $X2=0
+ $Y2=0
cc_909 N_A_39_481#_c_1367_n N_VPWR_c_1389_n 0.0200611f $X=2.08 $Y=2.55 $X2=0
+ $Y2=0
cc_910 N_A_39_481#_c_1367_n A_208_481# 0.00179114f $X=2.08 $Y=2.55 $X2=-0.19
+ $Y2=1.655
cc_911 N_A_39_481#_c_1367_n N_A_244_121#_M1018_d 0.00328212f $X=2.08 $Y=2.55
+ $X2=0 $Y2=0
cc_912 N_A_39_481#_M1033_d N_A_244_121#_c_1563_n 0.00330823f $X=1.94 $Y=2.405
+ $X2=0 $Y2=0
cc_913 N_A_39_481#_c_1367_n N_A_244_121#_c_1563_n 0.0490665f $X=2.08 $Y=2.55
+ $X2=0 $Y2=0
cc_914 N_A_39_481#_c_1367_n N_A_244_121#_c_1565_n 0.0201139f $X=2.08 $Y=2.55
+ $X2=0 $Y2=0
cc_915 N_VPWR_c_1390_n N_A_244_121#_c_1563_n 0.00451626f $X=0.75 $Y=2.92 $X2=0
+ $Y2=0
cc_916 N_VPWR_c_1391_n N_A_244_121#_c_1563_n 0.0226147f $X=2.93 $Y=2.465 $X2=0
+ $Y2=0
cc_917 N_VPWR_c_1400_n N_A_244_121#_c_1563_n 0.0776493f $X=2.765 $Y=3.33 $X2=0
+ $Y2=0
cc_918 N_VPWR_c_1389_n N_A_244_121#_c_1563_n 0.0436693f $X=15.12 $Y=3.33 $X2=0
+ $Y2=0
cc_919 N_VPWR_c_1391_n N_A_244_121#_c_1565_n 0.0400342f $X=2.93 $Y=2.465 $X2=0
+ $Y2=0
cc_920 N_VPWR_c_1391_n N_A_244_121#_c_1566_n 0.0209251f $X=2.93 $Y=2.465 $X2=0
+ $Y2=0
cc_921 N_VPWR_M1014_s N_A_244_121#_c_1567_n 0.00521084f $X=2.795 $Y=2.31 $X2=0
+ $Y2=0
cc_922 N_VPWR_c_1391_n N_A_244_121#_c_1567_n 0.0375009f $X=2.93 $Y=2.465 $X2=0
+ $Y2=0
cc_923 N_VPWR_c_1411_n N_A_244_121#_c_1568_n 0.0300459f $X=4.5 $Y=3.33 $X2=0
+ $Y2=0
cc_924 N_VPWR_c_1389_n N_A_244_121#_c_1568_n 0.0274738f $X=15.12 $Y=3.33 $X2=0
+ $Y2=0
cc_925 N_VPWR_M1014_s N_A_244_121#_c_1569_n 0.00166402f $X=2.795 $Y=2.31 $X2=0
+ $Y2=0
cc_926 N_VPWR_c_1391_n N_A_244_121#_c_1569_n 0.0143026f $X=2.93 $Y=2.465 $X2=0
+ $Y2=0
cc_927 N_VPWR_c_1411_n N_A_244_121#_c_1569_n 0.0071719f $X=4.5 $Y=3.33 $X2=0
+ $Y2=0
cc_928 N_VPWR_c_1389_n N_A_244_121#_c_1569_n 0.00620582f $X=15.12 $Y=3.33 $X2=0
+ $Y2=0
cc_929 N_VPWR_M1020_d N_A_244_121#_c_1623_n 0.00230146f $X=4.525 $Y=2.415 $X2=0
+ $Y2=0
cc_930 N_VPWR_c_1392_n N_A_244_121#_c_1623_n 0.00768852f $X=4.665 $Y=2.93 $X2=0
+ $Y2=0
cc_931 N_VPWR_c_1411_n N_A_244_121#_c_1623_n 0.00239434f $X=4.5 $Y=3.33 $X2=0
+ $Y2=0
cc_932 N_VPWR_c_1389_n N_A_244_121#_c_1623_n 0.0050981f $X=15.12 $Y=3.33 $X2=0
+ $Y2=0
cc_933 N_VPWR_c_1389_n N_A_244_121#_c_1570_n 0.00572383f $X=15.12 $Y=3.33 $X2=0
+ $Y2=0
cc_934 N_VPWR_c_1411_n N_A_244_121#_c_1611_n 0.00681871f $X=4.5 $Y=3.33 $X2=0
+ $Y2=0
cc_935 N_VPWR_c_1389_n N_A_244_121#_c_1611_n 0.0060866f $X=15.12 $Y=3.33 $X2=0
+ $Y2=0
cc_936 N_VPWR_M1020_d N_A_244_121#_c_1573_n 0.00221858f $X=4.525 $Y=2.415 $X2=0
+ $Y2=0
cc_937 N_VPWR_c_1392_n N_A_244_121#_c_1573_n 0.00877092f $X=4.665 $Y=2.93 $X2=0
+ $Y2=0
cc_938 N_VPWR_c_1389_n N_A_244_121#_c_1573_n 7.42495e-19 $X=15.12 $Y=3.33 $X2=0
+ $Y2=0
cc_939 N_VPWR_c_1394_n N_A_1781_379#_c_1699_n 0.0015231f $X=8.615 $Y=2.24 $X2=0
+ $Y2=0
cc_940 N_VPWR_c_1406_n N_A_1781_379#_c_1699_n 0.00674548f $X=11.53 $Y=3.33 $X2=0
+ $Y2=0
cc_941 N_VPWR_c_1389_n N_A_1781_379#_c_1699_n 0.00812916f $X=15.12 $Y=3.33 $X2=0
+ $Y2=0
cc_942 N_VPWR_c_1395_n N_A_1888_463#_c_1733_n 0.0147663f $X=11.655 $Y=2.44 $X2=0
+ $Y2=0
cc_943 N_VPWR_c_1406_n N_A_1888_463#_c_1733_n 0.062108f $X=11.53 $Y=3.33 $X2=0
+ $Y2=0
cc_944 N_VPWR_c_1389_n N_A_1888_463#_c_1733_n 0.0515665f $X=15.12 $Y=3.33 $X2=0
+ $Y2=0
cc_945 N_VPWR_c_1395_n N_A_1888_463#_c_1734_n 0.016086f $X=11.655 $Y=2.44 $X2=0
+ $Y2=0
cc_946 N_VPWR_c_1394_n N_A_1888_463#_c_1735_n 0.00644165f $X=8.615 $Y=2.24 $X2=0
+ $Y2=0
cc_947 N_VPWR_c_1406_n N_A_1888_463#_c_1735_n 0.0131563f $X=11.53 $Y=3.33 $X2=0
+ $Y2=0
cc_948 N_VPWR_c_1389_n N_A_1888_463#_c_1735_n 0.0104251f $X=15.12 $Y=3.33 $X2=0
+ $Y2=0
cc_949 N_VPWR_c_1389_n N_Q_M1028_s 0.00501859f $X=15.12 $Y=3.33 $X2=0 $Y2=0
cc_950 N_VPWR_c_1413_n N_Q_c_1779_n 0.0128073f $X=14.76 $Y=3.33 $X2=0 $Y2=0
cc_951 N_VPWR_c_1389_n N_Q_c_1779_n 0.00769778f $X=15.12 $Y=3.33 $X2=0 $Y2=0
cc_952 N_VPWR_M1039_d N_Q_c_1761_n 0.00305454f $X=14.785 $Y=1.835 $X2=0 $Y2=0
cc_953 N_VPWR_c_1397_n N_Q_c_1761_n 0.0480501f $X=13.985 $Y=1.99 $X2=0 $Y2=0
cc_954 N_VPWR_c_1399_n N_Q_c_1761_n 0.0243971f $X=14.925 $Y=2.25 $X2=0 $Y2=0
cc_955 N_A_244_121#_c_1575_n N_VGND_c_1790_n 0.0110409f $X=1.36 $Y=0.815 $X2=0
+ $Y2=0
cc_956 N_A_244_121#_c_1575_n N_VGND_c_1791_n 0.0116218f $X=1.36 $Y=0.815 $X2=0
+ $Y2=0
cc_957 N_A_244_121#_c_1559_n N_VGND_c_1791_n 0.0491888f $X=2.425 $Y=1.277 $X2=0
+ $Y2=0
cc_958 N_A_244_121#_c_1575_n N_VGND_c_1806_n 0.00498781f $X=1.36 $Y=0.815 $X2=0
+ $Y2=0
cc_959 N_A_244_121#_c_1575_n N_VGND_c_1814_n 0.00845247f $X=1.36 $Y=0.815 $X2=0
+ $Y2=0
cc_960 N_A_1781_379#_c_1697_n N_A_1888_463#_M1032_s 0.00504151f $X=10.51 $Y=2.36
+ $X2=-0.19 $Y2=1.655
cc_961 N_A_1781_379#_c_1697_n N_A_1888_463#_c_1733_n 0.0282341f $X=10.51 $Y=2.36
+ $X2=0 $Y2=0
cc_962 N_A_1781_379#_c_1700_n N_A_1888_463#_c_1733_n 0.0213549f $X=10.675
+ $Y=2.36 $X2=0 $Y2=0
cc_963 N_A_1781_379#_c_1700_n N_A_1888_463#_c_1734_n 0.0234394f $X=10.675
+ $Y=2.36 $X2=0 $Y2=0
cc_964 N_A_1781_379#_c_1697_n N_A_1888_463#_c_1735_n 0.0253593f $X=10.51 $Y=2.36
+ $X2=0 $Y2=0
cc_965 N_A_1781_379#_c_1699_n N_A_1888_463#_c_1735_n 0.00996867f $X=9.062
+ $Y=2.36 $X2=0 $Y2=0
cc_966 N_Q_c_1759_n N_VGND_M1036_d 0.0031624f $X=14.832 $Y=1.135 $X2=0 $Y2=0
cc_967 N_Q_c_1759_n N_VGND_c_1796_n 0.00139572f $X=14.832 $Y=1.135 $X2=0 $Y2=0
cc_968 N_Q_c_1759_n N_VGND_c_1798_n 0.0243264f $X=14.832 $Y=1.135 $X2=0 $Y2=0
cc_969 N_Q_c_1787_p N_VGND_c_1809_n 0.0128073f $X=14.495 $Y=0.42 $X2=0 $Y2=0
cc_970 N_Q_M1021_s N_VGND_c_1814_n 0.00501859f $X=14.355 $Y=0.235 $X2=0 $Y2=0
cc_971 N_Q_c_1787_p N_VGND_c_1814_n 0.00769778f $X=14.495 $Y=0.42 $X2=0 $Y2=0
cc_972 N_VGND_c_1794_n A_1608_125# 0.00202734f $X=8.05 $Y=0.81 $X2=-0.19
+ $Y2=-0.245
cc_973 N_VGND_c_1859_n A_1608_125# 4.54916e-19 $X=8.135 $Y=0.91 $X2=-0.19
+ $Y2=-0.245
cc_974 N_VGND_c_1846_n A_1608_125# 0.0017598f $X=9.375 $Y=0.905 $X2=-0.19
+ $Y2=-0.245
