* File: sky130_fd_sc_lp__nand2_8.pex.spice
* Created: Fri Aug 28 10:47:26 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__NAND2_8%B 3 7 11 15 19 23 27 31 35 39 43 47 51 55 59
+ 63 75 78 79 104 106 109 114 116 122
c147 63 0 1.29724e-19 $X=3.485 $Y=2.465
c148 59 0 1.30471e-19 $X=3.485 $Y=0.745
c149 55 0 4.60864e-20 $X=3.055 $Y=2.465
r150 106 114 0.434254 $w=3.43e-07 $l=1.3e-08 $layer=LI1_cond $X=2.653 $Y=1.587
+ $X2=2.64 $Y2=1.587
r151 101 106 0.233829 $w=3.43e-07 $l=7e-09 $layer=LI1_cond $X=2.66 $Y=1.587
+ $X2=2.653 $Y2=1.587
r152 100 102 69.0702 $w=3.3e-07 $l=3.95e-07 $layer=POLY_cond $X=2.66 $Y=1.51
+ $X2=3.055 $Y2=1.51
r153 100 101 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.66
+ $Y=1.51 $X2=2.66 $Y2=1.51
r154 98 100 6.12014 $w=3.3e-07 $l=3.5e-08 $layer=POLY_cond $X=2.625 $Y=1.51
+ $X2=2.66 $Y2=1.51
r155 96 98 53.3327 $w=3.3e-07 $l=3.05e-07 $layer=POLY_cond $X=2.32 $Y=1.51
+ $X2=2.625 $Y2=1.51
r156 96 97 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.32
+ $Y=1.51 $X2=2.32 $Y2=1.51
r157 94 96 21.8577 $w=3.3e-07 $l=1.25e-07 $layer=POLY_cond $X=2.195 $Y=1.51
+ $X2=2.32 $Y2=1.51
r158 93 116 8.13615 $w=3.43e-07 $l=1.65e-07 $layer=LI1_cond $X=1.98 $Y=1.587
+ $X2=1.815 $Y2=1.587
r159 92 94 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=1.98 $Y=1.51
+ $X2=2.195 $Y2=1.51
r160 92 93 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.98
+ $Y=1.51 $X2=1.98 $Y2=1.51
r161 90 92 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=1.765 $Y=1.51
+ $X2=1.98 $Y2=1.51
r162 87 88 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=0.905 $Y=1.51
+ $X2=1.335 $Y2=1.51
r163 79 122 6.8518 $w=3.43e-07 $l=1.36e-07 $layer=LI1_cond $X=2.689 $Y=1.587
+ $X2=2.825 $Y2=1.587
r164 79 101 0.96872 $w=3.43e-07 $l=2.9e-08 $layer=LI1_cond $X=2.689 $Y=1.587
+ $X2=2.66 $Y2=1.587
r165 79 114 1.20255 $w=3.43e-07 $l=3.6e-08 $layer=LI1_cond $X=2.604 $Y=1.587
+ $X2=2.64 $Y2=1.587
r166 79 97 9.48678 $w=3.43e-07 $l=2.84e-07 $layer=LI1_cond $X=2.604 $Y=1.587
+ $X2=2.32 $Y2=1.587
r167 78 109 1.43638 $w=3.43e-07 $l=4.3e-08 $layer=LI1_cond $X=2.117 $Y=1.587
+ $X2=2.16 $Y2=1.587
r168 78 93 4.57637 $w=3.43e-07 $l=1.37e-07 $layer=LI1_cond $X=2.117 $Y=1.587
+ $X2=1.98 $Y2=1.587
r169 78 97 3.94169 $w=3.43e-07 $l=1.18e-07 $layer=LI1_cond $X=2.202 $Y=1.587
+ $X2=2.32 $Y2=1.587
r170 78 109 1.40297 $w=3.43e-07 $l=4.2e-08 $layer=LI1_cond $X=2.202 $Y=1.587
+ $X2=2.16 $Y2=1.587
r171 76 104 25.3549 $w=3.3e-07 $l=1.45e-07 $layer=POLY_cond $X=3.34 $Y=1.51
+ $X2=3.485 $Y2=1.51
r172 76 102 49.8355 $w=3.3e-07 $l=2.85e-07 $layer=POLY_cond $X=3.34 $Y=1.51
+ $X2=3.055 $Y2=1.51
r173 75 122 30.0622 $w=1.88e-07 $l=5.15e-07 $layer=LI1_cond $X=3.34 $Y=1.51
+ $X2=2.825 $Y2=1.51
r174 75 76 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.34
+ $Y=1.51 $X2=3.34 $Y2=1.51
r175 72 90 21.8577 $w=3.3e-07 $l=1.25e-07 $layer=POLY_cond $X=1.64 $Y=1.51
+ $X2=1.765 $Y2=1.51
r176 72 88 53.3327 $w=3.3e-07 $l=3.05e-07 $layer=POLY_cond $X=1.64 $Y=1.51
+ $X2=1.335 $Y2=1.51
r177 71 116 10.7828 $w=1.78e-07 $l=1.75e-07 $layer=LI1_cond $X=1.64 $Y=1.505
+ $X2=1.815 $Y2=1.505
r178 71 72 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.64
+ $Y=1.51 $X2=1.64 $Y2=1.51
r179 68 87 49.8355 $w=3.3e-07 $l=2.85e-07 $layer=POLY_cond $X=0.62 $Y=1.51
+ $X2=0.905 $Y2=1.51
r180 68 84 25.3549 $w=3.3e-07 $l=1.45e-07 $layer=POLY_cond $X=0.62 $Y=1.51
+ $X2=0.475 $Y2=1.51
r181 67 71 62.8485 $w=1.78e-07 $l=1.02e-06 $layer=LI1_cond $X=0.62 $Y=1.505
+ $X2=1.64 $Y2=1.505
r182 67 68 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.62
+ $Y=1.51 $X2=0.62 $Y2=1.51
r183 61 104 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.485 $Y=1.675
+ $X2=3.485 $Y2=1.51
r184 61 63 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.485 $Y=1.675
+ $X2=3.485 $Y2=2.465
r185 57 104 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.485 $Y=1.345
+ $X2=3.485 $Y2=1.51
r186 57 59 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=3.485 $Y=1.345
+ $X2=3.485 $Y2=0.745
r187 53 102 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.055 $Y=1.675
+ $X2=3.055 $Y2=1.51
r188 53 55 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.055 $Y=1.675
+ $X2=3.055 $Y2=2.465
r189 49 102 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.055 $Y=1.345
+ $X2=3.055 $Y2=1.51
r190 49 51 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=3.055 $Y=1.345
+ $X2=3.055 $Y2=0.745
r191 45 98 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.625 $Y=1.675
+ $X2=2.625 $Y2=1.51
r192 45 47 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.625 $Y=1.675
+ $X2=2.625 $Y2=2.465
r193 41 98 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.625 $Y=1.345
+ $X2=2.625 $Y2=1.51
r194 41 43 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=2.625 $Y=1.345
+ $X2=2.625 $Y2=0.745
r195 37 94 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.195 $Y=1.675
+ $X2=2.195 $Y2=1.51
r196 37 39 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.195 $Y=1.675
+ $X2=2.195 $Y2=2.465
r197 33 94 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.195 $Y=1.345
+ $X2=2.195 $Y2=1.51
r198 33 35 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=2.195 $Y=1.345
+ $X2=2.195 $Y2=0.745
r199 29 90 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.765 $Y=1.675
+ $X2=1.765 $Y2=1.51
r200 29 31 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.765 $Y=1.675
+ $X2=1.765 $Y2=2.465
r201 25 90 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.765 $Y=1.345
+ $X2=1.765 $Y2=1.51
r202 25 27 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=1.765 $Y=1.345
+ $X2=1.765 $Y2=0.745
r203 21 88 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.335 $Y=1.675
+ $X2=1.335 $Y2=1.51
r204 21 23 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.335 $Y=1.675
+ $X2=1.335 $Y2=2.465
r205 17 88 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.335 $Y=1.345
+ $X2=1.335 $Y2=1.51
r206 17 19 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=1.335 $Y=1.345
+ $X2=1.335 $Y2=0.745
r207 13 87 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.905 $Y=1.675
+ $X2=0.905 $Y2=1.51
r208 13 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=0.905 $Y=1.675
+ $X2=0.905 $Y2=2.465
r209 9 87 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.905 $Y=1.345
+ $X2=0.905 $Y2=1.51
r210 9 11 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=0.905 $Y=1.345
+ $X2=0.905 $Y2=0.745
r211 5 84 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=1.675
+ $X2=0.475 $Y2=1.51
r212 5 7 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=0.475 $Y=1.675
+ $X2=0.475 $Y2=2.465
r213 1 84 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=1.345
+ $X2=0.475 $Y2=1.51
r214 1 3 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=0.475 $Y=1.345 $X2=0.475
+ $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_LP__NAND2_8%A 3 7 11 15 19 23 25 29 33 37 41 45 49 53 57
+ 61 65 67 71 72 73 77 79 80 81 91 93
r147 93 94 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.275
+ $Y=1.51 $X2=5.275 $Y2=1.51
r148 90 91 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.615
+ $Y=1.51 $X2=5.615 $Y2=1.51
r149 88 93 10.9545 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=5.42 $Y=1.51
+ $X2=5.345 $Y2=1.51
r150 88 90 34.0979 $w=3.3e-07 $l=1.95e-07 $layer=POLY_cond $X=5.42 $Y=1.51
+ $X2=5.615 $Y2=1.51
r151 86 87 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.595
+ $Y=1.51 $X2=4.595 $Y2=1.51
r152 81 91 3.26812 $w=3.33e-07 $l=9.5e-08 $layer=LI1_cond $X=5.52 $Y=1.592
+ $X2=5.615 $Y2=1.592
r153 81 94 8.42831 $w=3.33e-07 $l=2.45e-07 $layer=LI1_cond $X=5.52 $Y=1.592
+ $X2=5.275 $Y2=1.592
r154 80 94 8.0843 $w=3.33e-07 $l=2.35e-07 $layer=LI1_cond $X=5.04 $Y=1.592
+ $X2=5.275 $Y2=1.592
r155 80 87 15.3086 $w=3.33e-07 $l=4.45e-07 $layer=LI1_cond $X=5.04 $Y=1.592
+ $X2=4.595 $Y2=1.592
r156 79 87 1.20404 $w=3.33e-07 $l=3.5e-08 $layer=LI1_cond $X=4.56 $Y=1.592
+ $X2=4.595 $Y2=1.592
r157 76 77 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=6.735 $Y=1.51
+ $X2=7.165 $Y2=1.51
r158 75 76 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=6.305 $Y=1.51
+ $X2=6.735 $Y2=1.51
r159 74 75 80.4362 $w=3.3e-07 $l=4.6e-07 $layer=POLY_cond $X=5.845 $Y=1.51
+ $X2=6.305 $Y2=1.51
r160 73 90 27.1035 $w=3.3e-07 $l=1.55e-07 $layer=POLY_cond $X=5.77 $Y=1.51
+ $X2=5.615 $Y2=1.51
r161 73 74 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=5.77 $Y=1.51
+ $X2=5.845 $Y2=1.51
r162 71 86 30.6007 $w=3.3e-07 $l=1.75e-07 $layer=POLY_cond $X=4.77 $Y=1.51
+ $X2=4.595 $Y2=1.51
r163 71 72 10.9545 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=4.77 $Y=1.51
+ $X2=4.845 $Y2=1.51
r164 68 70 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=3.915 $Y=1.51
+ $X2=4.345 $Y2=1.51
r165 67 86 30.6007 $w=3.3e-07 $l=1.75e-07 $layer=POLY_cond $X=4.42 $Y=1.51
+ $X2=4.595 $Y2=1.51
r166 67 70 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=4.42 $Y=1.51
+ $X2=4.345 $Y2=1.51
r167 63 77 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.165 $Y=1.675
+ $X2=7.165 $Y2=1.51
r168 63 65 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=7.165 $Y=1.675
+ $X2=7.165 $Y2=2.465
r169 59 77 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.165 $Y=1.345
+ $X2=7.165 $Y2=1.51
r170 59 61 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=7.165 $Y=1.345
+ $X2=7.165 $Y2=0.745
r171 55 76 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.735 $Y=1.675
+ $X2=6.735 $Y2=1.51
r172 55 57 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=6.735 $Y=1.675
+ $X2=6.735 $Y2=2.465
r173 51 76 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.735 $Y=1.345
+ $X2=6.735 $Y2=1.51
r174 51 53 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=6.735 $Y=1.345
+ $X2=6.735 $Y2=0.745
r175 47 75 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.305 $Y=1.675
+ $X2=6.305 $Y2=1.51
r176 47 49 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=6.305 $Y=1.675
+ $X2=6.305 $Y2=2.465
r177 43 75 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.305 $Y=1.345
+ $X2=6.305 $Y2=1.51
r178 43 45 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=6.305 $Y=1.345
+ $X2=6.305 $Y2=0.745
r179 39 74 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.845 $Y=1.675
+ $X2=5.845 $Y2=1.51
r180 39 41 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=5.845 $Y=1.675
+ $X2=5.845 $Y2=2.465
r181 35 74 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.845 $Y=1.345
+ $X2=5.845 $Y2=1.51
r182 35 37 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=5.845 $Y=1.345
+ $X2=5.845 $Y2=0.745
r183 31 93 53.02 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.345 $Y=1.675
+ $X2=5.345 $Y2=1.51
r184 31 33 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=5.345 $Y=1.675
+ $X2=5.345 $Y2=2.465
r185 27 93 53.02 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.345 $Y=1.345
+ $X2=5.345 $Y2=1.51
r186 27 29 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=5.345 $Y=1.345
+ $X2=5.345 $Y2=0.745
r187 26 72 10.9545 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=4.92 $Y=1.51
+ $X2=4.845 $Y2=1.51
r188 25 93 10.9545 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=5.27 $Y=1.51
+ $X2=5.345 $Y2=1.51
r189 25 26 61.2015 $w=3.3e-07 $l=3.5e-07 $layer=POLY_cond $X=5.27 $Y=1.51
+ $X2=4.92 $Y2=1.51
r190 21 72 53.02 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.845 $Y=1.675
+ $X2=4.845 $Y2=1.51
r191 21 23 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=4.845 $Y=1.675
+ $X2=4.845 $Y2=2.465
r192 17 72 53.02 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.845 $Y=1.345
+ $X2=4.845 $Y2=1.51
r193 17 19 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=4.845 $Y=1.345
+ $X2=4.845 $Y2=0.745
r194 13 70 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.345 $Y=1.675
+ $X2=4.345 $Y2=1.51
r195 13 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=4.345 $Y=1.675
+ $X2=4.345 $Y2=2.465
r196 9 70 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.345 $Y=1.345
+ $X2=4.345 $Y2=1.51
r197 9 11 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=4.345 $Y=1.345
+ $X2=4.345 $Y2=0.745
r198 5 68 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.915 $Y=1.675
+ $X2=3.915 $Y2=1.51
r199 5 7 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.915 $Y=1.675
+ $X2=3.915 $Y2=2.465
r200 1 68 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.915 $Y=1.345
+ $X2=3.915 $Y2=1.51
r201 1 3 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=3.915 $Y=1.345 $X2=3.915
+ $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_LP__NAND2_8%VPWR 1 2 3 4 5 6 7 8 9 28 30 36 42 46 48 52
+ 58 62 66 70 72 77 78 79 80 81 83 95 100 105 110 119 122 125 128 131 135
r131 134 135 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r132 131 132 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r133 128 129 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r134 125 126 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r135 122 123 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r136 119 120 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r137 116 117 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r138 114 135 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=7.44 $Y2=3.33
r139 114 132 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=6.48 $Y2=3.33
r140 113 114 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r141 111 131 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.685 $Y=3.33
+ $X2=6.52 $Y2=3.33
r142 111 113 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=6.685 $Y=3.33
+ $X2=6.96 $Y2=3.33
r143 110 134 3.63768 $w=1.7e-07 $l=2.02e-07 $layer=LI1_cond $X=7.275 $Y=3.33
+ $X2=7.477 $Y2=3.33
r144 110 113 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=7.275 $Y=3.33
+ $X2=6.96 $Y2=3.33
r145 109 132 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33
+ $X2=6.48 $Y2=3.33
r146 109 129 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33
+ $X2=5.52 $Y2=3.33
r147 108 109 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r148 106 128 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.76 $Y=3.33
+ $X2=5.595 $Y2=3.33
r149 106 108 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=5.76 $Y=3.33
+ $X2=6 $Y2=3.33
r150 105 131 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.355 $Y=3.33
+ $X2=6.52 $Y2=3.33
r151 105 108 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=6.355 $Y=3.33
+ $X2=6 $Y2=3.33
r152 104 129 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=5.52 $Y2=3.33
r153 104 126 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=4.56 $Y2=3.33
r154 103 104 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r155 101 125 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.76 $Y=3.33
+ $X2=4.595 $Y2=3.33
r156 101 103 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=4.76 $Y=3.33
+ $X2=5.04 $Y2=3.33
r157 100 128 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.43 $Y=3.33
+ $X2=5.595 $Y2=3.33
r158 100 103 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=5.43 $Y=3.33
+ $X2=5.04 $Y2=3.33
r159 99 126 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r160 98 99 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r161 96 122 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.865 $Y=3.33
+ $X2=3.7 $Y2=3.33
r162 96 98 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=3.865 $Y=3.33
+ $X2=4.08 $Y2=3.33
r163 95 125 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.43 $Y=3.33
+ $X2=4.595 $Y2=3.33
r164 95 98 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=4.43 $Y=3.33
+ $X2=4.08 $Y2=3.33
r165 94 123 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r166 93 94 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r167 91 94 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r168 91 120 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r169 90 91 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r170 88 119 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.285 $Y=3.33
+ $X2=1.12 $Y2=3.33
r171 88 90 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=1.285 $Y=3.33
+ $X2=1.68 $Y2=3.33
r172 87 120 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r173 87 117 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r174 86 87 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r175 84 116 4.78091 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=3.33
+ $X2=0.212 $Y2=3.33
r176 84 86 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.425 $Y=3.33
+ $X2=0.72 $Y2=3.33
r177 83 119 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.955 $Y=3.33
+ $X2=1.12 $Y2=3.33
r178 83 86 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=0.955 $Y=3.33
+ $X2=0.72 $Y2=3.33
r179 81 99 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.84 $Y=3.33
+ $X2=4.08 $Y2=3.33
r180 81 123 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.84 $Y=3.33
+ $X2=3.6 $Y2=3.33
r181 79 93 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=2.675 $Y=3.33
+ $X2=2.64 $Y2=3.33
r182 79 80 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.675 $Y=3.33
+ $X2=2.84 $Y2=3.33
r183 77 90 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=1.815 $Y=3.33
+ $X2=1.68 $Y2=3.33
r184 77 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.815 $Y=3.33
+ $X2=1.98 $Y2=3.33
r185 76 93 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=2.145 $Y=3.33
+ $X2=2.64 $Y2=3.33
r186 76 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.145 $Y=3.33
+ $X2=1.98 $Y2=3.33
r187 72 75 51.2294 $w=2.08e-07 $l=9.7e-07 $layer=LI1_cond $X=7.38 $Y=1.98
+ $X2=7.38 $Y2=2.95
r188 70 134 3.27751 $w=2.1e-07 $l=1.32868e-07 $layer=LI1_cond $X=7.38 $Y=3.245
+ $X2=7.477 $Y2=3.33
r189 70 75 15.5801 $w=2.08e-07 $l=2.95e-07 $layer=LI1_cond $X=7.38 $Y=3.245
+ $X2=7.38 $Y2=2.95
r190 66 69 26.8903 $w=3.28e-07 $l=7.7e-07 $layer=LI1_cond $X=6.52 $Y=2.18
+ $X2=6.52 $Y2=2.95
r191 64 131 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.52 $Y=3.245
+ $X2=6.52 $Y2=3.33
r192 64 69 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=6.52 $Y=3.245
+ $X2=6.52 $Y2=2.95
r193 60 128 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.595 $Y=3.245
+ $X2=5.595 $Y2=3.33
r194 60 62 31.081 $w=3.28e-07 $l=8.9e-07 $layer=LI1_cond $X=5.595 $Y=3.245
+ $X2=5.595 $Y2=2.355
r195 56 125 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.595 $Y=3.245
+ $X2=4.595 $Y2=3.33
r196 56 58 31.081 $w=3.28e-07 $l=8.9e-07 $layer=LI1_cond $X=4.595 $Y=3.245
+ $X2=4.595 $Y2=2.355
r197 52 55 26.8903 $w=3.28e-07 $l=7.7e-07 $layer=LI1_cond $X=3.7 $Y=2.2 $X2=3.7
+ $Y2=2.97
r198 50 122 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.7 $Y=3.245
+ $X2=3.7 $Y2=3.33
r199 50 55 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=3.7 $Y=3.245
+ $X2=3.7 $Y2=2.97
r200 49 80 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.005 $Y=3.33
+ $X2=2.84 $Y2=3.33
r201 48 122 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.535 $Y=3.33
+ $X2=3.7 $Y2=3.33
r202 48 49 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=3.535 $Y=3.33
+ $X2=3.005 $Y2=3.33
r203 44 80 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.84 $Y=3.245
+ $X2=2.84 $Y2=3.33
r204 44 46 31.081 $w=3.28e-07 $l=8.9e-07 $layer=LI1_cond $X=2.84 $Y=3.245
+ $X2=2.84 $Y2=2.355
r205 40 78 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.98 $Y=3.245
+ $X2=1.98 $Y2=3.33
r206 40 42 31.081 $w=3.28e-07 $l=8.9e-07 $layer=LI1_cond $X=1.98 $Y=3.245
+ $X2=1.98 $Y2=2.355
r207 36 39 26.5411 $w=3.28e-07 $l=7.6e-07 $layer=LI1_cond $X=1.12 $Y=2.19
+ $X2=1.12 $Y2=2.95
r208 34 119 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.12 $Y=3.245
+ $X2=1.12 $Y2=3.33
r209 34 39 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.12 $Y=3.245
+ $X2=1.12 $Y2=2.95
r210 30 33 33.7002 $w=3.28e-07 $l=9.65e-07 $layer=LI1_cond $X=0.26 $Y=1.985
+ $X2=0.26 $Y2=2.95
r211 28 116 2.98526 $w=3.3e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.26 $Y=3.245
+ $X2=0.212 $Y2=3.33
r212 28 33 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.26 $Y=3.245
+ $X2=0.26 $Y2=2.95
r213 9 75 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=7.24
+ $Y=1.835 $X2=7.38 $Y2=2.95
r214 9 72 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=7.24
+ $Y=1.835 $X2=7.38 $Y2=1.98
r215 8 69 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=6.38
+ $Y=1.835 $X2=6.52 $Y2=2.95
r216 8 66 400 $w=1.7e-07 $l=4.09054e-07 $layer=licon1_PDIFF $count=1 $X=6.38
+ $Y=1.835 $X2=6.52 $Y2=2.18
r217 7 62 300 $w=1.7e-07 $l=6.01166e-07 $layer=licon1_PDIFF $count=2 $X=5.42
+ $Y=1.835 $X2=5.595 $Y2=2.355
r218 6 58 300 $w=1.7e-07 $l=6.01166e-07 $layer=licon1_PDIFF $count=2 $X=4.42
+ $Y=1.835 $X2=4.595 $Y2=2.355
r219 5 55 400 $w=1.7e-07 $l=1.20297e-06 $layer=licon1_PDIFF $count=1 $X=3.56
+ $Y=1.835 $X2=3.7 $Y2=2.97
r220 5 52 400 $w=1.7e-07 $l=4.29331e-07 $layer=licon1_PDIFF $count=1 $X=3.56
+ $Y=1.835 $X2=3.7 $Y2=2.2
r221 4 46 300 $w=1.7e-07 $l=5.85833e-07 $layer=licon1_PDIFF $count=2 $X=2.7
+ $Y=1.835 $X2=2.84 $Y2=2.355
r222 3 42 300 $w=1.7e-07 $l=5.85833e-07 $layer=licon1_PDIFF $count=2 $X=1.84
+ $Y=1.835 $X2=1.98 $Y2=2.355
r223 2 39 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=0.98
+ $Y=1.835 $X2=1.12 $Y2=2.95
r224 2 36 400 $w=1.7e-07 $l=4.19196e-07 $layer=licon1_PDIFF $count=1 $X=0.98
+ $Y=1.835 $X2=1.12 $Y2=2.19
r225 1 33 400 $w=1.7e-07 $l=1.17584e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.835 $X2=0.26 $Y2=2.95
r226 1 30 400 $w=1.7e-07 $l=2.03101e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.835 $X2=0.26 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_LP__NAND2_8%Y 1 2 3 4 5 6 7 8 9 10 11 12 39 43 44 45 47
+ 49 53 55 59 61 63 65 67 69 73 77 79 81 85 89 93 97 106 107 119 120 125 127 128
+ 129 136 142
c154 128 0 2.83085e-19 $X=3.995 $Y=1.21
c155 107 0 1.29724e-19 $X=3.245 $Y=1.86
c156 61 0 4.60864e-20 $X=3.965 $Y=1.86
r157 140 142 1.56263 $w=2.93e-07 $l=4e-08 $layer=LI1_cond $X=4.112 $Y=1.255
+ $X2=4.112 $Y2=1.295
r158 128 134 3.03453 $w=3.12e-07 $l=8.5e-08 $layer=LI1_cond $X=4.13 $Y=1.17
+ $X2=4.13 $Y2=1.085
r159 128 140 3.03453 $w=3.12e-07 $l=9.35682e-08 $layer=LI1_cond $X=4.13 $Y=1.17
+ $X2=4.112 $Y2=1.255
r160 128 129 13.5949 $w=2.93e-07 $l=3.48e-07 $layer=LI1_cond $X=4.112 $Y=1.317
+ $X2=4.112 $Y2=1.665
r161 128 142 0.859449 $w=2.93e-07 $l=2.2e-08 $layer=LI1_cond $X=4.112 $Y=1.317
+ $X2=4.112 $Y2=1.295
r162 127 134 5.5876 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=4.13 $Y=0.925
+ $X2=4.13 $Y2=1.085
r163 127 136 7.85757 $w=3.28e-07 $l=2.25e-07 $layer=LI1_cond $X=4.13 $Y=0.925
+ $X2=4.13 $Y2=0.7
r164 124 125 13.0682 $w=8.01e-07 $l=8.58e-07 $layer=LI1_cond $X=6.092 $Y=1.587
+ $X2=6.95 $Y2=1.587
r165 123 124 0.0304619 $w=8.01e-07 $l=2e-09 $layer=LI1_cond $X=6.09 $Y=1.587
+ $X2=6.092 $Y2=1.587
r166 121 123 0.350312 $w=8.01e-07 $l=2.3e-08 $layer=LI1_cond $X=6.067 $Y=1.587
+ $X2=6.09 $Y2=1.587
r167 116 117 1.63602 $w=2.61e-07 $l=3.5e-08 $layer=LI1_cond $X=4.112 $Y=1.98
+ $X2=4.112 $Y2=2.015
r168 114 116 5.6092 $w=2.61e-07 $l=1.2e-07 $layer=LI1_cond $X=4.112 $Y=1.86
+ $X2=4.112 $Y2=1.98
r169 113 129 4.29725 $w=2.93e-07 $l=1.1e-07 $layer=LI1_cond $X=4.112 $Y=1.775
+ $X2=4.112 $Y2=1.665
r170 113 114 3.70728 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=4.112 $Y=1.775
+ $X2=4.112 $Y2=1.86
r171 111 112 4.6142 $w=2.38e-07 $l=8.5e-08 $layer=LI1_cond $X=3.245 $Y=2.015
+ $X2=3.245 $Y2=2.1
r172 110 111 1.68065 $w=2.38e-07 $l=3.5e-08 $layer=LI1_cond $X=3.245 $Y=1.98
+ $X2=3.245 $Y2=2.015
r173 107 110 5.76222 $w=2.38e-07 $l=1.2e-07 $layer=LI1_cond $X=3.245 $Y=1.86
+ $X2=3.245 $Y2=1.98
r174 103 104 2.30811 $w=1.85e-07 $l=3.5e-08 $layer=LI1_cond $X=1.55 $Y=1.98
+ $X2=1.55 $Y2=2.015
r175 101 103 8.57297 $w=1.85e-07 $l=1.3e-07 $layer=LI1_cond $X=1.55 $Y=1.85
+ $X2=1.55 $Y2=1.98
r176 97 99 51.5727 $w=1.98e-07 $l=9.3e-07 $layer=LI1_cond $X=6.955 $Y=1.98
+ $X2=6.955 $Y2=2.91
r177 95 125 0.0761548 $w=8.01e-07 $l=5e-09 $layer=LI1_cond $X=6.955 $Y=1.587
+ $X2=6.95 $Y2=1.587
r178 95 97 3.05 $w=1.98e-07 $l=5.5e-08 $layer=LI1_cond $X=6.955 $Y=1.925
+ $X2=6.955 $Y2=1.98
r179 91 125 5.96787 $w=3.3e-07 $l=4.32e-07 $layer=LI1_cond $X=6.95 $Y=1.155
+ $X2=6.95 $Y2=1.587
r180 91 93 15.8897 $w=3.28e-07 $l=4.55e-07 $layer=LI1_cond $X=6.95 $Y=1.155
+ $X2=6.95 $Y2=0.7
r181 87 124 7.57933 $w=2.55e-07 $l=5.12e-07 $layer=LI1_cond $X=6.092 $Y=1.075
+ $X2=6.092 $Y2=1.587
r182 87 89 12.2023 $w=2.53e-07 $l=2.7e-07 $layer=LI1_cond $X=6.092 $Y=1.075
+ $X2=6.092 $Y2=0.805
r183 83 121 8.10022 $w=2.35e-07 $l=5.13e-07 $layer=LI1_cond $X=6.067 $Y=2.1
+ $X2=6.067 $Y2=1.587
r184 83 85 17.4092 $w=2.33e-07 $l=3.55e-07 $layer=LI1_cond $X=6.067 $Y=2.1
+ $X2=6.067 $Y2=2.455
r185 82 120 8.43672 $w=1.75e-07 $l=1.65e-07 $layer=LI1_cond $X=5.295 $Y=1.165
+ $X2=5.13 $Y2=1.165
r186 81 121 4.44152 $w=4e-07 $l=4.76926e-07 $layer=LI1_cond $X=5.95 $Y=1.165
+ $X2=6.067 $Y2=1.587
r187 81 82 40.3586 $w=1.78e-07 $l=6.55e-07 $layer=LI1_cond $X=5.95 $Y=1.165
+ $X2=5.295 $Y2=1.165
r188 80 119 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.26 $Y=2.015
+ $X2=5.095 $Y2=2.015
r189 79 121 4.54752 $w=4e-07 $l=4.8297e-07 $layer=LI1_cond $X=5.95 $Y=2.015
+ $X2=6.067 $Y2=1.587
r190 79 80 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=5.95 $Y=2.015
+ $X2=5.26 $Y2=2.015
r191 75 120 0.806278 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=5.13 $Y=1.075
+ $X2=5.13 $Y2=1.165
r192 75 77 13.0959 $w=3.28e-07 $l=3.75e-07 $layer=LI1_cond $X=5.13 $Y=1.075
+ $X2=5.13 $Y2=0.7
r193 71 119 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.095 $Y=2.1
+ $X2=5.095 $Y2=2.015
r194 71 73 28.2872 $w=3.28e-07 $l=8.1e-07 $layer=LI1_cond $X=5.095 $Y=2.1
+ $X2=5.095 $Y2=2.91
r195 70 128 3.60271 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.295 $Y=1.17
+ $X2=4.13 $Y2=1.17
r196 69 120 8.43672 $w=1.75e-07 $l=1.67481e-07 $layer=LI1_cond $X=4.965 $Y=1.17
+ $X2=5.13 $Y2=1.165
r197 69 70 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.965 $Y=1.17
+ $X2=4.295 $Y2=1.17
r198 68 117 3.24614 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=4.26 $Y=2.015
+ $X2=4.112 $Y2=2.015
r199 67 119 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.93 $Y=2.015
+ $X2=5.095 $Y2=2.015
r200 67 68 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.93 $Y=2.015
+ $X2=4.26 $Y2=2.015
r201 63 117 4.23897 $w=2.61e-07 $l=1.00995e-07 $layer=LI1_cond $X=4.147 $Y=2.1
+ $X2=4.112 $Y2=2.015
r202 63 65 18.4391 $w=2.23e-07 $l=3.6e-07 $layer=LI1_cond $X=4.147 $Y=2.1
+ $X2=4.147 $Y2=2.46
r203 62 107 2.75731 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=3.365 $Y=1.86
+ $X2=3.245 $Y2=1.86
r204 61 114 3.24614 $w=1.7e-07 $l=1.47e-07 $layer=LI1_cond $X=3.965 $Y=1.86
+ $X2=4.112 $Y2=1.86
r205 61 62 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=3.965 $Y=1.86
+ $X2=3.365 $Y2=1.86
r206 59 112 21.0144 $w=1.88e-07 $l=3.6e-07 $layer=LI1_cond $X=3.27 $Y=2.46
+ $X2=3.27 $Y2=2.1
r207 56 106 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.505 $Y=2.015
+ $X2=2.41 $Y2=2.015
r208 55 111 2.75731 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=3.125 $Y=2.015
+ $X2=3.245 $Y2=2.015
r209 55 56 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=3.125 $Y=2.015
+ $X2=2.505 $Y2=2.015
r210 51 106 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=2.41 $Y=2.1
+ $X2=2.41 $Y2=2.015
r211 51 53 47.2823 $w=1.88e-07 $l=8.1e-07 $layer=LI1_cond $X=2.41 $Y=2.1
+ $X2=2.41 $Y2=2.91
r212 50 104 1.22693 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.645 $Y=2.015
+ $X2=1.55 $Y2=2.015
r213 49 106 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.315 $Y=2.015
+ $X2=2.41 $Y2=2.015
r214 49 50 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.315 $Y=2.015
+ $X2=1.645 $Y2=2.015
r215 45 104 5.45789 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.55 $Y=2.1
+ $X2=1.55 $Y2=2.015
r216 45 47 21.0144 $w=1.88e-07 $l=3.6e-07 $layer=LI1_cond $X=1.55 $Y=2.1
+ $X2=1.55 $Y2=2.46
r217 43 101 1.22693 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.455 $Y=1.85
+ $X2=1.55 $Y2=1.85
r218 43 44 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.455 $Y=1.85
+ $X2=0.785 $Y2=1.85
r219 39 41 54.2871 $w=1.88e-07 $l=9.3e-07 $layer=LI1_cond $X=0.69 $Y=1.98
+ $X2=0.69 $Y2=2.91
r220 37 44 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=0.69 $Y=1.935
+ $X2=0.785 $Y2=1.85
r221 37 39 2.62679 $w=1.88e-07 $l=4.5e-08 $layer=LI1_cond $X=0.69 $Y=1.935
+ $X2=0.69 $Y2=1.98
r222 12 99 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=6.81
+ $Y=1.835 $X2=6.95 $Y2=2.91
r223 12 97 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=6.81
+ $Y=1.835 $X2=6.95 $Y2=1.98
r224 11 123 600 $w=1.7e-07 $l=2.31409e-07 $layer=licon1_PDIFF $count=1 $X=5.92
+ $Y=1.835 $X2=6.09 $Y2=1.98
r225 11 85 300 $w=1.7e-07 $l=6.99857e-07 $layer=licon1_PDIFF $count=2 $X=5.92
+ $Y=1.835 $X2=6.09 $Y2=2.455
r226 10 119 400 $w=1.7e-07 $l=3.36303e-07 $layer=licon1_PDIFF $count=1 $X=4.92
+ $Y=1.835 $X2=5.095 $Y2=2.095
r227 10 73 400 $w=1.7e-07 $l=1.1592e-06 $layer=licon1_PDIFF $count=1 $X=4.92
+ $Y=1.835 $X2=5.095 $Y2=2.91
r228 9 116 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=3.99
+ $Y=1.835 $X2=4.13 $Y2=1.98
r229 9 65 300 $w=1.7e-07 $l=6.91466e-07 $layer=licon1_PDIFF $count=2 $X=3.99
+ $Y=1.835 $X2=4.13 $Y2=2.46
r230 8 110 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=3.13
+ $Y=1.835 $X2=3.27 $Y2=1.98
r231 8 59 300 $w=1.7e-07 $l=6.91466e-07 $layer=licon1_PDIFF $count=2 $X=3.13
+ $Y=1.835 $X2=3.27 $Y2=2.46
r232 7 106 400 $w=1.7e-07 $l=3.2249e-07 $layer=licon1_PDIFF $count=1 $X=2.27
+ $Y=1.835 $X2=2.41 $Y2=2.095
r233 7 53 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=2.27
+ $Y=1.835 $X2=2.41 $Y2=2.91
r234 6 103 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.41
+ $Y=1.835 $X2=1.55 $Y2=1.98
r235 6 47 300 $w=1.7e-07 $l=6.91466e-07 $layer=licon1_PDIFF $count=2 $X=1.41
+ $Y=1.835 $X2=1.55 $Y2=2.46
r236 5 41 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=1.835 $X2=0.69 $Y2=2.91
r237 5 39 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=1.835 $X2=0.69 $Y2=1.98
r238 4 93 91 $w=1.7e-07 $l=4.3946e-07 $layer=licon1_NDIFF $count=2 $X=6.81
+ $Y=0.325 $X2=6.95 $Y2=0.7
r239 3 89 182 $w=1.7e-07 $l=5.5857e-07 $layer=licon1_NDIFF $count=1 $X=5.92
+ $Y=0.325 $X2=6.09 $Y2=0.805
r240 2 77 91 $w=1.7e-07 $l=4.68375e-07 $layer=licon1_NDIFF $count=2 $X=4.92
+ $Y=0.325 $X2=5.13 $Y2=0.7
r241 1 136 91 $w=1.7e-07 $l=4.3946e-07 $layer=licon1_NDIFF $count=2 $X=3.99
+ $Y=0.325 $X2=4.13 $Y2=0.7
.ends

.subckt PM_SKY130_FD_SC_LP__NAND2_8%A_27_65# 1 2 3 4 5 6 7 8 9 30 32 33 36 38 42
+ 44 48 50 56 57 60 62 66 68 72 74 78 80 81 82 83 84 85
r132 76 78 1.55137 $w=2.58e-07 $l=3.5e-08 $layer=LI1_cond $X=7.415 $Y=0.435
+ $X2=7.415 $Y2=0.47
r133 75 85 6.19399 $w=1.8e-07 $l=1.13e-07 $layer=LI1_cond $X=6.615 $Y=0.345
+ $X2=6.502 $Y2=0.345
r134 74 76 7.11373 $w=1.8e-07 $l=1.69115e-07 $layer=LI1_cond $X=7.285 $Y=0.345
+ $X2=7.415 $Y2=0.435
r135 74 75 41.2828 $w=1.78e-07 $l=6.7e-07 $layer=LI1_cond $X=7.285 $Y=0.345
+ $X2=6.615 $Y2=0.345
r136 70 85 0.552779 $w=2.25e-07 $l=9e-08 $layer=LI1_cond $X=6.502 $Y=0.435
+ $X2=6.502 $Y2=0.345
r137 70 72 0.768295 $w=2.23e-07 $l=1.5e-08 $layer=LI1_cond $X=6.502 $Y=0.435
+ $X2=6.502 $Y2=0.45
r138 69 84 8.43672 $w=1.75e-07 $l=1.65e-07 $layer=LI1_cond $X=5.795 $Y=0.345
+ $X2=5.63 $Y2=0.345
r139 68 85 6.19399 $w=1.8e-07 $l=1.12e-07 $layer=LI1_cond $X=6.39 $Y=0.345
+ $X2=6.502 $Y2=0.345
r140 68 69 36.6616 $w=1.78e-07 $l=5.95e-07 $layer=LI1_cond $X=6.39 $Y=0.345
+ $X2=5.795 $Y2=0.345
r141 64 84 0.806278 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=5.63 $Y=0.435
+ $X2=5.63 $Y2=0.345
r142 64 66 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=5.63 $Y=0.435
+ $X2=5.63 $Y2=0.45
r143 63 83 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.795 $Y=0.34
+ $X2=4.63 $Y2=0.34
r144 62 84 8.43672 $w=1.75e-07 $l=1.67481e-07 $layer=LI1_cond $X=5.465 $Y=0.34
+ $X2=5.63 $Y2=0.345
r145 62 63 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.465 $Y=0.34
+ $X2=4.795 $Y2=0.34
r146 58 83 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.63 $Y=0.425
+ $X2=4.63 $Y2=0.34
r147 58 60 0.873063 $w=3.28e-07 $l=2.5e-08 $layer=LI1_cond $X=4.63 $Y=0.425
+ $X2=4.63 $Y2=0.45
r148 56 83 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.465 $Y=0.34
+ $X2=4.63 $Y2=0.34
r149 56 57 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.465 $Y=0.34
+ $X2=3.795 $Y2=0.34
r150 53 55 35.3158 $w=1.88e-07 $l=6.05e-07 $layer=LI1_cond $X=3.7 $Y=1.075
+ $X2=3.7 $Y2=0.47
r151 52 57 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=3.7 $Y=0.425
+ $X2=3.795 $Y2=0.34
r152 52 55 2.62679 $w=1.88e-07 $l=4.5e-08 $layer=LI1_cond $X=3.7 $Y=0.425
+ $X2=3.7 $Y2=0.47
r153 51 82 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.935 $Y=1.16
+ $X2=2.84 $Y2=1.16
r154 50 53 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=3.605 $Y=1.16
+ $X2=3.7 $Y2=1.075
r155 50 51 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.605 $Y=1.16
+ $X2=2.935 $Y2=1.16
r156 46 82 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=2.84 $Y=1.075
+ $X2=2.84 $Y2=1.16
r157 46 48 35.3158 $w=1.88e-07 $l=6.05e-07 $layer=LI1_cond $X=2.84 $Y=1.075
+ $X2=2.84 $Y2=0.47
r158 45 81 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.075 $Y=1.16
+ $X2=1.98 $Y2=1.16
r159 44 82 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.745 $Y=1.16
+ $X2=2.84 $Y2=1.16
r160 44 45 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.745 $Y=1.16
+ $X2=2.075 $Y2=1.16
r161 40 81 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.98 $Y=1.075
+ $X2=1.98 $Y2=1.16
r162 40 42 35.3158 $w=1.88e-07 $l=6.05e-07 $layer=LI1_cond $X=1.98 $Y=1.075
+ $X2=1.98 $Y2=0.47
r163 39 80 5.41628 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=1.205 $Y=1.16
+ $X2=1.115 $Y2=1.16
r164 38 81 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.885 $Y=1.16
+ $X2=1.98 $Y2=1.16
r165 38 39 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.885 $Y=1.16
+ $X2=1.205 $Y2=1.16
r166 34 80 1.13756 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=1.115 $Y=1.075
+ $X2=1.115 $Y2=1.16
r167 34 36 37.2778 $w=1.78e-07 $l=6.05e-07 $layer=LI1_cond $X=1.115 $Y=1.075
+ $X2=1.115 $Y2=0.47
r168 32 80 5.41628 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=1.025 $Y=1.16
+ $X2=1.115 $Y2=1.16
r169 32 33 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.025 $Y=1.16
+ $X2=0.355 $Y2=1.16
r170 28 33 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=0.225 $Y=1.075
+ $X2=0.355 $Y2=1.16
r171 28 30 26.8165 $w=2.58e-07 $l=6.05e-07 $layer=LI1_cond $X=0.225 $Y=1.075
+ $X2=0.225 $Y2=0.47
r172 9 78 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=7.24
+ $Y=0.325 $X2=7.38 $Y2=0.47
r173 8 72 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=6.38
+ $Y=0.325 $X2=6.52 $Y2=0.45
r174 7 66 91 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=2 $X=5.42
+ $Y=0.325 $X2=5.63 $Y2=0.45
r175 6 60 91 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=2 $X=4.42
+ $Y=0.325 $X2=4.63 $Y2=0.45
r176 5 55 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.56
+ $Y=0.325 $X2=3.7 $Y2=0.47
r177 4 48 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.7
+ $Y=0.325 $X2=2.84 $Y2=0.47
r178 3 42 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.84
+ $Y=0.325 $X2=1.98 $Y2=0.47
r179 2 36 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=0.98
+ $Y=0.325 $X2=1.12 $Y2=0.47
r180 1 30 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.325 $X2=0.26 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_LP__NAND2_8%VGND 1 2 3 4 15 19 23 25 29 32 33 34 35 36
+ 38 55 56 59 62
r101 62 63 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r102 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r103 55 56 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=7.44 $Y=0
+ $X2=7.44 $Y2=0
r104 53 63 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=3.12
+ $Y2=0
r105 52 55 250.524 $w=1.68e-07 $l=3.84e-06 $layer=LI1_cond $X=3.6 $Y=0 $X2=7.44
+ $Y2=0
r106 52 53 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=3.6 $Y=0
+ $X2=3.6 $Y2=0
r107 50 62 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.435 $Y=0 $X2=3.27
+ $Y2=0
r108 50 52 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=3.435 $Y=0 $X2=3.6
+ $Y2=0
r109 49 63 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r110 48 49 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r111 46 49 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r112 46 60 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r113 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r114 43 59 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.855 $Y=0 $X2=0.69
+ $Y2=0
r115 43 45 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.855 $Y=0 $X2=1.2
+ $Y2=0
r116 41 60 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r117 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r118 38 59 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.525 $Y=0 $X2=0.69
+ $Y2=0
r119 38 40 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.525 $Y=0
+ $X2=0.24 $Y2=0
r120 36 56 1.00344 $w=4.9e-07 $l=3.6e-06 $layer=MET1_cond $X=3.84 $Y=0 $X2=7.44
+ $Y2=0
r121 36 53 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.84 $Y=0 $X2=3.6
+ $Y2=0
r122 34 48 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=2.245 $Y=0 $X2=2.16
+ $Y2=0
r123 34 35 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.245 $Y=0 $X2=2.41
+ $Y2=0
r124 32 45 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=1.385 $Y=0 $X2=1.2
+ $Y2=0
r125 32 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.385 $Y=0 $X2=1.55
+ $Y2=0
r126 31 48 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=1.715 $Y=0
+ $X2=2.16 $Y2=0
r127 31 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.715 $Y=0 $X2=1.55
+ $Y2=0
r128 27 62 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.27 $Y=0.085
+ $X2=3.27 $Y2=0
r129 27 29 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=3.27 $Y=0.085
+ $X2=3.27 $Y2=0.45
r130 26 35 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.575 $Y=0 $X2=2.41
+ $Y2=0
r131 25 62 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.105 $Y=0 $X2=3.27
+ $Y2=0
r132 25 26 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=3.105 $Y=0
+ $X2=2.575 $Y2=0
r133 21 35 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.41 $Y=0.085
+ $X2=2.41 $Y2=0
r134 21 23 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=2.41 $Y=0.085
+ $X2=2.41 $Y2=0.45
r135 17 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.55 $Y=0.085
+ $X2=1.55 $Y2=0
r136 17 19 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=1.55 $Y=0.085
+ $X2=1.55 $Y2=0.45
r137 13 59 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=0.085
+ $X2=0.69 $Y2=0
r138 13 15 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=0.69 $Y=0.085
+ $X2=0.69 $Y2=0.47
r139 4 29 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=3.13
+ $Y=0.325 $X2=3.27 $Y2=0.45
r140 3 23 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=2.27
+ $Y=0.325 $X2=2.41 $Y2=0.45
r141 2 19 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=1.41
+ $Y=0.325 $X2=1.55 $Y2=0.45
r142 1 15 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=0.55
+ $Y=0.325 $X2=0.69 $Y2=0.47
.ends

