* File: sky130_fd_sc_lp__invlp_8.pex.spice
* Created: Fri Aug 28 10:40:11 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__INVLP_8%A 3 7 11 15 19 23 27 31 35 39 43 47 51 55 59
+ 63 67 71 75 79 83 87 91 95 99 103 107 111 115 119 123 127 134 135 137 138 139
+ 140 186 187 200
c312 135 0 1.28721e-19 $X=7.25 $Y=1.51
c313 123 0 1.66076e-19 $X=7.155 $Y=0.685
c314 11 0 1.4156e-19 $X=0.925 $Y=0.685
r315 182 183 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=6.725 $Y=1.51
+ $X2=7.155 $Y2=1.51
r316 181 182 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=6.655 $Y=1.51
+ $X2=6.725 $Y2=1.51
r317 180 181 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=6.225 $Y=1.51
+ $X2=6.655 $Y2=1.51
r318 179 180 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=6.155 $Y=1.51
+ $X2=6.225 $Y2=1.51
r319 178 179 62.9501 $w=3.3e-07 $l=3.6e-07 $layer=POLY_cond $X=5.795 $Y=1.51
+ $X2=6.155 $Y2=1.51
r320 177 178 24.4806 $w=3.3e-07 $l=1.4e-07 $layer=POLY_cond $X=5.655 $Y=1.51
+ $X2=5.795 $Y2=1.51
r321 176 177 50.7098 $w=3.3e-07 $l=2.9e-07 $layer=POLY_cond $X=5.365 $Y=1.51
+ $X2=5.655 $Y2=1.51
r322 175 176 24.4806 $w=3.3e-07 $l=1.4e-07 $layer=POLY_cond $X=5.225 $Y=1.51
+ $X2=5.365 $Y2=1.51
r323 174 175 50.7098 $w=3.3e-07 $l=2.9e-07 $layer=POLY_cond $X=4.935 $Y=1.51
+ $X2=5.225 $Y2=1.51
r324 173 174 24.4806 $w=3.3e-07 $l=1.4e-07 $layer=POLY_cond $X=4.795 $Y=1.51
+ $X2=4.935 $Y2=1.51
r325 172 173 50.7098 $w=3.3e-07 $l=2.9e-07 $layer=POLY_cond $X=4.505 $Y=1.51
+ $X2=4.795 $Y2=1.51
r326 171 172 24.4806 $w=3.3e-07 $l=1.4e-07 $layer=POLY_cond $X=4.365 $Y=1.51
+ $X2=4.505 $Y2=1.51
r327 170 171 50.7098 $w=3.3e-07 $l=2.9e-07 $layer=POLY_cond $X=4.075 $Y=1.51
+ $X2=4.365 $Y2=1.51
r328 169 170 24.4806 $w=3.3e-07 $l=1.4e-07 $layer=POLY_cond $X=3.935 $Y=1.51
+ $X2=4.075 $Y2=1.51
r329 168 169 50.7098 $w=3.3e-07 $l=2.9e-07 $layer=POLY_cond $X=3.645 $Y=1.51
+ $X2=3.935 $Y2=1.51
r330 165 166 50.7098 $w=3.3e-07 $l=2.9e-07 $layer=POLY_cond $X=3.215 $Y=1.51
+ $X2=3.505 $Y2=1.51
r331 164 200 2.42108 $w=4.33e-07 $l=6.5e-08 $layer=LI1_cond $X=3.17 $Y=1.562
+ $X2=3.235 $Y2=1.562
r332 163 165 7.86876 $w=3.3e-07 $l=4.5e-08 $layer=POLY_cond $X=3.17 $Y=1.51
+ $X2=3.215 $Y2=1.51
r333 163 164 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.17
+ $Y=1.51 $X2=3.17 $Y2=1.51
r334 161 163 16.6118 $w=3.3e-07 $l=9.5e-08 $layer=POLY_cond $X=3.075 $Y=1.51
+ $X2=3.17 $Y2=1.51
r335 160 161 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=2.645 $Y=1.51
+ $X2=3.075 $Y2=1.51
r336 158 160 27.1035 $w=3.3e-07 $l=1.55e-07 $layer=POLY_cond $X=2.49 $Y=1.51
+ $X2=2.645 $Y2=1.51
r337 158 159 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.49
+ $Y=1.51 $X2=2.49 $Y2=1.51
r338 156 158 48.0869 $w=3.3e-07 $l=2.75e-07 $layer=POLY_cond $X=2.215 $Y=1.51
+ $X2=2.49 $Y2=1.51
r339 155 187 5.45646 $w=4.35e-07 $l=1.9e-07 $layer=LI1_cond $X=1.81 $Y=1.562
+ $X2=2 $Y2=1.562
r340 154 156 70.8188 $w=3.3e-07 $l=4.05e-07 $layer=POLY_cond $X=1.81 $Y=1.51
+ $X2=2.215 $Y2=1.51
r341 154 155 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.81
+ $Y=1.51 $X2=1.81 $Y2=1.51
r342 152 154 4.37153 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=1.785 $Y=1.51
+ $X2=1.81 $Y2=1.51
r343 150 152 55.0813 $w=3.3e-07 $l=3.15e-07 $layer=POLY_cond $X=1.47 $Y=1.51
+ $X2=1.785 $Y2=1.51
r344 150 151 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.47
+ $Y=1.51 $X2=1.47 $Y2=1.51
r345 148 150 20.109 $w=3.3e-07 $l=1.15e-07 $layer=POLY_cond $X=1.355 $Y=1.51
+ $X2=1.47 $Y2=1.51
r346 147 148 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=0.925 $Y=1.51
+ $X2=1.355 $Y2=1.51
r347 145 147 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=0.495 $Y=1.51
+ $X2=0.925 $Y2=1.51
r348 140 164 1.32465 $w=4.33e-07 $l=5e-08 $layer=LI1_cond $X=3.12 $Y=1.562
+ $X2=3.17 $Y2=1.562
r349 140 186 2.70228 $w=4.33e-07 $l=1.02e-07 $layer=LI1_cond $X=3.12 $Y=1.562
+ $X2=3.018 $Y2=1.562
r350 139 186 10.0143 $w=4.33e-07 $l=3.78e-07 $layer=LI1_cond $X=2.64 $Y=1.562
+ $X2=3.018 $Y2=1.562
r351 139 159 3.97394 $w=4.33e-07 $l=1.5e-07 $layer=LI1_cond $X=2.64 $Y=1.562
+ $X2=2.49 $Y2=1.562
r352 138 159 8.74267 $w=4.33e-07 $l=3.3e-07 $layer=LI1_cond $X=2.16 $Y=1.562
+ $X2=2.49 $Y2=1.562
r353 138 187 4.23887 $w=4.33e-07 $l=1.6e-07 $layer=LI1_cond $X=2.16 $Y=1.562
+ $X2=2 $Y2=1.562
r354 137 155 4.01519 $w=3.95e-07 $l=1.3e-07 $layer=LI1_cond $X=1.68 $Y=1.562
+ $X2=1.81 $Y2=1.562
r355 137 151 6.48608 $w=3.95e-07 $l=2.1e-07 $layer=LI1_cond $X=1.68 $Y=1.562
+ $X2=1.47 $Y2=1.562
r356 135 183 16.6118 $w=3.3e-07 $l=9.5e-08 $layer=POLY_cond $X=7.25 $Y=1.51
+ $X2=7.155 $Y2=1.51
r357 134 135 24.2133 $w=1.7e-07 $l=1.02e-06 $layer=licon1_POLY $count=6 $X=7.25
+ $Y=1.51 $X2=7.25 $Y2=1.51
r358 132 168 23.6063 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=3.51 $Y=1.51
+ $X2=3.645 $Y2=1.51
r359 132 166 0.874306 $w=3.3e-07 $l=5e-09 $layer=POLY_cond $X=3.51 $Y=1.51
+ $X2=3.505 $Y2=1.51
r360 131 134 130.61 $w=3.28e-07 $l=3.74e-06 $layer=LI1_cond $X=3.51 $Y=1.51
+ $X2=7.25 $Y2=1.51
r361 131 200 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=3.51 $Y=1.51
+ $X2=3.235 $Y2=1.51
r362 131 132 24.2133 $w=1.7e-07 $l=1.02e-06 $layer=licon1_POLY $count=6 $X=3.51
+ $Y=1.51 $X2=3.51 $Y2=1.51
r363 125 183 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.155 $Y=1.675
+ $X2=7.155 $Y2=1.51
r364 125 127 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=7.155 $Y=1.675
+ $X2=7.155 $Y2=2.465
r365 121 183 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.155 $Y=1.345
+ $X2=7.155 $Y2=1.51
r366 121 123 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=7.155 $Y=1.345
+ $X2=7.155 $Y2=0.685
r367 117 182 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.725 $Y=1.675
+ $X2=6.725 $Y2=1.51
r368 117 119 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=6.725 $Y=1.675
+ $X2=6.725 $Y2=2.465
r369 113 181 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.655 $Y=1.345
+ $X2=6.655 $Y2=1.51
r370 113 115 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.655 $Y=1.345
+ $X2=6.655 $Y2=0.685
r371 109 180 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.225 $Y=1.675
+ $X2=6.225 $Y2=1.51
r372 109 111 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=6.225 $Y=1.675
+ $X2=6.225 $Y2=2.465
r373 105 179 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.155 $Y=1.345
+ $X2=6.155 $Y2=1.51
r374 105 107 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.155 $Y=1.345
+ $X2=6.155 $Y2=0.685
r375 101 178 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.795 $Y=1.675
+ $X2=5.795 $Y2=1.51
r376 101 103 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=5.795 $Y=1.675
+ $X2=5.795 $Y2=2.465
r377 97 177 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.655 $Y=1.345
+ $X2=5.655 $Y2=1.51
r378 97 99 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.655 $Y=1.345
+ $X2=5.655 $Y2=0.685
r379 93 176 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.365 $Y=1.675
+ $X2=5.365 $Y2=1.51
r380 93 95 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=5.365 $Y=1.675
+ $X2=5.365 $Y2=2.465
r381 89 175 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.225 $Y=1.345
+ $X2=5.225 $Y2=1.51
r382 89 91 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=5.225 $Y=1.345
+ $X2=5.225 $Y2=0.685
r383 85 174 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.935 $Y=1.675
+ $X2=4.935 $Y2=1.51
r384 85 87 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=4.935 $Y=1.675
+ $X2=4.935 $Y2=2.465
r385 81 173 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.795 $Y=1.345
+ $X2=4.795 $Y2=1.51
r386 81 83 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.795 $Y=1.345
+ $X2=4.795 $Y2=0.685
r387 77 172 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.505 $Y=1.675
+ $X2=4.505 $Y2=1.51
r388 77 79 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=4.505 $Y=1.675
+ $X2=4.505 $Y2=2.465
r389 73 171 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.365 $Y=1.345
+ $X2=4.365 $Y2=1.51
r390 73 75 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.365 $Y=1.345
+ $X2=4.365 $Y2=0.685
r391 69 170 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.075 $Y=1.675
+ $X2=4.075 $Y2=1.51
r392 69 71 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=4.075 $Y=1.675
+ $X2=4.075 $Y2=2.465
r393 65 169 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.935 $Y=1.345
+ $X2=3.935 $Y2=1.51
r394 65 67 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.935 $Y=1.345
+ $X2=3.935 $Y2=0.685
r395 61 168 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.645 $Y=1.675
+ $X2=3.645 $Y2=1.51
r396 61 63 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.645 $Y=1.675
+ $X2=3.645 $Y2=2.465
r397 57 166 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.505 $Y=1.345
+ $X2=3.505 $Y2=1.51
r398 57 59 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.505 $Y=1.345
+ $X2=3.505 $Y2=0.685
r399 53 165 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.215 $Y=1.675
+ $X2=3.215 $Y2=1.51
r400 53 55 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.215 $Y=1.675
+ $X2=3.215 $Y2=2.465
r401 49 161 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.075 $Y=1.345
+ $X2=3.075 $Y2=1.51
r402 49 51 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.075 $Y=1.345
+ $X2=3.075 $Y2=0.685
r403 45 160 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.645 $Y=1.675
+ $X2=2.645 $Y2=1.51
r404 45 47 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.645 $Y=1.675
+ $X2=2.645 $Y2=2.465
r405 41 160 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.645 $Y=1.345
+ $X2=2.645 $Y2=1.51
r406 41 43 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.645 $Y=1.345
+ $X2=2.645 $Y2=0.685
r407 37 156 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.215 $Y=1.675
+ $X2=2.215 $Y2=1.51
r408 37 39 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.215 $Y=1.675
+ $X2=2.215 $Y2=2.465
r409 33 156 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.215 $Y=1.345
+ $X2=2.215 $Y2=1.51
r410 33 35 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.215 $Y=1.345
+ $X2=2.215 $Y2=0.685
r411 29 152 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.785 $Y=1.675
+ $X2=1.785 $Y2=1.51
r412 29 31 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.785 $Y=1.675
+ $X2=1.785 $Y2=2.465
r413 25 152 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.785 $Y=1.345
+ $X2=1.785 $Y2=1.51
r414 25 27 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.785 $Y=1.345
+ $X2=1.785 $Y2=0.685
r415 21 148 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.355 $Y=1.675
+ $X2=1.355 $Y2=1.51
r416 21 23 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.355 $Y=1.675
+ $X2=1.355 $Y2=2.465
r417 17 148 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.355 $Y=1.345
+ $X2=1.355 $Y2=1.51
r418 17 19 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.355 $Y=1.345
+ $X2=1.355 $Y2=0.685
r419 13 147 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.925 $Y=1.675
+ $X2=0.925 $Y2=1.51
r420 13 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=0.925 $Y=1.675
+ $X2=0.925 $Y2=2.465
r421 9 147 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.925 $Y=1.345
+ $X2=0.925 $Y2=1.51
r422 9 11 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.925 $Y=1.345
+ $X2=0.925 $Y2=0.685
r423 5 145 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=1.675
+ $X2=0.495 $Y2=1.51
r424 5 7 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=0.495 $Y=1.675
+ $X2=0.495 $Y2=2.465
r425 1 145 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=1.345
+ $X2=0.495 $Y2=1.51
r426 1 3 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.495 $Y=1.345
+ $X2=0.495 $Y2=0.685
.ends

.subckt PM_SKY130_FD_SC_LP__INVLP_8%VPWR 1 2 3 4 5 16 18 24 28 32 34 36 41 42 44
+ 45 46 48 60 71 75
r110 74 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r111 71 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r112 68 69 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r113 66 75 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=7.44 $Y2=3.33
r114 65 66 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r115 62 65 250.524 $w=1.68e-07 $l=3.84e-06 $layer=LI1_cond $X=3.12 $Y=3.33
+ $X2=6.96 $Y2=3.33
r116 62 63 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r117 60 74 4.67153 $w=1.7e-07 $l=2.37e-07 $layer=LI1_cond $X=7.205 $Y=3.33
+ $X2=7.442 $Y2=3.33
r118 60 65 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=7.205 $Y=3.33
+ $X2=6.96 $Y2=3.33
r119 59 63 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r120 58 59 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r121 56 59 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r122 56 72 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r123 55 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r124 53 71 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.305 $Y=3.33
+ $X2=1.14 $Y2=3.33
r125 53 55 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.305 $Y=3.33
+ $X2=1.68 $Y2=3.33
r126 52 72 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r127 52 69 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r128 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r129 49 68 4.00981 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=0.365 $Y=3.33
+ $X2=0.182 $Y2=3.33
r130 49 51 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=0.365 $Y=3.33
+ $X2=0.72 $Y2=3.33
r131 48 71 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.975 $Y=3.33
+ $X2=1.14 $Y2=3.33
r132 48 51 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.975 $Y=3.33
+ $X2=0.72 $Y2=3.33
r133 46 66 0.869652 $w=4.9e-07 $l=3.12e-06 $layer=MET1_cond $X=3.84 $Y=3.33
+ $X2=6.96 $Y2=3.33
r134 46 63 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=3.84 $Y=3.33
+ $X2=3.12 $Y2=3.33
r135 44 58 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=2.765 $Y=3.33
+ $X2=2.64 $Y2=3.33
r136 44 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.765 $Y=3.33
+ $X2=2.93 $Y2=3.33
r137 43 62 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=3.095 $Y=3.33
+ $X2=3.12 $Y2=3.33
r138 43 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.095 $Y=3.33
+ $X2=2.93 $Y2=3.33
r139 41 55 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=1.835 $Y=3.33
+ $X2=1.68 $Y2=3.33
r140 41 42 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.835 $Y=3.33
+ $X2=1.96 $Y2=3.33
r141 40 58 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=2.085 $Y=3.33
+ $X2=2.64 $Y2=3.33
r142 40 42 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.085 $Y=3.33
+ $X2=1.96 $Y2=3.33
r143 36 39 32.8272 $w=3.28e-07 $l=9.4e-07 $layer=LI1_cond $X=7.37 $Y=2.01
+ $X2=7.37 $Y2=2.95
r144 34 74 3.09464 $w=3.3e-07 $l=1.15521e-07 $layer=LI1_cond $X=7.37 $Y=3.245
+ $X2=7.442 $Y2=3.33
r145 34 39 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=7.37 $Y=3.245
+ $X2=7.37 $Y2=2.95
r146 30 45 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.93 $Y=3.245
+ $X2=2.93 $Y2=3.33
r147 30 32 13.0959 $w=3.28e-07 $l=3.75e-07 $layer=LI1_cond $X=2.93 $Y=3.245
+ $X2=2.93 $Y2=2.87
r148 26 42 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.96 $Y=3.245
+ $X2=1.96 $Y2=3.33
r149 26 28 17.2866 $w=2.48e-07 $l=3.75e-07 $layer=LI1_cond $X=1.96 $Y=3.245
+ $X2=1.96 $Y2=2.87
r150 22 71 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.14 $Y=3.245
+ $X2=1.14 $Y2=3.33
r151 22 24 13.0959 $w=3.28e-07 $l=3.75e-07 $layer=LI1_cond $X=1.14 $Y=3.245
+ $X2=1.14 $Y2=2.87
r152 18 21 44.7148 $w=2.48e-07 $l=9.7e-07 $layer=LI1_cond $X=0.24 $Y=1.98
+ $X2=0.24 $Y2=2.95
r153 16 68 3.13335 $w=2.5e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.24 $Y=3.245
+ $X2=0.182 $Y2=3.33
r154 16 21 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=0.24 $Y=3.245
+ $X2=0.24 $Y2=2.95
r155 5 39 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=7.23
+ $Y=1.835 $X2=7.37 $Y2=2.95
r156 5 36 400 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_PDIFF $count=1 $X=7.23
+ $Y=1.835 $X2=7.37 $Y2=2.01
r157 4 32 600 $w=1.7e-07 $l=1.13515e-06 $layer=licon1_PDIFF $count=1 $X=2.72
+ $Y=1.835 $X2=2.93 $Y2=2.87
r158 3 28 600 $w=1.7e-07 $l=1.10278e-06 $layer=licon1_PDIFF $count=1 $X=1.86
+ $Y=1.835 $X2=2 $Y2=2.87
r159 2 24 600 $w=1.7e-07 $l=1.10278e-06 $layer=licon1_PDIFF $count=1 $X=1
+ $Y=1.835 $X2=1.14 $Y2=2.87
r160 1 21 400 $w=1.7e-07 $l=1.18528e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.835 $X2=0.28 $Y2=2.95
r161 1 18 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.835 $X2=0.28 $Y2=1.98
.ends

.subckt PM_SKY130_FD_SC_LP__INVLP_8%A_114_367# 1 2 3 4 5 6 7 8 27 31 33 37 41 43
+ 44 45 46 49 51 55 57 61 63 65 67 69 71 73 76 77 78
c114 33 0 1.28721e-19 $X=1.485 $Y=2.375
r115 65 80 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.94 $Y=2.905
+ $X2=6.94 $Y2=2.99
r116 65 67 58.3904 $w=1.68e-07 $l=8.95e-07 $layer=LI1_cond $X=6.94 $Y=2.905
+ $X2=6.94 $Y2=2.01
r117 64 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.175 $Y=2.99
+ $X2=6.01 $Y2=2.99
r118 63 80 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.855 $Y=2.99
+ $X2=6.94 $Y2=2.99
r119 63 64 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=6.855 $Y=2.99
+ $X2=6.175 $Y2=2.99
r120 59 78 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.01 $Y=2.905
+ $X2=6.01 $Y2=2.99
r121 59 61 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=6.01 $Y=2.905
+ $X2=6.01 $Y2=2.27
r122 58 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.315 $Y=2.99
+ $X2=5.15 $Y2=2.99
r123 57 78 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.845 $Y=2.99
+ $X2=6.01 $Y2=2.99
r124 57 58 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=5.845 $Y=2.99
+ $X2=5.315 $Y2=2.99
r125 53 77 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.15 $Y=2.905
+ $X2=5.15 $Y2=2.99
r126 53 55 19.382 $w=3.28e-07 $l=5.55e-07 $layer=LI1_cond $X=5.15 $Y=2.905
+ $X2=5.15 $Y2=2.35
r127 52 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.455 $Y=2.99
+ $X2=4.29 $Y2=2.99
r128 51 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.985 $Y=2.99
+ $X2=5.15 $Y2=2.99
r129 51 52 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=4.985 $Y=2.99
+ $X2=4.455 $Y2=2.99
r130 47 76 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.29 $Y=2.905
+ $X2=4.29 $Y2=2.99
r131 47 49 19.382 $w=3.28e-07 $l=5.55e-07 $layer=LI1_cond $X=4.29 $Y=2.905
+ $X2=4.29 $Y2=2.35
r132 45 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.125 $Y=2.99
+ $X2=4.29 $Y2=2.99
r133 45 46 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=4.125 $Y=2.99
+ $X2=3.595 $Y2=2.99
r134 44 46 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.43 $Y=2.905
+ $X2=3.595 $Y2=2.99
r135 43 75 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.43 $Y=2.46 $X2=3.43
+ $Y2=2.375
r136 43 44 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=3.43 $Y=2.46
+ $X2=3.43 $Y2=2.905
r137 42 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.595 $Y=2.375
+ $X2=2.43 $Y2=2.375
r138 41 75 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.265 $Y=2.375
+ $X2=3.43 $Y2=2.375
r139 41 42 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.265 $Y=2.375
+ $X2=2.595 $Y2=2.375
r140 38 71 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.655 $Y=2.375
+ $X2=1.57 $Y2=2.375
r141 37 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.265 $Y=2.375
+ $X2=2.43 $Y2=2.375
r142 37 38 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=2.265 $Y=2.375
+ $X2=1.655 $Y2=2.375
r143 34 69 2.76166 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.795 $Y=2.375
+ $X2=0.67 $Y2=2.375
r144 33 71 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.485 $Y=2.375
+ $X2=1.57 $Y2=2.375
r145 33 34 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.485 $Y=2.375
+ $X2=0.795 $Y2=2.375
r146 29 69 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.67 $Y=2.46
+ $X2=0.67 $Y2=2.375
r147 29 31 2.30489 $w=2.48e-07 $l=5e-08 $layer=LI1_cond $X=0.67 $Y=2.46 $X2=0.67
+ $Y2=2.51
r148 25 69 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.67 $Y=2.29
+ $X2=0.67 $Y2=2.375
r149 25 27 8.0671 $w=2.48e-07 $l=1.75e-07 $layer=LI1_cond $X=0.67 $Y=2.29
+ $X2=0.67 $Y2=2.115
r150 8 80 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=6.8
+ $Y=1.835 $X2=6.94 $Y2=2.91
r151 8 67 400 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_PDIFF $count=1 $X=6.8
+ $Y=1.835 $X2=6.94 $Y2=2.01
r152 7 61 300 $w=1.7e-07 $l=5.00125e-07 $layer=licon1_PDIFF $count=2 $X=5.87
+ $Y=1.835 $X2=6.01 $Y2=2.27
r153 6 55 300 $w=1.7e-07 $l=5.80797e-07 $layer=licon1_PDIFF $count=2 $X=5.01
+ $Y=1.835 $X2=5.15 $Y2=2.35
r154 5 49 300 $w=1.7e-07 $l=5.80797e-07 $layer=licon1_PDIFF $count=2 $X=4.15
+ $Y=1.835 $X2=4.29 $Y2=2.35
r155 4 75 300 $w=1.7e-07 $l=6.8644e-07 $layer=licon1_PDIFF $count=2 $X=3.29
+ $Y=1.835 $X2=3.43 $Y2=2.455
r156 3 73 300 $w=1.7e-07 $l=6.8644e-07 $layer=licon1_PDIFF $count=2 $X=2.29
+ $Y=1.835 $X2=2.43 $Y2=2.455
r157 2 71 300 $w=1.7e-07 $l=6.8644e-07 $layer=licon1_PDIFF $count=2 $X=1.43
+ $Y=1.835 $X2=1.57 $Y2=2.455
r158 1 31 300 $w=1.7e-07 $l=7.41704e-07 $layer=licon1_PDIFF $count=2 $X=0.57
+ $Y=1.835 $X2=0.71 $Y2=2.51
r159 1 27 600 $w=1.7e-07 $l=3.42929e-07 $layer=licon1_PDIFF $count=1 $X=0.57
+ $Y=1.835 $X2=0.71 $Y2=2.115
.ends

.subckt PM_SKY130_FD_SC_LP__INVLP_8%Y 1 2 3 4 5 6 7 8 26 28 29 30 31 32 35 39 41
+ 43 47 51 53 57 61 63 67 71 72 73 75 76 78 79 81 83 84
c175 67 0 1.66076e-19 $X=6.44 $Y=0.82
r176 71 84 12.276 $w=2.28e-07 $l=2.45e-07 $layer=LI1_cond $X=0.965 $Y=1.665
+ $X2=0.72 $Y2=1.665
r177 71 72 0.280307 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.965 $Y=1.665
+ $X2=1.05 $Y2=1.665
r178 65 67 6.46067 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=6.44 $Y=1.005
+ $X2=6.44 $Y2=0.82
r179 64 81 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.665 $Y=1.93
+ $X2=5.58 $Y2=1.93
r180 63 83 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.345 $Y=1.93
+ $X2=6.51 $Y2=1.93
r181 63 64 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=6.345 $Y=1.93
+ $X2=5.665 $Y2=1.93
r182 62 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.605 $Y=1.09
+ $X2=5.44 $Y2=1.09
r183 61 65 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.275 $Y=1.09
+ $X2=6.44 $Y2=1.005
r184 61 62 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=6.275 $Y=1.09
+ $X2=5.605 $Y2=1.09
r185 55 79 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.44 $Y=1.005
+ $X2=5.44 $Y2=1.09
r186 55 57 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=5.44 $Y=1.005
+ $X2=5.44 $Y2=0.86
r187 54 78 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.805 $Y=1.93
+ $X2=4.72 $Y2=1.93
r188 53 81 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.495 $Y=1.93
+ $X2=5.58 $Y2=1.93
r189 53 54 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=5.495 $Y=1.93
+ $X2=4.805 $Y2=1.93
r190 52 76 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.745 $Y=1.09
+ $X2=4.62 $Y2=1.09
r191 51 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.275 $Y=1.09
+ $X2=5.44 $Y2=1.09
r192 51 52 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=5.275 $Y=1.09
+ $X2=4.745 $Y2=1.09
r193 45 76 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.62 $Y=1.005
+ $X2=4.62 $Y2=1.09
r194 45 47 6.68417 $w=2.48e-07 $l=1.45e-07 $layer=LI1_cond $X=4.62 $Y=1.005
+ $X2=4.62 $Y2=0.86
r195 44 75 5.16603 $w=1.7e-07 $l=1.07912e-07 $layer=LI1_cond $X=3.945 $Y=1.93
+ $X2=3.86 $Y2=1.982
r196 43 78 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.635 $Y=1.93
+ $X2=4.72 $Y2=1.93
r197 43 44 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=4.635 $Y=1.93
+ $X2=3.945 $Y2=1.93
r198 42 73 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.805 $Y=1.09
+ $X2=3.68 $Y2=1.09
r199 41 76 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.495 $Y=1.09
+ $X2=4.62 $Y2=1.09
r200 41 42 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=4.495 $Y=1.09
+ $X2=3.805 $Y2=1.09
r201 37 75 1.34256 $w=1.7e-07 $l=1.38e-07 $layer=LI1_cond $X=3.86 $Y=2.12
+ $X2=3.86 $Y2=1.982
r202 37 39 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=3.86 $Y=2.12
+ $X2=3.86 $Y2=2.57
r203 33 73 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.68 $Y=1.005
+ $X2=3.68 $Y2=1.09
r204 33 35 6.68417 $w=2.48e-07 $l=1.45e-07 $layer=LI1_cond $X=3.68 $Y=1.005
+ $X2=3.68 $Y2=0.86
r205 31 75 5.16603 $w=1.7e-07 $l=1.08305e-07 $layer=LI1_cond $X=3.775 $Y=2.035
+ $X2=3.86 $Y2=1.982
r206 31 32 172.235 $w=1.68e-07 $l=2.64e-06 $layer=LI1_cond $X=3.775 $Y=2.035
+ $X2=1.135 $Y2=2.035
r207 29 73 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.555 $Y=1.09
+ $X2=3.68 $Y2=1.09
r208 29 30 157.882 $w=1.68e-07 $l=2.42e-06 $layer=LI1_cond $X=3.555 $Y=1.09
+ $X2=1.135 $Y2=1.09
r209 28 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.05 $Y=1.95
+ $X2=1.135 $Y2=2.035
r210 27 72 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=1.05 $Y=1.78
+ $X2=1.05 $Y2=1.665
r211 27 28 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.05 $Y=1.78
+ $X2=1.05 $Y2=1.95
r212 26 72 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=1.05 $Y=1.55
+ $X2=1.05 $Y2=1.665
r213 25 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.05 $Y=1.175
+ $X2=1.135 $Y2=1.09
r214 25 26 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.05 $Y=1.175
+ $X2=1.05 $Y2=1.55
r215 8 83 300 $w=1.7e-07 $l=2.84341e-07 $layer=licon1_PDIFF $count=2 $X=6.3
+ $Y=1.835 $X2=6.51 $Y2=2.01
r216 7 81 300 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_PDIFF $count=2 $X=5.44
+ $Y=1.835 $X2=5.58 $Y2=2.01
r217 6 78 300 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_PDIFF $count=2 $X=4.58
+ $Y=1.835 $X2=4.72 $Y2=2.01
r218 5 75 600 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_PDIFF $count=1 $X=3.72
+ $Y=1.835 $X2=3.86 $Y2=2.01
r219 5 39 600 $w=1.7e-07 $l=8.01951e-07 $layer=licon1_PDIFF $count=1 $X=3.72
+ $Y=1.835 $X2=3.86 $Y2=2.57
r220 4 67 182 $w=1.7e-07 $l=6.51594e-07 $layer=licon1_NDIFF $count=1 $X=6.23
+ $Y=0.265 $X2=6.44 $Y2=0.82
r221 3 57 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=5.3
+ $Y=0.265 $X2=5.44 $Y2=0.86
r222 2 47 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=4.44
+ $Y=0.265 $X2=4.58 $Y2=0.86
r223 1 35 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=3.58
+ $Y=0.265 $X2=3.72 $Y2=0.86
.ends

.subckt PM_SKY130_FD_SC_LP__INVLP_8%VGND 1 2 3 4 5 16 18 22 26 30 32 34 37 38 40
+ 41 42 44 56 67 71
r115 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r116 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r117 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r118 62 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0 $X2=7.44
+ $Y2=0
r119 61 62 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=6.96 $Y=0
+ $X2=6.96 $Y2=0
r120 58 61 250.524 $w=1.68e-07 $l=3.84e-06 $layer=LI1_cond $X=3.12 $Y=0 $X2=6.96
+ $Y2=0
r121 58 59 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=3.12 $Y=0
+ $X2=3.12 $Y2=0
r122 56 70 3.97515 $w=1.7e-07 $l=1.97e-07 $layer=LI1_cond $X=7.285 $Y=0
+ $X2=7.482 $Y2=0
r123 56 61 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=7.285 $Y=0
+ $X2=6.96 $Y2=0
r124 55 59 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r125 54 55 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r126 52 55 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r127 52 68 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r128 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r129 49 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.305 $Y=0 $X2=1.14
+ $Y2=0
r130 49 51 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.305 $Y=0
+ $X2=1.68 $Y2=0
r131 48 68 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r132 48 65 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r133 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r134 45 64 4.00981 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=0.365 $Y=0
+ $X2=0.182 $Y2=0
r135 45 47 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=0.365 $Y=0
+ $X2=0.72 $Y2=0
r136 44 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.975 $Y=0 $X2=1.14
+ $Y2=0
r137 44 47 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.975 $Y=0
+ $X2=0.72 $Y2=0
r138 42 62 0.869652 $w=4.9e-07 $l=3.12e-06 $layer=MET1_cond $X=3.84 $Y=0
+ $X2=6.96 $Y2=0
r139 42 59 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=3.84 $Y=0 $X2=3.12
+ $Y2=0
r140 40 54 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=2.695 $Y=0 $X2=2.64
+ $Y2=0
r141 40 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.695 $Y=0 $X2=2.86
+ $Y2=0
r142 39 58 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=3.025 $Y=0 $X2=3.12
+ $Y2=0
r143 39 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.025 $Y=0 $X2=2.86
+ $Y2=0
r144 37 51 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=1.835 $Y=0
+ $X2=1.68 $Y2=0
r145 37 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.835 $Y=0 $X2=2
+ $Y2=0
r146 36 54 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=2.165 $Y=0
+ $X2=2.64 $Y2=0
r147 36 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.165 $Y=0 $X2=2
+ $Y2=0
r148 32 70 3.16801 $w=2.5e-07 $l=1.15521e-07 $layer=LI1_cond $X=7.41 $Y=0.085
+ $X2=7.482 $Y2=0
r149 32 34 14.9818 $w=2.48e-07 $l=3.25e-07 $layer=LI1_cond $X=7.41 $Y=0.085
+ $X2=7.41 $Y2=0.41
r150 28 41 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.86 $Y=0.085
+ $X2=2.86 $Y2=0
r151 28 30 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=2.86 $Y=0.085
+ $X2=2.86 $Y2=0.41
r152 24 38 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2 $Y=0.085 $X2=2
+ $Y2=0
r153 24 26 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=2 $Y=0.085 $X2=2
+ $Y2=0.41
r154 20 67 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.14 $Y=0.085
+ $X2=1.14 $Y2=0
r155 20 22 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=1.14 $Y=0.085
+ $X2=1.14 $Y2=0.41
r156 16 64 3.13335 $w=2.5e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.24 $Y=0.085
+ $X2=0.182 $Y2=0
r157 16 18 14.9818 $w=2.48e-07 $l=3.25e-07 $layer=LI1_cond $X=0.24 $Y=0.085
+ $X2=0.24 $Y2=0.41
r158 5 34 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=7.23
+ $Y=0.265 $X2=7.37 $Y2=0.41
r159 4 30 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=2.72
+ $Y=0.265 $X2=2.86 $Y2=0.41
r160 3 26 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=1.86
+ $Y=0.265 $X2=2 $Y2=0.41
r161 2 22 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=1
+ $Y=0.265 $X2=1.14 $Y2=0.41
r162 1 18 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.265 $X2=0.28 $Y2=0.41
.ends

.subckt PM_SKY130_FD_SC_LP__INVLP_8%A_114_53# 1 2 3 4 5 6 7 8 27 31 33 37 39 43
+ 45 51 52 55 57 61 63 67 71 72 73 74 75 77 79
c131 31 0 1.4156e-19 $X=0.71 $Y=0.96
r132 68 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.105 $Y=0.34
+ $X2=5.94 $Y2=0.34
r133 67 79 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.775 $Y=0.34
+ $X2=6.94 $Y2=0.34
r134 67 68 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=6.775 $Y=0.34
+ $X2=6.105 $Y2=0.34
r135 64 75 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.095 $Y=0.34
+ $X2=5.01 $Y2=0.34
r136 63 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.775 $Y=0.34
+ $X2=5.94 $Y2=0.34
r137 63 64 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=5.775 $Y=0.34
+ $X2=5.095 $Y2=0.34
r138 59 75 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.01 $Y=0.425
+ $X2=5.01 $Y2=0.34
r139 59 61 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=5.01 $Y=0.425
+ $X2=5.01 $Y2=0.545
r140 58 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.315 $Y=0.34
+ $X2=4.15 $Y2=0.34
r141 57 75 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.925 $Y=0.34
+ $X2=5.01 $Y2=0.34
r142 57 58 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=4.925 $Y=0.34
+ $X2=4.315 $Y2=0.34
r143 53 74 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.15 $Y=0.425
+ $X2=4.15 $Y2=0.34
r144 53 55 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=4.15 $Y=0.425
+ $X2=4.15 $Y2=0.545
r145 51 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.985 $Y=0.34
+ $X2=4.15 $Y2=0.34
r146 51 52 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=3.985 $Y=0.34
+ $X2=3.375 $Y2=0.34
r147 48 50 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=3.29 $Y=0.665
+ $X2=3.29 $Y2=0.545
r148 47 52 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.29 $Y=0.425
+ $X2=3.375 $Y2=0.34
r149 47 50 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=3.29 $Y=0.425
+ $X2=3.29 $Y2=0.545
r150 46 73 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.515 $Y=0.75
+ $X2=2.43 $Y2=0.75
r151 45 48 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.205 $Y=0.75
+ $X2=3.29 $Y2=0.665
r152 45 46 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.205 $Y=0.75
+ $X2=2.515 $Y2=0.75
r153 41 73 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.43 $Y=0.665
+ $X2=2.43 $Y2=0.75
r154 41 43 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=2.43 $Y=0.665
+ $X2=2.43 $Y2=0.545
r155 40 72 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.655 $Y=0.75
+ $X2=1.57 $Y2=0.75
r156 39 73 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.345 $Y=0.75
+ $X2=2.43 $Y2=0.75
r157 39 40 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.345 $Y=0.75
+ $X2=1.655 $Y2=0.75
r158 35 72 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.57 $Y=0.665
+ $X2=1.57 $Y2=0.75
r159 35 37 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=1.57 $Y=0.665
+ $X2=1.57 $Y2=0.545
r160 34 71 2.76166 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.795 $Y=0.75
+ $X2=0.67 $Y2=0.75
r161 33 72 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.485 $Y=0.75
+ $X2=1.57 $Y2=0.75
r162 33 34 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.485 $Y=0.75
+ $X2=0.795 $Y2=0.75
r163 29 71 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.67 $Y=0.835
+ $X2=0.67 $Y2=0.75
r164 29 31 5.76222 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=0.67 $Y=0.835
+ $X2=0.67 $Y2=0.96
r165 25 71 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.67 $Y=0.665
+ $X2=0.67 $Y2=0.75
r166 25 27 11.2939 $w=2.48e-07 $l=2.45e-07 $layer=LI1_cond $X=0.67 $Y=0.665
+ $X2=0.67 $Y2=0.42
r167 8 79 91 $w=1.7e-07 $l=2.76857e-07 $layer=licon1_NDIFF $count=2 $X=6.73
+ $Y=0.265 $X2=6.94 $Y2=0.42
r168 7 77 91 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=2 $X=5.73
+ $Y=0.265 $X2=5.94 $Y2=0.41
r169 6 61 182 $w=1.7e-07 $l=3.42929e-07 $layer=licon1_NDIFF $count=1 $X=4.87
+ $Y=0.265 $X2=5.01 $Y2=0.545
r170 5 55 182 $w=1.7e-07 $l=3.42929e-07 $layer=licon1_NDIFF $count=1 $X=4.01
+ $Y=0.265 $X2=4.15 $Y2=0.545
r171 4 50 182 $w=1.7e-07 $l=3.42929e-07 $layer=licon1_NDIFF $count=1 $X=3.15
+ $Y=0.265 $X2=3.29 $Y2=0.545
r172 3 43 182 $w=1.7e-07 $l=3.42929e-07 $layer=licon1_NDIFF $count=1 $X=2.29
+ $Y=0.265 $X2=2.43 $Y2=0.545
r173 2 37 182 $w=1.7e-07 $l=3.42929e-07 $layer=licon1_NDIFF $count=1 $X=1.43
+ $Y=0.265 $X2=1.57 $Y2=0.545
r174 1 31 182 $w=1.7e-07 $l=7.61791e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.265 $X2=0.71 $Y2=0.96
r175 1 27 182 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.265 $X2=0.71 $Y2=0.42
.ends

