* File: sky130_fd_sc_lp__and4b_1.spice
* Created: Wed Sep  2 09:33:27 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__and4b_1.pex.spice"
.subckt sky130_fd_sc_lp__and4b_1  VNB VPB A_N B C D VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* D	D
* C	C
* B	B
* A_N	A_N
* VPB	VPB
* VNB	VNB
MM1005 N_VGND_M1005_d N_A_N_M1005_g N_A_27_49#_M1005_s VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.1113 PD=1.37 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1001 A_300_47# N_A_27_49#_M1001_g N_A_215_367#_M1001_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.1113 PD=0.63 PS=1.37 NRD=14.28 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75002.1 A=0.063 P=1.14 MULT=1
MM1003 A_372_47# N_B_M1003_g A_300_47# VNB NSHORT L=0.15 W=0.42 AD=0.0441
+ AS=0.0441 PD=0.63 PS=0.63 NRD=14.28 NRS=14.28 M=1 R=2.8 SA=75000.6 SB=75001.7
+ A=0.063 P=1.14 MULT=1
MM1004 A_444_47# N_C_M1004_g A_372_47# VNB NSHORT L=0.15 W=0.42 AD=0.0441
+ AS=0.0441 PD=0.63 PS=0.63 NRD=14.28 NRS=14.28 M=1 R=2.8 SA=75000.9 SB=75001.4
+ A=0.063 P=1.14 MULT=1
MM1011 N_VGND_M1011_d N_D_M1011_g A_444_47# VNB NSHORT L=0.15 W=0.42 AD=0.1288
+ AS=0.0441 PD=0.996667 PS=0.63 NRD=71.904 NRS=14.28 M=1 R=2.8 SA=75001.3
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1006 N_X_M1006_d N_A_215_367#_M1006_g N_VGND_M1011_d VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.2576 PD=2.21 PS=1.99333 NRD=0 NRS=0 M=1 R=5.6 SA=75001.1
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1010 N_VPWR_M1010_d N_A_N_M1010_g N_A_27_49#_M1010_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0672 AS=0.1113 PD=0.74 PS=1.37 NRD=9.3772 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75003 A=0.063 P=1.14 MULT=1
MM1008 N_A_215_367#_M1008_d N_A_27_49#_M1008_g N_VPWR_M1010_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0588 AS=0.0672 PD=0.7 PS=0.74 NRD=0 NRS=9.3772 M=1 R=2.8
+ SA=75000.7 SB=75002.5 A=0.063 P=1.14 MULT=1
MM1002 N_VPWR_M1002_d N_B_M1002_g N_A_215_367#_M1008_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.1659 AS=0.0588 PD=1.21 PS=0.7 NRD=49.25 NRS=0 M=1 R=2.8 SA=75001.1
+ SB=75002.1 A=0.063 P=1.14 MULT=1
MM1009 N_A_215_367#_M1009_d N_C_M1009_g N_VPWR_M1002_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0588 AS=0.1659 PD=0.7 PS=1.21 NRD=0 NRS=0 M=1 R=2.8 SA=75002 SB=75001.1
+ A=0.063 P=1.14 MULT=1
MM1007 N_VPWR_M1007_d N_D_M1007_g N_A_215_367#_M1009_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.095025 AS=0.0588 PD=0.8175 PS=0.7 NRD=23.443 NRS=0 M=1 R=2.8 SA=75002.5
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1000 N_X_M1000_d N_A_215_367#_M1000_g N_VPWR_M1007_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.285075 PD=3.05 PS=2.4525 NRD=0 NRS=2.3443 M=1 R=8.4 SA=75001.1
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX12_noxref VNB VPB NWDIODE A=7.8703 P=12.17
*
.include "sky130_fd_sc_lp__and4b_1.pxi.spice"
*
.ends
*
*
