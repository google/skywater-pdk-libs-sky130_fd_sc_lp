* File: sky130_fd_sc_lp__dfxtp_2.spice
* Created: Fri Aug 28 10:24:21 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__dfxtp_2.pex.spice"
.subckt sky130_fd_sc_lp__dfxtp_2  VNB VPB CLK D VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* D	D
* CLK	CLK
* VPB	VPB
* VNB	VNB
MM1023 N_A_110_62#_M1023_d N_CLK_M1023_g N_VGND_M1023_s VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.1113 PD=1.37 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1009 N_VGND_M1009_d N_A_110_62#_M1009_g N_A_240_443#_M1009_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0588 AS=0.1197 PD=0.7 PS=1.41 NRD=0 NRS=5.712 M=1 R=2.8 SA=75000.2
+ SB=75005.2 A=0.063 P=1.14 MULT=1
MM1012 N_A_432_119#_M1012_d N_D_M1012_g N_VGND_M1009_d VNB NSHORT L=0.15 W=0.42
+ AD=0.09345 AS=0.0588 PD=0.865 PS=0.7 NRD=25.704 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75004.7 A=0.063 P=1.14 MULT=1
MM1015 N_A_551_119#_M1015_d N_A_110_62#_M1015_g N_A_432_119#_M1012_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.0588 AS=0.09345 PD=0.7 PS=0.865 NRD=0 NRS=21.42 M=1 R=2.8
+ SA=75001.2 SB=75004.1 A=0.063 P=1.14 MULT=1
MM1004 A_637_119# N_A_240_443#_M1004_g N_A_551_119#_M1015_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75001.7
+ SB=75003.7 A=0.063 P=1.14 MULT=1
MM1024 N_VGND_M1024_d N_A_679_93#_M1024_g A_637_119# VNB NSHORT L=0.15 W=0.42
+ AD=0.170457 AS=0.0441 PD=1.20057 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75002
+ SB=75003.4 A=0.063 P=1.14 MULT=1
MM1000 N_A_679_93#_M1000_d N_A_551_119#_M1000_g N_VGND_M1024_d VNB NSHORT L=0.15
+ W=0.64 AD=0.130294 AS=0.259743 PD=1.22566 PS=1.82943 NRD=0 NRS=3.744 M=1
+ R=4.26667 SA=75002.1 SB=75001.6 A=0.096 P=1.58 MULT=1
MM1018 N_A_1004_379#_M1018_d N_A_240_443#_M1018_g N_A_679_93#_M1000_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.0882 AS=0.0855057 PD=0.84 PS=0.80434 NRD=21.42 NRS=27.852
+ M=1 R=2.8 SA=75003.6 SB=75001.8 A=0.063 P=1.14 MULT=1
MM1006 A_1133_119# N_A_110_62#_M1006_g N_A_1004_379#_M1018_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.0882 PD=0.63 PS=0.84 NRD=14.28 NRS=18.564 M=1 R=2.8
+ SA=75004.1 SB=75001.2 A=0.063 P=1.14 MULT=1
MM1001 N_VGND_M1001_d N_A_1175_93#_M1001_g A_1133_119# VNB NSHORT L=0.15 W=0.42
+ AD=0.121681 AS=0.0441 PD=0.935094 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75004.5
+ SB=75000.9 A=0.063 P=1.14 MULT=1
MM1003 N_A_1175_93#_M1003_d N_A_1004_379#_M1003_g N_VGND_M1001_d VNB NSHORT
+ L=0.15 W=0.64 AD=0.1696 AS=0.185419 PD=1.81 PS=1.42491 NRD=0 NRS=24.372 M=1
+ R=4.26667 SA=75003.5 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1016 N_Q_M1016_d N_A_1175_93#_M1016_g N_VGND_M1016_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1025 N_Q_M1016_d N_A_1175_93#_M1025_g N_VGND_M1025_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1021 N_A_110_62#_M1021_d N_CLK_M1021_g N_VPWR_M1021_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1696 AS=0.1696 PD=1.81 PS=1.81 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1013 N_VPWR_M1013_d N_A_110_62#_M1013_g N_A_240_443#_M1013_s VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.197615 AS=0.1696 PD=1.53358 PS=1.81 NRD=0 NRS=0 M=1
+ R=4.26667 SA=75000.2 SB=75002.8 A=0.096 P=1.58 MULT=1
MM1010 N_A_432_119#_M1010_d N_D_M1010_g N_VPWR_M1013_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0588 AS=0.129685 PD=0.7 PS=1.00642 NRD=0 NRS=164.16 M=1 R=2.8 SA=75001
+ SB=75003.4 A=0.063 P=1.14 MULT=1
MM1022 N_A_551_119#_M1022_d N_A_240_443#_M1022_g N_A_432_119#_M1010_d VPB
+ PHIGHVT L=0.15 W=0.42 AD=0.1155 AS=0.0588 PD=0.97 PS=0.7 NRD=126.632 NRS=0 M=1
+ R=2.8 SA=75001.4 SB=75003 A=0.063 P=1.14 MULT=1
MM1002 A_705_443# N_A_110_62#_M1002_g N_A_551_119#_M1022_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0441 AS=0.1155 PD=0.63 PS=0.97 NRD=23.443 NRS=0 M=1 R=2.8
+ SA=75002.1 SB=75002.3 A=0.063 P=1.14 MULT=1
MM1005 N_VPWR_M1005_d N_A_679_93#_M1005_g A_705_443# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.128233 AS=0.0441 PD=0.95 PS=0.63 NRD=117.392 NRS=23.443 M=1 R=2.8
+ SA=75002.5 SB=75001.9 A=0.063 P=1.14 MULT=1
MM1011 N_A_679_93#_M1011_d N_A_551_119#_M1011_g N_VPWR_M1005_d VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.1512 AS=0.256467 PD=1.2 PS=1.9 NRD=0 NRS=19.9167 M=1 R=5.6
+ SA=75001.7 SB=75001.7 A=0.126 P=1.98 MULT=1
MM1014 N_A_1004_379#_M1014_d N_A_110_62#_M1014_g N_A_679_93#_M1011_d VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.3304 AS=0.1512 PD=1.98 PS=1.2 NRD=63.3158 NRS=18.7544 M=1
+ R=5.6 SA=75002.2 SB=75001.2 A=0.126 P=1.98 MULT=1
MM1017 A_1163_379# N_A_240_443#_M1017_g N_A_1004_379#_M1014_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0441 AS=0.1652 PD=0.63 PS=0.99 NRD=23.443 NRS=44.5417 M=1 R=2.8
+ SA=75002.3 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1020 N_VPWR_M1020_d N_A_1175_93#_M1020_g A_1163_379# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0917 AS=0.0441 PD=0.82 PS=0.63 NRD=0 NRS=23.443 M=1 R=2.8 SA=75002.6
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1007 N_A_1175_93#_M1007_d N_A_1004_379#_M1007_g N_VPWR_M1020_d VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.2226 AS=0.1834 PD=2.21 PS=1.64 NRD=0 NRS=12.8838 M=1 R=5.6
+ SA=75001.7 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1008 N_Q_M1008_d N_A_1175_93#_M1008_g N_VPWR_M1008_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1019 N_Q_M1008_d N_A_1175_93#_M1019_g N_VPWR_M1019_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX26_noxref VNB VPB NWDIODE A=16.8223 P=21.77
*
.include "sky130_fd_sc_lp__dfxtp_2.pxi.spice"
*
.ends
*
*
