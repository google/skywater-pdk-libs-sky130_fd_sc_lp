* File: sky130_fd_sc_lp__a31oi_0.pxi.spice
* Created: Wed Sep  2 09:26:50 2020
* 
x_PM_SKY130_FD_SC_LP__A31OI_0%A3 N_A3_c_55_n N_A3_M1005_g N_A3_c_56_n
+ N_A3_M1002_g N_A3_c_57_n N_A3_c_58_n N_A3_c_63_n A3 A3 A3 N_A3_c_60_n
+ PM_SKY130_FD_SC_LP__A31OI_0%A3
x_PM_SKY130_FD_SC_LP__A31OI_0%A2 N_A2_M1001_g N_A2_M1007_g N_A2_c_97_n
+ N_A2_c_101_n A2 A2 A2 A2 N_A2_c_99_n PM_SKY130_FD_SC_LP__A31OI_0%A2
x_PM_SKY130_FD_SC_LP__A31OI_0%A1 N_A1_M1000_g N_A1_M1006_g N_A1_c_140_n
+ N_A1_c_141_n A1 A1 A1 N_A1_c_143_n PM_SKY130_FD_SC_LP__A31OI_0%A1
x_PM_SKY130_FD_SC_LP__A31OI_0%B1 N_B1_c_178_n N_B1_M1004_g N_B1_M1003_g B1 B1 B1
+ PM_SKY130_FD_SC_LP__A31OI_0%B1
x_PM_SKY130_FD_SC_LP__A31OI_0%VPWR N_VPWR_M1005_s N_VPWR_M1001_d N_VPWR_c_209_n
+ N_VPWR_c_210_n N_VPWR_c_211_n N_VPWR_c_212_n N_VPWR_c_213_n VPWR
+ N_VPWR_c_214_n N_VPWR_c_208_n PM_SKY130_FD_SC_LP__A31OI_0%VPWR
x_PM_SKY130_FD_SC_LP__A31OI_0%A_110_473# N_A_110_473#_M1005_d
+ N_A_110_473#_M1006_d N_A_110_473#_c_256_n N_A_110_473#_c_257_n
+ N_A_110_473#_c_258_n N_A_110_473#_c_259_n
+ PM_SKY130_FD_SC_LP__A31OI_0%A_110_473#
x_PM_SKY130_FD_SC_LP__A31OI_0%Y N_Y_M1000_d N_Y_M1004_d N_Y_c_282_n Y Y Y
+ N_Y_c_278_n PM_SKY130_FD_SC_LP__A31OI_0%Y
x_PM_SKY130_FD_SC_LP__A31OI_0%VGND N_VGND_M1002_s N_VGND_M1003_d N_VGND_c_310_n
+ N_VGND_c_311_n N_VGND_c_312_n N_VGND_c_313_n VGND N_VGND_c_314_n
+ N_VGND_c_315_n PM_SKY130_FD_SC_LP__A31OI_0%VGND
cc_1 VNB N_A3_c_55_n 0.00162933f $X=-0.19 $Y=-0.245 $X2=0.36 $Y2=2.065
cc_2 VNB N_A3_c_56_n 0.0219034f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=0.765
cc_3 VNB N_A3_c_57_n 0.0256434f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.46
cc_4 VNB N_A3_c_58_n 0.0175475f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.625
cc_5 VNB A3 0.0418827f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_6 VNB N_A3_c_60_n 0.0478306f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.12
cc_7 VNB N_A2_M1007_g 0.0343172f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=0.765
cc_8 VNB N_A2_c_97_n 0.0215832f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB A2 0.00694218f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.46
cc_10 VNB N_A2_c_99_n 0.0157583f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A1_M1000_g 0.0210765f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.215
cc_12 VNB N_A1_M1006_g 0.00661765f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=0.765
cc_13 VNB N_A1_c_140_n 0.0217578f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A1_c_141_n 0.0176281f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=0.765
cc_15 VNB A1 0.0103209f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.46
cc_16 VNB N_A1_c_143_n 0.0156416f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_17 VNB N_B1_c_178_n 0.0810186f $X=-0.19 $Y=-0.245 $X2=0.36 $Y2=1.625
cc_18 VNB N_B1_M1003_g 0.034558f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=0.765
cc_19 VNB B1 0.0340273f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=0.445
cc_20 VNB N_VPWR_c_208_n 0.103974f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.12
cc_21 VNB N_Y_c_278_n 0.00654561f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_VGND_c_310_n 0.0123757f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=0.765
cc_23 VNB N_VGND_c_311_n 0.0202617f $X=-0.19 $Y=-0.245 $X2=0.54 $Y2=0.445
cc_24 VNB N_VGND_c_312_n 0.0109108f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_313_n 0.0201869f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.46
cc_26 VNB N_VGND_c_314_n 0.04322f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.14
cc_27 VNB N_VGND_c_315_n 0.147359f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VPB N_A3_c_55_n 0.0286204f $X=-0.19 $Y=1.655 $X2=0.36 $Y2=2.065
cc_29 VPB N_A3_M1005_g 0.0211175f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.685
cc_30 VPB N_A3_c_63_n 0.01763f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.14
cc_31 VPB A3 0.00956296f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_32 VPB N_A2_M1001_g 0.0389159f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.215
cc_33 VPB N_A2_c_101_n 0.0157952f $X=-0.19 $Y=1.655 $X2=0.54 $Y2=0.765
cc_34 VPB A2 0.00297825f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.46
cc_35 VPB N_A1_M1006_g 0.0473477f $X=-0.19 $Y=1.655 $X2=0.54 $Y2=0.765
cc_36 VPB A1 0.00565184f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.46
cc_37 VPB N_B1_c_178_n 0.024845f $X=-0.19 $Y=1.655 $X2=0.36 $Y2=1.625
cc_38 VPB N_B1_M1004_g 0.0408039f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.215
cc_39 VPB B1 0.00812737f $X=-0.19 $Y=1.655 $X2=0.54 $Y2=0.445
cc_40 VPB N_VPWR_c_209_n 0.0108797f $X=-0.19 $Y=1.655 $X2=0.54 $Y2=0.445
cc_41 VPB N_VPWR_c_210_n 0.0430706f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.12
cc_42 VPB N_VPWR_c_211_n 0.0182558f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_43 VPB N_VPWR_c_212_n 0.00832033f $X=-0.19 $Y=1.655 $X2=0.54 $Y2=0.765
cc_44 VPB N_VPWR_c_213_n 0.00407598f $X=-0.19 $Y=1.655 $X2=0.36 $Y2=2.14
cc_45 VPB N_VPWR_c_214_n 0.0513432f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_46 VPB N_VPWR_c_208_n 0.0542428f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.12
cc_47 VPB N_A_110_473#_c_256_n 0.00257792f $X=-0.19 $Y=1.655 $X2=0.54 $Y2=0.445
cc_48 VPB N_A_110_473#_c_257_n 0.00484332f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_49 VPB N_A_110_473#_c_258_n 0.0025304f $X=-0.19 $Y=1.655 $X2=0.54 $Y2=0.765
cc_50 VPB N_A_110_473#_c_259_n 0.0085294f $X=-0.19 $Y=1.655 $X2=0.36 $Y2=2.14
cc_51 VPB Y 0.018475f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.625
cc_52 VPB Y 0.0459526f $X=-0.19 $Y=1.655 $X2=0.36 $Y2=2.14
cc_53 VPB N_Y_c_278_n 0.00403722f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_54 N_A3_c_55_n N_A2_M1001_g 0.00827396f $X=0.36 $Y=2.065 $X2=0 $Y2=0
cc_55 N_A3_c_63_n N_A2_M1001_g 0.0184544f $X=0.475 $Y=2.14 $X2=0 $Y2=0
cc_56 N_A3_c_56_n N_A2_M1007_g 0.0422071f $X=0.54 $Y=0.765 $X2=0 $Y2=0
cc_57 A3 N_A2_M1007_g 6.68743e-19 $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_58 N_A3_c_60_n N_A2_M1007_g 0.00615564f $X=0.27 $Y=1.12 $X2=0 $Y2=0
cc_59 N_A3_c_58_n N_A2_c_97_n 0.0122248f $X=0.27 $Y=1.625 $X2=0 $Y2=0
cc_60 N_A3_c_55_n N_A2_c_101_n 0.0122248f $X=0.36 $Y=2.065 $X2=0 $Y2=0
cc_61 N_A3_c_56_n A2 0.00532347f $X=0.54 $Y=0.765 $X2=0 $Y2=0
cc_62 A3 A2 0.0873333f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_63 N_A3_c_60_n A2 0.00299087f $X=0.27 $Y=1.12 $X2=0 $Y2=0
cc_64 N_A3_c_57_n N_A2_c_99_n 0.0122248f $X=0.27 $Y=1.46 $X2=0 $Y2=0
cc_65 A3 N_A2_c_99_n 0.00203596f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_66 N_A3_M1005_g N_VPWR_c_210_n 0.00831873f $X=0.475 $Y=2.685 $X2=0 $Y2=0
cc_67 N_A3_c_63_n N_VPWR_c_210_n 0.00483136f $X=0.475 $Y=2.14 $X2=0 $Y2=0
cc_68 N_A3_c_55_n N_VPWR_c_211_n 0.00192287f $X=0.36 $Y=2.065 $X2=0 $Y2=0
cc_69 N_A3_c_63_n N_VPWR_c_211_n 0.0113988f $X=0.475 $Y=2.14 $X2=0 $Y2=0
cc_70 A3 N_VPWR_c_211_n 0.00488717f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_71 N_A3_c_55_n N_VPWR_c_212_n 0.00347761f $X=0.36 $Y=2.065 $X2=0 $Y2=0
cc_72 N_A3_c_58_n N_VPWR_c_212_n 8.99341e-19 $X=0.27 $Y=1.625 $X2=0 $Y2=0
cc_73 N_A3_c_63_n N_VPWR_c_212_n 0.00280745f $X=0.475 $Y=2.14 $X2=0 $Y2=0
cc_74 A3 N_VPWR_c_212_n 0.0261185f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_75 N_A3_M1005_g N_VPWR_c_214_n 0.00499542f $X=0.475 $Y=2.685 $X2=0 $Y2=0
cc_76 N_A3_M1005_g N_VPWR_c_208_n 0.0100747f $X=0.475 $Y=2.685 $X2=0 $Y2=0
cc_77 N_A3_M1005_g N_A_110_473#_c_258_n 6.1781e-19 $X=0.475 $Y=2.685 $X2=0 $Y2=0
cc_78 A3 N_VGND_c_310_n 6.17286e-19 $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_79 N_A3_c_56_n N_VGND_c_311_n 0.00496033f $X=0.54 $Y=0.765 $X2=0 $Y2=0
cc_80 A3 N_VGND_c_311_n 0.026511f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_81 N_A3_c_60_n N_VGND_c_311_n 0.00197757f $X=0.27 $Y=1.12 $X2=0 $Y2=0
cc_82 N_A3_c_56_n N_VGND_c_314_n 0.00585385f $X=0.54 $Y=0.765 $X2=0 $Y2=0
cc_83 N_A3_c_56_n N_VGND_c_315_n 0.0115375f $X=0.54 $Y=0.765 $X2=0 $Y2=0
cc_84 A3 N_VGND_c_315_n 0.00239164f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_85 N_A2_M1007_g N_A1_M1000_g 0.0241012f $X=0.93 $Y=0.445 $X2=0 $Y2=0
cc_86 A2 N_A1_M1000_g 0.00222999f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_87 N_A2_M1001_g N_A1_M1006_g 0.0386692f $X=0.905 $Y=2.685 $X2=0 $Y2=0
cc_88 N_A2_c_97_n N_A1_M1006_g 0.0150507f $X=0.84 $Y=1.66 $X2=0 $Y2=0
cc_89 A2 N_A1_M1006_g 2.6786e-19 $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_90 N_A2_c_97_n N_A1_c_140_n 0.0241012f $X=0.84 $Y=1.66 $X2=0 $Y2=0
cc_91 N_A2_M1007_g A1 0.00734785f $X=0.93 $Y=0.445 $X2=0 $Y2=0
cc_92 A2 A1 0.0830633f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_93 N_A2_c_99_n N_A1_c_143_n 0.0241012f $X=0.84 $Y=1.32 $X2=0 $Y2=0
cc_94 N_A2_M1001_g N_VPWR_c_211_n 0.0166326f $X=0.905 $Y=2.685 $X2=0 $Y2=0
cc_95 N_A2_c_101_n N_VPWR_c_211_n 0.00220291f $X=0.84 $Y=1.825 $X2=0 $Y2=0
cc_96 A2 N_VPWR_c_211_n 0.023686f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_97 N_A2_M1001_g N_VPWR_c_213_n 0.00278677f $X=0.905 $Y=2.685 $X2=0 $Y2=0
cc_98 N_A2_M1001_g N_VPWR_c_214_n 0.00302501f $X=0.905 $Y=2.685 $X2=0 $Y2=0
cc_99 N_A2_M1001_g N_VPWR_c_208_n 0.0043662f $X=0.905 $Y=2.685 $X2=0 $Y2=0
cc_100 N_A2_M1001_g N_A_110_473#_c_257_n 0.0125362f $X=0.905 $Y=2.685 $X2=0
+ $Y2=0
cc_101 N_A2_M1007_g N_Y_c_282_n 0.00114759f $X=0.93 $Y=0.445 $X2=0 $Y2=0
cc_102 A2 N_Y_c_282_n 0.0078114f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_103 N_A2_M1007_g N_VGND_c_314_n 0.00492889f $X=0.93 $Y=0.445 $X2=0 $Y2=0
cc_104 A2 N_VGND_c_314_n 0.00920537f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_105 N_A2_M1007_g N_VGND_c_315_n 0.00830938f $X=0.93 $Y=0.445 $X2=0 $Y2=0
cc_106 A2 N_VGND_c_315_n 0.0103984f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_107 A2 A_123_47# 0.00165151f $X=0.635 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_108 N_A1_M1006_g N_B1_c_178_n 0.0378741f $X=1.335 $Y=2.685 $X2=-0.19
+ $Y2=-0.245
cc_109 N_A1_c_140_n N_B1_c_178_n 0.0174494f $X=1.41 $Y=1.345 $X2=-0.19
+ $Y2=-0.245
cc_110 A1 N_B1_c_178_n 9.51571e-19 $X=1.115 $Y=0.84 $X2=-0.19 $Y2=-0.245
cc_111 N_A1_M1000_g N_B1_M1003_g 0.0194807f $X=1.32 $Y=0.445 $X2=0 $Y2=0
cc_112 A1 N_B1_M1003_g 7.45043e-19 $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_113 N_A1_c_143_n N_B1_M1003_g 0.0174494f $X=1.41 $Y=1.005 $X2=0 $Y2=0
cc_114 N_A1_M1006_g N_VPWR_c_211_n 0.00239543f $X=1.335 $Y=2.685 $X2=0 $Y2=0
cc_115 A1 N_VPWR_c_211_n 0.0144294f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_116 N_A1_M1006_g N_VPWR_c_213_n 0.00275572f $X=1.335 $Y=2.685 $X2=0 $Y2=0
cc_117 N_A1_M1006_g N_VPWR_c_214_n 0.00302501f $X=1.335 $Y=2.685 $X2=0 $Y2=0
cc_118 N_A1_M1006_g N_VPWR_c_208_n 0.0043662f $X=1.335 $Y=2.685 $X2=0 $Y2=0
cc_119 N_A1_M1006_g N_A_110_473#_c_257_n 0.0125303f $X=1.335 $Y=2.685 $X2=0
+ $Y2=0
cc_120 A1 N_A_110_473#_c_259_n 0.00356597f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_121 N_A1_M1000_g N_Y_c_282_n 0.0111679f $X=1.32 $Y=0.445 $X2=0 $Y2=0
cc_122 A1 N_Y_c_282_n 0.00842484f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_123 N_A1_c_143_n N_Y_c_282_n 0.00350603f $X=1.41 $Y=1.005 $X2=0 $Y2=0
cc_124 N_A1_M1000_g N_Y_c_278_n 0.00342686f $X=1.32 $Y=0.445 $X2=0 $Y2=0
cc_125 N_A1_M1006_g N_Y_c_278_n 0.00573508f $X=1.335 $Y=2.685 $X2=0 $Y2=0
cc_126 A1 N_Y_c_278_n 0.0809654f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_127 N_A1_c_143_n N_Y_c_278_n 0.00436826f $X=1.41 $Y=1.005 $X2=0 $Y2=0
cc_128 N_A1_M1000_g N_VGND_c_314_n 0.00555741f $X=1.32 $Y=0.445 $X2=0 $Y2=0
cc_129 N_A1_M1000_g N_VGND_c_315_n 0.00653426f $X=1.32 $Y=0.445 $X2=0 $Y2=0
cc_130 A1 N_VGND_c_315_n 0.0107885f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_131 N_B1_M1004_g N_VPWR_c_214_n 0.00499542f $X=1.765 $Y=2.685 $X2=0 $Y2=0
cc_132 N_B1_M1004_g N_VPWR_c_208_n 0.0103203f $X=1.765 $Y=2.685 $X2=0 $Y2=0
cc_133 N_B1_M1004_g N_A_110_473#_c_257_n 0.00183415f $X=1.765 $Y=2.685 $X2=0
+ $Y2=0
cc_134 N_B1_M1003_g N_Y_c_282_n 0.00931971f $X=1.89 $Y=0.445 $X2=0 $Y2=0
cc_135 N_B1_c_178_n Y 0.0100936f $X=1.765 $Y=1.9 $X2=0 $Y2=0
cc_136 N_B1_M1004_g Y 0.016727f $X=1.765 $Y=2.685 $X2=0 $Y2=0
cc_137 B1 Y 0.0279205f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_138 N_B1_M1004_g Y 0.00630023f $X=1.765 $Y=2.685 $X2=0 $Y2=0
cc_139 N_B1_c_178_n N_Y_c_278_n 0.0287774f $X=1.765 $Y=1.9 $X2=0 $Y2=0
cc_140 N_B1_M1004_g N_Y_c_278_n 0.00150136f $X=1.765 $Y=2.685 $X2=0 $Y2=0
cc_141 N_B1_M1003_g N_Y_c_278_n 0.0135671f $X=1.89 $Y=0.445 $X2=0 $Y2=0
cc_142 B1 N_Y_c_278_n 0.0676712f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_143 N_B1_c_178_n N_VGND_c_313_n 0.00150452f $X=1.765 $Y=1.9 $X2=0 $Y2=0
cc_144 N_B1_M1003_g N_VGND_c_313_n 0.00483577f $X=1.89 $Y=0.445 $X2=0 $Y2=0
cc_145 B1 N_VGND_c_313_n 0.0193389f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_146 N_B1_M1003_g N_VGND_c_314_n 0.00540919f $X=1.89 $Y=0.445 $X2=0 $Y2=0
cc_147 N_B1_M1003_g N_VGND_c_315_n 0.011116f $X=1.89 $Y=0.445 $X2=0 $Y2=0
cc_148 B1 N_VGND_c_315_n 0.00196923f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_149 N_VPWR_c_210_n N_A_110_473#_c_256_n 0.00153963f $X=0.26 $Y=2.51 $X2=0
+ $Y2=0
cc_150 N_VPWR_c_211_n N_A_110_473#_c_256_n 0.0209251f $X=0.99 $Y=2.08 $X2=0
+ $Y2=0
cc_151 N_VPWR_c_213_n N_A_110_473#_c_256_n 0.00152491f $X=1.12 $Y=2.57 $X2=0
+ $Y2=0
cc_152 N_VPWR_M1001_d N_A_110_473#_c_257_n 0.00176461f $X=0.98 $Y=2.365 $X2=0
+ $Y2=0
cc_153 N_VPWR_c_213_n N_A_110_473#_c_257_n 0.0126348f $X=1.12 $Y=2.57 $X2=0
+ $Y2=0
cc_154 N_VPWR_c_214_n N_A_110_473#_c_257_n 0.0559995f $X=2.16 $Y=3.33 $X2=0
+ $Y2=0
cc_155 N_VPWR_c_208_n N_A_110_473#_c_257_n 0.0310993f $X=2.16 $Y=3.33 $X2=0
+ $Y2=0
cc_156 N_VPWR_c_210_n N_A_110_473#_c_258_n 0.00605088f $X=0.26 $Y=2.51 $X2=0
+ $Y2=0
cc_157 N_VPWR_c_214_n N_A_110_473#_c_258_n 0.0186386f $X=2.16 $Y=3.33 $X2=0
+ $Y2=0
cc_158 N_VPWR_c_208_n N_A_110_473#_c_258_n 0.0101082f $X=2.16 $Y=3.33 $X2=0
+ $Y2=0
cc_159 N_VPWR_c_213_n N_A_110_473#_c_259_n 0.00152267f $X=1.12 $Y=2.57 $X2=0
+ $Y2=0
cc_160 N_VPWR_c_211_n Y 0.00831987f $X=0.99 $Y=2.08 $X2=0 $Y2=0
cc_161 N_VPWR_c_213_n Y 4.34201e-19 $X=1.12 $Y=2.57 $X2=0 $Y2=0
cc_162 N_VPWR_c_213_n Y 0.00586667f $X=1.12 $Y=2.57 $X2=0 $Y2=0
cc_163 N_VPWR_c_214_n Y 0.02546f $X=2.16 $Y=3.33 $X2=0 $Y2=0
cc_164 N_VPWR_c_208_n Y 0.0177378f $X=2.16 $Y=3.33 $X2=0 $Y2=0
cc_165 N_A_110_473#_c_257_n Y 0.00172312f $X=1.42 $Y=2.99 $X2=0 $Y2=0
cc_166 N_A_110_473#_c_259_n Y 0.00159409f $X=1.55 $Y=2.51 $X2=0 $Y2=0
cc_167 N_Y_c_282_n N_VGND_c_314_n 0.0237998f $X=1.76 $Y=0.447 $X2=0 $Y2=0
cc_168 N_Y_M1000_d N_VGND_c_315_n 0.00341334f $X=1.395 $Y=0.235 $X2=0 $Y2=0
cc_169 N_Y_c_282_n N_VGND_c_315_n 0.0174624f $X=1.76 $Y=0.447 $X2=0 $Y2=0
cc_170 N_VGND_c_315_n A_123_47# 0.00245497f $X=2.16 $Y=0 $X2=-0.19 $Y2=-0.245
cc_171 N_VGND_c_315_n A_201_47# 0.00595894f $X=2.16 $Y=0 $X2=-0.19 $Y2=-0.245
