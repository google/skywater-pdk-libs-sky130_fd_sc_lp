* File: sky130_fd_sc_lp__nor4b_m.spice
* Created: Wed Sep  2 10:11:24 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__nor4b_m.pex.spice"
.subckt sky130_fd_sc_lp__nor4b_m  VNB VPB D_N A B C VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* C	C
* B	B
* A	A
* D_N	D_N
* VPB	VPB
* VNB	VNB
MM1008 N_VGND_M1008_d N_D_N_M1008_g N_A_33_68#_M1008_s VNB NSHORT L=0.15 W=0.42
+ AD=0.1365 AS=0.1113 PD=1.07 PS=1.37 NRD=99.996 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.4 A=0.063 P=1.14 MULT=1
MM1000 N_Y_M1000_d N_A_M1000_g N_VGND_M1008_d VNB NSHORT L=0.15 W=0.42 AD=0.0588
+ AS=0.1365 PD=0.7 PS=1.07 NRD=0 NRS=5.712 M=1 R=2.8 SA=75001 SB=75001.6 A=0.063
+ P=1.14 MULT=1
MM1004 N_VGND_M1004_d N_B_M1004_g N_Y_M1000_d VNB NSHORT L=0.15 W=0.42 AD=0.0756
+ AS=0.0588 PD=0.78 PS=0.7 NRD=5.712 NRS=0 M=1 R=2.8 SA=75001.4 SB=75001.1
+ A=0.063 P=1.14 MULT=1
MM1009 N_Y_M1009_d N_C_M1009_g N_VGND_M1004_d VNB NSHORT L=0.15 W=0.42 AD=0.0588
+ AS=0.0756 PD=0.7 PS=0.78 NRD=0 NRS=17.136 M=1 R=2.8 SA=75001.9 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1002 N_VGND_M1002_d N_A_33_68#_M1002_g N_Y_M1009_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75002.4 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1001 N_VPWR_M1001_d N_D_N_M1001_g N_A_33_68#_M1001_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0819 AS=0.1113 PD=0.81 PS=1.37 NRD=9.3772 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002 A=0.063 P=1.14 MULT=1
MM1005 A_312_496# N_A_M1005_g N_VPWR_M1001_d VPB PHIGHVT L=0.15 W=0.42 AD=0.0441
+ AS=0.0819 PD=0.63 PS=0.81 NRD=23.443 NRS=42.1974 M=1 R=2.8 SA=75000.7
+ SB=75001.5 A=0.063 P=1.14 MULT=1
MM1006 A_384_496# N_B_M1006_g A_312_496# VPB PHIGHVT L=0.15 W=0.42 AD=0.0441
+ AS=0.0441 PD=0.63 PS=0.63 NRD=23.443 NRS=23.443 M=1 R=2.8 SA=75001.1
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1007 A_456_496# N_C_M1007_g A_384_496# VPB PHIGHVT L=0.15 W=0.42 AD=0.0441
+ AS=0.0441 PD=0.63 PS=0.63 NRD=23.443 NRS=23.443 M=1 R=2.8 SA=75001.4
+ SB=75000.8 A=0.063 P=1.14 MULT=1
MM1003 N_Y_M1003_d N_A_33_68#_M1003_g A_456_496# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.2016 AS=0.0441 PD=1.8 PS=0.63 NRD=100.844 NRS=23.443 M=1 R=2.8 SA=75001.8
+ SB=75000.4 A=0.063 P=1.14 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9751 P=11.21
*
.include "sky130_fd_sc_lp__nor4b_m.pxi.spice"
*
.ends
*
*
