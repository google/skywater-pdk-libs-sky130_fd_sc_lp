* File: sky130_fd_sc_lp__xor3_lp.pex.spice
* Created: Wed Sep  2 10:41:52 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__XOR3_LP%A 3 7 11 13 20 21
r40 19 21 0.874306 $w=3.3e-07 $l=5e-09 $layer=POLY_cond $X=1 $Y=1.77 $X2=1.005
+ $Y2=1.77
r41 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1 $Y=1.77
+ $X2=1 $Y2=1.77
r42 17 19 42.841 $w=3.3e-07 $l=2.45e-07 $layer=POLY_cond $X=0.755 $Y=1.77 $X2=1
+ $Y2=1.77
r43 15 17 19.2347 $w=3.3e-07 $l=1.1e-07 $layer=POLY_cond $X=0.645 $Y=1.77
+ $X2=0.755 $Y2=1.77
r44 13 20 6.60335 $w=4.78e-07 $l=2.65e-07 $layer=LI1_cond $X=1.075 $Y=2.035
+ $X2=1.075 $Y2=1.77
r45 9 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.005 $Y=1.605
+ $X2=1.005 $Y2=1.77
r46 9 11 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=1.005 $Y=1.605
+ $X2=1.005 $Y2=0.775
r47 5 17 9.34494 $w=2.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.755 $Y=1.935
+ $X2=0.755 $Y2=1.77
r48 5 7 163.979 $w=2.5e-07 $l=6.6e-07 $layer=POLY_cond $X=0.755 $Y=1.935
+ $X2=0.755 $Y2=2.595
r49 1 15 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.645 $Y=1.605
+ $X2=0.645 $Y2=1.77
r50 1 3 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=0.645 $Y=1.605
+ $X2=0.645 $Y2=0.775
.ends

.subckt PM_SKY130_FD_SC_LP__XOR3_LP%A_57_113# 1 2 3 4 15 17 19 20 21 22 24 27 32
+ 35 37 40 41 42 44 45 46 49 51 52 56
c135 15 0 2.45354e-19 $X=1.815 $Y=2.595
r136 56 59 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=3.985 $Y=0.35
+ $X2=3.985 $Y2=0.495
r137 55 62 42.3262 $w=2.79e-07 $l=2.45e-07 $layer=POLY_cond $X=1.57 $Y=1.26
+ $X2=1.815 $Y2=1.26
r138 54 55 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.57
+ $Y=1.26 $X2=1.57 $Y2=1.26
r139 47 49 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=3.675 $Y=2.895
+ $X2=3.675 $Y2=2.745
r140 45 56 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.82 $Y=0.35
+ $X2=3.985 $Y2=0.35
r141 45 46 136.027 $w=1.68e-07 $l=2.085e-06 $layer=LI1_cond $X=3.82 $Y=0.35
+ $X2=1.735 $Y2=0.35
r142 44 54 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.65 $Y=1.095
+ $X2=1.65 $Y2=1.26
r143 43 46 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.65 $Y=0.435
+ $X2=1.735 $Y2=0.35
r144 43 44 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=1.65 $Y=0.435
+ $X2=1.65 $Y2=1.095
r145 41 47 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.51 $Y=2.98
+ $X2=3.675 $Y2=2.895
r146 41 42 128.85 $w=1.68e-07 $l=1.975e-06 $layer=LI1_cond $X=3.51 $Y=2.98
+ $X2=1.535 $Y2=2.98
r147 40 42 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.45 $Y=2.895
+ $X2=1.535 $Y2=2.98
r148 39 40 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=1.45 $Y=2.5
+ $X2=1.45 $Y2=2.895
r149 38 52 4.4465 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=0.655 $Y=2.415
+ $X2=0.46 $Y2=2.415
r150 37 39 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.365 $Y=2.415
+ $X2=1.45 $Y2=2.5
r151 37 38 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=1.365 $Y=2.415
+ $X2=0.655 $Y2=2.415
r152 36 51 1.65768 $w=3.3e-07 $l=1.95e-07 $layer=LI1_cond $X=0.655 $Y=1.26
+ $X2=0.46 $Y2=1.26
r153 35 54 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.565 $Y=1.26
+ $X2=1.65 $Y2=1.26
r154 35 36 31.7795 $w=3.28e-07 $l=9.1e-07 $layer=LI1_cond $X=1.565 $Y=1.26
+ $X2=0.655 $Y2=1.26
r155 30 52 2.47594 $w=3.9e-07 $l=8.5e-08 $layer=LI1_cond $X=0.46 $Y=2.33
+ $X2=0.46 $Y2=2.415
r156 30 32 2.65948 $w=3.88e-07 $l=9e-08 $layer=LI1_cond $X=0.46 $Y=2.33 $X2=0.46
+ $Y2=2.24
r157 29 51 4.80229 $w=3.6e-07 $l=1.65e-07 $layer=LI1_cond $X=0.46 $Y=1.425
+ $X2=0.46 $Y2=1.26
r158 29 32 24.0831 $w=3.88e-07 $l=8.15e-07 $layer=LI1_cond $X=0.46 $Y=1.425
+ $X2=0.46 $Y2=2.24
r159 25 51 4.80229 $w=3.6e-07 $l=1.79374e-07 $layer=LI1_cond $X=0.43 $Y=1.095
+ $X2=0.46 $Y2=1.26
r160 25 27 11.1752 $w=3.28e-07 $l=3.2e-07 $layer=LI1_cond $X=0.43 $Y=1.095
+ $X2=0.43 $Y2=0.775
r161 22 24 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.465 $Y=1.095
+ $X2=2.465 $Y2=0.775
r162 20 22 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.39 $Y=1.17
+ $X2=2.465 $Y2=1.095
r163 20 21 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=2.39 $Y=1.17
+ $X2=2.15 $Y2=1.17
r164 17 21 23.196 $w=2.79e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.075 $Y=1.095
+ $X2=2.15 $Y2=1.17
r165 17 62 44.9176 $w=2.79e-07 $l=3.32415e-07 $layer=POLY_cond $X=2.075 $Y=1.095
+ $X2=1.815 $Y2=1.26
r166 17 19 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.075 $Y=1.095
+ $X2=2.075 $Y2=0.775
r167 13 62 5.44115 $w=2.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.815 $Y=1.425
+ $X2=1.815 $Y2=1.26
r168 13 15 290.691 $w=2.5e-07 $l=1.17e-06 $layer=POLY_cond $X=1.815 $Y=1.425
+ $X2=1.815 $Y2=2.595
r169 4 49 600 $w=1.7e-07 $l=7.16589e-07 $layer=licon1_PDIFF $count=1 $X=3.535
+ $Y=2.095 $X2=3.675 $Y2=2.745
r170 3 32 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=0.345
+ $Y=2.095 $X2=0.49 $Y2=2.24
r171 2 59 182 $w=1.7e-07 $l=2.77489e-07 $layer=licon1_NDIFF $count=1 $X=3.765
+ $Y=0.625 $X2=3.985 $Y2=0.495
r172 1 27 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.285
+ $Y=0.565 $X2=0.43 $Y2=0.775
.ends

.subckt PM_SKY130_FD_SC_LP__XOR3_LP%B 3 7 10 14 15 16 18 19 23 27 29 33 35 36 37
+ 38 42 43 47 48 50 51 54 58 61 67
c171 48 0 1.30871e-19 $X=4.32 $Y=1.73
c172 43 0 2.42794e-20 $X=3.78 $Y=1.32
c173 38 0 1.12683e-19 $X=3.615 $Y=1.73
c174 35 0 1.96436e-19 $X=2.47 $Y=1.73
c175 16 0 1.29442e-19 $X=4.79 $Y=1.09
r176 54 55 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.88
+ $Y=1.73 $X2=2.88 $Y2=1.73
r177 51 67 3.84148 $w=3.43e-07 $l=1.15e-07 $layer=LI1_cond $X=3.12 $Y=1.722
+ $X2=3.235 $Y2=1.722
r178 51 55 8.01699 $w=3.43e-07 $l=2.4e-07 $layer=LI1_cond $X=3.12 $Y=1.722
+ $X2=2.88 $Y2=1.722
r179 48 62 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.32 $Y=1.73
+ $X2=4.32 $Y2=1.895
r180 48 61 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.32 $Y=1.73
+ $X2=4.32 $Y2=1.565
r181 47 48 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.32
+ $Y=1.73 $X2=4.32 $Y2=1.73
r182 45 50 5.16603 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=3.945 $Y=1.73
+ $X2=3.78 $Y2=1.73
r183 45 47 13.0959 $w=3.28e-07 $l=3.75e-07 $layer=LI1_cond $X=3.945 $Y=1.73
+ $X2=4.32 $Y2=1.73
r184 43 58 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.78 $Y=1.32
+ $X2=3.78 $Y2=1.155
r185 42 43 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.78
+ $Y=1.32 $X2=3.78 $Y2=1.32
r186 40 50 1.34256 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=3.78 $Y=1.565
+ $X2=3.78 $Y2=1.73
r187 40 42 8.55602 $w=3.28e-07 $l=2.45e-07 $layer=LI1_cond $X=3.78 $Y=1.565
+ $X2=3.78 $Y2=1.32
r188 38 50 5.16603 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=3.615 $Y=1.73
+ $X2=3.78 $Y2=1.73
r189 38 67 13.2706 $w=3.28e-07 $l=3.8e-07 $layer=LI1_cond $X=3.615 $Y=1.73
+ $X2=3.235 $Y2=1.73
r190 35 54 71.6931 $w=3.3e-07 $l=4.1e-07 $layer=POLY_cond $X=2.47 $Y=1.73
+ $X2=2.88 $Y2=1.73
r191 31 33 223.053 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.51 $Y=1.09
+ $X2=6.51 $Y2=0.655
r192 30 37 15.684 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=6.225 $Y=1.165
+ $X2=6.05 $Y2=1.165
r193 29 31 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.435 $Y=1.165
+ $X2=6.51 $Y2=1.09
r194 29 30 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=6.435 $Y=1.165
+ $X2=6.225 $Y2=1.165
r195 25 37 8.77658 $w=1.5e-07 $l=1.32288e-07 $layer=POLY_cond $X=6.15 $Y=1.09
+ $X2=6.05 $Y2=1.165
r196 25 27 223.053 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.15 $Y=1.09
+ $X2=6.15 $Y2=0.655
r197 21 37 8.77658 $w=2.5e-07 $l=9.68246e-08 $layer=POLY_cond $X=6 $Y=1.24
+ $X2=6.05 $Y2=1.165
r198 21 23 308.082 $w=2.5e-07 $l=1.24e-06 $layer=POLY_cond $X=6 $Y=1.24 $X2=6
+ $Y2=2.48
r199 20 36 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.865 $Y=1.165
+ $X2=4.79 $Y2=1.165
r200 19 37 15.684 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=5.875 $Y=1.165
+ $X2=6.05 $Y2=1.165
r201 19 20 517.894 $w=1.5e-07 $l=1.01e-06 $layer=POLY_cond $X=5.875 $Y=1.165
+ $X2=4.865 $Y2=1.165
r202 16 36 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.79 $Y=1.09
+ $X2=4.79 $Y2=1.165
r203 16 18 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=4.79 $Y=1.09
+ $X2=4.79 $Y2=0.805
r204 14 36 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.715 $Y=1.165
+ $X2=4.79 $Y2=1.165
r205 14 15 117.936 $w=1.5e-07 $l=2.3e-07 $layer=POLY_cond $X=4.715 $Y=1.165
+ $X2=4.485 $Y2=1.165
r206 12 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.41 $Y=1.24
+ $X2=4.485 $Y2=1.165
r207 12 61 166.649 $w=1.5e-07 $l=3.25e-07 $layer=POLY_cond $X=4.41 $Y=1.24
+ $X2=4.41 $Y2=1.565
r208 10 62 173.918 $w=2.5e-07 $l=7e-07 $layer=POLY_cond $X=4.28 $Y=2.595
+ $X2=4.28 $Y2=1.895
r209 7 58 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=3.69 $Y=0.835
+ $X2=3.69 $Y2=1.155
r210 1 35 27.6025 $w=3.3e-07 $l=2.18746e-07 $layer=POLY_cond $X=2.345 $Y=1.895
+ $X2=2.47 $Y2=1.73
r211 1 3 173.918 $w=2.5e-07 $l=7e-07 $layer=POLY_cond $X=2.345 $Y=1.895
+ $X2=2.345 $Y2=2.595
.ends

.subckt PM_SKY130_FD_SC_LP__XOR3_LP%A_580_21# 1 2 10 11 12 13 14 19 21 23 24 26
+ 28 31 32 33 34 35 36 40 43 46 49 53 54
c147 53 0 8.21899e-20 $X=5.515 $Y=0.43
c148 34 0 3.57353e-19 $X=3.395 $Y=1.875
c149 26 0 1.95972e-19 $X=4.82 $Y=2.08
c150 14 0 9.95572e-20 $X=3.05 $Y=1.195
c151 13 0 1.12683e-19 $X=3.255 $Y=1.195
c152 11 0 1.64741e-20 $X=4.125 $Y=0.18
r153 54 56 7.70806 $w=4.59e-07 $l=2.9e-07 $layer=LI1_cond $X=5.645 $Y=0.575
+ $X2=5.935 $Y2=0.575
r154 52 54 3.45534 $w=4.59e-07 $l=1.3e-07 $layer=LI1_cond $X=5.515 $Y=0.575
+ $X2=5.645 $Y2=0.575
r155 52 53 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.515
+ $Y=0.43 $X2=5.515 $Y2=0.43
r156 48 49 1.3969 $w=3.28e-07 $l=4e-08 $layer=LI1_cond $X=5.605 $Y=1.615
+ $X2=5.645 $Y2=1.615
r157 46 61 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=5.47 $Y=1.615
+ $X2=5.47 $Y2=1.705
r158 45 48 4.71454 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=5.47 $Y=1.615
+ $X2=5.605 $Y2=1.615
r159 45 46 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.47
+ $Y=1.615 $X2=5.47 $Y2=1.615
r160 43 49 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.645 $Y=1.45
+ $X2=5.645 $Y2=1.615
r161 42 54 6.62291 $w=1.7e-07 $l=3.1e-07 $layer=LI1_cond $X=5.645 $Y=0.885
+ $X2=5.645 $Y2=0.575
r162 42 43 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=5.645 $Y=0.885
+ $X2=5.645 $Y2=1.45
r163 38 48 2.36532 $w=2.5e-07 $l=1.65e-07 $layer=LI1_cond $X=5.605 $Y=1.78
+ $X2=5.605 $Y2=1.615
r164 38 40 15.9037 $w=2.48e-07 $l=3.45e-07 $layer=LI1_cond $X=5.605 $Y=1.78
+ $X2=5.605 $Y2=2.125
r165 37 53 30.6007 $w=3.3e-07 $l=1.75e-07 $layer=POLY_cond $X=5.515 $Y=0.255
+ $X2=5.515 $Y2=0.43
r166 33 34 47.1291 $w=2.5e-07 $l=1.5e-07 $layer=POLY_cond $X=3.395 $Y=1.725
+ $X2=3.395 $Y2=1.875
r167 31 61 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.305 $Y=1.705
+ $X2=5.47 $Y2=1.705
r168 31 32 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=5.305 $Y=1.705
+ $X2=4.945 $Y2=1.705
r169 29 32 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.87 $Y=1.78
+ $X2=4.945 $Y2=1.705
r170 29 36 89.734 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=4.87 $Y=1.78
+ $X2=4.87 $Y2=1.955
r171 26 36 40.9178 $w=2.5e-07 $l=1.25e-07 $layer=POLY_cond $X=4.82 $Y=2.08
+ $X2=4.82 $Y2=1.955
r172 26 28 99.292 $w=2.5e-07 $l=5.15e-07 $layer=POLY_cond $X=4.82 $Y=2.08
+ $X2=4.82 $Y2=2.595
r173 25 35 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.275 $Y=0.18
+ $X2=4.2 $Y2=0.18
r174 24 37 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=5.35 $Y=0.18
+ $X2=5.515 $Y2=0.255
r175 24 25 551.223 $w=1.5e-07 $l=1.075e-06 $layer=POLY_cond $X=5.35 $Y=0.18
+ $X2=4.275 $Y2=0.18
r176 21 35 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.2 $Y=0.255
+ $X2=4.2 $Y2=0.18
r177 21 23 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=4.2 $Y=0.255 $X2=4.2
+ $Y2=0.54
r178 19 34 178.887 $w=2.5e-07 $l=7.2e-07 $layer=POLY_cond $X=3.41 $Y=2.595
+ $X2=3.41 $Y2=1.875
r179 15 33 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=3.33 $Y=1.27
+ $X2=3.33 $Y2=1.725
r180 13 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.255 $Y=1.195
+ $X2=3.33 $Y2=1.27
r181 13 14 105.117 $w=1.5e-07 $l=2.05e-07 $layer=POLY_cond $X=3.255 $Y=1.195
+ $X2=3.05 $Y2=1.195
r182 11 35 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.125 $Y=0.18
+ $X2=4.2 $Y2=0.18
r183 11 12 551.223 $w=1.5e-07 $l=1.075e-06 $layer=POLY_cond $X=4.125 $Y=0.18
+ $X2=3.05 $Y2=0.18
r184 8 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.975 $Y=1.12
+ $X2=3.05 $Y2=1.195
r185 8 10 176.904 $w=1.5e-07 $l=3.45e-07 $layer=POLY_cond $X=2.975 $Y=1.12
+ $X2=2.975 $Y2=0.775
r186 7 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.975 $Y=0.255
+ $X2=3.05 $Y2=0.18
r187 7 10 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=2.975 $Y=0.255
+ $X2=2.975 $Y2=0.775
r188 2 40 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=5.5
+ $Y=1.98 $X2=5.645 $Y2=2.125
r189 1 56 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=5.79
+ $Y=0.445 $X2=5.935 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__XOR3_LP%A_1393_300# 1 2 9 13 17 20 22 24 28 32 46 48
r85 46 48 171.777 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=8.195 $Y=1.31
+ $X2=8.53 $Y2=1.31
r86 32 48 60.2004 $w=3.3e-07 $l=2.45e-07 $layer=POLY_cond $X=8.775 $Y=1.4
+ $X2=8.53 $Y2=1.4
r87 31 34 23.337 $w=3.98e-07 $l=8.1e-07 $layer=LI1_cond $X=8.865 $Y=1.4
+ $X2=8.865 $Y2=2.21
r88 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.775
+ $Y=1.4 $X2=8.775 $Y2=1.4
r89 28 31 13.9734 $w=3.98e-07 $l=4.85e-07 $layer=LI1_cond $X=8.865 $Y=0.915
+ $X2=8.865 $Y2=1.4
r90 25 46 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.03 $Y=1.4
+ $X2=8.195 $Y2=1.4
r91 25 43 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=8.03 $Y=1.4 $X2=8.01
+ $Y2=1.4
r92 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.03
+ $Y=1.4 $X2=8.03 $Y2=1.4
r93 22 24 13.6198 $w=3.28e-07 $l=3.9e-07 $layer=LI1_cond $X=7.64 $Y=1.4 $X2=8.03
+ $Y2=1.4
r94 20 42 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.13 $Y=1.665
+ $X2=7.13 $Y2=1.83
r95 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.13
+ $Y=1.665 $X2=7.13 $Y2=1.665
r96 17 22 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=7.555 $Y=1.665
+ $X2=7.555 $Y2=1.4
r97 17 19 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=7.47 $Y=1.665
+ $X2=7.13 $Y2=1.665
r98 11 43 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.01 $Y=1.235
+ $X2=8.01 $Y2=1.4
r99 11 13 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=8.01 $Y=1.235
+ $X2=8.01 $Y2=0.825
r100 9 42 173.918 $w=2.5e-07 $l=7e-07 $layer=POLY_cond $X=7.17 $Y=2.53 $X2=7.17
+ $Y2=1.83
r101 2 34 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=8.755
+ $Y=2.065 $X2=8.9 $Y2=2.21
r102 1 28 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=8.755
+ $Y=0.705 $X2=8.9 $Y2=0.915
.ends

.subckt PM_SKY130_FD_SC_LP__XOR3_LP%C 3 5 6 8 9 11 13 14 16 18 19 21 22 23 24 26
+ 28 29 35
c90 35 0 1.86955e-19 $X=9.495 $Y=1.4
c91 23 0 2.48255e-19 $X=7.565 $Y=1.26
c92 19 0 1.33731e-19 $X=9.585 $Y=1.235
c93 11 0 1.75882e-19 $X=9.165 $Y=1.955
r94 35 37 16.3083 $w=2.66e-07 $l=9e-08 $layer=POLY_cond $X=9.495 $Y=1.4
+ $X2=9.585 $Y2=1.4
r95 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.495
+ $Y=1.4 $X2=9.495 $Y2=1.4
r96 33 35 16.3083 $w=2.66e-07 $l=9e-08 $layer=POLY_cond $X=9.405 $Y=1.4
+ $X2=9.495 $Y2=1.4
r97 29 36 10.3271 $w=3.83e-07 $l=3.45e-07 $layer=LI1_cond $X=9.84 $Y=1.372
+ $X2=9.495 $Y2=1.372
r98 28 36 4.04103 $w=3.83e-07 $l=1.35e-07 $layer=LI1_cond $X=9.36 $Y=1.372
+ $X2=9.495 $Y2=1.372
r99 22 23 58.3064 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=7.565 $Y=1.11
+ $X2=7.565 $Y2=1.26
r100 19 37 16.1576 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.585 $Y=1.235
+ $X2=9.585 $Y2=1.4
r101 19 21 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=9.585 $Y=1.235
+ $X2=9.585 $Y2=0.915
r102 18 26 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.405 $Y=1.805
+ $X2=9.405 $Y2=1.88
r103 17 33 16.1576 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.405 $Y=1.565
+ $X2=9.405 $Y2=1.4
r104 17 18 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=9.405 $Y=1.565
+ $X2=9.405 $Y2=1.805
r105 14 33 32.6165 $w=2.66e-07 $l=2.49199e-07 $layer=POLY_cond $X=9.225 $Y=1.235
+ $X2=9.405 $Y2=1.4
r106 14 16 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=9.225 $Y=1.235
+ $X2=9.225 $Y2=0.915
r107 11 26 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=9.165 $Y=1.88
+ $X2=9.405 $Y2=1.88
r108 11 13 117.608 $w=2.5e-07 $l=6.1e-07 $layer=POLY_cond $X=9.165 $Y=1.955
+ $X2=9.165 $Y2=2.565
r109 10 24 9.46703 $w=1.5e-07 $l=1.6e-07 $layer=POLY_cond $X=7.825 $Y=1.88
+ $X2=7.665 $Y2=1.88
r110 9 11 64.0957 $w=1.5e-07 $l=1.25e-07 $layer=POLY_cond $X=9.04 $Y=1.88
+ $X2=9.165 $Y2=1.88
r111 9 10 623.011 $w=1.5e-07 $l=1.215e-06 $layer=POLY_cond $X=9.04 $Y=1.88
+ $X2=7.825 $Y2=1.88
r112 6 24 15.9654 $w=2e-07 $l=9.08295e-08 $layer=POLY_cond $X=7.7 $Y=1.955
+ $X2=7.665 $Y2=1.88
r113 6 8 110.86 $w=2.5e-07 $l=5.75e-07 $layer=POLY_cond $X=7.7 $Y=1.955 $X2=7.7
+ $Y2=2.53
r114 5 24 15.9654 $w=2e-07 $l=1.16619e-07 $layer=POLY_cond $X=7.58 $Y=1.805
+ $X2=7.665 $Y2=1.88
r115 5 23 279.457 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=7.58 $Y=1.805
+ $X2=7.58 $Y2=1.26
r116 3 22 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=7.55 $Y=0.825
+ $X2=7.55 $Y2=1.11
.ends

.subckt PM_SKY130_FD_SC_LP__XOR3_LP%A_1459_406# 1 2 9 14 15 17 20 24 25 28 30 31
+ 33 34 35 38 39 49
c110 39 0 6.45953e-20 $X=10.3 $Y=1.4
c111 38 0 1.86955e-19 $X=10.3 $Y=1.4
c112 30 0 1.33731e-19 $X=9.87 $Y=0.35
r113 51 52 11.2294 $w=5.58e-07 $l=1.3e-07 $layer=POLY_cond $X=10.025 $Y=1.57
+ $X2=10.155 $Y2=1.57
r114 45 49 20.9834 $w=3.3e-07 $l=1.2e-07 $layer=POLY_cond $X=10.035 $Y=0.43
+ $X2=10.155 $Y2=0.43
r115 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.035
+ $Y=0.43 $X2=10.035 $Y2=0.43
r116 39 52 12.5251 $w=5.58e-07 $l=1.45e-07 $layer=POLY_cond $X=10.3 $Y=1.57
+ $X2=10.155 $Y2=1.57
r117 38 39 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=10.3
+ $Y=1.4 $X2=10.3 $Y2=1.4
r118 36 38 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=10.3 $Y=1.745
+ $X2=10.3 $Y2=1.4
r119 34 36 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=10.135 $Y=1.83
+ $X2=10.3 $Y2=1.745
r120 34 35 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=10.135 $Y=1.83
+ $X2=9.415 $Y2=1.83
r121 32 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.33 $Y=1.915
+ $X2=9.415 $Y2=1.83
r122 32 33 63.9358 $w=1.68e-07 $l=9.8e-07 $layer=LI1_cond $X=9.33 $Y=1.915
+ $X2=9.33 $Y2=2.895
r123 30 44 3.35256 $w=2.73e-07 $l=8e-08 $layer=LI1_cond $X=10.007 $Y=0.35
+ $X2=10.007 $Y2=0.43
r124 30 31 124.61 $w=1.68e-07 $l=1.91e-06 $layer=LI1_cond $X=9.87 $Y=0.35
+ $X2=7.96 $Y2=0.35
r125 26 31 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=7.795 $Y=0.435
+ $X2=7.96 $Y2=0.35
r126 26 28 13.6198 $w=3.28e-07 $l=3.9e-07 $layer=LI1_cond $X=7.795 $Y=0.435
+ $X2=7.795 $Y2=0.825
r127 24 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.245 $Y=2.98
+ $X2=9.33 $Y2=2.895
r128 24 25 107.321 $w=1.68e-07 $l=1.645e-06 $layer=LI1_cond $X=9.245 $Y=2.98
+ $X2=7.6 $Y2=2.98
r129 20 23 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=7.435 $Y=2.175
+ $X2=7.435 $Y2=2.885
r130 18 25 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=7.435 $Y=2.895
+ $X2=7.6 $Y2=2.98
r131 18 23 0.349225 $w=3.28e-07 $l=1e-08 $layer=LI1_cond $X=7.435 $Y=2.895
+ $X2=7.435 $Y2=2.885
r132 15 39 21.1631 $w=5.58e-07 $l=4.40795e-07 $layer=POLY_cond $X=10.545
+ $Y=1.235 $X2=10.3 $Y2=1.57
r133 15 17 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=10.545 $Y=1.235
+ $X2=10.545 $Y2=0.915
r134 12 52 34.2028 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=10.155 $Y=1.235
+ $X2=10.155 $Y2=1.57
r135 12 14 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=10.155 $Y=1.235
+ $X2=10.155 $Y2=0.915
r136 11 49 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.155 $Y=0.595
+ $X2=10.155 $Y2=0.43
r137 11 14 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=10.155 $Y=0.595
+ $X2=10.155 $Y2=0.915
r138 7 51 21.5669 $w=2.5e-07 $l=3.35e-07 $layer=POLY_cond $X=10.025 $Y=1.905
+ $X2=10.025 $Y2=1.57
r139 7 9 163.979 $w=2.5e-07 $l=6.6e-07 $layer=POLY_cond $X=10.025 $Y=1.905
+ $X2=10.025 $Y2=2.565
r140 2 23 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=7.295
+ $Y=2.03 $X2=7.435 $Y2=2.885
r141 2 20 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=7.295
+ $Y=2.03 $X2=7.435 $Y2=2.175
r142 1 28 182 $w=1.7e-07 $l=2.82489e-07 $layer=licon1_NDIFF $count=1 $X=7.625
+ $Y=0.615 $X2=7.795 $Y2=0.825
.ends

.subckt PM_SKY130_FD_SC_LP__XOR3_LP%VPWR 1 2 3 12 16 22 25 26 28 29 30 42 51 52
+ 55
r88 55 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r89 52 56 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=10.8 $Y=3.33
+ $X2=9.84 $Y2=3.33
r90 51 52 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.8 $Y=3.33
+ $X2=10.8 $Y2=3.33
r91 49 55 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.925 $Y=3.33
+ $X2=9.76 $Y2=3.33
r92 49 51 57.0856 $w=1.68e-07 $l=8.75e-07 $layer=LI1_cond $X=9.925 $Y=3.33
+ $X2=10.8 $Y2=3.33
r93 48 56 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=9.84 $Y2=3.33
r94 47 48 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r95 45 48 0.802756 $w=4.9e-07 $l=2.88e-06 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=9.36 $Y2=3.33
r96 44 47 187.893 $w=1.68e-07 $l=2.88e-06 $layer=LI1_cond $X=6.48 $Y=3.33
+ $X2=9.36 $Y2=3.33
r97 44 45 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r98 42 55 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.595 $Y=3.33
+ $X2=9.76 $Y2=3.33
r99 42 47 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=9.595 $Y=3.33
+ $X2=9.36 $Y2=3.33
r100 41 45 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=6.48
+ $Y2=3.33
r101 40 41 1.69091 $w=1.7e-07 $l=9.35e-07 $layer=mcon $count=5 $X=6 $Y=3.33
+ $X2=6 $Y2=3.33
r102 37 40 313.155 $w=1.68e-07 $l=4.8e-06 $layer=LI1_cond $X=1.2 $Y=3.33 $X2=6
+ $Y2=3.33
r103 37 38 1.69091 $w=1.7e-07 $l=9.35e-07 $layer=mcon $count=5 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r104 34 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r105 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r106 30 41 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33 $X2=6
+ $Y2=3.33
r107 30 38 1.20413 $w=4.9e-07 $l=4.32e-06 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=1.2 $Y2=3.33
r108 28 40 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=6.26 $Y=3.33 $X2=6
+ $Y2=3.33
r109 28 29 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.26 $Y=3.33
+ $X2=6.345 $Y2=3.33
r110 27 44 3.26203 $w=1.68e-07 $l=5e-08 $layer=LI1_cond $X=6.43 $Y=3.33 $X2=6.48
+ $Y2=3.33
r111 27 29 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.43 $Y=3.33
+ $X2=6.345 $Y2=3.33
r112 25 33 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=0.855 $Y=3.33
+ $X2=0.72 $Y2=3.33
r113 25 26 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.855 $Y=3.33
+ $X2=1.02 $Y2=3.33
r114 24 37 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=1.185 $Y=3.33
+ $X2=1.2 $Y2=3.33
r115 24 26 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.185 $Y=3.33
+ $X2=1.02 $Y2=3.33
r116 20 55 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.76 $Y=3.245
+ $X2=9.76 $Y2=3.33
r117 20 22 34.3987 $w=3.28e-07 $l=9.85e-07 $layer=LI1_cond $X=9.76 $Y=3.245
+ $X2=9.76 $Y2=2.26
r118 16 19 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=6.345 $Y=2.125
+ $X2=6.345 $Y2=2.835
r119 14 29 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.345 $Y=3.245
+ $X2=6.345 $Y2=3.33
r120 14 19 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=6.345 $Y=3.245
+ $X2=6.345 $Y2=2.835
r121 10 26 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.02 $Y=3.245
+ $X2=1.02 $Y2=3.33
r122 10 12 12.2229 $w=3.28e-07 $l=3.5e-07 $layer=LI1_cond $X=1.02 $Y=3.245
+ $X2=1.02 $Y2=2.895
r123 3 22 300 $w=1.7e-07 $l=5.59062e-07 $layer=licon1_PDIFF $count=2 $X=9.29
+ $Y=2.065 $X2=9.76 $Y2=2.26
r124 2 19 400 $w=1.7e-07 $l=9.5871e-07 $layer=licon1_PDIFF $count=1 $X=6.125
+ $Y=1.98 $X2=6.345 $Y2=2.835
r125 2 16 400 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_PDIFF $count=1 $X=6.125
+ $Y=1.98 $X2=6.345 $Y2=2.125
r126 1 12 600 $w=1.7e-07 $l=8.67179e-07 $layer=licon1_PDIFF $count=1 $X=0.88
+ $Y=2.095 $X2=1.02 $Y2=2.895
.ends

.subckt PM_SKY130_FD_SC_LP__XOR3_LP%A_388_419# 1 2 3 4 13 15 17 19 21 23 26 30
+ 31 32 38
c117 38 0 2.51578e-19 $X=5.04 $Y=0.925
c118 32 0 1.96436e-19 $X=2.305 $Y=0.925
c119 31 0 4.07535e-20 $X=4.895 $Y=0.925
c120 19 0 1.89925e-19 $X=5.04 $Y=1.04
c121 15 0 9.95572e-20 $X=2.08 $Y=2.395
c122 13 0 1.81544e-19 $X=2.08 $Y=1.005
r123 38 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0.925
+ $X2=5.04 $Y2=0.925
r124 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0.925
+ $X2=2.16 $Y2=0.925
r125 32 34 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.305 $Y=0.925
+ $X2=2.16 $Y2=0.925
r126 31 38 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.895 $Y=0.925
+ $X2=5.04 $Y2=0.925
r127 31 32 3.20544 $w=1.4e-07 $l=2.59e-06 $layer=MET1_cond $X=4.895 $Y=0.925
+ $X2=2.305 $Y2=0.925
r128 26 28 4.60977 $w=3.28e-07 $l=1.32e-07 $layer=LI1_cond $X=2.68 $Y=0.775
+ $X2=2.68 $Y2=0.907
r129 21 30 7.79447 $w=2.93e-07 $l=1.47e-07 $layer=LI1_cond $X=5.102 $Y=2.107
+ $X2=5.102 $Y2=1.96
r130 21 23 11.251 $w=2.93e-07 $l=2.88e-07 $layer=LI1_cond $X=5.102 $Y=2.107
+ $X2=5.102 $Y2=2.395
r131 19 43 11.5608 $w=3.28e-07 $l=2.51893e-07 $layer=LI1_cond $X=5.04 $Y=1.04
+ $X2=5.005 $Y2=0.805
r132 19 30 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=5.04 $Y=1.04
+ $X2=5.04 $Y2=1.96
r133 18 35 4.65494 $w=1.95e-07 $l=1.65e-07 $layer=LI1_cond $X=2.245 $Y=0.907
+ $X2=2.08 $Y2=0.907
r134 17 28 3.83364 $w=1.95e-07 $l=1.65e-07 $layer=LI1_cond $X=2.515 $Y=0.907
+ $X2=2.68 $Y2=0.907
r135 17 18 15.3566 $w=1.93e-07 $l=2.7e-07 $layer=LI1_cond $X=2.515 $Y=0.907
+ $X2=2.245 $Y2=0.907
r136 13 35 2.76475 $w=3.3e-07 $l=9.8e-08 $layer=LI1_cond $X=2.08 $Y=1.005
+ $X2=2.08 $Y2=0.907
r137 13 15 48.5423 $w=3.28e-07 $l=1.39e-06 $layer=LI1_cond $X=2.08 $Y=1.005
+ $X2=2.08 $Y2=2.395
r138 4 23 600 $w=1.7e-07 $l=3.63318e-07 $layer=licon1_PDIFF $count=1 $X=4.945
+ $Y=2.095 $X2=5.085 $Y2=2.395
r139 3 15 600 $w=1.7e-07 $l=3.63318e-07 $layer=licon1_PDIFF $count=1 $X=1.94
+ $Y=2.095 $X2=2.08 $Y2=2.395
r140 2 43 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=4.865
+ $Y=0.595 $X2=5.005 $Y2=0.805
r141 1 26 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.54
+ $Y=0.565 $X2=2.68 $Y2=0.775
.ends

.subckt PM_SKY130_FD_SC_LP__XOR3_LP%A_494_419# 1 2 3 4 14 17 19 20 21 25 28 29
+ 30 32 33 34 39 41 43 44 46 47 49
c145 49 0 1.95889e-19 $X=7.285 $Y=0.825
c146 43 0 8.60881e-20 $X=2.6 $Y=2.16
c147 21 0 3.38679e-19 $X=4.02 $Y=2.16
c148 19 0 1.61987e-19 $X=3.105 $Y=1.27
c149 17 0 1.59266e-19 $X=2.61 $Y=2.395
r150 49 50 18.4576 $w=2.71e-07 $l=4.1e-07 $layer=LI1_cond $X=7.285 $Y=0.825
+ $X2=7.285 $Y2=1.235
r151 46 47 9.25191 $w=4.53e-07 $l=1.65e-07 $layer=LI1_cond $X=6.842 $Y=2.175
+ $X2=6.842 $Y2=2.01
r152 42 44 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.785 $Y=1.235
+ $X2=6.7 $Y2=1.235
r153 41 50 3.46554 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.12 $Y=1.235
+ $X2=7.285 $Y2=1.235
r154 41 42 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=7.12 $Y=1.235
+ $X2=6.785 $Y2=1.235
r155 37 46 1.62982 $w=4.53e-07 $l=6.2e-08 $layer=LI1_cond $X=6.842 $Y=2.237
+ $X2=6.842 $Y2=2.175
r156 37 39 17.0343 $w=4.53e-07 $l=6.48e-07 $layer=LI1_cond $X=6.842 $Y=2.237
+ $X2=6.842 $Y2=2.885
r157 35 44 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.7 $Y=1.32 $X2=6.7
+ $Y2=1.235
r158 35 47 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=6.7 $Y=1.32 $X2=6.7
+ $Y2=2.01
r159 33 44 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.615 $Y=1.235
+ $X2=6.7 $Y2=1.235
r160 33 34 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=6.615 $Y=1.235
+ $X2=6.08 $Y2=1.235
r161 31 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.995 $Y=1.32
+ $X2=6.08 $Y2=1.235
r162 31 32 102.754 $w=1.68e-07 $l=1.575e-06 $layer=LI1_cond $X=5.995 $Y=1.32
+ $X2=5.995 $Y2=2.895
r163 29 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.91 $Y=2.98
+ $X2=5.995 $Y2=2.895
r164 29 30 112.214 $w=1.68e-07 $l=1.72e-06 $layer=LI1_cond $X=5.91 $Y=2.98
+ $X2=4.19 $Y2=2.98
r165 28 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.105 $Y=2.895
+ $X2=4.19 $Y2=2.98
r166 27 28 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=4.105 $Y=2.245
+ $X2=4.105 $Y2=2.895
r167 23 25 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=3.27 $Y=1.185
+ $X2=3.27 $Y2=0.84
r168 22 43 2.90867 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=2.775 $Y=2.16
+ $X2=2.6 $Y2=2.16
r169 21 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.02 $Y=2.16
+ $X2=4.105 $Y2=2.245
r170 21 22 81.2246 $w=1.68e-07 $l=1.245e-06 $layer=LI1_cond $X=4.02 $Y=2.16
+ $X2=2.775 $Y2=2.16
r171 19 23 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.105 $Y=1.27
+ $X2=3.27 $Y2=1.185
r172 19 20 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=3.105 $Y=1.27
+ $X2=2.595 $Y2=1.27
r173 15 43 3.58051 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=2.6 $Y=2.245 $X2=2.6
+ $Y2=2.16
r174 15 17 4.93904 $w=3.48e-07 $l=1.5e-07 $layer=LI1_cond $X=2.6 $Y=2.245
+ $X2=2.6 $Y2=2.395
r175 14 43 3.58051 $w=2.6e-07 $l=1.25499e-07 $layer=LI1_cond $X=2.51 $Y=2.075
+ $X2=2.6 $Y2=2.16
r176 13 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.51 $Y=1.355
+ $X2=2.595 $Y2=1.27
r177 13 14 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=2.51 $Y=1.355
+ $X2=2.51 $Y2=2.075
r178 4 46 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=6.76
+ $Y=2.03 $X2=6.905 $Y2=2.175
r179 4 39 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=6.76
+ $Y=2.03 $X2=6.905 $Y2=2.885
r180 3 17 600 $w=1.7e-07 $l=3.63318e-07 $layer=licon1_PDIFF $count=1 $X=2.47
+ $Y=2.095 $X2=2.61 $Y2=2.395
r181 2 49 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=7.14
+ $Y=0.615 $X2=7.285 $Y2=0.825
r182 1 25 182 $w=1.7e-07 $l=3.68951e-07 $layer=licon1_NDIFF $count=1 $X=3.05
+ $Y=0.565 $X2=3.27 $Y2=0.84
.ends

.subckt PM_SKY130_FD_SC_LP__XOR3_LP%A_855_66# 1 2 3 4 15 18 20 22 23 26 29 32 33
+ 39
c105 26 0 1.8353e-19 $X=4.69 $Y=1.3
c106 22 0 2.28248e-19 $X=8.4 $Y=2.01
c107 18 0 2.29871e-19 $X=4.415 $Y=1.215
r108 40 50 0.763454 $w=7.03e-07 $l=4.5e-08 $layer=LI1_cond $X=7.92 $Y=2.362
+ $X2=7.965 $Y2=2.362
r109 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=2.405
+ $X2=7.92 $Y2=2.405
r110 35 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=2.405
+ $X2=4.56 $Y2=2.405
r111 33 35 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.705 $Y=2.405
+ $X2=4.56 $Y2=2.405
r112 32 39 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.775 $Y=2.405
+ $X2=7.92 $Y2=2.405
r113 32 33 3.7995 $w=1.4e-07 $l=3.07e-06 $layer=MET1_cond $X=7.775 $Y=2.405
+ $X2=4.705 $Y2=2.405
r114 29 31 10.3166 $w=3.43e-07 $l=2.2e-07 $layer=LI1_cond $X=8.312 $Y=0.835
+ $X2=8.312 $Y2=1.055
r115 24 26 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=4.415 $Y=1.3
+ $X2=4.69 $Y2=1.3
r116 22 50 7.38006 $w=7.03e-07 $l=4.35e-07 $layer=LI1_cond $X=8.4 $Y=2.362
+ $X2=7.965 $Y2=2.362
r117 22 31 62.3048 $w=1.68e-07 $l=9.55e-07 $layer=LI1_cond $X=8.4 $Y=2.01
+ $X2=8.4 $Y2=1.055
r118 20 43 3.84148 $w=4.03e-07 $l=1.35e-07 $layer=LI1_cond $X=4.69 $Y=2.512
+ $X2=4.555 $Y2=2.512
r119 19 26 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.69 $Y=1.385
+ $X2=4.69 $Y2=1.3
r120 19 20 60.3476 $w=1.68e-07 $l=9.25e-07 $layer=LI1_cond $X=4.69 $Y=1.385
+ $X2=4.69 $Y2=2.31
r121 18 24 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.415 $Y=1.215
+ $X2=4.415 $Y2=1.3
r122 18 23 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=4.415 $Y=1.215
+ $X2=4.415 $Y2=1.035
r123 13 23 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=4.495 $Y=0.87
+ $X2=4.495 $Y2=1.035
r124 13 15 13.7944 $w=3.28e-07 $l=3.95e-07 $layer=LI1_cond $X=4.495 $Y=0.87
+ $X2=4.495 $Y2=0.475
r125 4 50 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=7.825
+ $Y=2.03 $X2=7.965 $Y2=2.175
r126 3 43 600 $w=1.7e-07 $l=4.84226e-07 $layer=licon1_PDIFF $count=1 $X=4.405
+ $Y=2.095 $X2=4.555 $Y2=2.51
r127 2 29 182 $w=1.7e-07 $l=3.11127e-07 $layer=licon1_NDIFF $count=1 $X=8.085
+ $Y=0.615 $X2=8.305 $Y2=0.835
r128 1 15 91 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_NDIFF $count=2 $X=4.275
+ $Y=0.33 $X2=4.495 $Y2=0.475
.ends

.subckt PM_SKY130_FD_SC_LP__XOR3_LP%X 1 2 9 12 13 14 15 16 17 26 34
c24 9 0 6.45953e-20 $X=10.675 $Y=2.18
r25 24 34 2.76586 $w=2.48e-07 $l=6e-08 $layer=LI1_cond $X=10.8 $Y=2.095 $X2=10.8
+ $Y2=2.035
r26 16 17 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=10.8 $Y=2.405
+ $X2=10.8 $Y2=2.775
r27 16 35 6.45368 $w=2.48e-07 $l=1.4e-07 $layer=LI1_cond $X=10.8 $Y=2.405
+ $X2=10.8 $Y2=2.265
r28 15 24 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=10.8 $Y=2.18 $X2=10.8
+ $Y2=2.095
r29 15 35 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=10.8 $Y=2.18 $X2=10.8
+ $Y2=2.265
r30 15 34 0.59927 $w=2.48e-07 $l=1.3e-08 $layer=LI1_cond $X=10.8 $Y=2.022
+ $X2=10.8 $Y2=2.035
r31 14 15 16.4569 $w=2.48e-07 $l=3.57e-07 $layer=LI1_cond $X=10.8 $Y=1.665
+ $X2=10.8 $Y2=2.022
r32 13 14 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=10.8 $Y=1.295
+ $X2=10.8 $Y2=1.665
r33 13 26 17.5171 $w=2.48e-07 $l=3.8e-07 $layer=LI1_cond $X=10.8 $Y=1.295
+ $X2=10.8 $Y2=0.915
r34 10 12 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.455 $Y=2.18
+ $X2=10.29 $Y2=2.18
r35 9 15 2.76166 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.675 $Y=2.18
+ $X2=10.8 $Y2=2.18
r36 9 10 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=10.675 $Y=2.18
+ $X2=10.455 $Y2=2.18
r37 2 12 300 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_PDIFF $count=2 $X=10.15
+ $Y=2.065 $X2=10.29 $Y2=2.26
r38 1 26 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=10.62
+ $Y=0.705 $X2=10.76 $Y2=0.915
.ends

.subckt PM_SKY130_FD_SC_LP__XOR3_LP%VGND 1 2 3 12 16 18 23 25 26 28 29 30 32 51
+ 52 55
r84 55 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r85 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=0 $X2=10.8
+ $Y2=0
r86 49 52 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=0 $X2=10.8
+ $Y2=0
r87 48 49 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=10.32 $Y=0
+ $X2=10.32 $Y2=0
r88 46 49 0.936549 $w=4.9e-07 $l=3.36e-06 $layer=MET1_cond $X=6.96 $Y=0
+ $X2=10.32 $Y2=0
r89 45 48 219.209 $w=1.68e-07 $l=3.36e-06 $layer=LI1_cond $X=6.96 $Y=0 $X2=10.32
+ $Y2=0
r90 45 46 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=6.96 $Y=0 $X2=6.96
+ $Y2=0
r91 43 46 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6.96
+ $Y2=0
r92 42 43 1.69091 $w=1.7e-07 $l=9.35e-07 $layer=mcon $count=5 $X=6.48 $Y=0
+ $X2=6.48 $Y2=0
r93 40 56 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r94 39 42 313.155 $w=1.68e-07 $l=4.8e-06 $layer=LI1_cond $X=1.68 $Y=0 $X2=6.48
+ $Y2=0
r95 39 40 1.69091 $w=1.7e-07 $l=9.35e-07 $layer=mcon $count=5 $X=1.68 $Y=0
+ $X2=1.68 $Y2=0
r96 37 55 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.385 $Y=0 $X2=1.22
+ $Y2=0
r97 37 39 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.385 $Y=0 $X2=1.68
+ $Y2=0
r98 35 56 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r99 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r100 32 55 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.055 $Y=0 $X2=1.22
+ $Y2=0
r101 32 34 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.055 $Y=0
+ $X2=0.72 $Y2=0
r102 30 43 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=6.48
+ $Y2=0
r103 30 40 1.07034 $w=4.9e-07 $l=3.84e-06 $layer=MET1_cond $X=5.52 $Y=0 $X2=1.68
+ $Y2=0
r104 28 48 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=10.325 $Y=0
+ $X2=10.32 $Y2=0
r105 28 29 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.325 $Y=0
+ $X2=10.41 $Y2=0
r106 27 51 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=10.495 $Y=0
+ $X2=10.8 $Y2=0
r107 27 29 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.495 $Y=0
+ $X2=10.41 $Y2=0
r108 25 42 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=6.56 $Y=0 $X2=6.48
+ $Y2=0
r109 25 26 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.56 $Y=0 $X2=6.725
+ $Y2=0
r110 24 45 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=6.89 $Y=0 $X2=6.96
+ $Y2=0
r111 24 26 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.89 $Y=0 $X2=6.725
+ $Y2=0
r112 22 29 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.41 $Y=0.085
+ $X2=10.41 $Y2=0
r113 22 23 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=10.41 $Y=0.085
+ $X2=10.41 $Y2=0.775
r114 18 23 6.9898 $w=2.25e-07 $l=1.4854e-07 $layer=LI1_cond $X=10.325 $Y=0.887
+ $X2=10.41 $Y2=0.775
r115 18 20 19.7196 $w=2.23e-07 $l=3.85e-07 $layer=LI1_cond $X=10.325 $Y=0.887
+ $X2=9.94 $Y2=0.887
r116 14 26 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.725 $Y=0.085
+ $X2=6.725 $Y2=0
r117 14 16 19.9058 $w=3.28e-07 $l=5.7e-07 $layer=LI1_cond $X=6.725 $Y=0.085
+ $X2=6.725 $Y2=0.655
r118 10 55 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.22 $Y=0.085
+ $X2=1.22 $Y2=0
r119 10 12 22.525 $w=3.28e-07 $l=6.45e-07 $layer=LI1_cond $X=1.22 $Y=0.085
+ $X2=1.22 $Y2=0.73
r120 3 20 182 $w=1.7e-07 $l=3.58887e-07 $layer=licon1_NDIFF $count=1 $X=9.66
+ $Y=0.705 $X2=9.94 $Y2=0.885
r121 2 16 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=6.585
+ $Y=0.445 $X2=6.725 $Y2=0.655
r122 1 12 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=1.08
+ $Y=0.565 $X2=1.22 $Y2=0.73
.ends

