* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__and4b_lp A_N B C D VGND VNB VPB VPWR X
X0 a_114_47# a_84_21# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 X a_84_21# a_114_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 X a_84_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X3 a_354_47# B a_432_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 a_432_47# a_480_21# a_84_21# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 VPWR D a_84_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X6 VGND A_N a_708_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 a_276_47# C a_354_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 VPWR A_N a_480_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X9 a_84_21# a_480_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X10 a_708_47# A_N a_480_21# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X11 a_84_21# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X12 VPWR B a_84_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X13 VGND D a_276_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
