* File: sky130_fd_sc_lp__dfxbp_1.pex.spice
* Created: Fri Aug 28 10:23:41 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__DFXBP_1%CLK 2 5 8 10 11 12 13 14 20 22
r28 20 22 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=0.362 $Y=1.105
+ $X2=0.362 $Y2=0.94
r29 20 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.34
+ $Y=1.105 $X2=0.34 $Y2=1.105
r30 13 14 12.5413 $w=3.38e-07 $l=3.7e-07 $layer=LI1_cond $X=0.255 $Y=1.665
+ $X2=0.255 $Y2=2.035
r31 12 13 12.5413 $w=3.38e-07 $l=3.7e-07 $layer=LI1_cond $X=0.255 $Y=1.295
+ $X2=0.255 $Y2=1.665
r32 12 21 6.44012 $w=3.38e-07 $l=1.9e-07 $layer=LI1_cond $X=0.255 $Y=1.295
+ $X2=0.255 $Y2=1.105
r33 11 21 6.10117 $w=3.38e-07 $l=1.8e-07 $layer=LI1_cond $X=0.255 $Y=0.925
+ $X2=0.255 $Y2=1.105
r34 8 10 538.404 $w=1.5e-07 $l=1.05e-06 $layer=POLY_cond $X=0.475 $Y=2.66
+ $X2=0.475 $Y2=1.61
r35 5 22 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.475 $Y=0.62
+ $X2=0.475 $Y2=0.94
r36 2 10 48.4185 $w=3.75e-07 $l=1.87e-07 $layer=POLY_cond $X=0.362 $Y=1.423
+ $X2=0.362 $Y2=1.61
r37 1 20 3.26277 $w=3.75e-07 $l=2.2e-08 $layer=POLY_cond $X=0.362 $Y=1.127
+ $X2=0.362 $Y2=1.105
r38 1 2 43.8991 $w=3.75e-07 $l=2.96e-07 $layer=POLY_cond $X=0.362 $Y=1.127
+ $X2=0.362 $Y2=1.423
.ends

.subckt PM_SKY130_FD_SC_LP__DFXBP_1%D 3 7 12 15 16 17 18 23
c42 3 0 9.09583e-20 $X=2.125 $Y=2.525
r43 23 24 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.99
+ $Y=1.375 $X2=1.99 $Y2=1.375
r44 17 18 9.12472 $w=4.83e-07 $l=3.7e-07 $layer=LI1_cond $X=1.832 $Y=1.665
+ $X2=1.832 $Y2=2.035
r45 17 24 7.15181 $w=4.83e-07 $l=2.9e-07 $layer=LI1_cond $X=1.832 $Y=1.665
+ $X2=1.832 $Y2=1.375
r46 16 24 1.97291 $w=4.83e-07 $l=8e-08 $layer=LI1_cond $X=1.832 $Y=1.295
+ $X2=1.832 $Y2=1.375
r47 14 23 47.1618 $w=3.75e-07 $l=3.18e-07 $layer=POLY_cond $X=2.012 $Y=1.693
+ $X2=2.012 $Y2=1.375
r48 14 15 48.4185 $w=3.75e-07 $l=1.87e-07 $layer=POLY_cond $X=2.012 $Y=1.693
+ $X2=2.012 $Y2=1.88
r49 10 23 2.22462 $w=3.75e-07 $l=1.5e-08 $layer=POLY_cond $X=2.012 $Y=1.36
+ $X2=2.012 $Y2=1.375
r50 10 12 168.187 $w=1.5e-07 $l=3.28e-07 $layer=POLY_cond $X=2.012 $Y=1.285
+ $X2=2.34 $Y2=1.285
r51 5 12 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.34 $Y=1.21 $X2=2.34
+ $Y2=1.285
r52 5 7 207.67 $w=1.5e-07 $l=4.05e-07 $layer=POLY_cond $X=2.34 $Y=1.21 $X2=2.34
+ $Y2=0.805
r53 3 15 330.734 $w=1.5e-07 $l=6.45e-07 $layer=POLY_cond $X=2.125 $Y=2.525
+ $X2=2.125 $Y2=1.88
.ends

.subckt PM_SKY130_FD_SC_LP__DFXBP_1%A_217_463# 1 2 9 13 17 19 23 25 26 32 34 37
+ 38 39 41 43 44 47 49 54 56 58 59
c167 58 0 1.87194e-19 $X=5 $Y=1.39
c168 49 0 9.09583e-20 $X=1.21 $Y=2.46
r169 59 65 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=5 $Y=1.39 $X2=5
+ $Y2=1.48
r170 59 64 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5 $Y=1.39 $X2=5
+ $Y2=1.225
r171 58 61 9.07524 $w=2.28e-07 $l=1.65e-07 $layer=LI1_cond $X=4.98 $Y=1.39
+ $X2=4.98 $Y2=1.555
r172 58 59 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5 $Y=1.39
+ $X2=5 $Y2=1.39
r173 51 54 4.6541 $w=2.58e-07 $l=1.05e-07 $layer=LI1_cond $X=3.11 $Y=2.025
+ $X2=3.215 $Y2=2.025
r174 51 52 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.11
+ $Y=1.99 $X2=3.11 $Y2=1.99
r175 47 61 56.107 $w=1.68e-07 $l=8.6e-07 $layer=LI1_cond $X=4.95 $Y=2.415
+ $X2=4.95 $Y2=1.555
r176 45 56 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.3 $Y=2.5 $X2=3.215
+ $Y2=2.5
r177 44 47 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.865 $Y=2.5
+ $X2=4.95 $Y2=2.415
r178 44 45 102.102 $w=1.68e-07 $l=1.565e-06 $layer=LI1_cond $X=4.865 $Y=2.5
+ $X2=3.3 $Y2=2.5
r179 42 56 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.215 $Y=2.585
+ $X2=3.215 $Y2=2.5
r180 42 43 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=3.215 $Y=2.585
+ $X2=3.215 $Y2=2.865
r181 41 56 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.215 $Y=2.415
+ $X2=3.215 $Y2=2.5
r182 40 54 3.22376 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.215 $Y=2.155
+ $X2=3.215 $Y2=2.025
r183 40 41 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=3.215 $Y=2.155
+ $X2=3.215 $Y2=2.415
r184 38 43 6.91519 $w=2.1e-07 $l=1.41244e-07 $layer=LI1_cond $X=3.13 $Y=2.97
+ $X2=3.215 $Y2=2.865
r185 38 39 55.7186 $w=2.08e-07 $l=1.055e-06 $layer=LI1_cond $X=3.13 $Y=2.97
+ $X2=2.075 $Y2=2.97
r186 37 39 6.91519 $w=2.1e-07 $l=1.41244e-07 $layer=LI1_cond $X=1.99 $Y=2.865
+ $X2=2.075 $Y2=2.97
r187 36 37 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=1.99 $Y=2.485
+ $X2=1.99 $Y2=2.865
r188 35 49 2.68609 $w=1.7e-07 $l=1.92935e-07 $layer=LI1_cond $X=1.42 $Y=2.4
+ $X2=1.232 $Y2=2.39
r189 34 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.905 $Y=2.4
+ $X2=1.99 $Y2=2.485
r190 34 35 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=1.905 $Y=2.4
+ $X2=1.42 $Y2=2.4
r191 30 49 3.77418 $w=2.45e-07 $l=1.30038e-07 $layer=LI1_cond $X=1.315 $Y=2.295
+ $X2=1.232 $Y2=2.39
r192 30 32 78.6926 $w=2.08e-07 $l=1.49e-06 $layer=LI1_cond $X=1.315 $Y=2.295
+ $X2=1.315 $Y2=0.805
r193 26 52 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=3.125 $Y=1.99
+ $X2=3.11 $Y2=1.99
r194 25 52 83.9334 $w=3.3e-07 $l=4.8e-07 $layer=POLY_cond $X=2.63 $Y=1.99
+ $X2=3.11 $Y2=1.99
r195 21 27 10.146 $w=1.5e-07 $l=1.3e-07 $layer=POLY_cond $X=5.61 $Y=1.665
+ $X2=5.61 $Y2=1.535
r196 21 23 225.617 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=5.61 $Y=1.665
+ $X2=5.61 $Y2=2.105
r197 20 65 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.165 $Y=1.48
+ $X2=5 $Y2=1.48
r198 19 27 56.4625 $w=2.05e-07 $l=2.50998e-07 $layer=POLY_cond $X=5.385 $Y=1.48
+ $X2=5.61 $Y2=1.535
r199 19 20 112.809 $w=1.5e-07 $l=2.2e-07 $layer=POLY_cond $X=5.385 $Y=1.48
+ $X2=5.165 $Y2=1.48
r200 17 64 215.362 $w=1.5e-07 $l=4.2e-07 $layer=POLY_cond $X=4.91 $Y=0.805
+ $X2=4.91 $Y2=1.225
r201 11 26 32.1775 $w=3.3e-07 $l=1.98997e-07 $layer=POLY_cond $X=3.2 $Y=1.825
+ $X2=3.125 $Y2=1.99
r202 11 13 523.021 $w=1.5e-07 $l=1.02e-06 $layer=POLY_cond $X=3.2 $Y=1.825
+ $X2=3.2 $Y2=0.805
r203 7 25 32.1775 $w=3.3e-07 $l=1.98997e-07 $layer=POLY_cond $X=2.555 $Y=2.155
+ $X2=2.63 $Y2=1.99
r204 7 9 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=2.555 $Y=2.155
+ $X2=2.555 $Y2=2.525
r205 2 49 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=1.085
+ $Y=2.315 $X2=1.21 $Y2=2.46
r206 1 32 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=1.2
+ $Y=0.595 $X2=1.325 $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_LP__DFXBP_1%A_697_93# 1 2 7 9 12 18 21 23 27 29 36 41
c70 27 0 8.14738e-20 $X=4.6 $Y=0.75
r71 33 41 6.99445 $w=3.3e-07 $l=4e-08 $layer=POLY_cond $X=3.71 $Y=1.29 $X2=3.75
+ $Y2=1.29
r72 33 38 26.2292 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=3.71 $Y=1.29
+ $X2=3.56 $Y2=1.29
r73 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.71
+ $Y=1.29 $X2=3.71 $Y2=1.29
r74 29 32 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=3.71 $Y=1.17 $X2=3.71
+ $Y2=1.29
r75 25 27 19.555 $w=1.88e-07 $l=3.35e-07 $layer=LI1_cond $X=4.6 $Y=1.085 $X2=4.6
+ $Y2=0.75
r76 24 29 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.875 $Y=1.17
+ $X2=3.71 $Y2=1.17
r77 23 25 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=4.505 $Y=1.17
+ $X2=4.6 $Y2=1.085
r78 23 24 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=4.505 $Y=1.17
+ $X2=3.875 $Y2=1.17
r79 18 37 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.66 $Y=1.99
+ $X2=3.66 $Y2=2.155
r80 18 36 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.66 $Y=1.99
+ $X2=3.66 $Y2=1.825
r81 17 21 31.8617 $w=3.38e-07 $l=9.4e-07 $layer=LI1_cond $X=3.66 $Y=2.065
+ $X2=4.6 $Y2=2.065
r82 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.66
+ $Y=1.99 $X2=3.66 $Y2=1.99
r83 14 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.75 $Y=1.455
+ $X2=3.75 $Y2=1.29
r84 14 36 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=3.75 $Y=1.455
+ $X2=3.75 $Y2=1.825
r85 12 37 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=3.685 $Y=2.525
+ $X2=3.685 $Y2=2.155
r86 7 38 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.56 $Y=1.125
+ $X2=3.56 $Y2=1.29
r87 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=3.56 $Y=1.125 $X2=3.56
+ $Y2=0.805
r88 2 21 600 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_PDIFF $count=1 $X=4.46
+ $Y=1.895 $X2=4.6 $Y2=2.07
r89 1 27 91 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=2 $X=4.46
+ $Y=0.595 $X2=4.6 $Y2=0.75
.ends

.subckt PM_SKY130_FD_SC_LP__DFXBP_1%A_526_463# 1 2 9 13 16 19 22 29 32 33 34
c82 34 0 3.12341e-20 $X=4.13 $Y=1.575
c83 33 0 1.55547e-19 $X=4.295 $Y=1.57
c84 9 0 8.14738e-20 $X=4.385 $Y=0.915
r85 33 38 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.295 $Y=1.57
+ $X2=4.295 $Y2=1.735
r86 33 37 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.295 $Y=1.57
+ $X2=4.295 $Y2=1.405
r87 32 34 8.48463 $w=2.98e-07 $l=1.65e-07 $layer=LI1_cond $X=4.295 $Y=1.575
+ $X2=4.13 $Y2=1.575
r88 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.295
+ $Y=1.57 $X2=4.295 $Y2=1.57
r89 26 29 6.11144 $w=3.28e-07 $l=1.75e-07 $layer=LI1_cond $X=2.69 $Y=2.53
+ $X2=2.865 $Y2=2.53
r90 22 34 63.2834 $w=1.68e-07 $l=9.7e-07 $layer=LI1_cond $X=3.16 $Y=1.64
+ $X2=4.13 $Y2=1.64
r91 17 22 9.65561 $w=1.68e-07 $l=1.48e-07 $layer=LI1_cond $X=3.012 $Y=1.64
+ $X2=3.16 $Y2=1.64
r92 17 23 21.0075 $w=1.68e-07 $l=3.22e-07 $layer=LI1_cond $X=3.012 $Y=1.64
+ $X2=2.69 $Y2=1.64
r93 17 19 29.4947 $w=2.93e-07 $l=7.55e-07 $layer=LI1_cond $X=3.012 $Y=1.555
+ $X2=3.012 $Y2=0.8
r94 16 26 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.69 $Y=2.365
+ $X2=2.69 $Y2=2.53
r95 15 23 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.69 $Y=1.725
+ $X2=2.69 $Y2=1.64
r96 15 16 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=2.69 $Y=1.725
+ $X2=2.69 $Y2=2.365
r97 13 38 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=4.385 $Y=2.315
+ $X2=4.385 $Y2=1.735
r98 9 37 251.255 $w=1.5e-07 $l=4.9e-07 $layer=POLY_cond $X=4.385 $Y=0.915
+ $X2=4.385 $Y2=1.405
r99 2 29 600 $w=1.7e-07 $l=3.25192e-07 $layer=licon1_PDIFF $count=1 $X=2.63
+ $Y=2.315 $X2=2.865 $Y2=2.53
r100 1 19 182 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_NDIFF $count=1 $X=2.845
+ $Y=0.595 $X2=2.985 $Y2=0.8
.ends

.subckt PM_SKY130_FD_SC_LP__DFXBP_1%A_110_82# 1 2 7 8 12 16 17 18 19 20 23 25 29
+ 31 35 39 43 45 46 47 49 53 56 59 61 62 64
c138 56 0 4.113e-20 $X=0.817 $Y=1.663
r139 61 63 5.84975 $w=4.43e-07 $l=1.65e-07 $layer=LI1_cond $X=0.817 $Y=1.38
+ $X2=0.817 $Y2=1.215
r140 61 62 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.955
+ $Y=1.38 $X2=0.955 $Y2=1.38
r141 59 64 24.1227 $w=1.98e-07 $l=4.35e-07 $layer=LI1_cond $X=0.695 $Y=2.32
+ $X2=0.695 $Y2=1.885
r142 56 64 9.28731 $w=4.43e-07 $l=2.22e-07 $layer=LI1_cond $X=0.817 $Y=1.663
+ $X2=0.817 $Y2=1.885
r143 55 61 1.47616 $w=4.43e-07 $l=5.7e-08 $layer=LI1_cond $X=0.817 $Y=1.437
+ $X2=0.817 $Y2=1.38
r144 55 56 5.85286 $w=4.43e-07 $l=2.26e-07 $layer=LI1_cond $X=0.817 $Y=1.437
+ $X2=0.817 $Y2=1.663
r145 53 63 24.6952 $w=2.78e-07 $l=6e-07 $layer=LI1_cond $X=0.735 $Y=0.615
+ $X2=0.735 $Y2=1.215
r146 47 59 6.02628 $w=2.33e-07 $l=1.17e-07 $layer=LI1_cond $X=0.677 $Y=2.437
+ $X2=0.677 $Y2=2.32
r147 47 49 2.35393 $w=2.33e-07 $l=4.8e-08 $layer=LI1_cond $X=0.677 $Y=2.437
+ $X2=0.677 $Y2=2.485
r148 42 43 58.9681 $w=1.5e-07 $l=1.15e-07 $layer=POLY_cond $X=1.425 $Y=1.29
+ $X2=1.54 $Y2=1.29
r149 41 62 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=0.955 $Y=1.365
+ $X2=0.955 $Y2=1.38
r150 37 39 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=5.45 $Y=0.255
+ $X2=5.45 $Y2=0.805
r151 33 35 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=5.085 $Y=3.075
+ $X2=5.085 $Y2=2.315
r152 32 46 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.25 $Y=3.15
+ $X2=3.175 $Y2=3.15
r153 31 33 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.01 $Y=3.15
+ $X2=5.085 $Y2=3.075
r154 31 32 902.468 $w=1.5e-07 $l=1.76e-06 $layer=POLY_cond $X=5.01 $Y=3.15
+ $X2=3.25 $Y2=3.15
r155 27 46 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.175 $Y=3.075
+ $X2=3.175 $Y2=3.15
r156 27 29 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=3.175 $Y=3.075
+ $X2=3.175 $Y2=2.705
r157 26 45 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.845 $Y=0.18
+ $X2=2.77 $Y2=0.18
r158 25 37 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.375 $Y=0.18
+ $X2=5.45 $Y2=0.255
r159 25 26 1297.3 $w=1.5e-07 $l=2.53e-06 $layer=POLY_cond $X=5.375 $Y=0.18
+ $X2=2.845 $Y2=0.18
r160 21 45 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.77 $Y=0.255
+ $X2=2.77 $Y2=0.18
r161 21 23 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=2.77 $Y=0.255
+ $X2=2.77 $Y2=0.805
r162 19 45 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.695 $Y=0.18
+ $X2=2.77 $Y2=0.18
r163 19 20 553.787 $w=1.5e-07 $l=1.08e-06 $layer=POLY_cond $X=2.695 $Y=0.18
+ $X2=1.615 $Y2=0.18
r164 17 46 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.1 $Y=3.15
+ $X2=3.175 $Y2=3.15
r165 17 18 820.426 $w=1.5e-07 $l=1.6e-06 $layer=POLY_cond $X=3.1 $Y=3.15 $X2=1.5
+ $Y2=3.15
r166 14 43 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.54 $Y=1.215
+ $X2=1.54 $Y2=1.29
r167 14 16 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=1.54 $Y=1.215
+ $X2=1.54 $Y2=0.805
r168 13 20 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.54 $Y=0.255
+ $X2=1.615 $Y2=0.18
r169 13 16 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=1.54 $Y=0.255
+ $X2=1.54 $Y2=0.805
r170 10 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.425 $Y=3.075
+ $X2=1.5 $Y2=3.15
r171 10 12 225.617 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=1.425 $Y=3.075
+ $X2=1.425 $Y2=2.635
r172 9 42 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.425 $Y=1.365
+ $X2=1.425 $Y2=1.29
r173 9 12 651.213 $w=1.5e-07 $l=1.27e-06 $layer=POLY_cond $X=1.425 $Y=1.365
+ $X2=1.425 $Y2=2.635
r174 8 41 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=1.12 $Y=1.29
+ $X2=0.955 $Y2=1.365
r175 7 42 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.35 $Y=1.29
+ $X2=1.425 $Y2=1.29
r176 7 8 117.936 $w=1.5e-07 $l=2.3e-07 $layer=POLY_cond $X=1.35 $Y=1.29 $X2=1.12
+ $Y2=1.29
r177 2 49 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=0.55
+ $Y=2.34 $X2=0.69 $Y2=2.485
r178 1 53 182 $w=1.7e-07 $l=2.73542e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.41 $X2=0.71 $Y2=0.615
.ends

.subckt PM_SKY130_FD_SC_LP__DFXBP_1%A_1149_93# 1 2 7 9 10 12 14 16 19 21 23 26
+ 28 29 30 35 36 37 38 39 42 46 54 63
c122 28 0 1.16669e-19 $X=7.545 $Y=1.485
c123 19 0 6.36774e-20 $X=7.64 $Y=2.155
c124 10 0 3.16466e-20 $X=5.97 $Y=1.735
r125 56 57 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.17
+ $Y=1.485 $X2=7.17 $Y2=1.485
r126 54 56 8.91694 $w=3.01e-07 $l=2.2e-07 $layer=LI1_cond $X=6.95 $Y=1.562
+ $X2=7.17 $Y2=1.562
r127 46 49 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=6.06 $Y=1.57
+ $X2=6.06 $Y2=1.72
r128 46 47 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.06
+ $Y=1.57 $X2=6.06 $Y2=1.57
r129 43 63 41.9667 $w=3.3e-07 $l=2.4e-07 $layer=POLY_cond $X=8.885 $Y=1.51
+ $X2=9.125 $Y2=1.51
r130 42 43 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.885
+ $Y=1.51 $X2=8.885 $Y2=1.51
r131 40 42 30.208 $w=3.28e-07 $l=8.65e-07 $layer=LI1_cond $X=8.885 $Y=2.375
+ $X2=8.885 $Y2=1.51
r132 38 40 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=8.72 $Y=2.46
+ $X2=8.885 $Y2=2.375
r133 38 39 109.93 $w=1.68e-07 $l=1.685e-06 $layer=LI1_cond $X=8.72 $Y=2.46
+ $X2=7.035 $Y2=2.46
r134 37 54 4.08057 $w=1.7e-07 $l=2.42e-07 $layer=LI1_cond $X=6.95 $Y=1.32
+ $X2=6.95 $Y2=1.562
r135 36 52 17.6853 $w=3.83e-07 $l=5.07893e-07 $layer=LI1_cond $X=6.95 $Y=0.955
+ $X2=6.792 $Y2=0.52
r136 36 37 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=6.95 $Y=0.955
+ $X2=6.95 $Y2=1.32
r137 33 39 13.1494 $w=2.1e-07 $l=2.6714e-07 $layer=LI1_cond $X=6.807 $Y=2.375
+ $X2=7.035 $Y2=2.46
r138 33 35 8.80629 $w=4.53e-07 $l=3.35e-07 $layer=LI1_cond $X=6.807 $Y=2.375
+ $X2=6.807 $Y2=2.04
r139 32 54 5.79601 $w=3.01e-07 $l=3.06265e-07 $layer=LI1_cond $X=6.807 $Y=1.805
+ $X2=6.95 $Y2=1.562
r140 32 35 6.17755 $w=4.53e-07 $l=2.35e-07 $layer=LI1_cond $X=6.807 $Y=1.805
+ $X2=6.807 $Y2=2.04
r141 31 49 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.225 $Y=1.72
+ $X2=6.06 $Y2=1.72
r142 30 32 11.4926 $w=3.01e-07 $l=2.66128e-07 $layer=LI1_cond $X=6.58 $Y=1.72
+ $X2=6.807 $Y2=1.805
r143 30 31 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=6.58 $Y=1.72
+ $X2=6.225 $Y2=1.72
r144 28 57 65.573 $w=3.3e-07 $l=3.75e-07 $layer=POLY_cond $X=7.545 $Y=1.485
+ $X2=7.17 $Y2=1.485
r145 28 29 5.03009 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.545 $Y=1.485
+ $X2=7.545 $Y2=1.32
r146 24 63 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.125 $Y=1.675
+ $X2=9.125 $Y2=1.51
r147 24 26 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=9.125 $Y=1.675
+ $X2=9.125 $Y2=2.465
r148 21 63 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.125 $Y=1.345
+ $X2=9.125 $Y2=1.51
r149 21 23 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=9.125 $Y=1.345
+ $X2=9.125 $Y2=0.815
r150 17 29 37.0704 $w=1.5e-07 $l=3.745e-07 $layer=POLY_cond $X=7.64 $Y=1.65
+ $X2=7.545 $Y2=1.32
r151 17 19 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=7.64 $Y=1.65
+ $X2=7.64 $Y2=2.155
r152 14 29 37.0704 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.62 $Y=1.32
+ $X2=7.545 $Y2=1.32
r153 14 16 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=7.62 $Y=1.32
+ $X2=7.62 $Y2=1
r154 10 47 38.561 $w=2.98e-07 $l=1.72337e-07 $layer=POLY_cond $X=5.97 $Y=1.735
+ $X2=5.985 $Y2=1.57
r155 10 12 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=5.97 $Y=1.735
+ $X2=5.97 $Y2=2.105
r156 7 47 83.8496 $w=2.98e-07 $l=5.21009e-07 $layer=POLY_cond $X=5.82 $Y=1.125
+ $X2=5.985 $Y2=1.57
r157 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=5.82 $Y=1.125
+ $X2=5.82 $Y2=0.805
r158 2 35 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=6.585
+ $Y=1.895 $X2=6.725 $Y2=2.04
r159 1 52 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.585
+ $Y=0.375 $X2=6.725 $Y2=0.52
.ends

.subckt PM_SKY130_FD_SC_LP__DFXBP_1%A_997_119# 1 2 9 12 14 16 20 22 27 28 32 35
c72 28 0 1.16669e-19 $X=6.56 $Y=1.21
r73 32 36 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.6 $Y=1.29 $X2=6.6
+ $Y2=1.455
r74 32 35 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.6 $Y=1.29 $X2=6.6
+ $Y2=1.125
r75 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.6
+ $Y=1.29 $X2=6.6 $Y2=1.29
r76 28 31 3.68782 $w=2.48e-07 $l=8e-08 $layer=LI1_cond $X=6.56 $Y=1.21 $X2=6.56
+ $Y2=1.29
r77 23 25 15.6857 $w=3.15e-07 $l=5.06325e-07 $layer=LI1_cond $X=5.465 $Y=1.21
+ $X2=5.237 $Y2=0.805
r78 22 28 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.435 $Y=1.21
+ $X2=6.56 $Y2=1.21
r79 22 23 63.2834 $w=1.68e-07 $l=9.7e-07 $layer=LI1_cond $X=6.435 $Y=1.21
+ $X2=5.465 $Y2=1.21
r80 20 23 4.91151 $w=3.15e-07 $l=1.36015e-07 $layer=LI1_cond $X=5.365 $Y=1.295
+ $X2=5.465 $Y2=1.21
r81 20 27 32.1636 $w=1.98e-07 $l=5.8e-07 $layer=LI1_cond $X=5.365 $Y=1.295
+ $X2=5.365 $Y2=1.875
r82 16 18 24.157 $w=2.58e-07 $l=5.45e-07 $layer=LI1_cond $X=5.335 $Y=2.04
+ $X2=5.335 $Y2=2.585
r83 14 27 6.4054 $w=2.58e-07 $l=1.3e-07 $layer=LI1_cond $X=5.335 $Y=2.005
+ $X2=5.335 $Y2=1.875
r84 14 16 1.55137 $w=2.58e-07 $l=3.5e-08 $layer=LI1_cond $X=5.335 $Y=2.005
+ $X2=5.335 $Y2=2.04
r85 12 36 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=6.51 $Y=2.315
+ $X2=6.51 $Y2=1.455
r86 9 35 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=6.51 $Y=0.695
+ $X2=6.51 $Y2=1.125
r87 2 18 600 $w=1.7e-07 $l=7.56769e-07 $layer=licon1_PDIFF $count=1 $X=5.16
+ $Y=1.895 $X2=5.3 $Y2=2.585
r88 2 16 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=5.16
+ $Y=1.895 $X2=5.3 $Y2=2.04
r89 1 25 182 $w=1.7e-07 $l=2.89828e-07 $layer=licon1_NDIFF $count=1 $X=4.985
+ $Y=0.595 $X2=5.175 $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_LP__DFXBP_1%A_1401_22# 1 2 7 8 11 13 17 19 22 24 30 35
r64 33 35 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=7.425 $Y=2.04
+ $X2=7.52 $Y2=2.04
r65 29 30 6.07359 $w=2.08e-07 $l=1.15e-07 $layer=LI1_cond $X=7.405 $Y=0.935
+ $X2=7.52 $Y2=0.935
r66 26 29 5.54545 $w=2.08e-07 $l=1.05e-07 $layer=LI1_cond $X=7.3 $Y=0.935
+ $X2=7.405 $Y2=0.935
r67 21 24 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=7.17 $Y=0.43 $X2=7.3
+ $Y2=0.43
r68 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.17
+ $Y=0.43 $X2=7.17 $Y2=0.43
r69 19 35 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.52 $Y=1.875
+ $X2=7.52 $Y2=2.04
r70 18 30 1.9771 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=7.52 $Y=1.04 $X2=7.52
+ $Y2=0.935
r71 18 19 54.4759 $w=1.68e-07 $l=8.35e-07 $layer=LI1_cond $X=7.52 $Y=1.04
+ $X2=7.52 $Y2=1.875
r72 17 26 1.9771 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=7.3 $Y=0.83 $X2=7.3
+ $Y2=0.935
r73 16 24 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.3 $Y=0.595 $X2=7.3
+ $Y2=0.43
r74 16 17 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=7.3 $Y=0.595
+ $X2=7.3 $Y2=0.83
r75 15 22 29.7264 $w=3.3e-07 $l=1.7e-07 $layer=POLY_cond $X=7.17 $Y=0.26
+ $X2=7.17 $Y2=0.43
r76 11 13 858.883 $w=1.5e-07 $l=1.675e-06 $layer=POLY_cond $X=8.165 $Y=0.79
+ $X2=8.165 $Y2=2.465
r77 9 11 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=8.165 $Y=0.26
+ $X2=8.165 $Y2=0.79
r78 8 15 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=7.335 $Y=0.185
+ $X2=7.17 $Y2=0.26
r79 7 9 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.09 $Y=0.185
+ $X2=8.165 $Y2=0.26
r80 7 8 387.138 $w=1.5e-07 $l=7.55e-07 $layer=POLY_cond $X=8.09 $Y=0.185
+ $X2=7.335 $Y2=0.185
r81 2 33 600 $w=1.7e-07 $l=2.60096e-07 $layer=licon1_PDIFF $count=1 $X=7.3
+ $Y=1.835 $X2=7.425 $Y2=2.04
r82 1 29 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=7.28
+ $Y=0.79 $X2=7.405 $Y2=0.935
.ends

.subckt PM_SKY130_FD_SC_LP__DFXBP_1%VPWR 1 2 3 4 5 6 19 21 25 29 33 39 41 45 48
+ 49 50 52 57 69 78 79 85 88 91 94
r98 94 95 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r99 92 95 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=8.88 $Y2=3.33
r100 91 92 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r101 88 89 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r102 85 86 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r103 82 83 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r104 79 95 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=8.88 $Y2=3.33
r105 78 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r106 76 94 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=9.015 $Y=3.33
+ $X2=8.91 $Y2=3.33
r107 76 78 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=9.015 $Y=3.33
+ $X2=9.36 $Y2=3.33
r108 75 92 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=7.92 $Y2=3.33
r109 74 75 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r110 72 75 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=7.44 $Y2=3.33
r111 71 74 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=6.48 $Y=3.33
+ $X2=7.44 $Y2=3.33
r112 71 72 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r113 69 91 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.785 $Y=3.33
+ $X2=7.95 $Y2=3.33
r114 69 74 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=7.785 $Y=3.33
+ $X2=7.44 $Y2=3.33
r115 68 72 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=6.48
+ $Y2=3.33
r116 67 68 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r117 65 89 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=4.08 $Y2=3.33
r118 64 67 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=4.56 $Y=3.33 $X2=6
+ $Y2=3.33
r119 64 65 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r120 62 88 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.275 $Y=3.33
+ $X2=4.11 $Y2=3.33
r121 62 64 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=4.275 $Y=3.33
+ $X2=4.56 $Y2=3.33
r122 61 89 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r123 61 86 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=1.68 $Y2=3.33
r124 60 61 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r125 58 85 6.81202 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=1.735 $Y=3.33
+ $X2=1.615 $Y2=3.33
r126 58 60 121.674 $w=1.68e-07 $l=1.865e-06 $layer=LI1_cond $X=1.735 $Y=3.33
+ $X2=3.6 $Y2=3.33
r127 57 88 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.945 $Y=3.33
+ $X2=4.11 $Y2=3.33
r128 57 60 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=3.945 $Y=3.33
+ $X2=3.6 $Y2=3.33
r129 56 86 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r130 56 83 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.24 $Y2=3.33
r131 55 56 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r132 53 82 4.45907 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=0.39 $Y=3.33
+ $X2=0.195 $Y2=3.33
r133 53 55 52.8449 $w=1.68e-07 $l=8.1e-07 $layer=LI1_cond $X=0.39 $Y=3.33
+ $X2=1.2 $Y2=3.33
r134 52 85 6.81202 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=1.495 $Y=3.33
+ $X2=1.615 $Y2=3.33
r135 52 55 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.495 $Y=3.33
+ $X2=1.2 $Y2=3.33
r136 50 68 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=4.8 $Y=3.33 $X2=6
+ $Y2=3.33
r137 50 65 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.8 $Y=3.33
+ $X2=4.56 $Y2=3.33
r138 48 67 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=6.08 $Y=3.33 $X2=6
+ $Y2=3.33
r139 48 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.08 $Y=3.33
+ $X2=6.245 $Y2=3.33
r140 47 71 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=6.41 $Y=3.33 $X2=6.48
+ $Y2=3.33
r141 47 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.41 $Y=3.33
+ $X2=6.245 $Y2=3.33
r142 43 94 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=8.91 $Y=3.245
+ $X2=8.91 $Y2=3.33
r143 43 45 15.5801 $w=2.08e-07 $l=2.95e-07 $layer=LI1_cond $X=8.91 $Y=3.245
+ $X2=8.91 $Y2=2.95
r144 42 91 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.115 $Y=3.33
+ $X2=7.95 $Y2=3.33
r145 41 94 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=8.805 $Y=3.33
+ $X2=8.91 $Y2=3.33
r146 41 42 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=8.805 $Y=3.33
+ $X2=8.115 $Y2=3.33
r147 37 91 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.95 $Y=3.245
+ $X2=7.95 $Y2=3.33
r148 37 39 14.1436 $w=3.28e-07 $l=4.05e-07 $layer=LI1_cond $X=7.95 $Y=3.245
+ $X2=7.95 $Y2=2.84
r149 33 36 18.3343 $w=3.28e-07 $l=5.25e-07 $layer=LI1_cond $X=6.245 $Y=2.065
+ $X2=6.245 $Y2=2.59
r150 31 49 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.245 $Y=3.245
+ $X2=6.245 $Y2=3.33
r151 31 36 22.8742 $w=3.28e-07 $l=6.55e-07 $layer=LI1_cond $X=6.245 $Y=3.245
+ $X2=6.245 $Y2=2.59
r152 27 88 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.11 $Y=3.245
+ $X2=4.11 $Y2=3.33
r153 27 29 13.7944 $w=3.28e-07 $l=3.95e-07 $layer=LI1_cond $X=4.11 $Y=3.245
+ $X2=4.11 $Y2=2.85
r154 23 85 0.135687 $w=2.4e-07 $l=8.5e-08 $layer=LI1_cond $X=1.615 $Y=3.245
+ $X2=1.615 $Y2=3.33
r155 23 25 20.4078 $w=2.38e-07 $l=4.25e-07 $layer=LI1_cond $X=1.615 $Y=3.245
+ $X2=1.615 $Y2=2.82
r156 19 82 3.01845 $w=2.95e-07 $l=1.05924e-07 $layer=LI1_cond $X=0.242 $Y=3.245
+ $X2=0.195 $Y2=3.33
r157 19 21 29.6901 $w=2.93e-07 $l=7.6e-07 $layer=LI1_cond $X=0.242 $Y=3.245
+ $X2=0.242 $Y2=2.485
r158 6 45 600 $w=1.7e-07 $l=1.17584e-06 $layer=licon1_PDIFF $count=1 $X=8.785
+ $Y=1.835 $X2=8.91 $Y2=2.95
r159 5 39 600 $w=1.7e-07 $l=1.11633e-06 $layer=licon1_PDIFF $count=1 $X=7.715
+ $Y=1.835 $X2=7.95 $Y2=2.84
r160 4 36 600 $w=1.7e-07 $l=8.10417e-07 $layer=licon1_PDIFF $count=1 $X=6.045
+ $Y=1.895 $X2=6.295 $Y2=2.59
r161 4 33 600 $w=1.7e-07 $l=2.72029e-07 $layer=licon1_PDIFF $count=1 $X=6.045
+ $Y=1.895 $X2=6.245 $Y2=2.065
r162 3 29 600 $w=1.7e-07 $l=6.88095e-07 $layer=licon1_PDIFF $count=1 $X=3.76
+ $Y=2.315 $X2=4.11 $Y2=2.85
r163 2 25 600 $w=1.7e-07 $l=5.70723e-07 $layer=licon1_PDIFF $count=1 $X=1.5
+ $Y=2.315 $X2=1.64 $Y2=2.82
r164 1 21 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.34 $X2=0.26 $Y2=2.485
.ends

.subckt PM_SKY130_FD_SC_LP__DFXBP_1%A_440_463# 1 2 9 14
r19 11 14 7.50834 $w=3.28e-07 $l=2.15e-07 $layer=LI1_cond $X=2.34 $Y=0.8
+ $X2=2.555 $Y2=0.8
r20 7 11 3.96751 $w=1.9e-07 $l=1.65e-07 $layer=LI1_cond $X=2.34 $Y=0.965
+ $X2=2.34 $Y2=0.8
r21 7 9 91.3541 $w=1.88e-07 $l=1.565e-06 $layer=LI1_cond $X=2.34 $Y=0.965
+ $X2=2.34 $Y2=2.53
r22 2 9 600 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_PDIFF $count=1 $X=2.2
+ $Y=2.315 $X2=2.34 $Y2=2.53
r23 1 14 182 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_NDIFF $count=1 $X=2.415
+ $Y=0.595 $X2=2.555 $Y2=0.8
.ends

.subckt PM_SKY130_FD_SC_LP__DFXBP_1%Q_N 1 2 7 8 9 10 16
r14 9 10 14.7036 $w=2.88e-07 $l=3.7e-07 $layer=LI1_cond $X=8.4 $Y=1.665 $X2=8.4
+ $Y2=2.035
r15 8 9 14.7036 $w=2.88e-07 $l=3.7e-07 $layer=LI1_cond $X=8.4 $Y=1.295 $X2=8.4
+ $Y2=1.665
r16 7 8 14.7036 $w=2.88e-07 $l=3.7e-07 $layer=LI1_cond $X=8.4 $Y=0.925 $X2=8.4
+ $Y2=1.295
r17 7 16 16.0945 $w=2.88e-07 $l=4.05e-07 $layer=LI1_cond $X=8.4 $Y=0.925 $X2=8.4
+ $Y2=0.52
r18 2 10 600 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=1 $X=8.24
+ $Y=1.835 $X2=8.38 $Y2=2.04
r19 1 16 91 $w=1.7e-07 $l=2.08567e-07 $layer=licon1_NDIFF $count=2 $X=8.24
+ $Y=0.37 $X2=8.38 $Y2=0.52
.ends

.subckt PM_SKY130_FD_SC_LP__DFXBP_1%Q 1 2 7 8 9 10 11 12 13
r10 13 39 5.76222 $w=2.68e-07 $l=1.35e-07 $layer=LI1_cond $X=9.37 $Y=2.775
+ $X2=9.37 $Y2=2.91
r11 12 13 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=9.37 $Y=2.405
+ $X2=9.37 $Y2=2.775
r12 11 12 18.1403 $w=2.68e-07 $l=4.25e-07 $layer=LI1_cond $X=9.37 $Y=1.98
+ $X2=9.37 $Y2=2.405
r13 10 11 13.4452 $w=2.68e-07 $l=3.15e-07 $layer=LI1_cond $X=9.37 $Y=1.665
+ $X2=9.37 $Y2=1.98
r14 9 10 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=9.37 $Y=1.295
+ $X2=9.37 $Y2=1.665
r15 8 9 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=9.37 $Y=0.925 $X2=9.37
+ $Y2=1.295
r16 7 8 16.433 $w=2.68e-07 $l=3.85e-07 $layer=LI1_cond $X=9.37 $Y=0.54 $X2=9.37
+ $Y2=0.925
r17 2 39 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=9.2
+ $Y=1.835 $X2=9.34 $Y2=2.91
r18 2 11 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=9.2
+ $Y=1.835 $X2=9.34 $Y2=1.98
r19 1 7 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=9.2
+ $Y=0.395 $X2=9.34 $Y2=0.54
.ends

.subckt PM_SKY130_FD_SC_LP__DFXBP_1%VGND 1 2 3 4 5 6 19 21 25 29 33 37 43 46 47
+ 49 50 51 60 74 81 88 89 95 98 101
c109 29 0 3.12341e-20 $X=4.17 $Y=0.785
r110 101 102 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=0
+ $X2=8.88 $Y2=0
r111 98 99 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r112 95 96 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r113 92 93 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r114 89 102 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=0
+ $X2=8.88 $Y2=0
r115 88 89 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=0 $X2=9.36
+ $Y2=0
r116 86 101 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=9.015 $Y=0
+ $X2=8.88 $Y2=0
r117 86 88 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=9.015 $Y=0 $X2=9.36
+ $Y2=0
r118 85 102 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=0 $X2=8.88
+ $Y2=0
r119 85 99 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=0 $X2=7.92
+ $Y2=0
r120 84 85 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r121 82 98 8.23795 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=8.085 $Y=0 $X2=7.93
+ $Y2=0
r122 82 84 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=8.085 $Y=0 $X2=8.4
+ $Y2=0
r123 81 101 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=8.745 $Y=0
+ $X2=8.88 $Y2=0
r124 81 84 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=8.745 $Y=0 $X2=8.4
+ $Y2=0
r125 80 99 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0 $X2=7.92
+ $Y2=0
r126 79 80 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r127 77 80 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=7.44
+ $Y2=0
r128 76 79 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=6.48 $Y=0 $X2=7.44
+ $Y2=0
r129 76 77 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r130 74 98 8.23795 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=7.775 $Y=0 $X2=7.93
+ $Y2=0
r131 74 79 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=7.775 $Y=0
+ $X2=7.44 $Y2=0
r132 73 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.48
+ $Y2=0
r133 72 73 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=0 $X2=6 $Y2=0
r134 70 96 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=4.08
+ $Y2=0
r135 69 72 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=4.56 $Y=0 $X2=6
+ $Y2=0
r136 69 70 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r137 67 95 13.9156 $w=1.7e-07 $l=3.63e-07 $layer=LI1_cond $X=4.335 $Y=0
+ $X2=3.972 $Y2=0
r138 67 69 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=4.335 $Y=0
+ $X2=4.56 $Y2=0
r139 66 96 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r140 65 66 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r141 63 66 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.6
+ $Y2=0
r142 62 65 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=2.16 $Y=0 $X2=3.6
+ $Y2=0
r143 62 63 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r144 60 95 13.9156 $w=1.7e-07 $l=3.62e-07 $layer=LI1_cond $X=3.61 $Y=0 $X2=3.972
+ $Y2=0
r145 60 65 0.652406 $w=1.68e-07 $l=1e-08 $layer=LI1_cond $X=3.61 $Y=0 $X2=3.6
+ $Y2=0
r146 59 63 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r147 58 59 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r148 56 59 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r149 56 93 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r150 55 58 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r151 55 56 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r152 53 92 4.78091 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=0
+ $X2=0.212 $Y2=0
r153 53 55 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.425 $Y=0 $X2=0.72
+ $Y2=0
r154 51 73 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=4.8 $Y=0 $X2=6
+ $Y2=0
r155 51 70 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.8 $Y=0 $X2=4.56
+ $Y2=0
r156 49 72 3.26203 $w=1.68e-07 $l=5e-08 $layer=LI1_cond $X=6.05 $Y=0 $X2=6 $Y2=0
r157 49 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.05 $Y=0 $X2=6.215
+ $Y2=0
r158 48 76 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=6.38 $Y=0 $X2=6.48
+ $Y2=0
r159 48 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.38 $Y=0 $X2=6.215
+ $Y2=0
r160 46 58 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=1.755 $Y=0 $X2=1.68
+ $Y2=0
r161 46 47 8.42608 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=1.755 $Y=0 $X2=1.915
+ $Y2=0
r162 45 62 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=2.075 $Y=0 $X2=2.16
+ $Y2=0
r163 45 47 8.42608 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=2.075 $Y=0 $X2=1.915
+ $Y2=0
r164 41 101 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.88 $Y=0.085
+ $X2=8.88 $Y2=0
r165 41 43 19.4208 $w=2.68e-07 $l=4.55e-07 $layer=LI1_cond $X=8.88 $Y=0.085
+ $X2=8.88 $Y2=0.54
r166 37 39 21.1901 $w=3.08e-07 $l=5.7e-07 $layer=LI1_cond $X=7.93 $Y=0.495
+ $X2=7.93 $Y2=1.065
r167 35 98 0.701276 $w=3.1e-07 $l=8.5e-08 $layer=LI1_cond $X=7.93 $Y=0.085
+ $X2=7.93 $Y2=0
r168 35 37 15.242 $w=3.08e-07 $l=4.1e-07 $layer=LI1_cond $X=7.93 $Y=0.085
+ $X2=7.93 $Y2=0.495
r169 31 50 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.215 $Y=0.085
+ $X2=6.215 $Y2=0
r170 31 33 15.1913 $w=3.28e-07 $l=4.35e-07 $layer=LI1_cond $X=6.215 $Y=0.085
+ $X2=6.215 $Y2=0.52
r171 27 95 2.93543 $w=7.25e-07 $l=8.5e-08 $layer=LI1_cond $X=3.972 $Y=0.085
+ $X2=3.972 $Y2=0
r172 27 29 11.5483 $w=7.23e-07 $l=7e-07 $layer=LI1_cond $X=3.972 $Y=0.085
+ $X2=3.972 $Y2=0.785
r173 23 47 0.800721 $w=3.2e-07 $l=8.5e-08 $layer=LI1_cond $X=1.915 $Y=0.085
+ $X2=1.915 $Y2=0
r174 23 25 26.11 $w=3.18e-07 $l=7.25e-07 $layer=LI1_cond $X=1.915 $Y=0.085
+ $X2=1.915 $Y2=0.81
r175 19 92 2.98526 $w=3.3e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.212 $Y2=0
r176 19 21 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.26 $Y2=0.565
r177 6 43 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=8.785
+ $Y=0.395 $X2=8.91 $Y2=0.54
r178 5 39 182 $w=1.7e-07 $l=3.67083e-07 $layer=licon1_NDIFF $count=1 $X=7.695
+ $Y=0.79 $X2=7.91 $Y2=1.065
r179 5 37 182 $w=1.7e-07 $l=4.02803e-07 $layer=licon1_NDIFF $count=1 $X=7.695
+ $Y=0.79 $X2=7.95 $Y2=0.495
r180 4 33 91 $w=1.7e-07 $l=3.55528e-07 $layer=licon1_NDIFF $count=2 $X=5.895
+ $Y=0.595 $X2=6.215 $Y2=0.52
r181 3 29 91 $w=1.7e-07 $l=6.22796e-07 $layer=licon1_NDIFF $count=2 $X=3.635
+ $Y=0.595 $X2=4.17 $Y2=0.785
r182 2 25 182 $w=1.7e-07 $l=3.98246e-07 $layer=licon1_NDIFF $count=1 $X=1.615
+ $Y=0.595 $X2=1.92 $Y2=0.81
r183 1 21 182 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.41 $X2=0.26 $Y2=0.565
.ends

