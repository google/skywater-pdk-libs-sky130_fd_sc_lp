* File: sky130_fd_sc_lp__nor2_m.pxi.spice
* Created: Fri Aug 28 10:54:16 2020
* 
x_PM_SKY130_FD_SC_LP__NOR2_M%A N_A_c_29_n N_A_M1003_g N_A_M1001_g N_A_c_31_n A A
+ A A N_A_c_33_n N_A_c_34_n PM_SKY130_FD_SC_LP__NOR2_M%A
x_PM_SKY130_FD_SC_LP__NOR2_M%B N_B_M1002_g N_B_M1000_g B B B B N_B_c_56_n
+ N_B_c_57_n PM_SKY130_FD_SC_LP__NOR2_M%B
x_PM_SKY130_FD_SC_LP__NOR2_M%VPWR N_VPWR_M1001_s N_VPWR_c_80_n N_VPWR_c_81_n
+ VPWR N_VPWR_c_82_n N_VPWR_c_79_n PM_SKY130_FD_SC_LP__NOR2_M%VPWR
x_PM_SKY130_FD_SC_LP__NOR2_M%Y N_Y_M1003_d N_Y_M1002_d Y Y Y Y Y N_Y_c_94_n
+ N_Y_c_96_n PM_SKY130_FD_SC_LP__NOR2_M%Y
x_PM_SKY130_FD_SC_LP__NOR2_M%VGND N_VGND_M1003_s N_VGND_M1000_d N_VGND_c_113_n
+ N_VGND_c_114_n N_VGND_c_115_n N_VGND_c_116_n VGND N_VGND_c_117_n
+ N_VGND_c_118_n PM_SKY130_FD_SC_LP__NOR2_M%VGND
cc_1 VNB N_A_c_29_n 0.0241981f $X=-0.19 $Y=-0.245 $X2=0.402 $Y2=1.353
cc_2 VNB N_A_M1001_g 0.00643673f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=2.625
cc_3 VNB N_A_c_31_n 0.0243911f $X=-0.19 $Y=-0.245 $X2=0.402 $Y2=1.55
cc_4 VNB A 0.0336651f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_5 VNB N_A_c_33_n 0.0243625f $X=-0.19 $Y=-0.245 $X2=0.37 $Y2=1.045
cc_6 VNB N_A_c_34_n 0.0207887f $X=-0.19 $Y=-0.245 $X2=0.402 $Y2=0.88
cc_7 VNB N_B_M1002_g 0.00510295f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=0.88
cc_8 VNB B 0.00788317f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=2.625
cc_9 VNB N_B_c_56_n 0.103364f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_B_c_57_n 0.0197697f $X=-0.19 $Y=-0.245 $X2=0.402 $Y2=1.045
cc_11 VNB N_VPWR_c_79_n 0.0641695f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_12 VNB N_Y_c_94_n 0.00844517f $X=-0.19 $Y=-0.245 $X2=0.402 $Y2=0.88
cc_13 VNB N_VGND_c_113_n 0.0127795f $X=-0.19 $Y=-0.245 $X2=0.525 $Y2=2.625
cc_14 VNB N_VGND_c_114_n 0.0100635f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_VGND_c_115_n 0.0115035f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_16 VNB N_VGND_c_116_n 0.0100561f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_17 VNB N_VGND_c_117_n 0.0185872f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_VGND_c_118_n 0.116382f $X=-0.19 $Y=-0.245 $X2=0.305 $Y2=1.295
cc_19 VPB N_A_M1001_g 0.0635505f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=2.625
cc_20 VPB A 0.0246537f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_21 VPB N_B_M1002_g 0.0587023f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=0.88
cc_22 VPB B 0.0256898f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=2.625
cc_23 VPB N_VPWR_c_80_n 0.0127536f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=0.56
cc_24 VPB N_VPWR_c_81_n 0.0242582f $X=-0.19 $Y=1.655 $X2=0.525 $Y2=1.55
cc_25 VPB N_VPWR_c_82_n 0.0311146f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_26 VPB N_VPWR_c_79_n 0.0637672f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_27 VPB N_Y_c_94_n 0.00600257f $X=-0.19 $Y=1.655 $X2=0.402 $Y2=0.88
cc_28 VPB N_Y_c_96_n 0.0117477f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_29 N_A_c_31_n N_B_M1002_g 0.0524855f $X=0.402 $Y=1.55 $X2=0 $Y2=0
cc_30 A N_B_c_56_n 8.98218e-19 $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_31 N_A_c_33_n N_B_c_56_n 0.0524855f $X=0.37 $Y=1.045 $X2=0 $Y2=0
cc_32 N_A_c_34_n N_B_c_57_n 0.0131374f $X=0.402 $Y=0.88 $X2=0 $Y2=0
cc_33 N_A_M1001_g N_VPWR_c_81_n 0.00567057f $X=0.525 $Y=2.625 $X2=0 $Y2=0
cc_34 A N_VPWR_c_81_n 0.0135673f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_35 N_A_M1001_g N_VPWR_c_82_n 0.00490845f $X=0.525 $Y=2.625 $X2=0 $Y2=0
cc_36 N_A_M1001_g N_VPWR_c_79_n 0.00506877f $X=0.525 $Y=2.625 $X2=0 $Y2=0
cc_37 A N_Y_c_94_n 0.0941117f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_38 N_A_c_34_n N_Y_c_94_n 0.0192172f $X=0.402 $Y=0.88 $X2=0 $Y2=0
cc_39 N_A_M1001_g N_Y_c_96_n 0.00220013f $X=0.525 $Y=2.625 $X2=0 $Y2=0
cc_40 A N_VGND_c_114_n 0.0168964f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_41 N_A_c_33_n N_VGND_c_114_n 0.00139532f $X=0.37 $Y=1.045 $X2=0 $Y2=0
cc_42 N_A_c_34_n N_VGND_c_114_n 0.00355398f $X=0.402 $Y=0.88 $X2=0 $Y2=0
cc_43 N_A_c_34_n N_VGND_c_117_n 0.00478016f $X=0.402 $Y=0.88 $X2=0 $Y2=0
cc_44 A N_VGND_c_118_n 0.00429626f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_45 N_A_c_34_n N_VGND_c_118_n 0.00939134f $X=0.402 $Y=0.88 $X2=0 $Y2=0
cc_46 N_B_M1002_g N_VPWR_c_82_n 0.00363612f $X=0.915 $Y=2.625 $X2=0 $Y2=0
cc_47 N_B_M1002_g N_VPWR_c_79_n 0.00506877f $X=0.915 $Y=2.625 $X2=0 $Y2=0
cc_48 N_B_M1002_g N_Y_c_94_n 0.0257793f $X=0.915 $Y=2.625 $X2=0 $Y2=0
cc_49 B N_Y_c_94_n 0.0817758f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_50 N_B_c_56_n N_Y_c_94_n 0.018981f $X=1.17 $Y=1.045 $X2=0 $Y2=0
cc_51 N_B_c_57_n N_Y_c_94_n 0.0127892f $X=1.087 $Y=0.88 $X2=0 $Y2=0
cc_52 N_B_M1002_g N_Y_c_96_n 0.0188594f $X=0.915 $Y=2.625 $X2=0 $Y2=0
cc_53 B N_Y_c_96_n 0.0096619f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_54 B N_VGND_c_116_n 0.0160482f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_55 N_B_c_56_n N_VGND_c_116_n 0.00131325f $X=1.17 $Y=1.045 $X2=0 $Y2=0
cc_56 N_B_c_57_n N_VGND_c_116_n 0.00354189f $X=1.087 $Y=0.88 $X2=0 $Y2=0
cc_57 N_B_c_57_n N_VGND_c_117_n 0.00473265f $X=1.087 $Y=0.88 $X2=0 $Y2=0
cc_58 B N_VGND_c_118_n 0.00109783f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_59 N_B_c_56_n N_VGND_c_118_n 0.00214977f $X=1.17 $Y=1.045 $X2=0 $Y2=0
cc_60 N_B_c_57_n N_VGND_c_118_n 0.00938468f $X=1.087 $Y=0.88 $X2=0 $Y2=0
cc_61 N_VPWR_c_81_n N_Y_c_96_n 0.0022613f $X=0.31 $Y=2.64 $X2=0 $Y2=0
cc_62 N_VPWR_c_82_n N_Y_c_96_n 0.0168794f $X=1.2 $Y=3.33 $X2=0 $Y2=0
cc_63 N_VPWR_c_79_n N_Y_c_96_n 0.0200116f $X=1.2 $Y=3.33 $X2=0 $Y2=0
cc_64 N_Y_c_94_n N_VGND_c_114_n 0.00124848f $X=0.74 $Y=0.495 $X2=0 $Y2=0
cc_65 N_Y_c_94_n N_VGND_c_116_n 0.0120439f $X=0.74 $Y=0.495 $X2=0 $Y2=0
cc_66 N_Y_c_94_n N_VGND_c_117_n 0.012017f $X=0.74 $Y=0.495 $X2=0 $Y2=0
cc_67 N_Y_c_94_n N_VGND_c_118_n 0.00924902f $X=0.74 $Y=0.495 $X2=0 $Y2=0
