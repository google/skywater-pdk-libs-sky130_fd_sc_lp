# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__o2bb2a_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_lp__o2bb2a_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.680000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1_N
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.645000 1.085000 5.170000 1.255000 ;
        RECT 3.645000 1.255000 4.175000 1.515000 ;
        RECT 4.920000 1.255000 5.170000 1.515000 ;
    END
  END A1_N
  PIN A2_N
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.345000 1.425000 4.750000 1.760000 ;
    END
  END A2_N
  PIN B1
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.330000 1.405000 0.815000 1.645000 ;
        RECT 0.625000 1.645000 0.815000 2.310000 ;
        RECT 0.625000 2.310000 2.025000 2.500000 ;
        RECT 1.845000 1.345000 2.095000 1.650000 ;
        RECT 1.845000 1.650000 2.025000 2.310000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.985000 1.405000 1.315000 1.760000 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  1.176000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.680000 1.745000 7.595000 1.925000 ;
        RECT 5.680000 1.925000 5.870000 3.075000 ;
        RECT 5.875000 0.255000 6.135000 1.045000 ;
        RECT 5.875000 1.045000 7.595000 1.235000 ;
        RECT 6.540000 1.925000 6.720000 3.075000 ;
        RECT 6.805000 0.255000 6.995000 1.045000 ;
        RECT 7.345000 1.235000 7.595000 1.745000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 7.680000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 7.680000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.680000 0.085000 ;
      RECT 0.000000  3.245000 7.680000 3.415000 ;
      RECT 0.205000  0.255000 0.465000 1.065000 ;
      RECT 0.205000  1.065000 1.315000 1.235000 ;
      RECT 0.205000  1.815000 0.455000 3.245000 ;
      RECT 0.625000  2.670000 1.765000 3.000000 ;
      RECT 0.635000  0.085000 0.965000 0.895000 ;
      RECT 0.985000  1.930000 1.665000 2.140000 ;
      RECT 1.135000  0.255000 1.325000 0.655000 ;
      RECT 1.135000  0.655000 2.335000 0.825000 ;
      RECT 1.135000  0.825000 1.315000 1.065000 ;
      RECT 1.485000  0.995000 2.760000 1.175000 ;
      RECT 1.485000  1.175000 1.665000 1.930000 ;
      RECT 1.495000  0.085000 1.825000 0.485000 ;
      RECT 1.935000  2.670000 2.420000 3.245000 ;
      RECT 2.005000  0.255000 3.125000 0.435000 ;
      RECT 2.005000  0.435000 2.335000 0.655000 ;
      RECT 2.195000  1.795000 2.420000 2.670000 ;
      RECT 2.505000  0.605000 2.760000 0.995000 ;
      RECT 2.590000  1.175000 2.760000 1.730000 ;
      RECT 2.590000  1.730000 2.930000 2.430000 ;
      RECT 2.590000  2.430000 5.510000 2.610000 ;
      RECT 2.590000  2.610000 2.860000 3.075000 ;
      RECT 2.930000  0.435000 3.125000 1.015000 ;
      RECT 2.930000  1.185000 3.475000 1.515000 ;
      RECT 3.030000  2.780000 3.700000 3.245000 ;
      RECT 3.295000  0.725000 4.575000 0.915000 ;
      RECT 3.295000  0.915000 3.475000 1.185000 ;
      RECT 3.295000  1.515000 3.475000 1.930000 ;
      RECT 3.295000  1.930000 4.945000 2.260000 ;
      RECT 3.385000  0.085000 3.645000 0.555000 ;
      RECT 3.815000  0.255000 5.005000 0.485000 ;
      RECT 4.230000  2.780000 4.560000 3.245000 ;
      RECT 4.245000  0.655000 4.575000 0.725000 ;
      RECT 4.745000  0.485000 5.005000 0.915000 ;
      RECT 5.105000  2.780000 5.435000 3.245000 ;
      RECT 5.175000  0.085000 5.705000 0.915000 ;
      RECT 5.340000  1.405000 7.175000 1.575000 ;
      RECT 5.340000  1.575000 5.510000 2.430000 ;
      RECT 6.040000  2.095000 6.370000 3.245000 ;
      RECT 6.305000  0.085000 6.635000 0.875000 ;
      RECT 6.900000  2.095000 7.230000 3.245000 ;
      RECT 7.165000  0.085000 7.495000 0.875000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
  END
END sky130_fd_sc_lp__o2bb2a_4
END LIBRARY
