* File: sky130_fd_sc_lp__dfbbp_1.spice
* Created: Wed Sep  2 09:43:07 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__dfbbp_1.pex.spice"
.subckt sky130_fd_sc_lp__dfbbp_1  VNB VPB CLK D SET_B RESET_B VPWR Q_N Q VGND
* 
* VGND	VGND
* Q	Q
* Q_N	Q_N
* VPWR	VPWR
* RESET_B	RESET_B
* SET_B	SET_B
* D	D
* CLK	CLK
* VPB	VPB
* VNB	VNB
MM1018 N_A_114_57#_M1018_d N_CLK_M1018_g N_VGND_M1018_s VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.1197 PD=1.41 PS=1.41 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1008 N_VGND_M1008_d N_A_114_57#_M1008_g N_A_225_47#_M1008_s VNB NSHORT L=0.15
+ W=0.42 AD=0.19845 AS=0.1197 PD=1.365 PS=1.41 NRD=65.712 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75004.3 A=0.063 P=1.14 MULT=1
MM1002 N_A_531_47#_M1002_d N_D_M1002_g N_VGND_M1008_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.19845 PD=0.7 PS=1.365 NRD=0 NRS=124.284 M=1 R=2.8 SA=75001.3
+ SB=75003.2 A=0.063 P=1.14 MULT=1
MM1021 N_A_617_47#_M1021_d N_A_114_57#_M1021_g N_A_531_47#_M1002_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.0756 AS=0.0588 PD=0.78 PS=0.7 NRD=22.848 NRS=0 M=1 R=2.8
+ SA=75001.7 SB=75002.7 A=0.063 P=1.14 MULT=1
MM1031 A_719_47# N_A_225_47#_M1031_g N_A_617_47#_M1021_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0504 AS=0.0756 PD=0.66 PS=0.78 NRD=18.564 NRS=0 M=1 R=2.8
+ SA=75002.2 SB=75002.2 A=0.063 P=1.14 MULT=1
MM1028 N_VGND_M1028_d N_A_767_21#_M1028_g A_719_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.106704 AS=0.0504 PD=0.863774 PS=0.66 NRD=25.704 NRS=18.564 M=1 R=2.8
+ SA=75002.6 SB=75001.8 A=0.063 P=1.14 MULT=1
MM1003 N_A_917_47#_M1003_d N_SET_B_M1003_g N_VGND_M1028_d VNB NSHORT L=0.15
+ W=0.64 AD=0.0896 AS=0.162596 PD=0.92 PS=1.31623 NRD=0 NRS=14.988 M=1 R=4.26667
+ SA=75002.2 SB=75001.2 A=0.096 P=1.58 MULT=1
MM1023 N_A_767_21#_M1023_d N_A_617_47#_M1023_g N_A_917_47#_M1003_d VNB NSHORT
+ L=0.15 W=0.64 AD=0.1408 AS=0.0896 PD=1.08 PS=0.92 NRD=14.988 NRS=0 M=1
+ R=4.26667 SA=75002.7 SB=75000.8 A=0.096 P=1.58 MULT=1
MM1019 N_A_917_47#_M1019_d N_A_1091_21#_M1019_g N_A_767_21#_M1023_d VNB NSHORT
+ L=0.15 W=0.64 AD=0.1824 AS=0.1408 PD=1.85 PS=1.08 NRD=0 NRS=14.988 M=1
+ R=4.26667 SA=75003.2 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1012 A_1319_54# N_A_767_21#_M1012_g N_VGND_M1012_s VNB NSHORT L=0.15 W=0.64
+ AD=0.0768 AS=0.1824 PD=0.88 PS=1.85 NRD=12.18 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75002.3 A=0.096 P=1.58 MULT=1
MM1013 N_A_1307_428#_M1013_d N_A_225_47#_M1013_g A_1319_54# VNB NSHORT L=0.15
+ W=0.64 AD=0.129147 AS=0.0768 PD=1.20755 PS=0.88 NRD=0 NRS=12.18 M=1 R=4.26667
+ SA=75000.6 SB=75001.9 A=0.096 P=1.58 MULT=1
MM1004 A_1499_98# N_A_114_57#_M1004_g N_A_1307_428#_M1013_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0504 AS=0.0847528 PD=0.66 PS=0.792453 NRD=18.564 NRS=22.848 M=1
+ R=2.8 SA=75001.1 SB=75002.2 A=0.063 P=1.14 MULT=1
MM1005 N_VGND_M1005_d N_A_1545_332#_M1005_g A_1499_98# VNB NSHORT L=0.15 W=0.42
+ AD=0.11336 AS=0.0504 PD=0.895472 PS=0.66 NRD=38.568 NRS=18.564 M=1 R=2.8
+ SA=75001.5 SB=75001.9 A=0.063 P=1.14 MULT=1
MM1020 N_A_1705_54#_M1020_d N_SET_B_M1020_g N_VGND_M1005_d VNB NSHORT L=0.15
+ W=0.64 AD=0.0896 AS=0.17274 PD=0.92 PS=1.36453 NRD=0 NRS=14.988 M=1 R=4.26667
+ SA=75001.5 SB=75001.2 A=0.096 P=1.58 MULT=1
MM1029 N_A_1545_332#_M1029_d N_A_1307_428#_M1029_g N_A_1705_54#_M1020_d VNB
+ NSHORT L=0.15 W=0.64 AD=0.214012 AS=0.0896 PD=1.6 PS=0.92 NRD=52.38 NRS=0 M=1
+ R=4.26667 SA=75001.9 SB=75000.8 A=0.096 P=1.58 MULT=1
MM1014 N_A_1705_54#_M1014_d N_A_1091_21#_M1014_g N_A_1545_332#_M1029_d VNB
+ NSHORT L=0.15 W=0.64 AD=0.1792 AS=0.214012 PD=1.84 PS=1.6 NRD=0 NRS=52.38 M=1
+ R=4.26667 SA=75002.5 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1035 N_VGND_M1035_d N_RESET_B_M1035_g N_A_1091_21#_M1035_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0903 AS=0.1197 PD=0.8 PS=1.41 NRD=22.848 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1037 N_Q_N_M1037_d N_A_1545_332#_M1037_g N_VGND_M1035_d VNB NSHORT L=0.15
+ W=0.84 AD=0.2394 AS=0.1806 PD=2.25 PS=1.6 NRD=0 NRS=0 M=1 R=5.6 SA=75000.5
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1000 N_VGND_M1000_d N_A_1545_332#_M1000_g N_A_2317_367#_M1000_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.0903 AS=0.1176 PD=0.8 PS=1.4 NRD=22.848 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1039 N_Q_M1039_d N_A_2317_367#_M1039_g N_VGND_M1000_d VNB NSHORT L=0.15 W=0.84
+ AD=0.2394 AS=0.1806 PD=2.25 PS=1.6 NRD=0 NRS=0 M=1 R=5.6 SA=75000.5 SB=75000.2
+ A=0.126 P=1.98 MULT=1
MM1033 N_A_114_57#_M1033_d N_CLK_M1033_g N_VPWR_M1033_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1824 AS=0.2336 PD=1.85 PS=2.01 NRD=0 NRS=24.6053 M=1 R=4.26667
+ SA=75000.3 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1011 N_VPWR_M1011_d N_A_114_57#_M1011_g N_A_225_47#_M1011_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.295728 AS=0.1824 PD=1.95019 PS=1.85 NRD=24.6053 NRS=0 M=1
+ R=4.26667 SA=75000.2 SB=75004.2 A=0.096 P=1.58 MULT=1
MM1006 N_A_531_47#_M1006_d N_D_M1006_g N_VPWR_M1011_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0588 AS=0.194072 PD=0.7 PS=1.27981 NRD=0 NRS=190.932 M=1 R=2.8 SA=75001.3
+ SB=75005.1 A=0.063 P=1.14 MULT=1
MM1032 N_A_617_47#_M1032_d N_A_225_47#_M1032_g N_A_531_47#_M1006_d VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.0756 AS=0.0588 PD=0.78 PS=0.7 NRD=37.5088 NRS=0 M=1 R=2.8
+ SA=75001.8 SB=75004.7 A=0.063 P=1.14 MULT=1
MM1034 A_755_463# N_A_114_57#_M1034_g N_A_617_47#_M1032_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0504 AS=0.0756 PD=0.66 PS=0.78 NRD=30.4759 NRS=0 M=1 R=2.8
+ SA=75002.3 SB=75004.2 A=0.063 P=1.14 MULT=1
MM1009 N_VPWR_M1009_d N_A_767_21#_M1009_g A_755_463# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.14365 AS=0.0504 PD=1.05333 PS=0.66 NRD=134.61 NRS=30.4759 M=1 R=2.8
+ SA=75002.7 SB=75003.8 A=0.063 P=1.14 MULT=1
MM1030 N_A_767_21#_M1030_d N_SET_B_M1030_g N_VPWR_M1009_d VPB PHIGHVT L=0.15
+ W=0.84 AD=0.1176 AS=0.2873 PD=1.12 PS=2.10667 NRD=0 NRS=67.2952 M=1 R=5.6
+ SA=75001.8 SB=75002.4 A=0.126 P=1.98 MULT=1
MM1015 A_1046_379# N_A_617_47#_M1015_g N_A_767_21#_M1030_d VPB PHIGHVT L=0.15
+ W=0.84 AD=0.1008 AS=0.1176 PD=1.08 PS=1.12 NRD=15.2281 NRS=0 M=1 R=5.6
+ SA=75002.2 SB=75002 A=0.126 P=1.98 MULT=1
MM1016 N_VPWR_M1016_d N_A_1091_21#_M1016_g A_1046_379# VPB PHIGHVT L=0.15 W=0.84
+ AD=0.1218 AS=0.1008 PD=1.13 PS=1.08 NRD=0 NRS=15.2281 M=1 R=5.6 SA=75002.6
+ SB=75001.6 A=0.126 P=1.98 MULT=1
MM1026 A_1212_379# N_A_767_21#_M1026_g N_VPWR_M1016_d VPB PHIGHVT L=0.15 W=0.84
+ AD=0.157937 AS=0.1218 PD=1.41 PS=1.13 NRD=31.1851 NRS=2.3443 M=1 R=5.6
+ SA=75003.1 SB=75001.1 A=0.126 P=1.98 MULT=1
MM1017 N_A_1307_428#_M1017_d N_A_114_57#_M1017_g A_1212_379# VPB PHIGHVT L=0.15
+ W=0.84 AD=0.1848 AS=0.157937 PD=1.66667 PS=1.41 NRD=30.4759 NRS=31.1851 M=1
+ R=5.6 SA=75003 SB=75001.7 A=0.126 P=1.98 MULT=1
MM1007 A_1419_512# N_A_225_47#_M1007_g N_A_1307_428#_M1017_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1344 AS=0.0924 PD=1.06 PS=0.833333 NRD=124.287 NRS=0 M=1 R=2.8
+ SA=75002.8 SB=75002.6 A=0.063 P=1.14 MULT=1
MM1036 N_VPWR_M1036_d N_A_1545_332#_M1036_g A_1419_512# VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1183 AS=0.1344 PD=0.933333 PS=1.06 NRD=131.32 NRS=124.287 M=1
+ R=2.8 SA=75003.5 SB=75001.8 A=0.063 P=1.14 MULT=1
MM1010 N_A_1545_332#_M1010_d N_SET_B_M1010_g N_VPWR_M1036_d VPB PHIGHVT L=0.15
+ W=0.84 AD=0.1554 AS=0.2366 PD=1.21 PS=1.86667 NRD=21.0987 NRS=0 M=1 R=5.6
+ SA=75002.2 SB=75001.1 A=0.126 P=1.98 MULT=1
MM1038 A_1823_430# N_A_1307_428#_M1038_g N_A_1545_332#_M1010_d VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.1092 AS=0.1554 PD=1.1 PS=1.21 NRD=17.5724 NRS=0 M=1 R=5.6
+ SA=75002.8 SB=75000.6 A=0.126 P=1.98 MULT=1
MM1001 N_VPWR_M1001_d N_A_1091_21#_M1001_g A_1823_430# VPB PHIGHVT L=0.15 W=0.84
+ AD=0.2394 AS=0.1092 PD=2.25 PS=1.1 NRD=0 NRS=17.5724 M=1 R=5.6 SA=75003.2
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1025 N_VPWR_M1025_d N_RESET_B_M1025_g N_A_1091_21#_M1025_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.137128 AS=0.1824 PD=1.09137 PS=1.85 NRD=49.0136 NRS=0 M=1
+ R=4.26667 SA=75000.2 SB=75000.7 A=0.096 P=1.58 MULT=1
MM1027 N_Q_N_M1027_d N_A_1545_332#_M1027_g N_VPWR_M1025_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3591 AS=0.269972 PD=3.09 PS=2.14863 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.5 SB=75000.2 A=0.189 P=2.82 MULT=1
MM1022 N_VPWR_M1022_d N_A_1545_332#_M1022_g N_A_2317_367#_M1022_s VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.137128 AS=0.1824 PD=1.09137 PS=1.85 NRD=25.3933 NRS=0 M=1
+ R=4.26667 SA=75000.2 SB=75000.7 A=0.096 P=1.58 MULT=1
MM1024 N_Q_M1024_d N_A_2317_367#_M1024_g N_VPWR_M1022_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3591 AS=0.269972 PD=3.09 PS=2.14863 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.5 SB=75000.2 A=0.189 P=2.82 MULT=1
DX40_noxref VNB VPB NWDIODE A=24.6998 P=31.28
c_145 VNB 0 2.46682e-19 $X=0 $Y=0
c_258 VPB 0 9.67699e-20 $X=0 $Y=3.085
c_1856 A_755_463# 0 1.19365e-19 $X=3.775 $Y=2.315
*
.include "sky130_fd_sc_lp__dfbbp_1.pxi.spice"
*
.ends
*
*
