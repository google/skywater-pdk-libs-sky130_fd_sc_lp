* File: sky130_fd_sc_lp__a32o_0.spice
* Created: Fri Aug 28 10:00:47 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__a32o_0.pex.spice"
.subckt sky130_fd_sc_lp__a32o_0  VNB VPB A3 A2 A1 B1 B2 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* B2	B2
* B1	B1
* A1	A1
* A2	A2
* A3	A3
* VPB	VPB
* VNB	VNB
MM1005 N_VGND_M1005_d N_A_80_21#_M1005_g N_X_M1005_s VNB NSHORT L=0.15 W=0.42
+ AD=0.14175 AS=0.1113 PD=1.095 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75003 A=0.063 P=1.14 MULT=1
MM1004 A_275_47# N_A3_M1004_g N_VGND_M1005_d VNB NSHORT L=0.15 W=0.42 AD=0.0609
+ AS=0.14175 PD=0.71 PS=1.095 NRD=25.704 NRS=0 M=1 R=2.8 SA=75001 SB=75002.2
+ A=0.063 P=1.14 MULT=1
MM1000 A_363_47# N_A2_M1000_g A_275_47# VNB NSHORT L=0.15 W=0.42 AD=0.0651
+ AS=0.0609 PD=0.73 PS=0.71 NRD=28.56 NRS=25.704 M=1 R=2.8 SA=75001.5 SB=75001.7
+ A=0.063 P=1.14 MULT=1
MM1007 N_A_80_21#_M1007_d N_A1_M1007_g A_363_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.0819 AS=0.0651 PD=0.81 PS=0.73 NRD=14.28 NRS=28.56 M=1 R=2.8 SA=75001.9
+ SB=75001.3 A=0.063 P=1.14 MULT=1
MM1010 A_563_47# N_B1_M1010_g N_A_80_21#_M1007_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0819 AS=0.0819 PD=0.81 PS=0.81 NRD=39.996 NRS=17.136 M=1 R=2.8 SA=75002.5
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1002 N_VGND_M1002_d N_B2_M1002_g A_563_47# VNB NSHORT L=0.15 W=0.42 AD=0.1176
+ AS=0.0819 PD=1.4 PS=0.81 NRD=4.284 NRS=39.996 M=1 R=2.8 SA=75003 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1009 N_VPWR_M1009_d N_A_80_21#_M1009_g N_X_M1009_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0896 AS=0.1696 PD=0.92 PS=1.81 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75002.6 A=0.096 P=1.58 MULT=1
MM1006 N_A_269_429#_M1006_d N_A3_M1006_g N_VPWR_M1009_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.12 AS=0.0896 PD=1.015 PS=0.92 NRD=16.9223 NRS=0 M=1 R=4.26667
+ SA=75000.6 SB=75002.1 A=0.096 P=1.58 MULT=1
MM1003 N_VPWR_M1003_d N_A2_M1003_g N_A_269_429#_M1006_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.12 AS=0.12 PD=1.015 PS=1.015 NRD=6.1464 NRS=12.2928 M=1 R=4.26667
+ SA=75001.1 SB=75001.6 A=0.096 P=1.58 MULT=1
MM1011 N_A_269_429#_M1011_d N_A1_M1011_g N_VPWR_M1003_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.096 AS=0.12 PD=0.94 PS=1.015 NRD=0 NRS=23.0687 M=1 R=4.26667
+ SA=75001.7 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1001 N_A_80_21#_M1001_d N_B1_M1001_g N_A_269_429#_M1011_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.0896 AS=0.096 PD=0.92 PS=0.94 NRD=0 NRS=6.1464 M=1 R=4.26667
+ SA=75002.1 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1008 N_A_269_429#_M1008_d N_B2_M1008_g N_A_80_21#_M1001_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1696 AS=0.0896 PD=1.81 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75002.6 SB=75000.2 A=0.096 P=1.58 MULT=1
DX12_noxref VNB VPB NWDIODE A=7.8703 P=12.17
*
.include "sky130_fd_sc_lp__a32o_0.pxi.spice"
*
.ends
*
*
