* File: sky130_fd_sc_lp__o211ai_0.pex.spice
* Created: Wed Sep  2 10:14:22 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O211AI_0%A1 1 3 7 10 11 12 13 18
c34 18 0 6.75121e-20 $X=0.49 $Y=1.245
r35 17 18 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.49
+ $Y=1.245 $X2=0.49 $Y2=1.245
r36 12 13 9.03161 $w=4.88e-07 $l=3.7e-07 $layer=LI1_cond $X=0.33 $Y=1.295
+ $X2=0.33 $Y2=1.665
r37 12 18 1.22049 $w=4.88e-07 $l=5e-08 $layer=LI1_cond $X=0.33 $Y=1.295 $X2=0.33
+ $Y2=1.245
r38 10 17 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.49 $Y=1.585
+ $X2=0.49 $Y2=1.245
r39 10 11 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.49 $Y=1.585
+ $X2=0.49 $Y2=1.75
r40 7 11 458.926 $w=1.5e-07 $l=8.95e-07 $layer=POLY_cond $X=0.58 $Y=2.645
+ $X2=0.58 $Y2=1.75
r41 1 17 58.9111 $w=2.7e-07 $l=3.44674e-07 $layer=POLY_cond $X=0.52 $Y=0.915
+ $X2=0.49 $Y2=1.245
r42 1 3 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=0.52 $Y=0.915 $X2=0.52
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__O211AI_0%A2 2 5 9 11 12 15 17 18 22 24
c49 24 0 6.75121e-20 $X=1.045 $Y=1.155
r50 22 24 46.5827 $w=3.6e-07 $l=1.65e-07 $layer=POLY_cond $X=1.045 $Y=1.32
+ $X2=1.045 $Y2=1.155
r51 22 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.06
+ $Y=1.32 $X2=1.06 $Y2=1.32
r52 18 23 9.93982 $w=3.98e-07 $l=3.45e-07 $layer=LI1_cond $X=1.095 $Y=1.665
+ $X2=1.095 $Y2=1.32
r53 17 23 0.720277 $w=3.98e-07 $l=2.5e-08 $layer=LI1_cond $X=1.095 $Y=1.295
+ $X2=1.095 $Y2=1.32
r54 13 15 71.7872 $w=1.5e-07 $l=1.4e-07 $layer=POLY_cond $X=1.15 $Y=0.845
+ $X2=1.29 $Y2=0.845
r55 9 15 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.29 $Y=0.77 $X2=1.29
+ $Y2=0.845
r56 9 11 104.433 $w=1.5e-07 $l=3.25e-07 $layer=POLY_cond $X=1.29 $Y=0.77
+ $X2=1.29 $Y2=0.445
r57 7 13 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.15 $Y=0.92 $X2=1.15
+ $Y2=0.845
r58 7 24 120.5 $w=1.5e-07 $l=2.35e-07 $layer=POLY_cond $X=1.15 $Y=0.92 $X2=1.15
+ $Y2=1.155
r59 5 12 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=0.94 $Y=2.645
+ $X2=0.94 $Y2=1.825
r60 2 12 48.987 $w=3.6e-07 $l=1.8e-07 $layer=POLY_cond $X=1.045 $Y=1.645
+ $X2=1.045 $Y2=1.825
r61 1 22 2.40434 $w=3.6e-07 $l=1.5e-08 $layer=POLY_cond $X=1.045 $Y=1.335
+ $X2=1.045 $Y2=1.32
r62 1 2 49.6898 $w=3.6e-07 $l=3.1e-07 $layer=POLY_cond $X=1.045 $Y=1.335
+ $X2=1.045 $Y2=1.645
.ends

.subckt PM_SKY130_FD_SC_LP__O211AI_0%B1 1 3 5 8 12 16 17 18 19 23
r51 18 19 11.3708 $w=3.73e-07 $l=3.7e-07 $layer=LI1_cond $X=1.652 $Y=1.295
+ $X2=1.652 $Y2=1.665
r52 18 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.63
+ $Y=1.325 $X2=1.63 $Y2=1.325
r53 16 23 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.63 $Y=1.665
+ $X2=1.63 $Y2=1.325
r54 16 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.63 $Y=1.665
+ $X2=1.63 $Y2=1.83
r55 15 23 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.63 $Y=1.16
+ $X2=1.63 $Y2=1.325
r56 10 12 87.1702 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=1.37 $Y=2.14
+ $X2=1.54 $Y2=2.14
r57 8 15 366.628 $w=1.5e-07 $l=7.15e-07 $layer=POLY_cond $X=1.72 $Y=0.445
+ $X2=1.72 $Y2=1.16
r58 5 12 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.54 $Y=2.065
+ $X2=1.54 $Y2=2.14
r59 5 17 120.5 $w=1.5e-07 $l=2.35e-07 $layer=POLY_cond $X=1.54 $Y=2.065 $X2=1.54
+ $Y2=1.83
r60 1 10 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.37 $Y=2.215
+ $X2=1.37 $Y2=2.14
r61 1 3 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=1.37 $Y=2.215 $X2=1.37
+ $Y2=2.645
.ends

.subckt PM_SKY130_FD_SC_LP__O211AI_0%C1 3 5 7 9 10 11
r28 16 17 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.485
+ $Y=1.005 $X2=2.485 $Y2=1.005
r29 10 11 10.795 $w=3.93e-07 $l=3.7e-07 $layer=LI1_cond $X=2.597 $Y=1.295
+ $X2=2.597 $Y2=1.665
r30 10 17 8.46097 $w=3.93e-07 $l=2.9e-07 $layer=LI1_cond $X=2.597 $Y=1.295
+ $X2=2.597 $Y2=1.005
r31 9 17 2.33406 $w=3.93e-07 $l=8e-08 $layer=LI1_cond $X=2.597 $Y=0.925
+ $X2=2.597 $Y2=1.005
r32 5 16 71.5532 $w=6.2e-07 $l=5.91151e-07 $layer=POLY_cond $X=2.14 $Y=1.51
+ $X2=2.327 $Y2=1.005
r33 5 7 581.989 $w=1.5e-07 $l=1.135e-06 $layer=POLY_cond $X=2.14 $Y=1.51
+ $X2=2.14 $Y2=2.645
r34 1 16 45.1209 $w=6.2e-07 $l=3.19005e-07 $layer=POLY_cond $X=2.08 $Y=0.84
+ $X2=2.327 $Y2=1.005
r35 1 3 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=2.08 $Y=0.84 $X2=2.08
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__O211AI_0%VPWR 1 2 7 9 13 15 17 24 25 31
r32 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r33 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r34 25 32 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=1.68 $Y2=3.33
r35 24 25 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r36 22 31 12.4404 $w=1.7e-07 $l=2.95e-07 $layer=LI1_cond $X=2.05 $Y=3.33
+ $X2=1.755 $Y2=3.33
r37 22 24 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=2.05 $Y=3.33 $X2=2.64
+ $Y2=3.33
r38 21 29 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.24 $Y2=3.33
r39 20 21 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r40 18 28 4.57341 $w=1.7e-07 $l=2.65e-07 $layer=LI1_cond $X=0.53 $Y=3.33
+ $X2=0.265 $Y2=3.33
r41 18 20 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=0.53 $Y=3.33 $X2=1.2
+ $Y2=3.33
r42 17 31 12.4404 $w=1.7e-07 $l=2.95e-07 $layer=LI1_cond $X=1.46 $Y=3.33
+ $X2=1.755 $Y2=3.33
r43 17 20 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=1.46 $Y=3.33 $X2=1.2
+ $Y2=3.33
r44 15 32 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=1.68 $Y2=3.33
r45 15 21 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=1.2 $Y2=3.33
r46 11 31 2.48142 $w=5.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.755 $Y=3.245
+ $X2=1.755 $Y2=3.33
r47 11 13 15.7112 $w=5.88e-07 $l=7.75e-07 $layer=LI1_cond $X=1.755 $Y=3.245
+ $X2=1.755 $Y2=2.47
r48 7 28 3.19276 $w=3.3e-07 $l=1.36015e-07 $layer=LI1_cond $X=0.365 $Y=3.245
+ $X2=0.265 $Y2=3.33
r49 7 9 27.0649 $w=3.28e-07 $l=7.75e-07 $layer=LI1_cond $X=0.365 $Y=3.245
+ $X2=0.365 $Y2=2.47
r50 2 13 150 $w=1.7e-07 $l=5.47723e-07 $layer=licon1_PDIFF $count=4 $X=1.445
+ $Y=2.325 $X2=1.925 $Y2=2.47
r51 1 9 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.24
+ $Y=2.325 $X2=0.365 $Y2=2.47
.ends

.subckt PM_SKY130_FD_SC_LP__O211AI_0%Y 1 2 3 10 12 18 20 21 22 24 25 33
r47 25 41 6.34442 $w=5.73e-07 $l=3.05e-07 $layer=LI1_cond $X=2.507 $Y=2.775
+ $X2=2.507 $Y2=2.47
r48 24 41 1.35209 $w=5.73e-07 $l=6.5e-08 $layer=LI1_cond $X=2.507 $Y=2.405
+ $X2=2.507 $Y2=2.47
r49 24 37 5.61637 $w=5.73e-07 $l=2.7e-07 $layer=LI1_cond $X=2.507 $Y=2.405
+ $X2=2.507 $Y2=2.135
r50 22 33 4.14799 $w=1.85e-07 $l=3.92e-07 $layer=LI1_cond $X=2.402 $Y=2.042
+ $X2=2.01 $Y2=2.042
r51 22 37 2.66143 $w=3.92e-07 $l=1.44187e-07 $layer=LI1_cond $X=2.402 $Y=2.042
+ $X2=2.507 $Y2=2.135
r52 21 33 19.7838 $w=1.83e-07 $l=3.3e-07 $layer=LI1_cond $X=1.68 $Y=2.042
+ $X2=2.01 $Y2=2.042
r53 21 34 23.3808 $w=1.83e-07 $l=3.9e-07 $layer=LI1_cond $X=1.68 $Y=2.042
+ $X2=1.29 $Y2=2.042
r54 20 34 4.52293 $w=1.85e-07 $l=1.5e-07 $layer=LI1_cond $X=1.14 $Y=2.042
+ $X2=1.29 $Y2=2.042
r55 15 22 44.5673 $w=3.53e-07 $l=1.335e-06 $layer=LI1_cond $X=2.115 $Y=0.615
+ $X2=2.115 $Y2=1.95
r56 14 18 6.19223 $w=3.33e-07 $l=1.8e-07 $layer=LI1_cond $X=2.115 $Y=0.447
+ $X2=2.295 $Y2=0.447
r57 14 15 3.46964 $w=2.1e-07 $l=1.68e-07 $layer=LI1_cond $X=2.115 $Y=0.447
+ $X2=2.115 $Y2=0.615
r58 10 20 2.80421 $w=3e-07 $l=9.3e-08 $layer=LI1_cond $X=1.14 $Y=2.135 $X2=1.14
+ $Y2=2.042
r59 10 12 12.8689 $w=2.98e-07 $l=3.35e-07 $layer=LI1_cond $X=1.14 $Y=2.135
+ $X2=1.14 $Y2=2.47
r60 3 41 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=2.215
+ $Y=2.325 $X2=2.355 $Y2=2.47
r61 2 12 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=1.015
+ $Y=2.325 $X2=1.155 $Y2=2.47
r62 1 18 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.155
+ $Y=0.235 $X2=2.295 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__O211AI_0%A_36_47# 1 2 9 11 12 15
r34 13 15 13.0758 $w=2.58e-07 $l=2.95e-07 $layer=LI1_cond $X=1.54 $Y=0.74
+ $X2=1.54 $Y2=0.445
r35 11 13 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=1.41 $Y=0.825
+ $X2=1.54 $Y2=0.74
r36 11 12 65.8931 $w=1.68e-07 $l=1.01e-06 $layer=LI1_cond $X=1.41 $Y=0.825
+ $X2=0.4 $Y2=0.825
r37 7 12 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=0.27 $Y=0.74
+ $X2=0.4 $Y2=0.825
r38 7 9 13.0758 $w=2.58e-07 $l=2.95e-07 $layer=LI1_cond $X=0.27 $Y=0.74 $X2=0.27
+ $Y2=0.445
r39 2 15 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.365
+ $Y=0.235 $X2=1.505 $Y2=0.445
r40 1 9 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.18
+ $Y=0.235 $X2=0.305 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__O211AI_0%VGND 1 4 13 14 19 25
r31 23 25 8.23183 $w=6.53e-07 $l=4e-08 $layer=LI1_cond $X=1.2 $Y=0.242 $X2=1.24
+ $Y2=0.242
r32 23 24 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r33 21 23 2.28259 $w=6.53e-07 $l=1.25e-07 $layer=LI1_cond $X=1.075 $Y=0.242
+ $X2=1.2 $Y2=0.242
r34 18 24 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r35 17 21 6.48256 $w=6.53e-07 $l=3.55e-07 $layer=LI1_cond $X=0.72 $Y=0.242
+ $X2=1.075 $Y2=0.242
r36 17 19 10.2405 $w=6.53e-07 $l=1.5e-07 $layer=LI1_cond $X=0.72 $Y=0.242
+ $X2=0.57 $Y2=0.242
r37 17 18 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r38 13 25 91.3369 $w=1.68e-07 $l=1.4e-06 $layer=LI1_cond $X=2.64 $Y=0 $X2=1.24
+ $Y2=0
r39 13 14 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r40 9 18 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r41 8 19 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=0.24 $Y=0 $X2=0.57
+ $Y2=0
r42 8 9 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r43 4 14 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=1.44 $Y=0 $X2=2.64
+ $Y2=0
r44 4 24 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=1.2
+ $Y2=0
r45 1 21 91 $w=1.7e-07 $l=5.755e-07 $layer=licon1_NDIFF $count=2 $X=0.595
+ $Y=0.235 $X2=1.075 $Y2=0.445
.ends

