* File: sky130_fd_sc_lp__dlxtn_2.pxi.spice
* Created: Wed Sep  2 09:48:31 2020
* 
x_PM_SKY130_FD_SC_LP__DLXTN_2%D N_D_M1007_g N_D_M1010_g D D D N_D_c_140_n
+ N_D_c_141_n PM_SKY130_FD_SC_LP__DLXTN_2%D
x_PM_SKY130_FD_SC_LP__DLXTN_2%GATE_N N_GATE_N_c_174_n N_GATE_N_M1017_g
+ N_GATE_N_M1002_g N_GATE_N_c_176_n N_GATE_N_c_177_n N_GATE_N_c_178_n GATE_N
+ GATE_N GATE_N N_GATE_N_c_180_n PM_SKY130_FD_SC_LP__DLXTN_2%GATE_N
x_PM_SKY130_FD_SC_LP__DLXTN_2%A_242_130# N_A_242_130#_M1017_d
+ N_A_242_130#_M1002_d N_A_242_130#_M1011_g N_A_242_130#_c_219_n
+ N_A_242_130#_c_220_n N_A_242_130#_c_221_n N_A_242_130#_M1006_g
+ N_A_242_130#_M1014_g N_A_242_130#_M1003_g N_A_242_130#_c_223_n
+ N_A_242_130#_c_224_n N_A_242_130#_c_233_n N_A_242_130#_c_234_n
+ N_A_242_130#_c_235_n N_A_242_130#_c_258_p N_A_242_130#_c_236_n
+ N_A_242_130#_c_237_n N_A_242_130#_c_225_n N_A_242_130#_c_226_n
+ N_A_242_130#_c_238_n N_A_242_130#_c_239_n N_A_242_130#_c_240_n
+ N_A_242_130#_c_227_n N_A_242_130#_c_228_n N_A_242_130#_c_229_n
+ N_A_242_130#_c_230_n PM_SKY130_FD_SC_LP__DLXTN_2%A_242_130#
x_PM_SKY130_FD_SC_LP__DLXTN_2%A_57_130# N_A_57_130#_M1007_s N_A_57_130#_M1010_s
+ N_A_57_130#_M1015_g N_A_57_130#_c_367_n N_A_57_130#_c_368_n
+ N_A_57_130#_M1019_g N_A_57_130#_c_374_n N_A_57_130#_c_370_n
+ N_A_57_130#_c_375_n N_A_57_130#_c_376_n N_A_57_130#_c_371_n
+ N_A_57_130#_c_377_n N_A_57_130#_c_412_n N_A_57_130#_c_372_n
+ PM_SKY130_FD_SC_LP__DLXTN_2%A_57_130#
x_PM_SKY130_FD_SC_LP__DLXTN_2%A_349_481# N_A_349_481#_M1006_s
+ N_A_349_481#_M1011_s N_A_349_481#_M1016_g N_A_349_481#_c_446_n
+ N_A_349_481#_c_447_n N_A_349_481#_M1004_g N_A_349_481#_c_449_n
+ N_A_349_481#_c_457_n N_A_349_481#_c_458_n N_A_349_481#_c_459_n
+ N_A_349_481#_c_460_n N_A_349_481#_c_450_n N_A_349_481#_c_451_n
+ N_A_349_481#_c_452_n N_A_349_481#_c_496_n N_A_349_481#_c_453_n
+ N_A_349_481#_c_454_n N_A_349_481#_c_455_n
+ PM_SKY130_FD_SC_LP__DLXTN_2%A_349_481#
x_PM_SKY130_FD_SC_LP__DLXTN_2%A_849_419# N_A_849_419#_M1005_d
+ N_A_849_419#_M1000_d N_A_849_419#_M1013_g N_A_849_419#_M1008_g
+ N_A_849_419#_c_560_n N_A_849_419#_M1001_g N_A_849_419#_M1012_g
+ N_A_849_419#_c_562_n N_A_849_419#_M1009_g N_A_849_419#_M1018_g
+ N_A_849_419#_c_578_n N_A_849_419#_c_565_n N_A_849_419#_c_566_n
+ N_A_849_419#_c_567_n N_A_849_419#_c_580_n N_A_849_419#_c_568_n
+ N_A_849_419#_c_581_n N_A_849_419#_c_569_n N_A_849_419#_c_570_n
+ N_A_849_419#_c_571_n N_A_849_419#_c_572_n N_A_849_419#_c_573_n
+ N_A_849_419#_c_574_n PM_SKY130_FD_SC_LP__DLXTN_2%A_849_419#
x_PM_SKY130_FD_SC_LP__DLXTN_2%A_663_481# N_A_663_481#_M1014_d
+ N_A_663_481#_M1016_d N_A_663_481#_M1005_g N_A_663_481#_M1000_g
+ N_A_663_481#_c_685_n N_A_663_481#_c_692_n N_A_663_481#_c_677_n
+ N_A_663_481#_c_678_n N_A_663_481#_c_698_n N_A_663_481#_c_679_n
+ N_A_663_481#_c_680_n N_A_663_481#_c_681_n N_A_663_481#_c_682_n
+ N_A_663_481#_c_683_n PM_SKY130_FD_SC_LP__DLXTN_2%A_663_481#
x_PM_SKY130_FD_SC_LP__DLXTN_2%VPWR N_VPWR_M1010_d N_VPWR_M1011_d N_VPWR_M1013_d
+ N_VPWR_M1012_d N_VPWR_M1018_d N_VPWR_c_777_n N_VPWR_c_778_n N_VPWR_c_824_n
+ N_VPWR_c_779_n N_VPWR_c_780_n N_VPWR_c_781_n N_VPWR_c_782_n N_VPWR_c_783_n
+ VPWR N_VPWR_c_784_n N_VPWR_c_785_n N_VPWR_c_786_n N_VPWR_c_787_n
+ N_VPWR_c_788_n N_VPWR_c_789_n N_VPWR_c_790_n N_VPWR_c_776_n
+ PM_SKY130_FD_SC_LP__DLXTN_2%VPWR
x_PM_SKY130_FD_SC_LP__DLXTN_2%Q N_Q_M1001_s N_Q_M1012_s Q Q Q Q Q Q Q
+ N_Q_c_864_n PM_SKY130_FD_SC_LP__DLXTN_2%Q
x_PM_SKY130_FD_SC_LP__DLXTN_2%VGND N_VGND_M1007_d N_VGND_M1006_d N_VGND_M1008_d
+ N_VGND_M1001_d N_VGND_M1009_d N_VGND_c_884_n N_VGND_c_885_n N_VGND_c_886_n
+ N_VGND_c_887_n N_VGND_c_888_n N_VGND_c_889_n N_VGND_c_900_n VGND
+ N_VGND_c_890_n N_VGND_c_891_n N_VGND_c_892_n N_VGND_c_893_n N_VGND_c_894_n
+ N_VGND_c_895_n N_VGND_c_896_n N_VGND_c_897_n N_VGND_c_898_n
+ PM_SKY130_FD_SC_LP__DLXTN_2%VGND
cc_1 VNB N_D_M1010_g 0.00861086f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=2.725
cc_2 VNB D 0.0167257f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.21
cc_3 VNB N_D_c_140_n 0.03533f $X=-0.19 $Y=-0.245 $X2=0.655 $Y2=1.345
cc_4 VNB N_D_c_141_n 0.0216145f $X=-0.19 $Y=-0.245 $X2=0.655 $Y2=1.18
cc_5 VNB N_GATE_N_c_174_n 0.0169132f $X=-0.19 $Y=-0.245 $X2=0.625 $Y2=1.18
cc_6 VNB N_GATE_N_M1002_g 0.0224851f $X=-0.19 $Y=-0.245 $X2=0.705 $Y2=2.725
cc_7 VNB N_GATE_N_c_176_n 0.0275503f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_8 VNB N_GATE_N_c_177_n 0.0382281f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_GATE_N_c_178_n 0.00426637f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB GATE_N 0.0247185f $X=-0.19 $Y=-0.245 $X2=0.655 $Y2=1.345
cc_11 VNB N_GATE_N_c_180_n 0.0486359f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_242_130#_M1011_g 0.0143233f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.21
cc_13 VNB N_A_242_130#_c_219_n 0.0357786f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_242_130#_c_220_n 0.0167563f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_242_130#_c_221_n 0.0193752f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_242_130#_M1014_g 0.023268f $X=-0.19 $Y=-0.245 $X2=0.655 $Y2=1.51
cc_17 VNB N_A_242_130#_c_223_n 0.017846f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_242_130#_c_224_n 0.007537f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_242_130#_c_225_n 0.0154953f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_242_130#_c_226_n 0.00176681f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_242_130#_c_227_n 0.00167841f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_242_130#_c_228_n 0.0341125f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_242_130#_c_229_n 0.028882f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_242_130#_c_230_n 0.0104999f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_57_130#_c_367_n 0.0284726f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_57_130#_c_368_n 0.0130551f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_57_130#_M1019_g 0.0350086f $X=-0.19 $Y=-0.245 $X2=0.655 $Y2=1.345
cc_28 VNB N_A_57_130#_c_370_n 0.0307877f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_57_130#_c_371_n 0.0165451f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_57_130#_c_372_n 0.036193f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_349_481#_c_446_n 0.049797f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_349_481#_c_447_n 0.0152174f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_349_481#_M1004_g 0.0211807f $X=-0.19 $Y=-0.245 $X2=0.655 $Y2=1.345
cc_34 VNB N_A_349_481#_c_449_n 0.00819705f $X=-0.19 $Y=-0.245 $X2=0.655 $Y2=1.51
cc_35 VNB N_A_349_481#_c_450_n 0.0038358f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_349_481#_c_451_n 0.00756068f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_349_481#_c_452_n 0.0048873f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_349_481#_c_453_n 0.0014517f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_349_481#_c_454_n 0.00116594f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_349_481#_c_455_n 0.0447739f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_849_419#_M1008_g 0.0577416f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_849_419#_c_560_n 0.0193477f $X=-0.19 $Y=-0.245 $X2=0.655 $Y2=1.345
cc_43 VNB N_A_849_419#_M1012_g 0.0033143f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_849_419#_c_562_n 0.0101534f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=1.345
cc_45 VNB N_A_849_419#_M1009_g 0.0328955f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_849_419#_M1018_g 0.0067324f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_849_419#_c_565_n 0.0386657f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_849_419#_c_566_n 0.00833898f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_849_419#_c_567_n 0.0106787f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_849_419#_c_568_n 0.00842015f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_849_419#_c_569_n 0.0045782f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_849_419#_c_570_n 0.00480765f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_849_419#_c_571_n 2.88537e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_849_419#_c_572_n 0.00824041f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_849_419#_c_573_n 0.00442376f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_849_419#_c_574_n 0.00254859f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_663_481#_c_677_n 0.0021717f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_663_481#_c_678_n 0.00951232f $X=-0.19 $Y=-0.245 $X2=1.68 $Y2=1.345
cc_59 VNB N_A_663_481#_c_679_n 0.00437834f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_663_481#_c_680_n 0.00844279f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_A_663_481#_c_681_n 0.0307839f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_A_663_481#_c_682_n 2.95047e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_A_663_481#_c_683_n 0.0209056f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_VPWR_c_776_n 0.302998f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_Q_c_864_n 0.00911762f $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=1.345
cc_66 VNB N_VGND_c_884_n 0.0192378f $X=-0.19 $Y=-0.245 $X2=0.655 $Y2=1.345
cc_67 VNB N_VGND_c_885_n 4.89148e-19 $X=-0.19 $Y=-0.245 $X2=1.2 $Y2=1.345
cc_68 VNB N_VGND_c_886_n 0.00680918f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_VGND_c_887_n 0.0147016f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_VGND_c_888_n 0.0111284f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_VGND_c_889_n 0.0471788f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_VGND_c_890_n 0.0493572f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_VGND_c_891_n 0.0417359f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_VGND_c_892_n 0.0199105f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_VGND_c_893_n 0.0169228f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_VGND_c_894_n 0.0254935f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_VGND_c_895_n 0.00436214f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_VGND_c_896_n 0.00432412f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_VGND_c_897_n 0.00567425f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_VGND_c_898_n 0.384999f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VPB N_D_M1010_g 0.0563099f $X=-0.19 $Y=1.655 $X2=0.705 $Y2=2.725
cc_82 VPB N_GATE_N_M1002_g 0.0631246f $X=-0.19 $Y=1.655 $X2=0.705 $Y2=2.725
cc_83 VPB N_A_242_130#_M1011_g 0.068529f $X=-0.19 $Y=1.655 $X2=1.115 $Y2=1.21
cc_84 VPB N_A_242_130#_M1003_g 0.0195035f $X=-0.19 $Y=1.655 $X2=1.2 $Y2=1.345
cc_85 VPB N_A_242_130#_c_233_n 0.00984336f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_86 VPB N_A_242_130#_c_234_n 0.013192f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_87 VPB N_A_242_130#_c_235_n 0.00287821f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_88 VPB N_A_242_130#_c_236_n 0.0148188f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_89 VPB N_A_242_130#_c_237_n 0.0013623f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_90 VPB N_A_242_130#_c_238_n 4.79405e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_91 VPB N_A_242_130#_c_239_n 8.26269e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_92 VPB N_A_242_130#_c_240_n 0.0343217f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_93 VPB N_A_242_130#_c_230_n 0.00375492f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_94 VPB N_A_57_130#_M1015_g 0.0387345f $X=-0.19 $Y=1.655 $X2=1.115 $Y2=1.21
cc_95 VPB N_A_57_130#_c_374_n 0.0190315f $X=-0.19 $Y=1.655 $X2=0.655 $Y2=1.345
cc_96 VPB N_A_57_130#_c_375_n 0.0702846f $X=-0.19 $Y=1.655 $X2=1.68 $Y2=1.345
cc_97 VPB N_A_57_130#_c_376_n 0.0412951f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_98 VPB N_A_57_130#_c_377_n 0.0135949f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_99 VPB N_A_57_130#_c_372_n 0.00730654f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_100 VPB N_A_349_481#_M1016_g 0.0239155f $X=-0.19 $Y=1.655 $X2=1.115 $Y2=1.21
cc_101 VPB N_A_349_481#_c_457_n 0.0142734f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_102 VPB N_A_349_481#_c_458_n 0.00865373f $X=-0.19 $Y=1.655 $X2=1.68 $Y2=1.345
cc_103 VPB N_A_349_481#_c_459_n 0.0269118f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_104 VPB N_A_349_481#_c_460_n 0.0057335f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_105 VPB N_A_349_481#_c_453_n 0.0281985f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_106 VPB N_A_849_419#_M1013_g 0.0214578f $X=-0.19 $Y=1.655 $X2=1.115 $Y2=1.21
cc_107 VPB N_A_849_419#_M1012_g 0.0242146f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_108 VPB N_A_849_419#_M1018_g 0.0272177f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_109 VPB N_A_849_419#_c_578_n 0.0653335f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_110 VPB N_A_849_419#_c_565_n 0.00303978f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_111 VPB N_A_849_419#_c_580_n 0.00891742f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_112 VPB N_A_849_419#_c_581_n 0.0131452f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_113 VPB N_A_849_419#_c_570_n 0.00480765f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_114 VPB N_A_849_419#_c_571_n 0.00482704f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_115 VPB N_A_849_419#_c_572_n 0.00948869f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_116 VPB N_A_849_419#_c_574_n 0.00564441f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_117 VPB N_A_663_481#_M1000_g 0.0223718f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_118 VPB N_A_663_481#_c_685_n 0.00857277f $X=-0.19 $Y=1.655 $X2=0.655
+ $Y2=1.345
cc_119 VPB N_A_663_481#_c_677_n 0.00836224f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_120 VPB N_A_663_481#_c_681_n 0.00730964f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_121 VPB N_VPWR_c_777_n 0.00650519f $X=-0.19 $Y=1.655 $X2=0.655 $Y2=1.51
cc_122 VPB N_VPWR_c_778_n 0.00666604f $X=-0.19 $Y=1.655 $X2=1.2 $Y2=1.345
cc_123 VPB N_VPWR_c_779_n 0.0187917f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_124 VPB N_VPWR_c_780_n 0.0111025f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_125 VPB N_VPWR_c_781_n 0.0585137f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_126 VPB N_VPWR_c_782_n 0.023072f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_127 VPB N_VPWR_c_783_n 0.0047828f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_128 VPB N_VPWR_c_784_n 0.0350337f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_129 VPB N_VPWR_c_785_n 0.0459789f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_130 VPB N_VPWR_c_786_n 0.0188074f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_131 VPB N_VPWR_c_787_n 0.0167145f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_132 VPB N_VPWR_c_788_n 0.00497591f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_133 VPB N_VPWR_c_789_n 0.0329073f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_134 VPB N_VPWR_c_790_n 0.00564836f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_135 VPB N_VPWR_c_776_n 0.0920018f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_136 VPB N_Q_c_864_n 0.00409125f $X=-0.19 $Y=1.655 $X2=1.2 $Y2=1.345
cc_137 N_D_c_141_n N_GATE_N_c_174_n 0.0152635f $X=0.655 $Y=1.18 $X2=-0.19
+ $Y2=-0.245
cc_138 N_D_M1010_g N_GATE_N_M1002_g 0.0475023f $X=0.705 $Y=2.725 $X2=0 $Y2=0
cc_139 D N_GATE_N_M1002_g 0.0096594f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_140 D N_GATE_N_c_176_n 0.0210205f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_141 D N_GATE_N_c_178_n 0.00688774f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_142 N_D_c_140_n N_GATE_N_c_178_n 0.0185618f $X=0.655 $Y=1.345 $X2=0 $Y2=0
cc_143 D GATE_N 0.00514857f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_144 N_D_c_141_n GATE_N 3.61926e-19 $X=0.655 $Y=1.18 $X2=0 $Y2=0
cc_145 D N_A_242_130#_c_224_n 0.0481923f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_146 D N_A_242_130#_c_227_n 0.024173f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_147 D N_A_242_130#_c_228_n 0.00475445f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_148 N_D_M1010_g N_A_57_130#_c_370_n 0.00434712f $X=0.705 $Y=2.725 $X2=0 $Y2=0
cc_149 D N_A_57_130#_c_370_n 0.0220364f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_150 N_D_c_140_n N_A_57_130#_c_370_n 0.00356598f $X=0.655 $Y=1.345 $X2=0 $Y2=0
cc_151 N_D_c_141_n N_A_57_130#_c_370_n 0.00443646f $X=0.655 $Y=1.18 $X2=0 $Y2=0
cc_152 N_D_M1010_g N_A_57_130#_c_375_n 0.0257194f $X=0.705 $Y=2.725 $X2=0 $Y2=0
cc_153 N_D_M1010_g N_A_57_130#_c_376_n 0.0181134f $X=0.705 $Y=2.725 $X2=0 $Y2=0
cc_154 D N_A_57_130#_c_376_n 0.0949205f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_155 N_D_c_140_n N_A_57_130#_c_376_n 0.00105396f $X=0.655 $Y=1.345 $X2=0 $Y2=0
cc_156 D N_A_57_130#_c_371_n 2.97449e-19 $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_157 D N_A_57_130#_c_377_n 0.0112849f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_158 N_D_c_140_n N_A_57_130#_c_377_n 0.00352386f $X=0.655 $Y=1.345 $X2=0 $Y2=0
cc_159 N_D_M1010_g N_VPWR_c_777_n 0.00294295f $X=0.705 $Y=2.725 $X2=0 $Y2=0
cc_160 N_D_M1010_g N_VPWR_c_782_n 0.0053602f $X=0.705 $Y=2.725 $X2=0 $Y2=0
cc_161 N_D_M1010_g N_VPWR_c_776_n 0.0109701f $X=0.705 $Y=2.725 $X2=0 $Y2=0
cc_162 N_D_c_141_n N_VGND_c_884_n 0.0107779f $X=0.655 $Y=1.18 $X2=0 $Y2=0
cc_163 D N_VGND_c_900_n 0.0224578f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_164 N_D_c_140_n N_VGND_c_900_n 0.00294168f $X=0.655 $Y=1.345 $X2=0 $Y2=0
cc_165 N_D_c_141_n N_VGND_c_900_n 0.00272292f $X=0.655 $Y=1.18 $X2=0 $Y2=0
cc_166 N_D_c_141_n N_VGND_c_894_n 0.00334468f $X=0.655 $Y=1.18 $X2=0 $Y2=0
cc_167 N_D_c_141_n N_VGND_c_898_n 0.00388565f $X=0.655 $Y=1.18 $X2=0 $Y2=0
cc_168 N_GATE_N_c_177_n N_A_242_130#_c_220_n 0.0116784f $X=1.625 $Y=1.18 $X2=0
+ $Y2=0
cc_169 GATE_N N_A_242_130#_c_220_n 0.00790284f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_170 N_GATE_N_c_174_n N_A_242_130#_c_224_n 0.00300291f $X=1.135 $Y=1.18 $X2=0
+ $Y2=0
cc_171 N_GATE_N_c_176_n N_A_242_130#_c_224_n 0.00315043f $X=1.55 $Y=1.255 $X2=0
+ $Y2=0
cc_172 N_GATE_N_c_177_n N_A_242_130#_c_224_n 0.013037f $X=1.625 $Y=1.18 $X2=0
+ $Y2=0
cc_173 GATE_N N_A_242_130#_c_224_n 0.0626884f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_174 N_GATE_N_c_180_n N_A_242_130#_c_224_n 9.68147e-19 $X=1.715 $Y=0.36 $X2=0
+ $Y2=0
cc_175 N_GATE_N_M1002_g N_A_242_130#_c_233_n 2.93193e-19 $X=1.135 $Y=2.725 $X2=0
+ $Y2=0
cc_176 N_GATE_N_M1002_g N_A_242_130#_c_235_n 7.32615e-19 $X=1.135 $Y=2.725 $X2=0
+ $Y2=0
cc_177 N_GATE_N_c_177_n N_A_242_130#_c_227_n 0.00102553f $X=1.625 $Y=1.18 $X2=0
+ $Y2=0
cc_178 GATE_N N_A_242_130#_c_227_n 0.0217927f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_179 N_GATE_N_c_176_n N_A_242_130#_c_228_n 0.0116784f $X=1.55 $Y=1.255 $X2=0
+ $Y2=0
cc_180 N_GATE_N_M1002_g N_A_57_130#_c_376_n 0.0184334f $X=1.135 $Y=2.725 $X2=0
+ $Y2=0
cc_181 N_GATE_N_c_176_n N_A_57_130#_c_376_n 0.00235361f $X=1.55 $Y=1.255 $X2=0
+ $Y2=0
cc_182 N_GATE_N_M1002_g N_A_349_481#_c_458_n 0.00532598f $X=1.135 $Y=2.725 $X2=0
+ $Y2=0
cc_183 N_GATE_N_M1002_g N_A_349_481#_c_460_n 0.00496909f $X=1.135 $Y=2.725 $X2=0
+ $Y2=0
cc_184 GATE_N N_A_349_481#_c_450_n 0.0315731f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_185 N_GATE_N_c_180_n N_A_349_481#_c_450_n 7.80396e-19 $X=1.715 $Y=0.36 $X2=0
+ $Y2=0
cc_186 N_GATE_N_M1002_g N_VPWR_c_777_n 0.00255955f $X=1.135 $Y=2.725 $X2=0 $Y2=0
cc_187 N_GATE_N_M1002_g N_VPWR_c_784_n 0.0053602f $X=1.135 $Y=2.725 $X2=0 $Y2=0
cc_188 N_GATE_N_M1002_g N_VPWR_c_776_n 0.0111156f $X=1.135 $Y=2.725 $X2=0 $Y2=0
cc_189 N_GATE_N_c_174_n N_VGND_c_884_n 0.0038382f $X=1.135 $Y=1.18 $X2=0 $Y2=0
cc_190 GATE_N N_VGND_c_884_n 0.030657f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_191 N_GATE_N_c_174_n N_VGND_c_890_n 5.22141e-19 $X=1.135 $Y=1.18 $X2=0 $Y2=0
cc_192 GATE_N N_VGND_c_890_n 0.0760047f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_193 N_GATE_N_c_180_n N_VGND_c_890_n 0.00642834f $X=1.715 $Y=0.36 $X2=0 $Y2=0
cc_194 GATE_N N_VGND_c_898_n 0.0467157f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_195 N_GATE_N_c_180_n N_VGND_c_898_n 0.00965717f $X=1.715 $Y=0.36 $X2=0 $Y2=0
cc_196 N_A_242_130#_M1011_g N_A_57_130#_M1015_g 0.0178075f $X=2.085 $Y=2.725
+ $X2=0 $Y2=0
cc_197 N_A_242_130#_c_258_p N_A_57_130#_M1015_g 0.00294614f $X=2.22 $Y=2.905
+ $X2=0 $Y2=0
cc_198 N_A_242_130#_c_236_n N_A_57_130#_M1015_g 0.0126033f $X=3.705 $Y=2.46
+ $X2=0 $Y2=0
cc_199 N_A_242_130#_c_225_n N_A_57_130#_c_367_n 0.0158075f $X=3.705 $Y=1.08
+ $X2=0 $Y2=0
cc_200 N_A_242_130#_c_229_n N_A_57_130#_c_367_n 0.0370453f $X=3.72 $Y=1.08 $X2=0
+ $Y2=0
cc_201 N_A_242_130#_c_230_n N_A_57_130#_c_367_n 0.00145518f $X=3.835 $Y=1.915
+ $X2=0 $Y2=0
cc_202 N_A_242_130#_c_219_n N_A_57_130#_c_368_n 0.0143813f $X=2.765 $Y=0.84
+ $X2=0 $Y2=0
cc_203 N_A_242_130#_c_225_n N_A_57_130#_c_368_n 0.00783949f $X=3.705 $Y=1.08
+ $X2=0 $Y2=0
cc_204 N_A_242_130#_c_227_n N_A_57_130#_c_368_n 0.00177825f $X=2.175 $Y=0.985
+ $X2=0 $Y2=0
cc_205 N_A_242_130#_c_228_n N_A_57_130#_c_368_n 0.0099832f $X=2.175 $Y=0.985
+ $X2=0 $Y2=0
cc_206 N_A_242_130#_c_221_n N_A_57_130#_M1019_g 0.0234435f $X=2.84 $Y=0.765
+ $X2=0 $Y2=0
cc_207 N_A_242_130#_M1014_g N_A_57_130#_M1019_g 0.0370453f $X=3.63 $Y=0.445
+ $X2=0 $Y2=0
cc_208 N_A_242_130#_c_225_n N_A_57_130#_M1019_g 0.00815259f $X=3.705 $Y=1.08
+ $X2=0 $Y2=0
cc_209 N_A_242_130#_c_233_n N_A_57_130#_c_375_n 3.17626e-19 $X=1.35 $Y=2.56
+ $X2=0 $Y2=0
cc_210 N_A_242_130#_M1011_g N_A_57_130#_c_376_n 0.0148844f $X=2.085 $Y=2.725
+ $X2=0 $Y2=0
cc_211 N_A_242_130#_c_223_n N_A_57_130#_c_376_n 0.00125756f $X=2.175 $Y=1.49
+ $X2=0 $Y2=0
cc_212 N_A_242_130#_c_224_n N_A_57_130#_c_376_n 0.0051708f $X=2.025 $Y=0.92
+ $X2=0 $Y2=0
cc_213 N_A_242_130#_c_233_n N_A_57_130#_c_376_n 0.0113731f $X=1.35 $Y=2.56 $X2=0
+ $Y2=0
cc_214 N_A_242_130#_c_225_n N_A_57_130#_c_376_n 0.00924654f $X=3.705 $Y=1.08
+ $X2=0 $Y2=0
cc_215 N_A_242_130#_c_227_n N_A_57_130#_c_376_n 0.024655f $X=2.175 $Y=0.985
+ $X2=0 $Y2=0
cc_216 N_A_242_130#_M1011_g N_A_57_130#_c_412_n 0.00107563f $X=2.085 $Y=2.725
+ $X2=0 $Y2=0
cc_217 N_A_242_130#_c_223_n N_A_57_130#_c_412_n 5.46087e-19 $X=2.175 $Y=1.49
+ $X2=0 $Y2=0
cc_218 N_A_242_130#_c_225_n N_A_57_130#_c_412_n 0.0239682f $X=3.705 $Y=1.08
+ $X2=0 $Y2=0
cc_219 N_A_242_130#_c_227_n N_A_57_130#_c_412_n 0.00784252f $X=2.175 $Y=0.985
+ $X2=0 $Y2=0
cc_220 N_A_242_130#_M1011_g N_A_57_130#_c_372_n 0.0128672f $X=2.085 $Y=2.725
+ $X2=0 $Y2=0
cc_221 N_A_242_130#_c_223_n N_A_57_130#_c_372_n 0.0057122f $X=2.175 $Y=1.49
+ $X2=0 $Y2=0
cc_222 N_A_242_130#_c_234_n N_A_349_481#_M1011_s 0.00286504f $X=2.135 $Y=2.99
+ $X2=0 $Y2=0
cc_223 N_A_242_130#_c_236_n N_A_349_481#_M1016_g 0.0115575f $X=3.705 $Y=2.46
+ $X2=0 $Y2=0
cc_224 N_A_242_130#_c_239_n N_A_349_481#_M1016_g 9.77395e-19 $X=3.87 $Y=2.08
+ $X2=0 $Y2=0
cc_225 N_A_242_130#_c_240_n N_A_349_481#_M1016_g 0.0195964f $X=3.87 $Y=2.08
+ $X2=0 $Y2=0
cc_226 N_A_242_130#_c_225_n N_A_349_481#_c_446_n 8.19067e-19 $X=3.705 $Y=1.08
+ $X2=0 $Y2=0
cc_227 N_A_242_130#_c_238_n N_A_349_481#_c_446_n 2.42701e-19 $X=3.835 $Y=2.045
+ $X2=0 $Y2=0
cc_228 N_A_242_130#_c_240_n N_A_349_481#_c_446_n 0.0154481f $X=3.87 $Y=2.08
+ $X2=0 $Y2=0
cc_229 N_A_242_130#_c_229_n N_A_349_481#_c_446_n 0.0189872f $X=3.72 $Y=1.08
+ $X2=0 $Y2=0
cc_230 N_A_242_130#_c_230_n N_A_349_481#_c_446_n 0.0143116f $X=3.835 $Y=1.915
+ $X2=0 $Y2=0
cc_231 N_A_242_130#_c_225_n N_A_349_481#_c_447_n 0.00596708f $X=3.705 $Y=1.08
+ $X2=0 $Y2=0
cc_232 N_A_242_130#_M1014_g N_A_349_481#_M1004_g 0.0201243f $X=3.63 $Y=0.445
+ $X2=0 $Y2=0
cc_233 N_A_242_130#_c_236_n N_A_349_481#_c_457_n 0.00125196f $X=3.705 $Y=2.46
+ $X2=0 $Y2=0
cc_234 N_A_242_130#_M1011_g N_A_349_481#_c_458_n 0.00755395f $X=2.085 $Y=2.725
+ $X2=0 $Y2=0
cc_235 N_A_242_130#_c_233_n N_A_349_481#_c_458_n 0.0254545f $X=1.35 $Y=2.56
+ $X2=0 $Y2=0
cc_236 N_A_242_130#_c_234_n N_A_349_481#_c_458_n 0.0189554f $X=2.135 $Y=2.99
+ $X2=0 $Y2=0
cc_237 N_A_242_130#_c_237_n N_A_349_481#_c_458_n 0.00795389f $X=2.305 $Y=2.46
+ $X2=0 $Y2=0
cc_238 N_A_242_130#_M1011_g N_A_349_481#_c_459_n 0.0171055f $X=2.085 $Y=2.725
+ $X2=0 $Y2=0
cc_239 N_A_242_130#_c_236_n N_A_349_481#_c_459_n 0.0893352f $X=3.705 $Y=2.46
+ $X2=0 $Y2=0
cc_240 N_A_242_130#_c_237_n N_A_349_481#_c_459_n 0.0141853f $X=2.305 $Y=2.46
+ $X2=0 $Y2=0
cc_241 N_A_242_130#_c_238_n N_A_349_481#_c_459_n 0.0111889f $X=3.835 $Y=2.045
+ $X2=0 $Y2=0
cc_242 N_A_242_130#_c_240_n N_A_349_481#_c_459_n 5.90248e-19 $X=3.87 $Y=2.08
+ $X2=0 $Y2=0
cc_243 N_A_242_130#_c_219_n N_A_349_481#_c_451_n 0.00363137f $X=2.765 $Y=0.84
+ $X2=0 $Y2=0
cc_244 N_A_242_130#_c_221_n N_A_349_481#_c_451_n 0.00864507f $X=2.84 $Y=0.765
+ $X2=0 $Y2=0
cc_245 N_A_242_130#_M1014_g N_A_349_481#_c_451_n 0.0119373f $X=3.63 $Y=0.445
+ $X2=0 $Y2=0
cc_246 N_A_242_130#_c_225_n N_A_349_481#_c_451_n 0.0681241f $X=3.705 $Y=1.08
+ $X2=0 $Y2=0
cc_247 N_A_242_130#_c_226_n N_A_349_481#_c_451_n 0.0170154f $X=3.815 $Y=1.165
+ $X2=0 $Y2=0
cc_248 N_A_242_130#_c_229_n N_A_349_481#_c_451_n 0.00440581f $X=3.72 $Y=1.08
+ $X2=0 $Y2=0
cc_249 N_A_242_130#_c_219_n N_A_349_481#_c_452_n 0.0111978f $X=2.765 $Y=0.84
+ $X2=0 $Y2=0
cc_250 N_A_242_130#_c_225_n N_A_349_481#_c_452_n 0.0195335f $X=3.705 $Y=1.08
+ $X2=0 $Y2=0
cc_251 N_A_242_130#_c_227_n N_A_349_481#_c_452_n 4.23254e-19 $X=2.175 $Y=0.985
+ $X2=0 $Y2=0
cc_252 N_A_242_130#_c_225_n N_A_349_481#_c_496_n 0.0138767f $X=3.705 $Y=1.08
+ $X2=0 $Y2=0
cc_253 N_A_242_130#_c_240_n N_A_349_481#_c_496_n 4.17313e-19 $X=3.87 $Y=2.08
+ $X2=0 $Y2=0
cc_254 N_A_242_130#_c_230_n N_A_349_481#_c_496_n 0.0318393f $X=3.835 $Y=1.915
+ $X2=0 $Y2=0
cc_255 N_A_242_130#_c_238_n N_A_349_481#_c_453_n 5.25462e-19 $X=3.835 $Y=2.045
+ $X2=0 $Y2=0
cc_256 N_A_242_130#_c_240_n N_A_349_481#_c_453_n 0.0179739f $X=3.87 $Y=2.08
+ $X2=0 $Y2=0
cc_257 N_A_242_130#_c_230_n N_A_349_481#_c_453_n 0.00613434f $X=3.835 $Y=1.915
+ $X2=0 $Y2=0
cc_258 N_A_242_130#_M1014_g N_A_349_481#_c_454_n 6.85545e-19 $X=3.63 $Y=0.445
+ $X2=0 $Y2=0
cc_259 N_A_242_130#_c_226_n N_A_349_481#_c_454_n 0.00885499f $X=3.815 $Y=1.165
+ $X2=0 $Y2=0
cc_260 N_A_242_130#_c_229_n N_A_349_481#_c_454_n 6.91667e-19 $X=3.72 $Y=1.08
+ $X2=0 $Y2=0
cc_261 N_A_242_130#_c_226_n N_A_349_481#_c_455_n 0.002417f $X=3.815 $Y=1.165
+ $X2=0 $Y2=0
cc_262 N_A_242_130#_c_229_n N_A_349_481#_c_455_n 0.0210414f $X=3.72 $Y=1.08
+ $X2=0 $Y2=0
cc_263 N_A_242_130#_c_230_n N_A_349_481#_c_455_n 0.00708664f $X=3.835 $Y=1.915
+ $X2=0 $Y2=0
cc_264 N_A_242_130#_M1003_g N_A_849_419#_M1013_g 0.0199364f $X=3.78 $Y=2.615
+ $X2=0 $Y2=0
cc_265 N_A_242_130#_c_236_n N_A_849_419#_M1013_g 5.68128e-19 $X=3.705 $Y=2.46
+ $X2=0 $Y2=0
cc_266 N_A_242_130#_c_239_n N_A_849_419#_M1013_g 3.6538e-19 $X=3.87 $Y=2.08
+ $X2=0 $Y2=0
cc_267 N_A_242_130#_c_240_n N_A_849_419#_c_578_n 0.012872f $X=3.87 $Y=2.08 $X2=0
+ $Y2=0
cc_268 N_A_242_130#_c_236_n N_A_663_481#_M1016_d 0.00311814f $X=3.705 $Y=2.46
+ $X2=0 $Y2=0
cc_269 N_A_242_130#_M1003_g N_A_663_481#_c_685_n 0.0151308f $X=3.78 $Y=2.615
+ $X2=0 $Y2=0
cc_270 N_A_242_130#_c_236_n N_A_663_481#_c_685_n 0.0382176f $X=3.705 $Y=2.46
+ $X2=0 $Y2=0
cc_271 N_A_242_130#_c_240_n N_A_663_481#_c_685_n 0.00243308f $X=3.87 $Y=2.08
+ $X2=0 $Y2=0
cc_272 N_A_242_130#_M1014_g N_A_663_481#_c_692_n 0.00339307f $X=3.63 $Y=0.445
+ $X2=0 $Y2=0
cc_273 N_A_242_130#_M1003_g N_A_663_481#_c_677_n 0.00401791f $X=3.78 $Y=2.615
+ $X2=0 $Y2=0
cc_274 N_A_242_130#_c_236_n N_A_663_481#_c_677_n 0.0139234f $X=3.705 $Y=2.46
+ $X2=0 $Y2=0
cc_275 N_A_242_130#_c_238_n N_A_663_481#_c_677_n 0.0343923f $X=3.835 $Y=2.045
+ $X2=0 $Y2=0
cc_276 N_A_242_130#_c_240_n N_A_663_481#_c_677_n 0.00260809f $X=3.87 $Y=2.08
+ $X2=0 $Y2=0
cc_277 N_A_242_130#_c_230_n N_A_663_481#_c_677_n 0.0293968f $X=3.835 $Y=1.915
+ $X2=0 $Y2=0
cc_278 N_A_242_130#_c_230_n N_A_663_481#_c_698_n 0.0124554f $X=3.835 $Y=1.915
+ $X2=0 $Y2=0
cc_279 N_A_242_130#_c_234_n N_VPWR_M1011_d 0.00138006f $X=2.135 $Y=2.99 $X2=0
+ $Y2=0
cc_280 N_A_242_130#_c_258_p N_VPWR_M1011_d 0.00439327f $X=2.22 $Y=2.905 $X2=0
+ $Y2=0
cc_281 N_A_242_130#_c_236_n N_VPWR_M1011_d 0.00840917f $X=3.705 $Y=2.46 $X2=0
+ $Y2=0
cc_282 N_A_242_130#_c_235_n N_VPWR_c_777_n 0.00251363f $X=1.515 $Y=2.99 $X2=0
+ $Y2=0
cc_283 N_A_242_130#_M1011_g N_VPWR_c_778_n 0.00264791f $X=2.085 $Y=2.725 $X2=0
+ $Y2=0
cc_284 N_A_242_130#_c_234_n N_VPWR_c_778_n 0.0143348f $X=2.135 $Y=2.99 $X2=0
+ $Y2=0
cc_285 N_A_242_130#_c_258_p N_VPWR_c_778_n 0.0142172f $X=2.22 $Y=2.905 $X2=0
+ $Y2=0
cc_286 N_A_242_130#_c_236_n N_VPWR_c_778_n 0.0204744f $X=3.705 $Y=2.46 $X2=0
+ $Y2=0
cc_287 N_A_242_130#_M1011_g N_VPWR_c_784_n 0.00325872f $X=2.085 $Y=2.725 $X2=0
+ $Y2=0
cc_288 N_A_242_130#_c_234_n N_VPWR_c_784_n 0.0516455f $X=2.135 $Y=2.99 $X2=0
+ $Y2=0
cc_289 N_A_242_130#_c_235_n N_VPWR_c_784_n 0.021506f $X=1.515 $Y=2.99 $X2=0
+ $Y2=0
cc_290 N_A_242_130#_M1003_g N_VPWR_c_785_n 7.10185e-19 $X=3.78 $Y=2.615 $X2=0
+ $Y2=0
cc_291 N_A_242_130#_M1011_g N_VPWR_c_776_n 0.00623479f $X=2.085 $Y=2.725 $X2=0
+ $Y2=0
cc_292 N_A_242_130#_c_234_n N_VPWR_c_776_n 0.0292342f $X=2.135 $Y=2.99 $X2=0
+ $Y2=0
cc_293 N_A_242_130#_c_235_n N_VPWR_c_776_n 0.0116633f $X=1.515 $Y=2.99 $X2=0
+ $Y2=0
cc_294 N_A_242_130#_c_236_n N_VPWR_c_776_n 0.0258868f $X=3.705 $Y=2.46 $X2=0
+ $Y2=0
cc_295 N_A_242_130#_c_236_n A_591_481# 0.00183853f $X=3.705 $Y=2.46 $X2=-0.19
+ $Y2=-0.245
cc_296 N_A_242_130#_c_236_n A_771_481# 0.00183677f $X=3.705 $Y=2.46 $X2=-0.19
+ $Y2=-0.245
cc_297 N_A_242_130#_c_221_n N_VGND_c_885_n 0.00870097f $X=2.84 $Y=0.765 $X2=0
+ $Y2=0
cc_298 N_A_242_130#_M1014_g N_VGND_c_885_n 0.00187081f $X=3.63 $Y=0.445 $X2=0
+ $Y2=0
cc_299 N_A_242_130#_c_219_n N_VGND_c_890_n 7.47573e-19 $X=2.765 $Y=0.84 $X2=0
+ $Y2=0
cc_300 N_A_242_130#_c_220_n N_VGND_c_890_n 0.00299783f $X=2.34 $Y=0.84 $X2=0
+ $Y2=0
cc_301 N_A_242_130#_c_221_n N_VGND_c_890_n 0.00354752f $X=2.84 $Y=0.765 $X2=0
+ $Y2=0
cc_302 N_A_242_130#_M1014_g N_VGND_c_891_n 0.00426565f $X=3.63 $Y=0.445 $X2=0
+ $Y2=0
cc_303 N_A_242_130#_c_220_n N_VGND_c_898_n 0.00391593f $X=2.34 $Y=0.84 $X2=0
+ $Y2=0
cc_304 N_A_242_130#_c_221_n N_VGND_c_898_n 0.00559858f $X=2.84 $Y=0.765 $X2=0
+ $Y2=0
cc_305 N_A_242_130#_M1014_g N_VGND_c_898_n 0.00616897f $X=3.63 $Y=0.445 $X2=0
+ $Y2=0
cc_306 N_A_57_130#_c_367_n N_A_349_481#_c_447_n 0.0124615f $X=3.195 $Y=1.2 $X2=0
+ $Y2=0
cc_307 N_A_57_130#_c_412_n N_A_349_481#_c_447_n 0.00147234f $X=2.76 $Y=1.43
+ $X2=0 $Y2=0
cc_308 N_A_57_130#_c_372_n N_A_349_481#_c_447_n 0.0358085f $X=2.76 $Y=1.43 $X2=0
+ $Y2=0
cc_309 N_A_57_130#_M1015_g N_A_349_481#_c_457_n 0.0358085f $X=2.88 $Y=2.725
+ $X2=0 $Y2=0
cc_310 N_A_57_130#_M1015_g N_A_349_481#_c_459_n 0.0123288f $X=2.88 $Y=2.725
+ $X2=0 $Y2=0
cc_311 N_A_57_130#_c_374_n N_A_349_481#_c_459_n 0.00597251f $X=2.775 $Y=1.935
+ $X2=0 $Y2=0
cc_312 N_A_57_130#_c_376_n N_A_349_481#_c_459_n 0.045593f $X=2.595 $Y=1.757
+ $X2=0 $Y2=0
cc_313 N_A_57_130#_c_412_n N_A_349_481#_c_459_n 0.0240811f $X=2.76 $Y=1.43 $X2=0
+ $Y2=0
cc_314 N_A_57_130#_c_376_n N_A_349_481#_c_460_n 0.0205161f $X=2.595 $Y=1.757
+ $X2=0 $Y2=0
cc_315 N_A_57_130#_c_368_n N_A_349_481#_c_451_n 0.00154699f $X=2.955 $Y=1.2
+ $X2=0 $Y2=0
cc_316 N_A_57_130#_M1019_g N_A_349_481#_c_451_n 0.0111159f $X=3.27 $Y=0.445
+ $X2=0 $Y2=0
cc_317 N_A_57_130#_c_367_n N_A_349_481#_c_496_n 6.80333e-19 $X=3.195 $Y=1.2
+ $X2=0 $Y2=0
cc_318 N_A_57_130#_c_412_n N_A_349_481#_c_496_n 0.0181736f $X=2.76 $Y=1.43 $X2=0
+ $Y2=0
cc_319 N_A_57_130#_c_372_n N_A_349_481#_c_496_n 0.00239084f $X=2.76 $Y=1.43
+ $X2=0 $Y2=0
cc_320 N_A_57_130#_c_374_n N_A_349_481#_c_453_n 0.0358085f $X=2.775 $Y=1.935
+ $X2=0 $Y2=0
cc_321 N_A_57_130#_M1015_g N_A_663_481#_c_685_n 9.91921e-19 $X=2.88 $Y=2.725
+ $X2=0 $Y2=0
cc_322 N_A_57_130#_c_375_n N_VPWR_c_777_n 7.55893e-19 $X=0.49 $Y=2.55 $X2=0
+ $Y2=0
cc_323 N_A_57_130#_c_376_n N_VPWR_c_777_n 0.00723332f $X=2.595 $Y=1.757 $X2=0
+ $Y2=0
cc_324 N_A_57_130#_M1015_g N_VPWR_c_778_n 0.00848238f $X=2.88 $Y=2.725 $X2=0
+ $Y2=0
cc_325 N_A_57_130#_c_375_n N_VPWR_c_782_n 0.0307335f $X=0.49 $Y=2.55 $X2=0 $Y2=0
cc_326 N_A_57_130#_M1015_g N_VPWR_c_785_n 0.0053602f $X=2.88 $Y=2.725 $X2=0
+ $Y2=0
cc_327 N_A_57_130#_M1015_g N_VPWR_c_776_n 0.00612193f $X=2.88 $Y=2.725 $X2=0
+ $Y2=0
cc_328 N_A_57_130#_c_375_n N_VPWR_c_776_n 0.0185968f $X=0.49 $Y=2.55 $X2=0 $Y2=0
cc_329 N_A_57_130#_M1019_g N_VGND_c_885_n 0.00933457f $X=3.27 $Y=0.445 $X2=0
+ $Y2=0
cc_330 N_A_57_130#_M1019_g N_VGND_c_891_n 0.00354752f $X=3.27 $Y=0.445 $X2=0
+ $Y2=0
cc_331 N_A_57_130#_c_371_n N_VGND_c_894_n 0.0058201f $X=0.41 $Y=0.86 $X2=0 $Y2=0
cc_332 N_A_57_130#_M1019_g N_VGND_c_898_n 0.00404424f $X=3.27 $Y=0.445 $X2=0
+ $Y2=0
cc_333 N_A_57_130#_c_371_n N_VGND_c_898_n 0.00994318f $X=0.41 $Y=0.86 $X2=0
+ $Y2=0
cc_334 N_A_349_481#_M1004_g N_A_849_419#_M1008_g 0.0216861f $X=4.17 $Y=0.445
+ $X2=0 $Y2=0
cc_335 N_A_349_481#_c_449_n N_A_849_419#_M1008_g 0.00660924f $X=4.17 $Y=1.485
+ $X2=0 $Y2=0
cc_336 N_A_349_481#_c_454_n N_A_849_419#_M1008_g 0.00101405f $X=4.26 $Y=0.73
+ $X2=0 $Y2=0
cc_337 N_A_349_481#_c_455_n N_A_849_419#_M1008_g 0.0310152f $X=4.26 $Y=1.005
+ $X2=0 $Y2=0
cc_338 N_A_349_481#_c_446_n N_A_849_419#_c_572_n 0.00321344f $X=4.095 $Y=1.56
+ $X2=0 $Y2=0
cc_339 N_A_349_481#_c_451_n N_A_663_481#_M1014_d 0.00305317f $X=4.095 $Y=0.73
+ $X2=-0.19 $Y2=-0.245
cc_340 N_A_349_481#_M1016_g N_A_663_481#_c_685_n 0.0070696f $X=3.24 $Y=2.725
+ $X2=0 $Y2=0
cc_341 N_A_349_481#_M1004_g N_A_663_481#_c_692_n 0.0096768f $X=4.17 $Y=0.445
+ $X2=0 $Y2=0
cc_342 N_A_349_481#_c_451_n N_A_663_481#_c_692_n 0.0174644f $X=4.095 $Y=0.73
+ $X2=0 $Y2=0
cc_343 N_A_349_481#_c_454_n N_A_663_481#_c_692_n 0.0198687f $X=4.26 $Y=0.73
+ $X2=0 $Y2=0
cc_344 N_A_349_481#_c_455_n N_A_663_481#_c_692_n 7.16339e-19 $X=4.26 $Y=1.005
+ $X2=0 $Y2=0
cc_345 N_A_349_481#_c_446_n N_A_663_481#_c_677_n 0.00745226f $X=4.095 $Y=1.56
+ $X2=0 $Y2=0
cc_346 N_A_349_481#_c_449_n N_A_663_481#_c_677_n 8.10217e-19 $X=4.17 $Y=1.485
+ $X2=0 $Y2=0
cc_347 N_A_349_481#_c_454_n N_A_663_481#_c_678_n 0.008769f $X=4.26 $Y=0.73 $X2=0
+ $Y2=0
cc_348 N_A_349_481#_c_455_n N_A_663_481#_c_678_n 0.00488328f $X=4.26 $Y=1.005
+ $X2=0 $Y2=0
cc_349 N_A_349_481#_c_449_n N_A_663_481#_c_698_n 0.00370052f $X=4.17 $Y=1.485
+ $X2=0 $Y2=0
cc_350 N_A_349_481#_c_454_n N_A_663_481#_c_698_n 0.0139639f $X=4.26 $Y=0.73
+ $X2=0 $Y2=0
cc_351 N_A_349_481#_c_455_n N_A_663_481#_c_698_n 0.00544946f $X=4.26 $Y=1.005
+ $X2=0 $Y2=0
cc_352 N_A_349_481#_M1004_g N_A_663_481#_c_679_n 4.30596e-19 $X=4.17 $Y=0.445
+ $X2=0 $Y2=0
cc_353 N_A_349_481#_c_454_n N_A_663_481#_c_679_n 0.0331504f $X=4.26 $Y=0.73
+ $X2=0 $Y2=0
cc_354 N_A_349_481#_c_455_n N_A_663_481#_c_679_n 0.00458488f $X=4.26 $Y=1.005
+ $X2=0 $Y2=0
cc_355 N_A_349_481#_c_455_n N_A_663_481#_c_682_n 2.6958e-19 $X=4.26 $Y=1.005
+ $X2=0 $Y2=0
cc_356 N_A_349_481#_M1016_g N_VPWR_c_785_n 0.00501304f $X=3.24 $Y=2.725 $X2=0
+ $Y2=0
cc_357 N_A_349_481#_M1016_g N_VPWR_c_776_n 0.00647292f $X=3.24 $Y=2.725 $X2=0
+ $Y2=0
cc_358 N_A_349_481#_c_451_n N_VGND_M1006_d 0.00169923f $X=4.095 $Y=0.73 $X2=0
+ $Y2=0
cc_359 N_A_349_481#_c_451_n N_VGND_c_885_n 0.0160487f $X=4.095 $Y=0.73 $X2=0
+ $Y2=0
cc_360 N_A_349_481#_c_450_n N_VGND_c_890_n 0.0155308f $X=2.625 $Y=0.44 $X2=0
+ $Y2=0
cc_361 N_A_349_481#_c_451_n N_VGND_c_890_n 0.00241405f $X=4.095 $Y=0.73 $X2=0
+ $Y2=0
cc_362 N_A_349_481#_M1004_g N_VGND_c_891_n 0.00357877f $X=4.17 $Y=0.445 $X2=0
+ $Y2=0
cc_363 N_A_349_481#_c_451_n N_VGND_c_891_n 0.00812722f $X=4.095 $Y=0.73 $X2=0
+ $Y2=0
cc_364 N_A_349_481#_M1006_s N_VGND_c_898_n 0.0023132f $X=2.5 $Y=0.235 $X2=0
+ $Y2=0
cc_365 N_A_349_481#_M1004_g N_VGND_c_898_n 0.00590678f $X=4.17 $Y=0.445 $X2=0
+ $Y2=0
cc_366 N_A_349_481#_c_450_n N_VGND_c_898_n 0.0098703f $X=2.625 $Y=0.44 $X2=0
+ $Y2=0
cc_367 N_A_349_481#_c_451_n N_VGND_c_898_n 0.0210126f $X=4.095 $Y=0.73 $X2=0
+ $Y2=0
cc_368 N_A_349_481#_c_451_n A_669_47# 0.00169092f $X=4.095 $Y=0.73 $X2=-0.19
+ $Y2=-0.245
cc_369 N_A_349_481#_c_454_n A_849_47# 0.00137569f $X=4.26 $Y=0.73 $X2=-0.19
+ $Y2=-0.245
cc_370 N_A_849_419#_M1008_g N_A_663_481#_M1000_g 0.00169627f $X=4.71 $Y=0.445
+ $X2=0 $Y2=0
cc_371 N_A_849_419#_c_580_n N_A_663_481#_M1000_g 0.0154086f $X=5.415 $Y=1.705
+ $X2=0 $Y2=0
cc_372 N_A_849_419#_c_581_n N_A_663_481#_M1000_g 0.00431747f $X=5.55 $Y=1.825
+ $X2=0 $Y2=0
cc_373 N_A_849_419#_c_571_n N_A_663_481#_M1000_g 6.7383e-19 $X=4.65 $Y=1.74
+ $X2=0 $Y2=0
cc_374 N_A_849_419#_c_572_n N_A_663_481#_M1000_g 0.0125726f $X=4.65 $Y=1.74
+ $X2=0 $Y2=0
cc_375 N_A_849_419#_M1013_g N_A_663_481#_c_685_n 0.00775407f $X=4.32 $Y=2.615
+ $X2=0 $Y2=0
cc_376 N_A_849_419#_M1008_g N_A_663_481#_c_692_n 0.00844691f $X=4.71 $Y=0.445
+ $X2=0 $Y2=0
cc_377 N_A_849_419#_M1013_g N_A_663_481#_c_677_n 0.0176812f $X=4.32 $Y=2.615
+ $X2=0 $Y2=0
cc_378 N_A_849_419#_M1008_g N_A_663_481#_c_677_n 0.00222474f $X=4.71 $Y=0.445
+ $X2=0 $Y2=0
cc_379 N_A_849_419#_c_578_n N_A_663_481#_c_677_n 0.00937203f $X=4.65 $Y=2.095
+ $X2=0 $Y2=0
cc_380 N_A_849_419#_c_571_n N_A_663_481#_c_677_n 0.0450841f $X=4.65 $Y=1.74
+ $X2=0 $Y2=0
cc_381 N_A_849_419#_c_572_n N_A_663_481#_c_677_n 0.00204574f $X=4.65 $Y=1.74
+ $X2=0 $Y2=0
cc_382 N_A_849_419#_c_578_n N_A_663_481#_c_678_n 0.00418763f $X=4.65 $Y=2.095
+ $X2=0 $Y2=0
cc_383 N_A_849_419#_c_571_n N_A_663_481#_c_678_n 0.00952692f $X=4.65 $Y=1.74
+ $X2=0 $Y2=0
cc_384 N_A_849_419#_c_572_n N_A_663_481#_c_678_n 0.00328354f $X=4.65 $Y=1.74
+ $X2=0 $Y2=0
cc_385 N_A_849_419#_M1008_g N_A_663_481#_c_679_n 0.0185978f $X=4.71 $Y=0.445
+ $X2=0 $Y2=0
cc_386 N_A_849_419#_M1008_g N_A_663_481#_c_680_n 0.00259971f $X=4.71 $Y=0.445
+ $X2=0 $Y2=0
cc_387 N_A_849_419#_c_580_n N_A_663_481#_c_680_n 0.0393492f $X=5.415 $Y=1.705
+ $X2=0 $Y2=0
cc_388 N_A_849_419#_c_569_n N_A_663_481#_c_680_n 6.523e-19 $X=5.62 $Y=1.27 $X2=0
+ $Y2=0
cc_389 N_A_849_419#_c_571_n N_A_663_481#_c_680_n 0.00312872f $X=4.65 $Y=1.74
+ $X2=0 $Y2=0
cc_390 N_A_849_419#_c_572_n N_A_663_481#_c_680_n 8.22402e-19 $X=4.65 $Y=1.74
+ $X2=0 $Y2=0
cc_391 N_A_849_419#_c_573_n N_A_663_481#_c_680_n 0.00113769f $X=5.522 $Y=1.09
+ $X2=0 $Y2=0
cc_392 N_A_849_419#_c_574_n N_A_663_481#_c_680_n 0.0151873f $X=5.415 $Y=1.62
+ $X2=0 $Y2=0
cc_393 N_A_849_419#_M1008_g N_A_663_481#_c_681_n 0.0187415f $X=4.71 $Y=0.445
+ $X2=0 $Y2=0
cc_394 N_A_849_419#_c_565_n N_A_663_481#_c_681_n 0.00773195f $X=6.21 $Y=1.435
+ $X2=0 $Y2=0
cc_395 N_A_849_419#_c_580_n N_A_663_481#_c_681_n 0.00606335f $X=5.415 $Y=1.705
+ $X2=0 $Y2=0
cc_396 N_A_849_419#_c_569_n N_A_663_481#_c_681_n 0.00307271f $X=5.62 $Y=1.27
+ $X2=0 $Y2=0
cc_397 N_A_849_419#_c_573_n N_A_663_481#_c_681_n 0.00236959f $X=5.522 $Y=1.09
+ $X2=0 $Y2=0
cc_398 N_A_849_419#_c_574_n N_A_663_481#_c_681_n 0.00709019f $X=5.415 $Y=1.62
+ $X2=0 $Y2=0
cc_399 N_A_849_419#_M1008_g N_A_663_481#_c_682_n 0.00686132f $X=4.71 $Y=0.445
+ $X2=0 $Y2=0
cc_400 N_A_849_419#_c_571_n N_A_663_481#_c_682_n 0.0144338f $X=4.65 $Y=1.74
+ $X2=0 $Y2=0
cc_401 N_A_849_419#_c_572_n N_A_663_481#_c_682_n 8.49234e-19 $X=4.65 $Y=1.74
+ $X2=0 $Y2=0
cc_402 N_A_849_419#_M1008_g N_A_663_481#_c_683_n 0.0186243f $X=4.71 $Y=0.445
+ $X2=0 $Y2=0
cc_403 N_A_849_419#_c_569_n N_A_663_481#_c_683_n 0.00326401f $X=5.62 $Y=1.27
+ $X2=0 $Y2=0
cc_404 N_A_849_419#_c_573_n N_A_663_481#_c_683_n 0.0026681f $X=5.522 $Y=1.09
+ $X2=0 $Y2=0
cc_405 N_A_849_419#_c_580_n N_VPWR_M1013_d 0.00406504f $X=5.415 $Y=1.705 $X2=0
+ $Y2=0
cc_406 N_A_849_419#_M1013_g N_VPWR_c_824_n 0.00522606f $X=4.32 $Y=2.615 $X2=0
+ $Y2=0
cc_407 N_A_849_419#_c_578_n N_VPWR_c_824_n 0.00244917f $X=4.65 $Y=2.095 $X2=0
+ $Y2=0
cc_408 N_A_849_419#_c_580_n N_VPWR_c_824_n 0.015214f $X=5.415 $Y=1.705 $X2=0
+ $Y2=0
cc_409 N_A_849_419#_c_571_n N_VPWR_c_824_n 0.0189569f $X=4.65 $Y=1.74 $X2=0
+ $Y2=0
cc_410 N_A_849_419#_M1012_g N_VPWR_c_779_n 0.0074362f $X=6.285 $Y=2.465 $X2=0
+ $Y2=0
cc_411 N_A_849_419#_c_565_n N_VPWR_c_779_n 0.00733316f $X=6.21 $Y=1.435 $X2=0
+ $Y2=0
cc_412 N_A_849_419#_c_581_n N_VPWR_c_779_n 0.0835233f $X=5.55 $Y=1.825 $X2=0
+ $Y2=0
cc_413 N_A_849_419#_c_570_n N_VPWR_c_779_n 0.0183201f $X=6 $Y=1.435 $X2=0 $Y2=0
cc_414 N_A_849_419#_M1018_g N_VPWR_c_781_n 0.00737621f $X=6.715 $Y=2.465 $X2=0
+ $Y2=0
cc_415 N_A_849_419#_M1013_g N_VPWR_c_785_n 0.0031907f $X=4.32 $Y=2.615 $X2=0
+ $Y2=0
cc_416 N_A_849_419#_c_581_n N_VPWR_c_786_n 0.0118947f $X=5.55 $Y=1.825 $X2=0
+ $Y2=0
cc_417 N_A_849_419#_M1012_g N_VPWR_c_787_n 0.00585385f $X=6.285 $Y=2.465 $X2=0
+ $Y2=0
cc_418 N_A_849_419#_M1018_g N_VPWR_c_787_n 0.00585385f $X=6.715 $Y=2.465 $X2=0
+ $Y2=0
cc_419 N_A_849_419#_M1013_g N_VPWR_c_789_n 0.00410802f $X=4.32 $Y=2.615 $X2=0
+ $Y2=0
cc_420 N_A_849_419#_c_578_n N_VPWR_c_789_n 0.00283741f $X=4.65 $Y=2.095 $X2=0
+ $Y2=0
cc_421 N_A_849_419#_c_581_n N_VPWR_c_789_n 0.00165723f $X=5.55 $Y=1.825 $X2=0
+ $Y2=0
cc_422 N_A_849_419#_c_571_n N_VPWR_c_789_n 0.0211346f $X=4.65 $Y=1.74 $X2=0
+ $Y2=0
cc_423 N_A_849_419#_M1013_g N_VPWR_c_776_n 0.00302331f $X=4.32 $Y=2.615 $X2=0
+ $Y2=0
cc_424 N_A_849_419#_M1012_g N_VPWR_c_776_n 0.0118221f $X=6.285 $Y=2.465 $X2=0
+ $Y2=0
cc_425 N_A_849_419#_M1018_g N_VPWR_c_776_n 0.011478f $X=6.715 $Y=2.465 $X2=0
+ $Y2=0
cc_426 N_A_849_419#_c_581_n N_VPWR_c_776_n 0.0105077f $X=5.55 $Y=1.825 $X2=0
+ $Y2=0
cc_427 N_A_849_419#_c_560_n N_Q_c_864_n 0.00409767f $X=6.285 $Y=1.27 $X2=0 $Y2=0
cc_428 N_A_849_419#_c_562_n N_Q_c_864_n 0.016912f $X=6.64 $Y=1.495 $X2=0 $Y2=0
cc_429 N_A_849_419#_M1009_g N_Q_c_864_n 0.00770444f $X=6.715 $Y=0.74 $X2=0 $Y2=0
cc_430 N_A_849_419#_M1018_g N_Q_c_864_n 0.007731f $X=6.715 $Y=2.465 $X2=0 $Y2=0
cc_431 N_A_849_419#_c_566_n N_Q_c_864_n 0.00453207f $X=6.285 $Y=1.435 $X2=0
+ $Y2=0
cc_432 N_A_849_419#_c_581_n N_Q_c_864_n 7.56995e-19 $X=5.55 $Y=1.825 $X2=0 $Y2=0
cc_433 N_A_849_419#_c_569_n N_Q_c_864_n 0.00410486f $X=5.62 $Y=1.27 $X2=0 $Y2=0
cc_434 N_A_849_419#_c_570_n N_Q_c_864_n 0.0227521f $X=6 $Y=1.435 $X2=0 $Y2=0
cc_435 N_A_849_419#_c_574_n N_Q_c_864_n 0.00622403f $X=5.415 $Y=1.62 $X2=0 $Y2=0
cc_436 N_A_849_419#_M1008_g N_VGND_c_886_n 0.00859366f $X=4.71 $Y=0.445 $X2=0
+ $Y2=0
cc_437 N_A_849_419#_c_573_n N_VGND_c_886_n 0.00114103f $X=5.522 $Y=1.09 $X2=0
+ $Y2=0
cc_438 N_A_849_419#_c_560_n N_VGND_c_887_n 0.00518514f $X=6.285 $Y=1.27 $X2=0
+ $Y2=0
cc_439 N_A_849_419#_c_565_n N_VGND_c_887_n 0.00668546f $X=6.21 $Y=1.435 $X2=0
+ $Y2=0
cc_440 N_A_849_419#_c_568_n N_VGND_c_887_n 0.0626174f $X=5.47 $Y=0.42 $X2=0
+ $Y2=0
cc_441 N_A_849_419#_c_570_n N_VGND_c_887_n 0.0209182f $X=6 $Y=1.435 $X2=0 $Y2=0
cc_442 N_A_849_419#_M1009_g N_VGND_c_889_n 0.00721079f $X=6.715 $Y=0.74 $X2=0
+ $Y2=0
cc_443 N_A_849_419#_M1008_g N_VGND_c_891_n 0.00372849f $X=4.71 $Y=0.445 $X2=0
+ $Y2=0
cc_444 N_A_849_419#_c_568_n N_VGND_c_892_n 0.024071f $X=5.47 $Y=0.42 $X2=0 $Y2=0
cc_445 N_A_849_419#_c_560_n N_VGND_c_893_n 0.00503963f $X=6.285 $Y=1.27 $X2=0
+ $Y2=0
cc_446 N_A_849_419#_M1009_g N_VGND_c_893_n 0.00503963f $X=6.715 $Y=0.74 $X2=0
+ $Y2=0
cc_447 N_A_849_419#_M1005_d N_VGND_c_898_n 0.00249946f $X=5.33 $Y=0.235 $X2=0
+ $Y2=0
cc_448 N_A_849_419#_M1008_g N_VGND_c_898_n 0.00637924f $X=4.71 $Y=0.445 $X2=0
+ $Y2=0
cc_449 N_A_849_419#_c_560_n N_VGND_c_898_n 0.0103261f $X=6.285 $Y=1.27 $X2=0
+ $Y2=0
cc_450 N_A_849_419#_M1009_g N_VGND_c_898_n 0.010187f $X=6.715 $Y=0.74 $X2=0
+ $Y2=0
cc_451 N_A_849_419#_c_568_n N_VGND_c_898_n 0.0141126f $X=5.47 $Y=0.42 $X2=0
+ $Y2=0
cc_452 N_A_663_481#_c_685_n N_VPWR_c_778_n 0.0111063f $X=4.135 $Y=2.89 $X2=0
+ $Y2=0
cc_453 N_A_663_481#_M1000_g N_VPWR_c_779_n 0.00364492f $X=5.335 $Y=2.31 $X2=0
+ $Y2=0
cc_454 N_A_663_481#_c_685_n N_VPWR_c_785_n 0.0651921f $X=4.135 $Y=2.89 $X2=0
+ $Y2=0
cc_455 N_A_663_481#_M1000_g N_VPWR_c_786_n 0.00563421f $X=5.335 $Y=2.31 $X2=0
+ $Y2=0
cc_456 N_A_663_481#_M1000_g N_VPWR_c_789_n 0.00412713f $X=5.335 $Y=2.31 $X2=0
+ $Y2=0
cc_457 N_A_663_481#_c_685_n N_VPWR_c_789_n 0.031371f $X=4.135 $Y=2.89 $X2=0
+ $Y2=0
cc_458 N_A_663_481#_c_677_n N_VPWR_c_789_n 0.017252f $X=4.22 $Y=2.715 $X2=0
+ $Y2=0
cc_459 N_A_663_481#_M1000_g N_VPWR_c_776_n 0.00539454f $X=5.335 $Y=2.31 $X2=0
+ $Y2=0
cc_460 N_A_663_481#_c_685_n N_VPWR_c_776_n 0.0385629f $X=4.135 $Y=2.89 $X2=0
+ $Y2=0
cc_461 N_A_663_481#_c_685_n A_771_481# 0.00594588f $X=4.135 $Y=2.89 $X2=-0.19
+ $Y2=-0.245
cc_462 N_A_663_481#_c_677_n A_771_481# 0.00335448f $X=4.22 $Y=2.715 $X2=-0.19
+ $Y2=-0.245
cc_463 N_A_663_481#_c_692_n N_VGND_c_885_n 0.00695402f $X=4.605 $Y=0.365 $X2=0
+ $Y2=0
cc_464 N_A_663_481#_c_692_n N_VGND_c_886_n 0.0176361f $X=4.605 $Y=0.365 $X2=0
+ $Y2=0
cc_465 N_A_663_481#_c_679_n N_VGND_c_886_n 0.0441213f $X=4.69 $Y=1.26 $X2=0
+ $Y2=0
cc_466 N_A_663_481#_c_680_n N_VGND_c_886_n 0.0184252f $X=5.19 $Y=1.355 $X2=0
+ $Y2=0
cc_467 N_A_663_481#_c_681_n N_VGND_c_886_n 0.00365212f $X=5.19 $Y=1.355 $X2=0
+ $Y2=0
cc_468 N_A_663_481#_c_683_n N_VGND_c_886_n 0.0043333f $X=5.217 $Y=1.19 $X2=0
+ $Y2=0
cc_469 N_A_663_481#_c_683_n N_VGND_c_887_n 0.00316215f $X=5.217 $Y=1.19 $X2=0
+ $Y2=0
cc_470 N_A_663_481#_c_692_n N_VGND_c_891_n 0.0587343f $X=4.605 $Y=0.365 $X2=0
+ $Y2=0
cc_471 N_A_663_481#_c_683_n N_VGND_c_892_n 0.00585385f $X=5.217 $Y=1.19 $X2=0
+ $Y2=0
cc_472 N_A_663_481#_M1014_d N_VGND_c_898_n 0.00345569f $X=3.705 $Y=0.235 $X2=0
+ $Y2=0
cc_473 N_A_663_481#_c_692_n N_VGND_c_898_n 0.0360229f $X=4.605 $Y=0.365 $X2=0
+ $Y2=0
cc_474 N_A_663_481#_c_683_n N_VGND_c_898_n 0.0120995f $X=5.217 $Y=1.19 $X2=0
+ $Y2=0
cc_475 N_A_663_481#_c_692_n A_849_47# 0.0101442f $X=4.605 $Y=0.365 $X2=-0.19
+ $Y2=-0.245
cc_476 N_VPWR_c_776_n N_Q_M1012_s 0.0027574f $X=6.96 $Y=3.33 $X2=0 $Y2=0
cc_477 N_VPWR_c_779_n N_Q_c_864_n 0.00154184f $X=6.07 $Y=1.98 $X2=0 $Y2=0
cc_478 N_VPWR_c_781_n N_Q_c_864_n 0.00153983f $X=6.93 $Y=1.98 $X2=0 $Y2=0
cc_479 N_VPWR_c_787_n N_Q_c_864_n 0.0151136f $X=6.805 $Y=3.33 $X2=0 $Y2=0
cc_480 N_VPWR_c_776_n N_Q_c_864_n 0.0102248f $X=6.96 $Y=3.33 $X2=0 $Y2=0
cc_481 N_VPWR_c_781_n N_VGND_c_889_n 0.0107079f $X=6.93 $Y=1.98 $X2=0 $Y2=0
cc_482 N_Q_c_864_n N_VGND_c_887_n 0.00154184f $X=6.5 $Y=0.465 $X2=0 $Y2=0
cc_483 N_Q_c_864_n N_VGND_c_889_n 0.00307966f $X=6.5 $Y=0.465 $X2=0 $Y2=0
cc_484 N_Q_c_864_n N_VGND_c_893_n 0.0146631f $X=6.5 $Y=0.465 $X2=0 $Y2=0
cc_485 N_Q_c_864_n N_VGND_c_898_n 0.00999513f $X=6.5 $Y=0.465 $X2=0 $Y2=0
cc_486 N_VGND_c_898_n A_669_47# 0.00247238f $X=6.96 $Y=0 $X2=-0.19 $Y2=-0.245
cc_487 N_VGND_c_898_n A_849_47# 0.00313854f $X=6.96 $Y=0 $X2=-0.19 $Y2=-0.245
