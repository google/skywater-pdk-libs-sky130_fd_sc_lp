* File: sky130_fd_sc_lp__sleep_pargate_plv_7.pxi.spice
* Created: Wed Sep  2 10:37:57 2020
* 
x_PM_SKY130_FD_SC_LP__SLEEP_PARGATE_PLV_7%SLEEP N_SLEEP_c_31_n N_SLEEP_M1000_g
+ SLEEP SLEEP SLEEP SLEEP SLEEP N_SLEEP_c_33_n
+ PM_SKY130_FD_SC_LP__SLEEP_PARGATE_PLV_7%SLEEP
x_PM_SKY130_FD_SC_LP__SLEEP_PARGATE_PLV_7%VPWR N_VPWR_M1000_s VPWR N_VPWR_c_54_n
+ N_VPWR_c_55_n N_VPWR_c_56_n N_VPWR_c_57_n N_VPWR_c_58_n N_VPWR_c_59_n
+ N_VPWR_c_53_n PM_SKY130_FD_SC_LP__SLEEP_PARGATE_PLV_7%VPWR
x_PM_SKY130_FD_SC_LP__SLEEP_PARGATE_PLV_7%VIRTPWR N_VIRTPWR_M1000_d
+ N_VIRTPWR_c_110_n N_VIRTPWR_c_111_n VIRTPWR N_VIRTPWR_c_112_n
+ N_VIRTPWR_c_101_n N_VIRTPWR_c_102_n N_VIRTPWR_c_103_n N_VIRTPWR_c_104_n
+ N_VIRTPWR_c_113_n N_VIRTPWR_c_105_n N_VIRTPWR_c_115_n N_VIRTPWR_c_106_n
+ N_VIRTPWR_c_107_n N_VIRTPWR_c_108_n VIRTPWR N_VIRTPWR_c_109_n
+ PM_SKY130_FD_SC_LP__SLEEP_PARGATE_PLV_7%VIRTPWR
cc_1 noxref_1 SLEEP 0.0599664f $X=-0.19 $Y=-0.007 $X2=8.315 $Y2=0.84
cc_2 noxref_1 N_VPWR_c_53_n 0.677152f $X=-0.19 $Y=-0.007 $X2=0 $Y2=0
cc_3 noxref_1 N_VIRTPWR_c_101_n 0.0262405f $X=-0.19 $Y=-0.007 $X2=8.52 $Y2=1.985
cc_4 noxref_1 N_VIRTPWR_c_102_n 0.0262405f $X=-0.19 $Y=-0.007 $X2=0 $Y2=0
cc_5 noxref_1 N_VIRTPWR_c_103_n 0.0262405f $X=-0.19 $Y=-0.007 $X2=0 $Y2=0
cc_6 noxref_1 N_VIRTPWR_c_104_n 0.0270802f $X=-0.19 $Y=-0.007 $X2=0 $Y2=0
cc_7 noxref_1 N_VIRTPWR_c_105_n 0.0836651f $X=-0.19 $Y=-0.007 $X2=0 $Y2=0
cc_8 noxref_1 N_VIRTPWR_c_106_n 0.0786895f $X=-0.19 $Y=-0.007 $X2=0 $Y2=0
cc_9 noxref_1 N_VIRTPWR_c_107_n 0.038478f $X=-0.19 $Y=-0.007 $X2=0 $Y2=0
cc_10 noxref_1 N_VIRTPWR_c_108_n 0.038478f $X=-0.19 $Y=-0.007 $X2=0 $Y2=0
cc_11 noxref_1 N_VIRTPWR_c_109_n 0.038478f $X=-0.19 $Y=-0.007 $X2=0 $Y2=0
cc_12 VPB N_SLEEP_c_31_n 0.0516733f $X=-0.19 $Y=1.655 $X2=8.17 $Y2=2.755
cc_13 VPB SLEEP 0.030975f $X=-0.19 $Y=1.655 $X2=8.315 $Y2=0.84
cc_14 VPB N_SLEEP_c_33_n 0.107893f $X=-0.19 $Y=1.655 $X2=8.42 $Y2=1.985
cc_15 VPB N_VPWR_c_54_n 0.115615f $X=-0.19 $Y=1.655 $X2=8.52 $Y2=0.925
cc_16 VPB N_VPWR_c_55_n 0.0107573f $X=-0.19 $Y=1.655 $X2=8.52 $Y2=1.665
cc_17 VPB N_VPWR_c_56_n 0.00806873f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_18 VPB N_VPWR_c_57_n 0.00806873f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_19 VPB N_VPWR_c_58_n 0.00806873f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_20 VPB N_VPWR_c_59_n 0.00806873f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_21 VPB N_VPWR_c_53_n 0.168806f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_22 VPB N_VIRTPWR_c_110_n 0.0130323f $X=-0.19 $Y=1.655 $X2=8.377 $Y2=2.68
cc_23 VPB N_VIRTPWR_c_111_n 0.0357155f $X=-0.19 $Y=1.655 $X2=8.315 $Y2=1.95
cc_24 VPB N_VIRTPWR_c_112_n 0.15875f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_25 VPB N_VIRTPWR_c_113_n 0.0329627f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_26 VPB N_VIRTPWR_c_105_n 0.0405705f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_27 VPB N_VIRTPWR_c_115_n 0.0130323f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_28 VPB N_VIRTPWR_c_106_n 0.0404102f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_29 N_SLEEP_c_31_n N_VPWR_c_54_n 0.011857f $X=8.17 $Y=2.755 $X2=0 $Y2=0
cc_30 SLEEP N_VPWR_c_54_n 0.0112305f $X=8.315 $Y=0.84 $X2=0 $Y2=0
cc_31 N_SLEEP_c_33_n N_VPWR_c_54_n 0.00525497f $X=8.42 $Y=1.985 $X2=0 $Y2=0
cc_32 N_SLEEP_c_31_n N_VPWR_c_55_n 0.00302781f $X=8.17 $Y=2.755 $X2=0 $Y2=0
cc_33 SLEEP N_VPWR_c_59_n 0.0033926f $X=8.315 $Y=0.84 $X2=0 $Y2=0
cc_34 N_SLEEP_c_31_n N_VPWR_c_53_n 0.0125423f $X=8.17 $Y=2.755 $X2=0 $Y2=0
cc_35 SLEEP N_VPWR_c_53_n 0.108262f $X=8.315 $Y=0.84 $X2=0 $Y2=0
cc_36 N_SLEEP_c_33_n N_VPWR_c_53_n 0.0112731f $X=8.42 $Y=1.985 $X2=0 $Y2=0
cc_37 N_SLEEP_c_31_n N_VIRTPWR_c_110_n 0.0158929f $X=8.17 $Y=2.755 $X2=0 $Y2=0
cc_38 N_SLEEP_c_31_n N_VIRTPWR_c_111_n 0.00259154f $X=8.17 $Y=2.755 $X2=0 $Y2=0
cc_39 N_SLEEP_c_31_n N_VIRTPWR_c_101_n 0.00927999f $X=8.17 $Y=2.755 $X2=0 $Y2=0
cc_40 N_SLEEP_c_31_n N_VIRTPWR_c_102_n 0.00927999f $X=8.17 $Y=2.755 $X2=0 $Y2=0
cc_41 N_SLEEP_c_31_n N_VIRTPWR_c_103_n 0.00927999f $X=8.17 $Y=2.755 $X2=0 $Y2=0
cc_42 N_SLEEP_c_31_n N_VIRTPWR_c_104_n 0.00957695f $X=8.17 $Y=2.755 $X2=0 $Y2=0
cc_43 N_SLEEP_c_31_n N_VIRTPWR_c_113_n 0.00576677f $X=8.17 $Y=2.755 $X2=0 $Y2=0
cc_44 SLEEP N_VIRTPWR_c_113_n 0.0165417f $X=8.315 $Y=0.84 $X2=0 $Y2=0
cc_45 N_SLEEP_c_31_n N_VIRTPWR_c_105_n 0.0037323f $X=8.17 $Y=2.755 $X2=0 $Y2=0
cc_46 SLEEP N_VIRTPWR_c_105_n 0.0123629f $X=8.315 $Y=0.84 $X2=0 $Y2=0
cc_47 N_SLEEP_c_31_n N_VIRTPWR_c_106_n 0.00224979f $X=8.17 $Y=2.755 $X2=0 $Y2=0
cc_48 N_VPWR_c_54_n N_VIRTPWR_c_110_n 0.267892f $X=7.785 $Y=2.54 $X2=0 $Y2=0
cc_49 N_VPWR_c_55_n N_VIRTPWR_c_110_n 0.00538617f $X=1.545 $Y=2.54 $X2=0 $Y2=0
cc_50 N_VPWR_c_53_n N_VIRTPWR_c_110_n 0.00611837f $X=7.775 $Y=2.54 $X2=0 $Y2=0
cc_51 N_VPWR_c_56_n N_VIRTPWR_c_112_n 0.00538893f $X=3.09 $Y=2.54 $X2=0 $Y2=0
cc_52 N_VPWR_c_57_n N_VIRTPWR_c_112_n 0.00538893f $X=4.645 $Y=2.54 $X2=0 $Y2=0
cc_53 N_VPWR_c_58_n N_VIRTPWR_c_112_n 0.00538893f $X=6.2 $Y=2.54 $X2=0 $Y2=0
cc_54 N_VPWR_c_59_n N_VIRTPWR_c_112_n 0.00538617f $X=7.775 $Y=2.54 $X2=0 $Y2=0
cc_55 N_VPWR_c_53_n N_VIRTPWR_c_112_n 0.0186573f $X=7.775 $Y=2.54 $X2=0 $Y2=0
cc_56 N_VPWR_c_54_n N_VIRTPWR_c_101_n 0.0138562f $X=7.785 $Y=2.54 $X2=0 $Y2=0
cc_57 N_VPWR_c_53_n N_VIRTPWR_c_101_n 0.123829f $X=7.775 $Y=2.54 $X2=0 $Y2=0
cc_58 N_VPWR_c_54_n N_VIRTPWR_c_102_n 0.0138562f $X=7.785 $Y=2.54 $X2=0 $Y2=0
cc_59 N_VPWR_c_53_n N_VIRTPWR_c_102_n 0.123829f $X=7.775 $Y=2.54 $X2=0 $Y2=0
cc_60 N_VPWR_c_54_n N_VIRTPWR_c_103_n 0.0138562f $X=7.785 $Y=2.54 $X2=0 $Y2=0
cc_61 N_VPWR_c_53_n N_VIRTPWR_c_103_n 0.123829f $X=7.775 $Y=2.54 $X2=0 $Y2=0
cc_62 N_VPWR_c_54_n N_VIRTPWR_c_104_n 0.0142996f $X=7.785 $Y=2.54 $X2=0 $Y2=0
cc_63 N_VPWR_c_53_n N_VIRTPWR_c_104_n 0.127311f $X=7.775 $Y=2.54 $X2=0 $Y2=0
cc_64 N_VPWR_c_54_n N_VIRTPWR_c_105_n 0.00290716f $X=7.785 $Y=2.54 $X2=0 $Y2=0
cc_65 N_VPWR_c_59_n N_VIRTPWR_c_105_n 0.0256157f $X=7.775 $Y=2.54 $X2=0 $Y2=0
cc_66 N_VPWR_c_53_n N_VIRTPWR_c_105_n 0.227442f $X=7.775 $Y=2.54 $X2=0 $Y2=0
cc_67 N_VPWR_c_53_n N_VIRTPWR_c_115_n 0.00787277f $X=7.775 $Y=2.54 $X2=0 $Y2=0
cc_68 N_VPWR_c_54_n N_VIRTPWR_c_106_n 0.00285709f $X=7.785 $Y=2.54 $X2=0 $Y2=0
cc_69 N_VPWR_c_55_n N_VIRTPWR_c_106_n 0.0256157f $X=1.545 $Y=2.54 $X2=0 $Y2=0
cc_70 N_VPWR_c_53_n N_VIRTPWR_c_106_n 0.212348f $X=7.775 $Y=2.54 $X2=0 $Y2=0
cc_71 N_VPWR_c_54_n N_VIRTPWR_c_107_n 0.00424894f $X=7.785 $Y=2.54 $X2=0 $Y2=0
cc_72 N_VPWR_c_56_n N_VIRTPWR_c_107_n 0.0256093f $X=3.09 $Y=2.54 $X2=0 $Y2=0
cc_73 N_VPWR_c_53_n N_VIRTPWR_c_107_n 0.110096f $X=7.775 $Y=2.54 $X2=0 $Y2=0
cc_74 N_VPWR_c_54_n N_VIRTPWR_c_108_n 0.00424894f $X=7.785 $Y=2.54 $X2=0 $Y2=0
cc_75 N_VPWR_c_57_n N_VIRTPWR_c_108_n 0.0256093f $X=4.645 $Y=2.54 $X2=0 $Y2=0
cc_76 N_VPWR_c_53_n N_VIRTPWR_c_108_n 0.110096f $X=7.775 $Y=2.54 $X2=0 $Y2=0
cc_77 N_VPWR_c_54_n N_VIRTPWR_c_109_n 0.00424894f $X=7.785 $Y=2.54 $X2=0 $Y2=0
cc_78 N_VPWR_c_58_n N_VIRTPWR_c_109_n 0.0256093f $X=6.2 $Y=2.54 $X2=0 $Y2=0
cc_79 N_VPWR_c_53_n N_VIRTPWR_c_109_n 0.110096f $X=7.775 $Y=2.54 $X2=0 $Y2=0
