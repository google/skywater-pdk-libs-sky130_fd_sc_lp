* File: sky130_fd_sc_lp__or4bb_lp.pxi.spice
* Created: Fri Aug 28 11:26:57 2020
* 
x_PM_SKY130_FD_SC_LP__OR4BB_LP%A_86_21# N_A_86_21#_M1013_d N_A_86_21#_M1004_d
+ N_A_86_21#_M1019_d N_A_86_21#_M1012_g N_A_86_21#_c_157_n N_A_86_21#_c_158_n
+ N_A_86_21#_M1002_g N_A_86_21#_M1009_g N_A_86_21#_c_160_n N_A_86_21#_c_161_n
+ N_A_86_21#_c_162_n N_A_86_21#_c_163_n N_A_86_21#_c_164_n N_A_86_21#_c_165_n
+ N_A_86_21#_c_166_n N_A_86_21#_c_196_p N_A_86_21#_c_167_n N_A_86_21#_c_168_n
+ N_A_86_21#_c_169_n N_A_86_21#_c_170_n N_A_86_21#_c_171_n N_A_86_21#_c_172_n
+ N_A_86_21#_c_173_n N_A_86_21#_c_174_n PM_SKY130_FD_SC_LP__OR4BB_LP%A_86_21#
x_PM_SKY130_FD_SC_LP__OR4BB_LP%C_N N_C_N_c_291_n N_C_N_M1015_g N_C_N_M1000_g
+ N_C_N_c_292_n N_C_N_c_293_n N_C_N_c_294_n N_C_N_M1017_g N_C_N_c_295_n
+ N_C_N_c_296_n C_N N_C_N_c_298_n PM_SKY130_FD_SC_LP__OR4BB_LP%C_N
x_PM_SKY130_FD_SC_LP__OR4BB_LP%A_318_409# N_A_318_409#_M1017_d
+ N_A_318_409#_M1000_d N_A_318_409#_c_348_n N_A_318_409#_c_349_n
+ N_A_318_409#_c_363_n N_A_318_409#_M1014_g N_A_318_409#_c_350_n
+ N_A_318_409#_M1016_g N_A_318_409#_c_352_n N_A_318_409#_c_353_n
+ N_A_318_409#_M1008_g N_A_318_409#_c_355_n N_A_318_409#_c_356_n
+ N_A_318_409#_c_357_n N_A_318_409#_c_358_n N_A_318_409#_c_366_n
+ N_A_318_409#_c_367_n N_A_318_409#_c_359_n N_A_318_409#_c_368_n
+ N_A_318_409#_c_425_n N_A_318_409#_c_360_n N_A_318_409#_c_369_n
+ N_A_318_409#_c_370_n N_A_318_409#_c_371_n N_A_318_409#_c_372_n
+ PM_SKY130_FD_SC_LP__OR4BB_LP%A_318_409#
x_PM_SKY130_FD_SC_LP__OR4BB_LP%A_654_355# N_A_654_355#_M1006_d
+ N_A_654_355#_M1001_d N_A_654_355#_M1019_g N_A_654_355#_c_488_n
+ N_A_654_355#_c_489_n N_A_654_355#_c_500_n N_A_654_355#_c_501_n
+ N_A_654_355#_c_490_n N_A_654_355#_M1010_g N_A_654_355#_c_491_n
+ N_A_654_355#_c_492_n N_A_654_355#_c_493_n N_A_654_355#_M1004_g
+ N_A_654_355#_c_502_n N_A_654_355#_c_494_n N_A_654_355#_c_503_n
+ N_A_654_355#_c_504_n N_A_654_355#_c_495_n N_A_654_355#_c_506_n
+ N_A_654_355#_c_507_n N_A_654_355#_c_508_n N_A_654_355#_c_509_n
+ N_A_654_355#_c_496_n PM_SKY130_FD_SC_LP__OR4BB_LP%A_654_355#
x_PM_SKY130_FD_SC_LP__OR4BB_LP%B N_B_c_603_n N_B_M1007_g N_B_c_604_n N_B_c_605_n
+ N_B_c_606_n N_B_c_607_n N_B_c_608_n N_B_M1005_g N_B_M1011_g N_B_c_609_n B
+ PM_SKY130_FD_SC_LP__OR4BB_LP%B
x_PM_SKY130_FD_SC_LP__OR4BB_LP%A N_A_M1013_g N_A_c_665_n N_A_c_666_n N_A_M1020_g
+ N_A_M1018_g A N_A_c_669_n N_A_c_670_n PM_SKY130_FD_SC_LP__OR4BB_LP%A
x_PM_SKY130_FD_SC_LP__OR4BB_LP%D_N N_D_N_c_730_n N_D_N_M1001_g N_D_N_M1003_g
+ N_D_N_M1006_g D_N D_N PM_SKY130_FD_SC_LP__OR4BB_LP%D_N
x_PM_SKY130_FD_SC_LP__OR4BB_LP%X N_X_M1012_s N_X_M1009_s X X X X X X X
+ N_X_c_768_n X PM_SKY130_FD_SC_LP__OR4BB_LP%X
x_PM_SKY130_FD_SC_LP__OR4BB_LP%VPWR N_VPWR_M1009_d N_VPWR_M1020_d N_VPWR_c_791_n
+ N_VPWR_c_792_n VPWR N_VPWR_c_793_n N_VPWR_c_794_n N_VPWR_c_795_n
+ N_VPWR_c_790_n N_VPWR_c_797_n N_VPWR_c_798_n PM_SKY130_FD_SC_LP__OR4BB_LP%VPWR
x_PM_SKY130_FD_SC_LP__OR4BB_LP%A_505_400# N_A_505_400#_M1014_s
+ N_A_505_400#_M1011_s N_A_505_400#_c_848_n N_A_505_400#_c_849_n
+ PM_SKY130_FD_SC_LP__OR4BB_LP%A_505_400#
x_PM_SKY130_FD_SC_LP__OR4BB_LP%VGND N_VGND_M1002_d N_VGND_M1008_d N_VGND_M1005_d
+ N_VGND_M1003_s N_VGND_c_884_n N_VGND_c_885_n N_VGND_c_886_n N_VGND_c_887_n
+ N_VGND_c_888_n N_VGND_c_889_n N_VGND_c_890_n VGND N_VGND_c_891_n
+ N_VGND_c_892_n N_VGND_c_893_n N_VGND_c_894_n N_VGND_c_895_n N_VGND_c_896_n
+ N_VGND_c_897_n PM_SKY130_FD_SC_LP__OR4BB_LP%VGND
x_PM_SKY130_FD_SC_LP__OR4BB_LP%A_476_125# N_A_476_125#_M1013_s
+ N_A_476_125#_M1018_d N_A_476_125#_c_972_n N_A_476_125#_c_973_n
+ N_A_476_125#_c_982_n N_A_476_125#_c_1010_n N_A_476_125#_c_974_n
+ N_A_476_125#_c_975_n N_A_476_125#_c_976_n N_A_476_125#_c_977_n
+ N_A_476_125#_c_985_n N_A_476_125#_c_986_n N_A_476_125#_c_978_n
+ N_A_476_125#_c_979_n N_A_476_125#_c_980_n
+ PM_SKY130_FD_SC_LP__OR4BB_LP%A_476_125#
cc_1 VNB N_A_86_21#_M1012_g 0.0357312f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=0.445
cc_2 VNB N_A_86_21#_c_157_n 0.0125553f $X=-0.19 $Y=-0.245 $X2=0.79 $Y2=1.2
cc_3 VNB N_A_86_21#_c_158_n 0.0124933f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=1.2
cc_4 VNB N_A_86_21#_M1002_g 0.0349044f $X=-0.19 $Y=-0.245 $X2=0.865 $Y2=0.445
cc_5 VNB N_A_86_21#_c_160_n 0.0136741f $X=-0.19 $Y=-0.245 $X2=0.96 $Y2=1.2
cc_6 VNB N_A_86_21#_c_161_n 0.00228944f $X=-0.19 $Y=-0.245 $X2=0.96 $Y2=1.795
cc_7 VNB N_A_86_21#_c_162_n 0.0222452f $X=-0.19 $Y=-0.245 $X2=1.775 $Y2=1.21
cc_8 VNB N_A_86_21#_c_163_n 0.00795158f $X=-0.19 $Y=-0.245 $X2=1.86 $Y2=1.125
cc_9 VNB N_A_86_21#_c_164_n 0.0235143f $X=-0.19 $Y=-0.245 $X2=2.87 $Y2=0.86
cc_10 VNB N_A_86_21#_c_165_n 0.00360548f $X=-0.19 $Y=-0.245 $X2=1.945 $Y2=0.86
cc_11 VNB N_A_86_21#_c_166_n 0.00277677f $X=-0.19 $Y=-0.245 $X2=3.035 $Y2=0.945
cc_12 VNB N_A_86_21#_c_167_n 0.00784971f $X=-0.19 $Y=-0.245 $X2=3.495 $Y2=1.2
cc_13 VNB N_A_86_21#_c_168_n 0.00455286f $X=-0.19 $Y=-0.245 $X2=3.2 $Y2=1.2
cc_14 VNB N_A_86_21#_c_169_n 0.00789736f $X=-0.19 $Y=-0.245 $X2=3.66 $Y2=2.145
cc_15 VNB N_A_86_21#_c_170_n 0.00542636f $X=-0.19 $Y=-0.245 $X2=4.17 $Y2=1.2
cc_16 VNB N_A_86_21#_c_171_n 0.00180932f $X=-0.19 $Y=-0.245 $X2=0.965 $Y2=1.29
cc_17 VNB N_A_86_21#_c_172_n 0.0305017f $X=-0.19 $Y=-0.245 $X2=0.965 $Y2=1.29
cc_18 VNB N_A_86_21#_c_173_n 0.00296709f $X=-0.19 $Y=-0.245 $X2=3.66 $Y2=1.2
cc_19 VNB N_A_86_21#_c_174_n 0.00857527f $X=-0.19 $Y=-0.245 $X2=4.615 $Y2=0.835
cc_20 VNB N_C_N_c_291_n 0.0137164f $X=-0.19 $Y=-0.245 $X2=2.895 $Y2=0.625
cc_21 VNB N_C_N_c_292_n 0.00875756f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_C_N_c_293_n 0.00877538f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_C_N_c_294_n 0.0182972f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.125
cc_24 VNB N_C_N_c_295_n 0.0358686f $X=-0.19 $Y=-0.245 $X2=0.79 $Y2=1.2
cc_25 VNB N_C_N_c_296_n 0.0073149f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=1.2
cc_26 VNB C_N 0.00929242f $X=-0.19 $Y=-0.245 $X2=0.865 $Y2=1.125
cc_27 VNB N_C_N_c_298_n 0.0220212f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_318_409#_c_348_n 0.0147889f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_318_409#_c_349_n 0.0205262f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_318_409#_c_350_n 0.0155871f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_318_409#_M1016_g 0.0261989f $X=-0.19 $Y=-0.245 $X2=0.865 $Y2=1.125
cc_32 VNB N_A_318_409#_c_352_n 0.0136208f $X=-0.19 $Y=-0.245 $X2=0.865 $Y2=0.445
cc_33 VNB N_A_318_409#_c_353_n 0.0285773f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_318_409#_M1008_g 0.0222523f $X=-0.19 $Y=-0.245 $X2=0.935 $Y2=2.545
cc_35 VNB N_A_318_409#_c_355_n 0.00505023f $X=-0.19 $Y=-0.245 $X2=0.96 $Y2=1.2
cc_36 VNB N_A_318_409#_c_356_n 0.00873682f $X=-0.19 $Y=-0.245 $X2=1.775 $Y2=1.21
cc_37 VNB N_A_318_409#_c_357_n 0.0125506f $X=-0.19 $Y=-0.245 $X2=1.13 $Y2=1.21
cc_38 VNB N_A_318_409#_c_358_n 0.00182737f $X=-0.19 $Y=-0.245 $X2=1.86 $Y2=0.945
cc_39 VNB N_A_318_409#_c_359_n 6.72053e-19 $X=-0.19 $Y=-0.245 $X2=3.495 $Y2=1.2
cc_40 VNB N_A_318_409#_c_360_n 0.0137618f $X=-0.19 $Y=-0.245 $X2=3.825 $Y2=1.2
cc_41 VNB N_A_654_355#_c_488_n 0.0135884f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=0.445
cc_42 VNB N_A_654_355#_c_489_n 0.00637342f $X=-0.19 $Y=-0.245 $X2=0.505
+ $Y2=0.445
cc_43 VNB N_A_654_355#_c_490_n 0.0117728f $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=1.2
cc_44 VNB N_A_654_355#_c_491_n 0.0309594f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_654_355#_c_492_n 0.0196125f $X=-0.19 $Y=-0.245 $X2=0.935 $Y2=1.795
cc_46 VNB N_A_654_355#_c_493_n 0.0121942f $X=-0.19 $Y=-0.245 $X2=0.935 $Y2=2.545
cc_47 VNB N_A_654_355#_c_494_n 0.00438508f $X=-0.19 $Y=-0.245 $X2=0.96 $Y2=1.795
cc_48 VNB N_A_654_355#_c_495_n 0.0468372f $X=-0.19 $Y=-0.245 $X2=1.945 $Y2=0.86
cc_49 VNB N_A_654_355#_c_496_n 0.0209565f $X=-0.19 $Y=-0.245 $X2=0.965 $Y2=1.29
cc_50 VNB N_B_c_603_n 0.0125783f $X=-0.19 $Y=-0.245 $X2=2.895 $Y2=0.625
cc_51 VNB N_B_c_604_n 0.0353161f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_B_c_605_n 0.0202579f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_B_c_606_n 0.0196419f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_B_c_607_n 0.0104464f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_B_c_608_n 0.0138046f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.125
cc_56 VNB N_B_c_609_n 0.00535423f $X=-0.19 $Y=-0.245 $X2=0.865 $Y2=0.445
cc_57 VNB B 0.0028724f $X=-0.19 $Y=-0.245 $X2=0.865 $Y2=0.445
cc_58 VNB N_A_M1013_g 0.0498548f $X=-0.19 $Y=-0.245 $X2=3.52 $Y2=2
cc_59 VNB N_A_c_665_n 0.220075f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_c_666_n 0.012806f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_A_M1020_g 0.00250726f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_A_M1018_g 0.0568541f $X=-0.19 $Y=-0.245 $X2=0.79 $Y2=1.2
cc_63 VNB N_A_c_669_n 0.0339248f $X=-0.19 $Y=-0.245 $X2=0.865 $Y2=0.445
cc_64 VNB N_A_c_670_n 0.00689105f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_D_N_c_730_n 0.0768845f $X=-0.19 $Y=-0.245 $X2=2.895 $Y2=0.625
cc_66 VNB N_D_N_M1001_g 6.32853e-19 $X=-0.19 $Y=-0.245 $X2=3.52 $Y2=2
cc_67 VNB N_D_N_M1003_g 0.0349851f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_D_N_M1006_g 0.0367157f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=0.445
cc_69 VNB D_N 0.00191571f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB X 0.0510816f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_X_c_768_n 0.0126766f $X=-0.19 $Y=-0.245 $X2=3.66 $Y2=1.285
cc_72 VNB N_VPWR_c_790_n 0.302998f $X=-0.19 $Y=-0.245 $X2=1.86 $Y2=1.125
cc_73 VNB N_VGND_c_884_n 4.89148e-19 $X=-0.19 $Y=-0.245 $X2=0.58 $Y2=1.2
cc_74 VNB N_VGND_c_885_n 0.0183781f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_VGND_c_886_n 0.0280391f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_VGND_c_887_n 0.00891349f $X=-0.19 $Y=-0.245 $X2=0.96 $Y2=1.2
cc_77 VNB N_VGND_c_888_n 0.00957833f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_VGND_c_889_n 0.0675139f $X=-0.19 $Y=-0.245 $X2=1.86 $Y2=0.945
cc_79 VNB N_VGND_c_890_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=1.86 $Y2=1.125
cc_80 VNB N_VGND_c_891_n 0.0271715f $X=-0.19 $Y=-0.245 $X2=3.035 $Y2=0.945
cc_81 VNB N_VGND_c_892_n 0.0386067f $X=-0.19 $Y=-0.245 $X2=3.825 $Y2=1.2
cc_82 VNB N_VGND_c_893_n 0.0268694f $X=-0.19 $Y=-0.245 $X2=4.17 $Y2=1.2
cc_83 VNB N_VGND_c_894_n 0.364089f $X=-0.19 $Y=-0.245 $X2=0.96 $Y2=1.29
cc_84 VNB N_VGND_c_895_n 0.00436868f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_VGND_c_896_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_VGND_c_897_n 0.00513431f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_A_476_125#_c_972_n 0.00890684f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_A_476_125#_c_973_n 0.00613306f $X=-0.19 $Y=-0.245 $X2=0.505
+ $Y2=0.445
cc_89 VNB N_A_476_125#_c_974_n 0.00249415f $X=-0.19 $Y=-0.245 $X2=0.865
+ $Y2=1.125
cc_90 VNB N_A_476_125#_c_975_n 0.020174f $X=-0.19 $Y=-0.245 $X2=0.865 $Y2=0.445
cc_91 VNB N_A_476_125#_c_976_n 3.79193e-19 $X=-0.19 $Y=-0.245 $X2=0.865
+ $Y2=0.445
cc_92 VNB N_A_476_125#_c_977_n 0.00174095f $X=-0.19 $Y=-0.245 $X2=0.935
+ $Y2=1.795
cc_93 VNB N_A_476_125#_c_978_n 0.00798392f $X=-0.19 $Y=-0.245 $X2=0.96 $Y2=1.275
cc_94 VNB N_A_476_125#_c_979_n 0.00798776f $X=-0.19 $Y=-0.245 $X2=0.96 $Y2=1.625
cc_95 VNB N_A_476_125#_c_980_n 0.017413f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_96 VPB N_A_86_21#_M1009_g 0.035148f $X=-0.19 $Y=1.655 $X2=0.935 $Y2=2.545
cc_97 VPB N_A_86_21#_c_161_n 0.0131801f $X=-0.19 $Y=1.655 $X2=0.96 $Y2=1.795
cc_98 VPB N_A_86_21#_c_169_n 0.00272191f $X=-0.19 $Y=1.655 $X2=3.66 $Y2=2.145
cc_99 VPB N_A_86_21#_c_171_n 6.60545e-19 $X=-0.19 $Y=1.655 $X2=0.965 $Y2=1.29
cc_100 VPB N_C_N_M1000_g 0.0342252f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_101 VPB N_C_N_c_298_n 0.0162683f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_102 VPB N_A_318_409#_c_348_n 0.0141725f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_103 VPB N_A_318_409#_c_349_n 0.00565056f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_104 VPB N_A_318_409#_c_363_n 0.0234518f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_105 VPB N_A_318_409#_c_355_n 0.00457817f $X=-0.19 $Y=1.655 $X2=0.96 $Y2=1.2
cc_106 VPB N_A_318_409#_c_356_n 0.00719818f $X=-0.19 $Y=1.655 $X2=1.775 $Y2=1.21
cc_107 VPB N_A_318_409#_c_366_n 0.00219754f $X=-0.19 $Y=1.655 $X2=2.87 $Y2=0.86
cc_108 VPB N_A_318_409#_c_367_n 0.00408807f $X=-0.19 $Y=1.655 $X2=1.945 $Y2=0.86
cc_109 VPB N_A_318_409#_c_368_n 0.0164873f $X=-0.19 $Y=1.655 $X2=3.66 $Y2=2.145
cc_110 VPB N_A_318_409#_c_369_n 0.00410959f $X=-0.19 $Y=1.655 $X2=0.965 $Y2=1.29
cc_111 VPB N_A_318_409#_c_370_n 0.00367154f $X=-0.19 $Y=1.655 $X2=0.965 $Y2=1.29
cc_112 VPB N_A_318_409#_c_371_n 0.0269825f $X=-0.19 $Y=1.655 $X2=3.035 $Y2=0.835
cc_113 VPB N_A_318_409#_c_372_n 0.0500643f $X=-0.19 $Y=1.655 $X2=4.615 $Y2=0.835
cc_114 VPB N_A_654_355#_M1019_g 0.00618134f $X=-0.19 $Y=1.655 $X2=0.505
+ $Y2=1.125
cc_115 VPB N_A_654_355#_c_488_n 0.0248346f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=0.445
cc_116 VPB N_A_654_355#_c_489_n 0.00458038f $X=-0.19 $Y=1.655 $X2=0.505
+ $Y2=0.445
cc_117 VPB N_A_654_355#_c_500_n 0.0664844f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_118 VPB N_A_654_355#_c_501_n 0.0163736f $X=-0.19 $Y=1.655 $X2=0.79 $Y2=1.2
cc_119 VPB N_A_654_355#_c_502_n 0.0317113f $X=-0.19 $Y=1.655 $X2=0.96 $Y2=1.625
cc_120 VPB N_A_654_355#_c_503_n 0.00357627f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_121 VPB N_A_654_355#_c_504_n 0.0274462f $X=-0.19 $Y=1.655 $X2=1.86 $Y2=0.945
cc_122 VPB N_A_654_355#_c_495_n 0.0215179f $X=-0.19 $Y=1.655 $X2=1.945 $Y2=0.86
cc_123 VPB N_A_654_355#_c_506_n 0.0369839f $X=-0.19 $Y=1.655 $X2=3.495 $Y2=1.2
cc_124 VPB N_A_654_355#_c_507_n 0.00810489f $X=-0.19 $Y=1.655 $X2=3.66 $Y2=1.285
cc_125 VPB N_A_654_355#_c_508_n 0.0156464f $X=-0.19 $Y=1.655 $X2=3.66 $Y2=2.145
cc_126 VPB N_A_654_355#_c_509_n 0.0187087f $X=-0.19 $Y=1.655 $X2=3.825 $Y2=1.2
cc_127 VPB N_B_c_606_n 0.0100626f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_128 VPB N_B_c_607_n 0.0361057f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_129 VPB N_B_M1011_g 0.0248071f $X=-0.19 $Y=1.655 $X2=0.58 $Y2=1.2
cc_130 VPB B 0.00222787f $X=-0.19 $Y=1.655 $X2=0.865 $Y2=0.445
cc_131 VPB N_A_M1020_g 0.0262042f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_132 VPB N_D_N_c_730_n 0.0156098f $X=-0.19 $Y=1.655 $X2=2.895 $Y2=0.625
cc_133 VPB N_D_N_M1001_g 0.0305528f $X=-0.19 $Y=1.655 $X2=3.52 $Y2=2
cc_134 VPB D_N 0.00283076f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_135 VPB X 0.0341876f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_136 VPB X 0.0538654f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_137 VPB N_VPWR_c_791_n 0.00177638f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_138 VPB N_VPWR_c_792_n 4.89148e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_139 VPB N_VPWR_c_793_n 0.0278297f $X=-0.19 $Y=1.655 $X2=0.865 $Y2=0.445
cc_140 VPB N_VPWR_c_794_n 0.112284f $X=-0.19 $Y=1.655 $X2=0.935 $Y2=2.545
cc_141 VPB N_VPWR_c_795_n 0.0299095f $X=-0.19 $Y=1.655 $X2=1.86 $Y2=0.945
cc_142 VPB N_VPWR_c_790_n 0.0889423f $X=-0.19 $Y=1.655 $X2=1.86 $Y2=1.125
cc_143 VPB N_VPWR_c_797_n 0.00497896f $X=-0.19 $Y=1.655 $X2=3.035 $Y2=0.945
cc_144 VPB N_VPWR_c_798_n 0.00436768f $X=-0.19 $Y=1.655 $X2=3.2 $Y2=1.2
cc_145 VPB N_A_505_400#_c_848_n 0.0253175f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_146 VPB N_A_505_400#_c_849_n 0.00782961f $X=-0.19 $Y=1.655 $X2=0.505
+ $Y2=0.445
cc_147 VPB N_A_476_125#_c_973_n 0.00115015f $X=-0.19 $Y=1.655 $X2=0.505
+ $Y2=0.445
cc_148 VPB N_A_476_125#_c_982_n 0.00870189f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_149 VPB N_A_476_125#_c_974_n 0.0159976f $X=-0.19 $Y=1.655 $X2=0.865 $Y2=1.125
cc_150 VPB N_A_476_125#_c_977_n 0.00136576f $X=-0.19 $Y=1.655 $X2=0.935
+ $Y2=1.795
cc_151 VPB N_A_476_125#_c_985_n 0.00838226f $X=-0.19 $Y=1.655 $X2=0.935
+ $Y2=2.545
cc_152 VPB N_A_476_125#_c_986_n 2.51035e-19 $X=-0.19 $Y=1.655 $X2=0.935
+ $Y2=2.545
cc_153 VPB N_A_476_125#_c_978_n 0.00133865f $X=-0.19 $Y=1.655 $X2=0.96 $Y2=1.275
cc_154 N_A_86_21#_M1002_g N_C_N_c_291_n 0.0189395f $X=0.865 $Y=0.445 $X2=-0.19
+ $Y2=-0.245
cc_155 N_A_86_21#_c_162_n N_C_N_c_293_n 0.00150396f $X=1.775 $Y=1.21 $X2=0 $Y2=0
cc_156 N_A_86_21#_M1002_g N_C_N_c_295_n 0.00365984f $X=0.865 $Y=0.445 $X2=0
+ $Y2=0
cc_157 N_A_86_21#_c_160_n N_C_N_c_295_n 0.00658013f $X=0.96 $Y=1.2 $X2=0 $Y2=0
cc_158 N_A_86_21#_c_162_n N_C_N_c_295_n 0.0140586f $X=1.775 $Y=1.21 $X2=0 $Y2=0
cc_159 N_A_86_21#_c_163_n N_C_N_c_295_n 0.00723204f $X=1.86 $Y=1.125 $X2=0 $Y2=0
cc_160 N_A_86_21#_c_171_n N_C_N_c_295_n 4.97623e-19 $X=0.965 $Y=1.29 $X2=0 $Y2=0
cc_161 N_A_86_21#_c_165_n N_C_N_c_296_n 0.0051689f $X=1.945 $Y=0.86 $X2=0 $Y2=0
cc_162 N_A_86_21#_c_162_n C_N 0.0282442f $X=1.775 $Y=1.21 $X2=0 $Y2=0
cc_163 N_A_86_21#_c_171_n C_N 0.0165746f $X=0.965 $Y=1.29 $X2=0 $Y2=0
cc_164 N_A_86_21#_c_172_n C_N 0.0010193f $X=0.965 $Y=1.29 $X2=0 $Y2=0
cc_165 N_A_86_21#_M1009_g N_C_N_c_298_n 0.0312205f $X=0.935 $Y=2.545 $X2=0 $Y2=0
cc_166 N_A_86_21#_c_162_n N_C_N_c_298_n 0.00356525f $X=1.775 $Y=1.21 $X2=0 $Y2=0
cc_167 N_A_86_21#_c_171_n N_C_N_c_298_n 0.00120485f $X=0.965 $Y=1.29 $X2=0 $Y2=0
cc_168 N_A_86_21#_c_172_n N_C_N_c_298_n 0.0199797f $X=0.965 $Y=1.29 $X2=0 $Y2=0
cc_169 N_A_86_21#_c_169_n N_A_318_409#_c_350_n 0.00670572f $X=3.66 $Y=2.145
+ $X2=0 $Y2=0
cc_170 N_A_86_21#_c_166_n N_A_318_409#_M1016_g 0.00621342f $X=3.035 $Y=0.945
+ $X2=0 $Y2=0
cc_171 N_A_86_21#_c_196_p N_A_318_409#_M1016_g 0.00389259f $X=3.035 $Y=1.115
+ $X2=0 $Y2=0
cc_172 N_A_86_21#_c_167_n N_A_318_409#_M1016_g 0.0124196f $X=3.495 $Y=1.2 $X2=0
+ $Y2=0
cc_173 N_A_86_21#_c_168_n N_A_318_409#_M1016_g 0.0044825f $X=3.2 $Y=1.2 $X2=0
+ $Y2=0
cc_174 N_A_86_21#_c_169_n N_A_318_409#_M1016_g 0.00225434f $X=3.66 $Y=2.145
+ $X2=0 $Y2=0
cc_175 N_A_86_21#_c_167_n N_A_318_409#_c_352_n 0.00110828f $X=3.495 $Y=1.2 $X2=0
+ $Y2=0
cc_176 N_A_86_21#_c_169_n N_A_318_409#_c_352_n 0.0125278f $X=3.66 $Y=2.145 $X2=0
+ $Y2=0
cc_177 N_A_86_21#_c_168_n N_A_318_409#_c_353_n 0.0128431f $X=3.2 $Y=1.2 $X2=0
+ $Y2=0
cc_178 N_A_86_21#_c_166_n N_A_318_409#_M1008_g 9.46627e-19 $X=3.035 $Y=0.945
+ $X2=0 $Y2=0
cc_179 N_A_86_21#_c_196_p N_A_318_409#_M1008_g 8.46384e-19 $X=3.035 $Y=1.115
+ $X2=0 $Y2=0
cc_180 N_A_86_21#_c_169_n N_A_318_409#_M1008_g 0.0023254f $X=3.66 $Y=2.145 $X2=0
+ $Y2=0
cc_181 N_A_86_21#_c_173_n N_A_318_409#_M1008_g 0.012533f $X=3.66 $Y=1.2 $X2=0
+ $Y2=0
cc_182 N_A_86_21#_c_168_n N_A_318_409#_c_355_n 0.00107259f $X=3.2 $Y=1.2 $X2=0
+ $Y2=0
cc_183 N_A_86_21#_c_169_n N_A_318_409#_c_355_n 0.00203754f $X=3.66 $Y=2.145
+ $X2=0 $Y2=0
cc_184 N_A_86_21#_M1012_g N_A_318_409#_c_356_n 0.00329838f $X=0.505 $Y=0.445
+ $X2=0 $Y2=0
cc_185 N_A_86_21#_c_157_n N_A_318_409#_c_356_n 0.0056593f $X=0.79 $Y=1.2 $X2=0
+ $Y2=0
cc_186 N_A_86_21#_c_158_n N_A_318_409#_c_356_n 0.00401358f $X=0.58 $Y=1.2 $X2=0
+ $Y2=0
cc_187 N_A_86_21#_M1002_g N_A_318_409#_c_356_n 0.00380893f $X=0.865 $Y=0.445
+ $X2=0 $Y2=0
cc_188 N_A_86_21#_M1009_g N_A_318_409#_c_356_n 0.00675352f $X=0.935 $Y=2.545
+ $X2=0 $Y2=0
cc_189 N_A_86_21#_c_171_n N_A_318_409#_c_356_n 0.0478287f $X=0.965 $Y=1.29 $X2=0
+ $Y2=0
cc_190 N_A_86_21#_c_172_n N_A_318_409#_c_356_n 0.0125413f $X=0.965 $Y=1.29 $X2=0
+ $Y2=0
cc_191 N_A_86_21#_c_157_n N_A_318_409#_c_357_n 8.29573e-19 $X=0.79 $Y=1.2 $X2=0
+ $Y2=0
cc_192 N_A_86_21#_M1002_g N_A_318_409#_c_357_n 0.0138432f $X=0.865 $Y=0.445
+ $X2=0 $Y2=0
cc_193 N_A_86_21#_c_160_n N_A_318_409#_c_357_n 0.00130612f $X=0.96 $Y=1.2 $X2=0
+ $Y2=0
cc_194 N_A_86_21#_c_162_n N_A_318_409#_c_357_n 0.0349229f $X=1.775 $Y=1.21 $X2=0
+ $Y2=0
cc_195 N_A_86_21#_c_165_n N_A_318_409#_c_357_n 0.0144687f $X=1.945 $Y=0.86 $X2=0
+ $Y2=0
cc_196 N_A_86_21#_c_171_n N_A_318_409#_c_357_n 0.0206963f $X=0.965 $Y=1.29 $X2=0
+ $Y2=0
cc_197 N_A_86_21#_M1012_g N_A_318_409#_c_358_n 0.00592256f $X=0.505 $Y=0.445
+ $X2=0 $Y2=0
cc_198 N_A_86_21#_c_162_n N_A_318_409#_c_360_n 0.00452428f $X=1.775 $Y=1.21
+ $X2=0 $Y2=0
cc_199 N_A_86_21#_c_164_n N_A_318_409#_c_360_n 0.0064714f $X=2.87 $Y=0.86 $X2=0
+ $Y2=0
cc_200 N_A_86_21#_c_165_n N_A_318_409#_c_360_n 0.0128789f $X=1.945 $Y=0.86 $X2=0
+ $Y2=0
cc_201 N_A_86_21#_M1009_g N_A_318_409#_c_369_n 0.0213822f $X=0.935 $Y=2.545
+ $X2=0 $Y2=0
cc_202 N_A_86_21#_c_161_n N_A_318_409#_c_369_n 8.2121e-19 $X=0.96 $Y=1.795 $X2=0
+ $Y2=0
cc_203 N_A_86_21#_c_171_n N_A_318_409#_c_369_n 0.0200865f $X=0.965 $Y=1.29 $X2=0
+ $Y2=0
cc_204 N_A_86_21#_M1009_g N_A_318_409#_c_370_n 0.00292253f $X=0.935 $Y=2.545
+ $X2=0 $Y2=0
cc_205 N_A_86_21#_c_161_n N_A_318_409#_c_370_n 4.76756e-19 $X=0.96 $Y=1.795
+ $X2=0 $Y2=0
cc_206 N_A_86_21#_M1009_g N_A_318_409#_c_371_n 7.06436e-19 $X=0.935 $Y=2.545
+ $X2=0 $Y2=0
cc_207 N_A_86_21#_c_169_n N_A_654_355#_M1019_g 0.00618603f $X=3.66 $Y=2.145
+ $X2=0 $Y2=0
cc_208 N_A_86_21#_c_169_n N_A_654_355#_c_488_n 0.01746f $X=3.66 $Y=2.145 $X2=0
+ $Y2=0
cc_209 N_A_86_21#_c_170_n N_A_654_355#_c_488_n 0.00340128f $X=4.17 $Y=1.2 $X2=0
+ $Y2=0
cc_210 N_A_86_21#_c_167_n N_A_654_355#_c_489_n 0.00237285f $X=3.495 $Y=1.2 $X2=0
+ $Y2=0
cc_211 N_A_86_21#_c_169_n N_A_654_355#_c_489_n 0.00314391f $X=3.66 $Y=2.145
+ $X2=0 $Y2=0
cc_212 N_A_86_21#_c_170_n N_A_654_355#_c_490_n 0.00574613f $X=4.17 $Y=1.2 $X2=0
+ $Y2=0
cc_213 N_A_86_21#_c_174_n N_A_654_355#_c_490_n 0.00299589f $X=4.615 $Y=0.835
+ $X2=0 $Y2=0
cc_214 N_A_86_21#_c_169_n N_A_654_355#_c_491_n 0.00967686f $X=3.66 $Y=2.145
+ $X2=0 $Y2=0
cc_215 N_A_86_21#_c_170_n N_A_654_355#_c_491_n 0.00377086f $X=4.17 $Y=1.2 $X2=0
+ $Y2=0
cc_216 N_A_86_21#_c_170_n N_A_654_355#_c_492_n 0.00149568f $X=4.17 $Y=1.2 $X2=0
+ $Y2=0
cc_217 N_A_86_21#_c_174_n N_A_654_355#_c_492_n 0.00799789f $X=4.615 $Y=0.835
+ $X2=0 $Y2=0
cc_218 N_A_86_21#_c_174_n N_A_654_355#_c_493_n 0.0149324f $X=4.615 $Y=0.835
+ $X2=0 $Y2=0
cc_219 N_A_86_21#_c_170_n N_A_654_355#_c_494_n 0.00390272f $X=4.17 $Y=1.2 $X2=0
+ $Y2=0
cc_220 N_A_86_21#_c_174_n N_B_c_603_n 0.0107687f $X=4.615 $Y=0.835 $X2=-0.19
+ $Y2=-0.245
cc_221 N_A_86_21#_c_174_n N_B_c_604_n 3.67374e-19 $X=4.615 $Y=0.835 $X2=0 $Y2=0
cc_222 N_A_86_21#_c_174_n N_B_c_608_n 0.0013073f $X=4.615 $Y=0.835 $X2=0 $Y2=0
cc_223 N_A_86_21#_c_164_n N_A_M1013_g 0.0136182f $X=2.87 $Y=0.86 $X2=0 $Y2=0
cc_224 N_A_86_21#_c_166_n N_A_M1013_g 0.00873064f $X=3.035 $Y=0.945 $X2=0 $Y2=0
cc_225 N_A_86_21#_c_196_p N_A_M1013_g 0.0082691f $X=3.035 $Y=1.115 $X2=0 $Y2=0
cc_226 N_A_86_21#_c_168_n N_A_M1013_g 0.00202154f $X=3.2 $Y=1.2 $X2=0 $Y2=0
cc_227 N_A_86_21#_c_166_n N_A_c_665_n 0.00383072f $X=3.035 $Y=0.945 $X2=0 $Y2=0
cc_228 N_A_86_21#_c_174_n N_A_c_665_n 0.00878848f $X=4.615 $Y=0.835 $X2=0 $Y2=0
cc_229 N_A_86_21#_M1012_g X 0.017758f $X=0.505 $Y=0.445 $X2=0 $Y2=0
cc_230 N_A_86_21#_M1009_g X 0.00525175f $X=0.935 $Y=2.545 $X2=0 $Y2=0
cc_231 N_A_86_21#_M1012_g N_X_c_768_n 0.00660176f $X=0.505 $Y=0.445 $X2=0 $Y2=0
cc_232 N_A_86_21#_M1002_g N_X_c_768_n 8.94139e-19 $X=0.865 $Y=0.445 $X2=0 $Y2=0
cc_233 N_A_86_21#_M1009_g X 0.0142655f $X=0.935 $Y=2.545 $X2=0 $Y2=0
cc_234 N_A_86_21#_M1009_g N_VPWR_c_791_n 0.0181886f $X=0.935 $Y=2.545 $X2=0
+ $Y2=0
cc_235 N_A_86_21#_M1009_g N_VPWR_c_793_n 0.00769046f $X=0.935 $Y=2.545 $X2=0
+ $Y2=0
cc_236 N_A_86_21#_M1009_g N_VPWR_c_790_n 0.0143431f $X=0.935 $Y=2.545 $X2=0
+ $Y2=0
cc_237 N_A_86_21#_M1019_d N_A_505_400#_c_848_n 0.00385398f $X=3.52 $Y=2 $X2=0
+ $Y2=0
cc_238 N_A_86_21#_M1012_g N_VGND_c_884_n 0.00218427f $X=0.505 $Y=0.445 $X2=0
+ $Y2=0
cc_239 N_A_86_21#_M1002_g N_VGND_c_884_n 0.0108815f $X=0.865 $Y=0.445 $X2=0
+ $Y2=0
cc_240 N_A_86_21#_c_166_n N_VGND_c_885_n 0.0113788f $X=3.035 $Y=0.945 $X2=0
+ $Y2=0
cc_241 N_A_86_21#_c_170_n N_VGND_c_885_n 0.0103214f $X=4.17 $Y=1.2 $X2=0 $Y2=0
cc_242 N_A_86_21#_c_173_n N_VGND_c_885_n 0.01178f $X=3.66 $Y=1.2 $X2=0 $Y2=0
cc_243 N_A_86_21#_c_174_n N_VGND_c_885_n 0.00972526f $X=4.615 $Y=0.835 $X2=0
+ $Y2=0
cc_244 N_A_86_21#_c_174_n N_VGND_c_886_n 0.00764838f $X=4.615 $Y=0.835 $X2=0
+ $Y2=0
cc_245 N_A_86_21#_c_166_n N_VGND_c_889_n 0.00699628f $X=3.035 $Y=0.945 $X2=0
+ $Y2=0
cc_246 N_A_86_21#_M1012_g N_VGND_c_891_n 0.00547815f $X=0.505 $Y=0.445 $X2=0
+ $Y2=0
cc_247 N_A_86_21#_M1002_g N_VGND_c_891_n 0.00486043f $X=0.865 $Y=0.445 $X2=0
+ $Y2=0
cc_248 N_A_86_21#_c_174_n N_VGND_c_892_n 0.00679357f $X=4.615 $Y=0.835 $X2=0
+ $Y2=0
cc_249 N_A_86_21#_M1012_g N_VGND_c_894_n 0.00842675f $X=0.505 $Y=0.445 $X2=0
+ $Y2=0
cc_250 N_A_86_21#_M1002_g N_VGND_c_894_n 0.00427207f $X=0.865 $Y=0.445 $X2=0
+ $Y2=0
cc_251 N_A_86_21#_c_164_n N_VGND_c_894_n 0.0297869f $X=2.87 $Y=0.86 $X2=0 $Y2=0
cc_252 N_A_86_21#_c_166_n N_VGND_c_894_n 0.00885524f $X=3.035 $Y=0.945 $X2=0
+ $Y2=0
cc_253 N_A_86_21#_c_174_n N_VGND_c_894_n 0.00869867f $X=4.615 $Y=0.835 $X2=0
+ $Y2=0
cc_254 N_A_86_21#_c_164_n N_A_476_125#_M1013_s 0.0109183f $X=2.87 $Y=0.86
+ $X2=-0.19 $Y2=-0.245
cc_255 N_A_86_21#_c_162_n N_A_476_125#_c_972_n 0.00809759f $X=1.775 $Y=1.21
+ $X2=0 $Y2=0
cc_256 N_A_86_21#_c_164_n N_A_476_125#_c_972_n 0.0252954f $X=2.87 $Y=0.86 $X2=0
+ $Y2=0
cc_257 N_A_86_21#_c_168_n N_A_476_125#_c_972_n 0.0133612f $X=3.2 $Y=1.2 $X2=0
+ $Y2=0
cc_258 N_A_86_21#_M1019_d N_A_476_125#_c_982_n 0.00582286f $X=3.52 $Y=2 $X2=0
+ $Y2=0
cc_259 N_A_86_21#_c_169_n N_A_476_125#_c_982_n 0.02102f $X=3.66 $Y=2.145 $X2=0
+ $Y2=0
cc_260 N_A_86_21#_c_169_n N_A_476_125#_c_974_n 0.0435217f $X=3.66 $Y=2.145 $X2=0
+ $Y2=0
cc_261 N_A_86_21#_c_174_n N_A_476_125#_c_975_n 0.031509f $X=4.615 $Y=0.835 $X2=0
+ $Y2=0
cc_262 N_A_86_21#_c_169_n N_A_476_125#_c_976_n 0.0136596f $X=3.66 $Y=2.145 $X2=0
+ $Y2=0
cc_263 N_A_86_21#_c_170_n N_A_476_125#_c_976_n 0.0124251f $X=4.17 $Y=1.2 $X2=0
+ $Y2=0
cc_264 N_A_86_21#_c_174_n N_A_476_125#_c_976_n 4.31638e-19 $X=4.615 $Y=0.835
+ $X2=0 $Y2=0
cc_265 N_A_86_21#_c_174_n A_823_125# 0.00183662f $X=4.615 $Y=0.835 $X2=-0.19
+ $Y2=-0.245
cc_266 N_C_N_M1000_g N_A_318_409#_c_349_n 0.010974f $X=1.465 $Y=2.545 $X2=0
+ $Y2=0
cc_267 C_N N_A_318_409#_c_349_n 6.98448e-19 $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_268 N_C_N_c_298_n N_A_318_409#_c_349_n 0.00125544f $X=1.655 $Y=1.64 $X2=0
+ $Y2=0
cc_269 N_C_N_c_292_n N_A_318_409#_c_357_n 0.00542644f $X=1.58 $Y=0.805 $X2=0
+ $Y2=0
cc_270 N_C_N_c_293_n N_A_318_409#_c_357_n 0.00797978f $X=1.37 $Y=0.805 $X2=0
+ $Y2=0
cc_271 N_C_N_c_295_n N_A_318_409#_c_357_n 8.85328e-19 $X=1.655 $Y=1.475 $X2=0
+ $Y2=0
cc_272 N_C_N_c_296_n N_A_318_409#_c_357_n 0.00108502f $X=1.655 $Y=0.805 $X2=0
+ $Y2=0
cc_273 N_C_N_M1000_g N_A_318_409#_c_367_n 0.0195254f $X=1.465 $Y=2.545 $X2=0
+ $Y2=0
cc_274 C_N N_A_318_409#_c_367_n 0.0112228f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_275 N_C_N_c_291_n N_A_318_409#_c_359_n 0.0018904f $X=1.295 $Y=0.73 $X2=0
+ $Y2=0
cc_276 N_C_N_c_292_n N_A_318_409#_c_359_n 0.00202101f $X=1.58 $Y=0.805 $X2=0
+ $Y2=0
cc_277 N_C_N_c_294_n N_A_318_409#_c_359_n 0.00602462f $X=1.655 $Y=0.73 $X2=0
+ $Y2=0
cc_278 N_C_N_c_296_n N_A_318_409#_c_359_n 0.00173995f $X=1.655 $Y=0.805 $X2=0
+ $Y2=0
cc_279 N_C_N_M1000_g N_A_318_409#_c_368_n 0.0102692f $X=1.465 $Y=2.545 $X2=0
+ $Y2=0
cc_280 N_C_N_c_294_n N_A_318_409#_c_425_n 0.00250803f $X=1.655 $Y=0.73 $X2=0
+ $Y2=0
cc_281 N_C_N_c_294_n N_A_318_409#_c_360_n 0.00881787f $X=1.655 $Y=0.73 $X2=0
+ $Y2=0
cc_282 N_C_N_M1000_g N_A_318_409#_c_370_n 2.66868e-19 $X=1.465 $Y=2.545 $X2=0
+ $Y2=0
cc_283 N_C_N_M1000_g N_A_318_409#_c_371_n 0.00928588f $X=1.465 $Y=2.545 $X2=0
+ $Y2=0
cc_284 C_N N_A_318_409#_c_371_n 0.0187365f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_285 N_C_N_c_298_n N_A_318_409#_c_371_n 0.00379157f $X=1.655 $Y=1.64 $X2=0
+ $Y2=0
cc_286 N_C_N_M1000_g N_VPWR_c_791_n 0.0181144f $X=1.465 $Y=2.545 $X2=0 $Y2=0
cc_287 N_C_N_M1000_g N_VPWR_c_794_n 0.00769046f $X=1.465 $Y=2.545 $X2=0 $Y2=0
cc_288 N_C_N_M1000_g N_VPWR_c_790_n 0.0143431f $X=1.465 $Y=2.545 $X2=0 $Y2=0
cc_289 N_C_N_c_291_n N_VGND_c_884_n 0.00899674f $X=1.295 $Y=0.73 $X2=0 $Y2=0
cc_290 N_C_N_c_294_n N_VGND_c_884_n 0.00154134f $X=1.655 $Y=0.73 $X2=0 $Y2=0
cc_291 N_C_N_c_291_n N_VGND_c_889_n 0.00486043f $X=1.295 $Y=0.73 $X2=0 $Y2=0
cc_292 N_C_N_c_294_n N_VGND_c_889_n 0.00359944f $X=1.655 $Y=0.73 $X2=0 $Y2=0
cc_293 N_C_N_c_291_n N_VGND_c_894_n 0.00427207f $X=1.295 $Y=0.73 $X2=0 $Y2=0
cc_294 N_C_N_c_294_n N_VGND_c_894_n 0.00644174f $X=1.655 $Y=0.73 $X2=0 $Y2=0
cc_295 N_C_N_c_295_n N_A_476_125#_c_972_n 0.00302501f $X=1.655 $Y=1.475 $X2=0
+ $Y2=0
cc_296 C_N N_A_476_125#_c_979_n 0.00587354f $X=1.595 $Y=1.58 $X2=0 $Y2=0
cc_297 N_C_N_c_298_n N_A_476_125#_c_979_n 0.00311163f $X=1.655 $Y=1.64 $X2=0
+ $Y2=0
cc_298 N_A_318_409#_c_363_n N_A_654_355#_M1019_g 0.0463544f $X=2.935 $Y=1.925
+ $X2=0 $Y2=0
cc_299 N_A_318_409#_c_352_n N_A_654_355#_c_488_n 0.0128685f $X=3.535 $Y=1.46
+ $X2=0 $Y2=0
cc_300 N_A_318_409#_c_353_n N_A_654_355#_c_489_n 0.0128685f $X=3.325 $Y=1.46
+ $X2=0 $Y2=0
cc_301 N_A_318_409#_c_355_n N_A_654_355#_c_489_n 0.0463544f $X=2.935 $Y=1.85
+ $X2=0 $Y2=0
cc_302 N_A_318_409#_M1008_g N_A_654_355#_c_490_n 0.0152955f $X=3.61 $Y=0.835
+ $X2=0 $Y2=0
cc_303 N_A_318_409#_c_352_n N_A_654_355#_c_494_n 0.0152955f $X=3.535 $Y=1.46
+ $X2=0 $Y2=0
cc_304 N_A_318_409#_c_348_n N_A_M1013_g 0.00437433f $X=2.81 $Y=1.85 $X2=0 $Y2=0
cc_305 N_A_318_409#_M1016_g N_A_M1013_g 0.0136973f $X=3.25 $Y=0.835 $X2=0 $Y2=0
cc_306 N_A_318_409#_M1016_g N_A_c_665_n 0.00894493f $X=3.25 $Y=0.835 $X2=0 $Y2=0
cc_307 N_A_318_409#_M1008_g N_A_c_665_n 0.00894529f $X=3.61 $Y=0.835 $X2=0 $Y2=0
cc_308 N_A_318_409#_c_366_n N_X_M1009_s 0.0022818f $X=0.675 $Y=2.06 $X2=0 $Y2=0
cc_309 N_A_318_409#_c_369_n N_X_M1009_s 8.384e-19 $X=1.05 $Y=2.065 $X2=0 $Y2=0
cc_310 N_A_318_409#_c_356_n X 0.0740678f $X=0.59 $Y=1.975 $X2=0 $Y2=0
cc_311 N_A_318_409#_c_358_n X 0.0131605f $X=0.675 $Y=0.86 $X2=0 $Y2=0
cc_312 N_A_318_409#_c_366_n X 0.0139452f $X=0.675 $Y=2.06 $X2=0 $Y2=0
cc_313 N_A_318_409#_c_366_n X 0.0147089f $X=0.675 $Y=2.06 $X2=0 $Y2=0
cc_314 N_A_318_409#_c_369_n X 0.00775102f $X=1.05 $Y=2.065 $X2=0 $Y2=0
cc_315 N_A_318_409#_c_367_n N_VPWR_M1009_d 6.75075e-19 $X=1.565 $Y=2.07
+ $X2=-0.19 $Y2=-0.245
cc_316 N_A_318_409#_c_370_n N_VPWR_M1009_d 0.00112348f $X=1.22 $Y=2.065
+ $X2=-0.19 $Y2=-0.245
cc_317 N_A_318_409#_c_368_n N_VPWR_c_791_n 0.0381836f $X=1.73 $Y=2.9 $X2=0 $Y2=0
cc_318 N_A_318_409#_c_369_n N_VPWR_c_791_n 9.43903e-19 $X=1.05 $Y=2.065 $X2=0
+ $Y2=0
cc_319 N_A_318_409#_c_370_n N_VPWR_c_791_n 0.015332f $X=1.22 $Y=2.065 $X2=0
+ $Y2=0
cc_320 N_A_318_409#_c_371_n N_VPWR_c_791_n 0.0105054f $X=1.73 $Y=2.19 $X2=0
+ $Y2=0
cc_321 N_A_318_409#_c_363_n N_VPWR_c_794_n 0.00510529f $X=2.935 $Y=1.925 $X2=0
+ $Y2=0
cc_322 N_A_318_409#_c_368_n N_VPWR_c_794_n 0.0220321f $X=1.73 $Y=2.9 $X2=0 $Y2=0
cc_323 N_A_318_409#_c_363_n N_VPWR_c_790_n 0.00714516f $X=2.935 $Y=1.925 $X2=0
+ $Y2=0
cc_324 N_A_318_409#_c_368_n N_VPWR_c_790_n 0.0125808f $X=1.73 $Y=2.9 $X2=0 $Y2=0
cc_325 N_A_318_409#_c_371_n N_VPWR_c_790_n 0.0169786f $X=1.73 $Y=2.19 $X2=0
+ $Y2=0
cc_326 N_A_318_409#_c_363_n N_A_505_400#_c_848_n 0.0115234f $X=2.935 $Y=1.925
+ $X2=0 $Y2=0
cc_327 N_A_318_409#_c_363_n N_A_505_400#_c_849_n 0.00412617f $X=2.935 $Y=1.925
+ $X2=0 $Y2=0
cc_328 N_A_318_409#_c_368_n N_A_505_400#_c_849_n 0.00941491f $X=1.73 $Y=2.9
+ $X2=0 $Y2=0
cc_329 N_A_318_409#_c_357_n N_VGND_c_884_n 0.0198622f $X=1.425 $Y=0.86 $X2=0
+ $Y2=0
cc_330 N_A_318_409#_M1016_g N_VGND_c_885_n 0.00144941f $X=3.25 $Y=0.835 $X2=0
+ $Y2=0
cc_331 N_A_318_409#_M1008_g N_VGND_c_885_n 0.00925952f $X=3.61 $Y=0.835 $X2=0
+ $Y2=0
cc_332 N_A_318_409#_c_425_n N_VGND_c_889_n 0.00927824f $X=1.595 $Y=0.43 $X2=0
+ $Y2=0
cc_333 N_A_318_409#_c_360_n N_VGND_c_889_n 0.0254844f $X=1.87 $Y=0.43 $X2=0
+ $Y2=0
cc_334 N_A_318_409#_M1017_d N_VGND_c_894_n 0.00232217f $X=1.73 $Y=0.235 $X2=0
+ $Y2=0
cc_335 N_A_318_409#_M1016_g N_VGND_c_894_n 9.49986e-19 $X=3.25 $Y=0.835 $X2=0
+ $Y2=0
cc_336 N_A_318_409#_M1008_g N_VGND_c_894_n 7.97988e-19 $X=3.61 $Y=0.835 $X2=0
+ $Y2=0
cc_337 N_A_318_409#_c_357_n N_VGND_c_894_n 0.0145523f $X=1.425 $Y=0.86 $X2=0
+ $Y2=0
cc_338 N_A_318_409#_c_358_n N_VGND_c_894_n 0.00651511f $X=0.675 $Y=0.86 $X2=0
+ $Y2=0
cc_339 N_A_318_409#_c_425_n N_VGND_c_894_n 0.00649785f $X=1.595 $Y=0.43 $X2=0
+ $Y2=0
cc_340 N_A_318_409#_c_360_n N_VGND_c_894_n 0.0160028f $X=1.87 $Y=0.43 $X2=0
+ $Y2=0
cc_341 N_A_318_409#_c_425_n A_274_47# 9.59731e-19 $X=1.595 $Y=0.43 $X2=-0.19
+ $Y2=-0.245
cc_342 N_A_318_409#_M1016_g N_A_476_125#_c_972_n 0.00309831f $X=3.25 $Y=0.835
+ $X2=0 $Y2=0
cc_343 N_A_318_409#_c_353_n N_A_476_125#_c_972_n 0.00334419f $X=3.325 $Y=1.46
+ $X2=0 $Y2=0
cc_344 N_A_318_409#_c_348_n N_A_476_125#_c_973_n 0.016115f $X=2.81 $Y=1.85 $X2=0
+ $Y2=0
cc_345 N_A_318_409#_c_363_n N_A_476_125#_c_973_n 0.0122412f $X=2.935 $Y=1.925
+ $X2=0 $Y2=0
cc_346 N_A_318_409#_c_350_n N_A_476_125#_c_973_n 0.00565312f $X=2.985 $Y=1.775
+ $X2=0 $Y2=0
cc_347 N_A_318_409#_c_371_n N_A_476_125#_c_973_n 0.0437783f $X=1.73 $Y=2.19
+ $X2=0 $Y2=0
cc_348 N_A_318_409#_c_372_n N_A_476_125#_c_973_n 0.00175892f $X=2.2 $Y=1.98
+ $X2=0 $Y2=0
cc_349 N_A_318_409#_c_363_n N_A_476_125#_c_982_n 0.0235474f $X=2.935 $Y=1.925
+ $X2=0 $Y2=0
cc_350 N_A_318_409#_c_368_n N_A_476_125#_c_1010_n 0.00308874f $X=1.73 $Y=2.9
+ $X2=0 $Y2=0
cc_351 N_A_318_409#_c_371_n N_A_476_125#_c_1010_n 0.00626907f $X=1.73 $Y=2.19
+ $X2=0 $Y2=0
cc_352 N_A_318_409#_c_372_n N_A_476_125#_c_1010_n 3.3884e-19 $X=2.2 $Y=1.98
+ $X2=0 $Y2=0
cc_353 N_A_318_409#_c_349_n N_A_476_125#_c_979_n 0.00814725f $X=2.365 $Y=1.85
+ $X2=0 $Y2=0
cc_354 N_A_318_409#_c_353_n N_A_476_125#_c_979_n 0.00565312f $X=3.325 $Y=1.46
+ $X2=0 $Y2=0
cc_355 N_A_654_355#_c_493_n N_B_c_603_n 0.00972807f $X=4.4 $Y=1.12 $X2=-0.19
+ $Y2=-0.245
cc_356 N_A_654_355#_c_491_n N_B_c_604_n 0.00915914f $X=4.04 $Y=1.775 $X2=0 $Y2=0
cc_357 N_A_654_355#_c_488_n N_B_c_607_n 0.00617829f $X=3.965 $Y=1.85 $X2=0 $Y2=0
cc_358 N_A_654_355#_c_492_n N_B_c_607_n 0.00200612f $X=4.325 $Y=1.195 $X2=0
+ $Y2=0
cc_359 N_A_654_355#_c_503_n N_B_c_607_n 0.0059056f $X=6.395 $Y=2.49 $X2=0 $Y2=0
cc_360 N_A_654_355#_c_506_n N_B_c_607_n 0.0213356f $X=4.52 $Y=2.52 $X2=0 $Y2=0
cc_361 N_A_654_355#_c_507_n N_B_c_607_n 4.09747e-19 $X=4.685 $Y=2.52 $X2=0 $Y2=0
cc_362 N_A_654_355#_c_502_n N_B_M1011_g 0.00729837f $X=4.43 $Y=3.075 $X2=0 $Y2=0
cc_363 N_A_654_355#_c_503_n N_B_M1011_g 0.0182986f $X=6.395 $Y=2.49 $X2=0 $Y2=0
cc_364 N_A_654_355#_c_506_n N_B_M1011_g 0.00780546f $X=4.52 $Y=2.52 $X2=0 $Y2=0
cc_365 N_A_654_355#_c_507_n N_B_M1011_g 9.40379e-19 $X=4.685 $Y=2.52 $X2=0 $Y2=0
cc_366 N_A_654_355#_c_492_n N_B_c_609_n 0.00972807f $X=4.325 $Y=1.195 $X2=0
+ $Y2=0
cc_367 N_A_654_355#_c_506_n B 0.00195982f $X=4.52 $Y=2.52 $X2=0 $Y2=0
cc_368 N_A_654_355#_c_507_n B 0.0226851f $X=4.685 $Y=2.52 $X2=0 $Y2=0
cc_369 N_A_654_355#_c_490_n N_A_c_665_n 0.00894529f $X=4.04 $Y=1.12 $X2=0 $Y2=0
cc_370 N_A_654_355#_c_493_n N_A_c_665_n 0.00861922f $X=4.4 $Y=1.12 $X2=0 $Y2=0
cc_371 N_A_654_355#_c_503_n N_A_M1020_g 0.017497f $X=6.395 $Y=2.49 $X2=0 $Y2=0
cc_372 N_A_654_355#_c_508_n N_A_M1020_g 0.00166537f $X=6.56 $Y=2.16 $X2=0 $Y2=0
cc_373 N_A_654_355#_c_504_n N_D_N_c_730_n 0.00199732f $X=6.915 $Y=2.16 $X2=-0.19
+ $Y2=-0.245
cc_374 N_A_654_355#_c_495_n N_D_N_c_730_n 0.0075942f $X=7 $Y=2.075 $X2=-0.19
+ $Y2=-0.245
cc_375 N_A_654_355#_c_508_n N_D_N_c_730_n 0.00222881f $X=6.56 $Y=2.16 $X2=-0.19
+ $Y2=-0.245
cc_376 N_A_654_355#_c_503_n N_D_N_M1001_g 0.0204085f $X=6.395 $Y=2.49 $X2=0
+ $Y2=0
cc_377 N_A_654_355#_c_508_n N_D_N_M1001_g 0.010667f $X=6.56 $Y=2.16 $X2=0 $Y2=0
cc_378 N_A_654_355#_c_509_n N_D_N_M1001_g 0.0119428f $X=6.56 $Y=2.49 $X2=0 $Y2=0
cc_379 N_A_654_355#_c_496_n N_D_N_M1003_g 0.00111595f $X=6.92 $Y=0.47 $X2=0
+ $Y2=0
cc_380 N_A_654_355#_c_495_n N_D_N_M1006_g 0.0327249f $X=7 $Y=2.075 $X2=0 $Y2=0
cc_381 N_A_654_355#_c_496_n N_D_N_M1006_g 0.00850743f $X=6.92 $Y=0.47 $X2=0
+ $Y2=0
cc_382 N_A_654_355#_c_495_n D_N 0.0463087f $X=7 $Y=2.075 $X2=0 $Y2=0
cc_383 N_A_654_355#_c_508_n D_N 0.019204f $X=6.56 $Y=2.16 $X2=0 $Y2=0
cc_384 N_A_654_355#_c_503_n N_VPWR_M1020_d 0.0040089f $X=6.395 $Y=2.49 $X2=0
+ $Y2=0
cc_385 N_A_654_355#_c_503_n N_VPWR_c_792_n 0.0158375f $X=6.395 $Y=2.49 $X2=0
+ $Y2=0
cc_386 N_A_654_355#_c_509_n N_VPWR_c_792_n 0.0189303f $X=6.56 $Y=2.49 $X2=0
+ $Y2=0
cc_387 N_A_654_355#_c_501_n N_VPWR_c_794_n 0.0276595f $X=3.52 $Y=3.15 $X2=0
+ $Y2=0
cc_388 N_A_654_355#_c_503_n N_VPWR_c_794_n 0.00816968f $X=6.395 $Y=2.49 $X2=0
+ $Y2=0
cc_389 N_A_654_355#_c_503_n N_VPWR_c_795_n 0.0027514f $X=6.395 $Y=2.49 $X2=0
+ $Y2=0
cc_390 N_A_654_355#_c_509_n N_VPWR_c_795_n 0.019758f $X=6.56 $Y=2.49 $X2=0 $Y2=0
cc_391 N_A_654_355#_M1001_d N_VPWR_c_790_n 0.0023218f $X=6.42 $Y=2.095 $X2=0
+ $Y2=0
cc_392 N_A_654_355#_c_500_n N_VPWR_c_790_n 0.0250335f $X=4.355 $Y=3.15 $X2=0
+ $Y2=0
cc_393 N_A_654_355#_c_501_n N_VPWR_c_790_n 0.00801311f $X=3.52 $Y=3.15 $X2=0
+ $Y2=0
cc_394 N_A_654_355#_c_503_n N_VPWR_c_790_n 0.0228535f $X=6.395 $Y=2.49 $X2=0
+ $Y2=0
cc_395 N_A_654_355#_c_509_n N_VPWR_c_790_n 0.012508f $X=6.56 $Y=2.49 $X2=0 $Y2=0
cc_396 N_A_654_355#_c_503_n N_A_505_400#_M1011_s 0.0060424f $X=6.395 $Y=2.49
+ $X2=0 $Y2=0
cc_397 N_A_654_355#_M1019_g N_A_505_400#_c_848_n 0.0155089f $X=3.395 $Y=2.5
+ $X2=0 $Y2=0
cc_398 N_A_654_355#_c_500_n N_A_505_400#_c_848_n 0.0150315f $X=4.355 $Y=3.15
+ $X2=0 $Y2=0
cc_399 N_A_654_355#_c_502_n N_A_505_400#_c_848_n 0.0134022f $X=4.43 $Y=3.075
+ $X2=0 $Y2=0
cc_400 N_A_654_355#_c_503_n N_A_505_400#_c_848_n 0.0184421f $X=6.395 $Y=2.49
+ $X2=0 $Y2=0
cc_401 N_A_654_355#_c_506_n N_A_505_400#_c_848_n 0.00400978f $X=4.52 $Y=2.52
+ $X2=0 $Y2=0
cc_402 N_A_654_355#_c_507_n N_A_505_400#_c_848_n 0.0218436f $X=4.685 $Y=2.52
+ $X2=0 $Y2=0
cc_403 N_A_654_355#_M1019_g N_A_505_400#_c_849_n 5.12042e-19 $X=3.395 $Y=2.5
+ $X2=0 $Y2=0
cc_404 N_A_654_355#_c_503_n A_1076_419# 0.00386135f $X=6.395 $Y=2.49 $X2=-0.19
+ $Y2=-0.245
cc_405 N_A_654_355#_c_490_n N_VGND_c_885_n 0.00903154f $X=4.04 $Y=1.12 $X2=0
+ $Y2=0
cc_406 N_A_654_355#_c_493_n N_VGND_c_885_n 0.00137204f $X=4.4 $Y=1.12 $X2=0
+ $Y2=0
cc_407 N_A_654_355#_c_496_n N_VGND_c_888_n 0.0137175f $X=6.92 $Y=0.47 $X2=0
+ $Y2=0
cc_408 N_A_654_355#_c_496_n N_VGND_c_893_n 0.0195507f $X=6.92 $Y=0.47 $X2=0
+ $Y2=0
cc_409 N_A_654_355#_M1006_d N_VGND_c_894_n 0.00232985f $X=6.78 $Y=0.235 $X2=0
+ $Y2=0
cc_410 N_A_654_355#_c_490_n N_VGND_c_894_n 7.97988e-19 $X=4.04 $Y=1.12 $X2=0
+ $Y2=0
cc_411 N_A_654_355#_c_493_n N_VGND_c_894_n 9.49986e-19 $X=4.4 $Y=1.12 $X2=0
+ $Y2=0
cc_412 N_A_654_355#_c_496_n N_VGND_c_894_n 0.0124998f $X=6.92 $Y=0.47 $X2=0
+ $Y2=0
cc_413 N_A_654_355#_c_489_n N_A_476_125#_c_973_n 5.90928e-19 $X=3.52 $Y=1.85
+ $X2=0 $Y2=0
cc_414 N_A_654_355#_M1019_g N_A_476_125#_c_982_n 0.0238953f $X=3.395 $Y=2.5
+ $X2=0 $Y2=0
cc_415 N_A_654_355#_c_488_n N_A_476_125#_c_982_n 0.00567633f $X=3.965 $Y=1.85
+ $X2=0 $Y2=0
cc_416 N_A_654_355#_c_506_n N_A_476_125#_c_982_n 0.0013355f $X=4.52 $Y=2.52
+ $X2=0 $Y2=0
cc_417 N_A_654_355#_c_507_n N_A_476_125#_c_982_n 0.0144906f $X=4.685 $Y=2.52
+ $X2=0 $Y2=0
cc_418 N_A_654_355#_M1019_g N_A_476_125#_c_974_n 0.00318434f $X=3.395 $Y=2.5
+ $X2=0 $Y2=0
cc_419 N_A_654_355#_c_488_n N_A_476_125#_c_974_n 0.00708912f $X=3.965 $Y=1.85
+ $X2=0 $Y2=0
cc_420 N_A_654_355#_c_491_n N_A_476_125#_c_974_n 0.00379544f $X=4.04 $Y=1.775
+ $X2=0 $Y2=0
cc_421 N_A_654_355#_c_506_n N_A_476_125#_c_974_n 3.73707e-19 $X=4.52 $Y=2.52
+ $X2=0 $Y2=0
cc_422 N_A_654_355#_c_507_n N_A_476_125#_c_974_n 0.00389017f $X=4.685 $Y=2.52
+ $X2=0 $Y2=0
cc_423 N_A_654_355#_c_492_n N_A_476_125#_c_975_n 0.00300777f $X=4.325 $Y=1.195
+ $X2=0 $Y2=0
cc_424 N_A_654_355#_c_491_n N_A_476_125#_c_976_n 0.00781592f $X=4.04 $Y=1.775
+ $X2=0 $Y2=0
cc_425 N_A_654_355#_c_492_n N_A_476_125#_c_976_n 4.62928e-19 $X=4.325 $Y=1.195
+ $X2=0 $Y2=0
cc_426 N_A_654_355#_c_503_n N_A_476_125#_c_985_n 0.0604667f $X=6.395 $Y=2.49
+ $X2=0 $Y2=0
cc_427 N_A_654_355#_c_508_n N_A_476_125#_c_985_n 0.0114341f $X=6.56 $Y=2.16
+ $X2=0 $Y2=0
cc_428 N_A_654_355#_c_503_n N_A_476_125#_c_986_n 0.0132521f $X=6.395 $Y=2.49
+ $X2=0 $Y2=0
cc_429 N_B_c_603_n N_A_c_665_n 0.00894493f $X=4.83 $Y=1.12 $X2=0 $Y2=0
cc_430 N_B_c_608_n N_A_c_665_n 0.00907339f $X=5.19 $Y=1.12 $X2=0 $Y2=0
cc_431 N_B_c_606_n N_A_M1020_g 0.0792423f $X=5.13 $Y=1.89 $X2=0 $Y2=0
cc_432 N_B_c_608_n N_A_M1018_g 0.0139357f $X=5.19 $Y=1.12 $X2=0 $Y2=0
cc_433 N_B_c_604_n N_A_c_669_n 0.00184011f $X=4.83 $Y=1.815 $X2=0 $Y2=0
cc_434 N_B_c_606_n N_A_c_669_n 0.00392977f $X=5.13 $Y=1.89 $X2=0 $Y2=0
cc_435 N_B_c_604_n N_A_c_670_n 6.90103e-19 $X=4.83 $Y=1.815 $X2=0 $Y2=0
cc_436 N_B_c_606_n N_A_c_670_n 7.28704e-19 $X=5.13 $Y=1.89 $X2=0 $Y2=0
cc_437 N_B_M1011_g N_VPWR_c_792_n 0.0023756f $X=5.255 $Y=2.595 $X2=0 $Y2=0
cc_438 N_B_M1011_g N_VPWR_c_794_n 0.00723832f $X=5.255 $Y=2.595 $X2=0 $Y2=0
cc_439 N_B_M1011_g N_VPWR_c_790_n 0.00975423f $X=5.255 $Y=2.595 $X2=0 $Y2=0
cc_440 N_B_M1011_g N_A_505_400#_c_848_n 0.00426005f $X=5.255 $Y=2.595 $X2=0
+ $Y2=0
cc_441 N_B_c_606_n N_VGND_c_886_n 0.00212528f $X=5.13 $Y=1.89 $X2=0 $Y2=0
cc_442 N_B_c_608_n N_VGND_c_886_n 0.0126295f $X=5.19 $Y=1.12 $X2=0 $Y2=0
cc_443 N_B_c_603_n N_VGND_c_894_n 9.49986e-19 $X=4.83 $Y=1.12 $X2=0 $Y2=0
cc_444 N_B_c_608_n N_VGND_c_894_n 9.49986e-19 $X=5.19 $Y=1.12 $X2=0 $Y2=0
cc_445 N_B_c_604_n N_A_476_125#_c_974_n 0.00274974f $X=4.83 $Y=1.815 $X2=0 $Y2=0
cc_446 N_B_c_607_n N_A_476_125#_c_974_n 0.0057545f $X=4.905 $Y=1.89 $X2=0 $Y2=0
cc_447 B N_A_476_125#_c_974_n 0.0241369f $X=4.475 $Y=1.95 $X2=0 $Y2=0
cc_448 N_B_c_604_n N_A_476_125#_c_975_n 0.0189881f $X=4.83 $Y=1.815 $X2=0 $Y2=0
cc_449 N_B_c_605_n N_A_476_125#_c_975_n 0.00402814f $X=5.115 $Y=1.195 $X2=0
+ $Y2=0
cc_450 N_B_c_607_n N_A_476_125#_c_975_n 0.00432525f $X=4.905 $Y=1.89 $X2=0 $Y2=0
cc_451 B N_A_476_125#_c_975_n 0.0237494f $X=4.475 $Y=1.95 $X2=0 $Y2=0
cc_452 N_B_c_604_n N_A_476_125#_c_977_n 0.0085922f $X=4.83 $Y=1.815 $X2=0 $Y2=0
cc_453 N_B_c_606_n N_A_476_125#_c_977_n 0.00898979f $X=5.13 $Y=1.89 $X2=0 $Y2=0
cc_454 N_B_c_607_n N_A_476_125#_c_977_n 0.00415425f $X=4.905 $Y=1.89 $X2=0 $Y2=0
cc_455 N_B_M1011_g N_A_476_125#_c_977_n 0.00225096f $X=5.255 $Y=2.595 $X2=0
+ $Y2=0
cc_456 B N_A_476_125#_c_977_n 0.0166748f $X=4.475 $Y=1.95 $X2=0 $Y2=0
cc_457 N_B_c_606_n N_A_476_125#_c_985_n 0.00351081f $X=5.13 $Y=1.89 $X2=0 $Y2=0
cc_458 N_B_M1011_g N_A_476_125#_c_985_n 0.0217704f $X=5.255 $Y=2.595 $X2=0 $Y2=0
cc_459 N_B_c_607_n N_A_476_125#_c_986_n 8.1196e-19 $X=4.905 $Y=1.89 $X2=0 $Y2=0
cc_460 B N_A_476_125#_c_986_n 0.00759712f $X=4.475 $Y=1.95 $X2=0 $Y2=0
cc_461 N_A_M1020_g N_D_N_c_730_n 0.0425487f $X=5.745 $Y=2.595 $X2=-0.19
+ $Y2=-0.245
cc_462 N_A_M1018_g N_D_N_c_730_n 0.0129353f $X=5.78 $Y=1.135 $X2=-0.19
+ $Y2=-0.245
cc_463 N_A_c_669_n N_D_N_c_730_n 0.0116634f $X=5.755 $Y=1.71 $X2=-0.19
+ $Y2=-0.245
cc_464 N_A_c_665_n N_D_N_M1003_g 0.0129353f $X=5.705 $Y=0.18 $X2=0 $Y2=0
cc_465 N_A_M1020_g N_VPWR_c_792_n 0.0120934f $X=5.745 $Y=2.595 $X2=0 $Y2=0
cc_466 N_A_M1020_g N_VPWR_c_794_n 0.00661993f $X=5.745 $Y=2.595 $X2=0 $Y2=0
cc_467 N_A_M1020_g N_VPWR_c_790_n 0.00743555f $X=5.745 $Y=2.595 $X2=0 $Y2=0
cc_468 N_A_M1020_g N_A_505_400#_c_848_n 7.19588e-19 $X=5.745 $Y=2.595 $X2=0
+ $Y2=0
cc_469 N_A_c_665_n N_VGND_c_885_n 0.0253836f $X=5.705 $Y=0.18 $X2=0 $Y2=0
cc_470 N_A_c_665_n N_VGND_c_886_n 0.0229725f $X=5.705 $Y=0.18 $X2=0 $Y2=0
cc_471 N_A_M1018_g N_VGND_c_886_n 0.0189417f $X=5.78 $Y=1.135 $X2=0 $Y2=0
cc_472 N_A_c_669_n N_VGND_c_886_n 0.00148082f $X=5.755 $Y=1.71 $X2=0 $Y2=0
cc_473 N_A_c_670_n N_VGND_c_886_n 0.0204813f $X=5.755 $Y=1.71 $X2=0 $Y2=0
cc_474 N_A_c_665_n N_VGND_c_887_n 0.00796123f $X=5.705 $Y=0.18 $X2=0 $Y2=0
cc_475 N_A_c_665_n N_VGND_c_888_n 0.00572682f $X=5.705 $Y=0.18 $X2=0 $Y2=0
cc_476 N_A_c_666_n N_VGND_c_889_n 0.0295252f $X=2.895 $Y=0.18 $X2=0 $Y2=0
cc_477 N_A_c_665_n N_VGND_c_892_n 0.0432832f $X=5.705 $Y=0.18 $X2=0 $Y2=0
cc_478 N_A_c_665_n N_VGND_c_894_n 0.0925341f $X=5.705 $Y=0.18 $X2=0 $Y2=0
cc_479 N_A_c_666_n N_VGND_c_894_n 0.00692425f $X=2.895 $Y=0.18 $X2=0 $Y2=0
cc_480 N_A_M1013_g N_A_476_125#_c_972_n 0.0011274f $X=2.82 $Y=0.835 $X2=0 $Y2=0
cc_481 N_A_M1018_g N_A_476_125#_c_975_n 0.00195421f $X=5.78 $Y=1.135 $X2=0 $Y2=0
cc_482 N_A_c_669_n N_A_476_125#_c_975_n 3.34773e-19 $X=5.755 $Y=1.71 $X2=0 $Y2=0
cc_483 N_A_c_670_n N_A_476_125#_c_975_n 0.00470995f $X=5.755 $Y=1.71 $X2=0 $Y2=0
cc_484 N_A_M1020_g N_A_476_125#_c_977_n 3.18719e-19 $X=5.745 $Y=2.595 $X2=0
+ $Y2=0
cc_485 N_A_c_669_n N_A_476_125#_c_977_n 6.81758e-19 $X=5.755 $Y=1.71 $X2=0 $Y2=0
cc_486 N_A_c_670_n N_A_476_125#_c_977_n 0.0111371f $X=5.755 $Y=1.71 $X2=0 $Y2=0
cc_487 N_A_M1020_g N_A_476_125#_c_985_n 0.0149583f $X=5.745 $Y=2.595 $X2=0 $Y2=0
cc_488 N_A_c_669_n N_A_476_125#_c_985_n 0.00252644f $X=5.755 $Y=1.71 $X2=0 $Y2=0
cc_489 N_A_c_670_n N_A_476_125#_c_985_n 0.0329605f $X=5.755 $Y=1.71 $X2=0 $Y2=0
cc_490 N_A_M1020_g N_A_476_125#_c_978_n 0.00379441f $X=5.745 $Y=2.595 $X2=0
+ $Y2=0
cc_491 N_A_M1018_g N_A_476_125#_c_978_n 0.00384843f $X=5.78 $Y=1.135 $X2=0 $Y2=0
cc_492 N_A_c_669_n N_A_476_125#_c_978_n 0.00248633f $X=5.755 $Y=1.71 $X2=0 $Y2=0
cc_493 N_A_c_670_n N_A_476_125#_c_978_n 0.0243331f $X=5.755 $Y=1.71 $X2=0 $Y2=0
cc_494 N_A_M1018_g N_A_476_125#_c_980_n 0.00743077f $X=5.78 $Y=1.135 $X2=0 $Y2=0
cc_495 N_A_c_669_n N_A_476_125#_c_980_n 0.00257741f $X=5.755 $Y=1.71 $X2=0 $Y2=0
cc_496 N_A_c_670_n N_A_476_125#_c_980_n 0.00255596f $X=5.755 $Y=1.71 $X2=0 $Y2=0
cc_497 N_D_N_M1001_g N_VPWR_c_792_n 0.0105481f $X=6.295 $Y=2.595 $X2=0 $Y2=0
cc_498 N_D_N_M1001_g N_VPWR_c_795_n 0.00708727f $X=6.295 $Y=2.595 $X2=0 $Y2=0
cc_499 N_D_N_M1001_g N_VPWR_c_790_n 0.00922111f $X=6.295 $Y=2.595 $X2=0 $Y2=0
cc_500 N_D_N_M1003_g N_VGND_c_888_n 0.0139571f $X=6.345 $Y=0.445 $X2=0 $Y2=0
cc_501 N_D_N_M1006_g N_VGND_c_888_n 0.00239794f $X=6.705 $Y=0.445 $X2=0 $Y2=0
cc_502 N_D_N_M1003_g N_VGND_c_893_n 0.00486043f $X=6.345 $Y=0.445 $X2=0 $Y2=0
cc_503 N_D_N_M1006_g N_VGND_c_893_n 0.00549284f $X=6.705 $Y=0.445 $X2=0 $Y2=0
cc_504 N_D_N_M1003_g N_VGND_c_894_n 0.00814425f $X=6.345 $Y=0.445 $X2=0 $Y2=0
cc_505 N_D_N_M1006_g N_VGND_c_894_n 0.010905f $X=6.705 $Y=0.445 $X2=0 $Y2=0
cc_506 N_D_N_M1001_g N_A_476_125#_c_985_n 0.00657695f $X=6.295 $Y=2.595 $X2=0
+ $Y2=0
cc_507 N_D_N_c_730_n N_A_476_125#_c_978_n 0.0138658f $X=6.295 $Y=1.905 $X2=0
+ $Y2=0
cc_508 N_D_N_M1001_g N_A_476_125#_c_978_n 0.00745999f $X=6.295 $Y=2.595 $X2=0
+ $Y2=0
cc_509 N_D_N_M1003_g N_A_476_125#_c_980_n 0.00657717f $X=6.345 $Y=0.445 $X2=0
+ $Y2=0
cc_510 D_N N_A_476_125#_c_980_n 0.0494035f $X=6.395 $Y=1.21 $X2=0 $Y2=0
cc_511 X N_VPWR_c_791_n 0.0510876f $X=0.24 $Y=2.405 $X2=0 $Y2=0
cc_512 X N_VPWR_c_793_n 0.0476534f $X=0.24 $Y=2.405 $X2=0 $Y2=0
cc_513 X N_VPWR_c_790_n 0.0272842f $X=0.24 $Y=2.405 $X2=0 $Y2=0
cc_514 N_X_c_768_n N_VGND_c_884_n 0.0109996f $X=0.29 $Y=0.43 $X2=0 $Y2=0
cc_515 N_X_c_768_n N_VGND_c_891_n 0.0188684f $X=0.29 $Y=0.43 $X2=0 $Y2=0
cc_516 N_X_M1012_s N_VGND_c_894_n 0.00232217f $X=0.145 $Y=0.235 $X2=0 $Y2=0
cc_517 N_X_c_768_n N_VGND_c_894_n 0.0123379f $X=0.29 $Y=0.43 $X2=0 $Y2=0
cc_518 N_VPWR_c_790_n N_A_505_400#_M1011_s 0.0023412f $X=6.96 $Y=3.33 $X2=0
+ $Y2=0
cc_519 N_VPWR_c_794_n N_A_505_400#_c_848_n 0.116216f $X=5.845 $Y=3.33 $X2=0
+ $Y2=0
cc_520 N_VPWR_c_790_n N_A_505_400#_c_848_n 0.0786091f $X=6.96 $Y=3.33 $X2=0
+ $Y2=0
cc_521 N_VPWR_c_794_n N_A_505_400#_c_849_n 0.0174975f $X=5.845 $Y=3.33 $X2=0
+ $Y2=0
cc_522 N_VPWR_c_790_n N_A_505_400#_c_849_n 0.0120749f $X=6.96 $Y=3.33 $X2=0
+ $Y2=0
cc_523 N_VPWR_c_790_n A_1076_419# 0.00321616f $X=6.96 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_524 N_VPWR_c_790_n N_A_476_125#_c_982_n 0.00302344f $X=6.96 $Y=3.33 $X2=0
+ $Y2=0
cc_525 N_VPWR_M1020_d N_A_476_125#_c_985_n 0.00204972f $X=5.87 $Y=2.095 $X2=0
+ $Y2=0
cc_526 N_A_505_400#_c_848_n A_612_400# 0.00129482f $X=4.99 $Y=2.95 $X2=-0.19
+ $Y2=1.655
cc_527 N_A_505_400#_M1014_s N_A_476_125#_c_973_n 0.0100549f $X=2.525 $Y=2 $X2=0
+ $Y2=0
cc_528 N_A_505_400#_M1014_s N_A_476_125#_c_982_n 0.0016529f $X=2.525 $Y=2 $X2=0
+ $Y2=0
cc_529 N_A_505_400#_c_848_n N_A_476_125#_c_982_n 0.05192f $X=4.99 $Y=2.95 $X2=0
+ $Y2=0
cc_530 N_A_505_400#_c_849_n N_A_476_125#_c_982_n 0.00414392f $X=2.67 $Y=2.85
+ $X2=0 $Y2=0
cc_531 N_A_505_400#_M1014_s N_A_476_125#_c_1010_n 0.00540198f $X=2.525 $Y=2
+ $X2=0 $Y2=0
cc_532 N_A_505_400#_c_849_n N_A_476_125#_c_1010_n 0.0131037f $X=2.67 $Y=2.85
+ $X2=0 $Y2=0
cc_533 N_A_505_400#_M1011_s N_A_476_125#_c_985_n 4.03818e-19 $X=4.845 $Y=2.095
+ $X2=0 $Y2=0
cc_534 N_A_505_400#_M1011_s N_A_476_125#_c_986_n 0.00619517f $X=4.845 $Y=2.095
+ $X2=0 $Y2=0
cc_535 A_612_400# N_A_476_125#_c_982_n 0.00491832f $X=3.06 $Y=2 $X2=0 $Y2=0
cc_536 A_1076_419# N_A_476_125#_c_985_n 0.00137516f $X=5.38 $Y=2.095 $X2=4.115
+ $Y2=1.195
cc_537 A_116_47# N_VGND_c_894_n 0.00287567f $X=0.58 $Y=0.235 $X2=6.96 $Y2=0
cc_538 N_VGND_c_894_n A_274_47# 0.00200144f $X=6.96 $Y=0 $X2=-0.19 $Y2=-0.245
cc_539 N_VGND_c_886_n N_A_476_125#_c_980_n 0.018399f $X=5.485 $Y=0.77 $X2=0
+ $Y2=0
cc_540 N_VGND_c_888_n N_A_476_125#_c_980_n 0.0185998f $X=6.13 $Y=0.445 $X2=0
+ $Y2=0
cc_541 N_VGND_c_894_n A_1284_47# 0.00899413f $X=6.96 $Y=0 $X2=-0.19 $Y2=-0.245
