* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__or4bb_2 A B C_N D_N VGND VNB VPB VPWR X
X0 VGND a_40_47# a_276_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 X a_276_47# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X2 a_40_47# C_N VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 a_276_47# a_462_351# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 VGND D_N a_462_351# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 VPWR D_N a_462_351# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X6 a_348_403# a_40_47# a_420_403# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X7 a_420_403# a_462_351# a_276_47# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X8 VPWR a_276_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X9 a_40_47# C_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X10 VPWR A a_276_403# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X11 a_276_403# B a_348_403# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X12 VGND a_276_47# X VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X13 VGND A a_276_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X14 a_276_47# B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X15 X a_276_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
.ends
