* File: sky130_fd_sc_lp__dfbbn_2.pex.spice
* Created: Fri Aug 28 10:21:17 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__DFBBN_2%CLK_N 2 5 7 9 12 14 17 19 20 21 26 27
r34 26 27 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.27
+ $Y=1.075 $X2=0.27 $Y2=1.075
r35 20 21 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.27 $Y=1.665
+ $X2=0.27 $Y2=2.035
r36 19 20 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.27 $Y=1.295
+ $X2=0.27 $Y2=1.665
r37 19 27 7.68295 $w=3.28e-07 $l=2.2e-07 $layer=LI1_cond $X=0.27 $Y=1.295
+ $X2=0.27 $Y2=1.075
r38 15 17 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=0.36 $Y=2.255
+ $X2=0.6 $Y2=2.255
r39 13 26 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.27 $Y=1.415
+ $X2=0.27 $Y2=1.075
r40 13 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.27 $Y=1.415
+ $X2=0.27 $Y2=1.58
r41 12 26 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=0.27 $Y=1.06
+ $X2=0.27 $Y2=1.075
r42 11 12 43.5886 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=0.335 $Y=0.91
+ $X2=0.335 $Y2=1.06
r43 7 17 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.6 $Y=2.33 $X2=0.6
+ $Y2=2.255
r44 7 9 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.6 $Y=2.33 $X2=0.6
+ $Y2=2.725
r45 5 11 212.798 $w=1.5e-07 $l=4.15e-07 $layer=POLY_cond $X=0.49 $Y=0.495
+ $X2=0.49 $Y2=0.91
r46 2 15 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.36 $Y=2.18 $X2=0.36
+ $Y2=2.255
r47 2 14 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=0.36 $Y=2.18 $X2=0.36
+ $Y2=1.58
.ends

.subckt PM_SKY130_FD_SC_LP__DFBBN_2%D 2 3 5 7 8 10 13 15 17 21
c55 21 0 1.13211e-19 $X=1.92 $Y=1.345
c56 17 0 3.67314e-20 $X=1.92 $Y=1.165
r57 20 22 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.92 $Y=1.345
+ $X2=1.92 $Y2=1.51
r58 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.92
+ $Y=1.345 $X2=1.92 $Y2=1.345
r59 17 20 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=1.92 $Y=1.165
+ $X2=1.92 $Y2=1.345
r60 15 21 8.3814 $w=3.28e-07 $l=2.4e-07 $layer=LI1_cond $X=1.68 $Y=1.345
+ $X2=1.92 $Y2=1.345
r61 11 13 133.319 $w=1.5e-07 $l=2.6e-07 $layer=POLY_cond $X=1.98 $Y=2.095
+ $X2=2.24 $Y2=2.095
r62 8 10 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.395 $Y=1.09
+ $X2=2.395 $Y2=0.805
r63 5 13 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.24 $Y=2.17 $X2=2.24
+ $Y2=2.095
r64 5 7 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.24 $Y=2.17 $X2=2.24
+ $Y2=2.455
r65 4 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.085 $Y=1.165
+ $X2=1.92 $Y2=1.165
r66 3 8 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.32 $Y=1.165
+ $X2=2.395 $Y2=1.09
r67 3 4 120.5 $w=1.5e-07 $l=2.35e-07 $layer=POLY_cond $X=2.32 $Y=1.165 $X2=2.085
+ $Y2=1.165
r68 2 11 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.98 $Y=2.02 $X2=1.98
+ $Y2=2.095
r69 2 22 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=1.98 $Y=2.02 $X2=1.98
+ $Y2=1.51
.ends

.subckt PM_SKY130_FD_SC_LP__DFBBN_2%A_113_57# 1 2 7 8 9 10 14 18 19 20 21 22 25
+ 30 33 34 36 44 50 54 55 57 58 60 61 62 64 65 66 68 69 70 73 74 77 81 82 83 84
+ 88 96
c248 96 0 1.71827e-19 $X=7.61 $Y=1.345
c249 88 0 2.25888e-20 $X=7.61 $Y=1.51
c250 73 0 1.23337e-19 $X=8.51 $Y=1.865
c251 54 0 9.08694e-20 $X=3.54 $Y=1.255
c252 7 0 2.98096e-20 $X=1.395 $Y=1.375
r253 88 96 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.61 $Y=1.51
+ $X2=7.61 $Y2=1.345
r254 87 89 8.83531 $w=4.38e-07 $l=1.65e-07 $layer=LI1_cond $X=7.555 $Y=1.51
+ $X2=7.555 $Y2=1.675
r255 87 88 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.61
+ $Y=1.51 $X2=7.61 $Y2=1.51
r256 84 87 8.90524 $w=4.38e-07 $l=3.4e-07 $layer=LI1_cond $X=7.555 $Y=1.17
+ $X2=7.555 $Y2=1.51
r257 81 83 7.01288 $w=3.53e-07 $l=1.65e-07 $layer=LI1_cond $X=0.827 $Y=1.465
+ $X2=0.827 $Y2=1.3
r258 81 82 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.84
+ $Y=1.465 $X2=0.84 $Y2=1.465
r259 79 83 30.1207 $w=2.18e-07 $l=5.75e-07 $layer=LI1_cond $X=0.76 $Y=0.725
+ $X2=0.76 $Y2=1.3
r260 77 79 9.31567 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=0.705 $Y=0.495
+ $X2=0.705 $Y2=0.725
r261 73 74 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=8.51
+ $Y=1.865 $X2=8.51 $Y2=1.865
r262 71 73 43.9636 $w=2.68e-07 $l=1.03e-06 $layer=LI1_cond $X=8.48 $Y=2.895
+ $X2=8.48 $Y2=1.865
r263 69 71 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=8.345 $Y=2.98
+ $X2=8.48 $Y2=2.895
r264 69 70 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=8.345 $Y=2.98
+ $X2=7.505 $Y2=2.98
r265 68 70 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.42 $Y=2.895
+ $X2=7.505 $Y2=2.98
r266 68 89 79.5936 $w=1.68e-07 $l=1.22e-06 $layer=LI1_cond $X=7.42 $Y=2.895
+ $X2=7.42 $Y2=1.675
r267 65 84 6.36164 $w=1.7e-07 $l=2.2e-07 $layer=LI1_cond $X=7.335 $Y=1.17
+ $X2=7.555 $Y2=1.17
r268 65 66 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=7.335 $Y=1.17
+ $X2=6.68 $Y2=1.17
r269 64 66 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.595 $Y=1.085
+ $X2=6.68 $Y2=1.17
r270 63 64 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=6.595 $Y=0.435
+ $X2=6.595 $Y2=1.085
r271 61 63 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.51 $Y=0.35
+ $X2=6.595 $Y2=0.435
r272 61 62 106.016 $w=1.68e-07 $l=1.625e-06 $layer=LI1_cond $X=6.51 $Y=0.35
+ $X2=4.885 $Y2=0.35
r273 59 62 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.8 $Y=0.435
+ $X2=4.885 $Y2=0.35
r274 59 60 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=4.8 $Y=0.435
+ $X2=4.8 $Y2=1.055
r275 57 60 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.715 $Y=1.14
+ $X2=4.8 $Y2=1.055
r276 57 58 70.1337 $w=1.68e-07 $l=1.075e-06 $layer=LI1_cond $X=4.715 $Y=1.14
+ $X2=3.64 $Y2=1.14
r277 54 55 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.54
+ $Y=1.255 $X2=3.54 $Y2=1.255
r278 52 58 6.87494 $w=1.7e-07 $l=1.36015e-07 $layer=LI1_cond $X=3.54 $Y=1.225
+ $X2=3.64 $Y2=1.14
r279 52 54 1.66364 $w=1.98e-07 $l=3e-08 $layer=LI1_cond $X=3.54 $Y=1.225
+ $X2=3.54 $Y2=1.255
r280 48 81 0.389558 $w=3.53e-07 $l=1.2e-08 $layer=LI1_cond $X=0.827 $Y=1.477
+ $X2=0.827 $Y2=1.465
r281 48 50 34.833 $w=3.53e-07 $l=1.073e-06 $layer=LI1_cond $X=0.827 $Y=1.477
+ $X2=0.827 $Y2=2.55
r282 44 74 76.939 $w=3.3e-07 $l=4.4e-07 $layer=POLY_cond $X=8.51 $Y=2.305
+ $X2=8.51 $Y2=1.865
r283 41 44 187.16 $w=1.5e-07 $l=3.65e-07 $layer=POLY_cond $X=8.145 $Y=2.38
+ $X2=8.51 $Y2=2.38
r284 40 55 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.54 $Y=1.09
+ $X2=3.54 $Y2=1.255
r285 38 82 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=0.84 $Y=1.82
+ $X2=0.84 $Y2=1.465
r286 37 82 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=0.84 $Y=1.45
+ $X2=0.84 $Y2=1.465
r287 34 41 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.145 $Y=2.455
+ $X2=8.145 $Y2=2.38
r288 34 36 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=8.145 $Y=2.455
+ $X2=8.145 $Y2=2.74
r289 33 96 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=7.67 $Y=0.915
+ $X2=7.67 $Y2=1.345
r290 30 40 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=3.45 $Y=0.73
+ $X2=3.45 $Y2=1.09
r291 27 30 243.564 $w=1.5e-07 $l=4.75e-07 $layer=POLY_cond $X=3.45 $Y=0.255
+ $X2=3.45 $Y2=0.73
r292 23 25 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=2.67 $Y=3.005
+ $X2=2.67 $Y2=2.455
r293 21 23 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.595 $Y=3.08
+ $X2=2.67 $Y2=3.005
r294 21 22 476.872 $w=1.5e-07 $l=9.3e-07 $layer=POLY_cond $X=2.595 $Y=3.08
+ $X2=1.665 $Y2=3.08
r295 19 27 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.375 $Y=0.18
+ $X2=3.45 $Y2=0.255
r296 19 20 938.362 $w=1.5e-07 $l=1.83e-06 $layer=POLY_cond $X=3.375 $Y=0.18
+ $X2=1.545 $Y2=0.18
r297 16 22 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.59 $Y=3.005
+ $X2=1.665 $Y2=3.08
r298 16 18 225.617 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=1.59 $Y=3.005
+ $X2=1.59 $Y2=2.565
r299 15 18 305.096 $w=1.5e-07 $l=5.95e-07 $layer=POLY_cond $X=1.59 $Y=1.97
+ $X2=1.59 $Y2=2.565
r300 12 14 253.819 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=1.47 $Y=1.3
+ $X2=1.47 $Y2=0.805
r301 11 20 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.47 $Y=0.255
+ $X2=1.545 $Y2=0.18
r302 11 14 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=1.47 $Y=0.255
+ $X2=1.47 $Y2=0.805
r303 10 38 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=1.005 $Y=1.895
+ $X2=0.84 $Y2=1.82
r304 9 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.515 $Y=1.895
+ $X2=1.59 $Y2=1.97
r305 9 10 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=1.515 $Y=1.895
+ $X2=1.005 $Y2=1.895
r306 8 37 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=1.005 $Y=1.375
+ $X2=0.84 $Y2=1.45
r307 7 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.395 $Y=1.375
+ $X2=1.47 $Y2=1.3
r308 7 8 199.979 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=1.395 $Y=1.375
+ $X2=1.005 $Y2=1.375
r309 2 50 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=0.675
+ $Y=2.405 $X2=0.815 $Y2=2.55
r310 1 77 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.565
+ $Y=0.285 $X2=0.705 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__DFBBN_2%A_789_78# 1 2 9 13 17 21 25 26 29 30 33 35
+ 40 41 43 45 47 48 49
c131 41 0 1.52357e-19 $X=5.47 $Y=2.532
c132 35 0 1.76227e-19 $X=5.97 $Y=2.31
r133 48 57 45.9078 $w=4.1e-07 $l=1.65e-07 $layer=POLY_cond $X=7.03 $Y=1.57
+ $X2=7.03 $Y2=1.735
r134 48 56 45.9078 $w=4.1e-07 $l=1.65e-07 $layer=POLY_cond $X=7.03 $Y=1.57
+ $X2=7.03 $Y2=1.405
r135 47 49 8.48463 $w=2.98e-07 $l=1.65e-07 $layer=LI1_cond $X=6.99 $Y=1.585
+ $X2=6.825 $Y2=1.585
r136 47 48 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.99
+ $Y=1.57 $X2=6.99 $Y2=1.57
r137 43 44 10.0214 $w=2.8e-07 $l=2.3e-07 $layer=LI1_cond $X=5.74 $Y=1.13
+ $X2=5.97 $Y2=1.13
r138 39 41 8.86124 $w=4.43e-07 $l=1.65e-07 $layer=LI1_cond $X=5.305 $Y=2.532
+ $X2=5.47 $Y2=2.532
r139 39 40 8.86124 $w=4.43e-07 $l=1.65e-07 $layer=LI1_cond $X=5.305 $Y=2.532
+ $X2=5.14 $Y2=2.532
r140 37 45 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.055 $Y=1.52
+ $X2=5.97 $Y2=1.52
r141 37 49 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=6.055 $Y=1.52
+ $X2=6.825 $Y2=1.52
r142 34 45 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.97 $Y=1.605
+ $X2=5.97 $Y2=1.52
r143 34 35 45.9947 $w=1.68e-07 $l=7.05e-07 $layer=LI1_cond $X=5.97 $Y=1.605
+ $X2=5.97 $Y2=2.31
r144 33 45 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.97 $Y=1.435
+ $X2=5.97 $Y2=1.52
r145 32 44 3.65648 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.97 $Y=1.295
+ $X2=5.97 $Y2=1.13
r146 32 33 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=5.97 $Y=1.295
+ $X2=5.97 $Y2=1.435
r147 30 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.885 $Y=2.395
+ $X2=5.97 $Y2=2.31
r148 30 41 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=5.885 $Y=2.395
+ $X2=5.47 $Y2=2.395
r149 29 40 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=4.37 $Y=2.395
+ $X2=5.14 $Y2=2.395
r150 26 51 43.7153 $w=3.3e-07 $l=2.5e-07 $layer=POLY_cond $X=4.27 $Y=1.92
+ $X2=4.02 $Y2=1.92
r151 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.27
+ $Y=1.92 $X2=4.27 $Y2=1.92
r152 23 29 6.87494 $w=1.7e-07 $l=1.36015e-07 $layer=LI1_cond $X=4.27 $Y=2.31
+ $X2=4.37 $Y2=2.395
r153 23 25 21.6273 $w=1.98e-07 $l=3.9e-07 $layer=LI1_cond $X=4.27 $Y=2.31
+ $X2=4.27 $Y2=1.92
r154 21 57 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=7.16 $Y=2.315
+ $X2=7.16 $Y2=1.735
r155 17 56 251.255 $w=1.5e-07 $l=4.9e-07 $layer=POLY_cond $X=7.16 $Y=0.915
+ $X2=7.16 $Y2=1.405
r156 11 51 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.02 $Y=2.085
+ $X2=4.02 $Y2=1.92
r157 11 13 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=4.02 $Y=2.085
+ $X2=4.02 $Y2=2.455
r158 7 51 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.02 $Y=1.755
+ $X2=4.02 $Y2=1.92
r159 7 9 525.585 $w=1.5e-07 $l=1.025e-06 $layer=POLY_cond $X=4.02 $Y=1.755
+ $X2=4.02 $Y2=0.73
r160 2 39 600 $w=1.7e-07 $l=7.01516e-07 $layer=licon1_PDIFF $count=1 $X=5.165
+ $Y=1.895 $X2=5.305 $Y2=2.53
r161 1 43 182 $w=1.7e-07 $l=9.31316e-07 $layer=licon1_NDIFF $count=1 $X=5.525
+ $Y=0.3 $X2=5.74 $Y2=1.13
.ends

.subckt PM_SKY130_FD_SC_LP__DFBBN_2%SET_B 3 7 11 13 15 16 18 19 25 29 30
c127 30 0 7.79776e-20 $X=5 $Y=1.57
c128 18 0 1.31498e-19 $X=8.735 $Y=1.665
r129 29 32 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5 $Y=1.57 $X2=5
+ $Y2=1.735
r130 29 31 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5 $Y=1.57 $X2=5
+ $Y2=1.405
r131 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5 $Y=1.57
+ $X2=5 $Y2=1.57
r132 25 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=1.665
+ $X2=8.88 $Y2=1.665
r133 21 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=1.665
+ $X2=5.04 $Y2=1.665
r134 19 21 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.185 $Y=1.665
+ $X2=5.04 $Y2=1.665
r135 18 25 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.735 $Y=1.665
+ $X2=8.88 $Y2=1.665
r136 18 19 4.39356 $w=1.4e-07 $l=3.55e-06 $layer=MET1_cond $X=8.735 $Y=1.665
+ $X2=5.185 $Y2=1.665
r137 16 26 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=9.36 $Y=1.635
+ $X2=8.88 $Y2=1.635
r138 16 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.41
+ $Y=1.635 $X2=9.41 $Y2=1.635
r139 13 34 79.8686 $w=3.09e-07 $l=5.23775e-07 $layer=POLY_cond $X=9.735 $Y=2.065
+ $X2=9.527 $Y2=1.635
r140 13 15 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=9.735 $Y=2.065
+ $X2=9.735 $Y2=2.56
r141 9 34 38.532 $w=3.09e-07 $l=1.87029e-07 $layer=POLY_cond $X=9.48 $Y=1.47
+ $X2=9.527 $Y2=1.635
r142 9 11 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=9.48 $Y=1.47
+ $X2=9.48 $Y2=0.915
r143 7 32 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=5.09 $Y=2.315
+ $X2=5.09 $Y2=1.735
r144 3 31 402.521 $w=1.5e-07 $l=7.85e-07 $layer=POLY_cond $X=5.015 $Y=0.62
+ $X2=5.015 $Y2=1.405
.ends

.subckt PM_SKY130_FD_SC_LP__DFBBN_2%A_549_449# 1 2 9 13 17 20 21 24 25 26 28 29
+ 30 33 34 36 41
c139 34 0 1.52357e-19 $X=5.54 $Y=1.57
c140 13 0 7.79776e-20 $X=5.52 $Y=2.315
r141 40 41 9.2801 $w=4.58e-07 $l=1.65e-07 $layer=LI1_cond $X=3.255 $Y=2.455
+ $X2=3.42 $Y2=2.455
r142 37 40 2.08014 $w=4.58e-07 $l=8e-08 $layer=LI1_cond $X=3.175 $Y=2.455
+ $X2=3.255 $Y2=2.455
r143 34 44 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.54 $Y=1.57
+ $X2=5.54 $Y2=1.735
r144 34 43 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.54 $Y=1.57
+ $X2=5.54 $Y2=1.405
r145 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.54
+ $Y=1.57 $X2=5.54 $Y2=1.57
r146 31 33 13.6198 $w=3.28e-07 $l=3.9e-07 $layer=LI1_cond $X=5.54 $Y=1.96
+ $X2=5.54 $Y2=1.57
r147 29 31 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.375 $Y=2.045
+ $X2=5.54 $Y2=1.96
r148 29 30 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=5.375 $Y=2.045
+ $X2=4.72 $Y2=2.045
r149 28 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.635 $Y=1.96
+ $X2=4.72 $Y2=2.045
r150 27 28 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=4.635 $Y=1.575
+ $X2=4.635 $Y2=1.96
r151 25 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.55 $Y=1.49
+ $X2=4.635 $Y2=1.575
r152 25 26 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=4.55 $Y=1.49
+ $X2=3.99 $Y2=1.49
r153 23 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.905 $Y=1.575
+ $X2=3.99 $Y2=1.49
r154 23 24 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=3.905 $Y=1.575
+ $X2=3.905 $Y2=2.225
r155 21 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.82 $Y=2.31
+ $X2=3.905 $Y2=2.225
r156 21 41 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=3.82 $Y=2.31 $X2=3.42
+ $Y2=2.31
r157 20 37 6.6364 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=3.175 $Y=2.225
+ $X2=3.175 $Y2=2.455
r158 20 36 83.1818 $w=1.68e-07 $l=1.275e-06 $layer=LI1_cond $X=3.175 $Y=2.225
+ $X2=3.175 $Y2=0.95
r159 15 36 6.45221 $w=2.23e-07 $l=1.12e-07 $layer=LI1_cond $X=3.147 $Y=0.838
+ $X2=3.147 $Y2=0.95
r160 15 17 5.78782 $w=2.23e-07 $l=1.13e-07 $layer=LI1_cond $X=3.147 $Y=0.838
+ $X2=3.147 $Y2=0.725
r161 13 44 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=5.52 $Y=2.315
+ $X2=5.52 $Y2=1.735
r162 9 43 402.521 $w=1.5e-07 $l=7.85e-07 $layer=POLY_cond $X=5.45 $Y=0.62
+ $X2=5.45 $Y2=1.405
r163 2 40 600 $w=1.7e-07 $l=6.0597e-07 $layer=licon1_PDIFF $count=1 $X=2.745
+ $Y=2.245 $X2=3.255 $Y2=2.455
r164 1 17 182 $w=1.7e-07 $l=2.77489e-07 $layer=licon1_NDIFF $count=1 $X=2.9
+ $Y=0.595 $X2=3.12 $Y2=0.725
.ends

.subckt PM_SKY130_FD_SC_LP__DFBBN_2%A_223_119# 1 2 9 12 13 14 18 19 20 24 25 26
+ 28 29 30 31 33 34 35 38 41 43 47 51 54
c169 47 0 3.67314e-20 $X=2.46 $Y=1.645
c170 43 0 2.98096e-20 $X=2.295 $Y=1.96
c171 35 0 9.08694e-20 $X=2.825 $Y=1.66
c172 34 0 1.13211e-19 $X=2.75 $Y=1.645
c173 24 0 1.23337e-19 $X=7.635 $Y=2.56
r174 51 53 10.2083 $w=3.28e-07 $l=2.15e-07 $layer=LI1_cond $X=1.255 $Y=0.785
+ $X2=1.255 $Y2=1
r175 47 48 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.46
+ $Y=1.645 $X2=2.46 $Y2=1.645
r176 45 47 10.0023 $w=2.63e-07 $l=2.3e-07 $layer=LI1_cond $X=2.427 $Y=1.875
+ $X2=2.427 $Y2=1.645
r177 44 54 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.54 $Y=1.96
+ $X2=1.375 $Y2=1.96
r178 43 45 7.24806 $w=1.7e-07 $l=1.69245e-07 $layer=LI1_cond $X=2.295 $Y=1.96
+ $X2=2.427 $Y2=1.875
r179 43 44 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=2.295 $Y=1.96
+ $X2=1.54 $Y2=1.96
r180 39 54 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.375 $Y=2.045
+ $X2=1.375 $Y2=1.96
r181 39 41 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=1.375 $Y=2.045
+ $X2=1.375 $Y2=2.39
r182 38 54 3.70735 $w=2.5e-07 $l=1.18427e-07 $layer=LI1_cond $X=1.295 $Y=1.875
+ $X2=1.375 $Y2=1.96
r183 38 53 57.0856 $w=1.68e-07 $l=8.75e-07 $layer=LI1_cond $X=1.295 $Y=1.875
+ $X2=1.295 $Y2=1
r184 35 36 51.4864 $w=2.2e-07 $l=2.35e-07 $layer=POLY_cond $X=2.825 $Y=1.66
+ $X2=3.06 $Y2=1.66
r185 34 48 50.7098 $w=3.3e-07 $l=2.9e-07 $layer=POLY_cond $X=2.75 $Y=1.645
+ $X2=2.46 $Y2=1.645
r186 34 35 16.3226 $w=3.3e-07 $l=8.21584e-08 $layer=POLY_cond $X=2.75 $Y=1.645
+ $X2=2.825 $Y2=1.66
r187 31 33 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=8.415 $Y=1.31
+ $X2=8.415 $Y2=1.025
r188 29 31 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.34 $Y=1.385
+ $X2=8.415 $Y2=1.31
r189 29 30 105.117 $w=1.5e-07 $l=2.05e-07 $layer=POLY_cond $X=8.34 $Y=1.385
+ $X2=8.135 $Y2=1.385
r190 27 30 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.06 $Y=1.46
+ $X2=8.135 $Y2=1.385
r191 27 28 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=8.06 $Y=1.46
+ $X2=8.06 $Y2=1.915
r192 25 28 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.985 $Y=1.99
+ $X2=8.06 $Y2=1.915
r193 25 26 141.011 $w=1.5e-07 $l=2.75e-07 $layer=POLY_cond $X=7.985 $Y=1.99
+ $X2=7.71 $Y2=1.99
r194 22 24 264.074 $w=1.5e-07 $l=5.15e-07 $layer=POLY_cond $X=7.635 $Y=3.075
+ $X2=7.635 $Y2=2.56
r195 21 26 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.635 $Y=2.065
+ $X2=7.71 $Y2=1.99
r196 21 24 253.819 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=7.635 $Y=2.065
+ $X2=7.635 $Y2=2.56
r197 19 22 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.56 $Y=3.15
+ $X2=7.635 $Y2=3.075
r198 19 20 2058.76 $w=1.5e-07 $l=4.015e-06 $layer=POLY_cond $X=7.56 $Y=3.15
+ $X2=3.545 $Y2=3.15
r199 16 20 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.47 $Y=3.075
+ $X2=3.545 $Y2=3.15
r200 16 18 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=3.47 $Y=3.075
+ $X2=3.47 $Y2=2.455
r201 15 18 156.394 $w=1.5e-07 $l=3.05e-07 $layer=POLY_cond $X=3.47 $Y=2.15
+ $X2=3.47 $Y2=2.455
r202 13 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.395 $Y=2.075
+ $X2=3.47 $Y2=2.15
r203 13 14 133.319 $w=1.5e-07 $l=2.6e-07 $layer=POLY_cond $X=3.395 $Y=2.075
+ $X2=3.135 $Y2=2.075
r204 12 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.06 $Y=2
+ $X2=3.135 $Y2=2.075
r205 11 36 11.7719 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=3.06 $Y=1.81
+ $X2=3.06 $Y2=1.66
r206 11 12 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=3.06 $Y=1.81
+ $X2=3.06 $Y2=2
r207 7 35 11.7719 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=2.825 $Y=1.48
+ $X2=2.825 $Y2=1.66
r208 7 9 346.117 $w=1.5e-07 $l=6.75e-07 $layer=POLY_cond $X=2.825 $Y=1.48
+ $X2=2.825 $Y2=0.805
r209 2 41 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=1.23
+ $Y=2.245 $X2=1.375 $Y2=2.39
r210 1 51 182 $w=1.7e-07 $l=2.504e-07 $layer=licon1_NDIFF $count=1 $X=1.115
+ $Y=0.595 $X2=1.255 $Y2=0.785
.ends

.subckt PM_SKY130_FD_SC_LP__DFBBN_2%A_1746_137# 1 2 7 9 14 18 22 23 27 29 31 32
+ 34 36 39 43 45 46 47 51 55 58 59 62 64 65 70 71 72 74 79 81 82
c178 82 0 1.68582e-19 $X=11.96 $Y=1.185
c179 62 0 1.38329e-19 $X=11.88 $Y=2.2
c180 46 0 1.41247e-19 $X=13.45 $Y=1.26
c181 43 0 1.31498e-19 $X=8.96 $Y=1.385
r182 81 82 30.474 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=11.96 $Y=1.26
+ $X2=11.96 $Y2=1.185
r183 75 84 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=11.96 $Y=1.35
+ $X2=11.96 $Y2=1.515
r184 75 81 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=11.96 $Y=1.35
+ $X2=11.96 $Y2=1.26
r185 74 77 8.65224 $w=2.63e-07 $l=1.65e-07 $layer=LI1_cond $X=11.927 $Y=1.35
+ $X2=11.927 $Y2=1.515
r186 74 75 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.96
+ $Y=1.35 $X2=11.96 $Y2=1.35
r187 65 80 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=9.05 $Y=2.205
+ $X2=9.05 $Y2=2.37
r188 65 79 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=9.05 $Y=2.205
+ $X2=9.05 $Y2=2.04
r189 64 67 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=9.05 $Y=2.205 $X2=9.05
+ $Y2=2.285
r190 64 65 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.05
+ $Y=2.205 $X2=9.05 $Y2=2.205
r191 62 77 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=11.88 $Y=2.2
+ $X2=11.88 $Y2=1.515
r192 60 72 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.475 $Y=2.285
+ $X2=10.39 $Y2=2.285
r193 59 62 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=11.795 $Y=2.285
+ $X2=11.88 $Y2=2.2
r194 59 60 86.1176 $w=1.68e-07 $l=1.32e-06 $layer=LI1_cond $X=11.795 $Y=2.285
+ $X2=10.475 $Y2=2.285
r195 58 72 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.39 $Y=2.2
+ $X2=10.39 $Y2=2.285
r196 58 71 67.5241 $w=1.68e-07 $l=1.035e-06 $layer=LI1_cond $X=10.39 $Y=2.2
+ $X2=10.39 $Y2=1.165
r197 53 71 8.64139 $w=3.38e-07 $l=1.7e-07 $layer=LI1_cond $X=10.305 $Y=0.995
+ $X2=10.305 $Y2=1.165
r198 53 55 3.55902 $w=3.38e-07 $l=1.05e-07 $layer=LI1_cond $X=10.305 $Y=0.995
+ $X2=10.305 $Y2=0.89
r199 52 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.115 $Y=2.285
+ $X2=9.95 $Y2=2.285
r200 51 72 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.305 $Y=2.285
+ $X2=10.39 $Y2=2.285
r201 51 52 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=10.305 $Y=2.285
+ $X2=10.115 $Y2=2.285
r202 48 67 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.215 $Y=2.285
+ $X2=9.05 $Y2=2.285
r203 47 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.785 $Y=2.285
+ $X2=9.95 $Y2=2.285
r204 47 48 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=9.785 $Y=2.285
+ $X2=9.215 $Y2=2.285
r205 41 43 79.4787 $w=1.5e-07 $l=1.55e-07 $layer=POLY_cond $X=8.805 $Y=1.385
+ $X2=8.96 $Y2=1.385
r206 37 46 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=13.45 $Y=1.335
+ $X2=13.45 $Y2=1.26
r207 37 39 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=13.45 $Y=1.335
+ $X2=13.45 $Y2=2.155
r208 34 46 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=13.45 $Y=1.185
+ $X2=13.45 $Y2=1.26
r209 34 36 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=13.45 $Y=1.185
+ $X2=13.45 $Y2=0.865
r210 33 45 12.05 $w=1.5e-07 $l=8e-08 $layer=POLY_cond $X=12.535 $Y=1.26
+ $X2=12.455 $Y2=1.26
r211 32 46 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=13.375 $Y=1.26
+ $X2=13.45 $Y2=1.26
r212 32 33 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=13.375 $Y=1.26
+ $X2=12.535 $Y2=1.26
r213 29 45 12.05 $w=1.5e-07 $l=7.74597e-08 $layer=POLY_cond $X=12.46 $Y=1.185
+ $X2=12.455 $Y2=1.26
r214 29 31 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=12.46 $Y=1.185
+ $X2=12.46 $Y2=0.655
r215 25 45 12.05 $w=1.5e-07 $l=7.74597e-08 $layer=POLY_cond $X=12.45 $Y=1.335
+ $X2=12.455 $Y2=1.26
r216 25 27 515.33 $w=1.5e-07 $l=1.005e-06 $layer=POLY_cond $X=12.45 $Y=1.335
+ $X2=12.45 $Y2=2.34
r217 24 81 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=12.125 $Y=1.26
+ $X2=11.96 $Y2=1.26
r218 23 45 12.05 $w=1.5e-07 $l=8e-08 $layer=POLY_cond $X=12.375 $Y=1.26
+ $X2=12.455 $Y2=1.26
r219 23 24 128.191 $w=1.5e-07 $l=2.5e-07 $layer=POLY_cond $X=12.375 $Y=1.26
+ $X2=12.125 $Y2=1.26
r220 22 82 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=12.03 $Y=0.655
+ $X2=12.03 $Y2=1.185
r221 18 84 423.032 $w=1.5e-07 $l=8.25e-07 $layer=POLY_cond $X=12.02 $Y=2.34
+ $X2=12.02 $Y2=1.515
r222 14 80 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=8.99 $Y=2.74
+ $X2=8.99 $Y2=2.37
r223 10 43 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.96 $Y=1.46
+ $X2=8.96 $Y2=1.385
r224 10 79 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=8.96 $Y=1.46
+ $X2=8.96 $Y2=2.04
r225 7 41 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.805 $Y=1.31
+ $X2=8.805 $Y2=1.385
r226 7 9 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=8.805 $Y=1.31
+ $X2=8.805 $Y2=1.025
r227 2 70 300 $w=1.7e-07 $l=2.86575e-07 $layer=licon1_PDIFF $count=2 $X=9.81
+ $Y=2.14 $X2=9.95 $Y2=2.365
r228 1 55 182 $w=1.7e-07 $l=3.89776e-07 $layer=licon1_NDIFF $count=1 $X=10
+ $Y=0.595 $X2=10.22 $Y2=0.89
.ends

.subckt PM_SKY130_FD_SC_LP__DFBBN_2%A_1542_428# 1 2 7 9 14 15 16 19 23 26 27 29
+ 30 37
c96 30 0 9.01378e-20 $X=9.955 $Y=1.205
c97 27 0 1.71827e-19 $X=7.905 $Y=2.12
c98 26 0 2.25888e-20 $X=7.85 $Y=2.415
r99 33 37 28.8521 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=9.96 $Y=1.51
+ $X2=10.125 $Y2=1.51
r100 33 34 6.12014 $w=3.3e-07 $l=3.5e-08 $layer=POLY_cond $X=9.96 $Y=1.51
+ $X2=9.925 $Y2=1.51
r101 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.96
+ $Y=1.51 $X2=9.96 $Y2=1.51
r102 30 32 13.7306 $w=2.71e-07 $l=3.05e-07 $layer=LI1_cond $X=9.955 $Y=1.205
+ $X2=9.955 $Y2=1.51
r103 26 27 12.2403 $w=4.38e-07 $l=2.95e-07 $layer=LI1_cond $X=7.905 $Y=2.415
+ $X2=7.905 $Y2=2.12
r104 24 29 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.285 $Y=1.205
+ $X2=8.12 $Y2=1.205
r105 23 30 3.46554 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=9.785 $Y=1.205
+ $X2=9.955 $Y2=1.205
r106 23 24 97.861 $w=1.68e-07 $l=1.5e-06 $layer=LI1_cond $X=9.785 $Y=1.205
+ $X2=8.285 $Y2=1.205
r107 21 29 3.70735 $w=2.5e-07 $l=1.18427e-07 $layer=LI1_cond $X=8.04 $Y=1.29
+ $X2=8.12 $Y2=1.205
r108 21 27 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=8.04 $Y=1.29
+ $X2=8.04 $Y2=2.12
r109 17 29 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=8.12 $Y=1.12
+ $X2=8.12 $Y2=1.205
r110 17 19 13.2706 $w=3.28e-07 $l=3.8e-07 $layer=LI1_cond $X=8.12 $Y=1.12
+ $X2=8.12 $Y2=0.74
r111 15 16 53.9552 $w=1.9e-07 $l=1.5e-07 $layer=POLY_cond $X=10.145 $Y=1.915
+ $X2=10.145 $Y2=2.065
r112 14 16 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=10.165 $Y=2.56
+ $X2=10.165 $Y2=2.065
r113 10 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.125 $Y=1.675
+ $X2=10.125 $Y2=1.51
r114 10 15 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=10.125 $Y=1.675
+ $X2=10.125 $Y2=1.915
r115 7 34 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.925 $Y=1.345
+ $X2=9.925 $Y2=1.51
r116 7 9 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=9.925 $Y=1.345
+ $X2=9.925 $Y2=0.915
r117 2 26 600 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=1 $X=7.71
+ $Y=2.14 $X2=7.85 $Y2=2.415
r118 1 19 91 $w=1.7e-07 $l=4.41588e-07 $layer=licon1_NDIFF $count=2 $X=7.745
+ $Y=0.595 $X2=8.12 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_LP__DFBBN_2%A_1191_21# 1 2 9 11 13 14 18 21 26 27 28 29
+ 30 32 36
c110 30 0 6.64683e-20 $X=10.985 $Y=1.855
c111 26 0 7.76368e-20 $X=10.82 $Y=1.51
c112 9 0 1.70135e-19 $X=6.03 $Y=0.955
r113 38 40 1.74861 $w=3.3e-07 $l=1e-08 $layer=POLY_cond $X=10.515 $Y=1.51
+ $X2=10.525 $Y2=1.51
r114 34 36 16.5952 $w=2.48e-07 $l=3.6e-07 $layer=LI1_cond $X=11.345 $Y=0.83
+ $X2=11.345 $Y2=0.47
r115 30 32 10.826 $w=3.28e-07 $l=3.1e-07 $layer=LI1_cond $X=10.985 $Y=1.855
+ $X2=11.295 $Y2=1.855
r116 28 34 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=11.22 $Y=0.915
+ $X2=11.345 $Y2=0.83
r117 28 29 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=11.22 $Y=0.915
+ $X2=10.985 $Y2=0.915
r118 27 40 51.5841 $w=3.3e-07 $l=2.95e-07 $layer=POLY_cond $X=10.82 $Y=1.51
+ $X2=10.525 $Y2=1.51
r119 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.82
+ $Y=1.51 $X2=10.82 $Y2=1.51
r120 24 30 6.71475 $w=3.35e-07 $l=4.04166e-07 $layer=LI1_cond $X=10.82 $Y=1.525
+ $X2=10.985 $Y2=1.855
r121 24 26 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=10.82 $Y=1.525
+ $X2=10.82 $Y2=1.51
r122 23 29 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=10.82 $Y=1
+ $X2=10.985 $Y2=0.915
r123 23 26 17.8105 $w=3.28e-07 $l=5.1e-07 $layer=LI1_cond $X=10.82 $Y=1
+ $X2=10.82 $Y2=1.51
r124 19 40 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.525 $Y=1.675
+ $X2=10.525 $Y2=1.51
r125 19 21 453.798 $w=1.5e-07 $l=8.85e-07 $layer=POLY_cond $X=10.525 $Y=1.675
+ $X2=10.525 $Y2=2.56
r126 16 38 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.515 $Y=1.345
+ $X2=10.515 $Y2=1.51
r127 16 18 351.245 $w=1.5e-07 $l=6.85e-07 $layer=POLY_cond $X=10.515 $Y=1.345
+ $X2=10.515 $Y2=0.66
r128 15 18 207.67 $w=1.5e-07 $l=4.05e-07 $layer=POLY_cond $X=10.515 $Y=0.255
+ $X2=10.515 $Y2=0.66
r129 13 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=10.44 $Y=0.18
+ $X2=10.515 $Y2=0.255
r130 13 14 2222.84 $w=1.5e-07 $l=4.335e-06 $layer=POLY_cond $X=10.44 $Y=0.18
+ $X2=6.105 $Y2=0.18
r131 9 11 697.362 $w=1.5e-07 $l=1.36e-06 $layer=POLY_cond $X=6.03 $Y=0.955
+ $X2=6.03 $Y2=2.315
r132 7 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.03 $Y=0.255
+ $X2=6.105 $Y2=0.18
r133 7 9 358.936 $w=1.5e-07 $l=7e-07 $layer=POLY_cond $X=6.03 $Y=0.255 $X2=6.03
+ $Y2=0.955
r134 2 32 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=11.155
+ $Y=1.71 $X2=11.295 $Y2=1.855
r135 1 36 182 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_NDIFF $count=1 $X=11.16
+ $Y=0.235 $X2=11.305 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_LP__DFBBN_2%RESET_B 2 5 9 13 15 21 22
c38 22 0 1.68582e-19 $X=11.51 $Y=1.345
c39 5 0 7.76368e-20 $X=11.51 $Y=2.03
r40 20 22 20.109 $w=3.3e-07 $l=1.15e-07 $layer=POLY_cond $X=11.395 $Y=1.345
+ $X2=11.51 $Y2=1.345
r41 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.395
+ $Y=1.345 $X2=11.395 $Y2=1.345
r42 17 20 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=11.305 $Y=1.345
+ $X2=11.395 $Y2=1.345
r43 15 21 4.01609 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=11.28 $Y=1.345
+ $X2=11.395 $Y2=1.345
r44 11 13 110.245 $w=1.5e-07 $l=2.15e-07 $layer=POLY_cond $X=11.305 $Y=0.87
+ $X2=11.52 $Y2=0.87
r45 7 13 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=11.52 $Y=0.795
+ $X2=11.52 $Y2=0.87
r46 7 9 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=11.52 $Y=0.795
+ $X2=11.52 $Y2=0.445
r47 3 22 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=11.51 $Y=1.51
+ $X2=11.51 $Y2=1.345
r48 3 5 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=11.51 $Y=1.51
+ $X2=11.51 $Y2=2.03
r49 2 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=11.305 $Y=1.18
+ $X2=11.305 $Y2=1.345
r50 1 11 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=11.305 $Y=0.945
+ $X2=11.305 $Y2=0.87
r51 1 2 120.5 $w=1.5e-07 $l=2.35e-07 $layer=POLY_cond $X=11.305 $Y=0.945
+ $X2=11.305 $Y2=1.18
.ends

.subckt PM_SKY130_FD_SC_LP__DFBBN_2%A_2618_131# 1 2 9 13 15 19 23 25 28 32 36 39
+ 40
c76 39 0 1.41247e-19 $X=13.235 $Y=1.44
r77 40 41 30.474 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=13.93 $Y=1.35
+ $X2=13.93 $Y2=1.275
r78 37 43 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=13.93 $Y=1.44
+ $X2=13.93 $Y2=1.605
r79 37 40 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=13.93 $Y=1.44
+ $X2=13.93 $Y2=1.35
r80 36 37 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=13.93
+ $Y=1.44 $X2=13.93 $Y2=1.44
r81 34 39 1.34256 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=13.4 $Y=1.44
+ $X2=13.235 $Y2=1.44
r82 34 36 18.5089 $w=3.28e-07 $l=5.3e-07 $layer=LI1_cond $X=13.4 $Y=1.44
+ $X2=13.93 $Y2=1.44
r83 30 39 5.16603 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=13.235 $Y=1.605
+ $X2=13.235 $Y2=1.44
r84 30 32 13.0959 $w=3.28e-07 $l=3.75e-07 $layer=LI1_cond $X=13.235 $Y=1.605
+ $X2=13.235 $Y2=1.98
r85 26 39 5.16603 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=13.235 $Y=1.275
+ $X2=13.235 $Y2=1.44
r86 26 28 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=13.235 $Y=1.275
+ $X2=13.235 $Y2=0.865
r87 21 25 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=14.39 $Y=1.425
+ $X2=14.39 $Y2=1.35
r88 21 23 533.277 $w=1.5e-07 $l=1.04e-06 $layer=POLY_cond $X=14.39 $Y=1.425
+ $X2=14.39 $Y2=2.465
r89 17 25 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=14.39 $Y=1.275
+ $X2=14.39 $Y2=1.35
r90 17 19 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=14.39 $Y=1.275
+ $X2=14.39 $Y2=0.655
r91 16 40 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=14.095 $Y=1.35
+ $X2=13.93 $Y2=1.35
r92 15 25 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=14.315 $Y=1.35
+ $X2=14.39 $Y2=1.35
r93 15 16 112.809 $w=1.5e-07 $l=2.2e-07 $layer=POLY_cond $X=14.315 $Y=1.35
+ $X2=14.095 $Y2=1.35
r94 13 43 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=13.96 $Y=2.465
+ $X2=13.96 $Y2=1.605
r95 9 41 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=13.96 $Y=0.655
+ $X2=13.96 $Y2=1.275
r96 2 32 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=13.09
+ $Y=1.835 $X2=13.235 $Y2=1.98
r97 1 28 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=13.09
+ $Y=0.655 $X2=13.235 $Y2=0.865
.ends

.subckt PM_SKY130_FD_SC_LP__DFBBN_2%VPWR 1 2 3 4 5 6 7 8 9 10 31 33 37 41 45 49
+ 53 57 61 67 71 73 76 77 79 80 81 96 103 108 113 118 123 128 137 140 143 146
+ 149 152 156
r154 155 156 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.64 $Y=3.33
+ $X2=14.64 $Y2=3.33
r155 152 153 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.68 $Y=3.33
+ $X2=13.68 $Y2=3.33
r156 149 150 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.72 $Y=3.33
+ $X2=12.72 $Y2=3.33
r157 146 147 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.76 $Y=3.33
+ $X2=11.76 $Y2=3.33
r158 143 144 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=3.33
+ $X2=10.8 $Y2=3.33
r159 140 141 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r160 137 138 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r161 134 135 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r162 132 156 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=14.16 $Y=3.33
+ $X2=14.64 $Y2=3.33
r163 132 153 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=14.16 $Y=3.33
+ $X2=13.68 $Y2=3.33
r164 131 132 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.16 $Y=3.33
+ $X2=14.16 $Y2=3.33
r165 129 152 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=13.83 $Y=3.33
+ $X2=13.705 $Y2=3.33
r166 129 131 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=13.83 $Y=3.33
+ $X2=14.16 $Y2=3.33
r167 128 155 4.01803 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=14.52 $Y=3.33
+ $X2=14.7 $Y2=3.33
r168 128 131 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=14.52 $Y=3.33
+ $X2=14.16 $Y2=3.33
r169 127 153 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.2 $Y=3.33
+ $X2=13.68 $Y2=3.33
r170 127 150 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.2 $Y=3.33
+ $X2=12.72 $Y2=3.33
r171 126 127 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.2 $Y=3.33
+ $X2=13.2 $Y2=3.33
r172 124 149 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=12.84 $Y=3.33
+ $X2=12.715 $Y2=3.33
r173 124 126 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=12.84 $Y=3.33
+ $X2=13.2 $Y2=3.33
r174 123 152 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=13.58 $Y=3.33
+ $X2=13.705 $Y2=3.33
r175 123 126 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=13.58 $Y=3.33
+ $X2=13.2 $Y2=3.33
r176 122 150 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.24 $Y=3.33
+ $X2=12.72 $Y2=3.33
r177 122 147 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.24 $Y=3.33
+ $X2=11.76 $Y2=3.33
r178 121 122 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.24 $Y=3.33
+ $X2=12.24 $Y2=3.33
r179 119 146 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.97 $Y=3.33
+ $X2=11.805 $Y2=3.33
r180 119 121 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=11.97 $Y=3.33
+ $X2=12.24 $Y2=3.33
r181 118 149 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=12.59 $Y=3.33
+ $X2=12.715 $Y2=3.33
r182 118 121 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=12.59 $Y=3.33
+ $X2=12.24 $Y2=3.33
r183 117 147 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=3.33
+ $X2=11.76 $Y2=3.33
r184 117 144 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=3.33
+ $X2=10.8 $Y2=3.33
r185 116 117 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.28 $Y=3.33
+ $X2=11.28 $Y2=3.33
r186 114 143 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.905 $Y=3.33
+ $X2=10.74 $Y2=3.33
r187 114 116 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=10.905 $Y=3.33
+ $X2=11.28 $Y2=3.33
r188 113 146 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.64 $Y=3.33
+ $X2=11.805 $Y2=3.33
r189 113 116 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=11.64 $Y=3.33
+ $X2=11.28 $Y2=3.33
r190 112 144 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=3.33
+ $X2=10.8 $Y2=3.33
r191 112 141 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=10.32 $Y=3.33
+ $X2=9.36 $Y2=3.33
r192 111 112 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.32 $Y=3.33
+ $X2=10.32 $Y2=3.33
r193 109 140 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.605 $Y=3.33
+ $X2=9.48 $Y2=3.33
r194 109 111 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=9.605 $Y=3.33
+ $X2=10.32 $Y2=3.33
r195 108 143 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.575 $Y=3.33
+ $X2=10.74 $Y2=3.33
r196 108 111 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=10.575 $Y=3.33
+ $X2=10.32 $Y2=3.33
r197 107 138 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=6.48 $Y2=3.33
r198 106 107 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r199 104 137 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.565 $Y=3.33
+ $X2=6.4 $Y2=3.33
r200 104 106 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=6.565 $Y=3.33
+ $X2=6.96 $Y2=3.33
r201 103 140 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.355 $Y=3.33
+ $X2=9.48 $Y2=3.33
r202 103 106 156.251 $w=1.68e-07 $l=2.395e-06 $layer=LI1_cond $X=9.355 $Y=3.33
+ $X2=6.96 $Y2=3.33
r203 102 138 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33
+ $X2=6.48 $Y2=3.33
r204 101 102 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r205 99 102 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=6 $Y2=3.33
r206 98 101 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=5.04 $Y=3.33 $X2=6
+ $Y2=3.33
r207 98 99 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r208 96 137 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.235 $Y=3.33
+ $X2=6.4 $Y2=3.33
r209 96 101 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=6.235 $Y=3.33
+ $X2=6 $Y2=3.33
r210 95 99 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.04 $Y2=3.33
r211 94 95 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r212 92 95 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=4.56 $Y2=3.33
r213 91 94 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=2.16 $Y=3.33
+ $X2=4.56 $Y2=3.33
r214 91 92 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r215 89 92 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r216 88 89 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r217 86 89 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r218 86 135 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r219 85 88 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r220 85 86 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r221 83 134 4.67962 $w=1.7e-07 $l=2.35e-07 $layer=LI1_cond $X=0.47 $Y=3.33
+ $X2=0.235 $Y2=3.33
r222 83 85 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=0.47 $Y=3.33
+ $X2=0.72 $Y2=3.33
r223 81 141 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=9.36 $Y2=3.33
r224 81 107 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=6.96 $Y2=3.33
r225 79 94 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=4.63 $Y=3.33 $X2=4.56
+ $Y2=3.33
r226 79 80 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.63 $Y=3.33
+ $X2=4.795 $Y2=3.33
r227 78 98 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=4.96 $Y=3.33 $X2=5.04
+ $Y2=3.33
r228 78 80 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.96 $Y=3.33
+ $X2=4.795 $Y2=3.33
r229 76 88 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=1.72 $Y=3.33 $X2=1.68
+ $Y2=3.33
r230 76 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.72 $Y=3.33
+ $X2=1.885 $Y2=3.33
r231 75 91 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=2.05 $Y=3.33
+ $X2=2.16 $Y2=3.33
r232 75 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.05 $Y=3.33
+ $X2=1.885 $Y2=3.33
r233 71 155 3.12513 $w=2.5e-07 $l=1.09087e-07 $layer=LI1_cond $X=14.645 $Y=3.245
+ $X2=14.7 $Y2=3.33
r234 71 73 43.5623 $w=2.48e-07 $l=9.45e-07 $layer=LI1_cond $X=14.645 $Y=3.245
+ $X2=14.645 $Y2=2.3
r235 67 70 22.3574 $w=2.48e-07 $l=4.85e-07 $layer=LI1_cond $X=13.705 $Y=1.98
+ $X2=13.705 $Y2=2.465
r236 65 152 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=13.705 $Y=3.245
+ $X2=13.705 $Y2=3.33
r237 65 70 35.9562 $w=2.48e-07 $l=7.8e-07 $layer=LI1_cond $X=13.705 $Y=3.245
+ $X2=13.705 $Y2=2.465
r238 61 64 44.7148 $w=2.48e-07 $l=9.7e-07 $layer=LI1_cond $X=12.715 $Y=1.855
+ $X2=12.715 $Y2=2.825
r239 59 149 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=12.715 $Y=3.245
+ $X2=12.715 $Y2=3.33
r240 59 64 19.361 $w=2.48e-07 $l=4.2e-07 $layer=LI1_cond $X=12.715 $Y=3.245
+ $X2=12.715 $Y2=2.825
r241 55 146 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=11.805 $Y=3.245
+ $X2=11.805 $Y2=3.33
r242 55 57 16.5882 $w=3.28e-07 $l=4.75e-07 $layer=LI1_cond $X=11.805 $Y=3.245
+ $X2=11.805 $Y2=2.77
r243 51 143 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.74 $Y=3.245
+ $X2=10.74 $Y2=3.33
r244 51 53 16.4136 $w=3.28e-07 $l=4.7e-07 $layer=LI1_cond $X=10.74 $Y=3.245
+ $X2=10.74 $Y2=2.775
r245 47 140 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=9.48 $Y=3.245
+ $X2=9.48 $Y2=3.33
r246 47 49 21.6659 $w=2.48e-07 $l=4.7e-07 $layer=LI1_cond $X=9.48 $Y=3.245
+ $X2=9.48 $Y2=2.775
r247 43 137 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.4 $Y=3.245
+ $X2=6.4 $Y2=3.33
r248 43 45 42.0816 $w=3.28e-07 $l=1.205e-06 $layer=LI1_cond $X=6.4 $Y=3.245
+ $X2=6.4 $Y2=2.04
r249 39 80 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.795 $Y=3.245
+ $X2=4.795 $Y2=3.33
r250 39 41 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=4.795 $Y=3.245
+ $X2=4.795 $Y2=2.825
r251 35 77 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.885 $Y=3.245
+ $X2=1.885 $Y2=3.33
r252 35 37 29.8588 $w=3.28e-07 $l=8.55e-07 $layer=LI1_cond $X=1.885 $Y=3.245
+ $X2=1.885 $Y2=2.39
r253 31 134 3.08656 $w=3.3e-07 $l=1.14782e-07 $layer=LI1_cond $X=0.305 $Y=3.245
+ $X2=0.235 $Y2=3.33
r254 31 33 24.2711 $w=3.28e-07 $l=6.95e-07 $layer=LI1_cond $X=0.305 $Y=3.245
+ $X2=0.305 $Y2=2.55
r255 10 73 300 $w=1.7e-07 $l=5.30401e-07 $layer=licon1_PDIFF $count=2 $X=14.465
+ $Y=1.835 $X2=14.605 $Y2=2.3
r256 9 70 300 $w=1.7e-07 $l=7.31779e-07 $layer=licon1_PDIFF $count=2 $X=13.525
+ $Y=1.835 $X2=13.745 $Y2=2.465
r257 9 67 600 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_PDIFF $count=1 $X=13.525
+ $Y=1.835 $X2=13.745 $Y2=1.98
r258 8 64 400 $w=1.7e-07 $l=1.18763e-06 $layer=licon1_PDIFF $count=1 $X=12.525
+ $Y=1.71 $X2=12.675 $Y2=2.825
r259 8 61 400 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=12.525
+ $Y=1.71 $X2=12.675 $Y2=1.855
r260 7 57 600 $w=1.7e-07 $l=1.16482e-06 $layer=licon1_PDIFF $count=1 $X=11.585
+ $Y=1.71 $X2=11.805 $Y2=2.77
r261 6 53 600 $w=1.7e-07 $l=7.01516e-07 $layer=licon1_PDIFF $count=1 $X=10.6
+ $Y=2.14 $X2=10.74 $Y2=2.775
r262 5 49 600 $w=1.7e-07 $l=5.64358e-07 $layer=licon1_PDIFF $count=1 $X=9.065
+ $Y=2.53 $X2=9.52 $Y2=2.775
r263 4 45 300 $w=1.7e-07 $l=3.60278e-07 $layer=licon1_PDIFF $count=2 $X=6.105
+ $Y=1.895 $X2=6.4 $Y2=2.04
r264 3 41 600 $w=1.7e-07 $l=9.46573e-07 $layer=licon1_PDIFF $count=1 $X=4.095
+ $Y=2.245 $X2=4.795 $Y2=2.825
r265 2 37 300 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_PDIFF $count=2 $X=1.665
+ $Y=2.245 $X2=1.885 $Y2=2.39
r266 1 33 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=0.16
+ $Y=2.405 $X2=0.305 $Y2=2.55
.ends

.subckt PM_SKY130_FD_SC_LP__DFBBN_2%A_463_449# 1 2 9 12 14 17
r45 16 17 8.63679 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=2.677 $Y=1.13
+ $X2=2.677 $Y2=1.3
r46 12 14 16.0641 $w=2.81e-07 $l=4.55192e-07 $layer=LI1_cond $X=2.825 $Y=2.305
+ $X2=2.455 $Y2=2.495
r47 12 17 65.5668 $w=1.68e-07 $l=1.005e-06 $layer=LI1_cond $X=2.825 $Y=2.305
+ $X2=2.825 $Y2=1.3
r48 9 16 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=2.61 $Y=0.805
+ $X2=2.61 $Y2=1.13
r49 2 14 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=2.315
+ $Y=2.245 $X2=2.455 $Y2=2.455
r50 1 9 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.47
+ $Y=0.595 $X2=2.61 $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_LP__DFBBN_2%Q_N 1 2 7 9 16 17 18 21
r34 18 21 4.36531 $w=3.28e-07 $l=1.25e-07 $layer=LI1_cond $X=12.245 $Y=0.555
+ $X2=12.245 $Y2=0.43
r35 16 17 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=12.325 $Y=1.005
+ $X2=12.325 $Y2=1.695
r36 15 18 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=12.245 $Y=0.84
+ $X2=12.245 $Y2=0.555
r37 15 16 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=12.245 $Y=0.84
+ $X2=12.245 $Y2=1.005
r38 9 11 42.7734 $w=2.58e-07 $l=9.65e-07 $layer=LI1_cond $X=12.28 $Y=1.86
+ $X2=12.28 $Y2=2.825
r39 7 17 7.14225 $w=2.58e-07 $l=1.3e-07 $layer=LI1_cond $X=12.28 $Y=1.825
+ $X2=12.28 $Y2=1.695
r40 7 9 1.55137 $w=2.58e-07 $l=3.5e-08 $layer=LI1_cond $X=12.28 $Y=1.825
+ $X2=12.28 $Y2=1.86
r41 2 11 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=12.095
+ $Y=1.71 $X2=12.235 $Y2=2.825
r42 2 9 400 $w=1.7e-07 $l=2.08567e-07 $layer=licon1_PDIFF $count=1 $X=12.095
+ $Y=1.71 $X2=12.235 $Y2=1.86
r43 1 21 91 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_NDIFF $count=2 $X=12.105
+ $Y=0.235 $X2=12.245 $Y2=0.43
.ends

.subckt PM_SKY130_FD_SC_LP__DFBBN_2%Q 1 2 9 15 16 17 18 24 30
r35 18 35 7.82962 $w=4.33e-07 $l=1.28e-07 $layer=LI1_cond $X=14.227 $Y=0.967
+ $X2=14.227 $Y2=1.095
r36 18 30 1.1127 $w=4.33e-07 $l=4.2e-08 $layer=LI1_cond $X=14.227 $Y=0.967
+ $X2=14.227 $Y2=0.925
r37 18 30 1.50167 $w=3.28e-07 $l=4.3e-08 $layer=LI1_cond $X=14.175 $Y=0.882
+ $X2=14.175 $Y2=0.925
r38 17 18 11.4197 $w=3.28e-07 $l=3.27e-07 $layer=LI1_cond $X=14.175 $Y=0.555
+ $X2=14.175 $Y2=0.882
r39 17 24 4.36531 $w=3.28e-07 $l=1.25e-07 $layer=LI1_cond $X=14.175 $Y=0.555
+ $X2=14.175 $Y2=0.43
r40 15 16 8.63679 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=14.227 $Y=1.785
+ $X2=14.227 $Y2=1.955
r41 15 35 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=14.36 $Y=1.785
+ $X2=14.36 $Y2=1.095
r42 9 11 32.1287 $w=3.28e-07 $l=9.2e-07 $layer=LI1_cond $X=14.175 $Y=1.98
+ $X2=14.175 $Y2=2.9
r43 9 16 0.873063 $w=3.28e-07 $l=2.5e-08 $layer=LI1_cond $X=14.175 $Y=1.98
+ $X2=14.175 $Y2=1.955
r44 2 11 400 $w=1.7e-07 $l=1.13284e-06 $layer=licon1_PDIFF $count=1 $X=14.035
+ $Y=1.835 $X2=14.175 $Y2=2.9
r45 2 9 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=14.035
+ $Y=1.835 $X2=14.175 $Y2=1.98
r46 1 24 91 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_NDIFF $count=2 $X=14.035
+ $Y=0.235 $X2=14.175 $Y2=0.43
.ends

.subckt PM_SKY130_FD_SC_LP__DFBBN_2%VGND 1 2 3 4 5 6 7 8 9 28 30 34 38 42 46 50
+ 56 60 64 66 69 70 71 73 85 92 100 105 110 115 124 127 130 133 136 139 143
r148 142 143 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.64 $Y=0
+ $X2=14.64 $Y2=0
r149 139 140 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.68 $Y=0
+ $X2=13.68 $Y2=0
r150 136 137 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.72 $Y=0
+ $X2=12.72 $Y2=0
r151 133 134 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.76 $Y=0
+ $X2=11.76 $Y2=0
r152 130 131 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=9.36 $Y=0
+ $X2=9.36 $Y2=0
r153 127 128 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=0
+ $X2=6.96 $Y2=0
r154 124 125 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0
+ $X2=1.68 $Y2=0
r155 121 122 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0
+ $X2=0.24 $Y2=0
r156 119 143 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=14.16 $Y=0
+ $X2=14.64 $Y2=0
r157 119 140 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=14.16 $Y=0
+ $X2=13.68 $Y2=0
r158 118 119 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.16 $Y=0
+ $X2=14.16 $Y2=0
r159 116 139 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=13.83 $Y=0
+ $X2=13.705 $Y2=0
r160 116 118 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=13.83 $Y=0
+ $X2=14.16 $Y2=0
r161 115 142 4.01803 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=14.52 $Y=0
+ $X2=14.7 $Y2=0
r162 115 118 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=14.52 $Y=0
+ $X2=14.16 $Y2=0
r163 114 140 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.2 $Y=0
+ $X2=13.68 $Y2=0
r164 114 137 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.2 $Y=0
+ $X2=12.72 $Y2=0
r165 113 114 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.2 $Y=0
+ $X2=13.2 $Y2=0
r166 111 136 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=12.84 $Y=0
+ $X2=12.715 $Y2=0
r167 111 113 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=12.84 $Y=0
+ $X2=13.2 $Y2=0
r168 110 139 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=13.58 $Y=0
+ $X2=13.705 $Y2=0
r169 110 113 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=13.58 $Y=0
+ $X2=13.2 $Y2=0
r170 109 137 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.24 $Y=0
+ $X2=12.72 $Y2=0
r171 109 134 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.24 $Y=0
+ $X2=11.76 $Y2=0
r172 108 109 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.24 $Y=0
+ $X2=12.24 $Y2=0
r173 106 133 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=11.9 $Y=0
+ $X2=11.775 $Y2=0
r174 106 108 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=11.9 $Y=0
+ $X2=12.24 $Y2=0
r175 105 136 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=12.59 $Y=0
+ $X2=12.715 $Y2=0
r176 105 108 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=12.59 $Y=0
+ $X2=12.24 $Y2=0
r177 104 134 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=0
+ $X2=11.76 $Y2=0
r178 104 131 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=11.28 $Y=0
+ $X2=9.36 $Y2=0
r179 103 104 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=11.28 $Y=0
+ $X2=11.28 $Y2=0
r180 101 130 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.365 $Y=0
+ $X2=9.2 $Y2=0
r181 101 103 124.936 $w=1.68e-07 $l=1.915e-06 $layer=LI1_cond $X=9.365 $Y=0
+ $X2=11.28 $Y2=0
r182 100 133 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=11.65 $Y=0
+ $X2=11.775 $Y2=0
r183 100 103 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=11.65 $Y=0
+ $X2=11.28 $Y2=0
r184 99 131 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=0
+ $X2=9.36 $Y2=0
r185 98 99 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.88 $Y=0 $X2=8.88
+ $Y2=0
r186 95 98 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=7.44 $Y=0 $X2=8.88
+ $Y2=0
r187 93 127 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.11 $Y=0
+ $X2=6.985 $Y2=0
r188 93 95 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=7.11 $Y=0 $X2=7.44
+ $Y2=0
r189 92 130 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.035 $Y=0 $X2=9.2
+ $Y2=0
r190 92 98 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=9.035 $Y=0
+ $X2=8.88 $Y2=0
r191 91 128 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0
+ $X2=6.96 $Y2=0
r192 90 91 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.48 $Y=0
+ $X2=6.48 $Y2=0
r193 88 91 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=4.56 $Y=0
+ $X2=6.48 $Y2=0
r194 87 90 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=4.56 $Y=0 $X2=6.48
+ $Y2=0
r195 87 88 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.56 $Y=0
+ $X2=4.56 $Y2=0
r196 85 127 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.86 $Y=0
+ $X2=6.985 $Y2=0
r197 85 90 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=6.86 $Y=0 $X2=6.48
+ $Y2=0
r198 84 88 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=4.56
+ $Y2=0
r199 83 84 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.08 $Y=0
+ $X2=4.08 $Y2=0
r200 81 84 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=2.16 $Y=0
+ $X2=4.08 $Y2=0
r201 81 125 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0
+ $X2=1.68 $Y2=0
r202 80 83 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=2.16 $Y=0 $X2=4.08
+ $Y2=0
r203 80 81 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.16 $Y=0
+ $X2=2.16 $Y2=0
r204 78 124 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.93 $Y=0
+ $X2=1.765 $Y2=0
r205 78 80 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=1.93 $Y=0 $X2=2.16
+ $Y2=0
r206 77 125 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0
+ $X2=1.68 $Y2=0
r207 77 122 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0
+ $X2=0.24 $Y2=0
r208 76 77 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r209 74 121 4.01803 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=0.36 $Y=0 $X2=0.18
+ $Y2=0
r210 74 76 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=0.36 $Y=0 $X2=0.72
+ $Y2=0
r211 73 124 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.6 $Y=0 $X2=1.765
+ $Y2=0
r212 73 76 57.4118 $w=1.68e-07 $l=8.8e-07 $layer=LI1_cond $X=1.6 $Y=0 $X2=0.72
+ $Y2=0
r213 71 99 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=7.44 $Y=0
+ $X2=8.88 $Y2=0
r214 71 128 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0
+ $X2=6.96 $Y2=0
r215 71 95 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r216 69 83 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=4.205 $Y=0
+ $X2=4.08 $Y2=0
r217 69 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.205 $Y=0 $X2=4.37
+ $Y2=0
r218 68 87 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=4.535 $Y=0 $X2=4.56
+ $Y2=0
r219 68 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.535 $Y=0 $X2=4.37
+ $Y2=0
r220 64 142 3.12513 $w=2.5e-07 $l=1.09087e-07 $layer=LI1_cond $X=14.645 $Y=0.085
+ $X2=14.7 $Y2=0
r221 64 66 18.2086 $w=2.48e-07 $l=3.95e-07 $layer=LI1_cond $X=14.645 $Y=0.085
+ $X2=14.645 $Y2=0.48
r222 60 62 25.3537 $w=2.48e-07 $l=5.5e-07 $layer=LI1_cond $X=13.705 $Y=0.38
+ $X2=13.705 $Y2=0.93
r223 58 139 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=13.705 $Y=0.085
+ $X2=13.705 $Y2=0
r224 58 60 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=13.705 $Y=0.085
+ $X2=13.705 $Y2=0.38
r225 54 136 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=12.715 $Y=0.085
+ $X2=12.715 $Y2=0
r226 54 56 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=12.715 $Y=0.085
+ $X2=12.715 $Y2=0.38
r227 50 52 20.9745 $w=2.48e-07 $l=4.55e-07 $layer=LI1_cond $X=11.775 $Y=0.38
+ $X2=11.775 $Y2=0.835
r228 48 133 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=11.775 $Y=0.085
+ $X2=11.775 $Y2=0
r229 48 50 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=11.775 $Y=0.085
+ $X2=11.775 $Y2=0.38
r230 44 130 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.2 $Y=0.085
+ $X2=9.2 $Y2=0
r231 44 46 23.3981 $w=3.28e-07 $l=6.7e-07 $layer=LI1_cond $X=9.2 $Y=0.085
+ $X2=9.2 $Y2=0.755
r232 40 127 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.985 $Y=0.085
+ $X2=6.985 $Y2=0
r233 40 42 30.194 $w=2.48e-07 $l=6.55e-07 $layer=LI1_cond $X=6.985 $Y=0.085
+ $X2=6.985 $Y2=0.74
r234 36 70 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.37 $Y=0.085
+ $X2=4.37 $Y2=0
r235 36 38 17.112 $w=3.28e-07 $l=4.9e-07 $layer=LI1_cond $X=4.37 $Y=0.085
+ $X2=4.37 $Y2=0.575
r236 32 124 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.765 $Y=0.085
+ $X2=1.765 $Y2=0
r237 32 34 24.4458 $w=3.28e-07 $l=7e-07 $layer=LI1_cond $X=1.765 $Y=0.085
+ $X2=1.765 $Y2=0.785
r238 28 121 3.12513 $w=2.5e-07 $l=1.09087e-07 $layer=LI1_cond $X=0.235 $Y=0.085
+ $X2=0.18 $Y2=0
r239 28 30 18.9001 $w=2.48e-07 $l=4.1e-07 $layer=LI1_cond $X=0.235 $Y=0.085
+ $X2=0.235 $Y2=0.495
r240 9 66 182 $w=1.7e-07 $l=3.07124e-07 $layer=licon1_NDIFF $count=1 $X=14.465
+ $Y=0.235 $X2=14.605 $Y2=0.48
r241 8 62 182 $w=1.7e-07 $l=3.68951e-07 $layer=licon1_NDIFF $count=1 $X=13.525
+ $Y=0.655 $X2=13.745 $Y2=0.93
r242 8 60 182 $w=1.7e-07 $l=3.68951e-07 $layer=licon1_NDIFF $count=1 $X=13.525
+ $Y=0.655 $X2=13.745 $Y2=0.38
r243 7 56 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=12.535
+ $Y=0.235 $X2=12.675 $Y2=0.38
r244 6 52 182 $w=1.7e-07 $l=7.01427e-07 $layer=licon1_NDIFF $count=1 $X=11.595
+ $Y=0.235 $X2=11.815 $Y2=0.835
r245 6 50 182 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_NDIFF $count=1 $X=11.595
+ $Y=0.235 $X2=11.815 $Y2=0.38
r246 5 46 182 $w=1.7e-07 $l=3.48712e-07 $layer=licon1_NDIFF $count=1 $X=8.88
+ $Y=0.815 $X2=9.2 $Y2=0.755
r247 4 42 182 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=1 $X=6.8
+ $Y=0.595 $X2=6.945 $Y2=0.74
r248 3 38 182 $w=1.7e-07 $l=3.01247e-07 $layer=licon1_NDIFF $count=1 $X=4.095
+ $Y=0.52 $X2=4.37 $Y2=0.575
r249 2 34 182 $w=1.7e-07 $l=3.00333e-07 $layer=licon1_NDIFF $count=1 $X=1.545
+ $Y=0.595 $X2=1.765 $Y2=0.785
r250 1 30 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.285 $X2=0.275 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__DFBBN_2%A_1018_60# 1 2 7 12 15
c22 15 0 1.70135e-19 $X=6.245 $Y=0.78
r23 10 12 8.4794 $w=3.43e-07 $l=1.65e-07 $layer=LI1_cond $X=5.23 $Y=0.787
+ $X2=5.395 $Y2=0.787
r24 7 15 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.16 $Y=0.7 $X2=6.245
+ $Y2=0.7
r25 7 12 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=6.16 $Y=0.7
+ $X2=5.395 $Y2=0.7
r26 2 15 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=6.105
+ $Y=0.635 $X2=6.245 $Y2=0.78
r27 1 10 182 $w=1.7e-07 $l=5.10221e-07 $layer=licon1_NDIFF $count=1 $X=5.09
+ $Y=0.3 $X2=5.23 $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_LP__DFBBN_2%A_1911_119# 1 2 9 11 12 13
c32 1 0 9.01378e-20 $X=9.555 $Y=0.595
r33 13 16 6.22319 $w=2.48e-07 $l=1.35e-07 $layer=LI1_cond $X=10.78 $Y=0.35
+ $X2=10.78 $Y2=0.485
r34 11 13 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.655 $Y=0.35
+ $X2=10.78 $Y2=0.35
r35 11 12 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=10.655 $Y=0.35
+ $X2=9.875 $Y2=0.35
r36 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=9.71 $Y=0.435
+ $X2=9.875 $Y2=0.35
r37 7 9 11.1752 $w=3.28e-07 $l=3.2e-07 $layer=LI1_cond $X=9.71 $Y=0.435 $X2=9.71
+ $Y2=0.755
r38 2 16 182 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_NDIFF $count=1 $X=10.59
+ $Y=0.34 $X2=10.74 $Y2=0.485
r39 1 9 182 $w=1.7e-07 $l=2.24499e-07 $layer=licon1_NDIFF $count=1 $X=9.555
+ $Y=0.595 $X2=9.71 $Y2=0.755
.ends

