* File: sky130_fd_sc_lp__a41o_4.pxi.spice
* Created: Fri Aug 28 10:02:54 2020
* 
x_PM_SKY130_FD_SC_LP__A41O_4%A_100_23# N_A_100_23#_M1013_d N_A_100_23#_M1017_s
+ N_A_100_23#_M1007_d N_A_100_23#_M1002_g N_A_100_23#_M1000_g
+ N_A_100_23#_M1004_g N_A_100_23#_M1006_g N_A_100_23#_M1016_g
+ N_A_100_23#_M1015_g N_A_100_23#_M1024_g N_A_100_23#_M1020_g
+ N_A_100_23#_c_131_n N_A_100_23#_c_227_p N_A_100_23#_c_132_n
+ N_A_100_23#_c_140_n N_A_100_23#_c_133_n N_A_100_23#_c_148_p
+ N_A_100_23#_c_134_n N_A_100_23#_c_135_n PM_SKY130_FD_SC_LP__A41O_4%A_100_23#
x_PM_SKY130_FD_SC_LP__A41O_4%B1 N_B1_c_243_n N_B1_M1013_g N_B1_c_244_n
+ N_B1_M1022_g N_B1_M1007_g N_B1_M1023_g B1 B1 N_B1_c_248_n
+ PM_SKY130_FD_SC_LP__A41O_4%B1
x_PM_SKY130_FD_SC_LP__A41O_4%A1 N_A1_c_294_n N_A1_M1017_g N_A1_M1001_g
+ N_A1_c_296_n N_A1_M1025_g N_A1_M1012_g A1 A1 N_A1_c_299_n
+ PM_SKY130_FD_SC_LP__A41O_4%A1
x_PM_SKY130_FD_SC_LP__A41O_4%A2 N_A2_c_344_n N_A2_M1003_g N_A2_M1008_g
+ N_A2_c_346_n N_A2_M1018_g N_A2_M1027_g A2 N_A2_c_349_n
+ PM_SKY130_FD_SC_LP__A41O_4%A2
x_PM_SKY130_FD_SC_LP__A41O_4%A3 N_A3_M1005_g N_A3_M1014_g N_A3_c_391_n
+ N_A3_M1011_g N_A3_c_392_n N_A3_c_393_n N_A3_c_394_n N_A3_M1026_g A3 A3
+ PM_SKY130_FD_SC_LP__A41O_4%A3
x_PM_SKY130_FD_SC_LP__A41O_4%A4 N_A4_M1010_g N_A4_c_442_n N_A4_c_443_n
+ N_A4_M1021_g N_A4_M1009_g N_A4_M1019_g A4 A4 A4 N_A4_c_447_n
+ PM_SKY130_FD_SC_LP__A41O_4%A4
x_PM_SKY130_FD_SC_LP__A41O_4%VPWR N_VPWR_M1000_s N_VPWR_M1006_s N_VPWR_M1020_s
+ N_VPWR_M1001_s N_VPWR_M1008_d N_VPWR_M1005_s N_VPWR_M1010_s N_VPWR_c_489_n
+ N_VPWR_c_490_n N_VPWR_c_491_n N_VPWR_c_492_n N_VPWR_c_493_n N_VPWR_c_494_n
+ N_VPWR_c_495_n N_VPWR_c_496_n N_VPWR_c_497_n N_VPWR_c_498_n N_VPWR_c_499_n
+ N_VPWR_c_500_n N_VPWR_c_501_n VPWR N_VPWR_c_502_n N_VPWR_c_503_n
+ N_VPWR_c_504_n N_VPWR_c_505_n N_VPWR_c_488_n N_VPWR_c_507_n N_VPWR_c_508_n
+ N_VPWR_c_509_n N_VPWR_c_510_n PM_SKY130_FD_SC_LP__A41O_4%VPWR
x_PM_SKY130_FD_SC_LP__A41O_4%X N_X_M1002_s N_X_M1016_s N_X_M1000_d N_X_M1015_d
+ N_X_c_608_n N_X_c_613_n N_X_c_614_n N_X_c_661_p N_X_c_646_n N_X_c_609_n
+ N_X_c_615_n N_X_c_660_p N_X_c_651_n N_X_c_610_n N_X_c_616_n X X N_X_c_611_n X
+ PM_SKY130_FD_SC_LP__A41O_4%X
x_PM_SKY130_FD_SC_LP__A41O_4%A_495_367# N_A_495_367#_M1007_s
+ N_A_495_367#_M1023_s N_A_495_367#_M1012_d N_A_495_367#_M1027_s
+ N_A_495_367#_M1014_d N_A_495_367#_M1021_d N_A_495_367#_c_666_n
+ N_A_495_367#_c_667_n N_A_495_367#_c_681_n N_A_495_367#_c_726_n
+ N_A_495_367#_c_668_n N_A_495_367#_c_669_n N_A_495_367#_c_730_n
+ N_A_495_367#_c_670_n N_A_495_367#_c_734_n N_A_495_367#_c_671_n
+ N_A_495_367#_c_738_n N_A_495_367#_c_672_n N_A_495_367#_c_673_n
+ N_A_495_367#_c_674_n N_A_495_367#_c_675_n N_A_495_367#_c_676_n
+ PM_SKY130_FD_SC_LP__A41O_4%A_495_367#
x_PM_SKY130_FD_SC_LP__A41O_4%VGND N_VGND_M1002_d N_VGND_M1004_d N_VGND_M1024_d
+ N_VGND_M1022_s N_VGND_M1009_s N_VGND_c_744_n N_VGND_c_745_n N_VGND_c_746_n
+ N_VGND_c_747_n N_VGND_c_748_n N_VGND_c_749_n N_VGND_c_750_n N_VGND_c_751_n
+ N_VGND_c_752_n N_VGND_c_753_n VGND N_VGND_c_754_n N_VGND_c_755_n
+ N_VGND_c_756_n N_VGND_c_757_n N_VGND_c_758_n N_VGND_c_759_n
+ PM_SKY130_FD_SC_LP__A41O_4%VGND
x_PM_SKY130_FD_SC_LP__A41O_4%A_667_47# N_A_667_47#_M1017_d N_A_667_47#_M1025_d
+ N_A_667_47#_M1018_d N_A_667_47#_c_849_n N_A_667_47#_c_856_n
+ N_A_667_47#_c_857_n N_A_667_47#_c_850_n PM_SKY130_FD_SC_LP__A41O_4%A_667_47#
x_PM_SKY130_FD_SC_LP__A41O_4%A_922_47# N_A_922_47#_M1003_s N_A_922_47#_M1011_s
+ N_A_922_47#_c_878_n PM_SKY130_FD_SC_LP__A41O_4%A_922_47#
x_PM_SKY130_FD_SC_LP__A41O_4%A_1115_47# N_A_1115_47#_M1011_d
+ N_A_1115_47#_M1026_d N_A_1115_47#_M1019_d N_A_1115_47#_c_894_n
+ N_A_1115_47#_c_902_n N_A_1115_47#_c_895_n N_A_1115_47#_c_896_n
+ N_A_1115_47#_c_904_n PM_SKY130_FD_SC_LP__A41O_4%A_1115_47#
cc_1 VNB N_A_100_23#_M1002_g 0.025885f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=0.665
cc_2 VNB N_A_100_23#_M1004_g 0.0213918f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=0.665
cc_3 VNB N_A_100_23#_M1016_g 0.0214129f $X=-0.19 $Y=-0.245 $X2=1.435 $Y2=0.665
cc_4 VNB N_A_100_23#_M1024_g 0.0232093f $X=-0.19 $Y=-0.245 $X2=1.865 $Y2=0.665
cc_5 VNB N_A_100_23#_c_131_n 0.0119992f $X=-0.19 $Y=-0.245 $X2=2.38 $Y2=1.49
cc_6 VNB N_A_100_23#_c_132_n 0.001949f $X=-0.19 $Y=-0.245 $X2=2.487 $Y2=1.405
cc_7 VNB N_A_100_23#_c_133_n 0.00830635f $X=-0.19 $Y=-0.245 $X2=3.89 $Y2=0.85
cc_8 VNB N_A_100_23#_c_134_n 0.00330644f $X=-0.19 $Y=-0.245 $X2=2.487 $Y2=1.49
cc_9 VNB N_A_100_23#_c_135_n 0.0729016f $X=-0.19 $Y=-0.245 $X2=1.865 $Y2=1.49
cc_10 VNB N_B1_c_243_n 0.0163189f $X=-0.19 $Y=-0.245 $X2=2.37 $Y2=0.245
cc_11 VNB N_B1_c_244_n 0.0207798f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_B1_M1007_g 0.00710979f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_B1_M1023_g 0.00669585f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB B1 0.00932786f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=2.465
cc_15 VNB N_B1_c_248_n 0.0829188f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=2.465
cc_16 VNB N_A1_c_294_n 0.0220814f $X=-0.19 $Y=-0.245 $X2=2.37 $Y2=0.245
cc_17 VNB N_A1_M1001_g 0.00718273f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A1_c_296_n 0.0164438f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A1_M1012_g 0.00662607f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB A1 0.00853535f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=2.465
cc_21 VNB N_A1_c_299_n 0.0375659f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=2.465
cc_22 VNB N_A2_c_344_n 0.0164438f $X=-0.19 $Y=-0.245 $X2=2.37 $Y2=0.245
cc_23 VNB N_A2_M1008_g 0.00687517f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A2_c_346_n 0.0220814f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A2_M1027_g 0.0075388f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB A2 0.00429511f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=2.465
cc_27 VNB N_A2_c_349_n 0.0431489f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=2.465
cc_28 VNB N_A3_M1005_g 0.00719465f $X=-0.19 $Y=-0.245 $X2=2.89 $Y2=1.835
cc_29 VNB N_A3_M1014_g 0.00740305f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A3_c_391_n 0.0220814f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A3_c_392_n 0.0209416f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=0.665
cc_32 VNB N_A3_c_393_n 0.0475032f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A3_c_394_n 0.0164438f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=1.655
cc_34 VNB A3 0.00812944f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=1.325
cc_35 VNB N_A4_c_442_n 0.0105119f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A4_c_443_n 0.00651937f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A4_M1009_g 0.0224738f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A4_M1019_g 0.0305917f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB A4 0.0377083f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A4_c_447_n 0.0426962f $X=-0.19 $Y=-0.245 $X2=1.435 $Y2=0.665
cc_41 VNB N_VPWR_c_488_n 0.322901f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_X_c_608_n 0.00144554f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_X_c_609_n 0.00660942f $X=-0.19 $Y=-0.245 $X2=1.435 $Y2=0.665
cc_44 VNB N_X_c_610_n 0.00147023f $X=-0.19 $Y=-0.245 $X2=2.38 $Y2=1.49
cc_45 VNB N_X_c_611_n 0.012488f $X=-0.19 $Y=-0.245 $X2=1.775 $Y2=1.49
cc_46 VNB X 0.0235437f $X=-0.19 $Y=-0.245 $X2=2.492 $Y2=0.42
cc_47 VNB N_VGND_c_744_n 0.0136313f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=2.465
cc_48 VNB N_VGND_c_745_n 0.0281524f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=1.325
cc_49 VNB N_VGND_c_746_n 4.81113e-19 $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=1.655
cc_50 VNB N_VGND_c_747_n 0.00760854f $X=-0.19 $Y=-0.245 $X2=1.435 $Y2=1.325
cc_51 VNB N_VGND_c_748_n 0.00587642f $X=-0.19 $Y=-0.245 $X2=1.435 $Y2=1.655
cc_52 VNB N_VGND_c_749_n 4.89148e-19 $X=-0.19 $Y=-0.245 $X2=1.865 $Y2=1.325
cc_53 VNB N_VGND_c_750_n 0.0148369f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_751_n 0.00500104f $X=-0.19 $Y=-0.245 $X2=1.865 $Y2=1.655
cc_55 VNB N_VGND_c_752_n 0.0141444f $X=-0.19 $Y=-0.245 $X2=1.865 $Y2=2.465
cc_56 VNB N_VGND_c_753_n 0.00518002f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_VGND_c_754_n 0.0130715f $X=-0.19 $Y=-0.245 $X2=0.755 $Y2=1.49
cc_58 VNB N_VGND_c_755_n 0.0880428f $X=-0.19 $Y=-0.245 $X2=2.865 $Y2=1.79
cc_59 VNB N_VGND_c_756_n 0.0153759f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_757_n 0.376953f $X=-0.19 $Y=-0.245 $X2=2.492 $Y2=0.85
cc_61 VNB N_VGND_c_758_n 0.00451663f $X=-0.19 $Y=-0.245 $X2=0.755 $Y2=1.49
cc_62 VNB N_VGND_c_759_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=1.775 $Y2=1.49
cc_63 VNB N_A_667_47#_c_849_n 0.00287018f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=1.325
cc_64 VNB N_A_667_47#_c_850_n 0.00401681f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=1.325
cc_65 VNB N_A_922_47#_c_878_n 0.00878641f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=0.665
cc_66 VNB N_A_1115_47#_c_894_n 0.00322959f $X=-0.19 $Y=-0.245 $X2=0.575
+ $Y2=1.325
cc_67 VNB N_A_1115_47#_c_895_n 0.00770748f $X=-0.19 $Y=-0.245 $X2=1.005
+ $Y2=1.325
cc_68 VNB N_A_1115_47#_c_896_n 0.0233935f $X=-0.19 $Y=-0.245 $X2=1.005 $Y2=1.655
cc_69 VPB N_A_100_23#_M1000_g 0.0224142f $X=-0.19 $Y=1.655 $X2=0.575 $Y2=2.465
cc_70 VPB N_A_100_23#_M1006_g 0.0188421f $X=-0.19 $Y=1.655 $X2=1.005 $Y2=2.465
cc_71 VPB N_A_100_23#_M1015_g 0.0188632f $X=-0.19 $Y=1.655 $X2=1.435 $Y2=2.465
cc_72 VPB N_A_100_23#_M1020_g 0.0240585f $X=-0.19 $Y=1.655 $X2=1.865 $Y2=2.465
cc_73 VPB N_A_100_23#_c_140_n 0.0036987f $X=-0.19 $Y=1.655 $X2=2.865 $Y2=1.79
cc_74 VPB N_A_100_23#_c_134_n 0.00546575f $X=-0.19 $Y=1.655 $X2=2.487 $Y2=1.49
cc_75 VPB N_A_100_23#_c_135_n 0.00700947f $X=-0.19 $Y=1.655 $X2=1.865 $Y2=1.49
cc_76 VPB N_B1_M1007_g 0.0235119f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_77 VPB N_B1_M1023_g 0.0195866f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_78 VPB N_A1_M1001_g 0.0191404f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_79 VPB N_A1_M1012_g 0.0191445f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_80 VPB N_A2_M1008_g 0.0196923f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_81 VPB N_A2_M1027_g 0.0198821f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_82 VPB N_A3_M1005_g 0.0191445f $X=-0.19 $Y=1.655 $X2=2.89 $Y2=1.835
cc_83 VPB N_A3_M1014_g 0.0191445f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_84 VPB N_A4_M1010_g 0.0169897f $X=-0.19 $Y=1.655 $X2=2.89 $Y2=1.835
cc_85 VPB N_A4_c_442_n 0.00331001f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_86 VPB N_A4_c_443_n 0.00143884f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_87 VPB N_A4_M1021_g 0.0224511f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_88 VPB N_A4_c_447_n 0.0217197f $X=-0.19 $Y=1.655 $X2=1.435 $Y2=0.665
cc_89 VPB N_VPWR_c_489_n 0.0135296f $X=-0.19 $Y=1.655 $X2=1.005 $Y2=1.655
cc_90 VPB N_VPWR_c_490_n 0.0415885f $X=-0.19 $Y=1.655 $X2=1.005 $Y2=2.465
cc_91 VPB N_VPWR_c_491_n 3.15212e-19 $X=-0.19 $Y=1.655 $X2=1.435 $Y2=1.655
cc_92 VPB N_VPWR_c_492_n 0.0199349f $X=-0.19 $Y=1.655 $X2=1.865 $Y2=0.665
cc_93 VPB N_VPWR_c_493_n 4.02668e-19 $X=-0.19 $Y=1.655 $X2=2.38 $Y2=1.49
cc_94 VPB N_VPWR_c_494_n 0.0021878f $X=-0.19 $Y=1.655 $X2=1.775 $Y2=1.49
cc_95 VPB N_VPWR_c_495_n 0.014594f $X=-0.19 $Y=1.655 $X2=2.51 $Y2=0.42
cc_96 VPB N_VPWR_c_496_n 3.13512e-19 $X=-0.19 $Y=1.655 $X2=2.865 $Y2=1.79
cc_97 VPB N_VPWR_c_497_n 3.99129e-19 $X=-0.19 $Y=1.655 $X2=3.03 $Y2=1.875
cc_98 VPB N_VPWR_c_498_n 0.0355025f $X=-0.19 $Y=1.655 $X2=2.51 $Y2=0.96
cc_99 VPB N_VPWR_c_499_n 0.00436868f $X=-0.19 $Y=1.655 $X2=2.487 $Y2=1.49
cc_100 VPB N_VPWR_c_500_n 0.0135762f $X=-0.19 $Y=1.655 $X2=2.487 $Y2=1.79
cc_101 VPB N_VPWR_c_501_n 0.00522677f $X=-0.19 $Y=1.655 $X2=0.575 $Y2=1.49
cc_102 VPB N_VPWR_c_502_n 0.0129398f $X=-0.19 $Y=1.655 $X2=1.005 $Y2=1.49
cc_103 VPB N_VPWR_c_503_n 0.0147711f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_104 VPB N_VPWR_c_504_n 0.0129398f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_105 VPB N_VPWR_c_505_n 0.0304913f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_106 VPB N_VPWR_c_488_n 0.077254f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_107 VPB N_VPWR_c_507_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_108 VPB N_VPWR_c_508_n 0.00545601f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_109 VPB N_VPWR_c_509_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_110 VPB N_VPWR_c_510_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_111 VPB N_X_c_613_n 0.00144554f $X=-0.19 $Y=1.655 $X2=0.575 $Y2=2.465
cc_112 VPB N_X_c_614_n 0.0122586f $X=-0.19 $Y=1.655 $X2=0.575 $Y2=2.465
cc_113 VPB N_X_c_615_n 0.00585698f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_114 VPB N_X_c_616_n 0.00147023f $X=-0.19 $Y=1.655 $X2=0.755 $Y2=1.49
cc_115 VPB X 0.00545686f $X=-0.19 $Y=1.655 $X2=2.492 $Y2=0.42
cc_116 VPB N_A_495_367#_c_666_n 0.00185093f $X=-0.19 $Y=1.655 $X2=1.005
+ $Y2=0.665
cc_117 VPB N_A_495_367#_c_667_n 0.00804019f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_118 VPB N_A_495_367#_c_668_n 0.00542755f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_119 VPB N_A_495_367#_c_669_n 0.00255678f $X=-0.19 $Y=1.655 $X2=1.435
+ $Y2=1.655
cc_120 VPB N_A_495_367#_c_670_n 0.00442372f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_121 VPB N_A_495_367#_c_671_n 0.00439679f $X=-0.19 $Y=1.655 $X2=0.755 $Y2=1.49
cc_122 VPB N_A_495_367#_c_672_n 0.012044f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_123 VPB N_A_495_367#_c_673_n 0.0435297f $X=-0.19 $Y=1.655 $X2=2.595 $Y2=1.79
cc_124 VPB N_A_495_367#_c_674_n 0.00178419f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_125 VPB N_A_495_367#_c_675_n 0.0066185f $X=-0.19 $Y=1.655 $X2=2.492 $Y2=0.85
cc_126 VPB N_A_495_367#_c_676_n 0.00208404f $X=-0.19 $Y=1.655 $X2=2.51 $Y2=0.96
cc_127 N_A_100_23#_M1024_g N_B1_c_243_n 0.0166514f $X=1.865 $Y=0.665 $X2=-0.19
+ $Y2=-0.245
cc_128 N_A_100_23#_c_132_n N_B1_c_243_n 0.00140738f $X=2.487 $Y=1.405 $X2=-0.19
+ $Y2=-0.245
cc_129 N_A_100_23#_c_132_n N_B1_c_244_n 0.00272908f $X=2.487 $Y=1.405 $X2=0
+ $Y2=0
cc_130 N_A_100_23#_c_133_n N_B1_c_244_n 0.022365f $X=3.89 $Y=0.85 $X2=0 $Y2=0
cc_131 N_A_100_23#_c_140_n N_B1_M1007_g 0.015675f $X=2.865 $Y=1.79 $X2=0 $Y2=0
cc_132 N_A_100_23#_c_148_p N_B1_M1007_g 0.0142118f $X=3.03 $Y=1.98 $X2=0 $Y2=0
cc_133 N_A_100_23#_c_134_n N_B1_M1007_g 0.00654326f $X=2.487 $Y=1.49 $X2=0 $Y2=0
cc_134 N_A_100_23#_c_140_n N_B1_M1023_g 0.00411143f $X=2.865 $Y=1.79 $X2=0 $Y2=0
cc_135 N_A_100_23#_c_148_p N_B1_M1023_g 0.0118885f $X=3.03 $Y=1.98 $X2=0 $Y2=0
cc_136 N_A_100_23#_c_132_n B1 0.016147f $X=2.487 $Y=1.405 $X2=0 $Y2=0
cc_137 N_A_100_23#_c_140_n B1 0.0359448f $X=2.865 $Y=1.79 $X2=0 $Y2=0
cc_138 N_A_100_23#_c_133_n B1 0.0678893f $X=3.89 $Y=0.85 $X2=0 $Y2=0
cc_139 N_A_100_23#_c_134_n B1 0.0109181f $X=2.487 $Y=1.49 $X2=0 $Y2=0
cc_140 N_A_100_23#_c_131_n N_B1_c_248_n 0.0126225f $X=2.38 $Y=1.49 $X2=0 $Y2=0
cc_141 N_A_100_23#_c_132_n N_B1_c_248_n 0.0128988f $X=2.487 $Y=1.405 $X2=0 $Y2=0
cc_142 N_A_100_23#_c_140_n N_B1_c_248_n 0.00670738f $X=2.865 $Y=1.79 $X2=0 $Y2=0
cc_143 N_A_100_23#_c_133_n N_B1_c_248_n 0.0133489f $X=3.89 $Y=0.85 $X2=0 $Y2=0
cc_144 N_A_100_23#_c_134_n N_B1_c_248_n 0.00850164f $X=2.487 $Y=1.49 $X2=0 $Y2=0
cc_145 N_A_100_23#_c_135_n N_B1_c_248_n 0.0166514f $X=1.865 $Y=1.49 $X2=0 $Y2=0
cc_146 N_A_100_23#_c_133_n N_A1_c_294_n 0.0177725f $X=3.89 $Y=0.85 $X2=-0.19
+ $Y2=-0.245
cc_147 N_A_100_23#_c_140_n N_A1_M1001_g 3.12761e-19 $X=2.865 $Y=1.79 $X2=0 $Y2=0
cc_148 N_A_100_23#_c_133_n A1 0.00626342f $X=3.89 $Y=0.85 $X2=0 $Y2=0
cc_149 N_A_100_23#_c_133_n N_A1_c_299_n 0.00317756f $X=3.89 $Y=0.85 $X2=0 $Y2=0
cc_150 N_A_100_23#_M1000_g N_VPWR_c_490_n 0.0152824f $X=0.575 $Y=2.465 $X2=0
+ $Y2=0
cc_151 N_A_100_23#_M1006_g N_VPWR_c_490_n 7.27171e-19 $X=1.005 $Y=2.465 $X2=0
+ $Y2=0
cc_152 N_A_100_23#_M1000_g N_VPWR_c_491_n 7.27171e-19 $X=0.575 $Y=2.465 $X2=0
+ $Y2=0
cc_153 N_A_100_23#_M1006_g N_VPWR_c_491_n 0.0142189f $X=1.005 $Y=2.465 $X2=0
+ $Y2=0
cc_154 N_A_100_23#_M1015_g N_VPWR_c_491_n 0.0142995f $X=1.435 $Y=2.465 $X2=0
+ $Y2=0
cc_155 N_A_100_23#_M1020_g N_VPWR_c_491_n 7.4139e-19 $X=1.865 $Y=2.465 $X2=0
+ $Y2=0
cc_156 N_A_100_23#_M1020_g N_VPWR_c_492_n 0.00767653f $X=1.865 $Y=2.465 $X2=0
+ $Y2=0
cc_157 N_A_100_23#_c_131_n N_VPWR_c_492_n 0.0187678f $X=2.38 $Y=1.49 $X2=0 $Y2=0
cc_158 N_A_100_23#_c_148_p N_VPWR_c_492_n 0.00490926f $X=3.03 $Y=1.98 $X2=0
+ $Y2=0
cc_159 N_A_100_23#_c_134_n N_VPWR_c_492_n 0.00525255f $X=2.487 $Y=1.49 $X2=0
+ $Y2=0
cc_160 N_A_100_23#_M1000_g N_VPWR_c_502_n 0.00486043f $X=0.575 $Y=2.465 $X2=0
+ $Y2=0
cc_161 N_A_100_23#_M1006_g N_VPWR_c_502_n 0.00486043f $X=1.005 $Y=2.465 $X2=0
+ $Y2=0
cc_162 N_A_100_23#_M1015_g N_VPWR_c_503_n 0.00486043f $X=1.435 $Y=2.465 $X2=0
+ $Y2=0
cc_163 N_A_100_23#_M1020_g N_VPWR_c_503_n 0.00585385f $X=1.865 $Y=2.465 $X2=0
+ $Y2=0
cc_164 N_A_100_23#_M1007_d N_VPWR_c_488_n 0.00225186f $X=2.89 $Y=1.835 $X2=0
+ $Y2=0
cc_165 N_A_100_23#_M1000_g N_VPWR_c_488_n 0.00824727f $X=0.575 $Y=2.465 $X2=0
+ $Y2=0
cc_166 N_A_100_23#_M1006_g N_VPWR_c_488_n 0.00824727f $X=1.005 $Y=2.465 $X2=0
+ $Y2=0
cc_167 N_A_100_23#_M1015_g N_VPWR_c_488_n 0.00824727f $X=1.435 $Y=2.465 $X2=0
+ $Y2=0
cc_168 N_A_100_23#_M1020_g N_VPWR_c_488_n 0.0118221f $X=1.865 $Y=2.465 $X2=0
+ $Y2=0
cc_169 N_A_100_23#_M1002_g N_X_c_608_n 0.0165646f $X=0.575 $Y=0.665 $X2=0 $Y2=0
cc_170 N_A_100_23#_c_131_n N_X_c_608_n 0.00693257f $X=2.38 $Y=1.49 $X2=0 $Y2=0
cc_171 N_A_100_23#_M1000_g N_X_c_613_n 0.0158423f $X=0.575 $Y=2.465 $X2=0 $Y2=0
cc_172 N_A_100_23#_c_131_n N_X_c_613_n 0.00693257f $X=2.38 $Y=1.49 $X2=0 $Y2=0
cc_173 N_A_100_23#_M1004_g N_X_c_609_n 0.0139493f $X=1.005 $Y=0.665 $X2=0 $Y2=0
cc_174 N_A_100_23#_M1016_g N_X_c_609_n 0.0137142f $X=1.435 $Y=0.665 $X2=0 $Y2=0
cc_175 N_A_100_23#_M1024_g N_X_c_609_n 0.00221459f $X=1.865 $Y=0.665 $X2=0 $Y2=0
cc_176 N_A_100_23#_c_131_n N_X_c_609_n 0.0620995f $X=2.38 $Y=1.49 $X2=0 $Y2=0
cc_177 N_A_100_23#_c_132_n N_X_c_609_n 0.00409365f $X=2.487 $Y=1.405 $X2=0 $Y2=0
cc_178 N_A_100_23#_c_135_n N_X_c_609_n 0.00500423f $X=1.865 $Y=1.49 $X2=0 $Y2=0
cc_179 N_A_100_23#_M1006_g N_X_c_615_n 0.013227f $X=1.005 $Y=2.465 $X2=0 $Y2=0
cc_180 N_A_100_23#_M1015_g N_X_c_615_n 0.0131144f $X=1.435 $Y=2.465 $X2=0 $Y2=0
cc_181 N_A_100_23#_M1020_g N_X_c_615_n 0.0012159f $X=1.865 $Y=2.465 $X2=0 $Y2=0
cc_182 N_A_100_23#_c_131_n N_X_c_615_n 0.0620995f $X=2.38 $Y=1.49 $X2=0 $Y2=0
cc_183 N_A_100_23#_c_134_n N_X_c_615_n 0.00223286f $X=2.487 $Y=1.49 $X2=0 $Y2=0
cc_184 N_A_100_23#_c_135_n N_X_c_615_n 0.00500423f $X=1.865 $Y=1.49 $X2=0 $Y2=0
cc_185 N_A_100_23#_c_131_n N_X_c_610_n 0.014687f $X=2.38 $Y=1.49 $X2=0 $Y2=0
cc_186 N_A_100_23#_c_135_n N_X_c_610_n 0.00255521f $X=1.865 $Y=1.49 $X2=0 $Y2=0
cc_187 N_A_100_23#_c_131_n N_X_c_616_n 0.014687f $X=2.38 $Y=1.49 $X2=0 $Y2=0
cc_188 N_A_100_23#_c_135_n N_X_c_616_n 0.00255521f $X=1.865 $Y=1.49 $X2=0 $Y2=0
cc_189 N_A_100_23#_M1002_g X 0.0209587f $X=0.575 $Y=0.665 $X2=0 $Y2=0
cc_190 N_A_100_23#_c_131_n X 0.0140636f $X=2.38 $Y=1.49 $X2=0 $Y2=0
cc_191 N_A_100_23#_c_140_n N_A_495_367#_M1007_s 9.24827e-19 $X=2.865 $Y=1.79
+ $X2=-0.19 $Y2=-0.245
cc_192 N_A_100_23#_c_134_n N_A_495_367#_M1007_s 0.00151614f $X=2.487 $Y=1.49
+ $X2=-0.19 $Y2=-0.245
cc_193 N_A_100_23#_c_140_n N_A_495_367#_c_667_n 0.00712307f $X=2.865 $Y=1.79
+ $X2=0 $Y2=0
cc_194 N_A_100_23#_c_134_n N_A_495_367#_c_667_n 0.0144736f $X=2.487 $Y=1.49
+ $X2=0 $Y2=0
cc_195 N_A_100_23#_M1007_d N_A_495_367#_c_681_n 0.00332344f $X=2.89 $Y=1.835
+ $X2=0 $Y2=0
cc_196 N_A_100_23#_c_148_p N_A_495_367#_c_681_n 0.0159805f $X=3.03 $Y=1.98 $X2=0
+ $Y2=0
cc_197 N_A_100_23#_c_140_n N_A_495_367#_c_669_n 0.00877753f $X=2.865 $Y=1.79
+ $X2=0 $Y2=0
cc_198 N_A_100_23#_c_133_n N_VGND_M1022_s 0.0055497f $X=3.89 $Y=0.85 $X2=0 $Y2=0
cc_199 N_A_100_23#_M1002_g N_VGND_c_745_n 0.0120262f $X=0.575 $Y=0.665 $X2=0
+ $Y2=0
cc_200 N_A_100_23#_M1004_g N_VGND_c_745_n 6.10117e-19 $X=1.005 $Y=0.665 $X2=0
+ $Y2=0
cc_201 N_A_100_23#_M1002_g N_VGND_c_746_n 6.10117e-19 $X=0.575 $Y=0.665 $X2=0
+ $Y2=0
cc_202 N_A_100_23#_M1004_g N_VGND_c_746_n 0.0110386f $X=1.005 $Y=0.665 $X2=0
+ $Y2=0
cc_203 N_A_100_23#_M1016_g N_VGND_c_746_n 0.0111138f $X=1.435 $Y=0.665 $X2=0
+ $Y2=0
cc_204 N_A_100_23#_M1024_g N_VGND_c_746_n 6.23351e-19 $X=1.865 $Y=0.665 $X2=0
+ $Y2=0
cc_205 N_A_100_23#_M1024_g N_VGND_c_747_n 0.00244279f $X=1.865 $Y=0.665 $X2=0
+ $Y2=0
cc_206 N_A_100_23#_c_131_n N_VGND_c_747_n 0.0146701f $X=2.38 $Y=1.49 $X2=0 $Y2=0
cc_207 N_A_100_23#_c_132_n N_VGND_c_747_n 0.00150325f $X=2.487 $Y=1.405 $X2=0
+ $Y2=0
cc_208 N_A_100_23#_c_133_n N_VGND_c_748_n 0.0218718f $X=3.89 $Y=0.85 $X2=0 $Y2=0
cc_209 N_A_100_23#_M1016_g N_VGND_c_750_n 0.00477554f $X=1.435 $Y=0.665 $X2=0
+ $Y2=0
cc_210 N_A_100_23#_M1024_g N_VGND_c_750_n 0.00575161f $X=1.865 $Y=0.665 $X2=0
+ $Y2=0
cc_211 N_A_100_23#_c_227_p N_VGND_c_752_n 0.0136943f $X=2.51 $Y=0.42 $X2=0 $Y2=0
cc_212 N_A_100_23#_c_133_n N_VGND_c_752_n 0.00228062f $X=3.89 $Y=0.85 $X2=0
+ $Y2=0
cc_213 N_A_100_23#_M1002_g N_VGND_c_754_n 0.00477554f $X=0.575 $Y=0.665 $X2=0
+ $Y2=0
cc_214 N_A_100_23#_M1004_g N_VGND_c_754_n 0.00477554f $X=1.005 $Y=0.665 $X2=0
+ $Y2=0
cc_215 N_A_100_23#_c_133_n N_VGND_c_755_n 0.00327417f $X=3.89 $Y=0.85 $X2=0
+ $Y2=0
cc_216 N_A_100_23#_M1013_d N_VGND_c_757_n 0.00276536f $X=2.37 $Y=0.245 $X2=0
+ $Y2=0
cc_217 N_A_100_23#_M1017_s N_VGND_c_757_n 0.00225186f $X=3.75 $Y=0.235 $X2=0
+ $Y2=0
cc_218 N_A_100_23#_M1002_g N_VGND_c_757_n 0.00825815f $X=0.575 $Y=0.665 $X2=0
+ $Y2=0
cc_219 N_A_100_23#_M1004_g N_VGND_c_757_n 0.00825815f $X=1.005 $Y=0.665 $X2=0
+ $Y2=0
cc_220 N_A_100_23#_M1016_g N_VGND_c_757_n 0.00825815f $X=1.435 $Y=0.665 $X2=0
+ $Y2=0
cc_221 N_A_100_23#_M1024_g N_VGND_c_757_n 0.0105607f $X=1.865 $Y=0.665 $X2=0
+ $Y2=0
cc_222 N_A_100_23#_c_227_p N_VGND_c_757_n 0.00866972f $X=2.51 $Y=0.42 $X2=0
+ $Y2=0
cc_223 N_A_100_23#_c_133_n N_VGND_c_757_n 0.0124195f $X=3.89 $Y=0.85 $X2=0 $Y2=0
cc_224 N_A_100_23#_c_133_n N_A_667_47#_M1017_d 0.00610451f $X=3.89 $Y=0.85
+ $X2=-0.19 $Y2=-0.245
cc_225 N_A_100_23#_M1017_s N_A_667_47#_c_849_n 0.00333397f $X=3.75 $Y=0.235
+ $X2=0 $Y2=0
cc_226 N_A_100_23#_c_133_n N_A_667_47#_c_849_n 0.039625f $X=3.89 $Y=0.85 $X2=0
+ $Y2=0
cc_227 N_B1_M1023_g N_A1_M1001_g 0.0207648f $X=3.245 $Y=2.465 $X2=0 $Y2=0
cc_228 B1 N_A1_M1001_g 0.00244676f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_229 B1 A1 0.0273854f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_230 B1 N_A1_c_299_n 0.0142794f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_231 N_B1_c_248_n N_A1_c_299_n 0.0207648f $X=2.86 $Y=1.36 $X2=0 $Y2=0
cc_232 N_B1_M1007_g N_VPWR_c_492_n 0.00619481f $X=2.815 $Y=2.465 $X2=0 $Y2=0
cc_233 N_B1_M1023_g N_VPWR_c_493_n 0.00109252f $X=3.245 $Y=2.465 $X2=0 $Y2=0
cc_234 N_B1_M1007_g N_VPWR_c_498_n 0.00357877f $X=2.815 $Y=2.465 $X2=0 $Y2=0
cc_235 N_B1_M1023_g N_VPWR_c_498_n 0.00357877f $X=3.245 $Y=2.465 $X2=0 $Y2=0
cc_236 N_B1_M1007_g N_VPWR_c_488_n 0.00665089f $X=2.815 $Y=2.465 $X2=0 $Y2=0
cc_237 N_B1_M1023_g N_VPWR_c_488_n 0.00537654f $X=3.245 $Y=2.465 $X2=0 $Y2=0
cc_238 N_B1_c_248_n N_A_495_367#_c_667_n 6.01138e-19 $X=2.86 $Y=1.36 $X2=0 $Y2=0
cc_239 N_B1_M1007_g N_A_495_367#_c_681_n 0.0114565f $X=2.815 $Y=2.465 $X2=0
+ $Y2=0
cc_240 N_B1_M1023_g N_A_495_367#_c_681_n 0.0115031f $X=3.245 $Y=2.465 $X2=0
+ $Y2=0
cc_241 B1 N_A_495_367#_c_668_n 0.00994467f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_242 N_B1_M1023_g N_A_495_367#_c_669_n 6.54275e-19 $X=3.245 $Y=2.465 $X2=0
+ $Y2=0
cc_243 B1 N_A_495_367#_c_669_n 0.0140497f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_244 N_B1_c_243_n N_VGND_c_747_n 0.00244313f $X=2.295 $Y=1.195 $X2=0 $Y2=0
cc_245 N_B1_c_243_n N_VGND_c_748_n 5.18675e-19 $X=2.295 $Y=1.195 $X2=0 $Y2=0
cc_246 N_B1_c_244_n N_VGND_c_748_n 0.00795518f $X=2.725 $Y=1.19 $X2=0 $Y2=0
cc_247 N_B1_c_243_n N_VGND_c_752_n 0.00575161f $X=2.295 $Y=1.195 $X2=0 $Y2=0
cc_248 N_B1_c_244_n N_VGND_c_752_n 0.00352442f $X=2.725 $Y=1.19 $X2=0 $Y2=0
cc_249 N_B1_c_243_n N_VGND_c_757_n 0.0105607f $X=2.295 $Y=1.195 $X2=0 $Y2=0
cc_250 N_B1_c_244_n N_VGND_c_757_n 0.00422979f $X=2.725 $Y=1.19 $X2=0 $Y2=0
cc_251 N_A1_c_296_n N_A2_c_344_n 0.0149293f $X=4.105 $Y=1.185 $X2=-0.19
+ $Y2=-0.245
cc_252 N_A1_M1012_g N_A2_M1008_g 0.0271327f $X=4.105 $Y=2.465 $X2=0 $Y2=0
cc_253 A1 N_A2_M1008_g 0.00428577f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_254 A1 N_A2_M1027_g 0.00173085f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_255 A1 A2 0.0241006f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_256 N_A1_c_299_n A2 2.02843e-19 $X=4.105 $Y=1.35 $X2=0 $Y2=0
cc_257 A1 N_A2_c_349_n 0.0179869f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_258 N_A1_c_299_n N_A2_c_349_n 0.0186568f $X=4.105 $Y=1.35 $X2=0 $Y2=0
cc_259 N_A1_M1001_g N_VPWR_c_493_n 0.0153918f $X=3.675 $Y=2.465 $X2=0 $Y2=0
cc_260 N_A1_M1012_g N_VPWR_c_493_n 0.0142653f $X=4.105 $Y=2.465 $X2=0 $Y2=0
cc_261 N_A1_M1012_g N_VPWR_c_494_n 7.27577e-19 $X=4.105 $Y=2.465 $X2=0 $Y2=0
cc_262 N_A1_M1001_g N_VPWR_c_498_n 0.00486043f $X=3.675 $Y=2.465 $X2=0 $Y2=0
cc_263 N_A1_M1012_g N_VPWR_c_500_n 0.00486043f $X=4.105 $Y=2.465 $X2=0 $Y2=0
cc_264 N_A1_M1001_g N_VPWR_c_488_n 0.0082726f $X=3.675 $Y=2.465 $X2=0 $Y2=0
cc_265 N_A1_M1012_g N_VPWR_c_488_n 0.0082726f $X=4.105 $Y=2.465 $X2=0 $Y2=0
cc_266 N_A1_M1001_g N_A_495_367#_c_668_n 0.0141589f $X=3.675 $Y=2.465 $X2=0
+ $Y2=0
cc_267 N_A1_M1012_g N_A_495_367#_c_668_n 0.013144f $X=4.105 $Y=2.465 $X2=0 $Y2=0
cc_268 A1 N_A_495_367#_c_668_n 0.0256027f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_269 N_A1_c_299_n N_A_495_367#_c_668_n 0.0022691f $X=4.105 $Y=1.35 $X2=0 $Y2=0
cc_270 A1 N_A_495_367#_c_670_n 0.0215987f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_271 A1 N_A_495_367#_c_674_n 0.0169627f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_272 N_A1_c_294_n N_VGND_c_748_n 0.00231444f $X=3.675 $Y=1.185 $X2=0 $Y2=0
cc_273 N_A1_c_294_n N_VGND_c_755_n 0.00357877f $X=3.675 $Y=1.185 $X2=0 $Y2=0
cc_274 N_A1_c_296_n N_VGND_c_755_n 0.00357842f $X=4.105 $Y=1.185 $X2=0 $Y2=0
cc_275 N_A1_c_294_n N_VGND_c_757_n 0.00665089f $X=3.675 $Y=1.185 $X2=0 $Y2=0
cc_276 N_A1_c_296_n N_VGND_c_757_n 0.00537652f $X=4.105 $Y=1.185 $X2=0 $Y2=0
cc_277 N_A1_c_294_n N_A_667_47#_c_849_n 0.0097922f $X=3.675 $Y=1.185 $X2=0 $Y2=0
cc_278 N_A1_c_296_n N_A_667_47#_c_849_n 0.0126605f $X=4.105 $Y=1.185 $X2=0 $Y2=0
cc_279 N_A1_c_296_n N_A_667_47#_c_856_n 7.70569e-19 $X=4.105 $Y=1.185 $X2=0
+ $Y2=0
cc_280 N_A1_c_294_n N_A_667_47#_c_857_n 8.15389e-19 $X=3.675 $Y=1.185 $X2=0
+ $Y2=0
cc_281 N_A1_c_296_n N_A_667_47#_c_857_n 0.00752504f $X=4.105 $Y=1.185 $X2=0
+ $Y2=0
cc_282 A1 N_A_667_47#_c_857_n 0.0177989f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_283 A1 N_A_667_47#_c_850_n 0.0155243f $X=4.475 $Y=1.21 $X2=0 $Y2=0
cc_284 N_A2_M1027_g N_A3_M1005_g 0.0273153f $X=5.01 $Y=2.465 $X2=0 $Y2=0
cc_285 A2 N_A3_c_393_n 0.00160792f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_286 N_A2_c_349_n N_A3_c_393_n 0.0216046f $X=5.01 $Y=1.35 $X2=0 $Y2=0
cc_287 A2 A3 0.0229306f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_288 N_A2_c_349_n A3 3.65643e-19 $X=5.01 $Y=1.35 $X2=0 $Y2=0
cc_289 N_A2_M1008_g N_VPWR_c_493_n 7.35335e-19 $X=4.535 $Y=2.465 $X2=0 $Y2=0
cc_290 N_A2_M1008_g N_VPWR_c_494_n 0.0123626f $X=4.535 $Y=2.465 $X2=0 $Y2=0
cc_291 N_A2_M1027_g N_VPWR_c_494_n 0.00168492f $X=5.01 $Y=2.465 $X2=0 $Y2=0
cc_292 N_A2_M1027_g N_VPWR_c_495_n 0.00583607f $X=5.01 $Y=2.465 $X2=0 $Y2=0
cc_293 N_A2_M1027_g N_VPWR_c_496_n 7.3736e-19 $X=5.01 $Y=2.465 $X2=0 $Y2=0
cc_294 N_A2_M1008_g N_VPWR_c_500_n 0.00564095f $X=4.535 $Y=2.465 $X2=0 $Y2=0
cc_295 N_A2_M1008_g N_VPWR_c_488_n 0.00950825f $X=4.535 $Y=2.465 $X2=0 $Y2=0
cc_296 N_A2_M1027_g N_VPWR_c_488_n 0.010626f $X=5.01 $Y=2.465 $X2=0 $Y2=0
cc_297 N_A2_M1008_g N_A_495_367#_c_670_n 0.0140089f $X=4.535 $Y=2.465 $X2=0
+ $Y2=0
cc_298 N_A2_M1027_g N_A_495_367#_c_670_n 0.0145935f $X=5.01 $Y=2.465 $X2=0 $Y2=0
cc_299 A2 N_A_495_367#_c_670_n 0.0133212f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_300 N_A2_c_349_n N_A_495_367#_c_670_n 0.00537831f $X=5.01 $Y=1.35 $X2=0 $Y2=0
cc_301 A2 N_A_495_367#_c_675_n 0.00391946f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_302 N_A2_c_349_n N_A_495_367#_c_675_n 3.41485e-19 $X=5.01 $Y=1.35 $X2=0 $Y2=0
cc_303 N_A2_c_344_n N_VGND_c_755_n 0.00562843f $X=4.535 $Y=1.185 $X2=0 $Y2=0
cc_304 N_A2_c_346_n N_VGND_c_755_n 0.00359964f $X=4.965 $Y=1.185 $X2=0 $Y2=0
cc_305 N_A2_c_344_n N_VGND_c_757_n 0.00613151f $X=4.535 $Y=1.185 $X2=0 $Y2=0
cc_306 N_A2_c_346_n N_VGND_c_757_n 0.00675254f $X=4.965 $Y=1.185 $X2=0 $Y2=0
cc_307 N_A2_c_344_n N_A_667_47#_c_850_n 0.0119264f $X=4.535 $Y=1.185 $X2=0 $Y2=0
cc_308 N_A2_c_346_n N_A_667_47#_c_850_n 0.0105736f $X=4.965 $Y=1.185 $X2=0 $Y2=0
cc_309 A2 N_A_667_47#_c_850_n 0.0194685f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_310 N_A2_c_349_n N_A_667_47#_c_850_n 0.00461157f $X=5.01 $Y=1.35 $X2=0 $Y2=0
cc_311 N_A2_c_344_n N_A_922_47#_c_878_n 0.00342256f $X=4.535 $Y=1.185 $X2=0
+ $Y2=0
cc_312 N_A2_c_346_n N_A_922_47#_c_878_n 0.0159537f $X=4.965 $Y=1.185 $X2=0 $Y2=0
cc_313 N_A3_M1014_g N_A4_c_443_n 0.0269089f $X=5.87 $Y=2.465 $X2=0 $Y2=0
cc_314 N_A3_c_392_n N_A4_c_443_n 0.014292f $X=6.27 $Y=1.26 $X2=0 $Y2=0
cc_315 N_A3_c_394_n N_A4_M1009_g 0.0110309f $X=6.345 $Y=1.185 $X2=0 $Y2=0
cc_316 N_A3_M1014_g A4 9.24756e-19 $X=5.87 $Y=2.465 $X2=0 $Y2=0
cc_317 N_A3_c_392_n A4 0.00484916f $X=6.27 $Y=1.26 $X2=0 $Y2=0
cc_318 N_A3_c_393_n A4 0.00102868f $X=5.99 $Y=1.26 $X2=0 $Y2=0
cc_319 A3 A4 0.0178645f $X=5.915 $Y=1.21 $X2=0 $Y2=0
cc_320 N_A3_c_392_n N_A4_c_447_n 0.0110309f $X=6.27 $Y=1.26 $X2=0 $Y2=0
cc_321 A3 N_A4_c_447_n 7.80859e-19 $X=5.915 $Y=1.21 $X2=0 $Y2=0
cc_322 N_A3_M1005_g N_VPWR_c_495_n 0.00486043f $X=5.44 $Y=2.465 $X2=0 $Y2=0
cc_323 N_A3_M1005_g N_VPWR_c_496_n 0.0142768f $X=5.44 $Y=2.465 $X2=0 $Y2=0
cc_324 N_A3_M1014_g N_VPWR_c_496_n 0.0142189f $X=5.87 $Y=2.465 $X2=0 $Y2=0
cc_325 N_A3_M1014_g N_VPWR_c_497_n 7.27171e-19 $X=5.87 $Y=2.465 $X2=0 $Y2=0
cc_326 N_A3_M1014_g N_VPWR_c_504_n 0.00486043f $X=5.87 $Y=2.465 $X2=0 $Y2=0
cc_327 N_A3_M1005_g N_VPWR_c_488_n 0.0082726f $X=5.44 $Y=2.465 $X2=0 $Y2=0
cc_328 N_A3_M1014_g N_VPWR_c_488_n 0.0082726f $X=5.87 $Y=2.465 $X2=0 $Y2=0
cc_329 N_A3_M1005_g N_A_495_367#_c_671_n 0.0135756f $X=5.44 $Y=2.465 $X2=0 $Y2=0
cc_330 N_A3_M1014_g N_A_495_367#_c_671_n 0.0135756f $X=5.87 $Y=2.465 $X2=0 $Y2=0
cc_331 N_A3_c_393_n N_A_495_367#_c_671_n 8.49466e-19 $X=5.99 $Y=1.26 $X2=0 $Y2=0
cc_332 A3 N_A_495_367#_c_671_n 0.0368787f $X=5.915 $Y=1.21 $X2=0 $Y2=0
cc_333 N_A3_c_392_n N_A_495_367#_c_672_n 0.00252353f $X=6.27 $Y=1.26 $X2=0 $Y2=0
cc_334 N_A3_c_392_n N_A_495_367#_c_676_n 0.00348732f $X=6.27 $Y=1.26 $X2=0 $Y2=0
cc_335 A3 N_A_495_367#_c_676_n 0.00666549f $X=5.915 $Y=1.21 $X2=0 $Y2=0
cc_336 N_A3_c_394_n N_VGND_c_749_n 0.00124765f $X=6.345 $Y=1.185 $X2=0 $Y2=0
cc_337 N_A3_c_391_n N_VGND_c_755_n 0.00359964f $X=5.915 $Y=1.185 $X2=0 $Y2=0
cc_338 N_A3_c_394_n N_VGND_c_755_n 0.00564131f $X=6.345 $Y=1.185 $X2=0 $Y2=0
cc_339 N_A3_c_391_n N_VGND_c_757_n 0.00675254f $X=5.915 $Y=1.185 $X2=0 $Y2=0
cc_340 N_A3_c_394_n N_VGND_c_757_n 0.00612225f $X=6.345 $Y=1.185 $X2=0 $Y2=0
cc_341 N_A3_c_391_n N_A_922_47#_c_878_n 0.0159537f $X=5.915 $Y=1.185 $X2=0 $Y2=0
cc_342 N_A3_c_393_n N_A_922_47#_c_878_n 0.00359757f $X=5.99 $Y=1.26 $X2=0 $Y2=0
cc_343 A3 N_A_922_47#_c_878_n 0.00506579f $X=5.915 $Y=1.21 $X2=0 $Y2=0
cc_344 N_A3_c_391_n N_A_1115_47#_c_894_n 0.0112176f $X=5.915 $Y=1.185 $X2=0
+ $Y2=0
cc_345 N_A3_c_392_n N_A_1115_47#_c_894_n 0.00363964f $X=6.27 $Y=1.26 $X2=0 $Y2=0
cc_346 N_A3_c_393_n N_A_1115_47#_c_894_n 0.00780731f $X=5.99 $Y=1.26 $X2=0 $Y2=0
cc_347 N_A3_c_394_n N_A_1115_47#_c_894_n 0.012163f $X=6.345 $Y=1.185 $X2=0 $Y2=0
cc_348 A3 N_A_1115_47#_c_894_n 0.0370601f $X=5.915 $Y=1.21 $X2=0 $Y2=0
cc_349 N_A3_c_391_n N_A_1115_47#_c_902_n 7.5319e-19 $X=5.915 $Y=1.185 $X2=0
+ $Y2=0
cc_350 N_A3_c_394_n N_A_1115_47#_c_902_n 0.00687753f $X=6.345 $Y=1.185 $X2=0
+ $Y2=0
cc_351 N_A3_c_394_n N_A_1115_47#_c_904_n 5.5611e-19 $X=6.345 $Y=1.185 $X2=0
+ $Y2=0
cc_352 N_A4_M1010_g N_VPWR_c_496_n 7.27171e-19 $X=6.3 $Y=2.465 $X2=0 $Y2=0
cc_353 N_A4_M1010_g N_VPWR_c_497_n 0.0142189f $X=6.3 $Y=2.465 $X2=0 $Y2=0
cc_354 N_A4_M1021_g N_VPWR_c_497_n 0.0161992f $X=6.73 $Y=2.465 $X2=0 $Y2=0
cc_355 N_A4_M1010_g N_VPWR_c_504_n 0.00486043f $X=6.3 $Y=2.465 $X2=0 $Y2=0
cc_356 N_A4_M1021_g N_VPWR_c_505_n 0.00486043f $X=6.73 $Y=2.465 $X2=0 $Y2=0
cc_357 N_A4_M1010_g N_VPWR_c_488_n 0.0082726f $X=6.3 $Y=2.465 $X2=0 $Y2=0
cc_358 N_A4_M1021_g N_VPWR_c_488_n 0.00954696f $X=6.73 $Y=2.465 $X2=0 $Y2=0
cc_359 N_A4_M1010_g N_A_495_367#_c_672_n 0.0134623f $X=6.3 $Y=2.465 $X2=0 $Y2=0
cc_360 N_A4_c_442_n N_A_495_367#_c_672_n 0.00219467f $X=6.655 $Y=1.62 $X2=0
+ $Y2=0
cc_361 N_A4_M1021_g N_A_495_367#_c_672_n 0.0139178f $X=6.73 $Y=2.465 $X2=0 $Y2=0
cc_362 A4 N_A_495_367#_c_672_n 0.0535151f $X=7.355 $Y=1.21 $X2=0 $Y2=0
cc_363 N_A4_c_447_n N_A_495_367#_c_672_n 0.00910745f $X=7.115 $Y=1.49 $X2=0
+ $Y2=0
cc_364 N_A4_M1009_g N_VGND_c_749_n 0.0112814f $X=6.775 $Y=0.655 $X2=0 $Y2=0
cc_365 N_A4_M1019_g N_VGND_c_749_n 0.011776f $X=7.205 $Y=0.655 $X2=0 $Y2=0
cc_366 N_A4_M1009_g N_VGND_c_755_n 0.00486043f $X=6.775 $Y=0.655 $X2=0 $Y2=0
cc_367 N_A4_M1019_g N_VGND_c_756_n 0.00486043f $X=7.205 $Y=0.655 $X2=0 $Y2=0
cc_368 N_A4_M1009_g N_VGND_c_757_n 0.0082726f $X=6.775 $Y=0.655 $X2=0 $Y2=0
cc_369 N_A4_M1019_g N_VGND_c_757_n 0.00917987f $X=7.205 $Y=0.655 $X2=0 $Y2=0
cc_370 N_A4_c_443_n N_A_1115_47#_c_894_n 5.30526e-19 $X=6.375 $Y=1.62 $X2=0
+ $Y2=0
cc_371 A4 N_A_1115_47#_c_894_n 7.09458e-19 $X=7.355 $Y=1.21 $X2=0 $Y2=0
cc_372 N_A4_M1009_g N_A_1115_47#_c_895_n 0.0122595f $X=6.775 $Y=0.655 $X2=0
+ $Y2=0
cc_373 N_A4_M1019_g N_A_1115_47#_c_895_n 0.0122595f $X=7.205 $Y=0.655 $X2=0
+ $Y2=0
cc_374 A4 N_A_1115_47#_c_895_n 0.0649944f $X=7.355 $Y=1.21 $X2=0 $Y2=0
cc_375 N_A4_c_447_n N_A_1115_47#_c_895_n 5.26104e-19 $X=7.115 $Y=1.49 $X2=0
+ $Y2=0
cc_376 N_A4_c_442_n N_A_1115_47#_c_904_n 8.07653e-19 $X=6.655 $Y=1.62 $X2=0
+ $Y2=0
cc_377 A4 N_A_1115_47#_c_904_n 0.0185905f $X=7.355 $Y=1.21 $X2=0 $Y2=0
cc_378 N_VPWR_c_488_n N_X_M1000_d 0.00536646f $X=7.44 $Y=3.33 $X2=0 $Y2=0
cc_379 N_VPWR_c_488_n N_X_M1015_d 0.0041489f $X=7.44 $Y=3.33 $X2=0 $Y2=0
cc_380 N_VPWR_M1000_s N_X_c_613_n 2.33864e-19 $X=0.235 $Y=1.835 $X2=0 $Y2=0
cc_381 N_VPWR_c_490_n N_X_c_613_n 0.00362085f $X=0.36 $Y=2.18 $X2=0 $Y2=0
cc_382 N_VPWR_M1000_s N_X_c_614_n 0.00247068f $X=0.235 $Y=1.835 $X2=0 $Y2=0
cc_383 N_VPWR_c_490_n N_X_c_614_n 0.0203341f $X=0.36 $Y=2.18 $X2=0 $Y2=0
cc_384 N_VPWR_c_502_n N_X_c_646_n 0.0124525f $X=1.055 $Y=3.33 $X2=0 $Y2=0
cc_385 N_VPWR_c_488_n N_X_c_646_n 0.00730901f $X=7.44 $Y=3.33 $X2=0 $Y2=0
cc_386 N_VPWR_M1006_s N_X_c_615_n 0.00176461f $X=1.08 $Y=1.835 $X2=0 $Y2=0
cc_387 N_VPWR_c_491_n N_X_c_615_n 0.0170777f $X=1.22 $Y=2.18 $X2=0 $Y2=0
cc_388 N_VPWR_c_492_n N_X_c_615_n 0.00166212f $X=2.08 $Y=1.98 $X2=0 $Y2=0
cc_389 N_VPWR_c_503_n N_X_c_651_n 0.0136943f $X=1.95 $Y=3.33 $X2=0 $Y2=0
cc_390 N_VPWR_c_488_n N_X_c_651_n 0.00866972f $X=7.44 $Y=3.33 $X2=0 $Y2=0
cc_391 N_VPWR_c_488_n N_A_495_367#_M1007_s 0.00215161f $X=7.44 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_392 N_VPWR_c_488_n N_A_495_367#_M1023_s 0.00376627f $X=7.44 $Y=3.33 $X2=0
+ $Y2=0
cc_393 N_VPWR_c_488_n N_A_495_367#_M1012_d 0.00536646f $X=7.44 $Y=3.33 $X2=0
+ $Y2=0
cc_394 N_VPWR_c_488_n N_A_495_367#_M1027_s 0.00467071f $X=7.44 $Y=3.33 $X2=0
+ $Y2=0
cc_395 N_VPWR_c_488_n N_A_495_367#_M1014_d 0.00536646f $X=7.44 $Y=3.33 $X2=0
+ $Y2=0
cc_396 N_VPWR_c_488_n N_A_495_367#_M1021_d 0.00371702f $X=7.44 $Y=3.33 $X2=0
+ $Y2=0
cc_397 N_VPWR_c_492_n N_A_495_367#_c_666_n 0.0132687f $X=2.08 $Y=1.98 $X2=0
+ $Y2=0
cc_398 N_VPWR_c_498_n N_A_495_367#_c_666_n 0.0179183f $X=3.725 $Y=3.33 $X2=0
+ $Y2=0
cc_399 N_VPWR_c_488_n N_A_495_367#_c_666_n 0.0101082f $X=7.44 $Y=3.33 $X2=0
+ $Y2=0
cc_400 N_VPWR_c_492_n N_A_495_367#_c_667_n 0.0620204f $X=2.08 $Y=1.98 $X2=0
+ $Y2=0
cc_401 N_VPWR_c_498_n N_A_495_367#_c_681_n 0.0361172f $X=3.725 $Y=3.33 $X2=0
+ $Y2=0
cc_402 N_VPWR_c_488_n N_A_495_367#_c_681_n 0.023676f $X=7.44 $Y=3.33 $X2=0 $Y2=0
cc_403 N_VPWR_c_498_n N_A_495_367#_c_726_n 0.0125234f $X=3.725 $Y=3.33 $X2=0
+ $Y2=0
cc_404 N_VPWR_c_488_n N_A_495_367#_c_726_n 0.00738676f $X=7.44 $Y=3.33 $X2=0
+ $Y2=0
cc_405 N_VPWR_M1001_s N_A_495_367#_c_668_n 0.00176461f $X=3.75 $Y=1.835 $X2=0
+ $Y2=0
cc_406 N_VPWR_c_493_n N_A_495_367#_c_668_n 0.0170777f $X=3.89 $Y=2.18 $X2=0
+ $Y2=0
cc_407 N_VPWR_c_500_n N_A_495_367#_c_730_n 0.0124525f $X=4.605 $Y=3.33 $X2=0
+ $Y2=0
cc_408 N_VPWR_c_488_n N_A_495_367#_c_730_n 0.00730901f $X=7.44 $Y=3.33 $X2=0
+ $Y2=0
cc_409 N_VPWR_M1008_d N_A_495_367#_c_670_n 0.00224297f $X=4.61 $Y=1.835 $X2=0
+ $Y2=0
cc_410 N_VPWR_c_494_n N_A_495_367#_c_670_n 0.0174292f $X=4.77 $Y=2.18 $X2=0
+ $Y2=0
cc_411 N_VPWR_c_495_n N_A_495_367#_c_734_n 0.0131621f $X=5.49 $Y=3.33 $X2=0
+ $Y2=0
cc_412 N_VPWR_c_488_n N_A_495_367#_c_734_n 0.00808656f $X=7.44 $Y=3.33 $X2=0
+ $Y2=0
cc_413 N_VPWR_M1005_s N_A_495_367#_c_671_n 0.00176461f $X=5.515 $Y=1.835 $X2=0
+ $Y2=0
cc_414 N_VPWR_c_496_n N_A_495_367#_c_671_n 0.0170777f $X=5.655 $Y=2.18 $X2=0
+ $Y2=0
cc_415 N_VPWR_c_504_n N_A_495_367#_c_738_n 0.0124525f $X=6.35 $Y=3.33 $X2=0
+ $Y2=0
cc_416 N_VPWR_c_488_n N_A_495_367#_c_738_n 0.00730901f $X=7.44 $Y=3.33 $X2=0
+ $Y2=0
cc_417 N_VPWR_M1010_s N_A_495_367#_c_672_n 0.00176461f $X=6.375 $Y=1.835 $X2=0
+ $Y2=0
cc_418 N_VPWR_c_497_n N_A_495_367#_c_672_n 0.0170777f $X=6.515 $Y=2.18 $X2=0
+ $Y2=0
cc_419 N_VPWR_c_505_n N_A_495_367#_c_673_n 0.0178111f $X=7.44 $Y=3.33 $X2=0
+ $Y2=0
cc_420 N_VPWR_c_488_n N_A_495_367#_c_673_n 0.0100304f $X=7.44 $Y=3.33 $X2=0
+ $Y2=0
cc_421 N_X_c_608_n N_VGND_M1002_d 2.33864e-19 $X=0.695 $Y=1.14 $X2=-0.19
+ $Y2=-0.245
cc_422 N_X_c_611_n N_VGND_M1002_d 0.0021884f $X=0.26 $Y=1.225 $X2=-0.19
+ $Y2=-0.245
cc_423 N_X_c_609_n N_VGND_M1004_d 0.00176461f $X=1.555 $Y=1.14 $X2=0 $Y2=0
cc_424 N_X_c_608_n N_VGND_c_745_n 0.00362085f $X=0.695 $Y=1.14 $X2=0 $Y2=0
cc_425 N_X_c_611_n N_VGND_c_745_n 0.0203341f $X=0.26 $Y=1.225 $X2=0 $Y2=0
cc_426 N_X_c_609_n N_VGND_c_746_n 0.0170777f $X=1.555 $Y=1.14 $X2=0 $Y2=0
cc_427 N_X_c_609_n N_VGND_c_747_n 0.0016514f $X=1.555 $Y=1.14 $X2=0 $Y2=0
cc_428 N_X_c_660_p N_VGND_c_750_n 0.0136943f $X=1.65 $Y=0.42 $X2=0 $Y2=0
cc_429 N_X_c_661_p N_VGND_c_754_n 0.0124525f $X=0.79 $Y=0.42 $X2=0 $Y2=0
cc_430 N_X_M1002_s N_VGND_c_757_n 0.00536646f $X=0.65 $Y=0.245 $X2=0 $Y2=0
cc_431 N_X_M1016_s N_VGND_c_757_n 0.0041489f $X=1.51 $Y=0.245 $X2=0 $Y2=0
cc_432 N_X_c_661_p N_VGND_c_757_n 0.00730901f $X=0.79 $Y=0.42 $X2=0 $Y2=0
cc_433 N_X_c_660_p N_VGND_c_757_n 0.00866972f $X=1.65 $Y=0.42 $X2=0 $Y2=0
cc_434 N_VGND_c_757_n N_A_667_47#_M1017_d 0.00215176f $X=7.44 $Y=0 $X2=-0.19
+ $Y2=-0.245
cc_435 N_VGND_c_757_n N_A_667_47#_M1025_d 0.00242289f $X=7.44 $Y=0 $X2=0 $Y2=0
cc_436 N_VGND_c_757_n N_A_667_47#_M1018_d 0.00216245f $X=7.44 $Y=0 $X2=0 $Y2=0
cc_437 N_VGND_c_748_n N_A_667_47#_c_849_n 0.0202776f $X=2.94 $Y=0.41 $X2=0 $Y2=0
cc_438 N_VGND_c_755_n N_A_667_47#_c_849_n 0.0503094f $X=6.825 $Y=0 $X2=0 $Y2=0
cc_439 N_VGND_c_757_n N_A_667_47#_c_849_n 0.0312779f $X=7.44 $Y=0 $X2=0 $Y2=0
cc_440 N_VGND_c_755_n N_A_667_47#_c_856_n 0.0161465f $X=6.825 $Y=0 $X2=0 $Y2=0
cc_441 N_VGND_c_757_n N_A_667_47#_c_856_n 0.0103094f $X=7.44 $Y=0 $X2=0 $Y2=0
cc_442 N_VGND_c_757_n N_A_667_47#_c_850_n 0.00663243f $X=7.44 $Y=0 $X2=0 $Y2=0
cc_443 N_VGND_c_757_n N_A_922_47#_M1003_s 0.00223855f $X=7.44 $Y=0 $X2=-0.19
+ $Y2=-0.245
cc_444 N_VGND_c_757_n N_A_922_47#_M1011_s 0.00242549f $X=7.44 $Y=0 $X2=0 $Y2=0
cc_445 N_VGND_c_755_n N_A_922_47#_c_878_n 0.0929611f $X=6.825 $Y=0 $X2=0 $Y2=0
cc_446 N_VGND_c_757_n N_A_922_47#_c_878_n 0.060579f $X=7.44 $Y=0 $X2=0 $Y2=0
cc_447 N_VGND_c_757_n N_A_1115_47#_M1011_d 0.00216245f $X=7.44 $Y=0 $X2=-0.19
+ $Y2=-0.245
cc_448 N_VGND_c_757_n N_A_1115_47#_M1026_d 0.00380103f $X=7.44 $Y=0 $X2=0 $Y2=0
cc_449 N_VGND_c_757_n N_A_1115_47#_M1019_d 0.00371702f $X=7.44 $Y=0 $X2=0 $Y2=0
cc_450 N_VGND_c_757_n N_A_1115_47#_c_894_n 0.00666184f $X=7.44 $Y=0 $X2=0 $Y2=0
cc_451 N_VGND_c_755_n N_A_1115_47#_c_902_n 0.0150063f $X=6.825 $Y=0 $X2=0 $Y2=0
cc_452 N_VGND_c_757_n N_A_1115_47#_c_902_n 0.00950443f $X=7.44 $Y=0 $X2=0 $Y2=0
cc_453 N_VGND_M1009_s N_A_1115_47#_c_895_n 0.00334223f $X=6.85 $Y=0.235 $X2=0
+ $Y2=0
cc_454 N_VGND_c_749_n N_A_1115_47#_c_895_n 0.0170777f $X=6.99 $Y=0.535 $X2=0
+ $Y2=0
cc_455 N_VGND_c_756_n N_A_1115_47#_c_896_n 0.0178111f $X=7.44 $Y=0 $X2=0 $Y2=0
cc_456 N_VGND_c_757_n N_A_1115_47#_c_896_n 0.0100304f $X=7.44 $Y=0 $X2=0 $Y2=0
cc_457 N_A_667_47#_c_850_n N_A_922_47#_M1003_s 0.00466546f $X=5.18 $Y=0.88
+ $X2=-0.19 $Y2=-0.245
cc_458 N_A_667_47#_M1018_d N_A_922_47#_c_878_n 0.00578783f $X=5.04 $Y=0.235
+ $X2=0 $Y2=0
cc_459 N_A_667_47#_c_850_n N_A_922_47#_c_878_n 0.043225f $X=5.18 $Y=0.88 $X2=0
+ $Y2=0
cc_460 N_A_667_47#_c_850_n N_A_1115_47#_c_894_n 0.0214676f $X=5.18 $Y=0.88 $X2=0
+ $Y2=0
cc_461 N_A_922_47#_c_878_n N_A_1115_47#_M1011_d 0.00564433f $X=6.13 $Y=0.43
+ $X2=-0.19 $Y2=-0.245
cc_462 N_A_922_47#_M1011_s N_A_1115_47#_c_894_n 0.00464204f $X=5.99 $Y=0.235
+ $X2=0 $Y2=0
cc_463 N_A_922_47#_c_878_n N_A_1115_47#_c_894_n 0.042484f $X=6.13 $Y=0.43 $X2=0
+ $Y2=0
