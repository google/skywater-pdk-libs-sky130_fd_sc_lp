* File: sky130_fd_sc_lp__xnor2_2.pxi.spice
* Created: Wed Sep  2 10:40:09 2020
* 
x_PM_SKY130_FD_SC_LP__XNOR2_2%A N_A_M1007_g N_A_M1014_g N_A_M1019_g N_A_M1011_g
+ N_A_M1000_g N_A_M1010_g N_A_M1008_g N_A_M1009_g N_A_c_117_n N_A_c_118_n
+ N_A_c_134_p N_A_c_119_n N_A_c_120_n N_A_c_162_p A A N_A_c_121_n N_A_c_122_n
+ N_A_c_123_n PM_SKY130_FD_SC_LP__XNOR2_2%A
x_PM_SKY130_FD_SC_LP__XNOR2_2%B N_B_M1002_g N_B_M1005_g N_B_M1018_g N_B_M1015_g
+ N_B_M1016_g N_B_M1001_g N_B_M1017_g N_B_M1006_g N_B_c_259_n N_B_c_260_n
+ N_B_c_261_n N_B_c_262_n N_B_c_263_n N_B_c_274_n N_B_c_275_n B B N_B_c_264_n
+ PM_SKY130_FD_SC_LP__XNOR2_2%B
x_PM_SKY130_FD_SC_LP__XNOR2_2%A_162_367# N_A_162_367#_M1002_s
+ N_A_162_367#_M1014_s N_A_162_367#_M1005_d N_A_162_367#_M1003_g
+ N_A_162_367#_M1004_g N_A_162_367#_M1012_g N_A_162_367#_M1013_g
+ N_A_162_367#_c_399_n N_A_162_367#_c_483_p N_A_162_367#_c_400_n
+ N_A_162_367#_c_401_n N_A_162_367#_c_426_n N_A_162_367#_c_430_n
+ N_A_162_367#_c_523_p N_A_162_367#_c_431_n N_A_162_367#_c_434_n
+ N_A_162_367#_c_435_n N_A_162_367#_c_407_n N_A_162_367#_c_408_n
+ N_A_162_367#_c_409_n N_A_162_367#_c_468_n N_A_162_367#_c_402_n
+ N_A_162_367#_c_439_n N_A_162_367#_c_410_n N_A_162_367#_c_403_n
+ PM_SKY130_FD_SC_LP__XNOR2_2%A_162_367#
x_PM_SKY130_FD_SC_LP__XNOR2_2%VPWR N_VPWR_M1014_d N_VPWR_M1019_d N_VPWR_M1015_s
+ N_VPWR_M1010_d N_VPWR_M1004_s N_VPWR_c_545_n N_VPWR_c_546_n N_VPWR_c_547_n
+ N_VPWR_c_548_n N_VPWR_c_549_n N_VPWR_c_550_n N_VPWR_c_551_n N_VPWR_c_552_n
+ N_VPWR_c_553_n N_VPWR_c_554_n N_VPWR_c_555_n N_VPWR_c_556_n N_VPWR_c_557_n
+ N_VPWR_c_558_n VPWR N_VPWR_c_559_n N_VPWR_c_560_n N_VPWR_c_544_n
+ N_VPWR_c_562_n VPWR PM_SKY130_FD_SC_LP__XNOR2_2%VPWR
x_PM_SKY130_FD_SC_LP__XNOR2_2%A_545_367# N_A_545_367#_M1000_s
+ N_A_545_367#_M1001_s N_A_545_367#_c_639_n N_A_545_367#_c_640_n
+ N_A_545_367#_c_641_n N_A_545_367#_c_642_n N_A_545_367#_c_645_n
+ N_A_545_367#_c_650_n PM_SKY130_FD_SC_LP__XNOR2_2%A_545_367#
x_PM_SKY130_FD_SC_LP__XNOR2_2%Y N_Y_M1003_d N_Y_M1001_d N_Y_M1006_d N_Y_M1013_d
+ N_Y_c_692_n N_Y_c_722_n N_Y_c_686_n N_Y_c_687_n N_Y_c_682_n N_Y_c_683_n
+ N_Y_c_688_n N_Y_c_689_n Y Y Y Y Y Y N_Y_c_714_n N_Y_c_684_n Y
+ PM_SKY130_FD_SC_LP__XNOR2_2%Y
x_PM_SKY130_FD_SC_LP__XNOR2_2%A_27_47# N_A_27_47#_M1007_s N_A_27_47#_M1011_s
+ N_A_27_47#_M1018_d N_A_27_47#_c_743_n N_A_27_47#_c_748_n N_A_27_47#_c_744_n
+ N_A_27_47#_c_752_n N_A_27_47#_c_754_n N_A_27_47#_c_756_n N_A_27_47#_c_745_n
+ PM_SKY130_FD_SC_LP__XNOR2_2%A_27_47#
x_PM_SKY130_FD_SC_LP__XNOR2_2%VGND N_VGND_M1007_d N_VGND_M1008_d N_VGND_M1016_s
+ N_VGND_c_795_n N_VGND_c_796_n N_VGND_c_797_n N_VGND_c_798_n N_VGND_c_799_n
+ N_VGND_c_800_n VGND N_VGND_c_801_n N_VGND_c_802_n N_VGND_c_803_n
+ N_VGND_c_804_n N_VGND_c_805_n VGND PM_SKY130_FD_SC_LP__XNOR2_2%VGND
x_PM_SKY130_FD_SC_LP__XNOR2_2%A_555_65# N_A_555_65#_M1008_s N_A_555_65#_M1009_s
+ N_A_555_65#_M1017_d N_A_555_65#_M1012_s N_A_555_65#_c_875_n
+ N_A_555_65#_c_876_n N_A_555_65#_c_877_n N_A_555_65#_c_878_n
+ N_A_555_65#_c_879_n N_A_555_65#_c_880_n N_A_555_65#_c_881_n
+ N_A_555_65#_c_882_n N_A_555_65#_c_883_n PM_SKY130_FD_SC_LP__XNOR2_2%A_555_65#
cc_1 VNB N_A_M1007_g 0.038175f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.655
cc_2 VNB N_A_M1011_g 0.0267013f $X=-0.19 $Y=-0.245 $X2=1.205 $Y2=0.655
cc_3 VNB N_A_M1008_g 0.0220108f $X=-0.19 $Y=-0.245 $X2=3.115 $Y2=0.745
cc_4 VNB N_A_M1009_g 0.0185546f $X=-0.19 $Y=-0.245 $X2=3.545 $Y2=0.745
cc_5 VNB N_A_c_117_n 0.00147624f $X=-0.19 $Y=-0.245 $X2=1.74 $Y2=1.425
cc_6 VNB N_A_c_118_n 0.016072f $X=-0.19 $Y=-0.245 $X2=2.465 $Y2=1.09
cc_7 VNB N_A_c_119_n 0.00288164f $X=-0.19 $Y=-0.245 $X2=2.55 $Y2=1.405
cc_8 VNB N_A_c_120_n 0.00106771f $X=-0.19 $Y=-0.245 $X2=2.635 $Y2=1.49
cc_9 VNB N_A_c_121_n 0.0712165f $X=-0.19 $Y=-0.245 $X2=1.185 $Y2=1.51
cc_10 VNB N_A_c_122_n 0.0712695f $X=-0.19 $Y=-0.245 $X2=3.545 $Y2=1.49
cc_11 VNB N_A_c_123_n 0.00249538f $X=-0.19 $Y=-0.245 $X2=1.655 $Y2=1.587
cc_12 VNB N_B_M1002_g 0.0236383f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.655
cc_13 VNB N_B_M1018_g 0.0287085f $X=-0.19 $Y=-0.245 $X2=1.165 $Y2=2.465
cc_14 VNB N_B_M1016_g 0.0231904f $X=-0.19 $Y=-0.245 $X2=2.65 $Y2=2.465
cc_15 VNB N_B_M1017_g 0.0231791f $X=-0.19 $Y=-0.245 $X2=3.115 $Y2=0.745
cc_16 VNB N_B_c_259_n 0.0124512f $X=-0.19 $Y=-0.245 $X2=1.74 $Y2=1.175
cc_17 VNB N_B_c_260_n 0.017526f $X=-0.19 $Y=-0.245 $X2=1.74 $Y2=1.425
cc_18 VNB N_B_c_261_n 0.0315881f $X=-0.19 $Y=-0.245 $X2=2.55 $Y2=1.175
cc_19 VNB N_B_c_262_n 0.00360381f $X=-0.19 $Y=-0.245 $X2=2.97 $Y2=1.49
cc_20 VNB N_B_c_263_n 0.035508f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_B_c_264_n 0.00194988f $X=-0.19 $Y=-0.245 $X2=1.185 $Y2=1.51
cc_22 VNB N_A_162_367#_M1003_g 0.0198045f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_162_367#_M1012_g 0.0230444f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_162_367#_c_399_n 0.00196408f $X=-0.19 $Y=-0.245 $X2=3.115
+ $Y2=0.745
cc_25 VNB N_A_162_367#_c_400_n 0.00868012f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_162_367#_c_401_n 0.00235142f $X=-0.19 $Y=-0.245 $X2=1.74 $Y2=1.175
cc_27 VNB N_A_162_367#_c_402_n 0.00536134f $X=-0.19 $Y=-0.245 $X2=1.185 $Y2=1.51
cc_28 VNB N_A_162_367#_c_403_n 0.0371913f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VPWR_c_544_n 0.263193f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_Y_c_682_n 0.00112945f $X=-0.19 $Y=-0.245 $X2=3.115 $Y2=1.325
cc_31 VNB N_Y_c_683_n 0.00228776f $X=-0.19 $Y=-0.245 $X2=3.115 $Y2=0.745
cc_32 VNB N_Y_c_684_n 0.00845287f $X=-0.19 $Y=-0.245 $X2=1.205 $Y2=1.51
cc_33 VNB Y 0.0219127f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_27_47#_c_743_n 0.0187593f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_27_47#_c_744_n 0.0270273f $X=-0.19 $Y=-0.245 $X2=1.205 $Y2=0.655
cc_36 VNB N_A_27_47#_c_745_n 0.00669919f $X=-0.19 $Y=-0.245 $X2=3.115 $Y2=1.325
cc_37 VNB N_VGND_c_795_n 0.00496753f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_796_n 0.00228974f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_797_n 0.0142738f $X=-0.19 $Y=-0.245 $X2=2.65 $Y2=2.465
cc_40 VNB N_VGND_c_798_n 0.00539181f $X=-0.19 $Y=-0.245 $X2=3.08 $Y2=2.465
cc_41 VNB N_VGND_c_799_n 0.0574593f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_800_n 0.00549308f $X=-0.19 $Y=-0.245 $X2=3.115 $Y2=1.325
cc_43 VNB N_VGND_c_801_n 0.0170187f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_802_n 0.0365291f $X=-0.19 $Y=-0.245 $X2=1.595 $Y2=1.58
cc_45 VNB N_VGND_c_803_n 0.337125f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_804_n 0.00420141f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.345
cc_47 VNB N_VGND_c_805_n 0.0135569f $X=-0.19 $Y=-0.245 $X2=1.185 $Y2=1.51
cc_48 VNB N_A_555_65#_c_875_n 0.00201769f $X=-0.19 $Y=-0.245 $X2=1.205 $Y2=0.655
cc_49 VNB N_A_555_65#_c_876_n 0.00396512f $X=-0.19 $Y=-0.245 $X2=2.65 $Y2=1.655
cc_50 VNB N_A_555_65#_c_877_n 0.00177925f $X=-0.19 $Y=-0.245 $X2=2.65 $Y2=2.465
cc_51 VNB N_A_555_65#_c_878_n 0.00191707f $X=-0.19 $Y=-0.245 $X2=3.08 $Y2=1.655
cc_52 VNB N_A_555_65#_c_879_n 0.00922926f $X=-0.19 $Y=-0.245 $X2=3.08 $Y2=2.465
cc_53 VNB N_A_555_65#_c_880_n 0.0125819f $X=-0.19 $Y=-0.245 $X2=3.545 $Y2=1.325
cc_54 VNB N_A_555_65#_c_881_n 0.00190976f $X=-0.19 $Y=-0.245 $X2=3.545 $Y2=0.745
cc_55 VNB N_A_555_65#_c_882_n 0.0185206f $X=-0.19 $Y=-0.245 $X2=1.74 $Y2=1.175
cc_56 VNB N_A_555_65#_c_883_n 0.00169939f $X=-0.19 $Y=-0.245 $X2=2.465 $Y2=1.09
cc_57 VPB N_A_M1014_g 0.0249125f $X=-0.19 $Y=1.655 $X2=0.735 $Y2=2.465
cc_58 VPB N_A_M1019_g 0.0185251f $X=-0.19 $Y=1.655 $X2=1.165 $Y2=2.465
cc_59 VPB N_A_M1000_g 0.020677f $X=-0.19 $Y=1.655 $X2=2.65 $Y2=2.465
cc_60 VPB N_A_M1010_g 0.0233882f $X=-0.19 $Y=1.655 $X2=3.08 $Y2=2.465
cc_61 VPB N_A_c_117_n 0.00162782f $X=-0.19 $Y=1.655 $X2=1.74 $Y2=1.425
cc_62 VPB N_A_c_121_n 0.00844488f $X=-0.19 $Y=1.655 $X2=1.185 $Y2=1.51
cc_63 VPB N_A_c_122_n 0.0178922f $X=-0.19 $Y=1.655 $X2=3.545 $Y2=1.49
cc_64 VPB N_A_c_123_n 0.00408535f $X=-0.19 $Y=1.655 $X2=1.655 $Y2=1.587
cc_65 VPB N_B_M1005_g 0.0185303f $X=-0.19 $Y=1.655 $X2=0.735 $Y2=2.465
cc_66 VPB N_B_M1015_g 0.0196343f $X=-0.19 $Y=1.655 $X2=1.205 $Y2=0.655
cc_67 VPB N_B_M1001_g 0.0247157f $X=-0.19 $Y=1.655 $X2=3.08 $Y2=2.465
cc_68 VPB N_B_M1006_g 0.0183698f $X=-0.19 $Y=1.655 $X2=3.545 $Y2=0.745
cc_69 VPB N_B_c_259_n 0.0071881f $X=-0.19 $Y=1.655 $X2=1.74 $Y2=1.175
cc_70 VPB N_B_c_260_n 0.0106545f $X=-0.19 $Y=1.655 $X2=1.74 $Y2=1.425
cc_71 VPB N_B_c_261_n 0.00428687f $X=-0.19 $Y=1.655 $X2=2.55 $Y2=1.175
cc_72 VPB N_B_c_262_n 9.65867e-19 $X=-0.19 $Y=1.655 $X2=2.97 $Y2=1.49
cc_73 VPB N_B_c_263_n 0.00787825f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_74 VPB N_B_c_274_n 0.00575273f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_75 VPB N_B_c_275_n 0.00811955f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_76 VPB N_B_c_264_n 0.00904355f $X=-0.19 $Y=1.655 $X2=1.185 $Y2=1.51
cc_77 VPB N_A_162_367#_M1004_g 0.0182105f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_78 VPB N_A_162_367#_M1013_g 0.0219065f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_79 VPB N_A_162_367#_c_399_n 0.00131982f $X=-0.19 $Y=1.655 $X2=3.115 $Y2=0.745
cc_80 VPB N_A_162_367#_c_407_n 0.00548555f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_81 VPB N_A_162_367#_c_408_n 0.0125315f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_82 VPB N_A_162_367#_c_409_n 0.0012563f $X=-0.19 $Y=1.655 $X2=1.165 $Y2=1.51
cc_83 VPB N_A_162_367#_c_410_n 0.0116158f $X=-0.19 $Y=1.655 $X2=1.655 $Y2=1.587
cc_84 VPB N_A_162_367#_c_403_n 0.00645697f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_85 VPB N_VPWR_c_545_n 0.00640596f $X=-0.19 $Y=1.655 $X2=2.65 $Y2=2.465
cc_86 VPB N_VPWR_c_546_n 0.00509083f $X=-0.19 $Y=1.655 $X2=3.08 $Y2=2.465
cc_87 VPB N_VPWR_c_547_n 3.35682e-19 $X=-0.19 $Y=1.655 $X2=3.115 $Y2=0.745
cc_88 VPB N_VPWR_c_548_n 0.00450326f $X=-0.19 $Y=1.655 $X2=3.545 $Y2=0.745
cc_89 VPB N_VPWR_c_549_n 0.00860907f $X=-0.19 $Y=1.655 $X2=1.74 $Y2=1.425
cc_90 VPB N_VPWR_c_550_n 4.89148e-19 $X=-0.19 $Y=1.655 $X2=2.55 $Y2=1.405
cc_91 VPB N_VPWR_c_551_n 0.0116899f $X=-0.19 $Y=1.655 $X2=1.115 $Y2=1.58
cc_92 VPB N_VPWR_c_552_n 0.0066101f $X=-0.19 $Y=1.655 $X2=1.595 $Y2=1.58
cc_93 VPB N_VPWR_c_553_n 0.0153314f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_94 VPB N_VPWR_c_554_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_95 VPB N_VPWR_c_555_n 0.0162887f $X=-0.19 $Y=1.655 $X2=0.735 $Y2=1.51
cc_96 VPB N_VPWR_c_556_n 0.0063201f $X=-0.19 $Y=1.655 $X2=1.165 $Y2=1.51
cc_97 VPB N_VPWR_c_557_n 0.0174662f $X=-0.19 $Y=1.655 $X2=1.185 $Y2=1.51
cc_98 VPB N_VPWR_c_558_n 0.00497021f $X=-0.19 $Y=1.655 $X2=1.185 $Y2=1.51
cc_99 VPB N_VPWR_c_559_n 0.046467f $X=-0.19 $Y=1.655 $X2=1.74 $Y2=1.587
cc_100 VPB N_VPWR_c_560_n 0.0152818f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_101 VPB N_VPWR_c_544_n 0.0583247f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_102 VPB N_VPWR_c_562_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_103 VPB N_A_545_367#_c_639_n 0.0104889f $X=-0.19 $Y=1.655 $X2=1.165 $Y2=1.675
cc_104 VPB N_A_545_367#_c_640_n 0.00808185f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_105 VPB N_A_545_367#_c_641_n 0.0124186f $X=-0.19 $Y=1.655 $X2=1.205 $Y2=1.345
cc_106 VPB N_A_545_367#_c_642_n 0.00430895f $X=-0.19 $Y=1.655 $X2=1.205
+ $Y2=0.655
cc_107 VPB N_Y_c_686_n 0.00307864f $X=-0.19 $Y=1.655 $X2=3.08 $Y2=2.465
cc_108 VPB N_Y_c_687_n 0.0021323f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_109 VPB N_Y_c_688_n 0.00964961f $X=-0.19 $Y=1.655 $X2=3.115 $Y2=0.745
cc_110 VPB N_Y_c_689_n 0.00742669f $X=-0.19 $Y=1.655 $X2=1.825 $Y2=1.09
cc_111 VPB Y 0.0434569f $X=-0.19 $Y=1.655 $X2=2.97 $Y2=1.49
cc_112 VPB Y 0.00605831f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_113 N_A_M1011_g N_B_M1002_g 0.03765f $X=1.205 $Y=0.655 $X2=0 $Y2=0
cc_114 N_A_c_117_n N_B_M1002_g 0.00385091f $X=1.74 $Y=1.425 $X2=0 $Y2=0
cc_115 N_A_c_134_p N_B_M1002_g 0.00495301f $X=1.825 $Y=1.09 $X2=0 $Y2=0
cc_116 N_A_M1019_g N_B_M1005_g 0.0320168f $X=1.165 $Y=2.465 $X2=0 $Y2=0
cc_117 N_A_c_117_n N_B_M1005_g 0.00166283f $X=1.74 $Y=1.425 $X2=0 $Y2=0
cc_118 N_A_c_123_n N_B_M1005_g 0.00286284f $X=1.655 $Y=1.587 $X2=0 $Y2=0
cc_119 N_A_c_117_n N_B_M1018_g 0.00174241f $X=1.74 $Y=1.425 $X2=0 $Y2=0
cc_120 N_A_c_118_n N_B_M1018_g 0.0139962f $X=2.465 $Y=1.09 $X2=0 $Y2=0
cc_121 N_A_c_119_n N_B_M1018_g 0.00300334f $X=2.55 $Y=1.405 $X2=0 $Y2=0
cc_122 N_A_c_122_n N_B_M1018_g 7.69394e-19 $X=3.545 $Y=1.49 $X2=0 $Y2=0
cc_123 N_A_M1000_g N_B_M1015_g 0.0360003f $X=2.65 $Y=2.465 $X2=0 $Y2=0
cc_124 N_A_c_117_n N_B_M1015_g 6.24055e-19 $X=1.74 $Y=1.425 $X2=0 $Y2=0
cc_125 N_A_M1009_g N_B_M1016_g 0.020027f $X=3.545 $Y=0.745 $X2=0 $Y2=0
cc_126 N_A_c_122_n N_B_c_259_n 0.0213871f $X=3.545 $Y=1.49 $X2=0 $Y2=0
cc_127 N_A_M1000_g N_B_c_262_n 0.00174942f $X=2.65 $Y=2.465 $X2=0 $Y2=0
cc_128 N_A_c_117_n N_B_c_262_n 0.0296132f $X=1.74 $Y=1.425 $X2=0 $Y2=0
cc_129 N_A_c_118_n N_B_c_262_n 0.02205f $X=2.465 $Y=1.09 $X2=0 $Y2=0
cc_130 N_A_c_119_n N_B_c_262_n 0.00428208f $X=2.55 $Y=1.405 $X2=0 $Y2=0
cc_131 N_A_c_120_n N_B_c_262_n 0.0135772f $X=2.635 $Y=1.49 $X2=0 $Y2=0
cc_132 N_A_c_122_n N_B_c_262_n 0.00276733f $X=3.545 $Y=1.49 $X2=0 $Y2=0
cc_133 N_A_M1000_g N_B_c_263_n 6.86117e-19 $X=2.65 $Y=2.465 $X2=0 $Y2=0
cc_134 N_A_c_117_n N_B_c_263_n 0.0117744f $X=1.74 $Y=1.425 $X2=0 $Y2=0
cc_135 N_A_c_118_n N_B_c_263_n 0.00361082f $X=2.465 $Y=1.09 $X2=0 $Y2=0
cc_136 N_A_c_121_n N_B_c_263_n 0.022528f $X=1.185 $Y=1.51 $X2=0 $Y2=0
cc_137 N_A_c_122_n N_B_c_263_n 0.020445f $X=3.545 $Y=1.49 $X2=0 $Y2=0
cc_138 N_A_c_123_n N_B_c_263_n 0.00715501f $X=1.655 $Y=1.587 $X2=0 $Y2=0
cc_139 N_A_M1000_g N_B_c_274_n 0.0111853f $X=2.65 $Y=2.465 $X2=0 $Y2=0
cc_140 N_A_M1010_g N_B_c_274_n 0.0120631f $X=3.08 $Y=2.465 $X2=0 $Y2=0
cc_141 N_A_c_118_n N_B_c_274_n 0.00421128f $X=2.465 $Y=1.09 $X2=0 $Y2=0
cc_142 N_A_c_120_n N_B_c_274_n 0.0130887f $X=2.635 $Y=1.49 $X2=0 $Y2=0
cc_143 N_A_c_162_p N_B_c_274_n 0.0349068f $X=2.97 $Y=1.49 $X2=0 $Y2=0
cc_144 N_A_c_122_n N_B_c_274_n 0.0084802f $X=3.545 $Y=1.49 $X2=0 $Y2=0
cc_145 N_A_M1010_g N_B_c_275_n 0.0035724f $X=3.08 $Y=2.465 $X2=0 $Y2=0
cc_146 N_A_c_162_p N_B_c_275_n 0.0142053f $X=2.97 $Y=1.49 $X2=0 $Y2=0
cc_147 N_A_c_122_n N_B_c_275_n 0.0158366f $X=3.545 $Y=1.49 $X2=0 $Y2=0
cc_148 N_A_c_122_n N_B_c_264_n 0.0100133f $X=3.545 $Y=1.49 $X2=0 $Y2=0
cc_149 N_A_c_118_n N_A_162_367#_M1002_s 0.00119515f $X=2.465 $Y=1.09 $X2=-0.19
+ $Y2=-0.245
cc_150 N_A_c_134_p N_A_162_367#_M1002_s 6.74726e-19 $X=1.825 $Y=1.09 $X2=-0.19
+ $Y2=-0.245
cc_151 N_A_M1007_g N_A_162_367#_c_399_n 0.00245293f $X=0.475 $Y=0.655 $X2=0
+ $Y2=0
cc_152 N_A_M1014_g N_A_162_367#_c_399_n 0.00927741f $X=0.735 $Y=2.465 $X2=0
+ $Y2=0
cc_153 N_A_M1019_g N_A_162_367#_c_399_n 0.0018136f $X=1.165 $Y=2.465 $X2=0 $Y2=0
cc_154 N_A_M1011_g N_A_162_367#_c_399_n 0.00202797f $X=1.205 $Y=0.655 $X2=0
+ $Y2=0
cc_155 N_A_c_121_n N_A_162_367#_c_399_n 0.0278882f $X=1.185 $Y=1.51 $X2=0 $Y2=0
cc_156 N_A_c_123_n N_A_162_367#_c_399_n 0.0252159f $X=1.655 $Y=1.587 $X2=0 $Y2=0
cc_157 N_A_M1011_g N_A_162_367#_c_400_n 0.0128736f $X=1.205 $Y=0.655 $X2=0 $Y2=0
cc_158 N_A_c_117_n N_A_162_367#_c_400_n 0.00561306f $X=1.74 $Y=1.425 $X2=0 $Y2=0
cc_159 N_A_c_134_p N_A_162_367#_c_400_n 0.00891437f $X=1.825 $Y=1.09 $X2=0 $Y2=0
cc_160 N_A_c_121_n N_A_162_367#_c_400_n 0.00770273f $X=1.185 $Y=1.51 $X2=0 $Y2=0
cc_161 N_A_c_123_n N_A_162_367#_c_400_n 0.034803f $X=1.655 $Y=1.587 $X2=0 $Y2=0
cc_162 N_A_M1007_g N_A_162_367#_c_401_n 0.00502091f $X=0.475 $Y=0.655 $X2=0
+ $Y2=0
cc_163 N_A_M1019_g N_A_162_367#_c_426_n 0.012943f $X=1.165 $Y=2.465 $X2=0 $Y2=0
cc_164 N_A_c_117_n N_A_162_367#_c_426_n 0.00578843f $X=1.74 $Y=1.425 $X2=0 $Y2=0
cc_165 N_A_c_121_n N_A_162_367#_c_426_n 5.25142e-19 $X=1.185 $Y=1.51 $X2=0 $Y2=0
cc_166 N_A_c_123_n N_A_162_367#_c_426_n 0.0392154f $X=1.655 $Y=1.587 $X2=0 $Y2=0
cc_167 N_A_c_134_p N_A_162_367#_c_430_n 0.00546539f $X=1.825 $Y=1.09 $X2=0 $Y2=0
cc_168 N_A_c_118_n N_A_162_367#_c_431_n 0.00881641f $X=2.465 $Y=1.09 $X2=0 $Y2=0
cc_169 N_A_c_134_p N_A_162_367#_c_431_n 0.00823273f $X=1.825 $Y=1.09 $X2=0 $Y2=0
cc_170 N_A_c_123_n N_A_162_367#_c_431_n 0.00389096f $X=1.655 $Y=1.587 $X2=0
+ $Y2=0
cc_171 N_A_c_117_n N_A_162_367#_c_434_n 0.00636257f $X=1.74 $Y=1.425 $X2=0 $Y2=0
cc_172 N_A_M1000_g N_A_162_367#_c_435_n 9.45037e-19 $X=2.65 $Y=2.465 $X2=0 $Y2=0
cc_173 N_A_M1000_g N_A_162_367#_c_407_n 0.0150283f $X=2.65 $Y=2.465 $X2=0 $Y2=0
cc_174 N_A_M1010_g N_A_162_367#_c_407_n 0.0123148f $X=3.08 $Y=2.465 $X2=0 $Y2=0
cc_175 N_A_c_122_n N_A_162_367#_c_407_n 0.00238084f $X=3.545 $Y=1.49 $X2=0 $Y2=0
cc_176 N_A_M1014_g N_A_162_367#_c_439_n 0.00980004f $X=0.735 $Y=2.465 $X2=0
+ $Y2=0
cc_177 N_A_c_121_n N_A_162_367#_c_439_n 0.00274074f $X=1.185 $Y=1.51 $X2=0 $Y2=0
cc_178 N_A_c_123_n N_A_162_367#_c_439_n 0.00246053f $X=1.655 $Y=1.587 $X2=0
+ $Y2=0
cc_179 N_A_M1010_g N_A_162_367#_c_410_n 0.00456339f $X=3.08 $Y=2.465 $X2=0 $Y2=0
cc_180 N_A_M1014_g N_VPWR_c_545_n 0.00922365f $X=0.735 $Y=2.465 $X2=0 $Y2=0
cc_181 N_A_c_121_n N_VPWR_c_545_n 0.0044942f $X=1.185 $Y=1.51 $X2=0 $Y2=0
cc_182 N_A_M1014_g N_VPWR_c_546_n 0.00531226f $X=0.735 $Y=2.465 $X2=0 $Y2=0
cc_183 N_A_M1014_g N_VPWR_c_547_n 6.69872e-19 $X=0.735 $Y=2.465 $X2=0 $Y2=0
cc_184 N_A_M1019_g N_VPWR_c_547_n 0.0130072f $X=1.165 $Y=2.465 $X2=0 $Y2=0
cc_185 N_A_M1000_g N_VPWR_c_548_n 0.00588516f $X=2.65 $Y=2.465 $X2=0 $Y2=0
cc_186 N_A_M1010_g N_VPWR_c_549_n 0.00327679f $X=3.08 $Y=2.465 $X2=0 $Y2=0
cc_187 N_A_M1014_g N_VPWR_c_553_n 0.00585385f $X=0.735 $Y=2.465 $X2=0 $Y2=0
cc_188 N_A_M1019_g N_VPWR_c_553_n 0.00564095f $X=1.165 $Y=2.465 $X2=0 $Y2=0
cc_189 N_A_M1000_g N_VPWR_c_557_n 0.0054895f $X=2.65 $Y=2.465 $X2=0 $Y2=0
cc_190 N_A_M1010_g N_VPWR_c_557_n 0.00426006f $X=3.08 $Y=2.465 $X2=0 $Y2=0
cc_191 N_A_M1014_g N_VPWR_c_544_n 0.0116391f $X=0.735 $Y=2.465 $X2=0 $Y2=0
cc_192 N_A_M1019_g N_VPWR_c_544_n 0.00948291f $X=1.165 $Y=2.465 $X2=0 $Y2=0
cc_193 N_A_M1000_g N_VPWR_c_544_n 0.0102673f $X=2.65 $Y=2.465 $X2=0 $Y2=0
cc_194 N_A_M1010_g N_VPWR_c_544_n 0.00710517f $X=3.08 $Y=2.465 $X2=0 $Y2=0
cc_195 N_A_M1010_g N_A_545_367#_c_639_n 0.0108475f $X=3.08 $Y=2.465 $X2=0 $Y2=0
cc_196 N_A_M1010_g N_A_545_367#_c_640_n 0.00256818f $X=3.08 $Y=2.465 $X2=0 $Y2=0
cc_197 N_A_M1000_g N_A_545_367#_c_645_n 0.00746658f $X=2.65 $Y=2.465 $X2=0 $Y2=0
cc_198 N_A_M1010_g N_A_545_367#_c_645_n 0.00790197f $X=3.08 $Y=2.465 $X2=0 $Y2=0
cc_199 N_A_c_118_n N_A_27_47#_M1018_d 0.00353704f $X=2.465 $Y=1.09 $X2=0 $Y2=0
cc_200 N_A_M1007_g N_A_27_47#_c_743_n 0.00889565f $X=0.475 $Y=0.655 $X2=0 $Y2=0
cc_201 N_A_M1007_g N_A_27_47#_c_748_n 0.0136669f $X=0.475 $Y=0.655 $X2=0 $Y2=0
cc_202 N_A_M1011_g N_A_27_47#_c_748_n 0.00514682f $X=1.205 $Y=0.655 $X2=0 $Y2=0
cc_203 N_A_c_121_n N_A_27_47#_c_748_n 0.00198223f $X=1.185 $Y=1.51 $X2=0 $Y2=0
cc_204 N_A_M1007_g N_A_27_47#_c_744_n 0.00983521f $X=0.475 $Y=0.655 $X2=0 $Y2=0
cc_205 N_A_M1007_g N_A_27_47#_c_752_n 0.00138166f $X=0.475 $Y=0.655 $X2=0 $Y2=0
cc_206 N_A_M1011_g N_A_27_47#_c_752_n 0.00756757f $X=1.205 $Y=0.655 $X2=0 $Y2=0
cc_207 N_A_M1011_g N_A_27_47#_c_754_n 0.0072419f $X=1.205 $Y=0.655 $X2=0 $Y2=0
cc_208 N_A_c_118_n N_A_27_47#_c_754_n 0.00320671f $X=2.465 $Y=1.09 $X2=0 $Y2=0
cc_209 N_A_M1011_g N_A_27_47#_c_756_n 0.00282553f $X=1.205 $Y=0.655 $X2=0 $Y2=0
cc_210 N_A_M1008_g N_A_27_47#_c_745_n 0.00114103f $X=3.115 $Y=0.745 $X2=0 $Y2=0
cc_211 N_A_c_118_n N_A_27_47#_c_745_n 0.0259298f $X=2.465 $Y=1.09 $X2=0 $Y2=0
cc_212 N_A_M1007_g N_VGND_c_795_n 0.00331076f $X=0.475 $Y=0.655 $X2=0 $Y2=0
cc_213 N_A_M1011_g N_VGND_c_795_n 0.00304214f $X=1.205 $Y=0.655 $X2=0 $Y2=0
cc_214 N_A_M1008_g N_VGND_c_796_n 0.0111934f $X=3.115 $Y=0.745 $X2=0 $Y2=0
cc_215 N_A_M1009_g N_VGND_c_796_n 0.00998341f $X=3.545 $Y=0.745 $X2=0 $Y2=0
cc_216 N_A_M1009_g N_VGND_c_797_n 0.00414769f $X=3.545 $Y=0.745 $X2=0 $Y2=0
cc_217 N_A_M1009_g N_VGND_c_798_n 4.95999e-19 $X=3.545 $Y=0.745 $X2=0 $Y2=0
cc_218 N_A_M1011_g N_VGND_c_799_n 0.00357856f $X=1.205 $Y=0.655 $X2=0 $Y2=0
cc_219 N_A_M1008_g N_VGND_c_799_n 0.00414769f $X=3.115 $Y=0.745 $X2=0 $Y2=0
cc_220 N_A_M1007_g N_VGND_c_801_n 0.00432561f $X=0.475 $Y=0.655 $X2=0 $Y2=0
cc_221 N_A_M1007_g N_VGND_c_803_n 0.00738357f $X=0.475 $Y=0.655 $X2=0 $Y2=0
cc_222 N_A_M1011_g N_VGND_c_803_n 0.0060181f $X=1.205 $Y=0.655 $X2=0 $Y2=0
cc_223 N_A_M1008_g N_VGND_c_803_n 0.00837493f $X=3.115 $Y=0.745 $X2=0 $Y2=0
cc_224 N_A_M1009_g N_VGND_c_803_n 0.0078848f $X=3.545 $Y=0.745 $X2=0 $Y2=0
cc_225 N_A_M1008_g N_A_555_65#_c_875_n 0.00365282f $X=3.115 $Y=0.745 $X2=0 $Y2=0
cc_226 N_A_c_118_n N_A_555_65#_c_875_n 0.00498735f $X=2.465 $Y=1.09 $X2=0 $Y2=0
cc_227 N_A_M1008_g N_A_555_65#_c_876_n 0.0140921f $X=3.115 $Y=0.745 $X2=0 $Y2=0
cc_228 N_A_M1009_g N_A_555_65#_c_876_n 0.0130264f $X=3.545 $Y=0.745 $X2=0 $Y2=0
cc_229 N_A_c_162_p N_A_555_65#_c_876_n 0.00961976f $X=2.97 $Y=1.49 $X2=0 $Y2=0
cc_230 N_A_c_122_n N_A_555_65#_c_876_n 0.00417303f $X=3.545 $Y=1.49 $X2=0 $Y2=0
cc_231 N_A_c_118_n N_A_555_65#_c_877_n 0.0101297f $X=2.465 $Y=1.09 $X2=0 $Y2=0
cc_232 N_A_c_119_n N_A_555_65#_c_877_n 0.0050297f $X=2.55 $Y=1.405 $X2=0 $Y2=0
cc_233 N_A_c_162_p N_A_555_65#_c_877_n 0.0153281f $X=2.97 $Y=1.49 $X2=0 $Y2=0
cc_234 N_A_c_122_n N_A_555_65#_c_877_n 0.00526567f $X=3.545 $Y=1.49 $X2=0 $Y2=0
cc_235 N_A_M1009_g N_A_555_65#_c_878_n 8.64821e-19 $X=3.545 $Y=0.745 $X2=0 $Y2=0
cc_236 N_B_M1017_g N_A_162_367#_M1003_g 0.0203867f $X=4.835 $Y=0.745 $X2=0 $Y2=0
cc_237 N_B_M1006_g N_A_162_367#_M1004_g 0.0186707f $X=4.905 $Y=2.465 $X2=0 $Y2=0
cc_238 N_B_M1002_g N_A_162_367#_c_400_n 0.00131507f $X=1.635 $Y=0.655 $X2=0
+ $Y2=0
cc_239 N_B_M1005_g N_A_162_367#_c_426_n 0.0129928f $X=1.635 $Y=2.465 $X2=0 $Y2=0
cc_240 N_B_M1002_g N_A_162_367#_c_430_n 0.00486726f $X=1.635 $Y=0.655 $X2=0
+ $Y2=0
cc_241 N_B_M1002_g N_A_162_367#_c_431_n 0.0100983f $X=1.635 $Y=0.655 $X2=0 $Y2=0
cc_242 N_B_M1018_g N_A_162_367#_c_431_n 0.00273619f $X=2.065 $Y=0.655 $X2=0
+ $Y2=0
cc_243 N_B_M1015_g N_A_162_367#_c_434_n 8.55391e-19 $X=2.065 $Y=2.465 $X2=0
+ $Y2=0
cc_244 N_B_c_262_n N_A_162_367#_c_434_n 7.8471e-19 $X=2.09 $Y=1.51 $X2=0 $Y2=0
cc_245 N_B_c_263_n N_A_162_367#_c_434_n 0.00323808f $X=2.09 $Y=1.51 $X2=0 $Y2=0
cc_246 N_B_M1015_g N_A_162_367#_c_435_n 0.0110002f $X=2.065 $Y=2.465 $X2=0 $Y2=0
cc_247 N_B_M1015_g N_A_162_367#_c_407_n 0.0126967f $X=2.065 $Y=2.465 $X2=0 $Y2=0
cc_248 N_B_c_262_n N_A_162_367#_c_407_n 0.012437f $X=2.09 $Y=1.51 $X2=0 $Y2=0
cc_249 N_B_c_263_n N_A_162_367#_c_407_n 3.89763e-19 $X=2.09 $Y=1.51 $X2=0 $Y2=0
cc_250 N_B_c_274_n N_A_162_367#_c_407_n 0.0703711f $X=3.305 $Y=1.66 $X2=0 $Y2=0
cc_251 N_B_c_264_n N_A_162_367#_c_407_n 0.00843205f $X=4.335 $Y=1.51 $X2=0 $Y2=0
cc_252 N_B_M1001_g N_A_162_367#_c_408_n 0.013762f $X=4.475 $Y=2.465 $X2=0 $Y2=0
cc_253 N_B_M1006_g N_A_162_367#_c_408_n 0.00411163f $X=4.905 $Y=2.465 $X2=0
+ $Y2=0
cc_254 N_B_c_259_n N_A_162_367#_c_408_n 0.00301802f $X=4.05 $Y=1.51 $X2=0 $Y2=0
cc_255 N_B_c_261_n N_A_162_367#_c_408_n 0.00159823f $X=4.905 $Y=1.51 $X2=0 $Y2=0
cc_256 N_B_c_264_n N_A_162_367#_c_408_n 0.0481042f $X=4.335 $Y=1.51 $X2=0 $Y2=0
cc_257 N_B_M1001_g N_A_162_367#_c_409_n 0.00412209f $X=4.475 $Y=2.465 $X2=0
+ $Y2=0
cc_258 N_B_M1006_g N_A_162_367#_c_409_n 0.00492387f $X=4.905 $Y=2.465 $X2=0
+ $Y2=0
cc_259 N_B_c_261_n N_A_162_367#_c_409_n 0.00421111f $X=4.905 $Y=1.51 $X2=0 $Y2=0
cc_260 N_B_c_264_n N_A_162_367#_c_409_n 0.0104549f $X=4.335 $Y=1.51 $X2=0 $Y2=0
cc_261 N_B_c_261_n N_A_162_367#_c_468_n 0.00867263f $X=4.905 $Y=1.51 $X2=0 $Y2=0
cc_262 N_B_c_264_n N_A_162_367#_c_468_n 0.015729f $X=4.335 $Y=1.51 $X2=0 $Y2=0
cc_263 N_B_c_261_n N_A_162_367#_c_402_n 0.00890874f $X=4.905 $Y=1.51 $X2=0 $Y2=0
cc_264 N_B_M1001_g N_A_162_367#_c_410_n 0.00401662f $X=4.475 $Y=2.465 $X2=0
+ $Y2=0
cc_265 N_B_c_264_n N_A_162_367#_c_410_n 0.0174786f $X=4.335 $Y=1.51 $X2=0 $Y2=0
cc_266 N_B_c_261_n N_A_162_367#_c_403_n 0.0234857f $X=4.905 $Y=1.51 $X2=0 $Y2=0
cc_267 N_B_c_262_n N_VPWR_M1015_s 9.70984e-19 $X=2.09 $Y=1.51 $X2=0 $Y2=0
cc_268 N_B_c_274_n N_VPWR_M1015_s 0.00273991f $X=3.305 $Y=1.66 $X2=0 $Y2=0
cc_269 N_B_c_274_n N_VPWR_M1010_d 0.00100313f $X=3.305 $Y=1.66 $X2=0 $Y2=0
cc_270 N_B_c_275_n N_VPWR_M1010_d 0.00194712f $X=3.475 $Y=1.66 $X2=0 $Y2=0
cc_271 N_B_M1005_g N_VPWR_c_547_n 0.0132783f $X=1.635 $Y=2.465 $X2=0 $Y2=0
cc_272 N_B_M1015_g N_VPWR_c_547_n 7.16162e-19 $X=2.065 $Y=2.465 $X2=0 $Y2=0
cc_273 N_B_M1015_g N_VPWR_c_548_n 0.00576643f $X=2.065 $Y=2.465 $X2=0 $Y2=0
cc_274 N_B_M1006_g N_VPWR_c_550_n 0.001275f $X=4.905 $Y=2.465 $X2=0 $Y2=0
cc_275 N_B_M1005_g N_VPWR_c_555_n 0.00564095f $X=1.635 $Y=2.465 $X2=0 $Y2=0
cc_276 N_B_M1015_g N_VPWR_c_555_n 0.0054895f $X=2.065 $Y=2.465 $X2=0 $Y2=0
cc_277 N_B_M1001_g N_VPWR_c_559_n 0.00361434f $X=4.475 $Y=2.465 $X2=0 $Y2=0
cc_278 N_B_M1006_g N_VPWR_c_559_n 0.00549284f $X=4.905 $Y=2.465 $X2=0 $Y2=0
cc_279 N_B_M1005_g N_VPWR_c_544_n 0.00948291f $X=1.635 $Y=2.465 $X2=0 $Y2=0
cc_280 N_B_M1015_g N_VPWR_c_544_n 0.010281f $X=2.065 $Y=2.465 $X2=0 $Y2=0
cc_281 N_B_M1001_g N_VPWR_c_544_n 0.00681415f $X=4.475 $Y=2.465 $X2=0 $Y2=0
cc_282 N_B_M1006_g N_VPWR_c_544_n 0.0100092f $X=4.905 $Y=2.465 $X2=0 $Y2=0
cc_283 N_B_c_274_n N_A_545_367#_M1000_s 0.00176891f $X=3.305 $Y=1.66 $X2=-0.19
+ $Y2=-0.245
cc_284 N_B_M1001_g N_A_545_367#_c_640_n 0.0040562f $X=4.475 $Y=2.465 $X2=0 $Y2=0
cc_285 N_B_M1001_g N_A_545_367#_c_641_n 0.0111082f $X=4.475 $Y=2.465 $X2=0 $Y2=0
cc_286 N_B_M1001_g N_A_545_367#_c_650_n 0.00937059f $X=4.475 $Y=2.465 $X2=0
+ $Y2=0
cc_287 N_B_M1006_g N_A_545_367#_c_650_n 0.0069768f $X=4.905 $Y=2.465 $X2=0 $Y2=0
cc_288 N_B_M1001_g N_Y_c_692_n 0.00963526f $X=4.475 $Y=2.465 $X2=0 $Y2=0
cc_289 N_B_M1006_g N_Y_c_692_n 0.0140412f $X=4.905 $Y=2.465 $X2=0 $Y2=0
cc_290 N_B_c_261_n N_Y_c_692_n 2.23325e-19 $X=4.905 $Y=1.51 $X2=0 $Y2=0
cc_291 N_B_M1006_g N_Y_c_687_n 4.90985e-19 $X=4.905 $Y=2.465 $X2=0 $Y2=0
cc_292 N_B_M1002_g N_A_27_47#_c_752_n 6.72995e-19 $X=1.635 $Y=0.655 $X2=0 $Y2=0
cc_293 N_B_M1002_g N_A_27_47#_c_754_n 0.0082158f $X=1.635 $Y=0.655 $X2=0 $Y2=0
cc_294 N_B_M1018_g N_A_27_47#_c_754_n 0.013826f $X=2.065 $Y=0.655 $X2=0 $Y2=0
cc_295 N_B_M1016_g N_VGND_c_796_n 4.93338e-19 $X=3.975 $Y=0.745 $X2=0 $Y2=0
cc_296 N_B_M1016_g N_VGND_c_797_n 0.00414769f $X=3.975 $Y=0.745 $X2=0 $Y2=0
cc_297 N_B_M1016_g N_VGND_c_798_n 0.0111902f $X=3.975 $Y=0.745 $X2=0 $Y2=0
cc_298 N_B_M1017_g N_VGND_c_798_n 0.0112864f $X=4.835 $Y=0.745 $X2=0 $Y2=0
cc_299 N_B_M1002_g N_VGND_c_799_n 0.00357877f $X=1.635 $Y=0.655 $X2=0 $Y2=0
cc_300 N_B_M1018_g N_VGND_c_799_n 0.00357877f $X=2.065 $Y=0.655 $X2=0 $Y2=0
cc_301 N_B_M1017_g N_VGND_c_802_n 0.00414769f $X=4.835 $Y=0.745 $X2=0 $Y2=0
cc_302 N_B_M1002_g N_VGND_c_803_n 0.00537654f $X=1.635 $Y=0.655 $X2=0 $Y2=0
cc_303 N_B_M1018_g N_VGND_c_803_n 0.0068216f $X=2.065 $Y=0.655 $X2=0 $Y2=0
cc_304 N_B_M1016_g N_VGND_c_803_n 0.0078848f $X=3.975 $Y=0.745 $X2=0 $Y2=0
cc_305 N_B_M1017_g N_VGND_c_803_n 0.0078848f $X=4.835 $Y=0.745 $X2=0 $Y2=0
cc_306 N_B_M1018_g N_A_555_65#_c_875_n 0.00479376f $X=2.065 $Y=0.655 $X2=0 $Y2=0
cc_307 N_B_c_274_n N_A_555_65#_c_876_n 0.00392282f $X=3.305 $Y=1.66 $X2=0 $Y2=0
cc_308 N_B_c_275_n N_A_555_65#_c_876_n 0.0270949f $X=3.475 $Y=1.66 $X2=0 $Y2=0
cc_309 N_B_M1018_g N_A_555_65#_c_877_n 4.17289e-19 $X=2.065 $Y=0.655 $X2=0 $Y2=0
cc_310 N_B_M1016_g N_A_555_65#_c_878_n 8.64821e-19 $X=3.975 $Y=0.745 $X2=0 $Y2=0
cc_311 N_B_M1016_g N_A_555_65#_c_879_n 0.0146446f $X=3.975 $Y=0.745 $X2=0 $Y2=0
cc_312 N_B_M1017_g N_A_555_65#_c_879_n 0.0144775f $X=4.835 $Y=0.745 $X2=0 $Y2=0
cc_313 N_B_c_259_n N_A_555_65#_c_879_n 0.00108047f $X=4.05 $Y=1.51 $X2=0 $Y2=0
cc_314 N_B_c_260_n N_A_555_65#_c_879_n 0.0164675f $X=4.4 $Y=1.51 $X2=0 $Y2=0
cc_315 N_B_c_261_n N_A_555_65#_c_879_n 0.00200127f $X=4.905 $Y=1.51 $X2=0 $Y2=0
cc_316 N_B_c_264_n N_A_555_65#_c_879_n 0.0479655f $X=4.335 $Y=1.51 $X2=0 $Y2=0
cc_317 N_B_M1017_g N_A_555_65#_c_881_n 5.73473e-19 $X=4.835 $Y=0.745 $X2=0 $Y2=0
cc_318 N_B_c_259_n N_A_555_65#_c_883_n 6.26322e-19 $X=4.05 $Y=1.51 $X2=0 $Y2=0
cc_319 N_B_c_264_n N_A_555_65#_c_883_n 0.0167573f $X=4.335 $Y=1.51 $X2=0 $Y2=0
cc_320 N_A_162_367#_c_426_n N_VPWR_M1019_d 0.00427624f $X=1.745 $Y=2.005 $X2=0
+ $Y2=0
cc_321 N_A_162_367#_c_407_n N_VPWR_M1015_s 0.00745115f $X=3.645 $Y=2.17 $X2=0
+ $Y2=0
cc_322 N_A_162_367#_c_407_n N_VPWR_M1010_d 0.00557361f $X=3.645 $Y=2.17 $X2=0
+ $Y2=0
cc_323 N_A_162_367#_c_399_n N_VPWR_c_545_n 0.00748789f $X=0.765 $Y=1.92 $X2=0
+ $Y2=0
cc_324 N_A_162_367#_c_439_n N_VPWR_c_545_n 0.0143242f $X=0.95 $Y=2.015 $X2=0
+ $Y2=0
cc_325 N_A_162_367#_c_426_n N_VPWR_c_547_n 0.017285f $X=1.745 $Y=2.005 $X2=0
+ $Y2=0
cc_326 N_A_162_367#_c_407_n N_VPWR_c_548_n 0.0250231f $X=3.645 $Y=2.17 $X2=0
+ $Y2=0
cc_327 N_A_162_367#_M1004_g N_VPWR_c_550_n 0.0152499f $X=5.335 $Y=2.465 $X2=0
+ $Y2=0
cc_328 N_A_162_367#_M1013_g N_VPWR_c_550_n 0.0160463f $X=5.765 $Y=2.465 $X2=0
+ $Y2=0
cc_329 N_A_162_367#_c_483_p N_VPWR_c_553_n 0.0145813f $X=0.95 $Y=2.475 $X2=0
+ $Y2=0
cc_330 N_A_162_367#_c_435_n N_VPWR_c_555_n 0.0160429f $X=1.85 $Y=2.91 $X2=0
+ $Y2=0
cc_331 N_A_162_367#_M1004_g N_VPWR_c_559_n 0.00486043f $X=5.335 $Y=2.465 $X2=0
+ $Y2=0
cc_332 N_A_162_367#_M1013_g N_VPWR_c_560_n 0.00486043f $X=5.765 $Y=2.465 $X2=0
+ $Y2=0
cc_333 N_A_162_367#_M1014_s N_VPWR_c_544_n 0.00327921f $X=0.81 $Y=1.835 $X2=0
+ $Y2=0
cc_334 N_A_162_367#_M1005_d N_VPWR_c_544_n 0.00345315f $X=1.71 $Y=1.835 $X2=0
+ $Y2=0
cc_335 N_A_162_367#_M1004_g N_VPWR_c_544_n 0.0082726f $X=5.335 $Y=2.465 $X2=0
+ $Y2=0
cc_336 N_A_162_367#_M1013_g N_VPWR_c_544_n 0.00917987f $X=5.765 $Y=2.465 $X2=0
+ $Y2=0
cc_337 N_A_162_367#_c_483_p N_VPWR_c_544_n 0.0096311f $X=0.95 $Y=2.475 $X2=0
+ $Y2=0
cc_338 N_A_162_367#_c_435_n N_VPWR_c_544_n 0.0102362f $X=1.85 $Y=2.91 $X2=0
+ $Y2=0
cc_339 N_A_162_367#_c_407_n N_A_545_367#_M1000_s 0.00343569f $X=3.645 $Y=2.17
+ $X2=-0.19 $Y2=-0.245
cc_340 N_A_162_367#_c_408_n N_A_545_367#_M1001_s 0.00358483f $X=4.685 $Y=2.005
+ $X2=0 $Y2=0
cc_341 N_A_162_367#_c_409_n N_A_545_367#_M1001_s 9.53615e-19 $X=4.77 $Y=1.92
+ $X2=0 $Y2=0
cc_342 N_A_162_367#_c_407_n N_A_545_367#_c_639_n 0.038847f $X=3.645 $Y=2.17
+ $X2=0 $Y2=0
cc_343 N_A_162_367#_c_410_n N_A_545_367#_c_639_n 0.0176587f $X=3.75 $Y=2.005
+ $X2=0 $Y2=0
cc_344 N_A_162_367#_c_407_n N_A_545_367#_c_645_n 0.0164161f $X=3.645 $Y=2.17
+ $X2=0 $Y2=0
cc_345 N_A_162_367#_c_408_n N_Y_M1001_d 0.00479121f $X=4.685 $Y=2.005 $X2=0
+ $Y2=0
cc_346 N_A_162_367#_c_408_n N_Y_c_692_n 0.0247445f $X=4.685 $Y=2.005 $X2=0 $Y2=0
cc_347 N_A_162_367#_c_402_n N_Y_c_692_n 0.00344099f $X=5.55 $Y=1.51 $X2=0 $Y2=0
cc_348 N_A_162_367#_M1004_g N_Y_c_686_n 0.0128162f $X=5.335 $Y=2.465 $X2=0 $Y2=0
cc_349 N_A_162_367#_M1013_g N_Y_c_686_n 0.0146735f $X=5.765 $Y=2.465 $X2=0 $Y2=0
cc_350 N_A_162_367#_c_402_n N_Y_c_686_n 0.0355003f $X=5.55 $Y=1.51 $X2=0 $Y2=0
cc_351 N_A_162_367#_c_403_n N_Y_c_686_n 0.00401774f $X=5.765 $Y=1.51 $X2=0 $Y2=0
cc_352 N_A_162_367#_c_409_n N_Y_c_687_n 0.00765392f $X=4.77 $Y=1.92 $X2=0 $Y2=0
cc_353 N_A_162_367#_c_402_n N_Y_c_687_n 0.0161304f $X=5.55 $Y=1.51 $X2=0 $Y2=0
cc_354 N_A_162_367#_c_403_n N_Y_c_687_n 7.40448e-19 $X=5.765 $Y=1.51 $X2=0 $Y2=0
cc_355 N_A_162_367#_M1012_g N_Y_c_682_n 0.0113653f $X=5.695 $Y=0.745 $X2=0 $Y2=0
cc_356 N_A_162_367#_c_402_n N_Y_c_682_n 0.0047708f $X=5.55 $Y=1.51 $X2=0 $Y2=0
cc_357 N_A_162_367#_c_403_n N_Y_c_682_n 0.00227732f $X=5.765 $Y=1.51 $X2=0 $Y2=0
cc_358 N_A_162_367#_M1003_g N_Y_c_683_n 0.00288365f $X=5.265 $Y=0.745 $X2=0
+ $Y2=0
cc_359 N_A_162_367#_M1012_g N_Y_c_683_n 0.00156191f $X=5.695 $Y=0.745 $X2=0
+ $Y2=0
cc_360 N_A_162_367#_c_402_n N_Y_c_683_n 0.0265505f $X=5.55 $Y=1.51 $X2=0 $Y2=0
cc_361 N_A_162_367#_c_403_n N_Y_c_683_n 0.00279085f $X=5.765 $Y=1.51 $X2=0 $Y2=0
cc_362 N_A_162_367#_c_408_n N_Y_c_688_n 0.019272f $X=4.685 $Y=2.005 $X2=0 $Y2=0
cc_363 N_A_162_367#_M1003_g N_Y_c_714_n 0.00506661f $X=5.265 $Y=0.745 $X2=0
+ $Y2=0
cc_364 N_A_162_367#_M1012_g N_Y_c_714_n 0.0108478f $X=5.695 $Y=0.745 $X2=0 $Y2=0
cc_365 N_A_162_367#_M1012_g Y 0.00418691f $X=5.695 $Y=0.745 $X2=0 $Y2=0
cc_366 N_A_162_367#_c_402_n Y 0.0163654f $X=5.55 $Y=1.51 $X2=0 $Y2=0
cc_367 N_A_162_367#_c_403_n Y 0.0165762f $X=5.765 $Y=1.51 $X2=0 $Y2=0
cc_368 N_A_162_367#_c_430_n N_A_27_47#_M1011_s 0.00289906f $X=1.4 $Y=1.075 $X2=0
+ $Y2=0
cc_369 N_A_162_367#_c_523_p N_A_27_47#_M1011_s 0.0020224f $X=1.485 $Y=0.715
+ $X2=0 $Y2=0
cc_370 N_A_162_367#_c_431_n N_A_27_47#_M1011_s 5.17671e-19 $X=1.85 $Y=0.71 $X2=0
+ $Y2=0
cc_371 N_A_162_367#_c_400_n N_A_27_47#_c_748_n 0.0205395f $X=1.315 $Y=1.16 $X2=0
+ $Y2=0
cc_372 N_A_162_367#_c_401_n N_A_27_47#_c_748_n 0.0138309f $X=0.85 $Y=1.16 $X2=0
+ $Y2=0
cc_373 N_A_162_367#_c_401_n N_A_27_47#_c_744_n 0.00125018f $X=0.85 $Y=1.16 $X2=0
+ $Y2=0
cc_374 N_A_162_367#_M1002_s N_A_27_47#_c_754_n 0.00333918f $X=1.71 $Y=0.235
+ $X2=0 $Y2=0
cc_375 N_A_162_367#_c_400_n N_A_27_47#_c_754_n 0.00359918f $X=1.315 $Y=1.16
+ $X2=0 $Y2=0
cc_376 N_A_162_367#_c_523_p N_A_27_47#_c_754_n 0.011337f $X=1.485 $Y=0.715 $X2=0
+ $Y2=0
cc_377 N_A_162_367#_c_431_n N_A_27_47#_c_754_n 0.0241955f $X=1.85 $Y=0.71 $X2=0
+ $Y2=0
cc_378 N_A_162_367#_c_401_n N_VGND_M1007_d 0.00188589f $X=0.85 $Y=1.16 $X2=-0.19
+ $Y2=-0.245
cc_379 N_A_162_367#_M1003_g N_VGND_c_798_n 5.37457e-19 $X=5.265 $Y=0.745 $X2=0
+ $Y2=0
cc_380 N_A_162_367#_M1003_g N_VGND_c_802_n 0.00302501f $X=5.265 $Y=0.745 $X2=0
+ $Y2=0
cc_381 N_A_162_367#_M1012_g N_VGND_c_802_n 0.00302501f $X=5.695 $Y=0.745 $X2=0
+ $Y2=0
cc_382 N_A_162_367#_M1002_s N_VGND_c_803_n 0.00225186f $X=1.71 $Y=0.235 $X2=0
+ $Y2=0
cc_383 N_A_162_367#_M1003_g N_VGND_c_803_n 0.00435646f $X=5.265 $Y=0.745 $X2=0
+ $Y2=0
cc_384 N_A_162_367#_M1012_g N_VGND_c_803_n 0.00472841f $X=5.695 $Y=0.745 $X2=0
+ $Y2=0
cc_385 N_A_162_367#_M1003_g N_A_555_65#_c_879_n 5.72e-19 $X=5.265 $Y=0.745 $X2=0
+ $Y2=0
cc_386 N_A_162_367#_c_468_n N_A_555_65#_c_879_n 0.0132395f $X=4.855 $Y=1.505
+ $X2=0 $Y2=0
cc_387 N_A_162_367#_c_402_n N_A_555_65#_c_879_n 0.0230901f $X=5.55 $Y=1.51 $X2=0
+ $Y2=0
cc_388 N_A_162_367#_M1003_g N_A_555_65#_c_880_n 0.0118056f $X=5.265 $Y=0.745
+ $X2=0 $Y2=0
cc_389 N_A_162_367#_M1012_g N_A_555_65#_c_880_n 0.0126954f $X=5.695 $Y=0.745
+ $X2=0 $Y2=0
cc_390 N_VPWR_c_544_n N_A_545_367#_M1000_s 0.00223559f $X=6 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_391 N_VPWR_c_544_n N_A_545_367#_M1001_s 0.0022543f $X=6 $Y=3.33 $X2=0 $Y2=0
cc_392 N_VPWR_M1010_d N_A_545_367#_c_639_n 0.00582806f $X=3.155 $Y=1.835 $X2=0
+ $Y2=0
cc_393 N_VPWR_c_549_n N_A_545_367#_c_639_n 0.0193779f $X=3.295 $Y=2.94 $X2=0
+ $Y2=0
cc_394 N_VPWR_c_557_n N_A_545_367#_c_639_n 0.00200585f $X=3.2 $Y=3.33 $X2=0
+ $Y2=0
cc_395 N_VPWR_c_559_n N_A_545_367#_c_639_n 0.00256966f $X=5.385 $Y=3.33 $X2=0
+ $Y2=0
cc_396 N_VPWR_c_544_n N_A_545_367#_c_639_n 0.00940983f $X=6 $Y=3.33 $X2=0 $Y2=0
cc_397 N_VPWR_c_549_n N_A_545_367#_c_640_n 0.00949429f $X=3.295 $Y=2.94 $X2=0
+ $Y2=0
cc_398 N_VPWR_c_559_n N_A_545_367#_c_641_n 0.0384694f $X=5.385 $Y=3.33 $X2=0
+ $Y2=0
cc_399 N_VPWR_c_544_n N_A_545_367#_c_641_n 0.0244636f $X=6 $Y=3.33 $X2=0 $Y2=0
cc_400 N_VPWR_c_549_n N_A_545_367#_c_642_n 0.0147863f $X=3.295 $Y=2.94 $X2=0
+ $Y2=0
cc_401 N_VPWR_c_559_n N_A_545_367#_c_642_n 0.0150834f $X=5.385 $Y=3.33 $X2=0
+ $Y2=0
cc_402 N_VPWR_c_544_n N_A_545_367#_c_642_n 0.00868788f $X=6 $Y=3.33 $X2=0 $Y2=0
cc_403 N_VPWR_c_557_n N_A_545_367#_c_645_n 0.0188581f $X=3.2 $Y=3.33 $X2=0 $Y2=0
cc_404 N_VPWR_c_544_n N_A_545_367#_c_645_n 0.0123659f $X=6 $Y=3.33 $X2=0 $Y2=0
cc_405 N_VPWR_c_559_n N_A_545_367#_c_650_n 0.0174777f $X=5.385 $Y=3.33 $X2=0
+ $Y2=0
cc_406 N_VPWR_c_544_n N_A_545_367#_c_650_n 0.0123432f $X=6 $Y=3.33 $X2=0 $Y2=0
cc_407 N_VPWR_c_544_n N_Y_M1001_d 0.00216245f $X=6 $Y=3.33 $X2=0 $Y2=0
cc_408 N_VPWR_c_544_n N_Y_M1006_d 0.00536646f $X=6 $Y=3.33 $X2=0 $Y2=0
cc_409 N_VPWR_c_544_n N_Y_M1013_d 0.00371702f $X=6 $Y=3.33 $X2=0 $Y2=0
cc_410 N_VPWR_c_559_n N_Y_c_722_n 0.0124525f $X=5.385 $Y=3.33 $X2=0 $Y2=0
cc_411 N_VPWR_c_544_n N_Y_c_722_n 0.00730901f $X=6 $Y=3.33 $X2=0 $Y2=0
cc_412 N_VPWR_M1004_s N_Y_c_686_n 0.00176461f $X=5.41 $Y=1.835 $X2=0 $Y2=0
cc_413 N_VPWR_c_550_n N_Y_c_686_n 0.0170777f $X=5.55 $Y=2.2 $X2=0 $Y2=0
cc_414 N_VPWR_c_560_n Y 0.018528f $X=6 $Y=3.33 $X2=0 $Y2=0
cc_415 N_VPWR_c_544_n Y 0.0104192f $X=6 $Y=3.33 $X2=0 $Y2=0
cc_416 N_A_545_367#_c_641_n N_Y_M1001_d 0.00546453f $X=4.525 $Y=2.98 $X2=0 $Y2=0
cc_417 N_A_545_367#_M1001_s N_Y_c_692_n 0.00342676f $X=4.55 $Y=1.835 $X2=0 $Y2=0
cc_418 N_A_545_367#_c_641_n N_Y_c_692_n 0.00372874f $X=4.525 $Y=2.98 $X2=0 $Y2=0
cc_419 N_A_545_367#_c_650_n N_Y_c_692_n 0.0165605f $X=4.69 $Y=2.725 $X2=0 $Y2=0
cc_420 N_A_545_367#_c_639_n N_Y_c_688_n 0.0116101f $X=3.63 $Y=2.52 $X2=0 $Y2=0
cc_421 N_A_545_367#_c_640_n N_Y_c_688_n 0.00184295f $X=3.742 $Y=2.895 $X2=0
+ $Y2=0
cc_422 N_A_545_367#_c_641_n N_Y_c_688_n 0.0126403f $X=4.525 $Y=2.98 $X2=0 $Y2=0
cc_423 N_Y_c_682_n N_A_555_65#_M1012_s 6.05921e-19 $X=5.885 $Y=1.15 $X2=0 $Y2=0
cc_424 N_Y_c_684_n N_A_555_65#_M1012_s 0.0032925f $X=6.02 $Y=1.235 $X2=0 $Y2=0
cc_425 N_Y_c_683_n N_A_555_65#_c_879_n 0.0104256f $X=5.645 $Y=1.15 $X2=0 $Y2=0
cc_426 N_Y_M1003_d N_A_555_65#_c_880_n 0.00176461f $X=5.34 $Y=0.325 $X2=0 $Y2=0
cc_427 N_Y_c_682_n N_A_555_65#_c_880_n 0.00280043f $X=5.885 $Y=1.15 $X2=0 $Y2=0
cc_428 N_Y_c_714_n N_A_555_65#_c_880_n 0.0159058f $X=5.48 $Y=0.68 $X2=0 $Y2=0
cc_429 N_Y_c_682_n N_A_555_65#_c_882_n 0.00465902f $X=5.885 $Y=1.15 $X2=0 $Y2=0
cc_430 N_Y_c_684_n N_A_555_65#_c_882_n 0.0233844f $X=6.02 $Y=1.235 $X2=0 $Y2=0
cc_431 N_A_27_47#_c_748_n N_VGND_M1007_d 0.012905f $X=0.975 $Y=0.82 $X2=-0.19
+ $Y2=-0.245
cc_432 N_A_27_47#_c_752_n N_VGND_M1007_d 0.00354625f $X=1.06 $Y=0.735 $X2=-0.19
+ $Y2=-0.245
cc_433 N_A_27_47#_c_756_n N_VGND_M1007_d 0.00278279f $X=1.145 $Y=0.35 $X2=-0.19
+ $Y2=-0.245
cc_434 N_A_27_47#_c_748_n N_VGND_c_795_n 0.0154494f $X=0.975 $Y=0.82 $X2=0 $Y2=0
cc_435 N_A_27_47#_c_752_n N_VGND_c_795_n 0.00885133f $X=1.06 $Y=0.735 $X2=0
+ $Y2=0
cc_436 N_A_27_47#_c_756_n N_VGND_c_795_n 0.0157311f $X=1.145 $Y=0.35 $X2=0 $Y2=0
cc_437 N_A_27_47#_c_745_n N_VGND_c_796_n 0.00137251f $X=2.35 $Y=0.38 $X2=0 $Y2=0
cc_438 N_A_27_47#_c_748_n N_VGND_c_799_n 0.00239315f $X=0.975 $Y=0.82 $X2=0
+ $Y2=0
cc_439 N_A_27_47#_c_754_n N_VGND_c_799_n 0.0577029f $X=2.185 $Y=0.35 $X2=0 $Y2=0
cc_440 N_A_27_47#_c_756_n N_VGND_c_799_n 0.00990952f $X=1.145 $Y=0.35 $X2=0
+ $Y2=0
cc_441 N_A_27_47#_c_745_n N_VGND_c_799_n 0.022581f $X=2.35 $Y=0.38 $X2=0 $Y2=0
cc_442 N_A_27_47#_c_743_n N_VGND_c_801_n 0.0203649f $X=0.26 $Y=0.42 $X2=0 $Y2=0
cc_443 N_A_27_47#_c_748_n N_VGND_c_801_n 0.00188649f $X=0.975 $Y=0.82 $X2=0
+ $Y2=0
cc_444 N_A_27_47#_M1007_s N_VGND_c_803_n 0.00215158f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_445 N_A_27_47#_M1011_s N_VGND_c_803_n 0.00223577f $X=1.28 $Y=0.235 $X2=0
+ $Y2=0
cc_446 N_A_27_47#_M1018_d N_VGND_c_803_n 0.00274611f $X=2.14 $Y=0.235 $X2=0
+ $Y2=0
cc_447 N_A_27_47#_c_743_n N_VGND_c_803_n 0.0122259f $X=0.26 $Y=0.42 $X2=0 $Y2=0
cc_448 N_A_27_47#_c_748_n N_VGND_c_803_n 0.00890918f $X=0.975 $Y=0.82 $X2=0
+ $Y2=0
cc_449 N_A_27_47#_c_744_n N_VGND_c_803_n 2.22564e-19 $X=0.425 $Y=0.82 $X2=0
+ $Y2=0
cc_450 N_A_27_47#_c_754_n N_VGND_c_803_n 0.0370643f $X=2.185 $Y=0.35 $X2=0 $Y2=0
cc_451 N_A_27_47#_c_756_n N_VGND_c_803_n 0.00653273f $X=1.145 $Y=0.35 $X2=0
+ $Y2=0
cc_452 N_A_27_47#_c_745_n N_VGND_c_803_n 0.0127769f $X=2.35 $Y=0.38 $X2=0 $Y2=0
cc_453 N_A_27_47#_c_745_n N_A_555_65#_c_875_n 0.0292265f $X=2.35 $Y=0.38 $X2=0
+ $Y2=0
cc_454 N_VGND_c_796_n N_A_555_65#_c_875_n 0.0232442f $X=3.33 $Y=0.45 $X2=0 $Y2=0
cc_455 N_VGND_c_799_n N_A_555_65#_c_875_n 0.0104816f $X=3.165 $Y=0 $X2=0 $Y2=0
cc_456 N_VGND_c_803_n N_A_555_65#_c_875_n 0.00714481f $X=6 $Y=0 $X2=0 $Y2=0
cc_457 N_VGND_M1008_d N_A_555_65#_c_876_n 0.00176461f $X=3.19 $Y=0.325 $X2=0
+ $Y2=0
cc_458 N_VGND_c_796_n N_A_555_65#_c_876_n 0.0170777f $X=3.33 $Y=0.45 $X2=0 $Y2=0
cc_459 N_VGND_c_796_n N_A_555_65#_c_878_n 0.0232442f $X=3.33 $Y=0.45 $X2=0 $Y2=0
cc_460 N_VGND_c_797_n N_A_555_65#_c_878_n 0.0104816f $X=4.025 $Y=0 $X2=0 $Y2=0
cc_461 N_VGND_c_798_n N_A_555_65#_c_878_n 0.0258638f $X=4.62 $Y=0.45 $X2=0 $Y2=0
cc_462 N_VGND_c_803_n N_A_555_65#_c_878_n 0.00714481f $X=6 $Y=0 $X2=0 $Y2=0
cc_463 N_VGND_M1016_s N_A_555_65#_c_879_n 0.00825348f $X=4.05 $Y=0.325 $X2=0
+ $Y2=0
cc_464 N_VGND_c_798_n N_A_555_65#_c_879_n 0.0520618f $X=4.62 $Y=0.45 $X2=0 $Y2=0
cc_465 N_VGND_c_802_n N_A_555_65#_c_880_n 0.0657775f $X=6 $Y=0 $X2=0 $Y2=0
cc_466 N_VGND_c_803_n N_A_555_65#_c_880_n 0.0366266f $X=6 $Y=0 $X2=0 $Y2=0
cc_467 N_VGND_c_798_n N_A_555_65#_c_881_n 0.0103779f $X=4.62 $Y=0.45 $X2=0 $Y2=0
cc_468 N_VGND_c_802_n N_A_555_65#_c_881_n 0.0136205f $X=6 $Y=0 $X2=0 $Y2=0
cc_469 N_VGND_c_803_n N_A_555_65#_c_881_n 0.00738676f $X=6 $Y=0 $X2=0 $Y2=0
