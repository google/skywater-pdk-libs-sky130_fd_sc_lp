* NGSPICE file created from sky130_fd_sc_lp__sdfxbp_2.ext - technology: sky130A

.subckt sky130_fd_sc_lp__sdfxbp_2 CLK D SCD SCE VGND VNB VPB VPWR Q Q_N
M1000 VGND a_2122_329# a_2097_122# VNB nshort w=420000u l=150000u
+  ad=2.1442e+12p pd=1.874e+07u as=8.82e+10p ps=1.26e+06u
M1001 a_1188_93# CLK VPWR VPB phighvt w=640000u l=150000u
+  ad=1.824e+11p pd=1.85e+06u as=2.7553e+12p ps=2.403e+07u
M1002 Q a_2122_329# VGND VNB nshort w=840000u l=150000u
+  ad=2.352e+11p pd=2.24e+06u as=0p ps=0u
M1003 a_332_94# SCE VGND VNB nshort w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1004 VPWR a_733_21# a_778_399# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=6.131e+11p ps=4.99e+06u
M1005 VPWR SCE a_332_94# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=2.976e+11p ps=2.21e+06u
M1006 a_268_120# D a_182_120# VNB nshort w=420000u l=150000u
+  ad=1.344e+11p pd=1.48e+06u as=2.289e+11p ps=2.77e+06u
M1007 a_2710_56# a_2122_329# VPWR VPB phighvt w=640000u l=150000u
+  ad=1.696e+11p pd=1.81e+06u as=0p ps=0u
M1008 VPWR a_2710_56# Q_N VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=3.528e+11p ps=3.08e+06u
M1009 a_204_489# SCE VPWR VPB phighvt w=640000u l=150000u
+  ad=1.344e+11p pd=1.7e+06u as=0p ps=0u
M1010 a_182_120# a_1188_93# a_733_21# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.176e+11p ps=1.4e+06u
M1011 a_2008_122# a_1188_93# a_778_399# VPB phighvt w=840000u l=150000u
+  ad=2.709e+11p pd=2.4e+06u as=0p ps=0u
M1012 Q_N a_2710_56# VGND VNB nshort w=840000u l=150000u
+  ad=2.352e+11p pd=2.24e+06u as=0p ps=0u
M1013 VGND a_733_21# a_778_399# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=2.809e+11p ps=3.18e+06u
M1014 a_182_120# D a_204_489# VPB phighvt w=640000u l=150000u
+  ad=3.325e+11p pd=3.41e+06u as=0p ps=0u
M1015 a_2097_122# a_1188_93# a_2008_122# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.239e+11p ps=1.43e+06u
M1016 VGND a_1188_93# a_1102_93# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1017 a_733_21# a_1102_93# a_1060_119# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1018 a_1188_93# CLK VGND VNB nshort w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1019 VGND a_2122_329# Q VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_182_120# SCE a_110_120# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1021 a_2008_122# a_1102_93# a_778_399# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VPWR a_2122_329# Q VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=3.528e+11p ps=3.08e+06u
M1023 VPWR SCD a_27_489# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=3.392e+11p ps=3.62e+06u
M1024 a_993_425# a_1188_93# a_733_21# VPB phighvt w=420000u l=150000u
+  ad=3.785e+11p pd=3.97e+06u as=1.176e+11p ps=1.4e+06u
M1025 a_2122_329# a_2008_122# VPWR VPB phighvt w=840000u l=150000u
+  ad=2.226e+11p pd=2.21e+06u as=0p ps=0u
M1026 VGND a_332_94# a_268_120# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 VPWR a_1188_93# a_1102_93# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=2.56e+11p ps=2.08e+06u
M1028 Q_N a_2710_56# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 a_2710_56# a_2122_329# VGND VNB nshort w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1030 VGND a_2710_56# Q_N VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_1060_119# a_778_399# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 a_2122_329# a_2008_122# VGND VNB nshort w=640000u l=150000u
+  ad=1.696e+11p pd=1.81e+06u as=0p ps=0u
M1033 a_993_425# a_778_399# VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1034 a_2116_463# a_1102_93# a_2008_122# VPB phighvt w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1035 a_110_120# SCD VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1036 VPWR a_2122_329# a_2116_463# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1037 Q a_2122_329# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1038 a_27_489# a_332_94# a_182_120# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1039 a_733_21# a_1102_93# a_182_120# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

