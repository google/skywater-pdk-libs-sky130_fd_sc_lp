* File: sky130_fd_sc_lp__nand4_2.pxi.spice
* Created: Wed Sep  2 10:05:35 2020
* 
x_PM_SKY130_FD_SC_LP__NAND4_2%D N_D_M1004_g N_D_c_77_n N_D_M1000_g N_D_M1011_g
+ N_D_c_78_n N_D_M1005_g D D N_D_c_76_n PM_SKY130_FD_SC_LP__NAND4_2%D
x_PM_SKY130_FD_SC_LP__NAND4_2%C N_C_c_114_n N_C_M1009_g N_C_M1002_g N_C_c_116_n
+ N_C_M1014_g N_C_M1010_g C C N_C_c_119_n PM_SKY130_FD_SC_LP__NAND4_2%C
x_PM_SKY130_FD_SC_LP__NAND4_2%B N_B_M1003_g N_B_c_167_n N_B_c_168_n N_B_M1007_g
+ N_B_M1015_g N_B_M1013_g B N_B_c_171_n N_B_c_175_n
+ PM_SKY130_FD_SC_LP__NAND4_2%B
x_PM_SKY130_FD_SC_LP__NAND4_2%A N_A_M1001_g N_A_M1006_g N_A_M1008_g N_A_M1012_g
+ A A A N_A_c_226_n PM_SKY130_FD_SC_LP__NAND4_2%A
x_PM_SKY130_FD_SC_LP__NAND4_2%VPWR N_VPWR_M1000_d N_VPWR_M1005_d N_VPWR_M1010_d
+ N_VPWR_M1015_s N_VPWR_M1008_d N_VPWR_c_268_n N_VPWR_c_269_n N_VPWR_c_270_n
+ N_VPWR_c_271_n N_VPWR_c_272_n N_VPWR_c_273_n N_VPWR_c_274_n N_VPWR_c_275_n
+ N_VPWR_c_276_n N_VPWR_c_277_n N_VPWR_c_278_n N_VPWR_c_279_n N_VPWR_c_280_n
+ N_VPWR_c_281_n VPWR N_VPWR_c_282_n N_VPWR_c_267_n
+ PM_SKY130_FD_SC_LP__NAND4_2%VPWR
x_PM_SKY130_FD_SC_LP__NAND4_2%Y N_Y_M1006_s N_Y_M1000_s N_Y_M1002_s N_Y_M1003_d
+ N_Y_M1001_s N_Y_c_404_n N_Y_c_345_n N_Y_c_346_n N_Y_c_408_n N_Y_c_365_n
+ N_Y_c_341_n N_Y_c_342_n N_Y_c_371_n N_Y_c_343_n N_Y_c_394_n N_Y_c_379_n
+ N_Y_c_380_n Y PM_SKY130_FD_SC_LP__NAND4_2%Y
x_PM_SKY130_FD_SC_LP__NAND4_2%A_69_47# N_A_69_47#_M1004_d N_A_69_47#_M1011_d
+ N_A_69_47#_M1014_s N_A_69_47#_c_433_n N_A_69_47#_c_434_n N_A_69_47#_c_435_n
+ N_A_69_47#_c_454_p N_A_69_47#_c_443_n N_A_69_47#_c_436_n
+ PM_SKY130_FD_SC_LP__NAND4_2%A_69_47#
x_PM_SKY130_FD_SC_LP__NAND4_2%VGND N_VGND_M1004_s N_VGND_c_468_n N_VGND_c_469_n
+ N_VGND_c_470_n VGND N_VGND_c_471_n N_VGND_c_472_n
+ PM_SKY130_FD_SC_LP__NAND4_2%VGND
x_PM_SKY130_FD_SC_LP__NAND4_2%A_330_47# N_A_330_47#_M1009_d N_A_330_47#_M1007_s
+ N_A_330_47#_c_512_n N_A_330_47#_c_516_n PM_SKY130_FD_SC_LP__NAND4_2%A_330_47#
x_PM_SKY130_FD_SC_LP__NAND4_2%A_523_67# N_A_523_67#_M1007_d N_A_523_67#_M1013_d
+ N_A_523_67#_M1012_d N_A_523_67#_c_537_n N_A_523_67#_c_550_n
+ N_A_523_67#_c_538_n N_A_523_67#_c_539_n N_A_523_67#_c_540_n
+ PM_SKY130_FD_SC_LP__NAND4_2%A_523_67#
cc_1 VNB N_D_M1004_g 0.0329127f $X=-0.19 $Y=-0.245 $X2=0.685 $Y2=0.655
cc_2 VNB N_D_M1011_g 0.0243008f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=0.655
cc_3 VNB D 0.0119013f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_4 VNB N_D_c_76_n 0.0483006f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.535
cc_5 VNB N_C_c_114_n 0.01661f $X=-0.19 $Y=-0.245 $X2=0.685 $Y2=1.345
cc_6 VNB N_C_M1002_g 0.0165887f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=2.465
cc_7 VNB N_C_c_116_n 0.0198092f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.345
cc_8 VNB N_C_M1010_g 0.00718714f $X=-0.19 $Y=-0.245 $X2=1.285 $Y2=2.465
cc_9 VNB C 0.0117221f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.95
cc_10 VNB N_C_c_119_n 0.0554562f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.51
cc_11 VNB N_B_M1003_g 0.00709603f $X=-0.19 $Y=-0.245 $X2=0.685 $Y2=0.655
cc_12 VNB N_B_c_167_n 0.0116644f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=1.725
cc_13 VNB N_B_c_168_n 0.00847204f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=2.465
cc_14 VNB N_B_M1007_g 0.0225578f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=0.655
cc_15 VNB N_B_M1013_g 0.0188568f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_B_c_171_n 0.0309136f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=1.535
cc_17 VNB N_A_M1006_g 0.018874f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=2.465
cc_18 VNB N_A_M1012_g 0.0257996f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_19 VNB A 0.0201883f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_c_226_n 0.0419958f $X=-0.19 $Y=-0.245 $X2=0.715 $Y2=2.035
cc_21 VNB N_VPWR_c_267_n 0.203486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_Y_c_341_n 0.00769669f $X=-0.19 $Y=-0.245 $X2=0.715 $Y2=1.507
cc_23 VNB N_Y_c_342_n 0.00321513f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.507
cc_24 VNB N_Y_c_343_n 0.00852371f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB Y 0.00464141f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_69_47#_c_433_n 0.0277218f $X=-0.19 $Y=-0.245 $X2=1.285 $Y2=1.725
cc_27 VNB N_A_69_47#_c_434_n 0.00789982f $X=-0.19 $Y=-0.245 $X2=1.285 $Y2=2.465
cc_28 VNB N_A_69_47#_c_435_n 0.0141668f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_29 VNB N_A_69_47#_c_436_n 0.00335617f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.51
cc_30 VNB N_VGND_c_468_n 4.89148e-19 $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=2.465
cc_31 VNB N_VGND_c_469_n 0.0220585f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=0.655
cc_32 VNB N_VGND_c_470_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=0.655
cc_33 VNB N_VGND_c_471_n 0.0882887f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.535
cc_34 VNB N_VGND_c_472_n 0.272818f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.51
cc_35 VNB N_A_330_47#_c_512_n 0.0117349f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=0.655
cc_36 VNB N_A_523_67#_c_537_n 0.00749711f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=0.655
cc_37 VNB N_A_523_67#_c_538_n 0.0119396f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_523_67#_c_539_n 0.0319139f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.51
cc_39 VNB N_A_523_67#_c_540_n 0.00136752f $X=-0.19 $Y=-0.245 $X2=0.855 $Y2=1.535
cc_40 VPB N_D_c_77_n 0.0191474f $X=-0.19 $Y=1.655 $X2=0.855 $Y2=1.725
cc_41 VPB N_D_c_78_n 0.0153475f $X=-0.19 $Y=1.655 $X2=1.285 $Y2=1.725
cc_42 VPB D 0.00383842f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_43 VPB N_D_c_76_n 0.0200777f $X=-0.19 $Y=1.655 $X2=1.115 $Y2=1.535
cc_44 VPB N_C_M1002_g 0.0190638f $X=-0.19 $Y=1.655 $X2=0.855 $Y2=2.465
cc_45 VPB N_C_M1010_g 0.0192499f $X=-0.19 $Y=1.655 $X2=1.285 $Y2=2.465
cc_46 VPB N_B_M1003_g 0.0192456f $X=-0.19 $Y=1.655 $X2=0.685 $Y2=0.655
cc_47 VPB N_B_M1015_g 0.0205683f $X=-0.19 $Y=1.655 $X2=1.285 $Y2=2.465
cc_48 VPB N_B_c_171_n 0.0106615f $X=-0.19 $Y=1.655 $X2=0.855 $Y2=1.535
cc_49 VPB N_B_c_175_n 0.00258925f $X=-0.19 $Y=1.655 $X2=1.115 $Y2=1.535
cc_50 VPB N_A_M1001_g 0.02062f $X=-0.19 $Y=1.655 $X2=0.685 $Y2=0.655
cc_51 VPB N_A_M1008_g 0.0235869f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_52 VPB A 0.0186885f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_53 VPB N_A_c_226_n 0.00762096f $X=-0.19 $Y=1.655 $X2=0.715 $Y2=2.035
cc_54 VPB N_VPWR_c_268_n 0.0282008f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_55 VPB N_VPWR_c_269_n 0.042045f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=1.535
cc_56 VPB N_VPWR_c_270_n 3.16879e-19 $X=-0.19 $Y=1.655 $X2=0.855 $Y2=1.535
cc_57 VPB N_VPWR_c_271_n 0.0049741f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_58 VPB N_VPWR_c_272_n 0.00509424f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_59 VPB N_VPWR_c_273_n 0.0144866f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_60 VPB N_VPWR_c_274_n 0.0483836f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_61 VPB N_VPWR_c_275_n 0.0140974f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_62 VPB N_VPWR_c_276_n 0.0129398f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_63 VPB N_VPWR_c_277_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_64 VPB N_VPWR_c_278_n 0.0154998f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_279_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_280_n 0.0190096f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_67 VPB N_VPWR_c_281_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_282_n 0.0171783f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_69 VPB N_VPWR_c_267_n 0.0507015f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_70 VPB N_Y_c_345_n 0.00635217f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=1.51
cc_71 VPB N_Y_c_346_n 0.00291477f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=1.51
cc_72 VPB N_Y_c_343_n 0.00429918f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_73 N_D_M1011_g N_C_c_114_n 0.0205675f $X=1.115 $Y=0.655 $X2=-0.19 $Y2=-0.245
cc_74 N_D_M1011_g N_C_M1002_g 0.00758172f $X=1.115 $Y=0.655 $X2=0 $Y2=0
cc_75 N_D_c_76_n N_C_M1002_g 0.0255988f $X=1.115 $Y=1.535 $X2=0 $Y2=0
cc_76 N_D_M1011_g C 0.00319828f $X=1.115 $Y=0.655 $X2=0 $Y2=0
cc_77 D N_VPWR_M1000_d 0.00412896f $X=0.635 $Y=1.58 $X2=-0.19 $Y2=-0.245
cc_78 N_D_c_77_n N_VPWR_c_268_n 0.00453612f $X=0.855 $Y=1.725 $X2=0 $Y2=0
cc_79 D N_VPWR_c_268_n 0.0234052f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_80 N_D_c_77_n N_VPWR_c_269_n 0.0123252f $X=0.855 $Y=1.725 $X2=0 $Y2=0
cc_81 N_D_c_77_n N_VPWR_c_270_n 7.27171e-19 $X=0.855 $Y=1.725 $X2=0 $Y2=0
cc_82 N_D_c_78_n N_VPWR_c_270_n 0.0141832f $X=1.285 $Y=1.725 $X2=0 $Y2=0
cc_83 N_D_c_77_n N_VPWR_c_275_n 0.00372254f $X=0.855 $Y=1.725 $X2=0 $Y2=0
cc_84 N_D_c_78_n N_VPWR_c_275_n 6.83371e-19 $X=1.285 $Y=1.725 $X2=0 $Y2=0
cc_85 D N_VPWR_c_275_n 0.0125738f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_86 N_D_c_76_n N_VPWR_c_275_n 0.00181406f $X=1.115 $Y=1.535 $X2=0 $Y2=0
cc_87 N_D_c_77_n N_VPWR_c_276_n 0.00486043f $X=0.855 $Y=1.725 $X2=0 $Y2=0
cc_88 N_D_c_78_n N_VPWR_c_276_n 0.00486043f $X=1.285 $Y=1.725 $X2=0 $Y2=0
cc_89 N_D_c_77_n N_VPWR_c_267_n 0.00824727f $X=0.855 $Y=1.725 $X2=0 $Y2=0
cc_90 N_D_c_78_n N_VPWR_c_267_n 0.00824727f $X=1.285 $Y=1.725 $X2=0 $Y2=0
cc_91 N_D_c_78_n N_Y_c_345_n 0.013904f $X=1.285 $Y=1.725 $X2=0 $Y2=0
cc_92 N_D_c_77_n N_Y_c_346_n 6.55961e-19 $X=0.855 $Y=1.725 $X2=0 $Y2=0
cc_93 D N_Y_c_346_n 0.0095228f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_94 N_D_c_76_n N_Y_c_346_n 0.00400907f $X=1.115 $Y=1.535 $X2=0 $Y2=0
cc_95 N_D_M1004_g N_A_69_47#_c_434_n 0.0139356f $X=0.685 $Y=0.655 $X2=0 $Y2=0
cc_96 N_D_M1011_g N_A_69_47#_c_434_n 0.0149225f $X=1.115 $Y=0.655 $X2=0 $Y2=0
cc_97 D N_A_69_47#_c_434_n 0.0195314f $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_98 N_D_c_76_n N_A_69_47#_c_434_n 0.00844534f $X=1.115 $Y=1.535 $X2=0 $Y2=0
cc_99 D N_A_69_47#_c_435_n 7.78284e-19 $X=0.635 $Y=1.58 $X2=0 $Y2=0
cc_100 N_D_M1004_g N_VGND_c_468_n 0.0116286f $X=0.685 $Y=0.655 $X2=0 $Y2=0
cc_101 N_D_M1011_g N_VGND_c_468_n 0.0110862f $X=1.115 $Y=0.655 $X2=0 $Y2=0
cc_102 N_D_M1004_g N_VGND_c_469_n 0.00486043f $X=0.685 $Y=0.655 $X2=0 $Y2=0
cc_103 N_D_M1011_g N_VGND_c_471_n 0.00486043f $X=1.115 $Y=0.655 $X2=0 $Y2=0
cc_104 N_D_M1004_g N_VGND_c_472_n 0.0093271f $X=0.685 $Y=0.655 $X2=0 $Y2=0
cc_105 N_D_M1011_g N_VGND_c_472_n 0.00834351f $X=1.115 $Y=0.655 $X2=0 $Y2=0
cc_106 N_C_M1010_g N_B_M1003_g 0.0304718f $X=2.145 $Y=2.465 $X2=0 $Y2=0
cc_107 N_C_c_119_n N_B_c_168_n 0.00870365f $X=2.145 $Y=1.335 $X2=0 $Y2=0
cc_108 N_C_c_119_n N_B_M1007_g 0.00224572f $X=2.145 $Y=1.335 $X2=0 $Y2=0
cc_109 N_C_M1002_g N_VPWR_c_270_n 0.0142862f $X=1.715 $Y=2.465 $X2=0 $Y2=0
cc_110 N_C_M1010_g N_VPWR_c_270_n 7.45395e-19 $X=2.145 $Y=2.465 $X2=0 $Y2=0
cc_111 N_C_M1010_g N_VPWR_c_271_n 0.00272546f $X=2.145 $Y=2.465 $X2=0 $Y2=0
cc_112 N_C_M1002_g N_VPWR_c_278_n 0.00486043f $X=1.715 $Y=2.465 $X2=0 $Y2=0
cc_113 N_C_M1010_g N_VPWR_c_278_n 0.00585385f $X=2.145 $Y=2.465 $X2=0 $Y2=0
cc_114 N_C_M1002_g N_VPWR_c_267_n 0.00824727f $X=1.715 $Y=2.465 $X2=0 $Y2=0
cc_115 N_C_M1010_g N_VPWR_c_267_n 0.0107559f $X=2.145 $Y=2.465 $X2=0 $Y2=0
cc_116 N_C_M1002_g N_Y_c_345_n 0.0140082f $X=1.715 $Y=2.465 $X2=0 $Y2=0
cc_117 C N_Y_c_345_n 0.0113645f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_118 N_C_c_119_n N_Y_c_345_n 0.00321502f $X=2.145 $Y=1.335 $X2=0 $Y2=0
cc_119 N_C_c_116_n N_Y_c_342_n 0.00295673f $X=2.005 $Y=1.185 $X2=0 $Y2=0
cc_120 C N_Y_c_342_n 0.00712948f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_121 N_C_c_119_n N_Y_c_342_n 2.85736e-19 $X=2.145 $Y=1.335 $X2=0 $Y2=0
cc_122 N_C_M1002_g N_Y_c_343_n 0.00387184f $X=1.715 $Y=2.465 $X2=0 $Y2=0
cc_123 N_C_M1010_g N_Y_c_343_n 0.0249584f $X=2.145 $Y=2.465 $X2=0 $Y2=0
cc_124 C N_Y_c_343_n 0.0349885f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_125 N_C_c_119_n N_Y_c_343_n 0.00583617f $X=2.145 $Y=1.335 $X2=0 $Y2=0
cc_126 N_C_M1010_g Y 0.00190511f $X=2.145 $Y=2.465 $X2=0 $Y2=0
cc_127 C Y 0.0158361f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_128 N_C_c_119_n Y 0.00266381f $X=2.145 $Y=1.335 $X2=0 $Y2=0
cc_129 N_C_c_114_n N_A_69_47#_c_434_n 0.00465881f $X=1.575 $Y=1.185 $X2=0 $Y2=0
cc_130 N_C_c_114_n N_A_69_47#_c_443_n 0.00465062f $X=1.575 $Y=1.185 $X2=0 $Y2=0
cc_131 N_C_c_114_n N_A_69_47#_c_436_n 0.0142044f $X=1.575 $Y=1.185 $X2=0 $Y2=0
cc_132 N_C_c_116_n N_A_69_47#_c_436_n 0.0107715f $X=2.005 $Y=1.185 $X2=0 $Y2=0
cc_133 C N_A_69_47#_c_436_n 0.00100059f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_134 N_C_c_114_n N_VGND_c_468_n 0.00104858f $X=1.575 $Y=1.185 $X2=0 $Y2=0
cc_135 N_C_c_114_n N_VGND_c_471_n 0.00357877f $X=1.575 $Y=1.185 $X2=0 $Y2=0
cc_136 N_C_c_116_n N_VGND_c_471_n 0.00357877f $X=2.005 $Y=1.185 $X2=0 $Y2=0
cc_137 N_C_c_114_n N_VGND_c_472_n 0.00544745f $X=1.575 $Y=1.185 $X2=0 $Y2=0
cc_138 N_C_c_116_n N_VGND_c_472_n 0.00665089f $X=2.005 $Y=1.185 $X2=0 $Y2=0
cc_139 N_C_c_116_n N_A_330_47#_c_512_n 0.0105596f $X=2.005 $Y=1.185 $X2=0 $Y2=0
cc_140 C N_A_330_47#_c_512_n 0.019008f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_141 N_C_c_119_n N_A_330_47#_c_512_n 0.0013981f $X=2.145 $Y=1.335 $X2=0 $Y2=0
cc_142 N_C_c_114_n N_A_330_47#_c_516_n 0.00375432f $X=1.575 $Y=1.185 $X2=0 $Y2=0
cc_143 N_C_c_116_n N_A_330_47#_c_516_n 0.00496338f $X=2.005 $Y=1.185 $X2=0 $Y2=0
cc_144 C N_A_330_47#_c_516_n 0.0213806f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_145 N_C_c_119_n N_A_330_47#_c_516_n 6.92408e-19 $X=2.145 $Y=1.335 $X2=0 $Y2=0
cc_146 N_B_M1015_g N_A_M1001_g 0.0264449f $X=3.085 $Y=2.465 $X2=0 $Y2=0
cc_147 N_B_M1013_g N_A_M1006_g 0.0340606f $X=3.405 $Y=0.755 $X2=0 $Y2=0
cc_148 N_B_M1015_g A 2.29991e-19 $X=3.085 $Y=2.465 $X2=0 $Y2=0
cc_149 N_B_c_171_n A 0.00218081f $X=3.17 $Y=1.51 $X2=0 $Y2=0
cc_150 N_B_c_175_n A 0.0275411f $X=3.17 $Y=1.51 $X2=0 $Y2=0
cc_151 N_B_c_171_n N_A_c_226_n 0.0226962f $X=3.17 $Y=1.51 $X2=0 $Y2=0
cc_152 N_B_M1003_g N_VPWR_c_271_n 0.00433557f $X=2.655 $Y=2.465 $X2=0 $Y2=0
cc_153 N_B_M1015_g N_VPWR_c_272_n 0.0118569f $X=3.085 $Y=2.465 $X2=0 $Y2=0
cc_154 N_B_M1003_g N_VPWR_c_280_n 0.00585385f $X=2.655 $Y=2.465 $X2=0 $Y2=0
cc_155 N_B_M1015_g N_VPWR_c_280_n 0.0054895f $X=3.085 $Y=2.465 $X2=0 $Y2=0
cc_156 N_B_M1003_g N_VPWR_c_267_n 0.0107286f $X=2.655 $Y=2.465 $X2=0 $Y2=0
cc_157 N_B_M1015_g N_VPWR_c_267_n 0.0105734f $X=3.085 $Y=2.465 $X2=0 $Y2=0
cc_158 N_B_M1015_g N_Y_c_365_n 0.0147237f $X=3.085 $Y=2.465 $X2=0 $Y2=0
cc_159 N_B_c_167_n N_Y_c_341_n 0.00168762f $X=2.9 $Y=1.42 $X2=0 $Y2=0
cc_160 N_B_M1007_g N_Y_c_341_n 0.0127803f $X=2.975 $Y=0.755 $X2=0 $Y2=0
cc_161 N_B_M1013_g N_Y_c_341_n 0.0135704f $X=3.405 $Y=0.755 $X2=0 $Y2=0
cc_162 N_B_c_171_n N_Y_c_341_n 0.0025327f $X=3.17 $Y=1.51 $X2=0 $Y2=0
cc_163 N_B_c_175_n N_Y_c_341_n 0.023516f $X=3.17 $Y=1.51 $X2=0 $Y2=0
cc_164 N_B_M1015_g N_Y_c_371_n 0.0121862f $X=3.085 $Y=2.465 $X2=0 $Y2=0
cc_165 N_B_c_171_n N_Y_c_371_n 0.00505882f $X=3.17 $Y=1.51 $X2=0 $Y2=0
cc_166 N_B_c_175_n N_Y_c_371_n 0.0204607f $X=3.17 $Y=1.51 $X2=0 $Y2=0
cc_167 N_B_M1003_g N_Y_c_343_n 0.0209039f $X=2.655 $Y=2.465 $X2=0 $Y2=0
cc_168 N_B_c_167_n N_Y_c_343_n 0.00352364f $X=2.9 $Y=1.42 $X2=0 $Y2=0
cc_169 N_B_M1015_g N_Y_c_343_n 0.00540097f $X=3.085 $Y=2.465 $X2=0 $Y2=0
cc_170 N_B_c_171_n N_Y_c_343_n 5.13115e-19 $X=3.17 $Y=1.51 $X2=0 $Y2=0
cc_171 N_B_c_175_n N_Y_c_343_n 0.0146651f $X=3.17 $Y=1.51 $X2=0 $Y2=0
cc_172 N_B_M1015_g N_Y_c_379_n 8.94977e-19 $X=3.085 $Y=2.465 $X2=0 $Y2=0
cc_173 N_B_M1013_g N_Y_c_380_n 8.49133e-19 $X=3.405 $Y=0.755 $X2=0 $Y2=0
cc_174 N_B_M1003_g Y 0.00291602f $X=2.655 $Y=2.465 $X2=0 $Y2=0
cc_175 N_B_c_167_n Y 0.0106165f $X=2.9 $Y=1.42 $X2=0 $Y2=0
cc_176 N_B_c_168_n Y 0.0057802f $X=2.73 $Y=1.42 $X2=0 $Y2=0
cc_177 N_B_M1007_g Y 0.00298733f $X=2.975 $Y=0.755 $X2=0 $Y2=0
cc_178 N_B_c_171_n Y 7.49744e-19 $X=3.17 $Y=1.51 $X2=0 $Y2=0
cc_179 N_B_c_175_n Y 0.0139332f $X=3.17 $Y=1.51 $X2=0 $Y2=0
cc_180 N_B_M1007_g N_A_69_47#_c_436_n 7.43698e-19 $X=2.975 $Y=0.755 $X2=0 $Y2=0
cc_181 N_B_M1007_g N_VGND_c_471_n 0.00296932f $X=2.975 $Y=0.755 $X2=0 $Y2=0
cc_182 N_B_M1013_g N_VGND_c_471_n 0.00296932f $X=3.405 $Y=0.755 $X2=0 $Y2=0
cc_183 N_B_M1007_g N_VGND_c_472_n 0.00456657f $X=2.975 $Y=0.755 $X2=0 $Y2=0
cc_184 N_B_M1013_g N_VGND_c_472_n 0.00417446f $X=3.405 $Y=0.755 $X2=0 $Y2=0
cc_185 N_B_c_168_n N_A_330_47#_c_512_n 9.8351e-19 $X=2.73 $Y=1.42 $X2=0 $Y2=0
cc_186 N_B_M1007_g N_A_330_47#_c_512_n 0.0112377f $X=2.975 $Y=0.755 $X2=0 $Y2=0
cc_187 N_B_M1013_g N_A_330_47#_c_512_n 0.00252495f $X=3.405 $Y=0.755 $X2=0 $Y2=0
cc_188 N_B_M1007_g N_A_523_67#_c_537_n 0.0120247f $X=2.975 $Y=0.755 $X2=0 $Y2=0
cc_189 N_B_M1013_g N_A_523_67#_c_537_n 0.0151128f $X=3.405 $Y=0.755 $X2=0 $Y2=0
cc_190 N_A_M1001_g N_VPWR_c_272_n 0.0103844f $X=3.765 $Y=2.465 $X2=0 $Y2=0
cc_191 N_A_M1001_g N_VPWR_c_274_n 8.53014e-19 $X=3.765 $Y=2.465 $X2=0 $Y2=0
cc_192 N_A_M1008_g N_VPWR_c_274_n 0.0206595f $X=4.195 $Y=2.465 $X2=0 $Y2=0
cc_193 A N_VPWR_c_274_n 0.025707f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_194 N_A_c_226_n N_VPWR_c_274_n 4.32447e-19 $X=4.265 $Y=1.51 $X2=0 $Y2=0
cc_195 N_A_M1001_g N_VPWR_c_282_n 0.0054895f $X=3.765 $Y=2.465 $X2=0 $Y2=0
cc_196 N_A_M1008_g N_VPWR_c_282_n 0.00486043f $X=4.195 $Y=2.465 $X2=0 $Y2=0
cc_197 N_A_M1001_g N_VPWR_c_267_n 0.0105734f $X=3.765 $Y=2.465 $X2=0 $Y2=0
cc_198 N_A_M1008_g N_VPWR_c_267_n 0.00824727f $X=4.195 $Y=2.465 $X2=0 $Y2=0
cc_199 N_A_M1001_g N_Y_c_365_n 8.93495e-19 $X=3.765 $Y=2.465 $X2=0 $Y2=0
cc_200 N_A_M1006_g N_Y_c_341_n 0.0107689f $X=3.835 $Y=0.755 $X2=0 $Y2=0
cc_201 N_A_M1012_g N_Y_c_341_n 0.00482563f $X=4.265 $Y=0.755 $X2=0 $Y2=0
cc_202 A N_Y_c_341_n 0.053895f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_203 N_A_c_226_n N_Y_c_341_n 0.0048565f $X=4.265 $Y=1.51 $X2=0 $Y2=0
cc_204 N_A_M1001_g N_Y_c_371_n 0.0121913f $X=3.765 $Y=2.465 $X2=0 $Y2=0
cc_205 A N_Y_c_371_n 0.021215f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_206 N_A_M1001_g N_Y_c_394_n 7.32094e-19 $X=3.765 $Y=2.465 $X2=0 $Y2=0
cc_207 A N_Y_c_394_n 0.019204f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_208 N_A_c_226_n N_Y_c_394_n 6.47713e-19 $X=4.265 $Y=1.51 $X2=0 $Y2=0
cc_209 N_A_M1001_g N_Y_c_379_n 0.0139882f $X=3.765 $Y=2.465 $X2=0 $Y2=0
cc_210 N_A_M1006_g N_Y_c_380_n 0.00653973f $X=3.835 $Y=0.755 $X2=0 $Y2=0
cc_211 N_A_M1012_g N_Y_c_380_n 0.0054303f $X=4.265 $Y=0.755 $X2=0 $Y2=0
cc_212 N_A_M1006_g N_VGND_c_471_n 0.00296932f $X=3.835 $Y=0.755 $X2=0 $Y2=0
cc_213 N_A_M1012_g N_VGND_c_471_n 0.00296932f $X=4.265 $Y=0.755 $X2=0 $Y2=0
cc_214 N_A_M1006_g N_VGND_c_472_n 0.00417446f $X=3.835 $Y=0.755 $X2=0 $Y2=0
cc_215 N_A_M1012_g N_VGND_c_472_n 0.00446962f $X=4.265 $Y=0.755 $X2=0 $Y2=0
cc_216 N_A_M1006_g N_A_523_67#_c_538_n 0.0111282f $X=3.835 $Y=0.755 $X2=0 $Y2=0
cc_217 N_A_M1012_g N_A_523_67#_c_538_n 0.0127094f $X=4.265 $Y=0.755 $X2=0 $Y2=0
cc_218 N_A_M1012_g N_A_523_67#_c_539_n 0.00354524f $X=4.265 $Y=0.755 $X2=0 $Y2=0
cc_219 A N_A_523_67#_c_539_n 0.0184375f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_220 N_VPWR_c_267_n N_Y_M1000_s 0.00536646f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_221 N_VPWR_c_267_n N_Y_M1002_s 0.00571434f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_222 N_VPWR_c_267_n N_Y_M1003_d 0.00258346f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_223 N_VPWR_c_267_n N_Y_M1001_s 0.00380103f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_224 N_VPWR_c_276_n N_Y_c_404_n 0.0124525f $X=1.335 $Y=3.33 $X2=0 $Y2=0
cc_225 N_VPWR_c_267_n N_Y_c_404_n 0.00730901f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_226 N_VPWR_M1005_d N_Y_c_345_n 0.00176461f $X=1.36 $Y=1.835 $X2=0 $Y2=0
cc_227 N_VPWR_c_270_n N_Y_c_345_n 0.0170777f $X=1.5 $Y=2.18 $X2=0 $Y2=0
cc_228 N_VPWR_c_278_n N_Y_c_408_n 0.0120977f $X=2.24 $Y=3.33 $X2=0 $Y2=0
cc_229 N_VPWR_c_267_n N_Y_c_408_n 0.00691495f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_230 N_VPWR_c_272_n N_Y_c_365_n 0.0505935f $X=3.425 $Y=2.38 $X2=0 $Y2=0
cc_231 N_VPWR_c_280_n N_Y_c_365_n 0.0169299f $X=3.26 $Y=3.33 $X2=0 $Y2=0
cc_232 N_VPWR_c_267_n N_Y_c_365_n 0.0112082f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_233 N_VPWR_M1015_s N_Y_c_371_n 0.0134234f $X=3.16 $Y=1.835 $X2=0 $Y2=0
cc_234 N_VPWR_c_272_n N_Y_c_371_n 0.0266856f $X=3.425 $Y=2.38 $X2=0 $Y2=0
cc_235 N_VPWR_M1010_d N_Y_c_343_n 0.00269699f $X=2.22 $Y=1.835 $X2=0 $Y2=0
cc_236 N_VPWR_c_271_n N_Y_c_343_n 0.0216883f $X=2.405 $Y=2.38 $X2=0 $Y2=0
cc_237 N_VPWR_c_272_n N_Y_c_379_n 0.0501328f $X=3.425 $Y=2.38 $X2=0 $Y2=0
cc_238 N_VPWR_c_282_n N_Y_c_379_n 0.015688f $X=4.245 $Y=3.33 $X2=0 $Y2=0
cc_239 N_VPWR_c_267_n N_Y_c_379_n 0.00984745f $X=4.56 $Y=3.33 $X2=0 $Y2=0
cc_240 N_VPWR_c_268_n N_A_69_47#_c_435_n 0.00538344f $X=0.3 $Y=1.98 $X2=0 $Y2=0
cc_241 N_Y_c_345_n N_A_69_47#_c_434_n 0.00780745f $X=1.835 $Y=1.84 $X2=0 $Y2=0
cc_242 N_Y_c_346_n N_A_69_47#_c_434_n 0.00615998f $X=1.165 $Y=1.84 $X2=0 $Y2=0
cc_243 N_Y_c_341_n N_A_330_47#_M1007_s 0.00176891f $X=3.885 $Y=1.16 $X2=0 $Y2=0
cc_244 N_Y_c_341_n N_A_330_47#_c_512_n 0.0246032f $X=3.885 $Y=1.16 $X2=0 $Y2=0
cc_245 N_Y_c_342_n N_A_330_47#_c_512_n 0.0278209f $X=2.835 $Y=1.16 $X2=0 $Y2=0
cc_246 N_Y_c_342_n N_A_523_67#_M1007_d 0.00296362f $X=2.835 $Y=1.16 $X2=-0.19
+ $Y2=-0.245
cc_247 N_Y_c_341_n N_A_523_67#_M1013_d 0.00176461f $X=3.885 $Y=1.16 $X2=0 $Y2=0
cc_248 N_Y_c_341_n N_A_523_67#_c_537_n 0.00348248f $X=3.885 $Y=1.16 $X2=0 $Y2=0
cc_249 N_Y_c_341_n N_A_523_67#_c_550_n 0.0134558f $X=3.885 $Y=1.16 $X2=0 $Y2=0
cc_250 N_Y_M1006_s N_A_523_67#_c_538_n 0.00176461f $X=3.91 $Y=0.335 $X2=0 $Y2=0
cc_251 N_Y_c_341_n N_A_523_67#_c_538_n 0.00275981f $X=3.885 $Y=1.16 $X2=0 $Y2=0
cc_252 N_Y_c_380_n N_A_523_67#_c_538_n 0.0159249f $X=4.05 $Y=0.68 $X2=0 $Y2=0
cc_253 N_Y_c_341_n N_A_523_67#_c_539_n 0.00582057f $X=3.885 $Y=1.16 $X2=0 $Y2=0
cc_254 N_A_69_47#_c_434_n N_VGND_M1004_s 0.00180746f $X=1.235 $Y=1.07 $X2=-0.19
+ $Y2=-0.245
cc_255 N_A_69_47#_c_434_n N_VGND_c_468_n 0.0163515f $X=1.235 $Y=1.07 $X2=0 $Y2=0
cc_256 N_A_69_47#_c_433_n N_VGND_c_469_n 0.0178111f $X=0.47 $Y=0.42 $X2=0 $Y2=0
cc_257 N_A_69_47#_c_454_p N_VGND_c_471_n 0.0122383f $X=1.325 $Y=0.545 $X2=0
+ $Y2=0
cc_258 N_A_69_47#_c_436_n N_VGND_c_471_n 0.0561763f $X=2.22 $Y=0.41 $X2=0 $Y2=0
cc_259 N_A_69_47#_M1004_d N_VGND_c_472_n 0.00371702f $X=0.345 $Y=0.235 $X2=0
+ $Y2=0
cc_260 N_A_69_47#_M1011_d N_VGND_c_472_n 0.00400755f $X=1.19 $Y=0.235 $X2=0
+ $Y2=0
cc_261 N_A_69_47#_M1014_s N_VGND_c_472_n 0.00215176f $X=2.08 $Y=0.235 $X2=0
+ $Y2=0
cc_262 N_A_69_47#_c_433_n N_VGND_c_472_n 0.0100304f $X=0.47 $Y=0.42 $X2=0 $Y2=0
cc_263 N_A_69_47#_c_454_p N_VGND_c_472_n 0.00699798f $X=1.325 $Y=0.545 $X2=0
+ $Y2=0
cc_264 N_A_69_47#_c_436_n N_VGND_c_472_n 0.0353857f $X=2.22 $Y=0.41 $X2=0 $Y2=0
cc_265 N_A_69_47#_c_436_n N_A_330_47#_M1009_d 0.0032998f $X=2.22 $Y=0.41
+ $X2=-0.19 $Y2=-0.245
cc_266 N_A_69_47#_M1014_s N_A_330_47#_c_512_n 0.00563706f $X=2.08 $Y=0.235 $X2=0
+ $Y2=0
cc_267 N_A_69_47#_c_434_n N_A_330_47#_c_516_n 6.33961e-19 $X=1.235 $Y=1.07 $X2=0
+ $Y2=0
cc_268 N_A_69_47#_c_443_n N_A_330_47#_c_516_n 0.0176879f $X=1.33 $Y=0.93 $X2=0
+ $Y2=0
cc_269 N_A_69_47#_c_436_n N_A_330_47#_c_516_n 0.0427735f $X=2.22 $Y=0.41 $X2=0
+ $Y2=0
cc_270 N_A_69_47#_c_436_n N_A_523_67#_c_537_n 0.0232308f $X=2.22 $Y=0.41 $X2=0
+ $Y2=0
cc_271 N_VGND_c_472_n N_A_330_47#_M1009_d 0.00225186f $X=4.56 $Y=0 $X2=-0.19
+ $Y2=-0.245
cc_272 N_VGND_c_471_n N_A_330_47#_c_512_n 0.00328236f $X=4.56 $Y=0 $X2=0 $Y2=0
cc_273 N_VGND_c_472_n N_A_330_47#_c_516_n 0.00824483f $X=4.56 $Y=0 $X2=0 $Y2=0
cc_274 N_VGND_c_471_n N_A_523_67#_c_537_n 0.061227f $X=4.56 $Y=0 $X2=0 $Y2=0
cc_275 N_VGND_c_472_n N_A_523_67#_c_537_n 0.034007f $X=4.56 $Y=0 $X2=0 $Y2=0
cc_276 N_VGND_c_471_n N_A_523_67#_c_538_n 0.0608672f $X=4.56 $Y=0 $X2=0 $Y2=0
cc_277 N_VGND_c_472_n N_A_523_67#_c_538_n 0.0339255f $X=4.56 $Y=0 $X2=0 $Y2=0
cc_278 N_VGND_c_471_n N_A_523_67#_c_540_n 0.0135745f $X=4.56 $Y=0 $X2=0 $Y2=0
cc_279 N_VGND_c_472_n N_A_523_67#_c_540_n 0.00737808f $X=4.56 $Y=0 $X2=0 $Y2=0
cc_280 N_A_330_47#_c_512_n N_A_523_67#_M1007_d 0.00557614f $X=3.19 $Y=0.81
+ $X2=-0.19 $Y2=-0.245
cc_281 N_A_330_47#_M1007_s N_A_523_67#_c_537_n 0.00179825f $X=3.05 $Y=0.335
+ $X2=0 $Y2=0
cc_282 N_A_330_47#_c_512_n N_A_523_67#_c_537_n 0.0423195f $X=3.19 $Y=0.81 $X2=0
+ $Y2=0
