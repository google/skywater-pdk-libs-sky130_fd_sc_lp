* File: sky130_fd_sc_lp__a32o_m.spice
* Created: Fri Aug 28 10:01:23 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__a32o_m.pex.spice"
.subckt sky130_fd_sc_lp__a32o_m  VNB VPB A3 A2 A1 B1 B2 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* B2	B2
* B1	B1
* A1	A1
* A2	A2
* A3	A3
* VPB	VPB
* VNB	VNB
MM1001 N_VGND_M1001_d N_A_84_153#_M1001_g N_X_M1001_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0819 AS=0.1197 PD=0.81 PS=1.41 NRD=0 NRS=5.712 M=1 R=2.8 SA=75000.2
+ SB=75002.5 A=0.063 P=1.14 MULT=1
MM1003 A_228_47# N_A3_M1003_g N_VGND_M1001_d VNB NSHORT L=0.15 W=0.42 AD=0.0441
+ AS=0.0819 PD=0.63 PS=0.81 NRD=14.28 NRS=31.428 M=1 R=2.8 SA=75000.7 SB=75002
+ A=0.063 P=1.14 MULT=1
MM1000 A_300_47# N_A2_M1000_g A_228_47# VNB NSHORT L=0.15 W=0.42 AD=0.0819
+ AS=0.0441 PD=0.81 PS=0.63 NRD=39.996 NRS=14.28 M=1 R=2.8 SA=75001.1 SB=75001.6
+ A=0.063 P=1.14 MULT=1
MM1007 N_A_84_153#_M1007_d N_A1_M1007_g A_300_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.0819 AS=0.0819 PD=0.81 PS=0.81 NRD=31.428 NRS=39.996 M=1 R=2.8 SA=75001.6
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1009 A_516_47# N_B1_M1009_g N_A_84_153#_M1007_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0819 PD=0.63 PS=0.81 NRD=14.28 NRS=0 M=1 R=2.8 SA=75002.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1010 N_VGND_M1010_d N_B2_M1010_g A_516_47# VNB NSHORT L=0.15 W=0.42 AD=0.1113
+ AS=0.0441 PD=1.37 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75002.6 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1006 N_VPWR_M1006_d N_A_84_153#_M1006_g N_X_M1006_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0756 AS=0.1113 PD=0.78 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.4 A=0.063 P=1.14 MULT=1
MM1004 N_A_228_385#_M1004_d N_A3_M1004_g N_VPWR_M1006_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0588 AS=0.0756 PD=0.7 PS=0.78 NRD=0 NRS=37.5088 M=1 R=2.8
+ SA=75000.7 SB=75001.9 A=0.063 P=1.14 MULT=1
MM1011 N_VPWR_M1011_d N_A2_M1011_g N_A_228_385#_M1004_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.1
+ SB=75001.5 A=0.063 P=1.14 MULT=1
MM1005 N_A_228_385#_M1005_d N_A1_M1005_g N_VPWR_M1011_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.6
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1002 N_A_84_153#_M1002_d N_B1_M1002_g N_A_228_385#_M1005_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75002
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1008 N_A_228_385#_M1008_d N_B2_M1008_g N_A_84_153#_M1002_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1197 AS=0.0588 PD=1.41 PS=0.7 NRD=9.3772 NRS=0 M=1 R=2.8
+ SA=75002.4 SB=75000.2 A=0.063 P=1.14 MULT=1
DX12_noxref VNB VPB NWDIODE A=6.9751 P=11.21
*
.include "sky130_fd_sc_lp__a32o_m.pxi.spice"
*
.ends
*
*
