* File: sky130_fd_sc_lp__o21bai_m.pex.spice
* Created: Fri Aug 28 11:07:08 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O21BAI_M%B1_N 3 6 9 10 11 12 13 17
c36 9 0 1.84066e-19 $X=0.59 $Y=0.84
r37 17 18 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.59
+ $Y=1.005 $X2=0.59 $Y2=1.005
r38 13 18 11.1403 $w=2.98e-07 $l=2.9e-07 $layer=LI1_cond $X=0.655 $Y=1.295
+ $X2=0.655 $Y2=1.005
r39 12 18 3.07318 $w=2.98e-07 $l=8e-08 $layer=LI1_cond $X=0.655 $Y=0.925
+ $X2=0.655 $Y2=1.005
r40 10 17 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.59 $Y=1.345
+ $X2=0.59 $Y2=1.005
r41 10 11 41.8716 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.59 $Y=1.345
+ $X2=0.59 $Y2=1.51
r42 9 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.59 $Y=0.84
+ $X2=0.59 $Y2=1.005
r43 6 11 705.053 $w=1.5e-07 $l=1.375e-06 $layer=POLY_cond $X=0.53 $Y=2.885
+ $X2=0.53 $Y2=1.51
r44 3 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.5 $Y=0.52 $X2=0.5
+ $Y2=0.84
.ends

.subckt PM_SKY130_FD_SC_LP__O21BAI_M%A_32_62# 1 2 11 13 14 15 17 19 20 21 23 26
+ 28 33 36 38 39
c59 38 0 8.56146e-20 $X=0.98 $Y=1.915
c60 11 0 1.28946e-19 $X=1.07 $Y=2.885
r61 38 39 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.98
+ $Y=1.915 $X2=0.98 $Y2=1.915
r62 33 35 8.91885 $w=2.38e-07 $l=1.65e-07 $layer=LI1_cond $X=0.27 $Y=0.495
+ $X2=0.27 $Y2=0.66
r63 29 36 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.48 $Y=1.835
+ $X2=0.315 $Y2=1.835
r64 28 38 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.895 $Y=1.835
+ $X2=0.98 $Y2=1.835
r65 28 29 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=0.895 $Y=1.835
+ $X2=0.48 $Y2=1.835
r66 24 36 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.315 $Y=1.92
+ $X2=0.315 $Y2=1.835
r67 24 26 31.4303 $w=3.28e-07 $l=9e-07 $layer=LI1_cond $X=0.315 $Y=1.92
+ $X2=0.315 $Y2=2.82
r68 23 36 3.70735 $w=2.5e-07 $l=1.18427e-07 $layer=LI1_cond $X=0.235 $Y=1.75
+ $X2=0.315 $Y2=1.835
r69 23 35 71.1123 $w=1.68e-07 $l=1.09e-06 $layer=LI1_cond $X=0.235 $Y=1.75
+ $X2=0.235 $Y2=0.66
r70 20 39 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.98 $Y=2.255
+ $X2=0.98 $Y2=1.915
r71 20 21 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.98 $Y=2.255
+ $X2=0.98 $Y2=2.42
r72 19 39 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.98 $Y=1.75
+ $X2=0.98 $Y2=1.915
r73 15 17 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.525 $Y=0.92
+ $X2=1.525 $Y2=0.6
r74 13 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.45 $Y=0.995
+ $X2=1.525 $Y2=0.92
r75 13 14 156.394 $w=1.5e-07 $l=3.05e-07 $layer=POLY_cond $X=1.45 $Y=0.995
+ $X2=1.145 $Y2=0.995
r76 11 21 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.07 $Y=2.885
+ $X2=1.07 $Y2=2.42
r77 7 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.07 $Y=1.07
+ $X2=1.145 $Y2=0.995
r78 7 19 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=1.07 $Y=1.07 $X2=1.07
+ $Y2=1.75
r79 2 26 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.19
+ $Y=2.675 $X2=0.315 $Y2=2.82
r80 1 33 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=0.16
+ $Y=0.31 $X2=0.285 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__O21BAI_M%A2 3 7 9 10 11 16
c34 3 0 8.56146e-20 $X=1.5 $Y=2.885
r35 16 19 79.7055 $w=6.05e-07 $l=5.05e-07 $layer=POLY_cond $X=1.727 $Y=1.475
+ $X2=1.727 $Y2=1.98
r36 16 18 49.6377 $w=6.05e-07 $l=1.65e-07 $layer=POLY_cond $X=1.727 $Y=1.475
+ $X2=1.727 $Y2=1.31
r37 16 17 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.68
+ $Y=1.475 $X2=1.68 $Y2=1.475
r38 10 11 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=1.68 $Y=1.665
+ $X2=1.68 $Y2=2.035
r39 10 17 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=1.68 $Y=1.665
+ $X2=1.68 $Y2=1.475
r40 9 17 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=1.68 $Y=1.295
+ $X2=1.68 $Y2=1.475
r41 7 18 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=1.955 $Y=0.6
+ $X2=1.955 $Y2=1.31
r42 3 19 464.053 $w=1.5e-07 $l=9.05e-07 $layer=POLY_cond $X=1.5 $Y=2.885 $X2=1.5
+ $Y2=1.98
.ends

.subckt PM_SKY130_FD_SC_LP__O21BAI_M%A1 3 5 6 9 13 14 15 16 17 23
r31 23 24 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.475
+ $Y=1.74 $X2=2.475 $Y2=1.74
r32 16 17 12.7285 $w=3.33e-07 $l=3.7e-07 $layer=LI1_cond $X=2.557 $Y=2.035
+ $X2=2.557 $Y2=2.405
r33 16 24 10.1484 $w=3.33e-07 $l=2.95e-07 $layer=LI1_cond $X=2.557 $Y=2.035
+ $X2=2.557 $Y2=1.74
r34 15 24 2.5801 $w=3.33e-07 $l=7.5e-08 $layer=LI1_cond $X=2.557 $Y=1.665
+ $X2=2.557 $Y2=1.74
r35 14 15 12.7285 $w=3.33e-07 $l=3.7e-07 $layer=LI1_cond $X=2.557 $Y=1.295
+ $X2=2.557 $Y2=1.665
r36 13 23 83.9334 $w=3.3e-07 $l=4.8e-07 $layer=POLY_cond $X=2.475 $Y=2.22
+ $X2=2.475 $Y2=1.74
r37 12 23 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.475 $Y=1.575
+ $X2=2.475 $Y2=1.74
r38 9 12 499.947 $w=1.5e-07 $l=9.75e-07 $layer=POLY_cond $X=2.385 $Y=0.6
+ $X2=2.385 $Y2=1.575
r39 5 13 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=2.31 $Y=2.295
+ $X2=2.475 $Y2=2.22
r40 5 6 192.287 $w=1.5e-07 $l=3.75e-07 $layer=POLY_cond $X=2.31 $Y=2.295
+ $X2=1.935 $Y2=2.295
r41 1 6 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.86 $Y=2.37
+ $X2=1.935 $Y2=2.295
r42 1 3 264.074 $w=1.5e-07 $l=5.15e-07 $layer=POLY_cond $X=1.86 $Y=2.37 $X2=1.86
+ $Y2=2.885
.ends

.subckt PM_SKY130_FD_SC_LP__O21BAI_M%VPWR 1 2 11 15 18 19 20 27 28 31
r30 31 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r31 27 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r32 25 28 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r33 24 25 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r34 22 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.99 $Y=3.33
+ $X2=0.825 $Y2=3.33
r35 22 24 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=0.99 $Y=3.33 $X2=1.68
+ $Y2=3.33
r36 20 25 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=1.68 $Y2=3.33
r37 20 32 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=0.72 $Y2=3.33
r38 18 24 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=1.97 $Y=3.33
+ $X2=1.68 $Y2=3.33
r39 18 19 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.97 $Y=3.33
+ $X2=2.075 $Y2=3.33
r40 17 27 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=2.18 $Y=3.33
+ $X2=2.64 $Y2=3.33
r41 17 19 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=2.18 $Y=3.33
+ $X2=2.075 $Y2=3.33
r42 13 19 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=2.075 $Y=3.245
+ $X2=2.075 $Y2=3.33
r43 13 15 14.5238 $w=2.08e-07 $l=2.75e-07 $layer=LI1_cond $X=2.075 $Y=3.245
+ $X2=2.075 $Y2=2.97
r44 9 31 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.825 $Y=3.245
+ $X2=0.825 $Y2=3.33
r45 9 11 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.825 $Y=3.245
+ $X2=0.825 $Y2=2.95
r46 2 15 600 $w=1.7e-07 $l=3.58225e-07 $layer=licon1_PDIFF $count=1 $X=1.935
+ $Y=2.675 $X2=2.075 $Y2=2.97
r47 1 11 600 $w=1.7e-07 $l=3.68951e-07 $layer=licon1_PDIFF $count=1 $X=0.605
+ $Y=2.675 $X2=0.825 $Y2=2.95
.ends

.subckt PM_SKY130_FD_SC_LP__O21BAI_M%Y 1 2 8 10 13 14
c31 14 0 1.28946e-19 $X=1.68 $Y=2.775
c32 8 0 1.84066e-19 $X=1.33 $Y=2.32
r33 14 22 1.52818 $w=4.79e-07 $l=6e-08 $layer=LI1_cond $X=1.472 $Y=2.775
+ $X2=1.472 $Y2=2.835
r34 13 14 9.4238 $w=4.79e-07 $l=3.7e-07 $layer=LI1_cond $X=1.472 $Y=2.405
+ $X2=1.472 $Y2=2.775
r35 10 12 9.14916 $w=2.08e-07 $l=1.65e-07 $layer=LI1_cond $X=1.31 $Y=0.665
+ $X2=1.31 $Y2=0.83
r36 8 13 7.54064 $w=4.79e-07 $l=1.79538e-07 $layer=LI1_cond $X=1.33 $Y=2.32
+ $X2=1.472 $Y2=2.405
r37 8 12 97.2086 $w=1.68e-07 $l=1.49e-06 $layer=LI1_cond $X=1.33 $Y=2.32
+ $X2=1.33 $Y2=0.83
r38 2 22 600 $w=1.7e-07 $l=2.19089e-07 $layer=licon1_PDIFF $count=1 $X=1.145
+ $Y=2.675 $X2=1.285 $Y2=2.835
r39 1 10 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=1.185
+ $Y=0.39 $X2=1.31 $Y2=0.665
.ends

.subckt PM_SKY130_FD_SC_LP__O21BAI_M%VGND 1 2 9 13 15 17 22 29 30 33 36
r34 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r35 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r36 30 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=2.16
+ $Y2=0
r37 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r38 27 36 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=2.275 $Y=0 $X2=2.17
+ $Y2=0
r39 27 29 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=2.275 $Y=0 $X2=2.64
+ $Y2=0
r40 26 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r41 25 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r42 23 33 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=0.82 $Y=0 $X2=0.715
+ $Y2=0
r43 23 25 56.107 $w=1.68e-07 $l=8.6e-07 $layer=LI1_cond $X=0.82 $Y=0 $X2=1.68
+ $Y2=0
r44 22 36 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=2.065 $Y=0 $X2=2.17
+ $Y2=0
r45 22 25 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=2.065 $Y=0 $X2=1.68
+ $Y2=0
r46 20 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r47 19 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r48 17 33 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=0.61 $Y=0 $X2=0.715
+ $Y2=0
r49 17 19 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.61 $Y=0 $X2=0.24
+ $Y2=0
r50 15 26 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=1.68
+ $Y2=0
r51 15 34 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=0.72
+ $Y2=0
r52 11 36 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=2.17 $Y=0.085
+ $X2=2.17 $Y2=0
r53 11 13 22.71 $w=2.08e-07 $l=4.3e-07 $layer=LI1_cond $X=2.17 $Y=0.085 $X2=2.17
+ $Y2=0.515
r54 7 33 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=0.715 $Y=0.085
+ $X2=0.715 $Y2=0
r55 7 9 19.5411 $w=2.08e-07 $l=3.7e-07 $layer=LI1_cond $X=0.715 $Y=0.085
+ $X2=0.715 $Y2=0.455
r56 2 13 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=2.03
+ $Y=0.39 $X2=2.17 $Y2=0.515
r57 1 9 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=0.575
+ $Y=0.31 $X2=0.715 $Y2=0.455
.ends

.subckt PM_SKY130_FD_SC_LP__O21BAI_M%A_320_78# 1 2 9 11 12 15
r23 13 15 10.2987 $w=2.08e-07 $l=1.95e-07 $layer=LI1_cond $X=2.6 $Y=0.86 $X2=2.6
+ $Y2=0.665
r24 11 13 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=2.495 $Y=0.945
+ $X2=2.6 $Y2=0.86
r25 11 12 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=2.495 $Y=0.945
+ $X2=1.845 $Y2=0.945
r26 7 12 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=1.74 $Y=0.86
+ $X2=1.845 $Y2=0.945
r27 7 9 9.24242 $w=2.08e-07 $l=1.75e-07 $layer=LI1_cond $X=1.74 $Y=0.86 $X2=1.74
+ $Y2=0.685
r28 2 15 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=2.46
+ $Y=0.39 $X2=2.6 $Y2=0.665
r29 1 9 182 $w=1.7e-07 $l=3.58225e-07 $layer=licon1_NDIFF $count=1 $X=1.6
+ $Y=0.39 $X2=1.74 $Y2=0.685
.ends

