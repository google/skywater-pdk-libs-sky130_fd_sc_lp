* File: sky130_fd_sc_lp__dfrbp_2.spice
* Created: Wed Sep  2 09:43:21 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__dfrbp_2.pex.spice"
.subckt sky130_fd_sc_lp__dfrbp_2  VNB VPB CLK D RESET_B VPWR Q_N Q VGND
* 
* VGND	VGND
* Q	Q
* Q_N	Q_N
* VPWR	VPWR
* RESET_B	RESET_B
* D	D
* CLK	CLK
* VPB	VPB
* VNB	VNB
MM1033 N_VGND_M1033_d N_CLK_M1033_g N_A_27_79#_M1033_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1006 N_A_196_79#_M1006_d N_A_27_79#_M1006_g N_VGND_M1033_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1001 A_427_191# N_RESET_B_M1001_g N_VGND_M1001_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.32025 PD=0.63 PS=2.69 NRD=14.28 NRS=202.14 M=1 R=2.8 SA=75000.3
+ SB=75004.7 A=0.063 P=1.14 MULT=1
MM1027 N_A_308_463#_M1027_d N_D_M1027_g A_427_191# VNB NSHORT L=0.15 W=0.42
+ AD=0.1134 AS=0.0441 PD=0.96 PS=0.63 NRD=74.28 NRS=14.28 M=1 R=2.8 SA=75000.7
+ SB=75004.3 A=0.063 P=1.14 MULT=1
MM1028 N_A_637_191#_M1028_d N_A_27_79#_M1028_g N_A_308_463#_M1027_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.12285 AS=0.1134 PD=1.005 PS=0.96 NRD=87.132 NRS=0 M=1 R=2.8
+ SA=75001.4 SB=75003.6 A=0.063 P=1.14 MULT=1
MM1002 A_784_191# N_A_196_79#_M1002_g N_A_637_191#_M1028_d VNB NSHORT L=0.15
+ W=0.42 AD=0.04935 AS=0.12285 PD=0.655 PS=1.005 NRD=17.856 NRS=0 M=1 R=2.8
+ SA=75002.1 SB=75002.9 A=0.063 P=1.14 MULT=1
MM1034 A_861_191# N_A_811_341#_M1034_g A_784_191# VNB NSHORT L=0.15 W=0.42
+ AD=0.05775 AS=0.04935 PD=0.695 PS=0.655 NRD=23.568 NRS=17.856 M=1 R=2.8
+ SA=75002.5 SB=75002.5 A=0.063 P=1.14 MULT=1
MM1032 N_VGND_M1032_d N_RESET_B_M1032_g A_861_191# VNB NSHORT L=0.15 W=0.42
+ AD=0.23625 AS=0.05775 PD=1.56906 PS=0.695 NRD=144.996 NRS=23.568 M=1 R=2.8
+ SA=75002.9 SB=75002.1 A=0.063 P=1.14 MULT=1
MM1007 N_A_811_341#_M1007_d N_A_637_191#_M1007_g N_VGND_M1032_d VNB NSHORT
+ L=0.15 W=0.64 AD=0.1264 AS=0.36 PD=1.035 PS=2.39094 NRD=0 NRS=95.148 M=1
+ R=4.26667 SA=75002.3 SB=75002.1 A=0.096 P=1.58 MULT=1
MM1013 N_A_1272_128#_M1013_d N_A_196_79#_M1013_g N_A_811_341#_M1007_d VNB NSHORT
+ L=0.15 W=0.64 AD=0.221102 AS=0.1264 PD=1.50943 PS=1.035 NRD=44.052 NRS=21.552
+ M=1 R=4.26667 SA=75002.8 SB=75001.5 A=0.096 P=1.58 MULT=1
MM1015 A_1424_128# N_A_27_79#_M1015_g N_A_1272_128#_M1013_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.145098 PD=0.63 PS=0.990566 NRD=14.28 NRS=27.132 M=1
+ R=2.8 SA=75002.7 SB=75001.3 A=0.063 P=1.14 MULT=1
MM1037 N_VGND_M1037_d N_A_1444_320#_M1037_g A_1424_128# VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75003 SB=75001
+ A=0.063 P=1.14 MULT=1
MM1003 A_1582_128# N_RESET_B_M1003_g N_VGND_M1037_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75003.4
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1029 N_A_1444_320#_M1029_d N_A_1272_128#_M1029_g A_1582_128# VNB NSHORT L=0.15
+ W=0.42 AD=0.1113 AS=0.0441 PD=1.37 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8
+ SA=75003.8 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1010 N_Q_N_M1010_d N_A_1272_128#_M1010_g N_VGND_M1010_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1022 N_Q_N_M1010_d N_A_1272_128#_M1022_g N_VGND_M1022_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1004 N_VGND_M1004_d N_A_1272_128#_M1004_g N_A_2028_367#_M1004_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.0896 AS=0.1113 PD=0.81 PS=1.37 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1021 N_Q_M1021_d N_A_2028_367#_M1021_g N_VGND_M1004_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1792 PD=1.12 PS=1.62 NRD=0 NRS=6.78 M=1 R=5.6 SA=75000.5
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1030 N_Q_M1021_d N_A_2028_367#_M1030_g N_VGND_M1030_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.9
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1005 N_VPWR_M1005_d N_CLK_M1005_g N_A_27_79#_M1005_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0896 AS=0.1696 PD=0.92 PS=1.81 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75000.6 A=0.096 P=1.58 MULT=1
MM1020 N_A_196_79#_M1020_d N_A_27_79#_M1020_g N_VPWR_M1005_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1696 AS=0.0896 PD=1.81 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.6 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1016 N_VPWR_M1016_d N_RESET_B_M1016_g N_A_308_463#_M1016_s VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1125 AS=0.1113 PD=1.02 PS=1.37 NRD=35.1645 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1008 N_A_308_463#_M1008_d N_D_M1008_g N_VPWR_M1016_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.1197 AS=0.1125 PD=1.41 PS=1.02 NRD=0 NRS=35.1645 M=1 R=2.8 SA=75000.8
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1019 N_A_637_191#_M1019_d N_A_196_79#_M1019_g N_A_308_463#_M1019_s VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.0588 AS=0.1155 PD=0.7 PS=1.39 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.5 A=0.063 P=1.14 MULT=1
MM1035 A_793_463# N_A_27_79#_M1035_g N_A_637_191#_M1019_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=23.443 NRS=0 M=1 R=2.8
+ SA=75000.6 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1000 N_VPWR_M1000_d N_A_811_341#_M1000_g A_793_463# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.1065 AS=0.0441 PD=1 PS=0.63 NRD=30.4759 NRS=23.443 M=1 R=2.8 SA=75001
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1012 N_A_637_191#_M1012_d N_RESET_B_M1012_g N_VPWR_M1000_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1113 AS=0.1065 PD=1.37 PS=1 NRD=0 NRS=30.4759 M=1 R=2.8 SA=75001.5
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1025 N_A_811_341#_M1025_d N_A_637_191#_M1025_g N_VPWR_M1025_s VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.241012 AS=0.2226 PD=1.515 PS=2.21 NRD=22.655 NRS=0 M=1
+ R=5.6 SA=75000.2 SB=75001.7 A=0.126 P=1.98 MULT=1
MM1024 N_A_1272_128#_M1024_d N_A_27_79#_M1024_g N_A_811_341#_M1025_d VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.1792 AS=0.241012 PD=1.62 PS=1.515 NRD=0 NRS=32.0322 M=1
+ R=5.6 SA=75000.8 SB=75001.7 A=0.126 P=1.98 MULT=1
MM1031 A_1402_496# N_A_196_79#_M1031_g N_A_1272_128#_M1024_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0441 AS=0.0896 PD=0.63 PS=0.81 NRD=23.443 NRS=44.5417 M=1 R=2.8
+ SA=75001.2 SB=75002.8 A=0.063 P=1.14 MULT=1
MM1036 N_VPWR_M1036_d N_A_1444_320#_M1036_g A_1402_496# VPB PHIGHVT L=0.15
+ W=0.42 AD=0.13965 AS=0.0441 PD=1.085 PS=0.63 NRD=0 NRS=23.443 M=1 R=2.8
+ SA=75001.5 SB=75002.4 A=0.063 P=1.14 MULT=1
MM1011 N_A_1444_320#_M1011_d N_RESET_B_M1011_g N_VPWR_M1036_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0588 AS=0.13965 PD=0.7 PS=1.085 NRD=0 NRS=0 M=1 R=2.8 SA=75002.4
+ SB=75001.6 A=0.063 P=1.14 MULT=1
MM1017 N_VPWR_M1017_d N_A_1272_128#_M1017_g N_A_1444_320#_M1011_d VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.095025 AS=0.0588 PD=0.8175 PS=0.7 NRD=45.7237 NRS=0 M=1
+ R=2.8 SA=75002.8 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1009 N_VPWR_M1017_d N_A_1272_128#_M1009_g N_Q_N_M1009_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.285075 AS=0.1764 PD=2.4525 PS=1.54 NRD=0 NRS=0 M=1 R=8.4
+ SA=75001.2 SB=75000.6 A=0.189 P=2.82 MULT=1
MM1023 N_VPWR_M1023_d N_A_1272_128#_M1023_g N_Q_N_M1009_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.7
+ SB=75000.2 A=0.189 P=2.82 MULT=1
MM1014 N_VPWR_M1014_d N_A_1272_128#_M1014_g N_A_2028_367#_M1014_s VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.14912 AS=0.1696 PD=1.14189 PS=1.81 NRD=24.625 NRS=0 M=1
+ R=4.26667 SA=75000.2 SB=75001.2 A=0.096 P=1.58 MULT=1
MM1018 N_VPWR_M1014_d N_A_2028_367#_M1018_g N_Q_M1018_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.29358 AS=0.1764 PD=2.24811 PS=1.54 NRD=8.077 NRS=0 M=1 R=8.4
+ SA=75000.5 SB=75000.6 A=0.189 P=2.82 MULT=1
MM1026 N_VPWR_M1026_d N_A_2028_367#_M1026_g N_Q_M1018_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.9
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX38_noxref VNB VPB NWDIODE A=23.3096 P=29
*
.include "sky130_fd_sc_lp__dfrbp_2.pxi.spice"
*
.ends
*
*
