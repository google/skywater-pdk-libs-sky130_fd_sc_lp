* File: sky130_fd_sc_lp__nand2_4.pex.spice
* Created: Fri Aug 28 10:47:16 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__NAND2_4%B 3 7 11 15 19 23 27 31 33 34 35 36 54
c75 27 0 8.01629e-20 $X=1.945 $Y=0.745
r76 52 54 21.8577 $w=3.3e-07 $l=1.25e-07 $layer=POLY_cond $X=1.82 $Y=1.51
+ $X2=1.945 $Y2=1.51
r77 52 53 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.82
+ $Y=1.51 $X2=1.82 $Y2=1.51
r78 50 52 53.3327 $w=3.3e-07 $l=3.05e-07 $layer=POLY_cond $X=1.515 $Y=1.51
+ $X2=1.82 $Y2=1.51
r79 48 50 6.12014 $w=3.3e-07 $l=3.5e-08 $layer=POLY_cond $X=1.48 $Y=1.51
+ $X2=1.515 $Y2=1.51
r80 48 49 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.48
+ $Y=1.51 $X2=1.48 $Y2=1.51
r81 46 48 69.0702 $w=3.3e-07 $l=3.95e-07 $layer=POLY_cond $X=1.085 $Y=1.51
+ $X2=1.48 $Y2=1.51
r82 44 46 49.8355 $w=3.3e-07 $l=2.85e-07 $layer=POLY_cond $X=0.8 $Y=1.51
+ $X2=1.085 $Y2=1.51
r83 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.8
+ $Y=1.51 $X2=0.8 $Y2=1.51
r84 41 44 25.3549 $w=3.3e-07 $l=1.45e-07 $layer=POLY_cond $X=0.655 $Y=1.51
+ $X2=0.8 $Y2=1.51
r85 36 53 11.6964 $w=3.33e-07 $l=3.4e-07 $layer=LI1_cond $X=2.16 $Y=1.592
+ $X2=1.82 $Y2=1.592
r86 35 53 4.81618 $w=3.33e-07 $l=1.4e-07 $layer=LI1_cond $X=1.68 $Y=1.592
+ $X2=1.82 $Y2=1.592
r87 35 49 6.88026 $w=3.33e-07 $l=2e-07 $layer=LI1_cond $X=1.68 $Y=1.592 $X2=1.48
+ $Y2=1.592
r88 34 49 9.63236 $w=3.33e-07 $l=2.8e-07 $layer=LI1_cond $X=1.2 $Y=1.592
+ $X2=1.48 $Y2=1.592
r89 34 45 13.7605 $w=3.33e-07 $l=4e-07 $layer=LI1_cond $X=1.2 $Y=1.592 $X2=0.8
+ $Y2=1.592
r90 33 45 2.7521 $w=3.33e-07 $l=8e-08 $layer=LI1_cond $X=0.72 $Y=1.592 $X2=0.8
+ $Y2=1.592
r91 29 54 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.945 $Y=1.675
+ $X2=1.945 $Y2=1.51
r92 29 31 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.945 $Y=1.675
+ $X2=1.945 $Y2=2.465
r93 25 54 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.945 $Y=1.345
+ $X2=1.945 $Y2=1.51
r94 25 27 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=1.945 $Y=1.345
+ $X2=1.945 $Y2=0.745
r95 21 50 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.515 $Y=1.675
+ $X2=1.515 $Y2=1.51
r96 21 23 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.515 $Y=1.675
+ $X2=1.515 $Y2=2.465
r97 17 50 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.515 $Y=1.345
+ $X2=1.515 $Y2=1.51
r98 17 19 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=1.515 $Y=1.345
+ $X2=1.515 $Y2=0.745
r99 13 46 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.085 $Y=1.675
+ $X2=1.085 $Y2=1.51
r100 13 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.085 $Y=1.675
+ $X2=1.085 $Y2=2.465
r101 9 46 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.085 $Y=1.345
+ $X2=1.085 $Y2=1.51
r102 9 11 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=1.085 $Y=1.345
+ $X2=1.085 $Y2=0.745
r103 5 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.655 $Y=1.675
+ $X2=0.655 $Y2=1.51
r104 5 7 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=0.655 $Y=1.675
+ $X2=0.655 $Y2=2.465
r105 1 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.655 $Y=1.345
+ $X2=0.655 $Y2=1.51
r106 1 3 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=0.655 $Y=1.345 $X2=0.655
+ $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_LP__NAND2_4%A 3 7 11 15 19 23 27 31 33 37 38 41 49
r85 47 49 69.0702 $w=3.3e-07 $l=3.95e-07 $layer=POLY_cond $X=3.43 $Y=1.51
+ $X2=3.825 $Y2=1.51
r86 47 48 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.43
+ $Y=1.51 $X2=3.43 $Y2=1.51
r87 45 47 6.12014 $w=3.3e-07 $l=3.5e-08 $layer=POLY_cond $X=3.395 $Y=1.51
+ $X2=3.43 $Y2=1.51
r88 43 44 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.09
+ $Y=1.51 $X2=3.09 $Y2=1.51
r89 41 45 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=3.32 $Y=1.51
+ $X2=3.395 $Y2=1.51
r90 41 43 40.2181 $w=3.3e-07 $l=2.3e-07 $layer=POLY_cond $X=3.32 $Y=1.51
+ $X2=3.09 $Y2=1.51
r91 38 48 5.6787 $w=3.43e-07 $l=1.7e-07 $layer=LI1_cond $X=3.6 $Y=1.587 $X2=3.43
+ $Y2=1.587
r92 37 48 10.3553 $w=3.43e-07 $l=3.1e-07 $layer=LI1_cond $X=3.12 $Y=1.587
+ $X2=3.43 $Y2=1.587
r93 37 44 1.00212 $w=3.43e-07 $l=3e-08 $layer=LI1_cond $X=3.12 $Y=1.587 $X2=3.09
+ $Y2=1.587
r94 34 36 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=2.375 $Y=1.51
+ $X2=2.805 $Y2=1.51
r95 33 43 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=2.88 $Y=1.51
+ $X2=3.09 $Y2=1.51
r96 33 36 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=2.88 $Y=1.51
+ $X2=2.805 $Y2=1.51
r97 29 49 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.825 $Y=1.675
+ $X2=3.825 $Y2=1.51
r98 29 31 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.825 $Y=1.675
+ $X2=3.825 $Y2=2.465
r99 25 49 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.825 $Y=1.345
+ $X2=3.825 $Y2=1.51
r100 25 27 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=3.825 $Y=1.345
+ $X2=3.825 $Y2=0.745
r101 21 45 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.395 $Y=1.675
+ $X2=3.395 $Y2=1.51
r102 21 23 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.395 $Y=1.675
+ $X2=3.395 $Y2=2.465
r103 17 45 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.395 $Y=1.345
+ $X2=3.395 $Y2=1.51
r104 17 19 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=3.395 $Y=1.345
+ $X2=3.395 $Y2=0.745
r105 13 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.805 $Y=1.675
+ $X2=2.805 $Y2=1.51
r106 13 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.805 $Y=1.675
+ $X2=2.805 $Y2=2.465
r107 9 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.805 $Y=1.345
+ $X2=2.805 $Y2=1.51
r108 9 11 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=2.805 $Y=1.345
+ $X2=2.805 $Y2=0.745
r109 5 34 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.375 $Y=1.675
+ $X2=2.375 $Y2=1.51
r110 5 7 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.375 $Y=1.675
+ $X2=2.375 $Y2=2.465
r111 1 34 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.375 $Y=1.345
+ $X2=2.375 $Y2=1.51
r112 1 3 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=2.375 $Y=1.345 $X2=2.375
+ $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_LP__NAND2_4%VPWR 1 2 3 4 5 16 18 22 26 30 34 36 38 42 44
+ 49 54 63 66 69 73
r67 72 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r68 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r69 63 64 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r70 61 64 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.2 $Y2=3.33
r71 60 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r72 58 73 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r73 58 70 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=3.12 $Y2=3.33
r74 57 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r75 55 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.25 $Y=3.33
+ $X2=3.085 $Y2=3.33
r76 55 57 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=3.25 $Y=3.33 $X2=3.6
+ $Y2=3.33
r77 54 72 4.13553 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.94 $Y=3.33 $X2=4.13
+ $Y2=3.33
r78 54 57 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=3.94 $Y=3.33 $X2=3.6
+ $Y2=3.33
r79 53 70 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r80 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r81 50 66 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.325 $Y=3.33
+ $X2=2.16 $Y2=3.33
r82 50 52 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=2.325 $Y=3.33
+ $X2=2.64 $Y2=3.33
r83 49 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.92 $Y=3.33
+ $X2=3.085 $Y2=3.33
r84 49 52 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=2.92 $Y=3.33
+ $X2=2.64 $Y2=3.33
r85 48 64 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r86 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r87 45 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.465 $Y=3.33
+ $X2=1.3 $Y2=3.33
r88 45 47 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=1.465 $Y=3.33
+ $X2=1.68 $Y2=3.33
r89 44 66 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.995 $Y=3.33
+ $X2=2.16 $Y2=3.33
r90 44 47 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=1.995 $Y=3.33
+ $X2=1.68 $Y2=3.33
r91 42 53 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r92 42 48 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r93 42 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r94 38 41 42.1838 $w=2.63e-07 $l=9.7e-07 $layer=LI1_cond $X=4.072 $Y=1.98
+ $X2=4.072 $Y2=2.95
r95 36 72 3.11253 $w=2.65e-07 $l=1.1025e-07 $layer=LI1_cond $X=4.072 $Y=3.245
+ $X2=4.13 $Y2=3.33
r96 36 41 12.8291 $w=2.63e-07 $l=2.95e-07 $layer=LI1_cond $X=4.072 $Y=3.245
+ $X2=4.072 $Y2=2.95
r97 32 69 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.085 $Y=3.245
+ $X2=3.085 $Y2=3.33
r98 32 34 29.6841 $w=3.28e-07 $l=8.5e-07 $layer=LI1_cond $X=3.085 $Y=3.245
+ $X2=3.085 $Y2=2.395
r99 28 66 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.16 $Y=3.245
+ $X2=2.16 $Y2=3.33
r100 28 30 29.6841 $w=3.28e-07 $l=8.5e-07 $layer=LI1_cond $X=2.16 $Y=3.245
+ $X2=2.16 $Y2=2.395
r101 24 63 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.3 $Y=3.245 $X2=1.3
+ $Y2=3.33
r102 24 26 29.6841 $w=3.28e-07 $l=8.5e-07 $layer=LI1_cond $X=1.3 $Y=3.245
+ $X2=1.3 $Y2=2.395
r103 23 60 4.80136 $w=1.7e-07 $l=2.33e-07 $layer=LI1_cond $X=0.465 $Y=3.33
+ $X2=0.232 $Y2=3.33
r104 22 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.135 $Y=3.33
+ $X2=1.3 $Y2=3.33
r105 22 23 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.135 $Y=3.33
+ $X2=0.465 $Y2=3.33
r106 18 21 33.2175 $w=3.38e-07 $l=9.8e-07 $layer=LI1_cond $X=0.295 $Y=1.97
+ $X2=0.295 $Y2=2.95
r107 16 60 3.04979 $w=3.4e-07 $l=1.12161e-07 $layer=LI1_cond $X=0.295 $Y=3.245
+ $X2=0.232 $Y2=3.33
r108 16 21 9.99914 $w=3.38e-07 $l=2.95e-07 $layer=LI1_cond $X=0.295 $Y=3.245
+ $X2=0.295 $Y2=2.95
r109 5 41 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=3.9
+ $Y=1.835 $X2=4.04 $Y2=2.95
r110 5 38 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=3.9
+ $Y=1.835 $X2=4.04 $Y2=1.98
r111 4 34 300 $w=1.7e-07 $l=6.54523e-07 $layer=licon1_PDIFF $count=2 $X=2.88
+ $Y=1.835 $X2=3.085 $Y2=2.395
r112 3 30 300 $w=1.7e-07 $l=6.26099e-07 $layer=licon1_PDIFF $count=2 $X=2.02
+ $Y=1.835 $X2=2.16 $Y2=2.395
r113 2 26 300 $w=1.7e-07 $l=6.26099e-07 $layer=licon1_PDIFF $count=2 $X=1.16
+ $Y=1.835 $X2=1.3 $Y2=2.395
r114 1 21 400 $w=1.7e-07 $l=1.21776e-06 $layer=licon1_PDIFF $count=1 $X=0.165
+ $Y=1.835 $X2=0.38 $Y2=2.95
r115 1 18 400 $w=1.7e-07 $l=2.74317e-07 $layer=licon1_PDIFF $count=1 $X=0.165
+ $Y=1.835 $X2=0.38 $Y2=1.97
.ends

.subckt PM_SKY130_FD_SC_LP__NAND2_4%Y 1 2 3 4 5 6 19 21 25 29 32 35 37 39 41 45
+ 47 48 49 50 51 52 53 54 63 68 72
c87 47 0 8.01629e-20 $X=2.59 $Y=1.16
r88 54 72 4.61608 $w=2.1e-07 $l=1.75e-07 $layer=LI1_cond $X=3.595 $Y=2.035
+ $X2=3.42 $Y2=2.035
r89 53 72 15.8442 $w=2.08e-07 $l=3e-07 $layer=LI1_cond $X=3.12 $Y=2.035 $X2=3.42
+ $Y2=2.035
r90 53 73 19.2771 $w=2.08e-07 $l=3.65e-07 $layer=LI1_cond $X=3.12 $Y=2.035
+ $X2=2.755 $Y2=2.035
r91 52 68 4.11612 $w=2.1e-07 $l=1.65e-07 $layer=LI1_cond $X=2.59 $Y=2.035
+ $X2=2.425 $Y2=2.035
r92 52 73 4.11612 $w=2.1e-07 $l=1.65e-07 $layer=LI1_cond $X=2.59 $Y=2.035
+ $X2=2.755 $Y2=2.035
r93 51 68 13.9957 $w=2.08e-07 $l=2.65e-07 $layer=LI1_cond $X=2.16 $Y=2.035
+ $X2=2.425 $Y2=2.035
r94 51 69 17.6926 $w=2.08e-07 $l=3.35e-07 $layer=LI1_cond $X=2.16 $Y=2.035
+ $X2=1.825 $Y2=2.035
r95 50 63 4.74942 $w=2.1e-07 $l=9.5e-08 $layer=LI1_cond $X=1.73 $Y=2.035
+ $X2=1.635 $Y2=2.035
r96 50 69 4.74942 $w=2.1e-07 $l=9.5e-08 $layer=LI1_cond $X=1.73 $Y=2.035
+ $X2=1.825 $Y2=2.035
r97 50 63 1.05628 $w=2.08e-07 $l=2e-08 $layer=LI1_cond $X=1.615 $Y=2.035
+ $X2=1.635 $Y2=2.035
r98 49 50 21.9177 $w=2.08e-07 $l=4.15e-07 $layer=LI1_cond $X=1.2 $Y=2.035
+ $X2=1.615 $Y2=2.035
r99 49 64 12.4113 $w=2.08e-07 $l=2.35e-07 $layer=LI1_cond $X=1.2 $Y=2.035
+ $X2=0.965 $Y2=2.035
r100 48 64 4.43891 $w=2.1e-07 $l=1.65e-07 $layer=LI1_cond $X=0.8 $Y=2.035
+ $X2=0.965 $Y2=2.035
r101 43 45 13.0497 $w=3.38e-07 $l=3.85e-07 $layer=LI1_cond $X=3.605 $Y=1.075
+ $X2=3.605 $Y2=0.69
r102 39 54 2.76965 $w=3.5e-07 $l=1.05e-07 $layer=LI1_cond $X=3.595 $Y=2.14
+ $X2=3.595 $Y2=2.035
r103 39 41 24.6952 $w=3.48e-07 $l=7.5e-07 $layer=LI1_cond $X=3.595 $Y=2.14
+ $X2=3.595 $Y2=2.89
r104 38 47 3.80956 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.755 $Y=1.16
+ $X2=2.59 $Y2=1.16
r105 37 43 7.85115 $w=1.7e-07 $l=2.08207e-07 $layer=LI1_cond $X=3.435 $Y=1.16
+ $X2=3.605 $Y2=1.075
r106 37 38 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=3.435 $Y=1.16
+ $X2=2.755 $Y2=1.16
r107 33 52 2.10475 $w=2.55e-07 $l=1.19937e-07 $layer=LI1_cond $X=2.622 $Y=2.14
+ $X2=2.59 $Y2=2.035
r108 33 35 33.8954 $w=2.53e-07 $l=7.5e-07 $layer=LI1_cond $X=2.622 $Y=2.14
+ $X2=2.622 $Y2=2.89
r109 32 52 2.10475 $w=3.3e-07 $l=1.05e-07 $layer=LI1_cond $X=2.59 $Y=1.93
+ $X2=2.59 $Y2=2.035
r110 31 47 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.59 $Y=1.245
+ $X2=2.59 $Y2=1.16
r111 31 32 23.9219 $w=3.28e-07 $l=6.85e-07 $layer=LI1_cond $X=2.59 $Y=1.245
+ $X2=2.59 $Y2=1.93
r112 27 47 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.59 $Y=1.075
+ $X2=2.59 $Y2=1.16
r113 27 29 13.0959 $w=3.28e-07 $l=3.75e-07 $layer=LI1_cond $X=2.59 $Y=1.075
+ $X2=2.59 $Y2=0.7
r114 23 50 1.70532 $w=1.9e-07 $l=1.05e-07 $layer=LI1_cond $X=1.73 $Y=2.14
+ $X2=1.73 $Y2=2.035
r115 23 25 43.7799 $w=1.88e-07 $l=7.5e-07 $layer=LI1_cond $X=1.73 $Y=2.14
+ $X2=1.73 $Y2=2.89
r116 19 48 2.82476 $w=3.3e-07 $l=1.05e-07 $layer=LI1_cond $X=0.8 $Y=2.14 $X2=0.8
+ $Y2=2.035
r117 19 21 26.1919 $w=3.28e-07 $l=7.5e-07 $layer=LI1_cond $X=0.8 $Y=2.14 $X2=0.8
+ $Y2=2.89
r118 6 54 400 $w=1.7e-07 $l=3.2249e-07 $layer=licon1_PDIFF $count=1 $X=3.47
+ $Y=1.835 $X2=3.61 $Y2=2.095
r119 6 41 400 $w=1.7e-07 $l=1.12282e-06 $layer=licon1_PDIFF $count=1 $X=3.47
+ $Y=1.835 $X2=3.61 $Y2=2.89
r120 5 52 400 $w=1.7e-07 $l=3.2249e-07 $layer=licon1_PDIFF $count=1 $X=2.45
+ $Y=1.835 $X2=2.59 $Y2=2.095
r121 5 35 400 $w=1.7e-07 $l=1.12282e-06 $layer=licon1_PDIFF $count=1 $X=2.45
+ $Y=1.835 $X2=2.59 $Y2=2.89
r122 4 50 400 $w=1.7e-07 $l=3.2249e-07 $layer=licon1_PDIFF $count=1 $X=1.59
+ $Y=1.835 $X2=1.73 $Y2=2.095
r123 4 25 400 $w=1.7e-07 $l=1.12282e-06 $layer=licon1_PDIFF $count=1 $X=1.59
+ $Y=1.835 $X2=1.73 $Y2=2.89
r124 3 48 400 $w=1.7e-07 $l=3.2249e-07 $layer=licon1_PDIFF $count=1 $X=0.73
+ $Y=1.835 $X2=0.87 $Y2=2.095
r125 3 21 400 $w=1.7e-07 $l=1.12282e-06 $layer=licon1_PDIFF $count=1 $X=0.73
+ $Y=1.835 $X2=0.87 $Y2=2.89
r126 2 45 91 $w=1.7e-07 $l=4.29331e-07 $layer=licon1_NDIFF $count=2 $X=3.47
+ $Y=0.325 $X2=3.61 $Y2=0.69
r127 1 29 91 $w=1.7e-07 $l=4.3946e-07 $layer=licon1_NDIFF $count=2 $X=2.45
+ $Y=0.325 $X2=2.59 $Y2=0.7
.ends

.subckt PM_SKY130_FD_SC_LP__NAND2_4%A_63_65# 1 2 3 4 5 18 20 21 24 26 32 33 36
+ 38 42 44 45
r64 40 42 1.55137 $w=2.58e-07 $l=3.5e-08 $layer=LI1_cond $X=4.075 $Y=0.435
+ $X2=4.075 $Y2=0.47
r65 39 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.265 $Y=0.35
+ $X2=3.1 $Y2=0.35
r66 38 40 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=3.945 $Y=0.35
+ $X2=4.075 $Y2=0.435
r67 38 39 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=3.945 $Y=0.35
+ $X2=3.265 $Y2=0.35
r68 34 45 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.1 $Y=0.435 $X2=3.1
+ $Y2=0.35
r69 34 36 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=3.1 $Y=0.435
+ $X2=3.1 $Y2=0.45
r70 32 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.935 $Y=0.35
+ $X2=3.1 $Y2=0.35
r71 32 33 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=2.935 $Y=0.35
+ $X2=2.255 $Y2=0.35
r72 29 31 35.8995 $w=1.88e-07 $l=6.15e-07 $layer=LI1_cond $X=2.16 $Y=1.085
+ $X2=2.16 $Y2=0.47
r73 28 33 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=2.16 $Y=0.435
+ $X2=2.255 $Y2=0.35
r74 28 31 2.04306 $w=1.88e-07 $l=3.5e-08 $layer=LI1_cond $X=2.16 $Y=0.435
+ $X2=2.16 $Y2=0.47
r75 27 44 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.395 $Y=1.17 $X2=1.3
+ $Y2=1.17
r76 26 29 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=2.065 $Y=1.17
+ $X2=2.16 $Y2=1.085
r77 26 27 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.065 $Y=1.17
+ $X2=1.395 $Y2=1.17
r78 22 44 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.3 $Y=1.085 $X2=1.3
+ $Y2=1.17
r79 22 24 35.8995 $w=1.88e-07 $l=6.15e-07 $layer=LI1_cond $X=1.3 $Y=1.085
+ $X2=1.3 $Y2=0.47
r80 20 44 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.205 $Y=1.17 $X2=1.3
+ $Y2=1.17
r81 20 21 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.205 $Y=1.17
+ $X2=0.535 $Y2=1.17
r82 16 21 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.41 $Y=1.085
+ $X2=0.535 $Y2=1.17
r83 16 18 28.3501 $w=2.48e-07 $l=6.15e-07 $layer=LI1_cond $X=0.41 $Y=1.085
+ $X2=0.41 $Y2=0.47
r84 5 42 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.9
+ $Y=0.325 $X2=4.04 $Y2=0.47
r85 4 36 91 $w=1.7e-07 $l=2.755e-07 $layer=licon1_NDIFF $count=2 $X=2.88
+ $Y=0.325 $X2=3.1 $Y2=0.45
r86 3 31 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.02
+ $Y=0.325 $X2=2.16 $Y2=0.47
r87 2 24 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.16
+ $Y=0.325 $X2=1.3 $Y2=0.47
r88 1 18 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.315
+ $Y=0.325 $X2=0.44 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_LP__NAND2_4%VGND 1 2 11 15 17 19 29 30 33 36
r50 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r51 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r52 29 30 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r53 26 29 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=2.16 $Y=0 $X2=4.08
+ $Y2=0
r54 24 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.895 $Y=0 $X2=1.73
+ $Y2=0
r55 24 26 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=1.895 $Y=0 $X2=2.16
+ $Y2=0
r56 23 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r57 23 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r58 22 23 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r59 20 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.035 $Y=0 $X2=0.87
+ $Y2=0
r60 20 22 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=1.035 $Y=0 $X2=1.2
+ $Y2=0
r61 19 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.565 $Y=0 $X2=1.73
+ $Y2=0
r62 19 22 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=1.565 $Y=0 $X2=1.2
+ $Y2=0
r63 17 30 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=2.16 $Y=0 $X2=4.08
+ $Y2=0
r64 17 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.68
+ $Y2=0
r65 17 26 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r66 13 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.73 $Y=0.085
+ $X2=1.73 $Y2=0
r67 13 15 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=1.73 $Y=0.085
+ $X2=1.73 $Y2=0.47
r68 9 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.87 $Y=0.085 $X2=0.87
+ $Y2=0
r69 9 11 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=0.87 $Y=0.085
+ $X2=0.87 $Y2=0.45
r70 2 15 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.59
+ $Y=0.325 $X2=1.73 $Y2=0.47
r71 1 11 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=0.73
+ $Y=0.325 $X2=0.87 $Y2=0.45
.ends

