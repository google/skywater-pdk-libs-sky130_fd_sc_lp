* File: sky130_fd_sc_lp__nand4_1.pex.spice
* Created: Wed Sep  2 10:05:28 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__NAND4_1%D 3 6 8 9 13 15
r25 13 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.5 $Y=1.35 $X2=0.5
+ $Y2=1.515
r26 13 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.5 $Y=1.35 $X2=0.5
+ $Y2=1.185
r27 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.5
+ $Y=1.35 $X2=0.5 $Y2=1.35
r28 9 14 11.2683 $w=2.23e-07 $l=2.2e-07 $layer=LI1_cond $X=0.72 $Y=1.322 $X2=0.5
+ $Y2=1.322
r29 8 14 13.3171 $w=2.23e-07 $l=2.6e-07 $layer=LI1_cond $X=0.24 $Y=1.322 $X2=0.5
+ $Y2=1.322
r30 6 16 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=0.59 $Y=2.465
+ $X2=0.59 $Y2=1.515
r31 3 15 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.59 $Y=0.655
+ $X2=0.59 $Y2=1.185
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4_1%C 3 6 8 9 10 15 17
r31 15 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.07 $Y=1.35
+ $X2=1.07 $Y2=1.515
r32 15 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.07 $Y=1.35
+ $X2=1.07 $Y2=1.185
r33 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.07
+ $Y=1.35 $X2=1.07 $Y2=1.35
r34 10 16 2.11281 $w=2.98e-07 $l=5.5e-08 $layer=LI1_cond $X=1.135 $Y=1.295
+ $X2=1.135 $Y2=1.35
r35 9 10 14.2135 $w=2.98e-07 $l=3.7e-07 $layer=LI1_cond $X=1.135 $Y=0.925
+ $X2=1.135 $Y2=1.295
r36 8 9 14.2135 $w=2.98e-07 $l=3.7e-07 $layer=LI1_cond $X=1.135 $Y=0.555
+ $X2=1.135 $Y2=0.925
r37 6 18 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=1.02 $Y=2.465
+ $X2=1.02 $Y2=1.515
r38 3 17 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.98 $Y=0.655
+ $X2=0.98 $Y2=1.185
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4_1%B 3 6 8 9 10 15 17
r32 15 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.64 $Y=1.35
+ $X2=1.64 $Y2=1.515
r33 15 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.64 $Y=1.35
+ $X2=1.64 $Y2=1.185
r34 10 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.64
+ $Y=1.35 $X2=1.64 $Y2=1.35
r35 9 10 19.5411 $w=2.08e-07 $l=3.7e-07 $layer=LI1_cond $X=1.66 $Y=0.925
+ $X2=1.66 $Y2=1.295
r36 8 9 19.5411 $w=2.08e-07 $l=3.7e-07 $layer=LI1_cond $X=1.66 $Y=0.555 $X2=1.66
+ $Y2=0.925
r37 6 18 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=1.69 $Y=2.465
+ $X2=1.69 $Y2=1.515
r38 3 17 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.55 $Y=0.655
+ $X2=1.55 $Y2=1.185
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4_1%A 3 6 8 9 10 15 17
r31 15 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.21 $Y=1.35
+ $X2=2.21 $Y2=1.515
r32 15 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.21 $Y=1.35
+ $X2=2.21 $Y2=1.185
r33 10 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.21
+ $Y=1.35 $X2=2.21 $Y2=1.35
r34 9 10 19.382 $w=2.18e-07 $l=3.7e-07 $layer=LI1_cond $X=2.185 $Y=0.925
+ $X2=2.185 $Y2=1.295
r35 8 9 19.382 $w=2.18e-07 $l=3.7e-07 $layer=LI1_cond $X=2.185 $Y=0.555
+ $X2=2.185 $Y2=0.925
r36 6 18 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=2.12 $Y=2.465
+ $X2=2.12 $Y2=1.515
r37 3 17 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.12 $Y=0.655
+ $X2=2.12 $Y2=1.185
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4_1%VPWR 1 2 3 10 12 16 20 22 24 28 30 39 43
r36 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r37 39 40 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r38 37 40 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.2 $Y2=3.33
r39 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r40 34 43 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r41 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r42 31 39 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.34 $Y=3.33
+ $X2=1.235 $Y2=3.33
r43 31 33 53.4973 $w=1.68e-07 $l=8.2e-07 $layer=LI1_cond $X=1.34 $Y=3.33
+ $X2=2.16 $Y2=3.33
r44 30 42 3.61693 $w=1.7e-07 $l=2.27e-07 $layer=LI1_cond $X=2.425 $Y=3.33
+ $X2=2.652 $Y2=3.33
r45 30 33 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=2.425 $Y=3.33
+ $X2=2.16 $Y2=3.33
r46 28 34 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=2.16 $Y2=3.33
r47 28 40 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=1.2 $Y2=3.33
r48 24 27 35.9134 $w=2.08e-07 $l=6.8e-07 $layer=LI1_cond $X=2.53 $Y=2.27
+ $X2=2.53 $Y2=2.95
r49 22 42 3.29826 $w=2.1e-07 $l=1.58915e-07 $layer=LI1_cond $X=2.53 $Y=3.245
+ $X2=2.652 $Y2=3.33
r50 22 27 15.5801 $w=2.08e-07 $l=2.95e-07 $layer=LI1_cond $X=2.53 $Y=3.245
+ $X2=2.53 $Y2=2.95
r51 18 39 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=1.235 $Y=3.245
+ $X2=1.235 $Y2=3.33
r52 18 20 33.5368 $w=2.08e-07 $l=6.35e-07 $layer=LI1_cond $X=1.235 $Y=3.245
+ $X2=1.235 $Y2=2.61
r53 17 36 3.6162 $w=1.7e-07 $l=2.28e-07 $layer=LI1_cond $X=0.455 $Y=3.33
+ $X2=0.227 $Y2=3.33
r54 16 39 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.13 $Y=3.33
+ $X2=1.235 $Y2=3.33
r55 16 17 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=1.13 $Y=3.33
+ $X2=0.455 $Y2=3.33
r56 12 15 35.9134 $w=2.08e-07 $l=6.8e-07 $layer=LI1_cond $X=0.35 $Y=2.27
+ $X2=0.35 $Y2=2.95
r57 10 36 3.29899 $w=2.1e-07 $l=1.5995e-07 $layer=LI1_cond $X=0.35 $Y=3.245
+ $X2=0.227 $Y2=3.33
r58 10 15 15.5801 $w=2.08e-07 $l=2.95e-07 $layer=LI1_cond $X=0.35 $Y=3.245
+ $X2=0.35 $Y2=2.95
r59 3 27 400 $w=1.7e-07 $l=1.27151e-06 $layer=licon1_PDIFF $count=1 $X=2.195
+ $Y=1.835 $X2=2.53 $Y2=2.95
r60 3 24 400 $w=1.7e-07 $l=5.78749e-07 $layer=licon1_PDIFF $count=1 $X=2.195
+ $Y=1.835 $X2=2.53 $Y2=2.27
r61 2 20 300 $w=1.7e-07 $l=8.42096e-07 $layer=licon1_PDIFF $count=2 $X=1.095
+ $Y=1.835 $X2=1.235 $Y2=2.61
r62 1 15 400 $w=1.7e-07 $l=1.17584e-06 $layer=licon1_PDIFF $count=1 $X=0.225
+ $Y=1.835 $X2=0.35 $Y2=2.95
r63 1 12 400 $w=1.7e-07 $l=4.93559e-07 $layer=licon1_PDIFF $count=1 $X=0.225
+ $Y=1.835 $X2=0.35 $Y2=2.27
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4_1%Y 1 2 3 10 14 16 17 18 19 26 34 39
r43 19 26 7.70743 $w=2.67e-07 $l=2.22e-07 $layer=LI1_cond $X=2.022 $Y=1.937
+ $X2=1.8 $Y2=1.937
r44 19 39 4.82393 $w=6.13e-07 $l=2e-07 $layer=LI1_cond $X=2.022 $Y=2.12
+ $X2=2.022 $Y2=2.32
r45 18 26 3.78885 $w=3.63e-07 $l=1.2e-07 $layer=LI1_cond $X=1.68 $Y=1.937
+ $X2=1.8 $Y2=1.937
r46 17 18 15.1554 $w=3.63e-07 $l=4.8e-07 $layer=LI1_cond $X=1.2 $Y=1.937
+ $X2=1.68 $Y2=1.937
r47 17 27 9.1564 $w=3.63e-07 $l=2.9e-07 $layer=LI1_cond $X=1.2 $Y=1.937 $X2=0.91
+ $Y2=1.937
r48 16 27 3.00646 $w=3.65e-07 $l=1.38e-07 $layer=LI1_cond $X=0.772 $Y=1.937
+ $X2=0.91 $Y2=1.937
r49 16 34 6.85085 $w=4.43e-07 $l=2e-07 $layer=LI1_cond $X=0.772 $Y=2.12
+ $X2=0.772 $Y2=2.32
r50 12 14 61.5281 $w=2.08e-07 $l=1.165e-06 $layer=LI1_cond $X=2.58 $Y=1.755
+ $X2=2.58 $Y2=0.59
r51 11 19 7.70743 $w=2.67e-07 $l=2.67133e-07 $layer=LI1_cond $X=2.245 $Y=1.84
+ $X2=2.022 $Y2=1.937
r52 10 12 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=2.475 $Y=1.84
+ $X2=2.58 $Y2=1.755
r53 10 11 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=2.475 $Y=1.84
+ $X2=2.245 $Y2=1.84
r54 3 19 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.765
+ $Y=1.835 $X2=1.905 $Y2=1.98
r55 3 39 300 $w=1.7e-07 $l=5.50568e-07 $layer=licon1_PDIFF $count=2 $X=1.765
+ $Y=1.835 $X2=1.905 $Y2=2.32
r56 2 16 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.665
+ $Y=1.835 $X2=0.805 $Y2=1.98
r57 2 34 300 $w=1.7e-07 $l=5.50568e-07 $layer=licon1_PDIFF $count=2 $X=0.665
+ $Y=1.835 $X2=0.805 $Y2=2.32
r58 1 14 91 $w=1.7e-07 $l=5.3376e-07 $layer=licon1_NDIFF $count=2 $X=2.195
+ $Y=0.235 $X2=2.58 $Y2=0.59
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4_1%VGND 1 4 6 8 15 16
r27 19 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r28 15 16 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r29 13 20 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r30 12 15 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=0.72 $Y=0 $X2=2.64
+ $Y2=0
r31 12 13 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r32 10 19 3.60793 $w=1.7e-07 $l=2.4e-07 $layer=LI1_cond $X=0.48 $Y=0 $X2=0.24
+ $Y2=0
r33 10 12 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=0.48 $Y=0 $X2=0.72
+ $Y2=0
r34 8 16 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=1.44 $Y=0 $X2=2.64
+ $Y2=0
r35 8 13 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=0.72
+ $Y2=0
r36 4 19 3.30727 $w=2.1e-07 $l=1.72337e-07 $layer=LI1_cond $X=0.375 $Y=0.085
+ $X2=0.24 $Y2=0
r37 4 6 15.5801 $w=2.08e-07 $l=2.95e-07 $layer=LI1_cond $X=0.375 $Y=0.085
+ $X2=0.375 $Y2=0.38
r38 1 6 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.25
+ $Y=0.235 $X2=0.375 $Y2=0.38
.ends

