* File: sky130_fd_sc_lp__sleep_sergate_plv_14.pex.spice
* Created: Fri Aug 28 11:32:37 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__SLEEP_SERGATE_PLV_14%SLEEP 2 3 4 6 7 9 11 12 13 14
+ 15 22
r38 22 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=8.42
+ $Y=1.835 $X2=8.42 $Y2=1.835
r39 14 15 8.34998 $w=5.28e-07 $l=3.7e-07 $layer=LI1_cond $X=8.52 $Y=2.035
+ $X2=8.52 $Y2=2.405
r40 14 23 4.5135 $w=5.28e-07 $l=2e-07 $layer=LI1_cond $X=8.52 $Y=2.035 $X2=8.52
+ $Y2=1.835
r41 13 23 3.83648 $w=5.28e-07 $l=1.7e-07 $layer=LI1_cond $X=8.52 $Y=1.665
+ $X2=8.52 $Y2=1.835
r42 12 13 8.34998 $w=5.28e-07 $l=3.7e-07 $layer=LI1_cond $X=8.52 $Y=1.295
+ $X2=8.52 $Y2=1.665
r43 11 12 8.34998 $w=5.28e-07 $l=3.7e-07 $layer=LI1_cond $X=8.52 $Y=0.925
+ $X2=8.52 $Y2=1.295
r44 10 22 55.6154 $w=4.15e-07 $l=4.15e-07 $layer=POLY_cond $X=8.377 $Y=2.25
+ $X2=8.377 $Y2=1.835
r45 7 9 1148.77 $w=1.5e-07 $l=3.575e-06 $layer=POLY_cond $X=0.98 $Y=2.755
+ $X2=4.555 $Y2=2.755
r46 4 6 1833.14 $w=1.5e-07 $l=3.575e-06 $layer=POLY_cond $X=0.98 $Y=2.325
+ $X2=4.555 $Y2=2.325
r47 3 10 35.4752 $w=1.5e-07 $l=2.41607e-07 $layer=POLY_cond $X=8.17 $Y=2.325
+ $X2=8.377 $Y2=2.25
r48 3 6 1853.65 $w=1.5e-07 $l=3.615e-06 $layer=POLY_cond $X=8.17 $Y=2.325
+ $X2=4.555 $Y2=2.325
r49 2 7 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.905 $Y=2.68
+ $X2=0.98 $Y2=2.755
r50 1 4 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.905 $Y=2.4
+ $X2=0.98 $Y2=2.325
r51 1 2 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=0.905 $Y=2.4 $X2=0.905
+ $Y2=2.68
.ends

.subckt PM_SKY130_FD_SC_LP__SLEEP_SERGATE_PLV_14%VIRTPWR 1 2 7 11 12 30 66 69 72
+ 75 77 81 82 89 90 95 99 104 105
c88 105 0 1.43534e-19 $X=6.51 $Y=3.33
c89 99 0 1.43534e-19 $X=4.955 $Y=3.33
c90 95 0 1.43534e-19 $X=3.4 $Y=3.33
c91 12 0 3.89769e-19 $X=0 $Y=3.085
c92 1 0 6.58418e-21 $X=1.055 $Y=1.985
r93 99 104 0.0432039 $w=4.9e-07 $l=1.55e-07 $layer=MET1_cond $X=4.955 $Y=3.33
+ $X2=4.8 $Y2=3.33
r94 88 109 0.213232 $w=4.9e-07 $l=7.65e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=7.155 $Y2=3.33
r95 87 89 9.36939 $w=5.73e-07 $l=1.35e-07 $layer=LI1_cond $X=7.92 $Y=3.127
+ $X2=8.055 $Y2=3.127
r96 87 88 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r97 85 87 2.80818 $w=5.73e-07 $l=1.35e-07 $layer=LI1_cond $X=7.785 $Y=3.127
+ $X2=7.92 $Y2=3.127
r98 81 89 53.8235 $w=1.68e-07 $l=8.25e-07 $layer=LI1_cond $X=8.88 $Y=3.33
+ $X2=8.055 $Y2=3.33
r99 81 82 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r100 74 77 34.5733 $w=2.58e-07 $l=7.8e-07 $layer=LI1_cond $X=7.005 $Y=2.11
+ $X2=7.785 $Y2=2.11
r101 74 75 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.005 $Y=2.11
+ $X2=7.005 $Y2=2.11
r102 71 74 68.925 $w=2.58e-07 $l=1.555e-06 $layer=LI1_cond $X=5.45 $Y=2.11
+ $X2=7.005 $Y2=2.11
r103 71 72 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.45 $Y=2.11
+ $X2=5.45 $Y2=2.11
r104 68 71 68.925 $w=2.58e-07 $l=1.555e-06 $layer=LI1_cond $X=3.895 $Y=2.11
+ $X2=5.45 $Y2=2.11
r105 68 69 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.895 $Y=2.11
+ $X2=3.895 $Y2=2.11
r106 65 68 68.925 $w=2.58e-07 $l=1.555e-06 $layer=LI1_cond $X=2.34 $Y=2.11
+ $X2=3.895 $Y2=2.11
r107 65 66 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.34 $Y=2.11
+ $X2=2.34 $Y2=2.11
r108 62 65 44.9896 $w=2.58e-07 $l=1.015e-06 $layer=LI1_cond $X=1.325 $Y=2.11
+ $X2=2.34 $Y2=2.11
r109 60 75 0.175043 $w=6.45e-07 $l=8.6e-07 $layer=MET1_cond $X=6.832 $Y=2.97
+ $X2=6.832 $Y2=2.11
r110 59 60 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=7.005 $Y=2.97
+ $X2=7.005 $Y2=2.97
r111 57 105 0.00836204 $w=4.9e-07 $l=3e-08 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=6.51 $Y2=3.33
r112 56 59 10.9207 $w=5.73e-07 $l=5.25e-07 $layer=LI1_cond $X=6.48 $Y=3.127
+ $X2=7.005 $Y2=3.127
r113 56 57 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r114 53 56 19.9693 $w=5.73e-07 $l=9.6e-07 $layer=LI1_cond $X=5.52 $Y=3.127
+ $X2=6.48 $Y2=3.127
r115 51 72 0.180644 $w=6.25e-07 $l=8.6e-07 $layer=MET1_cond $X=5.267 $Y=2.97
+ $X2=5.267 $Y2=2.11
r116 50 53 1.4561 $w=5.73e-07 $l=7e-08 $layer=LI1_cond $X=5.45 $Y=3.127 $X2=5.52
+ $Y2=3.127
r117 50 51 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=5.45 $Y=2.97
+ $X2=5.45 $Y2=2.97
r118 48 104 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=4.8 $Y2=3.33
r119 47 50 18.5132 $w=5.73e-07 $l=8.9e-07 $layer=LI1_cond $X=4.56 $Y=3.127
+ $X2=5.45 $Y2=3.127
r120 47 48 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r121 45 69 0.180644 $w=6.25e-07 $l=8.6e-07 $layer=MET1_cond $X=3.712 $Y=2.97
+ $X2=3.712 $Y2=2.11
r122 44 47 13.8329 $w=5.73e-07 $l=6.65e-07 $layer=LI1_cond $X=3.895 $Y=3.127
+ $X2=4.56 $Y2=3.127
r123 44 45 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.895 $Y=2.97
+ $X2=3.895 $Y2=2.97
r124 42 95 0.0780457 $w=4.9e-07 $l=2.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.4 $Y2=3.33
r125 41 44 16.1211 $w=5.73e-07 $l=7.75e-07 $layer=LI1_cond $X=3.12 $Y=3.127
+ $X2=3.895 $Y2=3.127
r126 41 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r127 38 41 16.2251 $w=5.73e-07 $l=7.8e-07 $layer=LI1_cond $X=2.34 $Y=3.127
+ $X2=3.12 $Y2=3.127
r128 36 66 0.180644 $w=6.25e-07 $l=8.6e-07 $layer=MET1_cond $X=2.157 $Y=2.97
+ $X2=2.157 $Y2=2.11
r129 36 38 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.34 $Y=2.97
+ $X2=2.34 $Y2=2.97
r130 35 38 7.48849 $w=5.73e-07 $l=3.6e-07 $layer=LI1_cond $X=1.98 $Y=3.127
+ $X2=2.34 $Y2=3.127
r131 35 36 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.98 $Y=2.97
+ $X2=1.98 $Y2=2.97
r132 33 90 0.0459912 $w=4.9e-07 $l=1.65e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.845 $Y2=3.33
r133 32 35 6.24041 $w=5.73e-07 $l=3e-07 $layer=LI1_cond $X=1.68 $Y=3.127
+ $X2=1.98 $Y2=3.127
r134 32 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r135 30 85 0.353623 $w=5.73e-07 $l=1.7e-08 $layer=LI1_cond $X=7.768 $Y=3.127
+ $X2=7.785 $Y2=3.127
r136 30 59 15.8714 $w=5.73e-07 $l=7.63e-07 $layer=LI1_cond $X=7.768 $Y=3.127
+ $X2=7.005 $Y2=3.127
r137 27 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r138 12 105 0.0661031 $w=4.9e-07 $l=3.22e-07 $layer=MET1_cond $X=6.832 $Y=3.33
+ $X2=6.51 $Y2=3.33
r139 12 109 0.0661031 $w=4.9e-07 $l=3.23e-07 $layer=MET1_cond $X=6.832 $Y=3.33
+ $X2=7.155 $Y2=3.33
r140 12 99 0.0644858 $w=4.9e-07 $l=3.12e-07 $layer=MET1_cond $X=5.267 $Y=3.33
+ $X2=4.955 $Y2=3.33
r141 12 106 0.0644858 $w=4.9e-07 $l=3.13e-07 $layer=MET1_cond $X=5.267 $Y=3.33
+ $X2=5.58 $Y2=3.33
r142 12 95 0.0644858 $w=4.9e-07 $l=3.12e-07 $layer=MET1_cond $X=3.712 $Y=3.33
+ $X2=3.4 $Y2=3.33
r143 12 100 0.0644858 $w=4.9e-07 $l=3.13e-07 $layer=MET1_cond $X=3.712 $Y=3.33
+ $X2=4.025 $Y2=3.33
r144 12 90 0.0644858 $w=4.9e-07 $l=3.12e-07 $layer=MET1_cond $X=2.157 $Y=3.33
+ $X2=1.845 $Y2=3.33
r145 12 96 0.0644858 $w=4.9e-07 $l=3.13e-07 $layer=MET1_cond $X=2.157 $Y=3.33
+ $X2=2.47 $Y2=3.33
r146 12 60 0.044502 $w=1.29e-06 $l=1.15e-07 $layer=MET1_cond $X=6.832 $Y=3.085
+ $X2=6.832 $Y2=2.97
r147 12 51 0.0448765 $w=1.25e-06 $l=1.15e-07 $layer=MET1_cond $X=5.267 $Y=3.085
+ $X2=5.267 $Y2=2.97
r148 12 45 0.0448765 $w=1.25e-06 $l=1.15e-07 $layer=MET1_cond $X=3.712 $Y=3.085
+ $X2=3.712 $Y2=2.97
r149 12 36 0.0448765 $w=1.25e-06 $l=1.15e-07 $layer=MET1_cond $X=2.157 $Y=3.085
+ $X2=2.157 $Y2=2.97
r150 12 82 0.2071 $w=4.9e-07 $l=7.43e-07 $layer=MET1_cond $X=8.137 $Y=3.33
+ $X2=8.88 $Y2=3.33
r151 12 88 0.0604854 $w=4.9e-07 $l=2.17e-07 $layer=MET1_cond $X=8.137 $Y=3.33
+ $X2=7.92 $Y2=3.33
r152 12 57 0.12125 $w=4.9e-07 $l=4.35e-07 $layer=MET1_cond $X=6.045 $Y=3.33
+ $X2=6.48 $Y2=3.33
r153 12 106 0.129612 $w=4.9e-07 $l=4.65e-07 $layer=MET1_cond $X=6.045 $Y=3.33
+ $X2=5.58 $Y2=3.33
r154 12 48 0.0195114 $w=4.9e-07 $l=7e-08 $layer=MET1_cond $X=4.49 $Y=3.33
+ $X2=4.56 $Y2=3.33
r155 12 100 0.129612 $w=4.9e-07 $l=4.65e-07 $layer=MET1_cond $X=4.49 $Y=3.33
+ $X2=4.025 $Y2=3.33
r156 12 42 0.0515659 $w=4.9e-07 $l=1.85e-07 $layer=MET1_cond $X=2.935 $Y=3.33
+ $X2=3.12 $Y2=3.33
r157 12 96 0.129612 $w=4.9e-07 $l=4.65e-07 $layer=MET1_cond $X=2.935 $Y=3.33
+ $X2=2.47 $Y2=3.33
r158 12 33 0.211281 $w=4.9e-07 $l=7.58e-07 $layer=MET1_cond $X=0.922 $Y=3.33
+ $X2=1.68 $Y2=3.33
r159 12 28 0.0563044 $w=4.9e-07 $l=2.02e-07 $layer=MET1_cond $X=0.922 $Y=3.33
+ $X2=0.72 $Y2=3.33
r160 12 53 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r161 11 27 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.055 $Y=3.33
+ $X2=0.72 $Y2=3.33
r162 10 11 12.1776 $w=5.73e-07 $l=2.7e-07 $layer=LI1_cond $X=1.325 $Y=3.127
+ $X2=1.055 $Y2=3.127
r163 7 32 7.03086 $w=5.73e-07 $l=3.38e-07 $layer=LI1_cond $X=1.342 $Y=3.127
+ $X2=1.68 $Y2=3.127
r164 7 10 0.353623 $w=5.73e-07 $l=1.7e-08 $layer=LI1_cond $X=1.342 $Y=3.127
+ $X2=1.325 $Y2=3.127
r165 2 85 60 $w=1.7e-07 $l=6.79964e-06 $layer=licon1_PDIFF $count=10 $X=1.055
+ $Y=2.83 $X2=7.785 $Y2=2.97
r166 2 10 60 $w=1.7e-07 $l=3.32716e-07 $layer=licon1_PDIFF $count=10 $X=1.055
+ $Y=2.83 $X2=1.325 $Y2=2.97
r167 1 77 60 $w=1.7e-07 $l=6.79221e-06 $layer=licon1_PDIFF $count=10 $X=1.055
+ $Y=1.985 $X2=7.785 $Y2=2.11
r168 1 62 60 $w=1.7e-07 $l=3.26573e-07 $layer=licon1_PDIFF $count=10 $X=1.055
+ $Y=1.985 $X2=1.325 $Y2=2.11
.ends

.subckt PM_SKY130_FD_SC_LP__SLEEP_SERGATE_PLV_14%VPWR 1 4 22 27 32 37 42 47 48
c69 48 0 6.58418e-21 $X=7.775 $Y=2.54
r70 47 48 2.25 $w=1.5e-07 $l=3e-07 $layer=via $count=2 $X=7.775 $Y=2.54
+ $X2=7.775 $Y2=2.54
r71 43 48 0.0591216 $w=3.33e-06 $l=1.575e-06 $layer=MET2_cond $X=6.2 $Y=1.665
+ $X2=7.775 $Y2=1.665
r72 42 43 2.25 $w=1.5e-07 $l=3e-07 $layer=via $count=2 $X=6.2 $Y=2.54 $X2=6.2
+ $Y2=2.54
r73 38 43 0.0583709 $w=3.33e-06 $l=1.555e-06 $layer=MET2_cond $X=4.645 $Y=1.665
+ $X2=6.2 $Y2=1.665
r74 37 38 2.25 $w=1.5e-07 $l=3e-07 $layer=via $count=2 $X=4.645 $Y=2.54
+ $X2=4.645 $Y2=2.54
r75 32 33 2.25 $w=1.5e-07 $l=3e-07 $layer=via $count=2 $X=3.09 $Y=2.54 $X2=3.09
+ $Y2=2.54
r76 28 33 0.0579955 $w=3.33e-06 $l=1.545e-06 $layer=MET2_cond $X=1.545 $Y=1.665
+ $X2=3.09 $Y2=1.665
r77 27 28 2.25 $w=1.5e-07 $l=3e-07 $layer=via $count=2 $X=1.545 $Y=2.54
+ $X2=1.545 $Y2=2.54
r78 22 47 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.8 $Y=2.54 $X2=7.8
+ $Y2=2.54
r79 19 22 69.1466 $w=2.58e-07 $l=1.56e-06 $layer=LI1_cond $X=6.225 $Y=2.54
+ $X2=7.785 $Y2=2.54
r80 19 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.225 $Y=2.54
+ $X2=6.225 $Y2=2.54
r81 16 19 68.925 $w=2.58e-07 $l=1.555e-06 $layer=LI1_cond $X=4.67 $Y=2.54
+ $X2=6.225 $Y2=2.54
r82 16 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.67 $Y=2.54
+ $X2=4.67 $Y2=2.54
r83 13 16 68.925 $w=2.58e-07 $l=1.555e-06 $layer=LI1_cond $X=3.115 $Y=2.54
+ $X2=4.67 $Y2=2.54
r84 13 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.115 $Y=2.54
+ $X2=3.115 $Y2=2.54
r85 10 13 68.925 $w=2.58e-07 $l=1.555e-06 $layer=LI1_cond $X=1.56 $Y=2.54
+ $X2=3.115 $Y2=2.54
r86 10 27 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.56 $Y=2.54
+ $X2=1.56 $Y2=2.54
r87 7 10 10.4163 $w=2.58e-07 $l=2.35e-07 $layer=LI1_cond $X=1.325 $Y=2.54
+ $X2=1.56 $Y2=2.54
r88 4 38 0.00319069 $w=3.33e-06 $l=8.5e-08 $layer=MET2_cond $X=4.56 $Y=1.665
+ $X2=4.645 $Y2=1.665
r89 4 33 0.0551802 $w=3.33e-06 $l=1.47e-06 $layer=MET2_cond $X=4.56 $Y=1.665
+ $X2=3.09 $Y2=1.665
r90 1 22 60 $w=1.7e-07 $l=6.79964e-06 $layer=licon1_PDIFF $count=10 $X=1.055
+ $Y=2.4 $X2=7.785 $Y2=2.54
r91 1 7 60 $w=1.7e-07 $l=3.32716e-07 $layer=licon1_PDIFF $count=10 $X=1.055
+ $Y=2.4 $X2=1.325 $Y2=2.54
.ends

