* NGSPICE file created from sky130_fd_sc_lp__sdfsbp_1.ext - technology: sky130A

.subckt sky130_fd_sc_lp__sdfsbp_1 CLK D SCD SCE SET_B VGND VNB VPB VPWR Q Q_N
M1000 a_1232_463# a_640_481# a_1146_463# VPB phighvt w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=1.176e+11p ps=1.4e+06u
M1001 VPWR a_2067_92# a_2025_488# VPB phighvt w=420000u l=150000u
+  ad=2.99083e+12p pd=2.169e+07u as=8.82e+10p ps=1.26e+06u
M1002 a_2582_150# a_1920_119# VGND VNB nshort w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=1.7578e+12p ps=1.526e+07u
M1003 a_1920_119# SET_B VPWR VPB phighvt w=420000u l=150000u
+  ad=3.801e+11p pd=3.8e+06u as=0p ps=0u
M1004 a_1274_401# a_1146_463# VPWR VPB phighvt w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=0p ps=0u
M1005 a_1575_119# a_1146_463# a_1274_401# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=1.113e+11p ps=1.37e+06u
M1006 a_478_47# SCE a_275_481# VNB nshort w=420000u l=150000u
+  ad=1.155e+11p pd=1.39e+06u as=3.717e+11p ps=3.45e+06u
M1007 Q_N a_1920_119# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=3.339e+11p pd=3.05e+06u as=0p ps=0u
M1008 a_383_481# a_34_481# a_275_481# VPB phighvt w=640000u l=150000u
+  ad=1.344e+11p pd=1.7e+06u as=3.609e+11p ps=3.43e+06u
M1009 a_640_481# CLK VPWR VPB phighvt w=640000u l=150000u
+  ad=1.696e+11p pd=1.81e+06u as=0p ps=0u
M1010 VPWR SET_B a_1274_401# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR SCD a_383_481# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_2025_488# a_901_441# a_1920_119# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VGND SCE a_34_481# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1014 a_275_481# D a_252_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1015 VGND a_1274_401# a_1245_119# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1016 VPWR a_1920_119# a_2067_92# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1017 a_901_441# a_640_481# VPWR VPB phighvt w=640000u l=150000u
+  ad=1.696e+11p pd=1.81e+06u as=0p ps=0u
M1018 a_1146_463# a_901_441# a_275_481# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_1818_379# a_1146_463# VPWR VPB phighvt w=840000u l=150000u
+  ad=3.199e+11p pd=2.65e+06u as=0p ps=0u
M1020 VGND a_2582_150# Q VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=2.394e+11p ps=2.25e+06u
M1021 Q_N a_1920_119# VGND VNB nshort w=840000u l=150000u
+  ad=2.226e+11p pd=2.21e+06u as=0p ps=0u
M1022 VPWR SCE a_34_481# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.696e+11p ps=1.81e+06u
M1023 a_640_481# CLK VGND VNB nshort w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1024 a_1146_463# a_640_481# a_275_481# VNB nshort w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=0p ps=0u
M1025 a_1245_119# a_901_441# a_1146_463# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_901_441# a_640_481# VGND VNB nshort w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1027 VPWR a_2582_150# Q VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=3.339e+11p ps=3.05e+06u
M1028 VGND SET_B a_2097_118# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1029 a_1848_119# a_1146_463# VGND VNB nshort w=640000u l=150000u
+  ad=1.344e+11p pd=1.7e+06u as=0p ps=0u
M1030 a_2025_118# a_640_481# a_1920_119# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=2.165e+11p ps=2.04e+06u
M1031 VPWR a_1274_401# a_1232_463# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 a_252_47# a_34_481# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 VGND a_1920_119# a_2067_92# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1034 a_203_481# SCE VPWR VPB phighvt w=640000u l=150000u
+  ad=1.344e+11p pd=1.7e+06u as=0p ps=0u
M1035 a_2097_118# a_2067_92# a_2025_118# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1036 VGND SCD a_478_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1037 a_2582_150# a_1920_119# VPWR VPB phighvt w=640000u l=150000u
+  ad=1.696e+11p pd=1.81e+06u as=0p ps=0u
M1038 a_1920_119# a_901_441# a_1848_119# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1039 a_275_481# D a_203_481# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1040 a_1920_119# a_640_481# a_1818_379# VPB phighvt w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1041 VGND SET_B a_1575_119# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

