* NGSPICE file created from sky130_fd_sc_lp__o41a_0.ext - technology: sky130A

.subckt sky130_fd_sc_lp__o41a_0 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
M1000 a_319_51# A3 VGND VNB nshort w=420000u l=150000u
+  ad=3.465e+11p pd=4.17e+06u as=3.717e+11p ps=4.29e+06u
M1001 VPWR A1 a_603_483# VPB phighvt w=640000u l=150000u
+  ad=3.488e+11p pd=3.65e+06u as=1.344e+11p ps=1.7e+06u
M1002 a_319_51# A1 VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 VGND a_80_21# X VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1004 VGND A2 a_319_51# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_80_21# B1 VPWR VPB phighvt w=640000u l=150000u
+  ad=5.12e+11p pd=2.88e+06u as=0p ps=0u
M1006 a_423_483# A4 a_80_21# VPB phighvt w=640000u l=150000u
+  ad=1.92e+11p pd=1.88e+06u as=0p ps=0u
M1007 a_319_51# B1 a_80_21# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1008 a_513_483# A3 a_423_483# VPB phighvt w=640000u l=150000u
+  ad=1.92e+11p pd=1.88e+06u as=0p ps=0u
M1009 VGND A4 a_319_51# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR a_80_21# X VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.696e+11p ps=1.81e+06u
M1011 a_603_483# A2 a_513_483# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

