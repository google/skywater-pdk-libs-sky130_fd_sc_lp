* File: sky130_fd_sc_lp__o22a_2.spice
* Created: Wed Sep  2 10:19:56 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__o22a_2.pex.spice"
.subckt sky130_fd_sc_lp__o22a_2  VNB VPB B1 B2 A2 A1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A1	A1
* A2	A2
* B2	B2
* B1	B1
* VPB	VPB
* VNB	VNB
MM1005 N_X_M1005_d N_A_80_23#_M1005_g N_VGND_M1005_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1007 N_X_M1005_d N_A_80_23#_M1007_g N_VGND_M1007_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1008 N_A_80_23#_M1008_d N_B1_M1008_g N_A_303_49#_M1008_s VNB NSHORT L=0.15
+ W=0.84 AD=0.126 AS=0.2226 PD=1.14 PS=2.21 NRD=2.856 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75001.6 A=0.126 P=1.98 MULT=1
MM1009 N_A_303_49#_M1009_d N_B2_M1009_g N_A_80_23#_M1008_d VNB NSHORT L=0.15
+ W=0.84 AD=0.1365 AS=0.126 PD=1.165 PS=1.14 NRD=2.856 NRS=0 M=1 R=5.6
+ SA=75000.6 SB=75001.2 A=0.126 P=1.98 MULT=1
MM1001 N_VGND_M1001_d N_A2_M1001_g N_A_303_49#_M1009_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1596 AS=0.1365 PD=1.22 PS=1.165 NRD=6.42 NRS=3.564 M=1 R=5.6 SA=75001.1
+ SB=75000.7 A=0.126 P=1.98 MULT=1
MM1002 N_A_303_49#_M1002_d N_A1_M1002_g N_VGND_M1001_d VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1596 PD=2.21 PS=1.22 NRD=0 NRS=7.848 M=1 R=5.6 SA=75001.6
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1000 N_X_M1000_d N_A_80_23#_M1000_g N_VPWR_M1000_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.3654 PD=1.54 PS=3.1 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2 SB=75002.9
+ A=0.189 P=2.82 MULT=1
MM1003 N_X_M1000_d N_A_80_23#_M1003_g N_VPWR_M1003_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.43785 PD=1.54 PS=1.955 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75002.5 A=0.189 P=2.82 MULT=1
MM1010 A_386_367# N_B1_M1010_g N_VPWR_M1003_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1323 AS=0.43785 PD=1.47 PS=1.955 NRD=7.8012 NRS=0 M=1 R=8.4 SA=75001.5
+ SB=75001.6 A=0.189 P=2.82 MULT=1
MM1011 N_A_80_23#_M1011_d N_B2_M1011_g A_386_367# VPB PHIGHVT L=0.15 W=1.26
+ AD=0.2457 AS=0.1323 PD=1.65 PS=1.47 NRD=7.8012 NRS=7.8012 M=1 R=8.4 SA=75001.9
+ SB=75001.3 A=0.189 P=2.82 MULT=1
MM1004 A_566_367# N_A2_M1004_g N_A_80_23#_M1011_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.25515 AS=0.2457 PD=1.665 PS=1.65 NRD=23.049 NRS=9.3772 M=1 R=8.4
+ SA=75002.4 SB=75000.7 A=0.189 P=2.82 MULT=1
MM1006 N_VPWR_M1006_d N_A1_M1006_g A_566_367# VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.25515 PD=3.05 PS=1.665 NRD=0 NRS=23.049 M=1 R=8.4 SA=75002.9
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX12_noxref VNB VPB NWDIODE A=7.8703 P=12.17
c_62 VPB 0 5.82976e-20 $X=0 $Y=3.085
*
.include "sky130_fd_sc_lp__o22a_2.pxi.spice"
*
.ends
*
*
