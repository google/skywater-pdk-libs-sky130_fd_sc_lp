* File: sky130_fd_sc_lp__o41a_lp.pxi.spice
* Created: Fri Aug 28 11:19:43 2020
* 
x_PM_SKY130_FD_SC_LP__O41A_LP%A1 N_A1_M1008_g N_A1_M1002_g N_A1_c_88_n
+ N_A1_c_93_n A1 N_A1_c_89_n N_A1_c_90_n PM_SKY130_FD_SC_LP__O41A_LP%A1
x_PM_SKY130_FD_SC_LP__O41A_LP%A2 N_A2_M1010_g N_A2_M1003_g N_A2_c_123_n
+ N_A2_c_128_n A2 A2 A2 A2 N_A2_c_124_n N_A2_c_125_n
+ PM_SKY130_FD_SC_LP__O41A_LP%A2
x_PM_SKY130_FD_SC_LP__O41A_LP%A3 N_A3_M1000_g N_A3_M1007_g N_A3_c_169_n
+ N_A3_c_174_n A3 A3 A3 A3 N_A3_c_170_n N_A3_c_171_n
+ PM_SKY130_FD_SC_LP__O41A_LP%A3
x_PM_SKY130_FD_SC_LP__O41A_LP%A4 N_A4_M1009_g N_A4_M1004_g N_A4_c_210_n
+ N_A4_c_211_n N_A4_c_212_n N_A4_c_213_n N_A4_c_218_n A4 A4 A4 A4 N_A4_c_214_n
+ N_A4_c_215_n PM_SKY130_FD_SC_LP__O41A_LP%A4
x_PM_SKY130_FD_SC_LP__O41A_LP%B1 N_B1_c_264_n N_B1_M1011_g N_B1_c_265_n
+ N_B1_c_266_n N_B1_M1012_g N_B1_c_267_n B1 PM_SKY130_FD_SC_LP__O41A_LP%B1
x_PM_SKY130_FD_SC_LP__O41A_LP%A_457_412# N_A_457_412#_M1011_d
+ N_A_457_412#_M1004_d N_A_457_412#_M1006_g N_A_457_412#_M1005_g
+ N_A_457_412#_M1001_g N_A_457_412#_c_321_n N_A_457_412#_c_329_n
+ N_A_457_412#_c_322_n N_A_457_412#_c_330_n N_A_457_412#_c_323_n
+ N_A_457_412#_c_324_n N_A_457_412#_c_331_n N_A_457_412#_c_332_n
+ N_A_457_412#_c_362_n N_A_457_412#_c_325_n N_A_457_412#_c_326_n
+ N_A_457_412#_c_327_n PM_SKY130_FD_SC_LP__O41A_LP%A_457_412#
x_PM_SKY130_FD_SC_LP__O41A_LP%VPWR N_VPWR_M1008_s N_VPWR_M1012_d N_VPWR_c_404_n
+ N_VPWR_c_405_n N_VPWR_c_406_n VPWR N_VPWR_c_407_n N_VPWR_c_408_n
+ N_VPWR_c_403_n N_VPWR_c_410_n PM_SKY130_FD_SC_LP__O41A_LP%VPWR
x_PM_SKY130_FD_SC_LP__O41A_LP%X N_X_M1001_d N_X_M1005_d X X X X X X X X
+ PM_SKY130_FD_SC_LP__O41A_LP%X
x_PM_SKY130_FD_SC_LP__O41A_LP%A_31_57# N_A_31_57#_M1002_s N_A_31_57#_M1003_d
+ N_A_31_57#_M1009_d N_A_31_57#_c_473_n N_A_31_57#_c_474_n N_A_31_57#_c_475_n
+ N_A_31_57#_c_476_n N_A_31_57#_c_477_n N_A_31_57#_c_478_n N_A_31_57#_c_479_n
+ PM_SKY130_FD_SC_LP__O41A_LP%A_31_57#
x_PM_SKY130_FD_SC_LP__O41A_LP%VGND N_VGND_M1002_d N_VGND_M1000_d N_VGND_M1006_s
+ N_VGND_c_527_n N_VGND_c_528_n N_VGND_c_529_n N_VGND_c_530_n VGND
+ N_VGND_c_531_n N_VGND_c_532_n N_VGND_c_533_n N_VGND_c_534_n N_VGND_c_535_n
+ N_VGND_c_536_n PM_SKY130_FD_SC_LP__O41A_LP%VGND
cc_1 VNB N_A1_M1002_g 0.0500794f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=0.495
cc_2 VNB N_A1_c_88_n 0.0224878f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.695
cc_3 VNB N_A1_c_89_n 0.0172544f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.355
cc_4 VNB N_A1_c_90_n 0.0253335f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.355
cc_5 VNB N_A2_M1003_g 0.0407224f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=0.495
cc_6 VNB N_A2_c_123_n 0.0166972f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.695
cc_7 VNB N_A2_c_124_n 0.015746f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A2_c_125_n 0.0049996f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A3_M1000_g 0.040155f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=2.56
cc_10 VNB N_A3_c_169_n 0.0179815f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.695
cc_11 VNB N_A3_c_170_n 0.0165643f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A3_c_171_n 0.00171403f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A4_c_210_n 0.0149537f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.19
cc_14 VNB N_A4_c_211_n 0.0115256f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.695
cc_15 VNB N_A4_c_212_n 0.0179575f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_16 VNB N_A4_c_213_n 0.0195436f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A4_c_214_n 0.0169915f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A4_c_215_n 0.00230296f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_B1_c_264_n 0.0179956f $X=-0.19 $Y=-0.245 $X2=0.56 $Y2=1.86
cc_20 VNB N_B1_c_265_n 0.0165072f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=1.19
cc_21 VNB N_B1_c_266_n 0.0440058f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=0.495
cc_22 VNB N_B1_c_267_n 0.031215f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.86
cc_23 VNB B1 0.00975793f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_457_412#_M1006_g 0.0406459f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.355
cc_25 VNB N_A_457_412#_M1001_g 0.0405641f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.355
cc_26 VNB N_A_457_412#_c_321_n 0.0219298f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.525
cc_27 VNB N_A_457_412#_c_322_n 0.00827128f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_457_412#_c_323_n 0.0184519f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_457_412#_c_324_n 0.00660311f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_457_412#_c_325_n 0.00121962f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_457_412#_c_326_n 0.026785f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_457_412#_c_327_n 0.00148984f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VPWR_c_403_n 0.183584f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB X 0.0182758f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=0.495
cc_35 VNB X 0.0502536f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_31_57#_c_473_n 0.024646f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.86
cc_37 VNB N_A_31_57#_c_474_n 0.0148956f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_31_57#_c_475_n 0.0103497f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.355
cc_39 VNB N_A_31_57#_c_476_n 0.00354044f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.525
cc_40 VNB N_A_31_57#_c_477_n 0.0163504f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_31_57#_c_478_n 0.0028297f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_31_57#_c_479_n 0.00832431f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_527_n 0.00712794f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_528_n 0.0188675f $X=-0.19 $Y=-0.245 $X2=0.52 $Y2=1.355
cc_45 VNB N_VGND_c_529_n 0.00651282f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_530_n 0.00687099f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_531_n 0.0318541f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_532_n 0.0268694f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_533_n 0.249f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_534_n 0.0259899f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_535_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_536_n 0.00513431f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VPB N_A1_M1008_g 0.0354235f $X=-0.19 $Y=1.655 $X2=0.56 $Y2=2.56
cc_54 VPB N_A1_c_88_n 0.00293319f $X=-0.19 $Y=1.655 $X2=0.52 $Y2=1.695
cc_55 VPB N_A1_c_93_n 0.0144588f $X=-0.19 $Y=1.655 $X2=0.52 $Y2=1.86
cc_56 VPB N_A1_c_90_n 0.0123187f $X=-0.19 $Y=1.655 $X2=0.52 $Y2=1.355
cc_57 VPB N_A2_M1010_g 0.0251795f $X=-0.19 $Y=1.655 $X2=0.56 $Y2=2.56
cc_58 VPB N_A2_c_123_n 0.00509297f $X=-0.19 $Y=1.655 $X2=0.52 $Y2=1.695
cc_59 VPB N_A2_c_128_n 0.0129268f $X=-0.19 $Y=1.655 $X2=0.52 $Y2=1.86
cc_60 VPB N_A2_c_125_n 0.00252273f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_61 VPB N_A3_M1007_g 0.0257022f $X=-0.19 $Y=1.655 $X2=0.515 $Y2=0.495
cc_62 VPB N_A3_c_169_n 0.00548472f $X=-0.19 $Y=1.655 $X2=0.52 $Y2=1.695
cc_63 VPB N_A3_c_174_n 0.0137104f $X=-0.19 $Y=1.655 $X2=0.52 $Y2=1.86
cc_64 VPB N_A3_c_171_n 0.00105896f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_65 VPB N_A4_M1004_g 0.0277199f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_66 VPB N_A4_c_213_n 0.0061492f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_67 VPB N_A4_c_218_n 0.015037f $X=-0.19 $Y=1.655 $X2=0.52 $Y2=1.355
cc_68 VPB N_A4_c_215_n 0.00117171f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_69 VPB N_B1_c_266_n 0.0034244f $X=-0.19 $Y=1.655 $X2=0.515 $Y2=0.495
cc_70 VPB N_B1_M1012_g 0.0402341f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_71 VPB N_A_457_412#_M1005_g 0.0337892f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_72 VPB N_A_457_412#_c_329_n 0.0174306f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_73 VPB N_A_457_412#_c_330_n 0.00452152f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_74 VPB N_A_457_412#_c_331_n 0.0143099f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_75 VPB N_A_457_412#_c_332_n 0.00807345f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_76 VPB N_A_457_412#_c_326_n 0.00223641f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_77 VPB N_VPWR_c_404_n 0.0117216f $X=-0.19 $Y=1.655 $X2=0.515 $Y2=0.495
cc_78 VPB N_VPWR_c_405_n 0.0459728f $X=-0.19 $Y=1.655 $X2=0.52 $Y2=1.355
cc_79 VPB N_VPWR_c_406_n 0.00692321f $X=-0.19 $Y=1.655 $X2=0.52 $Y2=1.355
cc_80 VPB N_VPWR_c_407_n 0.0716193f $X=-0.19 $Y=1.655 $X2=0.52 $Y2=1.525
cc_81 VPB N_VPWR_c_408_n 0.0268044f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_82 VPB N_VPWR_c_403_n 0.0907643f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_83 VPB N_VPWR_c_410_n 0.0053738f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_84 VPB X 0.0203786f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_85 VPB X 0.0165209f $X=-0.19 $Y=1.655 $X2=0.52 $Y2=1.695
cc_86 VPB X 0.0390027f $X=-0.19 $Y=1.655 $X2=0.52 $Y2=1.86
cc_87 N_A1_M1008_g N_A2_M1010_g 0.0264321f $X=0.56 $Y=2.56 $X2=0 $Y2=0
cc_88 N_A1_M1002_g N_A2_M1003_g 0.0241928f $X=0.515 $Y=0.495 $X2=0 $Y2=0
cc_89 N_A1_c_89_n N_A2_M1003_g 0.00127629f $X=0.52 $Y=1.355 $X2=0 $Y2=0
cc_90 N_A1_c_90_n N_A2_M1003_g 2.28806e-19 $X=0.52 $Y=1.355 $X2=0 $Y2=0
cc_91 N_A1_c_88_n N_A2_c_123_n 0.0264321f $X=0.52 $Y=1.695 $X2=0 $Y2=0
cc_92 N_A1_c_93_n N_A2_c_128_n 0.0264321f $X=0.52 $Y=1.86 $X2=0 $Y2=0
cc_93 N_A1_c_89_n N_A2_c_124_n 0.0264321f $X=0.52 $Y=1.355 $X2=0 $Y2=0
cc_94 N_A1_c_90_n N_A2_c_124_n 0.00230645f $X=0.52 $Y=1.355 $X2=0 $Y2=0
cc_95 N_A1_c_93_n N_A2_c_125_n 0.00461461f $X=0.52 $Y=1.86 $X2=0 $Y2=0
cc_96 N_A1_c_89_n N_A2_c_125_n 8.00194e-19 $X=0.52 $Y=1.355 $X2=0 $Y2=0
cc_97 N_A1_c_90_n N_A2_c_125_n 0.0378235f $X=0.52 $Y=1.355 $X2=0 $Y2=0
cc_98 N_A1_M1008_g N_VPWR_c_405_n 0.0258359f $X=0.56 $Y=2.56 $X2=0 $Y2=0
cc_99 N_A1_c_93_n N_VPWR_c_405_n 0.00213543f $X=0.52 $Y=1.86 $X2=0 $Y2=0
cc_100 N_A1_c_90_n N_VPWR_c_405_n 0.0287632f $X=0.52 $Y=1.355 $X2=0 $Y2=0
cc_101 N_A1_M1008_g N_VPWR_c_407_n 0.00823892f $X=0.56 $Y=2.56 $X2=0 $Y2=0
cc_102 N_A1_M1008_g N_VPWR_c_403_n 0.0143247f $X=0.56 $Y=2.56 $X2=0 $Y2=0
cc_103 N_A1_M1002_g N_A_31_57#_c_473_n 0.0117966f $X=0.515 $Y=0.495 $X2=0 $Y2=0
cc_104 N_A1_M1002_g N_A_31_57#_c_474_n 0.00942811f $X=0.515 $Y=0.495 $X2=0 $Y2=0
cc_105 N_A1_c_89_n N_A_31_57#_c_474_n 0.00248655f $X=0.52 $Y=1.355 $X2=0 $Y2=0
cc_106 N_A1_c_90_n N_A_31_57#_c_474_n 0.0162345f $X=0.52 $Y=1.355 $X2=0 $Y2=0
cc_107 N_A1_M1002_g N_A_31_57#_c_475_n 0.00420809f $X=0.515 $Y=0.495 $X2=0 $Y2=0
cc_108 N_A1_c_89_n N_A_31_57#_c_475_n 0.00227085f $X=0.52 $Y=1.355 $X2=0 $Y2=0
cc_109 N_A1_c_90_n N_A_31_57#_c_475_n 0.0289101f $X=0.52 $Y=1.355 $X2=0 $Y2=0
cc_110 N_A1_M1002_g N_A_31_57#_c_476_n 8.89782e-19 $X=0.515 $Y=0.495 $X2=0 $Y2=0
cc_111 N_A1_M1002_g N_VGND_c_527_n 0.00520075f $X=0.515 $Y=0.495 $X2=0 $Y2=0
cc_112 N_A1_M1002_g N_VGND_c_533_n 0.00658755f $X=0.515 $Y=0.495 $X2=0 $Y2=0
cc_113 N_A1_M1002_g N_VGND_c_534_n 0.00502664f $X=0.515 $Y=0.495 $X2=0 $Y2=0
cc_114 N_A2_M1003_g N_A3_M1000_g 0.0271092f $X=1.105 $Y=0.495 $X2=0 $Y2=0
cc_115 N_A2_M1010_g N_A3_M1007_g 0.0489607f $X=1.05 $Y=2.56 $X2=0 $Y2=0
cc_116 N_A2_c_123_n N_A3_c_169_n 0.0117523f $X=1.09 $Y=1.735 $X2=0 $Y2=0
cc_117 N_A2_c_128_n N_A3_c_174_n 0.0117523f $X=1.09 $Y=1.9 $X2=0 $Y2=0
cc_118 N_A2_c_124_n N_A3_c_170_n 0.0117523f $X=1.09 $Y=1.395 $X2=0 $Y2=0
cc_119 N_A2_c_125_n N_A3_c_170_n 0.0109318f $X=1.09 $Y=1.395 $X2=0 $Y2=0
cc_120 N_A2_M1010_g N_A3_c_171_n 0.00101253f $X=1.05 $Y=2.56 $X2=0 $Y2=0
cc_121 N_A2_c_124_n N_A3_c_171_n 7.56445e-19 $X=1.09 $Y=1.395 $X2=0 $Y2=0
cc_122 N_A2_c_125_n N_A3_c_171_n 0.126121f $X=1.09 $Y=1.395 $X2=0 $Y2=0
cc_123 N_A2_M1010_g N_VPWR_c_405_n 0.00367874f $X=1.05 $Y=2.56 $X2=0 $Y2=0
cc_124 N_A2_c_125_n N_VPWR_c_405_n 0.0285381f $X=1.09 $Y=1.395 $X2=0 $Y2=0
cc_125 N_A2_M1010_g N_VPWR_c_407_n 0.00613785f $X=1.05 $Y=2.56 $X2=0 $Y2=0
cc_126 N_A2_c_125_n N_VPWR_c_407_n 0.0110411f $X=1.09 $Y=1.395 $X2=0 $Y2=0
cc_127 N_A2_M1010_g N_VPWR_c_403_n 0.00787277f $X=1.05 $Y=2.56 $X2=0 $Y2=0
cc_128 N_A2_c_125_n N_VPWR_c_403_n 0.0122875f $X=1.09 $Y=1.395 $X2=0 $Y2=0
cc_129 N_A2_c_125_n A_235_412# 0.00844609f $X=1.09 $Y=1.395 $X2=-0.19 $Y2=-0.245
cc_130 N_A2_M1003_g N_A_31_57#_c_473_n 8.89782e-19 $X=1.105 $Y=0.495 $X2=0 $Y2=0
cc_131 N_A2_M1003_g N_A_31_57#_c_474_n 0.00961978f $X=1.105 $Y=0.495 $X2=0 $Y2=0
cc_132 N_A2_c_124_n N_A_31_57#_c_474_n 6.85766e-19 $X=1.09 $Y=1.395 $X2=0 $Y2=0
cc_133 N_A2_c_125_n N_A_31_57#_c_474_n 0.0145508f $X=1.09 $Y=1.395 $X2=0 $Y2=0
cc_134 N_A2_M1003_g N_A_31_57#_c_476_n 0.0101544f $X=1.105 $Y=0.495 $X2=0 $Y2=0
cc_135 N_A2_M1003_g N_A_31_57#_c_479_n 0.00430621f $X=1.105 $Y=0.495 $X2=0 $Y2=0
cc_136 N_A2_c_124_n N_A_31_57#_c_479_n 5.82966e-19 $X=1.09 $Y=1.395 $X2=0 $Y2=0
cc_137 N_A2_c_125_n N_A_31_57#_c_479_n 0.0137298f $X=1.09 $Y=1.395 $X2=0 $Y2=0
cc_138 N_A2_M1003_g N_VGND_c_527_n 0.00520075f $X=1.105 $Y=0.495 $X2=0 $Y2=0
cc_139 N_A2_M1003_g N_VGND_c_528_n 0.00502664f $X=1.105 $Y=0.495 $X2=0 $Y2=0
cc_140 N_A2_M1003_g N_VGND_c_533_n 0.00599173f $X=1.105 $Y=0.495 $X2=0 $Y2=0
cc_141 N_A3_M1007_g N_A4_M1004_g 0.0556338f $X=1.62 $Y=2.56 $X2=0 $Y2=0
cc_142 N_A3_c_171_n N_A4_M1004_g 0.00638395f $X=1.66 $Y=1.395 $X2=0 $Y2=0
cc_143 N_A3_M1000_g N_A4_c_210_n 0.0137654f $X=1.57 $Y=0.495 $X2=0 $Y2=0
cc_144 N_A3_M1000_g N_A4_c_212_n 0.0101786f $X=1.57 $Y=0.495 $X2=0 $Y2=0
cc_145 N_A3_c_169_n N_A4_c_213_n 0.0135694f $X=1.66 $Y=1.735 $X2=0 $Y2=0
cc_146 N_A3_c_174_n N_A4_c_218_n 0.0135694f $X=1.66 $Y=1.9 $X2=0 $Y2=0
cc_147 N_A3_c_170_n N_A4_c_214_n 0.0135694f $X=1.66 $Y=1.395 $X2=0 $Y2=0
cc_148 N_A3_c_171_n N_A4_c_214_n 0.00232658f $X=1.66 $Y=1.395 $X2=0 $Y2=0
cc_149 N_A3_M1007_g N_A4_c_215_n 0.00111514f $X=1.62 $Y=2.56 $X2=0 $Y2=0
cc_150 N_A3_c_170_n N_A4_c_215_n 0.00232658f $X=1.66 $Y=1.395 $X2=0 $Y2=0
cc_151 N_A3_c_171_n N_A4_c_215_n 0.10788f $X=1.66 $Y=1.395 $X2=0 $Y2=0
cc_152 N_A3_M1007_g N_VPWR_c_407_n 0.00613785f $X=1.62 $Y=2.56 $X2=0 $Y2=0
cc_153 N_A3_c_171_n N_VPWR_c_407_n 0.00914393f $X=1.66 $Y=1.395 $X2=0 $Y2=0
cc_154 N_A3_M1007_g N_VPWR_c_403_n 0.00797423f $X=1.62 $Y=2.56 $X2=0 $Y2=0
cc_155 N_A3_c_171_n N_VPWR_c_403_n 0.0101955f $X=1.66 $Y=1.395 $X2=0 $Y2=0
cc_156 N_A3_c_171_n A_349_412# 0.00811515f $X=1.66 $Y=1.395 $X2=-0.19 $Y2=-0.245
cc_157 N_A3_M1000_g N_A_31_57#_c_476_n 0.00241057f $X=1.57 $Y=0.495 $X2=0 $Y2=0
cc_158 N_A3_M1000_g N_A_31_57#_c_477_n 0.0156948f $X=1.57 $Y=0.495 $X2=0 $Y2=0
cc_159 N_A3_c_170_n N_A_31_57#_c_477_n 0.00123061f $X=1.66 $Y=1.395 $X2=0 $Y2=0
cc_160 N_A3_c_171_n N_A_31_57#_c_477_n 0.0245349f $X=1.66 $Y=1.395 $X2=0 $Y2=0
cc_161 N_A3_M1000_g N_A_31_57#_c_478_n 6.68475e-19 $X=1.57 $Y=0.495 $X2=0 $Y2=0
cc_162 N_A3_M1000_g N_A_31_57#_c_479_n 7.06433e-19 $X=1.57 $Y=0.495 $X2=0 $Y2=0
cc_163 N_A3_M1000_g N_VGND_c_528_n 0.0053602f $X=1.57 $Y=0.495 $X2=0 $Y2=0
cc_164 N_A3_M1000_g N_VGND_c_529_n 0.00293322f $X=1.57 $Y=0.495 $X2=0 $Y2=0
cc_165 N_A3_M1000_g N_VGND_c_533_n 0.0103767f $X=1.57 $Y=0.495 $X2=0 $Y2=0
cc_166 N_A4_c_210_n N_B1_c_264_n 0.0104142f $X=2.077 $Y=0.78 $X2=-0.19
+ $Y2=-0.245
cc_167 N_A4_c_212_n N_B1_c_265_n 0.00733432f $X=2.2 $Y=1.23 $X2=0 $Y2=0
cc_168 N_A4_c_213_n N_B1_c_266_n 0.00448348f $X=2.2 $Y=1.735 $X2=0 $Y2=0
cc_169 N_A4_c_214_n N_B1_c_266_n 0.0110836f $X=2.2 $Y=1.395 $X2=0 $Y2=0
cc_170 N_A4_c_215_n N_B1_c_266_n 0.00155096f $X=2.2 $Y=1.395 $X2=0 $Y2=0
cc_171 N_A4_M1004_g N_B1_M1012_g 0.0129327f $X=2.16 $Y=2.56 $X2=0 $Y2=0
cc_172 N_A4_c_218_n N_B1_M1012_g 0.00448348f $X=2.2 $Y=1.9 $X2=0 $Y2=0
cc_173 N_A4_c_215_n N_B1_M1012_g 0.00159783f $X=2.2 $Y=1.395 $X2=0 $Y2=0
cc_174 N_A4_c_211_n N_B1_c_267_n 0.00911908f $X=2.077 $Y=0.93 $X2=0 $Y2=0
cc_175 N_A4_c_212_n B1 2.60965e-19 $X=2.2 $Y=1.23 $X2=0 $Y2=0
cc_176 N_A4_c_214_n B1 0.00110872f $X=2.2 $Y=1.395 $X2=0 $Y2=0
cc_177 N_A4_c_215_n B1 0.0136965f $X=2.2 $Y=1.395 $X2=0 $Y2=0
cc_178 N_A4_c_215_n N_A_457_412#_M1004_d 0.00847063f $X=2.2 $Y=1.395 $X2=0 $Y2=0
cc_179 N_A4_c_210_n N_A_457_412#_c_322_n 2.09694e-19 $X=2.077 $Y=0.78 $X2=0
+ $Y2=0
cc_180 N_A4_M1004_g N_A_457_412#_c_330_n 0.00770847f $X=2.16 $Y=2.56 $X2=0 $Y2=0
cc_181 N_A4_c_218_n N_A_457_412#_c_330_n 3.54793e-19 $X=2.2 $Y=1.9 $X2=0 $Y2=0
cc_182 N_A4_c_215_n N_A_457_412#_c_330_n 0.0795921f $X=2.2 $Y=1.395 $X2=0 $Y2=0
cc_183 N_A4_c_212_n N_A_457_412#_c_324_n 2.22755e-19 $X=2.2 $Y=1.23 $X2=0 $Y2=0
cc_184 N_A4_c_213_n N_A_457_412#_c_332_n 0.0016013f $X=2.2 $Y=1.735 $X2=0 $Y2=0
cc_185 N_A4_c_215_n N_A_457_412#_c_332_n 0.0136967f $X=2.2 $Y=1.395 $X2=0 $Y2=0
cc_186 N_A4_M1004_g N_VPWR_c_407_n 0.00613785f $X=2.16 $Y=2.56 $X2=0 $Y2=0
cc_187 N_A4_c_215_n N_VPWR_c_407_n 0.00914393f $X=2.2 $Y=1.395 $X2=0 $Y2=0
cc_188 N_A4_M1004_g N_VPWR_c_403_n 0.00833758f $X=2.16 $Y=2.56 $X2=0 $Y2=0
cc_189 N_A4_c_215_n N_VPWR_c_403_n 0.0101955f $X=2.2 $Y=1.395 $X2=0 $Y2=0
cc_190 N_A4_c_211_n N_A_31_57#_c_477_n 0.00851489f $X=2.077 $Y=0.93 $X2=0 $Y2=0
cc_191 N_A4_c_212_n N_A_31_57#_c_477_n 0.00697084f $X=2.2 $Y=1.23 $X2=0 $Y2=0
cc_192 N_A4_c_214_n N_A_31_57#_c_477_n 0.00124283f $X=2.2 $Y=1.395 $X2=0 $Y2=0
cc_193 N_A4_c_215_n N_A_31_57#_c_477_n 0.0251906f $X=2.2 $Y=1.395 $X2=0 $Y2=0
cc_194 N_A4_c_210_n N_A_31_57#_c_478_n 0.00734944f $X=2.077 $Y=0.78 $X2=0 $Y2=0
cc_195 N_A4_c_211_n N_A_31_57#_c_478_n 0.00455806f $X=2.077 $Y=0.93 $X2=0 $Y2=0
cc_196 N_A4_c_210_n N_VGND_c_529_n 0.00275065f $X=2.077 $Y=0.78 $X2=0 $Y2=0
cc_197 N_A4_c_210_n N_VGND_c_531_n 0.00502664f $X=2.077 $Y=0.78 $X2=0 $Y2=0
cc_198 N_A4_c_210_n N_VGND_c_533_n 0.00952614f $X=2.077 $Y=0.78 $X2=0 $Y2=0
cc_199 N_B1_c_266_n N_A_457_412#_M1006_g 0.0114154f $X=2.975 $Y=1.705 $X2=0
+ $Y2=0
cc_200 N_B1_c_267_n N_A_457_412#_M1006_g 0.00720445f $X=2.745 $Y=0.855 $X2=0
+ $Y2=0
cc_201 B1 N_A_457_412#_M1006_g 0.00291824f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_202 N_B1_M1012_g N_A_457_412#_M1005_g 0.022205f $X=2.975 $Y=2.56 $X2=0 $Y2=0
cc_203 N_B1_M1012_g N_A_457_412#_c_329_n 0.00630933f $X=2.975 $Y=2.56 $X2=0
+ $Y2=0
cc_204 N_B1_c_264_n N_A_457_412#_c_322_n 0.00801512f $X=2.475 $Y=0.78 $X2=0
+ $Y2=0
cc_205 N_B1_c_267_n N_A_457_412#_c_322_n 0.00831754f $X=2.745 $Y=0.855 $X2=0
+ $Y2=0
cc_206 N_B1_M1012_g N_A_457_412#_c_330_n 0.0246139f $X=2.975 $Y=2.56 $X2=0 $Y2=0
cc_207 N_B1_c_266_n N_A_457_412#_c_323_n 0.00379299f $X=2.975 $Y=1.705 $X2=0
+ $Y2=0
cc_208 B1 N_A_457_412#_c_323_n 0.0282986f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_209 N_B1_c_265_n N_A_457_412#_c_324_n 0.00528764f $X=2.745 $Y=1.18 $X2=0
+ $Y2=0
cc_210 N_B1_c_266_n N_A_457_412#_c_324_n 8.30838e-19 $X=2.975 $Y=1.705 $X2=0
+ $Y2=0
cc_211 N_B1_c_267_n N_A_457_412#_c_324_n 0.00774343f $X=2.745 $Y=0.855 $X2=0
+ $Y2=0
cc_212 B1 N_A_457_412#_c_324_n 0.0142614f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_213 N_B1_c_266_n N_A_457_412#_c_331_n 0.0030484f $X=2.975 $Y=1.705 $X2=0
+ $Y2=0
cc_214 N_B1_M1012_g N_A_457_412#_c_331_n 0.0142636f $X=2.975 $Y=2.56 $X2=0 $Y2=0
cc_215 B1 N_A_457_412#_c_331_n 0.0260084f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_216 N_B1_c_266_n N_A_457_412#_c_332_n 0.00538223f $X=2.975 $Y=1.705 $X2=0
+ $Y2=0
cc_217 N_B1_M1012_g N_A_457_412#_c_332_n 0.00257798f $X=2.975 $Y=2.56 $X2=0
+ $Y2=0
cc_218 B1 N_A_457_412#_c_332_n 0.0164462f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_219 N_B1_c_266_n N_A_457_412#_c_362_n 0.00107073f $X=2.975 $Y=1.705 $X2=0
+ $Y2=0
cc_220 N_B1_c_266_n N_A_457_412#_c_326_n 0.00630933f $X=2.975 $Y=1.705 $X2=0
+ $Y2=0
cc_221 N_B1_c_265_n N_A_457_412#_c_327_n 8.81901e-19 $X=2.745 $Y=1.18 $X2=0
+ $Y2=0
cc_222 N_B1_c_266_n N_A_457_412#_c_327_n 2.85461e-19 $X=2.975 $Y=1.705 $X2=0
+ $Y2=0
cc_223 B1 N_A_457_412#_c_327_n 0.0259555f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_224 N_B1_M1012_g N_VPWR_c_406_n 0.0239184f $X=2.975 $Y=2.56 $X2=0 $Y2=0
cc_225 N_B1_M1012_g N_VPWR_c_407_n 0.00789732f $X=2.975 $Y=2.56 $X2=0 $Y2=0
cc_226 N_B1_M1012_g N_VPWR_c_403_n 0.013957f $X=2.975 $Y=2.56 $X2=0 $Y2=0
cc_227 N_B1_M1012_g X 3.10289e-19 $X=2.975 $Y=2.56 $X2=0 $Y2=0
cc_228 N_B1_c_265_n N_A_31_57#_c_477_n 0.00145769f $X=2.745 $Y=1.18 $X2=0 $Y2=0
cc_229 N_B1_c_267_n N_A_31_57#_c_477_n 4.12917e-19 $X=2.745 $Y=0.855 $X2=0 $Y2=0
cc_230 N_B1_c_264_n N_A_31_57#_c_478_n 0.0015556f $X=2.475 $Y=0.78 $X2=0 $Y2=0
cc_231 N_B1_c_264_n N_VGND_c_530_n 0.00258896f $X=2.475 $Y=0.78 $X2=0 $Y2=0
cc_232 N_B1_c_264_n N_VGND_c_531_n 0.00502664f $X=2.475 $Y=0.78 $X2=0 $Y2=0
cc_233 N_B1_c_267_n N_VGND_c_531_n 5.79469e-19 $X=2.745 $Y=0.855 $X2=0 $Y2=0
cc_234 N_B1_c_264_n N_VGND_c_533_n 0.010456f $X=2.475 $Y=0.78 $X2=0 $Y2=0
cc_235 N_A_457_412#_M1005_g N_VPWR_c_406_n 0.0142714f $X=3.62 $Y=2.56 $X2=0
+ $Y2=0
cc_236 N_A_457_412#_c_329_n N_VPWR_c_406_n 3.79157e-19 $X=3.567 $Y=1.86 $X2=0
+ $Y2=0
cc_237 N_A_457_412#_c_330_n N_VPWR_c_406_n 0.067538f $X=2.71 $Y=2.205 $X2=0
+ $Y2=0
cc_238 N_A_457_412#_c_331_n N_VPWR_c_406_n 0.0263485f $X=3.415 $Y=1.775 $X2=0
+ $Y2=0
cc_239 N_A_457_412#_c_330_n N_VPWR_c_407_n 0.0220321f $X=2.71 $Y=2.205 $X2=0
+ $Y2=0
cc_240 N_A_457_412#_M1005_g N_VPWR_c_408_n 0.00883132f $X=3.62 $Y=2.56 $X2=0
+ $Y2=0
cc_241 N_A_457_412#_M1005_g N_VPWR_c_403_n 0.0169736f $X=3.62 $Y=2.56 $X2=0
+ $Y2=0
cc_242 N_A_457_412#_c_330_n N_VPWR_c_403_n 0.0125808f $X=2.71 $Y=2.205 $X2=0
+ $Y2=0
cc_243 N_A_457_412#_M1006_g X 0.00117329f $X=3.465 $Y=0.445 $X2=0 $Y2=0
cc_244 N_A_457_412#_M1001_g X 0.00849951f $X=3.825 $Y=0.445 $X2=0 $Y2=0
cc_245 N_A_457_412#_M1005_g X 0.00640485f $X=3.62 $Y=2.56 $X2=0 $Y2=0
cc_246 N_A_457_412#_M1001_g X 0.0194486f $X=3.825 $Y=0.445 $X2=0 $Y2=0
cc_247 N_A_457_412#_c_329_n X 0.00116864f $X=3.567 $Y=1.86 $X2=0 $Y2=0
cc_248 N_A_457_412#_c_323_n X 0.00837902f $X=3.415 $Y=0.915 $X2=0 $Y2=0
cc_249 N_A_457_412#_c_331_n X 0.0114669f $X=3.415 $Y=1.775 $X2=0 $Y2=0
cc_250 N_A_457_412#_c_325_n X 0.0316948f $X=3.58 $Y=1.355 $X2=0 $Y2=0
cc_251 N_A_457_412#_c_326_n X 0.0077371f $X=3.58 $Y=1.355 $X2=0 $Y2=0
cc_252 N_A_457_412#_c_327_n X 0.0083481f $X=3.58 $Y=1.19 $X2=0 $Y2=0
cc_253 N_A_457_412#_M1005_g X 0.00466064f $X=3.62 $Y=2.56 $X2=0 $Y2=0
cc_254 N_A_457_412#_c_321_n X 0.00435084f $X=3.645 $Y=1.34 $X2=0 $Y2=0
cc_255 N_A_457_412#_c_331_n X 0.00193744f $X=3.415 $Y=1.775 $X2=0 $Y2=0
cc_256 N_A_457_412#_M1005_g X 0.012738f $X=3.62 $Y=2.56 $X2=0 $Y2=0
cc_257 N_A_457_412#_c_324_n N_A_31_57#_c_477_n 0.0105633f $X=2.855 $Y=0.915
+ $X2=0 $Y2=0
cc_258 N_A_457_412#_c_322_n N_A_31_57#_c_478_n 0.0256576f $X=2.69 $Y=0.495 $X2=0
+ $Y2=0
cc_259 N_A_457_412#_c_324_n N_A_31_57#_c_478_n 0.00389608f $X=2.855 $Y=0.915
+ $X2=0 $Y2=0
cc_260 N_A_457_412#_M1006_g N_VGND_c_530_n 0.0133964f $X=3.465 $Y=0.445 $X2=0
+ $Y2=0
cc_261 N_A_457_412#_M1001_g N_VGND_c_530_n 0.0023299f $X=3.825 $Y=0.445 $X2=0
+ $Y2=0
cc_262 N_A_457_412#_c_322_n N_VGND_c_530_n 0.0259561f $X=2.69 $Y=0.495 $X2=0
+ $Y2=0
cc_263 N_A_457_412#_c_323_n N_VGND_c_530_n 0.0227314f $X=3.415 $Y=0.915 $X2=0
+ $Y2=0
cc_264 N_A_457_412#_c_322_n N_VGND_c_531_n 0.0220321f $X=2.69 $Y=0.495 $X2=0
+ $Y2=0
cc_265 N_A_457_412#_M1006_g N_VGND_c_532_n 0.00486043f $X=3.465 $Y=0.445 $X2=0
+ $Y2=0
cc_266 N_A_457_412#_M1001_g N_VGND_c_532_n 0.00549284f $X=3.825 $Y=0.445 $X2=0
+ $Y2=0
cc_267 N_A_457_412#_M1006_g N_VGND_c_533_n 0.00436917f $X=3.465 $Y=0.445 $X2=0
+ $Y2=0
cc_268 N_A_457_412#_M1001_g N_VGND_c_533_n 0.010905f $X=3.825 $Y=0.445 $X2=0
+ $Y2=0
cc_269 N_A_457_412#_c_322_n N_VGND_c_533_n 0.0125808f $X=2.69 $Y=0.495 $X2=0
+ $Y2=0
cc_270 N_A_457_412#_c_323_n N_VGND_c_533_n 0.0149196f $X=3.415 $Y=0.915 $X2=0
+ $Y2=0
cc_271 N_VPWR_c_406_n X 0.0510219f $X=3.24 $Y=2.205 $X2=0 $Y2=0
cc_272 N_VPWR_c_408_n X 0.0324829f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_273 N_VPWR_c_403_n X 0.0185782f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_274 X N_VGND_c_530_n 0.0128811f $X=3.995 $Y=0.47 $X2=0 $Y2=0
cc_275 X N_VGND_c_532_n 0.0197155f $X=3.995 $Y=0.47 $X2=0 $Y2=0
cc_276 N_X_M1001_d N_VGND_c_533_n 0.00232985f $X=3.9 $Y=0.235 $X2=0 $Y2=0
cc_277 X N_VGND_c_533_n 0.0125355f $X=3.995 $Y=0.47 $X2=0 $Y2=0
cc_278 N_A_31_57#_c_473_n N_VGND_c_527_n 0.0149165f $X=0.3 $Y=0.495 $X2=0 $Y2=0
cc_279 N_A_31_57#_c_474_n N_VGND_c_527_n 0.0252399f $X=1.155 $Y=0.925 $X2=0
+ $Y2=0
cc_280 N_A_31_57#_c_476_n N_VGND_c_527_n 0.0149165f $X=1.32 $Y=0.495 $X2=0 $Y2=0
cc_281 N_A_31_57#_c_476_n N_VGND_c_528_n 0.0220321f $X=1.32 $Y=0.495 $X2=0 $Y2=0
cc_282 N_A_31_57#_c_476_n N_VGND_c_529_n 0.00148713f $X=1.32 $Y=0.495 $X2=0
+ $Y2=0
cc_283 N_A_31_57#_c_477_n N_VGND_c_529_n 0.0180776f $X=2.095 $Y=0.965 $X2=0
+ $Y2=0
cc_284 N_A_31_57#_c_478_n N_VGND_c_529_n 0.0156695f $X=2.26 $Y=0.495 $X2=0 $Y2=0
cc_285 N_A_31_57#_c_478_n N_VGND_c_531_n 0.0166382f $X=2.26 $Y=0.495 $X2=0 $Y2=0
cc_286 N_A_31_57#_c_473_n N_VGND_c_533_n 0.0125808f $X=0.3 $Y=0.495 $X2=0 $Y2=0
cc_287 N_A_31_57#_c_474_n N_VGND_c_533_n 0.0117708f $X=1.155 $Y=0.925 $X2=0
+ $Y2=0
cc_288 N_A_31_57#_c_476_n N_VGND_c_533_n 0.0125808f $X=1.32 $Y=0.495 $X2=0 $Y2=0
cc_289 N_A_31_57#_c_478_n N_VGND_c_533_n 0.00948536f $X=2.26 $Y=0.495 $X2=0
+ $Y2=0
cc_290 N_A_31_57#_c_473_n N_VGND_c_534_n 0.0220321f $X=0.3 $Y=0.495 $X2=0 $Y2=0
cc_291 N_VGND_c_533_n A_708_47# 0.00771977f $X=4.08 $Y=0 $X2=-0.19 $Y2=-0.245
