# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_lp__o2111ai_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  10.08000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.925000 1.375000 9.995000 1.760000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.010000 1.355000 7.665000 1.525000 ;
        RECT 7.135000 1.205000 7.665000 1.355000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.945000 1.355000 5.685000 1.750000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.085000 1.325000 3.775000 1.505000 ;
        RECT 3.115000 1.155000 3.775000 1.325000 ;
    END
  END C1
  PIN D1
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.525000 1.335000 1.875000 1.505000 ;
        RECT 0.945000 1.200000 1.685000 1.335000 ;
    END
  END D1
  PIN Y
    ANTENNADIFFAREA  4.036200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.985000 1.685000 1.030000 ;
        RECT 0.085000 1.030000 0.775000 1.155000 ;
        RECT 0.085000 1.155000 0.355000 1.675000 ;
        RECT 0.085000 1.675000 3.775000 1.845000 ;
        RECT 0.085000 1.845000 0.355000 3.075000 ;
        RECT 0.595000 0.700000 1.685000 0.985000 ;
        RECT 1.025000 1.845000 1.215000 3.075000 ;
        RECT 1.885000 1.845000 2.075000 3.075000 ;
        RECT 2.745000 1.845000 2.935000 3.075000 ;
        RECT 3.605000 1.845000 3.775000 1.920000 ;
        RECT 3.605000 1.920000 6.715000 2.100000 ;
        RECT 3.605000 2.100000 4.130000 3.075000 ;
        RECT 4.805000 2.100000 4.995000 3.075000 ;
        RECT 5.665000 2.100000 5.855000 3.075000 ;
        RECT 6.510000 1.705000 7.645000 1.875000 ;
        RECT 6.510000 1.875000 6.715000 1.920000 ;
        RECT 6.525000 2.100000 6.715000 2.725000 ;
        RECT 7.315000 1.875000 7.645000 2.155000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 10.080000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.500000 0.500000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.800000 0.500000 3.300000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 10.080000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 10.080000 0.085000 ;
      RECT 0.000000  3.245000 10.080000 3.415000 ;
      RECT 0.095000  0.255000  2.075000 0.530000 ;
      RECT 0.095000  0.530000  0.425000 0.815000 ;
      RECT 0.525000  2.015000  0.855000 3.245000 ;
      RECT 1.385000  2.015000  1.715000 3.245000 ;
      RECT 1.855000  0.530000  2.075000 0.985000 ;
      RECT 1.855000  0.985000  2.945000 1.155000 ;
      RECT 2.245000  0.255000  5.675000 0.425000 ;
      RECT 2.245000  0.425000  4.815000 0.485000 ;
      RECT 2.245000  0.485000  2.575000 0.815000 ;
      RECT 2.245000  2.015000  2.575000 3.245000 ;
      RECT 2.745000  0.655000  3.805000 0.985000 ;
      RECT 3.105000  2.015000  3.435000 3.245000 ;
      RECT 4.055000  0.655000  4.315000 1.015000 ;
      RECT 4.055000  1.015000  9.905000 1.035000 ;
      RECT 4.055000  1.035000  6.965000 1.185000 ;
      RECT 4.300000  2.270000  4.635000 3.245000 ;
      RECT 4.485000  0.485000  4.815000 0.845000 ;
      RECT 4.985000  0.595000  5.175000 1.015000 ;
      RECT 5.165000  2.270000  5.495000 3.245000 ;
      RECT 5.345000  0.425000  5.675000 0.845000 ;
      RECT 5.845000  0.255000  6.035000 1.015000 ;
      RECT 6.025000  2.270000  6.355000 2.895000 ;
      RECT 6.025000  2.895000  7.215000 3.075000 ;
      RECT 6.205000  0.085000  6.535000 0.845000 ;
      RECT 6.705000  0.255000  6.895000 0.865000 ;
      RECT 6.705000  0.865000  8.115000 1.005000 ;
      RECT 6.705000  1.005000  9.905000 1.015000 ;
      RECT 6.885000  2.045000  7.145000 2.325000 ;
      RECT 6.885000  2.325000  8.525000 2.495000 ;
      RECT 6.885000  2.495000  7.215000 2.895000 ;
      RECT 7.065000  0.085000  7.395000 0.695000 ;
      RECT 7.565000  0.255000  8.115000 0.865000 ;
      RECT 7.835000  1.035000  9.905000 1.175000 ;
      RECT 7.835000  2.665000  8.165000 3.245000 ;
      RECT 8.265000  1.930000  9.385000 2.100000 ;
      RECT 8.265000  2.100000  8.525000 2.325000 ;
      RECT 8.285000  0.085000  8.615000 0.835000 ;
      RECT 8.335000  2.495000  8.525000 3.075000 ;
      RECT 8.695000  2.270000  9.025000 3.245000 ;
      RECT 8.785000  0.255000  8.975000 1.005000 ;
      RECT 9.145000  0.085000  9.475000 0.835000 ;
      RECT 9.195000  2.100000  9.385000 3.075000 ;
      RECT 9.555000  1.930000  9.885000 3.245000 ;
      RECT 9.645000  0.255000  9.905000 1.005000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
      RECT 6.875000 -0.085000 7.045000 0.085000 ;
      RECT 6.875000  3.245000 7.045000 3.415000 ;
      RECT 7.355000 -0.085000 7.525000 0.085000 ;
      RECT 7.355000  3.245000 7.525000 3.415000 ;
      RECT 7.835000 -0.085000 8.005000 0.085000 ;
      RECT 7.835000  3.245000 8.005000 3.415000 ;
      RECT 8.315000 -0.085000 8.485000 0.085000 ;
      RECT 8.315000  3.245000 8.485000 3.415000 ;
      RECT 8.795000 -0.085000 8.965000 0.085000 ;
      RECT 8.795000  3.245000 8.965000 3.415000 ;
      RECT 9.275000 -0.085000 9.445000 0.085000 ;
      RECT 9.275000  3.245000 9.445000 3.415000 ;
      RECT 9.755000 -0.085000 9.925000 0.085000 ;
      RECT 9.755000  3.245000 9.925000 3.415000 ;
  END
END sky130_fd_sc_lp__o2111ai_4
END LIBRARY
