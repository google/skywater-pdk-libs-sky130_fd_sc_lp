* File: sky130_fd_sc_lp__nor4bb_m.pex.spice
* Created: Fri Aug 28 10:59:28 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__NOR4BB_M%D_N 3 7 11 13 14 15 19
c35 7 0 9.48991e-20 $X=0.595 $Y=0.835
r36 19 20 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.385
+ $Y=1.67 $X2=0.385 $Y2=1.67
r37 15 20 13.3537 $w=3.13e-07 $l=3.65e-07 $layer=LI1_cond $X=0.312 $Y=2.035
+ $X2=0.312 $Y2=1.67
r38 14 20 0.182927 $w=3.13e-07 $l=5e-09 $layer=LI1_cond $X=0.312 $Y=1.665
+ $X2=0.312 $Y2=1.67
r39 12 19 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.385 $Y=2.01
+ $X2=0.385 $Y2=1.67
r40 12 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.385 $Y=2.01
+ $X2=0.385 $Y2=2.175
r41 11 19 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=0.385 $Y=1.655
+ $X2=0.385 $Y2=1.67
r42 10 11 43.5886 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=0.445 $Y=1.505
+ $X2=0.445 $Y2=1.655
r43 7 10 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=0.595 $Y=0.835
+ $X2=0.595 $Y2=1.505
r44 3 13 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=0.475 $Y=2.745
+ $X2=0.475 $Y2=2.175
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4BB_M%A_27_507# 1 2 9 10 11 14 17 18 21 25 27 28
+ 30 32 37 38 40
c73 37 0 1.51217e-19 $X=1.045 $Y=1.32
c74 30 0 9.75149e-20 $X=0.89 $Y=1.585
r75 37 38 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.045
+ $Y=1.32 $X2=1.045 $Y2=1.32
r76 32 40 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=0.735 $Y=2.355
+ $X2=0.735 $Y2=1.825
r77 30 40 11.2652 $w=4.78e-07 $l=2.4e-07 $layer=LI1_cond $X=0.89 $Y=1.585
+ $X2=0.89 $Y2=1.825
r78 29 37 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=0.89 $Y=1.24
+ $X2=1.045 $Y2=1.24
r79 29 30 6.47876 $w=4.78e-07 $l=2.6e-07 $layer=LI1_cond $X=0.89 $Y=1.325
+ $X2=0.89 $Y2=1.585
r80 27 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.65 $Y=2.44
+ $X2=0.735 $Y2=2.355
r81 27 28 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.65 $Y=2.44
+ $X2=0.345 $Y2=2.44
r82 23 29 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=0.38 $Y=1.24
+ $X2=0.89 $Y2=1.24
r83 23 25 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=0.38 $Y=1.155
+ $X2=0.38 $Y2=0.9
r84 19 28 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=0.25 $Y=2.525
+ $X2=0.345 $Y2=2.44
r85 19 21 9.04785 $w=1.88e-07 $l=1.55e-07 $layer=LI1_cond $X=0.25 $Y=2.525
+ $X2=0.25 $Y2=2.68
r86 18 38 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=1.045 $Y=1.675
+ $X2=1.045 $Y2=1.32
r87 17 38 38.6168 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.045 $Y=1.155
+ $X2=1.045 $Y2=1.32
r88 12 14 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=1.475 $Y=1.825
+ $X2=1.475 $Y2=2.195
r89 11 18 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=1.21 $Y=1.75
+ $X2=1.045 $Y2=1.675
r90 10 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.4 $Y=1.75
+ $X2=1.475 $Y2=1.825
r91 10 11 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=1.4 $Y=1.75 $X2=1.21
+ $Y2=1.75
r92 9 17 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.065 $Y=0.835
+ $X2=1.065 $Y2=1.155
r93 2 21 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.535 $X2=0.26 $Y2=2.68
r94 1 25 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=0.255
+ $Y=0.625 $X2=0.38 $Y2=0.9
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4BB_M%B 3 5 7 8 12
c34 3 0 1.91377e-19 $X=2.195 $Y=0.835
r35 12 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.175 $Y=0.35
+ $X2=2.175 $Y2=0.515
r36 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.175
+ $Y=0.35 $X2=2.175 $Y2=0.35
r37 8 13 14.2903 $w=3.73e-07 $l=4.65e-07 $layer=LI1_cond $X=2.64 $Y=0.452
+ $X2=2.175 $Y2=0.452
r38 7 13 0.460977 $w=3.73e-07 $l=1.5e-08 $layer=LI1_cond $X=2.16 $Y=0.452
+ $X2=2.175 $Y2=0.452
r39 3 5 697.362 $w=1.5e-07 $l=1.36e-06 $layer=POLY_cond $X=2.195 $Y=0.835
+ $X2=2.195 $Y2=2.195
r40 3 15 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.195 $Y=0.835
+ $X2=2.195 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4BB_M%A 3 7 9 10 11 12 13 17
c32 10 0 1.4009e-19 $X=2.645 $Y=1.66
c33 9 0 1.56674e-19 $X=2.645 $Y=1.155
r34 12 13 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=2.645 $Y=1.295
+ $X2=2.645 $Y2=1.665
r35 12 17 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.645
+ $Y=1.32 $X2=2.645 $Y2=1.32
r36 10 17 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.645 $Y=1.66
+ $X2=2.645 $Y2=1.32
r37 10 11 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.645 $Y=1.66
+ $X2=2.645 $Y2=1.825
r38 9 17 38.6168 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.645 $Y=1.155
+ $X2=2.645 $Y2=1.32
r39 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.625 $Y=0.835
+ $X2=2.625 $Y2=1.155
r40 3 11 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=2.555 $Y=2.195
+ $X2=2.555 $Y2=1.825
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4BB_M%A_284_99# 1 2 9 11 12 16 17 18 19 27 31 33
c58 31 0 1.56674e-19 $X=3.545 $Y=0.87
c59 12 0 1.11779e-19 $X=1.57 $Y=1.36
c60 9 0 1.51217e-19 $X=1.495 $Y=0.835
r61 29 31 6.60173 $w=2.08e-07 $l=1.25e-07 $layer=LI1_cond $X=3.42 $Y=0.87
+ $X2=3.545 $Y2=0.87
r62 25 27 42.3206 $w=1.88e-07 $l=7.25e-07 $layer=LI1_cond $X=3.545 $Y=2.855
+ $X2=3.545 $Y2=2.13
r63 24 31 1.31963 $w=1.9e-07 $l=1.05e-07 $layer=LI1_cond $X=3.545 $Y=0.975
+ $X2=3.545 $Y2=0.87
r64 24 27 67.4211 $w=1.88e-07 $l=1.155e-06 $layer=LI1_cond $X=3.545 $Y=0.975
+ $X2=3.545 $Y2=2.13
r65 22 33 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=3.2 $Y=2.94 $X2=3.2
+ $Y2=2.85
r66 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.2
+ $Y=2.94 $X2=3.2 $Y2=2.94
r67 19 25 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=3.45 $Y=2.94
+ $X2=3.545 $Y2=2.855
r68 19 21 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=3.45 $Y=2.94 $X2=3.2
+ $Y2=2.94
r69 17 33 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.035 $Y=2.85
+ $X2=3.2 $Y2=2.85
r70 17 18 576.862 $w=1.5e-07 $l=1.125e-06 $layer=POLY_cond $X=3.035 $Y=2.85
+ $X2=1.91 $Y2=2.85
r71 14 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.835 $Y=2.775
+ $X2=1.91 $Y2=2.85
r72 14 16 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=1.835 $Y=2.775
+ $X2=1.835 $Y2=2.195
r73 13 16 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=1.835 $Y=1.435
+ $X2=1.835 $Y2=2.195
r74 11 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.76 $Y=1.36
+ $X2=1.835 $Y2=1.435
r75 11 12 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=1.76 $Y=1.36
+ $X2=1.57 $Y2=1.36
r76 7 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.495 $Y=1.285
+ $X2=1.57 $Y2=1.36
r77 7 9 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=1.495 $Y=1.285
+ $X2=1.495 $Y2=0.835
r78 2 27 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=3.395
+ $Y=1.985 $X2=3.535 $Y2=2.13
r79 1 29 182 $w=1.7e-07 $l=3.07124e-07 $layer=licon1_NDIFF $count=1 $X=3.28
+ $Y=0.625 $X2=3.42 $Y2=0.87
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4BB_M%C_N 2 5 8 10 11 12 13 14 20 22
r36 20 22 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=3.207 $Y=1.32
+ $X2=3.207 $Y2=1.155
r37 13 14 18.1448 $w=2.33e-07 $l=3.7e-07 $layer=LI1_cond $X=3.152 $Y=2.035
+ $X2=3.152 $Y2=2.405
r38 12 13 18.1448 $w=2.33e-07 $l=3.7e-07 $layer=LI1_cond $X=3.152 $Y=1.665
+ $X2=3.152 $Y2=2.035
r39 11 12 18.1448 $w=2.33e-07 $l=3.7e-07 $layer=LI1_cond $X=3.152 $Y=1.295
+ $X2=3.152 $Y2=1.665
r40 11 20 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.185
+ $Y=1.32 $X2=3.185 $Y2=1.32
r41 8 10 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=3.32 $Y=2.195
+ $X2=3.32 $Y2=1.825
r42 5 22 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=3.205 $Y=0.835
+ $X2=3.205 $Y2=1.155
r43 2 10 48.4185 $w=3.75e-07 $l=1.87e-07 $layer=POLY_cond $X=3.207 $Y=1.638
+ $X2=3.207 $Y2=1.825
r44 1 20 3.26277 $w=3.75e-07 $l=2.2e-08 $layer=POLY_cond $X=3.207 $Y=1.342
+ $X2=3.207 $Y2=1.32
r45 1 2 43.8991 $w=3.75e-07 $l=2.96e-07 $layer=POLY_cond $X=3.207 $Y=1.342
+ $X2=3.207 $Y2=1.638
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4BB_M%VPWR 1 2 9 13 16 17 18 20 33 34 37
r34 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r35 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r36 31 34 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r37 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r38 28 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r39 27 30 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r40 27 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r41 25 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.855 $Y=3.33
+ $X2=0.69 $Y2=3.33
r42 25 27 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.855 $Y=3.33
+ $X2=1.2 $Y2=3.33
r43 23 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r44 22 23 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r45 20 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.525 $Y=3.33
+ $X2=0.69 $Y2=3.33
r46 20 22 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.525 $Y=3.33
+ $X2=0.24 $Y2=3.33
r47 18 31 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=2.64 $Y2=3.33
r48 18 28 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=1.2 $Y2=3.33
r49 16 30 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=2.665 $Y=3.33
+ $X2=2.64 $Y2=3.33
r50 16 17 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.665 $Y=3.33
+ $X2=2.76 $Y2=3.33
r51 15 33 48.6043 $w=1.68e-07 $l=7.45e-07 $layer=LI1_cond $X=2.855 $Y=3.33
+ $X2=3.6 $Y2=3.33
r52 15 17 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.855 $Y=3.33
+ $X2=2.76 $Y2=3.33
r53 11 17 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=2.76 $Y=3.245
+ $X2=2.76 $Y2=3.33
r54 11 13 56.3301 $w=1.88e-07 $l=9.65e-07 $layer=LI1_cond $X=2.76 $Y=3.245
+ $X2=2.76 $Y2=2.28
r55 7 37 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=3.245 $X2=0.69
+ $Y2=3.33
r56 7 9 15.1913 $w=3.28e-07 $l=4.35e-07 $layer=LI1_cond $X=0.69 $Y=3.245
+ $X2=0.69 $Y2=2.81
r57 2 13 600 $w=1.7e-07 $l=3.58225e-07 $layer=licon1_PDIFF $count=1 $X=2.63
+ $Y=1.985 $X2=2.77 $Y2=2.28
r58 1 9 600 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=2.535 $X2=0.69 $Y2=2.81
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4BB_M%Y 1 2 3 11 13 14 19 24 26 27 32
c58 27 0 2.39111e-20 $X=2.16 $Y=0.925
c59 24 0 1.49601e-19 $X=1.395 $Y=0.87
c60 19 0 1.42641e-20 $X=1.395 $Y=2.13
c61 11 0 1.36675e-19 $X=1.395 $Y=1.115
r62 38 39 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=2.16 $Y=0.93 $X2=2.16
+ $Y2=1.2
r63 27 38 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=2.16 $Y=0.925
+ $X2=2.16 $Y2=0.93
r64 27 38 0.0262452 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=2.245 $Y=0.93
+ $X2=2.16 $Y2=0.93
r65 27 32 7.83854 $w=3.58e-07 $l=1.65e-07 $layer=LI1_cond $X=2.245 $Y=0.93
+ $X2=2.41 $Y2=0.93
r66 22 24 6.07359 $w=2.08e-07 $l=1.15e-07 $layer=LI1_cond $X=1.28 $Y=0.87
+ $X2=1.395 $Y2=0.87
r67 17 19 7.12987 $w=2.08e-07 $l=1.35e-07 $layer=LI1_cond $X=1.26 $Y=2.13
+ $X2=1.395 $Y2=2.13
r68 15 26 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.48 $Y=1.2 $X2=1.395
+ $Y2=1.2
r69 14 39 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.075 $Y=1.2
+ $X2=2.16 $Y2=1.2
r70 14 15 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=2.075 $Y=1.2
+ $X2=1.48 $Y2=1.2
r71 13 19 1.9771 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.395 $Y=2.025
+ $X2=1.395 $Y2=2.13
r72 12 26 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.395 $Y=1.285
+ $X2=1.395 $Y2=1.2
r73 12 13 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=1.395 $Y=1.285
+ $X2=1.395 $Y2=2.025
r74 11 26 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.395 $Y=1.115
+ $X2=1.395 $Y2=1.2
r75 10 24 1.9771 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.395 $Y=0.975
+ $X2=1.395 $Y2=0.87
r76 10 11 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=1.395 $Y=0.975
+ $X2=1.395 $Y2=1.115
r77 3 17 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=1.135
+ $Y=1.985 $X2=1.26 $Y2=2.13
r78 2 32 182 $w=1.7e-07 $l=3.58225e-07 $layer=licon1_NDIFF $count=1 $X=2.27
+ $Y=0.625 $X2=2.41 $Y2=0.92
r79 1 22 182 $w=1.7e-07 $l=3.07124e-07 $layer=licon1_NDIFF $count=1 $X=1.14
+ $Y=0.625 $X2=1.28 $Y2=0.87
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4BB_M%VGND 1 2 3 12 14 18 22 24 25 27 28 29 40 41
+ 44
c45 22 0 2.39111e-20 $X=2.99 $Y=0.77
r46 44 45 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r47 40 41 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r48 38 41 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r49 37 38 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r50 35 44 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.83 $Y=0 $X2=1.745
+ $Y2=0
r51 35 37 52.8449 $w=1.68e-07 $l=8.1e-07 $layer=LI1_cond $X=1.83 $Y=0 $X2=2.64
+ $Y2=0
r52 33 45 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r53 32 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r54 29 38 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=2.64
+ $Y2=0
r55 29 45 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=1.68
+ $Y2=0
r56 27 37 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=2.905 $Y=0 $X2=2.64
+ $Y2=0
r57 27 28 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.905 $Y=0 $X2=2.99
+ $Y2=0
r58 26 40 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=3.075 $Y=0 $X2=3.6
+ $Y2=0
r59 26 28 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.075 $Y=0 $X2=2.99
+ $Y2=0
r60 24 32 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=0.725 $Y=0 $X2=0.72
+ $Y2=0
r61 24 25 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=0.725 $Y=0 $X2=0.83
+ $Y2=0
r62 20 28 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.99 $Y=0.085
+ $X2=2.99 $Y2=0
r63 20 22 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=2.99 $Y=0.085
+ $X2=2.99 $Y2=0.77
r64 16 44 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.745 $Y=0.085
+ $X2=1.745 $Y2=0
r65 16 18 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=1.745 $Y=0.085
+ $X2=1.745 $Y2=0.77
r66 15 25 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=0.935 $Y=0 $X2=0.83
+ $Y2=0
r67 14 44 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.66 $Y=0 $X2=1.745
+ $Y2=0
r68 14 15 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=1.66 $Y=0 $X2=0.935
+ $Y2=0
r69 10 25 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=0.83 $Y=0.085
+ $X2=0.83 $Y2=0
r70 10 12 36.1775 $w=2.08e-07 $l=6.85e-07 $layer=LI1_cond $X=0.83 $Y=0.085
+ $X2=0.83 $Y2=0.77
r71 3 22 182 $w=1.7e-07 $l=3.55176e-07 $layer=licon1_NDIFF $count=1 $X=2.7
+ $Y=0.625 $X2=2.99 $Y2=0.77
r72 2 18 182 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_NDIFF $count=1 $X=1.57
+ $Y=0.625 $X2=1.745 $Y2=0.77
r73 1 12 182 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_NDIFF $count=1 $X=0.67
+ $Y=0.625 $X2=0.83 $Y2=0.77
.ends

