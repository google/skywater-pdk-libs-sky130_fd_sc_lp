* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__mux2i_m A0 A1 S VGND VNB VPB VPWR Y
X0 a_55_125# S VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 a_256_497# A1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X2 a_55_125# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X3 VGND a_55_125# a_250_125# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 a_452_497# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X5 Y A1 a_416_125# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 a_416_125# S VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 VPWR a_55_125# a_256_497# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X8 a_250_125# A0 Y VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 Y A0 a_452_497# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
.ends
