# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__buf_lp
  CLASS CORE ;
  FOREIGN sky130_fd_sc_lp__buf_lp ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.400000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.376000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.465000 0.440000 1.795000 1.485000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.404700 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 0.265000 0.495000 1.835000 ;
        RECT 0.125000 1.835000 0.560000 2.890000 ;
        RECT 0.230000 2.890000 0.560000 3.055000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 2.400000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 2.400000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.400000 0.085000 ;
      RECT 0.000000  3.245000 2.400000 3.415000 ;
      RECT 0.740000  1.165000 1.070000 1.665000 ;
      RECT 0.740000  1.665000 2.225000 1.835000 ;
      RECT 0.760000  2.015000 1.090000 3.245000 ;
      RECT 0.955000  0.085000 1.285000 0.725000 ;
      RECT 1.535000  1.835000 1.865000 3.055000 ;
      RECT 1.975000  0.265000 2.225000 1.665000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
  END
END sky130_fd_sc_lp__buf_lp
END LIBRARY
