* File: sky130_fd_sc_lp__clkinvlp_8.pex.spice
* Created: Fri Aug 28 10:19:06 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__CLKINVLP_8%A 3 7 11 15 19 23 27 31 35 39 43 47 51 55
+ 57 59 63 65 66
r141 78 79 62.8061 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=1.625 $Y=1.407
+ $X2=2.055 $Y2=1.407
r142 73 74 45.2788 $w=3.3e-07 $l=3.1e-07 $layer=POLY_cond $X=0.525 $Y=1.407
+ $X2=0.835 $Y2=1.407
r143 72 73 7.30303 $w=3.3e-07 $l=5e-08 $layer=POLY_cond $X=0.475 $Y=1.407
+ $X2=0.525 $Y2=1.407
r144 70 72 22.6394 $w=3.3e-07 $l=1.55e-07 $layer=POLY_cond $X=0.32 $Y=1.407
+ $X2=0.475 $Y2=1.407
r145 70 71 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.32
+ $Y=1.415 $X2=0.32 $Y2=1.415
r146 66 71 8.1158 $w=3.53e-07 $l=2.5e-07 $layer=LI1_cond $X=0.277 $Y=1.665
+ $X2=0.277 $Y2=1.415
r147 65 71 3.89558 $w=3.53e-07 $l=1.2e-07 $layer=LI1_cond $X=0.277 $Y=1.295
+ $X2=0.277 $Y2=1.415
r148 61 63 227.335 $w=2.5e-07 $l=9.15e-07 $layer=POLY_cond $X=4.235 $Y=1.565
+ $X2=4.235 $Y2=2.48
r149 57 61 77.4121 $w=3.3e-07 $l=5.3e-07 $layer=POLY_cond $X=3.705 $Y=1.407
+ $X2=4.235 $Y2=1.407
r150 57 85 73.0303 $w=3.3e-07 $l=5e-07 $layer=POLY_cond $X=3.705 $Y=1.407
+ $X2=3.205 $Y2=1.407
r151 57 59 227.335 $w=2.5e-07 $l=9.15e-07 $layer=POLY_cond $X=3.705 $Y=1.565
+ $X2=3.705 $Y2=2.48
r152 53 85 21.2229 $w=1.5e-07 $l=1.72e-07 $layer=POLY_cond $X=3.205 $Y=1.235
+ $X2=3.205 $Y2=1.407
r153 53 55 320.479 $w=1.5e-07 $l=6.25e-07 $layer=POLY_cond $X=3.205 $Y=1.235
+ $X2=3.205 $Y2=0.61
r154 49 85 4.38182 $w=3.3e-07 $l=3e-08 $layer=POLY_cond $X=3.175 $Y=1.407
+ $X2=3.205 $Y2=1.407
r155 49 83 48.2 $w=3.3e-07 $l=3.3e-07 $layer=POLY_cond $X=3.175 $Y=1.407
+ $X2=2.845 $Y2=1.407
r156 49 51 227.335 $w=2.5e-07 $l=9.15e-07 $layer=POLY_cond $X=3.175 $Y=1.565
+ $X2=3.175 $Y2=2.48
r157 45 83 21.2229 $w=1.5e-07 $l=1.72e-07 $layer=POLY_cond $X=2.845 $Y=1.235
+ $X2=2.845 $Y2=1.407
r158 45 47 320.479 $w=1.5e-07 $l=6.25e-07 $layer=POLY_cond $X=2.845 $Y=1.235
+ $X2=2.845 $Y2=0.61
r159 41 83 29.2121 $w=3.3e-07 $l=2e-07 $layer=POLY_cond $X=2.645 $Y=1.407
+ $X2=2.845 $Y2=1.407
r160 41 81 33.5939 $w=3.3e-07 $l=2.3e-07 $layer=POLY_cond $X=2.645 $Y=1.407
+ $X2=2.415 $Y2=1.407
r161 41 43 227.335 $w=2.5e-07 $l=9.15e-07 $layer=POLY_cond $X=2.645 $Y=1.565
+ $X2=2.645 $Y2=2.48
r162 37 81 21.2229 $w=1.5e-07 $l=1.72e-07 $layer=POLY_cond $X=2.415 $Y=1.235
+ $X2=2.415 $Y2=1.407
r163 37 39 320.479 $w=1.5e-07 $l=6.25e-07 $layer=POLY_cond $X=2.415 $Y=1.235
+ $X2=2.415 $Y2=0.61
r164 33 81 43.8182 $w=3.3e-07 $l=3e-07 $layer=POLY_cond $X=2.115 $Y=1.407
+ $X2=2.415 $Y2=1.407
r165 33 79 8.76364 $w=3.3e-07 $l=6e-08 $layer=POLY_cond $X=2.115 $Y=1.407
+ $X2=2.055 $Y2=1.407
r166 33 35 227.335 $w=2.5e-07 $l=9.15e-07 $layer=POLY_cond $X=2.115 $Y=1.565
+ $X2=2.115 $Y2=2.48
r167 29 79 21.2229 $w=1.5e-07 $l=1.72e-07 $layer=POLY_cond $X=2.055 $Y=1.235
+ $X2=2.055 $Y2=1.407
r168 29 31 320.479 $w=1.5e-07 $l=6.25e-07 $layer=POLY_cond $X=2.055 $Y=1.235
+ $X2=2.055 $Y2=0.61
r169 25 78 21.2229 $w=1.5e-07 $l=1.72e-07 $layer=POLY_cond $X=1.625 $Y=1.235
+ $X2=1.625 $Y2=1.407
r170 25 27 320.479 $w=1.5e-07 $l=6.25e-07 $layer=POLY_cond $X=1.625 $Y=1.235
+ $X2=1.625 $Y2=0.61
r171 21 78 5.84242 $w=3.3e-07 $l=4e-08 $layer=POLY_cond $X=1.585 $Y=1.407
+ $X2=1.625 $Y2=1.407
r172 21 76 46.7394 $w=3.3e-07 $l=3.2e-07 $layer=POLY_cond $X=1.585 $Y=1.407
+ $X2=1.265 $Y2=1.407
r173 21 23 227.335 $w=2.5e-07 $l=9.15e-07 $layer=POLY_cond $X=1.585 $Y=1.565
+ $X2=1.585 $Y2=2.48
r174 17 76 21.2229 $w=1.5e-07 $l=1.72e-07 $layer=POLY_cond $X=1.265 $Y=1.235
+ $X2=1.265 $Y2=1.407
r175 17 19 320.479 $w=1.5e-07 $l=6.25e-07 $layer=POLY_cond $X=1.265 $Y=1.235
+ $X2=1.265 $Y2=0.61
r176 13 76 30.6727 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=1.055 $Y=1.407
+ $X2=1.265 $Y2=1.407
r177 13 74 32.1333 $w=3.3e-07 $l=2.2e-07 $layer=POLY_cond $X=1.055 $Y=1.407
+ $X2=0.835 $Y2=1.407
r178 13 15 227.335 $w=2.5e-07 $l=9.15e-07 $layer=POLY_cond $X=1.055 $Y=1.565
+ $X2=1.055 $Y2=2.48
r179 9 74 21.2229 $w=1.5e-07 $l=1.72e-07 $layer=POLY_cond $X=0.835 $Y=1.235
+ $X2=0.835 $Y2=1.407
r180 9 11 320.479 $w=1.5e-07 $l=6.25e-07 $layer=POLY_cond $X=0.835 $Y=1.235
+ $X2=0.835 $Y2=0.61
r181 5 73 9.34494 $w=2.5e-07 $l=1.73e-07 $layer=POLY_cond $X=0.525 $Y=1.58
+ $X2=0.525 $Y2=1.407
r182 5 7 223.608 $w=2.5e-07 $l=9e-07 $layer=POLY_cond $X=0.525 $Y=1.58 $X2=0.525
+ $Y2=2.48
r183 1 72 21.2229 $w=1.5e-07 $l=1.72e-07 $layer=POLY_cond $X=0.475 $Y=1.235
+ $X2=0.475 $Y2=1.407
r184 1 3 320.479 $w=1.5e-07 $l=6.25e-07 $layer=POLY_cond $X=0.475 $Y=1.235
+ $X2=0.475 $Y2=0.61
.ends

.subckt PM_SKY130_FD_SC_LP__CLKINVLP_8%VPWR 1 2 3 4 5 16 18 22 26 32 38 42 44 49
+ 50 52 53 54 63 71 75
r72 74 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r73 71 72 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r74 69 72 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.2 $Y2=3.33
r75 68 69 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r76 66 75 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r77 65 66 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r78 63 74 4.69206 $w=1.7e-07 $l=2.32e-07 $layer=LI1_cond $X=4.335 $Y=3.33
+ $X2=4.567 $Y2=3.33
r79 63 65 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=4.335 $Y=3.33
+ $X2=4.08 $Y2=3.33
r80 62 66 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=4.08 $Y2=3.33
r81 61 62 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r82 59 72 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.2 $Y2=3.33
r83 58 59 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r84 56 71 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.485 $Y=3.33
+ $X2=1.32 $Y2=3.33
r85 56 58 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=1.485 $Y=3.33
+ $X2=2.16 $Y2=3.33
r86 54 62 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.4 $Y=3.33
+ $X2=3.12 $Y2=3.33
r87 54 59 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.4 $Y=3.33
+ $X2=2.16 $Y2=3.33
r88 52 61 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=3.275 $Y=3.33
+ $X2=3.12 $Y2=3.33
r89 52 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.275 $Y=3.33
+ $X2=3.44 $Y2=3.33
r90 51 65 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=3.605 $Y=3.33
+ $X2=4.08 $Y2=3.33
r91 51 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.605 $Y=3.33
+ $X2=3.44 $Y2=3.33
r92 49 58 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=2.215 $Y=3.33
+ $X2=2.16 $Y2=3.33
r93 49 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.215 $Y=3.33
+ $X2=2.38 $Y2=3.33
r94 48 61 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=2.545 $Y=3.33
+ $X2=3.12 $Y2=3.33
r95 48 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.545 $Y=3.33
+ $X2=2.38 $Y2=3.33
r96 44 47 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=4.5 $Y=2.125 $X2=4.5
+ $Y2=2.835
r97 42 74 3.07411 $w=3.3e-07 $l=1.13666e-07 $layer=LI1_cond $X=4.5 $Y=3.245
+ $X2=4.567 $Y2=3.33
r98 42 47 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=4.5 $Y=3.245 $X2=4.5
+ $Y2=2.835
r99 38 41 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=3.44 $Y=2.125
+ $X2=3.44 $Y2=2.835
r100 36 53 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.44 $Y=3.245
+ $X2=3.44 $Y2=3.33
r101 36 41 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=3.44 $Y=3.245
+ $X2=3.44 $Y2=2.835
r102 32 35 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=2.38 $Y=2.125
+ $X2=2.38 $Y2=2.835
r103 30 50 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.38 $Y=3.245
+ $X2=2.38 $Y2=3.33
r104 30 35 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=2.38 $Y=3.245
+ $X2=2.38 $Y2=2.835
r105 26 29 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=1.32 $Y=2.125
+ $X2=1.32 $Y2=2.835
r106 24 71 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.32 $Y=3.245
+ $X2=1.32 $Y2=3.33
r107 24 29 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=1.32 $Y=3.245
+ $X2=1.32 $Y2=2.835
r108 23 68 4.78091 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=3.33
+ $X2=0.212 $Y2=3.33
r109 22 71 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.155 $Y=3.33
+ $X2=1.32 $Y2=3.33
r110 22 23 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=1.155 $Y=3.33
+ $X2=0.425 $Y2=3.33
r111 18 21 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=0.26 $Y=2.125
+ $X2=0.26 $Y2=2.835
r112 16 68 2.98526 $w=3.3e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.26 $Y=3.245
+ $X2=0.212 $Y2=3.33
r113 16 21 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=0.26 $Y=3.245
+ $X2=0.26 $Y2=2.835
r114 5 47 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=4.36
+ $Y=1.98 $X2=4.5 $Y2=2.835
r115 5 44 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=4.36
+ $Y=1.98 $X2=4.5 $Y2=2.125
r116 4 41 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=3.3
+ $Y=1.98 $X2=3.44 $Y2=2.835
r117 4 38 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=3.3
+ $Y=1.98 $X2=3.44 $Y2=2.125
r118 3 35 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=2.24
+ $Y=1.98 $X2=2.38 $Y2=2.835
r119 3 32 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.24
+ $Y=1.98 $X2=2.38 $Y2=2.125
r120 2 29 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=1.18
+ $Y=1.98 $X2=1.32 $Y2=2.835
r121 2 26 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.18
+ $Y=1.98 $X2=1.32 $Y2=2.125
r122 1 21 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.98 $X2=0.26 $Y2=2.835
r123 1 18 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.98 $X2=0.26 $Y2=2.125
.ends

.subckt PM_SKY130_FD_SC_LP__CLKINVLP_8%Y 1 2 3 4 5 6 19 23 27 31 35 39 40 43 51
+ 53 56 57 58 59 60 61
r94 60 61 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.79 $Y=2.405
+ $X2=0.79 $Y2=2.775
r95 60 77 9.7783 $w=3.28e-07 $l=2.8e-07 $layer=LI1_cond $X=0.79 $Y=2.405
+ $X2=0.79 $Y2=2.125
r96 59 77 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=0.79 $Y=2.035 $X2=0.79
+ $Y2=2.125
r97 58 59 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.79 $Y=1.665
+ $X2=0.79 $Y2=2.035
r98 58 71 3.49225 $w=3.28e-07 $l=1e-07 $layer=LI1_cond $X=0.79 $Y=1.665 $X2=0.79
+ $Y2=1.565
r99 57 68 5.67595 $w=3.3e-07 $l=1.85e-07 $layer=LI1_cond $X=0.79 $Y=1.38
+ $X2=0.79 $Y2=1.195
r100 57 71 5.67595 $w=3.3e-07 $l=1.85e-07 $layer=LI1_cond $X=0.79 $Y=1.38
+ $X2=0.79 $Y2=1.565
r101 56 68 9.42908 $w=3.28e-07 $l=2.7e-07 $layer=LI1_cond $X=0.79 $Y=0.925
+ $X2=0.79 $Y2=1.195
r102 54 55 8.72119 $w=3.68e-07 $l=2.8e-07 $layer=LI1_cond $X=2.63 $Y=1.38
+ $X2=2.91 $Y2=1.38
r103 48 56 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=0.79 $Y=0.78
+ $X2=0.79 $Y2=0.925
r104 47 51 6.68775 $w=4.63e-07 $l=2.6e-07 $layer=LI1_cond $X=0.79 $Y=0.547
+ $X2=1.05 $Y2=0.547
r105 47 48 2.74626 $w=3.3e-07 $l=2.33e-07 $layer=LI1_cond $X=0.79 $Y=0.547
+ $X2=0.79 $Y2=0.78
r106 43 45 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=3.97 $Y=2.125
+ $X2=3.97 $Y2=2.835
r107 41 43 19.5566 $w=3.28e-07 $l=5.6e-07 $layer=LI1_cond $X=3.97 $Y=1.565
+ $X2=3.97 $Y2=2.125
r108 40 55 5.13927 $w=3.68e-07 $l=1.65e-07 $layer=LI1_cond $X=3.075 $Y=1.38
+ $X2=2.91 $Y2=1.38
r109 39 41 6.84548 $w=3.7e-07 $l=2.5446e-07 $layer=LI1_cond $X=3.805 $Y=1.38
+ $X2=3.97 $Y2=1.565
r110 39 40 22.7374 $w=3.68e-07 $l=7.3e-07 $layer=LI1_cond $X=3.805 $Y=1.38
+ $X2=3.075 $Y2=1.38
r111 35 37 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=2.91 $Y=2.125
+ $X2=2.91 $Y2=2.835
r112 33 55 1.40494 $w=3.3e-07 $l=1.85e-07 $layer=LI1_cond $X=2.91 $Y=1.565
+ $X2=2.91 $Y2=1.38
r113 33 35 19.5566 $w=3.28e-07 $l=5.6e-07 $layer=LI1_cond $X=2.91 $Y=1.565
+ $X2=2.91 $Y2=2.125
r114 29 54 1.40494 $w=3.3e-07 $l=1.85e-07 $layer=LI1_cond $X=2.63 $Y=1.195
+ $X2=2.63 $Y2=1.38
r115 29 31 20.4297 $w=3.28e-07 $l=5.85e-07 $layer=LI1_cond $X=2.63 $Y=1.195
+ $X2=2.63 $Y2=0.61
r116 28 53 4.69202 $w=3.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.015 $Y=1.38
+ $X2=1.85 $Y2=1.38
r117 27 54 5.13927 $w=3.68e-07 $l=1.65e-07 $layer=LI1_cond $X=2.465 $Y=1.38
+ $X2=2.63 $Y2=1.38
r118 27 28 14.0162 $w=3.68e-07 $l=4.5e-07 $layer=LI1_cond $X=2.465 $Y=1.38
+ $X2=2.015 $Y2=1.38
r119 23 25 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=1.85 $Y=2.125
+ $X2=1.85 $Y2=2.835
r120 21 53 1.75761 $w=3.3e-07 $l=1.85e-07 $layer=LI1_cond $X=1.85 $Y=1.565
+ $X2=1.85 $Y2=1.38
r121 21 23 19.5566 $w=3.28e-07 $l=5.6e-07 $layer=LI1_cond $X=1.85 $Y=1.565
+ $X2=1.85 $Y2=2.125
r122 20 57 0.933993 $w=3.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.955 $Y=1.38
+ $X2=0.79 $Y2=1.38
r123 19 53 4.69202 $w=3.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.685 $Y=1.38
+ $X2=1.85 $Y2=1.38
r124 19 20 22.7374 $w=3.68e-07 $l=7.3e-07 $layer=LI1_cond $X=1.685 $Y=1.38
+ $X2=0.955 $Y2=1.38
r125 6 45 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=3.83
+ $Y=1.98 $X2=3.97 $Y2=2.835
r126 6 43 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=3.83
+ $Y=1.98 $X2=3.97 $Y2=2.125
r127 5 37 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=2.77
+ $Y=1.98 $X2=2.91 $Y2=2.835
r128 5 35 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.77
+ $Y=1.98 $X2=2.91 $Y2=2.125
r129 4 25 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=1.71
+ $Y=1.98 $X2=1.85 $Y2=2.835
r130 4 23 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.71
+ $Y=1.98 $X2=1.85 $Y2=2.125
r131 3 61 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=0.65
+ $Y=1.98 $X2=0.79 $Y2=2.835
r132 3 77 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.65
+ $Y=1.98 $X2=0.79 $Y2=2.125
r133 2 31 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=2.49
+ $Y=0.335 $X2=2.63 $Y2=0.61
r134 1 51 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.91
+ $Y=0.335 $X2=1.05 $Y2=0.545
.ends

.subckt PM_SKY130_FD_SC_LP__CLKINVLP_8%VGND 1 2 3 10 12 16 20 23 24 25 27 43 44
+ 50
r49 50 51 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r50 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r51 43 44 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r52 41 44 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.56
+ $Y2=0
r53 40 43 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=3.6 $Y=0 $X2=4.56
+ $Y2=0
r54 40 41 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r55 38 41 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r56 37 38 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r57 35 51 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.68
+ $Y2=0
r58 34 37 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r59 34 35 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r60 32 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.005 $Y=0 $X2=1.84
+ $Y2=0
r61 32 34 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=2.005 $Y=0 $X2=2.16
+ $Y2=0
r62 31 51 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r63 31 48 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r64 30 31 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r65 28 47 4.78091 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=0 $X2=0.212
+ $Y2=0
r66 28 30 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.425 $Y=0 $X2=0.72
+ $Y2=0
r67 27 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.675 $Y=0 $X2=1.84
+ $Y2=0
r68 27 30 62.3048 $w=1.68e-07 $l=9.55e-07 $layer=LI1_cond $X=1.675 $Y=0 $X2=0.72
+ $Y2=0
r69 25 38 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.4 $Y=0 $X2=3.12
+ $Y2=0
r70 25 35 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.4 $Y=0 $X2=2.16
+ $Y2=0
r71 23 37 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=3.255 $Y=0 $X2=3.12
+ $Y2=0
r72 23 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.255 $Y=0 $X2=3.42
+ $Y2=0
r73 22 40 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=3.585 $Y=0 $X2=3.6
+ $Y2=0
r74 22 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.585 $Y=0 $X2=3.42
+ $Y2=0
r75 18 24 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.42 $Y=0.085
+ $X2=3.42 $Y2=0
r76 18 20 18.3343 $w=3.28e-07 $l=5.25e-07 $layer=LI1_cond $X=3.42 $Y=0.085
+ $X2=3.42 $Y2=0.61
r77 14 50 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.84 $Y=0.085
+ $X2=1.84 $Y2=0
r78 14 16 18.3343 $w=3.28e-07 $l=5.25e-07 $layer=LI1_cond $X=1.84 $Y=0.085
+ $X2=1.84 $Y2=0.61
r79 10 47 2.98526 $w=3.3e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.212 $Y2=0
r80 10 12 18.3343 $w=3.28e-07 $l=5.25e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.26 $Y2=0.61
r81 3 20 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=3.28
+ $Y=0.335 $X2=3.42 $Y2=0.61
r82 2 16 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=1.7
+ $Y=0.335 $X2=1.84 $Y2=0.61
r83 1 12 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.335 $X2=0.26 $Y2=0.61
.ends

