* NGSPICE file created from sky130_fd_sc_lp__and2_m.ext - technology: sky130A

.subckt sky130_fd_sc_lp__and2_m A B VGND VNB VPB VPWR X
M1000 X a_34_141# VPWR VPB phighvt w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=2.688e+11p ps=2.96e+06u
M1001 VGND B a_117_141# VNB nshort w=420000u l=150000u
+  ad=1.785e+11p pd=1.69e+06u as=8.82e+10p ps=1.26e+06u
M1002 X a_34_141# VGND VNB nshort w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1003 a_34_141# A VPWR VPB phighvt w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=0p ps=0u
M1004 a_117_141# A a_34_141# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1005 VPWR B a_34_141# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

