* NGSPICE file created from sky130_fd_sc_lp__a221oi_1.ext - technology: sky130A

.subckt sky130_fd_sc_lp__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
M1000 VPWR A1 a_217_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=4.536e+11p pd=3.24e+06u as=1.0836e+12p ps=9.28e+06u
M1001 a_300_47# B2 VGND VNB nshort w=840000u l=150000u
+  ad=1.764e+11p pd=2.1e+06u as=7.56e+11p ps=5.16e+06u
M1002 a_217_367# A2 VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 Y B1 a_300_47# VNB nshort w=840000u l=150000u
+  ad=5.502e+11p pd=4.67e+06u as=0p ps=0u
M1004 a_110_367# B2 a_217_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=7.119e+11p pd=6.17e+06u as=0p ps=0u
M1005 a_480_47# A1 Y VNB nshort w=840000u l=150000u
+  ad=3.276e+11p pd=2.46e+06u as=0p ps=0u
M1006 a_217_367# B1 a_110_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND C1 Y VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND A2 a_480_47# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_110_367# C1 Y VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=3.339e+11p ps=3.05e+06u
.ends

