# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__or4_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_lp__or4_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.840000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.005000 1.355000 2.395000 1.675000 ;
        RECT 2.005000 1.675000 2.245000 2.345000 ;
        RECT 2.005000 2.345000 2.355000 2.960000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.520000 1.005000 1.835000 2.960000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.985000 1.075000 1.350000 2.960000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.760000 0.365000 1.750000 ;
    END
  END D
  PIN X
    ANTENNADIFFAREA  0.594300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.025000 1.105000 3.260000 3.075000 ;
        RECT 3.030000 0.255000 3.260000 1.105000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.840000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.840000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.840000 0.085000 ;
      RECT 0.000000  3.245000 3.840000 3.415000 ;
      RECT 0.300000  0.085000 0.630000 0.565000 ;
      RECT 0.320000  1.920000 0.705000 2.210000 ;
      RECT 0.535000  0.735000 2.285000 0.825000 ;
      RECT 0.535000  0.825000 0.980000 0.905000 ;
      RECT 0.535000  0.905000 0.705000 1.920000 ;
      RECT 0.800000  0.255000 1.090000 0.655000 ;
      RECT 0.800000  0.655000 2.285000 0.735000 ;
      RECT 1.260000  0.085000 1.590000 0.485000 ;
      RECT 1.760000  0.255000 2.020000 0.655000 ;
      RECT 2.005000  0.825000 2.285000 1.015000 ;
      RECT 2.005000  1.015000 2.745000 1.185000 ;
      RECT 2.190000  0.085000 2.860000 0.485000 ;
      RECT 2.415000  1.845000 2.855000 2.175000 ;
      RECT 2.455000  0.485000 2.860000 0.845000 ;
      RECT 2.525000  2.175000 2.855000 3.245000 ;
      RECT 2.575000  1.185000 2.745000 1.285000 ;
      RECT 2.575000  1.285000 2.855000 1.615000 ;
      RECT 3.430000  0.085000 3.720000 1.105000 ;
      RECT 3.430000  1.815000 3.720000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
  END
END sky130_fd_sc_lp__or4_2
END LIBRARY
