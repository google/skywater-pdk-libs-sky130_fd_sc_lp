* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__o221a_m A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
M1000 VGND A1 a_196_179# VNB nshort w=420000u l=150000u
+  ad=2.373e+11p pd=2.81e+06u as=3.225e+11p ps=3.24e+06u
M1001 a_110_179# C1 a_27_179# VNB nshort w=420000u l=150000u
+  ad=2.289e+11p pd=2.77e+06u as=1.113e+11p ps=1.37e+06u
M1002 X a_27_179# VPWR VPB phighvt w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=3.192e+11p ps=3.2e+06u
M1003 a_238_535# B1 VPWR VPB phighvt w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1004 VPWR A1 a_396_535# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.344e+11p ps=1.48e+06u
M1005 a_110_179# B2 a_196_179# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 X a_27_179# VGND VNB nshort w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1007 a_196_179# A2 VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_396_535# A2 a_27_179# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=2.289e+11p ps=2.77e+06u
M1009 a_196_179# B1 a_110_179# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR C1 a_27_179# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_27_179# B2 a_238_535# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
