* File: sky130_fd_sc_lp__a221oi_2.spice
* Created: Fri Aug 28 09:53:25 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__a221oi_2.pex.spice"
.subckt sky130_fd_sc_lp__a221oi_2  VNB VPB C1 B2 B1 A2 A1 Y VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Y	Y
* A1	A1
* A2	A2
* B1	B1
* B2	B2
* C1	C1
* VPB	VPB
* VNB	VNB
MM1003 N_Y_M1003_d N_C1_M1003_g N_VGND_M1003_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75004.6 A=0.126 P=1.98 MULT=1
MM1007 N_Y_M1003_d N_C1_M1007_g N_VGND_M1007_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2856 PD=1.12 PS=1.52 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75004.2 A=0.126 P=1.98 MULT=1
MM1004 N_A_384_47#_M1004_d N_B2_M1004_g N_VGND_M1007_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2856 PD=1.12 PS=1.52 NRD=0 NRS=2.856 M=1 R=5.6 SA=75001.4
+ SB=75003.4 A=0.126 P=1.98 MULT=1
MM1002 N_A_384_47#_M1004_d N_B1_M1002_g N_Y_M1002_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.9
+ SB=75002.9 A=0.126 P=1.98 MULT=1
MM1013 N_A_384_47#_M1013_d N_B1_M1013_g N_Y_M1002_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002.3
+ SB=75002.5 A=0.126 P=1.98 MULT=1
MM1010 N_A_384_47#_M1013_d N_B2_M1010_g N_VGND_M1010_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1848 PD=1.12 PS=1.28 NRD=0 NRS=10.704 M=1 R=5.6 SA=75002.7
+ SB=75002.1 A=0.126 P=1.98 MULT=1
MM1011 N_A_760_47#_M1011_d N_A2_M1011_g N_VGND_M1010_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1848 PD=1.12 PS=1.28 NRD=0 NRS=12.132 M=1 R=5.6 SA=75003.3
+ SB=75001.5 A=0.126 P=1.98 MULT=1
MM1001 N_Y_M1001_d N_A1_M1001_g N_A_760_47#_M1011_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75003.8
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1008 N_Y_M1001_d N_A1_M1008_g N_A_760_47#_M1008_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75004.2
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1015 N_A_760_47#_M1008_s N_A2_M1015_g N_VGND_M1015_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75004.6
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1005 N_A_27_367#_M1005_d N_C1_M1005_g N_Y_M1005_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1018 N_A_27_367#_M1018_d N_C1_M1018_g N_Y_M1005_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75000.2 A=0.189 P=2.82 MULT=1
MM1014 N_A_303_367#_M1014_d N_B2_M1014_g N_A_27_367#_M1014_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75003.3 A=0.189 P=2.82 MULT=1
MM1000 N_A_27_367#_M1014_s N_B1_M1000_g N_A_303_367#_M1000_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75002.9 A=0.189 P=2.82 MULT=1
MM1006 N_A_27_367#_M1006_d N_B1_M1006_g N_A_303_367#_M1000_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75002.5 A=0.189 P=2.82 MULT=1
MM1017 N_A_303_367#_M1017_d N_B2_M1017_g N_A_27_367#_M1006_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.2016 AS=0.1764 PD=1.58 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.5
+ SB=75002.1 A=0.189 P=2.82 MULT=1
MM1012 N_VPWR_M1012_d N_A2_M1012_g N_A_303_367#_M1017_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.2457 AS=0.2016 PD=1.65 PS=1.58 NRD=8.5892 NRS=6.2449 M=1 R=8.4
+ SA=75002 SB=75001.6 A=0.189 P=2.82 MULT=1
MM1009 N_VPWR_M1012_d N_A1_M1009_g N_A_303_367#_M1009_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.2457 AS=0.1764 PD=1.65 PS=1.54 NRD=8.5892 NRS=0 M=1 R=8.4
+ SA=75002.5 SB=75001.1 A=0.189 P=2.82 MULT=1
MM1019 N_VPWR_M1019_d N_A1_M1019_g N_A_303_367#_M1009_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.9
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1016 N_VPWR_M1019_d N_A2_M1016_g N_A_303_367#_M1016_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75003.3
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX20_noxref VNB VPB NWDIODE A=11.4511 P=16.01
*
.include "sky130_fd_sc_lp__a221oi_2.pxi.spice"
*
.ends
*
*
