* File: sky130_fd_sc_lp__dlrtp_lp.pex.spice
* Created: Fri Aug 28 10:27:37 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__DLRTP_LP%GATE 3 7 11 15 17 18 19 30
c31 11 0 1.1902e-19 $X=0.855 $Y=0.495
r32 30 31 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.585
+ $Y=1.345 $X2=0.585 $Y2=1.345
r33 18 19 6.23308 $w=7.08e-07 $l=3.7e-07 $layer=LI1_cond $X=0.48 $Y=1.665
+ $X2=0.48 $Y2=2.035
r34 18 31 5.39078 $w=7.08e-07 $l=3.2e-07 $layer=LI1_cond $X=0.48 $Y=1.665
+ $X2=0.48 $Y2=1.345
r35 17 31 0.842309 $w=7.08e-07 $l=5e-08 $layer=LI1_cond $X=0.48 $Y=1.295
+ $X2=0.48 $Y2=1.345
r36 13 30 97.1997 $w=2.55e-07 $l=5.88154e-07 $layer=POLY_cond $X=0.855 $Y=1.85
+ $X2=0.675 $Y2=1.345
r37 13 15 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=0.855 $Y=1.85
+ $X2=0.855 $Y2=2.67
r38 9 30 32.933 $w=2.55e-07 $l=2.49199e-07 $layer=POLY_cond $X=0.855 $Y=1.18
+ $X2=0.675 $Y2=1.345
r39 9 11 351.245 $w=1.5e-07 $l=6.85e-07 $layer=POLY_cond $X=0.855 $Y=1.18
+ $X2=0.855 $Y2=0.495
r40 5 30 97.1997 $w=2.55e-07 $l=5.88154e-07 $layer=POLY_cond $X=0.495 $Y=1.85
+ $X2=0.675 $Y2=1.345
r41 5 7 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=0.495 $Y=1.85
+ $X2=0.495 $Y2=2.67
r42 1 30 32.933 $w=2.55e-07 $l=1.8e-07 $layer=POLY_cond $X=0.495 $Y=1.345
+ $X2=0.675 $Y2=1.345
r43 1 3 351.245 $w=1.5e-07 $l=8.5e-07 $layer=POLY_cond $X=0.495 $Y=1.345
+ $X2=0.495 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__DLRTP_LP%A_186_57# 1 2 9 11 13 14 16 19 21 25 27 29
+ 31 32 35 39 44 46 47 48 49 51 52 54 57 62 63 67
c131 67 0 8.36941e-20 $X=3.76 $Y=1.06
c132 44 0 1.43074e-19 $X=2.145 $Y=1.59
c133 39 0 1.1902e-19 $X=1.98 $Y=0.35
c134 29 0 1.24286e-19 $X=4.785 $Y=1.035
c135 25 0 1.68694e-19 $X=4.36 $Y=2.035
r136 61 62 104.711 $w=1.68e-07 $l=1.605e-06 $layer=LI1_cond $X=1.15 $Y=0.725
+ $X2=1.15 $Y2=2.33
r137 60 61 10.7321 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=1.07 $Y=0.495
+ $X2=1.07 $Y2=0.725
r138 57 60 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=1.07 $Y=0.35
+ $X2=1.07 $Y2=0.495
r139 55 67 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.595 $Y=1.06
+ $X2=3.76 $Y2=1.06
r140 54 55 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.595
+ $Y=1.06 $X2=3.595 $Y2=1.06
r141 52 54 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=3.32 $Y=1.06
+ $X2=3.595 $Y2=1.06
r142 50 52 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.235 $Y=1.225
+ $X2=3.32 $Y2=1.06
r143 50 51 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=3.235 $Y=1.225
+ $X2=3.235 $Y2=1.59
r144 48 51 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.15 $Y=1.675
+ $X2=3.235 $Y2=1.59
r145 48 49 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=3.15 $Y=1.675
+ $X2=2.31 $Y2=1.675
r146 46 63 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=2.145 $Y=1.06
+ $X2=2.145 $Y2=0.895
r147 46 47 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.145
+ $Y=1.06 $X2=2.145 $Y2=1.06
r148 44 49 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.145 $Y=1.59
+ $X2=2.31 $Y2=1.675
r149 44 46 18.5089 $w=3.28e-07 $l=5.3e-07 $layer=LI1_cond $X=2.145 $Y=1.59
+ $X2=2.145 $Y2=1.06
r150 41 63 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=2.065 $Y=0.435
+ $X2=2.065 $Y2=0.895
r151 40 57 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.235 $Y=0.35
+ $X2=1.07 $Y2=0.35
r152 39 41 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.98 $Y=0.35
+ $X2=2.065 $Y2=0.435
r153 39 40 48.6043 $w=1.68e-07 $l=7.45e-07 $layer=LI1_cond $X=1.98 $Y=0.35
+ $X2=1.235 $Y2=0.35
r154 35 62 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=1.07 $Y=2.495
+ $X2=1.07 $Y2=2.33
r155 29 31 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=4.785 $Y=1.035
+ $X2=4.785 $Y2=0.715
r156 28 32 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.435 $Y=1.11
+ $X2=4.36 $Y2=1.11
r157 27 29 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.71 $Y=1.11
+ $X2=4.785 $Y2=1.035
r158 27 28 141.011 $w=1.5e-07 $l=2.75e-07 $layer=POLY_cond $X=4.71 $Y=1.11
+ $X2=4.435 $Y2=1.11
r159 23 32 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.36 $Y=1.185
+ $X2=4.36 $Y2=1.11
r160 23 25 435.851 $w=1.5e-07 $l=8.5e-07 $layer=POLY_cond $X=4.36 $Y=1.185
+ $X2=4.36 $Y2=2.035
r161 21 32 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.285 $Y=1.11
+ $X2=4.36 $Y2=1.11
r162 21 67 269.202 $w=1.5e-07 $l=5.25e-07 $layer=POLY_cond $X=4.285 $Y=1.11
+ $X2=3.76 $Y2=1.11
r163 17 47 79.2607 $w=3.2e-07 $l=6.19516e-07 $layer=POLY_cond $X=2.355 $Y=1.565
+ $X2=2.1 $Y2=1.06
r164 17 19 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.355 $Y=1.565
+ $X2=2.355 $Y2=2.045
r165 14 47 28.0482 $w=3.2e-07 $l=2.96226e-07 $layer=POLY_cond $X=2.325 $Y=0.895
+ $X2=2.1 $Y2=1.06
r166 14 16 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.325 $Y=0.895
+ $X2=2.325 $Y2=0.575
r167 11 47 28.0482 $w=3.2e-07 $l=2.22486e-07 $layer=POLY_cond $X=1.965 $Y=0.895
+ $X2=2.1 $Y2=1.06
r168 11 13 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.965 $Y=0.895
+ $X2=1.965 $Y2=0.575
r169 7 47 79.2607 $w=3.2e-07 $l=6.19516e-07 $layer=POLY_cond $X=1.845 $Y=1.565
+ $X2=2.1 $Y2=1.06
r170 7 9 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.845 $Y=1.565
+ $X2=1.845 $Y2=2.045
r171 2 35 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=0.93
+ $Y=2.35 $X2=1.07 $Y2=2.495
r172 1 60 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.93
+ $Y=0.285 $X2=1.07 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__DLRTP_LP%D 3 5 7 10 12 14 15 20 22
c42 20 0 8.36941e-20 $X=2.805 $Y=1.245
r43 21 22 15.0178 $w=3.37e-07 $l=1.05e-07 $layer=POLY_cond $X=3.01 $Y=1.347
+ $X2=3.115 $Y2=1.347
r44 19 21 29.3205 $w=3.37e-07 $l=2.05e-07 $layer=POLY_cond $X=2.805 $Y=1.347
+ $X2=3.01 $Y2=1.347
r45 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.805
+ $Y=1.245 $X2=2.805 $Y2=1.245
r46 17 19 7.15134 $w=3.37e-07 $l=5e-08 $layer=POLY_cond $X=2.755 $Y=1.347
+ $X2=2.805 $Y2=1.347
r47 15 20 5.76222 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=2.64 $Y=1.245
+ $X2=2.805 $Y2=1.245
r48 12 22 36.4718 $w=3.37e-07 $l=3.74385e-07 $layer=POLY_cond $X=3.37 $Y=1.615
+ $X2=3.115 $Y2=1.347
r49 12 14 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=3.37 $Y=1.615
+ $X2=3.37 $Y2=2.045
r50 8 22 21.7231 $w=1.5e-07 $l=2.67e-07 $layer=POLY_cond $X=3.115 $Y=1.08
+ $X2=3.115 $Y2=1.347
r51 8 10 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=3.115 $Y=1.08
+ $X2=3.115 $Y2=0.575
r52 5 21 21.7231 $w=1.5e-07 $l=2.68e-07 $layer=POLY_cond $X=3.01 $Y=1.615
+ $X2=3.01 $Y2=1.347
r53 5 7 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=3.01 $Y=1.615 $X2=3.01
+ $Y2=2.045
r54 1 17 21.7231 $w=1.5e-07 $l=2.67e-07 $layer=POLY_cond $X=2.755 $Y=1.08
+ $X2=2.755 $Y2=1.347
r55 1 3 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=2.755 $Y=1.08
+ $X2=2.755 $Y2=0.575
.ends

.subckt PM_SKY130_FD_SC_LP__DLRTP_LP%A_294_547# 1 2 7 12 13 14 17 20 28
c65 28 0 3.17905e-20 $X=1.635 $Y=2.81
c66 13 0 1.4542e-19 $X=5.14 $Y=1.53
c67 12 0 1.1902e-19 $X=4.905 $Y=1.925
r68 26 28 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=1.635 $Y=2.9 $X2=1.635
+ $Y2=2.81
r69 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.635
+ $Y=2.9 $X2=1.635 $Y2=2.9
r70 23 25 35.4333 $w=3.33e-07 $l=1.03e-06 $layer=LI1_cond $X=1.632 $Y=1.87
+ $X2=1.632 $Y2=2.9
r71 20 23 37.4974 $w=3.33e-07 $l=1.09e-06 $layer=LI1_cond $X=1.632 $Y=0.78
+ $X2=1.632 $Y2=1.87
r72 15 17 379.447 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=5.215 $Y=1.455
+ $X2=5.215 $Y2=0.715
r73 13 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.14 $Y=1.53
+ $X2=5.215 $Y2=1.455
r74 13 14 82.0426 $w=1.5e-07 $l=1.6e-07 $layer=POLY_cond $X=5.14 $Y=1.53
+ $X2=4.98 $Y2=1.53
r75 10 12 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=4.905 $Y=2.735
+ $X2=4.905 $Y2=1.925
r76 9 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.905 $Y=1.605
+ $X2=4.98 $Y2=1.53
r77 9 12 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=4.905 $Y=1.605
+ $X2=4.905 $Y2=1.925
r78 8 28 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.8 $Y=2.81
+ $X2=1.635 $Y2=2.81
r79 7 10 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.83 $Y=2.81
+ $X2=4.905 $Y2=2.735
r80 7 8 1553.68 $w=1.5e-07 $l=3.03e-06 $layer=POLY_cond $X=4.83 $Y=2.81 $X2=1.8
+ $Y2=2.81
r81 2 23 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=1.485
+ $Y=1.725 $X2=1.63 $Y2=1.87
r82 1 20 182 $w=1.7e-07 $l=4.82079e-07 $layer=licon1_NDIFF $count=1 $X=1.49
+ $Y=0.365 $X2=1.635 $Y2=0.78
.ends

.subckt PM_SKY130_FD_SC_LP__DLRTP_LP%A_638_73# 1 2 9 14 17 19 20 25 26 27 28 30
+ 34 36
c88 30 0 1.68694e-19 $X=5.6 $Y=2.9
r89 36 38 3.49225 $w=3.28e-07 $l=1e-07 $layer=LI1_cond $X=3.33 $Y=0.53 $X2=3.33
+ $Y2=0.63
r90 33 34 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=4.025 $Y=0.715
+ $X2=4.025 $Y2=1.405
r91 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.6 $Y=2.9
+ $X2=5.6 $Y2=2.9
r92 28 30 64.6067 $w=3.28e-07 $l=1.85e-06 $layer=LI1_cond $X=3.75 $Y=2.9 $X2=5.6
+ $Y2=2.9
r93 26 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.94 $Y=1.49
+ $X2=4.025 $Y2=1.405
r94 26 27 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=3.94 $Y=1.49
+ $X2=3.75 $Y2=1.49
r95 23 28 6.98653 $w=3.3e-07 $l=2.18746e-07 $layer=LI1_cond $X=3.625 $Y=2.735
+ $X2=3.75 $Y2=2.9
r96 23 25 39.8745 $w=2.48e-07 $l=8.65e-07 $layer=LI1_cond $X=3.625 $Y=2.735
+ $X2=3.625 $Y2=1.87
r97 22 27 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.625 $Y=1.575
+ $X2=3.75 $Y2=1.49
r98 22 25 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=3.625 $Y=1.575
+ $X2=3.625 $Y2=1.87
r99 21 38 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.495 $Y=0.63
+ $X2=3.33 $Y2=0.63
r100 20 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.94 $Y=0.63
+ $X2=4.025 $Y2=0.715
r101 20 21 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=3.94 $Y=0.63
+ $X2=3.495 $Y2=0.63
r102 19 31 38.4695 $w=3.3e-07 $l=2.2e-07 $layer=POLY_cond $X=5.82 $Y=2.9 $X2=5.6
+ $Y2=2.9
r103 15 17 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=5.605 $Y=1.5
+ $X2=5.895 $Y2=1.5
r104 12 19 32.1775 $w=3.3e-07 $l=1.98997e-07 $layer=POLY_cond $X=5.895 $Y=2.735
+ $X2=5.82 $Y2=2.9
r105 12 14 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=5.895 $Y=2.735
+ $X2=5.895 $Y2=2.255
r106 11 17 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.895 $Y=1.575
+ $X2=5.895 $Y2=1.5
r107 11 14 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=5.895 $Y=1.575
+ $X2=5.895 $Y2=2.255
r108 7 15 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.605 $Y=1.425
+ $X2=5.605 $Y2=1.5
r109 7 9 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=5.605 $Y=1.425
+ $X2=5.605 $Y2=0.715
r110 2 25 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=3.445
+ $Y=1.725 $X2=3.585 $Y2=1.87
r111 1 36 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=3.19
+ $Y=0.365 $X2=3.33 $Y2=0.53
.ends

.subckt PM_SKY130_FD_SC_LP__DLRTP_LP%A_1208_75# 1 2 7 9 10 11 14 16 18 20 21 23
+ 24 26 27 28 31 33 34 36 37 38 43 46 49 55 57
c123 38 0 1.19126e-20 $X=9.075 $Y=1.9
r124 56 63 36.9716 $w=3.52e-07 $l=2.7e-07 $layer=POLY_cond $X=9.3 $Y=1.455
+ $X2=9.57 $Y2=1.455
r125 56 61 12.3239 $w=3.52e-07 $l=9e-08 $layer=POLY_cond $X=9.3 $Y=1.455
+ $X2=9.21 $Y2=1.455
r126 55 58 8.60763 $w=3.88e-07 $l=1.65e-07 $layer=LI1_cond $X=9.27 $Y=1.35
+ $X2=9.27 $Y2=1.515
r127 55 57 8.60763 $w=3.88e-07 $l=1.65e-07 $layer=LI1_cond $X=9.27 $Y=1.35
+ $X2=9.27 $Y2=1.185
r128 55 56 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.3
+ $Y=1.35 $X2=9.3 $Y2=1.35
r129 49 52 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=8.465 $Y=1.9 $X2=8.465
+ $Y2=1.98
r130 45 48 8.51163 $w=6.02e-07 $l=4.2e-07 $layer=LI1_cond $X=6.84 $Y=0.6
+ $X2=7.26 $Y2=0.6
r131 45 46 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.84
+ $Y=0.43 $X2=6.84 $Y2=0.43
r132 43 58 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=9.16 $Y=1.815
+ $X2=9.16 $Y2=1.515
r133 40 57 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=9.16 $Y=0.815
+ $X2=9.16 $Y2=1.185
r134 39 49 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.63 $Y=1.9
+ $X2=8.465 $Y2=1.9
r135 38 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.075 $Y=1.9
+ $X2=9.16 $Y2=1.815
r136 38 39 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=9.075 $Y=1.9
+ $X2=8.63 $Y2=1.9
r137 37 48 10.3725 $w=6.02e-07 $l=2.20624e-07 $layer=LI1_cond $X=7.425 $Y=0.73
+ $X2=7.26 $Y2=0.6
r138 36 40 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.075 $Y=0.73
+ $X2=9.16 $Y2=0.815
r139 36 37 107.647 $w=1.68e-07 $l=1.65e-06 $layer=LI1_cond $X=9.075 $Y=0.73
+ $X2=7.425 $Y2=0.73
r140 34 46 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=6.84 $Y=0.77
+ $X2=6.84 $Y2=0.43
r141 34 35 54.9356 $w=3.3e-07 $l=3.47419e-07 $layer=POLY_cond $X=6.84 $Y=0.77
+ $X2=6.825 $Y2=1.11
r142 29 31 579.426 $w=1.5e-07 $l=1.13e-06 $layer=POLY_cond $X=10.06 $Y=1.335
+ $X2=10.06 $Y2=2.465
r143 27 29 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.985 $Y=1.26
+ $X2=10.06 $Y2=1.335
r144 27 28 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=9.985 $Y=1.26
+ $X2=9.645 $Y2=1.26
r145 24 28 19.6371 $w=3.52e-07 $l=4.77336e-07 $layer=POLY_cond $X=9.67 $Y=1.725
+ $X2=9.645 $Y2=1.26
r146 24 63 13.6932 $w=3.52e-07 $l=3.1607e-07 $layer=POLY_cond $X=9.67 $Y=1.725
+ $X2=9.57 $Y2=1.455
r147 24 26 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=9.67 $Y=1.725
+ $X2=9.67 $Y2=2.465
r148 21 63 22.7654 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=9.57 $Y=1.185
+ $X2=9.57 $Y2=1.455
r149 21 23 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=9.57 $Y=1.185
+ $X2=9.57 $Y2=0.655
r150 18 61 22.7654 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=9.21 $Y=1.185
+ $X2=9.21 $Y2=1.455
r151 18 20 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=9.21 $Y=1.185
+ $X2=9.21 $Y2=0.655
r152 17 33 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.515 $Y=1.11
+ $X2=6.44 $Y2=1.11
r153 16 35 11.8763 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=6.675 $Y=1.11
+ $X2=6.825 $Y2=1.11
r154 16 17 82.0426 $w=1.5e-07 $l=1.6e-07 $layer=POLY_cond $X=6.675 $Y=1.11
+ $X2=6.515 $Y2=1.11
r155 12 33 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.44 $Y=1.185
+ $X2=6.44 $Y2=1.11
r156 12 14 492.255 $w=1.5e-07 $l=9.6e-07 $layer=POLY_cond $X=6.44 $Y=1.185
+ $X2=6.44 $Y2=2.145
r157 10 33 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.365 $Y=1.11
+ $X2=6.44 $Y2=1.11
r158 10 11 89.734 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=6.365 $Y=1.11
+ $X2=6.19 $Y2=1.11
r159 7 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.115 $Y=1.035
+ $X2=6.19 $Y2=1.11
r160 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=6.115 $Y=1.035
+ $X2=6.115 $Y2=0.715
r161 2 52 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=8.325
+ $Y=1.835 $X2=8.465 $Y2=1.98
r162 1 48 182 $w=1.7e-07 $l=3.70473e-07 $layer=licon1_NDIFF $count=1 $X=7.115
+ $Y=0.235 $X2=7.26 $Y2=0.54
.ends

.subckt PM_SKY130_FD_SC_LP__DLRTP_LP%A_887_343# 1 2 9 13 16 20 24 26 27 29 30 31
+ 34 35 42 44
r119 42 45 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.385 $Y=1.35
+ $X2=7.385 $Y2=1.515
r120 42 44 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.385 $Y=1.35
+ $X2=7.385 $Y2=1.185
r121 41 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.385
+ $Y=1.35 $X2=7.385 $Y2=1.35
r122 35 48 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.73 $Y=1.46
+ $X2=8.73 $Y2=1.625
r123 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.73
+ $Y=1.46 $X2=8.73 $Y2=1.46
r124 32 34 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=8.73 $Y=1.165
+ $X2=8.73 $Y2=1.46
r125 30 32 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=8.565 $Y=1.08
+ $X2=8.73 $Y2=1.165
r126 30 31 66.2193 $w=1.68e-07 $l=1.015e-06 $layer=LI1_cond $X=8.565 $Y=1.08
+ $X2=7.55 $Y2=1.08
r127 29 41 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.385 $Y=1.345
+ $X2=7.385 $Y2=1.43
r128 28 31 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=7.385 $Y=1.165
+ $X2=7.55 $Y2=1.08
r129 28 29 6.28605 $w=3.28e-07 $l=1.8e-07 $layer=LI1_cond $X=7.385 $Y=1.165
+ $X2=7.385 $Y2=1.345
r130 26 41 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.22 $Y=1.43
+ $X2=7.385 $Y2=1.43
r131 26 27 139.289 $w=1.68e-07 $l=2.135e-06 $layer=LI1_cond $X=7.22 $Y=1.43
+ $X2=5.085 $Y2=1.43
r132 22 27 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=4.96 $Y=1.43
+ $X2=5.085 $Y2=1.43
r133 22 24 26.0452 $w=2.48e-07 $l=5.65e-07 $layer=LI1_cond $X=4.96 $Y=1.345
+ $X2=4.96 $Y2=0.78
r134 18 22 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=4.615 $Y=1.43
+ $X2=4.96 $Y2=1.43
r135 18 20 20.0525 $w=2.48e-07 $l=4.35e-07 $layer=LI1_cond $X=4.615 $Y=1.515
+ $X2=4.615 $Y2=1.95
r136 16 48 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=8.68 $Y=2.465
+ $X2=8.68 $Y2=1.625
r137 13 44 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=7.475 $Y=0.655
+ $X2=7.475 $Y2=1.185
r138 9 45 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=7.46 $Y=2.465
+ $X2=7.46 $Y2=1.515
r139 2 20 600 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_PDIFF $count=1 $X=4.435
+ $Y=1.715 $X2=4.575 $Y2=1.95
r140 1 24 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=4.86
+ $Y=0.505 $X2=5 $Y2=0.78
.ends

.subckt PM_SKY130_FD_SC_LP__DLRTP_LP%RESET_B 3 7 11 13 18 19
c45 18 0 1.33771e-19 $X=7.955 $Y=1.51
c46 11 0 1.19126e-20 $X=8.25 $Y=2.465
r47 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.955
+ $Y=1.51 $X2=7.955 $Y2=1.51
r48 16 18 12.0038 $w=2.61e-07 $l=6.5e-08 $layer=POLY_cond $X=7.89 $Y=1.51
+ $X2=7.955 $Y2=1.51
r49 15 16 4.61686 $w=2.61e-07 $l=2.5e-08 $layer=POLY_cond $X=7.865 $Y=1.51
+ $X2=7.89 $Y2=1.51
r50 13 19 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=7.955 $Y=1.665
+ $X2=7.955 $Y2=1.51
r51 9 18 54.4789 $w=2.61e-07 $l=3.68375e-07 $layer=POLY_cond $X=8.25 $Y=1.675
+ $X2=7.955 $Y2=1.51
r52 9 11 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=8.25 $Y=1.675
+ $X2=8.25 $Y2=2.465
r53 5 16 15.717 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.89 $Y=1.675
+ $X2=7.89 $Y2=1.51
r54 5 7 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=7.89 $Y=1.675 $X2=7.89
+ $Y2=2.465
r55 1 15 15.717 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.865 $Y=1.345
+ $X2=7.865 $Y2=1.51
r56 1 3 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=7.865 $Y=1.345
+ $X2=7.865 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__DLRTP_LP%VPWR 1 2 3 4 5 16 18 22 26 30 34 37 38 39
+ 41 49 61 67 68 74 77 80
c92 68 0 3.17905e-20 $X=10.32 $Y=3.33
r93 80 81 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r94 77 78 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r95 74 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r96 71 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r97 68 81 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=10.32 $Y=3.33
+ $X2=9.36 $Y2=3.33
r98 67 68 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.32 $Y=3.33
+ $X2=10.32 $Y2=3.33
r99 65 80 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.62 $Y=3.33
+ $X2=9.455 $Y2=3.33
r100 65 67 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=9.62 $Y=3.33
+ $X2=10.32 $Y2=3.33
r101 64 81 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=9.36 $Y2=3.33
r102 63 64 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r103 61 80 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.29 $Y=3.33
+ $X2=9.455 $Y2=3.33
r104 61 63 89.3797 $w=1.68e-07 $l=1.37e-06 $layer=LI1_cond $X=9.29 $Y=3.33
+ $X2=7.92 $Y2=3.33
r105 60 64 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=7.92 $Y2=3.33
r106 59 60 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r107 57 60 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=7.44 $Y2=3.33
r108 57 78 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33 $X2=6
+ $Y2=3.33
r109 56 59 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=6.48 $Y=3.33
+ $X2=7.44 $Y2=3.33
r110 56 57 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r111 54 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.275 $Y=3.33
+ $X2=6.11 $Y2=3.33
r112 54 56 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=6.275 $Y=3.33
+ $X2=6.48 $Y2=3.33
r113 53 75 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.64 $Y2=3.33
r114 52 53 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r115 50 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.735 $Y=3.33
+ $X2=2.57 $Y2=3.33
r116 50 52 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=2.735 $Y=3.33
+ $X2=3.12 $Y2=3.33
r117 49 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.945 $Y=3.33
+ $X2=6.11 $Y2=3.33
r118 49 52 184.305 $w=1.68e-07 $l=2.825e-06 $layer=LI1_cond $X=5.945 $Y=3.33
+ $X2=3.12 $Y2=3.33
r119 48 75 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r120 47 48 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r121 45 48 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=2.16 $Y2=3.33
r122 45 72 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r123 44 47 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=0.72 $Y=3.33
+ $X2=2.16 $Y2=3.33
r124 44 45 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r125 42 71 4.73185 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=3.33
+ $X2=0.222 $Y2=3.33
r126 42 44 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.445 $Y=3.33
+ $X2=0.72 $Y2=3.33
r127 41 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.405 $Y=3.33
+ $X2=2.57 $Y2=3.33
r128 41 47 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=2.405 $Y=3.33
+ $X2=2.16 $Y2=3.33
r129 39 78 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=5.28 $Y=3.33 $X2=6
+ $Y2=3.33
r130 39 53 0.602067 $w=4.9e-07 $l=2.16e-06 $layer=MET1_cond $X=5.28 $Y=3.33
+ $X2=3.12 $Y2=3.33
r131 37 59 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=7.59 $Y=3.33
+ $X2=7.44 $Y2=3.33
r132 37 38 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.59 $Y=3.33
+ $X2=7.715 $Y2=3.33
r133 36 63 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=7.84 $Y=3.33 $X2=7.92
+ $Y2=3.33
r134 36 38 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.84 $Y=3.33
+ $X2=7.715 $Y2=3.33
r135 32 80 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.455 $Y=3.245
+ $X2=9.455 $Y2=3.33
r136 32 34 31.9541 $w=3.28e-07 $l=9.15e-07 $layer=LI1_cond $X=9.455 $Y=3.245
+ $X2=9.455 $Y2=2.33
r137 28 38 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.715 $Y=3.245
+ $X2=7.715 $Y2=3.33
r138 28 30 16.1342 $w=2.48e-07 $l=3.5e-07 $layer=LI1_cond $X=7.715 $Y=3.245
+ $X2=7.715 $Y2=2.895
r139 24 77 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.11 $Y=3.245
+ $X2=6.11 $Y2=3.33
r140 24 26 32.3033 $w=3.28e-07 $l=9.25e-07 $layer=LI1_cond $X=6.11 $Y=3.245
+ $X2=6.11 $Y2=2.32
r141 20 74 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.57 $Y=3.245
+ $X2=2.57 $Y2=3.33
r142 20 22 37.8909 $w=3.28e-07 $l=1.085e-06 $layer=LI1_cond $X=2.57 $Y=3.245
+ $X2=2.57 $Y2=2.16
r143 16 71 3.03433 $w=3.3e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.222 $Y2=3.33
r144 16 18 26.1919 $w=3.28e-07 $l=7.5e-07 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.28 $Y2=2.495
r145 5 34 300 $w=1.7e-07 $l=5.6285e-07 $layer=licon1_PDIFF $count=2 $X=9.31
+ $Y=1.835 $X2=9.455 $Y2=2.33
r146 4 30 600 $w=1.7e-07 $l=1.12783e-06 $layer=licon1_PDIFF $count=1 $X=7.535
+ $Y=1.835 $X2=7.675 $Y2=2.895
r147 3 26 600 $w=1.7e-07 $l=4.49583e-07 $layer=licon1_PDIFF $count=1 $X=5.97
+ $Y=1.935 $X2=6.11 $Y2=2.32
r148 2 22 600 $w=1.7e-07 $l=5.00125e-07 $layer=licon1_PDIFF $count=1 $X=2.43
+ $Y=1.725 $X2=2.57 $Y2=2.16
r149 1 18 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.35 $X2=0.28 $Y2=2.495
.ends

.subckt PM_SKY130_FD_SC_LP__DLRTP_LP%A_800_343# 1 2 9 11 12 15
r24 13 15 3.91831 $w=2.48e-07 $l=8.5e-08 $layer=LI1_cond $X=5.64 $Y=2.385
+ $X2=5.64 $Y2=2.3
r25 11 13 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=5.515 $Y=2.47
+ $X2=5.64 $Y2=2.385
r26 11 12 78.615 $w=1.68e-07 $l=1.205e-06 $layer=LI1_cond $X=5.515 $Y=2.47
+ $X2=4.31 $Y2=2.47
r27 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.145 $Y=2.385
+ $X2=4.31 $Y2=2.47
r28 7 9 11.1752 $w=3.28e-07 $l=3.2e-07 $layer=LI1_cond $X=4.145 $Y=2.385
+ $X2=4.145 $Y2=2.065
r29 2 15 600 $w=1.7e-07 $l=4.31451e-07 $layer=licon1_PDIFF $count=1 $X=5.535
+ $Y=1.935 $X2=5.68 $Y2=2.3
r30 1 9 600 $w=1.7e-07 $l=4.16233e-07 $layer=licon1_PDIFF $count=1 $X=4 $Y=1.715
+ $X2=4.145 $Y2=2.065
.ends

.subckt PM_SKY130_FD_SC_LP__DLRTP_LP%A_996_343# 1 2 7 11 13
c25 7 0 2.6444e-19 $X=6.49 $Y=1.78
r26 13 16 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=5.12 $Y=1.78
+ $X2=5.12 $Y2=1.925
r27 9 11 9.7783 $w=3.28e-07 $l=2.8e-07 $layer=LI1_cond $X=6.655 $Y=1.865
+ $X2=6.655 $Y2=2.145
r28 8 13 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.285 $Y=1.78
+ $X2=5.12 $Y2=1.78
r29 7 9 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.49 $Y=1.78
+ $X2=6.655 $Y2=1.865
r30 7 8 78.615 $w=1.68e-07 $l=1.205e-06 $layer=LI1_cond $X=6.49 $Y=1.78
+ $X2=5.285 $Y2=1.78
r31 2 11 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=6.515
+ $Y=1.935 $X2=6.655 $Y2=2.145
r32 1 16 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=4.98
+ $Y=1.715 $X2=5.12 $Y2=1.925
.ends

.subckt PM_SKY130_FD_SC_LP__DLRTP_LP%A_1420_367# 1 2 9 13 15 17 19 21
c41 15 0 1.33771e-19 $X=8.81 $Y=2.41
r42 17 23 3.18546 $w=2.5e-07 $l=1.65e-07 $layer=LI1_cond $X=8.935 $Y=2.495
+ $X2=8.935 $Y2=2.33
r43 17 19 18.6696 $w=2.48e-07 $l=4.05e-07 $layer=LI1_cond $X=8.935 $Y=2.495
+ $X2=8.935 $Y2=2.9
r44 16 21 3.80956 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.41 $Y=2.41
+ $X2=7.245 $Y2=2.41
r45 15 23 3.9577 $w=1.7e-07 $l=1.60078e-07 $layer=LI1_cond $X=8.81 $Y=2.41
+ $X2=8.935 $Y2=2.33
r46 15 16 91.3369 $w=1.68e-07 $l=1.4e-06 $layer=LI1_cond $X=8.81 $Y=2.41
+ $X2=7.41 $Y2=2.41
r47 11 21 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.245 $Y=2.495
+ $X2=7.245 $Y2=2.41
r48 11 13 14.1436 $w=3.28e-07 $l=4.05e-07 $layer=LI1_cond $X=7.245 $Y=2.495
+ $X2=7.245 $Y2=2.9
r49 7 21 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.245 $Y=2.325
+ $X2=7.245 $Y2=2.41
r50 7 9 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=7.245 $Y=2.325
+ $X2=7.245 $Y2=1.98
r51 2 23 600 $w=1.7e-07 $l=5.60647e-07 $layer=licon1_PDIFF $count=1 $X=8.755
+ $Y=1.835 $X2=8.895 $Y2=2.33
r52 2 19 600 $w=1.7e-07 $l=1.13284e-06 $layer=licon1_PDIFF $count=1 $X=8.755
+ $Y=1.835 $X2=8.895 $Y2=2.9
r53 1 13 400 $w=1.7e-07 $l=1.13519e-06 $layer=licon1_PDIFF $count=1 $X=7.1
+ $Y=1.835 $X2=7.245 $Y2=2.9
r54 1 9 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=7.1
+ $Y=1.835 $X2=7.245 $Y2=1.98
.ends

.subckt PM_SKY130_FD_SC_LP__DLRTP_LP%Q 1 2 7 8 9 10 11 12 13 37
r19 13 34 4.36531 $w=3.28e-07 $l=1.25e-07 $layer=LI1_cond $X=10.275 $Y=2.775
+ $X2=10.275 $Y2=2.9
r20 12 13 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=10.275 $Y=2.405
+ $X2=10.275 $Y2=2.775
r21 11 12 14.8421 $w=3.28e-07 $l=4.25e-07 $layer=LI1_cond $X=10.275 $Y=1.98
+ $X2=10.275 $Y2=2.405
r22 10 11 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=10.275 $Y=1.665
+ $X2=10.275 $Y2=1.98
r23 9 10 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=10.275 $Y=1.295
+ $X2=10.275 $Y2=1.665
r24 9 43 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=10.275 $Y=1.295
+ $X2=10.275 $Y2=1.095
r25 8 43 6.75651 $w=7.93e-07 $l=1.7e-07 $layer=LI1_cond $X=10.042 $Y=0.925
+ $X2=10.042 $Y2=1.095
r26 7 8 5.56665 $w=7.93e-07 $l=3.7e-07 $layer=LI1_cond $X=10.042 $Y=0.555
+ $X2=10.042 $Y2=0.925
r27 7 37 1.88063 $w=7.93e-07 $l=1.25e-07 $layer=LI1_cond $X=10.042 $Y=0.555
+ $X2=10.042 $Y2=0.43
r28 2 34 400 $w=1.7e-07 $l=1.13284e-06 $layer=licon1_PDIFF $count=1 $X=10.135
+ $Y=1.835 $X2=10.275 $Y2=2.9
r29 2 11 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=10.135
+ $Y=1.835 $X2=10.275 $Y2=1.98
r30 1 37 91 $w=1.7e-07 $l=2.64953e-07 $layer=licon1_NDIFF $count=2 $X=9.645
+ $Y=0.235 $X2=9.81 $Y2=0.43
.ends

.subckt PM_SKY130_FD_SC_LP__DLRTP_LP%VGND 1 2 3 4 13 15 19 23 27 30 31 32 34 46
+ 55 56 62 65
r92 65 66 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r93 62 63 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=2.64 $Y=0
+ $X2=2.64 $Y2=0
r94 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r95 55 56 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=10.32 $Y=0
+ $X2=10.32 $Y2=0
r96 53 56 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=8.4 $Y=0 $X2=10.32
+ $Y2=0
r97 53 66 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=0 $X2=7.92
+ $Y2=0
r98 52 55 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=8.4 $Y=0 $X2=10.32
+ $Y2=0
r99 52 53 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r100 50 65 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.245 $Y=0 $X2=8.08
+ $Y2=0
r101 50 52 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=8.245 $Y=0 $X2=8.4
+ $Y2=0
r102 49 66 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=6 $Y=0 $X2=7.92
+ $Y2=0
r103 48 49 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6 $Y=0 $X2=6
+ $Y2=0
r104 46 65 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.915 $Y=0 $X2=8.08
+ $Y2=0
r105 46 48 124.936 $w=1.68e-07 $l=1.915e-06 $layer=LI1_cond $X=7.915 $Y=0 $X2=6
+ $Y2=0
r106 45 49 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=6
+ $Y2=0
r107 44 45 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=5.52 $Y=0
+ $X2=5.52 $Y2=0
r108 42 62 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.705 $Y=0 $X2=2.54
+ $Y2=0
r109 42 44 183.652 $w=1.68e-07 $l=2.815e-06 $layer=LI1_cond $X=2.705 $Y=0
+ $X2=5.52 $Y2=0
r110 41 63 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r111 40 41 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r112 38 41 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=0.72 $Y=0
+ $X2=2.16 $Y2=0
r113 38 60 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r114 37 40 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=0.72 $Y=0 $X2=2.16
+ $Y2=0
r115 37 38 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r116 35 59 4.73185 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=0
+ $X2=0.222 $Y2=0
r117 35 37 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.445 $Y=0
+ $X2=0.72 $Y2=0
r118 34 62 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.375 $Y=0 $X2=2.54
+ $Y2=0
r119 34 40 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=2.375 $Y=0
+ $X2=2.16 $Y2=0
r120 32 45 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=5.28 $Y=0
+ $X2=5.52 $Y2=0
r121 32 63 0.73586 $w=4.9e-07 $l=2.64e-06 $layer=MET1_cond $X=5.28 $Y=0 $X2=2.64
+ $Y2=0
r122 30 44 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=5.655 $Y=0
+ $X2=5.52 $Y2=0
r123 30 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.655 $Y=0 $X2=5.82
+ $Y2=0
r124 29 48 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=5.985 $Y=0 $X2=6
+ $Y2=0
r125 29 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.985 $Y=0 $X2=5.82
+ $Y2=0
r126 25 65 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.08 $Y=0.085
+ $X2=8.08 $Y2=0
r127 25 27 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=8.08 $Y=0.085
+ $X2=8.08 $Y2=0.38
r128 21 31 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.82 $Y=0.085
+ $X2=5.82 $Y2=0
r129 21 23 19.7312 $w=3.28e-07 $l=5.65e-07 $layer=LI1_cond $X=5.82 $Y=0.085
+ $X2=5.82 $Y2=0.65
r130 17 62 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.54 $Y=0.085
+ $X2=2.54 $Y2=0
r131 17 19 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=2.54 $Y=0.085
+ $X2=2.54 $Y2=0.53
r132 13 59 3.03433 $w=3.3e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.28 $Y=0.085
+ $X2=0.222 $Y2=0
r133 13 15 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=0.28 $Y=0.085
+ $X2=0.28 $Y2=0.495
r134 4 27 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=7.94
+ $Y=0.235 $X2=8.08 $Y2=0.38
r135 3 23 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=5.68
+ $Y=0.505 $X2=5.82 $Y2=0.65
r136 2 19 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=2.4
+ $Y=0.365 $X2=2.54 $Y2=0.53
r137 1 15 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.285 $X2=0.28 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__DLRTP_LP%A_862_101# 1 2 9 11 12 14 15 16 19
c49 16 0 1.24286e-19 $X=5.435 $Y=1.08
r50 17 19 9.7783 $w=3.28e-07 $l=2.8e-07 $layer=LI1_cond $X=6.33 $Y=0.995
+ $X2=6.33 $Y2=0.715
r51 15 17 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.165 $Y=1.08
+ $X2=6.33 $Y2=0.995
r52 15 16 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=6.165 $Y=1.08
+ $X2=5.435 $Y2=1.08
r53 14 16 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.35 $Y=0.995
+ $X2=5.435 $Y2=1.08
r54 13 14 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=5.35 $Y=0.435
+ $X2=5.35 $Y2=0.995
r55 11 13 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.265 $Y=0.35
+ $X2=5.35 $Y2=0.435
r56 11 12 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=5.265 $Y=0.35
+ $X2=4.62 $Y2=0.35
r57 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.455 $Y=0.435
+ $X2=4.62 $Y2=0.35
r58 7 9 9.7783 $w=3.28e-07 $l=2.8e-07 $layer=LI1_cond $X=4.455 $Y=0.435
+ $X2=4.455 $Y2=0.715
r59 2 19 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=6.19
+ $Y=0.505 $X2=6.33 $Y2=0.715
r60 1 9 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=4.31
+ $Y=0.505 $X2=4.455 $Y2=0.715
.ends

