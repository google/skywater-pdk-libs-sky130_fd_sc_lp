* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__ebufn_lp A TE_B VGND VNB VPB VPWR Z
X0 VPWR TE_B a_702_401# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X1 a_308_47# a_29_483# Z VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X2 Z a_29_483# a_515_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X3 VGND TE_B a_708_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 a_116_483# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X5 VGND a_242_237# a_308_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X6 a_702_401# TE_B a_242_237# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X7 a_708_47# TE_B a_242_237# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 a_122_131# A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 a_29_483# A a_122_131# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 a_29_483# A a_116_483# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X11 a_515_367# TE_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
.ends
