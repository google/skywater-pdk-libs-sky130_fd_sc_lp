* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__o2bb2a_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
M1000 a_300_21# A2_N VPWR VPB phighvt w=640000u l=150000u
+  ad=1.792e+11p pd=1.84e+06u as=1.6214e+12p ps=1.164e+07u
M1001 a_150_367# B1 VPWR VPB phighvt w=640000u l=150000u
+  ad=1.344e+11p pd=1.7e+06u as=0p ps=0u
M1002 X a_222_367# VGND VNB nshort w=840000u l=150000u
+  ad=2.352e+11p pd=2.24e+06u as=6.51e+11p ps=6.24e+06u
M1003 a_67_47# B2 VGND VNB nshort w=420000u l=150000u
+  ad=2.289e+11p pd=2.77e+06u as=0p ps=0u
M1004 VGND B1 a_67_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VPWR a_222_367# X VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=3.528e+11p ps=3.08e+06u
M1006 VGND a_222_367# X VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR a_300_21# a_222_367# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=2.496e+11p ps=2.06e+06u
M1008 VPWR A1_N a_300_21# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_222_367# a_300_21# a_67_47# VNB nshort w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1010 a_222_367# B2 a_150_367# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_585_47# A2_N a_300_21# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=1.113e+11p ps=1.37e+06u
M1012 VGND A1_N a_585_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 X a_222_367# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
