* File: sky130_fd_sc_lp__decapkapwr_12.spice
* Created: Fri Aug 28 10:20:20 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__decapkapwr_12.pex.spice"
.subckt sky130_fd_sc_lp__decapkapwr_12  VNB VPB VGND KAPWR VPWR
* 
* KAPWR	KAPWR
* VGND	VGND
* VPB	VPB
* VNB	VNB
MM1000 N_VGND_M1000_s N_KAPWR_M1000_g N_VGND_M1000_s VNB NSHORT L=4 W=1 AD=0.285
+ AS=0.265 PD=2.57 PS=2.53 NRD=0 NRS=0 M=1 R=0.25 SA=2e+06 SB=2e+06 A=4 P=10
+ MULT=1
MM1001 N_KAPWR_M1001_s N_VGND_M1001_g N_KAPWR_M1001_s VPB PHIGHVT L=4 W=1
+ AD=0.285 AS=0.275 PD=2.57 PS=2.55 NRD=0 NRS=1.9503 M=1 R=0.25 SA=2e+06
+ SB=2e+06 A=4 P=10 MULT=1
DX2_noxref VNB VPB NWDIODE A=11.4511 P=16.01
*
.include "sky130_fd_sc_lp__decapkapwr_12.pxi.spice"
*
.ends
*
*
