* File: sky130_fd_sc_lp__sdfstp_4.spice
* Created: Fri Aug 28 11:29:51 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__sdfstp_4.pex.spice"
.subckt sky130_fd_sc_lp__sdfstp_4  VNB VPB SCD D SCE CLK SET_B VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* SET_B	SET_B
* CLK	CLK
* SCE	SCE
* D	D
* SCD	SCD
* VPB	VPB
* VNB	VNB
MM1014 A_146_119# N_SCD_M1014_g N_VGND_M1014_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1113 PD=0.63 PS=1.37 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.8 A=0.063 P=1.14 MULT=1
MM1009 N_A_218_119#_M1009_d N_SCE_M1009_g A_146_119# VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1013 A_304_119# N_D_M1013_g N_A_218_119#_M1009_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75001 SB=75001
+ A=0.063 P=1.14 MULT=1
MM1000 N_VGND_M1000_d N_A_346_93#_M1000_g A_304_119# VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.3
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1001 N_A_346_93#_M1001_d N_SCE_M1001_g N_VGND_M1000_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.8 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1037 N_VGND_M1037_d N_CLK_M1037_g N_A_773_409#_M1037_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1005 N_A_961_491#_M1005_d N_A_773_409#_M1005_g N_VGND_M1037_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.6 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1041 N_A_1211_463#_M1041_d N_A_773_409#_M1041_g N_A_218_119#_M1041_s VNB
+ NSHORT L=0.15 W=0.42 AD=0.0588 AS=0.2667 PD=0.7 PS=2.11 NRD=0 NRS=97.14 M=1
+ R=2.8 SA=75000.6 SB=75001 A=0.063 P=1.14 MULT=1
MM1008 A_1315_81# N_A_961_491#_M1008_g N_A_1211_463#_M1041_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75001
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1011 N_VGND_M1011_d N_A_1339_331#_M1011_g A_1315_81# VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.0441 PD=1.37 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.3
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1027 A_1598_125# N_A_1211_463#_M1027_g N_A_1339_331#_M1027_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.1113 PD=0.63 PS=1.37 NRD=14.28 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75004.5 A=0.063 P=1.14 MULT=1
MM1032 N_VGND_M1032_d N_SET_B_M1032_g A_1598_125# VNB NSHORT L=0.15 W=0.42
+ AD=0.17953 AS=0.0441 PD=1.25208 PS=0.63 NRD=106.404 NRS=14.28 M=1 R=2.8
+ SA=75000.6 SB=75004.1 A=0.063 P=1.14 MULT=1
MM1028 A_1888_125# N_A_1211_463#_M1028_g N_VGND_M1032_d VNB NSHORT L=0.15 W=0.64
+ AD=0.0672 AS=0.27357 PD=0.85 PS=1.90792 NRD=9.372 NRS=69.828 M=1 R=4.26667
+ SA=75001.1 SB=75002.3 A=0.096 P=1.58 MULT=1
MM1035 N_A_1960_125#_M1035_d N_A_961_491#_M1035_g A_1888_125# VNB NSHORT L=0.15
+ W=0.64 AD=0.319638 AS=0.0672 PD=1.81736 PS=0.85 NRD=2.808 NRS=9.372 M=1
+ R=4.26667 SA=75001.5 SB=75002 A=0.096 P=1.58 MULT=1
MM1020 A_2163_125# N_A_773_409#_M1020_g N_A_1960_125#_M1035_d VNB NSHORT L=0.15
+ W=0.42 AD=0.05775 AS=0.209762 PD=0.695 PS=1.19264 NRD=23.568 NRS=28.56 M=1
+ R=2.8 SA=75003 SB=75001.6 A=0.063 P=1.14 MULT=1
MM1016 A_2248_125# N_A_2205_231#_M1016_g A_2163_125# VNB NSHORT L=0.15 W=0.42
+ AD=0.06825 AS=0.05775 PD=0.745 PS=0.695 NRD=30.708 NRS=23.568 M=1 R=2.8
+ SA=75003.4 SB=75001.2 A=0.063 P=1.14 MULT=1
MM1024 N_VGND_M1024_d N_SET_B_M1024_g A_2248_125# VNB NSHORT L=0.15 W=0.42
+ AD=0.0819 AS=0.06825 PD=0.81 PS=0.745 NRD=15.708 NRS=30.708 M=1 R=2.8
+ SA=75003.9 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1043 N_A_2205_231#_M1043_d N_A_1960_125#_M1043_g N_VGND_M1024_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.1113 AS=0.0819 PD=1.37 PS=0.81 NRD=0 NRS=15.708 M=1 R=2.8
+ SA=75004.5 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1007 N_VGND_M1007_d N_A_1960_125#_M1007_g N_A_2638_53#_M1007_s VNB NSHORT
+ L=0.15 W=0.84 AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6
+ SA=75000.2 SB=75001.9 A=0.126 P=1.98 MULT=1
MM1004 N_VGND_M1007_d N_A_2638_53#_M1004_g N_Q_M1004_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75001.5 A=0.126 P=1.98 MULT=1
MM1030 N_VGND_M1030_d N_A_2638_53#_M1030_g N_Q_M1004_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.1
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1036 N_VGND_M1030_d N_A_2638_53#_M1036_g N_Q_M1036_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.5
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1045 N_VGND_M1045_d N_A_2638_53#_M1045_g N_Q_M1036_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.9
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1038 N_VPWR_M1038_d N_SCD_M1038_g N_A_27_479#_M1038_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.0896 AS=0.1696 PD=0.92 PS=1.81 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75001.5 A=0.096 P=1.58 MULT=1
MM1012 A_196_479# N_SCE_M1012_g N_VPWR_M1038_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0672 AS=0.0896 PD=0.85 PS=0.92 NRD=15.3857 NRS=0 M=1 R=4.26667 SA=75000.6
+ SB=75001.1 A=0.096 P=1.58 MULT=1
MM1017 N_A_218_119#_M1017_d N_D_M1017_g A_196_479# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1248 AS=0.0672 PD=1.03 PS=0.85 NRD=16.9223 NRS=15.3857 M=1 R=4.26667
+ SA=75001 SB=75000.7 A=0.096 P=1.58 MULT=1
MM1031 N_A_27_479#_M1031_d N_A_346_93#_M1031_g N_A_218_119#_M1017_d VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.1696 AS=0.1248 PD=1.81 PS=1.03 NRD=0 NRS=16.9223 M=1
+ R=4.26667 SA=75001.5 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1039 N_A_346_93#_M1039_d N_SCE_M1039_g N_VPWR_M1039_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1696 AS=0.3424 PD=1.81 PS=2.35 NRD=0 NRS=83.0946 M=1 R=4.26667
+ SA=75000.5 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1042 N_VPWR_M1042_d N_CLK_M1042_g N_A_773_409#_M1042_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.0896 AS=0.3329 PD=0.92 PS=2.82 NRD=0 NRS=143.18 M=1 R=4.26667
+ SA=75000.3 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1023 N_A_961_491#_M1023_d N_A_773_409#_M1023_g N_VPWR_M1042_d VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.1696 AS=0.0896 PD=1.81 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.7 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1033 N_A_1211_463#_M1033_d N_A_961_491#_M1033_g N_A_218_119#_M1033_s VPB
+ PHIGHVT L=0.15 W=0.42 AD=0.0588 AS=0.2247 PD=0.7 PS=1.91 NRD=0 NRS=126.632 M=1
+ R=2.8 SA=75000.5 SB=75002.9 A=0.063 P=1.14 MULT=1
MM1022 A_1297_463# N_A_773_409#_M1022_g N_A_1211_463#_M1033_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=23.443 NRS=0 M=1 R=2.8
+ SA=75000.9 SB=75002.5 A=0.063 P=1.14 MULT=1
MM1025 N_VPWR_M1025_d N_A_1339_331#_M1025_g A_1297_463# VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1155 AS=0.0441 PD=0.97 PS=0.63 NRD=0 NRS=23.443 M=1 R=2.8
+ SA=75001.2 SB=75002.1 A=0.063 P=1.14 MULT=1
MM1029 N_A_1339_331#_M1029_d N_A_1211_463#_M1029_g N_VPWR_M1025_d VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.0672 AS=0.1155 PD=0.74 PS=0.97 NRD=0 NRS=126.632 M=1 R=2.8
+ SA=75001.9 SB=75001.4 A=0.063 P=1.14 MULT=1
MM1018 N_VPWR_M1018_d N_SET_B_M1018_g N_A_1339_331#_M1029_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1197 AS=0.0672 PD=0.953333 PS=0.74 NRD=145.386 NRS=18.7544 M=1
+ R=2.8 SA=75002.4 SB=75000.9 A=0.063 P=1.14 MULT=1
MM1010 N_A_1751_379#_M1010_d N_A_1211_463#_M1010_g N_VPWR_M1018_d VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.2226 AS=0.2394 PD=2.21 PS=1.90667 NRD=0 NRS=0 M=1 R=5.6
+ SA=75001.7 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1026 N_A_1960_125#_M1026_d N_A_961_491#_M1026_g N_A_1858_463#_M1026_s VPB
+ PHIGHVT L=0.15 W=0.42 AD=0.0896 AS=0.1887 PD=0.81 PS=1.86 NRD=74.2493
+ NRS=46.886 M=1 R=2.8 SA=75000.3 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1002 N_A_1751_379#_M1002_d N_A_773_409#_M1002_g N_A_1960_125#_M1026_d VPB
+ PHIGHVT L=0.15 W=0.84 AD=0.2226 AS=0.1792 PD=2.21 PS=1.62 NRD=0 NRS=0 M=1
+ R=5.6 SA=75000.5 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1019 N_VPWR_M1019_d N_A_2205_231#_M1019_g N_A_1858_463#_M1019_s VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1003 N_A_1960_125#_M1003_d N_SET_B_M1003_g N_VPWR_M1019_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1015 N_A_2205_231#_M1015_d N_A_1960_125#_M1015_g N_VPWR_M1015_s VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.1113 AS=0.1113 PD=1.37 PS=1.37 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1040 N_VPWR_M1040_d N_A_1960_125#_M1040_g N_A_2638_53#_M1040_s VPB PHIGHVT
+ L=0.15 W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.2 SB=75001.9 A=0.189 P=2.82 MULT=1
MM1006 N_VPWR_M1040_d N_A_2638_53#_M1006_g N_Q_M1006_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75001.5 A=0.189 P=2.82 MULT=1
MM1021 N_VPWR_M1021_d N_A_2638_53#_M1021_g N_Q_M1006_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1034 N_VPWR_M1021_d N_A_2638_53#_M1034_g N_Q_M1034_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.5
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1044 N_VPWR_M1044_d N_A_2638_53#_M1044_g N_Q_M1034_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.9
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX46_noxref VNB VPB NWDIODE A=30.2503 P=36.17
c_285 VPB 0 1.88632e-19 $X=0 $Y=3.085
c_2123 A_1598_125# 0 1.52906e-19 $X=7.99 $Y=0.625
*
.include "sky130_fd_sc_lp__sdfstp_4.pxi.spice"
*
.ends
*
*
