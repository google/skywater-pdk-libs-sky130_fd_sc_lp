* File: sky130_fd_sc_lp__nand4_lp.pex.spice
* Created: Wed Sep  2 10:05:48 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__NAND4_LP%D 3 7 9 12 13
r28 12 15 71.8729 $w=4.7e-07 $l=5.05e-07 $layer=POLY_cond $X=0.455 $Y=0.99
+ $X2=0.455 $Y2=1.495
r29 12 14 47.4991 $w=4.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.455 $Y=0.99
+ $X2=0.455 $Y2=0.825
r30 12 13 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.385
+ $Y=0.99 $X2=0.385 $Y2=0.99
r31 9 13 2.58853 $w=6.68e-07 $l=1.45e-07 $layer=LI1_cond $X=0.24 $Y=1.16
+ $X2=0.385 $Y2=1.16
r32 7 14 194.851 $w=1.5e-07 $l=3.8e-07 $layer=POLY_cond $X=0.585 $Y=0.445
+ $X2=0.585 $Y2=0.825
r33 3 15 260.876 $w=2.5e-07 $l=1.05e-06 $layer=POLY_cond $X=0.565 $Y=2.545
+ $X2=0.565 $Y2=1.495
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4_LP%C 3 6 9 10 11 12 13 14 19
c43 11 0 6.48616e-20 $X=1.065 $Y=1.435
r44 19 20 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.065
+ $Y=0.93 $X2=1.065 $Y2=0.93
r45 14 20 10.7857 $w=3.88e-07 $l=3.65e-07 $layer=LI1_cond $X=1.095 $Y=1.295
+ $X2=1.095 $Y2=0.93
r46 13 20 0.147749 $w=3.88e-07 $l=5e-09 $layer=LI1_cond $X=1.095 $Y=0.925
+ $X2=1.095 $Y2=0.93
r47 12 13 10.9334 $w=3.88e-07 $l=3.7e-07 $layer=LI1_cond $X=1.095 $Y=0.555
+ $X2=1.095 $Y2=0.925
r48 10 19 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.065 $Y=1.27
+ $X2=1.065 $Y2=0.93
r49 10 11 31.6748 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.065 $Y=1.27
+ $X2=1.065 $Y2=1.435
r50 9 19 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.065 $Y=0.765
+ $X2=1.065 $Y2=0.93
r51 6 11 275.784 $w=2.5e-07 $l=1.11e-06 $layer=POLY_cond $X=1.095 $Y=2.545
+ $X2=1.095 $Y2=1.435
r52 3 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.975 $Y=0.445
+ $X2=0.975 $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4_LP%B 3 4 6 9 10 11 12 13 18
c44 18 0 2.64121e-20 $X=1.635 $Y=0.93
c45 6 0 5.18852e-20 $X=1.635 $Y=2.545
r46 12 13 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.635 $Y=0.925
+ $X2=1.635 $Y2=1.295
r47 12 18 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.635
+ $Y=0.93 $X2=1.635 $Y2=0.93
r48 11 12 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.635 $Y=0.555
+ $X2=1.635 $Y2=0.925
r49 10 18 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.635 $Y=1.27
+ $X2=1.635 $Y2=0.93
r50 9 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.635 $Y=0.765
+ $X2=1.635 $Y2=0.93
r51 4 10 30.6163 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.635 $Y=1.435
+ $X2=1.635 $Y2=1.27
r52 4 6 275.784 $w=2.5e-07 $l=1.11e-06 $layer=POLY_cond $X=1.635 $Y=1.435
+ $X2=1.635 $Y2=2.545
r53 3 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.545 $Y=0.445
+ $X2=1.545 $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4_LP%A 3 7 9 10 14 15
c30 15 0 5.18852e-20 $X=2.495 $Y=1.275
r31 14 17 63.2352 $w=6.2e-07 $l=5.05e-07 $layer=POLY_cond $X=2.35 $Y=1.275
+ $X2=2.35 $Y2=1.78
r32 14 16 50.0851 $w=6.2e-07 $l=1.65e-07 $layer=POLY_cond $X=2.35 $Y=1.275
+ $X2=2.35 $Y2=1.11
r33 14 15 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.495
+ $Y=1.275 $X2=2.495 $Y2=1.275
r34 9 10 10.033 $w=4.23e-07 $l=3.7e-07 $layer=LI1_cond $X=2.542 $Y=1.295
+ $X2=2.542 $Y2=1.665
r35 9 15 0.542326 $w=4.23e-07 $l=2e-08 $layer=LI1_cond $X=2.542 $Y=1.295
+ $X2=2.542 $Y2=1.275
r36 7 17 190.067 $w=2.5e-07 $l=7.65e-07 $layer=POLY_cond $X=2.165 $Y=2.545
+ $X2=2.165 $Y2=1.78
r37 3 16 340.989 $w=1.5e-07 $l=6.65e-07 $layer=POLY_cond $X=2.115 $Y=0.445
+ $X2=2.115 $Y2=1.11
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4_LP%VPWR 1 2 3 10 12 16 20 24 26 30 32 41 45
r38 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r39 41 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r40 39 42 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.2 $Y2=3.33
r41 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r42 36 45 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r43 35 36 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r44 33 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.525 $Y=3.33
+ $X2=1.36 $Y2=3.33
r45 33 35 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=1.525 $Y=3.33
+ $X2=2.16 $Y2=3.33
r46 32 44 4.54404 $w=1.7e-07 $l=2.75e-07 $layer=LI1_cond $X=2.33 $Y=3.33
+ $X2=2.605 $Y2=3.33
r47 32 35 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=2.33 $Y=3.33
+ $X2=2.16 $Y2=3.33
r48 30 36 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=2.16 $Y2=3.33
r49 30 42 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.44 $Y=3.33
+ $X2=1.2 $Y2=3.33
r50 26 29 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=2.495 $Y=2.19
+ $X2=2.495 $Y2=2.9
r51 24 44 3.22214 $w=3.3e-07 $l=1.46458e-07 $layer=LI1_cond $X=2.495 $Y=3.245
+ $X2=2.605 $Y2=3.33
r52 24 29 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=2.495 $Y=3.245
+ $X2=2.495 $Y2=2.9
r53 20 23 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=1.36 $Y=2.19 $X2=1.36
+ $Y2=2.9
r54 18 41 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.36 $Y=3.245
+ $X2=1.36 $Y2=3.33
r55 18 23 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=1.36 $Y=3.245
+ $X2=1.36 $Y2=2.9
r56 17 38 4.68787 $w=1.7e-07 $l=2.33e-07 $layer=LI1_cond $X=0.465 $Y=3.33
+ $X2=0.232 $Y2=3.33
r57 16 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.195 $Y=3.33
+ $X2=1.36 $Y2=3.33
r58 16 17 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=1.195 $Y=3.33
+ $X2=0.465 $Y2=3.33
r59 12 15 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=0.3 $Y=2.19 $X2=0.3
+ $Y2=2.9
r60 10 38 3.0783 $w=3.3e-07 $l=1.14039e-07 $layer=LI1_cond $X=0.3 $Y=3.245
+ $X2=0.232 $Y2=3.33
r61 10 15 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=0.3 $Y=3.245
+ $X2=0.3 $Y2=2.9
r62 3 29 400 $w=1.7e-07 $l=9.51998e-07 $layer=licon1_PDIFF $count=1 $X=2.29
+ $Y=2.045 $X2=2.495 $Y2=2.9
r63 3 26 400 $w=1.7e-07 $l=2.67862e-07 $layer=licon1_PDIFF $count=1 $X=2.29
+ $Y=2.045 $X2=2.495 $Y2=2.19
r64 2 23 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=1.22
+ $Y=2.045 $X2=1.36 $Y2=2.9
r65 2 20 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.22
+ $Y=2.045 $X2=1.36 $Y2=2.19
r66 1 15 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.155
+ $Y=2.045 $X2=0.3 $Y2=2.9
r67 1 12 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.155
+ $Y=2.045 $X2=0.3 $Y2=2.19
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4_LP%Y 1 2 3 12 16 17 20 24 25 26 27 28 34
c56 25 0 1.89209e-19 $X=2.065 $Y=1.675
c57 24 0 1.38359e-19 $X=2.065 $Y=0.675
c58 16 0 6.48616e-20 $X=1.735 $Y=1.76
r59 32 34 0.281084 $w=4.08e-07 $l=1e-08 $layer=LI1_cond $X=2.15 $Y=0.47 $X2=2.16
+ $Y2=0.47
r60 28 37 8.71359 $w=4.08e-07 $l=3.1e-07 $layer=LI1_cond $X=2.64 $Y=0.47
+ $X2=2.33 $Y2=0.47
r61 27 32 2.47908 $w=4.1e-07 $l=8.5e-08 $layer=LI1_cond $X=2.065 $Y=0.47
+ $X2=2.15 $Y2=0.47
r62 27 37 3.73841 $w=4.08e-07 $l=1.33e-07 $layer=LI1_cond $X=2.197 $Y=0.47
+ $X2=2.33 $Y2=0.47
r63 27 34 1.04001 $w=4.08e-07 $l=3.7e-08 $layer=LI1_cond $X=2.197 $Y=0.47
+ $X2=2.16 $Y2=0.47
r64 25 26 3.22182 $w=2.92e-07 $l=1.5995e-07 $layer=LI1_cond $X=2.065 $Y=1.675
+ $X2=1.942 $Y2=1.76
r65 24 27 5.97895 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=2.065 $Y=0.675
+ $X2=2.065 $Y2=0.47
r66 24 25 65.2406 $w=1.68e-07 $l=1e-06 $layer=LI1_cond $X=2.065 $Y=0.675
+ $X2=2.065 $Y2=1.675
r67 20 22 19.7165 $w=4.13e-07 $l=7.1e-07 $layer=LI1_cond $X=1.942 $Y=2.19
+ $X2=1.942 $Y2=2.9
r68 18 26 3.22182 $w=2.92e-07 $l=8.5e-08 $layer=LI1_cond $X=1.942 $Y=1.845
+ $X2=1.942 $Y2=1.76
r69 18 20 9.58055 $w=4.13e-07 $l=3.45e-07 $layer=LI1_cond $X=1.942 $Y=1.845
+ $X2=1.942 $Y2=2.19
r70 16 26 3.35233 $w=1.7e-07 $l=2.07e-07 $layer=LI1_cond $X=1.735 $Y=1.76
+ $X2=1.942 $Y2=1.76
r71 16 17 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=1.735 $Y=1.76
+ $X2=0.995 $Y2=1.76
r72 12 14 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=0.83 $Y=2.19 $X2=0.83
+ $Y2=2.9
r73 10 17 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.83 $Y=1.845
+ $X2=0.995 $Y2=1.76
r74 10 12 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=0.83 $Y=1.845
+ $X2=0.83 $Y2=2.19
r75 3 22 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=1.76
+ $Y=2.045 $X2=1.9 $Y2=2.9
r76 3 20 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.76
+ $Y=2.045 $X2=1.9 $Y2=2.19
r77 2 14 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=0.69
+ $Y=2.045 $X2=0.83 $Y2=2.9
r78 2 12 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.69
+ $Y=2.045 $X2=0.83 $Y2=2.19
r79 1 37 182 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=1 $X=2.19
+ $Y=0.235 $X2=2.33 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_LP__NAND4_LP%VGND 1 4 6 8 15 16
c33 16 0 2.64121e-20 $X=2.64 $Y=0
r34 19 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r35 15 16 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r36 13 20 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r37 12 15 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=0.72 $Y=0 $X2=2.64
+ $Y2=0
r38 12 13 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r39 10 19 4.56433 $w=1.7e-07 $l=2.68e-07 $layer=LI1_cond $X=0.535 $Y=0 $X2=0.267
+ $Y2=0
r40 10 12 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=0.535 $Y=0 $X2=0.72
+ $Y2=0
r41 8 16 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=1.44 $Y=0 $X2=2.64
+ $Y2=0
r42 8 13 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.44 $Y=0 $X2=0.72
+ $Y2=0
r43 4 19 3.20184 $w=3.3e-07 $l=1.39155e-07 $layer=LI1_cond $X=0.37 $Y=0.085
+ $X2=0.267 $Y2=0
r44 4 6 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=0.37 $Y=0.085
+ $X2=0.37 $Y2=0.43
r45 1 6 182 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_NDIFF $count=1 $X=0.225
+ $Y=0.235 $X2=0.37 $Y2=0.43
.ends

