* File: sky130_fd_sc_lp__dlrtn_1.pex.spice
* Created: Wed Sep  2 09:46:50 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__DLRTN_1%D 3 5 8 10 11 12 13 14 20 22
r38 20 22 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=0.687 $Y=0.93
+ $X2=0.687 $Y2=0.765
r39 13 14 21.5981 $w=1.88e-07 $l=3.7e-07 $layer=LI1_cond $X=0.72 $Y=1.295
+ $X2=0.72 $Y2=1.665
r40 12 13 21.5981 $w=1.88e-07 $l=3.7e-07 $layer=LI1_cond $X=0.72 $Y=0.925
+ $X2=0.72 $Y2=1.295
r41 12 20 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.71
+ $Y=0.93 $X2=0.71 $Y2=0.93
r42 11 12 21.5981 $w=1.88e-07 $l=3.7e-07 $layer=LI1_cond $X=0.72 $Y=0.555
+ $X2=0.72 $Y2=0.925
r43 8 10 620.447 $w=1.5e-07 $l=1.21e-06 $layer=POLY_cond $X=0.575 $Y=2.645
+ $X2=0.575 $Y2=1.435
r44 5 10 48.4185 $w=3.75e-07 $l=1.87e-07 $layer=POLY_cond $X=0.687 $Y=1.248
+ $X2=0.687 $Y2=1.435
r45 4 20 3.26277 $w=3.75e-07 $l=2.2e-08 $layer=POLY_cond $X=0.687 $Y=0.952
+ $X2=0.687 $Y2=0.93
r46 4 5 43.8991 $w=3.75e-07 $l=2.96e-07 $layer=POLY_cond $X=0.687 $Y=0.952
+ $X2=0.687 $Y2=1.248
r47 3 22 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.575 $Y=0.445
+ $X2=0.575 $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_LP__DLRTN_1%GATE_N 2 3 5 6 8 11 13 14 15
c44 11 0 2.16337e-19 $X=1.285 $Y=0.84
r45 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.07
+ $Y=1.84 $X2=1.07 $Y2=1.84
r46 15 21 5.93169 $w=3.38e-07 $l=1.75e-07 $layer=LI1_cond $X=1.155 $Y=1.665
+ $X2=1.155 $Y2=1.84
r47 14 15 12.5413 $w=3.38e-07 $l=3.7e-07 $layer=LI1_cond $X=1.155 $Y=1.295
+ $X2=1.155 $Y2=1.665
r48 13 14 12.5413 $w=3.38e-07 $l=3.7e-07 $layer=LI1_cond $X=1.155 $Y=0.925
+ $X2=1.155 $Y2=1.295
r49 9 11 64.0957 $w=1.5e-07 $l=1.25e-07 $layer=POLY_cond $X=1.16 $Y=0.84
+ $X2=1.285 $Y2=0.84
r50 6 11 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.285 $Y=0.765
+ $X2=1.285 $Y2=0.84
r51 6 8 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.285 $Y=0.765
+ $X2=1.285 $Y2=0.445
r52 3 20 73.3907 $w=2.91e-07 $l=4.4286e-07 $layer=POLY_cond $X=1.275 $Y=2.215
+ $X2=1.127 $Y2=1.84
r53 3 5 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=1.275 $Y=2.215
+ $X2=1.275 $Y2=2.645
r54 2 20 38.6072 $w=2.91e-07 $l=1.80748e-07 $layer=POLY_cond $X=1.16 $Y=1.675
+ $X2=1.127 $Y2=1.84
r55 1 9 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.16 $Y=0.915 $X2=1.16
+ $Y2=0.84
r56 1 2 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=1.16 $Y=0.915 $X2=1.16
+ $Y2=1.675
.ends

.subckt PM_SKY130_FD_SC_LP__DLRTN_1%A_47_47# 1 2 9 13 17 21 23 26 27 28 30 31 32
+ 35 36 38
c97 35 0 1.19672e-19 $X=2.825 $Y=1.52
c98 13 0 1.09969e-19 $X=2.915 $Y=2.555
c99 9 0 1.17792e-20 $X=2.915 $Y=0.835
r100 36 41 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.825 $Y=1.52
+ $X2=2.825 $Y2=1.685
r101 36 40 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.825 $Y=1.52
+ $X2=2.825 $Y2=1.355
r102 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.825
+ $Y=1.52 $X2=2.825 $Y2=1.52
r103 33 35 27.7634 $w=3.28e-07 $l=7.95e-07 $layer=LI1_cond $X=2.825 $Y=2.315
+ $X2=2.825 $Y2=1.52
r104 31 33 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.66 $Y=2.4
+ $X2=2.825 $Y2=2.315
r105 31 32 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=2.66 $Y=2.4
+ $X2=2.045 $Y2=2.4
r106 29 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.96 $Y=2.485
+ $X2=2.045 $Y2=2.4
r107 29 30 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=1.96 $Y=2.485
+ $X2=1.96 $Y2=2.815
r108 27 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.875 $Y=2.9
+ $X2=1.96 $Y2=2.815
r109 27 28 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=1.875 $Y=2.9
+ $X2=1.235 $Y2=2.9
r110 26 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.15 $Y=2.815
+ $X2=1.235 $Y2=2.9
r111 25 26 30.6631 $w=1.68e-07 $l=4.7e-07 $layer=LI1_cond $X=1.15 $Y=2.345
+ $X2=1.15 $Y2=2.815
r112 24 38 2.98021 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=0.465 $Y=2.26
+ $X2=0.33 $Y2=2.26
r113 23 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.065 $Y=2.26
+ $X2=1.15 $Y2=2.345
r114 23 24 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=1.065 $Y=2.26
+ $X2=0.465 $Y2=2.26
r115 19 38 3.52026 $w=2.65e-07 $l=8.5e-08 $layer=LI1_cond $X=0.33 $Y=2.345
+ $X2=0.33 $Y2=2.26
r116 19 21 5.33538 $w=2.68e-07 $l=1.25e-07 $layer=LI1_cond $X=0.33 $Y=2.345
+ $X2=0.33 $Y2=2.47
r117 15 38 3.52026 $w=2.65e-07 $l=8.74643e-08 $layer=LI1_cond $X=0.325 $Y=2.175
+ $X2=0.33 $Y2=2.26
r118 15 17 75.7953 $w=2.58e-07 $l=1.71e-06 $layer=LI1_cond $X=0.325 $Y=2.175
+ $X2=0.325 $Y2=0.465
r119 13 41 446.106 $w=1.5e-07 $l=8.7e-07 $layer=POLY_cond $X=2.915 $Y=2.555
+ $X2=2.915 $Y2=1.685
r120 9 40 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=2.915 $Y=0.835
+ $X2=2.915 $Y2=1.355
r121 2 21 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.235
+ $Y=2.325 $X2=0.36 $Y2=2.47
r122 1 17 182 $w=1.7e-07 $l=2.85745e-07 $layer=licon1_NDIFF $count=1 $X=0.235
+ $Y=0.235 $X2=0.36 $Y2=0.465
.ends

.subckt PM_SKY130_FD_SC_LP__DLRTN_1%A_387_385# 1 2 9 13 16 20 22 25 26 28 29 31
+ 33 34 36 45
c99 31 0 1.77834e-19 $X=3.33 $Y=1.265
c100 20 0 1.09969e-19 $X=2.08 $Y=2.06
r101 34 42 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.365 $Y=1.91
+ $X2=3.365 $Y2=2.075
r102 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.365
+ $Y=1.91 $X2=3.365 $Y2=1.91
r103 31 33 28.5895 $w=2.58e-07 $l=6.45e-07 $layer=LI1_cond $X=3.33 $Y=1.265
+ $X2=3.33 $Y2=1.91
r104 29 45 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.725 $Y=0.35
+ $X2=3.725 $Y2=0.515
r105 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.725
+ $Y=0.35 $X2=3.725 $Y2=0.35
r106 26 28 27.8507 $w=2.38e-07 $l=5.8e-07 $layer=LI1_cond $X=3.145 $Y=0.375
+ $X2=3.725 $Y2=0.375
r107 25 31 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=3.035 $Y=1.18
+ $X2=3.33 $Y2=1.18
r108 24 26 6.83327 $w=2.4e-07 $l=1.66132e-07 $layer=LI1_cond $X=3.035 $Y=0.495
+ $X2=3.145 $Y2=0.375
r109 24 25 31.4303 $w=2.18e-07 $l=6e-07 $layer=LI1_cond $X=3.035 $Y=0.495
+ $X2=3.035 $Y2=1.095
r110 23 36 3.80956 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.245 $Y=1.18
+ $X2=2.08 $Y2=1.18
r111 22 25 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=2.925 $Y=1.18
+ $X2=3.035 $Y2=1.18
r112 22 23 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=2.925 $Y=1.18
+ $X2=2.245 $Y2=1.18
r113 18 36 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.08 $Y=1.265
+ $X2=2.08 $Y2=1.18
r114 18 20 27.7634 $w=3.28e-07 $l=7.95e-07 $layer=LI1_cond $X=2.08 $Y=1.265
+ $X2=2.08 $Y2=2.06
r115 14 36 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.08 $Y=1.095
+ $X2=2.08 $Y2=1.18
r116 14 16 8.55602 $w=3.28e-07 $l=2.45e-07 $layer=LI1_cond $X=2.08 $Y=1.095
+ $X2=2.08 $Y2=0.85
r117 13 45 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=3.705 $Y=0.835
+ $X2=3.705 $Y2=0.515
r118 9 42 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=3.275 $Y=2.555
+ $X2=3.275 $Y2=2.075
r119 2 20 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.935
+ $Y=1.925 $X2=2.08 $Y2=2.06
r120 1 16 182 $w=1.7e-07 $l=2.80624e-07 $layer=licon1_NDIFF $count=1 $X=2.015
+ $Y=0.625 $X2=2.14 $Y2=0.85
.ends

.subckt PM_SKY130_FD_SC_LP__DLRTN_1%A_270_465# 1 2 8 9 10 11 13 16 19 21 22 26
+ 32 37 40 45
c103 21 0 1.79834e-19 $X=3.275 $Y=0.835
c104 19 0 1.19672e-19 $X=3.275 $Y=1.155
r105 45 46 2.45203 $w=6.88e-07 $l=3.5e-08 $layer=POLY_cond $X=2.375 $Y=1.615
+ $X2=2.41 $Y2=1.615
r106 44 45 35.7297 $w=6.88e-07 $l=5.1e-07 $layer=POLY_cond $X=1.865 $Y=1.615
+ $X2=2.375 $Y2=1.615
r107 40 41 7.38866 $w=2.98e-07 $l=1.65e-07 $layer=LI1_cond $X=1.555 $Y=2.47
+ $X2=1.555 $Y2=2.305
r108 35 37 3.49225 $w=3.28e-07 $l=1e-07 $layer=LI1_cond $X=1.5 $Y=0.465 $X2=1.6
+ $Y2=0.465
r109 33 44 17.8648 $w=6.88e-07 $l=2.55e-07 $layer=POLY_cond $X=1.61 $Y=1.615
+ $X2=1.865 $Y2=1.615
r110 32 41 52.0216 $w=2.08e-07 $l=9.85e-07 $layer=LI1_cond $X=1.6 $Y=1.32
+ $X2=1.6 $Y2=2.305
r111 32 33 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.61
+ $Y=1.32 $X2=1.61 $Y2=1.32
r112 29 37 3.38185 $w=2.1e-07 $l=1.65e-07 $layer=LI1_cond $X=1.6 $Y=0.63 $X2=1.6
+ $Y2=0.465
r113 29 32 36.4416 $w=2.08e-07 $l=6.9e-07 $layer=LI1_cond $X=1.6 $Y=0.63 $X2=1.6
+ $Y2=1.32
r114 24 26 466.617 $w=1.5e-07 $l=9.1e-07 $layer=POLY_cond $X=3.815 $Y=1.535
+ $X2=3.815 $Y2=2.445
r115 23 28 4.52116 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.38 $Y=1.46 $X2=3.29
+ $Y2=1.46
r116 22 24 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.74 $Y=1.46
+ $X2=3.815 $Y2=1.535
r117 22 23 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=3.74 $Y=1.46
+ $X2=3.38 $Y2=1.46
r118 19 28 91.6059 $w=1.61e-07 $l=3.1241e-07 $layer=POLY_cond $X=3.275 $Y=1.155
+ $X2=3.29 $Y2=1.46
r119 19 21 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=3.275 $Y=1.155
+ $X2=3.275 $Y2=0.835
r120 18 21 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=3.275 $Y=0.255
+ $X2=3.275 $Y2=0.835
r121 14 46 39.6551 $w=1.5e-07 $l=4.6e-07 $layer=POLY_cond $X=2.41 $Y=2.075
+ $X2=2.41 $Y2=1.615
r122 14 16 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.41 $Y=2.075
+ $X2=2.41 $Y2=2.555
r123 11 45 39.6551 $w=1.5e-07 $l=4.6e-07 $layer=POLY_cond $X=2.375 $Y=1.155
+ $X2=2.375 $Y2=1.615
r124 11 13 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.375 $Y=1.155
+ $X2=2.375 $Y2=0.835
r125 9 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.2 $Y=0.18
+ $X2=3.275 $Y2=0.255
r126 9 10 646.085 $w=1.5e-07 $l=1.26e-06 $layer=POLY_cond $X=3.2 $Y=0.18
+ $X2=1.94 $Y2=0.18
r127 8 44 39.6551 $w=1.5e-07 $l=4.6e-07 $layer=POLY_cond $X=1.865 $Y=1.155
+ $X2=1.865 $Y2=1.615
r128 7 10 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.865 $Y=0.255
+ $X2=1.94 $Y2=0.18
r129 7 8 461.489 $w=1.5e-07 $l=9e-07 $layer=POLY_cond $X=1.865 $Y=0.255
+ $X2=1.865 $Y2=1.155
r130 2 40 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.35
+ $Y=2.325 $X2=1.49 $Y2=2.47
r131 1 35 182 $w=1.7e-07 $l=2.91719e-07 $layer=licon1_NDIFF $count=1 $X=1.36
+ $Y=0.235 $X2=1.5 $Y2=0.465
.ends

.subckt PM_SKY130_FD_SC_LP__DLRTN_1%A_820_99# 1 2 9 13 17 21 25 26 27 30 32 35
+ 39 40 43 44 49 52 54
c115 30 0 1.73265e-19 $X=5.165 $Y=1.685
c116 9 0 1.77834e-19 $X=4.175 $Y=0.835
r117 49 51 15.7453 $w=5.08e-07 $l=4.45e-07 $layer=LI1_cond $X=5 $Y=0.43 $X2=5
+ $Y2=0.875
r118 43 46 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=4.265 $Y=1.57
+ $X2=4.265 $Y2=1.77
r119 43 44 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.265
+ $Y=1.57 $X2=4.265 $Y2=1.57
r120 40 58 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.115 $Y=1.51
+ $X2=6.115 $Y2=1.675
r121 40 57 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.115 $Y=1.51
+ $X2=6.115 $Y2=1.345
r122 39 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.115
+ $Y=1.51 $X2=6.115 $Y2=1.51
r123 37 39 36.4172 $w=2.48e-07 $l=7.9e-07 $layer=LI1_cond $X=6.075 $Y=2.3
+ $X2=6.075 $Y2=1.51
r124 36 54 2.53056 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=5.385 $Y=2.385
+ $X2=5.235 $Y2=2.385
r125 35 37 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=5.95 $Y=2.385
+ $X2=6.075 $Y2=2.3
r126 35 36 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=5.95 $Y=2.385
+ $X2=5.385 $Y2=2.385
r127 32 54 3.91525 $w=2.35e-07 $l=1.12916e-07 $layer=LI1_cond $X=5.17 $Y=2.3
+ $X2=5.235 $Y2=2.385
r128 31 52 5.04255 $w=1.75e-07 $l=8.74643e-08 $layer=LI1_cond $X=5.17 $Y=1.855
+ $X2=5.165 $Y2=1.77
r129 31 32 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=5.17 $Y=1.855
+ $X2=5.17 $Y2=2.3
r130 30 52 5.04255 $w=1.75e-07 $l=8.5e-08 $layer=LI1_cond $X=5.165 $Y=1.685
+ $X2=5.165 $Y2=1.77
r131 30 51 49.9091 $w=1.78e-07 $l=8.1e-07 $layer=LI1_cond $X=5.165 $Y=1.685
+ $X2=5.165 $Y2=0.875
r132 28 46 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.43 $Y=1.77
+ $X2=4.265 $Y2=1.77
r133 27 52 1.44715 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=5.075 $Y=1.77
+ $X2=5.165 $Y2=1.77
r134 27 28 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=5.075 $Y=1.77
+ $X2=4.43 $Y2=1.77
r135 25 44 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=4.265 $Y=1.91
+ $X2=4.265 $Y2=1.57
r136 25 26 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.265 $Y=1.91
+ $X2=4.265 $Y2=2.075
r137 24 44 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.265 $Y=1.405
+ $X2=4.265 $Y2=1.57
r138 21 58 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=6.025 $Y=2.465
+ $X2=6.025 $Y2=1.675
r139 17 57 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=6.025 $Y=0.655
+ $X2=6.025 $Y2=1.345
r140 13 26 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=4.175 $Y=2.445
+ $X2=4.175 $Y2=2.075
r141 9 24 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=4.175 $Y=0.835
+ $X2=4.175 $Y2=1.405
r142 2 54 300 $w=1.7e-07 $l=6.96491e-07 $layer=licon1_PDIFF $count=2 $X=5.13
+ $Y=1.835 $X2=5.27 $Y2=2.465
r143 1 49 91 $w=1.7e-07 $l=2.498e-07 $layer=licon1_NDIFF $count=2 $X=4.785
+ $Y=0.235 $X2=4.91 $Y2=0.43
.ends

.subckt PM_SKY130_FD_SC_LP__DLRTN_1%A_670_125# 1 2 9 11 13 14 19 22 26 30 31 33
+ 35
c91 33 0 1.79834e-19 $X=3.715 $Y=1.15
c92 31 0 1.17792e-20 $X=3.57 $Y=2.245
c93 19 0 1.91944e-19 $X=3.715 $Y=1.065
r94 35 36 11.0261 $w=3.06e-07 $l=7e-08 $layer=POLY_cond $X=5.055 $Y=1.35
+ $X2=5.125 $Y2=1.35
r95 30 31 8.50005 $w=4.58e-07 $l=1.35e-07 $layer=LI1_cond $X=3.57 $Y=2.38
+ $X2=3.57 $Y2=2.245
r96 27 35 37.0163 $w=3.06e-07 $l=2.35e-07 $layer=POLY_cond $X=4.82 $Y=1.35
+ $X2=5.055 $Y2=1.35
r97 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.82
+ $Y=1.35 $X2=4.82 $Y2=1.35
r98 24 26 5.30124 $w=2.48e-07 $l=1.15e-07 $layer=LI1_cond $X=4.78 $Y=1.235
+ $X2=4.78 $Y2=1.35
r99 23 33 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.8 $Y=1.15 $X2=3.715
+ $Y2=1.15
r100 22 24 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=4.655 $Y=1.15
+ $X2=4.78 $Y2=1.235
r101 22 23 55.7807 $w=1.68e-07 $l=8.55e-07 $layer=LI1_cond $X=4.655 $Y=1.15
+ $X2=3.8 $Y2=1.15
r102 20 33 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.715 $Y=1.235
+ $X2=3.715 $Y2=1.15
r103 20 31 65.8931 $w=1.68e-07 $l=1.01e-06 $layer=LI1_cond $X=3.715 $Y=1.235
+ $X2=3.715 $Y2=2.245
r104 19 33 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.715 $Y=1.065
+ $X2=3.715 $Y2=1.15
r105 18 19 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=3.715 $Y=0.925
+ $X2=3.715 $Y2=1.065
r106 14 18 7.21222 $w=2.6e-07 $l=1.67183e-07 $layer=LI1_cond $X=3.63 $Y=0.795
+ $X2=3.715 $Y2=0.925
r107 14 16 6.20546 $w=2.58e-07 $l=1.4e-07 $layer=LI1_cond $X=3.63 $Y=0.795
+ $X2=3.49 $Y2=0.795
r108 11 36 19.4347 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.125 $Y=1.185
+ $X2=5.125 $Y2=1.35
r109 11 13 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=5.125 $Y=1.185
+ $X2=5.125 $Y2=0.655
r110 7 35 19.4347 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.055 $Y=1.515
+ $X2=5.055 $Y2=1.35
r111 7 9 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=5.055 $Y=1.515
+ $X2=5.055 $Y2=2.465
r112 2 30 300 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_PDIFF $count=2 $X=3.35
+ $Y=2.235 $X2=3.505 $Y2=2.38
r113 1 16 182 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=1 $X=3.35
+ $Y=0.625 $X2=3.49 $Y2=0.8
.ends

.subckt PM_SKY130_FD_SC_LP__DLRTN_1%RESET_B 3 6 8 9 10 11 17 19
r42 17 20 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.575 $Y=1.35
+ $X2=5.575 $Y2=1.515
r43 17 19 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.575 $Y=1.35
+ $X2=5.575 $Y2=1.185
r44 10 11 13.5366 $w=3.13e-07 $l=3.7e-07 $layer=LI1_cond $X=5.582 $Y=1.665
+ $X2=5.582 $Y2=2.035
r45 9 10 13.5366 $w=3.13e-07 $l=3.7e-07 $layer=LI1_cond $X=5.582 $Y=1.295
+ $X2=5.582 $Y2=1.665
r46 9 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.575
+ $Y=1.35 $X2=5.575 $Y2=1.35
r47 8 9 13.5366 $w=3.13e-07 $l=3.7e-07 $layer=LI1_cond $X=5.582 $Y=0.925
+ $X2=5.582 $Y2=1.295
r48 6 20 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=5.485 $Y=2.465
+ $X2=5.485 $Y2=1.515
r49 3 19 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=5.485 $Y=0.655
+ $X2=5.485 $Y2=1.185
.ends

.subckt PM_SKY130_FD_SC_LP__DLRTN_1%VPWR 1 2 3 4 17 21 23 26 29 34 35 36 38 46
+ 59 60 63 66 69
r84 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r85 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r86 63 64 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r87 59 60 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r88 57 60 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=6.48 $Y2=3.33
r89 57 70 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=4.56 $Y2=3.33
r90 56 57 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r91 54 69 12.7913 $w=1.7e-07 $l=3.1e-07 $layer=LI1_cond $X=4.915 $Y=3.33
+ $X2=4.605 $Y2=3.33
r92 54 56 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=4.915 $Y=3.33
+ $X2=5.52 $Y2=3.33
r93 53 70 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r94 52 53 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r95 50 67 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.64 $Y2=3.33
r96 49 52 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=3.12 $Y=3.33 $X2=4.08
+ $Y2=3.33
r97 49 50 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r98 47 66 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.83 $Y=3.33
+ $X2=2.665 $Y2=3.33
r99 47 49 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=2.83 $Y=3.33
+ $X2=3.12 $Y2=3.33
r100 46 69 12.7913 $w=1.7e-07 $l=3.1e-07 $layer=LI1_cond $X=4.295 $Y=3.33
+ $X2=4.605 $Y2=3.33
r101 46 52 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=4.295 $Y=3.33
+ $X2=4.08 $Y2=3.33
r102 45 67 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r103 44 45 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r104 42 45 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r105 42 64 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r106 41 44 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=3.33 $X2=2.16
+ $Y2=3.33
r107 41 42 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r108 39 63 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=0.895 $Y=3.33
+ $X2=0.79 $Y2=3.33
r109 39 41 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.895 $Y=3.33
+ $X2=1.2 $Y2=3.33
r110 38 66 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.5 $Y=3.33
+ $X2=2.665 $Y2=3.33
r111 38 44 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=2.5 $Y=3.33
+ $X2=2.16 $Y2=3.33
r112 36 53 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=3.36 $Y=3.33
+ $X2=4.08 $Y2=3.33
r113 36 50 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.36 $Y=3.33
+ $X2=3.12 $Y2=3.33
r114 34 56 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=5.575 $Y=3.33
+ $X2=5.52 $Y2=3.33
r115 34 35 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.575 $Y=3.33
+ $X2=5.74 $Y2=3.33
r116 33 59 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=5.905 $Y=3.33
+ $X2=6.48 $Y2=3.33
r117 33 35 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.905 $Y=3.33
+ $X2=5.74 $Y2=3.33
r118 27 35 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.74 $Y=3.245
+ $X2=5.74 $Y2=3.33
r119 27 29 16.5882 $w=3.28e-07 $l=4.75e-07 $layer=LI1_cond $X=5.74 $Y=3.245
+ $X2=5.74 $Y2=2.77
r120 24 69 2.59604 $w=6.2e-07 $l=8.5e-08 $layer=LI1_cond $X=4.605 $Y=3.245
+ $X2=4.605 $Y2=3.33
r121 24 26 12.2502 $w=6.18e-07 $l=6.35e-07 $layer=LI1_cond $X=4.605 $Y=3.245
+ $X2=4.605 $Y2=2.61
r122 23 32 8.82699 $w=6.2e-07 $l=4.99074e-07 $layer=LI1_cond $X=4.605 $Y=2.595
+ $X2=4.815 $Y2=2.19
r123 23 26 0.289374 $w=6.18e-07 $l=1.5e-08 $layer=LI1_cond $X=4.605 $Y=2.595
+ $X2=4.605 $Y2=2.61
r124 19 66 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.665 $Y=3.245
+ $X2=2.665 $Y2=3.33
r125 19 21 17.6359 $w=3.28e-07 $l=5.05e-07 $layer=LI1_cond $X=2.665 $Y=3.245
+ $X2=2.665 $Y2=2.74
r126 15 63 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=0.79 $Y=3.245
+ $X2=0.79 $Y2=3.33
r127 15 17 29.8398 $w=2.08e-07 $l=5.65e-07 $layer=LI1_cond $X=0.79 $Y=3.245
+ $X2=0.79 $Y2=2.68
r128 4 29 600 $w=1.7e-07 $l=1.02104e-06 $layer=licon1_PDIFF $count=1 $X=5.56
+ $Y=1.835 $X2=5.74 $Y2=2.77
r129 3 32 300 $w=1.7e-07 $l=5.87069e-07 $layer=licon1_PDIFF $count=2 $X=4.25
+ $Y=2.235 $X2=4.815 $Y2=2.19
r130 3 26 300 $w=1.7e-07 $l=7.28766e-07 $layer=licon1_PDIFF $count=2 $X=4.25
+ $Y=2.235 $X2=4.815 $Y2=2.61
r131 2 21 600 $w=1.7e-07 $l=5.88154e-07 $layer=licon1_PDIFF $count=1 $X=2.485
+ $Y=2.235 $X2=2.665 $Y2=2.74
r132 1 17 600 $w=1.7e-07 $l=4.2758e-07 $layer=licon1_PDIFF $count=1 $X=0.65
+ $Y=2.325 $X2=0.81 $Y2=2.68
.ends

.subckt PM_SKY130_FD_SC_LP__DLRTN_1%Q 1 2 10 13 14 15 16 17 18 27
r28 17 18 16.0907 $w=2.63e-07 $l=3.7e-07 $layer=LI1_cond $X=6.502 $Y=2.035
+ $X2=6.502 $Y2=2.405
r29 16 17 16.0907 $w=2.63e-07 $l=3.7e-07 $layer=LI1_cond $X=6.502 $Y=1.665
+ $X2=6.502 $Y2=2.035
r30 15 16 16.0907 $w=2.63e-07 $l=3.7e-07 $layer=LI1_cond $X=6.502 $Y=1.295
+ $X2=6.502 $Y2=1.665
r31 15 42 8.69768 $w=2.63e-07 $l=2e-07 $layer=LI1_cond $X=6.502 $Y=1.295
+ $X2=6.502 $Y2=1.095
r32 14 42 6.89526 $w=5.43e-07 $l=1.7e-07 $layer=LI1_cond $X=6.362 $Y=0.925
+ $X2=6.362 $Y2=1.095
r33 14 25 2.23853 $w=5.43e-07 $l=1.02e-07 $layer=LI1_cond $X=6.362 $Y=0.925
+ $X2=6.362 $Y2=0.823
r34 13 25 5.88163 $w=5.43e-07 $l=2.68e-07 $layer=LI1_cond $X=6.362 $Y=0.555
+ $X2=6.362 $Y2=0.823
r35 13 27 2.96276 $w=5.43e-07 $l=1.35e-07 $layer=LI1_cond $X=6.362 $Y=0.555
+ $X2=6.362 $Y2=0.42
r36 11 18 10.2198 $w=2.63e-07 $l=2.35e-07 $layer=LI1_cond $X=6.502 $Y=2.64
+ $X2=6.502 $Y2=2.405
r37 10 11 2.04284 $w=2.65e-07 $l=1.65e-07 $layer=LI1_cond $X=6.502 $Y=2.805
+ $X2=6.502 $Y2=2.64
r38 8 10 9.1497 $w=3.28e-07 $l=2.62e-07 $layer=LI1_cond $X=6.24 $Y=2.805
+ $X2=6.502 $Y2=2.805
r39 2 8 600 $w=1.7e-07 $l=1.03764e-06 $layer=licon1_PDIFF $count=1 $X=6.1
+ $Y=1.835 $X2=6.24 $Y2=2.805
r40 1 27 91 $w=1.7e-07 $l=2.52636e-07 $layer=licon1_NDIFF $count=2 $X=6.1
+ $Y=0.235 $X2=6.26 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__DLRTN_1%VGND 1 2 3 4 15 19 23 27 30 31 33 34 35 37
+ 42 61 62 65 68
c86 62 0 1.22634e-19 $X=6.48 $Y=0
c87 42 0 9.37026e-20 $X=2.425 $Y=0
r88 68 69 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r89 65 66 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r90 61 62 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r91 59 62 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=6.48
+ $Y2=0
r92 58 59 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r93 56 59 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.52
+ $Y2=0
r94 55 58 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=4.56 $Y=0 $X2=5.52
+ $Y2=0
r95 55 56 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r96 53 56 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=4.56
+ $Y2=0
r97 52 53 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r98 50 69 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.64
+ $Y2=0
r99 49 52 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=3.12 $Y=0 $X2=4.08
+ $Y2=0
r100 49 50 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r101 47 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.755 $Y=0 $X2=2.59
+ $Y2=0
r102 47 49 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=2.755 $Y=0
+ $X2=3.12 $Y2=0
r103 46 69 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r104 46 66 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.2
+ $Y2=0
r105 45 46 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r106 43 65 6.36606 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=1.205 $Y=0 $X2=1.095
+ $Y2=0
r107 43 45 62.3048 $w=1.68e-07 $l=9.55e-07 $layer=LI1_cond $X=1.205 $Y=0
+ $X2=2.16 $Y2=0
r108 42 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.425 $Y=0 $X2=2.59
+ $Y2=0
r109 42 45 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=2.425 $Y=0
+ $X2=2.16 $Y2=0
r110 40 66 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r111 39 40 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r112 37 65 6.36606 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=0.985 $Y=0 $X2=1.095
+ $Y2=0
r113 37 39 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.985 $Y=0
+ $X2=0.72 $Y2=0
r114 35 53 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=3.36 $Y=0 $X2=4.08
+ $Y2=0
r115 35 50 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.36 $Y=0
+ $X2=3.12 $Y2=0
r116 33 58 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=5.59 $Y=0 $X2=5.52
+ $Y2=0
r117 33 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.59 $Y=0 $X2=5.755
+ $Y2=0
r118 32 61 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=5.92 $Y=0 $X2=6.48
+ $Y2=0
r119 32 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.92 $Y=0 $X2=5.755
+ $Y2=0
r120 30 52 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=4.225 $Y=0
+ $X2=4.08 $Y2=0
r121 30 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.225 $Y=0 $X2=4.39
+ $Y2=0
r122 29 55 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=4.555 $Y=0 $X2=4.56
+ $Y2=0
r123 29 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.555 $Y=0 $X2=4.39
+ $Y2=0
r124 25 34 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.755 $Y=0.085
+ $X2=5.755 $Y2=0
r125 25 27 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=5.755 $Y=0.085
+ $X2=5.755 $Y2=0.535
r126 21 31 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.39 $Y=0.085
+ $X2=4.39 $Y2=0
r127 21 23 24.4458 $w=3.28e-07 $l=7e-07 $layer=LI1_cond $X=4.39 $Y=0.085
+ $X2=4.39 $Y2=0.785
r128 17 68 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.59 $Y=0.085
+ $X2=2.59 $Y2=0
r129 17 19 24.9696 $w=3.28e-07 $l=7.15e-07 $layer=LI1_cond $X=2.59 $Y=0.085
+ $X2=2.59 $Y2=0.8
r130 13 65 0.432806 $w=2.2e-07 $l=8.5e-08 $layer=LI1_cond $X=1.095 $Y=0.085
+ $X2=1.095 $Y2=0
r131 13 15 18.5962 $w=2.18e-07 $l=3.55e-07 $layer=LI1_cond $X=1.095 $Y=0.085
+ $X2=1.095 $Y2=0.44
r132 4 27 182 $w=1.7e-07 $l=3.85357e-07 $layer=licon1_NDIFF $count=1 $X=5.56
+ $Y=0.235 $X2=5.755 $Y2=0.535
r133 3 23 182 $w=1.7e-07 $l=2.19089e-07 $layer=licon1_NDIFF $count=1 $X=4.25
+ $Y=0.625 $X2=4.39 $Y2=0.785
r134 2 19 182 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=1 $X=2.45
+ $Y=0.625 $X2=2.59 $Y2=0.8
r135 1 15 182 $w=1.7e-07 $l=5.12348e-07 $layer=licon1_NDIFF $count=1 $X=0.65
+ $Y=0.235 $X2=1.07 $Y2=0.44
.ends

