# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__a2bb2o_0
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__a2bb2o_0 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.840000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.530000 0.780000 0.935000 1.760000 ;
    END
  END A1_N
  PIN A2_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.105000 1.145000 1.655000 1.750000 ;
    END
  END A2_N
  PIN B1
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.420000 0.400000 3.755000 2.195000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.760000 0.780000 3.250000 2.195000 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  0.293500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.280000 0.595000 0.610000 ;
        RECT 0.085000 0.610000 0.335000 2.430000 ;
        RECT 0.085000 2.430000 0.445000 3.075000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.840000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.840000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.840000 0.085000 ;
      RECT 0.000000  3.245000 3.840000 3.415000 ;
      RECT 0.505000  1.930000 1.310000 2.260000 ;
      RECT 0.615000  2.430000 0.970000 3.245000 ;
      RECT 0.765000  0.085000 1.025000 0.610000 ;
      RECT 1.140000  2.260000 1.310000 2.880000 ;
      RECT 1.140000  2.880000 2.420000 3.050000 ;
      RECT 1.195000  0.280000 1.465000 0.780000 ;
      RECT 1.195000  0.780000 2.005000 0.975000 ;
      RECT 1.480000  2.430000 2.005000 2.710000 ;
      RECT 1.660000  0.085000 1.990000 0.610000 ;
      RECT 1.835000  0.975000 2.005000 1.235000 ;
      RECT 1.835000  1.235000 2.155000 1.905000 ;
      RECT 1.835000  1.905000 2.005000 2.430000 ;
      RECT 2.160000  0.280000 2.495000 0.610000 ;
      RECT 2.185000  2.075000 2.495000 2.245000 ;
      RECT 2.185000  2.245000 2.420000 2.880000 ;
      RECT 2.325000  0.610000 2.495000 2.075000 ;
      RECT 2.590000  2.415000 3.745000 2.585000 ;
      RECT 2.590000  2.585000 2.825000 3.050000 ;
      RECT 2.980000  0.085000 3.250000 0.610000 ;
      RECT 3.020000  2.755000 3.285000 3.245000 ;
      RECT 3.455000  2.585000 3.745000 3.050000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
  END
END sky130_fd_sc_lp__a2bb2o_0
