* File: sky130_fd_sc_lp__a311oi_2.pex.spice
* Created: Fri Aug 28 09:58:26 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A311OI_2%A3 3 7 11 15 19 22 29 34
r45 26 34 8.46614 $w=3.33e-07 $l=1.65e-07 $layer=LI1_cond $X=0.385 $Y=1.582
+ $X2=0.55 $Y2=1.582
r46 25 27 30.8423 $w=3.36e-07 $l=2.15e-07 $layer=POLY_cond $X=0.385 $Y=1.505
+ $X2=0.6 $Y2=1.505
r47 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.385
+ $Y=1.51 $X2=0.385 $Y2=1.51
r48 22 26 4.98819 $w=3.33e-07 $l=1.45e-07 $layer=LI1_cond $X=0.24 $Y=1.582
+ $X2=0.385 $Y2=1.582
r49 20 29 12.9107 $w=3.36e-07 $l=9e-08 $layer=POLY_cond $X=0.94 $Y=1.505
+ $X2=1.03 $Y2=1.505
r50 20 27 48.7738 $w=3.36e-07 $l=3.4e-07 $layer=POLY_cond $X=0.94 $Y=1.505
+ $X2=0.6 $Y2=1.505
r51 19 34 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=0.94 $Y=1.5 $X2=0.55
+ $Y2=1.5
r52 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.94
+ $Y=1.5 $X2=0.94 $Y2=1.5
r53 13 29 21.6522 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=1.03 $Y=1.675
+ $X2=1.03 $Y2=1.505
r54 13 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.03 $Y=1.675
+ $X2=1.03 $Y2=2.465
r55 9 29 21.6522 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=1.03 $Y=1.335
+ $X2=1.03 $Y2=1.505
r56 9 11 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=1.03 $Y=1.335
+ $X2=1.03 $Y2=0.765
r57 5 27 21.6522 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=0.6 $Y=1.675 $X2=0.6
+ $Y2=1.505
r58 5 7 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=0.6 $Y=1.675 $X2=0.6
+ $Y2=2.465
r59 1 27 21.6522 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=0.6 $Y=1.335 $X2=0.6
+ $Y2=1.505
r60 1 3 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=0.6 $Y=1.335 $X2=0.6
+ $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_LP__A311OI_2%A2 3 7 11 15 22 23 28 32 37
c62 32 0 4.63826e-20 $X=2.275 $Y=1.582
r63 31 37 8.46614 $w=3.33e-07 $l=1.65e-07 $layer=LI1_cond $X=2.105 $Y=1.582
+ $X2=1.94 $Y2=1.582
r64 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.105
+ $Y=1.51 $X2=2.105 $Y2=1.51
r65 28 30 30.8423 $w=3.36e-07 $l=2.15e-07 $layer=POLY_cond $X=1.89 $Y=1.505
+ $X2=2.105 $Y2=1.505
r66 23 32 12.5565 $w=3.33e-07 $l=3.65e-07 $layer=LI1_cond $X=2.64 $Y=1.582
+ $X2=2.275 $Y2=1.582
r67 22 32 3.95615 $w=3.33e-07 $l=1.15e-07 $layer=LI1_cond $X=2.16 $Y=1.582
+ $X2=2.275 $Y2=1.582
r68 22 31 1.89207 $w=3.33e-07 $l=5.5e-08 $layer=LI1_cond $X=2.16 $Y=1.582
+ $X2=2.105 $Y2=1.582
r69 20 28 48.7738 $w=3.36e-07 $l=3.4e-07 $layer=POLY_cond $X=1.55 $Y=1.505
+ $X2=1.89 $Y2=1.505
r70 20 26 12.9107 $w=3.36e-07 $l=9e-08 $layer=POLY_cond $X=1.55 $Y=1.505
+ $X2=1.46 $Y2=1.505
r71 19 37 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=1.55 $Y=1.5 $X2=1.94
+ $Y2=1.5
r72 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.55
+ $Y=1.5 $X2=1.55 $Y2=1.5
r73 13 28 21.6522 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=1.89 $Y=1.675
+ $X2=1.89 $Y2=1.505
r74 13 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.89 $Y=1.675
+ $X2=1.89 $Y2=2.465
r75 9 28 21.6522 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=1.89 $Y=1.335
+ $X2=1.89 $Y2=1.505
r76 9 11 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=1.89 $Y=1.335
+ $X2=1.89 $Y2=0.765
r77 5 26 21.6522 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=1.46 $Y=1.675
+ $X2=1.46 $Y2=1.505
r78 5 7 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.46 $Y=1.675 $X2=1.46
+ $Y2=2.465
r79 1 26 21.6522 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=1.46 $Y=1.335
+ $X2=1.46 $Y2=1.505
r80 1 3 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=1.46 $Y=1.335 $X2=1.46
+ $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_LP__A311OI_2%A1 3 5 6 9 13 17 19 24 25
c67 24 0 1.86389e-19 $X=3.455 $Y=1.51
r68 24 26 14.6061 $w=2.97e-07 $l=9e-08 $layer=POLY_cond $X=3.455 $Y=1.51
+ $X2=3.545 $Y2=1.51
r69 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.455
+ $Y=1.51 $X2=3.455 $Y2=1.51
r70 22 24 55.1785 $w=2.97e-07 $l=3.4e-07 $layer=POLY_cond $X=3.115 $Y=1.51
+ $X2=3.455 $Y2=1.51
r71 19 25 4.52224 $w=3.93e-07 $l=1.55e-07 $layer=LI1_cond $X=3.487 $Y=1.665
+ $X2=3.487 $Y2=1.51
r72 15 26 18.7323 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.545 $Y=1.345
+ $X2=3.545 $Y2=1.51
r73 15 17 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=3.545 $Y=1.345
+ $X2=3.545 $Y2=0.745
r74 11 22 18.7323 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.115 $Y=1.345
+ $X2=3.115 $Y2=1.51
r75 11 13 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=3.115 $Y=1.345
+ $X2=3.115 $Y2=0.745
r76 7 22 21.0976 $w=2.97e-07 $l=2.20624e-07 $layer=POLY_cond $X=2.985 $Y=1.675
+ $X2=3.115 $Y2=1.51
r77 7 9 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.985 $Y=1.675
+ $X2=2.985 $Y2=2.465
r78 5 7 23.9601 $w=2.97e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.91 $Y=1.6
+ $X2=2.985 $Y2=1.675
r79 5 6 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.91 $Y=1.6 $X2=2.63
+ $Y2=1.6
r80 1 6 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.555 $Y=1.675
+ $X2=2.63 $Y2=1.6
r81 1 3 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.555 $Y=1.675
+ $X2=2.555 $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__A311OI_2%B1 3 7 11 15 17 23 24
c43 23 0 1.30901e-19 $X=4.065 $Y=1.51
c44 7 0 6.22842e-20 $X=3.975 $Y=2.465
c45 3 0 1.79852e-19 $X=3.975 $Y=0.745
r46 22 24 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=4.065 $Y=1.51
+ $X2=4.405 $Y2=1.51
r47 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.065
+ $Y=1.51 $X2=4.065 $Y2=1.51
r48 19 22 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=3.975 $Y=1.51
+ $X2=4.065 $Y2=1.51
r49 17 23 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=4.065 $Y=1.665
+ $X2=4.065 $Y2=1.51
r50 13 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.405 $Y=1.675
+ $X2=4.405 $Y2=1.51
r51 13 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=4.405 $Y=1.675
+ $X2=4.405 $Y2=2.465
r52 9 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.405 $Y=1.345
+ $X2=4.405 $Y2=1.51
r53 9 11 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=4.405 $Y=1.345 $X2=4.405
+ $Y2=0.745
r54 5 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.975 $Y=1.675
+ $X2=3.975 $Y2=1.51
r55 5 7 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.975 $Y=1.675
+ $X2=3.975 $Y2=2.465
r56 1 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.975 $Y=1.345
+ $X2=3.975 $Y2=1.51
r57 1 3 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=3.975 $Y=1.345 $X2=3.975
+ $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_LP__A311OI_2%C1 3 7 11 15 17 18 19 28
c41 28 0 1.30901e-19 $X=5.265 $Y=1.51
c42 19 0 6.22842e-20 $X=5.52 $Y=1.665
r43 26 28 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=5.175 $Y=1.51
+ $X2=5.265 $Y2=1.51
r44 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.175
+ $Y=1.51 $X2=5.175 $Y2=1.51
r45 23 26 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=4.835 $Y=1.51
+ $X2=5.175 $Y2=1.51
r46 19 27 12.2336 $w=3.23e-07 $l=3.45e-07 $layer=LI1_cond $X=5.52 $Y=1.587
+ $X2=5.175 $Y2=1.587
r47 18 27 4.78707 $w=3.23e-07 $l=1.35e-07 $layer=LI1_cond $X=5.04 $Y=1.587
+ $X2=5.175 $Y2=1.587
r48 17 18 17.0207 $w=3.23e-07 $l=4.8e-07 $layer=LI1_cond $X=4.56 $Y=1.587
+ $X2=5.04 $Y2=1.587
r49 13 28 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.265 $Y=1.675
+ $X2=5.265 $Y2=1.51
r50 13 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=5.265 $Y=1.675
+ $X2=5.265 $Y2=2.465
r51 9 28 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.265 $Y=1.345
+ $X2=5.265 $Y2=1.51
r52 9 11 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=5.265 $Y=1.345 $X2=5.265
+ $Y2=0.745
r53 5 23 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.835 $Y=1.675
+ $X2=4.835 $Y2=1.51
r54 5 7 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=4.835 $Y=1.675
+ $X2=4.835 $Y2=2.465
r55 1 23 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.835 $Y=1.345
+ $X2=4.835 $Y2=1.51
r56 1 3 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=4.835 $Y=1.345 $X2=4.835
+ $Y2=0.745
.ends

.subckt PM_SKY130_FD_SC_LP__A311OI_2%VPWR 1 2 3 4 13 15 21 27 31 33 35 40 45 55
+ 56 62 65 68
r80 68 69 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r81 65 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r82 62 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r83 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r84 55 56 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r85 53 56 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=5.52 $Y2=3.33
r86 53 69 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=3.12 $Y2=3.33
r87 52 55 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=3.6 $Y=3.33
+ $X2=5.52 $Y2=3.33
r88 52 53 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r89 50 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.365 $Y=3.33
+ $X2=3.2 $Y2=3.33
r90 50 52 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=3.365 $Y=3.33
+ $X2=3.6 $Y2=3.33
r91 49 66 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r92 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r93 46 65 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.39 $Y=3.33
+ $X2=2.225 $Y2=3.33
r94 46 48 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=2.39 $Y=3.33
+ $X2=2.64 $Y2=3.33
r95 45 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.035 $Y=3.33
+ $X2=3.2 $Y2=3.33
r96 45 48 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=3.035 $Y=3.33
+ $X2=2.64 $Y2=3.33
r97 44 66 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r98 44 63 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r99 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r100 41 62 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.41 $Y=3.33
+ $X2=1.245 $Y2=3.33
r101 41 43 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=1.41 $Y=3.33
+ $X2=1.68 $Y2=3.33
r102 40 65 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.06 $Y=3.33
+ $X2=2.225 $Y2=3.33
r103 40 43 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=2.06 $Y=3.33
+ $X2=1.68 $Y2=3.33
r104 39 63 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r105 39 60 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r106 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r107 36 59 4.54404 $w=1.7e-07 $l=2.75e-07 $layer=LI1_cond $X=0.55 $Y=3.33
+ $X2=0.275 $Y2=3.33
r108 36 38 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=0.55 $Y=3.33
+ $X2=0.72 $Y2=3.33
r109 35 62 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.08 $Y=3.33
+ $X2=1.245 $Y2=3.33
r110 35 38 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=1.08 $Y=3.33
+ $X2=0.72 $Y2=3.33
r111 33 69 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.88 $Y=3.33
+ $X2=3.12 $Y2=3.33
r112 33 49 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.88 $Y=3.33
+ $X2=2.64 $Y2=3.33
r113 29 68 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.2 $Y=3.245 $X2=3.2
+ $Y2=3.33
r114 29 31 16.9374 $w=3.28e-07 $l=4.85e-07 $layer=LI1_cond $X=3.2 $Y=3.245
+ $X2=3.2 $Y2=2.76
r115 25 65 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.225 $Y=3.245
+ $X2=2.225 $Y2=3.33
r116 25 27 16.9374 $w=3.28e-07 $l=4.85e-07 $layer=LI1_cond $X=2.225 $Y=3.245
+ $X2=2.225 $Y2=2.76
r117 21 24 26.8903 $w=3.28e-07 $l=7.7e-07 $layer=LI1_cond $X=1.245 $Y=2.18
+ $X2=1.245 $Y2=2.95
r118 19 62 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.245 $Y=3.245
+ $X2=1.245 $Y2=3.33
r119 19 24 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.245 $Y=3.245
+ $X2=1.245 $Y2=2.95
r120 15 18 33.0018 $w=3.28e-07 $l=9.45e-07 $layer=LI1_cond $X=0.385 $Y=2.005
+ $X2=0.385 $Y2=2.95
r121 13 59 3.22214 $w=3.3e-07 $l=1.46458e-07 $layer=LI1_cond $X=0.385 $Y=3.245
+ $X2=0.275 $Y2=3.33
r122 13 18 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.385 $Y=3.245
+ $X2=0.385 $Y2=2.95
r123 4 31 600 $w=1.7e-07 $l=9.92535e-07 $layer=licon1_PDIFF $count=1 $X=3.06
+ $Y=1.835 $X2=3.2 $Y2=2.76
r124 3 27 600 $w=1.7e-07 $l=1.04696e-06 $layer=licon1_PDIFF $count=1 $X=1.965
+ $Y=1.835 $X2=2.225 $Y2=2.76
r125 2 24 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=1.105
+ $Y=1.835 $X2=1.245 $Y2=2.95
r126 2 21 400 $w=1.7e-07 $l=4.09054e-07 $layer=licon1_PDIFF $count=1 $X=1.105
+ $Y=1.835 $X2=1.245 $Y2=2.18
r127 1 18 400 $w=1.7e-07 $l=1.17584e-06 $layer=licon1_PDIFF $count=1 $X=0.26
+ $Y=1.835 $X2=0.385 $Y2=2.95
r128 1 15 400 $w=1.7e-07 $l=2.23942e-07 $layer=licon1_PDIFF $count=1 $X=0.26
+ $Y=1.835 $X2=0.385 $Y2=2.005
.ends

.subckt PM_SKY130_FD_SC_LP__A311OI_2%A_135_367# 1 2 3 4 15 19 20 27 31 33 36 38
c53 33 0 1.86389e-19 $X=4.025 $Y=2.375
r54 34 38 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.865 $Y=2.375
+ $X2=2.735 $Y2=2.375
r55 33 42 3.12527 $w=2.93e-07 $l=8e-08 $layer=LI1_cond $X=4.172 $Y=2.375
+ $X2=4.172 $Y2=2.455
r56 33 34 75.6791 $w=1.68e-07 $l=1.16e-06 $layer=LI1_cond $X=4.025 $Y=2.375
+ $X2=2.865 $Y2=2.375
r57 29 38 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=2.735 $Y=2.46
+ $X2=2.735 $Y2=2.375
r58 29 31 19.9461 $w=2.58e-07 $l=4.5e-07 $layer=LI1_cond $X=2.735 $Y=2.46
+ $X2=2.735 $Y2=2.91
r59 28 36 2.36881 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.84 $Y=2.375
+ $X2=1.71 $Y2=2.375
r60 27 38 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.605 $Y=2.375
+ $X2=2.735 $Y2=2.375
r61 27 28 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=2.605 $Y=2.375
+ $X2=1.84 $Y2=2.375
r62 22 36 4.06715 $w=2.25e-07 $l=1.00995e-07 $layer=LI1_cond $X=1.675 $Y=2.29
+ $X2=1.71 $Y2=2.375
r63 22 24 18.0957 $w=1.88e-07 $l=3.1e-07 $layer=LI1_cond $X=1.675 $Y=2.29
+ $X2=1.675 $Y2=1.98
r64 21 24 3.21053 $w=1.88e-07 $l=5.5e-08 $layer=LI1_cond $X=1.675 $Y=1.925
+ $X2=1.675 $Y2=1.98
r65 19 21 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=1.58 $Y=1.84
+ $X2=1.675 $Y2=1.925
r66 19 20 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.58 $Y=1.84 $X2=0.9
+ $Y2=1.84
r67 15 17 57.303 $w=1.78e-07 $l=9.3e-07 $layer=LI1_cond $X=0.81 $Y=1.98 $X2=0.81
+ $Y2=2.91
r68 13 20 6.82373 $w=1.7e-07 $l=1.25499e-07 $layer=LI1_cond $X=0.81 $Y=1.925
+ $X2=0.9 $Y2=1.84
r69 13 15 3.38889 $w=1.78e-07 $l=5.5e-08 $layer=LI1_cond $X=0.81 $Y=1.925
+ $X2=0.81 $Y2=1.98
r70 4 42 600 $w=1.7e-07 $l=6.8644e-07 $layer=licon1_PDIFF $count=1 $X=4.05
+ $Y=1.835 $X2=4.19 $Y2=2.455
r71 3 38 600 $w=1.7e-07 $l=6.0597e-07 $layer=licon1_PDIFF $count=1 $X=2.63
+ $Y=1.835 $X2=2.77 $Y2=2.375
r72 3 31 600 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=2.63
+ $Y=1.835 $X2=2.77 $Y2=2.91
r73 2 36 300 $w=1.7e-07 $l=6.76387e-07 $layer=licon1_PDIFF $count=2 $X=1.535
+ $Y=1.835 $X2=1.675 $Y2=2.445
r74 2 24 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.535
+ $Y=1.835 $X2=1.675 $Y2=1.98
r75 1 17 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=0.675
+ $Y=1.835 $X2=0.815 $Y2=2.91
r76 1 15 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.675
+ $Y=1.835 $X2=0.815 $Y2=1.98
.ends

.subckt PM_SKY130_FD_SC_LP__A311OI_2%A_727_367# 1 2 3 10 16 18 20 22 25
r29 20 27 2.78046 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=5.505 $Y=2.905
+ $X2=5.505 $Y2=2.99
r30 20 22 33.7501 $w=2.78e-07 $l=8.2e-07 $layer=LI1_cond $X=5.505 $Y=2.905
+ $X2=5.505 $Y2=2.085
r31 19 25 5.8691 $w=2.22e-07 $l=1.5424e-07 $layer=LI1_cond $X=4.75 $Y=2.99
+ $X2=4.62 $Y2=2.937
r32 18 27 4.57959 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=5.365 $Y=2.99
+ $X2=5.505 $Y2=2.99
r33 18 19 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=5.365 $Y=2.99
+ $X2=4.75 $Y2=2.99
r34 14 25 0.788168 $w=2.6e-07 $l=1.37e-07 $layer=LI1_cond $X=4.62 $Y=2.8
+ $X2=4.62 $Y2=2.937
r35 14 16 15.292 $w=2.58e-07 $l=3.45e-07 $layer=LI1_cond $X=4.62 $Y=2.8 $X2=4.62
+ $Y2=2.455
r36 10 25 5.8691 $w=2.22e-07 $l=1.3e-07 $layer=LI1_cond $X=4.49 $Y=2.937
+ $X2=4.62 $Y2=2.937
r37 10 12 30.5921 $w=2.73e-07 $l=7.3e-07 $layer=LI1_cond $X=4.49 $Y=2.937
+ $X2=3.76 $Y2=2.937
r38 3 27 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=5.34
+ $Y=1.835 $X2=5.48 $Y2=2.91
r39 3 22 400 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_PDIFF $count=1 $X=5.34
+ $Y=1.835 $X2=5.48 $Y2=2.085
r40 2 25 600 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=4.48
+ $Y=1.835 $X2=4.62 $Y2=2.91
r41 2 16 600 $w=1.7e-07 $l=6.8644e-07 $layer=licon1_PDIFF $count=1 $X=4.48
+ $Y=1.835 $X2=4.62 $Y2=2.455
r42 1 12 600 $w=1.7e-07 $l=1.14079e-06 $layer=licon1_PDIFF $count=1 $X=3.635
+ $Y=1.835 $X2=3.76 $Y2=2.915
.ends

.subckt PM_SKY130_FD_SC_LP__A311OI_2%Y 1 2 3 4 5 18 21 22 26 28 32 34 40 42 43
+ 44 45 47 48 49 50 51 52 59 67
r101 65 67 2.49545 $w=1.98e-07 $l=4.5e-08 $layer=LI1_cond $X=3.075 $Y=2.02
+ $X2=3.12 $Y2=2.02
r102 51 52 26.6182 $w=1.98e-07 $l=4.8e-07 $layer=LI1_cond $X=3.6 $Y=2.02
+ $X2=4.08 $Y2=2.02
r103 50 59 4.50329 $w=2e-07 $l=8.5e-08 $layer=LI1_cond $X=2.99 $Y=2.02 $X2=2.905
+ $Y2=2.02
r104 50 65 4.50329 $w=2e-07 $l=8.5e-08 $layer=LI1_cond $X=2.99 $Y=2.02 $X2=3.075
+ $Y2=2.02
r105 50 51 25.5091 $w=1.98e-07 $l=4.6e-07 $layer=LI1_cond $X=3.14 $Y=2.02
+ $X2=3.6 $Y2=2.02
r106 50 67 1.10909 $w=1.98e-07 $l=2e-08 $layer=LI1_cond $X=3.14 $Y=2.02 $X2=3.12
+ $Y2=2.02
r107 49 59 14.6955 $w=1.98e-07 $l=2.65e-07 $layer=LI1_cond $X=2.64 $Y=2.02
+ $X2=2.905 $Y2=2.02
r108 48 49 26.6182 $w=1.98e-07 $l=4.8e-07 $layer=LI1_cond $X=2.16 $Y=2.02
+ $X2=2.64 $Y2=2.02
r109 45 52 46.5818 $w=1.98e-07 $l=8.4e-07 $layer=LI1_cond $X=4.92 $Y=2.02
+ $X2=4.08 $Y2=2.02
r110 45 47 4.06946 $w=2e-07 $l=1.37e-07 $layer=LI1_cond $X=4.92 $Y=2.02
+ $X2=5.057 $Y2=2.02
r111 38 40 25.3126 $w=2.78e-07 $l=6.15e-07 $layer=LI1_cond $X=5.525 $Y=1.085
+ $X2=5.525 $Y2=0.47
r112 35 44 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=4.715 $Y=1.17
+ $X2=4.62 $Y2=1.17
r113 34 38 7.36005 $w=1.7e-07 $l=1.77482e-07 $layer=LI1_cond $X=5.385 $Y=1.17
+ $X2=5.525 $Y2=1.085
r114 34 35 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.385 $Y=1.17
+ $X2=4.715 $Y2=1.17
r115 30 44 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=4.62 $Y=1.085
+ $X2=4.62 $Y2=1.17
r116 30 32 35.8995 $w=1.88e-07 $l=6.15e-07 $layer=LI1_cond $X=4.62 $Y=1.085
+ $X2=4.62 $Y2=0.47
r117 29 43 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=3.855 $Y=1.17
+ $X2=3.76 $Y2=1.17
r118 28 44 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=4.525 $Y=1.17
+ $X2=4.62 $Y2=1.17
r119 28 29 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.525 $Y=1.17
+ $X2=3.855 $Y2=1.17
r120 24 43 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=3.76 $Y=1.085
+ $X2=3.76 $Y2=1.17
r121 24 26 35.8995 $w=1.88e-07 $l=6.15e-07 $layer=LI1_cond $X=3.76 $Y=1.085
+ $X2=3.76 $Y2=0.47
r122 23 42 2.83584 $w=1.7e-07 $l=4.60543e-07 $layer=LI1_cond $X=3.075 $Y=1.17
+ $X2=2.655 $Y2=1.085
r123 22 43 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=3.665 $Y=1.17
+ $X2=3.76 $Y2=1.17
r124 22 23 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=3.665 $Y=1.17
+ $X2=3.075 $Y2=1.17
r125 21 50 1.93381 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=2.99 $Y=1.92 $X2=2.99
+ $Y2=2.02
r126 20 42 3.64284 $w=2.55e-07 $l=4.11309e-07 $layer=LI1_cond $X=2.99 $Y=1.255
+ $X2=2.655 $Y2=1.085
r127 20 21 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=2.99 $Y=1.255
+ $X2=2.99 $Y2=1.92
r128 16 42 3.64284 $w=2.55e-07 $l=1.7e-07 $layer=LI1_cond $X=2.825 $Y=1.085
+ $X2=2.655 $Y2=1.085
r129 16 18 13.7276 $w=3.38e-07 $l=4.05e-07 $layer=LI1_cond $X=2.825 $Y=1.085
+ $X2=2.825 $Y2=0.68
r130 5 47 300 $w=1.7e-07 $l=3.42929e-07 $layer=licon1_PDIFF $count=2 $X=4.91
+ $Y=1.835 $X2=5.05 $Y2=2.115
r131 4 40 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.34
+ $Y=0.325 $X2=5.48 $Y2=0.47
r132 3 32 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.48
+ $Y=0.325 $X2=4.62 $Y2=0.47
r133 2 26 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.62
+ $Y=0.325 $X2=3.76 $Y2=0.47
r134 1 18 91 $w=1.7e-07 $l=4.255e-07 $layer=licon1_NDIFF $count=2 $X=2.675
+ $Y=0.325 $X2=2.83 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_LP__A311OI_2%A_48_69# 1 2 3 12 14 15 18 20 24 26
r42 22 24 13.3887 $w=3.38e-07 $l=3.95e-07 $layer=LI1_cond $X=2.18 $Y=1.075
+ $X2=2.18 $Y2=0.68
r43 21 26 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.34 $Y=1.16
+ $X2=1.245 $Y2=1.16
r44 20 22 7.85115 $w=1.7e-07 $l=2.08207e-07 $layer=LI1_cond $X=2.01 $Y=1.16
+ $X2=2.18 $Y2=1.075
r45 20 21 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.01 $Y=1.16
+ $X2=1.34 $Y2=1.16
r46 16 26 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.245 $Y=1.075
+ $X2=1.245 $Y2=1.16
r47 16 18 34.1483 $w=1.88e-07 $l=5.85e-07 $layer=LI1_cond $X=1.245 $Y=1.075
+ $X2=1.245 $Y2=0.49
r48 14 26 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.15 $Y=1.16
+ $X2=1.245 $Y2=1.16
r49 14 15 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.15 $Y=1.16
+ $X2=0.48 $Y2=1.16
r50 10 15 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=0.35 $Y=1.075
+ $X2=0.48 $Y2=1.16
r51 10 12 25.93 $w=2.58e-07 $l=5.85e-07 $layer=LI1_cond $X=0.35 $Y=1.075
+ $X2=0.35 $Y2=0.49
r52 3 24 91 $w=1.7e-07 $l=4.27288e-07 $layer=licon1_NDIFF $count=2 $X=1.965
+ $Y=0.345 $X2=2.175 $Y2=0.68
r53 2 18 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.105
+ $Y=0.345 $X2=1.245 $Y2=0.49
r54 1 12 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.24
+ $Y=0.345 $X2=0.385 $Y2=0.49
.ends

.subckt PM_SKY130_FD_SC_LP__A311OI_2%VGND 1 2 3 14 18 22 24 26 31 38 39 42 45 48
r68 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r69 45 46 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=4.08 $Y=0
+ $X2=4.08 $Y2=0
r70 42 43 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r71 39 49 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=5.04
+ $Y2=0
r72 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r73 36 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.215 $Y=0 $X2=5.05
+ $Y2=0
r74 36 38 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=5.215 $Y=0 $X2=5.52
+ $Y2=0
r75 35 49 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.04
+ $Y2=0
r76 35 46 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=4.08
+ $Y2=0
r77 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r78 32 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.355 $Y=0 $X2=4.19
+ $Y2=0
r79 32 34 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=4.355 $Y=0 $X2=4.56
+ $Y2=0
r80 31 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.885 $Y=0 $X2=5.05
+ $Y2=0
r81 31 34 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=4.885 $Y=0 $X2=4.56
+ $Y2=0
r82 30 43 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r83 29 30 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=1.2 $Y=0
+ $X2=1.2 $Y2=0
r84 27 42 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.98 $Y=0 $X2=0.815
+ $Y2=0
r85 27 29 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=0.98 $Y=0 $X2=1.2
+ $Y2=0
r86 26 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.025 $Y=0 $X2=4.19
+ $Y2=0
r87 26 29 184.305 $w=1.68e-07 $l=2.825e-06 $layer=LI1_cond $X=4.025 $Y=0 $X2=1.2
+ $Y2=0
r88 24 46 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=2.88 $Y=0 $X2=4.08
+ $Y2=0
r89 24 30 0.468274 $w=4.9e-07 $l=1.68e-06 $layer=MET1_cond $X=2.88 $Y=0 $X2=1.2
+ $Y2=0
r90 20 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.05 $Y=0.085
+ $X2=5.05 $Y2=0
r91 20 22 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=5.05 $Y=0.085
+ $X2=5.05 $Y2=0.45
r92 16 45 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.19 $Y=0.085
+ $X2=4.19 $Y2=0
r93 16 18 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=4.19 $Y=0.085
+ $X2=4.19 $Y2=0.45
r94 12 42 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.815 $Y=0.085
+ $X2=0.815 $Y2=0
r95 12 14 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=0.815 $Y=0.085
+ $X2=0.815 $Y2=0.47
r96 3 22 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=4.91
+ $Y=0.325 $X2=5.05 $Y2=0.45
r97 2 18 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=4.05
+ $Y=0.325 $X2=4.19 $Y2=0.45
r98 1 14 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=0.675
+ $Y=0.345 $X2=0.815 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_LP__A311OI_2%A_307_69# 1 2 9 11 12 15
c31 11 0 1.79852e-19 $X=3.165 $Y=0.34
r32 13 15 0.873063 $w=3.28e-07 $l=2.5e-08 $layer=LI1_cond $X=3.33 $Y=0.425
+ $X2=3.33 $Y2=0.45
r33 11 13 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.165 $Y=0.34
+ $X2=3.33 $Y2=0.425
r34 11 12 86.4438 $w=1.68e-07 $l=1.325e-06 $layer=LI1_cond $X=3.165 $Y=0.34
+ $X2=1.84 $Y2=0.34
r35 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.675 $Y=0.425
+ $X2=1.84 $Y2=0.34
r36 7 9 1.57151 $w=3.28e-07 $l=4.5e-08 $layer=LI1_cond $X=1.675 $Y=0.425
+ $X2=1.675 $Y2=0.47
r37 2 15 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=3.19
+ $Y=0.325 $X2=3.33 $Y2=0.45
r38 1 9 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=1.535
+ $Y=0.345 $X2=1.675 $Y2=0.47
.ends

