# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__a41oi_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_lp__a41oi_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.240000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.115000 1.210000 1.900000 1.610000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.970000 1.425000 3.685000 1.830000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.105000 1.375000 4.785000 1.545000 ;
        RECT 4.400000 1.210000 4.730000 1.375000 ;
    END
  END A3
  PIN A4
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.250000 1.425000 6.155000 1.750000 ;
    END
  END A4
  PIN B1
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.210000 0.805000 1.750000 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  0.823200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.670000 0.255000 0.860000 0.870000 ;
        RECT 0.670000 0.870000 2.330000 1.040000 ;
        RECT 0.905000 1.890000 2.800000 1.950000 ;
        RECT 0.905000 1.950000 1.235000 2.725000 ;
        RECT 0.975000 1.780000 2.800000 1.890000 ;
        RECT 2.000000 0.595000 2.330000 0.870000 ;
        RECT 2.070000 1.040000 2.330000 1.425000 ;
        RECT 2.070000 1.425000 2.800000 1.780000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 6.240000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 6.240000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.240000 0.085000 ;
      RECT 0.000000  3.245000 6.240000 3.415000 ;
      RECT 0.170000  0.085000 0.500000 1.040000 ;
      RECT 0.475000  1.920000 0.735000 2.895000 ;
      RECT 0.475000  2.895000 1.665000 3.075000 ;
      RECT 1.030000  0.085000 1.360000 0.700000 ;
      RECT 1.335000  2.885000 1.665000 2.895000 ;
      RECT 1.405000  2.120000 4.130000 2.290000 ;
      RECT 1.405000  2.290000 1.665000 2.885000 ;
      RECT 1.550000  0.255000 2.690000 0.425000 ;
      RECT 1.550000  0.425000 1.830000 0.700000 ;
      RECT 1.845000  2.460000 2.175000 3.245000 ;
      RECT 2.360000  2.290000 4.130000 2.325000 ;
      RECT 2.360000  2.325000 2.690000 3.075000 ;
      RECT 2.500000  0.425000 2.690000 1.085000 ;
      RECT 2.500000  1.085000 3.690000 1.255000 ;
      RECT 2.860000  0.255000 4.730000 0.425000 ;
      RECT 2.860000  0.425000 3.190000 0.915000 ;
      RECT 2.860000  2.505000 3.700000 3.245000 ;
      RECT 3.360000  0.595000 3.690000 1.085000 ;
      RECT 3.855000  1.715000 5.080000 1.885000 ;
      RECT 3.855000  1.885000 4.130000 2.120000 ;
      RECT 3.870000  2.325000 4.130000 3.075000 ;
      RECT 3.900000  0.595000 4.230000 0.870000 ;
      RECT 3.900000  0.870000 5.090000 1.040000 ;
      RECT 3.900000  1.040000 4.230000 1.205000 ;
      RECT 4.315000  2.055000 4.645000 3.245000 ;
      RECT 4.400000  0.425000 4.730000 0.700000 ;
      RECT 4.830000  1.885000 5.080000 1.925000 ;
      RECT 4.830000  1.925000 6.020000 2.095000 ;
      RECT 4.830000  2.095000 5.090000 3.075000 ;
      RECT 4.900000  0.325000 5.090000 0.870000 ;
      RECT 4.910000  1.040000 5.090000 1.085000 ;
      RECT 4.910000  1.085000 6.020000 1.255000 ;
      RECT 5.260000  0.085000 5.590000 0.915000 ;
      RECT 5.260000  2.265000 5.590000 3.245000 ;
      RECT 5.760000  0.325000 6.020000 1.085000 ;
      RECT 5.760000  2.095000 6.020000 3.075000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
  END
END sky130_fd_sc_lp__a41oi_2
END LIBRARY
