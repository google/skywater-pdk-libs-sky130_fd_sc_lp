* NGSPICE file created from sky130_fd_sc_lp__and4b_lp.ext - technology: sky130A

.subckt sky130_fd_sc_lp__and4b_lp A_N B C D VGND VNB VPB VPWR X
M1000 a_276_47# D VGND VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=2.457e+11p ps=2.85e+06u
M1001 a_354_47# C a_276_47# VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1002 a_432_47# B a_354_47# VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1003 a_480_21# A_N a_708_47# VNB nshort w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=8.82e+10p ps=1.26e+06u
M1004 VPWR a_84_21# X VPB phighvt w=1e+06u l=250000u
+  ad=1.14e+12p pd=8.28e+06u as=2.85e+11p ps=2.57e+06u
M1005 a_480_21# A_N VPWR VPB phighvt w=1e+06u l=250000u
+  ad=2.85e+11p pd=2.57e+06u as=0p ps=0u
M1006 a_114_47# a_84_21# X VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=1.197e+11p ps=1.41e+06u
M1007 VPWR a_480_21# a_84_21# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=5.6e+11p ps=5.12e+06u
M1008 a_708_47# A_N VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR C a_84_21# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_84_21# a_480_21# a_432_47# VNB nshort w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=0p ps=0u
M1011 a_84_21# B VPWR VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VGND a_84_21# a_114_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_84_21# D VPWR VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
.ends

