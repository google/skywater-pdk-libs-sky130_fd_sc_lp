* File: sky130_fd_sc_lp__a2111oi_m.pxi.spice
* Created: Fri Aug 28 09:47:11 2020
* 
x_PM_SKY130_FD_SC_LP__A2111OI_M%D1 N_D1_M1009_g N_D1_M1000_g N_D1_c_71_n
+ N_D1_c_76_n D1 D1 D1 D1 D1 N_D1_c_73_n PM_SKY130_FD_SC_LP__A2111OI_M%D1
x_PM_SKY130_FD_SC_LP__A2111OI_M%C1 N_C1_M1007_g N_C1_M1003_g N_C1_c_107_n
+ N_C1_c_108_n C1 C1 C1 N_C1_c_109_n N_C1_c_110_n
+ PM_SKY130_FD_SC_LP__A2111OI_M%C1
x_PM_SKY130_FD_SC_LP__A2111OI_M%B1 N_B1_M1008_g N_B1_M1001_g N_B1_c_146_n B1 B1
+ B1 N_B1_c_148_n PM_SKY130_FD_SC_LP__A2111OI_M%B1
x_PM_SKY130_FD_SC_LP__A2111OI_M%A1 N_A1_c_194_n N_A1_M1004_g N_A1_M1005_g
+ N_A1_c_196_n A1 A1 A1 N_A1_c_193_n PM_SKY130_FD_SC_LP__A2111OI_M%A1
x_PM_SKY130_FD_SC_LP__A2111OI_M%A2 N_A2_M1002_g N_A2_c_239_n N_A2_M1006_g
+ N_A2_c_233_n N_A2_c_234_n N_A2_c_240_n N_A2_c_241_n N_A2_c_235_n N_A2_c_236_n
+ A2 A2 A2 A2 A2 N_A2_c_238_n PM_SKY130_FD_SC_LP__A2111OI_M%A2
x_PM_SKY130_FD_SC_LP__A2111OI_M%Y N_Y_M1009_d N_Y_M1001_d N_Y_M1000_s
+ N_Y_c_270_n N_Y_c_271_n N_Y_c_272_n N_Y_c_273_n N_Y_c_310_p Y N_Y_c_274_n
+ PM_SKY130_FD_SC_LP__A2111OI_M%Y
x_PM_SKY130_FD_SC_LP__A2111OI_M%A_299_533# N_A_299_533#_M1008_d
+ N_A_299_533#_M1006_d N_A_299_533#_c_323_n N_A_299_533#_c_320_n
+ N_A_299_533#_c_321_n N_A_299_533#_c_322_n
+ PM_SKY130_FD_SC_LP__A2111OI_M%A_299_533#
x_PM_SKY130_FD_SC_LP__A2111OI_M%VPWR N_VPWR_M1004_d N_VPWR_c_351_n VPWR
+ N_VPWR_c_352_n N_VPWR_c_353_n N_VPWR_c_350_n N_VPWR_c_355_n
+ PM_SKY130_FD_SC_LP__A2111OI_M%VPWR
x_PM_SKY130_FD_SC_LP__A2111OI_M%VGND N_VGND_M1009_s N_VGND_M1003_d
+ N_VGND_M1002_d N_VGND_c_389_n N_VGND_c_390_n N_VGND_c_391_n N_VGND_c_392_n
+ N_VGND_c_393_n VGND N_VGND_c_394_n N_VGND_c_395_n N_VGND_c_396_n
+ N_VGND_c_397_n N_VGND_c_398_n PM_SKY130_FD_SC_LP__A2111OI_M%VGND
cc_1 VNB N_D1_M1009_g 0.046155f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=0.445
cc_2 VNB N_D1_c_71_n 0.0191305f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.715
cc_3 VNB D1 0.00428674f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_4 VNB N_D1_c_73_n 0.016463f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.375
cc_5 VNB N_C1_M1007_g 0.00439882f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=0.445
cc_6 VNB N_C1_M1003_g 0.0236762f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=2.875
cc_7 VNB N_C1_c_107_n 0.0240788f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.715
cc_8 VNB N_C1_c_108_n 0.0163694f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.88
cc_9 VNB N_C1_c_109_n 0.0165614f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_C1_c_110_n 6.58274e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_B1_M1001_g 0.0452437f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=2.875
cc_12 VNB N_B1_c_146_n 0.0145094f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.88
cc_13 VNB B1 0.00109427f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=2.32
cc_14 VNB N_B1_c_148_n 0.0169766f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.375
cc_15 VNB N_A1_M1005_g 0.0596893f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=2.875
cc_16 VNB A1 0.00865124f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_17 VNB N_A1_c_193_n 0.0175904f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A2_M1002_g 0.0306166f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=0.445
cc_19 VNB N_A2_c_233_n 0.0598032f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A2_c_234_n 0.0132443f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.375
cc_21 VNB N_A2_c_235_n 0.00207687f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_22 VNB N_A2_c_236_n 0.025408f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=2.32
cc_23 VNB A2 0.0280692f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=2.69
cc_24 VNB N_A2_c_238_n 0.0392394f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_Y_c_270_n 0.0376448f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.88
cc_26 VNB N_Y_c_271_n 0.00904162f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_27 VNB N_Y_c_272_n 0.010412f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.95
cc_28 VNB N_Y_c_273_n 0.0191951f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=2.32
cc_29 VNB N_Y_c_274_n 0.00872407f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VPWR_c_350_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_389_n 0.0138712f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.21
cc_32 VNB N_VGND_c_390_n 0.00485511f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.88
cc_33 VNB N_VGND_c_391_n 0.0180839f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_34 VNB N_VGND_c_392_n 0.00295613f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_393_n 0.00495479f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_394_n 0.0313406f $X=-0.19 $Y=-0.245 $X2=0.665 $Y2=1.295
cc_37 VNB N_VGND_c_395_n 0.0180745f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_396_n 0.202095f $X=-0.19 $Y=-0.245 $X2=0.665 $Y2=2.405
cc_39 VNB N_VGND_c_397_n 0.00521838f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_398_n 0.00401177f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VPB N_D1_M1000_g 0.0558486f $X=-0.19 $Y=1.655 $X2=0.7 $Y2=2.875
cc_42 VPB N_D1_c_71_n 0.00404552f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=1.715
cc_43 VPB N_D1_c_76_n 0.0185838f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=1.88
cc_44 VPB D1 0.0158855f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_45 VPB N_C1_M1007_g 0.0571663f $X=-0.19 $Y=1.655 $X2=0.7 $Y2=0.445
cc_46 VPB N_C1_c_110_n 0.0105543f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_47 VPB N_B1_M1008_g 0.0487212f $X=-0.19 $Y=1.655 $X2=0.7 $Y2=0.445
cc_48 VPB N_B1_c_146_n 0.0444461f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=1.88
cc_49 VPB B1 0.00469355f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=2.32
cc_50 VPB N_A1_c_194_n 0.0545444f $X=-0.19 $Y=1.655 $X2=0.7 $Y2=1.21
cc_51 VPB N_A1_M1004_g 0.0302142f $X=-0.19 $Y=1.655 $X2=0.7 $Y2=0.445
cc_52 VPB N_A1_c_196_n 0.0276942f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=1.715
cc_53 VPB A1 0.00114206f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_54 VPB N_A1_c_193_n 0.00277856f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_55 VPB N_A2_c_239_n 0.0213622f $X=-0.19 $Y=1.655 $X2=0.7 $Y2=1.88
cc_56 VPB N_A2_c_240_n 0.0477572f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=1.21
cc_57 VPB N_A2_c_241_n 0.0143124f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=1.715
cc_58 VPB N_A2_c_235_n 0.0577506f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_59 VPB A2 0.0218042f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=2.69
cc_60 VPB N_Y_c_270_n 0.0486282f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=1.88
cc_61 VPB N_A_299_533#_c_320_n 0.0118052f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=1.715
cc_62 VPB N_A_299_533#_c_321_n 0.00459896f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=1.88
cc_63 VPB N_A_299_533#_c_322_n 0.0140462f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_64 VPB N_VPWR_c_351_n 0.00326684f $X=-0.19 $Y=1.655 $X2=0.7 $Y2=2.875
cc_65 VPB N_VPWR_c_352_n 0.0567345f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=1.21
cc_66 VPB N_VPWR_c_353_n 0.0339707f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_67 VPB N_VPWR_c_350_n 0.058117f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_355_n 0.00528984f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=1.375
cc_69 N_D1_c_76_n N_C1_M1007_g 0.0355002f $X=0.61 $Y=1.88 $X2=0 $Y2=0
cc_70 N_D1_M1009_g N_C1_M1003_g 0.0204171f $X=0.7 $Y=0.445 $X2=0 $Y2=0
cc_71 D1 N_C1_c_107_n 0.0171143f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_72 N_D1_c_73_n N_C1_c_107_n 0.0355002f $X=0.61 $Y=1.375 $X2=0 $Y2=0
cc_73 N_D1_c_71_n N_C1_c_108_n 0.0355002f $X=0.61 $Y=1.715 $X2=0 $Y2=0
cc_74 N_D1_M1009_g N_C1_c_109_n 0.0355002f $X=0.7 $Y=0.445 $X2=0 $Y2=0
cc_75 N_D1_M1009_g N_C1_c_110_n 9.42772e-19 $X=0.7 $Y=0.445 $X2=0 $Y2=0
cc_76 D1 N_C1_c_110_n 0.0680254f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_77 N_D1_c_73_n N_C1_c_110_n 0.0010756f $X=0.61 $Y=1.375 $X2=0 $Y2=0
cc_78 D1 N_Y_M1000_s 0.00277331f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_79 N_D1_M1009_g N_Y_c_270_n 0.00732638f $X=0.7 $Y=0.445 $X2=0 $Y2=0
cc_80 N_D1_M1000_g N_Y_c_270_n 0.00897795f $X=0.7 $Y=2.875 $X2=0 $Y2=0
cc_81 D1 N_Y_c_270_n 0.121676f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_82 N_D1_c_73_n N_Y_c_270_n 0.0164112f $X=0.61 $Y=1.375 $X2=0 $Y2=0
cc_83 N_D1_M1009_g N_Y_c_271_n 0.00427926f $X=0.7 $Y=0.445 $X2=0 $Y2=0
cc_84 D1 N_Y_c_271_n 0.00541828f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_85 N_D1_c_73_n N_Y_c_271_n 0.0034593f $X=0.61 $Y=1.375 $X2=0 $Y2=0
cc_86 N_D1_M1009_g N_Y_c_274_n 0.0223781f $X=0.7 $Y=0.445 $X2=0 $Y2=0
cc_87 D1 N_Y_c_274_n 0.00882626f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_88 N_D1_M1000_g N_VPWR_c_352_n 0.00390896f $X=0.7 $Y=2.875 $X2=0 $Y2=0
cc_89 D1 N_VPWR_c_352_n 0.00665758f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_90 N_D1_M1000_g N_VPWR_c_350_n 0.00648016f $X=0.7 $Y=2.875 $X2=0 $Y2=0
cc_91 D1 N_VPWR_c_350_n 0.0087435f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_92 N_D1_M1009_g N_VGND_c_390_n 0.0111409f $X=0.7 $Y=0.445 $X2=0 $Y2=0
cc_93 N_D1_M1009_g N_VGND_c_391_n 0.0037993f $X=0.7 $Y=0.445 $X2=0 $Y2=0
cc_94 N_D1_M1009_g N_VGND_c_392_n 0.00144619f $X=0.7 $Y=0.445 $X2=0 $Y2=0
cc_95 N_D1_M1009_g N_VGND_c_396_n 0.00672233f $X=0.7 $Y=0.445 $X2=0 $Y2=0
cc_96 N_C1_M1003_g N_B1_M1001_g 0.0164047f $X=1.13 $Y=0.445 $X2=0 $Y2=0
cc_97 N_C1_c_109_n N_B1_M1001_g 0.0162927f $X=1.15 $Y=1.06 $X2=0 $Y2=0
cc_98 N_C1_c_110_n N_B1_M1001_g 0.0015165f $X=1.15 $Y=1.06 $X2=0 $Y2=0
cc_99 N_C1_M1007_g N_B1_c_146_n 0.0941586f $X=1.06 $Y=2.875 $X2=0 $Y2=0
cc_100 N_C1_c_108_n N_B1_c_146_n 0.00861019f $X=1.15 $Y=1.565 $X2=0 $Y2=0
cc_101 N_C1_c_110_n N_B1_c_146_n 0.00499835f $X=1.15 $Y=1.06 $X2=0 $Y2=0
cc_102 N_C1_M1007_g B1 3.25521e-19 $X=1.06 $Y=2.875 $X2=0 $Y2=0
cc_103 N_C1_c_107_n B1 0.00136466f $X=1.15 $Y=1.4 $X2=0 $Y2=0
cc_104 N_C1_c_110_n B1 0.0469867f $X=1.15 $Y=1.06 $X2=0 $Y2=0
cc_105 N_C1_c_107_n N_B1_c_148_n 0.00861019f $X=1.15 $Y=1.4 $X2=0 $Y2=0
cc_106 N_C1_c_110_n N_B1_c_148_n 0.00102432f $X=1.15 $Y=1.06 $X2=0 $Y2=0
cc_107 N_C1_c_110_n N_Y_c_270_n 0.00644024f $X=1.15 $Y=1.06 $X2=0 $Y2=0
cc_108 N_C1_M1003_g N_Y_c_273_n 0.0119771f $X=1.13 $Y=0.445 $X2=0 $Y2=0
cc_109 N_C1_c_109_n N_Y_c_273_n 0.00413226f $X=1.15 $Y=1.06 $X2=0 $Y2=0
cc_110 N_C1_c_110_n N_Y_c_273_n 0.0218921f $X=1.15 $Y=1.06 $X2=0 $Y2=0
cc_111 N_C1_M1003_g N_Y_c_274_n 0.00245315f $X=1.13 $Y=0.445 $X2=0 $Y2=0
cc_112 N_C1_c_109_n N_Y_c_274_n 0.00104965f $X=1.15 $Y=1.06 $X2=0 $Y2=0
cc_113 N_C1_c_110_n N_Y_c_274_n 0.00281001f $X=1.15 $Y=1.06 $X2=0 $Y2=0
cc_114 N_C1_M1007_g N_VPWR_c_352_n 0.00575161f $X=1.06 $Y=2.875 $X2=0 $Y2=0
cc_115 N_C1_M1007_g N_VPWR_c_350_n 0.0105591f $X=1.06 $Y=2.875 $X2=0 $Y2=0
cc_116 N_C1_M1003_g N_VGND_c_391_n 0.00408791f $X=1.13 $Y=0.445 $X2=0 $Y2=0
cc_117 N_C1_M1003_g N_VGND_c_392_n 0.00715019f $X=1.13 $Y=0.445 $X2=0 $Y2=0
cc_118 N_C1_M1003_g N_VGND_c_396_n 0.00477058f $X=1.13 $Y=0.445 $X2=0 $Y2=0
cc_119 N_B1_M1008_g N_A1_c_194_n 0.0327306f $X=1.42 $Y=2.875 $X2=-0.19
+ $Y2=-0.245
cc_120 N_B1_c_146_n N_A1_c_194_n 0.00555098f $X=1.69 $Y=1.805 $X2=-0.19
+ $Y2=-0.245
cc_121 N_B1_M1001_g N_A1_M1005_g 0.0398442f $X=1.71 $Y=0.445 $X2=0 $Y2=0
cc_122 B1 N_A1_M1005_g 0.00223763f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_123 N_B1_c_148_n N_A1_M1005_g 0.0136161f $X=1.69 $Y=1.45 $X2=0 $Y2=0
cc_124 N_B1_M1008_g N_A1_c_196_n 0.0039012f $X=1.42 $Y=2.875 $X2=0 $Y2=0
cc_125 N_B1_c_146_n N_A1_c_196_n 0.0136161f $X=1.69 $Y=1.805 $X2=0 $Y2=0
cc_126 B1 N_A1_c_196_n 0.00145265f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_127 N_B1_M1008_g A1 4.28516e-19 $X=1.42 $Y=2.875 $X2=0 $Y2=0
cc_128 N_B1_M1001_g A1 2.47048e-19 $X=1.71 $Y=0.445 $X2=0 $Y2=0
cc_129 B1 A1 0.0409089f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_130 N_B1_c_148_n A1 0.00247762f $X=1.69 $Y=1.45 $X2=0 $Y2=0
cc_131 N_B1_c_146_n N_A1_c_193_n 0.0136161f $X=1.69 $Y=1.805 $X2=0 $Y2=0
cc_132 N_B1_M1001_g N_Y_c_273_n 0.0133206f $X=1.71 $Y=0.445 $X2=0 $Y2=0
cc_133 B1 N_Y_c_273_n 0.00691228f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_134 N_B1_c_148_n N_Y_c_273_n 0.00443848f $X=1.69 $Y=1.45 $X2=0 $Y2=0
cc_135 N_B1_M1008_g N_A_299_533#_c_323_n 2.1266e-19 $X=1.42 $Y=2.875 $X2=0 $Y2=0
cc_136 N_B1_c_146_n N_A_299_533#_c_320_n 4.94017e-19 $X=1.69 $Y=1.805 $X2=0
+ $Y2=0
cc_137 B1 N_A_299_533#_c_320_n 0.00166719f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_138 N_B1_M1008_g N_A_299_533#_c_321_n 0.00551383f $X=1.42 $Y=2.875 $X2=0
+ $Y2=0
cc_139 N_B1_c_146_n N_A_299_533#_c_321_n 0.00280893f $X=1.69 $Y=1.805 $X2=0
+ $Y2=0
cc_140 B1 N_A_299_533#_c_321_n 0.00773039f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_141 N_B1_M1008_g N_VPWR_c_351_n 0.00145858f $X=1.42 $Y=2.875 $X2=0 $Y2=0
cc_142 N_B1_M1008_g N_VPWR_c_352_n 0.00575161f $X=1.42 $Y=2.875 $X2=0 $Y2=0
cc_143 N_B1_M1008_g N_VPWR_c_350_n 0.0107404f $X=1.42 $Y=2.875 $X2=0 $Y2=0
cc_144 N_B1_M1001_g N_VGND_c_392_n 0.00670425f $X=1.71 $Y=0.445 $X2=0 $Y2=0
cc_145 N_B1_M1001_g N_VGND_c_394_n 0.0042361f $X=1.71 $Y=0.445 $X2=0 $Y2=0
cc_146 N_B1_M1001_g N_VGND_c_396_n 0.0063986f $X=1.71 $Y=0.445 $X2=0 $Y2=0
cc_147 N_A1_M1005_g N_A2_M1002_g 0.0646536f $X=2.14 $Y=0.445 $X2=0 $Y2=0
cc_148 N_A1_M1004_g N_A2_c_241_n 0.013561f $X=1.85 $Y=2.875 $X2=0 $Y2=0
cc_149 N_A1_c_194_n N_A2_c_235_n 0.00281326f $X=1.85 $Y=2.345 $X2=0 $Y2=0
cc_150 N_A1_c_196_n N_A2_c_235_n 0.0069306f $X=2.23 $Y=2.03 $X2=0 $Y2=0
cc_151 A1 N_A2_c_236_n 0.00315206f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_152 N_A1_c_193_n N_A2_c_236_n 0.0069306f $X=2.23 $Y=1.69 $X2=0 $Y2=0
cc_153 N_A1_c_193_n A2 0.00307118f $X=2.23 $Y=1.69 $X2=0 $Y2=0
cc_154 N_A1_M1005_g N_A2_c_238_n 0.00391664f $X=2.14 $Y=0.445 $X2=0 $Y2=0
cc_155 A1 N_A2_c_238_n 0.00506934f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_156 N_A1_M1005_g N_Y_c_273_n 0.00451277f $X=2.14 $Y=0.445 $X2=0 $Y2=0
cc_157 N_A1_M1004_g N_A_299_533#_c_323_n 2.1266e-19 $X=1.85 $Y=2.875 $X2=0 $Y2=0
cc_158 N_A1_c_194_n N_A_299_533#_c_320_n 0.0129628f $X=1.85 $Y=2.345 $X2=0 $Y2=0
cc_159 N_A1_M1004_g N_A_299_533#_c_320_n 0.014573f $X=1.85 $Y=2.875 $X2=0 $Y2=0
cc_160 A1 N_A_299_533#_c_320_n 0.0127206f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_161 N_A1_M1004_g N_A_299_533#_c_322_n 6.39991e-19 $X=1.85 $Y=2.875 $X2=0
+ $Y2=0
cc_162 N_A1_M1004_g N_VPWR_c_351_n 0.00762129f $X=1.85 $Y=2.875 $X2=0 $Y2=0
cc_163 N_A1_M1004_g N_VPWR_c_352_n 0.0040762f $X=1.85 $Y=2.875 $X2=0 $Y2=0
cc_164 N_A1_M1004_g N_VPWR_c_350_n 0.00483784f $X=1.85 $Y=2.875 $X2=0 $Y2=0
cc_165 N_A1_M1005_g N_VGND_c_394_n 0.00585385f $X=2.14 $Y=0.445 $X2=0 $Y2=0
cc_166 N_A1_M1005_g N_VGND_c_396_n 0.0108402f $X=2.14 $Y=0.445 $X2=0 $Y2=0
cc_167 N_A2_c_239_n N_A_299_533#_c_320_n 0.00617495f $X=2.5 $Y=2.555 $X2=0 $Y2=0
cc_168 N_A2_c_241_n N_A_299_533#_c_320_n 0.00717092f $X=2.575 $Y=2.48 $X2=0
+ $Y2=0
cc_169 N_A2_c_239_n N_A_299_533#_c_322_n 0.00804233f $X=2.5 $Y=2.555 $X2=0 $Y2=0
cc_170 N_A2_c_240_n N_A_299_533#_c_322_n 0.0239803f $X=2.92 $Y=2.48 $X2=0 $Y2=0
cc_171 N_A2_c_241_n N_A_299_533#_c_322_n 0.00137668f $X=2.575 $Y=2.48 $X2=0
+ $Y2=0
cc_172 N_A2_c_239_n N_VPWR_c_351_n 0.00758468f $X=2.5 $Y=2.555 $X2=0 $Y2=0
cc_173 N_A2_c_239_n N_VPWR_c_353_n 0.00416887f $X=2.5 $Y=2.555 $X2=0 $Y2=0
cc_174 N_A2_c_240_n N_VPWR_c_353_n 0.00434323f $X=2.92 $Y=2.48 $X2=0 $Y2=0
cc_175 N_A2_c_239_n N_VPWR_c_350_n 0.00767456f $X=2.5 $Y=2.555 $X2=0 $Y2=0
cc_176 N_A2_c_240_n N_VPWR_c_350_n 0.00484438f $X=2.92 $Y=2.48 $X2=0 $Y2=0
cc_177 N_A2_M1002_g N_VGND_c_393_n 0.00460896f $X=2.5 $Y=0.445 $X2=0 $Y2=0
cc_178 N_A2_c_233_n N_VGND_c_393_n 0.00613384f $X=2.92 $Y=1.03 $X2=0 $Y2=0
cc_179 A2 N_VGND_c_393_n 0.00548489f $X=3.035 $Y=0.47 $X2=0 $Y2=0
cc_180 N_A2_M1002_g N_VGND_c_394_n 0.00585385f $X=2.5 $Y=0.445 $X2=0 $Y2=0
cc_181 A2 N_VGND_c_395_n 0.00608642f $X=3.035 $Y=0.47 $X2=0 $Y2=0
cc_182 N_A2_M1002_g N_VGND_c_396_n 0.0118303f $X=2.5 $Y=0.445 $X2=0 $Y2=0
cc_183 A2 N_VGND_c_396_n 0.00693478f $X=3.035 $Y=0.47 $X2=0 $Y2=0
cc_184 N_Y_c_270_n N_VPWR_c_352_n 0.00799973f $X=0.26 $Y=2.81 $X2=0 $Y2=0
cc_185 N_Y_M1000_s N_VPWR_c_350_n 0.0112101f $X=0.135 $Y=2.665 $X2=0 $Y2=0
cc_186 N_Y_c_270_n N_VPWR_c_350_n 0.00692256f $X=0.26 $Y=2.81 $X2=0 $Y2=0
cc_187 N_Y_c_273_n N_VGND_M1003_d 0.00372411f $X=1.82 $Y=0.71 $X2=0 $Y2=0
cc_188 N_Y_c_272_n N_VGND_c_389_n 0.0018725f $X=0.345 $Y=0.81 $X2=0 $Y2=0
cc_189 N_Y_c_271_n N_VGND_c_390_n 0.00821663f $X=0.635 $Y=0.81 $X2=0 $Y2=0
cc_190 N_Y_c_272_n N_VGND_c_390_n 0.00662208f $X=0.345 $Y=0.81 $X2=0 $Y2=0
cc_191 N_Y_c_274_n N_VGND_c_390_n 0.0144853f $X=0.827 $Y=0.71 $X2=0 $Y2=0
cc_192 N_Y_c_271_n N_VGND_c_391_n 0.00270512f $X=0.635 $Y=0.81 $X2=0 $Y2=0
cc_193 N_Y_c_273_n N_VGND_c_391_n 0.00275886f $X=1.82 $Y=0.71 $X2=0 $Y2=0
cc_194 N_Y_c_274_n N_VGND_c_391_n 0.0148452f $X=0.827 $Y=0.71 $X2=0 $Y2=0
cc_195 N_Y_c_273_n N_VGND_c_392_n 0.0195102f $X=1.82 $Y=0.71 $X2=0 $Y2=0
cc_196 N_Y_c_273_n N_VGND_c_394_n 0.00427222f $X=1.82 $Y=0.71 $X2=0 $Y2=0
cc_197 N_Y_c_310_p N_VGND_c_394_n 0.00813208f $X=1.925 $Y=0.51 $X2=0 $Y2=0
cc_198 N_Y_M1009_d N_VGND_c_396_n 0.00244615f $X=0.775 $Y=0.235 $X2=0 $Y2=0
cc_199 N_Y_M1001_d N_VGND_c_396_n 0.00367929f $X=1.785 $Y=0.235 $X2=0 $Y2=0
cc_200 N_Y_c_271_n N_VGND_c_396_n 0.00520629f $X=0.635 $Y=0.81 $X2=0 $Y2=0
cc_201 N_Y_c_272_n N_VGND_c_396_n 0.00351912f $X=0.345 $Y=0.81 $X2=0 $Y2=0
cc_202 N_Y_c_273_n N_VGND_c_396_n 0.0136331f $X=1.82 $Y=0.71 $X2=0 $Y2=0
cc_203 N_Y_c_310_p N_VGND_c_396_n 0.00760156f $X=1.925 $Y=0.51 $X2=0 $Y2=0
cc_204 N_Y_c_274_n N_VGND_c_396_n 0.013426f $X=0.827 $Y=0.71 $X2=0 $Y2=0
cc_205 A_155_533# N_VPWR_c_350_n 0.00802611f $X=0.775 $Y=2.665 $X2=3.12 $Y2=3.33
cc_206 A_227_533# N_VPWR_c_350_n 0.00899413f $X=1.135 $Y=2.665 $X2=3.12 $Y2=3.33
cc_207 N_A_299_533#_c_320_n N_VPWR_c_351_n 0.0220107f $X=2.55 $Y=2.57 $X2=0
+ $Y2=0
cc_208 N_A_299_533#_c_322_n N_VPWR_c_351_n 0.00401826f $X=2.715 $Y=2.57 $X2=0
+ $Y2=0
cc_209 N_A_299_533#_c_323_n N_VPWR_c_352_n 0.00785054f $X=1.635 $Y=2.81 $X2=0
+ $Y2=0
cc_210 N_A_299_533#_c_320_n N_VPWR_c_352_n 0.00273212f $X=2.55 $Y=2.57 $X2=0
+ $Y2=0
cc_211 N_A_299_533#_c_320_n N_VPWR_c_353_n 0.00479132f $X=2.55 $Y=2.57 $X2=0
+ $Y2=0
cc_212 N_A_299_533#_c_322_n N_VPWR_c_353_n 0.0100292f $X=2.715 $Y=2.57 $X2=0
+ $Y2=0
cc_213 N_A_299_533#_M1008_d N_VPWR_c_350_n 0.00371762f $X=1.495 $Y=2.665 $X2=0
+ $Y2=0
cc_214 N_A_299_533#_M1006_d N_VPWR_c_350_n 0.00235368f $X=2.575 $Y=2.665 $X2=0
+ $Y2=0
cc_215 N_A_299_533#_c_323_n N_VPWR_c_350_n 0.00757496f $X=1.635 $Y=2.81 $X2=0
+ $Y2=0
cc_216 N_A_299_533#_c_320_n N_VPWR_c_350_n 0.013411f $X=2.55 $Y=2.57 $X2=0 $Y2=0
cc_217 N_A_299_533#_c_322_n N_VPWR_c_350_n 0.0113031f $X=2.715 $Y=2.57 $X2=0
+ $Y2=0
cc_218 N_VGND_c_396_n A_443_47# 0.00899413f $X=3.12 $Y=0 $X2=-0.19 $Y2=-0.245
