* NGSPICE file created from sky130_fd_sc_lp__dlrtp_lp2.ext - technology: sky130A

.subckt sky130_fd_sc_lp__dlrtp_lp2 D GATE RESET_B VGND VNB VPB VPWR Q
M1000 Q a_898_21# VPWR VPB phighvt w=1e+06u l=250000u
+  ad=2.85e+11p pd=2.57e+06u as=1.96225e+12p ps=1.204e+07u
M1001 VPWR a_256_405# a_413_47# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=2.85e+11p ps=2.57e+06u
M1002 a_1216_57# a_736_47# a_898_21# VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=1.197e+11p ps=1.41e+06u
M1003 VGND RESET_B a_1216_57# VNB nshort w=420000u l=150000u
+  ad=7.43925e+11p pd=7.27e+06u as=0p ps=0u
M1004 VGND D a_114_122# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1005 a_740_419# a_27_122# VPWR VPB phighvt w=1e+06u l=250000u
+  ad=2.4e+11p pd=2.48e+06u as=0p ps=0u
M1006 a_944_419# a_413_47# a_736_47# VPB phighvt w=1e+06u l=250000u
+  ad=2.5e+11p pd=2.5e+06u as=2.8e+11p ps=2.56e+06u
M1007 VPWR RESET_B a_898_21# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=2.8e+11p ps=2.56e+06u
M1008 a_256_405# GATE a_294_185# VNB nshort w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=8.82e+10p ps=1.26e+06u
M1009 VPWR a_898_21# a_944_419# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_658_47# a_27_122# VGND VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1011 a_736_47# a_413_47# a_658_47# VNB nshort w=420000u l=150000u
+  ad=1.764e+11p pd=1.68e+06u as=0p ps=0u
M1012 a_1380_57# a_898_21# VGND VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1013 Q a_898_21# a_1380_57# VNB nshort w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=0p ps=0u
M1014 a_256_405# GATE VPWR VPB phighvt w=1e+06u l=250000u
+  ad=2.85e+11p pd=2.57e+06u as=0p ps=0u
M1015 VGND a_898_21# a_850_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1016 a_114_122# D a_27_122# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1017 a_294_185# GATE VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_850_47# a_256_405# a_736_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_736_47# a_256_405# a_740_419# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_898_21# a_736_47# VPWR VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_500_47# a_256_405# a_413_47# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=1.197e+11p ps=1.41e+06u
M1022 VPWR D a_27_122# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=2.85e+11p ps=2.57e+06u
M1023 VGND a_256_405# a_500_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

