* File: sky130_fd_sc_lp__and4_2.pxi.spice
* Created: Fri Aug 28 10:07:38 2020
* 
x_PM_SKY130_FD_SC_LP__AND4_2%A N_A_c_67_n N_A_M1010_g N_A_M1009_g N_A_c_69_n A A
+ N_A_c_70_n N_A_c_71_n PM_SKY130_FD_SC_LP__AND4_2%A
x_PM_SKY130_FD_SC_LP__AND4_2%B N_B_M1007_g N_B_M1003_g N_B_c_100_n N_B_c_101_n B
+ N_B_c_103_n PM_SKY130_FD_SC_LP__AND4_2%B
x_PM_SKY130_FD_SC_LP__AND4_2%C N_C_M1001_g N_C_M1005_g N_C_c_140_n N_C_c_141_n C
+ N_C_c_142_n N_C_c_150_n PM_SKY130_FD_SC_LP__AND4_2%C
x_PM_SKY130_FD_SC_LP__AND4_2%D N_D_M1006_g N_D_M1000_g N_D_c_176_n N_D_c_177_n D
+ N_D_c_178_n N_D_c_179_n PM_SKY130_FD_SC_LP__AND4_2%D
x_PM_SKY130_FD_SC_LP__AND4_2%A_72_49# N_A_72_49#_M1010_s N_A_72_49#_M1009_d
+ N_A_72_49#_M1005_d N_A_72_49#_M1002_g N_A_72_49#_M1004_g N_A_72_49#_M1008_g
+ N_A_72_49#_M1011_g N_A_72_49#_c_216_n N_A_72_49#_c_217_n N_A_72_49#_c_218_n
+ N_A_72_49#_c_223_n N_A_72_49#_c_243_n N_A_72_49#_c_224_n N_A_72_49#_c_219_n
+ N_A_72_49#_c_225_n N_A_72_49#_c_226_n N_A_72_49#_c_220_n
+ PM_SKY130_FD_SC_LP__AND4_2%A_72_49#
x_PM_SKY130_FD_SC_LP__AND4_2%VPWR N_VPWR_M1009_s N_VPWR_M1003_d N_VPWR_M1000_d
+ N_VPWR_M1011_s N_VPWR_c_316_n N_VPWR_c_317_n N_VPWR_c_318_n N_VPWR_c_319_n
+ N_VPWR_c_320_n N_VPWR_c_321_n N_VPWR_c_322_n N_VPWR_c_323_n N_VPWR_c_324_n
+ VPWR N_VPWR_c_325_n N_VPWR_c_326_n N_VPWR_c_327_n N_VPWR_c_315_n
+ PM_SKY130_FD_SC_LP__AND4_2%VPWR
x_PM_SKY130_FD_SC_LP__AND4_2%X N_X_M1002_d N_X_M1004_d X X X X X X X N_X_c_356_n
+ PM_SKY130_FD_SC_LP__AND4_2%X
x_PM_SKY130_FD_SC_LP__AND4_2%VGND N_VGND_M1006_d N_VGND_M1008_s N_VGND_c_376_n
+ N_VGND_c_377_n N_VGND_c_378_n N_VGND_c_379_n N_VGND_c_380_n VGND
+ N_VGND_c_381_n N_VGND_c_382_n PM_SKY130_FD_SC_LP__AND4_2%VGND
cc_1 VNB N_A_c_67_n 0.0260287f $X=-0.19 $Y=-0.245 $X2=0.597 $Y2=1.498
cc_2 VNB N_A_M1010_g 0.0356607f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=0.455
cc_3 VNB N_A_c_69_n 0.013206f $X=-0.19 $Y=-0.245 $X2=0.597 $Y2=1.675
cc_4 VNB N_A_c_70_n 0.020507f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.17
cc_5 VNB N_A_c_71_n 0.0420725f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.17
cc_6 VNB N_B_M1007_g 0.0231842f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.005
cc_7 VNB N_B_M1003_g 0.00362747f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.675
cc_8 VNB N_B_c_100_n 0.0187158f $X=-0.19 $Y=-0.245 $X2=0.597 $Y2=1.675
cc_9 VNB N_B_c_101_n 0.0147112f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_10 VNB B 0.00770422f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_11 VNB N_B_c_103_n 0.014718f $X=-0.19 $Y=-0.245 $X2=0.597 $Y2=1.17
cc_12 VNB N_C_M1001_g 0.0258829f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.005
cc_13 VNB N_C_M1005_g 0.00363285f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.675
cc_14 VNB N_C_c_140_n 0.0230433f $X=-0.19 $Y=-0.245 $X2=0.597 $Y2=1.675
cc_15 VNB N_C_c_141_n 0.0158082f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_16 VNB N_C_c_142_n 0.0158082f $X=-0.19 $Y=-0.245 $X2=0.597 $Y2=1.17
cc_17 VNB N_D_M1006_g 0.0280166f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.005
cc_18 VNB N_D_M1000_g 0.00327845f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.675
cc_19 VNB N_D_c_176_n 0.020845f $X=-0.19 $Y=-0.245 $X2=0.597 $Y2=1.675
cc_20 VNB N_D_c_177_n 0.014707f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_21 VNB N_D_c_178_n 0.0160533f $X=-0.19 $Y=-0.245 $X2=0.597 $Y2=1.17
cc_22 VNB N_D_c_179_n 0.00748241f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.17
cc_23 VNB N_A_72_49#_M1002_g 0.0253493f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_24 VNB N_A_72_49#_M1008_g 0.0335493f $X=-0.19 $Y=-0.245 $X2=0.377 $Y2=1.17
cc_25 VNB N_A_72_49#_c_216_n 0.0147786f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_72_49#_c_217_n 0.046799f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_72_49#_c_218_n 0.00983942f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_72_49#_c_219_n 0.00183986f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_72_49#_c_220_n 0.058432f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VPWR_c_315_n 0.163682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_X_c_356_n 0.00450975f $X=-0.19 $Y=-0.245 $X2=0.377 $Y2=1.295
cc_32 VNB N_VGND_c_376_n 0.00602232f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=2.045
cc_33 VNB N_VGND_c_377_n 0.0117664f $X=-0.19 $Y=-0.245 $X2=0.597 $Y2=1.675
cc_34 VNB N_VGND_c_378_n 0.0505793f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_35 VNB N_VGND_c_379_n 0.0671958f $X=-0.19 $Y=-0.245 $X2=0.597 $Y2=1.17
cc_36 VNB N_VGND_c_380_n 0.00631622f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=1.17
cc_37 VNB N_VGND_c_381_n 0.0204928f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_382_n 0.218551f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VPB N_A_M1009_g 0.0275447f $X=-0.19 $Y=1.655 $X2=0.7 $Y2=2.045
cc_40 VPB N_A_c_69_n 0.0075696f $X=-0.19 $Y=1.655 $X2=0.597 $Y2=1.675
cc_41 VPB N_A_c_71_n 0.0167584f $X=-0.19 $Y=1.655 $X2=0.585 $Y2=1.17
cc_42 VPB N_B_M1003_g 0.0252724f $X=-0.19 $Y=1.655 $X2=0.7 $Y2=1.675
cc_43 VPB N_C_M1005_g 0.0253774f $X=-0.19 $Y=1.655 $X2=0.7 $Y2=1.675
cc_44 VPB N_D_M1000_g 0.0241773f $X=-0.19 $Y=1.655 $X2=0.7 $Y2=1.675
cc_45 VPB N_A_72_49#_M1004_g 0.0210269f $X=-0.19 $Y=1.655 $X2=0.597 $Y2=1.17
cc_46 VPB N_A_72_49#_M1011_g 0.0255346f $X=-0.19 $Y=1.655 $X2=0.377 $Y2=1.665
cc_47 VPB N_A_72_49#_c_223_n 0.00861667f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_48 VPB N_A_72_49#_c_224_n 0.0080783f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_49 VPB N_A_72_49#_c_225_n 0.0169688f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_50 VPB N_A_72_49#_c_226_n 0.00722547f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_51 VPB N_A_72_49#_c_220_n 0.0125093f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_52 VPB N_VPWR_c_316_n 0.0676358f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_53 VPB N_VPWR_c_317_n 0.0377459f $X=-0.19 $Y=1.655 $X2=0.597 $Y2=1.005
cc_54 VPB N_VPWR_c_318_n 0.021305f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_55 VPB N_VPWR_c_319_n 0.0117405f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_56 VPB N_VPWR_c_320_n 0.0653393f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_57 VPB N_VPWR_c_321_n 0.0123263f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_58 VPB N_VPWR_c_322_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_59 VPB N_VPWR_c_323_n 0.0199842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_60 VPB N_VPWR_c_324_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_61 VPB N_VPWR_c_325_n 0.0206207f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_62 VPB N_VPWR_c_326_n 0.0148832f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_63 VPB N_VPWR_c_327_n 0.0102056f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_64 VPB N_VPWR_c_315_n 0.106923f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_65 VPB N_X_c_356_n 0.00234245f $X=-0.19 $Y=1.655 $X2=0.377 $Y2=1.295
cc_66 N_A_M1010_g N_B_M1007_g 0.0237638f $X=0.7 $Y=0.455 $X2=0 $Y2=0
cc_67 N_A_c_69_n N_B_M1003_g 0.0178962f $X=0.597 $Y=1.675 $X2=0 $Y2=0
cc_68 N_A_c_71_n N_B_M1003_g 4.97281e-19 $X=0.585 $Y=1.17 $X2=0 $Y2=0
cc_69 N_A_c_67_n N_B_c_100_n 0.0237638f $X=0.597 $Y=1.498 $X2=0 $Y2=0
cc_70 N_A_c_69_n N_B_c_101_n 0.0237638f $X=0.597 $Y=1.675 $X2=0 $Y2=0
cc_71 N_A_c_71_n N_B_c_101_n 4.50813e-19 $X=0.585 $Y=1.17 $X2=0 $Y2=0
cc_72 N_A_c_70_n B 0.00192966f $X=0.585 $Y=1.17 $X2=0 $Y2=0
cc_73 N_A_c_71_n B 0.0245157f $X=0.585 $Y=1.17 $X2=0 $Y2=0
cc_74 N_A_c_70_n N_B_c_103_n 0.0237638f $X=0.585 $Y=1.17 $X2=0 $Y2=0
cc_75 N_A_c_71_n N_B_c_103_n 5.43311e-19 $X=0.585 $Y=1.17 $X2=0 $Y2=0
cc_76 N_A_M1010_g N_A_72_49#_c_216_n 0.00697863f $X=0.7 $Y=0.455 $X2=0 $Y2=0
cc_77 N_A_M1010_g N_A_72_49#_c_217_n 0.0113324f $X=0.7 $Y=0.455 $X2=0 $Y2=0
cc_78 N_A_c_71_n N_A_72_49#_c_217_n 0.00141328f $X=0.585 $Y=1.17 $X2=0 $Y2=0
cc_79 N_A_M1010_g N_A_72_49#_c_218_n 0.00415813f $X=0.7 $Y=0.455 $X2=0 $Y2=0
cc_80 N_A_c_70_n N_A_72_49#_c_218_n 0.00156669f $X=0.585 $Y=1.17 $X2=0 $Y2=0
cc_81 N_A_c_71_n N_A_72_49#_c_218_n 0.0292631f $X=0.585 $Y=1.17 $X2=0 $Y2=0
cc_82 N_A_M1009_g N_A_72_49#_c_225_n 0.00534714f $X=0.7 $Y=2.045 $X2=0 $Y2=0
cc_83 N_A_c_71_n N_A_72_49#_c_225_n 0.00570506f $X=0.585 $Y=1.17 $X2=0 $Y2=0
cc_84 N_A_M1009_g N_VPWR_c_316_n 0.00967789f $X=0.7 $Y=2.045 $X2=0 $Y2=0
cc_85 N_A_c_69_n N_VPWR_c_316_n 0.00117248f $X=0.597 $Y=1.675 $X2=0 $Y2=0
cc_86 N_A_c_71_n N_VPWR_c_316_n 0.0274351f $X=0.585 $Y=1.17 $X2=0 $Y2=0
cc_87 N_A_M1010_g N_VGND_c_379_n 0.00411983f $X=0.7 $Y=0.455 $X2=0 $Y2=0
cc_88 N_A_M1010_g N_VGND_c_382_n 0.00679885f $X=0.7 $Y=0.455 $X2=0 $Y2=0
cc_89 N_B_M1007_g N_C_M1001_g 0.0285467f $X=1.06 $Y=0.455 $X2=0 $Y2=0
cc_90 N_B_M1003_g N_C_M1005_g 0.0146288f $X=1.13 $Y=2.045 $X2=0 $Y2=0
cc_91 N_B_c_100_n N_C_c_140_n 0.0145549f $X=1.15 $Y=1.43 $X2=0 $Y2=0
cc_92 N_B_c_101_n N_C_c_141_n 0.0145549f $X=1.15 $Y=1.595 $X2=0 $Y2=0
cc_93 B N_C_c_142_n 0.00289107f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_94 N_B_c_103_n N_C_c_142_n 0.0145549f $X=1.15 $Y=1.09 $X2=0 $Y2=0
cc_95 B N_C_c_150_n 0.0406944f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_96 N_B_c_103_n N_C_c_150_n 5.82269e-19 $X=1.15 $Y=1.09 $X2=0 $Y2=0
cc_97 N_B_M1007_g N_A_72_49#_c_216_n 0.00187772f $X=1.06 $Y=0.455 $X2=0 $Y2=0
cc_98 N_B_M1007_g N_A_72_49#_c_217_n 0.0120044f $X=1.06 $Y=0.455 $X2=0 $Y2=0
cc_99 B N_A_72_49#_c_217_n 0.0283757f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_100 N_B_c_103_n N_A_72_49#_c_217_n 0.00516293f $X=1.15 $Y=1.09 $X2=0 $Y2=0
cc_101 N_B_M1003_g N_A_72_49#_c_223_n 0.0118175f $X=1.13 $Y=2.045 $X2=0 $Y2=0
cc_102 N_B_c_101_n N_A_72_49#_c_223_n 0.00313676f $X=1.15 $Y=1.595 $X2=0 $Y2=0
cc_103 B N_A_72_49#_c_223_n 0.0210507f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_104 N_B_M1003_g N_A_72_49#_c_243_n 7.81681e-19 $X=1.13 $Y=2.045 $X2=0 $Y2=0
cc_105 N_B_M1003_g N_A_72_49#_c_225_n 0.00988818f $X=1.13 $Y=2.045 $X2=0 $Y2=0
cc_106 N_B_c_101_n N_A_72_49#_c_225_n 0.00208596f $X=1.15 $Y=1.595 $X2=0 $Y2=0
cc_107 B N_A_72_49#_c_225_n 0.00803702f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_108 N_B_M1003_g N_VPWR_c_316_n 4.80874e-19 $X=1.13 $Y=2.045 $X2=0 $Y2=0
cc_109 N_B_M1003_g N_VPWR_c_317_n 0.0043959f $X=1.13 $Y=2.045 $X2=0 $Y2=0
cc_110 N_B_M1007_g N_VGND_c_379_n 0.00421031f $X=1.06 $Y=0.455 $X2=0 $Y2=0
cc_111 N_B_M1007_g N_VGND_c_382_n 0.00609929f $X=1.06 $Y=0.455 $X2=0 $Y2=0
cc_112 N_C_M1001_g N_D_M1006_g 0.0275597f $X=1.6 $Y=0.455 $X2=0 $Y2=0
cc_113 N_C_M1005_g N_D_M1000_g 0.0179728f $X=1.78 $Y=2.045 $X2=0 $Y2=0
cc_114 N_C_c_140_n N_D_c_176_n 0.0145549f $X=1.69 $Y=1.43 $X2=0 $Y2=0
cc_115 N_C_c_141_n N_D_c_177_n 0.0145549f $X=1.69 $Y=1.595 $X2=0 $Y2=0
cc_116 N_C_c_142_n N_D_c_178_n 0.0145549f $X=1.69 $Y=1.09 $X2=0 $Y2=0
cc_117 N_C_c_150_n N_D_c_178_n 5.82269e-19 $X=1.69 $Y=1.09 $X2=0 $Y2=0
cc_118 N_C_c_142_n N_D_c_179_n 0.00289107f $X=1.69 $Y=1.09 $X2=0 $Y2=0
cc_119 N_C_c_150_n N_D_c_179_n 0.0406944f $X=1.69 $Y=1.09 $X2=0 $Y2=0
cc_120 N_C_M1001_g N_A_72_49#_c_217_n 0.0130064f $X=1.6 $Y=0.455 $X2=0 $Y2=0
cc_121 N_C_c_142_n N_A_72_49#_c_217_n 0.00521111f $X=1.69 $Y=1.09 $X2=0 $Y2=0
cc_122 N_C_c_150_n N_A_72_49#_c_217_n 0.0250619f $X=1.69 $Y=1.09 $X2=0 $Y2=0
cc_123 N_C_M1005_g N_A_72_49#_c_223_n 0.0118124f $X=1.78 $Y=2.045 $X2=0 $Y2=0
cc_124 N_C_c_141_n N_A_72_49#_c_223_n 0.00521111f $X=1.69 $Y=1.595 $X2=0 $Y2=0
cc_125 N_C_c_150_n N_A_72_49#_c_223_n 0.0232429f $X=1.69 $Y=1.09 $X2=0 $Y2=0
cc_126 N_C_M1005_g N_A_72_49#_c_243_n 0.00672015f $X=1.78 $Y=2.045 $X2=0 $Y2=0
cc_127 N_C_M1005_g N_A_72_49#_c_225_n 7.9114e-19 $X=1.78 $Y=2.045 $X2=0 $Y2=0
cc_128 N_C_M1005_g N_A_72_49#_c_226_n 0.00265346f $X=1.78 $Y=2.045 $X2=0 $Y2=0
cc_129 N_C_c_150_n N_A_72_49#_c_226_n 0.00195053f $X=1.69 $Y=1.09 $X2=0 $Y2=0
cc_130 N_C_M1005_g N_VPWR_c_317_n 0.00460817f $X=1.78 $Y=2.045 $X2=0 $Y2=0
cc_131 N_C_M1005_g N_VPWR_c_318_n 4.72952e-19 $X=1.78 $Y=2.045 $X2=0 $Y2=0
cc_132 N_C_M1001_g N_VGND_c_379_n 0.00421031f $X=1.6 $Y=0.455 $X2=0 $Y2=0
cc_133 N_C_M1001_g N_VGND_c_382_n 0.00652274f $X=1.6 $Y=0.455 $X2=0 $Y2=0
cc_134 N_D_M1006_g N_A_72_49#_M1002_g 0.0125545f $X=2.14 $Y=0.455 $X2=0 $Y2=0
cc_135 N_D_c_178_n N_A_72_49#_M1002_g 0.0101019f $X=2.23 $Y=1.09 $X2=0 $Y2=0
cc_136 N_D_c_179_n N_A_72_49#_M1002_g 3.17819e-19 $X=2.23 $Y=1.09 $X2=0 $Y2=0
cc_137 N_D_M1000_g N_A_72_49#_M1004_g 0.00944965f $X=2.21 $Y=2.045 $X2=0 $Y2=0
cc_138 N_D_M1006_g N_A_72_49#_c_217_n 0.0137823f $X=2.14 $Y=0.455 $X2=0 $Y2=0
cc_139 N_D_c_178_n N_A_72_49#_c_217_n 0.00516293f $X=2.23 $Y=1.09 $X2=0 $Y2=0
cc_140 N_D_c_179_n N_A_72_49#_c_217_n 0.0283757f $X=2.23 $Y=1.09 $X2=0 $Y2=0
cc_141 N_D_M1000_g N_A_72_49#_c_224_n 0.0150087f $X=2.21 $Y=2.045 $X2=0 $Y2=0
cc_142 N_D_c_177_n N_A_72_49#_c_224_n 0.00443672f $X=2.23 $Y=1.595 $X2=0 $Y2=0
cc_143 N_D_c_179_n N_A_72_49#_c_224_n 0.0231101f $X=2.23 $Y=1.09 $X2=0 $Y2=0
cc_144 N_D_M1006_g N_A_72_49#_c_219_n 0.00172705f $X=2.14 $Y=0.455 $X2=0 $Y2=0
cc_145 N_D_M1000_g N_A_72_49#_c_219_n 6.75623e-19 $X=2.21 $Y=2.045 $X2=0 $Y2=0
cc_146 N_D_c_176_n N_A_72_49#_c_219_n 2.13583e-19 $X=2.23 $Y=1.43 $X2=0 $Y2=0
cc_147 N_D_c_177_n N_A_72_49#_c_219_n 5.80416e-19 $X=2.23 $Y=1.595 $X2=0 $Y2=0
cc_148 N_D_c_178_n N_A_72_49#_c_219_n 0.00322536f $X=2.23 $Y=1.09 $X2=0 $Y2=0
cc_149 N_D_c_179_n N_A_72_49#_c_219_n 0.0331286f $X=2.23 $Y=1.09 $X2=0 $Y2=0
cc_150 N_D_c_177_n N_A_72_49#_c_226_n 7.43484e-19 $X=2.23 $Y=1.595 $X2=0 $Y2=0
cc_151 N_D_c_179_n N_A_72_49#_c_226_n 0.00571126f $X=2.23 $Y=1.09 $X2=0 $Y2=0
cc_152 N_D_M1000_g N_A_72_49#_c_220_n 0.00355803f $X=2.21 $Y=2.045 $X2=0 $Y2=0
cc_153 N_D_c_176_n N_A_72_49#_c_220_n 0.017097f $X=2.23 $Y=1.43 $X2=0 $Y2=0
cc_154 N_D_c_179_n N_A_72_49#_c_220_n 6.8244e-19 $X=2.23 $Y=1.09 $X2=0 $Y2=0
cc_155 N_D_M1000_g N_VPWR_c_318_n 0.00856564f $X=2.21 $Y=2.045 $X2=0 $Y2=0
cc_156 N_D_M1006_g N_VGND_c_376_n 0.00961203f $X=2.14 $Y=0.455 $X2=0 $Y2=0
cc_157 N_D_M1006_g N_VGND_c_379_n 0.00421031f $X=2.14 $Y=0.455 $X2=0 $Y2=0
cc_158 N_D_M1006_g N_VGND_c_382_n 0.00688986f $X=2.14 $Y=0.455 $X2=0 $Y2=0
cc_159 N_A_72_49#_c_223_n N_VPWR_M1003_d 0.00584696f $X=1.83 $Y=1.77 $X2=0 $Y2=0
cc_160 N_A_72_49#_c_224_n N_VPWR_M1000_d 0.00464424f $X=2.605 $Y=1.77 $X2=0
+ $Y2=0
cc_161 N_A_72_49#_c_225_n N_VPWR_c_316_n 0.0129796f $X=0.95 $Y=1.77 $X2=0 $Y2=0
cc_162 N_A_72_49#_c_223_n N_VPWR_c_317_n 0.0266856f $X=1.83 $Y=1.77 $X2=0 $Y2=0
cc_163 N_A_72_49#_c_243_n N_VPWR_c_317_n 0.011577f $X=1.995 $Y=2.045 $X2=0 $Y2=0
cc_164 N_A_72_49#_c_225_n N_VPWR_c_317_n 0.0158962f $X=0.95 $Y=1.77 $X2=0 $Y2=0
cc_165 N_A_72_49#_M1004_g N_VPWR_c_318_n 0.0230606f $X=2.905 $Y=2.465 $X2=0
+ $Y2=0
cc_166 N_A_72_49#_M1011_g N_VPWR_c_318_n 7.73703e-19 $X=3.335 $Y=2.465 $X2=0
+ $Y2=0
cc_167 N_A_72_49#_c_224_n N_VPWR_c_318_n 0.0403257f $X=2.605 $Y=1.77 $X2=0 $Y2=0
cc_168 N_A_72_49#_c_220_n N_VPWR_c_318_n 0.00104047f $X=3.335 $Y=1.51 $X2=0
+ $Y2=0
cc_169 N_A_72_49#_M1011_g N_VPWR_c_320_n 0.0076281f $X=3.335 $Y=2.465 $X2=0
+ $Y2=0
cc_170 N_A_72_49#_M1004_g N_VPWR_c_326_n 0.00486043f $X=2.905 $Y=2.465 $X2=0
+ $Y2=0
cc_171 N_A_72_49#_M1011_g N_VPWR_c_326_n 0.00585385f $X=3.335 $Y=2.465 $X2=0
+ $Y2=0
cc_172 N_A_72_49#_M1004_g N_VPWR_c_315_n 0.00824727f $X=2.905 $Y=2.465 $X2=0
+ $Y2=0
cc_173 N_A_72_49#_M1011_g N_VPWR_c_315_n 0.0114959f $X=3.335 $Y=2.465 $X2=0
+ $Y2=0
cc_174 N_A_72_49#_M1002_g N_X_c_356_n 0.00245966f $X=2.905 $Y=0.665 $X2=0 $Y2=0
cc_175 N_A_72_49#_M1004_g N_X_c_356_n 0.00180916f $X=2.905 $Y=2.465 $X2=0 $Y2=0
cc_176 N_A_72_49#_M1008_g N_X_c_356_n 0.00722653f $X=3.335 $Y=0.665 $X2=0 $Y2=0
cc_177 N_A_72_49#_M1011_g N_X_c_356_n 0.00462542f $X=3.335 $Y=2.465 $X2=0 $Y2=0
cc_178 N_A_72_49#_c_224_n N_X_c_356_n 0.013055f $X=2.605 $Y=1.77 $X2=0 $Y2=0
cc_179 N_A_72_49#_c_219_n N_X_c_356_n 0.0527337f $X=2.77 $Y=1.51 $X2=0 $Y2=0
cc_180 N_A_72_49#_c_220_n N_X_c_356_n 0.0296325f $X=3.335 $Y=1.51 $X2=0 $Y2=0
cc_181 N_A_72_49#_c_217_n N_VGND_M1006_d 0.00513639f $X=2.605 $Y=0.75 $X2=-0.19
+ $Y2=-0.245
cc_182 N_A_72_49#_c_219_n N_VGND_M1006_d 0.00365568f $X=2.77 $Y=1.51 $X2=-0.19
+ $Y2=-0.245
cc_183 N_A_72_49#_M1002_g N_VGND_c_376_n 0.00587184f $X=2.905 $Y=0.665 $X2=0
+ $Y2=0
cc_184 N_A_72_49#_c_217_n N_VGND_c_376_n 0.026125f $X=2.605 $Y=0.75 $X2=0 $Y2=0
cc_185 N_A_72_49#_M1008_g N_VGND_c_378_n 0.00844812f $X=3.335 $Y=0.665 $X2=0
+ $Y2=0
cc_186 N_A_72_49#_c_216_n N_VGND_c_379_n 0.0169541f $X=0.485 $Y=0.455 $X2=0
+ $Y2=0
cc_187 N_A_72_49#_c_217_n N_VGND_c_379_n 0.0281903f $X=2.605 $Y=0.75 $X2=0 $Y2=0
cc_188 N_A_72_49#_M1002_g N_VGND_c_381_n 0.00549449f $X=2.905 $Y=0.665 $X2=0
+ $Y2=0
cc_189 N_A_72_49#_M1008_g N_VGND_c_381_n 0.00575161f $X=3.335 $Y=0.665 $X2=0
+ $Y2=0
cc_190 N_A_72_49#_c_217_n N_VGND_c_381_n 0.00242794f $X=2.605 $Y=0.75 $X2=0
+ $Y2=0
cc_191 N_A_72_49#_M1010_s N_VGND_c_382_n 0.00214692f $X=0.36 $Y=0.245 $X2=0
+ $Y2=0
cc_192 N_A_72_49#_M1002_g N_VGND_c_382_n 0.0106452f $X=2.905 $Y=0.665 $X2=0
+ $Y2=0
cc_193 N_A_72_49#_M1008_g N_VGND_c_382_n 0.0115088f $X=3.335 $Y=0.665 $X2=0
+ $Y2=0
cc_194 N_A_72_49#_c_216_n N_VGND_c_382_n 0.0123289f $X=0.485 $Y=0.455 $X2=0
+ $Y2=0
cc_195 N_A_72_49#_c_217_n N_VGND_c_382_n 0.0511466f $X=2.605 $Y=0.75 $X2=0 $Y2=0
cc_196 N_VPWR_c_315_n N_X_M1004_d 0.00397496f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_197 N_VPWR_c_320_n N_X_c_356_n 0.00152359f $X=3.55 $Y=1.98 $X2=0 $Y2=0
cc_198 N_VPWR_c_326_n N_X_c_356_n 0.0138717f $X=3.425 $Y=3.33 $X2=0 $Y2=0
cc_199 N_VPWR_c_315_n N_X_c_356_n 0.00886411f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_200 N_X_c_356_n N_VGND_c_378_n 0.00152359f $X=3.12 $Y=0.42 $X2=0 $Y2=0
cc_201 N_X_c_356_n N_VGND_c_381_n 0.0138717f $X=3.12 $Y=0.42 $X2=0 $Y2=0
cc_202 N_X_M1002_d N_VGND_c_382_n 0.00397496f $X=2.98 $Y=0.245 $X2=0 $Y2=0
cc_203 N_X_c_356_n N_VGND_c_382_n 0.00886411f $X=3.12 $Y=0.42 $X2=0 $Y2=0
cc_204 A_155_49# N_VGND_c_382_n 0.00253354f $X=0.775 $Y=0.245 $X2=3.6 $Y2=0
cc_205 A_227_49# N_VGND_c_382_n 0.00470514f $X=1.135 $Y=0.245 $X2=3.6 $Y2=0
cc_206 A_335_49# N_VGND_c_382_n 0.00470514f $X=1.675 $Y=0.245 $X2=3.6 $Y2=0
