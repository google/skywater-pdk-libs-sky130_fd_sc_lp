* File: sky130_fd_sc_lp__nand3b_lp.spice
* Created: Wed Sep  2 10:05:06 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__nand3b_lp.pex.spice"
.subckt sky130_fd_sc_lp__nand3b_lp  VNB VPB B C A_N Y VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Y	Y
* A_N	A_N
* C	C
* B	B
* VPB	VPB
* VNB	VNB
MM1000 A_156_141# N_A_90_247#_M1000_g N_Y_M1000_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.1197 PD=0.66 PS=1.41 NRD=18.564 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.9 A=0.063 P=1.14 MULT=1
MM1005 A_234_141# N_B_M1005_g A_156_141# VNB NSHORT L=0.15 W=0.42 AD=0.0504
+ AS=0.0504 PD=0.66 PS=0.66 NRD=18.564 NRS=18.564 M=1 R=2.8 SA=75000.6
+ SB=75001.5 A=0.063 P=1.14 MULT=1
MM1002 N_VGND_M1002_d N_C_M1002_g A_234_141# VNB NSHORT L=0.15 W=0.42 AD=0.0819
+ AS=0.0504 PD=0.81 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75001 SB=75001.1
+ A=0.063 P=1.14 MULT=1
MM1006 A_420_141# N_A_N_M1006_g N_VGND_M1002_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0819 PD=0.63 PS=0.81 NRD=14.28 NRS=31.428 M=1 R=2.8 SA=75001.5
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1004 N_A_90_247#_M1004_d N_A_N_M1004_g A_420_141# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.9
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1007 N_VPWR_M1007_d N_A_90_247#_M1007_g N_Y_M1007_s VPB PHIGHVT L=0.25 W=1
+ AD=0.14 AS=0.285 PD=1.28 PS=2.57 NRD=0 NRS=0 M=1 R=4 SA=125000 SB=125002
+ A=0.25 P=2.5 MULT=1
MM1003 N_Y_M1003_d N_B_M1003_g N_VPWR_M1007_d VPB PHIGHVT L=0.25 W=1 AD=0.14
+ AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125001 SB=125001 A=0.25 P=2.5
+ MULT=1
MM1001 N_VPWR_M1001_d N_C_M1001_g N_Y_M1003_d VPB PHIGHVT L=0.25 W=1 AD=0.16
+ AS=0.14 PD=1.32 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125001 SB=125001 A=0.25 P=2.5
+ MULT=1
MM1008 N_A_90_247#_M1008_d N_A_N_M1008_g N_VPWR_M1001_d VPB PHIGHVT L=0.25 W=1
+ AD=0.285 AS=0.16 PD=2.57 PS=1.32 NRD=0 NRS=7.8603 M=1 R=4 SA=125002 SB=125000
+ A=0.25 P=2.5 MULT=1
DX9_noxref VNB VPB NWDIODE A=6.0799 P=10.25
*
.include "sky130_fd_sc_lp__nand3b_lp.pxi.spice"
*
.ends
*
*
