* File: sky130_fd_sc_lp__o2bb2ai_m.spice
* Created: Wed Sep  2 10:22:38 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__o2bb2ai_m.pex.spice"
.subckt sky130_fd_sc_lp__o2bb2ai_m  VNB VPB A1_N A2_N B2 B1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B1	B1
* B2	B2
* A2_N	A2_N
* A1_N	A1_N
* VPB	VPB
* VNB	VNB
MM1006 A_116_81# N_A1_N_M1006_g N_VGND_M1006_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1113 PD=0.63 PS=1.37 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1000 N_A_110_535#_M1000_d N_A2_N_M1000_g A_116_81# VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.0441 PD=1.37 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1003 N_A_410_78#_M1003_d N_A_110_535#_M1003_g N_Y_M1003_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1009 N_VGND_M1009_d N_B2_M1009_g N_A_410_78#_M1003_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1001 N_A_410_78#_M1001_d N_B1_M1001_g N_VGND_M1009_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.1 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1008 N_A_110_535#_M1008_d N_A1_N_M1008_g N_VPWR_M1008_s VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.9 A=0.063 P=1.14 MULT=1
MM1004 N_VPWR_M1004_d N_A2_N_M1004_g N_A_110_535#_M1008_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0819 AS=0.0588 PD=0.81 PS=0.7 NRD=9.3772 NRS=0 M=1 R=2.8
+ SA=75000.6 SB=75001.5 A=0.063 P=1.14 MULT=1
MM1007 N_Y_M1007_d N_A_110_535#_M1007_g N_VPWR_M1004_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0588 AS=0.0819 PD=0.7 PS=0.81 NRD=0 NRS=42.1974 M=1 R=2.8 SA=75001.2
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1002 A_390_535# N_B2_M1002_g N_Y_M1007_d VPB PHIGHVT L=0.15 W=0.42 AD=0.0441
+ AS=0.0588 PD=0.63 PS=0.7 NRD=23.443 NRS=0 M=1 R=2.8 SA=75001.6 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1005 N_VPWR_M1005_d N_B1_M1005_g A_390_535# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.1113 AS=0.0441 PD=1.37 PS=0.63 NRD=0 NRS=23.443 M=1 R=2.8 SA=75001.9
+ SB=75000.2 A=0.063 P=1.14 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9751 P=11.21
*
.include "sky130_fd_sc_lp__o2bb2ai_m.pxi.spice"
*
.ends
*
*
