* File: sky130_fd_sc_lp__nor2b_lp.pxi.spice
* Created: Wed Sep  2 10:08:34 2020
* 
x_PM_SKY130_FD_SC_LP__NOR2B_LP%A N_A_M1000_g N_A_M1004_g N_A_M1001_g N_A_c_67_n
+ N_A_c_68_n A A A N_A_c_70_n PM_SKY130_FD_SC_LP__NOR2B_LP%A
x_PM_SKY130_FD_SC_LP__NOR2B_LP%A_303_300# N_A_303_300#_M1007_d
+ N_A_303_300#_M1003_d N_A_303_300#_c_100_n N_A_303_300#_M1008_g
+ N_A_303_300#_M1005_g N_A_303_300#_c_103_n N_A_303_300#_M1002_g
+ N_A_303_300#_c_105_n N_A_303_300#_c_106_n N_A_303_300#_c_107_n
+ N_A_303_300#_c_108_n N_A_303_300#_c_109_n N_A_303_300#_c_110_n
+ N_A_303_300#_c_111_n N_A_303_300#_c_112_n N_A_303_300#_c_118_n
+ N_A_303_300#_c_113_n N_A_303_300#_c_119_n N_A_303_300#_c_114_n
+ PM_SKY130_FD_SC_LP__NOR2B_LP%A_303_300#
x_PM_SKY130_FD_SC_LP__NOR2B_LP%B_N N_B_N_c_189_n N_B_N_M1006_g N_B_N_c_190_n
+ N_B_N_c_191_n N_B_N_c_192_n N_B_N_M1003_g N_B_N_c_193_n N_B_N_M1007_g
+ N_B_N_c_199_n N_B_N_c_194_n B_N B_N N_B_N_c_196_n N_B_N_c_197_n
+ PM_SKY130_FD_SC_LP__NOR2B_LP%B_N
x_PM_SKY130_FD_SC_LP__NOR2B_LP%VPWR N_VPWR_M1004_s N_VPWR_M1003_s N_VPWR_c_239_n
+ N_VPWR_c_240_n N_VPWR_c_241_n N_VPWR_c_242_n VPWR N_VPWR_c_243_n
+ N_VPWR_c_238_n N_VPWR_c_245_n PM_SKY130_FD_SC_LP__NOR2B_LP%VPWR
x_PM_SKY130_FD_SC_LP__NOR2B_LP%Y N_Y_M1001_d N_Y_M1008_d Y Y Y Y Y Y Y
+ N_Y_c_268_n Y PM_SKY130_FD_SC_LP__NOR2B_LP%Y
x_PM_SKY130_FD_SC_LP__NOR2B_LP%VGND N_VGND_M1000_s N_VGND_M1002_d N_VGND_c_305_n
+ N_VGND_c_306_n VGND N_VGND_c_307_n N_VGND_c_308_n N_VGND_c_309_n
+ N_VGND_c_310_n N_VGND_c_311_n N_VGND_c_312_n PM_SKY130_FD_SC_LP__NOR2B_LP%VGND
cc_1 VNB N_A_M1000_g 0.0430814f $X=-0.19 $Y=-0.245 $X2=0.9 $Y2=0.495
cc_2 VNB N_A_M1001_g 0.0303456f $X=-0.19 $Y=-0.245 $X2=1.26 $Y2=0.495
cc_3 VNB N_A_c_67_n 0.0192252f $X=-0.19 $Y=-0.245 $X2=1.08 $Y2=1.26
cc_4 VNB N_A_c_68_n 0.00879153f $X=-0.19 $Y=-0.245 $X2=1.05 $Y2=1.78
cc_5 VNB A 0.0555865f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.21
cc_6 VNB N_A_c_70_n 0.0267173f $X=-0.19 $Y=-0.245 $X2=0.99 $Y2=1.275
cc_7 VNB N_A_303_300#_c_100_n 0.0110002f $X=-0.19 $Y=-0.245 $X2=1.15 $Y2=2.54
cc_8 VNB N_A_303_300#_M1008_g 0.00157364f $X=-0.19 $Y=-0.245 $X2=1.26 $Y2=1.11
cc_9 VNB N_A_303_300#_M1005_g 0.0286173f $X=-0.19 $Y=-0.245 $X2=1.05 $Y2=1.26
cc_10 VNB N_A_303_300#_c_103_n 0.00568422f $X=-0.19 $Y=-0.245 $X2=1.05 $Y2=1.78
cc_11 VNB N_A_303_300#_M1002_g 0.0336767f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_303_300#_c_105_n 0.00740747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_303_300#_c_106_n 0.00451996f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_303_300#_c_107_n 0.0132783f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_303_300#_c_108_n 0.00493453f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_303_300#_c_109_n 0.0224314f $X=-0.19 $Y=-0.245 $X2=1.05 $Y2=1.275
cc_17 VNB N_A_303_300#_c_110_n 0.00996019f $X=-0.19 $Y=-0.245 $X2=0.99 $Y2=1.275
cc_18 VNB N_A_303_300#_c_111_n 0.00271145f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.445
cc_19 VNB N_A_303_300#_c_112_n 0.024197f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_303_300#_c_113_n 0.0134429f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_303_300#_c_114_n 0.0309089f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_B_N_c_189_n 0.0138887f $X=-0.19 $Y=-0.245 $X2=0.9 $Y2=1.11
cc_23 VNB N_B_N_c_190_n 0.022028f $X=-0.19 $Y=-0.245 $X2=1.15 $Y2=1.78
cc_24 VNB N_B_N_c_191_n 0.00671294f $X=-0.19 $Y=-0.245 $X2=1.15 $Y2=2.54
cc_25 VNB N_B_N_c_192_n 0.00879792f $X=-0.19 $Y=-0.245 $X2=1.15 $Y2=2.54
cc_26 VNB N_B_N_c_193_n 0.0175316f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_B_N_c_194_n 0.00664349f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_28 VNB B_N 0.00479613f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_B_N_c_196_n 0.0164456f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_B_N_c_197_n 0.0133507f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VPWR_c_238_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB Y 0.0119793f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_Y_c_268_n 0.0115611f $X=-0.19 $Y=-0.245 $X2=0.99 $Y2=1.445
cc_34 VNB N_VGND_c_305_n 0.0261127f $X=-0.19 $Y=-0.245 $X2=1.26 $Y2=1.11
cc_35 VNB N_VGND_c_306_n 0.00177638f $X=-0.19 $Y=-0.245 $X2=1.05 $Y2=1.26
cc_36 VNB N_VGND_c_307_n 0.0186907f $X=-0.19 $Y=-0.245 $X2=1.05 $Y2=1.78
cc_37 VNB N_VGND_c_308_n 0.0338226f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.21
cc_38 VNB N_VGND_c_309_n 0.027948f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_310_n 0.2296f $X=-0.19 $Y=-0.245 $X2=1.05 $Y2=1.275
cc_40 VNB N_VGND_c_311_n 0.00551342f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.445
cc_41 VNB N_VGND_c_312_n 0.00500486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VPB N_A_M1004_g 0.0411747f $X=-0.19 $Y=1.655 $X2=1.15 $Y2=2.54
cc_43 VPB N_A_c_68_n 0.0164184f $X=-0.19 $Y=1.655 $X2=1.05 $Y2=1.78
cc_44 VPB A 0.0352665f $X=-0.19 $Y=1.655 $X2=1.115 $Y2=1.21
cc_45 VPB N_A_303_300#_M1008_g 0.0425515f $X=-0.19 $Y=1.655 $X2=1.26 $Y2=1.11
cc_46 VPB N_A_303_300#_c_108_n 0.0104598f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_47 VPB N_A_303_300#_c_109_n 0.0217862f $X=-0.19 $Y=1.655 $X2=1.05 $Y2=1.275
cc_48 VPB N_A_303_300#_c_118_n 0.0356992f $X=-0.19 $Y=1.655 $X2=0.99 $Y2=1.445
cc_49 VPB N_A_303_300#_c_119_n 0.0121631f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_50 VPB N_A_303_300#_c_114_n 0.0173944f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_51 VPB N_B_N_M1003_g 0.0406711f $X=-0.19 $Y=1.655 $X2=1.26 $Y2=0.495
cc_52 VPB N_B_N_c_199_n 0.0173713f $X=-0.19 $Y=1.655 $X2=1.05 $Y2=1.78
cc_53 VPB B_N 0.00276702f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_54 VPB N_VPWR_c_239_n 0.0469519f $X=-0.19 $Y=1.655 $X2=1.26 $Y2=0.495
cc_55 VPB N_VPWR_c_240_n 0.0221146f $X=-0.19 $Y=1.655 $X2=1.05 $Y2=1.78
cc_56 VPB N_VPWR_c_241_n 0.0363431f $X=-0.19 $Y=1.655 $X2=1.115 $Y2=1.21
cc_57 VPB N_VPWR_c_242_n 0.00548753f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_58 VPB N_VPWR_c_243_n 0.0196743f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_59 VPB N_VPWR_c_238_n 0.0975956f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_60 VPB N_VPWR_c_245_n 0.0305806f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_61 VPB Y 0.00752403f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_62 VPB Y 0.0101394f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_63 VPB Y 0.009877f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_64 A N_A_303_300#_c_100_n 0.00199926f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_65 N_A_c_70_n N_A_303_300#_c_100_n 0.0447229f $X=0.99 $Y=1.275 $X2=0 $Y2=0
cc_66 N_A_c_68_n N_A_303_300#_M1008_g 0.0447229f $X=1.05 $Y=1.78 $X2=0 $Y2=0
cc_67 N_A_M1001_g N_A_303_300#_M1005_g 0.0156127f $X=1.26 $Y=0.495 $X2=0 $Y2=0
cc_68 N_A_c_67_n N_A_303_300#_c_106_n 0.0156127f $X=1.08 $Y=1.26 $X2=0 $Y2=0
cc_69 A N_A_303_300#_c_106_n 9.85401e-19 $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_70 N_A_c_70_n N_A_303_300#_c_106_n 0.00838854f $X=0.99 $Y=1.275 $X2=0 $Y2=0
cc_71 N_A_M1004_g N_VPWR_c_239_n 0.0265299f $X=1.15 $Y=2.54 $X2=0 $Y2=0
cc_72 N_A_c_68_n N_VPWR_c_239_n 0.00521822f $X=1.05 $Y=1.78 $X2=0 $Y2=0
cc_73 A N_VPWR_c_239_n 0.0228311f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_74 N_A_M1004_g N_VPWR_c_241_n 0.00795364f $X=1.15 $Y=2.54 $X2=0 $Y2=0
cc_75 N_A_M1004_g N_VPWR_c_238_n 0.0142467f $X=1.15 $Y=2.54 $X2=0 $Y2=0
cc_76 N_A_M1001_g Y 0.00888454f $X=1.26 $Y=0.495 $X2=0 $Y2=0
cc_77 N_A_c_68_n Y 0.00262691f $X=1.05 $Y=1.78 $X2=0 $Y2=0
cc_78 A Y 0.0420964f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_79 N_A_c_70_n Y 0.00111773f $X=0.99 $Y=1.275 $X2=0 $Y2=0
cc_80 N_A_M1000_g N_Y_c_268_n 0.0012483f $X=0.9 $Y=0.495 $X2=0 $Y2=0
cc_81 N_A_M1001_g N_Y_c_268_n 0.00927375f $X=1.26 $Y=0.495 $X2=0 $Y2=0
cc_82 N_A_M1004_g Y 0.00262691f $X=1.15 $Y=2.54 $X2=0 $Y2=0
cc_83 N_A_M1000_g N_VGND_c_305_n 0.0142556f $X=0.9 $Y=0.495 $X2=0 $Y2=0
cc_84 N_A_M1001_g N_VGND_c_305_n 0.002112f $X=1.26 $Y=0.495 $X2=0 $Y2=0
cc_85 A N_VGND_c_305_n 0.0171088f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_86 N_A_M1000_g N_VGND_c_308_n 0.00445056f $X=0.9 $Y=0.495 $X2=0 $Y2=0
cc_87 N_A_M1001_g N_VGND_c_308_n 0.00502664f $X=1.26 $Y=0.495 $X2=0 $Y2=0
cc_88 N_A_M1000_g N_VGND_c_310_n 0.00796275f $X=0.9 $Y=0.495 $X2=0 $Y2=0
cc_89 N_A_M1001_g N_VGND_c_310_n 0.00942073f $X=1.26 $Y=0.495 $X2=0 $Y2=0
cc_90 N_A_303_300#_M1002_g N_B_N_c_189_n 0.0190851f $X=2.05 $Y=0.495 $X2=-0.19
+ $Y2=-0.245
cc_91 N_A_303_300#_c_112_n N_B_N_c_189_n 0.00170611f $X=3.055 $Y=0.495 $X2=-0.19
+ $Y2=-0.245
cc_92 N_A_303_300#_c_109_n N_B_N_c_190_n 0.0178703f $X=2.14 $Y=1.335 $X2=0 $Y2=0
cc_93 N_A_303_300#_c_110_n N_B_N_c_191_n 0.00773222f $X=2.89 $Y=0.91 $X2=0 $Y2=0
cc_94 N_A_303_300#_c_110_n N_B_N_c_192_n 0.00813947f $X=2.89 $Y=0.91 $X2=0 $Y2=0
cc_95 N_A_303_300#_c_118_n N_B_N_M1003_g 0.0158472f $X=3.055 $Y=2.9 $X2=0 $Y2=0
cc_96 N_A_303_300#_c_119_n N_B_N_M1003_g 0.00455769f $X=3.055 $Y=2.19 $X2=0
+ $Y2=0
cc_97 N_A_303_300#_c_112_n N_B_N_c_193_n 0.0110823f $X=3.055 $Y=0.495 $X2=0
+ $Y2=0
cc_98 N_A_303_300#_c_110_n N_B_N_c_194_n 0.00407103f $X=2.89 $Y=0.91 $X2=0 $Y2=0
cc_99 N_A_303_300#_c_112_n N_B_N_c_194_n 0.00296864f $X=3.055 $Y=0.495 $X2=0
+ $Y2=0
cc_100 N_A_303_300#_c_113_n N_B_N_c_194_n 0.00237652f $X=3.057 $Y=0.91 $X2=0
+ $Y2=0
cc_101 N_A_303_300#_c_107_n B_N 0.00415842f $X=2.14 $Y=1.245 $X2=0 $Y2=0
cc_102 N_A_303_300#_c_108_n B_N 0.0435845f $X=2.14 $Y=1.335 $X2=0 $Y2=0
cc_103 N_A_303_300#_c_110_n B_N 0.0262713f $X=2.89 $Y=0.91 $X2=0 $Y2=0
cc_104 N_A_303_300#_c_114_n B_N 0.0483743f $X=3.057 $Y=2.025 $X2=0 $Y2=0
cc_105 N_A_303_300#_c_107_n N_B_N_c_196_n 0.0178703f $X=2.14 $Y=1.245 $X2=0
+ $Y2=0
cc_106 N_A_303_300#_c_108_n N_B_N_c_196_n 8.16483e-19 $X=2.14 $Y=1.335 $X2=0
+ $Y2=0
cc_107 N_A_303_300#_c_110_n N_B_N_c_196_n 6.72787e-19 $X=2.89 $Y=0.91 $X2=0
+ $Y2=0
cc_108 N_A_303_300#_M1002_g N_B_N_c_197_n 7.8689e-19 $X=2.05 $Y=0.495 $X2=0
+ $Y2=0
cc_109 N_A_303_300#_c_108_n N_B_N_c_197_n 0.0012301f $X=2.14 $Y=1.335 $X2=0
+ $Y2=0
cc_110 N_A_303_300#_c_110_n N_B_N_c_197_n 0.0029312f $X=2.89 $Y=0.91 $X2=0 $Y2=0
cc_111 N_A_303_300#_c_113_n N_B_N_c_197_n 0.00274643f $X=3.057 $Y=0.91 $X2=0
+ $Y2=0
cc_112 N_A_303_300#_c_114_n N_B_N_c_197_n 0.0260795f $X=3.057 $Y=2.025 $X2=0
+ $Y2=0
cc_113 N_A_303_300#_M1008_g N_VPWR_c_239_n 0.00334008f $X=1.64 $Y=2.54 $X2=0
+ $Y2=0
cc_114 N_A_303_300#_M1008_g N_VPWR_c_240_n 0.0038838f $X=1.64 $Y=2.54 $X2=0
+ $Y2=0
cc_115 N_A_303_300#_c_119_n N_VPWR_c_240_n 0.0685723f $X=3.055 $Y=2.19 $X2=0
+ $Y2=0
cc_116 N_A_303_300#_M1008_g N_VPWR_c_241_n 0.00612332f $X=1.64 $Y=2.54 $X2=0
+ $Y2=0
cc_117 N_A_303_300#_c_118_n N_VPWR_c_243_n 0.0223692f $X=3.055 $Y=2.9 $X2=0
+ $Y2=0
cc_118 N_A_303_300#_M1008_g N_VPWR_c_238_n 0.0100408f $X=1.64 $Y=2.54 $X2=0
+ $Y2=0
cc_119 N_A_303_300#_c_118_n N_VPWR_c_238_n 0.0127743f $X=3.055 $Y=2.9 $X2=0
+ $Y2=0
cc_120 N_A_303_300#_c_100_n Y 0.00478542f $X=1.64 $Y=1.625 $X2=0 $Y2=0
cc_121 N_A_303_300#_M1008_g Y 0.0148301f $X=1.64 $Y=2.54 $X2=0 $Y2=0
cc_122 N_A_303_300#_M1005_g Y 0.00919972f $X=1.69 $Y=0.495 $X2=0 $Y2=0
cc_123 N_A_303_300#_c_103_n Y 0.00253815f $X=1.975 $Y=1.245 $X2=0 $Y2=0
cc_124 N_A_303_300#_M1002_g Y 0.00139845f $X=2.05 $Y=0.495 $X2=0 $Y2=0
cc_125 N_A_303_300#_c_105_n Y 0.00393291f $X=1.64 $Y=1.5 $X2=0 $Y2=0
cc_126 N_A_303_300#_c_106_n Y 0.00287871f $X=1.69 $Y=1.245 $X2=0 $Y2=0
cc_127 N_A_303_300#_c_108_n Y 0.0615677f $X=2.14 $Y=1.335 $X2=0 $Y2=0
cc_128 N_A_303_300#_c_109_n Y 0.00283088f $X=2.14 $Y=1.335 $X2=0 $Y2=0
cc_129 N_A_303_300#_c_111_n Y 0.0132974f $X=2.305 $Y=0.91 $X2=0 $Y2=0
cc_130 N_A_303_300#_M1008_g Y 0.0266734f $X=1.64 $Y=2.54 $X2=0 $Y2=0
cc_131 N_A_303_300#_M1005_g N_Y_c_268_n 0.0094252f $X=1.69 $Y=0.495 $X2=0 $Y2=0
cc_132 N_A_303_300#_M1002_g N_Y_c_268_n 0.003736f $X=2.05 $Y=0.495 $X2=0 $Y2=0
cc_133 N_A_303_300#_M1008_g Y 0.00829597f $X=1.64 $Y=2.54 $X2=0 $Y2=0
cc_134 N_A_303_300#_c_103_n Y 7.15443e-19 $X=1.975 $Y=1.245 $X2=0 $Y2=0
cc_135 N_A_303_300#_c_108_n Y 0.00793874f $X=2.14 $Y=1.335 $X2=0 $Y2=0
cc_136 N_A_303_300#_c_109_n Y 7.22101e-19 $X=2.14 $Y=1.335 $X2=0 $Y2=0
cc_137 N_A_303_300#_M1005_g N_VGND_c_306_n 0.00124485f $X=1.69 $Y=0.495 $X2=0
+ $Y2=0
cc_138 N_A_303_300#_M1002_g N_VGND_c_306_n 0.00951264f $X=2.05 $Y=0.495 $X2=0
+ $Y2=0
cc_139 N_A_303_300#_c_107_n N_VGND_c_306_n 5.87721e-19 $X=2.14 $Y=1.245 $X2=0
+ $Y2=0
cc_140 N_A_303_300#_c_110_n N_VGND_c_306_n 0.00688243f $X=2.89 $Y=0.91 $X2=0
+ $Y2=0
cc_141 N_A_303_300#_c_111_n N_VGND_c_306_n 0.0147604f $X=2.305 $Y=0.91 $X2=0
+ $Y2=0
cc_142 N_A_303_300#_c_112_n N_VGND_c_306_n 0.0127284f $X=3.055 $Y=0.495 $X2=0
+ $Y2=0
cc_143 N_A_303_300#_M1005_g N_VGND_c_308_n 0.00327544f $X=1.69 $Y=0.495 $X2=0
+ $Y2=0
cc_144 N_A_303_300#_M1002_g N_VGND_c_308_n 0.00445056f $X=2.05 $Y=0.495 $X2=0
+ $Y2=0
cc_145 N_A_303_300#_c_112_n N_VGND_c_309_n 0.0223692f $X=3.055 $Y=0.495 $X2=0
+ $Y2=0
cc_146 N_A_303_300#_M1005_g N_VGND_c_310_n 0.00475249f $X=1.69 $Y=0.495 $X2=0
+ $Y2=0
cc_147 N_A_303_300#_M1002_g N_VGND_c_310_n 0.0041935f $X=2.05 $Y=0.495 $X2=0
+ $Y2=0
cc_148 N_A_303_300#_c_110_n N_VGND_c_310_n 0.0139938f $X=2.89 $Y=0.91 $X2=0
+ $Y2=0
cc_149 N_A_303_300#_c_111_n N_VGND_c_310_n 0.00483194f $X=2.305 $Y=0.91 $X2=0
+ $Y2=0
cc_150 N_A_303_300#_c_112_n N_VGND_c_310_n 0.0127743f $X=3.055 $Y=0.495 $X2=0
+ $Y2=0
cc_151 N_B_N_M1003_g N_VPWR_c_240_n 0.0249766f $X=2.79 $Y=2.545 $X2=0 $Y2=0
cc_152 N_B_N_c_199_n N_VPWR_c_240_n 9.32746e-19 $X=2.73 $Y=1.845 $X2=0 $Y2=0
cc_153 B_N N_VPWR_c_240_n 0.0138772f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_154 N_B_N_M1003_g N_VPWR_c_243_n 0.00769046f $X=2.79 $Y=2.545 $X2=0 $Y2=0
cc_155 N_B_N_M1003_g N_VPWR_c_238_n 0.0140999f $X=2.79 $Y=2.545 $X2=0 $Y2=0
cc_156 N_B_N_M1003_g Y 0.00241917f $X=2.79 $Y=2.545 $X2=0 $Y2=0
cc_157 N_B_N_c_189_n N_VGND_c_306_n 0.0106455f $X=2.48 $Y=0.78 $X2=0 $Y2=0
cc_158 N_B_N_c_193_n N_VGND_c_306_n 0.00189426f $X=2.84 $Y=0.78 $X2=0 $Y2=0
cc_159 N_B_N_c_189_n N_VGND_c_309_n 0.00445056f $X=2.48 $Y=0.78 $X2=0 $Y2=0
cc_160 N_B_N_c_191_n N_VGND_c_309_n 4.57848e-19 $X=2.765 $Y=0.855 $X2=0 $Y2=0
cc_161 N_B_N_c_193_n N_VGND_c_309_n 0.00502664f $X=2.84 $Y=0.78 $X2=0 $Y2=0
cc_162 N_B_N_c_189_n N_VGND_c_310_n 0.0041956f $X=2.48 $Y=0.78 $X2=0 $Y2=0
cc_163 N_B_N_c_191_n N_VGND_c_310_n 6.33118e-19 $X=2.765 $Y=0.855 $X2=0 $Y2=0
cc_164 N_B_N_c_193_n N_VGND_c_310_n 0.00629305f $X=2.84 $Y=0.78 $X2=0 $Y2=0
cc_165 N_VPWR_c_241_n Y 0.0322497f $X=2.36 $Y=3.33 $X2=0 $Y2=0
cc_166 N_VPWR_c_238_n Y 0.0184956f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_167 N_VPWR_c_239_n Y 0.0325819f $X=0.885 $Y=2.185 $X2=0 $Y2=0
cc_168 N_VPWR_c_240_n Y 0.0614387f $X=2.525 $Y=2.19 $X2=0 $Y2=0
cc_169 N_Y_c_268_n N_VGND_c_305_n 0.0158572f $X=1.475 $Y=0.495 $X2=0 $Y2=0
cc_170 N_Y_c_268_n N_VGND_c_306_n 0.00949156f $X=1.475 $Y=0.495 $X2=0 $Y2=0
cc_171 N_Y_c_268_n N_VGND_c_308_n 0.0314759f $X=1.475 $Y=0.495 $X2=0 $Y2=0
cc_172 N_Y_c_268_n N_VGND_c_310_n 0.0177861f $X=1.475 $Y=0.495 $X2=0 $Y2=0
