* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__dfbbn_1 CLK_N D RESET_B SET_B VGND VNB VPB VPWR Q Q_N
X0 a_1013_66# a_546_449# a_755_398# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X1 a_1741_137# a_1531_428# a_2036_451# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X2 a_702_110# a_755_398# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 VGND a_2511_137# Q VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X4 a_1693_163# a_1741_137# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 a_1741_137# a_1186_21# a_1896_119# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X6 VPWR CLK_N a_113_67# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X7 a_707_449# a_755_398# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X8 VGND a_1741_137# Q_N VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X9 VPWR SET_B a_1741_137# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X10 a_2511_137# a_1741_137# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X11 a_223_119# a_113_67# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X12 a_223_119# a_113_67# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X13 a_1442_119# a_113_67# a_1531_428# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X14 a_2511_137# a_1741_137# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X15 a_1649_512# a_1741_137# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X16 a_1228_379# a_1186_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X17 VPWR a_755_398# a_1436_379# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X18 VGND a_755_398# a_1442_119# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X19 a_1436_379# a_223_119# a_1531_428# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X20 a_1186_21# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X21 a_1896_119# a_1531_428# a_1741_137# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X22 a_2036_451# a_1186_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X23 a_1531_428# a_113_67# a_1649_512# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X24 VGND D a_460_449# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X25 a_546_449# a_223_119# a_707_449# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X26 VGND SET_B a_1013_66# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X27 a_460_449# a_113_67# a_546_449# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X28 VPWR SET_B a_755_398# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X29 a_755_398# a_1186_21# a_1013_66# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X30 VPWR D a_460_449# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X31 a_1186_21# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X32 VGND CLK_N a_113_67# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X33 VPWR a_1741_137# Q_N VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X34 a_755_398# a_546_449# a_1228_379# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X35 a_460_449# a_223_119# a_546_449# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X36 VPWR a_2511_137# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X37 a_1531_428# a_223_119# a_1693_163# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X38 a_546_449# a_113_67# a_702_110# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X39 VGND SET_B a_1896_119# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
.ends
