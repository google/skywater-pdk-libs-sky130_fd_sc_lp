* File: sky130_fd_sc_lp__o31a_1.spice
* Created: Wed Sep  2 10:24:29 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__o31a_1.pex.spice"
.subckt sky130_fd_sc_lp__o31a_1  VNB VPB A1 A2 A3 B1 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* B1	B1
* A3	A3
* A2	A2
* A1	A1
* VPB	VPB
* VNB	VNB
MM1005 N_VGND_M1005_d N_A_86_23#_M1005_g N_X_M1005_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2709 AS=0.2226 PD=1.485 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75002.4 A=0.126 P=1.98 MULT=1
MM1002 N_A_275_49#_M1002_d N_A1_M1002_g N_VGND_M1005_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1281 AS=0.2709 PD=1.145 PS=1.485 NRD=3.564 NRS=0 M=1 R=5.6 SA=75001
+ SB=75001.6 A=0.126 P=1.98 MULT=1
MM1000 N_VGND_M1000_d N_A2_M1000_g N_A_275_49#_M1002_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1701 AS=0.1281 PD=1.245 PS=1.145 NRD=9.276 NRS=0 M=1 R=5.6 SA=75001.4
+ SB=75001.2 A=0.126 P=1.98 MULT=1
MM1004 N_A_275_49#_M1004_d N_A3_M1004_g N_VGND_M1000_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1701 PD=1.12 PS=1.245 NRD=0 NRS=8.568 M=1 R=5.6 SA=75002
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1008 N_A_86_23#_M1008_d N_B1_M1008_g N_A_275_49#_M1004_d VNB NSHORT L=0.15
+ W=0.84 AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002.4
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1003 N_VPWR_M1003_d N_A_86_23#_M1003_g N_X_M1003_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.40635 AS=0.3339 PD=1.905 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75002.4 A=0.189 P=2.82 MULT=1
MM1007 A_275_367# N_A1_M1007_g N_VPWR_M1003_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1953 AS=0.40635 PD=1.57 PS=1.905 NRD=15.6221 NRS=0 M=1 R=8.4 SA=75001
+ SB=75001.6 A=0.189 P=2.82 MULT=1
MM1009 A_367_367# N_A2_M1009_g A_275_367# VPB PHIGHVT L=0.15 W=1.26 AD=0.1827
+ AS=0.1953 PD=1.55 PS=1.57 NRD=14.0658 NRS=15.6221 M=1 R=8.4 SA=75001.4
+ SB=75001.2 A=0.189 P=2.82 MULT=1
MM1001 N_A_86_23#_M1001_d N_A3_M1001_g A_367_367# VPB PHIGHVT L=0.15 W=1.26
+ AD=0.2457 AS=0.1827 PD=1.65 PS=1.55 NRD=6.2449 NRS=14.0658 M=1 R=8.4
+ SA=75001.9 SB=75000.7 A=0.189 P=2.82 MULT=1
MM1006 N_VPWR_M1006_d N_B1_M1006_g N_A_86_23#_M1001_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.2457 PD=3.05 PS=1.65 NRD=0 NRS=10.9335 M=1 R=8.4 SA=75002.4
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9751 P=11.21
*
.include "sky130_fd_sc_lp__o31a_1.pxi.spice"
*
.ends
*
*
