* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__ha_0 A B VGND VNB VPB VPWR COUT SUM
M1000 VPWR a_80_60# SUM VPB phighvt w=640000u l=150000u
+  ad=7.804e+11p pd=6.54e+06u as=1.824e+11p ps=1.85e+06u
M1001 a_393_491# B a_80_60# VPB phighvt w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=2.709e+11p ps=2.13e+06u
M1002 a_687_135# B a_204_315# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=1.239e+11p ps=1.43e+06u
M1003 VGND a_80_60# SUM VNB nshort w=420000u l=150000u
+  ad=4.2e+11p pd=4.52e+06u as=1.113e+11p ps=1.37e+06u
M1004 VGND B a_307_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=2.289e+11p ps=2.77e+06u
M1005 VPWR A a_393_491# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR A a_204_315# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.176e+11p ps=1.4e+06u
M1007 COUT a_204_315# VGND VNB nshort w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1008 a_80_60# a_204_315# VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 COUT a_204_315# VPWR VPB phighvt w=640000u l=150000u
+  ad=1.696e+11p pd=1.81e+06u as=0p ps=0u
M1010 a_204_315# B VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND A a_687_135# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_307_47# A VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_307_47# a_204_315# a_80_60# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
.ends
