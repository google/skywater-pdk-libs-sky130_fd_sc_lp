* File: sky130_fd_sc_lp__a2bb2o_2.pex.spice
* Created: Wed Sep  2 09:23:49 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A2BB2O_2%B1 3 5 7 8 9 10 17
c25 8 0 1.80367e-19 $X=0.24 $Y=1.295
r26 15 17 35.5432 $w=2.78e-07 $l=2.05e-07 $layer=POLY_cond $X=0.27 $Y=1.35
+ $X2=0.475 $Y2=1.35
r27 9 10 13.755 $w=3.08e-07 $l=3.7e-07 $layer=LI1_cond $X=0.24 $Y=1.665 $X2=0.24
+ $Y2=2.035
r28 8 9 13.755 $w=3.08e-07 $l=3.7e-07 $layer=LI1_cond $X=0.24 $Y=1.295 $X2=0.24
+ $Y2=1.665
r29 8 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=1.35 $X2=0.27 $Y2=1.35
r30 5 17 31.2086 $w=2.78e-07 $l=2.49199e-07 $layer=POLY_cond $X=0.655 $Y=1.185
+ $X2=0.475 $Y2=1.35
r31 5 7 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.655 $Y=1.185
+ $X2=0.655 $Y2=0.865
r32 1 17 17.1848 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=1.515
+ $X2=0.475 $Y2=1.35
r33 1 3 620.447 $w=1.5e-07 $l=1.21e-06 $layer=POLY_cond $X=0.475 $Y=1.515
+ $X2=0.475 $Y2=2.725
.ends

.subckt PM_SKY130_FD_SC_LP__A2BB2O_2%B2 3 7 11 12 13 14 15 20
c35 7 0 1.80367e-19 $X=1.015 $Y=0.865
c36 3 0 1.50287e-19 $X=0.945 $Y=2.725
r37 20 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.925
+ $Y=1.71 $X2=0.925 $Y2=1.71
r38 15 21 8.54342 $w=4.53e-07 $l=3.25e-07 $layer=LI1_cond $X=0.792 $Y=2.035
+ $X2=0.792 $Y2=1.71
r39 14 21 1.18293 $w=4.53e-07 $l=4.5e-08 $layer=LI1_cond $X=0.792 $Y=1.665
+ $X2=0.792 $Y2=1.71
r40 13 14 9.72635 $w=4.53e-07 $l=3.7e-07 $layer=LI1_cond $X=0.792 $Y=1.295
+ $X2=0.792 $Y2=1.665
r41 11 20 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.925 $Y=2.05
+ $X2=0.925 $Y2=1.71
r42 11 12 38.6168 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.925 $Y=2.05
+ $X2=0.925 $Y2=2.215
r43 10 20 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.925 $Y=1.545
+ $X2=0.925 $Y2=1.71
r44 7 10 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=1.015 $Y=0.865
+ $X2=1.015 $Y2=1.545
r45 3 12 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=0.945 $Y=2.725
+ $X2=0.945 $Y2=2.215
.ends

.subckt PM_SKY130_FD_SC_LP__A2BB2O_2%A_260_341# 1 2 9 13 16 17 19 21 22 23 24 29
+ 34
c59 17 0 1.93085e-19 $X=1.545 $Y=1.855
c60 9 0 1.73044e-19 $X=1.375 $Y=2.725
r61 29 31 4.22511 $w=2.08e-07 $l=8e-08 $layer=LI1_cond $X=2.52 $Y=0.865 $X2=2.52
+ $Y2=0.945
r62 23 31 1.9771 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=2.415 $Y=0.945
+ $X2=2.52 $Y2=0.945
r63 23 24 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=2.415 $Y=0.945
+ $X2=1.79 $Y2=0.945
r64 22 34 46.1517 $w=4.2e-07 $l=1.65e-07 $layer=POLY_cond $X=1.58 $Y=1.35
+ $X2=1.58 $Y2=1.185
r65 21 22 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.625
+ $Y=1.35 $X2=1.625 $Y2=1.35
r66 19 27 18.866 $w=2.91e-07 $l=5.83652e-07 $layer=LI1_cond $X=1.66 $Y=1.685
+ $X2=2.11 $Y2=1.992
r67 19 21 14.8488 $w=2.58e-07 $l=3.35e-07 $layer=LI1_cond $X=1.66 $Y=1.685
+ $X2=1.66 $Y2=1.35
r68 18 24 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=1.66 $Y=1.03
+ $X2=1.79 $Y2=0.945
r69 18 21 14.1839 $w=2.58e-07 $l=3.2e-07 $layer=LI1_cond $X=1.66 $Y=1.03
+ $X2=1.66 $Y2=1.35
r70 16 17 44.1654 $w=4.2e-07 $l=1.5e-07 $layer=POLY_cond $X=1.545 $Y=1.705
+ $X2=1.545 $Y2=1.855
r71 14 22 5.95879 $w=4.2e-07 $l=4.5e-08 $layer=POLY_cond $X=1.58 $Y=1.395
+ $X2=1.58 $Y2=1.35
r72 14 16 41.0494 $w=4.2e-07 $l=3.1e-07 $layer=POLY_cond $X=1.58 $Y=1.395
+ $X2=1.58 $Y2=1.705
r73 13 34 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.445 $Y=0.865
+ $X2=1.445 $Y2=1.185
r74 9 17 446.106 $w=1.5e-07 $l=8.7e-07 $layer=POLY_cond $X=1.375 $Y=2.725
+ $X2=1.375 $Y2=1.855
r75 2 27 600 $w=1.7e-07 $l=2.23942e-07 $layer=licon1_PDIFF $count=1 $X=1.985
+ $Y=1.835 $X2=2.11 $Y2=2.005
r76 1 29 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.38
+ $Y=0.655 $X2=2.52 $Y2=0.865
.ends

.subckt PM_SKY130_FD_SC_LP__A2BB2O_2%A2_N 1 3 4 6 8
r33 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.21
+ $Y=1.35 $X2=2.21 $Y2=1.35
r34 4 11 38.7185 $w=3.44e-07 $l=2.10286e-07 $layer=POLY_cond $X=2.325 $Y=1.515
+ $X2=2.222 $Y2=1.35
r35 4 6 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=2.325 $Y=1.515
+ $X2=2.325 $Y2=2.155
r36 1 11 38.7185 $w=3.44e-07 $l=2.02287e-07 $layer=POLY_cond $X=2.305 $Y=1.185
+ $X2=2.222 $Y2=1.35
r37 1 3 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.305 $Y=1.185
+ $X2=2.305 $Y2=0.865
.ends

.subckt PM_SKY130_FD_SC_LP__A2BB2O_2%A1_N 3 7 9 10 11 16
c37 16 0 3.61887e-20 $X=2.775 $Y=1.375
r38 16 19 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.775 $Y=1.375
+ $X2=2.775 $Y2=1.54
r39 16 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.775 $Y=1.375
+ $X2=2.775 $Y2=1.21
r40 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.775
+ $Y=1.375 $X2=2.775 $Y2=1.375
r41 10 11 13.1201 $w=3.23e-07 $l=3.7e-07 $layer=LI1_cond $X=2.707 $Y=1.665
+ $X2=2.707 $Y2=2.035
r42 10 17 10.2833 $w=3.23e-07 $l=2.9e-07 $layer=LI1_cond $X=2.707 $Y=1.665
+ $X2=2.707 $Y2=1.375
r43 9 17 2.83678 $w=3.23e-07 $l=8e-08 $layer=LI1_cond $X=2.707 $Y=1.295
+ $X2=2.707 $Y2=1.375
r44 7 18 176.904 $w=1.5e-07 $l=3.45e-07 $layer=POLY_cond $X=2.735 $Y=0.865
+ $X2=2.735 $Y2=1.21
r45 3 19 315.351 $w=1.5e-07 $l=6.15e-07 $layer=POLY_cond $X=2.685 $Y=2.155
+ $X2=2.685 $Y2=1.54
.ends

.subckt PM_SKY130_FD_SC_LP__A2BB2O_2%A_218_131# 1 2 9 13 17 21 24 27 29 30 32 34
+ 42 48
c91 29 0 1.93085e-19 $X=3.04 $Y=2.385
r92 43 48 65.573 $w=3.3e-07 $l=3.75e-07 $layer=POLY_cond $X=3.315 $Y=1.505
+ $X2=3.69 $Y2=1.505
r93 43 45 9.61737 $w=3.3e-07 $l=5.5e-08 $layer=POLY_cond $X=3.315 $Y=1.505
+ $X2=3.26 $Y2=1.505
r94 42 43 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.315
+ $Y=1.505 $X2=3.315 $Y2=1.505
r95 39 42 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=3.125 $Y=1.505
+ $X2=3.315 $Y2=1.505
r96 34 36 8.49766 $w=2.93e-07 $l=1.65e-07 $layer=LI1_cond $X=1.212 $Y=0.85
+ $X2=1.212 $Y2=1.015
r97 31 39 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.125 $Y=1.67
+ $X2=3.125 $Y2=1.505
r98 31 32 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=3.125 $Y=1.67
+ $X2=3.125 $Y2=2.3
r99 30 38 8.32986 $w=2.76e-07 $l=2.02109e-07 $layer=LI1_cond $X=1.755 $Y=2.385
+ $X2=1.607 $Y2=2.257
r100 29 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.04 $Y=2.385
+ $X2=3.125 $Y2=2.3
r101 29 30 83.8342 $w=1.68e-07 $l=1.285e-06 $layer=LI1_cond $X=3.04 $Y=2.385
+ $X2=1.755 $Y2=2.385
r102 25 38 0.328487 $w=2.95e-07 $l=2.13e-07 $layer=LI1_cond $X=1.607 $Y=2.47
+ $X2=1.607 $Y2=2.257
r103 25 27 3.12527 $w=2.93e-07 $l=8e-08 $layer=LI1_cond $X=1.607 $Y=2.47
+ $X2=1.607 $Y2=2.55
r104 24 38 14.6754 $w=2.76e-07 $l=4.2498e-07 $layer=LI1_cond $X=1.275 $Y=2.045
+ $X2=1.607 $Y2=2.257
r105 24 36 67.1979 $w=1.68e-07 $l=1.03e-06 $layer=LI1_cond $X=1.275 $Y=2.045
+ $X2=1.275 $Y2=1.015
r106 19 48 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.69 $Y=1.67
+ $X2=3.69 $Y2=1.505
r107 19 21 407.649 $w=1.5e-07 $l=7.95e-07 $layer=POLY_cond $X=3.69 $Y=1.67
+ $X2=3.69 $Y2=2.465
r108 15 48 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.69 $Y=1.34
+ $X2=3.69 $Y2=1.505
r109 15 17 351.245 $w=1.5e-07 $l=6.85e-07 $layer=POLY_cond $X=3.69 $Y=1.34
+ $X2=3.69 $Y2=0.655
r110 11 45 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.26 $Y=1.67
+ $X2=3.26 $Y2=1.505
r111 11 13 407.649 $w=1.5e-07 $l=7.95e-07 $layer=POLY_cond $X=3.26 $Y=1.67
+ $X2=3.26 $Y2=2.465
r112 7 45 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.26 $Y=1.34
+ $X2=3.26 $Y2=1.505
r113 7 9 351.245 $w=1.5e-07 $l=6.85e-07 $layer=POLY_cond $X=3.26 $Y=1.34
+ $X2=3.26 $Y2=0.655
r114 2 27 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=1.45
+ $Y=2.405 $X2=1.59 $Y2=2.55
r115 1 34 182 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_NDIFF $count=1 $X=1.09
+ $Y=0.655 $X2=1.23 $Y2=0.85
.ends

.subckt PM_SKY130_FD_SC_LP__A2BB2O_2%A_27_481# 1 2 9 13 16
c22 13 0 1.50287e-19 $X=1.16 $Y=2.56
c23 9 0 1.73044e-19 $X=1.055 $Y=2.47
r24 11 13 0.245201 $w=2.33e-07 $l=5e-09 $layer=LI1_cond $X=1.172 $Y=2.555
+ $X2=1.172 $Y2=2.56
r25 10 16 4.47015 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=0.365 $Y=2.47
+ $X2=0.23 $Y2=2.47
r26 9 11 7.04737 $w=1.7e-07 $l=1.53734e-07 $layer=LI1_cond $X=1.055 $Y=2.47
+ $X2=1.172 $Y2=2.555
r27 9 10 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.055 $Y=2.47
+ $X2=0.365 $Y2=2.47
r28 2 13 300 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_PDIFF $count=2 $X=1.02
+ $Y=2.405 $X2=1.16 $Y2=2.56
r29 1 16 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.405 $X2=0.26 $Y2=2.55
.ends

.subckt PM_SKY130_FD_SC_LP__A2BB2O_2%VPWR 1 2 3 12 16 18 20 24 26 31 39 45 48 52
r51 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r52 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r53 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r54 43 52 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r55 43 49 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=3.12 $Y2=3.33
r56 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r57 40 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.21 $Y=3.33
+ $X2=3.045 $Y2=3.33
r58 40 42 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=3.21 $Y=3.33 $X2=3.6
+ $Y2=3.33
r59 39 51 3.63491 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=3.91 $Y=3.33
+ $X2=4.115 $Y2=3.33
r60 39 42 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=3.91 $Y=3.33 $X2=3.6
+ $Y2=3.33
r61 38 49 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r62 37 38 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r63 35 46 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r64 34 37 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r65 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r66 32 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.875 $Y=3.33
+ $X2=0.71 $Y2=3.33
r67 32 34 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.875 $Y=3.33
+ $X2=1.2 $Y2=3.33
r68 31 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.88 $Y=3.33
+ $X2=3.045 $Y2=3.33
r69 31 37 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=2.88 $Y=3.33
+ $X2=2.64 $Y2=3.33
r70 29 46 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r71 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r72 26 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.545 $Y=3.33
+ $X2=0.71 $Y2=3.33
r73 26 28 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.545 $Y=3.33
+ $X2=0.24 $Y2=3.33
r74 24 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r75 24 35 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.2 $Y2=3.33
r76 20 23 51.2294 $w=2.08e-07 $l=9.7e-07 $layer=LI1_cond $X=4.015 $Y=1.98
+ $X2=4.015 $Y2=2.95
r77 18 51 3.28028 $w=2.1e-07 $l=1.36015e-07 $layer=LI1_cond $X=4.015 $Y=3.245
+ $X2=4.115 $Y2=3.33
r78 18 23 15.5801 $w=2.08e-07 $l=2.95e-07 $layer=LI1_cond $X=4.015 $Y=3.245
+ $X2=4.015 $Y2=2.95
r79 14 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.045 $Y=3.245
+ $X2=3.045 $Y2=3.33
r80 14 16 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=3.045 $Y=3.245
+ $X2=3.045 $Y2=2.78
r81 10 45 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.71 $Y=3.245
+ $X2=0.71 $Y2=3.33
r82 10 12 13.7944 $w=3.28e-07 $l=3.95e-07 $layer=LI1_cond $X=0.71 $Y=3.245
+ $X2=0.71 $Y2=2.85
r83 3 23 400 $w=1.7e-07 $l=1.22461e-06 $layer=licon1_PDIFF $count=1 $X=3.765
+ $Y=1.835 $X2=3.995 $Y2=2.95
r84 3 20 400 $w=1.7e-07 $l=2.93684e-07 $layer=licon1_PDIFF $count=1 $X=3.765
+ $Y=1.835 $X2=3.995 $Y2=1.98
r85 2 16 600 $w=1.7e-07 $l=1.07812e-06 $layer=licon1_PDIFF $count=1 $X=2.76
+ $Y=1.835 $X2=3.045 $Y2=2.78
r86 1 12 600 $w=1.7e-07 $l=5.18869e-07 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=2.405 $X2=0.71 $Y2=2.85
.ends

.subckt PM_SKY130_FD_SC_LP__A2BB2O_2%X 1 2 9 13 14 15 16 23 33
c27 33 0 3.61887e-20 $X=3.56 $Y=1.85
r28 21 35 0.480185 $w=3.58e-07 $l=1.5e-08 $layer=LI1_cond $X=3.56 $Y=2.03
+ $X2=3.56 $Y2=2.015
r29 21 23 0.160062 $w=3.58e-07 $l=5e-09 $layer=LI1_cond $X=3.56 $Y=2.03 $X2=3.56
+ $Y2=2.035
r30 16 30 4.32166 $w=3.58e-07 $l=1.35e-07 $layer=LI1_cond $X=3.56 $Y=2.775
+ $X2=3.56 $Y2=2.91
r31 15 16 11.8446 $w=3.58e-07 $l=3.7e-07 $layer=LI1_cond $X=3.56 $Y=2.405
+ $X2=3.56 $Y2=2.775
r32 14 35 0.800308 $w=3.58e-07 $l=2.5e-08 $layer=LI1_cond $X=3.56 $Y=1.99
+ $X2=3.56 $Y2=2.015
r33 14 33 7.71072 $w=3.58e-07 $l=1.4e-07 $layer=LI1_cond $X=3.56 $Y=1.99
+ $X2=3.56 $Y2=1.85
r34 14 15 10.5641 $w=3.58e-07 $l=3.3e-07 $layer=LI1_cond $X=3.56 $Y=2.075
+ $X2=3.56 $Y2=2.405
r35 14 23 1.28049 $w=3.58e-07 $l=4e-08 $layer=LI1_cond $X=3.56 $Y=2.075 $X2=3.56
+ $Y2=2.035
r36 13 33 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=3.655 $Y=1.095
+ $X2=3.655 $Y2=1.85
r37 7 13 9.16175 $w=3.68e-07 $l=1.85e-07 $layer=LI1_cond $X=3.555 $Y=0.91
+ $X2=3.555 $Y2=1.095
r38 7 9 15.2621 $w=3.68e-07 $l=4.9e-07 $layer=LI1_cond $X=3.555 $Y=0.91
+ $X2=3.555 $Y2=0.42
r39 2 35 400 $w=1.7e-07 $l=2.4e-07 $layer=licon1_PDIFF $count=1 $X=3.335
+ $Y=1.835 $X2=3.475 $Y2=2.015
r40 2 30 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=3.335
+ $Y=1.835 $X2=3.475 $Y2=2.91
r41 1 9 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=3.335
+ $Y=0.235 $X2=3.475 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__A2BB2O_2%VGND 1 2 3 4 15 19 23 25 27 30 31 33 34 35
+ 40 48 53 57
r55 56 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r56 53 54 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r57 51 57 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r58 50 51 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r59 48 56 3.63491 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=3.91 $Y=0 $X2=4.115
+ $Y2=0
r60 48 50 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=3.91 $Y=0 $X2=3.6
+ $Y2=0
r61 47 51 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r62 46 47 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r63 44 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.94 $Y=0 $X2=1.775
+ $Y2=0
r64 44 46 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=1.94 $Y=0 $X2=2.64
+ $Y2=0
r65 43 54 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r66 42 43 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r67 40 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.61 $Y=0 $X2=1.775
+ $Y2=0
r68 40 42 58.0642 $w=1.68e-07 $l=8.9e-07 $layer=LI1_cond $X=1.61 $Y=0 $X2=0.72
+ $Y2=0
r69 39 43 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r70 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r71 35 47 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r72 35 54 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.68
+ $Y2=0
r73 33 46 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=2.94 $Y=0 $X2=2.64
+ $Y2=0
r74 33 34 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.94 $Y=0 $X2=3.035
+ $Y2=0
r75 32 50 30.6631 $w=1.68e-07 $l=4.7e-07 $layer=LI1_cond $X=3.13 $Y=0 $X2=3.6
+ $Y2=0
r76 32 34 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=3.13 $Y=0 $X2=3.035
+ $Y2=0
r77 30 38 2.51176 $w=1.7e-07 $l=3.5e-08 $layer=LI1_cond $X=0.275 $Y=0 $X2=0.24
+ $Y2=0
r78 30 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.275 $Y=0 $X2=0.44
+ $Y2=0
r79 29 42 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=0.605 $Y=0 $X2=0.72
+ $Y2=0
r80 29 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.605 $Y=0 $X2=0.44
+ $Y2=0
r81 25 56 3.28028 $w=2.1e-07 $l=1.36015e-07 $layer=LI1_cond $X=4.015 $Y=0.085
+ $X2=4.115 $Y2=0
r82 25 27 15.5801 $w=2.08e-07 $l=2.95e-07 $layer=LI1_cond $X=4.015 $Y=0.085
+ $X2=4.015 $Y2=0.38
r83 21 34 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=3.035 $Y=0.085
+ $X2=3.035 $Y2=0
r84 21 23 17.2201 $w=1.88e-07 $l=2.95e-07 $layer=LI1_cond $X=3.035 $Y=0.085
+ $X2=3.035 $Y2=0.38
r85 17 53 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.775 $Y=0.085
+ $X2=1.775 $Y2=0
r86 17 19 17.8105 $w=3.28e-07 $l=5.1e-07 $layer=LI1_cond $X=1.775 $Y=0.085
+ $X2=1.775 $Y2=0.595
r87 13 31 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.44 $Y=0.085
+ $X2=0.44 $Y2=0
r88 13 15 27.2396 $w=3.28e-07 $l=7.8e-07 $layer=LI1_cond $X=0.44 $Y=0.085
+ $X2=0.44 $Y2=0.865
r89 4 27 91 $w=1.7e-07 $l=2.93684e-07 $layer=licon1_NDIFF $count=2 $X=3.765
+ $Y=0.235 $X2=3.995 $Y2=0.38
r90 3 23 91 $w=1.7e-07 $l=3.745e-07 $layer=licon1_NDIFF $count=2 $X=2.81
+ $Y=0.655 $X2=3.045 $Y2=0.38
r91 2 19 182 $w=1.7e-07 $l=2.83417e-07 $layer=licon1_NDIFF $count=1 $X=1.52
+ $Y=0.655 $X2=1.775 $Y2=0.595
r92 1 15 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.315
+ $Y=0.655 $X2=0.44 $Y2=0.865
.ends

