* File: sky130_fd_sc_lp__dlybuf4s15kapwr_2.pxi.spice
* Created: Fri Aug 28 10:29:36 2020
* 
x_PM_SKY130_FD_SC_LP__DLYBUF4S15KAPWR_2%A N_A_M1005_g N_A_M1009_g A A N_A_c_63_n
+ PM_SKY130_FD_SC_LP__DLYBUF4S15KAPWR_2%A
x_PM_SKY130_FD_SC_LP__DLYBUF4S15KAPWR_2%A_27_52# N_A_27_52#_M1005_s
+ N_A_27_52#_M1009_s N_A_27_52#_c_97_n N_A_27_52#_M1002_g N_A_27_52#_c_98_n
+ N_A_27_52#_M1004_g N_A_27_52#_c_99_n N_A_27_52#_c_106_n N_A_27_52#_c_107_n
+ N_A_27_52#_c_100_n N_A_27_52#_c_101_n N_A_27_52#_c_108_n N_A_27_52#_c_102_n
+ N_A_27_52#_c_103_n PM_SKY130_FD_SC_LP__DLYBUF4S15KAPWR_2%A_27_52#
x_PM_SKY130_FD_SC_LP__DLYBUF4S15KAPWR_2%A_282_52# N_A_282_52#_M1002_d
+ N_A_282_52#_M1004_d N_A_282_52#_c_169_n N_A_282_52#_M1008_g
+ N_A_282_52#_M1003_g N_A_282_52#_c_170_n N_A_282_52#_c_171_n
+ N_A_282_52#_c_172_n N_A_282_52#_c_177_n N_A_282_52#_c_173_n
+ N_A_282_52#_c_174_n N_A_282_52#_c_179_n
+ PM_SKY130_FD_SC_LP__DLYBUF4S15KAPWR_2%A_282_52#
x_PM_SKY130_FD_SC_LP__DLYBUF4S15KAPWR_2%A_394_52# N_A_394_52#_M1008_s
+ N_A_394_52#_M1003_s N_A_394_52#_M1000_g N_A_394_52#_M1001_g
+ N_A_394_52#_M1006_g N_A_394_52#_M1007_g N_A_394_52#_c_249_n
+ N_A_394_52#_c_251_n N_A_394_52#_c_254_n N_A_394_52#_c_244_n
+ N_A_394_52#_c_245_n N_A_394_52#_c_239_n N_A_394_52#_c_240_n
+ N_A_394_52#_c_273_n N_A_394_52#_c_241_n
+ PM_SKY130_FD_SC_LP__DLYBUF4S15KAPWR_2%A_394_52#
x_PM_SKY130_FD_SC_LP__DLYBUF4S15KAPWR_2%KAPWR N_KAPWR_M1009_d N_KAPWR_M1003_d
+ N_KAPWR_M1007_s KAPWR N_KAPWR_c_329_n N_KAPWR_c_342_n N_KAPWR_c_327_n
+ N_KAPWR_c_328_n KAPWR PM_SKY130_FD_SC_LP__DLYBUF4S15KAPWR_2%KAPWR
x_PM_SKY130_FD_SC_LP__DLYBUF4S15KAPWR_2%X N_X_M1000_s N_X_M1001_d X X X X X X X
+ N_X_c_383_n N_X_c_373_n X PM_SKY130_FD_SC_LP__DLYBUF4S15KAPWR_2%X
x_PM_SKY130_FD_SC_LP__DLYBUF4S15KAPWR_2%VGND N_VGND_M1005_d N_VGND_M1008_d
+ N_VGND_M1006_d N_VGND_c_401_n N_VGND_c_402_n N_VGND_c_403_n N_VGND_c_404_n
+ N_VGND_c_405_n N_VGND_c_406_n VGND N_VGND_c_407_n N_VGND_c_408_n
+ N_VGND_c_409_n N_VGND_c_410_n VGND PM_SKY130_FD_SC_LP__DLYBUF4S15KAPWR_2%VGND
x_PM_SKY130_FD_SC_LP__DLYBUF4S15KAPWR_2%VPWR VPWR N_VPWR_c_444_n N_VPWR_c_443_n
+ VPWR PM_SKY130_FD_SC_LP__DLYBUF4S15KAPWR_2%VPWR
cc_1 VNB N_A_M1005_g 0.0662132f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.47
cc_2 VNB A 0.0208018f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_3 VNB N_A_c_63_n 0.0329868f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.5
cc_4 VNB N_A_27_52#_c_97_n 0.021995f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.465
cc_5 VNB N_A_27_52#_c_98_n 0.0450206f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_6 VNB N_A_27_52#_c_99_n 0.0205357f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.335
cc_7 VNB N_A_27_52#_c_100_n 0.0050785f $X=-0.19 $Y=-0.245 $X2=0.325 $Y2=1.665
cc_8 VNB N_A_27_52#_c_101_n 0.0115829f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_27_52#_c_102_n 0.00219081f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_27_52#_c_103_n 9.66126e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_282_52#_c_169_n 0.0231219f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.465
cc_12 VNB N_A_282_52#_c_170_n 0.0226671f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.5
cc_13 VNB N_A_282_52#_c_171_n 0.011676f $X=-0.19 $Y=-0.245 $X2=0.325 $Y2=1.295
cc_14 VNB N_A_282_52#_c_172_n 0.0150178f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_282_52#_c_173_n 0.0124045f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_282_52#_c_174_n 0.0253565f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_394_52#_M1000_g 0.0515472f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_18 VNB N_A_394_52#_M1001_g 0.00156615f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.5
cc_19 VNB N_A_394_52#_M1006_g 0.0486632f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.665
cc_20 VNB N_A_394_52#_M1007_g 0.00167754f $X=-0.19 $Y=-0.245 $X2=0.325 $Y2=1.5
cc_21 VNB N_A_394_52#_c_239_n 0.0120567f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_394_52#_c_240_n 4.63484e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_394_52#_c_241_n 0.0414915f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB X 0.0402718f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_401_n 0.00648262f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_402_n 0.00647681f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.335
cc_27 VNB N_VGND_c_403_n 0.0132299f $X=-0.19 $Y=-0.245 $X2=0.325 $Y2=1.295
cc_28 VNB N_VGND_c_404_n 0.0223869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_405_n 0.0512685f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_406_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_407_n 0.0179296f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_408_n 0.0223295f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_409_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_410_n 0.276227f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VPWR_c_443_n 0.183584f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_36 VPB N_A_M1009_g 0.0260335f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.465
cc_37 VPB A 0.00827303f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_38 VPB N_A_c_63_n 0.00600603f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.5
cc_39 VPB N_A_27_52#_c_98_n 0.0465565f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_40 VPB N_A_27_52#_M1004_g 0.0252599f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_41 VPB N_A_27_52#_c_106_n 0.00794922f $X=-0.19 $Y=1.655 $X2=0.325 $Y2=1.295
cc_42 VPB N_A_27_52#_c_107_n 0.0277028f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_43 VPB N_A_27_52#_c_108_n 0.00375793f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_44 VPB N_A_27_52#_c_102_n 0.00497175f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_45 VPB N_A_282_52#_M1003_g 0.0425656f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_46 VPB N_A_282_52#_c_170_n 0.00905426f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.5
cc_47 VPB N_A_282_52#_c_177_n 0.0102217f $X=-0.19 $Y=1.655 $X2=0.325 $Y2=1.5
cc_48 VPB N_A_282_52#_c_174_n 0.0109227f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_49 VPB N_A_282_52#_c_179_n 0.0129686f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_50 VPB N_A_394_52#_M1001_g 0.0230649f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.5
cc_51 VPB N_A_394_52#_M1007_g 0.0236223f $X=-0.19 $Y=1.655 $X2=0.325 $Y2=1.5
cc_52 VPB N_A_394_52#_c_244_n 0.0118207f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_53 VPB N_A_394_52#_c_245_n 0.00462806f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_54 VPB N_A_394_52#_c_240_n 0.00376479f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_55 VPB N_KAPWR_c_327_n 0.0519559f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_56 VPB N_KAPWR_c_328_n 0.032581f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_57 VPB X 0.00701467f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_58 VPB N_X_c_373_n 0.00541438f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_59 VPB N_VPWR_c_444_n 0.118517f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_60 VPB N_VPWR_c_443_n 0.0471062f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_61 A N_A_27_52#_M1009_s 0.00237131f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_62 N_A_M1005_g N_A_27_52#_c_97_n 0.0123925f $X=0.475 $Y=0.47 $X2=0 $Y2=0
cc_63 A N_A_27_52#_c_98_n 0.00135678f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_64 N_A_c_63_n N_A_27_52#_c_98_n 0.0175907f $X=0.385 $Y=1.5 $X2=0 $Y2=0
cc_65 N_A_M1009_g N_A_27_52#_M1004_g 0.0160792f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_66 N_A_M1005_g N_A_27_52#_c_99_n 0.013604f $X=0.475 $Y=0.47 $X2=0 $Y2=0
cc_67 N_A_M1009_g N_A_27_52#_c_106_n 7.4234e-19 $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_68 A N_A_27_52#_c_106_n 0.0239868f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_69 N_A_c_63_n N_A_27_52#_c_106_n 7.87914e-19 $X=0.385 $Y=1.5 $X2=0 $Y2=0
cc_70 N_A_M1009_g N_A_27_52#_c_107_n 0.0141802f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_71 N_A_M1005_g N_A_27_52#_c_100_n 0.0119525f $X=0.475 $Y=0.47 $X2=0 $Y2=0
cc_72 A N_A_27_52#_c_100_n 0.0106601f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_73 N_A_M1005_g N_A_27_52#_c_101_n 0.00435937f $X=0.475 $Y=0.47 $X2=0 $Y2=0
cc_74 A N_A_27_52#_c_101_n 0.0289379f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_75 N_A_c_63_n N_A_27_52#_c_101_n 0.00100334f $X=0.385 $Y=1.5 $X2=0 $Y2=0
cc_76 N_A_M1009_g N_A_27_52#_c_108_n 0.00997145f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_77 A N_A_27_52#_c_108_n 0.00941865f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_78 N_A_M1009_g N_A_27_52#_c_102_n 0.0022019f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_79 A N_A_27_52#_c_102_n 0.0114464f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_80 N_A_c_63_n N_A_27_52#_c_102_n 0.0013726f $X=0.385 $Y=1.5 $X2=0 $Y2=0
cc_81 N_A_M1005_g N_A_27_52#_c_103_n 0.00532732f $X=0.475 $Y=0.47 $X2=0 $Y2=0
cc_82 A N_A_27_52#_c_103_n 0.0179575f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_83 N_A_c_63_n N_A_27_52#_c_103_n 9.52655e-19 $X=0.385 $Y=1.5 $X2=0 $Y2=0
cc_84 N_A_M1009_g N_KAPWR_c_329_n 0.00635965f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_85 N_A_M1009_g N_KAPWR_c_328_n 0.00551004f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_86 N_A_M1005_g N_VGND_c_401_n 0.00373445f $X=0.475 $Y=0.47 $X2=0 $Y2=0
cc_87 N_A_M1005_g N_VGND_c_407_n 0.00547602f $X=0.475 $Y=0.47 $X2=0 $Y2=0
cc_88 N_A_M1005_g N_VGND_c_410_n 0.00742906f $X=0.475 $Y=0.47 $X2=0 $Y2=0
cc_89 N_A_M1009_g N_VPWR_c_444_n 0.0054895f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_90 N_A_M1009_g N_VPWR_c_443_n 0.00699065f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_91 N_A_27_52#_c_98_n N_A_282_52#_M1003_g 0.00262015f $X=1.335 $Y=1.93 $X2=0
+ $Y2=0
cc_92 N_A_27_52#_c_98_n N_A_282_52#_c_170_n 0.00552637f $X=1.335 $Y=1.93 $X2=0
+ $Y2=0
cc_93 N_A_27_52#_c_97_n N_A_282_52#_c_172_n 0.00510471f $X=1.335 $Y=1.37 $X2=0
+ $Y2=0
cc_94 N_A_27_52#_c_98_n N_A_282_52#_c_172_n 0.00414437f $X=1.335 $Y=1.93 $X2=0
+ $Y2=0
cc_95 N_A_27_52#_c_102_n N_A_282_52#_c_172_n 0.00828764f $X=1.087 $Y=1.6 $X2=0
+ $Y2=0
cc_96 N_A_27_52#_c_103_n N_A_282_52#_c_172_n 0.022177f $X=1.085 $Y=1.535 $X2=0
+ $Y2=0
cc_97 N_A_27_52#_c_98_n N_A_282_52#_c_177_n 0.00361912f $X=1.335 $Y=1.93 $X2=0
+ $Y2=0
cc_98 N_A_27_52#_M1004_g N_A_282_52#_c_177_n 0.00319298f $X=1.335 $Y=2.595 $X2=0
+ $Y2=0
cc_99 N_A_27_52#_c_102_n N_A_282_52#_c_177_n 0.0285056f $X=1.087 $Y=1.6 $X2=0
+ $Y2=0
cc_100 N_A_27_52#_c_98_n N_A_282_52#_c_179_n 0.00392394f $X=1.335 $Y=1.93 $X2=0
+ $Y2=0
cc_101 N_A_27_52#_M1004_g N_A_282_52#_c_179_n 0.0114869f $X=1.335 $Y=2.595 $X2=0
+ $Y2=0
cc_102 N_A_27_52#_c_102_n N_A_282_52#_c_179_n 0.00501863f $X=1.087 $Y=1.6 $X2=0
+ $Y2=0
cc_103 N_A_27_52#_c_108_n N_KAPWR_M1009_d 0.0114913f $X=0.91 $Y=2.117 $X2=-0.19
+ $Y2=-0.245
cc_104 N_A_27_52#_c_102_n N_KAPWR_M1009_d 0.00700712f $X=1.087 $Y=1.6 $X2=-0.19
+ $Y2=-0.245
cc_105 N_A_27_52#_M1004_g N_KAPWR_c_329_n 0.00612446f $X=1.335 $Y=2.595 $X2=0
+ $Y2=0
cc_106 N_A_27_52#_c_107_n N_KAPWR_c_329_n 0.0294215f $X=0.26 $Y=2.915 $X2=0
+ $Y2=0
cc_107 N_A_27_52#_c_108_n N_KAPWR_c_329_n 0.0233037f $X=0.91 $Y=2.117 $X2=0
+ $Y2=0
cc_108 N_A_27_52#_c_102_n N_KAPWR_c_329_n 0.00118774f $X=1.087 $Y=1.6 $X2=0
+ $Y2=0
cc_109 N_A_27_52#_M1004_g N_KAPWR_c_328_n 0.00935473f $X=1.335 $Y=2.595 $X2=0
+ $Y2=0
cc_110 N_A_27_52#_c_107_n N_KAPWR_c_328_n 0.0377828f $X=0.26 $Y=2.915 $X2=0
+ $Y2=0
cc_111 N_A_27_52#_c_108_n N_KAPWR_c_328_n 0.00642807f $X=0.91 $Y=2.117 $X2=0
+ $Y2=0
cc_112 N_A_27_52#_c_102_n N_KAPWR_c_328_n 0.0140651f $X=1.087 $Y=1.6 $X2=0 $Y2=0
cc_113 N_A_27_52#_c_100_n N_VGND_M1005_d 0.0229926f $X=0.91 $Y=0.92 $X2=-0.19
+ $Y2=-0.245
cc_114 N_A_27_52#_c_103_n N_VGND_M1005_d 0.00497587f $X=1.085 $Y=1.535 $X2=-0.19
+ $Y2=-0.245
cc_115 N_A_27_52#_c_97_n N_VGND_c_401_n 0.0061026f $X=1.335 $Y=1.37 $X2=0 $Y2=0
cc_116 N_A_27_52#_c_100_n N_VGND_c_401_n 0.0252704f $X=0.91 $Y=0.92 $X2=0 $Y2=0
cc_117 N_A_27_52#_c_97_n N_VGND_c_405_n 0.00560159f $X=1.335 $Y=1.37 $X2=0 $Y2=0
cc_118 N_A_27_52#_c_99_n N_VGND_c_407_n 0.0152237f $X=0.26 $Y=0.47 $X2=0 $Y2=0
cc_119 N_A_27_52#_c_97_n N_VGND_c_410_n 0.0123684f $X=1.335 $Y=1.37 $X2=0 $Y2=0
cc_120 N_A_27_52#_c_99_n N_VGND_c_410_n 0.0118277f $X=0.26 $Y=0.47 $X2=0 $Y2=0
cc_121 N_A_27_52#_c_100_n N_VGND_c_410_n 0.0203772f $X=0.91 $Y=0.92 $X2=0 $Y2=0
cc_122 N_A_27_52#_M1004_g N_VPWR_c_444_n 0.00547432f $X=1.335 $Y=2.595 $X2=0
+ $Y2=0
cc_123 N_A_27_52#_c_107_n N_VPWR_c_444_n 0.0210467f $X=0.26 $Y=2.915 $X2=0 $Y2=0
cc_124 N_A_27_52#_M1009_s N_VPWR_c_443_n 0.00111591f $X=0.135 $Y=1.835 $X2=0
+ $Y2=0
cc_125 N_A_27_52#_M1004_g N_VPWR_c_443_n 0.00735386f $X=1.335 $Y=2.595 $X2=0
+ $Y2=0
cc_126 N_A_27_52#_c_107_n N_VPWR_c_443_n 0.00308298f $X=0.26 $Y=2.915 $X2=0
+ $Y2=0
cc_127 N_A_282_52#_c_169_n N_A_394_52#_M1000_g 0.0154668f $X=2.31 $Y=1.37 $X2=0
+ $Y2=0
cc_128 N_A_282_52#_M1003_g N_A_394_52#_M1001_g 0.0159437f $X=2.31 $Y=2.595 $X2=0
+ $Y2=0
cc_129 N_A_282_52#_c_169_n N_A_394_52#_c_249_n 0.0245206f $X=2.31 $Y=1.37 $X2=0
+ $Y2=0
cc_130 N_A_282_52#_c_171_n N_A_394_52#_c_249_n 0.0577683f $X=1.55 $Y=0.435 $X2=0
+ $Y2=0
cc_131 N_A_282_52#_c_169_n N_A_394_52#_c_251_n 0.0148888f $X=2.31 $Y=1.37 $X2=0
+ $Y2=0
cc_132 N_A_282_52#_c_173_n N_A_394_52#_c_251_n 0.0291078f $X=2.52 $Y=1.535 $X2=0
+ $Y2=0
cc_133 N_A_282_52#_c_174_n N_A_394_52#_c_251_n 0.00813341f $X=2.52 $Y=1.535
+ $X2=0 $Y2=0
cc_134 N_A_282_52#_c_169_n N_A_394_52#_c_254_n 8.78991e-19 $X=2.31 $Y=1.37 $X2=0
+ $Y2=0
cc_135 N_A_282_52#_c_170_n N_A_394_52#_c_254_n 0.00503939f $X=2.2 $Y=1.535 $X2=0
+ $Y2=0
cc_136 N_A_282_52#_c_171_n N_A_394_52#_c_254_n 0.00858119f $X=1.55 $Y=0.435
+ $X2=0 $Y2=0
cc_137 N_A_282_52#_c_172_n N_A_394_52#_c_254_n 0.0121129f $X=1.755 $Y=1.655
+ $X2=0 $Y2=0
cc_138 N_A_282_52#_c_173_n N_A_394_52#_c_254_n 0.0177106f $X=2.52 $Y=1.535 $X2=0
+ $Y2=0
cc_139 N_A_282_52#_c_173_n N_A_394_52#_c_244_n 0.0106947f $X=2.52 $Y=1.535 $X2=0
+ $Y2=0
cc_140 N_A_282_52#_c_174_n N_A_394_52#_c_244_n 0.0048475f $X=2.52 $Y=1.535 $X2=0
+ $Y2=0
cc_141 N_A_282_52#_M1003_g N_A_394_52#_c_245_n 0.0205083f $X=2.31 $Y=2.595 $X2=0
+ $Y2=0
cc_142 N_A_282_52#_c_170_n N_A_394_52#_c_245_n 0.00459953f $X=2.2 $Y=1.535 $X2=0
+ $Y2=0
cc_143 N_A_282_52#_c_177_n N_A_394_52#_c_245_n 0.00990869f $X=1.755 $Y=2.1 $X2=0
+ $Y2=0
cc_144 N_A_282_52#_c_173_n N_A_394_52#_c_245_n 0.0276207f $X=2.52 $Y=1.535 $X2=0
+ $Y2=0
cc_145 N_A_282_52#_c_174_n N_A_394_52#_c_245_n 0.00373286f $X=2.52 $Y=1.535
+ $X2=0 $Y2=0
cc_146 N_A_282_52#_c_179_n N_A_394_52#_c_245_n 0.0129926f $X=1.55 $Y=2.265 $X2=0
+ $Y2=0
cc_147 N_A_282_52#_c_169_n N_A_394_52#_c_239_n 0.00289451f $X=2.31 $Y=1.37 $X2=0
+ $Y2=0
cc_148 N_A_282_52#_c_173_n N_A_394_52#_c_239_n 0.0207685f $X=2.52 $Y=1.535 $X2=0
+ $Y2=0
cc_149 N_A_282_52#_c_174_n N_A_394_52#_c_239_n 0.0027866f $X=2.52 $Y=1.535 $X2=0
+ $Y2=0
cc_150 N_A_282_52#_M1003_g N_A_394_52#_c_240_n 0.00210429f $X=2.31 $Y=2.595
+ $X2=0 $Y2=0
cc_151 N_A_282_52#_c_173_n N_A_394_52#_c_240_n 0.00227963f $X=2.52 $Y=1.535
+ $X2=0 $Y2=0
cc_152 N_A_282_52#_c_174_n N_A_394_52#_c_240_n 0.00140233f $X=2.52 $Y=1.535
+ $X2=0 $Y2=0
cc_153 N_A_282_52#_M1003_g N_A_394_52#_c_273_n 0.0184516f $X=2.31 $Y=2.595 $X2=0
+ $Y2=0
cc_154 N_A_282_52#_c_179_n N_A_394_52#_c_273_n 0.0651214f $X=1.55 $Y=2.265 $X2=0
+ $Y2=0
cc_155 N_A_282_52#_c_174_n N_A_394_52#_c_241_n 0.0101988f $X=2.52 $Y=1.535 $X2=0
+ $Y2=0
cc_156 N_A_282_52#_c_179_n N_KAPWR_c_329_n 0.020862f $X=1.55 $Y=2.265 $X2=0
+ $Y2=0
cc_157 N_A_282_52#_M1003_g N_KAPWR_c_342_n 0.00776393f $X=2.31 $Y=2.595 $X2=0
+ $Y2=0
cc_158 N_A_282_52#_M1003_g N_KAPWR_c_328_n 0.00571761f $X=2.31 $Y=2.595 $X2=0
+ $Y2=0
cc_159 N_A_282_52#_c_179_n N_KAPWR_c_328_n 0.049599f $X=1.55 $Y=2.265 $X2=0
+ $Y2=0
cc_160 N_A_282_52#_c_169_n N_VGND_c_402_n 0.00633549f $X=2.31 $Y=1.37 $X2=0
+ $Y2=0
cc_161 N_A_282_52#_c_169_n N_VGND_c_405_n 0.00525608f $X=2.31 $Y=1.37 $X2=0
+ $Y2=0
cc_162 N_A_282_52#_c_171_n N_VGND_c_405_n 0.0250858f $X=1.55 $Y=0.435 $X2=0
+ $Y2=0
cc_163 N_A_282_52#_c_169_n N_VGND_c_410_n 0.0116294f $X=2.31 $Y=1.37 $X2=0 $Y2=0
cc_164 N_A_282_52#_c_171_n N_VGND_c_410_n 0.0155553f $X=1.55 $Y=0.435 $X2=0
+ $Y2=0
cc_165 N_A_282_52#_M1003_g N_VPWR_c_444_n 0.0054895f $X=2.31 $Y=2.595 $X2=0
+ $Y2=0
cc_166 N_A_282_52#_c_179_n N_VPWR_c_444_n 0.0301474f $X=1.55 $Y=2.265 $X2=0
+ $Y2=0
cc_167 N_A_282_52#_M1004_d N_VPWR_c_443_n 0.00111591f $X=1.41 $Y=2.095 $X2=0
+ $Y2=0
cc_168 N_A_282_52#_M1003_g N_VPWR_c_443_n 0.00735774f $X=2.31 $Y=2.595 $X2=0
+ $Y2=0
cc_169 N_A_282_52#_c_179_n N_VPWR_c_443_n 0.00429274f $X=1.55 $Y=2.265 $X2=0
+ $Y2=0
cc_170 N_A_394_52#_c_244_n N_KAPWR_M1003_d 0.00502062f $X=2.855 $Y=1.91 $X2=0
+ $Y2=0
cc_171 N_A_394_52#_c_245_n N_KAPWR_M1003_d 0.00403229f $X=2.54 $Y=1.91 $X2=0
+ $Y2=0
cc_172 N_A_394_52#_M1001_g N_KAPWR_c_342_n 0.00818219f $X=3.17 $Y=2.465 $X2=0
+ $Y2=0
cc_173 N_A_394_52#_c_244_n N_KAPWR_c_342_n 0.027185f $X=2.855 $Y=1.91 $X2=0
+ $Y2=0
cc_174 N_A_394_52#_c_245_n N_KAPWR_c_342_n 0.00710046f $X=2.54 $Y=1.91 $X2=0
+ $Y2=0
cc_175 N_A_394_52#_c_239_n N_KAPWR_c_342_n 5.09408e-19 $X=2.94 $Y=1.625 $X2=0
+ $Y2=0
cc_176 N_A_394_52#_c_273_n N_KAPWR_c_342_n 0.0257788f $X=2.095 $Y=2.245 $X2=0
+ $Y2=0
cc_177 N_A_394_52#_M1007_g N_KAPWR_c_327_n 0.00838687f $X=3.6 $Y=2.465 $X2=0
+ $Y2=0
cc_178 N_A_394_52#_M1003_s N_KAPWR_c_328_n 0.00185431f $X=1.97 $Y=2.095 $X2=0
+ $Y2=0
cc_179 N_A_394_52#_M1001_g N_KAPWR_c_328_n 0.00976215f $X=3.17 $Y=2.465 $X2=0
+ $Y2=0
cc_180 N_A_394_52#_c_245_n N_KAPWR_c_328_n 0.0101491f $X=2.54 $Y=1.91 $X2=0
+ $Y2=0
cc_181 N_A_394_52#_c_273_n N_KAPWR_c_328_n 0.0304541f $X=2.095 $Y=2.245 $X2=0
+ $Y2=0
cc_182 N_A_394_52#_M1000_g X 0.00799384f $X=3.17 $Y=0.47 $X2=0 $Y2=0
cc_183 N_A_394_52#_M1001_g X 0.0014189f $X=3.17 $Y=2.465 $X2=0 $Y2=0
cc_184 N_A_394_52#_M1006_g X 0.021587f $X=3.6 $Y=0.47 $X2=0 $Y2=0
cc_185 N_A_394_52#_M1007_g X 0.00596988f $X=3.6 $Y=2.465 $X2=0 $Y2=0
cc_186 N_A_394_52#_c_239_n X 0.0370853f $X=2.94 $Y=1.625 $X2=0 $Y2=0
cc_187 N_A_394_52#_c_240_n X 0.00685385f $X=2.94 $Y=1.825 $X2=0 $Y2=0
cc_188 N_A_394_52#_c_241_n X 0.0142477f $X=3.6 $Y=1.46 $X2=0 $Y2=0
cc_189 N_A_394_52#_M1001_g X 0.0153824f $X=3.17 $Y=2.465 $X2=0 $Y2=0
cc_190 N_A_394_52#_M1007_g X 0.0322293f $X=3.6 $Y=2.465 $X2=0 $Y2=0
cc_191 N_A_394_52#_M1000_g N_X_c_383_n 0.00509113f $X=3.17 $Y=0.47 $X2=0 $Y2=0
cc_192 N_A_394_52#_M1006_g N_X_c_383_n 0.0114044f $X=3.6 $Y=0.47 $X2=0 $Y2=0
cc_193 N_A_394_52#_c_239_n N_X_c_383_n 0.00268957f $X=2.94 $Y=1.625 $X2=0 $Y2=0
cc_194 N_A_394_52#_c_241_n N_X_c_383_n 0.00225933f $X=3.6 $Y=1.46 $X2=0 $Y2=0
cc_195 N_A_394_52#_M1001_g N_X_c_373_n 0.00491728f $X=3.17 $Y=2.465 $X2=0 $Y2=0
cc_196 N_A_394_52#_M1007_g N_X_c_373_n 0.00698802f $X=3.6 $Y=2.465 $X2=0 $Y2=0
cc_197 N_A_394_52#_c_244_n N_X_c_373_n 0.0124458f $X=2.855 $Y=1.91 $X2=0 $Y2=0
cc_198 N_A_394_52#_c_239_n N_X_c_373_n 0.00881931f $X=2.94 $Y=1.625 $X2=0 $Y2=0
cc_199 N_A_394_52#_c_240_n N_X_c_373_n 6.38382e-19 $X=2.94 $Y=1.825 $X2=0 $Y2=0
cc_200 N_A_394_52#_c_241_n N_X_c_373_n 0.00399236f $X=3.6 $Y=1.46 $X2=0 $Y2=0
cc_201 N_A_394_52#_c_251_n N_VGND_M1008_d 0.0212625f $X=2.855 $Y=1.097 $X2=0
+ $Y2=0
cc_202 N_A_394_52#_c_239_n N_VGND_M1008_d 0.00400434f $X=2.94 $Y=1.625 $X2=0
+ $Y2=0
cc_203 N_A_394_52#_M1000_g N_VGND_c_402_n 0.00709289f $X=3.17 $Y=0.47 $X2=0
+ $Y2=0
cc_204 N_A_394_52#_c_249_n N_VGND_c_402_n 0.0143516f $X=2.095 $Y=0.435 $X2=0
+ $Y2=0
cc_205 N_A_394_52#_c_251_n N_VGND_c_402_n 0.0076609f $X=2.855 $Y=1.097 $X2=0
+ $Y2=0
cc_206 N_A_394_52#_c_239_n N_VGND_c_402_n 0.0103475f $X=2.94 $Y=1.625 $X2=0
+ $Y2=0
cc_207 N_A_394_52#_M1006_g N_VGND_c_404_n 0.00756872f $X=3.6 $Y=0.47 $X2=0 $Y2=0
cc_208 N_A_394_52#_c_249_n N_VGND_c_405_n 0.0140261f $X=2.095 $Y=0.435 $X2=0
+ $Y2=0
cc_209 N_A_394_52#_M1000_g N_VGND_c_408_n 0.0051159f $X=3.17 $Y=0.47 $X2=0 $Y2=0
cc_210 N_A_394_52#_M1006_g N_VGND_c_408_n 0.00352007f $X=3.6 $Y=0.47 $X2=0 $Y2=0
cc_211 N_A_394_52#_M1000_g N_VGND_c_410_n 0.00995643f $X=3.17 $Y=0.47 $X2=0
+ $Y2=0
cc_212 N_A_394_52#_M1006_g N_VGND_c_410_n 0.00613857f $X=3.6 $Y=0.47 $X2=0 $Y2=0
cc_213 N_A_394_52#_c_249_n N_VGND_c_410_n 0.00945114f $X=2.095 $Y=0.435 $X2=0
+ $Y2=0
cc_214 N_A_394_52#_M1001_g N_VPWR_c_444_n 0.00564131f $X=3.17 $Y=2.465 $X2=0
+ $Y2=0
cc_215 N_A_394_52#_M1007_g N_VPWR_c_444_n 0.00357668f $X=3.6 $Y=2.465 $X2=0
+ $Y2=0
cc_216 N_A_394_52#_c_273_n N_VPWR_c_444_n 0.0153681f $X=2.095 $Y=2.245 $X2=0
+ $Y2=0
cc_217 N_A_394_52#_M1003_s N_VPWR_c_443_n 0.00128324f $X=1.97 $Y=2.095 $X2=0
+ $Y2=0
cc_218 N_A_394_52#_M1001_g N_VPWR_c_443_n 0.00609677f $X=3.17 $Y=2.465 $X2=0
+ $Y2=0
cc_219 N_A_394_52#_M1007_g N_VPWR_c_443_n 0.00594354f $X=3.6 $Y=2.465 $X2=0
+ $Y2=0
cc_220 N_A_394_52#_c_273_n N_VPWR_c_443_n 0.00232024f $X=2.095 $Y=2.245 $X2=0
+ $Y2=0
cc_221 N_KAPWR_c_342_n X 0.0352577f $X=2.875 $Y=2.27 $X2=0 $Y2=0
cc_222 N_KAPWR_c_328_n X 0.0493321f $X=3.96 $Y=2.805 $X2=0 $Y2=0
cc_223 N_KAPWR_c_327_n N_X_c_373_n 0.0530223f $X=3.96 $Y=1.98 $X2=0 $Y2=0
cc_224 N_KAPWR_c_329_n N_VPWR_c_444_n 0.0227152f $X=0.76 $Y=2.49 $X2=0 $Y2=0
cc_225 N_KAPWR_c_342_n N_VPWR_c_444_n 0.0230277f $X=2.875 $Y=2.27 $X2=0 $Y2=0
cc_226 N_KAPWR_c_327_n N_VPWR_c_444_n 0.0174911f $X=3.96 $Y=1.98 $X2=0 $Y2=0
cc_227 N_KAPWR_c_328_n N_VPWR_c_444_n 0.0109138f $X=3.96 $Y=2.805 $X2=0 $Y2=0
cc_228 N_KAPWR_M1009_d N_VPWR_c_443_n 0.00460091f $X=0.55 $Y=1.835 $X2=0 $Y2=0
cc_229 N_KAPWR_M1003_d N_VPWR_c_443_n 0.00460091f $X=2.385 $Y=2.095 $X2=0 $Y2=0
cc_230 N_KAPWR_M1007_s N_VPWR_c_443_n 0.00246793f $X=3.675 $Y=1.835 $X2=0 $Y2=0
cc_231 N_KAPWR_c_329_n N_VPWR_c_443_n 0.00313462f $X=0.76 $Y=2.49 $X2=0 $Y2=0
cc_232 N_KAPWR_c_342_n N_VPWR_c_443_n 0.00312197f $X=2.875 $Y=2.27 $X2=0 $Y2=0
cc_233 N_KAPWR_c_327_n N_VPWR_c_443_n 0.0023645f $X=3.96 $Y=1.98 $X2=0 $Y2=0
cc_234 N_KAPWR_c_328_n N_VPWR_c_443_n 0.432008f $X=3.96 $Y=2.805 $X2=0 $Y2=0
cc_235 N_X_c_383_n N_VGND_c_408_n 0.0207025f $X=3.61 $Y=0.475 $X2=0 $Y2=0
cc_236 N_X_c_383_n N_VGND_c_410_n 0.0174088f $X=3.61 $Y=0.475 $X2=0 $Y2=0
cc_237 X N_VPWR_c_444_n 0.0278606f $X=3.515 $Y=1.95 $X2=0 $Y2=0
cc_238 N_X_M1001_d N_VPWR_c_443_n 0.001145f $X=3.245 $Y=1.835 $X2=0 $Y2=0
cc_239 X N_VPWR_c_443_n 0.0042941f $X=3.515 $Y=1.95 $X2=0 $Y2=0
