* File: sky130_fd_sc_lp__einvp_0.pex.spice
* Created: Fri Aug 28 10:33:35 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__EINVP_0%TE 1 3 6 10 13 15 16 17 18 23
c39 16 0 1.99867e-19 $X=0.72 $Y=0.925
r40 23 24 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.655
+ $Y=1.045 $X2=0.655 $Y2=1.045
r41 17 18 11.6823 $w=3.63e-07 $l=3.7e-07 $layer=LI1_cond $X=0.742 $Y=1.295
+ $X2=0.742 $Y2=1.665
r42 17 24 7.89345 $w=3.63e-07 $l=2.5e-07 $layer=LI1_cond $X=0.742 $Y=1.295
+ $X2=0.742 $Y2=1.045
r43 16 24 3.78885 $w=3.63e-07 $l=1.2e-07 $layer=LI1_cond $X=0.742 $Y=0.925
+ $X2=0.742 $Y2=1.045
r44 14 23 43.3659 $w=3.95e-07 $l=3.08e-07 $layer=POLY_cond $X=0.622 $Y=1.353
+ $X2=0.622 $Y2=1.045
r45 14 15 50.0695 $w=3.95e-07 $l=1.97e-07 $layer=POLY_cond $X=0.622 $Y=1.353
+ $X2=0.622 $Y2=1.55
r46 13 23 2.11198 $w=3.95e-07 $l=1.5e-08 $layer=POLY_cond $X=0.622 $Y=1.03
+ $X2=0.622 $Y2=1.045
r47 6 15 666.596 $w=1.5e-07 $l=1.3e-06 $layer=POLY_cond $X=0.5 $Y=2.85 $X2=0.5
+ $Y2=1.55
r48 1 13 24.4706 $w=3.95e-07 $l=1.5e-07 $layer=POLY_cond $X=0.715 $Y=0.88
+ $X2=0.715 $Y2=1.03
r49 1 10 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.93 $Y=0.88 $X2=0.93
+ $Y2=0.56
r50 1 3 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.5 $Y=0.88 $X2=0.5
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_LP__EINVP_0%A_32_70# 1 2 9 13 17 21 22 24
r36 22 27 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.95 $Y=2.095
+ $X2=0.95 $Y2=2.26
r37 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.95
+ $Y=2.095 $X2=0.95 $Y2=2.095
r38 19 24 0.94211 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=0.45 $Y=2.095
+ $X2=0.285 $Y2=2.095
r39 19 21 17.4613 $w=3.28e-07 $l=5e-07 $layer=LI1_cond $X=0.45 $Y=2.095 $X2=0.95
+ $Y2=2.095
r40 15 24 5.66538 $w=2.95e-07 $l=1.65e-07 $layer=LI1_cond $X=0.285 $Y=2.26
+ $X2=0.285 $Y2=2.095
r41 15 17 20.6043 $w=3.28e-07 $l=5.9e-07 $layer=LI1_cond $X=0.285 $Y=2.26
+ $X2=0.285 $Y2=2.85
r42 11 24 5.66538 $w=2.95e-07 $l=1.81659e-07 $layer=LI1_cond $X=0.25 $Y=1.93
+ $X2=0.285 $Y2=2.095
r43 11 13 60.7249 $w=2.58e-07 $l=1.37e-06 $layer=LI1_cond $X=0.25 $Y=1.93
+ $X2=0.25 $Y2=0.56
r44 9 27 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.025 $Y=2.74
+ $X2=1.025 $Y2=2.26
r45 2 17 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=0.16
+ $Y=2.64 $X2=0.285 $Y2=2.85
r46 1 13 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.16
+ $Y=0.35 $X2=0.285 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_LP__EINVP_0%A 3 6 8 9 10 11 17 19
c31 19 0 1.99867e-19 $X=1.53 $Y=0.88
r32 17 20 80.5075 $w=5.7e-07 $l=5.05e-07 $layer=POLY_cond $X=1.53 $Y=1.045
+ $X2=1.53 $Y2=1.55
r33 17 19 48.5934 $w=5.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.53 $Y=1.045
+ $X2=1.53 $Y2=0.88
r34 17 18 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.65
+ $Y=1.045 $X2=1.65 $Y2=1.045
r35 10 11 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=1.7 $Y=1.665 $X2=1.7
+ $Y2=2.035
r36 9 10 15.7927 $w=2.68e-07 $l=3.7e-07 $layer=LI1_cond $X=1.7 $Y=1.295 $X2=1.7
+ $Y2=1.665
r37 9 18 10.6708 $w=2.68e-07 $l=2.5e-07 $layer=LI1_cond $X=1.7 $Y=1.295 $X2=1.7
+ $Y2=1.045
r38 8 18 5.12197 $w=2.68e-07 $l=1.2e-07 $layer=LI1_cond $X=1.7 $Y=0.925 $X2=1.7
+ $Y2=1.045
r39 6 20 610.191 $w=1.5e-07 $l=1.19e-06 $layer=POLY_cond $X=1.415 $Y=2.74
+ $X2=1.415 $Y2=1.55
r40 3 19 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.32 $Y=0.56 $X2=1.32
+ $Y2=0.88
.ends

.subckt PM_SKY130_FD_SC_LP__EINVP_0%VPWR 1 6 8 10 17 18 21
r25 21 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r26 17 18 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r27 15 21 9.05715 $w=1.7e-07 $l=1.78e-07 $layer=LI1_cond $X=0.975 $Y=3.33
+ $X2=0.797 $Y2=3.33
r28 15 17 45.9947 $w=1.68e-07 $l=7.05e-07 $layer=LI1_cond $X=0.975 $Y=3.33
+ $X2=1.68 $Y2=3.33
r29 13 22 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r30 12 13 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r31 10 21 9.05715 $w=1.7e-07 $l=1.77e-07 $layer=LI1_cond $X=0.62 $Y=3.33
+ $X2=0.797 $Y2=3.33
r32 10 12 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=0.62 $Y=3.33
+ $X2=0.24 $Y2=3.33
r33 8 18 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=0.96 $Y=3.33
+ $X2=1.68 $Y2=3.33
r34 8 22 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=0.96 $Y=3.33
+ $X2=0.72 $Y2=3.33
r35 4 21 1.11826 $w=3.55e-07 $l=8.5e-08 $layer=LI1_cond $X=0.797 $Y=3.245
+ $X2=0.797 $Y2=3.33
r36 4 6 21.7503 $w=3.53e-07 $l=6.7e-07 $layer=LI1_cond $X=0.797 $Y=3.245
+ $X2=0.797 $Y2=2.575
r37 1 6 300 $w=1.7e-07 $l=2.65518e-07 $layer=licon1_PDIFF $count=2 $X=0.575
+ $Y=2.64 $X2=0.81 $Y2=2.575
.ends

.subckt PM_SKY130_FD_SC_LP__EINVP_0%Z 1 2 8 12 14 15 21
r34 15 21 7.16384 $w=3.68e-07 $l=2.3e-07 $layer=LI1_cond $X=1.65 $Y=2.775
+ $X2=1.65 $Y2=2.545
r35 14 26 19.6864 $w=1.98e-07 $l=3.55e-07 $layer=LI1_cond $X=1.65 $Y=2.39
+ $X2=1.295 $Y2=2.39
r36 14 21 2.41259 $w=5.38e-07 $l=5.5e-08 $layer=LI1_cond $X=1.65 $Y=2.49
+ $X2=1.65 $Y2=2.545
r37 9 12 8.3814 $w=3.28e-07 $l=2.4e-07 $layer=LI1_cond $X=1.295 $Y=0.505
+ $X2=1.535 $Y2=0.505
r38 8 26 1.35108 $w=1.8e-07 $l=1e-07 $layer=LI1_cond $X=1.295 $Y=2.29 $X2=1.295
+ $Y2=2.39
r39 7 9 4.28565 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=1.295 $Y=0.67
+ $X2=1.295 $Y2=0.505
r40 7 8 99.8182 $w=1.78e-07 $l=1.62e-06 $layer=LI1_cond $X=1.295 $Y=0.67
+ $X2=1.295 $Y2=2.29
r41 2 21 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=1.49
+ $Y=2.42 $X2=1.63 $Y2=2.545
r42 1 12 182 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=1 $X=1.395
+ $Y=0.35 $X2=1.535 $Y2=0.505
.ends

.subckt PM_SKY130_FD_SC_LP__EINVP_0%VGND 1 6 8 10 17 18 21
r21 21 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r22 17 18 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r23 15 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.88 $Y=0 $X2=0.715
+ $Y2=0
r24 15 17 52.1925 $w=1.68e-07 $l=8e-07 $layer=LI1_cond $X=0.88 $Y=0 $X2=1.68
+ $Y2=0
r25 13 22 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r26 12 13 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r27 10 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.55 $Y=0 $X2=0.715
+ $Y2=0
r28 10 12 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=0.55 $Y=0 $X2=0.24
+ $Y2=0
r29 8 18 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=0.96 $Y=0 $X2=1.68
+ $Y2=0
r30 8 22 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=0.96 $Y=0 $X2=0.72
+ $Y2=0
r31 4 21 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.715 $Y=0.085
+ $X2=0.715 $Y2=0
r32 4 6 16.0644 $w=3.28e-07 $l=4.6e-07 $layer=LI1_cond $X=0.715 $Y=0.085
+ $X2=0.715 $Y2=0.545
r33 1 6 182 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_NDIFF $count=1 $X=0.575
+ $Y=0.35 $X2=0.715 $Y2=0.545
.ends

