* File: sky130_fd_sc_lp__srdlxtp_1.spice
* Created: Fri Aug 28 11:33:22 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__srdlxtp_1.pex.spice"
.subckt sky130_fd_sc_lp__srdlxtp_1  VNB VPB D GATE SLEEP_B VPWR KAPWR Q VGND
* 
* VGND	VGND
* Q	Q
* KAPWR	KAPWR
* VPWR	VPWR
* SLEEP_B	SLEEP_B
* GATE	GATE
* D	D
* VPB	VPB
* VNB	VNB
MM1013 N_A_114_179#_M1013_d N_A_84_153#_M1013_g N_VGND_M1013_s VNB NSHORT L=0.15
+ W=0.42 AD=0.1197 AS=0.1197 PD=1.41 PS=1.41 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1014 N_VGND_M1014_d N_D_M1014_g N_A_226_491#_M1014_s VNB NSHORT L=0.15 W=0.42
+ AD=0.1426 AS=0.1197 PD=1.13 PS=1.41 NRD=67.14 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75004 A=0.063 P=1.14 MULT=1
MM1025 N_A_476_47#_M1025_d N_A_226_491#_M1025_g N_VGND_M1014_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0882 AS=0.1426 PD=0.84 PS=1.13 NRD=1.428 NRS=29.988 M=1 R=2.8
+ SA=75001 SB=75003.3 A=0.063 P=1.14 MULT=1
MM1002 A_590_47# N_A_114_179#_M1002_g N_A_476_47#_M1025_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.0882 PD=0.63 PS=0.84 NRD=14.28 NRS=38.568 M=1 R=2.8
+ SA=75001.5 SB=75002.7 A=0.063 P=1.14 MULT=1
MM1003 N_A_662_47#_M1003_d N_A_114_179#_M1003_g A_590_47# VNB NSHORT L=0.15
+ W=0.42 AD=0.09555 AS=0.0441 PD=0.875 PS=0.63 NRD=49.992 NRS=14.28 M=1 R=2.8
+ SA=75001.9 SB=75002.4 A=0.063 P=1.14 MULT=1
MM1006 A_783_47# N_A_84_153#_M1006_g N_A_662_47#_M1003_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0504 AS=0.09555 PD=0.66 PS=0.875 NRD=18.564 NRS=0 M=1 R=2.8
+ SA=75002.5 SB=75001.7 A=0.063 P=1.14 MULT=1
MM1007 A_861_47# N_A_831_21#_M1007_g A_783_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0504 PD=0.63 PS=0.66 NRD=14.28 NRS=18.564 M=1 R=2.8 SA=75002.9
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1009 N_VGND_M1009_d N_A_831_21#_M1009_g A_861_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75003.3
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1016 A_1019_47# N_A_662_47#_M1016_g N_VGND_M1009_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75003.7
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1005 N_A_831_21#_M1005_d N_A_662_47#_M1005_g A_1019_47# VNB NSHORT L=0.15
+ W=0.42 AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75004
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1023 A_1289_47# N_GATE_M1023_g N_A_84_153#_M1023_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1197 PD=0.63 PS=1.41 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.9 A=0.063 P=1.14 MULT=1
MM1017 A_1361_47# N_SLEEP_B_M1017_g A_1289_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0441 PD=0.63 PS=0.63 NRD=14.28 NRS=14.28 M=1 R=2.8 SA=75000.6
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1019 N_VGND_M1019_d N_SLEEP_B_M1019_g A_1361_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.9
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1011 N_VGND_M1011_d N_A_662_47#_M1011_g N_A_1530_367#_M1011_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.0952 AS=0.1197 PD=0.823333 PS=1.41 NRD=32.856 NRS=0 M=1
+ R=2.8 SA=75000.2 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1010 N_Q_M1010_d N_A_1530_367#_M1010_g N_VGND_M1011_d VNB NSHORT L=0.15 W=0.84
+ AD=0.2394 AS=0.1904 PD=2.25 PS=1.64667 NRD=0 NRS=0 M=1 R=5.6 SA=75000.5
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1004 N_A_114_179#_M1004_d N_A_84_153#_M1004_g N_VPWR_M1004_s VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.1824 AS=0.1824 PD=1.85 PS=1.85 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1022 N_VPWR_M1022_d N_D_M1022_g N_A_226_491#_M1022_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.3072 AS=0.1824 PD=1.6 PS=1.85 NRD=21.5321 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75003.4 A=0.096 P=1.58 MULT=1
MM1012 N_A_476_47#_M1012_d N_A_226_491#_M1012_g N_VPWR_M1022_d VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.0896 AS=0.3072 PD=0.92 PS=1.6 NRD=0 NRS=187.761 M=1
+ R=4.26667 SA=75001.3 SB=75002.3 A=0.096 P=1.58 MULT=1
MM1015 A_621_491# N_A_84_153#_M1015_g N_A_476_47#_M1012_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1104 AS=0.0896 PD=0.985 PS=0.92 NRD=36.1495 NRS=0 M=1 R=4.26667
+ SA=75001.8 SB=75001.8 A=0.096 P=1.58 MULT=1
MM1024 N_A_662_47#_M1024_d N_A_84_153#_M1024_g A_621_491# VPB PHIGHVT L=0.15
+ W=0.64 AD=0.138693 AS=0.1104 PD=1.08878 PS=0.985 NRD=36.9375 NRS=36.1495 M=1
+ R=4.26667 SA=75002.2 SB=75001.3 A=0.096 P=1.58 MULT=1
MM1020 A_849_419# N_A_114_179#_M1020_g N_A_662_47#_M1024_d VPB PHIGHVT L=0.25
+ W=1 AD=0.12 AS=0.216707 PD=1.24 PS=1.70122 NRD=12.7853 NRS=0 M=1 R=4 SA=125002
+ SB=125001 A=0.25 P=2.5 MULT=1
MM1001 N_KAPWR_M1001_d N_A_831_21#_M1001_g A_849_419# VPB PHIGHVT L=0.25 W=1
+ AD=0.285 AS=0.12 PD=2.57 PS=1.24 NRD=0 NRS=12.7853 M=1 R=4 SA=125002 SB=125000
+ A=0.25 P=2.5 MULT=1
MM1021 N_KAPWR_M1021_d N_A_662_47#_M1021_g N_A_831_21#_M1021_s VPB PHIGHVT
+ L=0.25 W=1 AD=0.216707 AS=0.285 PD=1.70122 PS=2.57 NRD=0 NRS=0 M=1 R=4
+ SA=125000 SB=125001 A=0.25 P=2.5 MULT=1
MM1026 N_A_84_153#_M1026_d N_GATE_M1026_g N_KAPWR_M1021_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1344 AS=0.138693 PD=1.06 PS=1.08878 NRD=43.0839 NRS=49.7622 M=1
+ R=4.26667 SA=75000.9 SB=75000.8 A=0.096 P=1.58 MULT=1
MM1018 N_KAPWR_M1018_d N_SLEEP_B_M1018_g N_A_84_153#_M1026_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.2272 AS=0.1344 PD=1.99 PS=1.06 NRD=21.5321 NRS=0 M=1 R=4.26667
+ SA=75001.4 SB=75000.3 A=0.096 P=1.58 MULT=1
MM1000 N_VPWR_M1000_d N_A_662_47#_M1000_g N_A_1530_367#_M1000_s VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.174383 AS=0.1824 PD=1.16211 PS=1.85 NRD=36.1495 NRS=0 M=1
+ R=4.26667 SA=75000.2 SB=75000.8 A=0.096 P=1.58 MULT=1
MM1008 N_Q_M1008_d N_A_1530_367#_M1008_g N_VPWR_M1000_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3591 AS=0.343317 PD=3.09 PS=2.28789 NRD=0 NRS=10.9335 M=1 R=8.4
+ SA=75000.6 SB=75000.2 A=0.189 P=2.82 MULT=1
DX27_noxref VNB VPB NWDIODE A=18.0959 P=23.05
*
.include "sky130_fd_sc_lp__srdlxtp_1.pxi.spice"
*
.ends
*
*
