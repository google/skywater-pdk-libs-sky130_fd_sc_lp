* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__fa_0 A B CIN VGND VNB VPB VPWR COUT SUM
X0 VGND A a_382_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 a_781_119# a_80_225# a_1059_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 a_781_457# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X3 a_224_119# B a_80_225# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 VPWR CIN a_781_457# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X5 a_781_119# B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 a_382_119# B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 a_1145_119# B a_1239_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 a_1059_119# CIN a_1161_457# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X9 VPWR A a_218_532# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X10 VGND A a_224_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X11 VPWR a_1059_119# SUM VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X12 a_1059_119# CIN a_1145_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X13 a_80_225# CIN a_382_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X14 a_1239_457# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X15 VGND CIN a_781_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X16 COUT a_80_225# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X17 a_1161_457# B a_1239_457# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X18 a_781_457# a_80_225# a_1059_119# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X19 VPWR A a_404_532# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X20 VGND a_1059_119# SUM VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X21 a_80_225# CIN a_404_532# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X22 COUT a_80_225# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X23 VGND A a_781_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X24 a_218_532# B a_80_225# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X25 VPWR A a_781_457# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X26 a_1239_119# A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X27 a_404_532# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
.ends
