* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__xor2_lp A B VGND VNB VPB VPWR X
M1000 a_272_119# B X VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=1.176e+11p ps=1.4e+06u
M1001 VPWR A a_159_419# VPB phighvt w=1e+06u l=250000u
+  ad=5.65e+11p pd=5.13e+06u as=5.65e+11p ps=5.13e+06u
M1002 a_114_119# a_84_93# VGND VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=4.35225e+11p ps=4.89e+06u
M1003 a_84_93# B a_446_68# VNB nshort w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=1.008e+11p ps=1.32e+06u
M1004 a_159_419# a_84_93# X VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=3e+11p ps=2.6e+06u
M1005 a_159_419# B VPWR VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND A a_272_119# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_446_68# B VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_610_68# A a_84_93# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1009 VGND A a_610_68# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_590_412# B a_84_93# VPB phighvt w=1e+06u l=250000u
+  ad=2.1e+11p pd=2.42e+06u as=2.85e+11p ps=2.57e+06u
M1011 VPWR A a_590_412# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1012 X a_84_93# a_114_119# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
