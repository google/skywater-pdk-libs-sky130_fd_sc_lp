* File: sky130_fd_sc_lp__sdfrtn_1.pex.spice
* Created: Fri Aug 28 11:28:11 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__SDFRTN_1%A_113_63# 1 2 7 9 12 15 16 18 21 25 32 33
+ 37 38
r80 38 43 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.26 $Y=1.12
+ $X2=3.26 $Y2=0.955
r81 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.26
+ $Y=1.12 $X2=3.26 $Y2=1.12
r82 31 33 9.39634 $w=4.78e-07 $l=1.65e-07 $layer=LI1_cond $X=1.26 $Y=2.205
+ $X2=1.425 $Y2=2.205
r83 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.26
+ $Y=2.13 $X2=1.26 $Y2=2.13
r84 22 25 1.40854 $w=2.68e-07 $l=3.3e-08 $layer=LI1_cond $X=0.672 $Y=0.43
+ $X2=0.705 $Y2=0.43
r85 21 34 3.3128 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=3.18 $Y=2.02 $X2=3.18
+ $Y2=2.195
r86 20 37 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.18 $Y=1.205
+ $X2=3.18 $Y2=1.12
r87 20 21 53.1711 $w=1.68e-07 $l=8.15e-07 $layer=LI1_cond $X=3.18 $Y=1.205
+ $X2=3.18 $Y2=2.02
r88 18 34 19.5655 $w=2.64e-07 $l=4.65242e-07 $layer=LI1_cond $X=2.79 $Y=2.36
+ $X2=3.18 $Y2=2.195
r89 18 33 89.0535 $w=1.68e-07 $l=1.365e-06 $layer=LI1_cond $X=2.79 $Y=2.36
+ $X2=1.425 $Y2=2.36
r90 17 28 2.71462 $w=4.8e-07 $l=1.40798e-07 $layer=LI1_cond $X=0.81 $Y=2.205
+ $X2=0.692 $Y2=2.155
r91 16 31 1.86887 $w=4.78e-07 $l=7.5e-08 $layer=LI1_cond $X=1.185 $Y=2.205
+ $X2=1.26 $Y2=2.205
r92 16 17 9.34436 $w=4.78e-07 $l=3.75e-07 $layer=LI1_cond $X=1.185 $Y=2.205
+ $X2=0.81 $Y2=2.205
r93 15 28 5.81704 $w=1.95e-07 $l=3.49857e-07 $layer=LI1_cond $X=0.672 $Y=1.815
+ $X2=0.692 $Y2=2.155
r94 14 22 2.66673 $w=1.95e-07 $l=1.35e-07 $layer=LI1_cond $X=0.672 $Y=0.565
+ $X2=0.672 $Y2=0.43
r95 14 15 71.0956 $w=1.93e-07 $l=1.25e-06 $layer=LI1_cond $X=0.672 $Y=0.565
+ $X2=0.672 $Y2=1.815
r96 12 43 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=3.17 $Y=0.505
+ $X2=3.17 $Y2=0.955
r97 7 32 34.6486 $w=3.13e-07 $l=3.05573e-07 $layer=POLY_cond $X=1.485 $Y=2.345
+ $X2=1.26 $Y2=2.155
r98 7 9 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=1.485 $Y=2.345
+ $X2=1.485 $Y2=2.775
r99 2 28 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.565
+ $Y=1.835 $X2=0.705 $Y2=1.98
r100 2 28 600 $w=1.7e-07 $l=5.60647e-07 $layer=licon1_PDIFF $count=1 $X=0.565
+ $Y=1.835 $X2=0.705 $Y2=2.33
r101 1 25 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=0.565
+ $Y=0.315 $X2=0.705 $Y2=0.46
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRTN_1%SCD 1 3 5 8 10 12 13 15 16 24 28
c52 12 0 8.49613e-20 $X=1.8 $Y=1.79
c53 10 0 1.41229e-20 $X=1.762 $Y=1.095
r54 21 24 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.115 $Y=0.83
+ $X2=1.28 $Y2=0.83
r55 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.115
+ $Y=0.83 $X2=1.115 $Y2=0.83
r56 16 28 2.91497 $w=3.5e-07 $l=1.22e-07 $layer=LI1_cond $X=1.762 $Y=0.92
+ $X2=1.64 $Y2=0.92
r57 16 28 0.75732 $w=3.48e-07 $l=2.3e-08 $layer=LI1_cond $X=1.617 $Y=0.92
+ $X2=1.64 $Y2=0.92
r58 15 16 13.7305 $w=3.48e-07 $l=4.17e-07 $layer=LI1_cond $X=1.2 $Y=0.92
+ $X2=1.617 $Y2=0.92
r59 15 22 2.79879 $w=3.48e-07 $l=8.5e-08 $layer=LI1_cond $X=1.2 $Y=0.92
+ $X2=1.115 $Y2=0.92
r60 13 27 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.8 $Y=1.79 $X2=1.8
+ $Y2=1.955
r61 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.8
+ $Y=1.79 $X2=1.8 $Y2=1.79
r62 10 16 4.1813 $w=2.45e-07 $l=1.75e-07 $layer=LI1_cond $X=1.762 $Y=1.095
+ $X2=1.762 $Y2=0.92
r63 10 12 32.6917 $w=2.43e-07 $l=6.95e-07 $layer=LI1_cond $X=1.762 $Y=1.095
+ $X2=1.762 $Y2=1.79
r64 8 27 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=1.845 $Y=2.775
+ $X2=1.845 $Y2=1.955
r65 3 5 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.73 $Y=0.825 $X2=1.73
+ $Y2=0.505
r66 1 3 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.655 $Y=0.9
+ $X2=1.73 $Y2=0.825
r67 1 24 192.287 $w=1.5e-07 $l=3.75e-07 $layer=POLY_cond $X=1.655 $Y=0.9
+ $X2=1.28 $Y2=0.9
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRTN_1%SCE 3 7 9 13 17 19 22 23 25 26 34
c72 34 0 8.49613e-20 $X=2.37 $Y=2.02
c73 22 0 8.69653e-20 $X=2.18 $Y=1.22
c74 9 0 9.05516e-21 $X=2.015 $Y=1.31
r75 35 39 4.47161 $w=4.72e-07 $l=1.73e-07 $layer=LI1_cond $X=2.37 $Y=1.84
+ $X2=2.197 $Y2=1.84
r76 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.37
+ $Y=2.02 $X2=2.37 $Y2=2.02
r77 26 35 6.97881 $w=4.72e-07 $l=2.7e-07 $layer=LI1_cond $X=2.64 $Y=1.84
+ $X2=2.37 $Y2=1.84
r78 25 39 0.956356 $w=4.72e-07 $l=3.7e-08 $layer=LI1_cond $X=2.16 $Y=1.84
+ $X2=2.197 $Y2=1.84
r79 23 31 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=2.18 $Y=1.22 $X2=2.18
+ $Y2=1.31
r80 23 30 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.18 $Y=1.22
+ $X2=2.18 $Y2=1.055
r81 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.18
+ $Y=1.22 $X2=2.18 $Y2=1.22
r82 20 39 3.70158 $w=2.85e-07 $l=2.65e-07 $layer=LI1_cond $X=2.197 $Y=1.575
+ $X2=2.197 $Y2=1.84
r83 20 22 14.355 $w=2.83e-07 $l=3.55e-07 $layer=LI1_cond $X=2.197 $Y=1.575
+ $X2=2.197 $Y2=1.22
r84 15 34 61.7298 $w=2.85e-07 $l=4.39829e-07 $layer=POLY_cond $X=2.735 $Y=2.185
+ $X2=2.37 $Y2=2.02
r85 15 17 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=2.735 $Y=2.185
+ $X2=2.735 $Y2=2.775
r86 13 30 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=2.09 $Y=0.505
+ $X2=2.09 $Y2=1.055
r87 10 19 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.565 $Y=1.31
+ $X2=0.49 $Y2=1.31
r88 9 31 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.015 $Y=1.31
+ $X2=2.18 $Y2=1.31
r89 9 10 743.511 $w=1.5e-07 $l=1.45e-06 $layer=POLY_cond $X=2.015 $Y=1.31
+ $X2=0.565 $Y2=1.31
r90 5 19 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.49 $Y=1.385
+ $X2=0.49 $Y2=1.31
r91 5 7 394.83 $w=1.5e-07 $l=7.7e-07 $layer=POLY_cond $X=0.49 $Y=1.385 $X2=0.49
+ $Y2=2.155
r92 1 19 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.49 $Y=1.235
+ $X2=0.49 $Y2=1.31
r93 1 3 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=0.49 $Y=1.235 $X2=0.49
+ $Y2=0.525
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRTN_1%D 3 5 7 9
c47 3 0 8.69653e-20 $X=2.75 $Y=0.505
r48 9 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.72
+ $Y=1.235 $X2=2.72 $Y2=1.235
r49 5 12 80.2256 $w=3.18e-07 $l=5.44169e-07 $layer=POLY_cond $X=3.095 $Y=1.675
+ $X2=2.862 $Y2=1.235
r50 5 7 564.043 $w=1.5e-07 $l=1.1e-06 $layer=POLY_cond $X=3.095 $Y=1.675
+ $X2=3.095 $Y2=2.775
r51 1 12 38.5432 $w=3.18e-07 $l=2.13787e-07 $layer=POLY_cond $X=2.75 $Y=1.07
+ $X2=2.862 $Y2=1.235
r52 1 3 289.713 $w=1.5e-07 $l=5.65e-07 $layer=POLY_cond $X=2.75 $Y=1.07 $X2=2.75
+ $Y2=0.505
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRTN_1%RESET_B 3 7 9 11 14 17 19 22 26 30 32 35 37
+ 38 41 42 43 44 46 47 48 51 52 56 57 61 62 68 69 72 73 78 79 89
c239 69 0 1.74942e-19 $X=7.92 $Y=2.035
c240 61 0 1.22969e-19 $X=7.775 $Y=2.035
c241 35 0 9.85956e-20 $X=7.83 $Y=2.46
c242 26 0 3.32213e-20 $X=11.055 $Y=0.845
r243 87 89 0.101363 $w=5.88e-07 $l=5e-09 $layer=LI1_cond $X=10.315 $Y=1.67
+ $X2=10.32 $Y2=1.67
r244 78 80 46.1517 $w=4.2e-07 $l=1.65e-07 $layer=POLY_cond $X=10.92 $Y=1.46
+ $X2=10.92 $Y2=1.295
r245 78 79 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=10.875
+ $Y=1.46 $X2=10.875 $Y2=1.46
r246 72 73 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.545
+ $Y=1.69 $X2=3.545 $Y2=1.69
r247 68 69 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=2.035
+ $X2=7.92 $Y2=2.035
r248 65 73 16.9188 $w=2.33e-07 $l=3.45e-07 $layer=LI1_cond $X=3.577 $Y=2.035
+ $X2=3.577 $Y2=1.69
r249 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=2.035
+ $X2=3.6 $Y2=2.035
r250 62 64 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.745 $Y=2.035
+ $X2=3.6 $Y2=2.035
r251 61 68 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.775 $Y=2.035
+ $X2=7.92 $Y2=2.035
r252 61 62 4.98761 $w=1.4e-07 $l=4.03e-06 $layer=MET1_cond $X=7.775 $Y=2.035
+ $X2=3.745 $Y2=2.035
r253 57 79 1.52044 $w=5.88e-07 $l=7.5e-08 $layer=LI1_cond $X=10.8 $Y=1.67
+ $X2=10.875 $Y2=1.67
r254 56 87 2.22928 $w=5.9e-07 $l=8.5e-08 $layer=LI1_cond $X=10.23 $Y=1.67
+ $X2=10.315 $Y2=1.67
r255 56 57 8.91991 $w=5.88e-07 $l=4.4e-07 $layer=LI1_cond $X=10.36 $Y=1.67
+ $X2=10.8 $Y2=1.67
r256 56 89 0.810901 $w=5.88e-07 $l=4e-08 $layer=LI1_cond $X=10.36 $Y=1.67
+ $X2=10.32 $Y2=1.67
r257 52 54 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=9.18 $Y=2.72
+ $X2=9.18 $Y2=2.99
r258 51 76 45.9078 $w=4.1e-07 $l=1.65e-07 $layer=POLY_cond $X=7.96 $Y=1.58
+ $X2=7.96 $Y2=1.745
r259 51 75 45.9078 $w=4.1e-07 $l=1.65e-07 $layer=POLY_cond $X=7.96 $Y=1.58
+ $X2=7.96 $Y2=1.415
r260 50 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8 $Y=1.58
+ $X2=8 $Y2=1.58
r261 48 69 12.3781 $w=2.68e-07 $l=2.9e-07 $layer=LI1_cond $X=7.89 $Y=1.745
+ $X2=7.89 $Y2=2.035
r262 48 50 3.70415 $w=2.7e-07 $l=1.58e-07 $layer=LI1_cond $X=7.89 $Y=1.745
+ $X2=7.89 $Y2=1.587
r263 46 56 7.7369 $w=1.7e-07 $l=2.95e-07 $layer=LI1_cond $X=10.23 $Y=1.965
+ $X2=10.23 $Y2=1.67
r264 46 47 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=10.23 $Y=1.965
+ $X2=10.23 $Y2=2.905
r265 45 54 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.265 $Y=2.99
+ $X2=9.18 $Y2=2.99
r266 44 47 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.145 $Y=2.99
+ $X2=10.23 $Y2=2.905
r267 44 45 57.4118 $w=1.68e-07 $l=8.8e-07 $layer=LI1_cond $X=10.145 $Y=2.99
+ $X2=9.265 $Y2=2.99
r268 42 52 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.095 $Y=2.72
+ $X2=9.18 $Y2=2.72
r269 42 43 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=9.095 $Y=2.72
+ $X2=8.715 $Y2=2.72
r270 41 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.63 $Y=2.635
+ $X2=8.715 $Y2=2.72
r271 40 41 58.0642 $w=1.68e-07 $l=8.9e-07 $layer=LI1_cond $X=8.63 $Y=1.745
+ $X2=8.63 $Y2=2.635
r272 39 50 3.16494 $w=3.15e-07 $l=1.35e-07 $layer=LI1_cond $X=8.025 $Y=1.587
+ $X2=7.89 $Y2=1.587
r273 38 40 7.64049 $w=3.15e-07 $l=1.95944e-07 $layer=LI1_cond $X=8.545 $Y=1.587
+ $X2=8.63 $Y2=1.745
r274 38 39 19.0245 $w=3.13e-07 $l=5.2e-07 $layer=LI1_cond $X=8.545 $Y=1.587
+ $X2=8.025 $Y2=1.587
r275 33 35 151.266 $w=1.5e-07 $l=2.95e-07 $layer=POLY_cond $X=7.535 $Y=2.46
+ $X2=7.83 $Y2=2.46
r276 31 72 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=3.545 $Y=2.03
+ $X2=3.545 $Y2=1.69
r277 31 32 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.545 $Y=2.03
+ $X2=3.545 $Y2=2.195
r278 30 72 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=3.545 $Y=1.675
+ $X2=3.545 $Y2=1.69
r279 29 30 43.5886 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=3.597 $Y=1.525
+ $X2=3.597 $Y2=1.675
r280 26 80 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=11.055 $Y=0.845
+ $X2=11.055 $Y2=1.295
r281 22 37 466.617 $w=1.5e-07 $l=9.1e-07 $layer=POLY_cond $X=11.03 $Y=2.875
+ $X2=11.03 $Y2=1.965
r282 19 37 48.3131 $w=4.2e-07 $l=2.1e-07 $layer=POLY_cond $X=10.92 $Y=1.755
+ $X2=10.92 $Y2=1.965
r283 18 78 5.95879 $w=4.2e-07 $l=4.5e-08 $layer=POLY_cond $X=10.92 $Y=1.505
+ $X2=10.92 $Y2=1.46
r284 18 19 33.1044 $w=4.2e-07 $l=2.5e-07 $layer=POLY_cond $X=10.92 $Y=1.505
+ $X2=10.92 $Y2=1.755
r285 17 35 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.83 $Y=2.385
+ $X2=7.83 $Y2=2.46
r286 17 76 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=7.83 $Y=2.385
+ $X2=7.83 $Y2=1.745
r287 14 75 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=7.83 $Y=0.845
+ $X2=7.83 $Y2=1.415
r288 9 33 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.535 $Y=2.535
+ $X2=7.535 $Y2=2.46
r289 9 11 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=7.535 $Y=2.535
+ $X2=7.535 $Y2=2.855
r290 7 29 523.021 $w=1.5e-07 $l=1.02e-06 $layer=POLY_cond $X=3.71 $Y=0.505
+ $X2=3.71 $Y2=1.525
r291 3 32 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=3.635 $Y=2.775
+ $X2=3.635 $Y2=2.195
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRTN_1%CLK_N 3 7 9 15 16
c41 3 0 1.50305e-20 $X=4.21 $Y=2.465
r42 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.56
+ $Y=1.51 $X2=4.56 $Y2=1.51
r43 13 15 39.3438 $w=3.3e-07 $l=2.25e-07 $layer=POLY_cond $X=4.335 $Y=1.51
+ $X2=4.56 $Y2=1.51
r44 11 13 21.8577 $w=3.3e-07 $l=1.25e-07 $layer=POLY_cond $X=4.21 $Y=1.51
+ $X2=4.335 $Y2=1.51
r45 9 16 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=4.56 $Y=1.665
+ $X2=4.56 $Y2=1.51
r46 5 13 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.335 $Y=1.345
+ $X2=4.335 $Y2=1.51
r47 5 7 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=4.335 $Y=1.345
+ $X2=4.335 $Y2=0.765
r48 1 11 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.21 $Y=1.675
+ $X2=4.21 $Y2=1.51
r49 1 3 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=4.21 $Y=1.675 $X2=4.21
+ $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRTN_1%A_1080_47# 1 2 9 12 16 20 22 23 27 30 31 32
+ 35 36 37 39 41 42 44 45 48 55 58 59 63 64 68 72 78
c175 63 0 1.9959e-19 $X=9.53 $Y=1.92
c176 32 0 1.98122e-19 $X=7.18 $Y=0.382
c177 12 0 7.01851e-20 $X=6.745 $Y=2.855
r178 64 75 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=9.53 $Y=1.92
+ $X2=9.53 $Y2=2.085
r179 63 64 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.53
+ $Y=1.92 $X2=9.53 $Y2=1.92
r180 60 63 5.76222 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=9.365 $Y=1.92
+ $X2=9.53 $Y2=1.92
r181 58 72 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.625 $Y=0.36
+ $X2=6.625 $Y2=0.525
r182 57 58 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.625
+ $Y=0.36 $X2=6.625 $Y2=0.36
r183 48 50 4.06745 $w=4.23e-07 $l=1.5e-07 $layer=LI1_cond $X=5.607 $Y=1.06
+ $X2=5.607 $Y2=1.21
r184 45 78 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=9.945 $Y=0.36
+ $X2=9.945 $Y2=0.525
r185 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.945
+ $Y=0.36 $X2=9.945 $Y2=0.36
r186 42 44 27.45 $w=1.98e-07 $l=4.95e-07 $layer=LI1_cond $X=9.45 $Y=0.355
+ $X2=9.945 $Y2=0.355
r187 41 60 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.365 $Y=1.755
+ $X2=9.365 $Y2=1.92
r188 40 59 4.27425 $w=2.12e-07 $l=1.04307e-07 $layer=LI1_cond $X=9.365 $Y=0.89
+ $X2=9.322 $Y2=0.805
r189 40 41 56.4332 $w=1.68e-07 $l=8.65e-07 $layer=LI1_cond $X=9.365 $Y=0.89
+ $X2=9.365 $Y2=1.755
r190 39 59 4.27425 $w=2.12e-07 $l=8.5e-08 $layer=LI1_cond $X=9.322 $Y=0.72
+ $X2=9.322 $Y2=0.805
r191 38 42 6.94684 $w=2e-07 $l=1.70833e-07 $layer=LI1_cond $X=9.322 $Y=0.455
+ $X2=9.45 $Y2=0.355
r192 38 39 11.9764 $w=2.53e-07 $l=2.65e-07 $layer=LI1_cond $X=9.322 $Y=0.455
+ $X2=9.322 $Y2=0.72
r193 36 59 2.15711 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=9.195 $Y=0.805
+ $X2=9.322 $Y2=0.805
r194 36 37 120.369 $w=1.68e-07 $l=1.845e-06 $layer=LI1_cond $X=9.195 $Y=0.805
+ $X2=7.35 $Y2=0.805
r195 35 37 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.265 $Y=0.72
+ $X2=7.35 $Y2=0.805
r196 34 35 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=7.265 $Y=0.51
+ $X2=7.265 $Y2=0.72
r197 33 57 2.86415 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=6.63 $Y=0.382
+ $X2=6.545 $Y2=0.382
r198 32 34 7.17723 $w=2.55e-07 $l=1.65118e-07 $layer=LI1_cond $X=7.18 $Y=0.382
+ $X2=7.265 $Y2=0.51
r199 32 33 24.8566 $w=2.53e-07 $l=5.5e-07 $layer=LI1_cond $X=7.18 $Y=0.382
+ $X2=6.63 $Y2=0.382
r200 30 57 4.31308 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=6.545 $Y=0.51
+ $X2=6.545 $Y2=0.382
r201 30 31 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=6.545 $Y=0.51
+ $X2=6.545 $Y2=1.125
r202 28 68 34.9723 $w=3.3e-07 $l=2e-07 $layer=POLY_cond $X=6.545 $Y=1.98
+ $X2=6.745 $Y2=1.98
r203 27 55 13.2445 $w=3.33e-07 $l=3.85e-07 $layer=LI1_cond $X=6.545 $Y=1.982
+ $X2=6.16 $Y2=1.982
r204 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.545
+ $Y=1.98 $X2=6.545 $Y2=1.98
r205 24 50 6.14847 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=5.82 $Y=1.21
+ $X2=5.607 $Y2=1.21
r206 23 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.46 $Y=1.21
+ $X2=6.545 $Y2=1.125
r207 23 24 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=6.46 $Y=1.21
+ $X2=5.82 $Y2=1.21
r208 22 55 15.052 $w=4.43e-07 $l=5.53e-07 $layer=LI1_cond $X=5.607 $Y=2.037
+ $X2=6.16 $Y2=2.037
r209 22 52 1.73514 $w=4.43e-07 $l=6.7e-08 $layer=LI1_cond $X=5.607 $Y=2.037
+ $X2=5.54 $Y2=2.037
r210 21 50 2.30489 $w=4.23e-07 $l=8.5e-08 $layer=LI1_cond $X=5.607 $Y=1.295
+ $X2=5.607 $Y2=1.21
r211 21 22 14.1005 $w=4.23e-07 $l=5.2e-07 $layer=LI1_cond $X=5.607 $Y=1.295
+ $X2=5.607 $Y2=1.815
r212 20 78 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=10.035 $Y=0.845
+ $X2=10.035 $Y2=0.525
r213 16 75 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=9.51 $Y=2.665
+ $X2=9.51 $Y2=2.085
r214 10 68 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.745 $Y=2.145
+ $X2=6.745 $Y2=1.98
r215 10 12 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=6.745 $Y=2.145
+ $X2=6.745 $Y2=2.855
r216 9 72 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=6.68 $Y=0.845
+ $X2=6.68 $Y2=0.525
r217 2 52 600 $w=1.7e-07 $l=3.2249e-07 $layer=licon1_PDIFF $count=1 $X=5.4
+ $Y=1.835 $X2=5.54 $Y2=2.095
r218 1 48 182 $w=1.7e-07 $l=9.43928e-07 $layer=licon1_NDIFF $count=1 $X=5.4
+ $Y=0.235 $X2=5.655 $Y2=1.06
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRTN_1%A_1406_399# 1 2 9 13 17 18 20 21 22 23 24
+ 26
c88 26 0 1.61208e-19 $X=9.295 $Y=2.37
c89 17 0 9.85956e-20 $X=7.38 $Y=1.98
c90 13 0 1.55293e-19 $X=7.47 $Y=0.845
c91 9 0 2.42299e-19 $X=7.105 $Y=2.855
r92 24 26 10.2591 $w=1.98e-07 $l=1.85e-07 $layer=LI1_cond $X=9.11 $Y=2.365
+ $X2=9.295 $Y2=2.365
r93 23 24 6.87494 $w=2e-07 $l=1.36015e-07 $layer=LI1_cond $X=9.025 $Y=2.265
+ $X2=9.11 $Y2=2.365
r94 22 29 3.71618 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=9.025 $Y=1.26 $X2=9.025
+ $Y2=1.16
r95 22 23 65.5668 $w=1.68e-07 $l=1.005e-06 $layer=LI1_cond $X=9.025 $Y=1.26
+ $X2=9.025 $Y2=2.265
r96 20 29 3.15876 $w=2e-07 $l=8.5e-08 $layer=LI1_cond $X=8.94 $Y=1.16 $X2=9.025
+ $Y2=1.16
r97 20 21 77.3591 $w=1.98e-07 $l=1.395e-06 $layer=LI1_cond $X=8.94 $Y=1.16
+ $X2=7.545 $Y2=1.16
r98 18 32 13.7278 $w=3.16e-07 $l=9e-08 $layer=POLY_cond $X=7.38 $Y=1.98 $X2=7.47
+ $Y2=1.98
r99 18 30 41.9462 $w=3.16e-07 $l=2.75e-07 $layer=POLY_cond $X=7.38 $Y=1.98
+ $X2=7.105 $Y2=1.98
r100 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.38
+ $Y=1.98 $X2=7.38 $Y2=1.98
r101 15 21 7.36389 $w=2e-07 $l=2.09105e-07 $layer=LI1_cond $X=7.38 $Y=1.26
+ $X2=7.545 $Y2=1.16
r102 15 17 25.1442 $w=3.28e-07 $l=7.2e-07 $layer=LI1_cond $X=7.38 $Y=1.26
+ $X2=7.38 $Y2=1.98
r103 11 32 20.1942 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.47 $Y=1.815
+ $X2=7.47 $Y2=1.98
r104 11 13 497.383 $w=1.5e-07 $l=9.7e-07 $layer=POLY_cond $X=7.47 $Y=1.815
+ $X2=7.47 $Y2=0.845
r105 7 30 20.1942 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.105 $Y=2.145
+ $X2=7.105 $Y2=1.98
r106 7 9 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=7.105 $Y=2.145
+ $X2=7.105 $Y2=2.855
r107 2 26 600 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=9.155
+ $Y=2.245 $X2=9.295 $Y2=2.37
r108 1 29 182 $w=1.7e-07 $l=6.34823e-07 $layer=licon1_NDIFF $count=1 $X=8.69
+ $Y=0.635 $X2=8.945 $Y2=1.155
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRTN_1%A_1278_529# 1 2 3 12 14 15 16 18 25 29 35
+ 36 41 44 48
c114 48 0 1.90325e-19 $X=8.285 $Y=2.685
r115 46 48 0.0892596 $w=6.68e-07 $l=5e-09 $layer=LI1_cond $X=8.28 $Y=2.685
+ $X2=8.285 $Y2=2.685
r116 46 47 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.28
+ $Y=2.49 $X2=8.28 $Y2=2.49
r117 43 46 9.46152 $w=6.68e-07 $l=5.3e-07 $layer=LI1_cond $X=7.75 $Y=2.685
+ $X2=8.28 $Y2=2.685
r118 43 44 9.89763 $w=6.68e-07 $l=1.25e-07 $layer=LI1_cond $X=7.75 $Y=2.685
+ $X2=7.625 $Y2=2.685
r119 41 44 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=7 $Y=2.435
+ $X2=7.625 $Y2=2.435
r120 40 41 5.8268 $w=1.98e-07 $l=1e-07 $layer=LI1_cond $X=6.9 $Y=2.42 $X2=7
+ $Y2=2.42
r121 36 47 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=8.28 $Y=2.15
+ $X2=8.28 $Y2=2.49
r122 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.28
+ $Y=2.15 $X2=8.28 $Y2=2.15
r123 33 48 8.66103 $w=1.8e-07 $l=3.35e-07 $layer=LI1_cond $X=8.285 $Y=2.35
+ $X2=8.285 $Y2=2.685
r124 33 35 12.3232 $w=1.78e-07 $l=2e-07 $layer=LI1_cond $X=8.285 $Y=2.35
+ $X2=8.285 $Y2=2.15
r125 27 40 0.716491 $w=2e-07 $l=1e-07 $layer=LI1_cond $X=6.9 $Y=2.32 $X2=6.9
+ $Y2=2.42
r126 27 29 81.7955 $w=1.98e-07 $l=1.475e-06 $layer=LI1_cond $X=6.9 $Y=2.32
+ $X2=6.9 $Y2=0.845
r127 23 40 19.4091 $w=1.98e-07 $l=3.5e-07 $layer=LI1_cond $X=6.55 $Y=2.42
+ $X2=6.9 $Y2=2.42
r128 23 25 13.3127 $w=2.88e-07 $l=3.35e-07 $layer=LI1_cond $X=6.55 $Y=2.52
+ $X2=6.55 $Y2=2.855
r129 20 36 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=8.28 $Y=2.135
+ $X2=8.28 $Y2=2.15
r130 20 22 171.777 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=8.28 $Y=2.06
+ $X2=8.615 $Y2=2.06
r131 16 18 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=9.08 $Y=2.135
+ $X2=9.08 $Y2=2.665
r132 15 22 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.69 $Y=2.06
+ $X2=8.615 $Y2=2.06
r133 14 16 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.005 $Y=2.06
+ $X2=9.08 $Y2=2.135
r134 14 15 161.521 $w=1.5e-07 $l=3.15e-07 $layer=POLY_cond $X=9.005 $Y=2.06
+ $X2=8.69 $Y2=2.06
r135 10 22 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.615 $Y=1.985
+ $X2=8.615 $Y2=2.06
r136 10 12 528.149 $w=1.5e-07 $l=1.03e-06 $layer=POLY_cond $X=8.615 $Y=1.985
+ $X2=8.615 $Y2=0.955
r137 3 43 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=7.61
+ $Y=2.645 $X2=7.75 $Y2=2.855
r138 2 25 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=6.39
+ $Y=2.645 $X2=6.53 $Y2=2.855
r139 1 29 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=6.755
+ $Y=0.635 $X2=6.895 $Y2=0.845
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRTN_1%A_857_367# 1 2 9 13 15 18 19 21 23 27 28 29
+ 33 34 35 38 40 43 45 49 56 61
c152 43 0 1.16957e-19 $X=6.315 $Y=2.46
c153 38 0 1.61208e-19 $X=10.035 $Y=2.875
c154 29 0 4.28297e-20 $X=7.185 $Y=0.18
r155 60 61 30.474 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=5.325 $Y=1.46
+ $X2=5.4 $Y2=1.46
r156 57 60 34.0979 $w=3.3e-07 $l=1.95e-07 $layer=POLY_cond $X=5.13 $Y=1.46
+ $X2=5.325 $Y2=1.46
r157 56 57 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.13
+ $Y=1.46 $X2=5.13 $Y2=1.46
r158 54 56 30.6631 $w=1.68e-07 $l=4.7e-07 $layer=LI1_cond $X=5.13 $Y=1.93
+ $X2=5.13 $Y2=1.46
r159 53 56 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=5.13 $Y=1.165
+ $X2=5.13 $Y2=1.46
r160 49 53 6.87494 $w=2e-07 $l=1.36015e-07 $layer=LI1_cond $X=5.045 $Y=1.065
+ $X2=5.13 $Y2=1.165
r161 49 51 27.45 $w=1.98e-07 $l=4.95e-07 $layer=LI1_cond $X=5.045 $Y=1.065
+ $X2=4.55 $Y2=1.065
r162 45 54 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.045 $Y=2.095
+ $X2=5.13 $Y2=1.93
r163 45 47 21.652 $w=3.28e-07 $l=6.2e-07 $layer=LI1_cond $X=5.045 $Y=2.095
+ $X2=4.425 $Y2=2.095
r164 41 43 128.191 $w=1.5e-07 $l=2.5e-07 $layer=POLY_cond $X=6.065 $Y=2.46
+ $X2=6.315 $Y2=2.46
r165 36 38 681.979 $w=1.5e-07 $l=1.33e-06 $layer=POLY_cond $X=10.035 $Y=1.545
+ $X2=10.035 $Y2=2.875
r166 34 36 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.96 $Y=1.47
+ $X2=10.035 $Y2=1.545
r167 34 35 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=9.96 $Y=1.47
+ $X2=9.35 $Y2=1.47
r168 31 35 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.275 $Y=1.395
+ $X2=9.35 $Y2=1.47
r169 31 33 225.617 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=9.275 $Y=1.395
+ $X2=9.275 $Y2=0.955
r170 30 33 358.936 $w=1.5e-07 $l=7e-07 $layer=POLY_cond $X=9.275 $Y=0.255
+ $X2=9.275 $Y2=0.955
r171 28 30 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.2 $Y=0.18
+ $X2=9.275 $Y2=0.255
r172 28 29 1033.22 $w=1.5e-07 $l=2.015e-06 $layer=POLY_cond $X=9.2 $Y=0.18
+ $X2=7.185 $Y2=0.18
r173 25 27 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=7.11 $Y=1.425
+ $X2=7.11 $Y2=0.845
r174 24 29 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.11 $Y=0.255
+ $X2=7.185 $Y2=0.18
r175 24 27 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=7.11 $Y=0.255
+ $X2=7.11 $Y2=0.845
r176 21 43 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.315 $Y=2.535
+ $X2=6.315 $Y2=2.46
r177 21 23 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=6.315 $Y=2.535
+ $X2=6.315 $Y2=2.855
r178 20 40 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.14 $Y=1.5
+ $X2=6.065 $Y2=1.5
r179 19 25 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.035 $Y=1.5
+ $X2=7.11 $Y2=1.425
r180 19 20 458.926 $w=1.5e-07 $l=8.95e-07 $layer=POLY_cond $X=7.035 $Y=1.5
+ $X2=6.14 $Y2=1.5
r181 18 41 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.065 $Y=2.385
+ $X2=6.065 $Y2=2.46
r182 17 40 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.065 $Y=1.575
+ $X2=6.065 $Y2=1.5
r183 17 18 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=6.065 $Y=1.575
+ $X2=6.065 $Y2=2.385
r184 15 40 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.99 $Y=1.5
+ $X2=6.065 $Y2=1.5
r185 15 61 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=5.99 $Y=1.5 $X2=5.4
+ $Y2=1.5
r186 11 60 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.325 $Y=1.625
+ $X2=5.325 $Y2=1.46
r187 11 13 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=5.325 $Y=1.625
+ $X2=5.325 $Y2=2.465
r188 7 60 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.325 $Y=1.295
+ $X2=5.325 $Y2=1.46
r189 7 9 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=5.325 $Y=1.295
+ $X2=5.325 $Y2=0.655
r190 2 47 600 $w=1.7e-07 $l=3.2249e-07 $layer=licon1_PDIFF $count=1 $X=4.285
+ $Y=1.835 $X2=4.425 $Y2=2.095
r191 1 51 182 $w=1.7e-07 $l=7.81873e-07 $layer=licon1_NDIFF $count=1 $X=4.41
+ $Y=0.345 $X2=4.55 $Y2=1.06
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRTN_1%A_2064_101# 1 2 9 13 15 18 22 25 26 27 28
+ 33 34
c91 33 0 3.32213e-20 $X=11.855 $Y=1.795
c92 28 0 4.6212e-20 $X=11.77 $Y=0.725
r93 32 33 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=11.855 $Y=0.855
+ $X2=11.855 $Y2=1.795
r94 28 32 7.21222 $w=2.6e-07 $l=1.67183e-07 $layer=LI1_cond $X=11.77 $Y=0.725
+ $X2=11.855 $Y2=0.855
r95 28 30 6.20546 $w=2.58e-07 $l=1.4e-07 $layer=LI1_cond $X=11.77 $Y=0.725
+ $X2=11.63 $Y2=0.725
r96 26 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=11.77 $Y=1.88
+ $X2=11.855 $Y2=1.795
r97 26 27 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=11.77 $Y=1.88
+ $X2=11.39 $Y2=1.88
r98 25 34 6.7841 $w=2.35e-07 $l=1.96914e-07 $layer=LI1_cond $X=11.305 $Y=2.175
+ $X2=11.235 $Y2=2.34
r99 24 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=11.305 $Y=1.965
+ $X2=11.39 $Y2=1.88
r100 24 25 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=11.305 $Y=1.965
+ $X2=11.305 $Y2=2.175
r101 20 34 6.7841 $w=2.35e-07 $l=1.67481e-07 $layer=LI1_cond $X=11.23 $Y=2.505
+ $X2=11.235 $Y2=2.34
r102 20 22 14.2135 $w=2.98e-07 $l=3.7e-07 $layer=LI1_cond $X=11.23 $Y=2.505
+ $X2=11.23 $Y2=2.875
r103 18 35 32.3493 $w=3.3e-07 $l=1.85e-07 $layer=POLY_cond $X=10.58 $Y=2.34
+ $X2=10.395 $Y2=2.34
r104 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.58
+ $Y=2.34 $X2=10.58 $Y2=2.34
r105 15 34 0.153733 $w=3.3e-07 $l=1.55e-07 $layer=LI1_cond $X=11.08 $Y=2.34
+ $X2=11.235 $Y2=2.34
r106 15 17 17.4613 $w=3.28e-07 $l=5e-07 $layer=LI1_cond $X=11.08 $Y=2.34
+ $X2=10.58 $Y2=2.34
r107 11 35 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.395 $Y=2.505
+ $X2=10.395 $Y2=2.34
r108 11 13 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=10.395 $Y=2.505
+ $X2=10.395 $Y2=2.875
r109 7 35 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.395 $Y=2.175
+ $X2=10.395 $Y2=2.34
r110 7 9 681.979 $w=1.5e-07 $l=1.33e-06 $layer=POLY_cond $X=10.395 $Y=2.175
+ $X2=10.395 $Y2=0.845
r111 2 22 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=11.105
+ $Y=2.665 $X2=11.245 $Y2=2.875
r112 1 30 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=11.49
+ $Y=0.635 $X2=11.63 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRTN_1%A_1870_127# 1 2 9 12 14 17 20 22 24 27 29
+ 32 35 36 40 43 47 49 50
c125 43 0 1.9959e-19 $X=9.792 $Y=1.16
c126 27 0 4.6212e-20 $X=12.44 $Y=0.92
c127 12 0 1.69115e-19 $X=11.46 $Y=2.875
r128 49 50 30.474 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=11.505 $Y=1.24
+ $X2=11.505 $Y2=1.165
r129 45 47 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=9.725 $Y=2.57
+ $X2=9.88 $Y2=2.57
r130 41 52 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=11.505 $Y=1.33
+ $X2=11.505 $Y2=1.495
r131 41 49 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=11.505 $Y=1.33
+ $X2=11.505 $Y2=1.24
r132 40 41 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.505
+ $Y=1.33 $X2=11.505 $Y2=1.33
r133 38 40 5.54059 $w=2.58e-07 $l=1.25e-07 $layer=LI1_cond $X=11.47 $Y=1.205
+ $X2=11.47 $Y2=1.33
r134 37 43 2.65845 $w=1.8e-07 $l=1.94201e-07 $layer=LI1_cond $X=9.965 $Y=1.115
+ $X2=9.792 $Y2=1.16
r135 36 38 7.11373 $w=1.8e-07 $l=1.69115e-07 $layer=LI1_cond $X=11.34 $Y=1.115
+ $X2=11.47 $Y2=1.205
r136 36 37 84.7222 $w=1.78e-07 $l=1.375e-06 $layer=LI1_cond $X=11.34 $Y=1.115
+ $X2=9.965 $Y2=1.115
r137 35 47 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.88 $Y=2.405
+ $X2=9.88 $Y2=2.57
r138 34 43 3.7989 $w=2.57e-07 $l=1.73508e-07 $layer=LI1_cond $X=9.88 $Y=1.295
+ $X2=9.792 $Y2=1.16
r139 34 35 72.4171 $w=1.68e-07 $l=1.11e-06 $layer=LI1_cond $X=9.88 $Y=1.295
+ $X2=9.88 $Y2=2.405
r140 30 43 3.7989 $w=2.57e-07 $l=1.35e-07 $layer=LI1_cond $X=9.792 $Y=1.025
+ $X2=9.792 $Y2=1.16
r141 30 32 7.84997 $w=3.43e-07 $l=2.35e-07 $layer=LI1_cond $X=9.792 $Y=1.025
+ $X2=9.792 $Y2=0.79
r142 25 27 128.191 $w=1.5e-07 $l=2.5e-07 $layer=POLY_cond $X=12.19 $Y=0.92
+ $X2=12.44 $Y2=0.92
r143 22 27 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=12.44 $Y=0.845
+ $X2=12.44 $Y2=0.92
r144 22 24 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=12.44 $Y=0.845
+ $X2=12.44 $Y2=0.525
r145 18 29 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=12.19 $Y=1.315
+ $X2=12.19 $Y2=1.24
r146 18 20 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=12.19 $Y=1.315
+ $X2=12.19 $Y2=2.075
r147 17 29 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=12.19 $Y=1.165
+ $X2=12.19 $Y2=1.24
r148 16 25 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=12.19 $Y=0.995
+ $X2=12.19 $Y2=0.92
r149 16 17 87.1702 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=12.19 $Y=0.995
+ $X2=12.19 $Y2=1.165
r150 15 49 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=11.67 $Y=1.24
+ $X2=11.505 $Y2=1.24
r151 14 29 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=12.115 $Y=1.24
+ $X2=12.19 $Y2=1.24
r152 14 15 228.181 $w=1.5e-07 $l=4.45e-07 $layer=POLY_cond $X=12.115 $Y=1.24
+ $X2=11.67 $Y2=1.24
r153 12 52 707.617 $w=1.5e-07 $l=1.38e-06 $layer=POLY_cond $X=11.46 $Y=2.875
+ $X2=11.46 $Y2=1.495
r154 9 50 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=11.415 $Y=0.845
+ $X2=11.415 $Y2=1.165
r155 2 45 600 $w=1.7e-07 $l=3.88748e-07 $layer=licon1_PDIFF $count=1 $X=9.585
+ $Y=2.245 $X2=9.725 $Y2=2.57
r156 1 32 91 $w=1.7e-07 $l=4.255e-07 $layer=licon1_NDIFF $count=2 $X=9.35
+ $Y=0.635 $X2=9.705 $Y2=0.79
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRTN_1%A_2370_351# 1 2 9 13 14 20 23 26 27 29 31
c60 23 0 1.69115e-19 $X=12.195 $Y=2.135
r61 27 32 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=12.852 $Y=1.43
+ $X2=12.852 $Y2=1.595
r62 27 31 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=12.852 $Y=1.43
+ $X2=12.852 $Y2=1.265
r63 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=12.83
+ $Y=1.43 $X2=12.83 $Y2=1.43
r64 24 29 0.261258 $w=3.3e-07 $l=1.23e-07 $layer=LI1_cond $X=12.355 $Y=1.43
+ $X2=12.232 $Y2=1.43
r65 24 26 16.5882 $w=3.28e-07 $l=4.75e-07 $layer=LI1_cond $X=12.355 $Y=1.43
+ $X2=12.83 $Y2=1.43
r66 22 29 7.45506 $w=2.07e-07 $l=1.82565e-07 $layer=LI1_cond $X=12.195 $Y=1.595
+ $X2=12.232 $Y2=1.43
r67 22 23 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=12.195 $Y=1.595
+ $X2=12.195 $Y2=2.135
r68 18 29 7.45506 $w=2.07e-07 $l=1.65e-07 $layer=LI1_cond $X=12.232 $Y=1.265
+ $X2=12.232 $Y2=1.43
r69 18 20 35.2789 $w=2.43e-07 $l=7.5e-07 $layer=LI1_cond $X=12.232 $Y=1.265
+ $X2=12.232 $Y2=0.515
r70 14 23 7.36005 $w=2.8e-07 $l=1.77482e-07 $layer=LI1_cond $X=12.11 $Y=2.275
+ $X2=12.195 $Y2=2.135
r71 14 16 5.55642 $w=2.78e-07 $l=1.35e-07 $layer=LI1_cond $X=12.11 $Y=2.275
+ $X2=11.975 $Y2=2.275
r72 13 31 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=12.965 $Y=0.735
+ $X2=12.965 $Y2=1.265
r73 9 32 446.106 $w=1.5e-07 $l=8.7e-07 $layer=POLY_cond $X=12.81 $Y=2.465
+ $X2=12.81 $Y2=1.595
r74 2 16 600 $w=1.7e-07 $l=5.53986e-07 $layer=licon1_PDIFF $count=1 $X=11.85
+ $Y=1.755 $X2=11.975 $Y2=2.25
r75 1 20 182 $w=1.7e-07 $l=2.54951e-07 $layer=licon1_NDIFF $count=1 $X=12.1
+ $Y=0.315 $X2=12.225 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRTN_1%VPWR 1 2 3 4 5 6 7 8 9 28 30 34 38 42 46 50
+ 52 55 58 61 62 64 65 67 68 71 72 73 90 94 102 118 119 126 132 134 137 140
c173 119 0 1.16957e-19 $X=13.2 $Y=3.33
r174 143 144 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r175 140 143 9.07985 $w=3.28e-07 $l=2.6e-07 $layer=LI1_cond $X=8.75 $Y=3.07
+ $X2=8.75 $Y2=3.33
r176 137 138 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r177 134 135 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r178 131 132 9.2801 $w=4.58e-07 $l=1.65e-07 $layer=LI1_cond $X=2.46 $Y=3.185
+ $X2=2.625 $Y2=3.185
r179 128 131 7.80051 $w=4.58e-07 $l=3e-07 $layer=LI1_cond $X=2.16 $Y=3.185
+ $X2=2.46 $Y2=3.185
r180 128 129 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r181 125 128 1.04007 $w=4.58e-07 $l=4e-08 $layer=LI1_cond $X=2.12 $Y=3.185
+ $X2=2.16 $Y2=3.185
r182 125 126 9.2801 $w=4.58e-07 $l=1.65e-07 $layer=LI1_cond $X=2.12 $Y=3.185
+ $X2=1.955 $Y2=3.185
r183 122 123 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r184 118 119 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=13.2 $Y=3.33
+ $X2=13.2 $Y2=3.33
r185 116 119 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=12.24 $Y=3.33
+ $X2=13.2 $Y2=3.33
r186 115 116 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=12.24 $Y=3.33
+ $X2=12.24 $Y2=3.33
r187 113 116 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=11.28 $Y=3.33
+ $X2=12.24 $Y2=3.33
r188 112 113 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.28 $Y=3.33
+ $X2=11.28 $Y2=3.33
r189 110 113 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=10.32 $Y=3.33
+ $X2=11.28 $Y2=3.33
r190 110 144 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=10.32 $Y=3.33
+ $X2=8.88 $Y2=3.33
r191 109 110 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.32 $Y=3.33
+ $X2=10.32 $Y2=3.33
r192 107 143 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.915 $Y=3.33
+ $X2=8.75 $Y2=3.33
r193 107 109 91.6631 $w=1.68e-07 $l=1.405e-06 $layer=LI1_cond $X=8.915 $Y=3.33
+ $X2=10.32 $Y2=3.33
r194 106 144 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=8.88 $Y2=3.33
r195 106 138 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=7.44 $Y2=3.33
r196 105 106 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r197 103 137 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=7.455 $Y=3.33
+ $X2=7.305 $Y2=3.33
r198 103 105 61.6524 $w=1.68e-07 $l=9.45e-07 $layer=LI1_cond $X=7.455 $Y=3.33
+ $X2=8.4 $Y2=3.33
r199 102 143 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.585 $Y=3.33
+ $X2=8.75 $Y2=3.33
r200 102 105 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=8.585 $Y=3.33
+ $X2=8.4 $Y2=3.33
r201 101 138 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=7.44 $Y2=3.33
r202 100 101 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r203 98 135 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=5.04 $Y2=3.33
r204 97 100 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=5.52 $Y=3.33
+ $X2=6.96 $Y2=3.33
r205 97 98 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r206 95 134 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.275 $Y=3.33
+ $X2=5.11 $Y2=3.33
r207 95 97 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=5.275 $Y=3.33
+ $X2=5.52 $Y2=3.33
r208 94 137 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=7.155 $Y=3.33
+ $X2=7.305 $Y2=3.33
r209 94 100 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=7.155 $Y=3.33
+ $X2=6.96 $Y2=3.33
r210 93 135 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.04 $Y2=3.33
r211 92 93 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r212 90 134 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.945 $Y=3.33
+ $X2=5.11 $Y2=3.33
r213 90 92 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=4.945 $Y=3.33
+ $X2=4.56 $Y2=3.33
r214 89 93 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.56 $Y2=3.33
r215 88 89 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r216 86 89 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r217 86 129 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r218 85 88 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.64 $Y=3.33 $X2=3.6
+ $Y2=3.33
r219 85 132 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=2.64 $Y=3.33
+ $X2=2.625 $Y2=3.33
r220 85 86 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r221 82 129 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r222 81 126 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=1.68 $Y=3.33
+ $X2=1.955 $Y2=3.33
r223 81 82 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r224 79 82 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r225 79 123 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r226 78 81 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r227 78 79 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r228 76 122 4.42547 $w=1.7e-07 $l=2.03e-07 $layer=LI1_cond $X=0.405 $Y=3.33
+ $X2=0.202 $Y2=3.33
r229 76 78 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.405 $Y=3.33
+ $X2=0.72 $Y2=3.33
r230 73 101 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=6.72 $Y=3.33
+ $X2=6.96 $Y2=3.33
r231 73 98 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=6.72 $Y=3.33
+ $X2=5.52 $Y2=3.33
r232 71 115 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=12.37 $Y=3.33
+ $X2=12.24 $Y2=3.33
r233 71 72 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=12.37 $Y=3.33
+ $X2=12.54 $Y2=3.33
r234 70 118 31.9679 $w=1.68e-07 $l=4.9e-07 $layer=LI1_cond $X=12.71 $Y=3.33
+ $X2=13.2 $Y2=3.33
r235 70 72 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=12.71 $Y=3.33
+ $X2=12.54 $Y2=3.33
r236 67 112 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=11.55 $Y=3.33
+ $X2=11.28 $Y2=3.33
r237 67 68 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=11.55 $Y=3.33
+ $X2=11.695 $Y2=3.33
r238 66 115 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=11.84 $Y=3.33
+ $X2=12.24 $Y2=3.33
r239 66 68 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=11.84 $Y=3.33
+ $X2=11.695 $Y2=3.33
r240 64 109 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=10.54 $Y=3.33
+ $X2=10.32 $Y2=3.33
r241 64 65 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.54 $Y=3.33
+ $X2=10.705 $Y2=3.33
r242 63 112 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=10.87 $Y=3.33
+ $X2=11.28 $Y2=3.33
r243 63 65 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.87 $Y=3.33
+ $X2=10.705 $Y2=3.33
r244 61 88 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=3.755 $Y=3.33
+ $X2=3.6 $Y2=3.33
r245 61 62 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.755 $Y=3.33
+ $X2=3.92 $Y2=3.33
r246 60 92 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=4.085 $Y=3.33
+ $X2=4.56 $Y2=3.33
r247 60 62 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.085 $Y=3.33
+ $X2=3.92 $Y2=3.33
r248 58 69 27.703 $w=2.58e-07 $l=6.25e-07 $layer=LI1_cond $X=12.58 $Y=1.96
+ $X2=12.58 $Y2=2.585
r249 53 72 0.987631 $w=3.4e-07 $l=8.5e-08 $layer=LI1_cond $X=12.54 $Y=3.245
+ $X2=12.54 $Y2=3.33
r250 53 55 9.99914 $w=3.38e-07 $l=2.95e-07 $layer=LI1_cond $X=12.54 $Y=3.245
+ $X2=12.54 $Y2=2.95
r251 52 69 6.42894 $w=3.38e-07 $l=1.7e-07 $layer=LI1_cond $X=12.54 $Y=2.755
+ $X2=12.54 $Y2=2.585
r252 52 55 6.6096 $w=3.38e-07 $l=1.95e-07 $layer=LI1_cond $X=12.54 $Y=2.755
+ $X2=12.54 $Y2=2.95
r253 48 68 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=11.695 $Y=3.245
+ $X2=11.695 $Y2=3.33
r254 48 50 14.7036 $w=2.88e-07 $l=3.7e-07 $layer=LI1_cond $X=11.695 $Y=3.245
+ $X2=11.695 $Y2=2.875
r255 44 65 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.705 $Y=3.245
+ $X2=10.705 $Y2=3.33
r256 44 46 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=10.705 $Y=3.245
+ $X2=10.705 $Y2=2.875
r257 40 137 0.597483 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.305 $Y=3.245
+ $X2=7.305 $Y2=3.33
r258 40 42 14.9818 $w=2.98e-07 $l=3.9e-07 $layer=LI1_cond $X=7.305 $Y=3.245
+ $X2=7.305 $Y2=2.855
r259 36 134 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.11 $Y=3.245
+ $X2=5.11 $Y2=3.33
r260 36 38 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=5.11 $Y=3.245
+ $X2=5.11 $Y2=2.88
r261 32 62 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.92 $Y=3.245
+ $X2=3.92 $Y2=3.33
r262 32 34 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=3.92 $Y=3.245
+ $X2=3.92 $Y2=2.88
r263 28 122 3.05205 $w=2.95e-07 $l=1.09087e-07 $layer=LI1_cond $X=0.257 $Y=3.245
+ $X2=0.202 $Y2=3.33
r264 28 30 49.4183 $w=2.93e-07 $l=1.265e-06 $layer=LI1_cond $X=0.257 $Y=3.245
+ $X2=0.257 $Y2=1.98
r265 9 58 300 $w=1.7e-07 $l=3.5812e-07 $layer=licon1_PDIFF $count=2 $X=12.265
+ $Y=1.755 $X2=12.535 $Y2=1.96
r266 9 55 600 $w=1.7e-07 $l=1.32313e-06 $layer=licon1_PDIFF $count=1 $X=12.265
+ $Y=1.755 $X2=12.535 $Y2=2.95
r267 8 50 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=11.535
+ $Y=2.665 $X2=11.675 $Y2=2.875
r268 7 46 600 $w=1.7e-07 $l=3.23381e-07 $layer=licon1_PDIFF $count=1 $X=10.47
+ $Y=2.665 $X2=10.705 $Y2=2.875
r269 6 140 600 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=8.605
+ $Y=2.245 $X2=8.75 $Y2=3.07
r270 5 42 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=7.18
+ $Y=2.645 $X2=7.32 $Y2=2.855
r271 4 38 600 $w=1.7e-07 $l=1.10574e-06 $layer=licon1_PDIFF $count=1 $X=4.985
+ $Y=1.835 $X2=5.11 $Y2=2.88
r272 3 34 600 $w=1.7e-07 $l=5.19495e-07 $layer=licon1_PDIFF $count=1 $X=3.71
+ $Y=2.455 $X2=3.92 $Y2=2.88
r273 2 131 600 $w=1.7e-07 $l=8.11249e-07 $layer=licon1_PDIFF $count=1 $X=1.92
+ $Y=2.455 $X2=2.46 $Y2=3.04
r274 2 125 600 $w=1.7e-07 $l=6.77661e-07 $layer=licon1_PDIFF $count=1 $X=1.92
+ $Y=2.455 $X2=2.12 $Y2=3.04
r275 1 30 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.15
+ $Y=1.835 $X2=0.275 $Y2=1.98
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRTN_1%A_229_491# 1 2 3 4 5 16 18 20 23 24 26 30
+ 32 40 41 47 48 49
c146 47 0 1.86933e-19 $X=3.95 $Y=0.74
c147 41 0 1.50305e-20 $X=3.36 $Y=2.482
c148 26 0 7.01851e-20 $X=5.915 $Y=2.515
r149 49 52 3.68782 $w=2.48e-07 $l=8e-08 $layer=LI1_cond $X=6.165 $Y=0.71
+ $X2=6.165 $Y2=0.79
r150 44 45 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=3.36 $Y=2.62 $X2=3.36
+ $Y2=2.7
r151 41 44 4.81931 $w=3.28e-07 $l=1.38e-07 $layer=LI1_cond $X=3.36 $Y=2.482
+ $X2=3.36 $Y2=2.62
r152 38 40 8.79328 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=2.42 $Y=0.73
+ $X2=2.585 $Y2=0.73
r153 32 35 3.49225 $w=3.28e-07 $l=1e-07 $layer=LI1_cond $X=1.27 $Y=2.7 $X2=1.27
+ $Y2=2.8
r154 28 30 9.18353 $w=3.18e-07 $l=2.55e-07 $layer=LI1_cond $X=6.075 $Y=2.6
+ $X2=6.075 $Y2=2.855
r155 27 48 4.45556 $w=2.02e-07 $l=1.0015e-07 $layer=LI1_cond $X=4.035 $Y=2.515
+ $X2=3.95 $Y2=2.482
r156 26 28 7.68211 $w=1.7e-07 $l=1.9799e-07 $layer=LI1_cond $X=5.915 $Y=2.515
+ $X2=6.075 $Y2=2.6
r157 26 27 122.652 $w=1.68e-07 $l=1.88e-06 $layer=LI1_cond $X=5.915 $Y=2.515
+ $X2=4.035 $Y2=2.515
r158 25 47 5.16603 $w=1.7e-07 $l=9.88686e-08 $layer=LI1_cond $X=4.035 $Y=0.71
+ $X2=3.95 $Y2=0.74
r159 24 49 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.04 $Y=0.71
+ $X2=6.165 $Y2=0.71
r160 24 25 130.807 $w=1.68e-07 $l=2.005e-06 $layer=LI1_cond $X=6.04 $Y=0.71
+ $X2=4.035 $Y2=0.71
r161 23 48 1.97946 $w=1.7e-07 $l=1.17e-07 $layer=LI1_cond $X=3.95 $Y=2.365
+ $X2=3.95 $Y2=2.482
r162 22 47 1.34256 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=3.95 $Y=0.855
+ $X2=3.95 $Y2=0.74
r163 22 23 98.5134 $w=1.68e-07 $l=1.51e-06 $layer=LI1_cond $X=3.95 $Y=0.855
+ $X2=3.95 $Y2=2.365
r164 21 41 2.74472 $w=2.35e-07 $l=1.65e-07 $layer=LI1_cond $X=3.525 $Y=2.482
+ $X2=3.36 $Y2=2.482
r165 20 48 4.45556 $w=2.02e-07 $l=8.5e-08 $layer=LI1_cond $X=3.865 $Y=2.482
+ $X2=3.95 $Y2=2.482
r166 20 21 16.6736 $w=2.33e-07 $l=3.4e-07 $layer=LI1_cond $X=3.865 $Y=2.482
+ $X2=3.525 $Y2=2.482
r167 18 47 5.16603 $w=1.7e-07 $l=9.88686e-08 $layer=LI1_cond $X=3.865 $Y=0.77
+ $X2=3.95 $Y2=0.74
r168 18 40 83.508 $w=1.68e-07 $l=1.28e-06 $layer=LI1_cond $X=3.865 $Y=0.77
+ $X2=2.585 $Y2=0.77
r169 17 32 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.435 $Y=2.7
+ $X2=1.27 $Y2=2.7
r170 16 45 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.195 $Y=2.7
+ $X2=3.36 $Y2=2.7
r171 16 17 114.824 $w=1.68e-07 $l=1.76e-06 $layer=LI1_cond $X=3.195 $Y=2.7
+ $X2=1.435 $Y2=2.7
r172 5 30 600 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=1 $X=5.955
+ $Y=2.645 $X2=6.1 $Y2=2.855
r173 4 44 300 $w=1.7e-07 $l=2.59711e-07 $layer=licon1_PDIFF $count=2 $X=3.17
+ $Y=2.455 $X2=3.36 $Y2=2.62
r174 3 35 600 $w=1.7e-07 $l=4.02679e-07 $layer=licon1_PDIFF $count=1 $X=1.145
+ $Y=2.455 $X2=1.27 $Y2=2.8
r175 2 52 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=6.07
+ $Y=0.635 $X2=6.205 $Y2=0.79
r176 1 38 182 $w=1.7e-07 $l=5.17011e-07 $layer=licon1_NDIFF $count=1 $X=2.165
+ $Y=0.295 $X2=2.42 $Y2=0.7
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRTN_1%Q 1 2 7 8 9 10 11 12 13 24 44 48
r19 44 45 6.55033 $w=4.63e-07 $l=1.65e-07 $layer=LI1_cond $X=13.112 $Y=1.98
+ $X2=13.112 $Y2=1.815
r20 34 48 0.308665 $w=4.63e-07 $l=1.2e-08 $layer=LI1_cond $X=13.112 $Y=2.047
+ $X2=13.112 $Y2=2.035
r21 13 41 3.47249 $w=4.63e-07 $l=1.35e-07 $layer=LI1_cond $X=13.112 $Y=2.775
+ $X2=13.112 $Y2=2.91
r22 12 13 9.51718 $w=4.63e-07 $l=3.7e-07 $layer=LI1_cond $X=13.112 $Y=2.405
+ $X2=13.112 $Y2=2.775
r23 11 48 0.951718 $w=4.63e-07 $l=3.7e-08 $layer=LI1_cond $X=13.112 $Y=1.998
+ $X2=13.112 $Y2=2.035
r24 11 44 0.462998 $w=4.63e-07 $l=1.8e-08 $layer=LI1_cond $X=13.112 $Y=1.998
+ $X2=13.112 $Y2=1.98
r25 11 12 8.28252 $w=4.63e-07 $l=3.22e-07 $layer=LI1_cond $X=13.112 $Y=2.083
+ $X2=13.112 $Y2=2.405
r26 11 34 0.925996 $w=4.63e-07 $l=3.6e-08 $layer=LI1_cond $X=13.112 $Y=2.083
+ $X2=13.112 $Y2=2.047
r27 10 45 6.64871 $w=2.58e-07 $l=1.5e-07 $layer=LI1_cond $X=13.215 $Y=1.665
+ $X2=13.215 $Y2=1.815
r28 9 10 16.4002 $w=2.58e-07 $l=3.7e-07 $layer=LI1_cond $X=13.215 $Y=1.295
+ $X2=13.215 $Y2=1.665
r29 8 9 16.4002 $w=2.58e-07 $l=3.7e-07 $layer=LI1_cond $X=13.215 $Y=0.925
+ $X2=13.215 $Y2=1.295
r30 7 8 16.4002 $w=2.58e-07 $l=3.7e-07 $layer=LI1_cond $X=13.215 $Y=0.555
+ $X2=13.215 $Y2=0.925
r31 7 24 4.21085 $w=2.58e-07 $l=9.5e-08 $layer=LI1_cond $X=13.215 $Y=0.555
+ $X2=13.215 $Y2=0.46
r32 2 44 400 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_PDIFF $count=1 $X=12.885
+ $Y=1.835 $X2=13.045 $Y2=1.98
r33 2 41 400 $w=1.7e-07 $l=1.15223e-06 $layer=licon1_PDIFF $count=1 $X=12.885
+ $Y=1.835 $X2=13.045 $Y2=2.91
r34 1 24 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=13.04
+ $Y=0.315 $X2=13.18 $Y2=0.46
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRTN_1%VGND 1 2 3 4 5 6 19 21 25 29 33 37 41 45 47
+ 55 60 68 73 83 84 90 93 96 99 102
c131 47 0 2.01056e-19 $X=3.875 $Y=0
r132 102 103 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.72 $Y=0
+ $X2=12.72 $Y2=0
r133 99 100 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.8 $Y=0 $X2=10.8
+ $Y2=0
r134 96 97 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r135 93 94 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r136 90 91 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r137 87 88 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r138 84 103 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.2 $Y=0
+ $X2=12.72 $Y2=0
r139 83 84 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.2 $Y=0 $X2=13.2
+ $Y2=0
r140 81 102 9.6488 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=12.915 $Y=0
+ $X2=12.72 $Y2=0
r141 81 83 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=12.915 $Y=0
+ $X2=13.2 $Y2=0
r142 80 103 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.24 $Y=0
+ $X2=12.72 $Y2=0
r143 79 80 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=12.24 $Y=0
+ $X2=12.24 $Y2=0
r144 77 80 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=11.28 $Y=0
+ $X2=12.24 $Y2=0
r145 77 100 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=0
+ $X2=10.8 $Y2=0
r146 76 79 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=11.28 $Y=0 $X2=12.24
+ $Y2=0
r147 76 77 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=11.28 $Y=0
+ $X2=11.28 $Y2=0
r148 74 99 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.89 $Y=0
+ $X2=10.725 $Y2=0
r149 74 76 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=10.89 $Y=0
+ $X2=11.28 $Y2=0
r150 73 102 9.6488 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=12.525 $Y=0
+ $X2=12.72 $Y2=0
r151 73 79 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=12.525 $Y=0
+ $X2=12.24 $Y2=0
r152 72 100 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=0
+ $X2=10.8 $Y2=0
r153 72 97 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=10.32 $Y=0
+ $X2=8.4 $Y2=0
r154 71 72 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=10.32 $Y=0
+ $X2=10.32 $Y2=0
r155 69 96 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.45 $Y=0 $X2=8.285
+ $Y2=0
r156 69 71 122 $w=1.68e-07 $l=1.87e-06 $layer=LI1_cond $X=8.45 $Y=0 $X2=10.32
+ $Y2=0
r157 68 99 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.56 $Y=0
+ $X2=10.725 $Y2=0
r158 68 71 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=10.56 $Y=0
+ $X2=10.32 $Y2=0
r159 67 97 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0 $X2=8.4
+ $Y2=0
r160 66 67 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r161 64 94 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=5.04
+ $Y2=0
r162 63 66 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=5.52 $Y=0 $X2=7.92
+ $Y2=0
r163 63 64 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r164 61 93 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.275 $Y=0 $X2=5.11
+ $Y2=0
r165 61 63 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=5.275 $Y=0 $X2=5.52
+ $Y2=0
r166 60 96 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.12 $Y=0 $X2=8.285
+ $Y2=0
r167 60 66 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=8.12 $Y=0 $X2=7.92
+ $Y2=0
r168 59 94 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.04
+ $Y2=0
r169 59 91 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=4.08
+ $Y2=0
r170 58 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r171 56 90 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.205 $Y=0 $X2=4.04
+ $Y2=0
r172 56 58 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=4.205 $Y=0
+ $X2=4.56 $Y2=0
r173 55 93 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.945 $Y=0 $X2=5.11
+ $Y2=0
r174 55 58 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=4.945 $Y=0
+ $X2=4.56 $Y2=0
r175 54 91 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r176 53 54 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=3.6 $Y=0
+ $X2=3.6 $Y2=0
r177 51 54 0.802756 $w=4.9e-07 $l=2.88e-06 $layer=MET1_cond $X=0.72 $Y=0 $X2=3.6
+ $Y2=0
r178 51 88 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r179 50 53 187.893 $w=1.68e-07 $l=2.88e-06 $layer=LI1_cond $X=0.72 $Y=0 $X2=3.6
+ $Y2=0
r180 50 51 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=0.72 $Y=0
+ $X2=0.72 $Y2=0
r181 48 87 4.42547 $w=1.7e-07 $l=2.03e-07 $layer=LI1_cond $X=0.405 $Y=0
+ $X2=0.202 $Y2=0
r182 48 50 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.405 $Y=0
+ $X2=0.72 $Y2=0
r183 47 90 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.875 $Y=0 $X2=4.04
+ $Y2=0
r184 47 53 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=3.875 $Y=0 $X2=3.6
+ $Y2=0
r185 45 67 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=6.72 $Y=0 $X2=7.92
+ $Y2=0
r186 45 64 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=6.72 $Y=0 $X2=5.52
+ $Y2=0
r187 41 43 15.6614 $w=3.88e-07 $l=5.3e-07 $layer=LI1_cond $X=12.72 $Y=0.46
+ $X2=12.72 $Y2=0.99
r188 39 102 1.39532 $w=3.9e-07 $l=8.5e-08 $layer=LI1_cond $X=12.72 $Y=0.085
+ $X2=12.72 $Y2=0
r189 39 41 11.0812 $w=3.88e-07 $l=3.75e-07 $layer=LI1_cond $X=12.72 $Y=0.085
+ $X2=12.72 $Y2=0.46
r190 35 99 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.725 $Y=0.085
+ $X2=10.725 $Y2=0
r191 35 37 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=10.725 $Y=0.085
+ $X2=10.725 $Y2=0.76
r192 31 96 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.285 $Y=0.085
+ $X2=8.285 $Y2=0
r193 31 33 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=8.285 $Y=0.085
+ $X2=8.285 $Y2=0.455
r194 27 93 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.11 $Y=0.085
+ $X2=5.11 $Y2=0
r195 27 29 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=5.11 $Y=0.085
+ $X2=5.11 $Y2=0.36
r196 23 90 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.04 $Y=0.085
+ $X2=4.04 $Y2=0
r197 23 25 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=4.04 $Y=0.085
+ $X2=4.04 $Y2=0.36
r198 19 87 3.05205 $w=2.95e-07 $l=1.09087e-07 $layer=LI1_cond $X=0.257 $Y=0.085
+ $X2=0.202 $Y2=0
r199 19 21 17.189 $w=2.93e-07 $l=4.4e-07 $layer=LI1_cond $X=0.257 $Y=0.085
+ $X2=0.257 $Y2=0.525
r200 6 43 182 $w=1.7e-07 $l=7.83741e-07 $layer=licon1_NDIFF $count=1 $X=12.515
+ $Y=0.315 $X2=12.75 $Y2=0.99
r201 6 41 182 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_NDIFF $count=1 $X=12.515
+ $Y=0.315 $X2=12.69 $Y2=0.46
r202 5 37 182 $w=1.7e-07 $l=3.11288e-07 $layer=licon1_NDIFF $count=1 $X=10.47
+ $Y=0.635 $X2=10.725 $Y2=0.76
r203 4 33 182 $w=1.7e-07 $l=4.61302e-07 $layer=licon1_NDIFF $count=1 $X=7.905
+ $Y=0.635 $X2=8.285 $Y2=0.455
r204 3 29 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=4.965
+ $Y=0.235 $X2=5.11 $Y2=0.36
r205 2 25 182 $w=1.7e-07 $l=2.85657e-07 $layer=licon1_NDIFF $count=1 $X=3.785
+ $Y=0.295 $X2=4.04 $Y2=0.36
r206 1 21 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.15
+ $Y=0.315 $X2=0.275 $Y2=0.525
.ends

.subckt PM_SKY130_FD_SC_LP__SDFRTN_1%noxref_24 1 2 9 15 16
c31 9 0 9.05516e-21 $X=1.515 $Y=0.35
r32 15 16 8.79328 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=3.385 $Y=0.39
+ $X2=3.22 $Y2=0.39
r33 9 12 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=1.515 $Y=0.35 $X2=1.515
+ $Y2=0.44
r34 8 9 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.68 $Y=0.35 $X2=1.515
+ $Y2=0.35
r35 8 16 100.471 $w=1.68e-07 $l=1.54e-06 $layer=LI1_cond $X=1.68 $Y=0.35
+ $X2=3.22 $Y2=0.35
r36 2 15 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=3.245
+ $Y=0.295 $X2=3.385 $Y2=0.42
r37 1 12 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=1.39
+ $Y=0.295 $X2=1.515 $Y2=0.44
.ends

