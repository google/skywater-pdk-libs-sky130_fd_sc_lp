* File: sky130_fd_sc_lp__and3b_2.pex.spice
* Created: Fri Aug 28 10:06:44 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__AND3B_2%A_N 3 6 8 9 13 15
c27 15 0 3.02108e-20 $X=0.577 $Y=1.215
r28 13 16 46.504 $w=3.55e-07 $l=1.65e-07 $layer=POLY_cond $X=0.577 $Y=1.38
+ $X2=0.577 $Y2=1.545
r29 13 15 46.504 $w=3.55e-07 $l=1.65e-07 $layer=POLY_cond $X=0.577 $Y=1.38
+ $X2=0.577 $Y2=1.215
r30 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.59
+ $Y=1.38 $X2=0.59 $Y2=1.38
r31 9 14 7.91437 $w=4.13e-07 $l=2.85e-07 $layer=LI1_cond $X=0.712 $Y=1.665
+ $X2=0.712 $Y2=1.38
r32 8 14 2.36043 $w=4.13e-07 $l=8.5e-08 $layer=LI1_cond $X=0.712 $Y=1.295
+ $X2=0.712 $Y2=1.38
r33 6 16 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=0.535 $Y=2.045
+ $X2=0.535 $Y2=1.545
r34 3 15 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.475 $Y=0.895
+ $X2=0.475 $Y2=1.215
.ends

.subckt PM_SKY130_FD_SC_LP__AND3B_2%A_204_27# 1 2 3 12 16 22 26 28 31 32 34 35
+ 36 40 44 47 50 52
c86 36 0 1.5437e-19 $X=3.4 $Y=1.74
r87 51 52 30.474 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=1.525 $Y=1.46
+ $X2=1.45 $Y2=1.46
r88 47 49 8.92177 $w=2.94e-07 $l=2.15e-07 $layer=LI1_cond $X=2.56 $Y=1.82
+ $X2=2.56 $Y2=2.035
r89 46 47 3.31973 $w=2.94e-07 $l=8e-08 $layer=LI1_cond $X=2.56 $Y=1.74 $X2=2.56
+ $Y2=1.82
r90 42 50 3.52026 $w=2.65e-07 $l=8.74643e-08 $layer=LI1_cond $X=3.54 $Y=1.825
+ $X2=3.535 $Y2=1.74
r91 42 44 9.30819 $w=2.58e-07 $l=2.1e-07 $layer=LI1_cond $X=3.54 $Y=1.825
+ $X2=3.54 $Y2=2.035
r92 38 50 3.52026 $w=2.65e-07 $l=8.5e-08 $layer=LI1_cond $X=3.535 $Y=1.655
+ $X2=3.535 $Y2=1.74
r93 38 40 32.4391 $w=2.68e-07 $l=7.6e-07 $layer=LI1_cond $X=3.535 $Y=1.655
+ $X2=3.535 $Y2=0.895
r94 37 46 3.94234 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=2.715 $Y=1.74
+ $X2=2.56 $Y2=1.74
r95 36 50 2.98021 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=3.4 $Y=1.74
+ $X2=3.535 $Y2=1.74
r96 36 37 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=3.4 $Y=1.74
+ $X2=2.715 $Y2=1.74
r97 34 47 2.70854 $w=2.1e-07 $l=1.55e-07 $layer=LI1_cond $X=2.405 $Y=1.82
+ $X2=2.56 $Y2=1.82
r98 34 35 29.0476 $w=2.08e-07 $l=5.5e-07 $layer=LI1_cond $X=2.405 $Y=1.82
+ $X2=1.855 $Y2=1.82
r99 32 51 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=1.74 $Y=1.46
+ $X2=1.525 $Y2=1.46
r100 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.74
+ $Y=1.46 $X2=1.74 $Y2=1.46
r101 29 35 6.81649 $w=2.1e-07 $l=1.48492e-07 $layer=LI1_cond $X=1.75 $Y=1.715
+ $X2=1.855 $Y2=1.82
r102 29 31 13.4675 $w=2.08e-07 $l=2.55e-07 $layer=LI1_cond $X=1.75 $Y=1.715
+ $X2=1.75 $Y2=1.46
r103 24 51 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.525 $Y=1.625
+ $X2=1.525 $Y2=1.46
r104 24 26 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=1.525 $Y=1.625
+ $X2=1.525 $Y2=2.465
r105 20 51 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.525 $Y=1.295
+ $X2=1.525 $Y2=1.46
r106 20 22 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.525 $Y=1.295
+ $X2=1.525 $Y2=0.685
r107 19 28 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.17 $Y=1.55
+ $X2=1.095 $Y2=1.55
r108 19 52 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=1.17 $Y=1.55
+ $X2=1.45 $Y2=1.55
r109 14 28 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.095 $Y=1.625
+ $X2=1.095 $Y2=1.55
r110 14 16 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=1.095 $Y=1.625
+ $X2=1.095 $Y2=2.465
r111 10 28 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.095 $Y=1.475
+ $X2=1.095 $Y2=1.55
r112 10 12 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.095 $Y=1.475
+ $X2=1.095 $Y2=0.685
r113 3 44 600 $w=1.7e-07 $l=2.60768e-07 $layer=licon1_PDIFF $count=1 $X=3.375
+ $Y=1.835 $X2=3.515 $Y2=2.035
r114 2 49 600 $w=1.7e-07 $l=2.60768e-07 $layer=licon1_PDIFF $count=1 $X=2.43
+ $Y=1.835 $X2=2.57 $Y2=2.035
r115 1 40 182 $w=1.7e-07 $l=2.78747e-07 $layer=licon1_NDIFF $count=1 $X=3.345
+ $Y=0.685 $X2=3.505 $Y2=0.895
.ends

.subckt PM_SKY130_FD_SC_LP__AND3B_2%C 3 7 8 11 12 13
c33 11 0 1.11559e-19 $X=2.28 $Y=1.38
r34 11 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.28 $Y=1.38
+ $X2=2.28 $Y2=1.545
r35 11 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.28 $Y=1.38
+ $X2=2.28 $Y2=1.215
r36 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.28
+ $Y=1.38 $X2=2.28 $Y2=1.38
r37 8 12 3.33237 $w=4.13e-07 $l=1.2e-07 $layer=LI1_cond $X=2.16 $Y=1.337
+ $X2=2.28 $Y2=1.337
r38 7 13 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.37 $Y=0.895
+ $X2=2.37 $Y2=1.215
r39 3 14 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=2.355 $Y=2.045
+ $X2=2.355 $Y2=1.545
.ends

.subckt PM_SKY130_FD_SC_LP__AND3B_2%B 3 6 8 9 13 15
r34 13 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.82 $Y=1.38
+ $X2=2.82 $Y2=1.545
r35 13 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.82 $Y=1.38
+ $X2=2.82 $Y2=1.215
r36 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.82
+ $Y=1.38 $X2=2.82 $Y2=1.38
r37 9 14 9.73895 $w=3.53e-07 $l=3e-07 $layer=LI1_cond $X=3.12 $Y=1.307 $X2=2.82
+ $Y2=1.307
r38 8 14 5.84337 $w=3.53e-07 $l=1.8e-07 $layer=LI1_cond $X=2.64 $Y=1.307
+ $X2=2.82 $Y2=1.307
r39 6 16 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=2.785 $Y=2.045
+ $X2=2.785 $Y2=1.545
r40 3 15 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.73 $Y=0.895
+ $X2=2.73 $Y2=1.215
.ends

.subckt PM_SKY130_FD_SC_LP__AND3B_2%A_27_137# 1 2 10 13 16 18 21 22 23 31 33 35
+ 36
c71 16 0 1.5437e-19 $X=3.285 $Y=1.365
r72 36 40 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.21 $Y=0.41
+ $X2=3.21 $Y2=0.575
r73 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.21
+ $Y=0.41 $X2=3.21 $Y2=0.41
r74 28 31 4.69514 $w=2.68e-07 $l=1.1e-07 $layer=LI1_cond $X=0.21 $Y=2.065
+ $X2=0.32 $Y2=2.065
r75 26 27 6.13416 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=0.26 $Y=0.895
+ $X2=0.26 $Y2=1.04
r76 23 26 9.25447 $w=3.28e-07 $l=2.65e-07 $layer=LI1_cond $X=0.26 $Y=0.63
+ $X2=0.26 $Y2=0.895
r77 22 33 8.35379 $w=3.23e-07 $l=1.62e-07 $layer=LI1_cond $X=1.807 $Y=0.707
+ $X2=1.645 $Y2=0.707
r78 21 35 14.1539 $w=2.56e-07 $l=2.97e-07 $layer=LI1_cond $X=3.21 $Y=0.707
+ $X2=3.21 $Y2=0.41
r79 21 22 43.8992 $w=3.23e-07 $l=1.238e-06 $layer=LI1_cond $X=3.045 $Y=0.707
+ $X2=1.807 $Y2=0.707
r80 20 23 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.425 $Y=0.63
+ $X2=0.26 $Y2=0.63
r81 20 33 79.5936 $w=1.68e-07 $l=1.22e-06 $layer=LI1_cond $X=0.425 $Y=0.63
+ $X2=1.645 $Y2=0.63
r82 18 28 1.67709 $w=2.3e-07 $l=1.35e-07 $layer=LI1_cond $X=0.21 $Y=1.93
+ $X2=0.21 $Y2=2.065
r83 18 27 44.5945 $w=2.28e-07 $l=8.9e-07 $layer=LI1_cond $X=0.21 $Y=1.93
+ $X2=0.21 $Y2=1.04
r84 15 16 58.3064 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=3.285 $Y=1.215
+ $X2=3.285 $Y2=1.365
r85 13 16 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=3.3 $Y=2.045 $X2=3.3
+ $Y2=1.365
r86 10 15 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=3.27 $Y=0.895
+ $X2=3.27 $Y2=1.215
r87 10 40 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=3.27 $Y=0.895
+ $X2=3.27 $Y2=0.575
r88 2 31 600 $w=1.7e-07 $l=2.54951e-07 $layer=licon1_PDIFF $count=1 $X=0.195
+ $Y=1.835 $X2=0.32 $Y2=2.035
r89 1 26 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.685 $X2=0.26 $Y2=0.895
.ends

.subckt PM_SKY130_FD_SC_LP__AND3B_2%VPWR 1 2 3 14 18 22 28 30 32 39 40 43 46 49
r34 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r35 46 47 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r36 44 47 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r37 43 44 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r38 40 50 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=3.12 $Y2=3.33
r39 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r40 37 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.225 $Y=3.33
+ $X2=3.06 $Y2=3.33
r41 37 39 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=3.225 $Y=3.33
+ $X2=3.6 $Y2=3.33
r42 36 50 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r43 35 36 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r44 33 46 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=1.925 $Y=3.33
+ $X2=1.785 $Y2=3.33
r45 33 35 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=1.925 $Y=3.33
+ $X2=2.64 $Y2=3.33
r46 32 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.895 $Y=3.33
+ $X2=3.06 $Y2=3.33
r47 32 35 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=2.895 $Y=3.33
+ $X2=2.64 $Y2=3.33
r48 30 36 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=2.64 $Y2=3.33
r49 30 47 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=1.68 $Y2=3.33
r50 26 49 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.06 $Y=3.245
+ $X2=3.06 $Y2=3.33
r51 26 28 39.6371 $w=3.28e-07 $l=1.135e-06 $layer=LI1_cond $X=3.06 $Y=3.245
+ $X2=3.06 $Y2=2.11
r52 22 25 28.3995 $w=2.78e-07 $l=6.9e-07 $layer=LI1_cond $X=1.785 $Y=2.26
+ $X2=1.785 $Y2=2.95
r53 20 46 0.375625 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=1.785 $Y=3.245
+ $X2=1.785 $Y2=3.33
r54 20 25 12.1418 $w=2.78e-07 $l=2.95e-07 $layer=LI1_cond $X=1.785 $Y=3.245
+ $X2=1.785 $Y2=2.95
r55 19 43 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=0.945 $Y=3.33
+ $X2=0.8 $Y2=3.33
r56 18 46 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=1.645 $Y=3.33
+ $X2=1.785 $Y2=3.33
r57 18 19 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=1.645 $Y=3.33
+ $X2=0.945 $Y2=3.33
r58 14 17 16.4919 $w=2.88e-07 $l=4.15e-07 $layer=LI1_cond $X=0.8 $Y=2.095
+ $X2=0.8 $Y2=2.51
r59 12 43 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=0.8 $Y=3.245 $X2=0.8
+ $Y2=3.33
r60 12 17 29.2085 $w=2.88e-07 $l=7.35e-07 $layer=LI1_cond $X=0.8 $Y=3.245
+ $X2=0.8 $Y2=2.51
r61 3 28 600 $w=1.7e-07 $l=3.61421e-07 $layer=licon1_PDIFF $count=1 $X=2.86
+ $Y=1.835 $X2=3.06 $Y2=2.11
r62 2 25 400 $w=1.7e-07 $l=1.19232e-06 $layer=licon1_PDIFF $count=1 $X=1.6
+ $Y=1.835 $X2=1.76 $Y2=2.95
r63 2 22 400 $w=1.7e-07 $l=4.98623e-07 $layer=licon1_PDIFF $count=1 $X=1.6
+ $Y=1.835 $X2=1.76 $Y2=2.26
r64 1 17 300 $w=1.7e-07 $l=7.85891e-07 $layer=licon1_PDIFF $count=2 $X=0.61
+ $Y=1.835 $X2=0.85 $Y2=2.51
r65 1 14 600 $w=1.7e-07 $l=3.2249e-07 $layer=licon1_PDIFF $count=1 $X=0.61
+ $Y=1.835 $X2=0.75 $Y2=2.095
.ends

.subckt PM_SKY130_FD_SC_LP__AND3B_2%X 1 2 7 8 9 10 11 18
c20 18 0 1.11559e-19 $X=1.31 $Y=0.98
r21 11 33 4.32166 $w=3.58e-07 $l=1.35e-07 $layer=LI1_cond $X=1.295 $Y=2.775
+ $X2=1.295 $Y2=2.91
r22 10 11 11.8446 $w=3.58e-07 $l=3.7e-07 $layer=LI1_cond $X=1.295 $Y=2.405
+ $X2=1.295 $Y2=2.775
r23 9 10 11.8446 $w=3.58e-07 $l=3.7e-07 $layer=LI1_cond $X=1.295 $Y=2.035
+ $X2=1.295 $Y2=2.405
r24 9 25 1.76068 $w=3.58e-07 $l=5.5e-08 $layer=LI1_cond $X=1.295 $Y=2.035
+ $X2=1.295 $Y2=1.98
r25 8 25 10.0839 $w=3.58e-07 $l=3.15e-07 $layer=LI1_cond $X=1.295 $Y=1.665
+ $X2=1.295 $Y2=1.98
r26 7 8 11.8446 $w=3.58e-07 $l=3.7e-07 $layer=LI1_cond $X=1.295 $Y=1.295
+ $X2=1.295 $Y2=1.665
r27 7 18 10.0839 $w=3.58e-07 $l=3.15e-07 $layer=LI1_cond $X=1.295 $Y=1.295
+ $X2=1.295 $Y2=0.98
r28 2 33 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=1.17
+ $Y=1.835 $X2=1.31 $Y2=2.91
r29 2 25 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.17
+ $Y=1.835 $X2=1.31 $Y2=1.98
r30 1 18 182 $w=1.7e-07 $l=7.81873e-07 $layer=licon1_NDIFF $count=1 $X=1.17
+ $Y=0.265 $X2=1.31 $Y2=0.98
.ends

.subckt PM_SKY130_FD_SC_LP__AND3B_2%VGND 1 2 7 8 14 16 29 30 34
c34 30 0 3.02108e-20 $X=3.6 $Y=0
r35 34 37 9.7783 $w=3.28e-07 $l=2.8e-07 $layer=LI1_cond $X=0.785 $Y=0 $X2=0.785
+ $Y2=0.28
r36 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r37 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r38 27 30 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.6
+ $Y2=0
r39 26 29 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=2.16 $Y=0 $X2=3.6
+ $Y2=0
r40 26 27 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r41 24 35 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=0.72
+ $Y2=0
r42 23 24 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r43 21 34 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.95 $Y=0 $X2=0.785
+ $Y2=0
r44 21 23 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=0.95 $Y=0 $X2=1.68
+ $Y2=0
r45 19 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r46 18 19 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r47 16 34 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.62 $Y=0 $X2=0.785
+ $Y2=0
r48 16 18 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=0.62 $Y=0 $X2=0.24
+ $Y2=0
r49 14 27 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=2.16
+ $Y2=0
r50 14 24 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=1.68
+ $Y2=0
r51 10 26 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=2.02 $Y=0 $X2=2.16
+ $Y2=0
r52 8 23 0.652406 $w=1.68e-07 $l=1e-08 $layer=LI1_cond $X=1.69 $Y=0 $X2=1.68
+ $Y2=0
r53 7 12 9.7783 $w=3.28e-07 $l=2.8e-07 $layer=LI1_cond $X=1.855 $Y=0 $X2=1.855
+ $Y2=0.28
r54 7 10 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.855 $Y=0 $X2=2.02
+ $Y2=0
r55 7 8 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.855 $Y=0 $X2=1.69
+ $Y2=0
r56 2 12 182 $w=1.7e-07 $l=2.62393e-07 $layer=licon1_NDIFF $count=1 $X=1.6
+ $Y=0.265 $X2=1.855 $Y2=0.28
r57 1 37 182 $w=1.7e-07 $l=5.09117e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.685 $X2=0.785 $Y2=0.28
.ends

