* File: sky130_fd_sc_lp__einvn_2.spice
* Created: Wed Sep  2 09:51:39 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__einvn_2.pex.spice"
.subckt sky130_fd_sc_lp__einvn_2  VNB VPB TE_B A VPWR Z VGND
* 
* VGND	VGND
* Z	Z
* VPWR	VPWR
* A	A
* TE_B	TE_B
* VPB	VPB
* VNB	VNB
MM1002 N_VGND_M1002_d N_TE_B_M1002_g N_A_28_62#_M1002_s VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.1197 PD=1.37 PS=1.41 NRD=0 NRS=5.712 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1004 N_VGND_M1004_d N_A_28_62#_M1004_g N_A_251_47#_M1004_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75001.5 A=0.126 P=1.98 MULT=1
MM1005 N_VGND_M1004_d N_A_28_62#_M1005_g N_A_251_47#_M1005_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1001 N_Z_M1001_d N_A_M1001_g N_A_251_47#_M1005_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.1
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1003 N_Z_M1001_d N_A_M1003_g N_A_251_47#_M1003_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75001.5
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1006 N_VPWR_M1006_d N_TE_B_M1006_g N_A_28_62#_M1006_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.136185 AS=0.1696 PD=1.10147 PS=1.81 NRD=63.0991 NRS=0 M=1
+ R=4.26667 SA=75000.2 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1007 N_VPWR_M1006_d N_TE_B_M1007_g N_A_220_367#_M1007_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.268115 AS=0.1764 PD=2.16853 PS=1.54 NRD=2.3443 NRS=0 M=1 R=8.4
+ SA=75000.5 SB=75000.6 A=0.189 P=2.82 MULT=1
MM1009 N_VPWR_M1009_d N_TE_B_M1009_g N_A_220_367#_M1007_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.9
+ SB=75000.2 A=0.189 P=2.82 MULT=1
MM1000 N_A_220_367#_M1000_d N_A_M1000_g N_Z_M1000_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1008 N_A_220_367#_M1000_d N_A_M1008_g N_Z_M1008_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9751 P=11.21
*
.include "sky130_fd_sc_lp__einvn_2.pxi.spice"
*
.ends
*
*
