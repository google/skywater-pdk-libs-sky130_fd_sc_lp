# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__dlclkp_1
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__dlclkp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.720000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN GATE
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.975000 1.160000 1.415000 1.390000 ;
    END
  END GATE
  PIN GCLK
    ANTENNADIFFAREA  0.556500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.365000 0.255000 6.625000 3.075000 ;
    END
  END GCLK
  PIN CLK
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 3.465000 1.420000 3.915000 1.765000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 6.720000 0.085000 ;
        RECT 0.745000  0.085000 1.075000 0.650000 ;
        RECT 2.790000  0.085000 3.040000 0.780000 ;
        RECT 4.440000  0.085000 4.770000 0.515000 ;
        RECT 5.865000  0.085000 6.195000 0.495000 ;
      LAYER mcon ;
        RECT 0.155000 -0.085000 0.325000 0.085000 ;
        RECT 0.635000 -0.085000 0.805000 0.085000 ;
        RECT 1.115000 -0.085000 1.285000 0.085000 ;
        RECT 1.595000 -0.085000 1.765000 0.085000 ;
        RECT 2.075000 -0.085000 2.245000 0.085000 ;
        RECT 2.555000 -0.085000 2.725000 0.085000 ;
        RECT 3.035000 -0.085000 3.205000 0.085000 ;
        RECT 3.515000 -0.085000 3.685000 0.085000 ;
        RECT 3.995000 -0.085000 4.165000 0.085000 ;
        RECT 4.475000 -0.085000 4.645000 0.085000 ;
        RECT 4.955000 -0.085000 5.125000 0.085000 ;
        RECT 5.435000 -0.085000 5.605000 0.085000 ;
        RECT 5.915000 -0.085000 6.085000 0.085000 ;
        RECT 6.395000 -0.085000 6.565000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 6.720000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 3.245000 6.720000 3.415000 ;
        RECT 0.605000 2.240000 0.805000 3.245000 ;
        RECT 2.715000 2.615000 3.045000 3.245000 ;
        RECT 4.695000 2.905000 5.025000 3.245000 ;
        RECT 5.635000 1.835000 6.195000 3.245000 ;
      LAYER mcon ;
        RECT 0.155000 3.245000 0.325000 3.415000 ;
        RECT 0.635000 3.245000 0.805000 3.415000 ;
        RECT 1.115000 3.245000 1.285000 3.415000 ;
        RECT 1.595000 3.245000 1.765000 3.415000 ;
        RECT 2.075000 3.245000 2.245000 3.415000 ;
        RECT 2.555000 3.245000 2.725000 3.415000 ;
        RECT 3.035000 3.245000 3.205000 3.415000 ;
        RECT 3.515000 3.245000 3.685000 3.415000 ;
        RECT 3.995000 3.245000 4.165000 3.415000 ;
        RECT 4.475000 3.245000 4.645000 3.415000 ;
        RECT 4.955000 3.245000 5.125000 3.415000 ;
        RECT 5.435000 3.245000 5.605000 3.415000 ;
        RECT 5.915000 3.245000 6.085000 3.415000 ;
        RECT 6.395000 3.245000 6.565000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 6.720000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.095000 0.255000 0.575000 0.820000 ;
      RECT 0.095000 0.820000 1.415000 0.990000 ;
      RECT 0.095000 0.990000 0.580000 1.095000 ;
      RECT 0.095000 1.095000 0.365000 1.900000 ;
      RECT 0.095000 1.900000 1.145000 2.070000 ;
      RECT 0.095000 2.070000 0.425000 3.075000 ;
      RECT 0.535000 1.345000 0.795000 1.560000 ;
      RECT 0.535000 1.560000 1.755000 1.730000 ;
      RECT 0.975000 2.070000 1.145000 2.905000 ;
      RECT 0.975000 2.905000 2.445000 3.075000 ;
      RECT 1.245000 0.255000 2.620000 0.425000 ;
      RECT 1.245000 0.425000 1.415000 0.820000 ;
      RECT 1.315000 1.730000 1.755000 1.740000 ;
      RECT 1.315000 1.740000 1.485000 2.485000 ;
      RECT 1.315000 2.485000 2.070000 2.735000 ;
      RECT 1.585000 0.595000 2.060000 0.795000 ;
      RECT 1.585000 0.795000 1.755000 1.560000 ;
      RECT 1.655000 1.910000 2.095000 1.935000 ;
      RECT 1.655000 1.935000 3.825000 2.105000 ;
      RECT 1.655000 2.105000 2.095000 2.240000 ;
      RECT 1.925000 0.965000 2.280000 1.295000 ;
      RECT 1.925000 1.295000 2.095000 1.910000 ;
      RECT 2.265000 1.505000 3.295000 1.765000 ;
      RECT 2.275000 2.275000 3.395000 2.445000 ;
      RECT 2.275000 2.445000 2.445000 2.905000 ;
      RECT 2.450000 0.425000 2.620000 0.950000 ;
      RECT 2.450000 0.950000 2.835000 1.265000 ;
      RECT 3.045000 1.025000 4.415000 1.250000 ;
      RECT 3.045000 1.250000 3.295000 1.505000 ;
      RECT 3.210000 0.445000 3.500000 0.685000 ;
      RECT 3.210000 0.685000 4.755000 0.855000 ;
      RECT 3.225000 2.445000 3.395000 2.565000 ;
      RECT 3.225000 2.565000 5.095000 2.735000 ;
      RECT 3.225000 2.735000 3.915000 2.745000 ;
      RECT 3.565000 2.105000 3.825000 2.225000 ;
      RECT 3.565000 2.225000 4.755000 2.395000 ;
      RECT 3.585000 2.745000 3.915000 3.075000 ;
      RECT 4.085000 1.250000 4.415000 2.055000 ;
      RECT 4.585000 0.855000 4.755000 2.225000 ;
      RECT 4.925000 1.005000 5.675000 1.325000 ;
      RECT 4.925000 1.325000 5.095000 2.565000 ;
      RECT 5.265000 1.495000 6.195000 1.665000 ;
      RECT 5.265000 1.665000 5.465000 2.495000 ;
      RECT 5.345000 0.440000 5.675000 0.665000 ;
      RECT 5.345000 0.665000 6.195000 0.835000 ;
      RECT 5.945000 0.835000 6.195000 1.495000 ;
  END
END sky130_fd_sc_lp__dlclkp_1
