* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__dlclkp_4 CLK GATE VGND VNB VPB VPWR GCLK
X0 a_411_81# a_27_367# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 a_295_55# CLK VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 VGND GATE a_253_81# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 a_253_81# a_295_55# a_73_269# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 VPWR GATE a_235_465# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X5 a_73_269# a_277_367# a_411_81# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 a_27_367# a_73_269# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X7 GCLK a_1078_367# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X8 VGND a_1078_367# GCLK VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X9 VPWR a_1078_367# GCLK VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X10 GCLK a_1078_367# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X11 VGND a_1078_367# GCLK VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X12 VPWR CLK a_1078_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X13 VGND CLK a_1026_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X14 GCLK a_1078_367# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X15 a_73_269# a_295_55# a_415_465# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X16 a_415_465# a_27_367# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X17 VPWR a_295_55# a_277_367# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X18 a_27_367# a_73_269# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X19 GCLK a_1078_367# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X20 a_1078_367# a_27_367# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X21 VGND a_295_55# a_277_367# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X22 a_235_465# a_277_367# a_73_269# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X23 a_295_55# CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X24 a_1026_47# a_27_367# a_1078_367# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X25 VPWR a_1078_367# GCLK VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
.ends
