* NGSPICE file created from sky130_fd_sc_lp__a32oi_m.ext - technology: sky130A

.subckt sky130_fd_sc_lp__a32oi_m A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
M1000 Y B2 a_40_500# VPB phighvt w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=4.137e+11p ps=4.49e+06u
M1001 a_319_47# A1 Y VNB nshort w=420000u l=150000u
+  ad=1.638e+11p pd=1.62e+06u as=1.365e+11p ps=1.49e+06u
M1002 a_40_500# B1 Y VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 VPWR A1 a_40_500# VPB phighvt w=420000u l=150000u
+  ad=2.625e+11p pd=2.93e+06u as=0p ps=0u
M1004 a_40_500# A2 VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_427_47# A2 a_319_47# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1006 VGND A3 a_427_47# VNB nshort w=420000u l=150000u
+  ad=2.982e+11p pd=3.1e+06u as=0p ps=0u
M1007 Y B1 a_152_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1008 VPWR A3 a_40_500# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_152_47# B2 VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

