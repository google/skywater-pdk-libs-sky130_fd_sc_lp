* File: sky130_fd_sc_lp__srsdfrtn_1.pex.spice
* Created: Wed Sep  2 10:39:07 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__SRSDFRTN_1%SCE 3 7 9 11 15 17 19 21 23 24 25 29
c57 7 0 1.2623e-20 $X=0.66 $Y=2.775
r58 24 25 14.1436 $w=3.28e-07 $l=4.05e-07 $layer=LI1_cond $X=0.75 $Y=1.26
+ $X2=0.75 $Y2=1.665
r59 24 29 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.75
+ $Y=1.26 $X2=0.75 $Y2=1.26
r60 22 29 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=0.75 $Y=1.615
+ $X2=0.75 $Y2=1.26
r61 22 23 13.5877 $w=2.4e-07 $l=7.5e-08 $layer=POLY_cond $X=0.75 $Y=1.615
+ $X2=0.75 $Y2=1.69
r62 20 29 16.6118 $w=3.3e-07 $l=9.5e-08 $layer=POLY_cond $X=0.75 $Y=1.165
+ $X2=0.75 $Y2=1.26
r63 20 21 13.5877 $w=2.4e-07 $l=1.19766e-07 $layer=POLY_cond $X=0.75 $Y=1.165
+ $X2=0.662 $Y2=1.09
r64 17 19 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.45 $Y=1.015
+ $X2=1.45 $Y2=0.695
r65 13 15 517.894 $w=1.5e-07 $l=1.01e-06 $layer=POLY_cond $X=1.16 $Y=1.765
+ $X2=1.16 $Y2=2.775
r66 12 23 12.1617 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.915 $Y=1.69
+ $X2=0.75 $Y2=1.69
r67 11 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.085 $Y=1.69
+ $X2=1.16 $Y2=1.765
r68 11 12 87.1702 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=1.085 $Y=1.69
+ $X2=0.915 $Y2=1.69
r69 10 21 12.1617 $w=1.5e-07 $l=2.53e-07 $layer=POLY_cond $X=0.915 $Y=1.09
+ $X2=0.662 $Y2=1.09
r70 9 17 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.375 $Y=1.09
+ $X2=1.45 $Y2=1.015
r71 9 10 235.872 $w=1.5e-07 $l=4.6e-07 $layer=POLY_cond $X=1.375 $Y=1.09
+ $X2=0.915 $Y2=1.09
r72 5 23 13.5877 $w=2.4e-07 $l=1.21861e-07 $layer=POLY_cond $X=0.66 $Y=1.765
+ $X2=0.75 $Y2=1.69
r73 5 7 517.894 $w=1.5e-07 $l=1.01e-06 $layer=POLY_cond $X=0.66 $Y=1.765
+ $X2=0.66 $Y2=2.775
r74 1 21 13.5877 $w=2.4e-07 $l=2.11197e-07 $layer=POLY_cond $X=0.485 $Y=1.015
+ $X2=0.662 $Y2=1.09
r75 1 3 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.485 $Y=1.015
+ $X2=0.485 $Y2=0.485
.ends

.subckt PM_SKY130_FD_SC_LP__SRSDFRTN_1%D 3 7 9 11 19
c45 11 0 1.06697e-19 $X=1.68 $Y=1.665
r46 19 21 36.7238 $w=3.15e-07 $l=2.4e-07 $layer=POLY_cond $X=1.64 $Y=1.54
+ $X2=1.88 $Y2=1.54
r47 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.64
+ $Y=1.54 $X2=1.64 $Y2=1.54
r48 17 19 13.7714 $w=3.15e-07 $l=9e-08 $layer=POLY_cond $X=1.55 $Y=1.54 $X2=1.64
+ $Y2=1.54
r49 11 20 0.797386 $w=5.98e-07 $l=4e-08 $layer=LI1_cond $X=1.68 $Y=1.48 $X2=1.64
+ $Y2=1.48
r50 9 20 8.77124 $w=5.98e-07 $l=4.4e-07 $layer=LI1_cond $X=1.2 $Y=1.48 $X2=1.64
+ $Y2=1.48
r51 5 21 20.1192 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.88 $Y=1.375
+ $X2=1.88 $Y2=1.54
r52 5 7 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=1.88 $Y=1.375 $X2=1.88
+ $Y2=0.695
r53 1 17 20.1192 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.55 $Y=1.705
+ $X2=1.55 $Y2=1.54
r54 1 3 548.66 $w=1.5e-07 $l=1.07e-06 $layer=POLY_cond $X=1.55 $Y=1.705 $X2=1.55
+ $Y2=2.775
.ends

.subckt PM_SKY130_FD_SC_LP__SRSDFRTN_1%A_27_55# 1 2 7 9 12 15 18 21 25 29 31 33
c79 31 0 1.46816e-19 $X=2.14 $Y=2.11
c80 18 0 9.4074e-20 $X=2.255 $Y=1.365
c81 15 0 1.55978e-19 $X=2.27 $Y=0.695
r82 31 33 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=2.14 $Y=2.11
+ $X2=1.975 $Y2=2.11
r83 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.14
+ $Y=2.11 $X2=2.14 $Y2=2.11
r84 28 29 4.32201 $w=1.7e-07 $l=2.53e-07 $layer=LI1_cond $X=0.61 $Y=2.035
+ $X2=0.357 $Y2=2.035
r85 28 33 89.0535 $w=1.68e-07 $l=1.365e-06 $layer=LI1_cond $X=0.61 $Y=2.035
+ $X2=1.975 $Y2=2.035
r86 23 29 2.55177 $w=3.77e-07 $l=8.5e-08 $layer=LI1_cond $X=0.357 $Y=2.12
+ $X2=0.357 $Y2=2.035
r87 23 25 15.0398 $w=5.03e-07 $l=6.35e-07 $layer=LI1_cond $X=0.357 $Y=2.12
+ $X2=0.357 $Y2=2.755
r88 19 29 2.55177 $w=3.77e-07 $l=1.64085e-07 $layer=LI1_cond $X=0.23 $Y=1.95
+ $X2=0.357 $Y2=2.035
r89 19 21 67.5332 $w=2.48e-07 $l=1.465e-06 $layer=LI1_cond $X=0.23 $Y=1.95
+ $X2=0.23 $Y2=0.485
r90 17 18 58.3064 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=2.255 $Y=1.215
+ $X2=2.255 $Y2=1.365
r91 15 17 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=2.27 $Y=0.695
+ $X2=2.27 $Y2=1.215
r92 12 32 66.1652 $w=3.14e-07 $l=4.04815e-07 $layer=POLY_cond $X=2.24 $Y=1.765
+ $X2=2.11 $Y2=2.11
r93 12 18 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=2.24 $Y=1.765 $X2=2.24
+ $Y2=1.365
r94 7 32 38.5347 $w=3.14e-07 $l=2.20624e-07 $layer=POLY_cond $X=1.98 $Y=2.275
+ $X2=2.11 $Y2=2.11
r95 7 9 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=1.98 $Y=2.275 $X2=1.98
+ $Y2=2.775
r96 2 25 600 $w=1.7e-07 $l=3.65377e-07 $layer=licon1_PDIFF $count=1 $X=0.3
+ $Y=2.455 $X2=0.445 $Y2=2.755
r97 1 21 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.275 $X2=0.27 $Y2=0.485
.ends

.subckt PM_SKY130_FD_SC_LP__SRSDFRTN_1%SCD 3 7 10 11 14 17 18
c41 11 0 1.46816e-19 $X=2.715 $Y=2.305
c42 7 0 3.39925e-20 $X=2.7 $Y=0.695
r43 17 18 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.72
+ $Y=1.77 $X2=2.72 $Y2=1.77
r44 14 18 8.8521 $w=3.43e-07 $l=2.65e-07 $layer=LI1_cond $X=2.697 $Y=2.035
+ $X2=2.697 $Y2=1.77
r45 13 17 38.6168 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.72 $Y=1.605
+ $X2=2.72 $Y2=1.77
r46 10 17 67.3216 $w=3.3e-07 $l=3.85e-07 $layer=POLY_cond $X=2.72 $Y=2.155
+ $X2=2.72 $Y2=1.77
r47 10 11 43.5886 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=2.715 $Y=2.155
+ $X2=2.715 $Y2=2.305
r48 7 13 466.617 $w=1.5e-07 $l=9.1e-07 $layer=POLY_cond $X=2.7 $Y=0.695 $X2=2.7
+ $Y2=1.605
r49 3 11 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=2.62 $Y=2.775 $X2=2.62
+ $Y2=2.305
.ends

.subckt PM_SKY130_FD_SC_LP__SRSDFRTN_1%RESET_B 1 3 6 9 13 16 18 19 22 24 25 29
+ 33 35 36 37 40 43 44 45 46 51 56
c182 45 0 1.86972e-19 $X=7.07 $Y=1.695
c183 43 0 3.9366e-21 $X=6.985 $Y=1.61
c184 37 0 2.87822e-20 $X=6.9 $Y=0.34
c185 36 0 2.70432e-19 $X=8.16 $Y=1.215
c186 33 0 1.81355e-19 $X=4.86 $Y=1.22
c187 6 0 1.41889e-19 $X=4.585 $Y=2.415
r188 50 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.975
+ $Y=1.38 $X2=7.975 $Y2=1.38
r189 46 56 2.63384 $w=3.35e-07 $l=8.5e-08 $layer=LI1_cond $X=7.972 $Y=1.695
+ $X2=7.972 $Y2=1.61
r190 46 56 0.516019 $w=3.33e-07 $l=1.5e-08 $layer=LI1_cond $X=7.972 $Y=1.595
+ $X2=7.972 $Y2=1.61
r191 46 51 7.39628 $w=3.33e-07 $l=2.15e-07 $layer=LI1_cond $X=7.972 $Y=1.595
+ $X2=7.972 $Y2=1.38
r192 44 46 5.17472 $w=1.7e-07 $l=1.67e-07 $layer=LI1_cond $X=7.805 $Y=1.695
+ $X2=7.972 $Y2=1.695
r193 44 45 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=7.805 $Y=1.695
+ $X2=7.07 $Y2=1.695
r194 43 45 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.985 $Y=1.61
+ $X2=7.07 $Y2=1.695
r195 42 43 77.3102 $w=1.68e-07 $l=1.185e-06 $layer=LI1_cond $X=6.985 $Y=0.425
+ $X2=6.985 $Y2=1.61
r196 40 55 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.77 $Y=0.34
+ $X2=4.77 $Y2=0.505
r197 39 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.77
+ $Y=0.34 $X2=4.77 $Y2=0.34
r198 37 42 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.9 $Y=0.34
+ $X2=6.985 $Y2=0.425
r199 37 39 138.963 $w=1.68e-07 $l=2.13e-06 $layer=LI1_cond $X=6.9 $Y=0.34
+ $X2=4.77 $Y2=0.34
r200 35 50 32.3493 $w=3.3e-07 $l=1.85e-07 $layer=POLY_cond $X=8.16 $Y=1.38
+ $X2=7.975 $Y2=1.38
r201 35 36 1.50692 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.16 $Y=1.38
+ $X2=8.16 $Y2=1.215
r202 32 33 141.011 $w=1.5e-07 $l=2.75e-07 $layer=POLY_cond $X=4.585 $Y=1.22
+ $X2=4.86 $Y2=1.22
r203 30 32 135.883 $w=1.5e-07 $l=2.65e-07 $layer=POLY_cond $X=4.32 $Y=1.22
+ $X2=4.585 $Y2=1.22
r204 27 29 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=15.825 $Y=3.075
+ $X2=15.825 $Y2=2.525
r205 26 29 492.255 $w=1.5e-07 $l=9.6e-07 $layer=POLY_cond $X=15.825 $Y=1.565
+ $X2=15.825 $Y2=2.525
r206 24 26 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=15.75 $Y=1.49
+ $X2=15.825 $Y2=1.565
r207 24 25 89.734 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=15.75 $Y=1.49
+ $X2=15.575 $Y2=1.49
r208 20 25 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=15.5 $Y=1.415
+ $X2=15.575 $Y2=1.49
r209 20 22 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=15.5 $Y=1.415
+ $X2=15.5 $Y2=0.705
r210 18 27 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=15.75 $Y=3.15
+ $X2=15.825 $Y2=3.075
r211 18 19 3763.7 $w=1.5e-07 $l=7.34e-06 $layer=POLY_cond $X=15.75 $Y=3.15
+ $X2=8.41 $Y2=3.15
r212 14 36 30.2679 $w=2e-07 $l=1.05e-07 $layer=POLY_cond $X=8.265 $Y=1.215
+ $X2=8.16 $Y2=1.215
r213 14 16 394.83 $w=1.5e-07 $l=7.7e-07 $layer=POLY_cond $X=8.265 $Y=1.215
+ $X2=8.265 $Y2=0.445
r214 11 19 29.1797 $w=1.5e-07 $l=1.58114e-07 $layer=POLY_cond $X=8.285 $Y=3.075
+ $X2=8.41 $Y2=3.15
r215 11 13 216.155 $w=2.5e-07 $l=8.7e-07 $layer=POLY_cond $X=8.285 $Y=3.075
+ $X2=8.285 $Y2=2.205
r216 10 36 30.2679 $w=2e-07 $l=3.87492e-07 $layer=POLY_cond $X=8.285 $Y=1.545
+ $X2=8.16 $Y2=1.215
r217 10 13 163.979 $w=2.5e-07 $l=6.6e-07 $layer=POLY_cond $X=8.285 $Y=1.545
+ $X2=8.285 $Y2=2.205
r218 9 33 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.86 $Y=1.145
+ $X2=4.86 $Y2=1.22
r219 9 55 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=4.86 $Y=1.145
+ $X2=4.86 $Y2=0.505
r220 4 32 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.585 $Y=1.295
+ $X2=4.585 $Y2=1.22
r221 4 6 574.298 $w=1.5e-07 $l=1.12e-06 $layer=POLY_cond $X=4.585 $Y=1.295
+ $X2=4.585 $Y2=2.415
r222 1 30 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.32 $Y=1.145
+ $X2=4.32 $Y2=1.22
r223 1 3 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=4.32 $Y=1.145
+ $X2=4.32 $Y2=0.825
.ends

.subckt PM_SKY130_FD_SC_LP__SRSDFRTN_1%A_742_63# 1 2 9 12 13 14 18 19 24 25 27
+ 30 32 35 38 40 42 43 46 48 50 51 52 54 55 56 58 59 60 61 66 67 68 70 73 75 76
+ 78 80 82 89 91 97 99
c300 99 0 6.73578e-20 $X=13.02 $Y=1.48
c301 97 0 1.98227e-19 $X=5.5 $Y=1.77
c302 89 0 4.1238e-20 $X=12.98 $Y=1.57
c303 82 0 1.92106e-19 $X=5.215 $Y=1.77
c304 60 0 1.07616e-19 $X=9.58 $Y=2.81
c305 46 0 5.16263e-20 $X=13.74 $Y=1.1
c306 24 0 1.55617e-19 $X=5.49 $Y=2.305
r307 96 97 1.74861 $w=3.3e-07 $l=1e-08 $layer=POLY_cond $X=5.49 $Y=1.77 $X2=5.5
+ $Y2=1.77
r308 90 102 45.9078 $w=4.1e-07 $l=1.65e-07 $layer=POLY_cond $X=13.02 $Y=1.57
+ $X2=13.02 $Y2=1.735
r309 90 99 12.2083 $w=4.1e-07 $l=9e-08 $layer=POLY_cond $X=13.02 $Y=1.57
+ $X2=13.02 $Y2=1.48
r310 89 91 10.5918 $w=3.58e-07 $l=2.3e-07 $layer=LI1_cond $X=12.98 $Y=1.555
+ $X2=12.75 $Y2=1.555
r311 89 90 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=12.98
+ $Y=1.57 $X2=12.98 $Y2=1.57
r312 83 96 48.0869 $w=3.3e-07 $l=2.75e-07 $layer=POLY_cond $X=5.215 $Y=1.77
+ $X2=5.49 $Y2=1.77
r313 83 93 14.8632 $w=3.3e-07 $l=8.5e-08 $layer=POLY_cond $X=5.215 $Y=1.77
+ $X2=5.13 $Y2=1.77
r314 82 85 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=5.215 $Y=1.77
+ $X2=5.215 $Y2=1.935
r315 82 83 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.215
+ $Y=1.77 $X2=5.215 $Y2=1.77
r316 80 91 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=12.08 $Y=1.46
+ $X2=12.75 $Y2=1.46
r317 77 80 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=11.995 $Y=1.545
+ $X2=12.08 $Y2=1.46
r318 77 78 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=11.995 $Y=1.545
+ $X2=11.995 $Y2=1.95
r319 75 78 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=11.91 $Y=2.035
+ $X2=11.995 $Y2=1.95
r320 75 76 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=11.91 $Y=2.035
+ $X2=11.445 $Y2=2.035
r321 71 76 8.05333 $w=1.95e-07 $l=1.39194e-07 $layer=LI1_cond $X=11.32 $Y=2.065
+ $X2=11.445 $Y2=2.035
r322 71 73 10.372 $w=2.48e-07 $l=2.25e-07 $layer=LI1_cond $X=11.32 $Y=2.18
+ $X2=11.32 $Y2=2.405
r323 70 71 23.7744 $w=1.95e-07 $l=3.8e-07 $layer=LI1_cond $X=10.94 $Y=2.065
+ $X2=11.32 $Y2=2.065
r324 69 70 48.6043 $w=1.68e-07 $l=7.45e-07 $layer=LI1_cond $X=10.94 $Y=1.265
+ $X2=10.94 $Y2=2.01
r325 67 70 5.55076 $w=1.95e-07 $l=9.88686e-08 $layer=LI1_cond $X=10.855 $Y=2.095
+ $X2=10.94 $Y2=2.065
r326 67 68 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=10.855 $Y=2.095
+ $X2=10.675 $Y2=2.095
r327 65 68 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.59 $Y=2.18
+ $X2=10.675 $Y2=2.095
r328 65 66 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=10.59 $Y=2.18
+ $X2=10.59 $Y2=2.725
r329 61 69 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=10.855 $Y=1.1
+ $X2=10.94 $Y2=1.265
r330 61 63 9.42908 $w=3.28e-07 $l=2.7e-07 $layer=LI1_cond $X=10.855 $Y=1.1
+ $X2=10.585 $Y2=1.1
r331 59 66 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.505 $Y=2.81
+ $X2=10.59 $Y2=2.725
r332 59 60 60.3476 $w=1.68e-07 $l=9.25e-07 $layer=LI1_cond $X=10.505 $Y=2.81
+ $X2=9.58 $Y2=2.81
r333 58 60 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.495 $Y=2.725
+ $X2=9.58 $Y2=2.81
r334 57 58 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=9.495 $Y=2.52
+ $X2=9.495 $Y2=2.725
r335 55 57 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.41 $Y=2.435
+ $X2=9.495 $Y2=2.52
r336 55 56 141.246 $w=1.68e-07 $l=2.165e-06 $layer=LI1_cond $X=9.41 $Y=2.435
+ $X2=7.245 $Y2=2.435
r337 53 56 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.16 $Y=2.52
+ $X2=7.245 $Y2=2.435
r338 53 54 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=7.16 $Y=2.52
+ $X2=7.16 $Y2=2.905
r339 51 54 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.075 $Y=2.99
+ $X2=7.16 $Y2=2.905
r340 51 52 110.583 $w=1.68e-07 $l=1.695e-06 $layer=LI1_cond $X=7.075 $Y=2.99
+ $X2=5.38 $Y2=2.99
r341 50 52 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.295 $Y=2.905
+ $X2=5.38 $Y2=2.99
r342 50 85 63.2834 $w=1.68e-07 $l=9.7e-07 $layer=LI1_cond $X=5.295 $Y=2.905
+ $X2=5.295 $Y2=1.935
r343 44 46 117.936 $w=1.5e-07 $l=2.3e-07 $layer=POLY_cond $X=13.51 $Y=1.1
+ $X2=13.74 $Y2=1.1
r344 40 46 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=13.74 $Y=1.025
+ $X2=13.74 $Y2=1.1
r345 40 42 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=13.74 $Y=1.025
+ $X2=13.74 $Y2=0.595
r346 36 48 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=13.51 $Y=1.555
+ $X2=13.51 $Y2=1.48
r347 36 38 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=13.51 $Y=1.555
+ $X2=13.51 $Y2=2.345
r348 35 48 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=13.51 $Y=1.405
+ $X2=13.51 $Y2=1.48
r349 34 44 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=13.51 $Y=1.175
+ $X2=13.51 $Y2=1.1
r350 34 35 117.936 $w=1.5e-07 $l=2.3e-07 $layer=POLY_cond $X=13.51 $Y=1.175
+ $X2=13.51 $Y2=1.405
r351 33 99 26.4667 $w=1.5e-07 $l=2.05e-07 $layer=POLY_cond $X=13.225 $Y=1.48
+ $X2=13.02 $Y2=1.48
r352 32 48 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=13.435 $Y=1.48
+ $X2=13.51 $Y2=1.48
r353 32 33 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=13.435 $Y=1.48
+ $X2=13.225 $Y2=1.48
r354 30 102 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=13.15 $Y=2.345
+ $X2=13.15 $Y2=1.735
r355 25 97 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.5 $Y=1.605
+ $X2=5.5 $Y2=1.77
r356 25 27 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=5.5 $Y=1.605
+ $X2=5.5 $Y2=1.285
r357 22 24 394.83 $w=1.5e-07 $l=7.7e-07 $layer=POLY_cond $X=5.49 $Y=3.075
+ $X2=5.49 $Y2=2.305
r358 21 96 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.49 $Y=1.935
+ $X2=5.49 $Y2=1.77
r359 21 24 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=5.49 $Y=1.935
+ $X2=5.49 $Y2=2.305
r360 20 43 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.205 $Y=3.15
+ $X2=5.13 $Y2=3.15
r361 19 22 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.415 $Y=3.15
+ $X2=5.49 $Y2=3.075
r362 19 20 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=5.415 $Y=3.15
+ $X2=5.205 $Y2=3.15
r363 16 43 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.13 $Y=3.075
+ $X2=5.13 $Y2=3.15
r364 16 18 394.83 $w=1.5e-07 $l=7.7e-07 $layer=POLY_cond $X=5.13 $Y=3.075
+ $X2=5.13 $Y2=2.305
r365 15 93 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.13 $Y=1.935
+ $X2=5.13 $Y2=1.77
r366 15 18 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=5.13 $Y=1.935
+ $X2=5.13 $Y2=2.305
r367 13 43 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.055 $Y=3.15
+ $X2=5.13 $Y2=3.15
r368 13 14 612.755 $w=1.5e-07 $l=1.195e-06 $layer=POLY_cond $X=5.055 $Y=3.15
+ $X2=3.86 $Y2=3.15
r369 9 12 902.468 $w=1.5e-07 $l=1.76e-06 $layer=POLY_cond $X=3.785 $Y=0.655
+ $X2=3.785 $Y2=2.415
r370 7 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.785 $Y=3.075
+ $X2=3.86 $Y2=3.15
r371 7 12 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=3.785 $Y=3.075
+ $X2=3.785 $Y2=2.415
r372 2 73 600 $w=1.7e-07 $l=3.73497e-07 $layer=licon1_PDIFF $count=1 $X=11.22
+ $Y=2.095 $X2=11.36 $Y2=2.405
r373 1 63 182 $w=1.7e-07 $l=6.83667e-07 $layer=licon1_NDIFF $count=1 $X=10.44
+ $Y=0.485 $X2=10.585 $Y2=1.1
.ends

.subckt PM_SKY130_FD_SC_LP__SRSDFRTN_1%A_666_89# 1 2 7 9 12 14 16 17 19 23 25 29
+ 33 38 42 43 44 45 48 54 55 59 62
c197 62 0 3.2762e-19 $X=6.32 $Y=1.77
c198 59 0 3.44653e-19 $X=6.29 $Y=1.77
c199 55 0 5.93087e-20 $X=14.16 $Y=2.035
c200 42 0 2.62237e-20 $X=6.335 $Y=2.035
c201 38 0 5.16263e-20 $X=14.22 $Y=1.29
c202 33 0 1.69305e-19 $X=3.465 $Y=1.43
r203 61 62 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.32
+ $Y=1.77 $X2=6.32 $Y2=1.77
r204 59 61 4.82 $w=3e-07 $l=3e-08 $layer=POLY_cond $X=6.29 $Y=1.77 $X2=6.32
+ $Y2=1.77
r205 58 59 32.9367 $w=3e-07 $l=2.05e-07 $layer=POLY_cond $X=6.085 $Y=1.77
+ $X2=6.29 $Y2=1.77
r206 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.16 $Y=2.035
+ $X2=14.16 $Y2=2.035
r207 52 62 7.44872 $w=4.08e-07 $l=2.65e-07 $layer=LI1_cond $X=6.36 $Y=2.035
+ $X2=6.36 $Y2=1.77
r208 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=2.035
+ $X2=6.48 $Y2=2.035
r209 48 67 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=3.61 $Y=2.035
+ $X2=3.61 $Y2=2.405
r210 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=2.035
+ $X2=3.6 $Y2=2.035
r211 45 51 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.625 $Y=2.035
+ $X2=6.48 $Y2=2.035
r212 44 54 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=14.015 $Y=2.035
+ $X2=14.16 $Y2=2.035
r213 44 45 9.14602 $w=1.4e-07 $l=7.39e-06 $layer=MET1_cond $X=14.015 $Y=2.035
+ $X2=6.625 $Y2=2.035
r214 43 47 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.745 $Y=2.035
+ $X2=3.6 $Y2=2.035
r215 42 51 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.335 $Y=2.035
+ $X2=6.48 $Y2=2.035
r216 42 43 3.20544 $w=1.4e-07 $l=2.59e-06 $layer=MET1_cond $X=6.335 $Y=2.035
+ $X2=3.745 $Y2=2.035
r217 41 55 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=14.16 $Y=1.455
+ $X2=14.16 $Y2=2.035
r218 39 63 11.6613 $w=3.72e-07 $l=9e-08 $layer=POLY_cond $X=14.177 $Y=1.29
+ $X2=14.177 $Y2=1.2
r219 38 41 8.53353 $w=2.83e-07 $l=1.65e-07 $layer=LI1_cond $X=14.217 $Y=1.29
+ $X2=14.217 $Y2=1.455
r220 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=14.22
+ $Y=1.29 $X2=14.22 $Y2=1.29
r221 35 48 20.283 $w=2.48e-07 $l=4.4e-07 $layer=LI1_cond $X=3.61 $Y=1.595
+ $X2=3.61 $Y2=2.035
r222 33 35 6.37886 $w=3.53e-07 $l=1.65e-07 $layer=LI1_cond $X=3.557 $Y=1.43
+ $X2=3.557 $Y2=1.595
r223 27 29 215.362 $w=1.5e-07 $l=4.2e-07 $layer=POLY_cond $X=14.68 $Y=1.125
+ $X2=14.68 $Y2=0.705
r224 26 63 24.0971 $w=1.5e-07 $l=2.18e-07 $layer=POLY_cond $X=14.395 $Y=1.2
+ $X2=14.177 $Y2=1.2
r225 25 27 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=14.605 $Y=1.2
+ $X2=14.68 $Y2=1.125
r226 25 26 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=14.605 $Y=1.2
+ $X2=14.395 $Y2=1.2
r227 21 63 27.4257 $w=3.72e-07 $l=1.76562e-07 $layer=POLY_cond $X=14.32 $Y=1.125
+ $X2=14.177 $Y2=1.2
r228 21 23 215.362 $w=1.5e-07 $l=4.2e-07 $layer=POLY_cond $X=14.32 $Y=1.125
+ $X2=14.32 $Y2=0.705
r229 17 39 53.3397 $w=3.72e-07 $l=3.38637e-07 $layer=POLY_cond $X=14.035
+ $Y=1.565 $X2=14.177 $Y2=1.29
r230 17 19 292.277 $w=1.5e-07 $l=5.7e-07 $layer=POLY_cond $X=14.035 $Y=1.565
+ $X2=14.035 $Y2=2.135
r231 14 59 18.9685 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.29 $Y=1.605
+ $X2=6.29 $Y2=1.77
r232 14 16 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=6.29 $Y=1.605
+ $X2=6.29 $Y2=1.285
r233 10 58 7.1379 $w=2.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.085 $Y=1.935
+ $X2=6.085 $Y2=1.77
r234 10 12 163.979 $w=2.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.085 $Y=1.935
+ $X2=6.085 $Y2=2.595
r235 7 58 24.9033 $w=3e-07 $l=2.29783e-07 $layer=POLY_cond $X=5.93 $Y=1.605
+ $X2=6.085 $Y2=1.77
r236 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=5.93 $Y=1.605
+ $X2=5.93 $Y2=1.285
r237 2 67 600 $w=1.7e-07 $l=3.75566e-07 $layer=licon1_PDIFF $count=1 $X=3.425
+ $Y=2.095 $X2=3.57 $Y2=2.405
r238 1 33 182 $w=1.7e-07 $l=1.05033e-06 $layer=licon1_NDIFF $count=1 $X=3.33
+ $Y=0.445 $X2=3.465 $Y2=1.43
.ends

.subckt PM_SKY130_FD_SC_LP__SRSDFRTN_1%A_1343_51# 1 2 3 4 15 17 20 24 26 27 30
+ 33 34 36 37 40 44 45 46 48 49 50 52 54 55 59 62 63 65 66 70 71 74 78
c217 59 0 2.79523e-20 $X=14.5 $Y=1.86
c218 55 0 1.89357e-19 $X=14.53 $Y=0.34
c219 45 0 1.44185e-19 $X=11.535 $Y=0.34
c220 26 0 1.3264e-19 $X=6.795 $Y=0.915
r221 72 74 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=14.5 $Y=1.71
+ $X2=14.615 $Y2=1.71
r222 69 71 8.51103 $w=3.58e-07 $l=1.65e-07 $layer=LI1_cond $X=13.49 $Y=0.435
+ $X2=13.655 $Y2=0.435
r223 69 70 8.51103 $w=3.58e-07 $l=1.65e-07 $layer=LI1_cond $X=13.49 $Y=0.435
+ $X2=13.325 $Y2=0.435
r224 65 66 8.79328 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=9.795 $Y=1.715
+ $X2=9.63 $Y2=1.715
r225 62 74 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=14.615 $Y=1.625
+ $X2=14.615 $Y2=1.71
r226 61 62 78.2888 $w=1.68e-07 $l=1.2e-06 $layer=LI1_cond $X=14.615 $Y=0.425
+ $X2=14.615 $Y2=1.625
r227 57 72 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=14.5 $Y=1.795
+ $X2=14.5 $Y2=1.71
r228 57 59 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=14.5 $Y=1.795
+ $X2=14.5 $Y2=1.86
r229 55 61 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=14.53 $Y=0.34
+ $X2=14.615 $Y2=0.425
r230 55 71 57.0856 $w=1.68e-07 $l=8.75e-07 $layer=LI1_cond $X=14.53 $Y=0.34
+ $X2=13.655 $Y2=0.34
r231 54 70 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=12.595 $Y=0.34
+ $X2=13.325 $Y2=0.34
r232 51 54 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=12.51 $Y=0.425
+ $X2=12.595 $Y2=0.34
r233 51 52 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=12.51 $Y=0.425
+ $X2=12.51 $Y2=0.615
r234 49 52 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=12.425 $Y=0.7
+ $X2=12.51 $Y2=0.615
r235 49 50 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=12.425 $Y=0.7
+ $X2=11.705 $Y2=0.7
r236 48 50 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=11.62 $Y=0.615
+ $X2=11.705 $Y2=0.7
r237 47 48 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=11.62 $Y=0.425
+ $X2=11.62 $Y2=0.615
r238 45 47 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=11.535 $Y=0.34
+ $X2=11.62 $Y2=0.425
r239 45 46 108.952 $w=1.68e-07 $l=1.67e-06 $layer=LI1_cond $X=11.535 $Y=0.34
+ $X2=9.865 $Y2=0.34
r240 42 44 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=9.7 $Y=0.875
+ $X2=9.7 $Y2=0.465
r241 41 46 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=9.7 $Y=0.425
+ $X2=9.865 $Y2=0.34
r242 41 44 1.3969 $w=3.28e-07 $l=4e-08 $layer=LI1_cond $X=9.7 $Y=0.425 $X2=9.7
+ $Y2=0.465
r243 40 66 72.0909 $w=1.68e-07 $l=1.105e-06 $layer=LI1_cond $X=8.525 $Y=1.755
+ $X2=9.63 $Y2=1.755
r244 38 63 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.525 $Y=0.96
+ $X2=8.44 $Y2=0.96
r245 37 42 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=9.535 $Y=0.96
+ $X2=9.7 $Y2=0.875
r246 37 38 65.8931 $w=1.68e-07 $l=1.01e-06 $layer=LI1_cond $X=9.535 $Y=0.96
+ $X2=8.525 $Y2=0.96
r247 36 40 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.44 $Y=1.67
+ $X2=8.525 $Y2=1.755
r248 35 63 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.44 $Y=1.045
+ $X2=8.44 $Y2=0.96
r249 35 36 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=8.44 $Y=1.045
+ $X2=8.44 $Y2=1.67
r250 33 63 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.355 $Y=0.96
+ $X2=8.44 $Y2=0.96
r251 33 34 51.2139 $w=1.68e-07 $l=7.85e-07 $layer=LI1_cond $X=8.355 $Y=0.96
+ $X2=7.57 $Y2=0.96
r252 31 78 40.7992 $w=2.54e-07 $l=2.15e-07 $layer=POLY_cond $X=7.405 $Y=1.282
+ $X2=7.19 $Y2=1.282
r253 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.405
+ $Y=1.275 $X2=7.405 $Y2=1.275
r254 28 34 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=7.405 $Y=1.045
+ $X2=7.57 $Y2=0.96
r255 28 30 8.03218 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=7.405 $Y=1.045
+ $X2=7.405 $Y2=1.275
r256 26 27 69.5192 $w=1.6e-07 $l=1.5e-07 $layer=POLY_cond $X=6.795 $Y=0.915
+ $X2=6.795 $Y2=1.065
r257 22 78 15.087 $w=1.5e-07 $l=1.72e-07 $layer=POLY_cond $X=7.19 $Y=1.11
+ $X2=7.19 $Y2=1.282
r258 22 24 264.074 $w=1.5e-07 $l=5.15e-07 $layer=POLY_cond $X=7.19 $Y=1.11
+ $X2=7.19 $Y2=0.595
r259 18 78 64.5197 $w=2.54e-07 $l=4.17636e-07 $layer=POLY_cond $X=6.85 $Y=1.455
+ $X2=7.19 $Y2=1.282
r260 18 20 283.237 $w=2.5e-07 $l=1.14e-06 $layer=POLY_cond $X=6.85 $Y=1.455
+ $X2=6.85 $Y2=2.595
r261 17 18 9.48819 $w=2.54e-07 $l=1.73205e-07 $layer=POLY_cond $X=6.8 $Y=1.305
+ $X2=6.85 $Y2=1.455
r262 17 27 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=6.8 $Y=1.305
+ $X2=6.8 $Y2=1.065
r263 15 26 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=6.79 $Y=0.595
+ $X2=6.79 $Y2=0.915
r264 4 59 300 $w=1.7e-07 $l=4.56782e-07 $layer=licon1_PDIFF $count=2 $X=14.11
+ $Y=1.715 $X2=14.5 $Y2=1.86
r265 3 65 600 $w=1.7e-07 $l=2.58795e-07 $layer=licon1_PDIFF $count=1 $X=9.56
+ $Y=1.705 $X2=9.795 $Y2=1.755
r266 2 69 182 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_NDIFF $count=1 $X=13.345
+ $Y=0.275 $X2=13.49 $Y2=0.435
r267 1 44 182 $w=1.7e-07 $l=2.91719e-07 $layer=licon1_NDIFF $count=1 $X=9.56
+ $Y=0.235 $X2=9.7 $Y2=0.465
.ends

.subckt PM_SKY130_FD_SC_LP__SRSDFRTN_1%A_1724_21# 1 2 9 13 15 18 19 20 22 23 24
+ 25 27 29 33 35 38 41 43 46
c154 43 0 9.16269e-20 $X=9.025 $Y=1.357
c155 27 0 7.79314e-20 $X=12.415 $Y=2.59
c156 25 0 2.05894e-19 $X=12.415 $Y=2.075
c157 19 0 1.87318e-19 $X=11.195 $Y=0.68
c158 13 0 1.07616e-19 $X=8.745 $Y=2.205
c159 9 0 3.01101e-20 $X=8.695 $Y=0.445
r160 41 49 30.7525 $w=4.05e-07 $l=1.65e-07 $layer=POLY_cond $X=8.822 $Y=1.355
+ $X2=8.822 $Y2=1.52
r161 41 48 45.79 $w=4.05e-07 $l=1.65e-07 $layer=POLY_cond $X=8.822 $Y=1.355
+ $X2=8.822 $Y2=1.19
r162 40 43 8.53353 $w=2.83e-07 $l=1.65e-07 $layer=LI1_cond $X=8.86 $Y=1.357
+ $X2=9.025 $Y2=1.357
r163 40 41 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.86
+ $Y=1.355 $X2=8.86 $Y2=1.355
r164 37 38 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=13.4 $Y=1.125
+ $X2=13.4 $Y2=1.905
r165 36 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.095 $Y=1.04
+ $X2=12.93 $Y2=1.04
r166 35 37 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=13.315 $Y=1.04
+ $X2=13.4 $Y2=1.125
r167 35 36 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=13.315 $Y=1.04
+ $X2=13.095 $Y2=1.04
r168 31 46 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=12.93 $Y=0.955
+ $X2=12.93 $Y2=1.04
r169 31 33 6.80989 $w=3.28e-07 $l=1.95e-07 $layer=LI1_cond $X=12.93 $Y=0.955
+ $X2=12.93 $Y2=0.76
r170 30 45 4.5891 $w=1.7e-07 $l=2.07123e-07 $layer=LI1_cond $X=12.58 $Y=1.99
+ $X2=12.415 $Y2=1.895
r171 29 38 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=13.315 $Y=1.99
+ $X2=13.4 $Y2=1.905
r172 29 30 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=13.315 $Y=1.99
+ $X2=12.58 $Y2=1.99
r173 25 45 3.17707 $w=3.3e-07 $l=1.8e-07 $layer=LI1_cond $X=12.415 $Y=2.075
+ $X2=12.415 $Y2=1.895
r174 25 27 17.9851 $w=3.28e-07 $l=5.15e-07 $layer=LI1_cond $X=12.415 $Y=2.075
+ $X2=12.415 $Y2=2.59
r175 23 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.765 $Y=1.04
+ $X2=12.93 $Y2=1.04
r176 23 24 91.3369 $w=1.68e-07 $l=1.4e-06 $layer=LI1_cond $X=12.765 $Y=1.04
+ $X2=11.365 $Y2=1.04
r177 22 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=11.28 $Y=0.955
+ $X2=11.365 $Y2=1.04
r178 21 22 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=11.28 $Y=0.765
+ $X2=11.28 $Y2=0.955
r179 19 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=11.195 $Y=0.68
+ $X2=11.28 $Y2=0.765
r180 19 20 64.5882 $w=1.68e-07 $l=9.9e-07 $layer=LI1_cond $X=11.195 $Y=0.68
+ $X2=10.205 $Y2=0.68
r181 17 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.12 $Y=0.765
+ $X2=10.205 $Y2=0.68
r182 17 18 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=10.12 $Y=0.765
+ $X2=10.12 $Y2=1.215
r183 15 18 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.035 $Y=1.3
+ $X2=10.12 $Y2=1.215
r184 15 43 65.8931 $w=1.68e-07 $l=1.01e-06 $layer=LI1_cond $X=10.035 $Y=1.3
+ $X2=9.025 $Y2=1.3
r185 13 49 170.191 $w=2.5e-07 $l=6.85e-07 $layer=POLY_cond $X=8.745 $Y=2.205
+ $X2=8.745 $Y2=1.52
r186 9 48 382.011 $w=1.5e-07 $l=7.45e-07 $layer=POLY_cond $X=8.695 $Y=0.445
+ $X2=8.695 $Y2=1.19
r187 2 45 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=12.275
+ $Y=1.735 $X2=12.415 $Y2=1.88
r188 2 27 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=12.275
+ $Y=1.735 $X2=12.415 $Y2=2.59
r189 1 33 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=12.79
+ $Y=0.485 $X2=12.93 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_LP__SRSDFRTN_1%A_1113_419# 1 2 3 10 12 15 17 19 20 21 23
+ 27 29 31 34 35 36 39 43 44 48
c144 29 0 1.59996e-19 $X=5.715 $Y=1.36
c145 15 0 9.59449e-20 $X=9.435 $Y=2.205
r146 44 49 30.6007 $w=3.3e-07 $l=1.75e-07 $layer=POLY_cond $X=10.245 $Y=2.39
+ $X2=10.07 $Y2=2.39
r147 43 44 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.245
+ $Y=2.39 $X2=10.245 $Y2=2.39
r148 41 43 9.49071 $w=2.53e-07 $l=2.1e-07 $layer=LI1_cond $X=10.207 $Y=2.18
+ $X2=10.207 $Y2=2.39
r149 39 41 7.17723 $w=1.7e-07 $l=1.64085e-07 $layer=LI1_cond $X=10.08 $Y=2.095
+ $X2=10.207 $Y2=2.18
r150 39 48 123.631 $w=1.68e-07 $l=1.895e-06 $layer=LI1_cond $X=10.08 $Y=2.095
+ $X2=8.185 $Y2=2.095
r151 36 38 55.8684 $w=2.28e-07 $l=1.115e-06 $layer=LI1_cond $X=6.905 $Y=2.065
+ $X2=8.02 $Y2=2.065
r152 35 48 6.56993 $w=2.28e-07 $l=1.15e-07 $layer=LI1_cond $X=8.07 $Y=2.065
+ $X2=8.185 $Y2=2.065
r153 35 38 2.50531 $w=2.28e-07 $l=5e-08 $layer=LI1_cond $X=8.07 $Y=2.065
+ $X2=8.02 $Y2=2.065
r154 33 36 7.01789 $w=2.3e-07 $l=1.51658e-07 $layer=LI1_cond $X=6.82 $Y=2.18
+ $X2=6.905 $Y2=2.065
r155 33 34 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=6.82 $Y=2.18
+ $X2=6.82 $Y2=2.32
r156 32 47 5.39226 $w=1.7e-07 $l=2.7225e-07 $layer=LI1_cond $X=5.985 $Y=2.405
+ $X2=5.767 $Y2=2.527
r157 31 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.735 $Y=2.405
+ $X2=6.82 $Y2=2.32
r158 31 32 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=6.735 $Y=2.405
+ $X2=5.985 $Y2=2.405
r159 27 47 3.28293 $w=4.35e-07 $l=2.07e-07 $layer=LI1_cond $X=5.767 $Y=2.32
+ $X2=5.767 $Y2=2.527
r160 27 29 25.4332 $w=4.33e-07 $l=9.6e-07 $layer=LI1_cond $X=5.767 $Y=2.32
+ $X2=5.767 $Y2=1.36
r161 25 26 10.8072 $w=2.23e-07 $l=5e-08 $layer=POLY_cond $X=9.435 $Y=0.915
+ $X2=9.485 $Y2=0.915
r162 24 25 67.0045 $w=2.23e-07 $l=3.1e-07 $layer=POLY_cond $X=9.125 $Y=0.915
+ $X2=9.435 $Y2=0.915
r163 23 49 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.07 $Y=2.225
+ $X2=10.07 $Y2=2.39
r164 22 23 594.809 $w=1.5e-07 $l=1.16e-06 $layer=POLY_cond $X=10.07 $Y=1.065
+ $X2=10.07 $Y2=2.225
r165 21 26 21.3961 $w=2.23e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.56 $Y=0.99
+ $X2=9.485 $Y2=0.915
r166 20 22 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.995 $Y=0.99
+ $X2=10.07 $Y2=1.065
r167 20 21 223.053 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=9.995 $Y=0.99
+ $X2=9.56 $Y2=0.99
r168 17 26 12.0837 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=9.485 $Y=0.765
+ $X2=9.485 $Y2=0.915
r169 17 19 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=9.485 $Y=0.765
+ $X2=9.485 $Y2=0.445
r170 13 25 0.0270875 $w=2.5e-07 $l=1.5e-07 $layer=POLY_cond $X=9.435 $Y=1.065
+ $X2=9.435 $Y2=0.915
r171 13 15 283.237 $w=2.5e-07 $l=1.14e-06 $layer=POLY_cond $X=9.435 $Y=1.065
+ $X2=9.435 $Y2=2.205
r172 10 24 12.0837 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=9.125 $Y=0.765
+ $X2=9.125 $Y2=0.915
r173 10 12 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=9.125 $Y=0.765
+ $X2=9.125 $Y2=0.445
r174 3 38 600 $w=1.7e-07 $l=4.17852e-07 $layer=licon1_PDIFF $count=1 $X=7.895
+ $Y=1.705 $X2=8.02 $Y2=2.065
r175 2 47 600 $w=1.7e-07 $l=4.18509e-07 $layer=licon1_PDIFF $count=1 $X=5.565
+ $Y=2.095 $X2=5.82 $Y2=2.405
r176 1 29 182 $w=1.7e-07 $l=3.4803e-07 $layer=licon1_NDIFF $count=1 $X=5.575
+ $Y=1.075 $X2=5.715 $Y2=1.36
.ends

.subckt PM_SKY130_FD_SC_LP__SRSDFRTN_1%CLK_N 3 5 7 9 10 14
r48 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.52
+ $Y=1.695 $X2=10.52 $Y2=1.695
r49 10 14 8.08732 $w=2.83e-07 $l=2e-07 $layer=LI1_cond $X=10.32 $Y=1.697
+ $X2=10.52 $Y2=1.697
r50 9 13 39.1141 $w=4.55e-07 $l=3.2e-07 $layer=POLY_cond $X=10.84 $Y=1.757
+ $X2=10.52 $Y2=1.757
r51 5 9 54.2108 $w=2.25e-07 $l=2.95506e-07 $layer=POLY_cond $X=11.145 $Y=1.985
+ $X2=10.99 $Y2=1.757
r52 5 7 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=11.145 $Y=1.985
+ $X2=11.145 $Y2=2.415
r53 1 9 53.9965 $w=2.25e-07 $l=2.61828e-07 $layer=POLY_cond $X=10.915 $Y=1.53
+ $X2=10.99 $Y2=1.757
r54 1 3 428.16 $w=1.5e-07 $l=8.35e-07 $layer=POLY_cond $X=10.915 $Y=1.53
+ $X2=10.915 $Y2=0.695
.ends

.subckt PM_SKY130_FD_SC_LP__SRSDFRTN_1%SLEEP_B 1 3 6 8 10 11 13 14 16 17 18 19
+ 21 22 27
c97 18 0 1.44185e-19 $X=12.4 $Y=1.09
c98 11 0 4.1238e-20 $X=12.15 $Y=1.625
c99 8 0 1.87318e-19 $X=11.665 $Y=1.015
c100 6 0 1.38537e-19 $X=11.575 $Y=2.415
r101 29 30 41.7446 $w=5.6e-07 $l=4.85e-07 $layer=POLY_cond $X=11.665 $Y=1.32
+ $X2=12.15 $Y2=1.32
r102 28 29 7.74643 $w=5.6e-07 $l=9e-08 $layer=POLY_cond $X=11.575 $Y=1.32
+ $X2=11.665 $Y2=1.32
r103 26 28 15.4929 $w=5.6e-07 $l=1.8e-07 $layer=POLY_cond $X=11.395 $Y=1.32
+ $X2=11.575 $Y2=1.32
r104 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.395
+ $Y=1.46 $X2=11.395 $Y2=1.46
r105 24 26 7.74643 $w=5.6e-07 $l=9e-08 $layer=POLY_cond $X=11.305 $Y=1.32
+ $X2=11.395 $Y2=1.32
r106 22 27 6.47263 $w=3.63e-07 $l=2.05e-07 $layer=LI1_cond $X=11.377 $Y=1.665
+ $X2=11.377 $Y2=1.46
r107 19 21 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=12.715 $Y=1.015
+ $X2=12.715 $Y2=0.695
r108 17 19 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=12.64 $Y=1.09
+ $X2=12.715 $Y2=1.015
r109 17 18 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=12.64 $Y=1.09
+ $X2=12.4 $Y2=1.09
r110 14 18 35.7626 $w=5.6e-07 $l=1.06066e-07 $layer=POLY_cond $X=12.325 $Y=1.015
+ $X2=12.4 $Y2=1.09
r111 14 30 15.0625 $w=5.6e-07 $l=3.82623e-07 $layer=POLY_cond $X=12.325 $Y=1.015
+ $X2=12.15 $Y2=1.32
r112 14 16 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=12.325 $Y=1.015
+ $X2=12.325 $Y2=0.695
r113 11 30 21.6522 $w=2.5e-07 $l=3.05e-07 $layer=POLY_cond $X=12.15 $Y=1.625
+ $X2=12.15 $Y2=1.32
r114 11 13 117.608 $w=2.5e-07 $l=6.1e-07 $layer=POLY_cond $X=12.15 $Y=1.625
+ $X2=12.15 $Y2=2.235
r115 8 29 34.2947 $w=1.5e-07 $l=3.05e-07 $layer=POLY_cond $X=11.665 $Y=1.015
+ $X2=11.665 $Y2=1.32
r116 8 10 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=11.665 $Y=1.015
+ $X2=11.665 $Y2=0.695
r117 4 28 34.2947 $w=1.5e-07 $l=3.05e-07 $layer=POLY_cond $X=11.575 $Y=1.625
+ $X2=11.575 $Y2=1.32
r118 4 6 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=11.575 $Y=1.625
+ $X2=11.575 $Y2=2.415
r119 1 24 34.2947 $w=1.5e-07 $l=3.05e-07 $layer=POLY_cond $X=11.305 $Y=1.015
+ $X2=11.305 $Y2=1.32
r120 1 3 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=11.305 $Y=1.015
+ $X2=11.305 $Y2=0.695
.ends

.subckt PM_SKY130_FD_SC_LP__SRSDFRTN_1%A_2999_73# 1 2 9 13 15 22 25 26 30 35
c74 15 0 2.79523e-20 $X=15.875 $Y=1.97
c75 13 0 1.19187e-19 $X=15.395 $Y=2.525
c76 9 0 1.89357e-19 $X=15.07 $Y=0.705
r77 27 30 3.38954 $w=3.38e-07 $l=1e-07 $layer=LI1_cond $X=16.12 $Y=0.765
+ $X2=16.22 $Y2=0.765
r78 25 26 6.46576 $w=2.5e-07 $l=2.0106e-07 $layer=LI1_cond $X=16.12 $Y=1.805
+ $X2=16.04 $Y2=1.97
r79 24 27 4.80115 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=16.12 $Y=0.935
+ $X2=16.12 $Y2=0.765
r80 24 25 56.7594 $w=1.68e-07 $l=8.7e-07 $layer=LI1_cond $X=16.12 $Y=0.935
+ $X2=16.12 $Y2=1.805
r81 20 26 6.46576 $w=2.5e-07 $l=1.65e-07 $layer=LI1_cond $X=16.04 $Y=2.135
+ $X2=16.04 $Y2=1.97
r82 20 22 13.6198 $w=3.28e-07 $l=3.9e-07 $layer=LI1_cond $X=16.04 $Y=2.135
+ $X2=16.04 $Y2=2.525
r83 18 35 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=15.375 $Y=1.97
+ $X2=15.395 $Y2=1.97
r84 18 32 53.3327 $w=3.3e-07 $l=3.05e-07 $layer=POLY_cond $X=15.375 $Y=1.97
+ $X2=15.07 $Y2=1.97
r85 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=15.375
+ $Y=1.97 $X2=15.375 $Y2=1.97
r86 15 26 0.364692 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=15.875 $Y=1.97
+ $X2=16.04 $Y2=1.97
r87 15 17 17.4613 $w=3.28e-07 $l=5e-07 $layer=LI1_cond $X=15.875 $Y=1.97
+ $X2=15.375 $Y2=1.97
r88 11 35 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=15.395 $Y=2.135
+ $X2=15.395 $Y2=1.97
r89 11 13 199.979 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=15.395 $Y=2.135
+ $X2=15.395 $Y2=2.525
r90 7 32 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=15.07 $Y=1.805
+ $X2=15.07 $Y2=1.97
r91 7 9 564.043 $w=1.5e-07 $l=1.1e-06 $layer=POLY_cond $X=15.07 $Y=1.805
+ $X2=15.07 $Y2=0.705
r92 2 22 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=15.9
+ $Y=2.315 $X2=16.04 $Y2=2.525
r93 1 30 182 $w=1.7e-07 $l=3.76497e-07 $layer=licon1_NDIFF $count=1 $X=15.965
+ $Y=0.495 $X2=16.22 $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_LP__SRSDFRTN_1%A_2717_427# 1 2 7 9 10 11 14 17 18 20 21
+ 24 28 30 33 36 37 39 41 42 43 45 46 47 52 60 62 65
c159 52 0 1.98676e-19 $X=16.645 $Y=1.06
c160 41 0 5.93087e-20 $X=14.955 $Y=1.965
r161 58 60 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=14.84 $Y=2.05
+ $X2=14.955 $Y2=2.05
r162 53 65 3.2901 $w=5.86e-07 $l=4e-08 $layer=POLY_cond $X=16.502 $Y=1.06
+ $X2=16.502 $Y2=1.1
r163 53 63 7.40273 $w=5.86e-07 $l=9e-08 $layer=POLY_cond $X=16.502 $Y=1.06
+ $X2=16.502 $Y2=0.97
r164 52 62 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=16.645 $Y=1.06
+ $X2=16.645 $Y2=0.895
r165 52 53 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=16.645
+ $Y=1.06 $X2=16.645 $Y2=1.06
r166 48 62 30.6631 $w=1.68e-07 $l=4.7e-07 $layer=LI1_cond $X=16.565 $Y=0.425
+ $X2=16.565 $Y2=0.895
r167 46 48 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=16.48 $Y=0.34
+ $X2=16.565 $Y2=0.425
r168 46 47 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=16.48 $Y=0.34
+ $X2=15.79 $Y2=0.34
r169 44 47 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=15.705 $Y=0.425
+ $X2=15.79 $Y2=0.34
r170 44 45 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=15.705 $Y=0.425
+ $X2=15.705 $Y2=1.105
r171 42 45 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=15.62 $Y=1.19
+ $X2=15.705 $Y2=1.105
r172 42 43 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=15.62 $Y=1.19
+ $X2=15.04 $Y2=1.19
r173 41 60 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=14.955 $Y=1.965
+ $X2=14.955 $Y2=2.05
r174 40 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=14.955 $Y=1.275
+ $X2=15.04 $Y2=1.19
r175 40 41 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=14.955 $Y=1.275
+ $X2=14.955 $Y2=1.965
r176 38 58 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=14.84 $Y=2.135
+ $X2=14.84 $Y2=2.05
r177 38 39 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=14.84 $Y=2.135
+ $X2=14.84 $Y2=2.565
r178 36 39 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=14.755 $Y=2.65
+ $X2=14.84 $Y2=2.565
r179 36 37 55.4545 $w=1.68e-07 $l=8.5e-07 $layer=LI1_cond $X=14.755 $Y=2.65
+ $X2=13.905 $Y2=2.65
r180 33 35 25.3537 $w=2.48e-07 $l=5.5e-07 $layer=LI1_cond $X=13.78 $Y=1.86
+ $X2=13.78 $Y2=2.41
r181 31 37 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=13.78 $Y=2.565
+ $X2=13.905 $Y2=2.65
r182 31 35 7.14515 $w=2.48e-07 $l=1.55e-07 $layer=LI1_cond $X=13.78 $Y=2.565
+ $X2=13.78 $Y2=2.41
r183 30 57 8.68475 $w=2.95e-07 $l=2.86182e-07 $layer=LI1_cond $X=13.78 $Y=0.955
+ $X2=13.99 $Y2=0.775
r184 30 33 41.7184 $w=2.48e-07 $l=9.05e-07 $layer=LI1_cond $X=13.78 $Y=0.955
+ $X2=13.78 $Y2=1.86
r185 26 28 379.447 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=17.22 $Y=2.035
+ $X2=17.22 $Y2=2.775
r186 22 24 205.106 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=17.2 $Y=0.895
+ $X2=17.2 $Y2=0.495
r187 20 26 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=17.145 $Y=1.96
+ $X2=17.22 $Y2=2.035
r188 20 21 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=17.145 $Y=1.96
+ $X2=16.825 $Y2=1.96
r189 19 63 35.4637 $w=1.5e-07 $l=3.23e-07 $layer=POLY_cond $X=16.825 $Y=0.97
+ $X2=16.502 $Y2=0.97
r190 18 22 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=17.125 $Y=0.97
+ $X2=17.2 $Y2=0.895
r191 18 19 153.83 $w=1.5e-07 $l=3e-07 $layer=POLY_cond $X=17.125 $Y=0.97
+ $X2=16.825 $Y2=0.97
r192 17 21 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=16.75 $Y=1.885
+ $X2=16.825 $Y2=1.96
r193 16 65 79.0899 $w=2.93e-07 $l=5.75799e-07 $layer=POLY_cond $X=16.75 $Y=1.565
+ $X2=16.502 $Y2=1.1
r194 16 17 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=16.75 $Y=1.565
+ $X2=16.75 $Y2=1.885
r195 12 65 79.0899 $w=2.93e-07 $l=5.75396e-07 $layer=POLY_cond $X=16.255
+ $Y=1.565 $X2=16.502 $Y2=1.1
r196 12 14 492.255 $w=1.5e-07 $l=9.6e-07 $layer=POLY_cond $X=16.255 $Y=1.565
+ $X2=16.255 $Y2=2.525
r197 10 65 35.4637 $w=1.5e-07 $l=3.22e-07 $layer=POLY_cond $X=16.18 $Y=1.1
+ $X2=16.502 $Y2=1.1
r198 10 11 110.245 $w=1.5e-07 $l=2.15e-07 $layer=POLY_cond $X=16.18 $Y=1.1
+ $X2=15.965 $Y2=1.1
r199 7 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=15.89 $Y=1.025
+ $X2=15.965 $Y2=1.1
r200 7 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=15.89 $Y=1.025
+ $X2=15.89 $Y2=0.705
r201 2 35 600 $w=1.7e-07 $l=3.745e-07 $layer=licon1_PDIFF $count=1 $X=13.585
+ $Y=2.135 $X2=13.82 $Y2=2.41
r202 2 33 600 $w=1.7e-07 $l=3.745e-07 $layer=licon1_PDIFF $count=1 $X=13.585
+ $Y=2.135 $X2=13.82 $Y2=1.86
r203 1 57 182 $w=1.7e-07 $l=5.70833e-07 $layer=licon1_NDIFF $count=1 $X=13.815
+ $Y=0.275 $X2=13.99 $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_LP__SRSDFRTN_1%A_3368_57# 1 2 9 13 15 16 17 19 22 27 31
+ 34 35
c64 15 0 1.98676e-19 $X=17.67 $Y=1.48
r65 31 33 10.7321 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=16.985 $Y=0.495
+ $X2=16.985 $Y2=0.725
r66 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=17.46
+ $Y=1.48 $X2=17.46 $Y2=1.48
r67 25 35 0.718145 $w=3.3e-07 $l=9.5e-08 $layer=LI1_cond $X=17.17 $Y=1.48
+ $X2=17.075 $Y2=1.48
r68 25 27 10.1275 $w=3.28e-07 $l=2.9e-07 $layer=LI1_cond $X=17.17 $Y=1.48
+ $X2=17.46 $Y2=1.48
r69 23 35 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=17.075 $Y=1.645
+ $X2=17.075 $Y2=1.48
r70 23 34 46.1148 $w=1.88e-07 $l=7.9e-07 $layer=LI1_cond $X=17.075 $Y=1.645
+ $X2=17.075 $Y2=2.435
r71 22 35 8.26956 $w=1.8e-07 $l=1.69926e-07 $layer=LI1_cond $X=17.065 $Y=1.315
+ $X2=17.075 $Y2=1.48
r72 22 33 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=17.065 $Y=1.315
+ $X2=17.065 $Y2=0.725
r73 17 34 7.81899 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=17.005 $Y=2.6
+ $X2=17.005 $Y2=2.435
r74 17 19 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=17.005 $Y=2.6
+ $X2=17.005 $Y2=2.755
r75 15 28 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=17.67 $Y=1.48
+ $X2=17.46 $Y2=1.48
r76 15 16 5.03009 $w=3.3e-07 $l=8e-08 $layer=POLY_cond $X=17.67 $Y=1.48
+ $X2=17.75 $Y2=1.48
r77 11 16 37.0704 $w=1.5e-07 $l=1.67481e-07 $layer=POLY_cond $X=17.755 $Y=1.645
+ $X2=17.75 $Y2=1.48
r78 11 13 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=17.755 $Y=1.645
+ $X2=17.755 $Y2=2.465
r79 7 16 37.0704 $w=1.5e-07 $l=1.67481e-07 $layer=POLY_cond $X=17.745 $Y=1.315
+ $X2=17.75 $Y2=1.48
r80 7 9 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=17.745 $Y=1.315
+ $X2=17.745 $Y2=0.705
r81 2 19 600 $w=1.7e-07 $l=3.61248e-07 $layer=licon1_PDIFF $count=1 $X=16.87
+ $Y=2.455 $X2=17.005 $Y2=2.755
r82 1 31 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=16.84
+ $Y=0.285 $X2=16.985 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__SRSDFRTN_1%VPWR 1 2 3 4 5 6 21 25 29 33 37 41 46 47
+ 49 50 52 53 55 56 57 75 86 92 93 96 99
c169 93 0 3.57021e-19 $X=18 $Y=3.33
r170 99 100 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=17.52 $Y=3.33
+ $X2=17.52 $Y2=3.33
r171 96 97 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=15.6 $Y=3.33
+ $X2=15.6 $Y2=3.33
r172 93 100 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=18 $Y=3.33
+ $X2=17.52 $Y2=3.33
r173 92 93 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=18 $Y=3.33 $X2=18
+ $Y2=3.33
r174 90 99 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=17.625 $Y=3.33
+ $X2=17.5 $Y2=3.33
r175 90 92 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=17.625 $Y=3.33
+ $X2=18 $Y2=3.33
r176 89 100 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=17.04 $Y=3.33
+ $X2=17.52 $Y2=3.33
r177 88 89 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=17.04 $Y=3.33
+ $X2=17.04 $Y2=3.33
r178 86 99 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=17.375 $Y=3.33
+ $X2=17.5 $Y2=3.33
r179 86 88 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=17.375 $Y=3.33
+ $X2=17.04 $Y2=3.33
r180 85 89 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=16.08 $Y=3.33
+ $X2=17.04 $Y2=3.33
r181 85 97 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=16.08 $Y=3.33
+ $X2=15.6 $Y2=3.33
r182 84 85 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=16.08 $Y=3.33
+ $X2=16.08 $Y2=3.33
r183 82 96 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=15.695 $Y=3.33
+ $X2=15.57 $Y2=3.33
r184 82 84 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=15.695 $Y=3.33
+ $X2=16.08 $Y2=3.33
r185 81 97 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=15.12 $Y=3.33
+ $X2=15.6 $Y2=3.33
r186 80 81 0.808696 $w=1.7e-07 $l=1.955e-06 $layer=mcon $count=11 $X=15.12
+ $Y=3.33 $X2=15.12 $Y2=3.33
r187 77 80 688.941 $w=1.68e-07 $l=1.056e-05 $layer=LI1_cond $X=4.56 $Y=3.33
+ $X2=15.12 $Y2=3.33
r188 77 78 0.808696 $w=1.7e-07 $l=1.955e-06 $layer=mcon $count=11 $X=4.56
+ $Y=3.33 $X2=4.56 $Y2=3.33
r189 75 96 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=15.445 $Y=3.33
+ $X2=15.57 $Y2=3.33
r190 75 80 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=15.445 $Y=3.33
+ $X2=15.12 $Y2=3.33
r191 74 78 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r192 73 74 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r193 71 74 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=4.08 $Y2=3.33
r194 70 73 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=3.12 $Y=3.33
+ $X2=4.08 $Y2=3.33
r195 70 71 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r196 68 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r197 67 68 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r198 65 68 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r199 64 67 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r200 64 65 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r201 61 65 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r202 60 61 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r203 57 81 1.67241 $w=4.9e-07 $l=6e-06 $layer=MET1_cond $X=9.12 $Y=3.33
+ $X2=15.12 $Y2=3.33
r204 57 78 1.27103 $w=4.9e-07 $l=4.56e-06 $layer=MET1_cond $X=9.12 $Y=3.33
+ $X2=4.56 $Y2=3.33
r205 55 84 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=16.385 $Y=3.33
+ $X2=16.08 $Y2=3.33
r206 55 56 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=16.385 $Y=3.33
+ $X2=16.51 $Y2=3.33
r207 54 88 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=16.635 $Y=3.33
+ $X2=17.04 $Y2=3.33
r208 54 56 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=16.635 $Y=3.33
+ $X2=16.51 $Y2=3.33
r209 52 73 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=4.285 $Y=3.33
+ $X2=4.08 $Y2=3.33
r210 52 53 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.285 $Y=3.33
+ $X2=4.37 $Y2=3.33
r211 51 77 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=4.455 $Y=3.33
+ $X2=4.56 $Y2=3.33
r212 51 53 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.455 $Y=3.33
+ $X2=4.37 $Y2=3.33
r213 49 67 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=2.67 $Y=3.33 $X2=2.64
+ $Y2=3.33
r214 49 50 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.67 $Y=3.33
+ $X2=2.795 $Y2=3.33
r215 48 70 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=2.92 $Y=3.33 $X2=3.12
+ $Y2=3.33
r216 48 50 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.92 $Y=3.33
+ $X2=2.795 $Y2=3.33
r217 46 60 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=0.78 $Y=3.33 $X2=0.72
+ $Y2=3.33
r218 46 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.78 $Y=3.33
+ $X2=0.945 $Y2=3.33
r219 45 64 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=1.11 $Y=3.33 $X2=1.2
+ $Y2=3.33
r220 45 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.11 $Y=3.33
+ $X2=0.945 $Y2=3.33
r221 41 44 44.7148 $w=2.48e-07 $l=9.7e-07 $layer=LI1_cond $X=17.5 $Y=1.98
+ $X2=17.5 $Y2=2.95
r222 39 99 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=17.5 $Y=3.245
+ $X2=17.5 $Y2=3.33
r223 39 44 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=17.5 $Y=3.245
+ $X2=17.5 $Y2=2.95
r224 35 56 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=16.51 $Y=3.245
+ $X2=16.51 $Y2=3.33
r225 35 37 33.1904 $w=2.48e-07 $l=7.2e-07 $layer=LI1_cond $X=16.51 $Y=3.245
+ $X2=16.51 $Y2=2.525
r226 31 96 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=15.57 $Y=3.245
+ $X2=15.57 $Y2=3.33
r227 31 33 32.9599 $w=2.48e-07 $l=7.15e-07 $layer=LI1_cond $X=15.57 $Y=3.245
+ $X2=15.57 $Y2=2.53
r228 27 53 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.37 $Y=3.245
+ $X2=4.37 $Y2=3.33
r229 27 29 65.5668 $w=1.68e-07 $l=1.005e-06 $layer=LI1_cond $X=4.37 $Y=3.245
+ $X2=4.37 $Y2=2.24
r230 23 50 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.795 $Y=3.245
+ $X2=2.795 $Y2=3.33
r231 23 25 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=2.795 $Y=3.245
+ $X2=2.795 $Y2=2.95
r232 19 47 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.945 $Y=3.245
+ $X2=0.945 $Y2=3.33
r233 19 21 22.525 $w=3.28e-07 $l=6.45e-07 $layer=LI1_cond $X=0.945 $Y=3.245
+ $X2=0.945 $Y2=2.6
r234 6 44 600 $w=1.7e-07 $l=6.05227e-07 $layer=licon1_PDIFF $count=1 $X=17.295
+ $Y=2.455 $X2=17.54 $Y2=2.95
r235 6 41 300 $w=1.7e-07 $l=5.84808e-07 $layer=licon1_PDIFF $count=2 $X=17.295
+ $Y=2.455 $X2=17.54 $Y2=1.98
r236 5 37 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=16.33
+ $Y=2.315 $X2=16.47 $Y2=2.525
r237 4 33 600 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_PDIFF $count=1 $X=15.47
+ $Y=2.315 $X2=15.61 $Y2=2.53
r238 3 29 300 $w=1.7e-07 $l=5.77971e-07 $layer=licon1_PDIFF $count=2 $X=3.86
+ $Y=2.095 $X2=4.37 $Y2=2.24
r239 2 25 600 $w=1.7e-07 $l=5.60647e-07 $layer=licon1_PDIFF $count=1 $X=2.695
+ $Y=2.455 $X2=2.835 $Y2=2.95
r240 1 21 300 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=2 $X=0.735
+ $Y=2.455 $X2=0.945 $Y2=2.6
.ends

.subckt PM_SKY130_FD_SC_LP__SRSDFRTN_1%A_305_97# 1 2 3 4 13 19 21 22 24 25 26 28
+ 30 31 32 34 35 36 38 41 43 45 46 48 49 50 51 52 53 54
c183 53 0 6.31736e-20 $X=4.8 $Y=2.105
c184 34 0 1.92529e-19 $X=4.03 $Y=2.905
r185 54 57 7.85757 $w=3.28e-07 $l=2.25e-07 $layer=LI1_cond $X=6.505 $Y=1.02
+ $X2=6.505 $Y2=1.245
r186 49 54 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.34 $Y=1.02
+ $X2=6.505 $Y2=1.02
r187 49 50 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=6.34 $Y=1.02
+ $X2=5.38 $Y2=1.02
r188 47 50 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.295 $Y=1.105
+ $X2=5.38 $Y2=1.02
r189 47 48 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=5.295 $Y=1.105
+ $X2=5.295 $Y2=1.265
r190 45 48 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.21 $Y=1.35
+ $X2=5.295 $Y2=1.265
r191 45 46 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=5.21 $Y=1.35
+ $X2=4.805 $Y2=1.35
r192 41 53 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=4.8 $Y=2.27
+ $X2=4.8 $Y2=2.105
r193 41 43 5.5876 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=4.8 $Y=2.27 $X2=4.8
+ $Y2=2.43
r194 39 52 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.72 $Y=1.905
+ $X2=4.72 $Y2=1.82
r195 39 53 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=4.72 $Y=1.905
+ $X2=4.72 $Y2=2.105
r196 38 52 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.72 $Y=1.735
+ $X2=4.72 $Y2=1.82
r197 37 46 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.72 $Y=1.435
+ $X2=4.805 $Y2=1.35
r198 37 38 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=4.72 $Y=1.435
+ $X2=4.72 $Y2=1.735
r199 35 52 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.635 $Y=1.82
+ $X2=4.72 $Y2=1.82
r200 35 36 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=4.635 $Y=1.82
+ $X2=4.115 $Y2=1.82
r201 33 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.03 $Y=1.905
+ $X2=4.115 $Y2=1.82
r202 33 34 65.2406 $w=1.68e-07 $l=1e-06 $layer=LI1_cond $X=4.03 $Y=1.905
+ $X2=4.03 $Y2=2.905
r203 31 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.945 $Y=2.99
+ $X2=4.03 $Y2=2.905
r204 31 32 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=3.945 $Y=2.99
+ $X2=3.26 $Y2=2.99
r205 30 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.175 $Y=2.905
+ $X2=3.26 $Y2=2.99
r206 29 51 5.16603 $w=1.7e-07 $l=9.66954e-08 $layer=LI1_cond $X=3.175 $Y=2.615
+ $X2=3.15 $Y2=2.53
r207 29 30 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=3.175 $Y=2.615
+ $X2=3.175 $Y2=2.905
r208 28 51 5.16603 $w=1.7e-07 $l=9.66954e-08 $layer=LI1_cond $X=3.125 $Y=2.445
+ $X2=3.15 $Y2=2.53
r209 27 28 65.8931 $w=1.68e-07 $l=1.01e-06 $layer=LI1_cond $X=3.125 $Y=1.435
+ $X2=3.125 $Y2=2.445
r210 25 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.04 $Y=1.35
+ $X2=3.125 $Y2=1.435
r211 25 26 58.3904 $w=1.68e-07 $l=8.95e-07 $layer=LI1_cond $X=3.04 $Y=1.35
+ $X2=2.145 $Y2=1.35
r212 24 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.06 $Y=1.265
+ $X2=2.145 $Y2=1.35
r213 23 24 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=2.06 $Y=0.925
+ $X2=2.06 $Y2=1.265
r214 21 51 1.34256 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=3.04 $Y=2.53
+ $X2=3.15 $Y2=2.53
r215 21 22 72.4171 $w=1.68e-07 $l=1.11e-06 $layer=LI1_cond $X=3.04 $Y=2.53
+ $X2=1.93 $Y2=2.53
r216 17 22 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.765 $Y=2.615
+ $X2=1.93 $Y2=2.53
r217 17 19 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=1.765 $Y=2.615
+ $X2=1.765 $Y2=2.76
r218 13 23 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.975 $Y=0.76
+ $X2=2.06 $Y2=0.925
r219 13 15 10.826 $w=3.28e-07 $l=3.1e-07 $layer=LI1_cond $X=1.975 $Y=0.76
+ $X2=1.665 $Y2=0.76
r220 4 43 600 $w=1.7e-07 $l=3.98905e-07 $layer=licon1_PDIFF $count=1 $X=4.66
+ $Y=2.095 $X2=4.8 $Y2=2.43
r221 3 19 600 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_PDIFF $count=1 $X=1.625
+ $Y=2.455 $X2=1.765 $Y2=2.76
r222 2 57 182 $w=1.7e-07 $l=2.29565e-07 $layer=licon1_NDIFF $count=1 $X=6.365
+ $Y=1.075 $X2=6.505 $Y2=1.245
r223 1 15 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=1.525
+ $Y=0.485 $X2=1.665 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_LP__SRSDFRTN_1%KAPWR 1 2 3 4 15 17 18 20 30 38 41 46 50
+ 52 61 62
c185 62 0 7.79314e-20 $X=11.905 $Y=2.802
r186 50 52 0.314267 $w=2.7e-07 $l=5.75e-07 $layer=MET1_cond $X=8.545 $Y=2.81
+ $X2=9.12 $Y2=2.81
r187 41 44 7.25612 $w=4.03e-07 $l=2.55e-07 $layer=LI1_cond $X=11.847 $Y=2.52
+ $X2=11.847 $Y2=2.775
r188 35 50 0.0645018 $w=2.81e-07 $l=1.48946e-07 $layer=MET1_cond $X=8.4 $Y=2.802
+ $X2=8.545 $Y2=2.81
r189 34 38 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=8.4 $Y=2.855
+ $X2=9.075 $Y2=2.855
r190 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=2.775
+ $X2=8.4 $Y2=2.775
r191 31 46 0.0645018 $w=2.81e-07 $l=1.48946e-07 $layer=MET1_cond $X=7.92
+ $Y=2.802 $X2=7.775 $Y2=2.81
r192 30 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=2.775
+ $X2=7.92 $Y2=2.775
r193 27 30 12.5721 $w=3.83e-07 $l=4.2e-07 $layer=LI1_cond $X=7.5 $Y=2.882
+ $X2=7.92 $Y2=2.882
r194 20 62 0.072812 $w=2.85e-07 $l=1.45e-07 $layer=MET1_cond $X=11.76 $Y=2.802
+ $X2=11.905 $Y2=2.802
r195 20 61 0.072812 $w=2.85e-07 $l=1.45e-07 $layer=MET1_cond $X=11.76 $Y=2.802
+ $X2=11.615 $Y2=2.802
r196 20 35 0.106762 $w=2.81e-07 $l=2.4e-07 $layer=MET1_cond $X=8.16 $Y=2.802
+ $X2=8.4 $Y2=2.802
r197 20 31 0.106762 $w=2.81e-07 $l=2.4e-07 $layer=MET1_cond $X=8.16 $Y=2.802
+ $X2=7.92 $Y2=2.802
r198 20 62 1.7118 $w=2.7e-07 $l=3.132e-06 $layer=MET1_cond $X=15.037 $Y=2.81
+ $X2=11.905 $Y2=2.81
r199 20 61 0.838957 $w=2.7e-07 $l=1.535e-06 $layer=MET1_cond $X=10.08 $Y=2.81
+ $X2=11.615 $Y2=2.81
r200 20 52 0.52469 $w=2.7e-07 $l=9.6e-07 $layer=MET1_cond $X=10.08 $Y=2.81
+ $X2=9.12 $Y2=2.81
r201 20 46 2.10586 $w=2.7e-07 $l=3.853e-06 $layer=MET1_cond $X=3.922 $Y=2.81
+ $X2=7.775 $Y2=2.81
r202 20 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.76 $Y=2.775
+ $X2=11.76 $Y2=2.775
r203 19 44 3.6992 $w=4.03e-07 $l=1.3e-07 $layer=LI1_cond $X=11.847 $Y=2.905
+ $X2=11.847 $Y2=2.775
r204 17 19 8.41448 $w=1.7e-07 $l=2.40778e-07 $layer=LI1_cond $X=11.645 $Y=2.99
+ $X2=11.847 $Y2=2.905
r205 17 18 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=11.645 $Y=2.99
+ $X2=11.015 $Y2=2.99
r206 13 18 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.93 $Y=2.905
+ $X2=11.015 $Y2=2.99
r207 13 15 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=10.93 $Y=2.905
+ $X2=10.93 $Y2=2.55
r208 4 41 600 $w=1.7e-07 $l=5.29622e-07 $layer=licon1_PDIFF $count=1 $X=11.65
+ $Y=2.095 $X2=11.885 $Y2=2.52
r209 3 15 600 $w=1.7e-07 $l=5.22494e-07 $layer=licon1_PDIFF $count=1 $X=10.785
+ $Y=2.095 $X2=10.93 $Y2=2.55
r210 2 38 600 $w=1.7e-07 $l=1.2483e-06 $layer=licon1_PDIFF $count=1 $X=8.87
+ $Y=1.705 $X2=9.075 $Y2=2.855
r211 1 27 600 $w=1.7e-07 $l=1.01408e-06 $layer=licon1_PDIFF $count=1 $X=6.975
+ $Y=2.095 $X2=7.5 $Y2=2.88
.ends

.subckt PM_SKY130_FD_SC_LP__SRSDFRTN_1%A_2562_427# 1 2 9 11 12 15
r35 13 15 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=15.18 $Y=2.905
+ $X2=15.18 $Y2=2.53
r36 11 13 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=15.095 $Y=2.99
+ $X2=15.18 $Y2=2.905
r37 11 12 130.155 $w=1.68e-07 $l=1.995e-06 $layer=LI1_cond $X=15.095 $Y=2.99
+ $X2=13.1 $Y2=2.99
r38 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=12.935 $Y=2.905
+ $X2=13.1 $Y2=2.99
r39 7 9 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=12.935 $Y=2.905
+ $X2=12.935 $Y2=2.41
r40 2 15 600 $w=1.7e-07 $l=2.78209e-07 $layer=licon1_PDIFF $count=1 $X=15.035
+ $Y=2.315 $X2=15.18 $Y2=2.53
r41 1 9 600 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_PDIFF $count=1 $X=12.81
+ $Y=2.135 $X2=12.935 $Y2=2.41
.ends

.subckt PM_SKY130_FD_SC_LP__SRSDFRTN_1%Q 1 2 7 8 9 10 11 18
r16 11 32 31.5227 $w=3.38e-07 $l=9.3e-07 $layer=LI1_cond $X=17.965 $Y=1.98
+ $X2=17.965 $Y2=2.91
r17 10 11 10.677 $w=3.38e-07 $l=3.15e-07 $layer=LI1_cond $X=17.965 $Y=1.665
+ $X2=17.965 $Y2=1.98
r18 9 10 12.5413 $w=3.38e-07 $l=3.7e-07 $layer=LI1_cond $X=17.965 $Y=1.295
+ $X2=17.965 $Y2=1.665
r19 8 9 12.5413 $w=3.38e-07 $l=3.7e-07 $layer=LI1_cond $X=17.965 $Y=0.925
+ $X2=17.965 $Y2=1.295
r20 7 8 12.5413 $w=3.38e-07 $l=3.7e-07 $layer=LI1_cond $X=17.965 $Y=0.555
+ $X2=17.965 $Y2=0.925
r21 7 18 4.23692 $w=3.38e-07 $l=1.25e-07 $layer=LI1_cond $X=17.965 $Y=0.555
+ $X2=17.965 $Y2=0.43
r22 2 32 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=17.83
+ $Y=1.835 $X2=17.97 $Y2=2.91
r23 2 11 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=17.83
+ $Y=1.835 $X2=17.97 $Y2=1.98
r24 1 18 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=17.82
+ $Y=0.285 $X2=17.96 $Y2=0.43
.ends

.subckt PM_SKY130_FD_SC_LP__SRSDFRTN_1%VGND 1 2 3 4 5 6 7 24 28 30 34 38 42 46
+ 51 52 53 55 60 68 83 87 97 98 101 104 108 114 117 120
c161 98 0 3.39925e-20 $X=18 $Y=0
r162 120 121 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=17.52 $Y=0
+ $X2=17.52 $Y2=0
r163 117 118 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=15.12 $Y=0
+ $X2=15.12 $Y2=0
r164 114 115 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.88 $Y=0
+ $X2=8.88 $Y2=0
r165 109 115 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.92 $Y=0
+ $X2=8.88 $Y2=0
r166 108 111 9.7783 $w=3.28e-07 $l=2.8e-07 $layer=LI1_cond $X=7.945 $Y=0
+ $X2=7.945 $Y2=0.28
r167 108 109 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=0
+ $X2=7.92 $Y2=0
r168 104 105 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0
+ $X2=4.08 $Y2=0
r169 101 102 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0
+ $X2=0.72 $Y2=0
r170 98 121 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=18 $Y=0 $X2=17.52
+ $Y2=0
r171 97 98 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=18 $Y=0 $X2=18
+ $Y2=0
r172 95 120 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=17.615 $Y=0
+ $X2=17.49 $Y2=0
r173 95 97 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=17.615 $Y=0 $X2=18
+ $Y2=0
r174 94 121 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=17.04 $Y=0
+ $X2=17.52 $Y2=0
r175 93 94 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=17.04 $Y=0
+ $X2=17.04 $Y2=0
r176 91 94 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=15.6 $Y=0
+ $X2=17.04 $Y2=0
r177 91 118 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=15.6 $Y=0
+ $X2=15.12 $Y2=0
r178 90 93 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=15.6 $Y=0
+ $X2=17.04 $Y2=0
r179 90 91 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=15.6 $Y=0 $X2=15.6
+ $Y2=0
r180 88 117 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=15.45 $Y=0
+ $X2=15.285 $Y2=0
r181 88 90 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=15.45 $Y=0 $X2=15.6
+ $Y2=0
r182 87 120 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=17.365 $Y=0
+ $X2=17.49 $Y2=0
r183 87 93 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=17.365 $Y=0
+ $X2=17.04 $Y2=0
r184 86 118 0.802756 $w=4.9e-07 $l=2.88e-06 $layer=MET1_cond $X=12.24 $Y=0
+ $X2=15.12 $Y2=0
r185 85 86 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=12.24 $Y=0
+ $X2=12.24 $Y2=0
r186 83 117 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=15.12 $Y=0
+ $X2=15.285 $Y2=0
r187 83 85 187.893 $w=1.68e-07 $l=2.88e-06 $layer=LI1_cond $X=15.12 $Y=0
+ $X2=12.24 $Y2=0
r188 82 86 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.76 $Y=0
+ $X2=12.24 $Y2=0
r189 81 82 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=11.76 $Y=0
+ $X2=11.76 $Y2=0
r190 79 82 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=9.36 $Y=0
+ $X2=11.76 $Y2=0
r191 78 81 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=9.36 $Y=0 $X2=11.76
+ $Y2=0
r192 78 79 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=9.36 $Y=0 $X2=9.36
+ $Y2=0
r193 76 114 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.075 $Y=0
+ $X2=8.95 $Y2=0
r194 76 78 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=9.075 $Y=0
+ $X2=9.36 $Y2=0
r195 75 109 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0
+ $X2=7.92 $Y2=0
r196 74 75 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=7.44 $Y=0
+ $X2=7.44 $Y2=0
r197 72 75 0.802756 $w=4.9e-07 $l=2.88e-06 $layer=MET1_cond $X=4.56 $Y=0
+ $X2=7.44 $Y2=0
r198 72 105 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0
+ $X2=4.08 $Y2=0
r199 71 74 187.893 $w=1.68e-07 $l=2.88e-06 $layer=LI1_cond $X=4.56 $Y=0 $X2=7.44
+ $Y2=0
r200 71 72 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=4.56 $Y=0
+ $X2=4.56 $Y2=0
r201 69 104 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.165 $Y=0 $X2=4
+ $Y2=0
r202 69 71 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=4.165 $Y=0
+ $X2=4.56 $Y2=0
r203 68 108 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.78 $Y=0
+ $X2=7.945 $Y2=0
r204 68 74 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=7.78 $Y=0 $X2=7.44
+ $Y2=0
r205 67 105 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r206 66 67 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r207 64 67 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=1.2 $Y=0 $X2=3.6
+ $Y2=0
r208 64 102 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r209 63 66 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=3.6
+ $Y2=0
r210 63 64 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r211 61 101 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.865 $Y=0 $X2=0.7
+ $Y2=0
r212 61 63 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=0.865 $Y=0 $X2=1.2
+ $Y2=0
r213 60 104 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.835 $Y=0 $X2=4
+ $Y2=0
r214 60 66 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=3.835 $Y=0 $X2=3.6
+ $Y2=0
r215 58 102 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0
+ $X2=0.72 $Y2=0
r216 57 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r217 55 101 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.535 $Y=0 $X2=0.7
+ $Y2=0
r218 55 57 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.535 $Y=0 $X2=0.24
+ $Y2=0
r219 53 79 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=9.12 $Y=0
+ $X2=9.36 $Y2=0
r220 53 115 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=9.12 $Y=0
+ $X2=8.88 $Y2=0
r221 51 81 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=11.91 $Y=0 $X2=11.76
+ $Y2=0
r222 51 52 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=11.91 $Y=0
+ $X2=12.035 $Y2=0
r223 50 85 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=12.16 $Y=0 $X2=12.24
+ $Y2=0
r224 50 52 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=12.16 $Y=0
+ $X2=12.035 $Y2=0
r225 46 48 25.3537 $w=2.48e-07 $l=5.5e-07 $layer=LI1_cond $X=17.49 $Y=0.43
+ $X2=17.49 $Y2=0.98
r226 44 120 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=17.49 $Y=0.085
+ $X2=17.49 $Y2=0
r227 44 46 15.9037 $w=2.48e-07 $l=3.45e-07 $layer=LI1_cond $X=17.49 $Y=0.085
+ $X2=17.49 $Y2=0.43
r228 40 117 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=15.285 $Y=0.085
+ $X2=15.285 $Y2=0
r229 40 42 21.652 $w=3.28e-07 $l=6.2e-07 $layer=LI1_cond $X=15.285 $Y=0.085
+ $X2=15.285 $Y2=0.705
r230 36 52 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=12.035 $Y=0.085
+ $X2=12.035 $Y2=0
r231 36 38 8.98906 $w=2.48e-07 $l=1.95e-07 $layer=LI1_cond $X=12.035 $Y=0.085
+ $X2=12.035 $Y2=0.28
r232 32 114 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=8.95 $Y=0.085
+ $X2=8.95 $Y2=0
r233 32 34 16.5952 $w=2.48e-07 $l=3.6e-07 $layer=LI1_cond $X=8.95 $Y=0.085
+ $X2=8.95 $Y2=0.445
r234 31 108 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.11 $Y=0
+ $X2=7.945 $Y2=0
r235 30 114 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.825 $Y=0
+ $X2=8.95 $Y2=0
r236 30 31 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=8.825 $Y=0
+ $X2=8.11 $Y2=0
r237 26 104 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4 $Y=0.085 $X2=4
+ $Y2=0
r238 26 28 17.6359 $w=3.28e-07 $l=5.05e-07 $layer=LI1_cond $X=4 $Y=0.085 $X2=4
+ $Y2=0.59
r239 22 101 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.7 $Y=0.085
+ $X2=0.7 $Y2=0
r240 22 24 13.969 $w=3.28e-07 $l=4e-07 $layer=LI1_cond $X=0.7 $Y=0.085 $X2=0.7
+ $Y2=0.485
r241 7 48 182 $w=1.7e-07 $l=8.12558e-07 $layer=licon1_NDIFF $count=1 $X=17.275
+ $Y=0.285 $X2=17.53 $Y2=0.98
r242 7 46 182 $w=1.7e-07 $l=3.19374e-07 $layer=licon1_NDIFF $count=1 $X=17.275
+ $Y=0.285 $X2=17.53 $Y2=0.43
r243 6 42 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=15.145
+ $Y=0.495 $X2=15.285 $Y2=0.705
r244 5 38 182 $w=1.7e-07 $l=3.42491e-07 $layer=licon1_NDIFF $count=1 $X=11.74
+ $Y=0.485 $X2=11.995 $Y2=0.28
r245 4 34 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=8.77
+ $Y=0.235 $X2=8.91 $Y2=0.445
r246 3 111 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=7.81
+ $Y=0.135 $X2=7.945 $Y2=0.28
r247 2 28 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=3.86
+ $Y=0.445 $X2=4 $Y2=0.59
r248 1 24 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.56
+ $Y=0.275 $X2=0.7 $Y2=0.485
.ends

.subckt PM_SKY130_FD_SC_LP__SRSDFRTN_1%noxref_30 1 2 9 11 12 13
r29 13 16 10.826 $w=3.28e-07 $l=3.1e-07 $layer=LI1_cond $X=2.915 $Y=0.34
+ $X2=2.915 $Y2=0.65
r30 11 13 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.75 $Y=0.34
+ $X2=2.915 $Y2=0.34
r31 11 12 93.2941 $w=1.68e-07 $l=1.43e-06 $layer=LI1_cond $X=2.75 $Y=0.34
+ $X2=1.32 $Y2=0.34
r32 7 12 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.195 $Y=0.425
+ $X2=1.32 $Y2=0.34
r33 7 9 12.4464 $w=2.48e-07 $l=2.7e-07 $layer=LI1_cond $X=1.195 $Y=0.425
+ $X2=1.195 $Y2=0.695
r34 2 16 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=2.775
+ $Y=0.485 $X2=2.915 $Y2=0.65
r35 1 9 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=1.1
+ $Y=0.485 $X2=1.235 $Y2=0.695
.ends

.subckt PM_SKY130_FD_SC_LP__SRSDFRTN_1%noxref_32 1 2 9 11 12 14
c35 9 0 1.55978e-19 $X=2.485 $Y=0.76
r36 14 16 6.46067 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=4.535 $Y=0.825
+ $X2=4.535 $Y2=1.01
r37 11 16 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.37 $Y=1.01
+ $X2=4.535 $Y2=1.01
r38 11 12 117.433 $w=1.68e-07 $l=1.8e-06 $layer=LI1_cond $X=4.37 $Y=1.01
+ $X2=2.57 $Y2=1.01
r39 7 12 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.485 $Y=0.925
+ $X2=2.57 $Y2=1.01
r40 7 9 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=2.485 $Y=0.925
+ $X2=2.485 $Y2=0.76
r41 2 14 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=4.395
+ $Y=0.615 $X2=4.535 $Y2=0.825
r42 1 9 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=2.345
+ $Y=0.485 $X2=2.485 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_LP__SRSDFRTN_1%A_1009_107# 1 2 11
r16 8 11 90.3583 $w=1.68e-07 $l=1.385e-06 $layer=LI1_cond $X=5.18 $Y=0.68
+ $X2=6.565 $Y2=0.68
r17 2 11 182 $w=1.7e-07 $l=3.60278e-07 $layer=licon1_NDIFF $count=1 $X=6.42
+ $Y=0.385 $X2=6.565 $Y2=0.68
r18 1 8 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=5.045
+ $Y=0.535 $X2=5.18 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_LP__SRSDFRTN_1%A_1453_77# 1 2 7 10 15
c28 15 0 1.78805e-19 $X=8.48 $Y=0.465
c29 10 0 1.3264e-19 $X=7.405 $Y=0.535
c30 7 0 3.01101e-20 $X=8.315 $Y=0.62
r31 15 17 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=8.48 $Y=0.465
+ $X2=8.48 $Y2=0.62
r32 10 12 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=7.405 $Y=0.535
+ $X2=7.405 $Y2=0.62
r33 8 12 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.57 $Y=0.62
+ $X2=7.405 $Y2=0.62
r34 7 17 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.315 $Y=0.62
+ $X2=8.48 $Y2=0.62
r35 7 8 48.6043 $w=1.68e-07 $l=7.45e-07 $layer=LI1_cond $X=8.315 $Y=0.62
+ $X2=7.57 $Y2=0.62
r36 2 15 182 $w=1.7e-07 $l=2.91719e-07 $layer=licon1_NDIFF $count=1 $X=8.34
+ $Y=0.235 $X2=8.48 $Y2=0.465
r37 1 10 182 $w=1.7e-07 $l=2.08567e-07 $layer=licon1_NDIFF $count=1 $X=7.265
+ $Y=0.385 $X2=7.405 $Y2=0.535
.ends

