* File: sky130_fd_sc_lp__decapkapwr_12.pex.spice
* Created: Wed Sep  2 09:42:20 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__DECAPKAPWR_12%VGND 1 7 9 15 18 23 28 32 36 46 47 50
+ 53
c33 23 0 8.49014e-20 $X=2.415 $Y=1.77
r34 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r35 50 51 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r36 47 54 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=5.04
+ $Y2=0
r37 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r38 44 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.26 $Y=0 $X2=5.095
+ $Y2=0
r39 44 46 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=5.26 $Y=0 $X2=5.52
+ $Y2=0
r40 43 54 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.04
+ $Y2=0
r41 42 43 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r42 40 51 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r43 39 42 219.209 $w=1.68e-07 $l=3.36e-06 $layer=LI1_cond $X=1.2 $Y=0 $X2=4.56
+ $Y2=0
r44 39 40 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r45 37 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.98 $Y=0 $X2=0.815
+ $Y2=0
r46 37 39 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=0.98 $Y=0 $X2=1.2
+ $Y2=0
r47 36 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.93 $Y=0 $X2=5.095
+ $Y2=0
r48 36 42 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=4.93 $Y=0 $X2=4.56
+ $Y2=0
r49 32 43 0.468274 $w=4.9e-07 $l=1.68e-06 $layer=MET1_cond $X=2.88 $Y=0 $X2=4.56
+ $Y2=0
r50 32 40 0.468274 $w=4.9e-07 $l=1.68e-06 $layer=MET1_cond $X=2.88 $Y=0 $X2=1.2
+ $Y2=0
r51 28 30 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=5.095 $Y=0.36
+ $X2=5.095 $Y2=1.04
r52 26 53 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.095 $Y=0.085
+ $X2=5.095 $Y2=0
r53 26 28 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=5.095 $Y=0.085
+ $X2=5.095 $Y2=0.36
r54 23 24 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=2.415
+ $Y=1.77 $X2=2.415 $Y2=1.77
r55 21 24 40.8678 $w=1.604e-06 $l=1.36e-06 $layer=POLY_cond $X=1.055 $Y=2.415
+ $X2=2.415 $Y2=2.415
r56 20 23 47.4946 $w=3.28e-07 $l=1.36e-06 $layer=LI1_cond $X=1.055 $Y=1.77
+ $X2=2.415 $Y2=1.77
r57 20 21 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=1.055
+ $Y=1.77 $X2=1.055 $Y2=1.77
r58 18 20 2.61919 $w=3.28e-07 $l=7.5e-08 $layer=LI1_cond $X=0.98 $Y=1.77
+ $X2=1.055 $Y2=1.77
r59 15 17 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=0.815 $Y=0.38
+ $X2=0.815 $Y2=1.06
r60 13 18 6.81649 $w=3.3e-07 $l=2.33345e-07 $layer=LI1_cond $X=0.815 $Y=1.605
+ $X2=0.98 $Y2=1.77
r61 13 17 19.0328 $w=3.28e-07 $l=5.45e-07 $layer=LI1_cond $X=0.815 $Y=1.605
+ $X2=0.815 $Y2=1.06
r62 12 50 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.815 $Y=0.085
+ $X2=0.815 $Y2=0
r63 12 15 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.815 $Y=0.085
+ $X2=0.815 $Y2=0.38
r64 7 24 6.40574 $w=1.604e-06 $l=2.24332e-07 $layer=POLY_cond $X=2.58 $Y=2.555
+ $X2=2.415 $Y2=2.415
r65 7 9 11.1507 $w=1.34e-06 $l=3.1e-07 $layer=POLY_cond $X=2.58 $Y=2.555
+ $X2=2.89 $Y2=2.555
r66 1 30 121.333 $w=1.7e-07 $l=8.72195e-07 $layer=licon1_NDIFF $count=1 $X=4.955
+ $Y=0.235 $X2=5.095 $Y2=1.04
r67 1 28 121.333 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=4.955
+ $Y=0.235 $X2=5.095 $Y2=0.36
r68 1 17 121.333 $w=1.7e-07 $l=8.85297e-07 $layer=licon1_NDIFF $count=1 $X=4.955
+ $Y=0.235 $X2=0.815 $Y2=1.06
r69 1 15 121.333 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=4.955
+ $Y=0.235 $X2=0.815 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_LP__DECAPKAPWR_12%KAPWR 1 9 11 13 15 22 24 26 27 30 41
c37 22 0 8.49014e-20 $X=4.79 $Y=1.51
r38 40 41 1.43077 $w=1.7e-07 $l=1.105e-06 $layer=mcon $count=6 $X=5.015 $Y=2.81
+ $X2=5.015 $Y2=2.81
r39 36 37 1.43077 $w=1.7e-07 $l=1.105e-06 $layer=mcon $count=6 $X=0.66 $Y=2.81
+ $X2=0.66 $Y2=2.81
r40 27 41 1.16689 $w=2.7e-07 $l=2.135e-06 $layer=MET1_cond $X=2.88 $Y=2.81
+ $X2=5.015 $Y2=2.81
r41 27 37 1.21335 $w=2.7e-07 $l=2.22e-06 $layer=MET1_cond $X=2.88 $Y=2.81
+ $X2=0.66 $Y2=2.81
r42 24 40 3.21187 $w=3.3e-07 $l=2e-07 $layer=LI1_cond $X=5.03 $Y=2.675 $X2=5.03
+ $Y2=2.875
r43 24 26 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=5.03 $Y=2.675
+ $X2=5.03 $Y2=2.29
r44 23 26 21.4773 $w=3.28e-07 $l=6.15e-07 $layer=LI1_cond $X=5.03 $Y=1.675
+ $X2=5.03 $Y2=2.29
r45 21 22 48.4267 $w=1.7e-07 $l=5.1e-07 $layer=licon1_POLY $count=3 $X=4.79
+ $Y=1.51 $X2=4.79 $Y2=1.51
r46 18 22 53.4994 $w=1.57e-06 $l=1.7e-06 $layer=POLY_cond $X=3.09 $Y=0.89
+ $X2=4.79 $Y2=0.89
r47 18 30 4.24848 $w=1.57e-06 $l=1.35e-07 $layer=POLY_cond $X=3.09 $Y=0.89
+ $X2=2.955 $Y2=0.89
r48 17 21 58.4822 $w=3.33e-07 $l=1.7e-06 $layer=LI1_cond $X=3.09 $Y=1.507
+ $X2=4.79 $Y2=1.507
r49 17 18 48.4267 $w=1.7e-07 $l=5.1e-07 $layer=licon1_POLY $count=3 $X=3.09
+ $Y=1.51 $X2=3.09 $Y2=1.51
r50 15 23 6.81699 $w=3.35e-07 $l=2.36525e-07 $layer=LI1_cond $X=4.865 $Y=1.507
+ $X2=5.03 $Y2=1.675
r51 15 21 2.5801 $w=3.33e-07 $l=7.5e-08 $layer=LI1_cond $X=4.865 $Y=1.507
+ $X2=4.79 $Y2=1.507
r52 14 36 3.69365 $w=2.7e-07 $l=1.94808e-07 $layer=LI1_cond $X=0.905 $Y=2.81
+ $X2=0.74 $Y2=2.875
r53 13 40 3.69365 $w=2.7e-07 $l=1.94808e-07 $layer=LI1_cond $X=4.865 $Y=2.81
+ $X2=5.03 $Y2=2.875
r54 13 14 169.025 $w=2.68e-07 $l=3.96e-06 $layer=LI1_cond $X=4.865 $Y=2.81
+ $X2=0.905 $Y2=2.81
r55 9 36 3.21187 $w=3.3e-07 $l=2e-07 $layer=LI1_cond $X=0.74 $Y=2.675 $X2=0.74
+ $Y2=2.875
r56 9 11 14.1436 $w=3.28e-07 $l=4.05e-07 $layer=LI1_cond $X=0.74 $Y=2.675
+ $X2=0.74 $Y2=2.27
r57 1 40 400 $w=1.7e-07 $l=9.42404e-07 $layer=licon1_PDIFF $count=1 $X=4.89
+ $Y=2.095 $X2=5.03 $Y2=2.97
r58 1 36 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=4.89
+ $Y=2.095 $X2=0.74 $Y2=2.95
r59 1 26 400 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_PDIFF $count=1 $X=4.89
+ $Y=2.095 $X2=5.03 $Y2=2.29
r60 1 11 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=4.89
+ $Y=2.095 $X2=0.74 $Y2=2.27
.ends

.subckt PM_SKY130_FD_SC_LP__DECAPKAPWR_12%VPWR 1 8 14
r14 5 14 0.00264757 $w=5.76e-06 $l=1.22e-07 $layer=MET1_cond $X=2.88 $Y=3.33
+ $X2=2.88 $Y2=3.208
r15 5 8 1.55 $w=1.7e-07 $l=1.02e-06 $layer=mcon $count=6 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r16 4 8 344.471 $w=1.68e-07 $l=5.28e-06 $layer=LI1_cond $X=0.24 $Y=3.33 $X2=5.52
+ $Y2=3.33
r17 4 5 1.55 $w=1.7e-07 $l=1.02e-06 $layer=mcon $count=6 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r18 1 14 2.17014e-05 $w=5.76e-06 $l=1e-09 $layer=MET1_cond $X=2.88 $Y=3.207
+ $X2=2.88 $Y2=3.208
.ends

