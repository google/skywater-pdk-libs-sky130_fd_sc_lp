* File: sky130_fd_sc_lp__and4bb_4.pxi.spice
* Created: Fri Aug 28 10:09:28 2020
* 
x_PM_SKY130_FD_SC_LP__AND4BB_4%B_N N_B_N_M1001_g N_B_N_M1012_g B_N B_N B_N B_N
+ B_N N_B_N_c_110_n N_B_N_c_111_n PM_SKY130_FD_SC_LP__AND4BB_4%B_N
x_PM_SKY130_FD_SC_LP__AND4BB_4%A_254_21# N_A_254_21#_M1019_d N_A_254_21#_M1011_d
+ N_A_254_21#_M1008_d N_A_254_21#_M1006_g N_A_254_21#_M1004_g
+ N_A_254_21#_M1007_g N_A_254_21#_M1009_g N_A_254_21#_M1013_g
+ N_A_254_21#_M1014_g N_A_254_21#_M1015_g N_A_254_21#_M1017_g
+ N_A_254_21#_c_234_p N_A_254_21#_c_143_n N_A_254_21#_c_144_n
+ N_A_254_21#_c_152_n N_A_254_21#_c_253_p N_A_254_21#_c_194_p
+ N_A_254_21#_c_161_p N_A_254_21#_c_145_n N_A_254_21#_c_146_n
+ N_A_254_21#_c_165_p N_A_254_21#_c_166_p PM_SKY130_FD_SC_LP__AND4BB_4%A_254_21#
x_PM_SKY130_FD_SC_LP__AND4BB_4%D N_D_M1011_g N_D_M1003_g D D N_D_c_284_n
+ PM_SKY130_FD_SC_LP__AND4BB_4%D
x_PM_SKY130_FD_SC_LP__AND4BB_4%C N_C_M1005_g N_C_M1000_g C C N_C_c_327_n
+ PM_SKY130_FD_SC_LP__AND4BB_4%C
x_PM_SKY130_FD_SC_LP__AND4BB_4%A_49_131# N_A_49_131#_M1001_s N_A_49_131#_M1012_s
+ N_A_49_131#_M1010_g N_A_49_131#_M1008_g N_A_49_131#_c_358_n
+ N_A_49_131#_c_364_n N_A_49_131#_c_365_n N_A_49_131#_c_359_n
+ N_A_49_131#_c_367_n N_A_49_131#_c_360_n N_A_49_131#_c_361_n
+ PM_SKY130_FD_SC_LP__AND4BB_4%A_49_131#
x_PM_SKY130_FD_SC_LP__AND4BB_4%A_929_21# N_A_929_21#_M1016_d N_A_929_21#_M1002_d
+ N_A_929_21#_M1019_g N_A_929_21#_M1018_g N_A_929_21#_c_447_n
+ N_A_929_21#_c_448_n N_A_929_21#_c_449_n N_A_929_21#_c_450_n
+ N_A_929_21#_c_451_n N_A_929_21#_c_452_n N_A_929_21#_c_456_n
+ N_A_929_21#_c_453_n N_A_929_21#_c_454_n PM_SKY130_FD_SC_LP__AND4BB_4%A_929_21#
x_PM_SKY130_FD_SC_LP__AND4BB_4%A_N N_A_N_M1002_g N_A_N_c_500_n N_A_N_c_501_n
+ N_A_N_M1016_g A_N N_A_N_c_503_n N_A_N_c_504_n PM_SKY130_FD_SC_LP__AND4BB_4%A_N
x_PM_SKY130_FD_SC_LP__AND4BB_4%VPWR N_VPWR_M1012_d N_VPWR_M1009_s N_VPWR_M1017_s
+ N_VPWR_M1000_d N_VPWR_M1018_d N_VPWR_c_531_n N_VPWR_c_532_n N_VPWR_c_533_n
+ N_VPWR_c_534_n N_VPWR_c_535_n N_VPWR_c_536_n N_VPWR_c_537_n N_VPWR_c_538_n
+ N_VPWR_c_539_n N_VPWR_c_540_n N_VPWR_c_541_n VPWR N_VPWR_c_542_n
+ N_VPWR_c_543_n N_VPWR_c_544_n N_VPWR_c_530_n N_VPWR_c_546_n N_VPWR_c_547_n
+ PM_SKY130_FD_SC_LP__AND4BB_4%VPWR
x_PM_SKY130_FD_SC_LP__AND4BB_4%X N_X_M1006_d N_X_M1013_d N_X_M1004_d N_X_M1014_d
+ N_X_c_612_n N_X_c_610_n N_X_c_606_n N_X_c_607_n N_X_c_608_n N_X_c_654_p X
+ PM_SKY130_FD_SC_LP__AND4BB_4%X
x_PM_SKY130_FD_SC_LP__AND4BB_4%VGND N_VGND_M1001_d N_VGND_M1007_s N_VGND_M1015_s
+ N_VGND_M1016_s N_VGND_c_659_n N_VGND_c_660_n N_VGND_c_661_n N_VGND_c_662_n
+ N_VGND_c_663_n N_VGND_c_664_n N_VGND_c_665_n N_VGND_c_666_n N_VGND_c_667_n
+ N_VGND_c_668_n VGND N_VGND_c_669_n N_VGND_c_670_n N_VGND_c_671_n
+ N_VGND_c_672_n PM_SKY130_FD_SC_LP__AND4BB_4%VGND
cc_1 VNB N_B_N_M1012_g 0.00825229f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=2.045
cc_2 VNB B_N 0.00759708f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.47
cc_3 VNB N_B_N_c_110_n 0.0408476f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.35
cc_4 VNB N_B_N_c_111_n 0.0220629f $X=-0.19 $Y=-0.245 $X2=0.707 $Y2=1.185
cc_5 VNB N_A_254_21#_M1006_g 0.0261781f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.95
cc_6 VNB N_A_254_21#_M1007_g 0.022171f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.35
cc_7 VNB N_A_254_21#_M1013_g 0.0221884f $X=-0.19 $Y=-0.245 $X2=0.74 $Y2=1.295
cc_8 VNB N_A_254_21#_M1015_g 0.024738f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_254_21#_c_143_n 0.0723734f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_254_21#_c_144_n 0.002754f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_254_21#_c_145_n 0.00815024f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_254_21#_c_146_n 0.00147516f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_D_M1011_g 0.00503888f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=0.865
cc_14 VNB N_D_M1003_g 0.0190863f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB D 0.00303518f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.84
cc_16 VNB N_D_c_284_n 0.0333657f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_C_M1005_g 0.0183128f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=0.865
cc_18 VNB N_C_M1000_g 0.00530854f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB C 0.00868354f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.84
cc_20 VNB N_C_c_327_n 0.0285648f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_49_131#_M1010_g 0.0275273f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.84
cc_22 VNB N_A_49_131#_c_358_n 0.0440301f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_49_131#_c_359_n 0.00825357f $X=-0.19 $Y=-0.245 $X2=0.74 $Y2=0.555
cc_24 VNB N_A_49_131#_c_360_n 0.00484635f $X=-0.19 $Y=-0.245 $X2=0.74 $Y2=1.295
cc_25 VNB N_A_49_131#_c_361_n 0.0250565f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_929_21#_M1018_g 0.00725809f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.95
cc_27 VNB N_A_929_21#_c_447_n 0.0195478f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_929_21#_c_448_n 0.0151413f $X=-0.19 $Y=-0.245 $X2=0.707 $Y2=1.35
cc_29 VNB N_A_929_21#_c_449_n 0.0149219f $X=-0.19 $Y=-0.245 $X2=0.707 $Y2=1.515
cc_30 VNB N_A_929_21#_c_450_n 3.11212e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_929_21#_c_451_n 0.0378507f $X=-0.19 $Y=-0.245 $X2=0.74 $Y2=1.295
cc_32 VNB N_A_929_21#_c_452_n 0.00410449f $X=-0.19 $Y=-0.245 $X2=0.74 $Y2=1.665
cc_33 VNB N_A_929_21#_c_453_n 0.00532032f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_929_21#_c_454_n 0.0212214f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_N_c_500_n 0.0139752f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=2.045
cc_36 VNB N_A_N_c_501_n 0.00941881f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=2.045
cc_37 VNB N_A_N_M1016_g 0.0387045f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=0.84
cc_38 VNB N_A_N_c_503_n 0.0311873f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_N_c_504_n 0.0100269f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_VPWR_c_530_n 0.263193f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_X_c_606_n 3.90791e-19 $X=-0.19 $Y=-0.245 $X2=0.707 $Y2=1.185
cc_42 VNB N_X_c_607_n 0.011344f $X=-0.19 $Y=-0.245 $X2=0.74 $Y2=0.555
cc_43 VNB N_X_c_608_n 0.0060857f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB X 0.00348055f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_659_n 0.0044254f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_660_n 3.3315e-19 $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.35
cc_47 VNB N_VGND_c_661_n 0.00507173f $X=-0.19 $Y=-0.245 $X2=0.74 $Y2=0.555
cc_48 VNB N_VGND_c_662_n 0.0252905f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_663_n 0.0323839f $X=-0.19 $Y=-0.245 $X2=0.74 $Y2=1.665
cc_50 VNB N_VGND_c_664_n 0.00442399f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_665_n 0.0148832f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_666_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_667_n 0.0173279f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_668_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_669_n 0.0561623f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_VGND_c_670_n 0.0178307f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_VGND_c_671_n 0.34783f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_672_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VPB N_B_N_M1012_g 0.0230383f $X=-0.19 $Y=1.655 $X2=0.605 $Y2=2.045
cc_60 VPB B_N 0.00142959f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=0.47
cc_61 VPB N_A_254_21#_M1004_g 0.0216624f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_62 VPB N_A_254_21#_M1009_g 0.018828f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_63 VPB N_A_254_21#_M1014_g 0.0188453f $X=-0.19 $Y=1.655 $X2=0.74 $Y2=2.035
cc_64 VPB N_A_254_21#_M1017_g 0.0200811f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_65 VPB N_A_254_21#_c_143_n 0.0121814f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_66 VPB N_A_254_21#_c_152_n 0.00132466f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_67 VPB N_D_M1011_g 0.0204083f $X=-0.19 $Y=1.655 $X2=0.605 $Y2=0.865
cc_68 VPB D 0.00299314f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=0.84
cc_69 VPB N_C_M1000_g 0.0201853f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_70 VPB C 0.00428197f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=0.84
cc_71 VPB N_A_49_131#_M1008_g 0.0209616f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_72 VPB N_A_49_131#_c_358_n 0.038393f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_73 VPB N_A_49_131#_c_364_n 0.022079f $X=-0.19 $Y=1.655 $X2=0.707 $Y2=1.185
cc_74 VPB N_A_49_131#_c_365_n 0.0124852f $X=-0.19 $Y=1.655 $X2=0.707 $Y2=1.515
cc_75 VPB N_A_49_131#_c_359_n 0.00407392f $X=-0.19 $Y=1.655 $X2=0.74 $Y2=0.555
cc_76 VPB N_A_49_131#_c_367_n 4.0033e-19 $X=-0.19 $Y=1.655 $X2=0.74 $Y2=0.925
cc_77 VPB N_A_49_131#_c_360_n 0.0020497f $X=-0.19 $Y=1.655 $X2=0.74 $Y2=1.295
cc_78 VPB N_A_49_131#_c_361_n 0.00651302f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_79 VPB N_A_929_21#_M1018_g 0.0222177f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.95
cc_80 VPB N_A_929_21#_c_456_n 0.0248056f $X=-0.19 $Y=1.655 $X2=0.74 $Y2=2.035
cc_81 VPB N_A_929_21#_c_453_n 0.0045803f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_82 VPB N_A_N_M1002_g 0.0287918f $X=-0.19 $Y=1.655 $X2=0.605 $Y2=0.865
cc_83 VPB N_A_N_c_500_n 0.0111873f $X=-0.19 $Y=1.655 $X2=0.605 $Y2=2.045
cc_84 VPB N_A_N_c_501_n 7.92945e-19 $X=-0.19 $Y=1.655 $X2=0.605 $Y2=2.045
cc_85 VPB N_A_N_c_503_n 0.0106695f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_86 VPB N_A_N_c_504_n 0.0213874f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_87 VPB N_VPWR_c_531_n 0.0137165f $X=-0.19 $Y=1.655 $X2=0.707 $Y2=1.35
cc_88 VPB N_VPWR_c_532_n 3.22457e-19 $X=-0.19 $Y=1.655 $X2=0.707 $Y2=1.515
cc_89 VPB N_VPWR_c_533_n 0.00447432f $X=-0.19 $Y=1.655 $X2=0.74 $Y2=0.925
cc_90 VPB N_VPWR_c_534_n 0.00507026f $X=-0.19 $Y=1.655 $X2=0.74 $Y2=1.665
cc_91 VPB N_VPWR_c_535_n 0.0150054f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_92 VPB N_VPWR_c_536_n 0.0125849f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_93 VPB N_VPWR_c_537_n 0.00436447f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_94 VPB N_VPWR_c_538_n 0.0158557f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_95 VPB N_VPWR_c_539_n 0.00631736f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_96 VPB N_VPWR_c_540_n 0.0181535f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_97 VPB N_VPWR_c_541_n 0.00631736f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_98 VPB N_VPWR_c_542_n 0.0297794f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_99 VPB N_VPWR_c_543_n 0.0180581f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_100 VPB N_VPWR_c_544_n 0.0384204f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_101 VPB N_VPWR_c_530_n 0.101348f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_102 VPB N_VPWR_c_546_n 0.0051042f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_103 VPB N_VPWR_c_547_n 0.0051042f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_104 VPB N_X_c_610_n 0.00663963f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_105 VPB X 0.00127125f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_106 B_N N_A_254_21#_M1006_g 0.002632f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_107 N_B_N_c_110_n N_A_254_21#_M1006_g 0.00927041f $X=0.72 $Y=1.35 $X2=0 $Y2=0
cc_108 N_B_N_c_111_n N_A_254_21#_M1006_g 0.00635095f $X=0.707 $Y=1.185 $X2=0
+ $Y2=0
cc_109 N_B_N_M1012_g N_A_254_21#_c_143_n 0.0149882f $X=0.605 $Y=2.045 $X2=0
+ $Y2=0
cc_110 B_N N_A_254_21#_c_143_n 0.00183793f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_111 B_N N_A_49_131#_c_358_n 0.106054f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_112 N_B_N_c_111_n N_A_49_131#_c_358_n 0.0282332f $X=0.707 $Y=1.185 $X2=0
+ $Y2=0
cc_113 N_B_N_M1012_g N_A_49_131#_c_364_n 0.00612833f $X=0.605 $Y=2.045 $X2=0
+ $Y2=0
cc_114 B_N N_A_49_131#_c_364_n 0.00971448f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_115 B_N N_VPWR_M1012_d 0.00496333f $X=0.635 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_116 N_B_N_M1012_g N_X_c_612_n 0.00133977f $X=0.605 $Y=2.045 $X2=0 $Y2=0
cc_117 B_N N_X_c_612_n 0.0185626f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_118 B_N N_X_c_608_n 0.0105216f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_119 N_B_N_c_110_n N_X_c_608_n 5.19588e-19 $X=0.72 $Y=1.35 $X2=0 $Y2=0
cc_120 N_B_N_c_111_n N_X_c_608_n 3.87434e-19 $X=0.707 $Y=1.185 $X2=0 $Y2=0
cc_121 N_B_N_M1012_g X 8.40695e-19 $X=0.605 $Y=2.045 $X2=0 $Y2=0
cc_122 B_N X 0.0316952f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_123 N_B_N_c_110_n X 0.00208168f $X=0.72 $Y=1.35 $X2=0 $Y2=0
cc_124 B_N N_VGND_M1001_d 0.00499564f $X=0.635 $Y=0.47 $X2=-0.19 $Y2=-0.245
cc_125 B_N N_VGND_c_659_n 0.0333217f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_126 N_B_N_c_111_n N_VGND_c_659_n 0.00102892f $X=0.707 $Y=1.185 $X2=0 $Y2=0
cc_127 B_N N_VGND_c_663_n 0.00683597f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_128 N_B_N_c_111_n N_VGND_c_663_n 0.00279135f $X=0.707 $Y=1.185 $X2=0 $Y2=0
cc_129 B_N N_VGND_c_671_n 0.00778882f $X=0.635 $Y=0.47 $X2=0 $Y2=0
cc_130 N_B_N_c_111_n N_VGND_c_671_n 0.00295181f $X=0.707 $Y=1.185 $X2=0 $Y2=0
cc_131 N_A_254_21#_M1017_g N_D_M1011_g 0.0412621f $X=2.635 $Y=2.465 $X2=0 $Y2=0
cc_132 N_A_254_21#_c_143_n N_D_M1011_g 0.00475386f $X=2.65 $Y=1.5 $X2=0 $Y2=0
cc_133 N_A_254_21#_c_152_n N_D_M1011_g 0.00368626f $X=2.77 $Y=1.965 $X2=0 $Y2=0
cc_134 N_A_254_21#_c_161_p N_D_M1011_g 0.0140176f $X=4.45 $Y=2.13 $X2=0 $Y2=0
cc_135 N_A_254_21#_c_146_n N_D_M1011_g 3.49556e-19 $X=2.77 $Y=1.53 $X2=0 $Y2=0
cc_136 N_A_254_21#_M1015_g N_D_M1003_g 0.0210974f $X=2.635 $Y=0.655 $X2=0 $Y2=0
cc_137 N_A_254_21#_c_144_n N_D_M1003_g 0.00308442f $X=2.77 $Y=1.415 $X2=0 $Y2=0
cc_138 N_A_254_21#_c_165_p N_D_M1003_g 0.0167879f $X=3.46 $Y=0.647 $X2=0 $Y2=0
cc_139 N_A_254_21#_c_166_p N_D_M1003_g 0.00909081f $X=4.405 $Y=0.647 $X2=0 $Y2=0
cc_140 N_A_254_21#_M1017_g D 3.5579e-19 $X=2.635 $Y=2.465 $X2=0 $Y2=0
cc_141 N_A_254_21#_c_143_n D 6.38219e-19 $X=2.65 $Y=1.5 $X2=0 $Y2=0
cc_142 N_A_254_21#_c_144_n D 0.0145189f $X=2.77 $Y=1.415 $X2=0 $Y2=0
cc_143 N_A_254_21#_c_152_n D 0.0112217f $X=2.77 $Y=1.965 $X2=0 $Y2=0
cc_144 N_A_254_21#_c_161_p D 0.0190947f $X=4.45 $Y=2.13 $X2=0 $Y2=0
cc_145 N_A_254_21#_c_146_n D 0.0187757f $X=2.77 $Y=1.53 $X2=0 $Y2=0
cc_146 N_A_254_21#_c_165_p D 0.0188661f $X=3.46 $Y=0.647 $X2=0 $Y2=0
cc_147 N_A_254_21#_M1015_g N_D_c_284_n 0.00454838f $X=2.635 $Y=0.655 $X2=0 $Y2=0
cc_148 N_A_254_21#_c_143_n N_D_c_284_n 0.0128694f $X=2.65 $Y=1.5 $X2=0 $Y2=0
cc_149 N_A_254_21#_c_144_n N_D_c_284_n 0.00127291f $X=2.77 $Y=1.415 $X2=0 $Y2=0
cc_150 N_A_254_21#_c_161_p N_D_c_284_n 0.00171426f $X=4.45 $Y=2.13 $X2=0 $Y2=0
cc_151 N_A_254_21#_c_146_n N_D_c_284_n 7.87297e-19 $X=2.77 $Y=1.53 $X2=0 $Y2=0
cc_152 N_A_254_21#_c_165_p N_D_c_284_n 0.00147363f $X=3.46 $Y=0.647 $X2=0 $Y2=0
cc_153 N_A_254_21#_c_166_p N_C_M1005_g 0.0305696f $X=4.405 $Y=0.647 $X2=0 $Y2=0
cc_154 N_A_254_21#_c_161_p N_C_M1000_g 0.0137588f $X=4.45 $Y=2.13 $X2=0 $Y2=0
cc_155 N_A_254_21#_c_161_p C 0.0295413f $X=4.45 $Y=2.13 $X2=0 $Y2=0
cc_156 N_A_254_21#_c_166_p C 0.0308072f $X=4.405 $Y=0.647 $X2=0 $Y2=0
cc_157 N_A_254_21#_c_161_p N_C_c_327_n 6.69329e-19 $X=4.45 $Y=2.13 $X2=0 $Y2=0
cc_158 N_A_254_21#_c_166_p N_C_c_327_n 0.0012502f $X=4.405 $Y=0.647 $X2=0 $Y2=0
cc_159 N_A_254_21#_c_166_p N_A_49_131#_M1010_g 0.0381628f $X=4.405 $Y=0.647
+ $X2=0 $Y2=0
cc_160 N_A_254_21#_c_161_p N_A_49_131#_M1008_g 0.0137616f $X=4.45 $Y=2.13 $X2=0
+ $Y2=0
cc_161 N_A_254_21#_M1011_d N_A_49_131#_c_364_n 0.00483346f $X=3.285 $Y=1.835
+ $X2=0 $Y2=0
cc_162 N_A_254_21#_M1008_d N_A_49_131#_c_364_n 0.00833193f $X=4.255 $Y=1.835
+ $X2=0 $Y2=0
cc_163 N_A_254_21#_M1004_g N_A_49_131#_c_364_n 0.0151707f $X=1.345 $Y=2.465
+ $X2=0 $Y2=0
cc_164 N_A_254_21#_M1009_g N_A_49_131#_c_364_n 0.0130289f $X=1.775 $Y=2.465
+ $X2=0 $Y2=0
cc_165 N_A_254_21#_M1014_g N_A_49_131#_c_364_n 0.0130289f $X=2.205 $Y=2.465
+ $X2=0 $Y2=0
cc_166 N_A_254_21#_M1017_g N_A_49_131#_c_364_n 0.0170093f $X=2.635 $Y=2.465
+ $X2=0 $Y2=0
cc_167 N_A_254_21#_c_194_p N_A_49_131#_c_364_n 0.0090121f $X=2.855 $Y=2.13 $X2=0
+ $Y2=0
cc_168 N_A_254_21#_c_161_p N_A_49_131#_c_364_n 0.104253f $X=4.45 $Y=2.13 $X2=0
+ $Y2=0
cc_169 N_A_254_21#_c_161_p N_A_49_131#_c_359_n 0.0114635f $X=4.45 $Y=2.13 $X2=0
+ $Y2=0
cc_170 N_A_254_21#_c_161_p N_A_49_131#_c_360_n 0.023963f $X=4.45 $Y=2.13 $X2=0
+ $Y2=0
cc_171 N_A_254_21#_c_145_n N_A_49_131#_c_360_n 0.00158702f $X=4.935 $Y=0.42
+ $X2=0 $Y2=0
cc_172 N_A_254_21#_c_166_p N_A_49_131#_c_360_n 0.0140048f $X=4.405 $Y=0.647
+ $X2=0 $Y2=0
cc_173 N_A_254_21#_c_161_p N_A_49_131#_c_361_n 8.86683e-19 $X=4.45 $Y=2.13 $X2=0
+ $Y2=0
cc_174 N_A_254_21#_c_166_p N_A_49_131#_c_361_n 8.75751e-19 $X=4.405 $Y=0.647
+ $X2=0 $Y2=0
cc_175 N_A_254_21#_c_145_n N_A_929_21#_c_447_n 0.0103224f $X=4.935 $Y=0.42 $X2=0
+ $Y2=0
cc_176 N_A_254_21#_M1019_d N_A_929_21#_c_450_n 0.0019492f $X=4.795 $Y=0.235
+ $X2=0 $Y2=0
cc_177 N_A_254_21#_c_145_n N_A_929_21#_c_450_n 0.0246871f $X=4.935 $Y=0.42 $X2=0
+ $Y2=0
cc_178 N_A_254_21#_c_145_n N_A_929_21#_c_451_n 9.29503e-19 $X=4.935 $Y=0.42
+ $X2=0 $Y2=0
cc_179 N_A_254_21#_c_145_n N_A_929_21#_c_454_n 0.0222615f $X=4.935 $Y=0.42 $X2=0
+ $Y2=0
cc_180 N_A_254_21#_c_166_p N_A_929_21#_c_454_n 0.00353208f $X=4.405 $Y=0.647
+ $X2=0 $Y2=0
cc_181 N_A_254_21#_c_145_n N_A_N_M1016_g 0.00115735f $X=4.935 $Y=0.42 $X2=0
+ $Y2=0
cc_182 N_A_254_21#_c_152_n N_VPWR_M1017_s 0.00163015f $X=2.77 $Y=1.965 $X2=0
+ $Y2=0
cc_183 N_A_254_21#_c_194_p N_VPWR_M1017_s 9.65132e-19 $X=2.855 $Y=2.13 $X2=0
+ $Y2=0
cc_184 N_A_254_21#_c_161_p N_VPWR_M1017_s 0.0111473f $X=4.45 $Y=2.13 $X2=0 $Y2=0
cc_185 N_A_254_21#_c_161_p N_VPWR_M1000_d 0.0108754f $X=4.45 $Y=2.13 $X2=0 $Y2=0
cc_186 N_A_254_21#_M1004_g N_VPWR_c_531_n 0.00991439f $X=1.345 $Y=2.465 $X2=0
+ $Y2=0
cc_187 N_A_254_21#_M1009_g N_VPWR_c_531_n 0.00125151f $X=1.775 $Y=2.465 $X2=0
+ $Y2=0
cc_188 N_A_254_21#_M1004_g N_VPWR_c_532_n 0.00125151f $X=1.345 $Y=2.465 $X2=0
+ $Y2=0
cc_189 N_A_254_21#_M1009_g N_VPWR_c_532_n 0.00885091f $X=1.775 $Y=2.465 $X2=0
+ $Y2=0
cc_190 N_A_254_21#_M1014_g N_VPWR_c_532_n 0.00935543f $X=2.205 $Y=2.465 $X2=0
+ $Y2=0
cc_191 N_A_254_21#_M1017_g N_VPWR_c_532_n 0.00130861f $X=2.635 $Y=2.465 $X2=0
+ $Y2=0
cc_192 N_A_254_21#_M1017_g N_VPWR_c_533_n 0.00336811f $X=2.635 $Y=2.465 $X2=0
+ $Y2=0
cc_193 N_A_254_21#_M1004_g N_VPWR_c_536_n 0.00359504f $X=1.345 $Y=2.465 $X2=0
+ $Y2=0
cc_194 N_A_254_21#_M1009_g N_VPWR_c_536_n 0.00359504f $X=1.775 $Y=2.465 $X2=0
+ $Y2=0
cc_195 N_A_254_21#_M1014_g N_VPWR_c_538_n 0.00359504f $X=2.205 $Y=2.465 $X2=0
+ $Y2=0
cc_196 N_A_254_21#_M1017_g N_VPWR_c_538_n 0.00432313f $X=2.635 $Y=2.465 $X2=0
+ $Y2=0
cc_197 N_A_254_21#_M1011_d N_VPWR_c_530_n 0.00346035f $X=3.285 $Y=1.835 $X2=0
+ $Y2=0
cc_198 N_A_254_21#_M1008_d N_VPWR_c_530_n 0.00482985f $X=4.255 $Y=1.835 $X2=0
+ $Y2=0
cc_199 N_A_254_21#_M1004_g N_VPWR_c_530_n 0.00429447f $X=1.345 $Y=2.465 $X2=0
+ $Y2=0
cc_200 N_A_254_21#_M1009_g N_VPWR_c_530_n 0.00429447f $X=1.775 $Y=2.465 $X2=0
+ $Y2=0
cc_201 N_A_254_21#_M1014_g N_VPWR_c_530_n 0.00429447f $X=2.205 $Y=2.465 $X2=0
+ $Y2=0
cc_202 N_A_254_21#_M1017_g N_VPWR_c_530_n 0.0063872f $X=2.635 $Y=2.465 $X2=0
+ $Y2=0
cc_203 N_A_254_21#_M1004_g N_X_c_612_n 0.00552872f $X=1.345 $Y=2.465 $X2=0 $Y2=0
cc_204 N_A_254_21#_M1004_g N_X_c_610_n 0.00967522f $X=1.345 $Y=2.465 $X2=0 $Y2=0
cc_205 N_A_254_21#_M1009_g N_X_c_610_n 0.0137166f $X=1.775 $Y=2.465 $X2=0 $Y2=0
cc_206 N_A_254_21#_M1014_g N_X_c_610_n 0.0137609f $X=2.205 $Y=2.465 $X2=0 $Y2=0
cc_207 N_A_254_21#_c_234_p N_X_c_610_n 0.0789829f $X=2.685 $Y=1.53 $X2=0 $Y2=0
cc_208 N_A_254_21#_c_143_n N_X_c_610_n 0.00699881f $X=2.65 $Y=1.5 $X2=0 $Y2=0
cc_209 N_A_254_21#_c_152_n N_X_c_610_n 0.00561822f $X=2.77 $Y=1.965 $X2=0 $Y2=0
cc_210 N_A_254_21#_M1007_g N_X_c_607_n 0.0142467f $X=1.775 $Y=0.655 $X2=0 $Y2=0
cc_211 N_A_254_21#_M1013_g N_X_c_607_n 0.0138902f $X=2.205 $Y=0.655 $X2=0 $Y2=0
cc_212 N_A_254_21#_M1015_g N_X_c_607_n 0.00139835f $X=2.635 $Y=0.655 $X2=0 $Y2=0
cc_213 N_A_254_21#_c_234_p N_X_c_607_n 0.0156385f $X=2.685 $Y=1.53 $X2=0 $Y2=0
cc_214 N_A_254_21#_c_143_n N_X_c_607_n 0.00503231f $X=2.65 $Y=1.5 $X2=0 $Y2=0
cc_215 N_A_254_21#_c_144_n N_X_c_607_n 0.0136674f $X=2.77 $Y=1.415 $X2=0 $Y2=0
cc_216 N_A_254_21#_M1006_g N_X_c_608_n 0.0163115f $X=1.345 $Y=0.655 $X2=0 $Y2=0
cc_217 N_A_254_21#_c_234_p N_X_c_608_n 0.0617032f $X=2.685 $Y=1.53 $X2=0 $Y2=0
cc_218 N_A_254_21#_c_143_n N_X_c_608_n 0.00246472f $X=2.65 $Y=1.5 $X2=0 $Y2=0
cc_219 N_A_254_21#_M1006_g X 0.00247746f $X=1.345 $Y=0.655 $X2=0 $Y2=0
cc_220 N_A_254_21#_M1004_g X 0.00446177f $X=1.345 $Y=2.465 $X2=0 $Y2=0
cc_221 N_A_254_21#_M1007_g X 4.37715e-19 $X=1.775 $Y=0.655 $X2=0 $Y2=0
cc_222 N_A_254_21#_M1009_g X 7.30045e-19 $X=1.775 $Y=2.465 $X2=0 $Y2=0
cc_223 N_A_254_21#_c_234_p X 0.0174366f $X=2.685 $Y=1.53 $X2=0 $Y2=0
cc_224 N_A_254_21#_c_143_n X 0.0120896f $X=2.65 $Y=1.5 $X2=0 $Y2=0
cc_225 N_A_254_21#_c_144_n N_VGND_M1015_s 4.57336e-19 $X=2.77 $Y=1.415 $X2=0
+ $Y2=0
cc_226 N_A_254_21#_c_253_p N_VGND_M1015_s 0.00179089f $X=2.855 $Y=0.955 $X2=0
+ $Y2=0
cc_227 N_A_254_21#_c_165_p N_VGND_M1015_s 0.0126015f $X=3.46 $Y=0.647 $X2=0
+ $Y2=0
cc_228 N_A_254_21#_M1006_g N_VGND_c_659_n 0.00332889f $X=1.345 $Y=0.655 $X2=0
+ $Y2=0
cc_229 N_A_254_21#_M1006_g N_VGND_c_660_n 6.50036e-19 $X=1.345 $Y=0.655 $X2=0
+ $Y2=0
cc_230 N_A_254_21#_M1007_g N_VGND_c_660_n 0.0114577f $X=1.775 $Y=0.655 $X2=0
+ $Y2=0
cc_231 N_A_254_21#_M1013_g N_VGND_c_660_n 0.0115986f $X=2.205 $Y=0.655 $X2=0
+ $Y2=0
cc_232 N_A_254_21#_M1015_g N_VGND_c_660_n 6.75532e-19 $X=2.635 $Y=0.655 $X2=0
+ $Y2=0
cc_233 N_A_254_21#_M1015_g N_VGND_c_661_n 0.0069408f $X=2.635 $Y=0.655 $X2=0
+ $Y2=0
cc_234 N_A_254_21#_c_253_p N_VGND_c_661_n 0.00577035f $X=2.855 $Y=0.955 $X2=0
+ $Y2=0
cc_235 N_A_254_21#_c_165_p N_VGND_c_661_n 0.0214422f $X=3.46 $Y=0.647 $X2=0
+ $Y2=0
cc_236 N_A_254_21#_c_166_p N_VGND_c_661_n 0.0226458f $X=4.405 $Y=0.647 $X2=0
+ $Y2=0
cc_237 N_A_254_21#_c_145_n N_VGND_c_662_n 0.0399752f $X=4.935 $Y=0.42 $X2=0
+ $Y2=0
cc_238 N_A_254_21#_M1006_g N_VGND_c_665_n 0.00585385f $X=1.345 $Y=0.655 $X2=0
+ $Y2=0
cc_239 N_A_254_21#_M1007_g N_VGND_c_665_n 0.00486043f $X=1.775 $Y=0.655 $X2=0
+ $Y2=0
cc_240 N_A_254_21#_M1013_g N_VGND_c_667_n 0.00486043f $X=2.205 $Y=0.655 $X2=0
+ $Y2=0
cc_241 N_A_254_21#_M1015_g N_VGND_c_667_n 0.00585385f $X=2.635 $Y=0.655 $X2=0
+ $Y2=0
cc_242 N_A_254_21#_c_166_p N_VGND_c_669_n 0.101631f $X=4.405 $Y=0.647 $X2=0
+ $Y2=0
cc_243 N_A_254_21#_M1019_d N_VGND_c_671_n 0.00215176f $X=4.795 $Y=0.235 $X2=0
+ $Y2=0
cc_244 N_A_254_21#_M1006_g N_VGND_c_671_n 0.0118358f $X=1.345 $Y=0.655 $X2=0
+ $Y2=0
cc_245 N_A_254_21#_M1007_g N_VGND_c_671_n 0.00824727f $X=1.775 $Y=0.655 $X2=0
+ $Y2=0
cc_246 N_A_254_21#_M1013_g N_VGND_c_671_n 0.00824727f $X=2.205 $Y=0.655 $X2=0
+ $Y2=0
cc_247 N_A_254_21#_M1015_g N_VGND_c_671_n 0.0113138f $X=2.635 $Y=0.655 $X2=0
+ $Y2=0
cc_248 N_A_254_21#_c_166_p N_VGND_c_671_n 0.0615566f $X=4.405 $Y=0.647 $X2=0
+ $Y2=0
cc_249 N_A_254_21#_c_165_p A_671_47# 0.00358662f $X=3.46 $Y=0.647 $X2=-0.19
+ $Y2=-0.245
cc_250 N_A_254_21#_c_166_p A_671_47# 0.00902033f $X=4.405 $Y=0.647 $X2=-0.19
+ $Y2=-0.245
cc_251 N_A_254_21#_c_166_p A_743_47# 0.0117834f $X=4.405 $Y=0.647 $X2=-0.19
+ $Y2=-0.245
cc_252 N_A_254_21#_c_145_n A_851_47# 0.00989928f $X=4.935 $Y=0.42 $X2=-0.19
+ $Y2=-0.245
cc_253 N_A_254_21#_c_166_p A_851_47# 0.00393552f $X=4.405 $Y=0.647 $X2=-0.19
+ $Y2=-0.245
cc_254 N_D_M1003_g N_C_M1005_g 0.0444145f $X=3.28 $Y=0.655 $X2=0 $Y2=0
cc_255 N_D_M1011_g N_C_M1000_g 0.0606683f $X=3.21 $Y=2.465 $X2=0 $Y2=0
cc_256 D N_C_M1000_g 7.98648e-19 $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_257 N_D_M1011_g C 8.63014e-19 $X=3.21 $Y=2.465 $X2=0 $Y2=0
cc_258 D C 0.0471975f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_259 N_D_c_284_n C 0.00208795f $X=3.19 $Y=1.375 $X2=0 $Y2=0
cc_260 D N_C_c_327_n 3.24284e-19 $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_261 N_D_c_284_n N_C_c_327_n 0.0444145f $X=3.19 $Y=1.375 $X2=0 $Y2=0
cc_262 N_D_M1011_g N_A_49_131#_c_364_n 0.0131245f $X=3.21 $Y=2.465 $X2=0 $Y2=0
cc_263 N_D_M1011_g N_VPWR_c_533_n 0.00354544f $X=3.21 $Y=2.465 $X2=0 $Y2=0
cc_264 N_D_M1011_g N_VPWR_c_540_n 0.00432313f $X=3.21 $Y=2.465 $X2=0 $Y2=0
cc_265 N_D_M1011_g N_VPWR_c_530_n 0.00637348f $X=3.21 $Y=2.465 $X2=0 $Y2=0
cc_266 N_D_M1003_g N_VGND_c_661_n 0.00882187f $X=3.28 $Y=0.655 $X2=0 $Y2=0
cc_267 N_D_M1003_g N_VGND_c_669_n 0.00585385f $X=3.28 $Y=0.655 $X2=0 $Y2=0
cc_268 N_D_M1003_g N_VGND_c_671_n 0.0112674f $X=3.28 $Y=0.655 $X2=0 $Y2=0
cc_269 N_C_M1005_g N_A_49_131#_M1010_g 0.0341548f $X=3.64 $Y=0.655 $X2=0 $Y2=0
cc_270 C N_A_49_131#_M1010_g 0.00622888f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_271 N_C_c_327_n N_A_49_131#_M1010_g 0.0202556f $X=3.73 $Y=1.375 $X2=0 $Y2=0
cc_272 N_C_M1000_g N_A_49_131#_c_364_n 0.012967f $X=3.64 $Y=2.465 $X2=0 $Y2=0
cc_273 N_C_M1000_g N_A_49_131#_c_360_n 2.40819e-19 $X=3.64 $Y=2.465 $X2=0 $Y2=0
cc_274 C N_A_49_131#_c_360_n 0.0308984f $X=3.515 $Y=1.21 $X2=0 $Y2=0
cc_275 N_C_c_327_n N_A_49_131#_c_360_n 2.4405e-19 $X=3.73 $Y=1.375 $X2=0 $Y2=0
cc_276 N_C_M1000_g N_A_49_131#_c_361_n 0.0470571f $X=3.64 $Y=2.465 $X2=0 $Y2=0
cc_277 N_C_M1000_g N_VPWR_c_534_n 0.0034189f $X=3.64 $Y=2.465 $X2=0 $Y2=0
cc_278 N_C_M1000_g N_VPWR_c_540_n 0.00432313f $X=3.64 $Y=2.465 $X2=0 $Y2=0
cc_279 N_C_M1000_g N_VPWR_c_530_n 0.00628719f $X=3.64 $Y=2.465 $X2=0 $Y2=0
cc_280 N_C_M1005_g N_VGND_c_669_n 0.00357877f $X=3.64 $Y=0.655 $X2=0 $Y2=0
cc_281 N_C_M1005_g N_VGND_c_671_n 0.00554206f $X=3.64 $Y=0.655 $X2=0 $Y2=0
cc_282 N_A_49_131#_M1008_g N_A_929_21#_M1018_g 0.0365159f $X=4.18 $Y=2.465 $X2=0
+ $Y2=0
cc_283 N_A_49_131#_c_364_n N_A_929_21#_M1018_g 0.0181188f $X=4.79 $Y=2.555 $X2=0
+ $Y2=0
cc_284 N_A_49_131#_c_359_n N_A_929_21#_M1018_g 0.0140491f $X=4.79 $Y=1.7 $X2=0
+ $Y2=0
cc_285 N_A_49_131#_c_367_n N_A_929_21#_M1018_g 0.0164506f $X=4.875 $Y=2.465
+ $X2=0 $Y2=0
cc_286 N_A_49_131#_M1010_g N_A_929_21#_c_450_n 0.00155568f $X=4.18 $Y=0.655
+ $X2=0 $Y2=0
cc_287 N_A_49_131#_c_359_n N_A_929_21#_c_450_n 0.0248946f $X=4.79 $Y=1.7 $X2=0
+ $Y2=0
cc_288 N_A_49_131#_c_360_n N_A_929_21#_c_450_n 0.00702397f $X=4.27 $Y=1.51 $X2=0
+ $Y2=0
cc_289 N_A_49_131#_c_359_n N_A_929_21#_c_451_n 0.00418157f $X=4.79 $Y=1.7 $X2=0
+ $Y2=0
cc_290 N_A_49_131#_c_360_n N_A_929_21#_c_451_n 0.00438473f $X=4.27 $Y=1.51 $X2=0
+ $Y2=0
cc_291 N_A_49_131#_c_361_n N_A_929_21#_c_451_n 0.0204625f $X=4.27 $Y=1.51 $X2=0
+ $Y2=0
cc_292 N_A_49_131#_c_359_n N_A_929_21#_c_453_n 0.00777817f $X=4.79 $Y=1.7 $X2=0
+ $Y2=0
cc_293 N_A_49_131#_c_367_n N_A_929_21#_c_453_n 0.0107368f $X=4.875 $Y=2.465
+ $X2=0 $Y2=0
cc_294 N_A_49_131#_M1010_g N_A_929_21#_c_454_n 0.0375744f $X=4.18 $Y=0.655 $X2=0
+ $Y2=0
cc_295 N_A_49_131#_c_367_n N_A_N_M1002_g 0.00637803f $X=4.875 $Y=2.465 $X2=0
+ $Y2=0
cc_296 N_A_49_131#_c_359_n N_A_N_c_501_n 0.00167544f $X=4.79 $Y=1.7 $X2=0 $Y2=0
cc_297 N_A_49_131#_c_364_n N_VPWR_M1012_d 0.00861232f $X=4.79 $Y=2.555 $X2=-0.19
+ $Y2=-0.245
cc_298 N_A_49_131#_c_364_n N_VPWR_M1009_s 0.00409097f $X=4.79 $Y=2.555 $X2=0
+ $Y2=0
cc_299 N_A_49_131#_c_364_n N_VPWR_M1017_s 0.00715823f $X=4.79 $Y=2.555 $X2=0
+ $Y2=0
cc_300 N_A_49_131#_c_364_n N_VPWR_M1000_d 0.00609136f $X=4.79 $Y=2.555 $X2=0
+ $Y2=0
cc_301 N_A_49_131#_c_364_n N_VPWR_M1018_d 0.00926781f $X=4.79 $Y=2.555 $X2=0
+ $Y2=0
cc_302 N_A_49_131#_c_367_n N_VPWR_M1018_d 0.00959818f $X=4.875 $Y=2.465 $X2=0
+ $Y2=0
cc_303 N_A_49_131#_c_364_n N_VPWR_c_531_n 0.0210041f $X=4.79 $Y=2.555 $X2=0
+ $Y2=0
cc_304 N_A_49_131#_c_364_n N_VPWR_c_532_n 0.0163012f $X=4.79 $Y=2.555 $X2=0
+ $Y2=0
cc_305 N_A_49_131#_c_364_n N_VPWR_c_533_n 0.0241559f $X=4.79 $Y=2.555 $X2=0
+ $Y2=0
cc_306 N_A_49_131#_M1008_g N_VPWR_c_534_n 0.00325112f $X=4.18 $Y=2.465 $X2=0
+ $Y2=0
cc_307 N_A_49_131#_c_364_n N_VPWR_c_534_n 0.0214374f $X=4.79 $Y=2.555 $X2=0
+ $Y2=0
cc_308 N_A_49_131#_M1008_g N_VPWR_c_535_n 0.00218158f $X=4.18 $Y=2.465 $X2=0
+ $Y2=0
cc_309 N_A_49_131#_c_364_n N_VPWR_c_535_n 0.0109009f $X=4.79 $Y=2.555 $X2=0
+ $Y2=0
cc_310 N_A_49_131#_c_364_n N_VPWR_c_536_n 0.00723404f $X=4.79 $Y=2.555 $X2=0
+ $Y2=0
cc_311 N_A_49_131#_c_364_n N_VPWR_c_538_n 0.00807238f $X=4.79 $Y=2.555 $X2=0
+ $Y2=0
cc_312 N_A_49_131#_c_364_n N_VPWR_c_540_n 0.00861f $X=4.79 $Y=2.555 $X2=0 $Y2=0
cc_313 N_A_49_131#_c_364_n N_VPWR_c_542_n 0.00840615f $X=4.79 $Y=2.555 $X2=0
+ $Y2=0
cc_314 N_A_49_131#_c_365_n N_VPWR_c_542_n 0.00456049f $X=0.455 $Y=2.555 $X2=0
+ $Y2=0
cc_315 N_A_49_131#_M1008_g N_VPWR_c_543_n 0.00432313f $X=4.18 $Y=2.465 $X2=0
+ $Y2=0
cc_316 N_A_49_131#_c_364_n N_VPWR_c_543_n 0.00954063f $X=4.79 $Y=2.555 $X2=0
+ $Y2=0
cc_317 N_A_49_131#_M1008_g N_VPWR_c_530_n 0.00642496f $X=4.18 $Y=2.465 $X2=0
+ $Y2=0
cc_318 N_A_49_131#_c_364_n N_VPWR_c_530_n 0.0833352f $X=4.79 $Y=2.555 $X2=0
+ $Y2=0
cc_319 N_A_49_131#_c_365_n N_VPWR_c_530_n 0.00729675f $X=0.455 $Y=2.555 $X2=0
+ $Y2=0
cc_320 N_A_49_131#_c_364_n N_X_M1004_d 0.00543856f $X=4.79 $Y=2.555 $X2=0 $Y2=0
cc_321 N_A_49_131#_c_364_n N_X_M1014_d 0.00543856f $X=4.79 $Y=2.555 $X2=0 $Y2=0
cc_322 N_A_49_131#_c_358_n N_X_c_612_n 7.4539e-19 $X=0.37 $Y=0.865 $X2=0 $Y2=0
cc_323 N_A_49_131#_c_364_n N_X_c_612_n 0.00614205f $X=4.79 $Y=2.555 $X2=0 $Y2=0
cc_324 N_A_49_131#_c_364_n N_X_c_610_n 0.042285f $X=4.79 $Y=2.555 $X2=0 $Y2=0
cc_325 N_A_49_131#_c_358_n N_VGND_c_663_n 0.00421272f $X=0.37 $Y=0.865 $X2=0
+ $Y2=0
cc_326 N_A_49_131#_M1010_g N_VGND_c_669_n 0.00357877f $X=4.18 $Y=0.655 $X2=0
+ $Y2=0
cc_327 N_A_49_131#_M1010_g N_VGND_c_671_n 0.00599809f $X=4.18 $Y=0.655 $X2=0
+ $Y2=0
cc_328 N_A_49_131#_c_358_n N_VGND_c_671_n 0.00717262f $X=0.37 $Y=0.865 $X2=0
+ $Y2=0
cc_329 N_A_929_21#_c_453_n N_A_N_M1002_g 0.00565699f $X=5.49 $Y=1.93 $X2=0 $Y2=0
cc_330 N_A_929_21#_c_448_n N_A_N_c_500_n 0.00544769f $X=5.885 $Y=1.16 $X2=0
+ $Y2=0
cc_331 N_A_929_21#_c_456_n N_A_N_c_500_n 0.00437629f $X=5.475 $Y=2.095 $X2=0
+ $Y2=0
cc_332 N_A_929_21#_c_453_n N_A_N_c_500_n 0.0144327f $X=5.49 $Y=1.93 $X2=0 $Y2=0
cc_333 N_A_929_21#_M1018_g N_A_N_c_501_n 0.023439f $X=4.72 $Y=2.465 $X2=0 $Y2=0
cc_334 N_A_929_21#_c_447_n N_A_N_c_501_n 0.00565616f $X=5.34 $Y=1.16 $X2=0 $Y2=0
cc_335 N_A_929_21#_c_448_n N_A_N_M1016_g 0.0173358f $X=5.885 $Y=1.16 $X2=0 $Y2=0
cc_336 N_A_929_21#_c_449_n N_A_N_M1016_g 5.62685e-19 $X=5.98 $Y=0.86 $X2=0 $Y2=0
cc_337 N_A_929_21#_c_451_n N_A_N_M1016_g 0.00320882f $X=4.81 $Y=1.35 $X2=0 $Y2=0
cc_338 N_A_929_21#_c_453_n N_A_N_M1016_g 0.00565643f $X=5.49 $Y=1.93 $X2=0 $Y2=0
cc_339 N_A_929_21#_c_448_n N_A_N_c_503_n 0.00451636f $X=5.885 $Y=1.16 $X2=0
+ $Y2=0
cc_340 N_A_929_21#_c_448_n N_A_N_c_504_n 0.0342204f $X=5.885 $Y=1.16 $X2=0 $Y2=0
cc_341 N_A_929_21#_c_453_n N_A_N_c_504_n 0.0245021f $X=5.49 $Y=1.93 $X2=0 $Y2=0
cc_342 N_A_929_21#_M1018_g N_VPWR_c_535_n 0.0117039f $X=4.72 $Y=2.465 $X2=0
+ $Y2=0
cc_343 N_A_929_21#_M1018_g N_VPWR_c_543_n 0.00359504f $X=4.72 $Y=2.465 $X2=0
+ $Y2=0
cc_344 N_A_929_21#_M1018_g N_VPWR_c_530_n 0.00458255f $X=4.72 $Y=2.465 $X2=0
+ $Y2=0
cc_345 N_A_929_21#_c_448_n N_VGND_c_662_n 0.0140741f $X=5.885 $Y=1.16 $X2=0
+ $Y2=0
cc_346 N_A_929_21#_c_452_n N_VGND_c_662_n 0.0114682f $X=5.425 $Y=1.16 $X2=0
+ $Y2=0
cc_347 N_A_929_21#_c_454_n N_VGND_c_662_n 0.00196769f $X=4.81 $Y=1.185 $X2=0
+ $Y2=0
cc_348 N_A_929_21#_c_454_n N_VGND_c_669_n 0.00357877f $X=4.81 $Y=1.185 $X2=0
+ $Y2=0
cc_349 N_A_929_21#_c_449_n N_VGND_c_670_n 0.00426314f $X=5.98 $Y=0.86 $X2=0
+ $Y2=0
cc_350 N_A_929_21#_c_449_n N_VGND_c_671_n 0.00741356f $X=5.98 $Y=0.86 $X2=0
+ $Y2=0
cc_351 N_A_929_21#_c_454_n N_VGND_c_671_n 0.00693897f $X=4.81 $Y=1.185 $X2=0
+ $Y2=0
cc_352 N_A_N_c_500_n N_VGND_c_662_n 5.78859e-19 $X=5.69 $Y=1.6 $X2=0 $Y2=0
cc_353 N_A_N_M1016_g N_VGND_c_662_n 0.0135467f $X=5.765 $Y=0.855 $X2=0 $Y2=0
cc_354 N_A_N_M1016_g N_VGND_c_670_n 0.00336585f $X=5.765 $Y=0.855 $X2=0 $Y2=0
cc_355 N_A_N_M1016_g N_VGND_c_671_n 0.00389709f $X=5.765 $Y=0.855 $X2=0 $Y2=0
cc_356 N_VPWR_c_530_n N_X_M1004_d 0.00346035f $X=6 $Y=3.33 $X2=0 $Y2=0
cc_357 N_VPWR_c_530_n N_X_M1014_d 0.00346035f $X=6 $Y=3.33 $X2=0 $Y2=0
cc_358 N_VPWR_M1012_d N_X_c_612_n 0.00518301f $X=0.68 $Y=1.835 $X2=0 $Y2=0
cc_359 N_VPWR_M1009_s N_X_c_610_n 0.00242422f $X=1.85 $Y=1.835 $X2=0 $Y2=0
cc_360 N_X_c_608_n N_VGND_c_659_n 0.00965371f $X=1.655 $Y=1.16 $X2=0 $Y2=0
cc_361 N_X_c_607_n N_VGND_c_660_n 0.0216087f $X=2.325 $Y=1.16 $X2=0 $Y2=0
cc_362 N_X_c_606_n N_VGND_c_665_n 0.0138717f $X=1.56 $Y=0.42 $X2=0 $Y2=0
cc_363 N_X_c_654_p N_VGND_c_667_n 0.0124525f $X=2.42 $Y=0.42 $X2=0 $Y2=0
cc_364 N_X_M1006_d N_VGND_c_671_n 0.00397496f $X=1.42 $Y=0.235 $X2=0 $Y2=0
cc_365 N_X_M1013_d N_VGND_c_671_n 0.00536646f $X=2.28 $Y=0.235 $X2=0 $Y2=0
cc_366 N_X_c_606_n N_VGND_c_671_n 0.00886411f $X=1.56 $Y=0.42 $X2=0 $Y2=0
cc_367 N_X_c_654_p N_VGND_c_671_n 0.00730901f $X=2.42 $Y=0.42 $X2=0 $Y2=0
cc_368 N_VGND_c_671_n A_671_47# 0.00534151f $X=6 $Y=0 $X2=-0.19 $Y2=-0.245
cc_369 N_VGND_c_671_n A_743_47# 0.0031466f $X=6 $Y=0 $X2=-0.19 $Y2=-0.245
cc_370 N_VGND_c_671_n A_851_47# 0.0031466f $X=6 $Y=0 $X2=-0.19 $Y2=-0.245
