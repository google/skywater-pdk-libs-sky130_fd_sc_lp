* File: sky130_fd_sc_lp__sdfsbp_lp.pex.spice
* Created: Wed Sep  2 10:35:29 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__SDFSBP_LP%SCE 3 7 9 13 17 22 24 25 26 28 29 30 34 36
+ 37 38 42 43 45 46 55 59
c109 34 0 1.88859e-19 $X=1.095 $Y=1.02
r110 46 59 8.06514 $w=4.68e-07 $l=1.15e-07 $layer=LI1_cond $X=2.16 $Y=1.045
+ $X2=2.275 $Y2=1.045
r111 45 55 4.00199 $w=4.68e-07 $l=1.15e-07 $layer=LI1_cond $X=1.68 $Y=1.045
+ $X2=1.565 $Y2=1.045
r112 42 43 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.675
+ $Y=1.285 $X2=2.675 $Y2=1.285
r113 40 42 0.177299 $w=3.23e-07 $l=5e-09 $layer=LI1_cond $X=2.672 $Y=1.28
+ $X2=2.672 $Y2=1.285
r114 38 40 7.72402 $w=1.7e-07 $l=2.00035e-07 $layer=LI1_cond $X=2.51 $Y=1.195
+ $X2=2.672 $Y2=1.28
r115 38 59 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=2.51 $Y=1.195
+ $X2=2.275 $Y2=1.195
r116 37 45 3.05382 $w=4.68e-07 $l=1.2e-07 $layer=LI1_cond $X=1.8 $Y=1.045
+ $X2=1.68 $Y2=1.045
r117 36 46 3.05382 $w=4.68e-07 $l=1.2e-07 $layer=LI1_cond $X=2.04 $Y=1.045
+ $X2=2.16 $Y2=1.045
r118 36 37 6.10763 $w=4.68e-07 $l=2.4e-07 $layer=LI1_cond $X=2.04 $Y=1.045
+ $X2=1.8 $Y2=1.045
r119 34 52 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=1.095 $Y=1.02
+ $X2=1.095 $Y2=1.11
r120 34 51 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.095 $Y=1.02
+ $X2=1.095 $Y2=0.855
r121 33 55 16.4136 $w=3.28e-07 $l=4.7e-07 $layer=LI1_cond $X=1.095 $Y=1.02
+ $X2=1.565 $Y2=1.02
r122 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.095
+ $Y=1.02 $X2=1.095 $Y2=1.02
r123 29 43 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.675 $Y=1.625
+ $X2=2.675 $Y2=1.285
r124 29 30 31.2043 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.675 $Y=1.625
+ $X2=2.675 $Y2=1.79
r125 28 43 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.675 $Y=1.12
+ $X2=2.675 $Y2=1.285
r126 26 28 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=2.585 $Y=0.88
+ $X2=2.585 $Y2=1.12
r127 25 26 58.3064 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=2.57 $Y=0.73
+ $X2=2.57 $Y2=0.88
r128 22 30 187.582 $w=2.5e-07 $l=7.55e-07 $layer=POLY_cond $X=2.655 $Y=2.545
+ $X2=2.655 $Y2=1.79
r129 17 25 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.555 $Y=0.445
+ $X2=2.555 $Y2=0.73
r130 13 51 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=1.005 $Y=0.445
+ $X2=1.005 $Y2=0.855
r131 10 24 9.46703 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.69 $Y=1.11
+ $X2=0.555 $Y2=1.11
r132 9 52 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.93 $Y=1.11
+ $X2=1.095 $Y2=1.11
r133 9 10 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=0.93 $Y=1.11
+ $X2=0.69 $Y2=1.11
r134 5 24 15.9654 $w=2e-07 $l=1.00623e-07 $layer=POLY_cond $X=0.615 $Y=1.035
+ $X2=0.555 $Y2=1.11
r135 5 7 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=0.615 $Y=1.035
+ $X2=0.615 $Y2=0.445
r136 1 24 15.9654 $w=2e-07 $l=7.98436e-08 $layer=POLY_cond $X=0.545 $Y=1.185
+ $X2=0.555 $Y2=1.11
r137 1 3 337.897 $w=2.5e-07 $l=1.36e-06 $layer=POLY_cond $X=0.545 $Y=1.185
+ $X2=0.545 $Y2=2.545
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSBP_LP%A_27_409# 1 2 9 12 13 15 16 17 20 24 28 34
+ 37
c67 34 0 2.24716e-19 $X=1.22 $Y=1.59
c68 24 0 1.88859e-19 $X=0.4 $Y=0.47
c69 20 0 1.96756e-19 $X=1.735 $Y=0.805
r70 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.22
+ $Y=1.59 $X2=1.22 $Y2=1.59
r71 32 37 1.95047 $w=3.3e-07 $l=2.25e-07 $layer=LI1_cond $X=0.565 $Y=1.59
+ $X2=0.34 $Y2=1.59
r72 32 34 22.8742 $w=3.28e-07 $l=6.55e-07 $layer=LI1_cond $X=0.565 $Y=1.59
+ $X2=1.22 $Y2=1.59
r73 28 30 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=0.28 $Y=2.19 $X2=0.28
+ $Y2=2.9
r74 26 37 4.48582 $w=3.9e-07 $l=1.92678e-07 $layer=LI1_cond $X=0.28 $Y=1.755
+ $X2=0.34 $Y2=1.59
r75 26 28 15.1913 $w=3.28e-07 $l=4.35e-07 $layer=LI1_cond $X=0.28 $Y=1.755
+ $X2=0.28 $Y2=2.19
r76 22 37 4.48582 $w=3.9e-07 $l=1.65e-07 $layer=LI1_cond $X=0.34 $Y=1.425
+ $X2=0.34 $Y2=1.59
r77 22 24 25.3834 $w=4.48e-07 $l=9.55e-07 $layer=LI1_cond $X=0.34 $Y=1.425
+ $X2=0.34 $Y2=0.47
r78 18 20 41.0213 $w=1.5e-07 $l=8e-08 $layer=POLY_cond $X=1.655 $Y=0.805
+ $X2=1.735 $Y2=0.805
r79 16 35 50.7098 $w=3.3e-07 $l=2.9e-07 $layer=POLY_cond $X=1.51 $Y=1.59
+ $X2=1.22 $Y2=1.59
r80 16 17 1.50692 $w=3.3e-07 $l=1.25e-07 $layer=POLY_cond $X=1.51 $Y=1.59
+ $X2=1.635 $Y2=1.59
r81 13 20 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.735 $Y=0.73
+ $X2=1.735 $Y2=0.805
r82 13 15 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=1.735 $Y=0.73
+ $X2=1.735 $Y2=0.445
r83 12 17 30.2679 $w=2e-07 $l=1.74714e-07 $layer=POLY_cond $X=1.655 $Y=1.425
+ $X2=1.635 $Y2=1.59
r84 11 18 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.655 $Y=0.88
+ $X2=1.655 $Y2=0.805
r85 11 12 279.457 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=1.655 $Y=0.88
+ $X2=1.655 $Y2=1.425
r86 7 17 30.2679 $w=2e-07 $l=1.65e-07 $layer=POLY_cond $X=1.635 $Y=1.755
+ $X2=1.635 $Y2=1.59
r87 7 9 196.278 $w=2.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.635 $Y=1.755
+ $X2=1.635 $Y2=2.545
r88 2 30 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.045 $X2=0.28 $Y2=2.9
r89 2 28 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.045 $X2=0.28 $Y2=2.19
r90 1 24 182 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_NDIFF $count=1 $X=0.255
+ $Y=0.235 $X2=0.4 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSBP_LP%D 3 7 9 10 14
c43 14 0 1.18806e-19 $X=2.135 $Y=1.625
c44 10 0 1.96756e-19 $X=2.16 $Y=1.665
c45 7 0 1.05911e-19 $X=2.125 $Y=0.445
r46 14 17 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.135 $Y=1.625
+ $X2=2.135 $Y2=1.79
r47 14 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.135 $Y=1.625
+ $X2=2.135 $Y2=1.46
r48 10 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.135
+ $Y=1.625 $X2=2.135 $Y2=1.625
r49 9 10 15.8897 $w=3.28e-07 $l=4.55e-07 $layer=LI1_cond $X=1.68 $Y=1.625
+ $X2=2.135 $Y2=1.625
r50 7 16 520.457 $w=1.5e-07 $l=1.015e-06 $layer=POLY_cond $X=2.125 $Y=0.445
+ $X2=2.125 $Y2=1.46
r51 3 17 187.582 $w=2.5e-07 $l=7.55e-07 $layer=POLY_cond $X=2.165 $Y=2.545
+ $X2=2.165 $Y2=1.79
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSBP_LP%SCD 1 3 6 12 14 15 19 21
c53 19 0 1.86498e-19 $X=3.525 $Y=1.275
c54 6 0 4.76528e-20 $X=3.185 $Y=2.545
r55 19 22 63.0283 $w=6.3e-07 $l=5.05e-07 $layer=POLY_cond $X=3.375 $Y=1.275
+ $X2=3.375 $Y2=1.78
r56 19 21 50.3829 $w=6.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.375 $Y=1.275
+ $X2=3.375 $Y2=1.11
r57 14 15 14.0454 $w=3.18e-07 $l=3.9e-07 $layer=LI1_cond $X=3.525 $Y=1.275
+ $X2=3.525 $Y2=1.665
r58 14 19 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.525
+ $Y=1.275 $X2=3.525 $Y2=1.275
r59 10 12 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=2.945 $Y=0.805
+ $X2=3.155 $Y2=0.805
r60 8 12 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.155 $Y=0.88
+ $X2=3.155 $Y2=0.805
r61 8 21 117.936 $w=1.5e-07 $l=2.3e-07 $layer=POLY_cond $X=3.155 $Y=0.88
+ $X2=3.155 $Y2=1.11
r62 6 22 190.067 $w=2.5e-07 $l=7.65e-07 $layer=POLY_cond $X=3.185 $Y=2.545
+ $X2=3.185 $Y2=1.78
r63 1 10 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.945 $Y=0.73
+ $X2=2.945 $Y2=0.805
r64 1 3 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.945 $Y=0.73 $X2=2.945
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSBP_LP%CLK 3 6 9 13 16 17 20
c53 9 0 2.10375e-19 $X=4.28 $Y=2.545
c54 6 0 1.66046e-19 $X=4.282 $Y=1.588
r55 20 22 30.6629 $w=3.85e-07 $l=1.65e-07 $layer=POLY_cond $X=4.282 $Y=1.615
+ $X2=4.282 $Y2=1.78
r56 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.31
+ $Y=1.615 $X2=4.31 $Y2=1.615
r57 17 21 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=4.56 $Y=1.615
+ $X2=4.31 $Y2=1.615
r58 9 22 190.067 $w=2.5e-07 $l=7.65e-07 $layer=POLY_cond $X=4.28 $Y=2.545
+ $X2=4.28 $Y2=1.78
r59 6 20 3.9003 $w=3.85e-07 $l=2.7e-08 $layer=POLY_cond $X=4.282 $Y=1.588
+ $X2=4.282 $Y2=1.615
r60 6 16 39.4364 $w=3.85e-07 $l=2.73e-07 $layer=POLY_cond $X=4.282 $Y=1.588
+ $X2=4.282 $Y2=1.315
r61 1 16 24.5286 $w=3.85e-07 $l=1.5e-07 $layer=POLY_cond $X=4.345 $Y=1.165
+ $X2=4.345 $Y2=1.315
r62 1 13 199.979 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=4.525 $Y=1.165
+ $X2=4.525 $Y2=0.775
r63 1 3 199.979 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=4.165 $Y=1.165
+ $X2=4.165 $Y2=0.775
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSBP_LP%A_987_409# 1 2 9 13 17 20 24 26 27 29 31
+ 34 35 37 40 41 42 45 46 49 50 55 61 63 64 65 70 79
c212 63 0 1.7417e-19 $X=6.13 $Y=1.54
c213 50 0 2.85022e-19 $X=10.715 $Y=1.69
c214 46 0 3.84399e-20 $X=9.98 $Y=1.32
c215 35 0 6.73817e-20 $X=6.74 $Y=1.465
c216 27 0 4.93603e-20 $X=5.24 $Y=2.98
c217 24 0 1.61015e-19 $X=5.075 $Y=2.475
r218 70 83 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=10.88 $Y=1.77
+ $X2=10.88 $Y2=1.935
r219 69 70 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.88
+ $Y=1.77 $X2=10.88 $Y2=1.77
r220 62 63 3.29577 $w=4.78e-07 $l=8.5e-08 $layer=LI1_cond $X=6.045 $Y=1.54
+ $X2=6.13 $Y2=1.54
r221 61 74 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.84 $Y=1.615
+ $X2=5.84 $Y2=1.78
r222 60 62 5.10825 $w=4.78e-07 $l=2.05e-07 $layer=LI1_cond $X=5.84 $Y=1.54
+ $X2=6.045 $Y2=1.54
r223 60 61 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.84
+ $Y=1.615 $X2=5.84 $Y2=1.615
r224 57 60 2.11806 $w=4.78e-07 $l=8.5e-08 $layer=LI1_cond $X=5.755 $Y=1.54
+ $X2=5.84 $Y2=1.54
r225 53 55 6.64871 $w=3.88e-07 $l=2.25e-07 $layer=LI1_cond $X=5.53 $Y=0.81
+ $X2=5.755 $Y2=0.81
r226 51 65 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.145 $Y=1.69
+ $X2=9.98 $Y2=1.69
r227 50 69 3.47907 $w=2.63e-07 $l=8e-08 $layer=LI1_cond $X=10.847 $Y=1.69
+ $X2=10.847 $Y2=1.77
r228 50 51 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=10.715 $Y=1.69
+ $X2=10.145 $Y2=1.69
r229 48 65 3.70735 $w=2.5e-07 $l=1.18427e-07 $layer=LI1_cond $X=9.9 $Y=1.775
+ $X2=9.98 $Y2=1.69
r230 48 49 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=9.9 $Y=1.775
+ $X2=9.9 $Y2=2.515
r231 46 79 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=9.98 $Y=1.32
+ $X2=9.98 $Y2=1.155
r232 45 46 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.98
+ $Y=1.32 $X2=9.98 $Y2=1.32
r233 43 65 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=9.98 $Y=1.605
+ $X2=9.98 $Y2=1.69
r234 43 45 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=9.98 $Y=1.605
+ $X2=9.98 $Y2=1.32
r235 41 49 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.815 $Y=2.6
+ $X2=9.9 $Y2=2.515
r236 41 42 147.118 $w=1.68e-07 $l=2.255e-06 $layer=LI1_cond $X=9.815 $Y=2.6
+ $X2=7.56 $Y2=2.6
r237 39 42 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.475 $Y=2.685
+ $X2=7.56 $Y2=2.6
r238 39 40 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=7.475 $Y=2.685
+ $X2=7.475 $Y2=2.895
r239 38 64 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.13 $Y=2.98
+ $X2=6.045 $Y2=2.98
r240 37 40 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.39 $Y=2.98
+ $X2=7.475 $Y2=2.895
r241 37 38 82.2032 $w=1.68e-07 $l=1.26e-06 $layer=LI1_cond $X=7.39 $Y=2.98
+ $X2=6.13 $Y2=2.98
r242 35 76 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.74 $Y=1.465
+ $X2=6.74 $Y2=1.3
r243 34 63 21.3027 $w=3.28e-07 $l=6.1e-07 $layer=LI1_cond $X=6.74 $Y=1.465
+ $X2=6.13 $Y2=1.465
r244 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.74
+ $Y=1.465 $X2=6.74 $Y2=1.465
r245 31 64 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.045 $Y=2.895
+ $X2=6.045 $Y2=2.98
r246 30 62 6.90116 $w=1.7e-07 $l=2.4e-07 $layer=LI1_cond $X=6.045 $Y=1.78
+ $X2=6.045 $Y2=1.54
r247 30 31 72.7433 $w=1.68e-07 $l=1.115e-06 $layer=LI1_cond $X=6.045 $Y=1.78
+ $X2=6.045 $Y2=2.895
r248 29 57 6.90116 $w=1.7e-07 $l=2.4e-07 $layer=LI1_cond $X=5.755 $Y=1.3
+ $X2=5.755 $Y2=1.54
r249 28 55 5.6248 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=5.755 $Y=1.005
+ $X2=5.755 $Y2=0.81
r250 28 29 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=5.755 $Y=1.005
+ $X2=5.755 $Y2=1.3
r251 26 64 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.96 $Y=2.98
+ $X2=6.045 $Y2=2.98
r252 26 27 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=5.96 $Y=2.98
+ $X2=5.24 $Y2=2.98
r253 22 27 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.075 $Y=2.895
+ $X2=5.24 $Y2=2.98
r254 22 24 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=5.075 $Y=2.895
+ $X2=5.075 $Y2=2.475
r255 20 83 163.979 $w=2.5e-07 $l=6.6e-07 $layer=POLY_cond $X=10.84 $Y=2.595
+ $X2=10.84 $Y2=1.935
r256 17 79 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=10.04 $Y=0.835
+ $X2=10.04 $Y2=1.155
r257 13 76 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=6.83 $Y=0.835
+ $X2=6.83 $Y2=1.3
r258 9 74 202.49 $w=2.5e-07 $l=8.15e-07 $layer=POLY_cond $X=5.88 $Y=2.595
+ $X2=5.88 $Y2=1.78
r259 2 24 300 $w=1.7e-07 $l=4.95076e-07 $layer=licon1_PDIFF $count=2 $X=4.935
+ $Y=2.045 $X2=5.075 $Y2=2.475
r260 1 53 182 $w=1.7e-07 $l=3.07124e-07 $layer=licon1_NDIFF $count=1 $X=5.39
+ $Y=0.565 $X2=5.53 $Y2=0.81
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSBP_LP%A_1423_99# 1 2 9 13 18 19 20 21 22 24 27
+ 31
c81 27 0 2.90644e-20 $X=8.18 $Y=1.225
c82 22 0 1.75395e-19 $X=7.765 $Y=2.21
c83 20 0 8.26509e-20 $X=8.095 $Y=1.31
r84 33 35 13.9889 $w=3.3e-07 $l=8e-08 $layer=POLY_cond $X=7.19 $Y=1.675 $X2=7.27
+ $Y2=1.675
r85 28 31 4.97969 $w=4.03e-07 $l=1.75e-07 $layer=LI1_cond $X=8.18 $Y=0.817
+ $X2=8.355 $Y2=0.817
r86 26 28 5.85399 $w=1.7e-07 $l=2.03e-07 $layer=LI1_cond $X=8.18 $Y=1.02
+ $X2=8.18 $Y2=0.817
r87 26 27 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=8.18 $Y=1.02
+ $X2=8.18 $Y2=1.225
r88 22 24 30.8855 $w=2.48e-07 $l=6.7e-07 $layer=LI1_cond $X=7.765 $Y=2.21
+ $X2=8.435 $Y2=2.21
r89 20 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.095 $Y=1.31
+ $X2=8.18 $Y2=1.225
r90 20 21 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=8.095 $Y=1.31
+ $X2=7.765 $Y2=1.31
r91 19 35 57.7042 $w=3.3e-07 $l=3.3e-07 $layer=POLY_cond $X=7.6 $Y=1.675
+ $X2=7.27 $Y2=1.675
r92 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.6
+ $Y=1.675 $X2=7.6 $Y2=1.675
r93 16 22 6.98653 $w=2.5e-07 $l=2.18746e-07 $layer=LI1_cond $X=7.6 $Y=2.085
+ $X2=7.765 $Y2=2.21
r94 16 18 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=7.6 $Y=2.085 $X2=7.6
+ $Y2=1.675
r95 15 21 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=7.6 $Y=1.395
+ $X2=7.765 $Y2=1.31
r96 15 18 9.7783 $w=3.28e-07 $l=2.8e-07 $layer=LI1_cond $X=7.6 $Y=1.395 $X2=7.6
+ $Y2=1.675
r97 11 35 9.34494 $w=2.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.27 $Y=1.84
+ $X2=7.27 $Y2=1.675
r98 11 13 187.582 $w=2.5e-07 $l=7.55e-07 $layer=POLY_cond $X=7.27 $Y=1.84
+ $X2=7.27 $Y2=2.595
r99 7 33 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.19 $Y=1.51
+ $X2=7.19 $Y2=1.675
r100 7 9 346.117 $w=1.5e-07 $l=6.75e-07 $layer=POLY_cond $X=7.19 $Y=1.51
+ $X2=7.19 $Y2=0.835
r101 2 24 600 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_PDIFF $count=1 $X=8.295
+ $Y=2.095 $X2=8.435 $Y2=2.25
r102 1 31 182 $w=1.7e-07 $l=2.5229e-07 $layer=licon1_NDIFF $count=1 $X=8.21
+ $Y=0.625 $X2=8.355 $Y2=0.815
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSBP_LP%A_1201_419# 1 2 9 13 14 15 17 20 24 28 29
+ 32 34 35 36 39 40 43 44 45 46 49 52 54 55 56 60 64 69 70 73
c198 69 0 1.82916e-19 $X=9.44 $Y=1.365
c199 60 0 8.29256e-20 $X=6.615 $Y=0.835
c200 35 0 6.73817e-20 $X=6.64 $Y=2.16
c201 20 0 6.26699e-20 $X=9.48 $Y=2.595
r202 69 70 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=9.44
+ $Y=1.365 $X2=9.44 $Y2=1.365
r203 65 67 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=8.53 $Y=1.285
+ $X2=8.785 $Y2=1.285
r204 60 62 4.36531 $w=3.28e-07 $l=1.25e-07 $layer=LI1_cond $X=6.615 $Y=0.835
+ $X2=6.615 $Y2=0.96
r205 56 67 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=8.87 $Y=1.285
+ $X2=8.785 $Y2=1.285
r206 55 69 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.275 $Y=1.285
+ $X2=9.44 $Y2=1.285
r207 55 56 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=9.275 $Y=1.285
+ $X2=8.87 $Y2=1.285
r208 54 67 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.785 $Y=1.2
+ $X2=8.785 $Y2=1.285
r209 53 54 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=8.785 $Y=0.435
+ $X2=8.785 $Y2=1.2
r210 51 65 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.53 $Y=1.37
+ $X2=8.53 $Y2=1.285
r211 51 52 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=8.53 $Y=1.37
+ $X2=8.53 $Y2=1.575
r212 49 73 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.17 $Y=1.74
+ $X2=8.17 $Y2=1.575
r213 48 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.17
+ $Y=1.74 $X2=8.17 $Y2=1.74
r214 46 52 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=8.445 $Y=1.74
+ $X2=8.53 $Y2=1.575
r215 46 48 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=8.445 $Y=1.74
+ $X2=8.17 $Y2=1.74
r216 44 53 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.7 $Y=0.35
+ $X2=8.785 $Y2=0.435
r217 44 45 51.2139 $w=1.68e-07 $l=7.85e-07 $layer=LI1_cond $X=8.7 $Y=0.35
+ $X2=7.915 $Y2=0.35
r218 42 45 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.83 $Y=0.435
+ $X2=7.915 $Y2=0.35
r219 42 43 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=7.83 $Y=0.435
+ $X2=7.83 $Y2=0.875
r220 41 64 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.255 $Y=0.96
+ $X2=7.17 $Y2=0.96
r221 40 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.745 $Y=0.96
+ $X2=7.83 $Y2=0.875
r222 40 41 31.9679 $w=1.68e-07 $l=4.9e-07 $layer=LI1_cond $X=7.745 $Y=0.96
+ $X2=7.255 $Y2=0.96
r223 38 64 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.17 $Y=1.045
+ $X2=7.17 $Y2=0.96
r224 38 39 67.1979 $w=1.68e-07 $l=1.03e-06 $layer=LI1_cond $X=7.17 $Y=1.045
+ $X2=7.17 $Y2=2.075
r225 37 62 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.78 $Y=0.96
+ $X2=6.615 $Y2=0.96
r226 36 64 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.085 $Y=0.96
+ $X2=7.17 $Y2=0.96
r227 36 37 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=7.085 $Y=0.96
+ $X2=6.78 $Y2=0.96
r228 34 39 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.085 $Y=2.16
+ $X2=7.17 $Y2=2.075
r229 34 35 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=7.085 $Y=2.16
+ $X2=6.64 $Y2=2.16
r230 30 35 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.475 $Y=2.245
+ $X2=6.64 $Y2=2.16
r231 30 32 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=6.475 $Y=2.245
+ $X2=6.475 $Y2=2.395
r232 28 70 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=9.44 $Y=1.705
+ $X2=9.44 $Y2=1.365
r233 28 29 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=9.44 $Y=1.705
+ $X2=9.44 $Y2=1.87
r234 27 70 41.8716 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=9.44 $Y=1.2
+ $X2=9.44 $Y2=1.365
r235 24 27 187.16 $w=1.5e-07 $l=3.65e-07 $layer=POLY_cond $X=9.5 $Y=0.835
+ $X2=9.5 $Y2=1.2
r236 20 29 180.129 $w=2.5e-07 $l=7.25e-07 $layer=POLY_cond $X=9.48 $Y=2.595
+ $X2=9.48 $Y2=1.87
r237 15 17 104.433 $w=1.5e-07 $l=3.25e-07 $layer=POLY_cond $X=8.57 $Y=1.16
+ $X2=8.57 $Y2=0.835
r238 13 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.495 $Y=1.235
+ $X2=8.57 $Y2=1.16
r239 13 14 82.0426 $w=1.5e-07 $l=1.6e-07 $layer=POLY_cond $X=8.495 $Y=1.235
+ $X2=8.335 $Y2=1.235
r240 11 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.26 $Y=1.31
+ $X2=8.335 $Y2=1.235
r241 11 73 135.883 $w=1.5e-07 $l=2.65e-07 $layer=POLY_cond $X=8.26 $Y=1.31
+ $X2=8.26 $Y2=1.575
r242 7 49 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.17 $Y=1.905
+ $X2=8.17 $Y2=1.74
r243 7 9 171.433 $w=2.5e-07 $l=6.9e-07 $layer=POLY_cond $X=8.17 $Y=1.905
+ $X2=8.17 $Y2=2.595
r244 2 32 600 $w=1.7e-07 $l=6.01581e-07 $layer=licon1_PDIFF $count=1 $X=6.005
+ $Y=2.095 $X2=6.475 $Y2=2.395
r245 1 60 182 $w=1.7e-07 $l=5.18459e-07 $layer=licon1_NDIFF $count=1 $X=6.395
+ $Y=0.415 $X2=6.615 $Y2=0.835
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSBP_LP%SET_B 3 7 9 11 12 13 18 20 21 24 26 33 36
+ 37 38
c129 37 0 8.27582e-20 $X=12.15 $Y=1.725
c130 24 0 6.26699e-20 $X=8.88 $Y=1.665
c131 20 0 3.84399e-20 $X=12.095 $Y=1.665
c132 7 0 1.11715e-19 $X=8.96 $Y=0.835
r133 36 39 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=12.15 $Y=1.725
+ $X2=12.15 $Y2=1.89
r134 36 38 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=12.15 $Y=1.725
+ $X2=12.15 $Y2=1.56
r135 36 37 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=12.15
+ $Y=1.725 $X2=12.15 $Y2=1.725
r136 31 33 10.4917 $w=3.3e-07 $l=6e-08 $layer=POLY_cond $X=8.9 $Y=1.715 $X2=8.96
+ $Y2=1.715
r137 28 31 34.9723 $w=3.3e-07 $l=2e-07 $layer=POLY_cond $X=8.7 $Y=1.715 $X2=8.9
+ $Y2=1.715
r138 26 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.24 $Y=1.665
+ $X2=12.24 $Y2=1.665
r139 24 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.9
+ $Y=1.715 $X2=8.9 $Y2=1.715
r140 23 24 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=1.665
+ $X2=8.88 $Y2=1.665
r141 21 23 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=9.025 $Y=1.665
+ $X2=8.88 $Y2=1.665
r142 20 26 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=12.095 $Y=1.665
+ $X2=12.24 $Y2=1.665
r143 20 21 3.7995 $w=1.4e-07 $l=3.07e-06 $layer=MET1_cond $X=12.095 $Y=1.665
+ $X2=9.025 $Y2=1.665
r144 18 39 175.16 $w=2.5e-07 $l=7.05e-07 $layer=POLY_cond $X=12.11 $Y=2.595
+ $X2=12.11 $Y2=1.89
r145 14 38 299.968 $w=1.5e-07 $l=5.85e-07 $layer=POLY_cond $X=12.06 $Y=0.975
+ $X2=12.06 $Y2=1.56
r146 12 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=11.985 $Y=0.9
+ $X2=12.06 $Y2=0.975
r147 12 13 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=11.985 $Y=0.9
+ $X2=11.615 $Y2=0.9
r148 9 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=11.54 $Y=0.825
+ $X2=11.615 $Y2=0.9
r149 9 11 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=11.54 $Y=0.825
+ $X2=11.54 $Y2=0.54
r150 5 33 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.96 $Y=1.55
+ $X2=8.96 $Y2=1.715
r151 5 7 366.628 $w=1.5e-07 $l=7.15e-07 $layer=POLY_cond $X=8.96 $Y=1.55
+ $X2=8.96 $Y2=0.835
r152 1 28 9.34494 $w=2.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.7 $Y=1.88 $X2=8.7
+ $Y2=1.715
r153 1 3 177.644 $w=2.5e-07 $l=7.15e-07 $layer=POLY_cond $X=8.7 $Y=1.88 $X2=8.7
+ $Y2=2.595
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSBP_LP%A_761_113# 1 2 9 11 13 15 16 18 20 21 23
+ 24 28 29 30 31 32 33 35 38 40 41 43 44 45 49 50 51 55 60 61 65 66 68 70
c211 65 0 1.66046e-19 $X=4.98 $Y=1.72
c212 50 0 1.55371e-19 $X=4.955 $Y=1.135
c213 43 0 1.07173e-19 $X=10.43 $Y=1.725
c214 41 0 1.82916e-19 $X=10.095 $Y=1.8
c215 40 0 1.65443e-19 $X=10.355 $Y=1.8
c216 23 0 8.29256e-20 $X=6.29 $Y=1.21
c217 15 0 1.7417e-19 $X=4.955 $Y=1.555
r218 73 75 25.3549 $w=3.3e-07 $l=1.45e-07 $layer=POLY_cond $X=4.81 $Y=1.72
+ $X2=4.955 $Y2=1.72
r219 70 72 10.1762 $w=2.48e-07 $l=1.95e-07 $layer=LI1_cond $X=3.99 $Y=0.81
+ $X2=3.99 $Y2=1.005
r220 66 75 4.37153 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=4.98 $Y=1.72
+ $X2=4.955 $Y2=1.72
r221 65 66 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.98
+ $Y=1.72 $X2=4.98 $Y2=1.72
r222 63 65 8.78052 $w=3.13e-07 $l=2.4e-07 $layer=LI1_cond $X=4.982 $Y=1.96
+ $X2=4.982 $Y2=1.72
r223 62 68 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.18 $Y=2.045
+ $X2=4.015 $Y2=2.045
r224 61 63 7.64049 $w=1.7e-07 $l=1.94921e-07 $layer=LI1_cond $X=4.825 $Y=2.045
+ $X2=4.982 $Y2=1.96
r225 61 62 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=4.825 $Y=2.045
+ $X2=4.18 $Y2=2.045
r226 60 68 3.70735 $w=2.5e-07 $l=1.12916e-07 $layer=LI1_cond $X=3.95 $Y=1.96
+ $X2=4.015 $Y2=2.045
r227 60 72 62.3048 $w=1.68e-07 $l=9.55e-07 $layer=LI1_cond $X=3.95 $Y=1.96
+ $X2=3.95 $Y2=1.005
r228 55 57 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=4.015 $Y=2.19
+ $X2=4.015 $Y2=2.9
r229 53 68 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.015 $Y=2.13
+ $X2=4.015 $Y2=2.045
r230 53 55 2.09535 $w=3.28e-07 $l=6e-08 $layer=LI1_cond $X=4.015 $Y=2.13
+ $X2=4.015 $Y2=2.19
r231 47 49 346.117 $w=1.5e-07 $l=6.75e-07 $layer=POLY_cond $X=10.785 $Y=1.215
+ $X2=10.785 $Y2=0.54
r232 46 49 146.138 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=10.785 $Y=0.255
+ $X2=10.785 $Y2=0.54
r233 44 47 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=10.71 $Y=1.29
+ $X2=10.785 $Y2=1.215
r234 44 45 105.117 $w=1.5e-07 $l=2.05e-07 $layer=POLY_cond $X=10.71 $Y=1.29
+ $X2=10.505 $Y2=1.29
r235 42 45 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=10.43 $Y=1.365
+ $X2=10.505 $Y2=1.29
r236 42 43 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=10.43 $Y=1.365
+ $X2=10.43 $Y2=1.725
r237 40 43 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=10.355 $Y=1.8
+ $X2=10.43 $Y2=1.725
r238 40 41 133.319 $w=1.5e-07 $l=2.6e-07 $layer=POLY_cond $X=10.355 $Y=1.8
+ $X2=10.095 $Y2=1.8
r239 36 41 29.1797 $w=1.5e-07 $l=1.58114e-07 $layer=POLY_cond $X=9.97 $Y=1.875
+ $X2=10.095 $Y2=1.8
r240 36 38 178.887 $w=2.5e-07 $l=7.2e-07 $layer=POLY_cond $X=9.97 $Y=1.875
+ $X2=9.97 $Y2=2.595
r241 33 35 110.86 $w=2.5e-07 $l=5.75e-07 $layer=POLY_cond $X=6.74 $Y=2.02
+ $X2=6.74 $Y2=2.595
r242 31 46 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=10.71 $Y=0.18
+ $X2=10.785 $Y2=0.255
r243 31 32 2212.59 $w=1.5e-07 $l=4.315e-06 $layer=POLY_cond $X=10.71 $Y=0.18
+ $X2=6.395 $Y2=0.18
r244 29 33 29.1797 $w=1.5e-07 $l=1.58114e-07 $layer=POLY_cond $X=6.615 $Y=1.945
+ $X2=6.74 $Y2=2.02
r245 29 30 128.191 $w=1.5e-07 $l=2.5e-07 $layer=POLY_cond $X=6.615 $Y=1.945
+ $X2=6.365 $Y2=1.945
r246 26 52 66.2216 $w=1.65e-07 $l=2.32379e-07 $layer=POLY_cond $X=6.32 $Y=0.91
+ $X2=6.305 $Y2=1.135
r247 26 28 146.138 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=6.32 $Y=0.91
+ $X2=6.32 $Y2=0.625
r248 25 32 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.32 $Y=0.255
+ $X2=6.395 $Y2=0.18
r249 25 28 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=6.32 $Y=0.255
+ $X2=6.32 $Y2=0.625
r250 24 30 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.29 $Y=1.87
+ $X2=6.365 $Y2=1.945
r251 23 52 22.4034 $w=1.65e-07 $l=8.21584e-08 $layer=POLY_cond $X=6.29 $Y=1.21
+ $X2=6.305 $Y2=1.135
r252 23 24 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=6.29 $Y=1.21
+ $X2=6.29 $Y2=1.87
r253 22 51 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.39 $Y=1.135
+ $X2=5.315 $Y2=1.135
r254 21 52 5.10115 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=6.215 $Y=1.135
+ $X2=6.305 $Y2=1.135
r255 21 22 423.032 $w=1.5e-07 $l=8.25e-07 $layer=POLY_cond $X=6.215 $Y=1.135
+ $X2=5.39 $Y2=1.135
r256 18 51 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.315 $Y=1.06
+ $X2=5.315 $Y2=1.135
r257 18 20 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=5.315 $Y=1.06
+ $X2=5.315 $Y2=0.775
r258 17 50 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.03 $Y=1.135
+ $X2=4.955 $Y2=1.135
r259 16 51 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.24 $Y=1.135
+ $X2=5.315 $Y2=1.135
r260 16 17 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=5.24 $Y=1.135
+ $X2=5.03 $Y2=1.135
r261 15 75 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.955 $Y=1.555
+ $X2=4.955 $Y2=1.72
r262 14 50 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.955 $Y=1.21
+ $X2=4.955 $Y2=1.135
r263 14 15 176.904 $w=1.5e-07 $l=3.45e-07 $layer=POLY_cond $X=4.955 $Y=1.21
+ $X2=4.955 $Y2=1.555
r264 11 50 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.955 $Y=1.06
+ $X2=4.955 $Y2=1.135
r265 11 13 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=4.955 $Y=1.06
+ $X2=4.955 $Y2=0.775
r266 7 73 9.34494 $w=2.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.81 $Y=1.885
+ $X2=4.81 $Y2=1.72
r267 7 9 163.979 $w=2.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.81 $Y=1.885
+ $X2=4.81 $Y2=2.545
r268 2 57 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=3.87
+ $Y=2.045 $X2=4.015 $Y2=2.9
r269 2 55 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=3.87
+ $Y=2.045 $X2=4.015 $Y2=2.19
r270 1 70 182 $w=1.7e-07 $l=3.09112e-07 $layer=licon1_NDIFF $count=1 $X=3.805
+ $Y=0.565 $X2=3.95 $Y2=0.81
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSBP_LP%A_2220_40# 1 2 9 11 13 17 20 21 24 31 34
+ 35
c87 13 0 2.10017e-19 $X=11.41 $Y=2.595
c88 11 0 2.21142e-20 $X=11.41 $Y=1.885
r89 34 35 8.55446 $w=3.73e-07 $l=1.65e-07 $layer=LI1_cond $X=12.827 $Y=2.185
+ $X2=12.827 $Y2=2.02
r90 26 31 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=12.725 $Y=1.37
+ $X2=12.725 $Y2=1.285
r91 26 35 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=12.725 $Y=1.37
+ $X2=12.725 $Y2=2.02
r92 22 31 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=12.33 $Y=1.285
+ $X2=12.725 $Y2=1.285
r93 22 24 24.6204 $w=3.28e-07 $l=7.05e-07 $layer=LI1_cond $X=12.33 $Y=1.2
+ $X2=12.33 $Y2=0.495
r94 20 22 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=12.165 $Y=1.285
+ $X2=12.33 $Y2=1.285
r95 20 21 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=12.165 $Y=1.285
+ $X2=11.775 $Y2=1.285
r96 17 18 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=11.61
+ $Y=1.38 $X2=11.61 $Y2=1.38
r97 15 21 7.24806 $w=1.7e-07 $l=1.70276e-07 $layer=LI1_cond $X=11.642 $Y=1.37
+ $X2=11.775 $Y2=1.285
r98 15 17 0.434884 $w=2.63e-07 $l=1e-08 $layer=LI1_cond $X=11.642 $Y=1.37
+ $X2=11.642 $Y2=1.38
r99 11 18 58.6276 $w=5.54e-07 $l=5.18324e-07 $layer=POLY_cond $X=11.41 $Y=1.885
+ $X2=11.437 $Y2=1.38
r100 11 13 176.402 $w=2.5e-07 $l=7.1e-07 $layer=POLY_cond $X=11.41 $Y=1.885
+ $X2=11.41 $Y2=2.595
r101 7 18 43.3485 $w=5.54e-07 $l=3.34476e-07 $layer=POLY_cond $X=11.175 $Y=1.215
+ $X2=11.437 $Y2=1.38
r102 7 9 346.117 $w=1.5e-07 $l=6.75e-07 $layer=POLY_cond $X=11.175 $Y=1.215
+ $X2=11.175 $Y2=0.54
r103 2 34 300 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_PDIFF $count=2 $X=12.79
+ $Y=2 $X2=12.93 $Y2=2.185
r104 1 24 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=12.185
+ $Y=0.285 $X2=12.33 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSBP_LP%A_2019_419# 1 2 3 12 14 15 18 22 24 26 27
+ 29 30 31 33 34 36 38 40 42 45 47 49 51 53 59 65 67 69 70 72 73 75 76 77 78 81
+ 82 85 87 88 91
c210 75 0 1.64566e-19 $X=12.335 $Y=2.285
c211 72 0 8.27582e-20 $X=11.245 $Y=2.115
c212 70 0 1.65443e-19 $X=10.655 $Y=1.035
c213 59 0 3.36421e-19 $X=15.04 $Y=0.94
r214 85 91 68.8289 $w=1.68e-07 $l=1.055e-06 $layer=LI1_cond $X=13.28 $Y=2.895
+ $X2=13.28 $Y2=1.84
r215 81 82 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=13.155
+ $Y=1.335 $X2=13.155 $Y2=1.335
r216 79 91 9.23056 $w=3.73e-07 $l=1.87e-07 $layer=LI1_cond $X=13.177 $Y=1.653
+ $X2=13.177 $Y2=1.84
r217 79 81 9.77272 $w=3.73e-07 $l=3.18e-07 $layer=LI1_cond $X=13.177 $Y=1.653
+ $X2=13.177 $Y2=1.335
r218 77 85 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=13.195 $Y=2.98
+ $X2=13.28 $Y2=2.895
r219 77 78 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=13.195 $Y=2.98
+ $X2=12.46 $Y2=2.98
r220 76 78 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=12.335 $Y=2.895
+ $X2=12.46 $Y2=2.98
r221 75 90 3.00013 $w=2.5e-07 $l=1.05e-07 $layer=LI1_cond $X=12.335 $Y=2.285
+ $X2=12.335 $Y2=2.18
r222 75 76 28.1196 $w=2.48e-07 $l=6.1e-07 $layer=LI1_cond $X=12.335 $Y=2.285
+ $X2=12.335 $Y2=2.895
r223 74 88 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.33 $Y=2.2
+ $X2=11.245 $Y2=2.2
r224 73 90 4.14303 $w=1.7e-07 $l=1.34629e-07 $layer=LI1_cond $X=12.21 $Y=2.2
+ $X2=12.335 $Y2=2.18
r225 73 74 57.4118 $w=1.68e-07 $l=8.8e-07 $layer=LI1_cond $X=12.21 $Y=2.2
+ $X2=11.33 $Y2=2.2
r226 72 88 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.245 $Y=2.115
+ $X2=11.245 $Y2=2.2
r227 71 72 64.9144 $w=1.68e-07 $l=9.95e-07 $layer=LI1_cond $X=11.245 $Y=1.12
+ $X2=11.245 $Y2=2.115
r228 69 71 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=11.16 $Y=1.035
+ $X2=11.245 $Y2=1.12
r229 69 70 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=11.16 $Y=1.035
+ $X2=10.655 $Y2=1.035
r230 68 87 4.95428 $w=1.7e-07 $l=1.74714e-07 $layer=LI1_cond $X=10.535 $Y=2.2
+ $X2=10.37 $Y2=2.18
r231 67 88 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.16 $Y=2.2
+ $X2=11.245 $Y2=2.2
r232 67 68 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=11.16 $Y=2.2
+ $X2=10.535 $Y2=2.2
r233 63 70 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=10.49 $Y=0.95
+ $X2=10.655 $Y2=1.035
r234 63 65 16.5882 $w=3.28e-07 $l=4.75e-07 $layer=LI1_cond $X=10.49 $Y=0.95
+ $X2=10.49 $Y2=0.475
r235 55 56 40.8361 $w=3.6e-07 $l=3.05e-07 $layer=POLY_cond $X=13.82 $Y=0.94
+ $X2=13.82 $Y2=1.245
r236 52 82 28.3893 $w=4.9e-07 $l=2.6e-07 $layer=POLY_cond $X=13.075 $Y=1.595
+ $X2=13.075 $Y2=1.335
r237 52 53 39.5539 $w=4.9e-07 $l=2.45e-07 $layer=POLY_cond $X=13.075 $Y=1.595
+ $X2=13.075 $Y2=1.84
r238 50 82 1.63785 $w=4.9e-07 $l=1.5e-08 $layer=POLY_cond $X=13.075 $Y=1.32
+ $X2=13.075 $Y2=1.335
r239 50 51 4.35086 $w=4.9e-07 $l=7.5e-08 $layer=POLY_cond $X=13.075 $Y=1.32
+ $X2=13.075 $Y2=1.245
r240 47 59 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=15.04 $Y=0.865
+ $X2=15.04 $Y2=0.94
r241 47 49 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=15.04 $Y=0.865
+ $X2=15.04 $Y2=0.58
r242 43 59 28.2021 $w=1.5e-07 $l=5.5e-08 $layer=POLY_cond $X=14.985 $Y=0.94
+ $X2=15.04 $Y2=0.94
r243 43 57 156.394 $w=1.5e-07 $l=3.05e-07 $layer=POLY_cond $X=14.985 $Y=0.94
+ $X2=14.68 $Y2=0.94
r244 43 45 336.655 $w=2.5e-07 $l=1.355e-06 $layer=POLY_cond $X=14.985 $Y=1.015
+ $X2=14.985 $Y2=2.37
r245 40 57 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=14.68 $Y=0.865
+ $X2=14.68 $Y2=0.94
r246 40 42 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=14.68 $Y=0.865
+ $X2=14.68 $Y2=0.58
r247 39 55 23.3057 $w=1.5e-07 $l=2e-07 $layer=POLY_cond $X=14.02 $Y=0.94
+ $X2=13.82 $Y2=0.94
r248 38 57 38.4574 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=14.605 $Y=0.94
+ $X2=14.68 $Y2=0.94
r249 38 39 299.968 $w=1.5e-07 $l=5.85e-07 $layer=POLY_cond $X=14.605 $Y=0.94
+ $X2=14.02 $Y2=0.94
r250 34 56 14.5895 $w=3.6e-07 $l=1.06066e-07 $layer=POLY_cond $X=13.895 $Y=1.32
+ $X2=13.82 $Y2=1.245
r251 34 36 293.175 $w=2.5e-07 $l=1.18e-06 $layer=POLY_cond $X=13.895 $Y=1.32
+ $X2=13.895 $Y2=2.5
r252 31 33 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=13.695 $Y=0.78
+ $X2=13.695 $Y2=0.495
r253 29 55 11.3806 $w=3.6e-07 $l=2.38747e-07 $layer=POLY_cond $X=13.62 $Y=0.855
+ $X2=13.82 $Y2=0.94
r254 29 31 26.8603 $w=3.6e-07 $l=1.06066e-07 $layer=POLY_cond $X=13.62 $Y=0.855
+ $X2=13.695 $Y2=0.78
r255 29 30 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=13.62 $Y=0.855
+ $X2=13.41 $Y2=0.855
r256 28 51 22.1783 $w=1.5e-07 $l=2.45e-07 $layer=POLY_cond $X=13.32 $Y=1.245
+ $X2=13.075 $Y2=1.245
r257 27 56 23.3057 $w=1.5e-07 $l=2e-07 $layer=POLY_cond $X=13.62 $Y=1.245
+ $X2=13.82 $Y2=1.245
r258 27 28 153.83 $w=1.5e-07 $l=3e-07 $layer=POLY_cond $X=13.62 $Y=1.245
+ $X2=13.32 $Y2=1.245
r259 24 30 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=13.335 $Y=0.78
+ $X2=13.41 $Y2=0.855
r260 24 26 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=13.335 $Y=0.78
+ $X2=13.335 $Y2=0.495
r261 22 53 163.979 $w=2.5e-07 $l=6.6e-07 $layer=POLY_cond $X=13.195 $Y=2.5
+ $X2=13.195 $Y2=1.84
r262 16 51 4.35086 $w=1.5e-07 $l=2.04083e-07 $layer=POLY_cond $X=12.905 $Y=1.17
+ $X2=13.075 $Y2=1.245
r263 16 18 346.117 $w=1.5e-07 $l=6.75e-07 $layer=POLY_cond $X=12.905 $Y=1.17
+ $X2=12.905 $Y2=0.495
r264 14 51 22.1783 $w=1.5e-07 $l=2.45e-07 $layer=POLY_cond $X=12.83 $Y=1.245
+ $X2=13.075 $Y2=1.245
r265 14 15 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=12.83 $Y=1.245
+ $X2=12.62 $Y2=1.245
r266 10 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=12.545 $Y=1.17
+ $X2=12.62 $Y2=1.245
r267 10 12 346.117 $w=1.5e-07 $l=6.75e-07 $layer=POLY_cond $X=12.545 $Y=1.17
+ $X2=12.545 $Y2=0.495
r268 3 90 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=12.235
+ $Y=2.095 $X2=12.375 $Y2=2.24
r269 2 87 300 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=2 $X=10.095
+ $Y=2.095 $X2=10.37 $Y2=2.24
r270 1 65 91 $w=1.7e-07 $l=4.43706e-07 $layer=licon1_NDIFF $count=2 $X=10.115
+ $Y=0.625 $X2=10.49 $Y2=0.475
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSBP_LP%A_2865_74# 1 2 7 9 12 16 18 23 26 29 33 37
+ 38 41 44
c69 44 0 7.8944e-20 $X=14.672 $Y=1.575
c70 37 0 1.85811e-19 $X=15.56 $Y=1.155
c71 33 0 1.5061e-19 $X=15.395 $Y=1.575
r72 41 43 10.7321 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=14.465 $Y=0.58
+ $X2=14.465 $Y2=0.81
r73 37 38 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=15.56
+ $Y=1.155 $X2=15.56 $Y2=1.155
r74 35 37 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=15.56 $Y=1.49
+ $X2=15.56 $Y2=1.155
r75 34 44 3.41642 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=14.885 $Y=1.575
+ $X2=14.672 $Y2=1.575
r76 33 35 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=15.395 $Y=1.575
+ $X2=15.56 $Y2=1.49
r77 33 34 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=15.395 $Y=1.575
+ $X2=14.885 $Y2=1.575
r78 29 31 19.2526 $w=4.23e-07 $l=7.1e-07 $layer=LI1_cond $X=14.672 $Y=2.015
+ $X2=14.672 $Y2=2.725
r79 27 44 3.17288 $w=2.97e-07 $l=8.5e-08 $layer=LI1_cond $X=14.672 $Y=1.66
+ $X2=14.672 $Y2=1.575
r80 27 29 9.62629 $w=4.23e-07 $l=3.55e-07 $layer=LI1_cond $X=14.672 $Y=1.66
+ $X2=14.672 $Y2=2.015
r81 26 44 3.17288 $w=2.97e-07 $l=1.64085e-07 $layer=LI1_cond $X=14.545 $Y=1.49
+ $X2=14.672 $Y2=1.575
r82 26 43 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=14.545 $Y=1.49
+ $X2=14.545 $Y2=0.81
r83 22 38 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=15.56 $Y=1.14
+ $X2=15.56 $Y2=1.155
r84 22 23 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=15.56 $Y=1.065
+ $X2=15.83 $Y2=1.065
r85 19 22 46.1489 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=15.47 $Y=1.065
+ $X2=15.56 $Y2=1.065
r86 18 38 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=15.56 $Y=1.495
+ $X2=15.56 $Y2=1.155
r87 14 23 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=15.83 $Y=0.99
+ $X2=15.83 $Y2=1.065
r88 14 16 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=15.83 $Y=0.99
+ $X2=15.83 $Y2=0.58
r89 10 19 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=15.47 $Y=0.99
+ $X2=15.47 $Y2=1.065
r90 10 12 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=15.47 $Y=0.99
+ $X2=15.47 $Y2=0.58
r91 7 18 47.383 $w=2.95e-07 $l=3.11689e-07 $layer=POLY_cond $X=15.515 $Y=1.785
+ $X2=15.56 $Y2=1.495
r92 7 9 112.788 $w=2.5e-07 $l=5.85e-07 $layer=POLY_cond $X=15.515 $Y=1.785
+ $X2=15.515 $Y2=2.37
r93 2 31 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=14.575
+ $Y=1.87 $X2=14.72 $Y2=2.725
r94 2 29 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=14.575
+ $Y=1.87 $X2=14.72 $Y2=2.015
r95 1 41 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=14.325
+ $Y=0.37 $X2=14.465 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSBP_LP%VPWR 1 2 3 4 5 6 7 8 29 35 39 43 45 49 53
+ 57 63 68 69 70 79 86 94 102 107 114 115 118 121 124 127 130 133 136
r169 136 137 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=15.12 $Y=3.33
+ $X2=15.12 $Y2=3.33
r170 133 134 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.68 $Y=3.33
+ $X2=13.68 $Y2=3.33
r171 130 131 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.76 $Y=3.33
+ $X2=11.76 $Y2=3.33
r172 127 128 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r173 124 125 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r174 121 122 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r175 118 119 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r176 115 137 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=16.08 $Y=3.33
+ $X2=15.12 $Y2=3.33
r177 114 115 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=16.08 $Y=3.33
+ $X2=16.08 $Y2=3.33
r178 112 136 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=15.415 $Y=3.33
+ $X2=15.25 $Y2=3.33
r179 112 114 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=15.415 $Y=3.33
+ $X2=16.08 $Y2=3.33
r180 111 137 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=14.16 $Y=3.33
+ $X2=15.12 $Y2=3.33
r181 111 134 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=14.16 $Y=3.33
+ $X2=13.68 $Y2=3.33
r182 110 111 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=14.16 $Y=3.33
+ $X2=14.16 $Y2=3.33
r183 108 133 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=13.795 $Y=3.33
+ $X2=13.67 $Y2=3.33
r184 108 110 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=13.795 $Y=3.33
+ $X2=14.16 $Y2=3.33
r185 107 136 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=15.085 $Y=3.33
+ $X2=15.25 $Y2=3.33
r186 107 110 60.3476 $w=1.68e-07 $l=9.25e-07 $layer=LI1_cond $X=15.085 $Y=3.33
+ $X2=14.16 $Y2=3.33
r187 106 134 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.2 $Y=3.33
+ $X2=13.68 $Y2=3.33
r188 106 131 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=13.2 $Y=3.33
+ $X2=11.76 $Y2=3.33
r189 105 106 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=13.2 $Y=3.33
+ $X2=13.2 $Y2=3.33
r190 103 130 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.84 $Y=3.33
+ $X2=11.675 $Y2=3.33
r191 103 105 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=11.84 $Y=3.33
+ $X2=13.2 $Y2=3.33
r192 102 133 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=13.545 $Y=3.33
+ $X2=13.67 $Y2=3.33
r193 102 105 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=13.545 $Y=3.33
+ $X2=13.2 $Y2=3.33
r194 101 131 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=3.33
+ $X2=11.76 $Y2=3.33
r195 100 101 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=11.28 $Y=3.33
+ $X2=11.28 $Y2=3.33
r196 98 101 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=11.28 $Y2=3.33
r197 98 128 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=8.88 $Y2=3.33
r198 97 100 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=9.36 $Y=3.33
+ $X2=11.28 $Y2=3.33
r199 97 98 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r200 95 127 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.13 $Y=3.33
+ $X2=8.965 $Y2=3.33
r201 95 97 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=9.13 $Y=3.33
+ $X2=9.36 $Y2=3.33
r202 94 130 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.51 $Y=3.33
+ $X2=11.675 $Y2=3.33
r203 94 100 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=11.51 $Y=3.33
+ $X2=11.28 $Y2=3.33
r204 93 125 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=7.92 $Y2=3.33
r205 92 93 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r206 90 93 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=7.44 $Y2=3.33
r207 90 122 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=4.56 $Y2=3.33
r208 89 92 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=5.04 $Y=3.33
+ $X2=7.44 $Y2=3.33
r209 89 90 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r210 87 121 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.71 $Y=3.33
+ $X2=4.545 $Y2=3.33
r211 87 89 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=4.71 $Y=3.33
+ $X2=5.04 $Y2=3.33
r212 86 124 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.74 $Y=3.33
+ $X2=7.905 $Y2=3.33
r213 86 92 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=7.74 $Y=3.33 $X2=7.44
+ $Y2=3.33
r214 85 122 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r215 84 85 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r216 82 85 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=4.08 $Y2=3.33
r217 81 84 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=3.12 $Y=3.33
+ $X2=4.08 $Y2=3.33
r218 81 82 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r219 79 121 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.38 $Y=3.33
+ $X2=4.545 $Y2=3.33
r220 79 84 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=4.38 $Y=3.33 $X2=4.08
+ $Y2=3.33
r221 78 82 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r222 77 78 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r223 75 78 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r224 75 119 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r225 74 77 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r226 74 75 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r227 72 118 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.975 $Y=3.33
+ $X2=0.81 $Y2=3.33
r228 72 74 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=0.975 $Y=3.33
+ $X2=1.2 $Y2=3.33
r229 70 128 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=8.16 $Y=3.33
+ $X2=8.88 $Y2=3.33
r230 70 125 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=8.16 $Y=3.33
+ $X2=7.92 $Y2=3.33
r231 68 77 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=2.755 $Y=3.33
+ $X2=2.64 $Y2=3.33
r232 68 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.755 $Y=3.33
+ $X2=2.92 $Y2=3.33
r233 67 81 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=3.085 $Y=3.33
+ $X2=3.12 $Y2=3.33
r234 67 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.085 $Y=3.33
+ $X2=2.92 $Y2=3.33
r235 63 66 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=15.25 $Y=2.015
+ $X2=15.25 $Y2=2.725
r236 61 136 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=15.25 $Y=3.245
+ $X2=15.25 $Y2=3.33
r237 61 66 18.1597 $w=3.28e-07 $l=5.2e-07 $layer=LI1_cond $X=15.25 $Y=3.245
+ $X2=15.25 $Y2=2.725
r238 57 60 32.7294 $w=2.48e-07 $l=7.1e-07 $layer=LI1_cond $X=13.67 $Y=2.145
+ $X2=13.67 $Y2=2.855
r239 55 133 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=13.67 $Y=3.245
+ $X2=13.67 $Y2=3.33
r240 55 60 17.9781 $w=2.48e-07 $l=3.9e-07 $layer=LI1_cond $X=13.67 $Y=3.245
+ $X2=13.67 $Y2=2.855
r241 51 130 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=11.675 $Y=3.245
+ $X2=11.675 $Y2=3.33
r242 51 53 21.4773 $w=3.28e-07 $l=6.15e-07 $layer=LI1_cond $X=11.675 $Y=3.245
+ $X2=11.675 $Y2=2.63
r243 47 127 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.965 $Y=3.245
+ $X2=8.965 $Y2=3.33
r244 47 49 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=8.965 $Y=3.245
+ $X2=8.965 $Y2=2.95
r245 46 124 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.07 $Y=3.33
+ $X2=7.905 $Y2=3.33
r246 45 127 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.8 $Y=3.33
+ $X2=8.965 $Y2=3.33
r247 45 46 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=8.8 $Y=3.33
+ $X2=8.07 $Y2=3.33
r248 41 124 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.905 $Y=3.245
+ $X2=7.905 $Y2=3.33
r249 41 43 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=7.905 $Y=3.245
+ $X2=7.905 $Y2=2.95
r250 37 121 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.545 $Y=3.245
+ $X2=4.545 $Y2=3.33
r251 37 39 26.8903 $w=3.28e-07 $l=7.7e-07 $layer=LI1_cond $X=4.545 $Y=3.245
+ $X2=4.545 $Y2=2.475
r252 33 69 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.92 $Y=3.245
+ $X2=2.92 $Y2=3.33
r253 33 35 13.2706 $w=3.28e-07 $l=3.8e-07 $layer=LI1_cond $X=2.92 $Y=3.245
+ $X2=2.92 $Y2=2.865
r254 29 32 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=0.81 $Y=2.19
+ $X2=0.81 $Y2=2.9
r255 27 118 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.81 $Y=3.245
+ $X2=0.81 $Y2=3.33
r256 27 32 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=0.81 $Y=3.245
+ $X2=0.81 $Y2=2.9
r257 8 66 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=15.11
+ $Y=1.87 $X2=15.25 $Y2=2.725
r258 8 63 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=15.11
+ $Y=1.87 $X2=15.25 $Y2=2.015
r259 7 60 400 $w=1.7e-07 $l=9.98036e-07 $layer=licon1_PDIFF $count=1 $X=13.32
+ $Y=2 $X2=13.63 $Y2=2.855
r260 7 57 400 $w=1.7e-07 $l=3.75566e-07 $layer=licon1_PDIFF $count=1 $X=13.32
+ $Y=2 $X2=13.63 $Y2=2.145
r261 6 53 300 $w=1.7e-07 $l=6.00937e-07 $layer=licon1_PDIFF $count=2 $X=11.535
+ $Y=2.095 $X2=11.675 $Y2=2.63
r262 5 49 600 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=8.825
+ $Y=2.095 $X2=8.965 $Y2=2.95
r263 4 43 600 $w=1.7e-07 $l=1.08031e-06 $layer=licon1_PDIFF $count=1 $X=7.395
+ $Y=2.095 $X2=7.905 $Y2=2.95
r264 3 39 300 $w=1.7e-07 $l=4.95076e-07 $layer=licon1_PDIFF $count=2 $X=4.405
+ $Y=2.045 $X2=4.545 $Y2=2.475
r265 2 35 600 $w=1.7e-07 $l=8.87243e-07 $layer=licon1_PDIFF $count=1 $X=2.78
+ $Y=2.045 $X2=2.92 $Y2=2.865
r266 1 32 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=0.67
+ $Y=2.045 $X2=0.81 $Y2=2.9
r267 1 29 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.67
+ $Y=2.045 $X2=0.81 $Y2=2.19
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSBP_LP%A_245_409# 1 2 7 9 11 14 15 16 22
c52 11 0 4.76528e-20 $X=2.405 $Y=2.98
r53 15 22 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.285 $Y=2.405
+ $X2=3.45 $Y2=2.405
r54 15 16 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=3.285 $Y=2.405
+ $X2=2.575 $Y2=2.405
r55 13 16 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.49 $Y=2.49
+ $X2=2.575 $Y2=2.405
r56 13 14 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=2.49 $Y=2.49
+ $X2=2.49 $Y2=2.895
r57 12 20 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.535 $Y=2.98
+ $X2=1.37 $Y2=2.98
r58 11 14 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.405 $Y=2.98
+ $X2=2.49 $Y2=2.895
r59 11 12 56.7594 $w=1.68e-07 $l=8.7e-07 $layer=LI1_cond $X=2.405 $Y=2.98
+ $X2=1.535 $Y2=2.98
r60 7 20 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.37 $Y=2.895 $X2=1.37
+ $Y2=2.98
r61 7 9 24.6204 $w=3.28e-07 $l=7.05e-07 $layer=LI1_cond $X=1.37 $Y=2.895
+ $X2=1.37 $Y2=2.19
r62 2 22 300 $w=1.7e-07 $l=5.05173e-07 $layer=licon1_PDIFF $count=2 $X=3.31
+ $Y=2.045 $X2=3.45 $Y2=2.485
r63 1 20 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=1.225
+ $Y=2.045 $X2=1.37 $Y2=2.9
r64 1 9 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=1.225
+ $Y=2.045 $X2=1.37 $Y2=2.19
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSBP_LP%A_352_409# 1 2 3 4 15 17 18 19 22 23 26 27
+ 28 30 31 32 34 35 36 41 45 48 50 51 53 54
c181 51 0 1.55371e-19 $X=5.1 $Y=1.227
c182 27 0 1.86498e-19 $X=4.295 $Y=0.35
r183 53 54 8.63679 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=5.55 $Y=1.96
+ $X2=5.55 $Y2=2.13
r184 51 52 18.605 $w=2e-07 $l=3.05e-07 $layer=LI1_cond $X=5.1 $Y=1.227 $X2=5.405
+ $Y2=1.227
r185 43 45 8.75857 $w=2.48e-07 $l=1.9e-07 $layer=LI1_cond $X=6.145 $Y=0.435
+ $X2=6.145 $Y2=0.625
r186 41 54 9.25447 $w=3.28e-07 $l=2.65e-07 $layer=LI1_cond $X=5.615 $Y=2.395
+ $X2=5.615 $Y2=2.13
r187 37 52 1.68994 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=5.405 $Y=1.355
+ $X2=5.405 $Y2=1.227
r188 37 53 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=5.405 $Y=1.355
+ $X2=5.405 $Y2=1.96
r189 35 43 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=6.02 $Y=0.35
+ $X2=6.145 $Y2=0.435
r190 35 36 54.4759 $w=1.68e-07 $l=8.35e-07 $layer=LI1_cond $X=6.02 $Y=0.35
+ $X2=5.185 $Y2=0.35
r191 34 51 1.68994 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=5.1 $Y=1.1 $X2=5.1
+ $Y2=1.227
r192 33 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.1 $Y=0.435
+ $X2=5.185 $Y2=0.35
r193 33 34 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=5.1 $Y=0.435
+ $X2=5.1 $Y2=1.1
r194 31 51 5.49448 $w=2e-07 $l=1.03899e-07 $layer=LI1_cond $X=5.015 $Y=1.185
+ $X2=5.1 $Y2=1.227
r195 31 32 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=5.015 $Y=1.185
+ $X2=4.465 $Y2=1.185
r196 30 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.38 $Y=1.1
+ $X2=4.465 $Y2=1.185
r197 29 30 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=4.38 $Y=0.435
+ $X2=4.38 $Y2=1.1
r198 27 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.295 $Y=0.35
+ $X2=4.38 $Y2=0.435
r199 27 28 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=4.295 $Y=0.35
+ $X2=3.675 $Y2=0.35
r200 25 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.59 $Y=0.435
+ $X2=3.675 $Y2=0.35
r201 25 26 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=3.59 $Y=0.435
+ $X2=3.59 $Y2=0.76
r202 24 50 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.185 $Y=0.845
+ $X2=3.1 $Y2=0.845
r203 23 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.505 $Y=0.845
+ $X2=3.59 $Y2=0.76
r204 23 24 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=3.505 $Y=0.845
+ $X2=3.185 $Y2=0.845
r205 21 50 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.1 $Y=0.93 $X2=3.1
+ $Y2=0.845
r206 21 22 67.8503 $w=1.68e-07 $l=1.04e-06 $layer=LI1_cond $X=3.1 $Y=0.93
+ $X2=3.1 $Y2=1.97
r207 20 48 15.1084 $w=3.23e-07 $l=5e-07 $layer=LI1_cond $X=2.625 $Y=0.845
+ $X2=2.4 $Y2=0.445
r208 19 50 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.015 $Y=0.845
+ $X2=3.1 $Y2=0.845
r209 19 20 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=3.015 $Y=0.845
+ $X2=2.625 $Y2=0.845
r210 17 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.015 $Y=2.055
+ $X2=3.1 $Y2=1.97
r211 17 18 61.9786 $w=1.68e-07 $l=9.5e-07 $layer=LI1_cond $X=3.015 $Y=2.055
+ $X2=2.065 $Y2=2.055
r212 13 18 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.9 $Y=2.14
+ $X2=2.065 $Y2=2.055
r213 13 15 1.74613 $w=3.28e-07 $l=5e-08 $layer=LI1_cond $X=1.9 $Y=2.14 $X2=1.9
+ $Y2=2.19
r214 4 41 600 $w=1.7e-07 $l=3.61248e-07 $layer=licon1_PDIFF $count=1 $X=5.48
+ $Y=2.095 $X2=5.615 $Y2=2.395
r215 3 15 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=1.76
+ $Y=2.045 $X2=1.9 $Y2=2.19
r216 2 45 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=5.96
+ $Y=0.415 $X2=6.105 $Y2=0.625
r217 1 48 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.2
+ $Y=0.235 $X2=2.34 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSBP_LP%Q_N 1 2 7 11 15 16 17 18 25 32
r43 18 25 2.9826 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=13.68 $Y=1.695
+ $X2=13.68 $Y2=1.61
r44 18 25 0.751593 $w=2.28e-07 $l=1.5e-08 $layer=LI1_cond $X=13.68 $Y=1.595
+ $X2=13.68 $Y2=1.61
r45 17 18 15.0319 $w=2.28e-07 $l=3e-07 $layer=LI1_cond $X=13.68 $Y=1.295
+ $X2=13.68 $Y2=1.595
r46 16 17 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=13.68 $Y=0.925
+ $X2=13.68 $Y2=1.295
r47 16 36 10.0212 $w=2.28e-07 $l=2e-07 $layer=LI1_cond $X=13.68 $Y=0.925
+ $X2=13.68 $Y2=0.725
r48 15 36 7.63653 $w=5.08e-07 $l=1.7e-07 $layer=LI1_cond $X=13.82 $Y=0.555
+ $X2=13.82 $Y2=0.725
r49 15 32 1.40715 $w=5.08e-07 $l=6e-08 $layer=LI1_cond $X=13.82 $Y=0.555
+ $X2=13.82 $Y2=0.495
r50 11 13 32.7294 $w=2.48e-07 $l=7.1e-07 $layer=LI1_cond $X=14.12 $Y=2.145
+ $X2=14.12 $Y2=2.855
r51 9 11 16.8257 $w=2.48e-07 $l=3.65e-07 $layer=LI1_cond $X=14.12 $Y=1.78
+ $X2=14.12 $Y2=2.145
r52 8 18 4.03528 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=13.795 $Y=1.695
+ $X2=13.68 $Y2=1.695
r53 7 9 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=13.995 $Y=1.695
+ $X2=14.12 $Y2=1.78
r54 7 8 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=13.995 $Y=1.695
+ $X2=13.795 $Y2=1.695
r55 2 13 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=14.02
+ $Y=2 $X2=14.16 $Y2=2.855
r56 2 11 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=14.02
+ $Y=2 $X2=14.16 $Y2=2.145
r57 1 32 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=13.77
+ $Y=0.285 $X2=13.91 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSBP_LP%Q 1 2 10 13 14 15 28 29
r23 28 29 10.1235 $w=5.93e-07 $l=1.65e-07 $layer=LI1_cond $X=15.912 $Y=2.015
+ $X2=15.912 $Y2=1.85
r24 15 23 1.00511 $w=5.93e-07 $l=5e-08 $layer=LI1_cond $X=15.912 $Y=2.775
+ $X2=15.912 $Y2=2.725
r25 14 23 6.43269 $w=5.93e-07 $l=3.2e-07 $layer=LI1_cond $X=15.912 $Y=2.405
+ $X2=15.912 $Y2=2.725
r26 14 19 5.18636 $w=5.93e-07 $l=2.58e-07 $layer=LI1_cond $X=15.912 $Y=2.405
+ $X2=15.912 $Y2=2.147
r27 13 19 2.25144 $w=5.93e-07 $l=1.12e-07 $layer=LI1_cond $X=15.912 $Y=2.035
+ $X2=15.912 $Y2=2.147
r28 13 28 0.402043 $w=5.93e-07 $l=2e-08 $layer=LI1_cond $X=15.912 $Y=2.035
+ $X2=15.912 $Y2=2.015
r29 12 29 67.8503 $w=1.68e-07 $l=1.04e-06 $layer=LI1_cond $X=16.125 $Y=0.81
+ $X2=16.125 $Y2=1.85
r30 10 12 10.7321 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=16.045 $Y=0.58
+ $X2=16.045 $Y2=0.81
r31 2 28 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=15.64
+ $Y=1.87 $X2=15.78 $Y2=2.015
r32 2 23 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=15.64
+ $Y=1.87 $X2=15.78 $Y2=2.725
r33 1 10 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=15.905
+ $Y=0.37 $X2=16.045 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSBP_LP%VGND 1 2 3 4 5 6 7 8 27 31 35 39 43 47 51
+ 55 58 59 60 62 67 82 89 97 102 107 114 115 118 121 124 127 130 133 136
c181 47 0 2.21142e-20 $X=11.755 $Y=0.54
r182 136 137 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=15.12 $Y=0
+ $X2=15.12 $Y2=0
r183 133 134 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.2 $Y=0
+ $X2=13.2 $Y2=0
r184 130 131 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.76 $Y=0
+ $X2=11.76 $Y2=0
r185 127 128 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=9.36 $Y=0
+ $X2=9.36 $Y2=0
r186 124 125 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=0
+ $X2=7.44 $Y2=0
r187 121 122 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0
+ $X2=3.12 $Y2=0
r188 118 119 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r189 115 137 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=16.08 $Y=0
+ $X2=15.12 $Y2=0
r190 114 115 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=16.08 $Y=0
+ $X2=16.08 $Y2=0
r191 112 136 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=15.42 $Y=0
+ $X2=15.255 $Y2=0
r192 112 114 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=15.42 $Y=0
+ $X2=16.08 $Y2=0
r193 111 137 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=13.68 $Y=0
+ $X2=15.12 $Y2=0
r194 111 134 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.68 $Y=0
+ $X2=13.2 $Y2=0
r195 110 111 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=13.68 $Y=0
+ $X2=13.68 $Y2=0
r196 108 133 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.285 $Y=0
+ $X2=13.12 $Y2=0
r197 108 110 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=13.285 $Y=0
+ $X2=13.68 $Y2=0
r198 107 136 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=15.09 $Y=0
+ $X2=15.255 $Y2=0
r199 107 110 91.9893 $w=1.68e-07 $l=1.41e-06 $layer=LI1_cond $X=15.09 $Y=0
+ $X2=13.68 $Y2=0
r200 106 134 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.72 $Y=0
+ $X2=13.2 $Y2=0
r201 106 131 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=12.72 $Y=0
+ $X2=11.76 $Y2=0
r202 105 106 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=12.72 $Y=0
+ $X2=12.72 $Y2=0
r203 103 130 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.92 $Y=0
+ $X2=11.755 $Y2=0
r204 103 105 52.1925 $w=1.68e-07 $l=8e-07 $layer=LI1_cond $X=11.92 $Y=0
+ $X2=12.72 $Y2=0
r205 102 133 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.955 $Y=0
+ $X2=13.12 $Y2=0
r206 102 105 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=12.955 $Y=0
+ $X2=12.72 $Y2=0
r207 101 131 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=0
+ $X2=11.76 $Y2=0
r208 101 128 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=11.28 $Y=0
+ $X2=9.36 $Y2=0
r209 100 101 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=11.28 $Y=0
+ $X2=11.28 $Y2=0
r210 98 127 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.38 $Y=0
+ $X2=9.215 $Y2=0
r211 98 100 123.957 $w=1.68e-07 $l=1.9e-06 $layer=LI1_cond $X=9.38 $Y=0
+ $X2=11.28 $Y2=0
r212 97 130 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.59 $Y=0
+ $X2=11.755 $Y2=0
r213 97 100 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=11.59 $Y=0
+ $X2=11.28 $Y2=0
r214 96 128 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=0
+ $X2=9.36 $Y2=0
r215 95 96 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.88 $Y=0 $X2=8.88
+ $Y2=0
r216 93 125 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0
+ $X2=7.44 $Y2=0
r217 92 95 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=7.92 $Y=0 $X2=8.88
+ $Y2=0
r218 92 93 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r219 90 124 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.565 $Y=0
+ $X2=7.44 $Y2=0
r220 90 92 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=7.565 $Y=0
+ $X2=7.92 $Y2=0
r221 89 127 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.05 $Y=0
+ $X2=9.215 $Y2=0
r222 89 95 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=9.05 $Y=0 $X2=8.88
+ $Y2=0
r223 88 125 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0
+ $X2=7.44 $Y2=0
r224 87 88 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.96 $Y=0
+ $X2=6.96 $Y2=0
r225 85 88 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=5.04 $Y=0
+ $X2=6.96 $Y2=0
r226 84 87 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=5.04 $Y=0 $X2=6.96
+ $Y2=0
r227 84 85 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.04 $Y=0
+ $X2=5.04 $Y2=0
r228 82 124 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.315 $Y=0
+ $X2=7.44 $Y2=0
r229 82 87 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=7.315 $Y=0
+ $X2=6.96 $Y2=0
r230 81 85 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.04
+ $Y2=0
r231 80 81 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r232 78 81 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.56
+ $Y2=0
r233 78 122 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=3.12
+ $Y2=0
r234 77 80 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=3.6 $Y=0 $X2=4.56
+ $Y2=0
r235 77 78 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r236 75 121 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.325 $Y=0
+ $X2=3.16 $Y2=0
r237 75 77 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=3.325 $Y=0 $X2=3.6
+ $Y2=0
r238 74 122 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0
+ $X2=3.12 $Y2=0
r239 73 74 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r240 71 74 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r241 71 119 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r242 70 73 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r243 70 71 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r244 68 118 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.385 $Y=0
+ $X2=1.22 $Y2=0
r245 68 70 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.385 $Y=0 $X2=1.68
+ $Y2=0
r246 67 121 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.995 $Y=0
+ $X2=3.16 $Y2=0
r247 67 73 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=2.995 $Y=0
+ $X2=2.64 $Y2=0
r248 65 119 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r249 64 65 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r250 62 118 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.055 $Y=0
+ $X2=1.22 $Y2=0
r251 62 64 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.055 $Y=0
+ $X2=0.72 $Y2=0
r252 60 96 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=8.16 $Y=0 $X2=8.88
+ $Y2=0
r253 60 93 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=8.16 $Y=0
+ $X2=7.92 $Y2=0
r254 58 80 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=4.655 $Y=0 $X2=4.56
+ $Y2=0
r255 58 59 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.655 $Y=0 $X2=4.74
+ $Y2=0
r256 57 84 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=4.825 $Y=0
+ $X2=5.04 $Y2=0
r257 57 59 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.825 $Y=0 $X2=4.74
+ $Y2=0
r258 53 136 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=15.255 $Y=0.085
+ $X2=15.255 $Y2=0
r259 53 55 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=15.255 $Y=0.085
+ $X2=15.255 $Y2=0.58
r260 49 133 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=13.12 $Y=0.085
+ $X2=13.12 $Y2=0
r261 49 51 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=13.12 $Y=0.085
+ $X2=13.12 $Y2=0.495
r262 45 130 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=11.755 $Y=0.085
+ $X2=11.755 $Y2=0
r263 45 47 15.8897 $w=3.28e-07 $l=4.55e-07 $layer=LI1_cond $X=11.755 $Y=0.085
+ $X2=11.755 $Y2=0.54
r264 41 127 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.215 $Y=0.085
+ $X2=9.215 $Y2=0
r265 41 43 25.3188 $w=3.28e-07 $l=7.25e-07 $layer=LI1_cond $X=9.215 $Y=0.085
+ $X2=9.215 $Y2=0.81
r266 37 124 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.44 $Y=0.085
+ $X2=7.44 $Y2=0
r267 37 39 20.5135 $w=2.48e-07 $l=4.45e-07 $layer=LI1_cond $X=7.44 $Y=0.085
+ $X2=7.44 $Y2=0.53
r268 33 59 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.74 $Y=0.085
+ $X2=4.74 $Y2=0
r269 33 35 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=4.74 $Y=0.085
+ $X2=4.74 $Y2=0.73
r270 29 121 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.16 $Y=0.085
+ $X2=3.16 $Y2=0
r271 29 31 10.826 $w=3.28e-07 $l=3.1e-07 $layer=LI1_cond $X=3.16 $Y=0.085
+ $X2=3.16 $Y2=0.395
r272 25 118 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.22 $Y=0.085
+ $X2=1.22 $Y2=0
r273 25 27 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=1.22 $Y=0.085
+ $X2=1.22 $Y2=0.445
r274 8 55 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=15.115
+ $Y=0.37 $X2=15.255 $Y2=0.58
r275 7 51 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=12.98
+ $Y=0.285 $X2=13.12 $Y2=0.495
r276 6 47 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=11.615
+ $Y=0.33 $X2=11.755 $Y2=0.54
r277 5 43 182 $w=1.7e-07 $l=2.59856e-07 $layer=licon1_NDIFF $count=1 $X=9.035
+ $Y=0.625 $X2=9.215 $Y2=0.81
r278 4 39 182 $w=1.7e-07 $l=2.58167e-07 $layer=licon1_NDIFF $count=1 $X=7.265
+ $Y=0.625 $X2=7.48 $Y2=0.53
r279 3 35 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=4.6
+ $Y=0.565 $X2=4.74 $Y2=0.73
r280 2 31 182 $w=1.7e-07 $l=2.19089e-07 $layer=licon1_NDIFF $count=1 $X=3.02
+ $Y=0.235 $X2=3.16 $Y2=0.395
r281 1 27 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.08
+ $Y=0.235 $X2=1.22 $Y2=0.445
.ends

