* File: sky130_fd_sc_lp__o22a_lp.pex.spice
* Created: Fri Aug 28 11:10:02 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O22A_LP%A1 1 3 6 8 12
c28 6 0 4.68906e-20 $X=0.51 $Y=1.075
r29 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.45
+ $Y=1.67 $X2=0.45 $Y2=1.67
r30 8 12 8.64492 $w=5.03e-07 $l=3.65e-07 $layer=LI1_cond $X=0.362 $Y=2.035
+ $X2=0.362 $Y2=1.67
r31 4 11 41.312 $w=2.8e-07 $l=1.95806e-07 $layer=POLY_cond $X=0.51 $Y=1.49
+ $X2=0.477 $Y2=1.67
r32 4 6 212.798 $w=1.5e-07 $l=4.15e-07 $layer=POLY_cond $X=0.51 $Y=1.49 $X2=0.51
+ $Y2=1.075
r33 1 11 72.9649 $w=2.8e-07 $l=4.52725e-07 $layer=POLY_cond $X=0.545 $Y=2.09
+ $X2=0.477 $Y2=1.67
r34 1 3 97.364 $w=2.5e-07 $l=5.05e-07 $layer=POLY_cond $X=0.545 $Y=2.09
+ $X2=0.545 $Y2=2.595
.ends

.subckt PM_SKY130_FD_SC_LP__O22A_LP%A2 1 3 7 9 13
c41 3 0 1.24939e-19 $X=1.035 $Y=2.595
r42 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.99
+ $Y=1.67 $X2=0.99 $Y2=1.67
r43 9 13 8.64492 $w=5.03e-07 $l=3.65e-07 $layer=LI1_cond $X=1.077 $Y=2.035
+ $X2=1.077 $Y2=1.67
r44 5 12 40.7976 $w=3.24e-07 $l=2.04793e-07 $layer=POLY_cond $X=1.045 $Y=1.49
+ $X2=0.992 $Y2=1.67
r45 5 7 212.798 $w=1.5e-07 $l=4.15e-07 $layer=POLY_cond $X=1.045 $Y=1.49
+ $X2=1.045 $Y2=1.075
r46 1 12 27.1854 $w=3.24e-07 $l=1.85257e-07 $layer=POLY_cond $X=1.035 $Y=1.835
+ $X2=0.992 $Y2=1.67
r47 1 3 188.825 $w=2.5e-07 $l=7.6e-07 $layer=POLY_cond $X=1.035 $Y=1.835
+ $X2=1.035 $Y2=2.595
.ends

.subckt PM_SKY130_FD_SC_LP__O22A_LP%B2 4 7 10 11 12 13 18
c47 10 0 1.41198e-19 $X=1.545 $Y=1.735
r48 18 21 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.565 $Y=0.49
+ $X2=1.565 $Y2=0.655
r49 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.565
+ $Y=0.49 $X2=1.565 $Y2=0.49
r50 12 13 16.034 $w=3.43e-07 $l=4.8e-07 $layer=LI1_cond $X=1.68 $Y=0.497
+ $X2=2.16 $Y2=0.497
r51 12 19 3.84148 $w=3.43e-07 $l=1.15e-07 $layer=LI1_cond $X=1.68 $Y=0.497
+ $X2=1.565 $Y2=0.497
r52 11 19 12.1925 $w=3.43e-07 $l=3.65e-07 $layer=LI1_cond $X=1.2 $Y=0.497
+ $X2=1.565 $Y2=0.497
r53 9 10 47.1291 $w=2.5e-07 $l=1.5e-07 $layer=POLY_cond $X=1.545 $Y=1.585
+ $X2=1.545 $Y2=1.735
r54 7 10 213.67 $w=2.5e-07 $l=8.6e-07 $layer=POLY_cond $X=1.565 $Y=2.595
+ $X2=1.565 $Y2=1.735
r55 4 9 261.511 $w=1.5e-07 $l=5.1e-07 $layer=POLY_cond $X=1.475 $Y=1.075
+ $X2=1.475 $Y2=1.585
r56 4 21 215.362 $w=1.5e-07 $l=4.2e-07 $layer=POLY_cond $X=1.475 $Y=1.075
+ $X2=1.475 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__O22A_LP%B1 3 7 9 15
c34 15 0 5.90387e-20 $X=2.28 $Y=1.615
c35 9 0 1.41198e-19 $X=2.64 $Y=1.665
r36 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.28
+ $Y=1.615 $X2=2.28 $Y2=1.615
r37 13 15 28.8521 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.115 $Y=1.615
+ $X2=2.28 $Y2=1.615
r38 11 13 8.74306 $w=3.3e-07 $l=5e-08 $layer=POLY_cond $X=2.065 $Y=1.615
+ $X2=2.115 $Y2=1.615
r39 9 16 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=2.64 $Y=1.615
+ $X2=2.28 $Y2=1.615
r40 5 13 9.34494 $w=2.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.115 $Y=1.78
+ $X2=2.115 $Y2=1.615
r41 5 7 202.49 $w=2.5e-07 $l=8.15e-07 $layer=POLY_cond $X=2.115 $Y=1.78
+ $X2=2.115 $Y2=2.595
r42 1 11 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.065 $Y=1.45
+ $X2=2.065 $Y2=1.615
r43 1 3 192.287 $w=1.5e-07 $l=3.75e-07 $layer=POLY_cond $X=2.065 $Y=1.45
+ $X2=2.065 $Y2=1.075
.ends

.subckt PM_SKY130_FD_SC_LP__O22A_LP%A_232_419# 1 2 9 13 17 21 23 26 30 33 34 38
+ 39 42 44 45 46
c81 46 0 5.90387e-20 $X=3.1 $Y=1.525
c82 45 0 1.24939e-19 $X=1.81 $Y=2.045
r83 42 46 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=3.02 $Y=1.96
+ $X2=3.02 $Y2=1.525
r84 38 39 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.1 $Y=1.02
+ $X2=3.1 $Y2=1.02
r85 36 46 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=3.1 $Y=1.36 $X2=3.1
+ $Y2=1.525
r86 36 38 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=3.1 $Y=1.36 $X2=3.1
+ $Y2=1.02
r87 35 45 2.11342 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.935 $Y=2.045
+ $X2=1.81 $Y2=2.045
r88 34 42 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.935 $Y=2.045
+ $X2=3.02 $Y2=1.96
r89 34 35 65.2406 $w=1.68e-07 $l=1e-06 $layer=LI1_cond $X=2.935 $Y=2.045
+ $X2=1.935 $Y2=2.045
r90 32 45 4.3182 $w=2.1e-07 $l=1.03078e-07 $layer=LI1_cond $X=1.77 $Y=2.13
+ $X2=1.81 $Y2=2.045
r91 32 33 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=1.77 $Y=2.13
+ $X2=1.77 $Y2=2.31
r92 28 45 4.3182 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=1.81 $Y=1.96 $X2=1.81
+ $Y2=2.045
r93 28 30 27.4281 $w=2.48e-07 $l=5.95e-07 $layer=LI1_cond $X=1.81 $Y=1.96
+ $X2=1.81 $Y2=1.365
r94 27 44 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.465 $Y=2.395
+ $X2=1.3 $Y2=2.395
r95 26 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.685 $Y=2.395
+ $X2=1.77 $Y2=2.31
r96 26 27 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=1.685 $Y=2.395
+ $X2=1.465 $Y2=2.395
r97 22 39 42.4067 $w=4e-07 $l=3.05e-07 $layer=POLY_cond $X=3.11 $Y=1.325
+ $X2=3.11 $Y2=1.02
r98 22 23 35.5859 $w=4e-07 $l=2e-07 $layer=POLY_cond $X=3.11 $Y=1.325 $X2=3.11
+ $Y2=1.525
r99 21 39 2.08558 $w=4e-07 $l=1.5e-08 $layer=POLY_cond $X=3.11 $Y=1.005 $X2=3.11
+ $Y2=1.02
r100 13 23 265.845 $w=2.5e-07 $l=1.07e-06 $layer=POLY_cond $X=3.185 $Y=2.595
+ $X2=3.185 $Y2=1.525
r101 7 21 24.4565 $w=4e-07 $l=1.5e-07 $layer=POLY_cond $X=3.165 $Y=0.855
+ $X2=3.165 $Y2=1.005
r102 7 17 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=3.345 $Y=0.855
+ $X2=3.345 $Y2=0.445
r103 7 9 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=2.985 $Y=0.855
+ $X2=2.985 $Y2=0.445
r104 2 44 300 $w=1.7e-07 $l=4.44522e-07 $layer=licon1_PDIFF $count=2 $X=1.16
+ $Y=2.095 $X2=1.3 $Y2=2.475
r105 1 30 182 $w=1.7e-07 $l=6e-07 $layer=licon1_NDIFF $count=1 $X=1.55 $Y=0.865
+ $X2=1.77 $Y2=1.365
.ends

.subckt PM_SKY130_FD_SC_LP__O22A_LP%VPWR 1 2 7 9 13 16 17 18 31 32
r37 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r38 31 32 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r39 29 32 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r40 28 31 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.64 $Y=3.33 $X2=3.6
+ $Y2=3.33
r41 28 29 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r42 26 29 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r43 25 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r44 23 36 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r45 22 25 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=0.72 $Y=3.33
+ $X2=2.16 $Y2=3.33
r46 22 23 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r47 20 35 4.73185 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=3.33
+ $X2=0.222 $Y2=3.33
r48 20 22 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.445 $Y=3.33
+ $X2=0.72 $Y2=3.33
r49 18 26 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=2.16 $Y2=3.33
r50 18 23 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=0.72 $Y2=3.33
r51 16 25 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=2.22 $Y=3.33 $X2=2.16
+ $Y2=3.33
r52 16 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.22 $Y=3.33
+ $X2=2.385 $Y2=3.33
r53 15 28 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=2.55 $Y=3.33 $X2=2.64
+ $Y2=3.33
r54 15 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.55 $Y=3.33
+ $X2=2.385 $Y2=3.33
r55 11 17 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.385 $Y=3.245
+ $X2=2.385 $Y2=3.33
r56 11 13 26.8903 $w=3.28e-07 $l=7.7e-07 $layer=LI1_cond $X=2.385 $Y=3.245
+ $X2=2.385 $Y2=2.475
r57 7 35 3.03433 $w=3.3e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.28 $Y=3.245
+ $X2=0.222 $Y2=3.33
r58 7 9 26.8903 $w=3.28e-07 $l=7.7e-07 $layer=LI1_cond $X=0.28 $Y=3.245 $X2=0.28
+ $Y2=2.475
r59 2 13 300 $w=1.7e-07 $l=4.46654e-07 $layer=licon1_PDIFF $count=2 $X=2.24
+ $Y=2.095 $X2=2.385 $Y2=2.475
r60 1 9 300 $w=1.7e-07 $l=4.46654e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.095 $X2=0.28 $Y2=2.475
.ends

.subckt PM_SKY130_FD_SC_LP__O22A_LP%X 1 2 7 8 9 10 11 12 13 32
r22 33 47 1.44055 $w=4.38e-07 $l=5.5e-08 $layer=LI1_cond $X=3.505 $Y=2.295
+ $X2=3.505 $Y2=2.24
r23 32 45 1.92074 $w=2.38e-07 $l=4e-08 $layer=LI1_cond $X=3.605 $Y=2.035
+ $X2=3.605 $Y2=2.075
r24 12 13 9.691 $w=4.38e-07 $l=3.7e-07 $layer=LI1_cond $X=3.505 $Y=2.405
+ $X2=3.505 $Y2=2.775
r25 12 33 2.88111 $w=4.38e-07 $l=1.1e-07 $layer=LI1_cond $X=3.505 $Y=2.405
+ $X2=3.505 $Y2=2.295
r26 11 47 3.74544 $w=4.38e-07 $l=1.43e-07 $layer=LI1_cond $X=3.505 $Y=2.097
+ $X2=3.505 $Y2=2.24
r27 11 45 2.94049 $w=4.38e-07 $l=2.2e-08 $layer=LI1_cond $X=3.505 $Y=2.097
+ $X2=3.505 $Y2=2.075
r28 11 32 1.10442 $w=2.38e-07 $l=2.3e-08 $layer=LI1_cond $X=3.605 $Y=2.012
+ $X2=3.605 $Y2=2.035
r29 10 11 16.6624 $w=2.38e-07 $l=3.47e-07 $layer=LI1_cond $X=3.605 $Y=1.665
+ $X2=3.605 $Y2=2.012
r30 9 10 17.7668 $w=2.38e-07 $l=3.7e-07 $layer=LI1_cond $X=3.605 $Y=1.295
+ $X2=3.605 $Y2=1.665
r31 8 9 17.7668 $w=2.38e-07 $l=3.7e-07 $layer=LI1_cond $X=3.605 $Y=0.925
+ $X2=3.605 $Y2=1.295
r32 8 43 12.0046 $w=2.38e-07 $l=2.5e-07 $layer=LI1_cond $X=3.605 $Y=0.925
+ $X2=3.605 $Y2=0.675
r33 7 43 8.03684 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=3.56 $Y=0.47
+ $X2=3.56 $Y2=0.675
r34 2 47 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=3.31
+ $Y=2.095 $X2=3.45 $Y2=2.24
r35 1 7 182 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=1 $X=3.42
+ $Y=0.235 $X2=3.56 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_LP__O22A_LP%A_30_173# 1 2 3 12 14 15 19 20 21 22
c47 21 0 4.68906e-20 $X=1.505 $Y=0.935
r48 22 25 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=2.28 $Y=0.935
+ $X2=2.28 $Y2=1.085
r49 20 22 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.115 $Y=0.935
+ $X2=2.28 $Y2=0.935
r50 20 21 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=2.115 $Y=0.935
+ $X2=1.505 $Y2=0.935
r51 17 19 6.0433 $w=4.08e-07 $l=2.15e-07 $layer=LI1_cond $X=1.3 $Y=1.245 $X2=1.3
+ $Y2=1.03
r52 16 21 8.45803 $w=1.7e-07 $l=2.43824e-07 $layer=LI1_cond $X=1.3 $Y=1.02
+ $X2=1.505 $Y2=0.935
r53 16 19 0.281084 $w=4.08e-07 $l=1e-08 $layer=LI1_cond $X=1.3 $Y=1.02 $X2=1.3
+ $Y2=1.03
r54 14 17 8.45803 $w=1.7e-07 $l=2.43824e-07 $layer=LI1_cond $X=1.095 $Y=1.33
+ $X2=1.3 $Y2=1.245
r55 14 15 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.095 $Y=1.33
+ $X2=0.405 $Y2=1.33
r56 10 15 7.32204 $w=1.7e-07 $l=1.75425e-07 $layer=LI1_cond $X=0.267 $Y=1.245
+ $X2=0.405 $Y2=1.33
r57 10 12 9.01001 $w=2.73e-07 $l=2.15e-07 $layer=LI1_cond $X=0.267 $Y=1.245
+ $X2=0.267 $Y2=1.03
r58 3 25 182 $w=1.7e-07 $l=2.81425e-07 $layer=licon1_NDIFF $count=1 $X=2.14
+ $Y=0.865 $X2=2.28 $Y2=1.085
r59 2 19 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=1.12
+ $Y=0.865 $X2=1.26 $Y2=1.03
r60 1 12 182 $w=1.7e-07 $l=2.26164e-07 $layer=licon1_NDIFF $count=1 $X=0.15
+ $Y=0.865 $X2=0.295 $Y2=1.03
.ends

.subckt PM_SKY130_FD_SC_LP__O22A_LP%VGND 1 2 9 13 15 17 22 29 30 33 36
r41 36 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r42 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r43 30 37 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=2.64
+ $Y2=0
r44 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r45 27 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.935 $Y=0 $X2=2.77
+ $Y2=0
r46 27 29 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=2.935 $Y=0 $X2=3.6
+ $Y2=0
r47 26 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r48 25 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r49 23 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.905 $Y=0 $X2=0.74
+ $Y2=0
r50 23 25 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.905 $Y=0 $X2=1.2
+ $Y2=0
r51 22 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.605 $Y=0 $X2=2.77
+ $Y2=0
r52 22 25 91.6631 $w=1.68e-07 $l=1.405e-06 $layer=LI1_cond $X=2.605 $Y=0 $X2=1.2
+ $Y2=0
r53 20 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r54 19 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r55 17 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.575 $Y=0 $X2=0.74
+ $Y2=0
r56 17 19 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=0.575 $Y=0 $X2=0.24
+ $Y2=0
r57 15 37 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=2.64
+ $Y2=0
r58 15 26 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=1.2
+ $Y2=0
r59 11 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.77 $Y=0.085
+ $X2=2.77 $Y2=0
r60 11 13 11.5244 $w=3.28e-07 $l=3.3e-07 $layer=LI1_cond $X=2.77 $Y=0.085
+ $X2=2.77 $Y2=0.415
r61 7 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.74 $Y=0.085 $X2=0.74
+ $Y2=0
r62 7 9 31.6049 $w=3.28e-07 $l=9.05e-07 $layer=LI1_cond $X=0.74 $Y=0.085
+ $X2=0.74 $Y2=0.99
r63 2 13 182 $w=1.7e-07 $l=2.41868e-07 $layer=licon1_NDIFF $count=1 $X=2.625
+ $Y=0.235 $X2=2.77 $Y2=0.415
r64 1 9 182 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=1 $X=0.585
+ $Y=0.865 $X2=0.74 $Y2=0.99
.ends

