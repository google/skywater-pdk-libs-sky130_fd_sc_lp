* File: sky130_fd_sc_lp__nor2_m.pex.spice
* Created: Fri Aug 28 10:54:16 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__NOR2_M%A 2 5 8 10 11 12 13 14 20 22
c25 11 0 2.78553e-20 $X=0.24 $Y=0.925
r26 20 22 45.5639 $w=3.95e-07 $l=1.65e-07 $layer=POLY_cond $X=0.402 $Y=1.045
+ $X2=0.402 $Y2=0.88
r27 20 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.37
+ $Y=1.045 $X2=0.37 $Y2=1.045
r28 13 14 14.2135 $w=2.98e-07 $l=3.7e-07 $layer=LI1_cond $X=0.305 $Y=1.665
+ $X2=0.305 $Y2=2.035
r29 12 13 14.2135 $w=2.98e-07 $l=3.7e-07 $layer=LI1_cond $X=0.305 $Y=1.295
+ $X2=0.305 $Y2=1.665
r30 12 21 9.60369 $w=2.98e-07 $l=2.5e-07 $layer=LI1_cond $X=0.305 $Y=1.295
+ $X2=0.305 $Y2=1.045
r31 11 21 4.60977 $w=2.98e-07 $l=1.2e-07 $layer=LI1_cond $X=0.305 $Y=0.925
+ $X2=0.305 $Y2=1.045
r32 8 10 551.223 $w=1.5e-07 $l=1.075e-06 $layer=POLY_cond $X=0.525 $Y=2.625
+ $X2=0.525 $Y2=1.55
r33 5 22 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.525 $Y=0.56
+ $X2=0.525 $Y2=0.88
r34 2 10 50.0695 $w=3.95e-07 $l=1.97e-07 $layer=POLY_cond $X=0.402 $Y=1.353
+ $X2=0.402 $Y2=1.55
r35 1 20 4.50555 $w=3.95e-07 $l=3.2e-08 $layer=POLY_cond $X=0.402 $Y=1.077
+ $X2=0.402 $Y2=1.045
r36 1 2 38.8604 $w=3.95e-07 $l=2.76e-07 $layer=POLY_cond $X=0.402 $Y=1.077
+ $X2=0.402 $Y2=1.353
.ends

.subckt PM_SKY130_FD_SC_LP__NOR2_M%B 3 7 8 9 10 11 17 19
c25 19 0 2.78553e-20 $X=1.087 $Y=0.88
r26 17 20 83.1449 $w=4.95e-07 $l=5.05e-07 $layer=POLY_cond $X=1.087 $Y=1.045
+ $X2=1.087 $Y2=1.55
r27 17 19 46.3954 $w=4.95e-07 $l=1.65e-07 $layer=POLY_cond $X=1.087 $Y=1.045
+ $X2=1.087 $Y2=0.88
r28 17 18 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.17
+ $Y=1.045 $X2=1.17 $Y2=1.045
r29 10 11 20.5182 $w=1.98e-07 $l=3.7e-07 $layer=LI1_cond $X=1.185 $Y=1.665
+ $X2=1.185 $Y2=2.035
r30 9 10 20.5182 $w=1.98e-07 $l=3.7e-07 $layer=LI1_cond $X=1.185 $Y=1.295
+ $X2=1.185 $Y2=1.665
r31 9 18 13.8636 $w=1.98e-07 $l=2.5e-07 $layer=LI1_cond $X=1.185 $Y=1.295
+ $X2=1.185 $Y2=1.045
r32 8 18 6.65455 $w=1.98e-07 $l=1.2e-07 $layer=LI1_cond $X=1.185 $Y=0.925
+ $X2=1.185 $Y2=1.045
r33 7 19 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.955 $Y=0.56
+ $X2=0.955 $Y2=0.88
r34 3 20 551.223 $w=1.5e-07 $l=1.075e-06 $layer=POLY_cond $X=0.915 $Y=2.625
+ $X2=0.915 $Y2=1.55
.ends

.subckt PM_SKY130_FD_SC_LP__NOR2_M%VPWR 1 4 6 8 12 13
r14 16 17 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r15 12 13 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r16 10 16 3.63222 $w=1.7e-07 $l=2.08e-07 $layer=LI1_cond $X=0.415 $Y=3.33
+ $X2=0.207 $Y2=3.33
r17 10 12 51.2139 $w=1.68e-07 $l=7.85e-07 $layer=LI1_cond $X=0.415 $Y=3.33
+ $X2=1.2 $Y2=3.33
r18 8 13 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33 $X2=1.2
+ $Y2=3.33
r19 8 17 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r20 4 16 3.28297 $w=2.1e-07 $l=1.39155e-07 $layer=LI1_cond $X=0.31 $Y=3.245
+ $X2=0.207 $Y2=3.33
r21 4 6 31.9524 $w=2.08e-07 $l=6.05e-07 $layer=LI1_cond $X=0.31 $Y=3.245
+ $X2=0.31 $Y2=2.64
r22 1 6 600 $w=1.7e-07 $l=2.80624e-07 $layer=licon1_PDIFF $count=1 $X=0.185
+ $Y=2.415 $X2=0.31 $Y2=2.64
.ends

.subckt PM_SKY130_FD_SC_LP__NOR2_M%Y 1 2 7 8 9 10 11 22 36
c19 36 0 6.97414e-20 $X=0.76 $Y=2.627
r20 36 38 9.89912 $w=4.56e-07 $l=3.7e-07 $layer=LI1_cond $X=0.76 $Y=2.627
+ $X2=1.13 $Y2=2.627
r21 20 36 4.25555 $w=2.5e-07 $l=2.32e-07 $layer=LI1_cond $X=0.76 $Y=2.395
+ $X2=0.76 $Y2=2.627
r22 11 36 1.07018 $w=4.56e-07 $l=4e-08 $layer=LI1_cond $X=0.72 $Y=2.627 $X2=0.76
+ $Y2=2.627
r23 11 20 1.75171 $w=2.48e-07 $l=3.8e-08 $layer=LI1_cond $X=0.76 $Y=2.357
+ $X2=0.76 $Y2=2.395
r24 10 11 14.8435 $w=2.48e-07 $l=3.22e-07 $layer=LI1_cond $X=0.76 $Y=2.035
+ $X2=0.76 $Y2=2.357
r25 9 10 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=0.76 $Y=1.665
+ $X2=0.76 $Y2=2.035
r26 8 9 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=0.76 $Y=1.295 $X2=0.76
+ $Y2=1.665
r27 7 8 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=0.76 $Y=0.925 $X2=0.76
+ $Y2=1.295
r28 7 22 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=0.76 $Y=0.925 $X2=0.76
+ $Y2=0.495
r29 2 38 600 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_PDIFF $count=1 $X=0.99
+ $Y=2.415 $X2=1.13 $Y2=2.63
r30 1 22 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=0.6
+ $Y=0.35 $X2=0.74 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__NOR2_M%VGND 1 2 7 9 11 13 15 17 27
r23 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r24 23 24 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r25 18 23 3.63222 $w=1.7e-07 $l=2.08e-07 $layer=LI1_cond $X=0.415 $Y=0 $X2=0.207
+ $Y2=0
r26 18 20 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.415 $Y=0 $X2=0.72
+ $Y2=0
r27 17 26 3.65294 $w=1.7e-07 $l=1.87e-07 $layer=LI1_cond $X=1.065 $Y=0 $X2=1.252
+ $Y2=0
r28 17 20 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.065 $Y=0 $X2=0.72
+ $Y2=0
r29 15 27 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r30 15 24 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r31 15 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r32 11 26 3.26225 $w=2.1e-07 $l=1.19143e-07 $layer=LI1_cond $X=1.17 $Y=0.085
+ $X2=1.252 $Y2=0
r33 11 13 21.6537 $w=2.08e-07 $l=4.1e-07 $layer=LI1_cond $X=1.17 $Y=0.085
+ $X2=1.17 $Y2=0.495
r34 7 23 3.28297 $w=2.1e-07 $l=1.39155e-07 $layer=LI1_cond $X=0.31 $Y=0.085
+ $X2=0.207 $Y2=0
r35 7 9 21.6537 $w=2.08e-07 $l=4.1e-07 $layer=LI1_cond $X=0.31 $Y=0.085 $X2=0.31
+ $Y2=0.495
r36 2 13 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=1.03
+ $Y=0.35 $X2=1.17 $Y2=0.495
r37 1 9 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.185
+ $Y=0.35 $X2=0.31 $Y2=0.495
.ends

