# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__a21bo_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_lp__a21bo_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.840000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.315000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.075000 1.210000 2.810000 1.460000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.315000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.020000 1.210000 3.755000 1.460000 ;
    END
  END A2
  PIN B1_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.005000 1.345000 1.285000 1.750000 ;
    END
  END B1_N
  PIN X
    ANTENNADIFFAREA  0.556500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.325000 0.365000 1.815000 ;
        RECT 0.085000 1.815000 0.465000 3.075000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.840000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.840000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.840000 0.085000 ;
      RECT 0.000000  3.245000 3.840000 3.415000 ;
      RECT 0.535000  1.295000 0.825000 1.625000 ;
      RECT 0.635000  2.660000 0.965000 3.245000 ;
      RECT 0.640000  0.085000 0.970000 0.465000 ;
      RECT 0.655000  0.635000 2.575000 0.805000 ;
      RECT 0.655000  0.805000 0.825000 1.295000 ;
      RECT 0.655000  1.625000 0.825000 2.320000 ;
      RECT 0.655000  2.320000 2.025000 2.490000 ;
      RECT 1.160000  1.930000 1.635000 2.140000 ;
      RECT 1.185000  0.975000 1.635000 1.175000 ;
      RECT 1.465000  1.175000 1.635000 1.345000 ;
      RECT 1.465000  1.345000 1.895000 1.675000 ;
      RECT 1.465000  1.675000 1.635000 1.930000 ;
      RECT 1.725000  0.085000 2.055000 0.465000 ;
      RECT 1.725000  2.490000 2.025000 3.075000 ;
      RECT 1.805000  1.845000 2.025000 2.320000 ;
      RECT 2.195000  1.630000 3.415000 1.800000 ;
      RECT 2.195000  1.800000 2.455000 3.075000 ;
      RECT 2.245000  0.255000 2.575000 0.635000 ;
      RECT 2.245000  0.805000 2.575000 1.040000 ;
      RECT 2.635000  1.970000 2.965000 3.245000 ;
      RECT 3.115000  0.085000 3.445000 1.040000 ;
      RECT 3.175000  1.800000 3.415000 3.075000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
  END
END sky130_fd_sc_lp__a21bo_1
END LIBRARY
