* File: sky130_fd_sc_lp__a311oi_m.spice
* Created: Fri Aug 28 09:58:51 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__a311oi_m.pex.spice"
.subckt sky130_fd_sc_lp__a311oi_m  VNB VPB A3 A2 A1 B1 C1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* C1	C1
* B1	B1
* A1	A1
* A2	A2
* A3	A3
* VPB	VPB
* VNB	VNB
MM1001 A_199_51# N_A3_M1001_g N_VGND_M1001_s VNB NSHORT L=0.15 W=0.42 AD=0.0441
+ AS=0.2982 PD=0.63 PS=2.26 NRD=14.28 NRS=127.14 M=1 R=2.8 SA=75000.6 SB=75001.8
+ A=0.063 P=1.14 MULT=1
MM1008 A_271_51# N_A2_M1008_g A_199_51# VNB NSHORT L=0.15 W=0.42 AD=0.0441
+ AS=0.0441 PD=0.63 PS=0.63 NRD=14.28 NRS=14.28 M=1 R=2.8 SA=75001 SB=75001.4
+ A=0.063 P=1.14 MULT=1
MM1009 N_Y_M1009_d N_A1_M1009_g A_271_51# VNB NSHORT L=0.15 W=0.42 AD=0.0588
+ AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.4 SB=75001.1
+ A=0.063 P=1.14 MULT=1
MM1002 N_VGND_M1002_d N_B1_M1002_g N_Y_M1009_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.8 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1005 N_Y_M1005_d N_C1_M1005_g N_VGND_M1002_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75002.2 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1006 N_A_191_535#_M1006_d N_A3_M1006_g N_VPWR_M1006_s VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0588 AS=0.2814 PD=0.7 PS=2.18 NRD=0 NRS=189.947 M=1 R=2.8
+ SA=75000.6 SB=75001.8 A=0.063 P=1.14 MULT=1
MM1004 N_VPWR_M1004_d N_A2_M1004_g N_A_191_535#_M1006_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1000 N_A_191_535#_M1000_d N_A1_M1000_g N_VPWR_M1004_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.5
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1007 A_449_535# N_B1_M1007_g N_A_191_535#_M1000_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=23.443 NRS=0 M=1 R=2.8 SA=75001.9
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1003 N_Y_M1003_d N_C1_M1003_g A_449_535# VPB PHIGHVT L=0.15 W=0.42 AD=0.1134
+ AS=0.0441 PD=1.38 PS=0.63 NRD=2.3443 NRS=23.443 M=1 R=2.8 SA=75002.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9751 P=11.21
c_38 VNB 0 1.60224e-19 $X=0 $Y=0
*
.include "sky130_fd_sc_lp__a311oi_m.pxi.spice"
*
.ends
*
*
