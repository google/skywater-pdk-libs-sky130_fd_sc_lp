* NGSPICE file created from sky130_fd_sc_lp__dlrbp_2.ext - technology: sky130A

.subckt sky130_fd_sc_lp__dlrbp_2 D GATE RESET_B VGND VNB VPB VPWR Q Q_N
M1000 a_823_25# a_1023_405# a_981_503# VPB phighvt w=420000u l=150000u
+  ad=2.158e+11p pd=2.03e+06u as=1.848e+11p ps=1.72e+06u
M1001 Q a_432_109# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=3.528e+11p pd=3.08e+06u as=2.5951e+12p ps=2.041e+07u
M1002 a_781_51# RESET_B VGND VNB nshort w=840000u l=150000u
+  ad=1.764e+11p pd=2.1e+06u as=1.4721e+12p ps=1.368e+07u
M1003 a_432_109# RESET_B VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=3.528e+11p pd=3.08e+06u as=0p ps=0u
M1004 VPWR a_1109_21# a_1023_405# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.696e+11p ps=1.81e+06u
M1005 a_432_109# a_823_25# a_781_51# VNB nshort w=840000u l=150000u
+  ad=2.394e+11p pd=2.25e+06u as=0p ps=0u
M1006 VPWR a_80_21# Q_N VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=3.591e+11p ps=3.09e+06u
M1007 Q_N a_80_21# VGND VNB nshort w=840000u l=150000u
+  ad=2.352e+11p pd=2.24e+06u as=0p ps=0u
M1008 a_1109_21# GATE VPWR VPB phighvt w=640000u l=150000u
+  ad=1.824e+11p pd=1.85e+06u as=0p ps=0u
M1009 VGND a_432_109# a_80_21# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1010 VGND a_1109_21# a_1023_405# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1011 Q a_432_109# VGND VNB nshort w=840000u l=150000u
+  ad=2.352e+11p pd=2.24e+06u as=0p ps=0u
M1012 VGND a_80_21# Q_N VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_823_25# a_1109_21# a_1067_119# VNB nshort w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=8.82e+10p ps=1.26e+06u
M1014 VPWR a_432_109# Q VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_981_503# a_432_109# VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_1204_459# a_1109_21# a_823_25# VPB phighvt w=640000u l=150000u
+  ad=1.344e+11p pd=1.7e+06u as=0p ps=0u
M1017 a_1246_339# D VPWR VPB phighvt w=640000u l=150000u
+  ad=1.824e+11p pd=1.85e+06u as=0p ps=0u
M1018 a_1225_119# a_1023_405# a_823_25# VNB nshort w=420000u l=150000u
+  ad=1.344e+11p pd=1.48e+06u as=0p ps=0u
M1019 a_1067_119# a_432_109# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_1109_21# GATE VGND VNB nshort w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1021 VPWR a_432_109# a_80_21# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.824e+11p ps=1.85e+06u
M1022 VPWR a_823_25# a_432_109# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 VPWR a_1246_339# a_1204_459# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 VGND a_1246_339# a_1225_119# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 VGND a_432_109# Q VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_1246_339# D VGND VNB nshort w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1027 Q_N a_80_21# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

