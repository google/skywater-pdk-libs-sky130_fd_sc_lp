* File: sky130_fd_sc_lp__clkbuf_2.pex.spice
* Created: Fri Aug 28 10:14:55 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__CLKBUF_2%A 3 6 8 11 13
r31 11 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.51 $Y=0.94
+ $X2=0.51 $Y2=1.105
r32 11 13 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.51 $Y=0.94
+ $X2=0.51 $Y2=0.775
r33 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.51
+ $Y=0.94 $X2=0.51 $Y2=0.94
r34 8 12 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=0.72 $Y=0.94 $X2=0.51
+ $Y2=0.94
r35 6 14 697.362 $w=1.5e-07 $l=1.36e-06 $layer=POLY_cond $X=0.475 $Y=2.465
+ $X2=0.475 $Y2=1.105
r36 3 13 106.04 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=0.475 $Y=0.445
+ $X2=0.475 $Y2=0.775
.ends

.subckt PM_SKY130_FD_SC_LP__CLKBUF_2%A_27_47# 1 2 9 13 17 21 24 27 33 39 41 45
r63 45 46 0.710914 $w=3.39e-07 $l=5e-09 $layer=POLY_cond $X=1.385 $Y=1.375
+ $X2=1.39 $Y2=1.375
r64 42 43 0.710914 $w=3.39e-07 $l=5e-09 $layer=POLY_cond $X=0.955 $Y=1.375
+ $X2=0.96 $Y2=1.375
r65 36 39 3.05058 $w=3.38e-07 $l=9e-08 $layer=LI1_cond $X=0.17 $Y=0.435 $X2=0.26
+ $Y2=0.435
r66 34 45 47.6313 $w=3.39e-07 $l=3.35e-07 $layer=POLY_cond $X=1.05 $Y=1.375
+ $X2=1.385 $Y2=1.375
r67 34 43 12.7965 $w=3.39e-07 $l=9e-08 $layer=POLY_cond $X=1.05 $Y=1.375
+ $X2=0.96 $Y2=1.375
r68 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.05
+ $Y=1.38 $X2=1.05 $Y2=1.38
r69 31 41 1.05597 $w=2.6e-07 $l=1.55e-07 $layer=LI1_cond $X=0.395 $Y=1.405
+ $X2=0.24 $Y2=1.405
r70 31 33 29.0327 $w=2.58e-07 $l=6.55e-07 $layer=LI1_cond $X=0.395 $Y=1.405
+ $X2=1.05 $Y2=1.405
r71 27 29 31.2275 $w=3.08e-07 $l=8.4e-07 $layer=LI1_cond $X=0.24 $Y=2.04
+ $X2=0.24 $Y2=2.88
r72 25 41 5.51899 $w=2.4e-07 $l=1.3e-07 $layer=LI1_cond $X=0.24 $Y=1.535
+ $X2=0.24 $Y2=1.405
r73 25 27 18.7737 $w=3.08e-07 $l=5.05e-07 $layer=LI1_cond $X=0.24 $Y=1.535
+ $X2=0.24 $Y2=2.04
r74 24 41 5.51899 $w=2.4e-07 $l=1.61245e-07 $layer=LI1_cond $X=0.17 $Y=1.275
+ $X2=0.24 $Y2=1.405
r75 23 36 4.80115 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=0.17 $Y=0.605
+ $X2=0.17 $Y2=0.435
r76 23 24 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=0.17 $Y=0.605
+ $X2=0.17 $Y2=1.275
r77 19 46 21.8644 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=1.39 $Y=1.205
+ $X2=1.39 $Y2=1.375
r78 19 21 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=1.39 $Y=1.205
+ $X2=1.39 $Y2=0.445
r79 15 45 21.8644 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=1.385 $Y=1.545
+ $X2=1.385 $Y2=1.375
r80 15 17 471.745 $w=1.5e-07 $l=9.2e-07 $layer=POLY_cond $X=1.385 $Y=1.545
+ $X2=1.385 $Y2=2.465
r81 11 43 21.8644 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=0.96 $Y=1.205
+ $X2=0.96 $Y2=1.375
r82 11 13 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=0.96 $Y=1.205
+ $X2=0.96 $Y2=0.445
r83 7 42 21.8644 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=0.955 $Y=1.545
+ $X2=0.955 $Y2=1.375
r84 7 9 471.745 $w=1.5e-07 $l=9.2e-07 $layer=POLY_cond $X=0.955 $Y=1.545
+ $X2=0.955 $Y2=2.465
r85 2 29 400 $w=1.7e-07 $l=1.10574e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.835 $X2=0.26 $Y2=2.88
r86 2 27 400 $w=1.7e-07 $l=2.60096e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.835 $X2=0.26 $Y2=2.04
r87 1 39 182 $w=1.7e-07 $l=2.60096e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.44
.ends

.subckt PM_SKY130_FD_SC_LP__CLKBUF_2%VPWR 1 2 9 13 15 19 21 26 32 36
r26 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r27 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r28 30 36 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r29 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r30 27 32 8.23795 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=0.875 $Y=3.33
+ $X2=0.72 $Y2=3.33
r31 27 29 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.875 $Y=3.33
+ $X2=1.2 $Y2=3.33
r32 26 35 3.96354 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=1.475 $Y=3.33
+ $X2=1.697 $Y2=3.33
r33 26 29 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=1.475 $Y=3.33
+ $X2=1.2 $Y2=3.33
r34 24 33 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r35 23 24 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r36 21 32 8.23795 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=0.565 $Y=3.33
+ $X2=0.72 $Y2=3.33
r37 21 23 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.565 $Y=3.33
+ $X2=0.24 $Y2=3.33
r38 19 30 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=0.96 $Y=3.33
+ $X2=1.2 $Y2=3.33
r39 19 33 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=0.96 $Y=3.33
+ $X2=0.72 $Y2=3.33
r40 15 18 31.6357 $w=2.53e-07 $l=7e-07 $layer=LI1_cond $X=1.602 $Y=2.23
+ $X2=1.602 $Y2=2.93
r41 13 35 3.21368 $w=2.55e-07 $l=1.30767e-07 $layer=LI1_cond $X=1.602 $Y=3.245
+ $X2=1.697 $Y2=3.33
r42 13 18 14.2361 $w=2.53e-07 $l=3.15e-07 $layer=LI1_cond $X=1.602 $Y=3.245
+ $X2=1.602 $Y2=2.93
r43 9 12 31.2275 $w=3.08e-07 $l=8.4e-07 $layer=LI1_cond $X=0.72 $Y=2.04 $X2=0.72
+ $Y2=2.88
r44 7 32 0.701276 $w=3.1e-07 $l=8.5e-08 $layer=LI1_cond $X=0.72 $Y=3.245
+ $X2=0.72 $Y2=3.33
r45 7 12 13.5691 $w=3.08e-07 $l=3.65e-07 $layer=LI1_cond $X=0.72 $Y=3.245
+ $X2=0.72 $Y2=2.88
r46 2 18 400 $w=1.7e-07 $l=1.1629e-06 $layer=licon1_PDIFF $count=1 $X=1.46
+ $Y=1.835 $X2=1.6 $Y2=2.93
r47 2 15 400 $w=1.7e-07 $l=4.59701e-07 $layer=licon1_PDIFF $count=1 $X=1.46
+ $Y=1.835 $X2=1.6 $Y2=2.23
r48 1 12 400 $w=1.7e-07 $l=1.1128e-06 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=1.835 $X2=0.69 $Y2=2.88
r49 1 9 400 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=1.835 $X2=0.69 $Y2=2.04
.ends

.subckt PM_SKY130_FD_SC_LP__CLKBUF_2%X 1 2 9 13 14 15 16 17 26 36
r33 31 36 1.60806 $w=4.28e-07 $l=6e-08 $layer=LI1_cond $X=1.6 $Y=1.725 $X2=1.6
+ $Y2=1.665
r34 17 31 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=1.68 $Y=1.81 $X2=1.6
+ $Y2=1.81
r35 17 36 0.348413 $w=4.28e-07 $l=1.3e-08 $layer=LI1_cond $X=1.6 $Y=1.652
+ $X2=1.6 $Y2=1.665
r36 16 17 9.56796 $w=4.28e-07 $l=3.57e-07 $layer=LI1_cond $X=1.6 $Y=1.295
+ $X2=1.6 $Y2=1.652
r37 16 30 5.09219 $w=4.28e-07 $l=1.9e-07 $layer=LI1_cond $X=1.6 $Y=1.295 $X2=1.6
+ $Y2=1.105
r38 15 30 2.83678 $w=3.23e-07 $l=8e-08 $layer=LI1_cond $X=1.68 $Y=0.942 $X2=1.6
+ $Y2=0.942
r39 14 30 14.1839 $w=3.23e-07 $l=4e-07 $layer=LI1_cond $X=1.2 $Y=0.942 $X2=1.6
+ $Y2=0.942
r40 14 24 0.886495 $w=3.23e-07 $l=2.5e-08 $layer=LI1_cond $X=1.2 $Y=0.942
+ $X2=1.175 $Y2=0.942
r41 13 24 9.97306 $w=2.58e-07 $l=2.25e-07 $layer=LI1_cond $X=1.175 $Y=0.555
+ $X2=1.175 $Y2=0.78
r42 13 26 5.09734 $w=2.58e-07 $l=1.15e-07 $layer=LI1_cond $X=1.175 $Y=0.555
+ $X2=1.175 $Y2=0.44
r43 9 11 37.2328 $w=2.58e-07 $l=8.4e-07 $layer=LI1_cond $X=1.175 $Y=2.04
+ $X2=1.175 $Y2=2.88
r44 7 31 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=1.175 $Y=1.81
+ $X2=1.6 $Y2=1.81
r45 7 9 6.42709 $w=2.58e-07 $l=1.45e-07 $layer=LI1_cond $X=1.175 $Y=1.895
+ $X2=1.175 $Y2=2.04
r46 2 11 400 $w=1.7e-07 $l=1.1128e-06 $layer=licon1_PDIFF $count=1 $X=1.03
+ $Y=1.835 $X2=1.17 $Y2=2.88
r47 2 9 400 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=1 $X=1.03
+ $Y=1.835 $X2=1.17 $Y2=2.04
r48 1 26 182 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_NDIFF $count=1 $X=1.035
+ $Y=0.235 $X2=1.175 $Y2=0.44
.ends

.subckt PM_SKY130_FD_SC_LP__CLKBUF_2%VGND 1 2 9 11 13 15 17 22 28 32
r29 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r30 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r31 26 32 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r32 25 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r33 23 28 7.54988 $w=1.7e-07 $l=1.38e-07 $layer=LI1_cond $X=0.83 $Y=0 $X2=0.692
+ $Y2=0
r34 23 25 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.83 $Y=0 $X2=1.2
+ $Y2=0
r35 22 31 3.96354 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=1.475 $Y=0 $X2=1.697
+ $Y2=0
r36 22 25 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=1.475 $Y=0 $X2=1.2
+ $Y2=0
r37 20 29 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r38 19 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r39 17 28 7.54988 $w=1.7e-07 $l=1.37e-07 $layer=LI1_cond $X=0.555 $Y=0 $X2=0.692
+ $Y2=0
r40 17 19 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.555 $Y=0 $X2=0.24
+ $Y2=0
r41 15 26 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=0.96 $Y=0 $X2=1.2
+ $Y2=0
r42 15 29 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=0.96 $Y=0 $X2=0.72
+ $Y2=0
r43 11 31 3.21368 $w=2.55e-07 $l=1.30767e-07 $layer=LI1_cond $X=1.602 $Y=0.085
+ $X2=1.697 $Y2=0
r44 11 13 16.2698 $w=2.53e-07 $l=3.6e-07 $layer=LI1_cond $X=1.602 $Y=0.085
+ $X2=1.602 $Y2=0.445
r45 7 28 0.316938 $w=2.75e-07 $l=8.5e-08 $layer=LI1_cond $X=0.692 $Y=0.085
+ $X2=0.692 $Y2=0
r46 7 9 14.877 $w=2.73e-07 $l=3.55e-07 $layer=LI1_cond $X=0.692 $Y=0.085
+ $X2=0.692 $Y2=0.44
r47 2 13 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.465
+ $Y=0.235 $X2=1.605 $Y2=0.445
r48 1 9 182 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.235 $X2=0.69 $Y2=0.44
.ends

