* File: sky130_fd_sc_lp__o2111ai_4.spice
* Created: Fri Aug 28 11:01:11 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__o2111ai_4.pex.spice"
.subckt sky130_fd_sc_lp__o2111ai_4  VNB VPB D1 C1 B1 A2 A1 Y VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Y	Y
* A1	A1
* A2	A2
* B1	B1
* C1	C1
* D1	D1
* VPB	VPB
* VNB	VNB
MM1010 N_Y_M1010_d N_D1_M1010_g N_A_27_47#_M1010_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75003.2 A=0.126 P=1.98 MULT=1
MM1017 N_Y_M1010_d N_D1_M1017_g N_A_27_47#_M1017_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75002.8 A=0.126 P=1.98 MULT=1
MM1019 N_Y_M1019_d N_D1_M1019_g N_A_27_47#_M1017_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.1
+ SB=75002.3 A=0.126 P=1.98 MULT=1
MM1037 N_Y_M1019_d N_D1_M1037_g N_A_27_47#_M1037_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.5
+ SB=75001.9 A=0.126 P=1.98 MULT=1
MM1007 N_A_27_47#_M1037_s N_C1_M1007_g N_A_454_47#_M1007_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.9
+ SB=75001.5 A=0.126 P=1.98 MULT=1
MM1013 N_A_27_47#_M1013_d N_C1_M1013_g N_A_454_47#_M1007_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002.3
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1029 N_A_27_47#_M1013_d N_C1_M1029_g N_A_454_47#_M1029_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002.8
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1031 N_A_27_47#_M1031_d N_C1_M1031_g N_A_454_47#_M1029_s VNB NSHORT L=0.15
+ W=0.84 AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75003.2
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1001 N_A_819_47#_M1001_d N_B1_M1001_g N_A_454_47#_M1001_s VNB NSHORT L=0.15
+ W=0.84 AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75005.3 A=0.126 P=1.98 MULT=1
MM1016 N_A_819_47#_M1016_d N_B1_M1016_g N_A_454_47#_M1001_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75004.9 A=0.126 P=1.98 MULT=1
MM1022 N_A_819_47#_M1016_d N_B1_M1022_g N_A_454_47#_M1022_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.1
+ SB=75004.4 A=0.126 P=1.98 MULT=1
MM1033 N_A_819_47#_M1033_d N_B1_M1033_g N_A_454_47#_M1022_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.5
+ SB=75004 A=0.126 P=1.98 MULT=1
MM1008 N_VGND_M1008_d N_A2_M1008_g N_A_819_47#_M1033_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.9
+ SB=75003.6 A=0.126 P=1.98 MULT=1
MM1020 N_VGND_M1008_d N_A2_M1020_g N_A_819_47#_M1020_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002.3
+ SB=75003.1 A=0.126 P=1.98 MULT=1
MM1021 N_VGND_M1021_d N_A2_M1021_g N_A_819_47#_M1020_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002.8
+ SB=75002.7 A=0.126 P=1.98 MULT=1
MM1038 N_VGND_M1021_d N_A2_M1038_g N_A_819_47#_M1038_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2688 PD=1.12 PS=1.48 NRD=0 NRS=0 M=1 R=5.6 SA=75003.2
+ SB=75002.3 A=0.126 P=1.98 MULT=1
MM1018 N_A_819_47#_M1038_s N_A1_M1018_g N_VGND_M1018_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2688 AS=0.1176 PD=1.48 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75004 SB=75001.5
+ A=0.126 P=1.98 MULT=1
MM1034 N_A_819_47#_M1034_d N_A1_M1034_g N_VGND_M1018_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75004.4
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1035 N_A_819_47#_M1034_d N_A1_M1035_g N_VGND_M1035_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75004.9
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1039 N_A_819_47#_M1039_d N_A1_M1039_g N_VGND_M1035_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75005.3
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1000 N_VPWR_M1000_d N_D1_M1000_g N_Y_M1000_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2 SB=75007
+ A=0.189 P=2.82 MULT=1
MM1011 N_VPWR_M1000_d N_D1_M1011_g N_Y_M1011_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75006.5 A=0.189 P=2.82 MULT=1
MM1024 N_VPWR_M1024_d N_D1_M1024_g N_Y_M1011_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75006.1 A=0.189 P=2.82 MULT=1
MM1036 N_VPWR_M1024_d N_D1_M1036_g N_Y_M1036_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.5
+ SB=75005.7 A=0.189 P=2.82 MULT=1
MM1004 N_VPWR_M1004_d N_C1_M1004_g N_Y_M1036_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.9
+ SB=75005.3 A=0.189 P=2.82 MULT=1
MM1009 N_VPWR_M1004_d N_C1_M1009_g N_Y_M1009_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.3
+ SB=75004.8 A=0.189 P=2.82 MULT=1
MM1025 N_VPWR_M1025_d N_C1_M1025_g N_Y_M1009_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.8
+ SB=75004.4 A=0.189 P=2.82 MULT=1
MM1030 N_VPWR_M1025_d N_C1_M1030_g N_Y_M1030_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.3906 PD=1.54 PS=1.88 NRD=0 NRS=0 M=1 R=8.4 SA=75003.2 SB=75004
+ A=0.189 P=2.82 MULT=1
MM1002 N_VPWR_M1002_d N_B1_M1002_g N_Y_M1030_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.3906 PD=1.54 PS=1.88 NRD=0 NRS=0 M=1 R=8.4 SA=75004 SB=75003.2
+ A=0.189 P=2.82 MULT=1
MM1005 N_VPWR_M1002_d N_B1_M1005_g N_Y_M1005_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75004.4
+ SB=75002.8 A=0.189 P=2.82 MULT=1
MM1014 N_VPWR_M1014_d N_B1_M1014_g N_Y_M1005_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75004.8
+ SB=75002.3 A=0.189 P=2.82 MULT=1
MM1032 N_VPWR_M1014_d N_B1_M1032_g N_Y_M1032_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75005.3
+ SB=75001.9 A=0.189 P=2.82 MULT=1
MM1003 N_A_1210_367#_M1003_d N_A2_M1003_g N_Y_M1032_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75005.7
+ SB=75001.5 A=0.189 P=2.82 MULT=1
MM1015 N_A_1210_367#_M1003_d N_A2_M1015_g N_Y_M1015_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75006.1
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1026 N_A_1210_367#_M1026_d N_A2_M1026_g N_Y_M1015_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75006.5
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1027 N_A_1210_367#_M1026_d N_A2_M1027_g N_Y_M1027_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75007 SB=75000.2
+ A=0.189 P=2.82 MULT=1
MM1006 N_A_1210_367#_M1006_d N_A1_M1006_g N_VPWR_M1006_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75001.5 A=0.189 P=2.82 MULT=1
MM1012 N_A_1210_367#_M1006_d N_A1_M1012_g N_VPWR_M1012_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1023 N_A_1210_367#_M1023_d N_A1_M1023_g N_VPWR_M1012_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1028 N_A_1210_367#_M1023_d N_A1_M1028_g N_VPWR_M1028_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75001.5
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX40_noxref VNB VPB NWDIODE A=19.5079 P=24.65
*
.include "sky130_fd_sc_lp__o2111ai_4.pxi.spice"
*
.ends
*
*
