* File: sky130_fd_sc_lp__busdrivernovlpsleep_20.pex.spice
* Created: Wed Sep  2 09:37:27 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__BUSDRIVERNOVLPSLEEP_20%SLEEP 3 7 11 15 19 23 27 31
+ 35 37 42 45 46 47 48 53 54 56 60 66 69 74
c226 60 0 1.07875e-19 $X=5.51 $Y=1.93
c227 53 0 1.92998e-19 $X=11.865 $Y=2.035
c228 48 0 1.73847e-19 $X=5.645 $Y=2.035
c229 47 0 2.97955e-19 $X=11.72 $Y=2.035
c230 46 0 6.74658e-20 $X=0.915 $Y=2.035
c231 42 0 9.84968e-20 $X=11.95 $Y=1.445
c232 37 0 4.91905e-20 $X=5.71 $Y=1.93
r233 69 70 63.3823 $w=3.27e-07 $l=4.3e-07 $layer=POLY_cond $X=1.325 $Y=1.415
+ $X2=1.755 $Y2=1.415
r234 68 69 38.3242 $w=3.27e-07 $l=2.6e-07 $layer=POLY_cond $X=1.065 $Y=1.415
+ $X2=1.325 $Y2=1.415
r235 67 68 33.9021 $w=3.27e-07 $l=2.3e-07 $layer=POLY_cond $X=0.835 $Y=1.415
+ $X2=1.065 $Y2=1.415
r236 66 79 21.652 $w=3.28e-07 $l=6.2e-07 $layer=LI1_cond $X=0.76 $Y=1.415
+ $X2=0.76 $Y2=2.035
r237 65 67 11.055 $w=3.27e-07 $l=7.5e-08 $layer=POLY_cond $X=0.76 $Y=1.415
+ $X2=0.835 $Y2=1.415
r238 65 66 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.76
+ $Y=1.415 $X2=0.76 $Y2=1.415
r239 63 65 34.6391 $w=3.27e-07 $l=2.35e-07 $layer=POLY_cond $X=0.525 $Y=1.415
+ $X2=0.76 $Y2=1.415
r240 62 63 7.37003 $w=3.27e-07 $l=5e-08 $layer=POLY_cond $X=0.475 $Y=1.415
+ $X2=0.525 $Y2=1.415
r241 59 60 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.51
+ $Y=1.93 $X2=5.51 $Y2=1.93
r242 56 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.77 $Y=2.035
+ $X2=0.77 $Y2=2.035
r243 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.865 $Y=2.035
+ $X2=11.865 $Y2=2.035
r244 50 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.5 $Y=2.035
+ $X2=5.5 $Y2=2.035
r245 48 50 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.645 $Y=2.035
+ $X2=5.5 $Y2=2.035
r246 47 53 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=11.72 $Y=2.035
+ $X2=11.865 $Y2=2.035
r247 47 48 5.84951 $w=1.7e-07 $l=6.075e-06 $layer=MET1_cond $X=11.72 $Y=2.035
+ $X2=5.645 $Y2=2.035
r248 46 56 0.135456 $w=2.3e-07 $l=1.95e-07 $layer=MET1_cond $X=0.915 $Y=2.035
+ $X2=0.72 $Y2=2.035
r249 45 50 0.103375 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.355 $Y=2.035
+ $X2=5.5 $Y2=2.035
r250 45 46 4.2752 $w=1.7e-07 $l=4.44e-06 $layer=MET1_cond $X=5.355 $Y=2.035
+ $X2=0.915 $Y2=2.035
r251 43 74 18.5385 $w=3.9e-07 $l=1.3e-07 $layer=POLY_cond $X=11.95 $Y=1.475
+ $X2=12.08 $Y2=1.475
r252 43 71 42.7811 $w=3.9e-07 $l=3e-07 $layer=POLY_cond $X=11.95 $Y=1.475
+ $X2=11.65 $Y2=1.475
r253 42 43 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=11.95
+ $Y=1.445 $X2=11.95 $Y2=1.445
r254 39 54 14.0297 $w=3.43e-07 $l=4.2e-07 $layer=LI1_cond $X=11.882 $Y=1.615
+ $X2=11.882 $Y2=2.035
r255 39 42 2.70228 $w=2.88e-07 $l=6.8e-08 $layer=LI1_cond $X=11.882 $Y=1.47
+ $X2=11.95 $Y2=1.47
r256 37 59 34.9723 $w=3.3e-07 $l=2e-07 $layer=POLY_cond $X=5.71 $Y=1.93 $X2=5.51
+ $Y2=1.93
r257 33 74 25.2441 $w=1.5e-07 $l=1.95e-07 $layer=POLY_cond $X=12.08 $Y=1.67
+ $X2=12.08 $Y2=1.475
r258 33 35 407.649 $w=1.5e-07 $l=7.95e-07 $layer=POLY_cond $X=12.08 $Y=1.67
+ $X2=12.08 $Y2=2.465
r259 29 71 25.2441 $w=1.5e-07 $l=1.95e-07 $layer=POLY_cond $X=11.65 $Y=1.67
+ $X2=11.65 $Y2=1.475
r260 29 31 407.649 $w=1.5e-07 $l=7.95e-07 $layer=POLY_cond $X=11.65 $Y=1.67
+ $X2=11.65 $Y2=2.465
r261 25 37 32.1775 $w=3.3e-07 $l=1.98997e-07 $layer=POLY_cond $X=5.785 $Y=2.095
+ $X2=5.71 $Y2=1.93
r262 25 27 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=5.785 $Y=2.095
+ $X2=5.785 $Y2=2.675
r263 21 70 21.0057 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.755 $Y=1.25
+ $X2=1.755 $Y2=1.415
r264 21 23 305.096 $w=1.5e-07 $l=5.95e-07 $layer=POLY_cond $X=1.755 $Y=1.25
+ $X2=1.755 $Y2=0.655
r265 17 69 21.0057 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.325 $Y=1.25
+ $X2=1.325 $Y2=1.415
r266 17 19 305.096 $w=1.5e-07 $l=5.95e-07 $layer=POLY_cond $X=1.325 $Y=1.25
+ $X2=1.325 $Y2=0.655
r267 13 68 21.0057 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.065 $Y=1.58
+ $X2=1.065 $Y2=1.415
r268 13 15 612.755 $w=1.5e-07 $l=1.195e-06 $layer=POLY_cond $X=1.065 $Y=1.58
+ $X2=1.065 $Y2=2.775
r269 9 67 21.0057 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.835 $Y=1.25
+ $X2=0.835 $Y2=1.415
r270 9 11 412.777 $w=1.5e-07 $l=8.05e-07 $layer=POLY_cond $X=0.835 $Y=1.25
+ $X2=0.835 $Y2=0.445
r271 5 63 9.13417 $w=2.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.525 $Y=1.58
+ $X2=0.525 $Y2=1.415
r272 5 7 252.18 $w=2.5e-07 $l=1.015e-06 $layer=POLY_cond $X=0.525 $Y=1.58
+ $X2=0.525 $Y2=2.595
r273 1 62 21.0057 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=1.25
+ $X2=0.475 $Y2=1.415
r274 1 3 412.777 $w=1.5e-07 $l=8.05e-07 $layer=POLY_cond $X=0.475 $Y=1.25
+ $X2=0.475 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__BUSDRIVERNOVLPSLEEP_20%TE_B 3 5 6 8 11 15 17 25
r59 23 25 54.1518 $w=3.8e-07 $l=3.7e-07 $layer=POLY_cond $X=2.245 $Y=1.395
+ $X2=2.615 $Y2=1.395
r60 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.245
+ $Y=1.42 $X2=2.245 $Y2=1.42
r61 21 23 8.78138 $w=3.8e-07 $l=6e-08 $layer=POLY_cond $X=2.185 $Y=1.395
+ $X2=2.245 $Y2=1.395
r62 19 21 4.39069 $w=3.8e-07 $l=3e-08 $layer=POLY_cond $X=2.155 $Y=1.395
+ $X2=2.185 $Y2=1.395
r63 17 24 3.79093 $w=3.78e-07 $l=1.25e-07 $layer=LI1_cond $X=2.225 $Y=1.295
+ $X2=2.225 $Y2=1.42
r64 13 25 24.6126 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=2.615 $Y=1.205
+ $X2=2.615 $Y2=1.395
r65 13 15 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=2.615 $Y=1.205
+ $X2=2.615 $Y2=0.655
r66 9 21 24.6126 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=2.185 $Y=1.205
+ $X2=2.185 $Y2=1.395
r67 9 11 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=2.185 $Y=1.205
+ $X2=2.185 $Y2=0.655
r68 7 19 24.6126 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=2.155 $Y=1.585
+ $X2=2.155 $Y2=1.395
r69 7 8 102.553 $w=1.5e-07 $l=2e-07 $layer=POLY_cond $X=2.155 $Y=1.585 $X2=2.155
+ $Y2=1.785
r70 5 8 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.08 $Y=1.86
+ $X2=2.155 $Y2=1.785
r71 5 6 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=2.08 $Y=1.86 $X2=1.5
+ $Y2=1.86
r72 1 6 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.425 $Y=1.935
+ $X2=1.5 $Y2=1.86
r73 1 3 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=1.425 $Y=1.935
+ $X2=1.425 $Y2=2.775
.ends

.subckt PM_SKY130_FD_SC_LP__BUSDRIVERNOVLPSLEEP_20%A_27_47# 1 2 9 13 15 16 22 26
+ 27 29
c88 27 0 4.91905e-20 $X=4.65 $Y=1.445
c89 22 0 2.93767e-19 $X=4.65 $Y=1.665
c90 15 0 1.60636e-20 $X=4.505 $Y=1.665
r91 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.65
+ $Y=1.445 $X2=4.65 $Y2=1.445
r92 23 27 7.68295 $w=3.28e-07 $l=2.2e-07 $layer=LI1_cond $X=4.65 $Y=1.665
+ $X2=4.65 $Y2=1.445
r93 22 23 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.65 $Y=1.665
+ $X2=4.65 $Y2=1.665
r94 19 33 31.6049 $w=3.28e-07 $l=9.05e-07 $layer=LI1_cond $X=0.26 $Y=1.665
+ $X2=0.26 $Y2=2.57
r95 19 29 43.4785 $w=3.28e-07 $l=1.245e-06 $layer=LI1_cond $X=0.26 $Y=1.665
+ $X2=0.26 $Y2=0.42
r96 18 19 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=1.665
+ $X2=0.24 $Y2=1.665
r97 16 18 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.385 $Y=1.665
+ $X2=0.24 $Y2=1.665
r98 15 22 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.505 $Y=1.665
+ $X2=4.65 $Y2=1.665
r99 15 16 5.099 $w=1.4e-07 $l=4.12e-06 $layer=MET1_cond $X=4.505 $Y=1.665
+ $X2=0.385 $Y2=1.665
r100 11 26 46.1532 $w=2.87e-07 $l=3.51426e-07 $layer=POLY_cond $X=4.835 $Y=1.705
+ $X2=4.62 $Y2=1.445
r101 11 13 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=4.835 $Y=1.705
+ $X2=4.835 $Y2=2.465
r102 7 26 46.1532 $w=2.87e-07 $l=3.51426e-07 $layer=POLY_cond $X=4.405 $Y=1.705
+ $X2=4.62 $Y2=1.445
r103 7 9 389.702 $w=1.5e-07 $l=7.6e-07 $layer=POLY_cond $X=4.405 $Y=1.705
+ $X2=4.405 $Y2=2.465
r104 2 33 300 $w=1.7e-07 $l=5.33854e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=2.095 $X2=0.26 $Y2=2.57
r105 1 29 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__BUSDRIVERNOVLPSLEEP_20%A_280_47# 1 2 3 12 14 15 17
+ 18 20 23 25 27 28 29 32 35 36 37 40 42 45 48 51 53 55 59 63 67 68
c179 68 0 6.74658e-20 $X=1.612 $Y=1.845
c180 40 0 1.02413e-19 $X=6.145 $Y=2.675
r181 72 73 31.6192 $w=6.25e-07 $l=4.1e-07 $layer=POLY_cond $X=3.565 $Y=1.317
+ $X2=3.975 $Y2=1.317
r182 71 72 8.8688 $w=6.25e-07 $l=1.15e-07 $layer=POLY_cond $X=3.45 $Y=1.317
+ $X2=3.565 $Y2=1.317
r183 64 71 29.6912 $w=6.25e-07 $l=3.85e-07 $layer=POLY_cond $X=3.065 $Y=1.317
+ $X2=3.45 $Y2=1.317
r184 64 69 6.9408 $w=6.25e-07 $l=9e-08 $layer=POLY_cond $X=3.065 $Y=1.317
+ $X2=2.975 $Y2=1.317
r185 63 64 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.065
+ $Y=1.51 $X2=3.065 $Y2=1.51
r186 61 63 10.8721 $w=2.63e-07 $l=2.5e-07 $layer=LI1_cond $X=3.032 $Y=1.76
+ $X2=3.032 $Y2=1.51
r187 57 59 20.6969 $w=2.43e-07 $l=4.4e-07 $layer=LI1_cond $X=2.427 $Y=0.86
+ $X2=2.427 $Y2=0.42
r188 56 68 3.01551 $w=1.7e-07 $l=1.93e-07 $layer=LI1_cond $X=1.805 $Y=1.845
+ $X2=1.612 $Y2=1.845
r189 55 61 7.24806 $w=1.7e-07 $l=1.69245e-07 $layer=LI1_cond $X=2.9 $Y=1.845
+ $X2=3.032 $Y2=1.76
r190 55 56 71.4385 $w=1.68e-07 $l=1.095e-06 $layer=LI1_cond $X=2.9 $Y=1.845
+ $X2=1.805 $Y2=1.845
r191 54 67 2.11342 $w=1.7e-07 $l=1.08e-07 $layer=LI1_cond $X=1.635 $Y=0.945
+ $X2=1.527 $Y2=0.945
r192 53 57 7.11011 $w=1.7e-07 $l=1.58915e-07 $layer=LI1_cond $X=2.305 $Y=0.945
+ $X2=2.427 $Y2=0.86
r193 53 54 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.305 $Y=0.945
+ $X2=1.635 $Y2=0.945
r194 49 68 3.49088 $w=2.67e-07 $l=9.80051e-08 $layer=LI1_cond $X=1.64 $Y=1.93
+ $X2=1.612 $Y2=1.845
r195 49 51 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=1.64 $Y=1.93
+ $X2=1.64 $Y2=2.61
r196 48 68 3.49088 $w=2.67e-07 $l=1.25499e-07 $layer=LI1_cond $X=1.522 $Y=1.76
+ $X2=1.612 $Y2=1.845
r197 47 67 4.3182 $w=2.1e-07 $l=8.74643e-08 $layer=LI1_cond $X=1.522 $Y=1.03
+ $X2=1.527 $Y2=0.945
r198 47 48 39.4945 $w=2.03e-07 $l=7.3e-07 $layer=LI1_cond $X=1.522 $Y=1.03
+ $X2=1.522 $Y2=1.76
r199 43 67 4.3182 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=1.527 $Y=0.86
+ $X2=1.527 $Y2=0.945
r200 43 45 23.5849 $w=2.13e-07 $l=4.4e-07 $layer=LI1_cond $X=1.527 $Y=0.86
+ $X2=1.527 $Y2=0.42
r201 38 40 574.298 $w=1.5e-07 $l=1.12e-06 $layer=POLY_cond $X=6.145 $Y=1.555
+ $X2=6.145 $Y2=2.675
r202 36 38 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.07 $Y=1.48
+ $X2=6.145 $Y2=1.555
r203 36 37 412.777 $w=1.5e-07 $l=8.05e-07 $layer=POLY_cond $X=6.07 $Y=1.48
+ $X2=5.265 $Y2=1.48
r204 35 37 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.19 $Y=1.405
+ $X2=5.265 $Y2=1.48
r205 34 42 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.19 $Y=1.07
+ $X2=5.19 $Y2=0.995
r206 34 35 171.777 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=5.19 $Y=1.07
+ $X2=5.19 $Y2=1.405
r207 30 42 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.19 $Y=0.92
+ $X2=5.19 $Y2=0.995
r208 30 32 243.564 $w=1.5e-07 $l=4.75e-07 $layer=POLY_cond $X=5.19 $Y=0.92
+ $X2=5.19 $Y2=0.445
r209 29 73 38.3143 $w=6.25e-07 $l=3.57539e-07 $layer=POLY_cond $X=4.05 $Y=0.995
+ $X2=3.975 $Y2=1.317
r210 28 42 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.115 $Y=0.995
+ $X2=5.19 $Y2=0.995
r211 28 29 546.096 $w=1.5e-07 $l=1.065e-06 $layer=POLY_cond $X=5.115 $Y=0.995
+ $X2=4.05 $Y2=0.995
r212 25 73 37.1359 $w=1.5e-07 $l=3.98e-07 $layer=POLY_cond $X=3.975 $Y=1.715
+ $X2=3.975 $Y2=1.317
r213 25 27 241 $w=1.5e-07 $l=7.5e-07 $layer=POLY_cond $X=3.975 $Y=1.715
+ $X2=3.975 $Y2=2.465
r214 21 72 37.1359 $w=1.5e-07 $l=3.97e-07 $layer=POLY_cond $X=3.565 $Y=0.92
+ $X2=3.565 $Y2=1.317
r215 21 23 243.564 $w=1.5e-07 $l=4.75e-07 $layer=POLY_cond $X=3.565 $Y=0.92
+ $X2=3.565 $Y2=0.445
r216 18 71 37.1359 $w=1.5e-07 $l=3.98e-07 $layer=POLY_cond $X=3.45 $Y=1.715
+ $X2=3.45 $Y2=1.317
r217 18 20 241 $w=1.5e-07 $l=7.5e-07 $layer=POLY_cond $X=3.45 $Y=1.715 $X2=3.45
+ $Y2=2.465
r218 16 69 37.1359 $w=1.5e-07 $l=3.98e-07 $layer=POLY_cond $X=2.975 $Y=1.715
+ $X2=2.975 $Y2=1.317
r219 16 17 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=2.975 $Y=1.715
+ $X2=2.975 $Y2=2.145
r220 14 17 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.9 $Y=2.22
+ $X2=2.975 $Y2=2.145
r221 14 15 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=2.9 $Y=2.22
+ $X2=2.45 $Y2=2.22
r222 10 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.375 $Y=2.295
+ $X2=2.45 $Y2=2.22
r223 10 12 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.375 $Y=2.295
+ $X2=2.375 $Y2=2.775
r224 3 51 300 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_PDIFF $count=2 $X=1.5
+ $Y=2.455 $X2=1.64 $Y2=2.61
r225 2 59 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=2.26
+ $Y=0.235 $X2=2.4 $Y2=0.42
r226 1 67 182 $w=1.7e-07 $l=7.81873e-07 $layer=licon1_NDIFF $count=1 $X=1.4
+ $Y=0.235 $X2=1.54 $Y2=0.95
r227 1 45 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=1.4
+ $Y=0.235 $X2=1.54 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__BUSDRIVERNOVLPSLEEP_20%A_705_367# 1 2 3 12 14 15 17
+ 18 20 22 24 25 26 27 29 30 32 34 35 37 39 40 42 44 45 47 49 50 52 54 55 57 59
+ 60 62 64 65 67 69 70 72 74 75 77 79 80 82 83 85 86 88 89 91 92 94 95 97 98 100
+ 101 103 104 105 106 107 108 109 110 111 112 113 116 120 121 123 125 128 130
+ 131 134 137 138 140 143 144 148 159 164 172 177 182 187 188 205
c554 144 0 3.14657e-19 $X=6.625 $Y=1.665
c555 143 0 1.29574e-19 $X=14.5 $Y=1.665
c556 104 0 6.17609e-20 $X=14.84 $Y=1.65
c557 26 0 3.58277e-20 $X=14.485 $Y=1.65
c558 17 0 1.51872e-19 $X=6.505 $Y=1.575
r559 187 189 40.8145 $w=3.72e-07 $l=3.15e-07 $layer=POLY_cond $X=22.265 $Y=1.535
+ $X2=22.58 $Y2=1.535
r560 187 188 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=22.265
+ $Y=1.51 $X2=22.265 $Y2=1.51
r561 185 187 14.9005 $w=3.72e-07 $l=1.15e-07 $layer=POLY_cond $X=22.15 $Y=1.535
+ $X2=22.265 $Y2=1.535
r562 184 185 55.7151 $w=3.72e-07 $l=4.3e-07 $layer=POLY_cond $X=21.72 $Y=1.535
+ $X2=22.15 $Y2=1.535
r563 183 184 55.7151 $w=3.72e-07 $l=4.3e-07 $layer=POLY_cond $X=21.29 $Y=1.535
+ $X2=21.72 $Y2=1.535
r564 181 183 29.1532 $w=3.72e-07 $l=2.25e-07 $layer=POLY_cond $X=21.065 $Y=1.535
+ $X2=21.29 $Y2=1.535
r565 181 182 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=21.065
+ $Y=1.51 $X2=21.065 $Y2=1.51
r566 179 181 26.5618 $w=3.72e-07 $l=2.05e-07 $layer=POLY_cond $X=20.86 $Y=1.535
+ $X2=21.065 $Y2=1.535
r567 178 179 55.7151 $w=3.72e-07 $l=4.3e-07 $layer=POLY_cond $X=20.43 $Y=1.535
+ $X2=20.86 $Y2=1.535
r568 176 178 29.1532 $w=3.72e-07 $l=2.25e-07 $layer=POLY_cond $X=20.205 $Y=1.535
+ $X2=20.43 $Y2=1.535
r569 176 177 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=20.205
+ $Y=1.51 $X2=20.205 $Y2=1.51
r570 174 176 26.5618 $w=3.72e-07 $l=2.05e-07 $layer=POLY_cond $X=20 $Y=1.535
+ $X2=20.205 $Y2=1.535
r571 173 174 55.7151 $w=3.72e-07 $l=4.3e-07 $layer=POLY_cond $X=19.57 $Y=1.535
+ $X2=20 $Y2=1.535
r572 171 173 29.1532 $w=3.72e-07 $l=2.25e-07 $layer=POLY_cond $X=19.345 $Y=1.535
+ $X2=19.57 $Y2=1.535
r573 171 172 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=19.345
+ $Y=1.51 $X2=19.345 $Y2=1.51
r574 164 205 7.84979 $w=3.53e-07 $l=1.45e-07 $layer=LI1_cond $X=6.48 $Y=1.727
+ $X2=6.335 $Y2=1.727
r575 164 167 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.595
+ $Y=1.74 $X2=6.595 $Y2=1.74
r576 163 164 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=1.665
+ $X2=6.48 $Y2=1.665
r577 159 188 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=22.285 $Y=1.665
+ $X2=22.285 $Y2=1.665
r578 156 159 0.782757 $w=2.3e-07 $l=1.22e-06 $layer=MET1_cond $X=21.065 $Y=1.665
+ $X2=22.285 $Y2=1.665
r579 156 182 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=21.065 $Y=1.665
+ $X2=21.065 $Y2=1.665
r580 153 156 0.55178 $w=2.3e-07 $l=8.6e-07 $layer=MET1_cond $X=20.205 $Y=1.665
+ $X2=21.065 $Y2=1.665
r581 153 177 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=20.205 $Y=1.665
+ $X2=20.205 $Y2=1.665
r582 150 153 0.55178 $w=2.3e-07 $l=8.6e-07 $layer=MET1_cond $X=19.345 $Y=1.665
+ $X2=20.205 $Y2=1.665
r583 150 172 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=19.345 $Y=1.665
+ $X2=19.345 $Y2=1.665
r584 147 150 2.99308 $w=2.3e-07 $l=4.665e-06 $layer=MET1_cond $X=14.68 $Y=1.665
+ $X2=19.345 $Y2=1.665
r585 147 148 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.68 $Y=1.665
+ $X2=14.68 $Y2=1.665
r586 145 147 0.0384963 $w=2.3e-07 $l=6e-08 $layer=MET1_cond $X=14.62 $Y=1.665
+ $X2=14.68 $Y2=1.665
r587 144 163 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.625 $Y=1.665
+ $X2=6.48 $Y2=1.665
r588 143 145 0.0657895 $w=2.28e-07 $l=1.2e-07 $layer=MET1_cond $X=14.5 $Y=1.665
+ $X2=14.62 $Y2=1.665
r589 143 144 9.74627 $w=1.4e-07 $l=7.875e-06 $layer=MET1_cond $X=14.5 $Y=1.665
+ $X2=6.625 $Y2=1.665
r590 140 148 15.5329 $w=2.28e-07 $l=3.1e-07 $layer=LI1_cond $X=14.37 $Y=1.665
+ $X2=14.68 $Y2=1.665
r591 140 141 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=14.285 $Y=1.665
+ $X2=14.285 $Y2=1.87
r592 137 140 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=14.285 $Y=1.55
+ $X2=14.285 $Y2=1.665
r593 137 138 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=14.285 $Y=1.55
+ $X2=14.285 $Y2=1.095
r594 132 138 7.79447 $w=2.93e-07 $l=1.47e-07 $layer=LI1_cond $X=14.222 $Y=0.948
+ $X2=14.222 $Y2=1.095
r595 132 134 5.19576 $w=2.93e-07 $l=1.33e-07 $layer=LI1_cond $X=14.222 $Y=0.948
+ $X2=14.222 $Y2=0.815
r596 130 141 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=14.2 $Y=1.87
+ $X2=14.285 $Y2=1.87
r597 130 131 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=14.2 $Y=1.87
+ $X2=13.41 $Y2=1.87
r598 126 131 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=13.28 $Y=1.955
+ $X2=13.41 $Y2=1.87
r599 126 128 1.10812 $w=2.58e-07 $l=2.5e-08 $layer=LI1_cond $X=13.28 $Y=1.955
+ $X2=13.28 $Y2=1.98
r600 125 205 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=6.015 $Y=1.635
+ $X2=6.335 $Y2=1.635
r601 123 125 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.93 $Y=1.55
+ $X2=6.015 $Y2=1.635
r602 122 123 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=5.93 $Y=1.155
+ $X2=5.93 $Y2=1.55
r603 120 122 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.845 $Y=1.07
+ $X2=5.93 $Y2=1.155
r604 120 121 127.219 $w=1.68e-07 $l=1.95e-06 $layer=LI1_cond $X=5.845 $Y=1.07
+ $X2=3.895 $Y2=1.07
r605 116 118 49.2407 $w=2.18e-07 $l=9.4e-07 $layer=LI1_cond $X=3.785 $Y=1.96
+ $X2=3.785 $Y2=2.9
r606 114 121 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=3.785 $Y=1.155
+ $X2=3.895 $Y2=1.07
r607 114 116 42.1689 $w=2.18e-07 $l=8.05e-07 $layer=LI1_cond $X=3.785 $Y=1.155
+ $X2=3.785 $Y2=1.96
r608 101 189 24.0971 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=22.58 $Y=1.725
+ $X2=22.58 $Y2=1.535
r609 101 103 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=22.58 $Y=1.725
+ $X2=22.58 $Y2=2.465
r610 98 185 24.0971 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=22.15 $Y=1.725
+ $X2=22.15 $Y2=1.535
r611 98 100 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=22.15 $Y=1.725
+ $X2=22.15 $Y2=2.465
r612 95 184 24.0971 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=21.72 $Y=1.725
+ $X2=21.72 $Y2=1.535
r613 95 97 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=21.72 $Y=1.725
+ $X2=21.72 $Y2=2.465
r614 92 183 24.0971 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=21.29 $Y=1.725
+ $X2=21.29 $Y2=1.535
r615 92 94 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=21.29 $Y=1.725
+ $X2=21.29 $Y2=2.465
r616 89 179 24.0971 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=20.86 $Y=1.725
+ $X2=20.86 $Y2=1.535
r617 89 91 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=20.86 $Y=1.725
+ $X2=20.86 $Y2=2.465
r618 86 178 24.0971 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=20.43 $Y=1.725
+ $X2=20.43 $Y2=1.535
r619 86 88 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=20.43 $Y=1.725
+ $X2=20.43 $Y2=2.465
r620 83 174 24.0971 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=20 $Y=1.725 $X2=20
+ $Y2=1.535
r621 83 85 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=20 $Y=1.725 $X2=20
+ $Y2=2.465
r622 80 173 24.0971 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=19.57 $Y=1.725
+ $X2=19.57 $Y2=1.535
r623 80 82 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=19.57 $Y=1.725
+ $X2=19.57 $Y2=2.465
r624 77 171 26.5618 $w=3.72e-07 $l=2.84561e-07 $layer=POLY_cond $X=19.14
+ $Y=1.725 $X2=19.345 $Y2=1.535
r625 77 79 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=19.14 $Y=1.725
+ $X2=19.14 $Y2=2.465
r626 76 113 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=18.785 $Y=1.65
+ $X2=18.71 $Y2=1.65
r627 75 77 27.4257 $w=3.72e-07 $l=1.06066e-07 $layer=POLY_cond $X=19.065 $Y=1.65
+ $X2=19.14 $Y2=1.725
r628 75 76 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=19.065 $Y=1.65
+ $X2=18.785 $Y2=1.65
r629 72 113 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=18.71 $Y=1.725
+ $X2=18.71 $Y2=1.65
r630 72 74 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=18.71 $Y=1.725
+ $X2=18.71 $Y2=2.465
r631 71 112 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=18.355 $Y=1.65
+ $X2=18.28 $Y2=1.65
r632 70 113 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=18.635 $Y=1.65
+ $X2=18.71 $Y2=1.65
r633 70 71 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=18.635 $Y=1.65
+ $X2=18.355 $Y2=1.65
r634 67 112 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=18.28 $Y=1.725
+ $X2=18.28 $Y2=1.65
r635 67 69 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=18.28 $Y=1.725
+ $X2=18.28 $Y2=2.465
r636 66 111 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=17.925 $Y=1.65
+ $X2=17.85 $Y2=1.65
r637 65 112 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=18.205 $Y=1.65
+ $X2=18.28 $Y2=1.65
r638 65 66 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=18.205 $Y=1.65
+ $X2=17.925 $Y2=1.65
r639 62 111 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=17.85 $Y=1.725
+ $X2=17.85 $Y2=1.65
r640 62 64 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=17.85 $Y=1.725
+ $X2=17.85 $Y2=2.465
r641 61 110 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=17.495 $Y=1.65
+ $X2=17.42 $Y2=1.65
r642 60 111 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=17.775 $Y=1.65
+ $X2=17.85 $Y2=1.65
r643 60 61 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=17.775 $Y=1.65
+ $X2=17.495 $Y2=1.65
r644 57 110 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=17.42 $Y=1.725
+ $X2=17.42 $Y2=1.65
r645 57 59 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=17.42 $Y=1.725
+ $X2=17.42 $Y2=2.465
r646 56 109 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=17.065 $Y=1.65
+ $X2=16.99 $Y2=1.65
r647 55 110 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=17.345 $Y=1.65
+ $X2=17.42 $Y2=1.65
r648 55 56 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=17.345 $Y=1.65
+ $X2=17.065 $Y2=1.65
r649 52 109 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=16.99 $Y=1.725
+ $X2=16.99 $Y2=1.65
r650 52 54 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=16.99 $Y=1.725
+ $X2=16.99 $Y2=2.465
r651 51 108 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=16.635 $Y=1.65
+ $X2=16.56 $Y2=1.65
r652 50 109 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=16.915 $Y=1.65
+ $X2=16.99 $Y2=1.65
r653 50 51 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=16.915 $Y=1.65
+ $X2=16.635 $Y2=1.65
r654 47 108 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=16.56 $Y=1.725
+ $X2=16.56 $Y2=1.65
r655 47 49 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=16.56 $Y=1.725
+ $X2=16.56 $Y2=2.465
r656 46 107 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=16.205 $Y=1.65
+ $X2=16.13 $Y2=1.65
r657 45 108 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=16.485 $Y=1.65
+ $X2=16.56 $Y2=1.65
r658 45 46 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=16.485 $Y=1.65
+ $X2=16.205 $Y2=1.65
r659 42 107 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=16.13 $Y=1.725
+ $X2=16.13 $Y2=1.65
r660 42 44 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=16.13 $Y=1.725
+ $X2=16.13 $Y2=2.465
r661 41 106 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=15.775 $Y=1.65
+ $X2=15.7 $Y2=1.65
r662 40 107 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=16.055 $Y=1.65
+ $X2=16.13 $Y2=1.65
r663 40 41 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=16.055 $Y=1.65
+ $X2=15.775 $Y2=1.65
r664 37 106 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=15.7 $Y=1.725
+ $X2=15.7 $Y2=1.65
r665 37 39 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=15.7 $Y=1.725
+ $X2=15.7 $Y2=2.465
r666 36 105 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=15.345 $Y=1.65
+ $X2=15.27 $Y2=1.65
r667 35 106 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=15.625 $Y=1.65
+ $X2=15.7 $Y2=1.65
r668 35 36 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=15.625 $Y=1.65
+ $X2=15.345 $Y2=1.65
r669 32 105 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=15.27 $Y=1.725
+ $X2=15.27 $Y2=1.65
r670 32 34 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=15.27 $Y=1.725
+ $X2=15.27 $Y2=2.465
r671 31 104 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=14.915 $Y=1.65
+ $X2=14.84 $Y2=1.65
r672 30 105 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=15.195 $Y=1.65
+ $X2=15.27 $Y2=1.65
r673 30 31 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=15.195 $Y=1.65
+ $X2=14.915 $Y2=1.65
r674 27 104 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=14.84 $Y=1.725
+ $X2=14.84 $Y2=1.65
r675 27 29 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=14.84 $Y=1.725
+ $X2=14.84 $Y2=2.465
r676 25 104 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=14.765 $Y=1.65
+ $X2=14.84 $Y2=1.65
r677 25 26 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=14.765 $Y=1.65
+ $X2=14.485 $Y2=1.65
r678 22 26 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=14.41 $Y=1.725
+ $X2=14.485 $Y2=1.65
r679 22 24 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=14.41 $Y=1.725
+ $X2=14.41 $Y2=2.465
r680 18 167 39.3224 $w=3.28e-07 $l=1.79722e-07 $layer=POLY_cond $X=6.575 $Y=1.91
+ $X2=6.595 $Y2=1.74
r681 18 20 392.266 $w=1.5e-07 $l=7.65e-07 $layer=POLY_cond $X=6.575 $Y=1.91
+ $X2=6.575 $Y2=2.675
r682 17 167 38.5876 $w=3.28e-07 $l=2.05122e-07 $layer=POLY_cond $X=6.505
+ $Y=1.575 $X2=6.595 $Y2=1.74
r683 16 17 194.851 $w=1.5e-07 $l=3.8e-07 $layer=POLY_cond $X=6.505 $Y=1.195
+ $X2=6.505 $Y2=1.575
r684 14 16 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.43 $Y=1.12
+ $X2=6.505 $Y2=1.195
r685 14 15 412.777 $w=1.5e-07 $l=8.05e-07 $layer=POLY_cond $X=6.43 $Y=1.12
+ $X2=5.625 $Y2=1.12
r686 10 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.55 $Y=1.045
+ $X2=5.625 $Y2=1.12
r687 10 12 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=5.55 $Y=1.045 $X2=5.55
+ $Y2=0.445
r688 3 128 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=13.105
+ $Y=1.835 $X2=13.245 $Y2=1.98
r689 2 118 400 $w=1.7e-07 $l=1.17665e-06 $layer=licon1_PDIFF $count=1 $X=3.525
+ $Y=1.835 $X2=3.76 $Y2=2.9
r690 2 116 400 $w=1.7e-07 $l=2.90861e-07 $layer=licon1_PDIFF $count=1 $X=3.525
+ $Y=1.835 $X2=3.76 $Y2=1.96
r691 1 134 182 $w=1.7e-07 $l=6.4622e-07 $layer=licon1_NDIFF $count=1 $X=14.03
+ $Y=0.235 $X2=14.17 $Y2=0.815
.ends

.subckt PM_SKY130_FD_SC_LP__BUSDRIVERNOVLPSLEEP_20%A_407_491# 1 2 8 9 10 11 13
+ 14 16 18 19 21 25 27 28 31 33 34 35 36 37 41 42 46 48 49 51 52 53 55 56 57 64
+ 66
c214 64 0 3.00155e-20 $X=10.15 $Y=1.16
c215 21 0 1.20891e-19 $X=10.09 $Y=2.285
c216 19 0 1.91794e-19 $X=10.09 $Y=1.33
c217 14 0 7.24991e-20 $X=7.96 $Y=1.26
r218 64 66 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=10.15 $Y=1.16
+ $X2=10.15 $Y2=0.995
r219 64 65 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.15
+ $Y=1.16 $X2=10.15 $Y2=1.16
r220 61 62 13.5556 $w=2.61e-07 $l=2.9e-07 $layer=LI1_cond $X=3.345 $Y=0.44
+ $X2=3.345 $Y2=0.73
r221 58 66 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=10.07 $Y=0.825
+ $X2=10.07 $Y2=0.995
r222 56 58 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.985 $Y=0.74
+ $X2=10.07 $Y2=0.825
r223 56 57 113.519 $w=1.68e-07 $l=1.74e-06 $layer=LI1_cond $X=9.985 $Y=0.74
+ $X2=8.245 $Y2=0.74
r224 55 57 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.16 $Y=0.655
+ $X2=8.245 $Y2=0.74
r225 54 55 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=8.16 $Y=0.435
+ $X2=8.16 $Y2=0.655
r226 52 54 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.075 $Y=0.35
+ $X2=8.16 $Y2=0.435
r227 52 53 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=8.075 $Y=0.35
+ $X2=7.565 $Y2=0.35
r228 50 53 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.48 $Y=0.435
+ $X2=7.565 $Y2=0.35
r229 50 51 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=7.48 $Y=0.435
+ $X2=7.48 $Y2=0.85
r230 48 51 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.395 $Y=0.935
+ $X2=7.48 $Y2=0.85
r231 48 49 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=7.395 $Y=0.935
+ $X2=6.695 $Y2=0.935
r232 46 47 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.61
+ $Y=0.67 $X2=6.61 $Y2=0.67
r233 44 49 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.61 $Y=0.85
+ $X2=6.695 $Y2=0.935
r234 44 46 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=6.61 $Y=0.85
+ $X2=6.61 $Y2=0.67
r235 43 46 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=6.61 $Y=0.435
+ $X2=6.61 $Y2=0.67
r236 41 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.525 $Y=0.35
+ $X2=6.61 $Y2=0.435
r237 41 42 69.8075 $w=1.68e-07 $l=1.07e-06 $layer=LI1_cond $X=6.525 $Y=0.35
+ $X2=5.455 $Y2=0.35
r238 39 42 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.37 $Y=0.435
+ $X2=5.455 $Y2=0.35
r239 39 40 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=5.37 $Y=0.435
+ $X2=5.37 $Y2=0.645
r240 38 62 3.24614 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=3.505 $Y=0.73
+ $X2=3.345 $Y2=0.73
r241 37 40 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.285 $Y=0.73
+ $X2=5.37 $Y2=0.645
r242 37 38 116.128 $w=1.68e-07 $l=1.78e-06 $layer=LI1_cond $X=5.285 $Y=0.73
+ $X2=3.505 $Y2=0.73
r243 35 62 5.45457 $w=2.61e-07 $l=1.16619e-07 $layer=LI1_cond $X=3.42 $Y=0.815
+ $X2=3.345 $Y2=0.73
r244 35 36 83.8342 $w=1.68e-07 $l=1.285e-06 $layer=LI1_cond $X=3.42 $Y=0.815
+ $X2=3.42 $Y2=2.1
r245 33 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.335 $Y=2.185
+ $X2=3.42 $Y2=2.1
r246 33 34 65.8931 $w=1.68e-07 $l=1.01e-06 $layer=LI1_cond $X=3.335 $Y=2.185
+ $X2=2.325 $Y2=2.185
r247 29 34 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.16 $Y=2.27
+ $X2=2.325 $Y2=2.185
r248 29 31 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=2.16 $Y=2.27
+ $X2=2.16 $Y2=2.61
r249 27 47 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=6.79 $Y=0.67
+ $X2=6.61 $Y2=0.67
r250 23 65 38.5938 $w=3.29e-07 $l=2.05122e-07 $layer=POLY_cond $X=10.24 $Y=0.995
+ $X2=10.15 $Y2=1.16
r251 23 25 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=10.24 $Y=0.995
+ $X2=10.24 $Y2=0.445
r252 19 65 39.3263 $w=3.29e-07 $l=1.97737e-07 $layer=POLY_cond $X=10.09 $Y=1.33
+ $X2=10.15 $Y2=1.16
r253 19 21 489.691 $w=1.5e-07 $l=9.55e-07 $layer=POLY_cond $X=10.09 $Y=1.33
+ $X2=10.09 $Y2=2.285
r254 16 18 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=8.035 $Y=1.185
+ $X2=8.035 $Y2=0.655
r255 15 28 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.43 $Y=1.26
+ $X2=7.355 $Y2=1.26
r256 14 16 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.96 $Y=1.26
+ $X2=8.035 $Y2=1.185
r257 14 15 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=7.96 $Y=1.26
+ $X2=7.43 $Y2=1.26
r258 11 28 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.355 $Y=1.185
+ $X2=7.355 $Y2=1.26
r259 11 13 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=7.355 $Y=1.185
+ $X2=7.355 $Y2=0.655
r260 9 28 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.28 $Y=1.26
+ $X2=7.355 $Y2=1.26
r261 9 10 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=7.28 $Y=1.26 $X2=6.94
+ $Y2=1.26
r262 8 10 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.865 $Y=1.185
+ $X2=6.94 $Y2=1.26
r263 7 27 32.1775 $w=3.3e-07 $l=1.98997e-07 $layer=POLY_cond $X=6.865 $Y=0.835
+ $X2=6.79 $Y2=0.67
r264 7 8 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=6.865 $Y=0.835
+ $X2=6.865 $Y2=1.185
r265 2 31 300 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_PDIFF $count=2 $X=2.035
+ $Y=2.455 $X2=2.16 $Y2=2.61
r266 1 61 182 $w=1.7e-07 $l=2.60096e-07 $layer=licon1_NDIFF $count=1 $X=3.225
+ $Y=0.235 $X2=3.35 $Y2=0.44
.ends

.subckt PM_SKY130_FD_SC_LP__BUSDRIVERNOVLPSLEEP_20%A_896_367# 1 2 3 10 12 14 15
+ 17 19 20 23 25 27 32 35 36 37 42 45 48 52 53
c155 48 0 3.35109e-19 $X=6.36 $Y=2.17
c156 45 0 2.01956e-19 $X=4.62 $Y=2.225
c157 37 0 2.55807e-19 $X=6.97 $Y=2.17
c158 32 0 1.51872e-19 $X=6.27 $Y=1.2
c159 15 0 8.51739e-20 $X=8.155 $Y=1.65
r160 51 52 0.349225 $w=3.28e-07 $l=1e-08 $layer=LI1_cond $X=6.36 $Y=2.4 $X2=6.36
+ $Y2=2.41
r161 48 51 8.03218 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=6.36 $Y=2.17
+ $X2=6.36 $Y2=2.4
r162 45 47 9.26965 $w=2.28e-07 $l=1.85e-07 $layer=LI1_cond $X=4.6 $Y=2.225
+ $X2=4.6 $Y2=2.41
r163 43 53 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=7.135 $Y=1.74
+ $X2=7.135 $Y2=1.65
r164 42 43 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.135
+ $Y=1.74 $X2=7.135 $Y2=1.74
r165 40 42 15.292 $w=2.58e-07 $l=3.45e-07 $layer=LI1_cond $X=7.1 $Y=2.085
+ $X2=7.1 $Y2=1.74
r166 39 42 16.4002 $w=2.58e-07 $l=3.7e-07 $layer=LI1_cond $X=7.1 $Y=1.37 $X2=7.1
+ $Y2=1.74
r167 38 48 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.525 $Y=2.17
+ $X2=6.36 $Y2=2.17
r168 37 40 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=6.97 $Y=2.17
+ $X2=7.1 $Y2=2.085
r169 37 38 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=6.97 $Y=2.17
+ $X2=6.525 $Y2=2.17
r170 35 39 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=6.97 $Y=1.285
+ $X2=7.1 $Y2=1.37
r171 35 36 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=6.97 $Y=1.285
+ $X2=6.355 $Y2=1.285
r172 32 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.27 $Y=1.2
+ $X2=6.355 $Y2=1.285
r173 31 32 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=6.27 $Y=0.815
+ $X2=6.27 $Y2=1.2
r174 27 31 6.91519 $w=2.1e-07 $l=1.41244e-07 $layer=LI1_cond $X=6.185 $Y=0.71
+ $X2=6.27 $Y2=0.815
r175 27 29 19.013 $w=2.08e-07 $l=3.6e-07 $layer=LI1_cond $X=6.185 $Y=0.71
+ $X2=5.825 $Y2=0.71
r176 26 47 2.50919 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=4.715 $Y=2.41
+ $X2=4.6 $Y2=2.41
r177 25 52 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.195 $Y=2.41
+ $X2=6.36 $Y2=2.41
r178 25 26 96.5562 $w=1.68e-07 $l=1.48e-06 $layer=LI1_cond $X=6.195 $Y=2.41
+ $X2=4.715 $Y2=2.41
r179 21 47 4.25903 $w=2.28e-07 $l=8.5e-08 $layer=LI1_cond $X=4.6 $Y=2.495
+ $X2=4.6 $Y2=2.41
r180 21 23 3.50744 $w=2.28e-07 $l=7e-08 $layer=LI1_cond $X=4.6 $Y=2.495 $X2=4.6
+ $Y2=2.565
r181 17 19 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=8.23 $Y=1.725
+ $X2=8.23 $Y2=2.465
r182 16 20 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.875 $Y=1.65
+ $X2=7.8 $Y2=1.65
r183 15 17 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.155 $Y=1.65
+ $X2=8.23 $Y2=1.725
r184 15 16 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=8.155 $Y=1.65
+ $X2=7.875 $Y2=1.65
r185 12 20 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.8 $Y=1.725
+ $X2=7.8 $Y2=1.65
r186 12 14 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=7.8 $Y=1.725
+ $X2=7.8 $Y2=2.465
r187 11 53 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.3 $Y=1.65
+ $X2=7.135 $Y2=1.65
r188 10 20 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.725 $Y=1.65
+ $X2=7.8 $Y2=1.65
r189 10 11 217.926 $w=1.5e-07 $l=4.25e-07 $layer=POLY_cond $X=7.725 $Y=1.65
+ $X2=7.3 $Y2=1.65
r190 3 51 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=6.22
+ $Y=2.255 $X2=6.36 $Y2=2.4
r191 2 45 600 $w=1.7e-07 $l=4.54643e-07 $layer=licon1_PDIFF $count=1 $X=4.48
+ $Y=1.835 $X2=4.62 $Y2=2.225
r192 2 23 300 $w=1.7e-07 $l=7.96932e-07 $layer=licon1_PDIFF $count=2 $X=4.48
+ $Y=1.835 $X2=4.62 $Y2=2.565
r193 1 29 182 $w=1.7e-07 $l=5.45917e-07 $layer=licon1_NDIFF $count=1 $X=5.625
+ $Y=0.235 $X2=5.825 $Y2=0.69
.ends

.subckt PM_SKY130_FD_SC_LP__BUSDRIVERNOVLPSLEEP_20%A_1486_47# 1 2 3 12 16 20 24
+ 28 32 34 36 37 39 40 42 43 45 46 47 48 50 51 53 55 56 58 60 61 63 65 66 68 70
+ 71 73 75 77 78 81 82 83 84 85 88 92 94 101 103 104 105 106 107 121 126 130 132
+ 134 137 142 147 152 157
c344 130 0 1.20377e-19 $X=10.57 $Y=1.295
c345 105 0 6.62192e-20 $X=14.92 $Y=1.295
c346 101 0 2.44822e-19 $X=8.11 $Y=1.11
c347 12 0 1.43917e-19 $X=10.45 $Y=2.285
r348 156 157 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=18.505
+ $Y=1.2 $X2=18.505 $Y2=1.2
r349 154 156 31.5262 $w=3.44e-07 $l=2.25e-07 $layer=POLY_cond $X=18.28 $Y=1.175
+ $X2=18.505 $Y2=1.175
r350 153 154 60.25 $w=3.44e-07 $l=4.3e-07 $layer=POLY_cond $X=17.85 $Y=1.175
+ $X2=18.28 $Y2=1.175
r351 151 153 28.7238 $w=3.44e-07 $l=2.05e-07 $layer=POLY_cond $X=17.645 $Y=1.175
+ $X2=17.85 $Y2=1.175
r352 151 152 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=17.645
+ $Y=1.2 $X2=17.645 $Y2=1.2
r353 149 151 31.5262 $w=3.44e-07 $l=2.25e-07 $layer=POLY_cond $X=17.42 $Y=1.175
+ $X2=17.645 $Y2=1.175
r354 146 147 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=16.765
+ $Y=1.2 $X2=16.765 $Y2=1.2
r355 141 142 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=15.925
+ $Y=1.2 $X2=15.925 $Y2=1.2
r356 136 137 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=15.065
+ $Y=1.2 $X2=15.065 $Y2=1.2
r357 134 136 97.9223 $w=3.3e-07 $l=5.6e-07 $layer=POLY_cond $X=15.625 $Y=1.2
+ $X2=15.065 $Y2=1.2
r358 130 132 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=10.69
+ $Y=1.16 $X2=10.69 $Y2=1.16
r359 129 130 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.57 $Y=1.295
+ $X2=10.57 $Y2=1.295
r360 125 126 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.6 $Y=1.295
+ $X2=9.6 $Y2=1.295
r361 121 157 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=18.505 $Y=1.295
+ $X2=18.505 $Y2=1.295
r362 118 121 0.55178 $w=2.3e-07 $l=8.6e-07 $layer=MET1_cond $X=17.645 $Y=1.295
+ $X2=18.505 $Y2=1.295
r363 118 152 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=17.645 $Y=1.295
+ $X2=17.645 $Y2=1.295
r364 115 118 0.55178 $w=2.3e-07 $l=8.6e-07 $layer=MET1_cond $X=16.785 $Y=1.295
+ $X2=17.645 $Y2=1.295
r365 115 147 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=16.785 $Y=1.295
+ $X2=16.785 $Y2=1.295
r366 112 115 0.55178 $w=2.3e-07 $l=8.6e-07 $layer=MET1_cond $X=15.925 $Y=1.295
+ $X2=16.785 $Y2=1.295
r367 112 142 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=15.925 $Y=1.295
+ $X2=15.925 $Y2=1.295
r368 109 112 0.55178 $w=2.3e-07 $l=8.6e-07 $layer=MET1_cond $X=15.065 $Y=1.295
+ $X2=15.925 $Y2=1.295
r369 109 137 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=15.065 $Y=1.295
+ $X2=15.065 $Y2=1.295
r370 107 109 0.0192481 $w=2.3e-07 $l=3e-08 $layer=MET1_cond $X=15.035 $Y=1.295
+ $X2=15.065 $Y2=1.295
r371 106 129 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=10.715 $Y=1.295
+ $X2=10.57 $Y2=1.295
r372 105 107 0.0850015 $w=2.3e-07 $l=1.15e-07 $layer=MET1_cond $X=14.92 $Y=1.295
+ $X2=15.035 $Y2=1.295
r373 105 106 5.2042 $w=1.4e-07 $l=4.205e-06 $layer=MET1_cond $X=14.92 $Y=1.295
+ $X2=10.715 $Y2=1.295
r374 104 125 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=9.745 $Y=1.295
+ $X2=9.6 $Y2=1.295
r375 103 129 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=10.425 $Y=1.295
+ $X2=10.57 $Y2=1.295
r376 103 104 0.841583 $w=1.4e-07 $l=6.8e-07 $layer=MET1_cond $X=10.425 $Y=1.295
+ $X2=9.745 $Y2=1.295
r377 102 126 5.16612 $w=2.88e-07 $l=1.3e-07 $layer=LI1_cond $X=9.6 $Y=1.165
+ $X2=9.6 $Y2=1.295
r378 100 101 5.5678 $w=2.28e-07 $l=9.5e-08 $layer=LI1_cond $X=8.015 $Y=1.11
+ $X2=8.11 $Y2=1.11
r379 98 100 9.77071 $w=2.28e-07 $l=1.95e-07 $layer=LI1_cond $X=7.82 $Y=1.11
+ $X2=8.015 $Y2=1.11
r380 97 101 62.9572 $w=1.68e-07 $l=9.65e-07 $layer=LI1_cond $X=9.075 $Y=1.08
+ $X2=8.11 $Y2=1.08
r381 94 102 7.43784 $w=1.7e-07 $l=1.8262e-07 $layer=LI1_cond $X=9.455 $Y=1.08
+ $X2=9.6 $Y2=1.165
r382 94 97 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=9.455 $Y=1.08
+ $X2=9.075 $Y2=1.08
r383 90 100 1.85809 $w=1.9e-07 $l=1.15e-07 $layer=LI1_cond $X=8.015 $Y=1.225
+ $X2=8.015 $Y2=1.11
r384 90 92 44.0718 $w=1.88e-07 $l=7.55e-07 $layer=LI1_cond $X=8.015 $Y=1.225
+ $X2=8.015 $Y2=1.98
r385 86 98 2.50919 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=7.82 $Y=0.995
+ $X2=7.82 $Y2=1.11
r386 86 88 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=7.82 $Y=0.995
+ $X2=7.82 $Y2=0.82
r387 80 132 38.6168 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=10.69 $Y=0.995
+ $X2=10.69 $Y2=1.16
r388 77 132 66.4473 $w=3.3e-07 $l=3.8e-07 $layer=POLY_cond $X=10.69 $Y=1.54
+ $X2=10.69 $Y2=1.16
r389 77 78 43.5886 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=10.615 $Y=1.54
+ $X2=10.615 $Y2=1.69
r390 73 75 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=21.29 $Y=0.985
+ $X2=21.29 $Y2=0.555
r391 72 85 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=20.935 $Y=1.06
+ $X2=20.86 $Y2=1.06
r392 71 73 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=21.215 $Y=1.06
+ $X2=21.29 $Y2=0.985
r393 71 72 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=21.215 $Y=1.06
+ $X2=20.935 $Y2=1.06
r394 68 85 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=20.86 $Y=0.985
+ $X2=20.86 $Y2=1.06
r395 68 70 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=20.86 $Y=0.985
+ $X2=20.86 $Y2=0.555
r396 67 84 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=20.505 $Y=1.06
+ $X2=20.43 $Y2=1.06
r397 66 85 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=20.785 $Y=1.06
+ $X2=20.86 $Y2=1.06
r398 66 67 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=20.785 $Y=1.06
+ $X2=20.505 $Y2=1.06
r399 63 84 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=20.43 $Y=0.985
+ $X2=20.43 $Y2=1.06
r400 63 65 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=20.43 $Y=0.985
+ $X2=20.43 $Y2=0.555
r401 62 83 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=20.075 $Y=1.06
+ $X2=20 $Y2=1.06
r402 61 84 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=20.355 $Y=1.06
+ $X2=20.43 $Y2=1.06
r403 61 62 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=20.355 $Y=1.06
+ $X2=20.075 $Y2=1.06
r404 58 83 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=20 $Y=0.985 $X2=20
+ $Y2=1.06
r405 58 60 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=20 $Y=0.985 $X2=20
+ $Y2=0.555
r406 57 82 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=19.645 $Y=1.06
+ $X2=19.57 $Y2=1.06
r407 56 83 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=19.925 $Y=1.06
+ $X2=20 $Y2=1.06
r408 56 57 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=19.925 $Y=1.06
+ $X2=19.645 $Y2=1.06
r409 53 82 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=19.57 $Y=0.985
+ $X2=19.57 $Y2=1.06
r410 53 55 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=19.57 $Y=0.985
+ $X2=19.57 $Y2=0.555
r411 52 81 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=19.215 $Y=1.06
+ $X2=19.14 $Y2=1.06
r412 51 82 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=19.495 $Y=1.06
+ $X2=19.57 $Y2=1.06
r413 51 52 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=19.495 $Y=1.06
+ $X2=19.215 $Y2=1.06
r414 48 81 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=19.14 $Y=0.985
+ $X2=19.14 $Y2=1.06
r415 48 50 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=19.14 $Y=0.985
+ $X2=19.14 $Y2=0.555
r416 46 81 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=19.065 $Y=1.06
+ $X2=19.14 $Y2=1.06
r417 46 47 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=19.065 $Y=1.06
+ $X2=18.785 $Y2=1.06
r418 43 47 26.108 $w=3.44e-07 $l=1.06066e-07 $layer=POLY_cond $X=18.71 $Y=0.985
+ $X2=18.785 $Y2=1.06
r419 43 156 28.7238 $w=3.44e-07 $l=2.84561e-07 $layer=POLY_cond $X=18.71
+ $Y=0.985 $X2=18.505 $Y2=1.175
r420 43 45 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=18.71 $Y=0.985
+ $X2=18.71 $Y2=0.555
r421 40 154 22.2144 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=18.28 $Y=0.985
+ $X2=18.28 $Y2=1.175
r422 40 42 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=18.28 $Y=0.985
+ $X2=18.28 $Y2=0.555
r423 37 153 22.2144 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=17.85 $Y=0.985
+ $X2=17.85 $Y2=1.175
r424 37 39 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=17.85 $Y=0.985
+ $X2=17.85 $Y2=0.555
r425 34 149 22.2144 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=17.42 $Y=0.985
+ $X2=17.42 $Y2=1.175
r426 34 36 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=17.42 $Y=0.985
+ $X2=17.42 $Y2=0.555
r427 30 149 60.25 $w=3.44e-07 $l=4.3e-07 $layer=POLY_cond $X=16.99 $Y=1.175
+ $X2=17.42 $Y2=1.175
r428 30 146 31.5262 $w=3.44e-07 $l=2.25e-07 $layer=POLY_cond $X=16.99 $Y=1.175
+ $X2=16.765 $Y2=1.175
r429 30 32 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=16.99 $Y=1.035
+ $X2=16.99 $Y2=0.555
r430 26 146 28.7238 $w=3.44e-07 $l=2.05e-07 $layer=POLY_cond $X=16.56 $Y=1.175
+ $X2=16.765 $Y2=1.175
r431 26 28 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=16.56 $Y=1.035
+ $X2=16.56 $Y2=0.555
r432 22 26 60.25 $w=3.44e-07 $l=4.3e-07 $layer=POLY_cond $X=16.13 $Y=1.175
+ $X2=16.56 $Y2=1.175
r433 22 141 28.7238 $w=3.44e-07 $l=2.05e-07 $layer=POLY_cond $X=16.13 $Y=1.175
+ $X2=15.925 $Y2=1.175
r434 22 24 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=16.13 $Y=1.035
+ $X2=16.13 $Y2=0.555
r435 18 141 31.5262 $w=3.44e-07 $l=2.25e-07 $layer=POLY_cond $X=15.7 $Y=1.175
+ $X2=15.925 $Y2=1.175
r436 18 134 10.5087 $w=3.44e-07 $l=8.66025e-08 $layer=POLY_cond $X=15.7 $Y=1.175
+ $X2=15.625 $Y2=1.2
r437 18 20 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=15.7 $Y=1.035
+ $X2=15.7 $Y2=0.555
r438 16 80 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=10.67 $Y=0.445
+ $X2=10.67 $Y2=0.995
r439 12 78 305.096 $w=1.5e-07 $l=5.95e-07 $layer=POLY_cond $X=10.45 $Y=2.285
+ $X2=10.45 $Y2=1.69
r440 3 92 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=7.875
+ $Y=1.835 $X2=8.015 $Y2=1.98
r441 2 97 182 $w=1.7e-07 $l=9.4194e-07 $layer=licon1_NDIFF $count=1 $X=8.87
+ $Y=0.235 $X2=9.075 $Y2=1.08
r442 1 88 182 $w=1.7e-07 $l=7.55232e-07 $layer=licon1_NDIFF $count=1 $X=7.43
+ $Y=0.235 $X2=7.82 $Y2=0.82
.ends

.subckt PM_SKY130_FD_SC_LP__BUSDRIVERNOVLPSLEEP_20%A 1 3 6 8 10 13 16 17 18 20
+ 24 26 27 28 31 33 35 36 40 42 44 48 50 51 52 53 54 55 56 57 58
c218 52 0 1.0911e-19 $X=11.647 $Y=0.687
c219 51 0 2.29614e-19 $X=11.15 $Y=1.725
c220 42 0 1.12422e-19 $X=13.46 $Y=1.725
c221 28 0 9.84968e-20 $X=12.515 $Y=1.65
r222 58 62 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=12.22
+ $Y=0.605 $X2=12.22 $Y2=0.605
r223 57 58 16.0644 $w=3.28e-07 $l=4.6e-07 $layer=LI1_cond $X=11.76 $Y=0.605
+ $X2=12.22 $Y2=0.605
r224 54 62 15.6726 $w=4.95e-07 $l=1.45e-07 $layer=POLY_cond $X=12.365 $Y=0.687
+ $X2=12.22 $Y2=0.687
r225 52 62 61.9337 $w=4.95e-07 $l=5.73e-07 $layer=POLY_cond $X=11.647 $Y=0.687
+ $X2=12.22 $Y2=0.687
r226 52 53 55.2585 $w=4.95e-07 $l=2.47e-07 $layer=POLY_cond $X=11.647 $Y=0.687
+ $X2=11.4 $Y2=0.687
r227 50 51 63.4211 $w=1.7e-07 $l=1.5e-07 $layer=POLY_cond $X=11.15 $Y=1.575
+ $X2=11.15 $Y2=1.725
r228 47 48 54.4194 $w=2.79e-07 $l=3.15e-07 $layer=POLY_cond $X=9.09 $Y=1.562
+ $X2=9.405 $Y2=1.562
r229 46 47 50.9642 $w=2.79e-07 $l=2.95e-07 $layer=POLY_cond $X=8.795 $Y=1.562
+ $X2=9.09 $Y2=1.562
r230 45 46 23.3226 $w=2.79e-07 $l=1.35e-07 $layer=POLY_cond $X=8.66 $Y=1.562
+ $X2=8.795 $Y2=1.562
r231 42 56 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=13.46 $Y=1.725
+ $X2=13.46 $Y2=1.65
r232 42 44 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=13.46 $Y=1.725
+ $X2=13.46 $Y2=2.465
r233 38 56 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=13.46 $Y=1.575
+ $X2=13.46 $Y2=1.65
r234 38 40 471.745 $w=1.5e-07 $l=9.2e-07 $layer=POLY_cond $X=13.46 $Y=1.575
+ $X2=13.46 $Y2=0.655
r235 37 55 12.05 $w=1.5e-07 $l=1.23e-07 $layer=POLY_cond $X=13.105 $Y=1.65
+ $X2=12.982 $Y2=1.65
r236 36 56 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=13.385 $Y=1.65
+ $X2=13.46 $Y2=1.65
r237 36 37 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=13.385 $Y=1.65
+ $X2=13.105 $Y2=1.65
r238 33 55 12.05 $w=1.5e-07 $l=9.60469e-08 $layer=POLY_cond $X=13.03 $Y=1.725
+ $X2=12.982 $Y2=1.65
r239 33 35 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=13.03 $Y=1.725
+ $X2=13.03 $Y2=2.465
r240 29 55 12.05 $w=1.5e-07 $l=9.56556e-08 $layer=POLY_cond $X=12.935 $Y=1.575
+ $X2=12.982 $Y2=1.65
r241 29 31 471.745 $w=1.5e-07 $l=9.2e-07 $layer=POLY_cond $X=12.935 $Y=1.575
+ $X2=12.935 $Y2=0.655
r242 27 55 12.05 $w=1.5e-07 $l=1.22e-07 $layer=POLY_cond $X=12.86 $Y=1.65
+ $X2=12.982 $Y2=1.65
r243 27 28 176.904 $w=1.5e-07 $l=3.45e-07 $layer=POLY_cond $X=12.86 $Y=1.65
+ $X2=12.515 $Y2=1.65
r244 26 28 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=12.44 $Y=1.575
+ $X2=12.515 $Y2=1.65
r245 25 54 38.4574 $w=4.95e-07 $l=2.83026e-07 $layer=POLY_cond $X=12.44 $Y=0.935
+ $X2=12.365 $Y2=0.687
r246 25 26 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=12.44 $Y=0.935
+ $X2=12.44 $Y2=1.575
r247 24 53 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=11.235 $Y=0.86
+ $X2=11.4 $Y2=0.86
r248 21 24 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=11.16 $Y=0.935
+ $X2=11.235 $Y2=0.86
r249 21 50 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=11.16 $Y=0.935
+ $X2=11.16 $Y2=1.575
r250 20 51 692.234 $w=1.5e-07 $l=1.35e-06 $layer=POLY_cond $X=11.14 $Y=3.075
+ $X2=11.14 $Y2=1.725
r251 17 20 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=11.065 $Y=3.15
+ $X2=11.14 $Y2=3.075
r252 17 18 723 $w=1.5e-07 $l=1.41e-06 $layer=POLY_cond $X=11.065 $Y=3.15
+ $X2=9.655 $Y2=3.15
r253 16 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.58 $Y=3.075
+ $X2=9.655 $Y2=3.15
r254 15 48 30.233 $w=2.79e-07 $l=2.39583e-07 $layer=POLY_cond $X=9.58 $Y=1.715
+ $X2=9.405 $Y2=1.562
r255 15 16 697.362 $w=1.5e-07 $l=1.36e-06 $layer=POLY_cond $X=9.58 $Y=1.715
+ $X2=9.58 $Y2=3.075
r256 11 48 17.2686 $w=1.5e-07 $l=1.52e-07 $layer=POLY_cond $X=9.405 $Y=1.41
+ $X2=9.405 $Y2=1.562
r257 11 13 387.138 $w=1.5e-07 $l=7.55e-07 $layer=POLY_cond $X=9.405 $Y=1.41
+ $X2=9.405 $Y2=0.655
r258 8 47 17.2686 $w=1.5e-07 $l=1.53e-07 $layer=POLY_cond $X=9.09 $Y=1.715
+ $X2=9.09 $Y2=1.562
r259 8 10 241 $w=1.5e-07 $l=7.5e-07 $layer=POLY_cond $X=9.09 $Y=1.715 $X2=9.09
+ $Y2=2.465
r260 4 46 17.2686 $w=1.5e-07 $l=1.52e-07 $layer=POLY_cond $X=8.795 $Y=1.41
+ $X2=8.795 $Y2=1.562
r261 4 6 387.138 $w=1.5e-07 $l=7.55e-07 $layer=POLY_cond $X=8.795 $Y=1.41
+ $X2=8.795 $Y2=0.655
r262 1 45 17.2686 $w=1.5e-07 $l=1.53e-07 $layer=POLY_cond $X=8.66 $Y=1.715
+ $X2=8.66 $Y2=1.562
r263 1 3 241 $w=1.5e-07 $l=7.5e-07 $layer=POLY_cond $X=8.66 $Y=1.715 $X2=8.66
+ $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__BUSDRIVERNOVLPSLEEP_20%A_2063_47# 1 2 9 10 12 14 17
+ 21 22 24 26 27 30 31 33 37 39 41 42 43
c146 41 0 3.00155e-20 $X=11.055 $Y=1.042
c147 39 0 1.92998e-19 $X=11.055 $Y=1.93
c148 33 0 3.13694e-20 $X=13.91 $Y=1.44
c149 26 0 1.88719e-19 $X=11.055 $Y=1.845
c150 12 0 8.57257e-20 $X=14.385 $Y=1.185
r151 42 43 30.474 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=13.91 $Y=1.26
+ $X2=13.91 $Y2=1.185
r152 37 39 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=10.665 $Y=1.93
+ $X2=11.055 $Y2=1.93
r153 34 42 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=13.91 $Y=1.44
+ $X2=13.91 $Y2=1.26
r154 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=13.91
+ $Y=1.44 $X2=13.91 $Y2=1.44
r155 31 33 50.8123 $w=3.28e-07 $l=1.455e-06 $layer=LI1_cond $X=12.455 $Y=1.44
+ $X2=13.91 $Y2=1.44
r156 30 31 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=12.37 $Y=1.275
+ $X2=12.455 $Y2=1.44
r157 29 30 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=12.37 $Y=1.13
+ $X2=12.37 $Y2=1.275
r158 28 41 1.23839 $w=1.75e-07 $l=8.5e-08 $layer=LI1_cond $X=11.14 $Y=1.042
+ $X2=11.055 $Y2=1.042
r159 27 29 6.81835 $w=1.75e-07 $l=1.23386e-07 $layer=LI1_cond $X=12.285 $Y=1.042
+ $X2=12.37 $Y2=1.13
r160 27 28 72.5662 $w=1.73e-07 $l=1.145e-06 $layer=LI1_cond $X=12.285 $Y=1.042
+ $X2=11.14 $Y2=1.042
r161 26 39 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.055 $Y=1.845
+ $X2=11.055 $Y2=1.93
r162 25 41 5.29182 $w=1.7e-07 $l=8.8e-08 $layer=LI1_cond $X=11.055 $Y=1.13
+ $X2=11.055 $Y2=1.042
r163 25 26 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=11.055 $Y=1.13
+ $X2=11.055 $Y2=1.845
r164 24 41 5.29182 $w=1.7e-07 $l=8.7e-08 $layer=LI1_cond $X=11.055 $Y=0.955
+ $X2=11.055 $Y2=1.042
r165 23 24 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=11.055 $Y=0.815
+ $X2=11.055 $Y2=0.955
r166 21 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.97 $Y=0.73
+ $X2=11.055 $Y2=0.815
r167 21 22 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=10.97 $Y=0.73
+ $X2=10.55 $Y2=0.73
r168 15 22 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=10.455 $Y=0.645
+ $X2=10.55 $Y2=0.73
r169 15 17 10.2153 $w=1.88e-07 $l=1.75e-07 $layer=LI1_cond $X=10.455 $Y=0.645
+ $X2=10.455 $Y2=0.47
r170 12 14 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=14.385 $Y=1.185
+ $X2=14.385 $Y2=0.655
r171 11 42 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=14.075 $Y=1.26
+ $X2=13.91 $Y2=1.26
r172 10 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=14.31 $Y=1.26
+ $X2=14.385 $Y2=1.185
r173 10 11 120.5 $w=1.5e-07 $l=2.35e-07 $layer=POLY_cond $X=14.31 $Y=1.26
+ $X2=14.075 $Y2=1.26
r174 9 43 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=13.955 $Y=0.655
+ $X2=13.955 $Y2=1.185
r175 2 37 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=10.525
+ $Y=1.865 $X2=10.665 $Y2=2.01
r176 1 17 182 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=1 $X=10.315
+ $Y=0.235 $X2=10.455 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_LP__BUSDRIVERNOVLPSLEEP_20%VPWR 1 2 3 4 5 6 7 8 9 10 11
+ 12 13 14 15 16 17 18 57 63 67 71 75 79 81 85 89 95 99 103 107 109 113 117 121
+ 125 129 133 136 137 139 140 142 143 145 146 147 148 150 151 153 154 156 157
+ 159 160 161 163 168 180 187 192 197 231 237 238 241 244 247 250 253 256 259
+ 262 265
c417 238 0 2.64808e-19 $X=23.28 $Y=3.33
c418 75 0 1.91794e-19 $X=9.875 $Y=2.01
r419 265 266 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=22.8 $Y=3.33
+ $X2=22.8 $Y2=3.33
r420 262 263 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=18.48 $Y=3.33
+ $X2=18.48 $Y2=3.33
r421 259 260 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.16 $Y=3.33
+ $X2=14.16 $Y2=3.33
r422 256 257 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=12.24 $Y=3.33
+ $X2=12.24 $Y2=3.33
r423 253 254 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=11.28 $Y=3.33
+ $X2=11.28 $Y2=3.33
r424 250 251 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r425 247 248 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r426 244 245 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r427 241 242 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r428 238 266 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=23.28 $Y=3.33
+ $X2=22.8 $Y2=3.33
r429 237 238 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=23.28 $Y=3.33
+ $X2=23.28 $Y2=3.33
r430 235 265 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=22.96 $Y=3.33
+ $X2=22.835 $Y2=3.33
r431 235 237 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=22.96 $Y=3.33
+ $X2=23.28 $Y2=3.33
r432 234 266 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=22.32 $Y=3.33
+ $X2=22.8 $Y2=3.33
r433 233 234 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=22.32 $Y=3.33
+ $X2=22.32 $Y2=3.33
r434 231 265 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=22.71 $Y=3.33
+ $X2=22.835 $Y2=3.33
r435 231 233 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=22.71 $Y=3.33
+ $X2=22.32 $Y2=3.33
r436 230 234 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=21.84 $Y=3.33
+ $X2=22.32 $Y2=3.33
r437 229 230 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=21.84 $Y=3.33
+ $X2=21.84 $Y2=3.33
r438 227 230 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=20.88 $Y=3.33
+ $X2=21.84 $Y2=3.33
r439 226 227 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=20.88 $Y=3.33
+ $X2=20.88 $Y2=3.33
r440 224 227 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=19.92 $Y=3.33
+ $X2=20.88 $Y2=3.33
r441 223 224 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=19.92 $Y=3.33
+ $X2=19.92 $Y2=3.33
r442 221 224 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=18.96 $Y=3.33
+ $X2=19.92 $Y2=3.33
r443 221 263 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=18.96 $Y=3.33
+ $X2=18.48 $Y2=3.33
r444 220 221 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=18.96 $Y=3.33
+ $X2=18.96 $Y2=3.33
r445 218 262 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=18.58 $Y=3.33
+ $X2=18.495 $Y2=3.33
r446 218 220 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=18.58 $Y=3.33
+ $X2=18.96 $Y2=3.33
r447 217 263 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=17.52 $Y=3.33
+ $X2=18.48 $Y2=3.33
r448 216 217 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=17.52 $Y=3.33
+ $X2=17.52 $Y2=3.33
r449 214 217 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=16.56 $Y=3.33
+ $X2=17.52 $Y2=3.33
r450 213 214 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=16.56 $Y=3.33
+ $X2=16.56 $Y2=3.33
r451 211 214 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=15.6 $Y=3.33
+ $X2=16.56 $Y2=3.33
r452 210 211 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=15.6 $Y=3.33
+ $X2=15.6 $Y2=3.33
r453 208 211 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=14.64 $Y=3.33
+ $X2=15.6 $Y2=3.33
r454 208 260 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=14.64 $Y=3.33
+ $X2=14.16 $Y2=3.33
r455 207 208 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.64 $Y=3.33
+ $X2=14.64 $Y2=3.33
r456 205 259 8.70163 $w=1.7e-07 $l=1.68e-07 $layer=LI1_cond $X=14.36 $Y=3.33
+ $X2=14.192 $Y2=3.33
r457 205 207 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=14.36 $Y=3.33
+ $X2=14.64 $Y2=3.33
r458 204 260 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.68 $Y=3.33
+ $X2=14.16 $Y2=3.33
r459 203 204 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=13.68 $Y=3.33
+ $X2=13.68 $Y2=3.33
r460 201 204 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=12.72 $Y=3.33
+ $X2=13.68 $Y2=3.33
r461 201 257 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.72 $Y=3.33
+ $X2=12.24 $Y2=3.33
r462 200 203 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=12.72 $Y=3.33
+ $X2=13.68 $Y2=3.33
r463 200 201 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=12.72 $Y=3.33
+ $X2=12.72 $Y2=3.33
r464 198 256 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=12.46 $Y=3.33
+ $X2=12.33 $Y2=3.33
r465 198 200 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=12.46 $Y=3.33
+ $X2=12.72 $Y2=3.33
r466 197 259 8.70163 $w=1.7e-07 $l=1.67e-07 $layer=LI1_cond $X=14.025 $Y=3.33
+ $X2=14.192 $Y2=3.33
r467 197 203 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=14.025 $Y=3.33
+ $X2=13.68 $Y2=3.33
r468 196 254 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=10.32 $Y=3.33
+ $X2=11.28 $Y2=3.33
r469 196 251 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=3.33
+ $X2=9.84 $Y2=3.33
r470 195 196 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=10.32 $Y=3.33
+ $X2=10.32 $Y2=3.33
r471 193 250 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.04 $Y=3.33
+ $X2=9.875 $Y2=3.33
r472 193 195 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=10.04 $Y=3.33
+ $X2=10.32 $Y2=3.33
r473 192 253 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=11.27 $Y=3.33
+ $X2=11.4 $Y2=3.33
r474 192 195 61.9786 $w=1.68e-07 $l=9.5e-07 $layer=LI1_cond $X=11.27 $Y=3.33
+ $X2=10.32 $Y2=3.33
r475 191 251 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=9.84 $Y2=3.33
r476 191 248 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=8.88 $Y2=3.33
r477 190 191 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r478 188 247 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=9.04 $Y=3.33
+ $X2=8.91 $Y2=3.33
r479 188 190 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=9.04 $Y=3.33
+ $X2=9.36 $Y2=3.33
r480 187 250 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.71 $Y=3.33
+ $X2=9.875 $Y2=3.33
r481 187 190 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=9.71 $Y=3.33
+ $X2=9.36 $Y2=3.33
r482 186 248 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=8.88 $Y2=3.33
r483 185 186 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r484 183 186 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=6.96 $Y=3.33
+ $X2=8.4 $Y2=3.33
r485 182 185 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=6.96 $Y=3.33
+ $X2=8.4 $Y2=3.33
r486 182 183 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.96 $Y=3.33
+ $X2=6.96 $Y2=3.33
r487 180 247 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=8.78 $Y=3.33
+ $X2=8.91 $Y2=3.33
r488 180 185 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=8.78 $Y=3.33
+ $X2=8.4 $Y2=3.33
r489 179 183 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=6.96 $Y2=3.33
r490 179 245 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=5.52 $Y2=3.33
r491 178 179 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r492 176 244 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.735 $Y=3.33
+ $X2=5.57 $Y2=3.33
r493 176 178 48.6043 $w=1.68e-07 $l=7.45e-07 $layer=LI1_cond $X=5.735 $Y=3.33
+ $X2=6.48 $Y2=3.33
r494 175 245 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=5.52 $Y2=3.33
r495 174 175 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r496 172 175 1.07034 $w=4.9e-07 $l=3.84e-06 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=5.04 $Y2=3.33
r497 172 242 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r498 171 174 250.524 $w=1.68e-07 $l=3.84e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=5.04 $Y2=3.33
r499 171 172 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r500 169 241 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.955 $Y=3.33
+ $X2=0.79 $Y2=3.33
r501 169 171 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=0.955 $Y=3.33
+ $X2=1.2 $Y2=3.33
r502 168 244 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.405 $Y=3.33
+ $X2=5.57 $Y2=3.33
r503 168 174 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=5.405 $Y=3.33
+ $X2=5.04 $Y2=3.33
r504 166 242 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r505 165 166 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r506 163 241 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.625 $Y=3.33
+ $X2=0.79 $Y2=3.33
r507 163 165 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=0.625 $Y=3.33
+ $X2=0.24 $Y2=3.33
r508 161 257 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.76 $Y=3.33
+ $X2=12.24 $Y2=3.33
r509 161 254 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.76 $Y=3.33
+ $X2=11.28 $Y2=3.33
r510 159 229 0.652406 $w=1.68e-07 $l=1e-08 $layer=LI1_cond $X=21.85 $Y=3.33
+ $X2=21.84 $Y2=3.33
r511 159 160 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=21.85 $Y=3.33
+ $X2=21.935 $Y2=3.33
r512 158 233 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=22.02 $Y=3.33
+ $X2=22.32 $Y2=3.33
r513 158 160 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=22.02 $Y=3.33
+ $X2=21.935 $Y2=3.33
r514 156 226 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=20.99 $Y=3.33
+ $X2=20.88 $Y2=3.33
r515 156 157 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=20.99 $Y=3.33
+ $X2=21.075 $Y2=3.33
r516 155 229 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=21.16 $Y=3.33
+ $X2=21.84 $Y2=3.33
r517 155 157 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=21.16 $Y=3.33
+ $X2=21.075 $Y2=3.33
r518 153 223 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=20.13 $Y=3.33
+ $X2=19.92 $Y2=3.33
r519 153 154 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=20.13 $Y=3.33
+ $X2=20.215 $Y2=3.33
r520 152 226 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=20.3 $Y=3.33
+ $X2=20.88 $Y2=3.33
r521 152 154 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=20.3 $Y=3.33
+ $X2=20.215 $Y2=3.33
r522 150 220 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=19.27 $Y=3.33
+ $X2=18.96 $Y2=3.33
r523 150 151 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=19.27 $Y=3.33
+ $X2=19.355 $Y2=3.33
r524 149 223 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=19.44 $Y=3.33
+ $X2=19.92 $Y2=3.33
r525 149 151 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=19.44 $Y=3.33
+ $X2=19.355 $Y2=3.33
r526 147 216 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=17.55 $Y=3.33
+ $X2=17.52 $Y2=3.33
r527 147 148 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=17.55 $Y=3.33
+ $X2=17.635 $Y2=3.33
r528 145 213 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=16.69 $Y=3.33
+ $X2=16.56 $Y2=3.33
r529 145 146 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=16.69 $Y=3.33
+ $X2=16.775 $Y2=3.33
r530 144 216 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=16.86 $Y=3.33
+ $X2=17.52 $Y2=3.33
r531 144 146 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=16.86 $Y=3.33
+ $X2=16.775 $Y2=3.33
r532 142 210 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=15.83 $Y=3.33
+ $X2=15.6 $Y2=3.33
r533 142 143 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=15.83 $Y=3.33
+ $X2=15.915 $Y2=3.33
r534 141 213 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=16 $Y=3.33
+ $X2=16.56 $Y2=3.33
r535 141 143 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=16 $Y=3.33
+ $X2=15.915 $Y2=3.33
r536 139 207 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=14.89 $Y=3.33
+ $X2=14.64 $Y2=3.33
r537 139 140 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=14.89 $Y=3.33
+ $X2=15.015 $Y2=3.33
r538 138 210 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=15.14 $Y=3.33
+ $X2=15.6 $Y2=3.33
r539 138 140 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=15.14 $Y=3.33
+ $X2=15.015 $Y2=3.33
r540 136 178 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=6.705 $Y=3.33
+ $X2=6.48 $Y2=3.33
r541 136 137 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.705 $Y=3.33
+ $X2=6.83 $Y2=3.33
r542 135 182 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=6.955 $Y=3.33
+ $X2=6.96 $Y2=3.33
r543 135 137 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.955 $Y=3.33
+ $X2=6.83 $Y2=3.33
r544 131 265 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=22.835 $Y=3.245
+ $X2=22.835 $Y2=3.33
r545 131 133 36.4172 $w=2.48e-07 $l=7.9e-07 $layer=LI1_cond $X=22.835 $Y=3.245
+ $X2=22.835 $Y2=2.455
r546 127 160 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=21.935 $Y=3.245
+ $X2=21.935 $Y2=3.33
r547 127 129 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=21.935 $Y=3.245
+ $X2=21.935 $Y2=2.455
r548 123 157 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=21.075 $Y=3.245
+ $X2=21.075 $Y2=3.33
r549 123 125 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=21.075 $Y=3.245
+ $X2=21.075 $Y2=2.455
r550 119 154 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=20.215 $Y=3.245
+ $X2=20.215 $Y2=3.33
r551 119 121 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=20.215 $Y=3.245
+ $X2=20.215 $Y2=2.455
r552 115 151 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=19.355 $Y=3.245
+ $X2=19.355 $Y2=3.33
r553 115 117 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=19.355 $Y=3.245
+ $X2=19.355 $Y2=2.455
r554 111 262 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=18.495 $Y=3.245
+ $X2=18.495 $Y2=3.33
r555 111 113 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=18.495 $Y=3.245
+ $X2=18.495 $Y2=2.455
r556 110 148 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=17.72 $Y=3.33
+ $X2=17.635 $Y2=3.33
r557 109 262 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=18.41 $Y=3.33
+ $X2=18.495 $Y2=3.33
r558 109 110 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=18.41 $Y=3.33
+ $X2=17.72 $Y2=3.33
r559 105 148 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=17.635 $Y=3.245
+ $X2=17.635 $Y2=3.33
r560 105 107 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=17.635 $Y=3.245
+ $X2=17.635 $Y2=2.455
r561 101 146 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=16.775 $Y=3.245
+ $X2=16.775 $Y2=3.33
r562 101 103 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=16.775 $Y=3.245
+ $X2=16.775 $Y2=2.455
r563 97 143 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=15.915 $Y=3.245
+ $X2=15.915 $Y2=3.33
r564 97 99 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=15.915 $Y=3.245
+ $X2=15.915 $Y2=2.455
r565 93 140 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=15.015 $Y=3.245
+ $X2=15.015 $Y2=3.33
r566 93 95 35.4952 $w=2.48e-07 $l=7.7e-07 $layer=LI1_cond $X=15.015 $Y=3.245
+ $X2=15.015 $Y2=2.475
r567 89 92 23.3929 $w=3.33e-07 $l=6.8e-07 $layer=LI1_cond $X=14.192 $Y=2.27
+ $X2=14.192 $Y2=2.95
r568 87 259 0.942324 $w=3.35e-07 $l=8.5e-08 $layer=LI1_cond $X=14.192 $Y=3.245
+ $X2=14.192 $Y2=3.33
r569 87 92 10.1484 $w=3.33e-07 $l=2.95e-07 $layer=LI1_cond $X=14.192 $Y=3.245
+ $X2=14.192 $Y2=2.95
r570 83 256 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=12.33 $Y=3.245
+ $X2=12.33 $Y2=3.33
r571 83 85 15.292 $w=2.58e-07 $l=3.45e-07 $layer=LI1_cond $X=12.33 $Y=3.245
+ $X2=12.33 $Y2=2.9
r572 82 253 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=11.53 $Y=3.33
+ $X2=11.4 $Y2=3.33
r573 81 256 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=12.2 $Y=3.33
+ $X2=12.33 $Y2=3.33
r574 81 82 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=12.2 $Y=3.33
+ $X2=11.53 $Y2=3.33
r575 77 253 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=11.4 $Y=3.245
+ $X2=11.4 $Y2=3.33
r576 77 79 33.6868 $w=2.58e-07 $l=7.6e-07 $layer=LI1_cond $X=11.4 $Y=3.245
+ $X2=11.4 $Y2=2.485
r577 73 250 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.875 $Y=3.245
+ $X2=9.875 $Y2=3.33
r578 73 75 43.1293 $w=3.28e-07 $l=1.235e-06 $layer=LI1_cond $X=9.875 $Y=3.245
+ $X2=9.875 $Y2=2.01
r579 69 247 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=8.91 $Y=3.245
+ $X2=8.91 $Y2=3.33
r580 69 71 18.1731 $w=2.58e-07 $l=4.1e-07 $layer=LI1_cond $X=8.91 $Y=3.245
+ $X2=8.91 $Y2=2.835
r581 65 137 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.83 $Y=3.245
+ $X2=6.83 $Y2=3.33
r582 65 67 29.733 $w=2.48e-07 $l=6.45e-07 $layer=LI1_cond $X=6.83 $Y=3.245
+ $X2=6.83 $Y2=2.6
r583 61 244 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.57 $Y=3.245
+ $X2=5.57 $Y2=3.33
r584 61 63 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=5.57 $Y=3.245
+ $X2=5.57 $Y2=2.83
r585 57 60 16.4136 $w=3.28e-07 $l=4.7e-07 $layer=LI1_cond $X=0.79 $Y=2.43
+ $X2=0.79 $Y2=2.9
r586 55 241 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.79 $Y=3.245
+ $X2=0.79 $Y2=3.33
r587 55 60 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=0.79 $Y=3.245
+ $X2=0.79 $Y2=2.9
r588 18 133 300 $w=1.7e-07 $l=6.8644e-07 $layer=licon1_PDIFF $count=2 $X=22.655
+ $Y=1.835 $X2=22.795 $Y2=2.455
r589 17 129 300 $w=1.7e-07 $l=6.8644e-07 $layer=licon1_PDIFF $count=2 $X=21.795
+ $Y=1.835 $X2=21.935 $Y2=2.455
r590 16 125 300 $w=1.7e-07 $l=6.8644e-07 $layer=licon1_PDIFF $count=2 $X=20.935
+ $Y=1.835 $X2=21.075 $Y2=2.455
r591 15 121 300 $w=1.7e-07 $l=6.8644e-07 $layer=licon1_PDIFF $count=2 $X=20.075
+ $Y=1.835 $X2=20.215 $Y2=2.455
r592 14 117 300 $w=1.7e-07 $l=6.8644e-07 $layer=licon1_PDIFF $count=2 $X=19.215
+ $Y=1.835 $X2=19.355 $Y2=2.455
r593 13 113 300 $w=1.7e-07 $l=6.8644e-07 $layer=licon1_PDIFF $count=2 $X=18.355
+ $Y=1.835 $X2=18.495 $Y2=2.455
r594 12 107 300 $w=1.7e-07 $l=6.8644e-07 $layer=licon1_PDIFF $count=2 $X=17.495
+ $Y=1.835 $X2=17.635 $Y2=2.455
r595 11 103 300 $w=1.7e-07 $l=6.8644e-07 $layer=licon1_PDIFF $count=2 $X=16.635
+ $Y=1.835 $X2=16.775 $Y2=2.455
r596 10 99 300 $w=1.7e-07 $l=6.8644e-07 $layer=licon1_PDIFF $count=2 $X=15.775
+ $Y=1.835 $X2=15.915 $Y2=2.455
r597 9 95 300 $w=1.7e-07 $l=7.06541e-07 $layer=licon1_PDIFF $count=2 $X=14.915
+ $Y=1.835 $X2=15.055 $Y2=2.475
r598 8 92 400 $w=1.7e-07 $l=1.17584e-06 $layer=licon1_PDIFF $count=1 $X=14.07
+ $Y=1.835 $X2=14.195 $Y2=2.95
r599 8 89 400 $w=1.7e-07 $l=4.93559e-07 $layer=licon1_PDIFF $count=1 $X=14.07
+ $Y=1.835 $X2=14.195 $Y2=2.27
r600 7 85 600 $w=1.7e-07 $l=1.13284e-06 $layer=licon1_PDIFF $count=1 $X=12.155
+ $Y=1.835 $X2=12.295 $Y2=2.9
r601 6 79 300 $w=1.7e-07 $l=7.09753e-07 $layer=licon1_PDIFF $count=2 $X=11.31
+ $Y=1.835 $X2=11.435 $Y2=2.485
r602 5 75 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=9.73
+ $Y=1.865 $X2=9.875 $Y2=2.01
r603 4 71 600 $w=1.7e-07 $l=1.06771e-06 $layer=licon1_PDIFF $count=1 $X=8.735
+ $Y=1.835 $X2=8.875 $Y2=2.835
r604 3 67 300 $w=1.7e-07 $l=4.09054e-07 $layer=licon1_PDIFF $count=2 $X=6.65
+ $Y=2.255 $X2=6.79 $Y2=2.6
r605 2 63 600 $w=1.7e-07 $l=6.34429e-07 $layer=licon1_PDIFF $count=1 $X=5.445
+ $Y=2.255 $X2=5.57 $Y2=2.83
r606 1 60 600 $w=1.7e-07 $l=8.72195e-07 $layer=licon1_PDIFF $count=1 $X=0.65
+ $Y=2.095 $X2=0.79 $Y2=2.9
r607 1 57 600 $w=1.7e-07 $l=3.98905e-07 $layer=licon1_PDIFF $count=1 $X=0.65
+ $Y=2.095 $X2=0.79 $Y2=2.43
.ends

.subckt PM_SKY130_FD_SC_LP__BUSDRIVERNOVLPSLEEP_20%KAPWR 1 2 3 10 21 25 33
r188 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=2.8
+ $X2=5.04 $Y2=2.8
r189 29 34 0.464569 $w=2.7e-07 $l=8.5e-07 $layer=MET1_cond $X=4.19 $Y=2.81
+ $X2=5.04 $Y2=2.81
r190 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.19 $Y=2.8
+ $X2=4.19 $Y2=2.8
r191 25 28 36.1867 $w=2.48e-07 $l=7.85e-07 $layer=LI1_cond $X=4.19 $Y=2.015
+ $X2=4.19 $Y2=2.8
r192 22 29 0.483698 $w=2.7e-07 $l=8.85e-07 $layer=MET1_cond $X=3.305 $Y=2.81
+ $X2=4.19 $Y2=2.81
r193 21 22 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.305 $Y=2.8
+ $X2=3.305 $Y2=2.8
r194 19 21 1.31851 $w=6.33e-07 $l=7e-08 $layer=LI1_cond $X=3.235 $Y=2.757
+ $X2=3.305 $Y2=2.757
r195 17 19 10.8306 $w=6.33e-07 $l=5.75e-07 $layer=LI1_cond $X=2.66 $Y=2.757
+ $X2=3.235 $Y2=2.757
r196 14 22 0.393517 $w=2.7e-07 $l=7.2e-07 $layer=MET1_cond $X=2.585 $Y=2.81
+ $X2=3.305 $Y2=2.81
r197 13 17 1.41269 $w=6.33e-07 $l=7.5e-08 $layer=LI1_cond $X=2.585 $Y=2.757
+ $X2=2.66 $Y2=2.757
r198 13 14 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.585 $Y=2.8
+ $X2=2.585 $Y2=2.8
r199 10 34 3.67283 $w=2.7e-07 $l=6.72e-06 $layer=MET1_cond $X=11.76 $Y=2.81
+ $X2=5.04 $Y2=2.81
r200 3 33 600 $w=1.7e-07 $l=1.02762e-06 $layer=licon1_PDIFF $count=1 $X=4.91
+ $Y=1.835 $X2=5.05 $Y2=2.795
r201 2 28 400 $w=1.7e-07 $l=1.1128e-06 $layer=licon1_PDIFF $count=1 $X=4.05
+ $Y=1.835 $X2=4.19 $Y2=2.88
r202 2 25 400 $w=1.7e-07 $l=2.4e-07 $layer=licon1_PDIFF $count=1 $X=4.05
+ $Y=1.835 $X2=4.19 $Y2=2.015
r203 1 19 300 $w=1.7e-07 $l=8.45192e-07 $layer=licon1_PDIFF $count=2 $X=2.45
+ $Y=2.455 $X2=3.235 $Y2=2.58
r204 1 17 300 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=2 $X=2.45
+ $Y=2.455 $X2=2.66 $Y2=2.58
.ends

.subckt PM_SKY130_FD_SC_LP__BUSDRIVERNOVLPSLEEP_20%A_1492_367# 1 2 3 10 12 14 18
+ 21 22 28 32
c67 12 0 2.32147e-19 $X=7.585 $Y=1.98
r68 23 28 3.59259 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=8.61 $Y=2.41
+ $X2=8.445 $Y2=2.41
r69 22 32 4.20357 $w=1.8e-07 $l=1.3e-07 $layer=LI1_cond $X=9.21 $Y=2.41 $X2=9.34
+ $Y2=2.41
r70 22 23 36.9697 $w=1.78e-07 $l=6e-07 $layer=LI1_cond $X=9.21 $Y=2.41 $X2=8.61
+ $Y2=2.41
r71 21 30 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.445 $Y=2.895
+ $X2=8.445 $Y2=2.98
r72 20 28 3.0419 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=8.445 $Y=2.5 $X2=8.445
+ $Y2=2.41
r73 20 21 13.7944 $w=3.28e-07 $l=3.95e-07 $layer=LI1_cond $X=8.445 $Y=2.5
+ $X2=8.445 $Y2=2.895
r74 16 28 3.0419 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=8.445 $Y=2.32 $X2=8.445
+ $Y2=2.41
r75 16 18 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=8.445 $Y=2.32
+ $X2=8.445 $Y2=1.98
r76 15 27 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.75 $Y=2.98
+ $X2=7.625 $Y2=2.98
r77 14 30 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.28 $Y=2.98
+ $X2=8.445 $Y2=2.98
r78 14 15 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=8.28 $Y=2.98
+ $X2=7.75 $Y2=2.98
r79 10 27 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.625 $Y=2.895
+ $X2=7.625 $Y2=2.98
r80 10 12 42.1794 $w=2.48e-07 $l=9.15e-07 $layer=LI1_cond $X=7.625 $Y=2.895
+ $X2=7.625 $Y2=1.98
r81 3 32 300 $w=1.7e-07 $l=7.16589e-07 $layer=licon1_PDIFF $count=2 $X=9.165
+ $Y=1.835 $X2=9.305 $Y2=2.485
r82 2 30 400 $w=1.7e-07 $l=1.13284e-06 $layer=licon1_PDIFF $count=1 $X=8.305
+ $Y=1.835 $X2=8.445 $Y2=2.9
r83 2 18 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=8.305
+ $Y=1.835 $X2=8.445 $Y2=1.98
r84 1 27 400 $w=1.7e-07 $l=1.12577e-06 $layer=licon1_PDIFF $count=1 $X=7.46
+ $Y=1.835 $X2=7.585 $Y2=2.9
r85 1 12 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=7.46
+ $Y=1.835 $X2=7.585 $Y2=1.98
.ends

.subckt PM_SKY130_FD_SC_LP__BUSDRIVERNOVLPSLEEP_20%A_2345_367# 1 2 3 12 14 15 16
+ 17 18 20 23
c61 23 0 1.29574e-19 $X=11.865 $Y=2.485
c62 14 0 1.12422e-19 $X=12.815 $Y=2.49
r63 18 27 3.75819 $w=2.5e-07 $l=1.5e-07 $layer=LI1_cond $X=13.715 $Y=2.775
+ $X2=13.715 $Y2=2.925
r64 18 20 19.5915 $w=2.48e-07 $l=4.25e-07 $layer=LI1_cond $X=13.715 $Y=2.775
+ $X2=13.715 $Y2=2.35
r65 16 27 3.13183 $w=3e-07 $l=1.25e-07 $layer=LI1_cond $X=13.59 $Y=2.925
+ $X2=13.715 $Y2=2.925
r66 16 17 23.433 $w=2.98e-07 $l=6.1e-07 $layer=LI1_cond $X=13.59 $Y=2.925
+ $X2=12.98 $Y2=2.925
r67 15 17 6.83662 $w=3e-07 $l=2.2798e-07 $layer=LI1_cond $X=12.815 $Y=2.775
+ $X2=12.98 $Y2=2.925
r68 14 25 3.0783 $w=3.3e-07 $l=1.53e-07 $layer=LI1_cond $X=12.815 $Y=2.49
+ $X2=12.815 $Y2=2.337
r69 14 15 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=12.815 $Y=2.49
+ $X2=12.815 $Y2=2.775
r70 13 23 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.03 $Y=2.405
+ $X2=11.865 $Y2=2.405
r71 12 25 4.68787 $w=1.7e-07 $l=1.96074e-07 $layer=LI1_cond $X=12.65 $Y=2.405
+ $X2=12.815 $Y2=2.337
r72 12 13 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=12.65 $Y=2.405
+ $X2=12.03 $Y2=2.405
r73 3 27 600 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=13.535
+ $Y=1.835 $X2=13.675 $Y2=2.91
r74 3 20 600 $w=1.7e-07 $l=5.80797e-07 $layer=licon1_PDIFF $count=1 $X=13.535
+ $Y=1.835 $X2=13.675 $Y2=2.35
r75 2 25 300 $w=1.7e-07 $l=5.74108e-07 $layer=licon1_PDIFF $count=2 $X=12.69
+ $Y=1.835 $X2=12.815 $Y2=2.35
r76 1 23 300 $w=1.7e-07 $l=7.16589e-07 $layer=licon1_PDIFF $count=2 $X=11.725
+ $Y=1.835 $X2=11.865 $Y2=2.485
.ends

.subckt PM_SKY130_FD_SC_LP__BUSDRIVERNOVLPSLEEP_20%Z 1 2 3 4 5 6 7 8 9 10 11 12
+ 13 14 15 16 17 18 55 57 59 63 67 69 72 82 92 102 112 122 132 142 143 154 168
r296 154 155 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=15.485 $Y=2.035
+ $X2=15.485 $Y2=2.035
r297 151 155 0.55178 $w=2.3e-07 $l=8.6e-07 $layer=MET1_cond $X=14.625 $Y=2.035
+ $X2=15.485 $Y2=2.035
r298 150 151 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.625 $Y=2.035
+ $X2=14.625 $Y2=2.035
r299 142 147 30.208 $w=3.28e-07 $l=8.65e-07 $layer=LI1_cond $X=22.365 $Y=2.035
+ $X2=22.365 $Y2=2.9
r300 142 143 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=22.365 $Y=2.035
+ $X2=22.365 $Y2=2.035
r301 136 143 0.55178 $w=2.3e-07 $l=8.6e-07 $layer=MET1_cond $X=21.505 $Y=2.035
+ $X2=22.365 $Y2=2.035
r302 136 168 0.413835 $w=2.3e-07 $l=6.45e-07 $layer=MET1_cond $X=21.505 $Y=2.035
+ $X2=20.86 $Y2=2.035
r303 135 139 30.208 $w=3.28e-07 $l=8.65e-07 $layer=LI1_cond $X=21.505 $Y=2.035
+ $X2=21.505 $Y2=2.9
r304 135 136 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=21.505 $Y=2.035
+ $X2=21.505 $Y2=2.035
r305 132 135 58.4952 $w=3.28e-07 $l=1.675e-06 $layer=LI1_cond $X=21.505 $Y=0.36
+ $X2=21.505 $Y2=2.035
r306 126 168 0.137945 $w=2.3e-07 $l=2.15e-07 $layer=MET1_cond $X=20.645 $Y=2.035
+ $X2=20.86 $Y2=2.035
r307 125 129 30.208 $w=3.28e-07 $l=8.65e-07 $layer=LI1_cond $X=20.645 $Y=2.035
+ $X2=20.645 $Y2=2.9
r308 125 126 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=20.645 $Y=2.035
+ $X2=20.645 $Y2=2.035
r309 122 125 58.4952 $w=3.28e-07 $l=1.675e-06 $layer=LI1_cond $X=20.645 $Y=0.36
+ $X2=20.645 $Y2=2.035
r310 116 126 0.55178 $w=2.3e-07 $l=8.6e-07 $layer=MET1_cond $X=19.785 $Y=2.035
+ $X2=20.645 $Y2=2.035
r311 115 119 30.208 $w=3.28e-07 $l=8.65e-07 $layer=LI1_cond $X=19.785 $Y=2.035
+ $X2=19.785 $Y2=2.9
r312 115 116 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=19.785 $Y=2.035
+ $X2=19.785 $Y2=2.035
r313 112 115 58.4952 $w=3.28e-07 $l=1.675e-06 $layer=LI1_cond $X=19.785 $Y=0.36
+ $X2=19.785 $Y2=2.035
r314 106 116 0.55178 $w=2.3e-07 $l=8.6e-07 $layer=MET1_cond $X=18.925 $Y=2.035
+ $X2=19.785 $Y2=2.035
r315 105 109 30.208 $w=3.28e-07 $l=8.65e-07 $layer=LI1_cond $X=18.925 $Y=2.035
+ $X2=18.925 $Y2=2.9
r316 105 106 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=18.925 $Y=2.035
+ $X2=18.925 $Y2=2.035
r317 102 105 58.4952 $w=3.28e-07 $l=1.675e-06 $layer=LI1_cond $X=18.925 $Y=0.36
+ $X2=18.925 $Y2=2.035
r318 95 99 30.208 $w=3.28e-07 $l=8.65e-07 $layer=LI1_cond $X=18.065 $Y=2.035
+ $X2=18.065 $Y2=2.9
r319 95 96 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=18.065 $Y=2.035
+ $X2=18.065 $Y2=2.035
r320 92 95 58.4952 $w=3.28e-07 $l=1.675e-06 $layer=LI1_cond $X=18.065 $Y=0.36
+ $X2=18.065 $Y2=2.035
r321 86 96 0.55178 $w=2.3e-07 $l=8.6e-07 $layer=MET1_cond $X=17.205 $Y=2.035
+ $X2=18.065 $Y2=2.035
r322 85 89 30.208 $w=3.28e-07 $l=8.65e-07 $layer=LI1_cond $X=17.205 $Y=2.035
+ $X2=17.205 $Y2=2.9
r323 85 86 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=17.205 $Y=2.035
+ $X2=17.205 $Y2=2.035
r324 82 85 58.4952 $w=3.28e-07 $l=1.675e-06 $layer=LI1_cond $X=17.205 $Y=0.36
+ $X2=17.205 $Y2=2.035
r325 76 86 0.55178 $w=2.3e-07 $l=8.6e-07 $layer=MET1_cond $X=16.345 $Y=2.035
+ $X2=17.205 $Y2=2.035
r326 76 155 0.55178 $w=2.3e-07 $l=8.6e-07 $layer=MET1_cond $X=16.345 $Y=2.035
+ $X2=15.485 $Y2=2.035
r327 75 79 30.208 $w=3.28e-07 $l=8.65e-07 $layer=LI1_cond $X=16.345 $Y=2.035
+ $X2=16.345 $Y2=2.9
r328 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=16.345 $Y=2.035
+ $X2=16.345 $Y2=2.035
r329 72 75 58.4952 $w=3.28e-07 $l=1.675e-06 $layer=LI1_cond $X=16.345 $Y=0.36
+ $X2=16.345 $Y2=2.035
r330 69 106 0.27589 $w=2.3e-07 $l=4.3e-07 $layer=MET1_cond $X=18.495 $Y=2.035
+ $X2=18.925 $Y2=2.035
r331 69 96 0.27589 $w=2.3e-07 $l=4.3e-07 $layer=MET1_cond $X=18.495 $Y=2.035
+ $X2=18.065 $Y2=2.035
r332 65 154 3.0419 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=15.485 $Y=2.13
+ $X2=15.485 $Y2=2.04
r333 65 67 26.8903 $w=3.28e-07 $l=7.7e-07 $layer=LI1_cond $X=15.485 $Y=2.13
+ $X2=15.485 $Y2=2.9
r334 61 154 3.0419 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=15.485 $Y=1.95
+ $X2=15.485 $Y2=2.04
r335 61 63 55.5268 $w=3.28e-07 $l=1.59e-06 $layer=LI1_cond $X=15.485 $Y=1.95
+ $X2=15.485 $Y2=0.36
r336 60 150 3.31438 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=14.71 $Y=2.04
+ $X2=14.625 $Y2=2.04
r337 59 154 3.59259 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=15.32 $Y=2.04
+ $X2=15.485 $Y2=2.04
r338 59 60 37.5859 $w=1.78e-07 $l=6.1e-07 $layer=LI1_cond $X=15.32 $Y=2.04
+ $X2=14.71 $Y2=2.04
r339 55 150 3.50935 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=14.625 $Y=2.13
+ $X2=14.625 $Y2=2.04
r340 55 57 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=14.625 $Y=2.13
+ $X2=14.625 $Y2=2.9
r341 18 147 400 $w=1.7e-07 $l=1.13284e-06 $layer=licon1_PDIFF $count=1 $X=22.225
+ $Y=1.835 $X2=22.365 $Y2=2.9
r342 18 142 400 $w=1.7e-07 $l=3.32716e-07 $layer=licon1_PDIFF $count=1 $X=22.225
+ $Y=1.835 $X2=22.365 $Y2=2.105
r343 17 139 400 $w=1.7e-07 $l=1.13284e-06 $layer=licon1_PDIFF $count=1 $X=21.365
+ $Y=1.835 $X2=21.505 $Y2=2.9
r344 17 135 400 $w=1.7e-07 $l=3.32716e-07 $layer=licon1_PDIFF $count=1 $X=21.365
+ $Y=1.835 $X2=21.505 $Y2=2.105
r345 16 129 400 $w=1.7e-07 $l=1.13284e-06 $layer=licon1_PDIFF $count=1 $X=20.505
+ $Y=1.835 $X2=20.645 $Y2=2.9
r346 16 125 400 $w=1.7e-07 $l=3.32716e-07 $layer=licon1_PDIFF $count=1 $X=20.505
+ $Y=1.835 $X2=20.645 $Y2=2.105
r347 15 119 400 $w=1.7e-07 $l=1.13284e-06 $layer=licon1_PDIFF $count=1 $X=19.645
+ $Y=1.835 $X2=19.785 $Y2=2.9
r348 15 115 400 $w=1.7e-07 $l=3.32716e-07 $layer=licon1_PDIFF $count=1 $X=19.645
+ $Y=1.835 $X2=19.785 $Y2=2.105
r349 14 109 400 $w=1.7e-07 $l=1.13284e-06 $layer=licon1_PDIFF $count=1 $X=18.785
+ $Y=1.835 $X2=18.925 $Y2=2.9
r350 14 105 400 $w=1.7e-07 $l=3.32716e-07 $layer=licon1_PDIFF $count=1 $X=18.785
+ $Y=1.835 $X2=18.925 $Y2=2.105
r351 13 99 400 $w=1.7e-07 $l=1.13284e-06 $layer=licon1_PDIFF $count=1 $X=17.925
+ $Y=1.835 $X2=18.065 $Y2=2.9
r352 13 95 400 $w=1.7e-07 $l=3.32716e-07 $layer=licon1_PDIFF $count=1 $X=17.925
+ $Y=1.835 $X2=18.065 $Y2=2.105
r353 12 89 400 $w=1.7e-07 $l=1.13284e-06 $layer=licon1_PDIFF $count=1 $X=17.065
+ $Y=1.835 $X2=17.205 $Y2=2.9
r354 12 85 400 $w=1.7e-07 $l=3.32716e-07 $layer=licon1_PDIFF $count=1 $X=17.065
+ $Y=1.835 $X2=17.205 $Y2=2.105
r355 11 79 400 $w=1.7e-07 $l=1.13284e-06 $layer=licon1_PDIFF $count=1 $X=16.205
+ $Y=1.835 $X2=16.345 $Y2=2.9
r356 11 75 400 $w=1.7e-07 $l=3.32716e-07 $layer=licon1_PDIFF $count=1 $X=16.205
+ $Y=1.835 $X2=16.345 $Y2=2.105
r357 10 154 400 $w=1.7e-07 $l=3.32716e-07 $layer=licon1_PDIFF $count=1 $X=15.345
+ $Y=1.835 $X2=15.485 $Y2=2.105
r358 10 67 400 $w=1.7e-07 $l=1.13284e-06 $layer=licon1_PDIFF $count=1 $X=15.345
+ $Y=1.835 $X2=15.485 $Y2=2.9
r359 9 150 400 $w=1.7e-07 $l=3.53129e-07 $layer=licon1_PDIFF $count=1 $X=14.485
+ $Y=1.835 $X2=14.625 $Y2=2.125
r360 9 57 400 $w=1.7e-07 $l=1.13284e-06 $layer=licon1_PDIFF $count=1 $X=14.485
+ $Y=1.835 $X2=14.625 $Y2=2.9
r361 8 132 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=21.365
+ $Y=0.235 $X2=21.505 $Y2=0.36
r362 7 122 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=20.505
+ $Y=0.235 $X2=20.645 $Y2=0.36
r363 6 112 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=19.645
+ $Y=0.235 $X2=19.785 $Y2=0.36
r364 5 102 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=18.785
+ $Y=0.235 $X2=18.925 $Y2=0.36
r365 4 92 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=17.925
+ $Y=0.235 $X2=18.065 $Y2=0.36
r366 3 82 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=17.065
+ $Y=0.235 $X2=17.205 $Y2=0.36
r367 2 72 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=16.205
+ $Y=0.235 $X2=16.345 $Y2=0.36
r368 1 63 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=15.34
+ $Y=0.235 $X2=15.485 $Y2=0.36
.ends

.subckt PM_SKY130_FD_SC_LP__BUSDRIVERNOVLPSLEEP_20%VGND 1 2 3 4 5 6 7 8 9 10 11
+ 12 13 14 15 16 51 57 61 65 69 71 75 79 83 87 91 93 97 101 105 109 112 113 115
+ 116 118 119 120 124 126 127 129 130 132 133 135 136 137 138 140 141 143 144
+ 146 147 148 163 181 216 217 224 228 231 233 236 239
c290 75 0 1.0911e-19 $X=10.885 $Y=0.38
r291 239 240 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=18.48 $Y=0
+ $X2=18.48 $Y2=0
r292 236 237 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.2 $Y=0
+ $X2=13.2 $Y2=0
r293 233 234 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.8 $Y=0
+ $X2=10.8 $Y2=0
r294 230 231 9.96101 $w=5.68e-07 $l=1.65e-07 $layer=LI1_cond $X=10.025 $Y=0.2
+ $X2=10.19 $Y2=0.2
r295 227 234 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=9.84 $Y=0
+ $X2=10.8 $Y2=0
r296 226 230 3.88201 $w=5.68e-07 $l=1.85e-07 $layer=LI1_cond $X=9.84 $Y=0.2
+ $X2=10.025 $Y2=0.2
r297 226 228 14.5775 $w=5.68e-07 $l=3.85e-07 $layer=LI1_cond $X=9.84 $Y=0.2
+ $X2=9.455 $Y2=0.2
r298 226 227 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=0
+ $X2=9.84 $Y2=0
r299 222 224 7.86729 $w=5.58e-07 $l=7e-08 $layer=LI1_cond $X=5.04 $Y=0.195
+ $X2=5.11 $Y2=0.195
r300 222 223 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.04 $Y=0
+ $X2=5.04 $Y2=0
r301 220 222 2.02906 $w=5.58e-07 $l=9.5e-08 $layer=LI1_cond $X=4.945 $Y=0.195
+ $X2=5.04 $Y2=0.195
r302 216 217 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=23.28 $Y=0
+ $X2=23.28 $Y2=0
r303 214 217 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=21.36 $Y=0
+ $X2=23.28 $Y2=0
r304 213 216 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=21.36 $Y=0
+ $X2=23.28 $Y2=0
r305 213 214 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=21.36 $Y=0
+ $X2=21.36 $Y2=0
r306 211 214 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=20.88 $Y=0
+ $X2=21.36 $Y2=0
r307 210 211 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=20.88 $Y=0
+ $X2=20.88 $Y2=0
r308 208 211 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=19.92 $Y=0
+ $X2=20.88 $Y2=0
r309 207 208 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=19.92 $Y=0
+ $X2=19.92 $Y2=0
r310 205 208 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=18.96 $Y=0
+ $X2=19.92 $Y2=0
r311 205 240 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=18.96 $Y=0
+ $X2=18.48 $Y2=0
r312 204 205 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=18.96 $Y=0
+ $X2=18.96 $Y2=0
r313 202 239 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=18.58 $Y=0
+ $X2=18.495 $Y2=0
r314 202 204 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=18.58 $Y=0
+ $X2=18.96 $Y2=0
r315 201 240 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=17.52 $Y=0
+ $X2=18.48 $Y2=0
r316 200 201 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=17.52 $Y=0
+ $X2=17.52 $Y2=0
r317 198 201 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=16.56 $Y=0
+ $X2=17.52 $Y2=0
r318 197 198 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=16.56 $Y=0
+ $X2=16.56 $Y2=0
r319 195 198 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=15.6 $Y=0
+ $X2=16.56 $Y2=0
r320 194 195 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=15.6 $Y=0
+ $X2=15.6 $Y2=0
r321 192 195 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=13.68 $Y=0
+ $X2=15.6 $Y2=0
r322 192 237 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.68 $Y=0
+ $X2=13.2 $Y2=0
r323 191 194 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=13.68 $Y=0
+ $X2=15.6 $Y2=0
r324 191 192 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=13.68 $Y=0
+ $X2=13.68 $Y2=0
r325 189 236 8.23795 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=13.365 $Y=0
+ $X2=13.21 $Y2=0
r326 189 191 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=13.365 $Y=0
+ $X2=13.68 $Y2=0
r327 188 237 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.72 $Y=0
+ $X2=13.2 $Y2=0
r328 187 188 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=12.72 $Y=0
+ $X2=12.72 $Y2=0
r329 185 234 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=0
+ $X2=10.8 $Y2=0
r330 184 187 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=11.28 $Y=0
+ $X2=12.72 $Y2=0
r331 184 185 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.28 $Y=0
+ $X2=11.28 $Y2=0
r332 182 233 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.05 $Y=0
+ $X2=10.885 $Y2=0
r333 182 184 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=11.05 $Y=0
+ $X2=11.28 $Y2=0
r334 181 236 8.23795 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=13.055 $Y=0
+ $X2=13.21 $Y2=0
r335 181 187 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=13.055 $Y=0
+ $X2=12.72 $Y2=0
r336 180 227 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=0
+ $X2=9.84 $Y2=0
r337 179 228 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=9.36 $Y=0
+ $X2=9.455 $Y2=0
r338 179 180 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.36 $Y=0
+ $X2=9.36 $Y2=0
r339 176 180 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=8.4 $Y=0
+ $X2=9.36 $Y2=0
r340 175 176 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r341 173 176 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.44 $Y=0
+ $X2=8.4 $Y2=0
r342 172 175 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=7.44 $Y=0 $X2=8.4
+ $Y2=0
r343 172 173 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=7.44 $Y=0
+ $X2=7.44 $Y2=0
r344 170 173 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0
+ $X2=7.44 $Y2=0
r345 170 223 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=6.96 $Y=0
+ $X2=5.04 $Y2=0
r346 169 224 120.695 $w=1.68e-07 $l=1.85e-06 $layer=LI1_cond $X=6.96 $Y=0
+ $X2=5.11 $Y2=0
r347 169 170 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.96 $Y=0
+ $X2=6.96 $Y2=0
r348 166 223 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0
+ $X2=5.04 $Y2=0
r349 165 166 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=0
+ $X2=4.56 $Y2=0
r350 163 220 2.45623 $w=5.58e-07 $l=1.15e-07 $layer=LI1_cond $X=4.83 $Y=0.195
+ $X2=4.945 $Y2=0.195
r351 163 165 5.76681 $w=5.58e-07 $l=2.7e-07 $layer=LI1_cond $X=4.83 $Y=0.195
+ $X2=4.56 $Y2=0.195
r352 162 166 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=0
+ $X2=4.56 $Y2=0
r353 161 162 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r354 159 162 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0
+ $X2=3.6 $Y2=0
r355 158 159 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0
+ $X2=2.64 $Y2=0
r356 156 159 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0
+ $X2=2.64 $Y2=0
r357 155 156 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0
+ $X2=1.68 $Y2=0
r358 152 156 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0
+ $X2=1.68 $Y2=0
r359 151 152 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0
+ $X2=0.72 $Y2=0
r360 148 188 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=11.76 $Y=0
+ $X2=12.72 $Y2=0
r361 148 185 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.76 $Y=0
+ $X2=11.28 $Y2=0
r362 146 210 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=20.99 $Y=0
+ $X2=20.88 $Y2=0
r363 146 147 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=20.99 $Y=0
+ $X2=21.075 $Y2=0
r364 145 213 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=21.16 $Y=0
+ $X2=21.36 $Y2=0
r365 145 147 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=21.16 $Y=0
+ $X2=21.075 $Y2=0
r366 143 207 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=20.13 $Y=0
+ $X2=19.92 $Y2=0
r367 143 144 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=20.13 $Y=0
+ $X2=20.215 $Y2=0
r368 142 210 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=20.3 $Y=0
+ $X2=20.88 $Y2=0
r369 142 144 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=20.3 $Y=0
+ $X2=20.215 $Y2=0
r370 140 204 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=19.27 $Y=0
+ $X2=18.96 $Y2=0
r371 140 141 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=19.27 $Y=0
+ $X2=19.355 $Y2=0
r372 139 207 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=19.44 $Y=0
+ $X2=19.92 $Y2=0
r373 139 141 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=19.44 $Y=0
+ $X2=19.355 $Y2=0
r374 137 200 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=17.55 $Y=0
+ $X2=17.52 $Y2=0
r375 137 138 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=17.55 $Y=0
+ $X2=17.635 $Y2=0
r376 135 197 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=16.69 $Y=0
+ $X2=16.56 $Y2=0
r377 135 136 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=16.69 $Y=0
+ $X2=16.775 $Y2=0
r378 134 200 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=16.86 $Y=0
+ $X2=17.52 $Y2=0
r379 134 136 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=16.86 $Y=0
+ $X2=16.775 $Y2=0
r380 132 194 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=15.83 $Y=0
+ $X2=15.6 $Y2=0
r381 132 133 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=15.83 $Y=0
+ $X2=15.915 $Y2=0
r382 131 197 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=16 $Y=0 $X2=16.56
+ $Y2=0
r383 131 133 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=16 $Y=0 $X2=15.915
+ $Y2=0
r384 129 175 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=8.415 $Y=0
+ $X2=8.4 $Y2=0
r385 129 130 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=8.415 $Y=0
+ $X2=8.6 $Y2=0
r386 128 179 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=8.785 $Y=0
+ $X2=9.36 $Y2=0
r387 128 130 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=8.785 $Y=0
+ $X2=8.6 $Y2=0
r388 126 169 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=6.975 $Y=0
+ $X2=6.96 $Y2=0
r389 126 127 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.975 $Y=0
+ $X2=7.1 $Y2=0
r390 125 172 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=7.225 $Y=0
+ $X2=7.44 $Y2=0
r391 125 127 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.225 $Y=0
+ $X2=7.1 $Y2=0
r392 124 161 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=3.675 $Y=0
+ $X2=3.6 $Y2=0
r393 123 124 9.89636 $w=5.58e-07 $l=1.65e-07 $layer=LI1_cond $X=3.84 $Y=0.195
+ $X2=3.675 $Y2=0.195
r394 120 165 6.94153 $w=5.58e-07 $l=3.25e-07 $layer=LI1_cond $X=4.235 $Y=0.195
+ $X2=4.56 $Y2=0.195
r395 120 123 8.43662 $w=5.58e-07 $l=3.95e-07 $layer=LI1_cond $X=4.235 $Y=0.195
+ $X2=3.84 $Y2=0.195
r396 118 158 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=2.72 $Y=0 $X2=2.64
+ $Y2=0
r397 118 119 7.54988 $w=1.7e-07 $l=1.37e-07 $layer=LI1_cond $X=2.72 $Y=0
+ $X2=2.857 $Y2=0
r398 117 161 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=2.995 $Y=0
+ $X2=3.6 $Y2=0
r399 117 119 7.54988 $w=1.7e-07 $l=1.38e-07 $layer=LI1_cond $X=2.995 $Y=0
+ $X2=2.857 $Y2=0
r400 115 155 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=1.805 $Y=0
+ $X2=1.68 $Y2=0
r401 115 116 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.805 $Y=0
+ $X2=1.97 $Y2=0
r402 114 158 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=2.135 $Y=0
+ $X2=2.64 $Y2=0
r403 114 116 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.135 $Y=0
+ $X2=1.97 $Y2=0
r404 112 151 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=0.945 $Y=0
+ $X2=0.72 $Y2=0
r405 112 113 8.14251 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=0.945 $Y=0
+ $X2=1.097 $Y2=0
r406 111 155 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=1.25 $Y=0
+ $X2=1.68 $Y2=0
r407 111 113 8.14251 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=1.25 $Y=0
+ $X2=1.097 $Y2=0
r408 107 147 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=21.075 $Y=0.085
+ $X2=21.075 $Y2=0
r409 107 109 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=21.075 $Y=0.085
+ $X2=21.075 $Y2=0.36
r410 103 144 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=20.215 $Y=0.085
+ $X2=20.215 $Y2=0
r411 103 105 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=20.215 $Y=0.085
+ $X2=20.215 $Y2=0.36
r412 99 141 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=19.355 $Y=0.085
+ $X2=19.355 $Y2=0
r413 99 101 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=19.355 $Y=0.085
+ $X2=19.355 $Y2=0.36
r414 95 239 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=18.495 $Y=0.085
+ $X2=18.495 $Y2=0
r415 95 97 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=18.495 $Y=0.085
+ $X2=18.495 $Y2=0.36
r416 94 138 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=17.72 $Y=0
+ $X2=17.635 $Y2=0
r417 93 239 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=18.41 $Y=0
+ $X2=18.495 $Y2=0
r418 93 94 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=18.41 $Y=0 $X2=17.72
+ $Y2=0
r419 89 138 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=17.635 $Y=0.085
+ $X2=17.635 $Y2=0
r420 89 91 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=17.635 $Y=0.085
+ $X2=17.635 $Y2=0.36
r421 85 136 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=16.775 $Y=0.085
+ $X2=16.775 $Y2=0
r422 85 87 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=16.775 $Y=0.085
+ $X2=16.775 $Y2=0.36
r423 81 133 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=15.915 $Y=0.085
+ $X2=15.915 $Y2=0
r424 81 83 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=15.915 $Y=0.085
+ $X2=15.915 $Y2=0.36
r425 77 236 0.701276 $w=3.1e-07 $l=8.5e-08 $layer=LI1_cond $X=13.21 $Y=0.085
+ $X2=13.21 $Y2=0
r426 77 79 18.7737 $w=3.08e-07 $l=5.05e-07 $layer=LI1_cond $X=13.21 $Y=0.085
+ $X2=13.21 $Y2=0.59
r427 73 233 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.885 $Y=0.085
+ $X2=10.885 $Y2=0
r428 73 75 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=10.885 $Y=0.085
+ $X2=10.885 $Y2=0.38
r429 71 233 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.72 $Y=0
+ $X2=10.885 $Y2=0
r430 71 231 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=10.72 $Y=0
+ $X2=10.19 $Y2=0
r431 67 130 1.24149 $w=3.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.6 $Y=0.085
+ $X2=8.6 $Y2=0
r432 67 69 9.1884 $w=3.68e-07 $l=2.95e-07 $layer=LI1_cond $X=8.6 $Y=0.085
+ $X2=8.6 $Y2=0.38
r433 63 127 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.1 $Y=0.085
+ $X2=7.1 $Y2=0
r434 63 65 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=7.1 $Y=0.085 $X2=7.1
+ $Y2=0.515
r435 59 119 0.316938 $w=2.75e-07 $l=8.5e-08 $layer=LI1_cond $X=2.857 $Y=0.085
+ $X2=2.857 $Y2=0
r436 59 61 12.5721 $w=2.73e-07 $l=3e-07 $layer=LI1_cond $X=2.857 $Y=0.085
+ $X2=2.857 $Y2=0.385
r437 55 116 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.97 $Y=0.085
+ $X2=1.97 $Y2=0
r438 55 57 15.3659 $w=3.28e-07 $l=4.4e-07 $layer=LI1_cond $X=1.97 $Y=0.085
+ $X2=1.97 $Y2=0.525
r439 51 53 18.7036 $w=3.03e-07 $l=4.95e-07 $layer=LI1_cond $X=1.097 $Y=0.36
+ $X2=1.097 $Y2=0.855
r440 49 113 0.649941 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.097 $Y=0.085
+ $X2=1.097 $Y2=0
r441 49 51 10.3909 $w=3.03e-07 $l=2.75e-07 $layer=LI1_cond $X=1.097 $Y=0.085
+ $X2=1.097 $Y2=0.36
r442 16 109 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=20.935
+ $Y=0.235 $X2=21.075 $Y2=0.36
r443 15 105 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=20.075
+ $Y=0.235 $X2=20.215 $Y2=0.36
r444 14 101 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=19.215
+ $Y=0.235 $X2=19.355 $Y2=0.36
r445 13 97 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=18.355
+ $Y=0.235 $X2=18.495 $Y2=0.36
r446 12 91 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=17.495
+ $Y=0.235 $X2=17.635 $Y2=0.36
r447 11 87 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=16.635
+ $Y=0.235 $X2=16.775 $Y2=0.36
r448 10 83 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=15.775
+ $Y=0.235 $X2=15.915 $Y2=0.36
r449 9 79 182 $w=1.7e-07 $l=4.41871e-07 $layer=licon1_NDIFF $count=1 $X=13.01
+ $Y=0.235 $X2=13.205 $Y2=0.59
r450 8 75 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=10.745
+ $Y=0.235 $X2=10.885 $Y2=0.38
r451 7 230 91 $w=1.7e-07 $l=6.04276e-07 $layer=licon1_NDIFF $count=2 $X=9.48
+ $Y=0.235 $X2=10.025 $Y2=0.36
r452 6 69 182 $w=1.7e-07 $l=5.37634e-07 $layer=licon1_NDIFF $count=1 $X=8.11
+ $Y=0.235 $X2=8.58 $Y2=0.38
r453 5 65 182 $w=1.7e-07 $l=3.36749e-07 $layer=licon1_NDIFF $count=1 $X=7.015
+ $Y=0.235 $X2=7.14 $Y2=0.515
r454 4 220 91 $w=1.7e-07 $l=1.36607e-06 $layer=licon1_NDIFF $count=2 $X=3.64
+ $Y=0.235 $X2=4.945 $Y2=0.36
r455 4 123 91 $w=1.7e-07 $l=2.54951e-07 $layer=licon1_NDIFF $count=2 $X=3.64
+ $Y=0.235 $X2=3.84 $Y2=0.36
r456 3 61 91 $w=1.7e-07 $l=2.08567e-07 $layer=licon1_NDIFF $count=2 $X=2.69
+ $Y=0.235 $X2=2.83 $Y2=0.385
r457 2 57 182 $w=1.7e-07 $l=3.53129e-07 $layer=licon1_NDIFF $count=1 $X=1.83
+ $Y=0.235 $X2=1.97 $Y2=0.525
r458 1 53 182 $w=1.7e-07 $l=7.13022e-07 $layer=licon1_NDIFF $count=1 $X=0.91
+ $Y=0.235 $X2=1.11 $Y2=0.855
r459 1 51 182 $w=1.7e-07 $l=2.54951e-07 $layer=licon1_NDIFF $count=1 $X=0.91
+ $Y=0.235 $X2=1.11 $Y2=0.36
.ends

.subckt PM_SKY130_FD_SC_LP__BUSDRIVERNOVLPSLEEP_20%A_2519_47# 1 2 3 11 12 13 14
+ 15 16 21 27
c53 12 0 8.57257e-20 $X=13.575 $Y=1.01
r54 17 25 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.905 $Y=0.35
+ $X2=13.74 $Y2=0.35
r55 16 27 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=14.54 $Y=0.35
+ $X2=14.665 $Y2=0.35
r56 16 17 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=14.54 $Y=0.35
+ $X2=13.905 $Y2=0.35
r57 14 25 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=13.74 $Y=0.435
+ $X2=13.74 $Y2=0.35
r58 14 15 17.112 $w=3.28e-07 $l=4.9e-07 $layer=LI1_cond $X=13.74 $Y=0.435
+ $X2=13.74 $Y2=0.925
r59 12 15 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=13.575 $Y=1.01
+ $X2=13.74 $Y2=0.925
r60 12 13 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=13.575 $Y=1.01
+ $X2=12.885 $Y2=1.01
r61 11 13 6.89401 $w=1.7e-07 $l=1.39155e-07 $layer=LI1_cond $X=12.782 $Y=0.925
+ $X2=12.885 $Y2=1.01
r62 11 21 24.8869 $w=2.03e-07 $l=4.6e-07 $layer=LI1_cond $X=12.782 $Y=0.925
+ $X2=12.782 $Y2=0.465
r63 3 27 91 $w=1.7e-07 $l=2.64953e-07 $layer=licon1_NDIFF $count=2 $X=14.46
+ $Y=0.235 $X2=14.625 $Y2=0.43
r64 2 25 91 $w=1.7e-07 $l=2.86356e-07 $layer=licon1_NDIFF $count=2 $X=13.535
+ $Y=0.235 $X2=13.74 $Y2=0.43
r65 1 21 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=12.595
+ $Y=0.235 $X2=12.72 $Y2=0.38
.ends

