* File: sky130_fd_sc_lp__a41oi_m.spice
* Created: Fri Aug 28 10:04:01 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__a41oi_m.pex.spice"
.subckt sky130_fd_sc_lp__a41oi_m  VNB VPB B1 A1 A2 A3 A4 Y VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Y	Y
* A4	A4
* A3	A3
* A2	A2
* A1	A1
* B1	B1
* VPB	VPB
* VNB	VNB
MM1008 N_Y_M1008_d N_B1_M1008_g N_VGND_M1008_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75001.8
+ A=0.063 P=1.14 MULT=1
MM1001 A_300_47# N_A1_M1001_g N_Y_M1008_d VNB NSHORT L=0.15 W=0.42 AD=0.0441
+ AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.6 SB=75001.4
+ A=0.063 P=1.14 MULT=1
MM1003 A_372_47# N_A2_M1003_g A_300_47# VNB NSHORT L=0.15 W=0.42 AD=0.0672
+ AS=0.0441 PD=0.74 PS=0.63 NRD=30 NRS=14.28 M=1 R=2.8 SA=75001 SB=75001 A=0.063
+ P=1.14 MULT=1
MM1002 A_466_47# N_A3_M1002_g A_372_47# VNB NSHORT L=0.15 W=0.42 AD=0.0441
+ AS=0.0672 PD=0.63 PS=0.74 NRD=14.28 NRS=30 M=1 R=2.8 SA=75001.4 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1004 N_VGND_M1004_d N_A4_M1004_g A_466_47# VNB NSHORT L=0.15 W=0.42 AD=0.1113
+ AS=0.0441 PD=1.37 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.8 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1007 N_A_186_531#_M1007_d N_B1_M1007_g N_Y_M1007_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0588 AS=0.2331 PD=0.7 PS=1.95 NRD=0 NRS=136.009 M=1 R=2.8 SA=75000.5
+ SB=75001.9 A=0.063 P=1.14 MULT=1
MM1005 N_VPWR_M1005_d N_A1_M1005_g N_A_186_531#_M1007_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.9
+ SB=75001.5 A=0.063 P=1.14 MULT=1
MM1009 N_A_186_531#_M1009_d N_A2_M1009_g N_VPWR_M1005_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.3
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1006 N_VPWR_M1006_d N_A3_M1006_g N_A_186_531#_M1009_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.8
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1000 N_A_186_531#_M1000_d N_A4_M1000_g N_VPWR_M1006_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75002.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9751 P=11.21
*
.include "sky130_fd_sc_lp__a41oi_m.pxi.spice"
*
.ends
*
*
