* File: sky130_fd_sc_lp__ebufn_lp.pxi.spice
* Created: Fri Aug 28 10:32:11 2020
* 
x_PM_SKY130_FD_SC_LP__EBUFN_LP%A N_A_M1010_g N_A_M1004_g N_A_M1000_g N_A_M1001_g
+ A A N_A_c_75_n N_A_c_76_n PM_SKY130_FD_SC_LP__EBUFN_LP%A
x_PM_SKY130_FD_SC_LP__EBUFN_LP%A_242_237# N_A_242_237#_M1003_d
+ N_A_242_237#_M1006_d N_A_242_237#_M1009_g N_A_242_237#_c_111_n
+ N_A_242_237#_c_112_n N_A_242_237#_c_113_n N_A_242_237#_c_114_n
+ N_A_242_237#_c_175_p N_A_242_237#_c_115_n N_A_242_237#_c_116_n
+ N_A_242_237#_c_117_n N_A_242_237#_c_118_n N_A_242_237#_c_122_n
+ N_A_242_237#_c_119_n N_A_242_237#_c_120_n N_A_242_237#_c_121_n
+ PM_SKY130_FD_SC_LP__EBUFN_LP%A_242_237#
x_PM_SKY130_FD_SC_LP__EBUFN_LP%A_29_483# N_A_29_483#_M1004_s N_A_29_483#_M1010_s
+ N_A_29_483#_M1008_g N_A_29_483#_c_187_n N_A_29_483#_M1002_g
+ N_A_29_483#_c_188_n N_A_29_483#_c_195_n N_A_29_483#_c_196_n
+ N_A_29_483#_c_197_n N_A_29_483#_c_198_n N_A_29_483#_c_189_n
+ N_A_29_483#_c_190_n N_A_29_483#_c_200_n N_A_29_483#_c_191_n
+ PM_SKY130_FD_SC_LP__EBUFN_LP%A_29_483#
x_PM_SKY130_FD_SC_LP__EBUFN_LP%TE_B N_TE_B_M1007_g N_TE_B_c_256_n N_TE_B_c_257_n
+ N_TE_B_M1011_g N_TE_B_M1005_g N_TE_B_c_260_n N_TE_B_M1003_g N_TE_B_c_266_n
+ N_TE_B_M1006_g N_TE_B_c_262_n N_TE_B_c_268_n TE_B TE_B
+ PM_SKY130_FD_SC_LP__EBUFN_LP%TE_B
x_PM_SKY130_FD_SC_LP__EBUFN_LP%VPWR N_VPWR_M1001_d N_VPWR_M1007_d N_VPWR_c_313_n
+ N_VPWR_c_314_n N_VPWR_c_315_n N_VPWR_c_316_n VPWR N_VPWR_c_317_n
+ N_VPWR_c_318_n N_VPWR_c_312_n N_VPWR_c_320_n PM_SKY130_FD_SC_LP__EBUFN_LP%VPWR
x_PM_SKY130_FD_SC_LP__EBUFN_LP%Z N_Z_M1008_d N_Z_M1002_s Z Z Z Z Z Z
+ PM_SKY130_FD_SC_LP__EBUFN_LP%Z
x_PM_SKY130_FD_SC_LP__EBUFN_LP%VGND N_VGND_M1000_d N_VGND_M1005_s N_VGND_c_388_n
+ N_VGND_c_389_n VGND N_VGND_c_390_n N_VGND_c_391_n N_VGND_c_392_n
+ N_VGND_c_393_n N_VGND_c_394_n N_VGND_c_395_n PM_SKY130_FD_SC_LP__EBUFN_LP%VGND
cc_1 VNB N_A_M1004_g 0.0244897f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=0.865
cc_2 VNB N_A_M1000_g 0.0205182f $X=-0.19 $Y=-0.245 $X2=0.895 $Y2=0.865
cc_3 VNB N_A_c_75_n 0.0477494f $X=-0.19 $Y=-0.245 $X2=0.655 $Y2=1.41
cc_4 VNB N_A_c_76_n 0.00122182f $X=-0.19 $Y=-0.245 $X2=0.655 $Y2=1.41
cc_5 VNB N_A_242_237#_c_111_n 0.00825926f $X=-0.19 $Y=-0.245 $X2=0.895 $Y2=0.865
cc_6 VNB N_A_242_237#_c_112_n 0.0317896f $X=-0.19 $Y=-0.245 $X2=0.895 $Y2=1.915
cc_7 VNB N_A_242_237#_c_113_n 0.00165187f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_242_237#_c_114_n 0.0207887f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_9 VNB N_A_242_237#_c_115_n 0.0150324f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_242_237#_c_116_n 0.0173745f $X=-0.19 $Y=-0.245 $X2=0.7 $Y2=1.41
cc_11 VNB N_A_242_237#_c_117_n 0.00684563f $X=-0.19 $Y=-0.245 $X2=0.655 $Y2=1.41
cc_12 VNB N_A_242_237#_c_118_n 0.0228189f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_242_237#_c_119_n 0.00919847f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_242_237#_c_120_n 0.0237347f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_242_237#_c_121_n 0.0185254f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_29_483#_M1008_g 0.0296093f $X=-0.19 $Y=-0.245 $X2=0.895 $Y2=1.245
cc_17 VNB N_A_29_483#_c_187_n 0.0152324f $X=-0.19 $Y=-0.245 $X2=0.895 $Y2=0.865
cc_18 VNB N_A_29_483#_c_188_n 0.0273873f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.95
cc_19 VNB N_A_29_483#_c_189_n 0.00283509f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_29_483#_c_190_n 0.0260212f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_29_483#_c_191_n 0.0395261f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_TE_B_M1007_g 0.0199465f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=2.735
cc_23 VNB N_TE_B_c_256_n 0.0217042f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=1.41
cc_24 VNB N_TE_B_c_257_n 0.0100615f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=0.865
cc_25 VNB N_TE_B_M1011_g 0.00863872f $X=-0.19 $Y=-0.245 $X2=0.895 $Y2=1.245
cc_26 VNB N_TE_B_M1005_g 0.0448129f $X=-0.19 $Y=-0.245 $X2=0.895 $Y2=1.915
cc_27 VNB N_TE_B_c_260_n 0.0533643f $X=-0.19 $Y=-0.245 $X2=0.895 $Y2=2.735
cc_28 VNB N_TE_B_M1003_g 0.0428421f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_29 VNB N_TE_B_c_262_n 0.0197591f $X=-0.19 $Y=-0.245 $X2=0.655 $Y2=1.41
cc_30 VNB TE_B 0.00137398f $X=-0.19 $Y=-0.245 $X2=0.662 $Y2=2.035
cc_31 VNB N_VPWR_c_312_n 0.183584f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB Z 0.0428125f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=0.865
cc_33 VNB N_VGND_c_388_n 0.0150983f $X=-0.19 $Y=-0.245 $X2=0.895 $Y2=1.245
cc_34 VNB N_VGND_c_389_n 0.00973205f $X=-0.19 $Y=-0.245 $X2=0.895 $Y2=2.735
cc_35 VNB N_VGND_c_390_n 0.03444f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_391_n 0.039836f $X=-0.19 $Y=-0.245 $X2=0.662 $Y2=1.41
cc_37 VNB N_VGND_c_392_n 0.0266819f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_393_n 0.25999f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_394_n 0.00525267f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_395_n 0.00513431f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VPB N_A_M1010_g 0.0401762f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=2.735
cc_42 VPB N_A_M1001_g 0.0383385f $X=-0.19 $Y=1.655 $X2=0.895 $Y2=2.735
cc_43 VPB N_A_c_75_n 0.0302667f $X=-0.19 $Y=1.655 $X2=0.655 $Y2=1.41
cc_44 VPB N_A_c_76_n 0.0025801f $X=-0.19 $Y=1.655 $X2=0.655 $Y2=1.41
cc_45 VPB N_A_242_237#_c_122_n 0.0314438f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_46 VPB N_A_242_237#_c_120_n 0.0119903f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_47 VPB N_A_29_483#_c_187_n 0.00573268f $X=-0.19 $Y=1.655 $X2=0.895 $Y2=0.865
cc_48 VPB N_A_29_483#_M1002_g 0.022024f $X=-0.19 $Y=1.655 $X2=0.895 $Y2=2.735
cc_49 VPB N_A_29_483#_c_188_n 0.0348875f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.95
cc_50 VPB N_A_29_483#_c_195_n 0.00374081f $X=-0.19 $Y=1.655 $X2=0.7 $Y2=1.41
cc_51 VPB N_A_29_483#_c_196_n 0.0246742f $X=-0.19 $Y=1.655 $X2=0.662 $Y2=1.41
cc_52 VPB N_A_29_483#_c_197_n 0.0384707f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_53 VPB N_A_29_483#_c_198_n 0.00634098f $X=-0.19 $Y=1.655 $X2=0.662 $Y2=1.665
cc_54 VPB N_A_29_483#_c_189_n 3.90621e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_55 VPB N_A_29_483#_c_200_n 0.0342361f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_56 VPB N_A_29_483#_c_191_n 0.0145503f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_57 VPB N_TE_B_M1007_g 0.0220816f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=2.735
cc_58 VPB N_TE_B_M1011_g 0.031378f $X=-0.19 $Y=1.655 $X2=0.895 $Y2=1.245
cc_59 VPB N_TE_B_c_266_n 0.0219031f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_60 VPB N_TE_B_c_262_n 0.00395679f $X=-0.19 $Y=1.655 $X2=0.655 $Y2=1.41
cc_61 VPB N_TE_B_c_268_n 0.0252384f $X=-0.19 $Y=1.655 $X2=0.662 $Y2=1.665
cc_62 VPB TE_B 0.010624f $X=-0.19 $Y=1.655 $X2=0.662 $Y2=2.035
cc_63 VPB N_VPWR_c_313_n 0.0224696f $X=-0.19 $Y=1.655 $X2=0.895 $Y2=1.245
cc_64 VPB N_VPWR_c_314_n 0.0250657f $X=-0.19 $Y=1.655 $X2=0.895 $Y2=1.915
cc_65 VPB N_VPWR_c_315_n 0.0417303f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_316_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0.7 $Y2=1.41
cc_67 VPB N_VPWR_c_317_n 0.0339091f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_318_n 0.0341808f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_69 VPB N_VPWR_c_312_n 0.101831f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_70 VPB N_VPWR_c_320_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_71 VPB Z 0.00318651f $X=-0.19 $Y=1.655 $X2=0.535 $Y2=0.865
cc_72 VPB Z 0.0255249f $X=-0.19 $Y=1.655 $X2=0.895 $Y2=0.865
cc_73 N_A_M1000_g N_A_242_237#_c_111_n 0.0015484f $X=0.895 $Y=0.865 $X2=0 $Y2=0
cc_74 N_A_c_76_n N_A_242_237#_c_111_n 0.0111442f $X=0.655 $Y=1.41 $X2=0 $Y2=0
cc_75 N_A_M1000_g N_A_242_237#_c_112_n 0.0179808f $X=0.895 $Y=0.865 $X2=0 $Y2=0
cc_76 N_A_c_76_n N_A_242_237#_c_112_n 2.82003e-19 $X=0.655 $Y=1.41 $X2=0 $Y2=0
cc_77 N_A_M1000_g N_A_242_237#_c_121_n 0.010363f $X=0.895 $Y=0.865 $X2=0 $Y2=0
cc_78 N_A_M1004_g N_A_29_483#_c_188_n 0.00411368f $X=0.535 $Y=0.865 $X2=0 $Y2=0
cc_79 N_A_c_75_n N_A_29_483#_c_188_n 0.0292061f $X=0.655 $Y=1.41 $X2=0 $Y2=0
cc_80 N_A_c_76_n N_A_29_483#_c_188_n 0.0615185f $X=0.655 $Y=1.41 $X2=0 $Y2=0
cc_81 N_A_M1010_g N_A_29_483#_c_195_n 0.0093864f $X=0.505 $Y=2.735 $X2=0 $Y2=0
cc_82 N_A_M1001_g N_A_29_483#_c_195_n 0.016689f $X=0.895 $Y=2.735 $X2=0 $Y2=0
cc_83 N_A_c_75_n N_A_29_483#_c_195_n 2.42696e-19 $X=0.655 $Y=1.41 $X2=0 $Y2=0
cc_84 N_A_c_76_n N_A_29_483#_c_195_n 0.0215412f $X=0.655 $Y=1.41 $X2=0 $Y2=0
cc_85 N_A_c_75_n N_A_29_483#_c_196_n 0.0167091f $X=0.655 $Y=1.41 $X2=0 $Y2=0
cc_86 N_A_c_76_n N_A_29_483#_c_196_n 0.0221681f $X=0.655 $Y=1.41 $X2=0 $Y2=0
cc_87 N_A_c_75_n N_A_29_483#_c_198_n 0.00514843f $X=0.655 $Y=1.41 $X2=0 $Y2=0
cc_88 N_A_c_76_n N_A_29_483#_c_198_n 0.0143781f $X=0.655 $Y=1.41 $X2=0 $Y2=0
cc_89 N_A_M1004_g N_A_29_483#_c_190_n 0.0104468f $X=0.535 $Y=0.865 $X2=0 $Y2=0
cc_90 N_A_M1000_g N_A_29_483#_c_190_n 0.00140201f $X=0.895 $Y=0.865 $X2=0 $Y2=0
cc_91 N_A_M1010_g N_A_29_483#_c_200_n 0.0115938f $X=0.505 $Y=2.735 $X2=0 $Y2=0
cc_92 N_A_M1001_g N_A_29_483#_c_200_n 0.00252509f $X=0.895 $Y=2.735 $X2=0 $Y2=0
cc_93 N_A_M1001_g N_VPWR_c_313_n 0.0182872f $X=0.895 $Y=2.735 $X2=0 $Y2=0
cc_94 N_A_M1010_g N_VPWR_c_315_n 0.00511358f $X=0.505 $Y=2.735 $X2=0 $Y2=0
cc_95 N_A_M1001_g N_VPWR_c_315_n 0.00545548f $X=0.895 $Y=2.735 $X2=0 $Y2=0
cc_96 N_A_M1010_g N_VPWR_c_312_n 0.00639603f $X=0.505 $Y=2.735 $X2=0 $Y2=0
cc_97 N_A_M1001_g N_VPWR_c_312_n 0.00682061f $X=0.895 $Y=2.735 $X2=0 $Y2=0
cc_98 N_A_M1000_g N_VGND_c_388_n 0.00834995f $X=0.895 $Y=0.865 $X2=0 $Y2=0
cc_99 N_A_M1004_g N_VGND_c_390_n 0.00385415f $X=0.535 $Y=0.865 $X2=0 $Y2=0
cc_100 N_A_M1000_g N_VGND_c_390_n 0.00399858f $X=0.895 $Y=0.865 $X2=0 $Y2=0
cc_101 N_A_M1004_g N_VGND_c_393_n 0.0046122f $X=0.535 $Y=0.865 $X2=0 $Y2=0
cc_102 N_A_M1000_g N_VGND_c_393_n 0.0046122f $X=0.895 $Y=0.865 $X2=0 $Y2=0
cc_103 N_A_242_237#_c_111_n N_A_29_483#_M1008_g 0.00390888f $X=1.565 $Y=1.35
+ $X2=0 $Y2=0
cc_104 N_A_242_237#_c_113_n N_A_29_483#_M1008_g 0.00320806f $X=1.65 $Y=1.185
+ $X2=0 $Y2=0
cc_105 N_A_242_237#_c_114_n N_A_29_483#_M1008_g 0.0149072f $X=2.745 $Y=0.34
+ $X2=0 $Y2=0
cc_106 N_A_242_237#_c_121_n N_A_29_483#_M1008_g 0.0334873f $X=1.375 $Y=1.185
+ $X2=0 $Y2=0
cc_107 N_A_242_237#_c_111_n N_A_29_483#_c_197_n 0.0411005f $X=1.565 $Y=1.35
+ $X2=0 $Y2=0
cc_108 N_A_242_237#_c_112_n N_A_29_483#_c_197_n 0.00798977f $X=1.375 $Y=1.35
+ $X2=0 $Y2=0
cc_109 N_A_242_237#_c_111_n N_A_29_483#_c_189_n 0.0140339f $X=1.565 $Y=1.35
+ $X2=0 $Y2=0
cc_110 N_A_242_237#_c_112_n N_A_29_483#_c_191_n 0.0334873f $X=1.375 $Y=1.35
+ $X2=0 $Y2=0
cc_111 N_A_242_237#_c_116_n N_TE_B_c_257_n 0.0180868f $X=3.875 $Y=0.92 $X2=0
+ $Y2=0
cc_112 N_A_242_237#_c_117_n N_TE_B_c_257_n 0.00483855f $X=2.915 $Y=0.92 $X2=0
+ $Y2=0
cc_113 N_A_242_237#_c_122_n N_TE_B_M1011_g 0.00202956f $X=4.04 $Y=2.15 $X2=0
+ $Y2=0
cc_114 N_A_242_237#_c_120_n N_TE_B_M1011_g 8.1286e-19 $X=4.04 $Y=1.985 $X2=0
+ $Y2=0
cc_115 N_A_242_237#_c_115_n N_TE_B_M1005_g 0.00458181f $X=2.83 $Y=0.835 $X2=0
+ $Y2=0
cc_116 N_A_242_237#_c_116_n N_TE_B_M1005_g 0.0147831f $X=3.875 $Y=0.92 $X2=0
+ $Y2=0
cc_117 N_A_242_237#_c_118_n N_TE_B_M1005_g 0.00196547f $X=4.04 $Y=0.465 $X2=0
+ $Y2=0
cc_118 N_A_242_237#_c_116_n N_TE_B_c_260_n 2.11484e-19 $X=3.875 $Y=0.92 $X2=0
+ $Y2=0
cc_119 N_A_242_237#_c_119_n N_TE_B_c_260_n 0.00573152f $X=4.04 $Y=0.92 $X2=0
+ $Y2=0
cc_120 N_A_242_237#_c_120_n N_TE_B_c_260_n 0.0118244f $X=4.04 $Y=1.985 $X2=0
+ $Y2=0
cc_121 N_A_242_237#_c_116_n N_TE_B_M1003_g 0.010909f $X=3.875 $Y=0.92 $X2=0
+ $Y2=0
cc_122 N_A_242_237#_c_118_n N_TE_B_M1003_g 0.013569f $X=4.04 $Y=0.465 $X2=0
+ $Y2=0
cc_123 N_A_242_237#_c_119_n N_TE_B_M1003_g 0.00501393f $X=4.04 $Y=0.92 $X2=0
+ $Y2=0
cc_124 N_A_242_237#_c_120_n N_TE_B_M1003_g 0.00424967f $X=4.04 $Y=1.985 $X2=0
+ $Y2=0
cc_125 N_A_242_237#_c_122_n N_TE_B_c_266_n 0.014206f $X=4.04 $Y=2.15 $X2=0 $Y2=0
cc_126 N_A_242_237#_c_120_n N_TE_B_c_266_n 0.00140486f $X=4.04 $Y=1.985 $X2=0
+ $Y2=0
cc_127 N_A_242_237#_c_120_n N_TE_B_c_262_n 0.0157287f $X=4.04 $Y=1.985 $X2=0
+ $Y2=0
cc_128 N_A_242_237#_c_122_n N_TE_B_c_268_n 0.00620649f $X=4.04 $Y=2.15 $X2=0
+ $Y2=0
cc_129 N_A_242_237#_c_120_n N_TE_B_c_268_n 0.00966862f $X=4.04 $Y=1.985 $X2=0
+ $Y2=0
cc_130 N_A_242_237#_c_116_n TE_B 0.0255304f $X=3.875 $Y=0.92 $X2=0 $Y2=0
cc_131 N_A_242_237#_c_120_n TE_B 0.0312739f $X=4.04 $Y=1.985 $X2=0 $Y2=0
cc_132 N_A_242_237#_c_122_n N_VPWR_c_314_n 0.0194249f $X=4.04 $Y=2.15 $X2=0
+ $Y2=0
cc_133 N_A_242_237#_c_122_n N_VPWR_c_318_n 0.00619475f $X=4.04 $Y=2.15 $X2=0
+ $Y2=0
cc_134 N_A_242_237#_c_122_n N_VPWR_c_312_n 0.00970591f $X=4.04 $Y=2.15 $X2=0
+ $Y2=0
cc_135 N_A_242_237#_c_114_n N_Z_M1008_d 0.0055411f $X=2.745 $Y=0.34 $X2=-0.19
+ $Y2=-0.245
cc_136 N_A_242_237#_c_111_n Z 0.00526815f $X=1.565 $Y=1.35 $X2=0 $Y2=0
cc_137 N_A_242_237#_c_113_n Z 0.027655f $X=1.65 $Y=1.185 $X2=0 $Y2=0
cc_138 N_A_242_237#_c_114_n Z 0.0398343f $X=2.745 $Y=0.34 $X2=0 $Y2=0
cc_139 N_A_242_237#_c_115_n Z 0.0121867f $X=2.83 $Y=0.835 $X2=0 $Y2=0
cc_140 N_A_242_237#_c_117_n Z 0.0105341f $X=2.915 $Y=0.92 $X2=0 $Y2=0
cc_141 N_A_242_237#_c_111_n N_VGND_c_388_n 0.0125835f $X=1.565 $Y=1.35 $X2=0
+ $Y2=0
cc_142 N_A_242_237#_c_112_n N_VGND_c_388_n 0.00401953f $X=1.375 $Y=1.35 $X2=0
+ $Y2=0
cc_143 N_A_242_237#_c_121_n N_VGND_c_388_n 0.0132553f $X=1.375 $Y=1.185 $X2=0
+ $Y2=0
cc_144 N_A_242_237#_c_114_n N_VGND_c_389_n 0.0150383f $X=2.745 $Y=0.34 $X2=0
+ $Y2=0
cc_145 N_A_242_237#_c_115_n N_VGND_c_389_n 0.0189907f $X=2.83 $Y=0.835 $X2=0
+ $Y2=0
cc_146 N_A_242_237#_c_116_n N_VGND_c_389_n 0.0268908f $X=3.875 $Y=0.92 $X2=0
+ $Y2=0
cc_147 N_A_242_237#_c_118_n N_VGND_c_389_n 0.0137175f $X=4.04 $Y=0.465 $X2=0
+ $Y2=0
cc_148 N_A_242_237#_c_114_n N_VGND_c_391_n 0.0735751f $X=2.745 $Y=0.34 $X2=0
+ $Y2=0
cc_149 N_A_242_237#_c_175_p N_VGND_c_391_n 0.0104206f $X=1.735 $Y=0.34 $X2=0
+ $Y2=0
cc_150 N_A_242_237#_c_121_n N_VGND_c_391_n 0.00564095f $X=1.375 $Y=1.185 $X2=0
+ $Y2=0
cc_151 N_A_242_237#_c_118_n N_VGND_c_392_n 0.0210519f $X=4.04 $Y=0.465 $X2=0
+ $Y2=0
cc_152 N_A_242_237#_M1003_d N_VGND_c_393_n 0.00232718f $X=3.9 $Y=0.235 $X2=0
+ $Y2=0
cc_153 N_A_242_237#_c_114_n N_VGND_c_393_n 0.0438924f $X=2.745 $Y=0.34 $X2=0
+ $Y2=0
cc_154 N_A_242_237#_c_175_p N_VGND_c_393_n 0.00660921f $X=1.735 $Y=0.34 $X2=0
+ $Y2=0
cc_155 N_A_242_237#_c_116_n N_VGND_c_393_n 0.0211587f $X=3.875 $Y=0.92 $X2=0
+ $Y2=0
cc_156 N_A_242_237#_c_118_n N_VGND_c_393_n 0.0126421f $X=4.04 $Y=0.465 $X2=0
+ $Y2=0
cc_157 N_A_242_237#_c_121_n N_VGND_c_393_n 0.00950947f $X=1.375 $Y=1.185 $X2=0
+ $Y2=0
cc_158 N_A_242_237#_c_113_n A_308_47# 0.00284462f $X=1.65 $Y=1.185 $X2=-0.19
+ $Y2=-0.245
cc_159 N_A_242_237#_c_175_p A_308_47# 0.00126025f $X=1.735 $Y=0.34 $X2=-0.19
+ $Y2=-0.245
cc_160 N_A_29_483#_c_187_n N_TE_B_M1007_g 0.084759f $X=2.425 $Y=1.6 $X2=0 $Y2=0
cc_161 N_A_29_483#_c_191_n N_TE_B_M1007_g 0.00226009f $X=2.235 $Y=1.51 $X2=0
+ $Y2=0
cc_162 N_A_29_483#_c_195_n A_116_483# 0.00236867f $X=1.005 $Y=2.48 $X2=-0.19
+ $Y2=-0.245
cc_163 N_A_29_483#_c_195_n N_VPWR_M1001_d 0.00515788f $X=1.005 $Y=2.48 $X2=-0.19
+ $Y2=-0.245
cc_164 N_A_29_483#_c_195_n N_VPWR_c_313_n 0.0145437f $X=1.005 $Y=2.48 $X2=0
+ $Y2=0
cc_165 N_A_29_483#_c_197_n N_VPWR_c_313_n 0.012401f $X=1.905 $Y=1.77 $X2=0 $Y2=0
cc_166 N_A_29_483#_M1002_g N_VPWR_c_314_n 0.00255107f $X=2.5 $Y=2.465 $X2=0
+ $Y2=0
cc_167 N_A_29_483#_c_200_n N_VPWR_c_315_n 0.0234289f $X=0.29 $Y=2.56 $X2=0 $Y2=0
cc_168 N_A_29_483#_M1002_g N_VPWR_c_317_n 0.00387413f $X=2.5 $Y=2.465 $X2=0
+ $Y2=0
cc_169 N_A_29_483#_M1002_g N_VPWR_c_312_n 0.00672174f $X=2.5 $Y=2.465 $X2=0
+ $Y2=0
cc_170 N_A_29_483#_c_195_n N_VPWR_c_312_n 0.0254408f $X=1.005 $Y=2.48 $X2=0
+ $Y2=0
cc_171 N_A_29_483#_c_200_n N_VPWR_c_312_n 0.0126421f $X=0.29 $Y=2.56 $X2=0 $Y2=0
cc_172 N_A_29_483#_c_197_n N_Z_M1002_s 0.00120658f $X=1.905 $Y=1.77 $X2=0 $Y2=0
cc_173 N_A_29_483#_M1008_g Z 0.0138848f $X=1.855 $Y=0.655 $X2=0 $Y2=0
cc_174 N_A_29_483#_c_187_n Z 0.0153994f $X=2.425 $Y=1.6 $X2=0 $Y2=0
cc_175 N_A_29_483#_M1002_g Z 0.0119307f $X=2.5 $Y=2.465 $X2=0 $Y2=0
cc_176 N_A_29_483#_c_197_n Z 0.0141781f $X=1.905 $Y=1.77 $X2=0 $Y2=0
cc_177 N_A_29_483#_c_189_n Z 0.0545535f $X=2.07 $Y=1.51 $X2=0 $Y2=0
cc_178 N_A_29_483#_c_191_n Z 0.00426042f $X=2.235 $Y=1.51 $X2=0 $Y2=0
cc_179 N_A_29_483#_M1002_g Z 0.0236349f $X=2.5 $Y=2.465 $X2=0 $Y2=0
cc_180 N_A_29_483#_c_197_n Z 0.0102225f $X=1.905 $Y=1.77 $X2=0 $Y2=0
cc_181 N_A_29_483#_c_191_n Z 0.00562815f $X=2.235 $Y=1.51 $X2=0 $Y2=0
cc_182 N_A_29_483#_M1008_g N_VGND_c_388_n 0.00144236f $X=1.855 $Y=0.655 $X2=0
+ $Y2=0
cc_183 N_A_29_483#_c_197_n N_VGND_c_388_n 0.00104901f $X=1.905 $Y=1.77 $X2=0
+ $Y2=0
cc_184 N_A_29_483#_c_198_n N_VGND_c_388_n 0.00368503f $X=1.175 $Y=1.77 $X2=0
+ $Y2=0
cc_185 N_A_29_483#_c_190_n N_VGND_c_388_n 0.0113338f $X=0.32 $Y=0.855 $X2=0
+ $Y2=0
cc_186 N_A_29_483#_c_190_n N_VGND_c_390_n 0.00707271f $X=0.32 $Y=0.855 $X2=0
+ $Y2=0
cc_187 N_A_29_483#_M1008_g N_VGND_c_391_n 0.00357877f $X=1.855 $Y=0.655 $X2=0
+ $Y2=0
cc_188 N_A_29_483#_M1008_g N_VGND_c_393_n 0.00674037f $X=1.855 $Y=0.655 $X2=0
+ $Y2=0
cc_189 N_A_29_483#_c_190_n N_VGND_c_393_n 0.0107231f $X=0.32 $Y=0.855 $X2=0
+ $Y2=0
cc_190 N_TE_B_M1007_g N_VPWR_c_314_n 0.0243337f $X=2.89 $Y=2.465 $X2=0 $Y2=0
cc_191 N_TE_B_c_256_n N_VPWR_c_314_n 0.00628708f $X=3.36 $Y=1.25 $X2=0 $Y2=0
cc_192 N_TE_B_M1011_g N_VPWR_c_314_n 0.0172891f $X=3.435 $Y=2.325 $X2=0 $Y2=0
cc_193 N_TE_B_M1007_g N_VPWR_c_317_n 0.00486043f $X=2.89 $Y=2.465 $X2=0 $Y2=0
cc_194 N_TE_B_M1011_g N_VPWR_c_318_n 0.00385058f $X=3.435 $Y=2.325 $X2=0 $Y2=0
cc_195 N_TE_B_c_266_n N_VPWR_c_318_n 0.00371502f $X=3.825 $Y=1.895 $X2=0 $Y2=0
cc_196 N_TE_B_M1007_g N_VPWR_c_312_n 0.00827383f $X=2.89 $Y=2.465 $X2=0 $Y2=0
cc_197 N_TE_B_M1011_g N_VPWR_c_312_n 0.00453162f $X=3.435 $Y=2.325 $X2=0 $Y2=0
cc_198 N_TE_B_c_266_n N_VPWR_c_312_n 0.00453162f $X=3.825 $Y=1.895 $X2=0 $Y2=0
cc_199 N_TE_B_M1007_g Z 0.0145925f $X=2.89 $Y=2.465 $X2=0 $Y2=0
cc_200 N_TE_B_c_257_n Z 0.00854093f $X=2.965 $Y=1.25 $X2=0 $Y2=0
cc_201 N_TE_B_M1007_g Z 0.00714162f $X=2.89 $Y=2.465 $X2=0 $Y2=0
cc_202 N_TE_B_M1005_g N_VGND_c_389_n 0.0139354f $X=3.465 $Y=0.445 $X2=0 $Y2=0
cc_203 N_TE_B_M1003_g N_VGND_c_389_n 0.00234778f $X=3.825 $Y=0.445 $X2=0 $Y2=0
cc_204 N_TE_B_M1005_g N_VGND_c_392_n 0.00486043f $X=3.465 $Y=0.445 $X2=0 $Y2=0
cc_205 N_TE_B_M1003_g N_VGND_c_392_n 0.0054895f $X=3.825 $Y=0.445 $X2=0 $Y2=0
cc_206 N_TE_B_M1005_g N_VGND_c_393_n 0.00439806f $X=3.465 $Y=0.445 $X2=0 $Y2=0
cc_207 N_TE_B_M1003_g N_VGND_c_393_n 0.00714213f $X=3.825 $Y=0.445 $X2=0 $Y2=0
cc_208 N_VPWR_c_312_n N_Z_M1002_s 0.00231914f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_209 N_VPWR_c_314_n Z 0.0153347f $X=3.105 $Y=1.98 $X2=0 $Y2=0
cc_210 N_VPWR_c_313_n Z 0.0302825f $X=1.51 $Y=2.56 $X2=0 $Y2=0
cc_211 N_VPWR_c_314_n Z 0.0724096f $X=3.105 $Y=1.98 $X2=0 $Y2=0
cc_212 N_VPWR_c_317_n Z 0.0297557f $X=2.94 $Y=3.33 $X2=0 $Y2=0
cc_213 N_VPWR_c_312_n Z 0.0226359f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_214 N_VPWR_c_312_n A_515_367# 0.00421247f $X=4.08 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_215 Z A_515_367# 0.00162456f $X=2.555 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_216 Z A_515_367# 0.00925121f $X=2.555 $Y=2.69 $X2=-0.19 $Y2=-0.245
cc_217 N_Z_M1008_d N_VGND_c_393_n 0.00232737f $X=1.93 $Y=0.235 $X2=0 $Y2=0
cc_218 N_VGND_c_393_n A_308_47# 0.00279972f $X=4.08 $Y=0 $X2=-0.19 $Y2=-0.245
cc_219 N_VGND_c_393_n A_708_47# 0.00306596f $X=4.08 $Y=0 $X2=-0.19 $Y2=-0.245
