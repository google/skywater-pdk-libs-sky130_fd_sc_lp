* File: sky130_fd_sc_lp__a221oi_2.pex.spice
* Created: Fri Aug 28 09:53:25 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A221OI_2%C1 3 7 11 15 17 18 26
r40 25 26 50.241 $w=3.07e-07 $l=3.2e-07 $layer=POLY_cond $X=0.585 $Y=1.375
+ $X2=0.905 $Y2=1.375
r41 24 25 17.2704 $w=3.07e-07 $l=1.1e-07 $layer=POLY_cond $X=0.475 $Y=1.375
+ $X2=0.585 $Y2=1.375
r42 22 24 16.4853 $w=3.07e-07 $l=1.05e-07 $layer=POLY_cond $X=0.37 $Y=1.375
+ $X2=0.475 $Y2=1.375
r43 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.37
+ $Y=1.375 $X2=0.37 $Y2=1.375
r44 18 23 8.79496 $w=3.78e-07 $l=2.9e-07 $layer=LI1_cond $X=0.275 $Y=1.665
+ $X2=0.275 $Y2=1.375
r45 17 23 2.4262 $w=3.78e-07 $l=8e-08 $layer=LI1_cond $X=0.275 $Y=1.295
+ $X2=0.275 $Y2=1.375
r46 13 26 17.2704 $w=3.07e-07 $l=2.13014e-07 $layer=POLY_cond $X=1.015 $Y=1.21
+ $X2=0.905 $Y2=1.375
r47 13 15 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=1.015 $Y=1.21
+ $X2=1.015 $Y2=0.655
r48 9 26 19.5117 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.905 $Y=1.54
+ $X2=0.905 $Y2=1.375
r49 9 11 474.309 $w=1.5e-07 $l=9.25e-07 $layer=POLY_cond $X=0.905 $Y=1.54
+ $X2=0.905 $Y2=2.465
r50 5 25 19.5117 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.585 $Y=1.21
+ $X2=0.585 $Y2=1.375
r51 5 7 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=0.585 $Y=1.21
+ $X2=0.585 $Y2=0.655
r52 1 24 19.5117 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=1.54
+ $X2=0.475 $Y2=1.375
r53 1 3 474.309 $w=1.5e-07 $l=9.25e-07 $layer=POLY_cond $X=0.475 $Y=1.54
+ $X2=0.475 $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__A221OI_2%B2 3 7 11 15 17 20 21 25 26 27 33 50
c83 20 0 1.40934e-19 $X=3.165 $Y=1.46
c84 15 0 1.73857e-19 $X=3.145 $Y=2.465
r85 33 36 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.825 $Y=1.51
+ $X2=1.825 $Y2=1.675
r86 33 35 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.825 $Y=1.51
+ $X2=1.825 $Y2=1.345
r87 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.825
+ $Y=1.51 $X2=1.825 $Y2=1.51
r88 27 50 6.27016 $w=3.58e-07 $l=9.5e-08 $layer=LI1_cond $X=2.16 $Y=1.605
+ $X2=2.255 $Y2=1.605
r89 27 34 6.87953 $w=5.28e-07 $l=2.5e-07 $layer=LI1_cond $X=2.075 $Y=1.605
+ $X2=1.825 $Y2=1.605
r90 26 34 4.64178 $w=3.58e-07 $l=1.45e-07 $layer=LI1_cond $X=1.68 $Y=1.605
+ $X2=1.825 $Y2=1.605
r91 25 26 15.3659 $w=3.58e-07 $l=4.8e-07 $layer=LI1_cond $X=1.2 $Y=1.605
+ $X2=1.68 $Y2=1.605
r92 21 39 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.165 $Y=1.46
+ $X2=3.165 $Y2=1.625
r93 21 38 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.165 $Y=1.46
+ $X2=3.165 $Y2=1.295
r94 20 23 8.3814 $w=3.28e-07 $l=2.4e-07 $layer=LI1_cond $X=3.165 $Y=1.46
+ $X2=3.165 $Y2=1.7
r95 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.165
+ $Y=1.46 $X2=3.165 $Y2=1.46
r96 17 23 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3 $Y=1.7 $X2=3.165
+ $Y2=1.7
r97 17 50 48.6043 $w=1.68e-07 $l=7.45e-07 $layer=LI1_cond $X=3 $Y=1.7 $X2=2.255
+ $Y2=1.7
r98 15 39 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=3.145 $Y=2.465
+ $X2=3.145 $Y2=1.625
r99 11 38 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=3.135 $Y=0.655
+ $X2=3.135 $Y2=1.295
r100 7 36 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.855 $Y=2.465
+ $X2=1.855 $Y2=1.675
r101 3 35 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.845 $Y=0.655
+ $X2=1.845 $Y2=1.345
.ends

.subckt PM_SKY130_FD_SC_LP__A221OI_2%B1 1 3 6 8 10 13 15 22
c52 13 0 1.40934e-19 $X=2.715 $Y=2.465
r53 22 23 1.47853 $w=3.26e-07 $l=1e-08 $layer=POLY_cond $X=2.705 $Y=1.35
+ $X2=2.715 $Y2=1.35
r54 20 22 17.0031 $w=3.26e-07 $l=1.15e-07 $layer=POLY_cond $X=2.59 $Y=1.35
+ $X2=2.705 $Y2=1.35
r55 18 20 45.0951 $w=3.26e-07 $l=3.05e-07 $layer=POLY_cond $X=2.285 $Y=1.35
+ $X2=2.59 $Y2=1.35
r56 17 18 1.47853 $w=3.26e-07 $l=1e-08 $layer=POLY_cond $X=2.275 $Y=1.35
+ $X2=2.285 $Y2=1.35
r57 15 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.59
+ $Y=1.35 $X2=2.59 $Y2=1.35
r58 11 23 20.933 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.715 $Y=1.515
+ $X2=2.715 $Y2=1.35
r59 11 13 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=2.715 $Y=1.515
+ $X2=2.715 $Y2=2.465
r60 8 22 20.933 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.705 $Y=1.185
+ $X2=2.705 $Y2=1.35
r61 8 10 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.705 $Y=1.185
+ $X2=2.705 $Y2=0.655
r62 4 18 20.933 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.285 $Y=1.515
+ $X2=2.285 $Y2=1.35
r63 4 6 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=2.285 $Y=1.515
+ $X2=2.285 $Y2=2.465
r64 1 17 20.933 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.275 $Y=1.185
+ $X2=2.275 $Y2=1.35
r65 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.275 $Y=1.185
+ $X2=2.275 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__A221OI_2%A2 3 7 11 15 18 19 22 23 27 28 33 39
c77 22 0 2.96718e-19 $X=3.705 $Y=1.51
c78 3 0 1.73468e-19 $X=3.615 $Y=2.465
r79 28 39 2.61705 $w=3.4e-07 $l=8.5e-08 $layer=LI1_cond $X=5.505 $Y=1.7
+ $X2=5.505 $Y2=1.615
r80 28 39 0.610117 $w=3.38e-07 $l=1.8e-08 $layer=LI1_cond $X=5.505 $Y=1.597
+ $X2=5.505 $Y2=1.615
r81 27 28 10.2364 $w=3.38e-07 $l=3.02e-07 $layer=LI1_cond $X=5.505 $Y=1.295
+ $X2=5.505 $Y2=1.597
r82 27 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.49
+ $Y=1.375 $X2=5.49 $Y2=1.375
r83 23 38 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.705 $Y=1.51
+ $X2=3.705 $Y2=1.675
r84 23 37 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.705 $Y=1.51
+ $X2=3.705 $Y2=1.345
r85 22 25 8.75857 $w=2.48e-07 $l=1.9e-07 $layer=LI1_cond $X=3.665 $Y=1.51
+ $X2=3.665 $Y2=1.7
r86 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.705
+ $Y=1.51 $X2=3.705 $Y2=1.51
r87 20 25 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.79 $Y=1.7
+ $X2=3.665 $Y2=1.7
r88 19 28 5.2341 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=5.335 $Y=1.7 $X2=5.505
+ $Y2=1.7
r89 19 20 100.797 $w=1.68e-07 $l=1.545e-06 $layer=LI1_cond $X=5.335 $Y=1.7
+ $X2=3.79 $Y2=1.7
r90 17 33 69.9445 $w=3.3e-07 $l=4e-07 $layer=POLY_cond $X=5.09 $Y=1.375 $X2=5.49
+ $Y2=1.375
r91 17 18 5.03009 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=5.09 $Y=1.375
+ $X2=5.015 $Y2=1.375
r92 13 18 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.015 $Y=1.54
+ $X2=5.015 $Y2=1.375
r93 13 15 474.309 $w=1.5e-07 $l=9.25e-07 $layer=POLY_cond $X=5.015 $Y=1.54
+ $X2=5.015 $Y2=2.465
r94 9 18 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.015 $Y=1.21
+ $X2=5.015 $Y2=1.375
r95 9 11 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=5.015 $Y=1.21
+ $X2=5.015 $Y2=0.655
r96 7 37 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.725 $Y=0.655
+ $X2=3.725 $Y2=1.345
r97 3 38 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.615 $Y=2.465
+ $X2=3.615 $Y2=1.675
.ends

.subckt PM_SKY130_FD_SC_LP__A221OI_2%A1 1 3 6 8 10 13 15 16 17 26
c52 6 0 1.22861e-19 $X=4.155 $Y=2.465
r53 24 26 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=4.245 $Y=1.35
+ $X2=4.585 $Y2=1.35
r54 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.245
+ $Y=1.35 $X2=4.245 $Y2=1.35
r55 21 24 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=4.155 $Y=1.35
+ $X2=4.245 $Y2=1.35
r56 16 17 23.5393 $w=2.33e-07 $l=4.8e-07 $layer=LI1_cond $X=4.56 $Y=1.327
+ $X2=5.04 $Y2=1.327
r57 16 25 15.4476 $w=2.33e-07 $l=3.15e-07 $layer=LI1_cond $X=4.56 $Y=1.327
+ $X2=4.245 $Y2=1.327
r58 15 25 8.09162 $w=2.33e-07 $l=1.65e-07 $layer=LI1_cond $X=4.08 $Y=1.327
+ $X2=4.245 $Y2=1.327
r59 11 26 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.585 $Y=1.515
+ $X2=4.585 $Y2=1.35
r60 11 13 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=4.585 $Y=1.515
+ $X2=4.585 $Y2=2.465
r61 8 26 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.585 $Y=1.185
+ $X2=4.585 $Y2=1.35
r62 8 10 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=4.585 $Y=1.185
+ $X2=4.585 $Y2=0.655
r63 4 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.155 $Y=1.515
+ $X2=4.155 $Y2=1.35
r64 4 6 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=4.155 $Y=1.515
+ $X2=4.155 $Y2=2.465
r65 1 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.155 $Y=1.185
+ $X2=4.155 $Y2=1.35
r66 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=4.155 $Y=1.185
+ $X2=4.155 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__A221OI_2%A_27_367# 1 2 3 4 13 15 17 19 20 21 25 36
+ 38
c50 38 0 1.73468e-19 $X=2.93 $Y=2.04
r51 26 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.235 $Y=2.04
+ $X2=2.07 $Y2=2.04
r52 25 38 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.765 $Y=2.04
+ $X2=2.93 $Y2=2.04
r53 25 26 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=2.765 $Y=2.04
+ $X2=2.235 $Y2=2.04
r54 22 32 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.285 $Y=2.04
+ $X2=1.155 $Y2=2.04
r55 21 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.905 $Y=2.04
+ $X2=2.07 $Y2=2.04
r56 21 22 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=1.905 $Y=2.04
+ $X2=1.285 $Y2=2.04
r57 20 34 2.85134 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=1.155 $Y=2.905
+ $X2=1.155 $Y2=2.99
r58 19 32 2.85134 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=1.155 $Y=2.125
+ $X2=1.155 $Y2=2.04
r59 19 20 34.5733 $w=2.58e-07 $l=7.8e-07 $layer=LI1_cond $X=1.155 $Y=2.125
+ $X2=1.155 $Y2=2.905
r60 18 30 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.355 $Y=2.99
+ $X2=0.225 $Y2=2.99
r61 17 34 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.025 $Y=2.99
+ $X2=1.155 $Y2=2.99
r62 17 18 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.025 $Y=2.99
+ $X2=0.355 $Y2=2.99
r63 13 30 2.85134 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=0.225 $Y=2.905
+ $X2=0.225 $Y2=2.99
r64 13 15 36.1247 $w=2.58e-07 $l=8.15e-07 $layer=LI1_cond $X=0.225 $Y=2.905
+ $X2=0.225 $Y2=2.09
r65 4 38 300 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=2 $X=2.79
+ $Y=1.835 $X2=2.93 $Y2=2.04
r66 3 36 300 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=2 $X=1.93
+ $Y=1.835 $X2=2.07 $Y2=2.04
r67 2 34 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=0.98
+ $Y=1.835 $X2=1.12 $Y2=2.91
r68 2 32 400 $w=1.7e-07 $l=3.4803e-07 $layer=licon1_PDIFF $count=1 $X=0.98
+ $Y=1.835 $X2=1.12 $Y2=2.12
r69 1 30 400 $w=1.7e-07 $l=1.13578e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.835 $X2=0.26 $Y2=2.91
r70 1 15 400 $w=1.7e-07 $l=3.11288e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.835 $X2=0.26 $Y2=2.09
.ends

.subckt PM_SKY130_FD_SC_LP__A221OI_2%Y 1 2 3 4 18 19 21 22 23 24 25 26
r55 25 45 2.37473 $w=3.28e-07 $l=6.8e-08 $layer=LI1_cond $X=0.69 $Y=2.017
+ $X2=0.69 $Y2=2.085
r56 25 53 4.67098 $w=3.28e-07 $l=9.7e-08 $layer=LI1_cond $X=0.69 $Y=2.017
+ $X2=0.69 $Y2=1.92
r57 25 26 10.5815 $w=3.28e-07 $l=3.03e-07 $layer=LI1_cond $X=0.69 $Y=2.102
+ $X2=0.69 $Y2=2.405
r58 25 45 0.593683 $w=3.28e-07 $l=1.7e-08 $layer=LI1_cond $X=0.69 $Y=2.102
+ $X2=0.69 $Y2=2.085
r59 24 53 13.3579 $w=2.18e-07 $l=2.55e-07 $layer=LI1_cond $X=0.745 $Y=1.665
+ $X2=0.745 $Y2=1.92
r60 23 24 19.382 $w=2.18e-07 $l=3.7e-07 $layer=LI1_cond $X=0.745 $Y=1.295
+ $X2=0.745 $Y2=1.665
r61 23 39 13.3579 $w=2.18e-07 $l=2.55e-07 $layer=LI1_cond $X=0.745 $Y=1.295
+ $X2=0.745 $Y2=1.04
r62 22 34 5.43174 $w=2.4e-07 $l=1.27e-07 $layer=LI1_cond $X=0.765 $Y=0.912
+ $X2=0.765 $Y2=0.785
r63 22 39 5.43174 $w=2.4e-07 $l=1.37637e-07 $layer=LI1_cond $X=0.765 $Y=0.912
+ $X2=0.745 $Y2=1.04
r64 21 34 13.0758 $w=2.58e-07 $l=2.95e-07 $layer=LI1_cond $X=0.765 $Y=0.49
+ $X2=0.765 $Y2=0.785
r65 18 19 6.2579 $w=3.73e-07 $l=1.65e-07 $layer=LI1_cond $X=4.37 $Y=0.852
+ $X2=4.205 $Y2=0.852
r66 16 19 77.5074 $w=2.53e-07 $l=1.715e-06 $layer=LI1_cond $X=2.49 $Y=0.912
+ $X2=4.205 $Y2=0.912
r67 14 22 1.12519 $w=2.55e-07 $l=1.3e-07 $layer=LI1_cond $X=0.895 $Y=0.912
+ $X2=0.765 $Y2=0.912
r68 14 16 72.0842 $w=2.53e-07 $l=1.595e-06 $layer=LI1_cond $X=0.895 $Y=0.912
+ $X2=2.49 $Y2=0.912
r69 4 25 300 $w=1.7e-07 $l=2.504e-07 $layer=licon1_PDIFF $count=2 $X=0.55
+ $Y=1.835 $X2=0.69 $Y2=2.025
r70 3 18 182 $w=1.7e-07 $l=6.61306e-07 $layer=licon1_NDIFF $count=1 $X=4.23
+ $Y=0.235 $X2=4.37 $Y2=0.83
r71 2 16 182 $w=1.7e-07 $l=7.21613e-07 $layer=licon1_NDIFF $count=1 $X=2.35
+ $Y=0.235 $X2=2.49 $Y2=0.89
r72 1 21 91 $w=1.7e-07 $l=3.17372e-07 $layer=licon1_NDIFF $count=2 $X=0.66
+ $Y=0.235 $X2=0.8 $Y2=0.49
.ends

.subckt PM_SKY130_FD_SC_LP__A221OI_2%A_303_367# 1 2 3 4 5 18 20 21 24 26 28 29
+ 30 34 36 38 40 42 48
r62 38 50 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.27 $Y=2.125
+ $X2=5.27 $Y2=2.04
r63 38 40 16.3647 $w=2.48e-07 $l=3.55e-07 $layer=LI1_cond $X=5.27 $Y=2.125
+ $X2=5.27 $Y2=2.48
r64 37 48 6.70225 $w=1.7e-07 $l=1.18e-07 $layer=LI1_cond $X=4.455 $Y=2.04
+ $X2=4.337 $Y2=2.04
r65 36 50 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.145 $Y=2.04
+ $X2=5.27 $Y2=2.04
r66 36 37 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=5.145 $Y=2.04
+ $X2=4.455 $Y2=2.04
r67 32 48 0.207053 $w=2.35e-07 $l=8.5e-08 $layer=LI1_cond $X=4.337 $Y=2.125
+ $X2=4.337 $Y2=2.04
r68 32 34 17.4092 $w=2.33e-07 $l=3.55e-07 $layer=LI1_cond $X=4.337 $Y=2.125
+ $X2=4.337 $Y2=2.48
r69 31 44 4.64039 $w=1.7e-07 $l=1.43e-07 $layer=LI1_cond $X=3.55 $Y=2.04
+ $X2=3.407 $Y2=2.04
r70 30 48 6.70225 $w=1.7e-07 $l=1.17e-07 $layer=LI1_cond $X=4.22 $Y=2.04
+ $X2=4.337 $Y2=2.04
r71 30 31 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.22 $Y=2.04
+ $X2=3.55 $Y2=2.04
r72 29 46 2.77043 $w=2.85e-07 $l=8.5e-08 $layer=LI1_cond $X=3.407 $Y=2.905
+ $X2=3.407 $Y2=2.99
r73 28 44 2.75828 $w=2.85e-07 $l=8.5e-08 $layer=LI1_cond $X=3.407 $Y=2.125
+ $X2=3.407 $Y2=2.04
r74 28 29 31.5405 $w=2.83e-07 $l=7.8e-07 $layer=LI1_cond $X=3.407 $Y=2.125
+ $X2=3.407 $Y2=2.905
r75 27 42 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.595 $Y=2.99 $X2=2.5
+ $Y2=2.99
r76 26 46 4.62824 $w=1.7e-07 $l=1.42e-07 $layer=LI1_cond $X=3.265 $Y=2.99
+ $X2=3.407 $Y2=2.99
r77 26 27 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.265 $Y=2.99
+ $X2=2.595 $Y2=2.99
r78 22 42 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=2.5 $Y=2.905 $X2=2.5
+ $Y2=2.99
r79 22 24 25.9761 $w=1.88e-07 $l=4.45e-07 $layer=LI1_cond $X=2.5 $Y=2.905
+ $X2=2.5 $Y2=2.46
r80 20 42 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.405 $Y=2.99 $X2=2.5
+ $Y2=2.99
r81 20 21 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.405 $Y=2.99
+ $X2=1.735 $Y2=2.99
r82 16 21 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=1.605 $Y=2.905
+ $X2=1.735 $Y2=2.99
r83 16 18 19.7245 $w=2.58e-07 $l=4.45e-07 $layer=LI1_cond $X=1.605 $Y=2.905
+ $X2=1.605 $Y2=2.46
r84 5 50 600 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=1 $X=5.09
+ $Y=1.835 $X2=5.23 $Y2=2.04
r85 5 40 300 $w=1.7e-07 $l=7.11565e-07 $layer=licon1_PDIFF $count=2 $X=5.09
+ $Y=1.835 $X2=5.23 $Y2=2.48
r86 4 48 600 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_PDIFF $count=1 $X=4.23
+ $Y=1.835 $X2=4.37 $Y2=2.04
r87 4 34 300 $w=1.7e-07 $l=7.11565e-07 $layer=licon1_PDIFF $count=2 $X=4.23
+ $Y=1.835 $X2=4.37 $Y2=2.48
r88 3 46 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=3.22
+ $Y=1.835 $X2=3.36 $Y2=2.91
r89 3 44 400 $w=1.7e-07 $l=3.4803e-07 $layer=licon1_PDIFF $count=1 $X=3.22
+ $Y=1.835 $X2=3.36 $Y2=2.12
r90 2 24 300 $w=1.7e-07 $l=6.91466e-07 $layer=licon1_PDIFF $count=2 $X=2.36
+ $Y=1.835 $X2=2.5 $Y2=2.46
r91 1 18 300 $w=1.7e-07 $l=6.84653e-07 $layer=licon1_PDIFF $count=2 $X=1.515
+ $Y=1.835 $X2=1.64 $Y2=2.46
.ends

.subckt PM_SKY130_FD_SC_LP__A221OI_2%VPWR 1 2 9 13 16 17 19 20 21 34 35
r68 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r69 32 35 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.52 $Y2=3.33
r70 31 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r71 29 32 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.56 $Y2=3.33
r72 28 29 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r73 24 28 219.209 $w=1.68e-07 $l=3.36e-06 $layer=LI1_cond $X=0.24 $Y=3.33
+ $X2=3.6 $Y2=3.33
r74 24 25 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r75 21 29 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.88 $Y=3.33
+ $X2=3.6 $Y2=3.33
r76 21 25 0.73586 $w=4.9e-07 $l=2.64e-06 $layer=MET1_cond $X=2.88 $Y=3.33
+ $X2=0.24 $Y2=3.33
r77 19 31 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=4.635 $Y=3.33
+ $X2=4.56 $Y2=3.33
r78 19 20 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.635 $Y=3.33
+ $X2=4.8 $Y2=3.33
r79 18 34 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=4.965 $Y=3.33
+ $X2=5.52 $Y2=3.33
r80 18 20 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.965 $Y=3.33
+ $X2=4.8 $Y2=3.33
r81 16 28 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=3.72 $Y=3.33 $X2=3.6
+ $Y2=3.33
r82 16 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.72 $Y=3.33
+ $X2=3.885 $Y2=3.33
r83 15 31 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=4.05 $Y=3.33
+ $X2=4.56 $Y2=3.33
r84 15 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.05 $Y=3.33
+ $X2=3.885 $Y2=3.33
r85 11 20 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.8 $Y=3.245 $X2=4.8
+ $Y2=3.33
r86 11 13 29.5095 $w=3.28e-07 $l=8.45e-07 $layer=LI1_cond $X=4.8 $Y=3.245
+ $X2=4.8 $Y2=2.4
r87 7 17 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.885 $Y=3.245
+ $X2=3.885 $Y2=3.33
r88 7 9 29.5095 $w=3.28e-07 $l=8.45e-07 $layer=LI1_cond $X=3.885 $Y=3.245
+ $X2=3.885 $Y2=2.4
r89 2 13 300 $w=1.7e-07 $l=6.3113e-07 $layer=licon1_PDIFF $count=2 $X=4.66
+ $Y=1.835 $X2=4.8 $Y2=2.4
r90 1 9 300 $w=1.7e-07 $l=6.55286e-07 $layer=licon1_PDIFF $count=2 $X=3.69
+ $Y=1.835 $X2=3.885 $Y2=2.4
.ends

.subckt PM_SKY130_FD_SC_LP__A221OI_2%VGND 1 2 3 4 13 15 19 23 26 27 29 30 31 52
+ 53 61 67
r67 65 67 9.60904 $w=6.98e-07 $l=9.5e-08 $layer=LI1_cond $X=1.68 $Y=0.265
+ $X2=1.775 $Y2=0.265
r68 65 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r69 63 65 1.19608 $w=6.98e-07 $l=7e-08 $layer=LI1_cond $X=1.61 $Y=0.265 $X2=1.68
+ $Y2=0.265
r70 60 66 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r71 59 63 7.0056 $w=6.98e-07 $l=4.1e-07 $layer=LI1_cond $X=1.2 $Y=0.265 $X2=1.61
+ $Y2=0.265
r72 59 61 10.2925 $w=6.98e-07 $l=1.35e-07 $layer=LI1_cond $X=1.2 $Y=0.265
+ $X2=1.065 $Y2=0.265
r73 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r74 56 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r75 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r76 50 53 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=5.52
+ $Y2=0
r77 49 50 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r78 47 50 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=3.6 $Y=0 $X2=5.04
+ $Y2=0
r79 46 49 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=3.6 $Y=0 $X2=5.04
+ $Y2=0
r80 46 47 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r81 44 47 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r82 43 44 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r83 41 66 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.68
+ $Y2=0
r84 40 43 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r85 40 67 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=2.16 $Y=0 $X2=1.775
+ $Y2=0
r86 40 41 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r87 37 60 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r88 37 57 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r89 36 61 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.72 $Y=0 $X2=1.065
+ $Y2=0
r90 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r91 34 56 3.99156 $w=1.7e-07 $l=2.33e-07 $layer=LI1_cond $X=0.465 $Y=0 $X2=0.232
+ $Y2=0
r92 34 36 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.465 $Y=0 $X2=0.72
+ $Y2=0
r93 31 44 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.88 $Y=0 $X2=3.12
+ $Y2=0
r94 31 41 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.88 $Y=0 $X2=2.16
+ $Y2=0
r95 29 49 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=5.135 $Y=0 $X2=5.04
+ $Y2=0
r96 29 30 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=5.135 $Y=0 $X2=5.265
+ $Y2=0
r97 28 52 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=5.395 $Y=0 $X2=5.52
+ $Y2=0
r98 28 30 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=5.395 $Y=0 $X2=5.265
+ $Y2=0
r99 26 43 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=3.26 $Y=0 $X2=3.12
+ $Y2=0
r100 26 27 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.26 $Y=0 $X2=3.425
+ $Y2=0
r101 25 46 0.652406 $w=1.68e-07 $l=1e-08 $layer=LI1_cond $X=3.59 $Y=0 $X2=3.6
+ $Y2=0
r102 25 27 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.59 $Y=0 $X2=3.425
+ $Y2=0
r103 21 30 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=5.265 $Y=0.085
+ $X2=5.265 $Y2=0
r104 21 23 13.0758 $w=2.58e-07 $l=2.95e-07 $layer=LI1_cond $X=5.265 $Y=0.085
+ $X2=5.265 $Y2=0.38
r105 17 27 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.425 $Y=0.085
+ $X2=3.425 $Y2=0
r106 17 19 13.7944 $w=3.28e-07 $l=3.95e-07 $layer=LI1_cond $X=3.425 $Y=0.085
+ $X2=3.425 $Y2=0.48
r107 13 56 3.22066 $w=2.6e-07 $l=1.39155e-07 $layer=LI1_cond $X=0.335 $Y=0.085
+ $X2=0.232 $Y2=0
r108 13 15 13.0758 $w=2.58e-07 $l=2.95e-07 $layer=LI1_cond $X=0.335 $Y=0.085
+ $X2=0.335 $Y2=0.38
r109 4 23 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.09
+ $Y=0.235 $X2=5.23 $Y2=0.38
r110 3 19 182 $w=1.7e-07 $l=3.35708e-07 $layer=licon1_NDIFF $count=1 $X=3.21
+ $Y=0.235 $X2=3.425 $Y2=0.48
r111 2 63 91 $w=1.7e-07 $l=6.34823e-07 $layer=licon1_NDIFF $count=2 $X=1.09
+ $Y=0.235 $X2=1.61 $Y2=0.49
r112 1 15 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.245
+ $Y=0.235 $X2=0.37 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_LP__A221OI_2%A_384_47# 1 2 11
r11 8 11 30.0334 $w=3.28e-07 $l=8.6e-07 $layer=LI1_cond $X=2.06 $Y=0.45 $X2=2.92
+ $Y2=0.45
r12 2 11 182 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_NDIFF $count=1 $X=2.78
+ $Y=0.235 $X2=2.92 $Y2=0.45
r13 1 8 182 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_NDIFF $count=1 $X=1.92
+ $Y=0.235 $X2=2.06 $Y2=0.45
.ends

.subckt PM_SKY130_FD_SC_LP__A221OI_2%A_760_47# 1 2 7 14
r18 7 14 4.18573 $w=2.3e-07 $l=1.65e-07 $layer=LI1_cond $X=4.635 $Y=0.37 $X2=4.8
+ $Y2=0.37
r19 7 9 34.8238 $w=2.28e-07 $l=6.95e-07 $layer=LI1_cond $X=4.635 $Y=0.37
+ $X2=3.94 $Y2=0.37
r20 2 14 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=4.66
+ $Y=0.235 $X2=4.8 $Y2=0.38
r21 1 9 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=3.8
+ $Y=0.235 $X2=3.94 $Y2=0.38
.ends

