* File: sky130_fd_sc_lp__a311o_2.spice
* Created: Fri Aug 28 09:57:38 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__a311o_2.pex.spice"
.subckt sky130_fd_sc_lp__a311o_2  VNB VPB A3 A2 A1 B1 C1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* C1	C1
* B1	B1
* A1	A1
* A2	A2
* A3	A3
* VPB	VPB
* VNB	VNB
MM1012 N_VGND_M1012_d N_A_85_21#_M1012_g N_X_M1012_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2394 AS=0.1176 PD=2.25 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75003.4 A=0.126 P=1.98 MULT=1
MM1013 N_VGND_M1013_d N_A_85_21#_M1013_g N_X_M1012_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2604 AS=0.1176 PD=1.46 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75002.9 A=0.126 P=1.98 MULT=1
MM1010 A_355_47# N_A3_M1010_g N_VGND_M1013_d VNB NSHORT L=0.15 W=0.84 AD=0.0882
+ AS=0.2604 PD=1.05 PS=1.46 NRD=7.14 NRS=0 M=1 R=5.6 SA=75001.4 SB=75002.2
+ A=0.126 P=1.98 MULT=1
MM1006 A_427_47# N_A2_M1006_g A_355_47# VNB NSHORT L=0.15 W=0.84 AD=0.1638
+ AS=0.0882 PD=1.23 PS=1.05 NRD=19.992 NRS=7.14 M=1 R=5.6 SA=75001.8 SB=75001.8
+ A=0.126 P=1.98 MULT=1
MM1000 N_A_85_21#_M1000_d N_A1_M1000_g A_427_47# VNB NSHORT L=0.15 W=0.84
+ AD=0.1638 AS=0.1638 PD=1.23 PS=1.23 NRD=7.848 NRS=19.992 M=1 R=5.6 SA=75002.3
+ SB=75001.3 A=0.126 P=1.98 MULT=1
MM1003 N_VGND_M1003_d N_B1_M1003_g N_A_85_21#_M1000_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1638 AS=0.1638 PD=1.23 PS=1.23 NRD=8.568 NRS=7.848 M=1 R=5.6 SA=75002.8
+ SB=75000.7 A=0.126 P=1.98 MULT=1
MM1008 N_A_85_21#_M1008_d N_C1_M1008_g N_VGND_M1003_d VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1638 PD=2.21 PS=1.23 NRD=0 NRS=7.14 M=1 R=5.6 SA=75003.4
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1001 N_X_M1001_d N_A_85_21#_M1001_g N_VPWR_M1001_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75003.3 A=0.189 P=2.82 MULT=1
MM1004 N_X_M1001_d N_A_85_21#_M1004_g N_VPWR_M1004_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.29925 PD=1.54 PS=1.735 NRD=0 NRS=14.8341 M=1 R=8.4 SA=75000.6
+ SB=75002.9 A=0.189 P=2.82 MULT=1
MM1005 N_A_341_367#_M1005_d N_A3_M1005_g N_VPWR_M1004_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.29925 PD=1.54 PS=1.735 NRD=0 NRS=15.6221 M=1 R=8.4
+ SA=75001.2 SB=75002.2 A=0.189 P=2.82 MULT=1
MM1009 N_VPWR_M1009_d N_A2_M1009_g N_A_341_367#_M1005_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3591 AS=0.1764 PD=1.83 PS=1.54 NRD=23.443 NRS=0 M=1 R=8.4
+ SA=75001.7 SB=75001.8 A=0.189 P=2.82 MULT=1
MM1011 N_A_341_367#_M1011_d N_A1_M1011_g N_VPWR_M1009_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.3591 PD=1.54 PS=1.83 NRD=0 NRS=21.8867 M=1 R=8.4
+ SA=75002.4 SB=75001.1 A=0.189 P=2.82 MULT=1
MM1007 A_657_367# N_B1_M1007_g N_A_341_367#_M1011_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.2016 AS=0.1764 PD=1.58 PS=1.54 NRD=16.4101 NRS=0 M=1 R=8.4 SA=75002.8
+ SB=75000.7 A=0.189 P=2.82 MULT=1
MM1002 N_A_85_21#_M1002_d N_C1_M1002_g A_657_367# VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.2016 PD=3.05 PS=1.58 NRD=0 NRS=16.4101 M=1 R=8.4 SA=75003.3
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX14_noxref VNB VPB NWDIODE A=8.7655 P=13.13
*
.include "sky130_fd_sc_lp__a311o_2.pxi.spice"
*
.ends
*
*
