# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__o31ai_0
  CLASS CORE ;
  FOREIGN sky130_fd_sc_lp__o31ai_0 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.880000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.840000 0.410000 2.225000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.580000 1.130000 1.005000 2.225000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.360000 1.105000 1.895000 1.810000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.065000 0.840000 2.255000 1.810000 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  0.433300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.485000 1.980000 2.790000 2.225000 ;
        RECT 1.485000 2.225000 1.815000 3.065000 ;
        RECT 2.065000 0.340000 2.790000 0.670000 ;
        RECT 2.425000 0.670000 2.790000 1.980000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 2.880000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 2.880000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.880000 0.085000 ;
      RECT 0.000000  3.245000 2.880000 3.415000 ;
      RECT 0.235000  0.085000 0.565000 0.670000 ;
      RECT 0.275000  2.395000 0.605000 3.245000 ;
      RECT 0.735000  0.370000 0.975000 0.765000 ;
      RECT 0.735000  0.765000 1.895000 0.935000 ;
      RECT 1.145000  0.085000 1.475000 0.595000 ;
      RECT 1.645000  0.370000 1.895000 0.765000 ;
      RECT 1.985000  2.395000 2.245000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
  END
END sky130_fd_sc_lp__o31ai_0
END LIBRARY
