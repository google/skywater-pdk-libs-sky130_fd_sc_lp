* File: sky130_fd_sc_lp__sdlclkp_lp.pxi.spice
* Created: Fri Aug 28 11:31:46 2020
* 
x_PM_SKY130_FD_SC_LP__SDLCLKP_LP%GATE N_GATE_c_165_n N_GATE_M1011_g
+ N_GATE_M1018_g N_GATE_c_166_n N_GATE_M1027_g GATE N_GATE_c_167_n
+ N_GATE_c_168_n PM_SKY130_FD_SC_LP__SDLCLKP_LP%GATE
x_PM_SKY130_FD_SC_LP__SDLCLKP_LP%SCE N_SCE_c_199_n N_SCE_M1019_g N_SCE_M1000_g
+ N_SCE_c_200_n N_SCE_c_201_n N_SCE_M1023_g N_SCE_c_202_n SCE SCE N_SCE_c_203_n
+ N_SCE_c_204_n N_SCE_c_205_n PM_SKY130_FD_SC_LP__SDLCLKP_LP%SCE
x_PM_SKY130_FD_SC_LP__SDLCLKP_LP%A_356_278# N_A_356_278#_M1017_s
+ N_A_356_278#_M1007_s N_A_356_278#_M1006_g N_A_356_278#_c_255_n
+ N_A_356_278#_M1015_g N_A_356_278#_c_256_n N_A_356_278#_c_257_n
+ N_A_356_278#_c_258_n N_A_356_278#_M1009_g N_A_356_278#_c_259_n
+ N_A_356_278#_c_260_n N_A_356_278#_c_261_n N_A_356_278#_M1013_g
+ N_A_356_278#_M1021_g N_A_356_278#_c_262_n N_A_356_278#_c_263_n
+ N_A_356_278#_c_264_n N_A_356_278#_c_265_n N_A_356_278#_c_293_p
+ N_A_356_278#_c_290_n N_A_356_278#_c_275_n N_A_356_278#_c_266_n
+ N_A_356_278#_c_277_n N_A_356_278#_c_295_p N_A_356_278#_c_267_n
+ N_A_356_278#_c_268_n N_A_356_278#_c_269_n N_A_356_278#_c_279_n
+ N_A_356_278#_c_270_n N_A_356_278#_c_271_n
+ PM_SKY130_FD_SC_LP__SDLCLKP_LP%A_356_278#
x_PM_SKY130_FD_SC_LP__SDLCLKP_LP%A_447_376# N_A_447_376#_M1009_d
+ N_A_447_376#_M1006_d N_A_447_376#_c_435_n N_A_447_376#_M1002_g
+ N_A_447_376#_c_436_n N_A_447_376#_M1026_g N_A_447_376#_c_438_n
+ N_A_447_376#_c_445_n N_A_447_376#_c_439_n N_A_447_376#_c_440_n
+ N_A_447_376#_c_441_n PM_SKY130_FD_SC_LP__SDLCLKP_LP%A_447_376#
x_PM_SKY130_FD_SC_LP__SDLCLKP_LP%A_860_21# N_A_860_21#_M1004_d
+ N_A_860_21#_M1003_d N_A_860_21#_M1024_g N_A_860_21#_M1008_g
+ N_A_860_21#_c_512_n N_A_860_21#_M1001_g N_A_860_21#_M1010_g
+ N_A_860_21#_c_514_n N_A_860_21#_c_526_n N_A_860_21#_c_515_n
+ N_A_860_21#_c_562_p N_A_860_21#_c_546_n N_A_860_21#_c_528_n
+ N_A_860_21#_c_516_n N_A_860_21#_c_517_n N_A_860_21#_c_529_n
+ N_A_860_21#_c_584_p N_A_860_21#_c_518_n N_A_860_21#_c_531_n
+ N_A_860_21#_c_532_n N_A_860_21#_c_519_n N_A_860_21#_c_520_n
+ N_A_860_21#_c_577_p N_A_860_21#_c_521_n N_A_860_21#_c_522_n
+ N_A_860_21#_c_523_n PM_SKY130_FD_SC_LP__SDLCLKP_LP%A_860_21#
x_PM_SKY130_FD_SC_LP__SDLCLKP_LP%A_698_405# N_A_698_405#_M1013_d
+ N_A_698_405#_M1002_d N_A_698_405#_M1003_g N_A_698_405#_c_679_n
+ N_A_698_405#_M1014_g N_A_698_405#_c_680_n N_A_698_405#_M1004_g
+ N_A_698_405#_c_681_n N_A_698_405#_c_682_n N_A_698_405#_c_683_n
+ N_A_698_405#_c_689_n N_A_698_405#_c_684_n N_A_698_405#_c_685_n
+ N_A_698_405#_c_686_n PM_SKY130_FD_SC_LP__SDLCLKP_LP%A_698_405#
x_PM_SKY130_FD_SC_LP__SDLCLKP_LP%CLK N_CLK_c_760_n N_CLK_c_761_n N_CLK_M1017_g
+ N_CLK_M1007_g N_CLK_c_763_n N_CLK_M1012_g N_CLK_c_764_n N_CLK_M1025_g
+ N_CLK_c_766_n N_CLK_M1016_g CLK CLK N_CLK_c_768_n
+ PM_SKY130_FD_SC_LP__SDLCLKP_LP%CLK
x_PM_SKY130_FD_SC_LP__SDLCLKP_LP%A_1384_416# N_A_1384_416#_M1001_d
+ N_A_1384_416#_M1025_d N_A_1384_416#_c_832_n N_A_1384_416#_M1020_g
+ N_A_1384_416#_c_840_n N_A_1384_416#_M1022_g N_A_1384_416#_c_833_n
+ N_A_1384_416#_M1005_g N_A_1384_416#_c_841_n N_A_1384_416#_c_842_n
+ N_A_1384_416#_c_834_n N_A_1384_416#_c_835_n N_A_1384_416#_c_836_n
+ N_A_1384_416#_c_837_n N_A_1384_416#_c_845_n N_A_1384_416#_c_838_n
+ N_A_1384_416#_c_839_n PM_SKY130_FD_SC_LP__SDLCLKP_LP%A_1384_416#
x_PM_SKY130_FD_SC_LP__SDLCLKP_LP%A_93_376# N_A_93_376#_M1027_d
+ N_A_93_376#_M1013_s N_A_93_376#_M1018_s N_A_93_376#_M1002_s
+ N_A_93_376#_c_916_n N_A_93_376#_c_909_n N_A_93_376#_c_924_n
+ N_A_93_376#_c_910_n N_A_93_376#_c_917_n N_A_93_376#_c_911_n
+ N_A_93_376#_c_912_n N_A_93_376#_c_913_n N_A_93_376#_c_918_n
+ N_A_93_376#_c_919_n N_A_93_376#_c_914_n N_A_93_376#_c_920_n
+ N_A_93_376#_c_915_n PM_SKY130_FD_SC_LP__SDLCLKP_LP%A_93_376#
x_PM_SKY130_FD_SC_LP__SDLCLKP_LP%VPWR N_VPWR_M1000_d N_VPWR_M1008_d
+ N_VPWR_M1007_d N_VPWR_M1010_d N_VPWR_c_1021_n N_VPWR_c_1022_n N_VPWR_c_1023_n
+ N_VPWR_c_1024_n N_VPWR_c_1025_n VPWR N_VPWR_c_1026_n N_VPWR_c_1027_n
+ N_VPWR_c_1028_n N_VPWR_c_1029_n N_VPWR_c_1020_n N_VPWR_c_1031_n
+ N_VPWR_c_1032_n N_VPWR_c_1033_n PM_SKY130_FD_SC_LP__SDLCLKP_LP%VPWR
x_PM_SKY130_FD_SC_LP__SDLCLKP_LP%GCLK N_GCLK_M1005_d N_GCLK_M1022_d GCLK GCLK
+ GCLK GCLK GCLK GCLK GCLK PM_SKY130_FD_SC_LP__SDLCLKP_LP%GCLK
x_PM_SKY130_FD_SC_LP__SDLCLKP_LP%VGND N_VGND_M1011_s N_VGND_M1023_d
+ N_VGND_M1024_d N_VGND_M1012_d N_VGND_M1020_s N_VGND_c_1139_n N_VGND_c_1140_n
+ N_VGND_c_1141_n N_VGND_c_1142_n N_VGND_c_1143_n N_VGND_c_1144_n
+ N_VGND_c_1145_n N_VGND_c_1146_n N_VGND_c_1147_n N_VGND_c_1148_n VGND
+ N_VGND_c_1149_n N_VGND_c_1150_n N_VGND_c_1151_n N_VGND_c_1152_n
+ N_VGND_c_1153_n N_VGND_c_1154_n PM_SKY130_FD_SC_LP__SDLCLKP_LP%VGND
cc_1 VNB N_GATE_c_165_n 0.020605f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.035
cc_2 VNB N_GATE_c_166_n 0.0150226f $X=-0.19 $Y=-0.245 $X2=0.885 $Y2=1.035
cc_3 VNB N_GATE_c_167_n 0.0247996f $X=-0.19 $Y=-0.245 $X2=0.39 $Y2=1.2
cc_4 VNB N_GATE_c_168_n 0.0878873f $X=-0.19 $Y=-0.245 $X2=0.875 $Y2=1.37
cc_5 VNB N_SCE_c_199_n 0.0137712f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.035
cc_6 VNB N_SCE_c_200_n 0.0165134f $X=-0.19 $Y=-0.245 $X2=0.885 $Y2=0.715
cc_7 VNB N_SCE_c_201_n 0.0135526f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_SCE_c_202_n 0.0043185f $X=-0.19 $Y=-0.245 $X2=0.39 $Y2=1.2
cc_9 VNB N_SCE_c_203_n 0.018815f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_SCE_c_204_n 0.00422896f $X=-0.19 $Y=-0.245 $X2=0.39 $Y2=1.37
cc_11 VNB N_SCE_c_205_n 0.0144257f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_356_278#_c_255_n 0.0135105f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_13 VNB N_A_356_278#_c_256_n 0.0177091f $X=-0.19 $Y=-0.245 $X2=0.39 $Y2=1.2
cc_14 VNB N_A_356_278#_c_257_n 0.00915008f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.37
cc_15 VNB N_A_356_278#_c_258_n 0.0150665f $X=-0.19 $Y=-0.245 $X2=0.885 $Y2=1.37
cc_16 VNB N_A_356_278#_c_259_n 0.0228867f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_356_278#_c_260_n 0.0269792f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_356_278#_c_261_n 0.0189567f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_356_278#_c_262_n 0.00465991f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_356_278#_c_263_n 0.00651024f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_356_278#_c_264_n 0.0250447f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_356_278#_c_265_n 0.00238432f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_356_278#_c_266_n 0.00795058f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_356_278#_c_267_n 0.00964304f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_356_278#_c_268_n 0.0333011f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_356_278#_c_269_n 0.00912181f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_356_278#_c_270_n 0.00570896f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_356_278#_c_271_n 0.0292961f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_447_376#_c_435_n 0.0299612f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_447_376#_c_436_n 0.0349448f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_31 VNB N_A_447_376#_M1026_g 0.0335594f $X=-0.19 $Y=-0.245 $X2=0.39 $Y2=1.2
cc_32 VNB N_A_447_376#_c_438_n 0.0196612f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.37
cc_33 VNB N_A_447_376#_c_439_n 0.00694158f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_447_376#_c_440_n 0.00874739f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_447_376#_c_441_n 0.00640987f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_860_21#_M1024_g 0.0610837f $X=-0.19 $Y=-0.245 $X2=0.885 $Y2=0.715
cc_37 VNB N_A_860_21#_c_512_n 0.0156717f $X=-0.19 $Y=-0.245 $X2=0.39 $Y2=1.2
cc_38 VNB N_A_860_21#_M1010_g 0.0079442f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_860_21#_c_514_n 0.00959351f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_860_21#_c_515_n 0.009395f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_860_21#_c_516_n 0.0182379f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_860_21#_c_517_n 0.00830358f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_860_21#_c_518_n 0.00114126f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_860_21#_c_519_n 0.0144277f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_860_21#_c_520_n 0.00116734f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_860_21#_c_521_n 0.00389184f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_860_21#_c_522_n 0.0305539f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_860_21#_c_523_n 0.0252788f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_698_405#_M1003_g 0.0302314f $X=-0.19 $Y=-0.245 $X2=0.885 $Y2=0.715
cc_50 VNB N_A_698_405#_c_679_n 0.0158652f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_51 VNB N_A_698_405#_c_680_n 0.0188781f $X=-0.19 $Y=-0.245 $X2=0.39 $Y2=1.2
cc_52 VNB N_A_698_405#_c_681_n 0.00523556f $X=-0.19 $Y=-0.245 $X2=0.885 $Y2=1.37
cc_53 VNB N_A_698_405#_c_682_n 0.00258484f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_698_405#_c_683_n 0.00732276f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_698_405#_c_684_n 0.00380776f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_698_405#_c_685_n 0.0611942f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_698_405#_c_686_n 0.0240846f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_CLK_c_760_n 0.0286762f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.035
cc_59 VNB N_CLK_c_761_n 0.0167906f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=0.715
cc_60 VNB N_CLK_M1007_g 0.00216806f $X=-0.19 $Y=-0.245 $X2=0.885 $Y2=1.035
cc_61 VNB N_CLK_c_763_n 0.0149407f $X=-0.19 $Y=-0.245 $X2=0.885 $Y2=0.715
cc_62 VNB N_CLK_c_764_n 0.0369541f $X=-0.19 $Y=-0.245 $X2=0.39 $Y2=1.37
cc_63 VNB N_CLK_M1025_g 0.00719531f $X=-0.19 $Y=-0.245 $X2=0.39 $Y2=1.2
cc_64 VNB N_CLK_c_766_n 0.0157525f $X=-0.19 $Y=-0.245 $X2=0.875 $Y2=1.37
cc_65 VNB CLK 0.00185325f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_CLK_c_768_n 0.0158315f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_A_1384_416#_c_832_n 0.0173651f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_A_1384_416#_c_833_n 0.0168121f $X=-0.19 $Y=-0.245 $X2=0.39 $Y2=1.37
cc_69 VNB N_A_1384_416#_c_834_n 0.0320132f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.37
cc_70 VNB N_A_1384_416#_c_835_n 0.00141796f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_A_1384_416#_c_836_n 0.00327253f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_A_1384_416#_c_837_n 0.00249621f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_A_1384_416#_c_838_n 0.00277722f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_A_1384_416#_c_839_n 0.081715f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_A_93_376#_c_909_n 0.00514557f $X=-0.19 $Y=-0.245 $X2=0.875 $Y2=1.37
cc_76 VNB N_A_93_376#_c_910_n 0.0171742f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_A_93_376#_c_911_n 0.00107242f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_A_93_376#_c_912_n 0.016101f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_A_93_376#_c_913_n 0.00267405f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_A_93_376#_c_914_n 0.00497436f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_A_93_376#_c_915_n 0.00697642f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_VPWR_c_1020_n 0.362705f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB GCLK 0.0639155f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_VGND_c_1139_n 0.0122168f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.37
cc_85 VNB N_VGND_c_1140_n 0.0351245f $X=-0.19 $Y=-0.245 $X2=0.885 $Y2=1.37
cc_86 VNB N_VGND_c_1141_n 0.0120462f $X=-0.19 $Y=-0.245 $X2=0.39 $Y2=1.37
cc_87 VNB N_VGND_c_1142_n 0.00619667f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_VGND_c_1143_n 0.0387534f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_VGND_c_1144_n 0.0110853f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_VGND_c_1145_n 0.0375052f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_VGND_c_1146_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_VGND_c_1147_n 0.0515662f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_93 VNB N_VGND_c_1148_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_94 VNB N_VGND_c_1149_n 0.0603227f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_95 VNB N_VGND_c_1150_n 0.0136198f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_96 VNB N_VGND_c_1151_n 0.0303284f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_97 VNB N_VGND_c_1152_n 0.47501f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_98 VNB N_VGND_c_1153_n 0.00513431f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_99 VNB N_VGND_c_1154_n 0.00528688f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_100 VPB N_GATE_M1018_g 0.031197f $X=-0.19 $Y=1.655 $X2=0.875 $Y2=2.38
cc_101 VPB N_GATE_c_167_n 0.00595129f $X=-0.19 $Y=1.655 $X2=0.39 $Y2=1.2
cc_102 VPB N_GATE_c_168_n 0.0265453f $X=-0.19 $Y=1.655 $X2=0.875 $Y2=1.37
cc_103 VPB N_SCE_M1000_g 0.0252032f $X=-0.19 $Y=1.655 $X2=0.885 $Y2=1.035
cc_104 VPB N_SCE_c_203_n 0.00636794f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_105 VPB N_SCE_c_204_n 0.00255333f $X=-0.19 $Y=1.655 $X2=0.39 $Y2=1.37
cc_106 VPB N_A_356_278#_M1006_g 0.0285111f $X=-0.19 $Y=1.655 $X2=0.885 $Y2=0.715
cc_107 VPB N_A_356_278#_M1021_g 0.0278157f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_108 VPB N_A_356_278#_c_265_n 0.00110614f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_109 VPB N_A_356_278#_c_275_n 0.0170506f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_110 VPB N_A_356_278#_c_266_n 0.00326884f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_111 VPB N_A_356_278#_c_277_n 0.00120828f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_112 VPB N_A_356_278#_c_267_n 0.0156777f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_113 VPB N_A_356_278#_c_279_n 0.00841556f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_114 VPB N_A_356_278#_c_270_n 0.00601076f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_115 VPB N_A_356_278#_c_271_n 0.0155637f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_116 VPB N_A_447_376#_c_435_n 0.00476372f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_117 VPB N_A_447_376#_M1002_g 0.0406972f $X=-0.19 $Y=1.655 $X2=0.885 $Y2=0.715
cc_118 VPB N_A_447_376#_c_438_n 0.026552f $X=-0.19 $Y=1.655 $X2=0.24 $Y2=1.37
cc_119 VPB N_A_447_376#_c_445_n 0.00855079f $X=-0.19 $Y=1.655 $X2=0.39 $Y2=1.37
cc_120 VPB N_A_447_376#_c_440_n 0.0128691f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_121 VPB N_A_860_21#_M1008_g 0.0253858f $X=-0.19 $Y=1.655 $X2=0.39 $Y2=1.37
cc_122 VPB N_A_860_21#_M1010_g 0.040715f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_123 VPB N_A_860_21#_c_526_n 0.00115338f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_124 VPB N_A_860_21#_c_515_n 0.0225197f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_125 VPB N_A_860_21#_c_528_n 0.0175635f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_126 VPB N_A_860_21#_c_529_n 0.00341465f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_127 VPB N_A_860_21#_c_518_n 0.00387523f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_128 VPB N_A_860_21#_c_531_n 0.00685109f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_129 VPB N_A_860_21#_c_532_n 0.0169931f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_130 VPB N_A_860_21#_c_520_n 6.48412e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_131 VPB N_A_698_405#_M1003_g 0.0455428f $X=-0.19 $Y=1.655 $X2=0.885 $Y2=0.715
cc_132 VPB N_A_698_405#_c_681_n 0.00311039f $X=-0.19 $Y=1.655 $X2=0.885 $Y2=1.37
cc_133 VPB N_A_698_405#_c_689_n 0.00693517f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_134 VPB N_CLK_M1007_g 0.040719f $X=-0.19 $Y=1.655 $X2=0.885 $Y2=1.035
cc_135 VPB N_CLK_M1025_g 0.0378927f $X=-0.19 $Y=1.655 $X2=0.39 $Y2=1.2
cc_136 VPB CLK 0.00724025f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_137 VPB N_CLK_c_768_n 0.0210201f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_138 VPB N_A_1384_416#_c_840_n 0.0240865f $X=-0.19 $Y=1.655 $X2=0.885
+ $Y2=0.715
cc_139 VPB N_A_1384_416#_c_841_n 0.0259318f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=1.37
cc_140 VPB N_A_1384_416#_c_842_n 0.0128631f $X=-0.19 $Y=1.655 $X2=0.875 $Y2=1.37
cc_141 VPB N_A_1384_416#_c_834_n 0.0120086f $X=-0.19 $Y=1.655 $X2=0.24 $Y2=1.37
cc_142 VPB N_A_1384_416#_c_835_n 0.00262795f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_143 VPB N_A_1384_416#_c_845_n 0.00930495f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_144 VPB N_A_93_376#_c_916_n 0.0341715f $X=-0.19 $Y=1.655 $X2=0.39 $Y2=1.2
cc_145 VPB N_A_93_376#_c_917_n 0.0156996f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_146 VPB N_A_93_376#_c_918_n 0.00920819f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_147 VPB N_A_93_376#_c_919_n 0.00597752f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_148 VPB N_A_93_376#_c_920_n 0.0017035f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_149 VPB N_VPWR_c_1021_n 0.00470917f $X=-0.19 $Y=1.655 $X2=0.39 $Y2=1.2
cc_150 VPB N_VPWR_c_1022_n 8.75318e-19 $X=-0.19 $Y=1.655 $X2=0.24 $Y2=1.37
cc_151 VPB N_VPWR_c_1023_n 0.00533208f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_152 VPB N_VPWR_c_1024_n 0.0214158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_153 VPB N_VPWR_c_1025_n 0.00631593f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_154 VPB N_VPWR_c_1026_n 0.045046f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_155 VPB N_VPWR_c_1027_n 0.0687569f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_156 VPB N_VPWR_c_1028_n 0.0402047f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_157 VPB N_VPWR_c_1029_n 0.02371f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_158 VPB N_VPWR_c_1020_n 0.112f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_159 VPB N_VPWR_c_1031_n 0.0170543f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_160 VPB N_VPWR_c_1032_n 0.00563917f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_161 VPB N_VPWR_c_1033_n 0.00454612f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_162 VPB GCLK 0.0173146f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_163 VPB GCLK 0.009439f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_164 VPB GCLK 0.0339839f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_165 N_GATE_c_166_n N_SCE_c_199_n 0.00979377f $X=0.885 $Y=1.035 $X2=-0.19
+ $Y2=-0.245
cc_166 N_GATE_c_168_n N_SCE_c_202_n 0.00979377f $X=0.875 $Y=1.37 $X2=0 $Y2=0
cc_167 N_GATE_M1018_g N_SCE_c_203_n 0.0509526f $X=0.875 $Y=2.38 $X2=0 $Y2=0
cc_168 N_GATE_c_168_n N_SCE_c_204_n 0.00593208f $X=0.875 $Y=1.37 $X2=0 $Y2=0
cc_169 N_GATE_c_168_n N_SCE_c_205_n 0.0509526f $X=0.875 $Y=1.37 $X2=0 $Y2=0
cc_170 N_GATE_M1018_g N_A_93_376#_c_916_n 0.0222518f $X=0.875 $Y=2.38 $X2=0
+ $Y2=0
cc_171 N_GATE_c_165_n N_A_93_376#_c_909_n 0.00741244f $X=0.495 $Y=1.035 $X2=0
+ $Y2=0
cc_172 N_GATE_c_166_n N_A_93_376#_c_909_n 0.0139334f $X=0.885 $Y=1.035 $X2=0
+ $Y2=0
cc_173 N_GATE_M1018_g N_A_93_376#_c_924_n 0.00896603f $X=0.875 $Y=2.38 $X2=0
+ $Y2=0
cc_174 N_GATE_M1018_g N_A_93_376#_c_918_n 0.00499348f $X=0.875 $Y=2.38 $X2=0
+ $Y2=0
cc_175 N_GATE_c_167_n N_A_93_376#_c_918_n 0.00909368f $X=0.39 $Y=1.2 $X2=0 $Y2=0
cc_176 N_GATE_c_168_n N_A_93_376#_c_918_n 0.0105393f $X=0.875 $Y=1.37 $X2=0
+ $Y2=0
cc_177 N_GATE_M1018_g N_A_93_376#_c_919_n 0.00631945f $X=0.875 $Y=2.38 $X2=0
+ $Y2=0
cc_178 N_GATE_c_167_n N_A_93_376#_c_919_n 0.0345636f $X=0.39 $Y=1.2 $X2=0 $Y2=0
cc_179 N_GATE_c_168_n N_A_93_376#_c_919_n 0.0198776f $X=0.875 $Y=1.37 $X2=0
+ $Y2=0
cc_180 N_GATE_c_167_n N_A_93_376#_c_914_n 0.0132756f $X=0.39 $Y=1.2 $X2=0 $Y2=0
cc_181 N_GATE_c_168_n N_A_93_376#_c_914_n 0.0141055f $X=0.875 $Y=1.37 $X2=0
+ $Y2=0
cc_182 N_GATE_M1018_g N_VPWR_c_1026_n 0.00649425f $X=0.875 $Y=2.38 $X2=0 $Y2=0
cc_183 N_GATE_M1018_g N_VPWR_c_1020_n 0.00867623f $X=0.875 $Y=2.38 $X2=0 $Y2=0
cc_184 N_GATE_c_165_n N_VGND_c_1140_n 0.0101424f $X=0.495 $Y=1.035 $X2=0 $Y2=0
cc_185 N_GATE_c_166_n N_VGND_c_1140_n 8.991e-19 $X=0.885 $Y=1.035 $X2=0 $Y2=0
cc_186 N_GATE_c_167_n N_VGND_c_1140_n 0.0244313f $X=0.39 $Y=1.2 $X2=0 $Y2=0
cc_187 N_GATE_c_168_n N_VGND_c_1140_n 0.00502558f $X=0.875 $Y=1.37 $X2=0 $Y2=0
cc_188 N_GATE_c_165_n N_VGND_c_1145_n 0.00402651f $X=0.495 $Y=1.035 $X2=0 $Y2=0
cc_189 N_GATE_c_166_n N_VGND_c_1145_n 0.00359585f $X=0.885 $Y=1.035 $X2=0 $Y2=0
cc_190 N_GATE_c_165_n N_VGND_c_1152_n 0.00423264f $X=0.495 $Y=1.035 $X2=0 $Y2=0
cc_191 N_GATE_c_166_n N_VGND_c_1152_n 0.00503886f $X=0.885 $Y=1.035 $X2=0 $Y2=0
cc_192 N_SCE_M1000_g N_A_356_278#_M1006_g 0.0286219f $X=1.365 $Y=2.38 $X2=0
+ $Y2=0
cc_193 N_SCE_c_204_n N_A_356_278#_M1006_g 0.00123175f $X=1.405 $Y=1.555 $X2=0
+ $Y2=0
cc_194 N_SCE_c_201_n N_A_356_278#_c_255_n 0.00970089f $X=1.675 $Y=1 $X2=0 $Y2=0
cc_195 N_SCE_c_205_n N_A_356_278#_c_256_n 0.00494918f $X=1.405 $Y=1.39 $X2=0
+ $Y2=0
cc_196 N_SCE_c_200_n N_A_356_278#_c_262_n 0.00970089f $X=1.6 $Y=1.075 $X2=0
+ $Y2=0
cc_197 N_SCE_M1000_g N_A_356_278#_c_265_n 0.0040909f $X=1.365 $Y=2.38 $X2=0
+ $Y2=0
cc_198 N_SCE_c_203_n N_A_356_278#_c_265_n 0.00114936f $X=1.405 $Y=1.555 $X2=0
+ $Y2=0
cc_199 N_SCE_c_204_n N_A_356_278#_c_265_n 0.0524477f $X=1.405 $Y=1.555 $X2=0
+ $Y2=0
cc_200 N_SCE_M1000_g N_A_356_278#_c_290_n 0.00434054f $X=1.365 $Y=2.38 $X2=0
+ $Y2=0
cc_201 N_SCE_c_203_n N_A_356_278#_c_271_n 0.0206108f $X=1.405 $Y=1.555 $X2=0
+ $Y2=0
cc_202 N_SCE_c_204_n N_A_356_278#_c_271_n 0.00121877f $X=1.405 $Y=1.555 $X2=0
+ $Y2=0
cc_203 N_SCE_M1000_g N_A_93_376#_c_916_n 0.00305219f $X=1.365 $Y=2.38 $X2=0
+ $Y2=0
cc_204 N_SCE_c_199_n N_A_93_376#_c_909_n 0.0102656f $X=1.315 $Y=1 $X2=0 $Y2=0
cc_205 N_SCE_c_201_n N_A_93_376#_c_909_n 0.00170895f $X=1.675 $Y=1 $X2=0 $Y2=0
cc_206 N_SCE_c_202_n N_A_93_376#_c_909_n 0.00235019f $X=1.315 $Y=1.075 $X2=0
+ $Y2=0
cc_207 N_SCE_M1000_g N_A_93_376#_c_924_n 0.0188296f $X=1.365 $Y=2.38 $X2=0 $Y2=0
cc_208 N_SCE_c_204_n N_A_93_376#_c_924_n 0.012982f $X=1.405 $Y=1.555 $X2=0 $Y2=0
cc_209 N_SCE_c_200_n N_A_93_376#_c_910_n 0.0231148f $X=1.6 $Y=1.075 $X2=0 $Y2=0
cc_210 N_SCE_c_202_n N_A_93_376#_c_910_n 0.00658743f $X=1.315 $Y=1.075 $X2=0
+ $Y2=0
cc_211 N_SCE_c_203_n N_A_93_376#_c_910_n 5.45825e-19 $X=1.405 $Y=1.555 $X2=0
+ $Y2=0
cc_212 N_SCE_c_204_n N_A_93_376#_c_910_n 0.0227565f $X=1.405 $Y=1.555 $X2=0
+ $Y2=0
cc_213 N_SCE_c_205_n N_A_93_376#_c_910_n 0.00357417f $X=1.405 $Y=1.39 $X2=0
+ $Y2=0
cc_214 N_SCE_M1000_g N_A_93_376#_c_918_n 3.18039e-19 $X=1.365 $Y=2.38 $X2=0
+ $Y2=0
cc_215 N_SCE_c_203_n N_A_93_376#_c_919_n 3.18039e-19 $X=1.405 $Y=1.555 $X2=0
+ $Y2=0
cc_216 N_SCE_c_204_n N_A_93_376#_c_919_n 0.057659f $X=1.405 $Y=1.555 $X2=0 $Y2=0
cc_217 N_SCE_c_205_n N_A_93_376#_c_919_n 9.51545e-19 $X=1.405 $Y=1.39 $X2=0
+ $Y2=0
cc_218 N_SCE_c_202_n N_A_93_376#_c_914_n 0.00156724f $X=1.315 $Y=1.075 $X2=0
+ $Y2=0
cc_219 N_SCE_c_204_n N_A_93_376#_c_914_n 0.0158731f $X=1.405 $Y=1.555 $X2=0
+ $Y2=0
cc_220 N_SCE_c_205_n N_A_93_376#_c_914_n 0.00116227f $X=1.405 $Y=1.39 $X2=0
+ $Y2=0
cc_221 N_SCE_M1000_g N_A_93_376#_c_920_n 0.00102723f $X=1.365 $Y=2.38 $X2=0
+ $Y2=0
cc_222 N_SCE_c_204_n A_200_376# 0.00409434f $X=1.405 $Y=1.555 $X2=-0.19
+ $Y2=-0.245
cc_223 N_SCE_c_204_n N_VPWR_M1000_d 0.00319188f $X=1.405 $Y=1.555 $X2=-0.19
+ $Y2=-0.245
cc_224 N_SCE_M1000_g N_VPWR_c_1026_n 0.00651444f $X=1.365 $Y=2.38 $X2=0 $Y2=0
cc_225 N_SCE_M1000_g N_VPWR_c_1020_n 0.00867623f $X=1.365 $Y=2.38 $X2=0 $Y2=0
cc_226 N_SCE_M1000_g N_VPWR_c_1031_n 0.00137428f $X=1.365 $Y=2.38 $X2=0 $Y2=0
cc_227 N_SCE_c_199_n N_VGND_c_1141_n 0.0015724f $X=1.315 $Y=1 $X2=0 $Y2=0
cc_228 N_SCE_c_201_n N_VGND_c_1141_n 0.0102638f $X=1.675 $Y=1 $X2=0 $Y2=0
cc_229 N_SCE_c_199_n N_VGND_c_1145_n 0.00464519f $X=1.315 $Y=1 $X2=0 $Y2=0
cc_230 N_SCE_c_201_n N_VGND_c_1145_n 0.00402651f $X=1.675 $Y=1 $X2=0 $Y2=0
cc_231 N_SCE_c_199_n N_VGND_c_1152_n 0.00503886f $X=1.315 $Y=1 $X2=0 $Y2=0
cc_232 N_SCE_c_201_n N_VGND_c_1152_n 0.00423264f $X=1.675 $Y=1 $X2=0 $Y2=0
cc_233 N_A_356_278#_c_293_p N_A_447_376#_M1006_d 0.00341813f $X=2.405 $Y=2.35
+ $X2=0 $Y2=0
cc_234 N_A_356_278#_c_275_n N_A_447_376#_M1006_d 0.00130239f $X=3.975 $Y=2.52
+ $X2=0 $Y2=0
cc_235 N_A_356_278#_c_295_p N_A_447_376#_M1006_d 0.0125549f $X=2.49 $Y=2.35
+ $X2=0 $Y2=0
cc_236 N_A_356_278#_c_260_n N_A_447_376#_c_435_n 0.0184679f $X=3.48 $Y=0.82
+ $X2=0 $Y2=0
cc_237 N_A_356_278#_c_264_n N_A_447_376#_c_435_n 0.00320021f $X=3.055 $Y=0.82
+ $X2=0 $Y2=0
cc_238 N_A_356_278#_c_266_n N_A_447_376#_c_435_n 0.00177428f $X=4.06 $Y=1.825
+ $X2=0 $Y2=0
cc_239 N_A_356_278#_c_267_n N_A_447_376#_c_435_n 0.0181559f $X=3.895 $Y=1.66
+ $X2=0 $Y2=0
cc_240 N_A_356_278#_M1021_g N_A_447_376#_M1002_g 0.0485073f $X=3.895 $Y=2.525
+ $X2=0 $Y2=0
cc_241 N_A_356_278#_c_275_n N_A_447_376#_M1002_g 0.0235467f $X=3.975 $Y=2.52
+ $X2=0 $Y2=0
cc_242 N_A_356_278#_c_277_n N_A_447_376#_M1002_g 8.06325e-19 $X=4.06 $Y=2.435
+ $X2=0 $Y2=0
cc_243 N_A_356_278#_c_295_p N_A_447_376#_M1002_g 0.00402421f $X=2.49 $Y=2.35
+ $X2=0 $Y2=0
cc_244 N_A_356_278#_c_266_n N_A_447_376#_c_436_n 0.0041815f $X=4.06 $Y=1.825
+ $X2=0 $Y2=0
cc_245 N_A_356_278#_c_267_n N_A_447_376#_c_436_n 0.0174905f $X=3.895 $Y=1.66
+ $X2=0 $Y2=0
cc_246 N_A_356_278#_c_261_n N_A_447_376#_M1026_g 0.0187178f $X=3.555 $Y=0.745
+ $X2=0 $Y2=0
cc_247 N_A_356_278#_c_259_n N_A_447_376#_c_438_n 0.0150517f $X=2.98 $Y=1.075
+ $X2=0 $Y2=0
cc_248 N_A_356_278#_c_260_n N_A_447_376#_c_438_n 0.00654725f $X=3.48 $Y=0.82
+ $X2=0 $Y2=0
cc_249 N_A_356_278#_c_271_n N_A_447_376#_c_438_n 0.00391708f $X=2.11 $Y=1.555
+ $X2=0 $Y2=0
cc_250 N_A_356_278#_M1006_g N_A_447_376#_c_445_n 0.00837638f $X=2.11 $Y=2.38
+ $X2=0 $Y2=0
cc_251 N_A_356_278#_c_265_n N_A_447_376#_c_445_n 0.0193998f $X=1.945 $Y=1.555
+ $X2=0 $Y2=0
cc_252 N_A_356_278#_c_293_p N_A_447_376#_c_445_n 0.00838038f $X=2.405 $Y=2.35
+ $X2=0 $Y2=0
cc_253 N_A_356_278#_c_275_n N_A_447_376#_c_445_n 0.00205938f $X=3.975 $Y=2.52
+ $X2=0 $Y2=0
cc_254 N_A_356_278#_c_295_p N_A_447_376#_c_445_n 0.0131611f $X=2.49 $Y=2.35
+ $X2=0 $Y2=0
cc_255 N_A_356_278#_c_256_n N_A_447_376#_c_439_n 0.00410395f $X=2.105 $Y=1.39
+ $X2=0 $Y2=0
cc_256 N_A_356_278#_c_258_n N_A_447_376#_c_439_n 4.41767e-19 $X=2.465 $Y=1 $X2=0
+ $Y2=0
cc_257 N_A_356_278#_c_259_n N_A_447_376#_c_439_n 0.0115466f $X=2.98 $Y=1.075
+ $X2=0 $Y2=0
cc_258 N_A_356_278#_c_264_n N_A_447_376#_c_439_n 7.34184e-19 $X=3.055 $Y=0.82
+ $X2=0 $Y2=0
cc_259 N_A_356_278#_c_257_n N_A_447_376#_c_440_n 7.10888e-19 $X=2.39 $Y=1.075
+ $X2=0 $Y2=0
cc_260 N_A_356_278#_c_259_n N_A_447_376#_c_440_n 0.00148662f $X=2.98 $Y=1.075
+ $X2=0 $Y2=0
cc_261 N_A_356_278#_c_260_n N_A_447_376#_c_440_n 3.73041e-19 $X=3.48 $Y=0.82
+ $X2=0 $Y2=0
cc_262 N_A_356_278#_c_263_n N_A_447_376#_c_440_n 0.0123433f $X=2.465 $Y=1.075
+ $X2=0 $Y2=0
cc_263 N_A_356_278#_c_265_n N_A_447_376#_c_440_n 0.0264912f $X=1.945 $Y=1.555
+ $X2=0 $Y2=0
cc_264 N_A_356_278#_c_271_n N_A_447_376#_c_440_n 0.00482329f $X=2.11 $Y=1.555
+ $X2=0 $Y2=0
cc_265 N_A_356_278#_c_258_n N_A_447_376#_c_441_n 0.00377315f $X=2.465 $Y=1 $X2=0
+ $Y2=0
cc_266 N_A_356_278#_c_259_n N_A_447_376#_c_441_n 0.00535332f $X=2.98 $Y=1.075
+ $X2=0 $Y2=0
cc_267 N_A_356_278#_c_261_n N_A_447_376#_c_441_n 0.00198385f $X=3.555 $Y=0.745
+ $X2=0 $Y2=0
cc_268 N_A_356_278#_c_264_n N_A_447_376#_c_441_n 0.00563069f $X=3.055 $Y=0.82
+ $X2=0 $Y2=0
cc_269 N_A_356_278#_c_266_n N_A_860_21#_M1024_g 0.00704817f $X=4.06 $Y=1.825
+ $X2=0 $Y2=0
cc_270 N_A_356_278#_c_267_n N_A_860_21#_M1024_g 0.0172874f $X=3.895 $Y=1.66
+ $X2=0 $Y2=0
cc_271 N_A_356_278#_c_268_n N_A_860_21#_M1024_g 0.0132113f $X=5.715 $Y=1.17
+ $X2=0 $Y2=0
cc_272 N_A_356_278#_c_275_n N_A_860_21#_M1008_g 0.00345416f $X=3.975 $Y=2.52
+ $X2=0 $Y2=0
cc_273 N_A_356_278#_M1021_g N_A_860_21#_c_526_n 5.01352e-19 $X=3.895 $Y=2.525
+ $X2=0 $Y2=0
cc_274 N_A_356_278#_c_266_n N_A_860_21#_c_526_n 0.0190054f $X=4.06 $Y=1.825
+ $X2=0 $Y2=0
cc_275 N_A_356_278#_c_277_n N_A_860_21#_c_526_n 0.035836f $X=4.06 $Y=2.435 $X2=0
+ $Y2=0
cc_276 N_A_356_278#_c_267_n N_A_860_21#_c_526_n 2.54027e-19 $X=3.895 $Y=1.66
+ $X2=0 $Y2=0
cc_277 N_A_356_278#_c_268_n N_A_860_21#_c_526_n 0.0246282f $X=5.715 $Y=1.17
+ $X2=0 $Y2=0
cc_278 N_A_356_278#_M1021_g N_A_860_21#_c_515_n 0.0608409f $X=3.895 $Y=2.525
+ $X2=0 $Y2=0
cc_279 N_A_356_278#_c_277_n N_A_860_21#_c_515_n 0.00381388f $X=4.06 $Y=2.435
+ $X2=0 $Y2=0
cc_280 N_A_356_278#_c_268_n N_A_860_21#_c_515_n 0.0052375f $X=5.715 $Y=1.17
+ $X2=0 $Y2=0
cc_281 N_A_356_278#_c_275_n N_A_860_21#_c_546_n 0.00543316f $X=3.975 $Y=2.52
+ $X2=0 $Y2=0
cc_282 N_A_356_278#_c_277_n N_A_860_21#_c_546_n 0.0078583f $X=4.06 $Y=2.435
+ $X2=0 $Y2=0
cc_283 N_A_356_278#_M1007_s N_A_860_21#_c_528_n 0.00758822f $X=5.855 $Y=2.08
+ $X2=0 $Y2=0
cc_284 N_A_356_278#_c_279_n N_A_860_21#_c_528_n 0.0206639f $X=6 $Y=2.225 $X2=0
+ $Y2=0
cc_285 N_A_356_278#_c_269_n N_A_860_21#_c_516_n 0.0160333f $X=5.94 $Y=1.17 $X2=0
+ $Y2=0
cc_286 N_A_356_278#_c_269_n N_A_860_21#_c_517_n 0.0185183f $X=5.94 $Y=1.17 $X2=0
+ $Y2=0
cc_287 N_A_356_278#_c_270_n N_A_860_21#_c_517_n 0.0120199f $X=6 $Y=2.06 $X2=0
+ $Y2=0
cc_288 N_A_356_278#_c_279_n N_A_860_21#_c_529_n 0.0170533f $X=6 $Y=2.225 $X2=0
+ $Y2=0
cc_289 N_A_356_278#_c_270_n N_A_860_21#_c_529_n 0.0147536f $X=6 $Y=2.06 $X2=0
+ $Y2=0
cc_290 N_A_356_278#_c_268_n N_A_860_21#_c_519_n 0.0094486f $X=5.715 $Y=1.17
+ $X2=0 $Y2=0
cc_291 N_A_356_278#_c_269_n N_A_860_21#_c_519_n 0.00377213f $X=5.94 $Y=1.17
+ $X2=0 $Y2=0
cc_292 N_A_356_278#_c_270_n N_A_860_21#_c_520_n 0.0117918f $X=6 $Y=2.06 $X2=0
+ $Y2=0
cc_293 N_A_356_278#_c_275_n N_A_698_405#_M1002_d 0.00497251f $X=3.975 $Y=2.52
+ $X2=0 $Y2=0
cc_294 N_A_356_278#_c_268_n N_A_698_405#_M1003_g 0.0192395f $X=5.715 $Y=1.17
+ $X2=0 $Y2=0
cc_295 N_A_356_278#_M1021_g N_A_698_405#_c_681_n 0.00142022f $X=3.895 $Y=2.525
+ $X2=0 $Y2=0
cc_296 N_A_356_278#_c_264_n N_A_698_405#_c_681_n 0.00163434f $X=3.055 $Y=0.82
+ $X2=0 $Y2=0
cc_297 N_A_356_278#_c_266_n N_A_698_405#_c_681_n 0.035487f $X=4.06 $Y=1.825
+ $X2=0 $Y2=0
cc_298 N_A_356_278#_c_277_n N_A_698_405#_c_681_n 0.00647858f $X=4.06 $Y=2.435
+ $X2=0 $Y2=0
cc_299 N_A_356_278#_c_267_n N_A_698_405#_c_681_n 0.00100913f $X=3.895 $Y=1.66
+ $X2=0 $Y2=0
cc_300 N_A_356_278#_c_261_n N_A_698_405#_c_682_n 0.00567533f $X=3.555 $Y=0.745
+ $X2=0 $Y2=0
cc_301 N_A_356_278#_c_260_n N_A_698_405#_c_683_n 0.0090824f $X=3.48 $Y=0.82
+ $X2=0 $Y2=0
cc_302 N_A_356_278#_c_264_n N_A_698_405#_c_683_n 0.00362009f $X=3.055 $Y=0.82
+ $X2=0 $Y2=0
cc_303 N_A_356_278#_c_266_n N_A_698_405#_c_683_n 0.00868865f $X=4.06 $Y=1.825
+ $X2=0 $Y2=0
cc_304 N_A_356_278#_M1021_g N_A_698_405#_c_689_n 0.00492906f $X=3.895 $Y=2.525
+ $X2=0 $Y2=0
cc_305 N_A_356_278#_c_275_n N_A_698_405#_c_689_n 0.0207709f $X=3.975 $Y=2.52
+ $X2=0 $Y2=0
cc_306 N_A_356_278#_c_266_n N_A_698_405#_c_689_n 0.00474393f $X=4.06 $Y=1.825
+ $X2=0 $Y2=0
cc_307 N_A_356_278#_c_277_n N_A_698_405#_c_689_n 0.017318f $X=4.06 $Y=2.435
+ $X2=0 $Y2=0
cc_308 N_A_356_278#_c_267_n N_A_698_405#_c_689_n 2.86873e-19 $X=3.895 $Y=1.66
+ $X2=0 $Y2=0
cc_309 N_A_356_278#_c_269_n N_A_698_405#_c_684_n 0.00436748f $X=5.94 $Y=1.17
+ $X2=0 $Y2=0
cc_310 N_A_356_278#_c_268_n N_A_698_405#_c_685_n 0.00886244f $X=5.715 $Y=1.17
+ $X2=0 $Y2=0
cc_311 N_A_356_278#_c_269_n N_A_698_405#_c_685_n 0.00543302f $X=5.94 $Y=1.17
+ $X2=0 $Y2=0
cc_312 N_A_356_278#_c_266_n N_A_698_405#_c_686_n 0.0130771f $X=4.06 $Y=1.825
+ $X2=0 $Y2=0
cc_313 N_A_356_278#_c_268_n N_A_698_405#_c_686_n 0.0784595f $X=5.715 $Y=1.17
+ $X2=0 $Y2=0
cc_314 N_A_356_278#_c_269_n N_CLK_c_760_n 0.00749784f $X=5.94 $Y=1.17 $X2=-0.19
+ $Y2=-0.245
cc_315 N_A_356_278#_c_270_n N_CLK_c_760_n 0.0134346f $X=6 $Y=2.06 $X2=-0.19
+ $Y2=-0.245
cc_316 N_A_356_278#_c_269_n N_CLK_c_761_n 0.00654503f $X=5.94 $Y=1.17 $X2=0
+ $Y2=0
cc_317 N_A_356_278#_c_270_n N_CLK_c_761_n 0.00167975f $X=6 $Y=2.06 $X2=0 $Y2=0
cc_318 N_A_356_278#_c_279_n N_CLK_M1007_g 0.00582324f $X=6 $Y=2.225 $X2=0 $Y2=0
cc_319 N_A_356_278#_c_270_n N_CLK_M1007_g 0.00684043f $X=6 $Y=2.06 $X2=0 $Y2=0
cc_320 N_A_356_278#_c_269_n N_CLK_c_763_n 3.59804e-19 $X=5.94 $Y=1.17 $X2=0
+ $Y2=0
cc_321 N_A_356_278#_c_279_n N_CLK_c_764_n 0.00330143f $X=6 $Y=2.225 $X2=0 $Y2=0
cc_322 N_A_356_278#_c_270_n N_CLK_c_764_n 0.00574672f $X=6 $Y=2.06 $X2=0 $Y2=0
cc_323 N_A_356_278#_c_268_n CLK 0.0550545f $X=5.715 $Y=1.17 $X2=0 $Y2=0
cc_324 N_A_356_278#_c_270_n CLK 0.0452319f $X=6 $Y=2.06 $X2=0 $Y2=0
cc_325 N_A_356_278#_c_268_n N_CLK_c_768_n 0.00645913f $X=5.715 $Y=1.17 $X2=0
+ $Y2=0
cc_326 N_A_356_278#_c_270_n N_CLK_c_768_n 6.92791e-19 $X=6 $Y=2.06 $X2=0 $Y2=0
cc_327 N_A_356_278#_c_275_n N_A_93_376#_M1002_s 0.0121002f $X=3.975 $Y=2.52
+ $X2=0 $Y2=0
cc_328 N_A_356_278#_M1006_g N_A_93_376#_c_924_n 0.00727788f $X=2.11 $Y=2.38
+ $X2=0 $Y2=0
cc_329 N_A_356_278#_c_290_n N_A_93_376#_c_924_n 0.0165861f $X=2.11 $Y=2.35 $X2=0
+ $Y2=0
cc_330 N_A_356_278#_c_256_n N_A_93_376#_c_910_n 0.00731758f $X=2.105 $Y=1.39
+ $X2=0 $Y2=0
cc_331 N_A_356_278#_c_257_n N_A_93_376#_c_910_n 0.00702722f $X=2.39 $Y=1.075
+ $X2=0 $Y2=0
cc_332 N_A_356_278#_c_262_n N_A_93_376#_c_910_n 0.0085808f $X=2.105 $Y=1.075
+ $X2=0 $Y2=0
cc_333 N_A_356_278#_c_263_n N_A_93_376#_c_910_n 0.00292563f $X=2.465 $Y=1.075
+ $X2=0 $Y2=0
cc_334 N_A_356_278#_c_265_n N_A_93_376#_c_910_n 0.0247989f $X=1.945 $Y=1.555
+ $X2=0 $Y2=0
cc_335 N_A_356_278#_c_271_n N_A_93_376#_c_910_n 0.00287998f $X=2.11 $Y=1.555
+ $X2=0 $Y2=0
cc_336 N_A_356_278#_M1006_g N_A_93_376#_c_917_n 0.00741896f $X=2.11 $Y=2.38
+ $X2=0 $Y2=0
cc_337 N_A_356_278#_M1021_g N_A_93_376#_c_917_n 0.00110056f $X=3.895 $Y=2.525
+ $X2=0 $Y2=0
cc_338 N_A_356_278#_c_293_p N_A_93_376#_c_917_n 0.00537843f $X=2.405 $Y=2.35
+ $X2=0 $Y2=0
cc_339 N_A_356_278#_c_275_n N_A_93_376#_c_917_n 0.0443931f $X=3.975 $Y=2.52
+ $X2=0 $Y2=0
cc_340 N_A_356_278#_c_295_p N_A_93_376#_c_917_n 0.0122106f $X=2.49 $Y=2.35 $X2=0
+ $Y2=0
cc_341 N_A_356_278#_c_255_n N_A_93_376#_c_911_n 0.00348793f $X=2.105 $Y=1 $X2=0
+ $Y2=0
cc_342 N_A_356_278#_c_257_n N_A_93_376#_c_911_n 0.00192385f $X=2.39 $Y=1.075
+ $X2=0 $Y2=0
cc_343 N_A_356_278#_c_258_n N_A_93_376#_c_911_n 0.0145568f $X=2.465 $Y=1 $X2=0
+ $Y2=0
cc_344 N_A_356_278#_c_263_n N_A_93_376#_c_911_n 8.99024e-19 $X=2.465 $Y=1.075
+ $X2=0 $Y2=0
cc_345 N_A_356_278#_c_258_n N_A_93_376#_c_912_n 0.0102609f $X=2.465 $Y=1 $X2=0
+ $Y2=0
cc_346 N_A_356_278#_c_264_n N_A_93_376#_c_912_n 0.00628993f $X=3.055 $Y=0.82
+ $X2=0 $Y2=0
cc_347 N_A_356_278#_c_255_n N_A_93_376#_c_913_n 4.39628e-19 $X=2.105 $Y=1 $X2=0
+ $Y2=0
cc_348 N_A_356_278#_c_258_n N_A_93_376#_c_913_n 6.78527e-19 $X=2.465 $Y=1 $X2=0
+ $Y2=0
cc_349 N_A_356_278#_M1006_g N_A_93_376#_c_920_n 0.0219837f $X=2.11 $Y=2.38 $X2=0
+ $Y2=0
cc_350 N_A_356_278#_c_293_p N_A_93_376#_c_920_n 0.00795121f $X=2.405 $Y=2.35
+ $X2=0 $Y2=0
cc_351 N_A_356_278#_c_290_n N_A_93_376#_c_920_n 0.00417655f $X=2.11 $Y=2.35
+ $X2=0 $Y2=0
cc_352 N_A_356_278#_c_258_n N_A_93_376#_c_915_n 0.00436159f $X=2.465 $Y=1 $X2=0
+ $Y2=0
cc_353 N_A_356_278#_c_260_n N_A_93_376#_c_915_n 0.0109457f $X=3.48 $Y=0.82 $X2=0
+ $Y2=0
cc_354 N_A_356_278#_c_261_n N_A_93_376#_c_915_n 0.00537328f $X=3.555 $Y=0.745
+ $X2=0 $Y2=0
cc_355 N_A_356_278#_c_265_n N_VPWR_M1000_d 0.00468157f $X=1.945 $Y=1.555
+ $X2=-0.19 $Y2=-0.245
cc_356 N_A_356_278#_c_290_n N_VPWR_M1000_d 0.00441009f $X=2.11 $Y=2.35 $X2=-0.19
+ $Y2=-0.245
cc_357 N_A_356_278#_M1021_g N_VPWR_c_1021_n 0.00219388f $X=3.895 $Y=2.525 $X2=0
+ $Y2=0
cc_358 N_A_356_278#_M1006_g N_VPWR_c_1027_n 0.00285527f $X=2.11 $Y=2.38 $X2=0
+ $Y2=0
cc_359 N_A_356_278#_M1021_g N_VPWR_c_1027_n 0.00635287f $X=3.895 $Y=2.525 $X2=0
+ $Y2=0
cc_360 N_A_356_278#_c_275_n N_VPWR_c_1027_n 0.0112036f $X=3.975 $Y=2.52 $X2=0
+ $Y2=0
cc_361 N_A_356_278#_M1006_g N_VPWR_c_1020_n 0.00249875f $X=2.11 $Y=2.38 $X2=0
+ $Y2=0
cc_362 N_A_356_278#_M1021_g N_VPWR_c_1020_n 0.00857631f $X=3.895 $Y=2.525 $X2=0
+ $Y2=0
cc_363 N_A_356_278#_c_275_n N_VPWR_c_1020_n 0.0225716f $X=3.975 $Y=2.52 $X2=0
+ $Y2=0
cc_364 N_A_356_278#_M1006_g N_VPWR_c_1031_n 4.45696e-19 $X=2.11 $Y=2.38 $X2=0
+ $Y2=0
cc_365 N_A_356_278#_c_275_n A_804_405# 0.00334823f $X=3.975 $Y=2.52 $X2=-0.19
+ $Y2=-0.245
cc_366 N_A_356_278#_c_277_n A_804_405# 0.00347854f $X=4.06 $Y=2.435 $X2=-0.19
+ $Y2=-0.245
cc_367 N_A_356_278#_c_255_n N_VGND_c_1141_n 0.00732974f $X=2.105 $Y=1 $X2=0
+ $Y2=0
cc_368 N_A_356_278#_c_258_n N_VGND_c_1141_n 3.8342e-19 $X=2.465 $Y=1 $X2=0 $Y2=0
cc_369 N_A_356_278#_c_255_n N_VGND_c_1149_n 0.00402651f $X=2.105 $Y=1 $X2=0
+ $Y2=0
cc_370 N_A_356_278#_c_258_n N_VGND_c_1149_n 7.27932e-19 $X=2.465 $Y=1 $X2=0
+ $Y2=0
cc_371 N_A_356_278#_c_260_n N_VGND_c_1149_n 2.80012e-19 $X=3.48 $Y=0.82 $X2=0
+ $Y2=0
cc_372 N_A_356_278#_c_261_n N_VGND_c_1149_n 0.00549284f $X=3.555 $Y=0.745 $X2=0
+ $Y2=0
cc_373 N_A_356_278#_c_255_n N_VGND_c_1152_n 0.00423264f $X=2.105 $Y=1 $X2=0
+ $Y2=0
cc_374 N_A_356_278#_c_261_n N_VGND_c_1152_n 0.0115186f $X=3.555 $Y=0.745 $X2=0
+ $Y2=0
cc_375 N_A_447_376#_M1026_g N_A_860_21#_M1024_g 0.0623602f $X=3.985 $Y=0.445
+ $X2=0 $Y2=0
cc_376 N_A_447_376#_c_435_n N_A_698_405#_c_681_n 0.0191959f $X=3.365 $Y=1.72
+ $X2=0 $Y2=0
cc_377 N_A_447_376#_M1002_g N_A_698_405#_c_681_n 0.0154127f $X=3.365 $Y=2.525
+ $X2=0 $Y2=0
cc_378 N_A_447_376#_c_436_n N_A_698_405#_c_681_n 0.00818566f $X=3.91 $Y=1.18
+ $X2=0 $Y2=0
cc_379 N_A_447_376#_M1026_g N_A_698_405#_c_681_n 0.00152495f $X=3.985 $Y=0.445
+ $X2=0 $Y2=0
cc_380 N_A_447_376#_c_439_n N_A_698_405#_c_681_n 0.012451f $X=2.885 $Y=1.39
+ $X2=0 $Y2=0
cc_381 N_A_447_376#_c_440_n N_A_698_405#_c_681_n 0.0238596f $X=3.035 $Y=1.555
+ $X2=0 $Y2=0
cc_382 N_A_447_376#_M1026_g N_A_698_405#_c_682_n 0.0128265f $X=3.985 $Y=0.445
+ $X2=0 $Y2=0
cc_383 N_A_447_376#_c_435_n N_A_698_405#_c_683_n 2.49984e-19 $X=3.365 $Y=1.72
+ $X2=0 $Y2=0
cc_384 N_A_447_376#_c_436_n N_A_698_405#_c_683_n 0.0103206f $X=3.91 $Y=1.18
+ $X2=0 $Y2=0
cc_385 N_A_447_376#_M1026_g N_A_698_405#_c_683_n 0.00453079f $X=3.985 $Y=0.445
+ $X2=0 $Y2=0
cc_386 N_A_447_376#_c_439_n N_A_698_405#_c_683_n 0.00456709f $X=2.885 $Y=1.39
+ $X2=0 $Y2=0
cc_387 N_A_447_376#_c_441_n N_A_698_405#_c_683_n 0.00298219f $X=2.885 $Y=0.78
+ $X2=0 $Y2=0
cc_388 N_A_447_376#_M1002_g N_A_698_405#_c_689_n 0.0151911f $X=3.365 $Y=2.525
+ $X2=0 $Y2=0
cc_389 N_A_447_376#_M1026_g N_A_698_405#_c_686_n 0.0108893f $X=3.985 $Y=0.445
+ $X2=0 $Y2=0
cc_390 N_A_447_376#_c_439_n N_A_93_376#_c_910_n 0.00706198f $X=2.885 $Y=1.39
+ $X2=0 $Y2=0
cc_391 N_A_447_376#_c_440_n N_A_93_376#_c_910_n 0.00976759f $X=3.035 $Y=1.555
+ $X2=0 $Y2=0
cc_392 N_A_447_376#_M1006_d N_A_93_376#_c_917_n 0.00480708f $X=2.235 $Y=1.88
+ $X2=0 $Y2=0
cc_393 N_A_447_376#_M1002_g N_A_93_376#_c_917_n 0.00665394f $X=3.365 $Y=2.525
+ $X2=0 $Y2=0
cc_394 N_A_447_376#_c_439_n N_A_93_376#_c_911_n 0.00343975f $X=2.885 $Y=1.39
+ $X2=0 $Y2=0
cc_395 N_A_447_376#_c_441_n N_A_93_376#_c_911_n 0.0109205f $X=2.885 $Y=0.78
+ $X2=0 $Y2=0
cc_396 N_A_447_376#_c_441_n N_A_93_376#_c_912_n 0.0261957f $X=2.885 $Y=0.78
+ $X2=0 $Y2=0
cc_397 N_A_447_376#_c_441_n N_A_93_376#_c_915_n 0.00436704f $X=2.885 $Y=0.78
+ $X2=0 $Y2=0
cc_398 N_A_447_376#_M1002_g N_VPWR_c_1027_n 0.00624975f $X=3.365 $Y=2.525 $X2=0
+ $Y2=0
cc_399 N_A_447_376#_M1002_g N_VPWR_c_1020_n 0.00913771f $X=3.365 $Y=2.525 $X2=0
+ $Y2=0
cc_400 N_A_447_376#_M1026_g N_VGND_c_1142_n 0.00239701f $X=3.985 $Y=0.445 $X2=0
+ $Y2=0
cc_401 N_A_447_376#_M1026_g N_VGND_c_1149_n 0.00549284f $X=3.985 $Y=0.445 $X2=0
+ $Y2=0
cc_402 N_A_447_376#_M1026_g N_VGND_c_1152_n 0.0100377f $X=3.985 $Y=0.445 $X2=0
+ $Y2=0
cc_403 N_A_860_21#_M1008_g N_A_698_405#_M1003_g 0.0358667f $X=4.425 $Y=2.525
+ $X2=0 $Y2=0
cc_404 N_A_860_21#_c_526_n N_A_698_405#_M1003_g 0.00728698f $X=4.49 $Y=1.7 $X2=0
+ $Y2=0
cc_405 N_A_860_21#_c_515_n N_A_698_405#_M1003_g 0.0205957f $X=4.49 $Y=1.7 $X2=0
+ $Y2=0
cc_406 N_A_860_21#_c_562_p N_A_698_405#_M1003_g 0.0164395f $X=5.09 $Y=2.415
+ $X2=0 $Y2=0
cc_407 N_A_860_21#_c_531_n N_A_698_405#_M1003_g 0.00455951f $X=5.255 $Y=2.415
+ $X2=0 $Y2=0
cc_408 N_A_860_21#_c_532_n N_A_698_405#_M1003_g 0.00609848f $X=5.255 $Y=2.575
+ $X2=0 $Y2=0
cc_409 N_A_860_21#_M1024_g N_A_698_405#_c_679_n 0.0184168f $X=4.375 $Y=0.445
+ $X2=0 $Y2=0
cc_410 N_A_860_21#_c_519_n N_A_698_405#_c_679_n 0.00203234f $X=5.61 $Y=0.47
+ $X2=0 $Y2=0
cc_411 N_A_860_21#_c_519_n N_A_698_405#_c_680_n 0.00851396f $X=5.61 $Y=0.47
+ $X2=0 $Y2=0
cc_412 N_A_860_21#_M1024_g N_A_698_405#_c_682_n 0.00218328f $X=4.375 $Y=0.445
+ $X2=0 $Y2=0
cc_413 N_A_860_21#_M1024_g N_A_698_405#_c_684_n 6.14756e-19 $X=4.375 $Y=0.445
+ $X2=0 $Y2=0
cc_414 N_A_860_21#_M1024_g N_A_698_405#_c_685_n 0.0144298f $X=4.375 $Y=0.445
+ $X2=0 $Y2=0
cc_415 N_A_860_21#_M1024_g N_A_698_405#_c_686_n 0.0150151f $X=4.375 $Y=0.445
+ $X2=0 $Y2=0
cc_416 N_A_860_21#_c_516_n N_CLK_c_761_n 0.00597177f $X=6.225 $Y=0.59 $X2=0
+ $Y2=0
cc_417 N_A_860_21#_c_517_n N_CLK_c_761_n 0.00449682f $X=6.31 $Y=1.58 $X2=0 $Y2=0
cc_418 N_A_860_21#_c_528_n N_CLK_M1007_g 0.0204741f $X=6.345 $Y=2.575 $X2=0
+ $Y2=0
cc_419 N_A_860_21#_c_529_n N_CLK_M1007_g 0.0229073f $X=6.43 $Y=2.49 $X2=0 $Y2=0
cc_420 N_A_860_21#_c_520_n N_CLK_M1007_g 0.0073588f $X=6.43 $Y=1.665 $X2=0 $Y2=0
cc_421 N_A_860_21#_c_577_p N_CLK_M1007_g 0.00357905f $X=6.43 $Y=2.575 $X2=0
+ $Y2=0
cc_422 N_A_860_21#_c_517_n N_CLK_c_763_n 0.0104414f $X=6.31 $Y=1.58 $X2=0 $Y2=0
cc_423 N_A_860_21#_c_514_n N_CLK_c_764_n 0.0205589f $X=7.325 $Y=1.53 $X2=0 $Y2=0
cc_424 N_A_860_21#_c_517_n N_CLK_c_764_n 0.0103026f $X=6.31 $Y=1.58 $X2=0 $Y2=0
cc_425 N_A_860_21#_c_520_n N_CLK_c_764_n 0.0109247f $X=6.43 $Y=1.665 $X2=0 $Y2=0
cc_426 N_A_860_21#_M1010_g N_CLK_M1025_g 0.0608318f $X=7.325 $Y=2.58 $X2=0 $Y2=0
cc_427 N_A_860_21#_c_529_n N_CLK_M1025_g 0.0126328f $X=6.43 $Y=2.49 $X2=0 $Y2=0
cc_428 N_A_860_21#_c_584_p N_CLK_M1025_g 0.0239177f $X=7.755 $Y=2.575 $X2=0
+ $Y2=0
cc_429 N_A_860_21#_c_520_n N_CLK_M1025_g 0.00343114f $X=6.43 $Y=1.665 $X2=0
+ $Y2=0
cc_430 N_A_860_21#_c_512_n N_CLK_c_766_n 0.0205589f $X=7.275 $Y=1.455 $X2=0
+ $Y2=0
cc_431 N_A_860_21#_c_517_n N_CLK_c_766_n 5.17572e-19 $X=6.31 $Y=1.58 $X2=0 $Y2=0
cc_432 N_A_860_21#_M1003_d CLK 0.00318129f $X=5.115 $Y=2.025 $X2=0 $Y2=0
cc_433 N_A_860_21#_M1008_g CLK 2.84609e-19 $X=4.425 $Y=2.525 $X2=0 $Y2=0
cc_434 N_A_860_21#_c_526_n CLK 0.0322719f $X=4.49 $Y=1.7 $X2=0 $Y2=0
cc_435 N_A_860_21#_c_515_n CLK 9.14216e-19 $X=4.49 $Y=1.7 $X2=0 $Y2=0
cc_436 N_A_860_21#_c_562_p CLK 0.0117706f $X=5.09 $Y=2.415 $X2=0 $Y2=0
cc_437 N_A_860_21#_c_528_n CLK 0.0120562f $X=6.345 $Y=2.575 $X2=0 $Y2=0
cc_438 N_A_860_21#_c_531_n CLK 0.0229823f $X=5.255 $Y=2.415 $X2=0 $Y2=0
cc_439 N_A_860_21#_c_528_n N_CLK_c_768_n 8.67584e-19 $X=6.345 $Y=2.575 $X2=0
+ $Y2=0
cc_440 N_A_860_21#_c_531_n N_CLK_c_768_n 4.0267e-19 $X=5.255 $Y=2.415 $X2=0
+ $Y2=0
cc_441 N_A_860_21#_c_584_p N_A_1384_416#_M1025_d 0.00481389f $X=7.755 $Y=2.575
+ $X2=0 $Y2=0
cc_442 N_A_860_21#_c_584_p N_A_1384_416#_c_840_n 0.00676895f $X=7.755 $Y=2.575
+ $X2=0 $Y2=0
cc_443 N_A_860_21#_c_518_n N_A_1384_416#_c_840_n 0.0135283f $X=7.84 $Y=2.49
+ $X2=0 $Y2=0
cc_444 N_A_860_21#_M1010_g N_A_1384_416#_c_842_n 0.0331657f $X=7.325 $Y=2.58
+ $X2=0 $Y2=0
cc_445 N_A_860_21#_c_518_n N_A_1384_416#_c_842_n 0.00541751f $X=7.84 $Y=2.49
+ $X2=0 $Y2=0
cc_446 N_A_860_21#_c_521_n N_A_1384_416#_c_842_n 0.00122569f $X=7.92 $Y=1.48
+ $X2=0 $Y2=0
cc_447 N_A_860_21#_c_522_n N_A_1384_416#_c_842_n 0.0129762f $X=7.92 $Y=1.48
+ $X2=0 $Y2=0
cc_448 N_A_860_21#_c_518_n N_A_1384_416#_c_834_n 6.71092e-19 $X=7.84 $Y=2.49
+ $X2=0 $Y2=0
cc_449 N_A_860_21#_c_521_n N_A_1384_416#_c_834_n 3.94517e-19 $X=7.92 $Y=1.48
+ $X2=0 $Y2=0
cc_450 N_A_860_21#_c_522_n N_A_1384_416#_c_834_n 0.0178856f $X=7.92 $Y=1.48
+ $X2=0 $Y2=0
cc_451 N_A_860_21#_c_512_n N_A_1384_416#_c_835_n 0.00684684f $X=7.275 $Y=1.455
+ $X2=0 $Y2=0
cc_452 N_A_860_21#_M1010_g N_A_1384_416#_c_835_n 0.0181925f $X=7.325 $Y=2.58
+ $X2=0 $Y2=0
cc_453 N_A_860_21#_c_514_n N_A_1384_416#_c_835_n 0.00627647f $X=7.325 $Y=1.53
+ $X2=0 $Y2=0
cc_454 N_A_860_21#_c_521_n N_A_1384_416#_c_835_n 0.0546271f $X=7.92 $Y=1.48
+ $X2=0 $Y2=0
cc_455 N_A_860_21#_c_522_n N_A_1384_416#_c_835_n 0.00137308f $X=7.92 $Y=1.48
+ $X2=0 $Y2=0
cc_456 N_A_860_21#_c_523_n N_A_1384_416#_c_835_n 0.00955949f $X=7.755 $Y=1.48
+ $X2=0 $Y2=0
cc_457 N_A_860_21#_c_521_n N_A_1384_416#_c_836_n 0.00129388f $X=7.92 $Y=1.48
+ $X2=0 $Y2=0
cc_458 N_A_860_21#_c_523_n N_A_1384_416#_c_836_n 0.00349763f $X=7.755 $Y=1.48
+ $X2=0 $Y2=0
cc_459 N_A_860_21#_c_512_n N_A_1384_416#_c_837_n 0.00367566f $X=7.275 $Y=1.455
+ $X2=0 $Y2=0
cc_460 N_A_860_21#_M1010_g N_A_1384_416#_c_845_n 0.0174598f $X=7.325 $Y=2.58
+ $X2=0 $Y2=0
cc_461 N_A_860_21#_c_529_n N_A_1384_416#_c_845_n 0.0103748f $X=6.43 $Y=2.49
+ $X2=0 $Y2=0
cc_462 N_A_860_21#_c_584_p N_A_1384_416#_c_845_n 0.0308954f $X=7.755 $Y=2.575
+ $X2=0 $Y2=0
cc_463 N_A_860_21#_c_518_n N_A_1384_416#_c_845_n 0.0157494f $X=7.84 $Y=2.49
+ $X2=0 $Y2=0
cc_464 N_A_860_21#_c_512_n N_A_1384_416#_c_838_n 5.55961e-19 $X=7.275 $Y=1.455
+ $X2=0 $Y2=0
cc_465 N_A_860_21#_c_521_n N_A_1384_416#_c_838_n 0.0202407f $X=7.92 $Y=1.48
+ $X2=0 $Y2=0
cc_466 N_A_860_21#_c_522_n N_A_1384_416#_c_838_n 3.89635e-19 $X=7.92 $Y=1.48
+ $X2=0 $Y2=0
cc_467 N_A_860_21#_c_512_n N_A_1384_416#_c_839_n 0.00777008f $X=7.275 $Y=1.455
+ $X2=0 $Y2=0
cc_468 N_A_860_21#_c_521_n N_A_1384_416#_c_839_n 3.84356e-19 $X=7.92 $Y=1.48
+ $X2=0 $Y2=0
cc_469 N_A_860_21#_c_522_n N_A_1384_416#_c_839_n 0.020691f $X=7.92 $Y=1.48 $X2=0
+ $Y2=0
cc_470 N_A_860_21#_c_523_n N_A_1384_416#_c_839_n 0.00233268f $X=7.755 $Y=1.48
+ $X2=0 $Y2=0
cc_471 N_A_860_21#_c_526_n N_VPWR_M1008_d 0.00362077f $X=4.49 $Y=1.7 $X2=0 $Y2=0
cc_472 N_A_860_21#_c_562_p N_VPWR_M1008_d 0.00743015f $X=5.09 $Y=2.415 $X2=0
+ $Y2=0
cc_473 N_A_860_21#_c_546_n N_VPWR_M1008_d 5.24955e-19 $X=4.655 $Y=2.415 $X2=0
+ $Y2=0
cc_474 N_A_860_21#_c_529_n N_VPWR_M1007_d 0.00472499f $X=6.43 $Y=2.49 $X2=0
+ $Y2=0
cc_475 N_A_860_21#_c_584_p N_VPWR_M1007_d 0.00472161f $X=7.755 $Y=2.575 $X2=0
+ $Y2=0
cc_476 N_A_860_21#_c_577_p N_VPWR_M1007_d 7.33924e-19 $X=6.43 $Y=2.575 $X2=0
+ $Y2=0
cc_477 N_A_860_21#_c_584_p N_VPWR_M1010_d 0.0118912f $X=7.755 $Y=2.575 $X2=0
+ $Y2=0
cc_478 N_A_860_21#_c_518_n N_VPWR_M1010_d 0.0048048f $X=7.84 $Y=2.49 $X2=0 $Y2=0
cc_479 N_A_860_21#_M1008_g N_VPWR_c_1021_n 0.0120899f $X=4.425 $Y=2.525 $X2=0
+ $Y2=0
cc_480 N_A_860_21#_c_562_p N_VPWR_c_1021_n 0.011574f $X=5.09 $Y=2.415 $X2=0
+ $Y2=0
cc_481 N_A_860_21#_c_546_n N_VPWR_c_1021_n 0.0058241f $X=4.655 $Y=2.415 $X2=0
+ $Y2=0
cc_482 N_A_860_21#_c_532_n N_VPWR_c_1021_n 0.0112035f $X=5.255 $Y=2.575 $X2=0
+ $Y2=0
cc_483 N_A_860_21#_M1010_g N_VPWR_c_1022_n 0.00186015f $X=7.325 $Y=2.58 $X2=0
+ $Y2=0
cc_484 N_A_860_21#_c_584_p N_VPWR_c_1022_n 0.00875035f $X=7.755 $Y=2.575 $X2=0
+ $Y2=0
cc_485 N_A_860_21#_c_577_p N_VPWR_c_1022_n 0.00723599f $X=6.43 $Y=2.575 $X2=0
+ $Y2=0
cc_486 N_A_860_21#_M1010_g N_VPWR_c_1023_n 0.00476977f $X=7.325 $Y=2.58 $X2=0
+ $Y2=0
cc_487 N_A_860_21#_c_584_p N_VPWR_c_1023_n 0.0244081f $X=7.755 $Y=2.575 $X2=0
+ $Y2=0
cc_488 N_A_860_21#_M1010_g N_VPWR_c_1024_n 0.00695957f $X=7.325 $Y=2.58 $X2=0
+ $Y2=0
cc_489 N_A_860_21#_c_584_p N_VPWR_c_1024_n 0.0113397f $X=7.755 $Y=2.575 $X2=0
+ $Y2=0
cc_490 N_A_860_21#_M1008_g N_VPWR_c_1027_n 0.00774619f $X=4.425 $Y=2.525 $X2=0
+ $Y2=0
cc_491 N_A_860_21#_c_528_n N_VPWR_c_1028_n 0.0146589f $X=6.345 $Y=2.575 $X2=0
+ $Y2=0
cc_492 N_A_860_21#_c_532_n N_VPWR_c_1028_n 0.0197499f $X=5.255 $Y=2.575 $X2=0
+ $Y2=0
cc_493 N_A_860_21#_c_577_p N_VPWR_c_1028_n 3.22416e-19 $X=6.43 $Y=2.575 $X2=0
+ $Y2=0
cc_494 N_A_860_21#_c_584_p N_VPWR_c_1029_n 0.00105582f $X=7.755 $Y=2.575 $X2=0
+ $Y2=0
cc_495 N_A_860_21#_M1008_g N_VPWR_c_1020_n 0.00824529f $X=4.425 $Y=2.525 $X2=0
+ $Y2=0
cc_496 N_A_860_21#_M1010_g N_VPWR_c_1020_n 0.00915201f $X=7.325 $Y=2.58 $X2=0
+ $Y2=0
cc_497 N_A_860_21#_c_562_p N_VPWR_c_1020_n 0.00727245f $X=5.09 $Y=2.415 $X2=0
+ $Y2=0
cc_498 N_A_860_21#_c_546_n N_VPWR_c_1020_n 0.00690593f $X=4.655 $Y=2.415 $X2=0
+ $Y2=0
cc_499 N_A_860_21#_c_528_n N_VPWR_c_1020_n 0.0246914f $X=6.345 $Y=2.575 $X2=0
+ $Y2=0
cc_500 N_A_860_21#_c_584_p N_VPWR_c_1020_n 0.0249569f $X=7.755 $Y=2.575 $X2=0
+ $Y2=0
cc_501 N_A_860_21#_c_532_n N_VPWR_c_1020_n 0.0124713f $X=5.255 $Y=2.575 $X2=0
+ $Y2=0
cc_502 N_A_860_21#_c_577_p N_VPWR_c_1020_n 0.00124515f $X=6.43 $Y=2.575 $X2=0
+ $Y2=0
cc_503 N_A_860_21#_c_518_n GCLK 0.0175754f $X=7.84 $Y=2.49 $X2=0 $Y2=0
cc_504 N_A_860_21#_c_521_n GCLK 0.0224717f $X=7.92 $Y=1.48 $X2=0 $Y2=0
cc_505 N_A_860_21#_c_522_n GCLK 0.00202814f $X=7.92 $Y=1.48 $X2=0 $Y2=0
cc_506 N_A_860_21#_c_518_n GCLK 0.0284642f $X=7.84 $Y=2.49 $X2=0 $Y2=0
cc_507 N_A_860_21#_M1010_g GCLK 8.8466e-19 $X=7.325 $Y=2.58 $X2=0 $Y2=0
cc_508 N_A_860_21#_c_584_p GCLK 0.012582f $X=7.755 $Y=2.575 $X2=0 $Y2=0
cc_509 N_A_860_21#_M1024_g N_VGND_c_1142_n 0.013565f $X=4.375 $Y=0.445 $X2=0
+ $Y2=0
cc_510 N_A_860_21#_c_512_n N_VGND_c_1143_n 0.00184127f $X=7.275 $Y=1.455 $X2=0
+ $Y2=0
cc_511 N_A_860_21#_c_516_n N_VGND_c_1143_n 0.01353f $X=6.225 $Y=0.59 $X2=0 $Y2=0
cc_512 N_A_860_21#_c_517_n N_VGND_c_1143_n 0.0342135f $X=6.31 $Y=1.58 $X2=0
+ $Y2=0
cc_513 N_A_860_21#_c_512_n N_VGND_c_1144_n 0.00364971f $X=7.275 $Y=1.455 $X2=0
+ $Y2=0
cc_514 N_A_860_21#_c_516_n N_VGND_c_1147_n 0.01575f $X=6.225 $Y=0.59 $X2=0 $Y2=0
cc_515 N_A_860_21#_c_519_n N_VGND_c_1147_n 0.0191504f $X=5.61 $Y=0.47 $X2=0
+ $Y2=0
cc_516 N_A_860_21#_M1024_g N_VGND_c_1149_n 0.00486043f $X=4.375 $Y=0.445 $X2=0
+ $Y2=0
cc_517 N_A_860_21#_M1004_d N_VGND_c_1152_n 0.00232985f $X=5.47 $Y=0.235 $X2=0
+ $Y2=0
cc_518 N_A_860_21#_M1024_g N_VGND_c_1152_n 0.00827383f $X=4.375 $Y=0.445 $X2=0
+ $Y2=0
cc_519 N_A_860_21#_c_512_n N_VGND_c_1152_n 0.00169847f $X=7.275 $Y=1.455 $X2=0
+ $Y2=0
cc_520 N_A_860_21#_c_516_n N_VGND_c_1152_n 0.0198723f $X=6.225 $Y=0.59 $X2=0
+ $Y2=0
cc_521 N_A_860_21#_c_519_n N_VGND_c_1152_n 0.0124135f $X=5.61 $Y=0.47 $X2=0
+ $Y2=0
cc_522 N_A_698_405#_c_685_n N_CLK_c_761_n 0.00166739f $X=5.1 $Y=0.93 $X2=0 $Y2=0
cc_523 N_A_698_405#_M1003_g CLK 0.0295788f $X=4.99 $Y=2.525 $X2=0 $Y2=0
cc_524 N_A_698_405#_M1003_g N_CLK_c_768_n 0.0219904f $X=4.99 $Y=2.525 $X2=0
+ $Y2=0
cc_525 N_A_698_405#_c_685_n N_CLK_c_768_n 0.00178711f $X=5.1 $Y=0.93 $X2=0 $Y2=0
cc_526 N_A_698_405#_c_682_n N_A_93_376#_c_915_n 0.0154229f $X=3.77 $Y=0.47 $X2=0
+ $Y2=0
cc_527 N_A_698_405#_c_683_n N_A_93_376#_c_915_n 0.00819257f $X=3.935 $Y=0.965
+ $X2=0 $Y2=0
cc_528 N_A_698_405#_M1003_g N_VPWR_c_1021_n 0.00311159f $X=4.99 $Y=2.525 $X2=0
+ $Y2=0
cc_529 N_A_698_405#_M1003_g N_VPWR_c_1028_n 0.00830671f $X=4.99 $Y=2.525 $X2=0
+ $Y2=0
cc_530 N_A_698_405#_M1003_g N_VPWR_c_1020_n 0.00932362f $X=4.99 $Y=2.525 $X2=0
+ $Y2=0
cc_531 N_A_698_405#_c_679_n N_VGND_c_1142_n 0.0135424f $X=5.005 $Y=0.735 $X2=0
+ $Y2=0
cc_532 N_A_698_405#_c_682_n N_VGND_c_1142_n 0.0127186f $X=3.77 $Y=0.47 $X2=0
+ $Y2=0
cc_533 N_A_698_405#_c_686_n N_VGND_c_1142_n 0.0240722f $X=4.935 $Y=0.907 $X2=0
+ $Y2=0
cc_534 N_A_698_405#_c_679_n N_VGND_c_1147_n 0.00585385f $X=5.005 $Y=0.735 $X2=0
+ $Y2=0
cc_535 N_A_698_405#_c_680_n N_VGND_c_1147_n 0.00549284f $X=5.395 $Y=0.735 $X2=0
+ $Y2=0
cc_536 N_A_698_405#_c_685_n N_VGND_c_1147_n 0.00110551f $X=5.1 $Y=0.93 $X2=0
+ $Y2=0
cc_537 N_A_698_405#_c_682_n N_VGND_c_1149_n 0.0143539f $X=3.77 $Y=0.47 $X2=0
+ $Y2=0
cc_538 N_A_698_405#_M1013_d N_VGND_c_1152_n 0.00420187f $X=3.63 $Y=0.235 $X2=0
+ $Y2=0
cc_539 N_A_698_405#_c_679_n N_VGND_c_1152_n 0.00684944f $X=5.005 $Y=0.735 $X2=0
+ $Y2=0
cc_540 N_A_698_405#_c_680_n N_VGND_c_1152_n 0.0113743f $X=5.395 $Y=0.735 $X2=0
+ $Y2=0
cc_541 N_A_698_405#_c_682_n N_VGND_c_1152_n 0.00945389f $X=3.77 $Y=0.47 $X2=0
+ $Y2=0
cc_542 N_A_698_405#_c_684_n N_VGND_c_1152_n 0.0110106f $X=5.1 $Y=0.93 $X2=0
+ $Y2=0
cc_543 N_A_698_405#_c_685_n N_VGND_c_1152_n 0.00146508f $X=5.1 $Y=0.93 $X2=0
+ $Y2=0
cc_544 N_CLK_M1025_g N_A_1384_416#_c_835_n 0.00234098f $X=6.795 $Y=2.58 $X2=0
+ $Y2=0
cc_545 N_CLK_c_766_n N_A_1384_416#_c_835_n 0.00198127f $X=6.885 $Y=1.455 $X2=0
+ $Y2=0
cc_546 N_CLK_c_766_n N_A_1384_416#_c_837_n 4.80837e-19 $X=6.885 $Y=1.455 $X2=0
+ $Y2=0
cc_547 N_CLK_M1007_g N_A_1384_416#_c_845_n 2.00158e-19 $X=6.265 $Y=2.58 $X2=0
+ $Y2=0
cc_548 N_CLK_c_764_n N_A_1384_416#_c_845_n 0.00127983f $X=6.795 $Y=1.605 $X2=0
+ $Y2=0
cc_549 N_CLK_M1025_g N_A_1384_416#_c_845_n 0.00601675f $X=6.795 $Y=2.58 $X2=0
+ $Y2=0
cc_550 N_CLK_M1007_g N_VPWR_c_1022_n 0.0161187f $X=6.265 $Y=2.58 $X2=0 $Y2=0
cc_551 N_CLK_M1025_g N_VPWR_c_1022_n 0.0101696f $X=6.795 $Y=2.58 $X2=0 $Y2=0
cc_552 N_CLK_M1025_g N_VPWR_c_1024_n 0.00625647f $X=6.795 $Y=2.58 $X2=0 $Y2=0
cc_553 N_CLK_M1007_g N_VPWR_c_1028_n 0.0062563f $X=6.265 $Y=2.58 $X2=0 $Y2=0
cc_554 N_CLK_M1007_g N_VPWR_c_1020_n 0.00840299f $X=6.265 $Y=2.58 $X2=0 $Y2=0
cc_555 N_CLK_M1025_g N_VPWR_c_1020_n 0.00715932f $X=6.795 $Y=2.58 $X2=0 $Y2=0
cc_556 N_CLK_c_763_n N_VGND_c_1143_n 0.00125495f $X=6.455 $Y=1.455 $X2=0 $Y2=0
cc_557 N_CLK_c_764_n N_VGND_c_1143_n 0.00548523f $X=6.795 $Y=1.605 $X2=0 $Y2=0
cc_558 N_CLK_c_766_n N_VGND_c_1143_n 0.0130087f $X=6.885 $Y=1.455 $X2=0 $Y2=0
cc_559 N_CLK_c_763_n N_VGND_c_1152_n 0.00348778f $X=6.455 $Y=1.455 $X2=0 $Y2=0
cc_560 N_CLK_c_766_n N_VGND_c_1152_n 0.00324254f $X=6.885 $Y=1.455 $X2=0 $Y2=0
cc_561 N_A_1384_416#_c_845_n N_VPWR_M1010_d 0.00232721f $X=7.06 $Y=2.225 $X2=0
+ $Y2=0
cc_562 N_A_1384_416#_c_840_n N_VPWR_c_1023_n 0.00476977f $X=8.015 $Y=2.005 $X2=0
+ $Y2=0
cc_563 N_A_1384_416#_c_840_n N_VPWR_c_1029_n 0.0087931f $X=8.015 $Y=2.005 $X2=0
+ $Y2=0
cc_564 N_A_1384_416#_c_840_n N_VPWR_c_1020_n 0.0161906f $X=8.015 $Y=2.005 $X2=0
+ $Y2=0
cc_565 N_A_1384_416#_c_832_n GCLK 9.02236e-19 $X=7.665 $Y=0.735 $X2=0 $Y2=0
cc_566 N_A_1384_416#_c_840_n GCLK 0.00131441f $X=8.015 $Y=2.005 $X2=0 $Y2=0
cc_567 N_A_1384_416#_c_833_n GCLK 0.0102863f $X=8.025 $Y=0.735 $X2=0 $Y2=0
cc_568 N_A_1384_416#_c_841_n GCLK 0.0136057f $X=8.325 $Y=1.93 $X2=0 $Y2=0
cc_569 N_A_1384_416#_c_834_n GCLK 0.0262036f $X=8.4 $Y=1.855 $X2=0 $Y2=0
cc_570 N_A_1384_416#_c_838_n GCLK 0.0248513f $X=7.94 $Y=0.94 $X2=0 $Y2=0
cc_571 N_A_1384_416#_c_839_n GCLK 0.0304719f $X=8.025 $Y=0.92 $X2=0 $Y2=0
cc_572 N_A_1384_416#_c_840_n GCLK 0.00486759f $X=8.015 $Y=2.005 $X2=0 $Y2=0
cc_573 N_A_1384_416#_c_841_n GCLK 0.00673816f $X=8.325 $Y=1.93 $X2=0 $Y2=0
cc_574 N_A_1384_416#_c_840_n GCLK 0.0205585f $X=8.015 $Y=2.005 $X2=0 $Y2=0
cc_575 N_A_1384_416#_c_835_n N_VGND_c_1143_n 0.00894133f $X=7.49 $Y=1.17 $X2=0
+ $Y2=0
cc_576 N_A_1384_416#_c_837_n N_VGND_c_1143_n 0.00541809f $X=7.575 $Y=1.02 $X2=0
+ $Y2=0
cc_577 N_A_1384_416#_c_832_n N_VGND_c_1144_n 0.0129599f $X=7.665 $Y=0.735 $X2=0
+ $Y2=0
cc_578 N_A_1384_416#_c_833_n N_VGND_c_1144_n 0.00247568f $X=8.025 $Y=0.735 $X2=0
+ $Y2=0
cc_579 N_A_1384_416#_c_836_n N_VGND_c_1144_n 0.00116079f $X=7.775 $Y=1.02 $X2=0
+ $Y2=0
cc_580 N_A_1384_416#_c_837_n N_VGND_c_1144_n 0.0174924f $X=7.575 $Y=1.02 $X2=0
+ $Y2=0
cc_581 N_A_1384_416#_c_832_n N_VGND_c_1151_n 0.00559147f $X=7.665 $Y=0.735 $X2=0
+ $Y2=0
cc_582 N_A_1384_416#_c_833_n N_VGND_c_1151_n 0.00542974f $X=8.025 $Y=0.735 $X2=0
+ $Y2=0
cc_583 N_A_1384_416#_c_839_n N_VGND_c_1151_n 5.55121e-19 $X=8.025 $Y=0.92 $X2=0
+ $Y2=0
cc_584 N_A_1384_416#_c_832_n N_VGND_c_1152_n 0.00936293f $X=7.665 $Y=0.735 $X2=0
+ $Y2=0
cc_585 N_A_1384_416#_c_833_n N_VGND_c_1152_n 0.00695377f $X=8.025 $Y=0.735 $X2=0
+ $Y2=0
cc_586 N_A_1384_416#_c_838_n N_VGND_c_1152_n 0.0101022f $X=7.94 $Y=0.94 $X2=0
+ $Y2=0
cc_587 N_A_1384_416#_c_839_n N_VGND_c_1152_n 7.35503e-19 $X=8.025 $Y=0.92 $X2=0
+ $Y2=0
cc_588 N_A_93_376#_c_924_n A_200_376# 0.00474891f $X=2.055 $Y=2.7 $X2=-0.19
+ $Y2=-0.245
cc_589 N_A_93_376#_c_924_n N_VPWR_M1000_d 0.0154205f $X=2.055 $Y=2.7 $X2=-0.19
+ $Y2=-0.245
cc_590 N_A_93_376#_c_916_n N_VPWR_c_1026_n 0.0139457f $X=0.675 $Y=2.615 $X2=0
+ $Y2=0
cc_591 N_A_93_376#_c_924_n N_VPWR_c_1026_n 0.0118398f $X=2.055 $Y=2.7 $X2=0
+ $Y2=0
cc_592 N_A_93_376#_c_924_n N_VPWR_c_1027_n 0.00327848f $X=2.055 $Y=2.7 $X2=0
+ $Y2=0
cc_593 N_A_93_376#_c_917_n N_VPWR_c_1027_n 0.0580227f $X=3.1 $Y=2.875 $X2=0
+ $Y2=0
cc_594 N_A_93_376#_c_920_n N_VPWR_c_1027_n 0.00978294f $X=2.14 $Y=2.7 $X2=0
+ $Y2=0
cc_595 N_A_93_376#_c_916_n N_VPWR_c_1020_n 0.0156198f $X=0.675 $Y=2.615 $X2=0
+ $Y2=0
cc_596 N_A_93_376#_c_924_n N_VPWR_c_1020_n 0.0265795f $X=2.055 $Y=2.7 $X2=0
+ $Y2=0
cc_597 N_A_93_376#_c_917_n N_VPWR_c_1020_n 0.0386722f $X=3.1 $Y=2.875 $X2=0
+ $Y2=0
cc_598 N_A_93_376#_c_920_n N_VPWR_c_1020_n 0.00635315f $X=2.14 $Y=2.7 $X2=0
+ $Y2=0
cc_599 N_A_93_376#_c_924_n N_VPWR_c_1031_n 0.0230277f $X=2.055 $Y=2.7 $X2=0
+ $Y2=0
cc_600 N_A_93_376#_c_920_n N_VPWR_c_1031_n 0.00592055f $X=2.14 $Y=2.7 $X2=0
+ $Y2=0
cc_601 N_A_93_376#_c_909_n N_VGND_c_1140_n 0.019842f $X=1.1 $Y=0.715 $X2=0 $Y2=0
cc_602 N_A_93_376#_c_909_n N_VGND_c_1141_n 0.0130179f $X=1.1 $Y=0.715 $X2=0
+ $Y2=0
cc_603 N_A_93_376#_c_910_n N_VGND_c_1141_n 0.0207154f $X=2.235 $Y=1.125 $X2=0
+ $Y2=0
cc_604 N_A_93_376#_c_911_n N_VGND_c_1141_n 0.0176897f $X=2.32 $Y=1.04 $X2=0
+ $Y2=0
cc_605 N_A_93_376#_c_913_n N_VGND_c_1141_n 0.0141902f $X=2.405 $Y=0.35 $X2=0
+ $Y2=0
cc_606 N_A_93_376#_c_909_n N_VGND_c_1145_n 0.014752f $X=1.1 $Y=0.715 $X2=0 $Y2=0
cc_607 N_A_93_376#_c_912_n N_VGND_c_1149_n 0.0466613f $X=3.175 $Y=0.35 $X2=0
+ $Y2=0
cc_608 N_A_93_376#_c_913_n N_VGND_c_1149_n 0.0114622f $X=2.405 $Y=0.35 $X2=0
+ $Y2=0
cc_609 N_A_93_376#_c_915_n N_VGND_c_1149_n 0.0191504f $X=3.34 $Y=0.35 $X2=0
+ $Y2=0
cc_610 N_A_93_376#_M1013_s N_VGND_c_1152_n 0.00232985f $X=3.195 $Y=0.235 $X2=0
+ $Y2=0
cc_611 N_A_93_376#_c_909_n N_VGND_c_1152_n 0.0176693f $X=1.1 $Y=0.715 $X2=0
+ $Y2=0
cc_612 N_A_93_376#_c_912_n N_VGND_c_1152_n 0.0287732f $X=3.175 $Y=0.35 $X2=0
+ $Y2=0
cc_613 N_A_93_376#_c_913_n N_VGND_c_1152_n 0.00657784f $X=2.405 $Y=0.35 $X2=0
+ $Y2=0
cc_614 N_A_93_376#_c_915_n N_VGND_c_1152_n 0.0124135f $X=3.34 $Y=0.35 $X2=0
+ $Y2=0
cc_615 N_A_93_376#_c_909_n A_114_101# 0.00469244f $X=1.1 $Y=0.715 $X2=-0.19
+ $Y2=-0.245
cc_616 N_VPWR_c_1029_n GCLK 0.0244777f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_617 N_VPWR_c_1020_n GCLK 0.015279f $X=8.4 $Y=3.33 $X2=0 $Y2=0
cc_618 GCLK N_VGND_c_1144_n 0.0108399f $X=8.315 $Y=0.47 $X2=0 $Y2=0
cc_619 GCLK N_VGND_c_1151_n 0.0258562f $X=8.315 $Y=0.47 $X2=0 $Y2=0
cc_620 N_GCLK_M1005_d N_VGND_c_1152_n 0.00228036f $X=8.1 $Y=0.24 $X2=0 $Y2=0
cc_621 GCLK N_VGND_c_1152_n 0.0165126f $X=8.315 $Y=0.47 $X2=0 $Y2=0
cc_622 N_VGND_c_1152_n A_812_47# 0.010279f $X=8.4 $Y=0 $X2=-0.19 $Y2=-0.245
cc_623 N_VGND_c_1152_n A_1016_47# 0.00486245f $X=8.4 $Y=0 $X2=-0.19 $Y2=-0.245
cc_624 N_VGND_c_1152_n A_1548_48# 0.00392312f $X=8.4 $Y=0 $X2=-0.19 $Y2=-0.245
