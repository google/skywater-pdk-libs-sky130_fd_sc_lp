* File: sky130_fd_sc_lp__o22a_lp.pxi.spice
* Created: Fri Aug 28 11:10:02 2020
* 
x_PM_SKY130_FD_SC_LP__O22A_LP%A1 N_A1_c_66_n N_A1_M1008_g N_A1_M1007_g A1
+ N_A1_c_68_n PM_SKY130_FD_SC_LP__O22A_LP%A1
x_PM_SKY130_FD_SC_LP__O22A_LP%A2 N_A2_c_94_n N_A2_M1001_g N_A2_M1004_g A2
+ N_A2_c_97_n PM_SKY130_FD_SC_LP__O22A_LP%A2
x_PM_SKY130_FD_SC_LP__O22A_LP%B2 N_B2_M1005_g N_B2_M1006_g N_B2_c_137_n B2 B2 B2
+ N_B2_c_139_n PM_SKY130_FD_SC_LP__O22A_LP%B2
x_PM_SKY130_FD_SC_LP__O22A_LP%B1 N_B1_M1003_g N_B1_M1009_g B1 N_B1_c_185_n
+ PM_SKY130_FD_SC_LP__O22A_LP%B1
x_PM_SKY130_FD_SC_LP__O22A_LP%A_232_419# N_A_232_419#_M1005_d
+ N_A_232_419#_M1001_d N_A_232_419#_M1010_g N_A_232_419#_M1002_g
+ N_A_232_419#_M1000_g N_A_232_419#_c_219_n N_A_232_419#_c_220_n
+ N_A_232_419#_c_239_n N_A_232_419#_c_221_n N_A_232_419#_c_233_n
+ N_A_232_419#_c_227_n N_A_232_419#_c_222_n N_A_232_419#_c_223_n
+ N_A_232_419#_c_224_n N_A_232_419#_c_229_n N_A_232_419#_c_237_n
+ N_A_232_419#_c_260_n PM_SKY130_FD_SC_LP__O22A_LP%A_232_419#
x_PM_SKY130_FD_SC_LP__O22A_LP%VPWR N_VPWR_M1008_s N_VPWR_M1009_d N_VPWR_c_298_n
+ N_VPWR_c_299_n N_VPWR_c_300_n N_VPWR_c_301_n N_VPWR_c_302_n VPWR
+ N_VPWR_c_303_n N_VPWR_c_297_n PM_SKY130_FD_SC_LP__O22A_LP%VPWR
x_PM_SKY130_FD_SC_LP__O22A_LP%X N_X_M1000_d N_X_M1002_d X X X X X X X X
+ PM_SKY130_FD_SC_LP__O22A_LP%X
x_PM_SKY130_FD_SC_LP__O22A_LP%A_30_173# N_A_30_173#_M1007_s N_A_30_173#_M1004_d
+ N_A_30_173#_M1003_d N_A_30_173#_c_362_n N_A_30_173#_c_363_n
+ N_A_30_173#_c_364_n N_A_30_173#_c_374_n N_A_30_173#_c_365_n
+ N_A_30_173#_c_366_n N_A_30_173#_c_367_n PM_SKY130_FD_SC_LP__O22A_LP%A_30_173#
x_PM_SKY130_FD_SC_LP__O22A_LP%VGND N_VGND_M1007_d N_VGND_M1010_s N_VGND_c_409_n
+ N_VGND_c_410_n VGND N_VGND_c_411_n N_VGND_c_412_n N_VGND_c_413_n
+ N_VGND_c_414_n N_VGND_c_415_n N_VGND_c_416_n PM_SKY130_FD_SC_LP__O22A_LP%VGND
cc_1 VNB N_A1_c_66_n 0.0194487f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=2.09
cc_2 VNB N_A1_M1007_g 0.0297238f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.075
cc_3 VNB N_A1_c_68_n 0.00495072f $X=-0.19 $Y=-0.245 $X2=0.45 $Y2=1.67
cc_4 VNB N_A2_c_94_n 0.0210239f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=2.09
cc_5 VNB N_A2_M1001_g 0.00252117f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=2.595
cc_6 VNB N_A2_M1004_g 0.0227159f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_A2_c_97_n 0.00415811f $X=-0.19 $Y=-0.245 $X2=0.362 $Y2=1.67
cc_8 VNB N_B2_M1005_g 0.0312581f $X=-0.19 $Y=-0.245 $X2=0.51 $Y2=1.49
cc_9 VNB N_B2_M1006_g 0.0107053f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_B2_c_137_n 0.0155202f $X=-0.19 $Y=-0.245 $X2=0.477 $Y2=1.67
cc_11 VNB B2 0.0296301f $X=-0.19 $Y=-0.245 $X2=0.362 $Y2=1.67
cc_12 VNB N_B2_c_139_n 0.0441679f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_B1_M1003_g 0.0289749f $X=-0.19 $Y=-0.245 $X2=0.545 $Y2=2.595
cc_14 VNB N_B1_M1009_g 0.0107205f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB B1 0.0138638f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_B1_c_185_n 0.0329753f $X=-0.19 $Y=-0.245 $X2=0.362 $Y2=2.035
cc_17 VNB N_A_232_419#_M1010_g 0.0270238f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_232_419#_M1002_g 0.00936211f $X=-0.19 $Y=-0.245 $X2=0.362 $Y2=1.67
cc_19 VNB N_A_232_419#_M1000_g 0.0233013f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_232_419#_c_219_n 0.0233607f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_232_419#_c_220_n 0.026149f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_232_419#_c_221_n 0.00634532f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_232_419#_c_222_n 6.19362e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_232_419#_c_223_n 0.0322071f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_232_419#_c_224_n 9.34566e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_VPWR_c_297_n 0.163682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB X 0.0182758f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB X 0.0500601f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.95
cc_29 VNB N_A_30_173#_c_362_n 0.0203502f $X=-0.19 $Y=-0.245 $X2=0.45 $Y2=1.67
cc_30 VNB N_A_30_173#_c_363_n 0.0119949f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_30_173#_c_364_n 0.00965289f $X=-0.19 $Y=-0.245 $X2=0.362 $Y2=2.035
cc_32 VNB N_A_30_173#_c_365_n 0.00341811f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_30_173#_c_366_n 0.00254323f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_30_173#_c_367_n 0.00950508f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_409_n 0.0373187f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_410_n 0.0119746f $X=-0.19 $Y=-0.245 $X2=0.362 $Y2=1.67
cc_37 VNB N_VGND_c_411_n 0.0204409f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_412_n 0.04429f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_413_n 0.0268694f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_414_n 0.242083f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_415_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_416_n 0.00510939f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VPB N_A1_c_66_n 0.0553968f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=2.09
cc_44 VPB N_A1_c_68_n 0.0198387f $X=-0.19 $Y=1.655 $X2=0.45 $Y2=1.67
cc_45 VPB N_A2_c_94_n 0.00833743f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=2.09
cc_46 VPB N_A2_M1001_g 0.0263938f $X=-0.19 $Y=1.655 $X2=0.545 $Y2=2.595
cc_47 VPB N_A2_c_97_n 0.00319161f $X=-0.19 $Y=1.655 $X2=0.362 $Y2=1.67
cc_48 VPB N_B2_M1006_g 0.0263851f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_49 VPB N_B1_M1009_g 0.0302431f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_50 VPB B1 0.00436383f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_51 VPB N_B1_c_185_n 0.0099238f $X=-0.19 $Y=1.655 $X2=0.362 $Y2=2.035
cc_52 VPB N_A_232_419#_M1002_g 0.0546048f $X=-0.19 $Y=1.655 $X2=0.362 $Y2=1.67
cc_53 VPB N_A_232_419#_c_221_n 4.19001e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_54 VPB N_A_232_419#_c_227_n 0.0139117f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_55 VPB N_A_232_419#_c_224_n 0.00360237f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_56 VPB N_VPWR_c_298_n 0.0108753f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_57 VPB N_VPWR_c_299_n 0.0325875f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_58 VPB N_VPWR_c_300_n 0.00287347f $X=-0.19 $Y=1.655 $X2=0.362 $Y2=1.67
cc_59 VPB N_VPWR_c_301_n 0.0513008f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_60 VPB N_VPWR_c_302_n 0.00513801f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_61 VPB N_VPWR_c_303_n 0.0391528f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_62 VPB N_VPWR_c_297_n 0.0469055f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_63 VPB X 0.0220378f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.95
cc_64 VPB X 0.0167475f $X=-0.19 $Y=1.655 $X2=0.45 $Y2=1.67
cc_65 VPB X 0.0343114f $X=-0.19 $Y=1.655 $X2=0.45 $Y2=1.67
cc_66 N_A1_c_66_n N_A2_c_94_n 0.0217699f $X=0.545 $Y=2.09 $X2=-0.19 $Y2=-0.245
cc_67 N_A1_c_68_n N_A2_c_94_n 8.36272e-19 $X=0.45 $Y=1.67 $X2=-0.19 $Y2=-0.245
cc_68 N_A1_c_66_n N_A2_M1001_g 0.0755139f $X=0.545 $Y=2.09 $X2=0 $Y2=0
cc_69 N_A1_c_68_n N_A2_M1001_g 3.19528e-19 $X=0.45 $Y=1.67 $X2=0 $Y2=0
cc_70 N_A1_M1007_g N_A2_M1004_g 0.0166842f $X=0.51 $Y=1.075 $X2=0 $Y2=0
cc_71 N_A1_c_66_n N_A2_c_97_n 0.00296978f $X=0.545 $Y=2.09 $X2=0 $Y2=0
cc_72 N_A1_c_68_n N_A2_c_97_n 0.0388486f $X=0.45 $Y=1.67 $X2=0 $Y2=0
cc_73 N_A1_c_66_n N_A_232_419#_c_229_n 0.00325465f $X=0.545 $Y=2.09 $X2=0 $Y2=0
cc_74 N_A1_c_68_n N_VPWR_M1008_s 0.00276905f $X=0.45 $Y=1.67 $X2=-0.19
+ $Y2=-0.245
cc_75 N_A1_c_66_n N_VPWR_c_299_n 0.0240068f $X=0.545 $Y=2.09 $X2=0 $Y2=0
cc_76 N_A1_c_68_n N_VPWR_c_299_n 0.0239637f $X=0.45 $Y=1.67 $X2=0 $Y2=0
cc_77 N_A1_c_66_n N_VPWR_c_301_n 0.008763f $X=0.545 $Y=2.09 $X2=0 $Y2=0
cc_78 N_A1_c_66_n N_VPWR_c_297_n 0.0144563f $X=0.545 $Y=2.09 $X2=0 $Y2=0
cc_79 N_A1_M1007_g N_A_30_173#_c_362_n 7.35003e-19 $X=0.51 $Y=1.075 $X2=0 $Y2=0
cc_80 N_A1_c_66_n N_A_30_173#_c_363_n 0.00323663f $X=0.545 $Y=2.09 $X2=0 $Y2=0
cc_81 N_A1_M1007_g N_A_30_173#_c_363_n 0.0163415f $X=0.51 $Y=1.075 $X2=0 $Y2=0
cc_82 N_A1_c_68_n N_A_30_173#_c_363_n 0.0158351f $X=0.45 $Y=1.67 $X2=0 $Y2=0
cc_83 N_A1_c_66_n N_A_30_173#_c_364_n 0.00305593f $X=0.545 $Y=2.09 $X2=0 $Y2=0
cc_84 N_A1_c_68_n N_A_30_173#_c_364_n 0.0244963f $X=0.45 $Y=1.67 $X2=0 $Y2=0
cc_85 N_A1_M1007_g N_A_30_173#_c_374_n 5.20836e-19 $X=0.51 $Y=1.075 $X2=0 $Y2=0
cc_86 N_A1_M1007_g N_VGND_c_409_n 0.00902878f $X=0.51 $Y=1.075 $X2=0 $Y2=0
cc_87 N_A1_M1007_g N_VGND_c_411_n 0.0028751f $X=0.51 $Y=1.075 $X2=0 $Y2=0
cc_88 N_A1_M1007_g N_VGND_c_414_n 0.00383429f $X=0.51 $Y=1.075 $X2=0 $Y2=0
cc_89 N_A2_c_94_n N_B2_M1005_g 0.0123738f $X=1.035 $Y=1.835 $X2=0 $Y2=0
cc_90 N_A2_M1004_g N_B2_M1005_g 0.0180785f $X=1.045 $Y=1.075 $X2=0 $Y2=0
cc_91 N_A2_c_94_n N_B2_M1006_g 0.0321648f $X=1.035 $Y=1.835 $X2=0 $Y2=0
cc_92 N_A2_c_97_n N_B2_M1006_g 0.00418744f $X=0.99 $Y=1.67 $X2=0 $Y2=0
cc_93 N_A2_c_94_n N_B2_c_137_n 5.15389e-19 $X=1.035 $Y=1.835 $X2=0 $Y2=0
cc_94 N_A2_c_97_n N_B2_c_137_n 0.00162694f $X=0.99 $Y=1.67 $X2=0 $Y2=0
cc_95 N_A2_M1004_g B2 0.00112309f $X=1.045 $Y=1.075 $X2=0 $Y2=0
cc_96 N_A2_c_97_n N_A_232_419#_M1001_d 0.00173842f $X=0.99 $Y=1.67 $X2=0 $Y2=0
cc_97 N_A2_c_94_n N_A_232_419#_c_221_n 2.70718e-19 $X=1.035 $Y=1.835 $X2=0 $Y2=0
cc_98 N_A2_c_97_n N_A_232_419#_c_221_n 0.0173975f $X=0.99 $Y=1.67 $X2=0 $Y2=0
cc_99 N_A2_M1001_g N_A_232_419#_c_233_n 6.58757e-19 $X=1.035 $Y=2.595 $X2=0
+ $Y2=0
cc_100 N_A2_c_97_n N_A_232_419#_c_233_n 4.17353e-19 $X=0.99 $Y=1.67 $X2=0 $Y2=0
cc_101 N_A2_M1001_g N_A_232_419#_c_229_n 0.0160831f $X=1.035 $Y=2.595 $X2=0
+ $Y2=0
cc_102 N_A2_c_97_n N_A_232_419#_c_229_n 0.01199f $X=0.99 $Y=1.67 $X2=0 $Y2=0
cc_103 N_A2_c_97_n N_A_232_419#_c_237_n 0.00842429f $X=0.99 $Y=1.67 $X2=0 $Y2=0
cc_104 N_A2_M1001_g N_VPWR_c_299_n 0.00429931f $X=1.035 $Y=2.595 $X2=0 $Y2=0
cc_105 N_A2_M1001_g N_VPWR_c_301_n 0.00939541f $X=1.035 $Y=2.595 $X2=0 $Y2=0
cc_106 N_A2_M1001_g N_VPWR_c_297_n 0.0161521f $X=1.035 $Y=2.595 $X2=0 $Y2=0
cc_107 N_A2_c_97_n A_134_419# 0.00160945f $X=0.99 $Y=1.67 $X2=-0.19 $Y2=-0.245
cc_108 N_A2_c_94_n N_A_30_173#_c_363_n 0.00493073f $X=1.035 $Y=1.835 $X2=0 $Y2=0
cc_109 N_A2_M1004_g N_A_30_173#_c_363_n 0.0139305f $X=1.045 $Y=1.075 $X2=0 $Y2=0
cc_110 N_A2_c_97_n N_A_30_173#_c_363_n 0.0415685f $X=0.99 $Y=1.67 $X2=0 $Y2=0
cc_111 N_A2_M1004_g N_A_30_173#_c_374_n 0.00423118f $X=1.045 $Y=1.075 $X2=0
+ $Y2=0
cc_112 N_A2_M1004_g N_A_30_173#_c_366_n 0.00220896f $X=1.045 $Y=1.075 $X2=0
+ $Y2=0
cc_113 N_A2_M1004_g N_VGND_c_409_n 0.00523555f $X=1.045 $Y=1.075 $X2=0 $Y2=0
cc_114 N_A2_M1004_g N_VGND_c_412_n 0.00239141f $X=1.045 $Y=1.075 $X2=0 $Y2=0
cc_115 N_A2_M1004_g N_VGND_c_414_n 0.00312726f $X=1.045 $Y=1.075 $X2=0 $Y2=0
cc_116 N_B2_M1005_g N_B1_M1003_g 0.0191965f $X=1.475 $Y=1.075 $X2=0 $Y2=0
cc_117 B2 N_B1_M1003_g 0.00458954f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_118 N_B2_M1006_g N_B1_M1009_g 0.0335761f $X=1.565 $Y=2.595 $X2=0 $Y2=0
cc_119 N_B2_c_137_n N_B1_c_185_n 0.0335761f $X=1.545 $Y=1.735 $X2=0 $Y2=0
cc_120 B2 N_A_232_419#_M1010_g 0.00209023f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_121 N_B2_M1006_g N_A_232_419#_c_239_n 0.0198602f $X=1.565 $Y=2.595 $X2=0
+ $Y2=0
cc_122 N_B2_M1005_g N_A_232_419#_c_221_n 0.0059562f $X=1.475 $Y=1.075 $X2=0
+ $Y2=0
cc_123 N_B2_M1006_g N_A_232_419#_c_221_n 0.00560487f $X=1.565 $Y=2.595 $X2=0
+ $Y2=0
cc_124 N_B2_c_137_n N_A_232_419#_c_221_n 0.00387297f $X=1.545 $Y=1.735 $X2=0
+ $Y2=0
cc_125 N_B2_M1006_g N_A_232_419#_c_233_n 0.00456218f $X=1.565 $Y=2.595 $X2=0
+ $Y2=0
cc_126 N_B2_M1006_g N_A_232_419#_c_229_n 0.0142731f $X=1.565 $Y=2.595 $X2=0
+ $Y2=0
cc_127 N_B2_M1006_g N_A_232_419#_c_237_n 0.00471591f $X=1.565 $Y=2.595 $X2=0
+ $Y2=0
cc_128 N_B2_M1006_g N_VPWR_c_300_n 0.00357372f $X=1.565 $Y=2.595 $X2=0 $Y2=0
cc_129 N_B2_M1006_g N_VPWR_c_301_n 0.00939541f $X=1.565 $Y=2.595 $X2=0 $Y2=0
cc_130 N_B2_M1006_g N_VPWR_c_297_n 0.00963314f $X=1.565 $Y=2.595 $X2=0 $Y2=0
cc_131 N_B2_M1005_g N_A_30_173#_c_363_n 0.00985339f $X=1.475 $Y=1.075 $X2=0
+ $Y2=0
cc_132 B2 N_A_30_173#_c_363_n 2.89014e-19 $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_133 N_B2_M1005_g N_A_30_173#_c_374_n 0.00536128f $X=1.475 $Y=1.075 $X2=0
+ $Y2=0
cc_134 N_B2_M1005_g N_A_30_173#_c_365_n 0.00599575f $X=1.475 $Y=1.075 $X2=0
+ $Y2=0
cc_135 N_B2_c_137_n N_A_30_173#_c_365_n 0.00308567f $X=1.545 $Y=1.735 $X2=0
+ $Y2=0
cc_136 B2 N_A_30_173#_c_365_n 0.0445379f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_137 N_B2_c_139_n N_A_30_173#_c_365_n 0.00120377f $X=1.565 $Y=0.49 $X2=0 $Y2=0
cc_138 N_B2_M1005_g N_A_30_173#_c_366_n 0.00338062f $X=1.475 $Y=1.075 $X2=0
+ $Y2=0
cc_139 B2 N_A_30_173#_c_366_n 0.0324503f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_140 N_B2_M1005_g N_A_30_173#_c_367_n 6.49093e-19 $X=1.475 $Y=1.075 $X2=0
+ $Y2=0
cc_141 B2 N_A_30_173#_c_367_n 0.0125838f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_142 N_B2_M1005_g N_VGND_c_409_n 0.00195367f $X=1.475 $Y=1.075 $X2=0 $Y2=0
cc_143 B2 N_VGND_c_409_n 0.0291367f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_144 N_B2_c_139_n N_VGND_c_409_n 0.00129136f $X=1.565 $Y=0.49 $X2=0 $Y2=0
cc_145 B2 N_VGND_c_410_n 0.0161204f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_146 B2 N_VGND_c_412_n 0.0549916f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_147 N_B2_c_139_n N_VGND_c_412_n 0.00738902f $X=1.565 $Y=0.49 $X2=0 $Y2=0
cc_148 B2 N_VGND_c_414_n 0.0434008f $X=2.075 $Y=0.47 $X2=0 $Y2=0
cc_149 N_B2_c_139_n N_VGND_c_414_n 0.0107124f $X=1.565 $Y=0.49 $X2=0 $Y2=0
cc_150 B1 N_A_232_419#_M1002_g 9.10511e-19 $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_151 N_B1_c_185_n N_A_232_419#_M1002_g 0.00331134f $X=2.28 $Y=1.615 $X2=0
+ $Y2=0
cc_152 B1 N_A_232_419#_c_220_n 7.3228e-19 $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_153 N_B1_c_185_n N_A_232_419#_c_220_n 0.00157106f $X=2.28 $Y=1.615 $X2=0
+ $Y2=0
cc_154 N_B1_M1009_g N_A_232_419#_c_239_n 0.00182997f $X=2.115 $Y=2.595 $X2=0
+ $Y2=0
cc_155 N_B1_M1003_g N_A_232_419#_c_221_n 0.0130933f $X=2.065 $Y=1.075 $X2=0
+ $Y2=0
cc_156 B1 N_A_232_419#_c_221_n 0.0256895f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_157 N_B1_M1009_g N_A_232_419#_c_233_n 0.0039751f $X=2.115 $Y=2.595 $X2=0
+ $Y2=0
cc_158 N_B1_M1009_g N_A_232_419#_c_227_n 0.0279257f $X=2.115 $Y=2.595 $X2=0
+ $Y2=0
cc_159 B1 N_A_232_419#_c_227_n 0.0468923f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_160 N_B1_c_185_n N_A_232_419#_c_227_n 0.0045667f $X=2.28 $Y=1.615 $X2=0 $Y2=0
cc_161 N_B1_M1009_g N_A_232_419#_c_224_n 0.00379086f $X=2.115 $Y=2.595 $X2=0
+ $Y2=0
cc_162 N_B1_c_185_n N_A_232_419#_c_224_n 5.02332e-19 $X=2.28 $Y=1.615 $X2=0
+ $Y2=0
cc_163 N_B1_M1009_g N_A_232_419#_c_229_n 0.00250591f $X=2.115 $Y=2.595 $X2=0
+ $Y2=0
cc_164 B1 N_A_232_419#_c_260_n 0.0264065f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_165 N_B1_M1009_g N_VPWR_c_300_n 0.0231558f $X=2.115 $Y=2.595 $X2=0 $Y2=0
cc_166 N_B1_M1009_g N_VPWR_c_301_n 0.00895812f $X=2.115 $Y=2.595 $X2=0 $Y2=0
cc_167 N_B1_M1009_g N_VPWR_c_297_n 0.0149261f $X=2.115 $Y=2.595 $X2=0 $Y2=0
cc_168 N_B1_M1003_g N_A_30_173#_c_374_n 6.46858e-19 $X=2.065 $Y=1.075 $X2=0
+ $Y2=0
cc_169 N_B1_M1003_g N_A_30_173#_c_365_n 0.0118287f $X=2.065 $Y=1.075 $X2=0 $Y2=0
cc_170 N_B1_M1003_g N_A_30_173#_c_367_n 0.00649129f $X=2.065 $Y=1.075 $X2=0
+ $Y2=0
cc_171 B1 N_A_30_173#_c_367_n 0.0225878f $X=2.555 $Y=1.58 $X2=0 $Y2=0
cc_172 N_B1_c_185_n N_A_30_173#_c_367_n 0.00716761f $X=2.28 $Y=1.615 $X2=0 $Y2=0
cc_173 N_A_232_419#_c_227_n N_VPWR_M1009_d 0.0213669f $X=2.935 $Y=2.045 $X2=0
+ $Y2=0
cc_174 N_A_232_419#_M1002_g N_VPWR_c_300_n 0.0235096f $X=3.185 $Y=2.595 $X2=0
+ $Y2=0
cc_175 N_A_232_419#_c_239_n N_VPWR_c_300_n 0.00783338f $X=1.685 $Y=2.395 $X2=0
+ $Y2=0
cc_176 N_A_232_419#_c_227_n N_VPWR_c_300_n 0.0209862f $X=2.935 $Y=2.045 $X2=0
+ $Y2=0
cc_177 N_A_232_419#_c_229_n N_VPWR_c_301_n 0.0177952f $X=1.3 $Y=2.475 $X2=0
+ $Y2=0
cc_178 N_A_232_419#_M1002_g N_VPWR_c_303_n 0.00939541f $X=3.185 $Y=2.595 $X2=0
+ $Y2=0
cc_179 N_A_232_419#_M1001_d N_VPWR_c_297_n 0.00223819f $X=1.16 $Y=2.095 $X2=0
+ $Y2=0
cc_180 N_A_232_419#_M1002_g N_VPWR_c_297_n 0.0186591f $X=3.185 $Y=2.595 $X2=0
+ $Y2=0
cc_181 N_A_232_419#_c_239_n N_VPWR_c_297_n 0.01253f $X=1.685 $Y=2.395 $X2=0
+ $Y2=0
cc_182 N_A_232_419#_c_229_n N_VPWR_c_297_n 0.0123247f $X=1.3 $Y=2.475 $X2=0
+ $Y2=0
cc_183 N_A_232_419#_c_239_n A_338_419# 0.00460496f $X=1.685 $Y=2.395 $X2=-0.19
+ $Y2=-0.245
cc_184 N_A_232_419#_c_233_n A_338_419# 0.00202076f $X=1.77 $Y=2.31 $X2=-0.19
+ $Y2=-0.245
cc_185 N_A_232_419#_c_237_n A_338_419# 0.00351862f $X=1.81 $Y=2.045 $X2=-0.19
+ $Y2=-0.245
cc_186 N_A_232_419#_M1010_g X 0.00125358f $X=2.985 $Y=0.445 $X2=0 $Y2=0
cc_187 N_A_232_419#_M1000_g X 0.00848459f $X=3.345 $Y=0.445 $X2=0 $Y2=0
cc_188 N_A_232_419#_M1000_g X 0.0114743f $X=3.345 $Y=0.445 $X2=0 $Y2=0
cc_189 N_A_232_419#_c_227_n X 0.0051207f $X=2.935 $Y=2.045 $X2=0 $Y2=0
cc_190 N_A_232_419#_c_222_n X 0.0425408f $X=3.1 $Y=1.02 $X2=0 $Y2=0
cc_191 N_A_232_419#_c_223_n X 0.0254518f $X=3.1 $Y=1.02 $X2=0 $Y2=0
cc_192 N_A_232_419#_c_224_n X 0.0175506f $X=3.02 $Y=1.96 $X2=0 $Y2=0
cc_193 N_A_232_419#_M1002_g X 0.0101731f $X=3.185 $Y=2.595 $X2=0 $Y2=0
cc_194 N_A_232_419#_c_227_n X 0.0042816f $X=2.935 $Y=2.045 $X2=0 $Y2=0
cc_195 N_A_232_419#_M1002_g X 0.0414486f $X=3.185 $Y=2.595 $X2=0 $Y2=0
cc_196 N_A_232_419#_c_221_n N_A_30_173#_c_363_n 0.0131328f $X=1.77 $Y=1.365
+ $X2=0 $Y2=0
cc_197 N_A_232_419#_c_221_n N_A_30_173#_c_374_n 0.00328956f $X=1.77 $Y=1.365
+ $X2=0 $Y2=0
cc_198 N_A_232_419#_M1005_d N_A_30_173#_c_365_n 0.00465811f $X=1.55 $Y=0.865
+ $X2=0 $Y2=0
cc_199 N_A_232_419#_c_221_n N_A_30_173#_c_365_n 0.0192545f $X=1.77 $Y=1.365
+ $X2=0 $Y2=0
cc_200 N_A_232_419#_M1010_g N_A_30_173#_c_367_n 0.0082654f $X=2.985 $Y=0.445
+ $X2=0 $Y2=0
cc_201 N_A_232_419#_c_222_n N_A_30_173#_c_367_n 0.0148595f $X=3.1 $Y=1.02 $X2=0
+ $Y2=0
cc_202 N_A_232_419#_M1010_g N_VGND_c_410_n 0.0133253f $X=2.985 $Y=0.445 $X2=0
+ $Y2=0
cc_203 N_A_232_419#_M1000_g N_VGND_c_410_n 0.00223463f $X=3.345 $Y=0.445 $X2=0
+ $Y2=0
cc_204 N_A_232_419#_M1010_g N_VGND_c_413_n 0.00486043f $X=2.985 $Y=0.445 $X2=0
+ $Y2=0
cc_205 N_A_232_419#_M1000_g N_VGND_c_413_n 0.00549284f $X=3.345 $Y=0.445 $X2=0
+ $Y2=0
cc_206 N_A_232_419#_M1010_g N_VGND_c_414_n 0.00440432f $X=2.985 $Y=0.445 $X2=0
+ $Y2=0
cc_207 N_A_232_419#_M1000_g N_VGND_c_414_n 0.010905f $X=3.345 $Y=0.445 $X2=0
+ $Y2=0
cc_208 N_A_232_419#_c_222_n N_VGND_c_414_n 0.0110078f $X=3.1 $Y=1.02 $X2=0 $Y2=0
cc_209 N_VPWR_c_297_n A_134_419# 0.010279f $X=3.6 $Y=3.33 $X2=-0.19 $Y2=-0.245
cc_210 N_VPWR_c_297_n A_338_419# 0.00822544f $X=3.6 $Y=3.33 $X2=-0.19 $Y2=-0.245
cc_211 N_VPWR_c_297_n N_X_M1002_d 0.0023218f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_212 N_VPWR_c_303_n X 0.0271747f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_213 N_VPWR_c_297_n X 0.0167643f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_214 X N_VGND_c_410_n 0.0117101f $X=3.515 $Y=0.47 $X2=0 $Y2=0
cc_215 X N_VGND_c_413_n 0.0197155f $X=3.515 $Y=0.47 $X2=0 $Y2=0
cc_216 N_X_M1000_d N_VGND_c_414_n 0.00232985f $X=3.42 $Y=0.235 $X2=0 $Y2=0
cc_217 X N_VGND_c_414_n 0.0125355f $X=3.515 $Y=0.47 $X2=0 $Y2=0
cc_218 N_A_30_173#_c_363_n N_VGND_M1007_d 0.00318248f $X=1.095 $Y=1.33 $X2=-0.19
+ $Y2=-0.245
cc_219 N_A_30_173#_c_362_n N_VGND_c_409_n 0.00900914f $X=0.295 $Y=1.03 $X2=0
+ $Y2=0
cc_220 N_A_30_173#_c_363_n N_VGND_c_409_n 0.0219594f $X=1.095 $Y=1.33 $X2=0
+ $Y2=0
cc_221 N_A_30_173#_c_374_n N_VGND_c_409_n 0.00394685f $X=1.26 $Y=1.03 $X2=0
+ $Y2=0
cc_222 N_A_30_173#_c_366_n N_VGND_c_409_n 0.0128719f $X=1.505 $Y=0.935 $X2=0
+ $Y2=0
cc_223 N_A_30_173#_c_362_n N_VGND_c_414_n 0.010476f $X=0.295 $Y=1.03 $X2=0 $Y2=0
cc_224 N_A_30_173#_c_367_n N_VGND_c_414_n 0.00657009f $X=2.28 $Y=0.935 $X2=0
+ $Y2=0
cc_225 N_VGND_c_414_n A_612_47# 0.00329326f $X=3.6 $Y=0 $X2=-0.19 $Y2=-0.245
