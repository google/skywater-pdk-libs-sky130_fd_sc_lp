* File: sky130_fd_sc_lp__o31a_2.pex.spice
* Created: Wed Sep  2 10:24:37 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O31A_2%A_85_21# 1 2 7 9 12 14 16 19 23 24 27 28 32
+ 36 38 40 41 43 44
r100 51 52 6.12014 $w=3.3e-07 $l=3.5e-08 $layer=POLY_cond $X=0.93 $Y=1.35
+ $X2=0.965 $Y2=1.35
r101 50 51 69.0702 $w=3.3e-07 $l=3.95e-07 $layer=POLY_cond $X=0.535 $Y=1.35
+ $X2=0.93 $Y2=1.35
r102 48 50 6.12014 $w=3.3e-07 $l=3.5e-08 $layer=POLY_cond $X=0.5 $Y=1.35
+ $X2=0.535 $Y2=1.35
r103 43 44 8.71334 $w=4.13e-07 $l=1.65e-07 $layer=LI1_cond $X=2.917 $Y=2.095
+ $X2=2.917 $Y2=1.93
r104 40 41 9.42727 $w=1.98e-07 $l=1.7e-07 $layer=LI1_cond $X=1.76 $Y=1.105
+ $X2=1.93 $Y2=1.105
r105 36 45 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=3.39 $Y=1.09
+ $X2=3.04 $Y2=1.09
r106 36 38 25.93 $w=2.58e-07 $l=5.85e-07 $layer=LI1_cond $X=3.39 $Y=1.005
+ $X2=3.39 $Y2=0.42
r107 34 45 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.04 $Y=1.175
+ $X2=3.04 $Y2=1.09
r108 34 44 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=3.04 $Y=1.175
+ $X2=3.04 $Y2=1.93
r109 30 43 1.16633 $w=4.13e-07 $l=4.2e-08 $layer=LI1_cond $X=2.917 $Y=2.137
+ $X2=2.917 $Y2=2.095
r110 30 32 21.466 $w=4.13e-07 $l=7.73e-07 $layer=LI1_cond $X=2.917 $Y=2.137
+ $X2=2.917 $Y2=2.91
r111 28 45 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=2.955 $Y=1.09
+ $X2=3.04 $Y2=1.09
r112 28 41 66.8717 $w=1.68e-07 $l=1.025e-06 $layer=LI1_cond $X=2.955 $Y=1.09
+ $X2=1.93 $Y2=1.09
r113 27 40 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=1.235 $Y=1.12
+ $X2=1.76 $Y2=1.12
r114 24 52 18.3604 $w=3.3e-07 $l=1.05e-07 $layer=POLY_cond $X=1.07 $Y=1.35
+ $X2=0.965 $Y2=1.35
r115 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.07
+ $Y=1.35 $X2=1.07 $Y2=1.35
r116 21 27 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.11 $Y=1.205
+ $X2=1.235 $Y2=1.12
r117 21 23 6.68417 $w=2.48e-07 $l=1.45e-07 $layer=LI1_cond $X=1.11 $Y=1.205
+ $X2=1.11 $Y2=1.35
r118 17 52 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.965 $Y=1.515
+ $X2=0.965 $Y2=1.35
r119 17 19 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=0.965 $Y=1.515
+ $X2=0.965 $Y2=2.465
r120 14 51 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.93 $Y=1.185
+ $X2=0.93 $Y2=1.35
r121 14 16 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.93 $Y=1.185
+ $X2=0.93 $Y2=0.655
r122 10 50 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.535 $Y=1.515
+ $X2=0.535 $Y2=1.35
r123 10 12 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=0.535 $Y=1.515
+ $X2=0.535 $Y2=2.465
r124 7 48 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.5 $Y=1.185
+ $X2=0.5 $Y2=1.35
r125 7 9 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.5 $Y=1.185 $X2=0.5
+ $Y2=0.655
r126 2 43 400 $w=1.7e-07 $l=3.45832e-07 $layer=licon1_PDIFF $count=1 $X=2.675
+ $Y=1.835 $X2=2.875 $Y2=2.095
r127 2 32 400 $w=1.7e-07 $l=1.17074e-06 $layer=licon1_PDIFF $count=1 $X=2.675
+ $Y=1.835 $X2=2.875 $Y2=2.91
r128 1 38 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=3.215
+ $Y=0.235 $X2=3.355 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__O31A_2%A1 3 7 9 10 11 12 19 20 36
r44 36 37 0.881781 $w=3.68e-07 $l=1e-08 $layer=LI1_cond $X=1.63 $Y=1.665
+ $X2=1.63 $Y2=1.675
r45 19 22 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.61 $Y=1.51
+ $X2=1.61 $Y2=1.675
r46 19 21 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.61 $Y=1.51
+ $X2=1.61 $Y2=1.345
r47 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.61
+ $Y=1.51 $X2=1.61 $Y2=1.51
r48 11 12 14.7036 $w=2.88e-07 $l=3.7e-07 $layer=LI1_cond $X=1.67 $Y=2.405
+ $X2=1.67 $Y2=2.775
r49 10 11 14.7036 $w=2.88e-07 $l=3.7e-07 $layer=LI1_cond $X=1.67 $Y=2.035
+ $X2=1.67 $Y2=2.405
r50 9 36 1.18359 $w=3.68e-07 $l=3.8e-08 $layer=LI1_cond $X=1.63 $Y=1.627
+ $X2=1.63 $Y2=1.665
r51 9 20 3.64421 $w=3.68e-07 $l=1.17e-07 $layer=LI1_cond $X=1.63 $Y=1.627
+ $X2=1.63 $Y2=1.51
r52 9 10 12.8358 $w=2.88e-07 $l=3.23e-07 $layer=LI1_cond $X=1.67 $Y=1.712
+ $X2=1.67 $Y2=2.035
r53 9 37 1.47036 $w=2.88e-07 $l=3.7e-08 $layer=LI1_cond $X=1.67 $Y=1.712
+ $X2=1.67 $Y2=1.675
r54 7 22 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.7 $Y=2.465 $X2=1.7
+ $Y2=1.675
r55 3 21 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.7 $Y=0.655 $X2=1.7
+ $Y2=1.345
.ends

.subckt PM_SKY130_FD_SC_LP__O31A_2%A2 3 7 9 10 11 12 18 19
c33 3 0 7.37998e-20 $X=2.06 $Y=2.465
r34 18 21 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.15 $Y=1.51
+ $X2=2.15 $Y2=1.675
r35 18 20 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.15 $Y=1.51
+ $X2=2.15 $Y2=1.345
r36 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.15
+ $Y=1.51 $X2=2.15 $Y2=1.51
r37 11 12 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=2.15 $Y=2.405
+ $X2=2.15 $Y2=2.775
r38 10 11 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=2.15 $Y=2.035
+ $X2=2.15 $Y2=2.405
r39 9 10 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=2.15 $Y=1.665
+ $X2=2.15 $Y2=2.035
r40 9 19 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=2.15 $Y=1.665
+ $X2=2.15 $Y2=1.51
r41 7 20 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.21 $Y=0.655
+ $X2=2.21 $Y2=1.345
r42 3 21 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.06 $Y=2.465
+ $X2=2.06 $Y2=1.675
.ends

.subckt PM_SKY130_FD_SC_LP__O31A_2%A3 3 7 9 12 13
c33 13 0 7.37998e-20 $X=2.69 $Y=1.51
r34 12 15 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.69 $Y=1.51
+ $X2=2.69 $Y2=1.675
r35 12 14 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.69 $Y=1.51
+ $X2=2.69 $Y2=1.345
r36 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.69
+ $Y=1.51 $X2=2.69 $Y2=1.51
r37 9 13 6.87033 $w=2.58e-07 $l=1.55e-07 $layer=LI1_cond $X=2.655 $Y=1.665
+ $X2=2.655 $Y2=1.51
r38 7 14 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.64 $Y=0.655
+ $X2=2.64 $Y2=1.345
r39 3 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.6 $Y=2.465 $X2=2.6
+ $Y2=1.675
.ends

.subckt PM_SKY130_FD_SC_LP__O31A_2%B1 3 7 9 14
r30 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.39
+ $Y=1.51 $X2=3.39 $Y2=1.51
r31 11 14 43.7153 $w=3.3e-07 $l=2.5e-07 $layer=POLY_cond $X=3.14 $Y=1.51
+ $X2=3.39 $Y2=1.51
r32 9 15 5.97563 $w=4.03e-07 $l=2.1e-07 $layer=LI1_cond $X=3.6 $Y=1.547 $X2=3.39
+ $Y2=1.547
r33 5 11 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.14 $Y=1.675
+ $X2=3.14 $Y2=1.51
r34 5 7 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.14 $Y=1.675 $X2=3.14
+ $Y2=2.465
r35 1 11 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.14 $Y=1.345
+ $X2=3.14 $Y2=1.51
r36 1 3 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.14 $Y=1.345 $X2=3.14
+ $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__O31A_2%VPWR 1 2 3 10 12 18 24 29 30 31 33 46 47 53
r49 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r50 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r51 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r52 44 47 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r53 43 44 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r54 41 54 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r55 40 43 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.68 $Y=3.33
+ $X2=3.12 $Y2=3.33
r56 40 41 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r57 38 53 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.355 $Y=3.33
+ $X2=1.23 $Y2=3.33
r58 38 40 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=1.355 $Y=3.33
+ $X2=1.68 $Y2=3.33
r59 37 54 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r60 37 51 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r61 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r62 34 50 4.1267 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=3.33
+ $X2=0.212 $Y2=3.33
r63 34 36 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.425 $Y=3.33
+ $X2=0.72 $Y2=3.33
r64 33 53 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.105 $Y=3.33
+ $X2=1.23 $Y2=3.33
r65 33 36 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=1.105 $Y=3.33
+ $X2=0.72 $Y2=3.33
r66 31 44 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=3.12 $Y2=3.33
r67 31 41 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=1.68 $Y2=3.33
r68 29 43 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=3.295 $Y=3.33
+ $X2=3.12 $Y2=3.33
r69 29 30 6.36606 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=3.295 $Y=3.33
+ $X2=3.405 $Y2=3.33
r70 28 46 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=3.515 $Y=3.33
+ $X2=3.6 $Y2=3.33
r71 28 30 6.36606 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=3.515 $Y=3.33
+ $X2=3.405 $Y2=3.33
r72 24 27 45.312 $w=2.18e-07 $l=8.65e-07 $layer=LI1_cond $X=3.405 $Y=2.085
+ $X2=3.405 $Y2=2.95
r73 22 30 0.432806 $w=2.2e-07 $l=8.5e-08 $layer=LI1_cond $X=3.405 $Y=3.245
+ $X2=3.405 $Y2=3.33
r74 22 27 15.4532 $w=2.18e-07 $l=2.95e-07 $layer=LI1_cond $X=3.405 $Y=3.245
+ $X2=3.405 $Y2=2.95
r75 18 21 44.4843 $w=2.48e-07 $l=9.65e-07 $layer=LI1_cond $X=1.23 $Y=1.985
+ $X2=1.23 $Y2=2.95
r76 16 53 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.23 $Y=3.245
+ $X2=1.23 $Y2=3.33
r77 16 21 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=1.23 $Y=3.245
+ $X2=1.23 $Y2=2.95
r78 12 15 41.4026 $w=2.68e-07 $l=9.7e-07 $layer=LI1_cond $X=0.29 $Y=1.98
+ $X2=0.29 $Y2=2.95
r79 10 50 3.15799 $w=2.7e-07 $l=1.17707e-07 $layer=LI1_cond $X=0.29 $Y=3.245
+ $X2=0.212 $Y2=3.33
r80 10 15 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.29 $Y=3.245
+ $X2=0.29 $Y2=2.95
r81 3 27 400 $w=1.7e-07 $l=1.19465e-06 $layer=licon1_PDIFF $count=1 $X=3.215
+ $Y=1.835 $X2=3.38 $Y2=2.95
r82 3 24 400 $w=1.7e-07 $l=3.22102e-07 $layer=licon1_PDIFF $count=1 $X=3.215
+ $Y=1.835 $X2=3.38 $Y2=2.085
r83 2 21 400 $w=1.7e-07 $l=1.22461e-06 $layer=licon1_PDIFF $count=1 $X=1.04
+ $Y=1.835 $X2=1.27 $Y2=2.95
r84 2 18 400 $w=1.7e-07 $l=2.95635e-07 $layer=licon1_PDIFF $count=1 $X=1.04
+ $Y=1.835 $X2=1.27 $Y2=1.985
r85 1 15 400 $w=1.7e-07 $l=1.17584e-06 $layer=licon1_PDIFF $count=1 $X=0.195
+ $Y=1.835 $X2=0.32 $Y2=2.95
r86 1 12 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.195
+ $Y=1.835 $X2=0.32 $Y2=1.98
.ends

.subckt PM_SKY130_FD_SC_LP__O31A_2%X 1 2 7 8 9 10 11 12 13 24 34
r25 34 47 1.57151 $w=2.18e-07 $l=3e-08 $layer=LI1_cond $X=0.705 $Y=1.665
+ $X2=0.705 $Y2=1.695
r26 13 44 4.86187 $w=3.18e-07 $l=1.35e-07 $layer=LI1_cond $X=0.755 $Y=2.775
+ $X2=0.755 $Y2=2.91
r27 12 13 13.3251 $w=3.18e-07 $l=3.7e-07 $layer=LI1_cond $X=0.755 $Y=2.405
+ $X2=0.755 $Y2=2.775
r28 11 12 15.3059 $w=3.18e-07 $l=4.25e-07 $layer=LI1_cond $X=0.755 $Y=1.98
+ $X2=0.755 $Y2=2.405
r29 11 35 4.50173 $w=3.18e-07 $l=1.25e-07 $layer=LI1_cond $X=0.755 $Y=1.98
+ $X2=0.755 $Y2=1.855
r30 10 35 4.78984 $w=3.18e-07 $l=1.33e-07 $layer=LI1_cond $X=0.755 $Y=1.722
+ $X2=0.755 $Y2=1.855
r31 10 47 2.10712 $w=3.18e-07 $l=2.7e-08 $layer=LI1_cond $X=0.755 $Y=1.722
+ $X2=0.755 $Y2=1.695
r32 10 34 1.46675 $w=2.18e-07 $l=2.8e-08 $layer=LI1_cond $X=0.705 $Y=1.637
+ $X2=0.705 $Y2=1.665
r33 9 10 17.9153 $w=2.18e-07 $l=3.42e-07 $layer=LI1_cond $X=0.705 $Y=1.295
+ $X2=0.705 $Y2=1.637
r34 8 9 19.382 $w=2.18e-07 $l=3.7e-07 $layer=LI1_cond $X=0.705 $Y=0.925
+ $X2=0.705 $Y2=1.295
r35 7 8 19.382 $w=2.18e-07 $l=3.7e-07 $layer=LI1_cond $X=0.705 $Y=0.555
+ $X2=0.705 $Y2=0.925
r36 7 24 7.07181 $w=2.18e-07 $l=1.35e-07 $layer=LI1_cond $X=0.705 $Y=0.555
+ $X2=0.705 $Y2=0.42
r37 2 44 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=0.61
+ $Y=1.835 $X2=0.75 $Y2=2.91
r38 2 11 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.61
+ $Y=1.835 $X2=0.75 $Y2=1.98
r39 1 24 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=0.575
+ $Y=0.235 $X2=0.715 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__O31A_2%VGND 1 2 3 10 12 16 20 23 24 25 27 40 41 47
r54 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r55 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r56 40 41 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r57 38 41 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r58 37 40 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r59 37 38 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r60 35 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r61 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r62 32 47 12.6176 $w=1.7e-07 $l=3.03e-07 $layer=LI1_cond $X=1.59 $Y=0 $X2=1.287
+ $Y2=0
r63 32 34 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=1.59 $Y=0 $X2=2.16
+ $Y2=0
r64 31 48 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r65 31 45 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r66 30 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r67 28 44 4.22672 $w=1.7e-07 $l=1.98e-07 $layer=LI1_cond $X=0.395 $Y=0 $X2=0.197
+ $Y2=0
r68 28 30 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.395 $Y=0 $X2=0.72
+ $Y2=0
r69 27 47 12.6176 $w=1.7e-07 $l=3.02e-07 $layer=LI1_cond $X=0.985 $Y=0 $X2=1.287
+ $Y2=0
r70 27 30 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.985 $Y=0 $X2=0.72
+ $Y2=0
r71 25 35 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=2.16
+ $Y2=0
r72 25 48 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=1.2
+ $Y2=0
r73 23 34 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=2.26 $Y=0 $X2=2.16
+ $Y2=0
r74 23 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.26 $Y=0 $X2=2.425
+ $Y2=0
r75 22 37 3.26203 $w=1.68e-07 $l=5e-08 $layer=LI1_cond $X=2.59 $Y=0 $X2=2.64
+ $Y2=0
r76 22 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.59 $Y=0 $X2=2.425
+ $Y2=0
r77 18 24 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.425 $Y=0.085
+ $X2=2.425 $Y2=0
r78 18 20 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=2.425 $Y=0.085
+ $X2=2.425 $Y2=0.37
r79 14 47 2.53987 $w=6.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.287 $Y=0.085
+ $X2=1.287 $Y2=0
r80 14 16 5.43672 $w=6.03e-07 $l=2.75e-07 $layer=LI1_cond $X=1.287 $Y=0.085
+ $X2=1.287 $Y2=0.36
r81 10 44 3.09532 $w=2.75e-07 $l=1.11018e-07 $layer=LI1_cond $X=0.257 $Y=0.085
+ $X2=0.197 $Y2=0
r82 10 12 12.3626 $w=2.73e-07 $l=2.95e-07 $layer=LI1_cond $X=0.257 $Y=0.085
+ $X2=0.257 $Y2=0.38
r83 3 20 182 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_NDIFF $count=1 $X=2.285
+ $Y=0.235 $X2=2.425 $Y2=0.37
r84 2 16 45.5 $w=1.7e-07 $l=5.38888e-07 $layer=licon1_NDIFF $count=4 $X=1.005
+ $Y=0.235 $X2=1.485 $Y2=0.36
r85 1 12 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.16
+ $Y=0.235 $X2=0.285 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_LP__O31A_2%A_355_47# 1 2 7 9 11 13 15
r24 13 20 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.925 $Y=0.665
+ $X2=2.925 $Y2=0.75
r25 13 15 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.925 $Y=0.665
+ $X2=2.925 $Y2=0.37
r26 12 18 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.09 $Y=0.75
+ $X2=1.925 $Y2=0.75
r27 11 20 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.76 $Y=0.75
+ $X2=2.925 $Y2=0.75
r28 11 12 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.76 $Y=0.75
+ $X2=2.09 $Y2=0.75
r29 7 18 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.925 $Y=0.665
+ $X2=1.925 $Y2=0.75
r30 7 9 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.925 $Y=0.665
+ $X2=1.925 $Y2=0.37
r31 2 20 182 $w=1.7e-07 $l=6.11044e-07 $layer=licon1_NDIFF $count=1 $X=2.715
+ $Y=0.235 $X2=2.925 $Y2=0.75
r32 2 15 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=2.715
+ $Y=0.235 $X2=2.925 $Y2=0.37
r33 1 18 182 $w=1.7e-07 $l=5.85214e-07 $layer=licon1_NDIFF $count=1 $X=1.775
+ $Y=0.235 $X2=1.925 $Y2=0.75
r34 1 9 182 $w=1.7e-07 $l=2.06761e-07 $layer=licon1_NDIFF $count=1 $X=1.775
+ $Y=0.235 $X2=1.925 $Y2=0.37
.ends

