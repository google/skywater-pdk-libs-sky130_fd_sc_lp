* File: sky130_fd_sc_lp__sdfbbn_1.pxi.spice
* Created: Wed Sep  2 10:33:42 2020
* 
x_PM_SKY130_FD_SC_LP__SDFBBN_1%SCD N_SCD_c_349_n N_SCD_M1024_g N_SCD_M1032_g
+ N_SCD_c_355_n SCD N_SCD_c_351_n N_SCD_c_352_n PM_SKY130_FD_SC_LP__SDFBBN_1%SCD
x_PM_SKY130_FD_SC_LP__SDFBBN_1%D N_D_M1046_g N_D_M1007_g N_D_c_382_n D D D
+ N_D_c_384_n PM_SKY130_FD_SC_LP__SDFBBN_1%D
x_PM_SKY130_FD_SC_LP__SDFBBN_1%A_328_429# N_A_328_429#_M1010_d
+ N_A_328_429#_M1047_d N_A_328_429#_c_439_n N_A_328_429#_M1031_g
+ N_A_328_429#_c_440_n N_A_328_429#_c_441_n N_A_328_429#_M1013_g
+ N_A_328_429#_c_431_n N_A_328_429#_c_432_n N_A_328_429#_c_433_n
+ N_A_328_429#_c_434_n N_A_328_429#_c_435_n N_A_328_429#_c_436_n
+ N_A_328_429#_c_437_n N_A_328_429#_c_438_n
+ PM_SKY130_FD_SC_LP__SDFBBN_1%A_328_429#
x_PM_SKY130_FD_SC_LP__SDFBBN_1%SCE N_SCE_M1012_g N_SCE_M1042_g N_SCE_c_505_n
+ N_SCE_c_506_n N_SCE_M1010_g N_SCE_M1047_g SCE N_SCE_c_508_n N_SCE_c_509_n
+ PM_SKY130_FD_SC_LP__SDFBBN_1%SCE
x_PM_SKY130_FD_SC_LP__SDFBBN_1%CLK_N N_CLK_N_M1015_g N_CLK_N_c_569_n
+ N_CLK_N_c_575_n N_CLK_N_M1029_g N_CLK_N_c_570_n N_CLK_N_c_571_n
+ N_CLK_N_c_576_n CLK_N N_CLK_N_c_572_n N_CLK_N_c_573_n
+ PM_SKY130_FD_SC_LP__SDFBBN_1%CLK_N
x_PM_SKY130_FD_SC_LP__SDFBBN_1%A_838_50# N_A_838_50#_M1015_d N_A_838_50#_M1029_d
+ N_A_838_50#_M1039_g N_A_838_50#_M1018_g N_A_838_50#_c_619_n
+ N_A_838_50#_c_620_n N_A_838_50#_c_641_n N_A_838_50#_c_642_n
+ N_A_838_50#_M1033_g N_A_838_50#_M1028_g N_A_838_50#_M1016_g
+ N_A_838_50#_c_644_n N_A_838_50#_M1026_g N_A_838_50#_c_622_n
+ N_A_838_50#_c_623_n N_A_838_50#_c_645_n N_A_838_50#_c_624_n
+ N_A_838_50#_c_625_n N_A_838_50#_c_626_n N_A_838_50#_c_627_n
+ N_A_838_50#_c_673_p N_A_838_50#_c_705_p N_A_838_50#_c_674_p
+ N_A_838_50#_c_628_n N_A_838_50#_c_629_n N_A_838_50#_c_630_n
+ N_A_838_50#_c_631_n N_A_838_50#_c_632_n N_A_838_50#_c_633_n
+ N_A_838_50#_c_648_n N_A_838_50#_c_649_n N_A_838_50#_c_650_n
+ N_A_838_50#_c_651_n N_A_838_50#_c_652_n N_A_838_50#_c_634_n
+ N_A_838_50#_c_635_n N_A_838_50#_c_636_n N_A_838_50#_c_637_n
+ N_A_838_50#_c_638_n N_A_838_50#_c_639_n PM_SKY130_FD_SC_LP__SDFBBN_1%A_838_50#
x_PM_SKY130_FD_SC_LP__SDFBBN_1%A_1445_324# N_A_1445_324#_M1000_d
+ N_A_1445_324#_M1030_d N_A_1445_324#_c_877_n N_A_1445_324#_M1009_g
+ N_A_1445_324#_c_866_n N_A_1445_324#_M1040_g N_A_1445_324#_M1027_g
+ N_A_1445_324#_M1043_g N_A_1445_324#_c_869_n N_A_1445_324#_c_870_n
+ N_A_1445_324#_c_912_p N_A_1445_324#_c_940_p N_A_1445_324#_c_871_n
+ N_A_1445_324#_c_882_n N_A_1445_324#_c_872_n N_A_1445_324#_c_873_n
+ N_A_1445_324#_c_874_n N_A_1445_324#_c_885_n N_A_1445_324#_c_875_n
+ N_A_1445_324#_c_876_n PM_SKY130_FD_SC_LP__SDFBBN_1%A_1445_324#
x_PM_SKY130_FD_SC_LP__SDFBBN_1%SET_B N_SET_B_M1035_g N_SET_B_M1030_g
+ N_SET_B_M1022_g N_SET_B_c_1017_n N_SET_B_M1011_g N_SET_B_c_1019_n SET_B
+ N_SET_B_c_1008_n N_SET_B_c_1009_n N_SET_B_c_1010_n N_SET_B_c_1011_n
+ N_SET_B_c_1012_n N_SET_B_c_1013_n N_SET_B_c_1014_n N_SET_B_c_1015_n
+ PM_SKY130_FD_SC_LP__SDFBBN_1%SET_B
x_PM_SKY130_FD_SC_LP__SDFBBN_1%A_1295_379# N_A_1295_379#_M1005_d
+ N_A_1295_379#_M1033_d N_A_1295_379#_M1000_g N_A_1295_379#_c_1147_n
+ N_A_1295_379#_c_1148_n N_A_1295_379#_M1001_g N_A_1295_379#_c_1149_n
+ N_A_1295_379#_c_1161_n N_A_1295_379#_c_1150_n N_A_1295_379#_c_1151_n
+ N_A_1295_379#_c_1152_n N_A_1295_379#_c_1153_n N_A_1295_379#_c_1154_n
+ N_A_1295_379#_c_1155_n N_A_1295_379#_c_1165_n N_A_1295_379#_c_1156_n
+ PM_SKY130_FD_SC_LP__SDFBBN_1%A_1295_379#
x_PM_SKY130_FD_SC_LP__SDFBBN_1%A_995_66# N_A_995_66#_M1039_s N_A_995_66#_M1018_s
+ N_A_995_66#_c_1275_n N_A_995_66#_M1005_g N_A_995_66#_c_1277_n
+ N_A_995_66#_c_1278_n N_A_995_66#_M1034_g N_A_995_66#_c_1289_n
+ N_A_995_66#_c_1290_n N_A_995_66#_M1038_g N_A_995_66#_c_1292_n
+ N_A_995_66#_c_1293_n N_A_995_66#_c_1279_n N_A_995_66#_c_1280_n
+ N_A_995_66#_M1014_g N_A_995_66#_c_1281_n N_A_995_66#_c_1282_n
+ N_A_995_66#_c_1283_n N_A_995_66#_c_1295_n N_A_995_66#_c_1284_n
+ N_A_995_66#_c_1285_n N_A_995_66#_c_1286_n
+ PM_SKY130_FD_SC_LP__SDFBBN_1%A_995_66#
x_PM_SKY130_FD_SC_LP__SDFBBN_1%A_2449_137# N_A_2449_137#_M1036_d
+ N_A_2449_137#_M1011_d N_A_2449_137#_c_1397_n N_A_2449_137#_M1025_g
+ N_A_2449_137#_c_1398_n N_A_2449_137#_c_1399_n N_A_2449_137#_M1037_g
+ N_A_2449_137#_M1020_g N_A_2449_137#_M1021_g N_A_2449_137#_c_1401_n
+ N_A_2449_137#_c_1402_n N_A_2449_137#_M1002_g N_A_2449_137#_M1041_g
+ N_A_2449_137#_c_1404_n N_A_2449_137#_c_1405_n N_A_2449_137#_c_1406_n
+ N_A_2449_137#_c_1416_n N_A_2449_137#_c_1417_n N_A_2449_137#_c_1453_n
+ N_A_2449_137#_c_1463_p N_A_2449_137#_c_1407_n N_A_2449_137#_c_1408_n
+ N_A_2449_137#_c_1419_n N_A_2449_137#_c_1420_n N_A_2449_137#_c_1454_n
+ N_A_2449_137#_c_1409_n N_A_2449_137#_c_1483_p N_A_2449_137#_c_1410_n
+ N_A_2449_137#_c_1411_n N_A_2449_137#_c_1412_n
+ PM_SKY130_FD_SC_LP__SDFBBN_1%A_2449_137#
x_PM_SKY130_FD_SC_LP__SDFBBN_1%A_2299_119# N_A_2299_119#_M1016_d
+ N_A_2299_119#_M1038_d N_A_2299_119#_M1036_g N_A_2299_119#_M1045_g
+ N_A_2299_119#_c_1615_n N_A_2299_119#_c_1584_n N_A_2299_119#_c_1590_n
+ N_A_2299_119#_c_1585_n N_A_2299_119#_c_1586_n N_A_2299_119#_c_1587_n
+ N_A_2299_119#_c_1588_n PM_SKY130_FD_SC_LP__SDFBBN_1%A_2299_119#
x_PM_SKY130_FD_SC_LP__SDFBBN_1%A_1926_21# N_A_1926_21#_M1006_s
+ N_A_1926_21#_M1019_s N_A_1926_21#_M1008_g N_A_1926_21#_c_1682_n
+ N_A_1926_21#_c_1683_n N_A_1926_21#_c_1684_n N_A_1926_21#_c_1685_n
+ N_A_1926_21#_M1003_g N_A_1926_21#_M1044_g N_A_1926_21#_M1017_g
+ N_A_1926_21#_c_1688_n N_A_1926_21#_c_1689_n N_A_1926_21#_c_1697_n
+ N_A_1926_21#_c_1690_n N_A_1926_21#_c_1691_n N_A_1926_21#_c_1692_n
+ N_A_1926_21#_c_1698_n N_A_1926_21#_c_1699_n N_A_1926_21#_c_1693_n
+ PM_SKY130_FD_SC_LP__SDFBBN_1%A_1926_21#
x_PM_SKY130_FD_SC_LP__SDFBBN_1%RESET_B N_RESET_B_M1019_g N_RESET_B_M1006_g
+ RESET_B N_RESET_B_c_1804_n N_RESET_B_c_1805_n
+ PM_SKY130_FD_SC_LP__SDFBBN_1%RESET_B
x_PM_SKY130_FD_SC_LP__SDFBBN_1%A_3279_367# N_A_3279_367#_M1041_s
+ N_A_3279_367#_M1002_s N_A_3279_367#_M1023_g N_A_3279_367#_M1004_g
+ N_A_3279_367#_c_1843_n N_A_3279_367#_c_1848_n N_A_3279_367#_c_1844_n
+ N_A_3279_367#_c_1845_n N_A_3279_367#_c_1846_n
+ PM_SKY130_FD_SC_LP__SDFBBN_1%A_3279_367#
x_PM_SKY130_FD_SC_LP__SDFBBN_1%A_27_474# N_A_27_474#_M1024_s N_A_27_474#_M1031_d
+ N_A_27_474#_c_1894_n N_A_27_474#_c_1895_n N_A_27_474#_c_1896_n
+ N_A_27_474#_c_1897_n N_A_27_474#_c_1898_n N_A_27_474#_c_1899_n
+ N_A_27_474#_c_1900_n PM_SKY130_FD_SC_LP__SDFBBN_1%A_27_474#
x_PM_SKY130_FD_SC_LP__SDFBBN_1%VPWR N_VPWR_M1024_d N_VPWR_M1047_s N_VPWR_M1029_s
+ N_VPWR_M1018_d N_VPWR_M1009_d N_VPWR_M1003_d N_VPWR_M1037_d N_VPWR_M1044_d
+ N_VPWR_M1019_d N_VPWR_M1002_d N_VPWR_c_1941_n N_VPWR_c_1942_n N_VPWR_c_1943_n
+ N_VPWR_c_1944_n N_VPWR_c_1945_n N_VPWR_c_1946_n N_VPWR_c_1947_n
+ N_VPWR_c_1948_n N_VPWR_c_1949_n N_VPWR_c_1950_n N_VPWR_c_1951_n
+ N_VPWR_c_1952_n N_VPWR_c_1953_n N_VPWR_c_1954_n N_VPWR_c_1955_n
+ N_VPWR_c_1956_n N_VPWR_c_1957_n N_VPWR_c_1958_n VPWR N_VPWR_c_1959_n
+ N_VPWR_c_1960_n N_VPWR_c_1961_n N_VPWR_c_1962_n N_VPWR_c_1963_n
+ N_VPWR_c_1964_n N_VPWR_c_1965_n N_VPWR_c_1940_n N_VPWR_c_1967_n
+ N_VPWR_c_1968_n N_VPWR_c_1969_n N_VPWR_c_1970_n N_VPWR_c_1971_n
+ N_VPWR_c_1972_n PM_SKY130_FD_SC_LP__SDFBBN_1%VPWR
x_PM_SKY130_FD_SC_LP__SDFBBN_1%A_200_119# N_A_200_119#_M1012_d
+ N_A_200_119#_M1005_s N_A_200_119#_M1046_d N_A_200_119#_M1033_s
+ N_A_200_119#_c_2126_n N_A_200_119#_c_2127_n N_A_200_119#_c_2128_n
+ N_A_200_119#_c_2132_n N_A_200_119#_c_2133_n N_A_200_119#_c_2134_n
+ N_A_200_119#_c_2129_n N_A_200_119#_c_2135_n N_A_200_119#_c_2136_n
+ N_A_200_119#_c_2137_n N_A_200_119#_c_2138_n N_A_200_119#_c_2139_n
+ N_A_200_119#_c_2140_n N_A_200_119#_c_2141_n N_A_200_119#_c_2142_n
+ N_A_200_119#_c_2143_n N_A_200_119#_c_2144_n N_A_200_119#_c_2145_n
+ N_A_200_119#_c_2146_n N_A_200_119#_c_2147_n N_A_200_119#_c_2148_n
+ N_A_200_119#_c_2149_n N_A_200_119#_c_2150_n N_A_200_119#_c_2151_n
+ N_A_200_119#_c_2130_n N_A_200_119#_c_2131_n
+ PM_SKY130_FD_SC_LP__SDFBBN_1%A_200_119#
x_PM_SKY130_FD_SC_LP__SDFBBN_1%Q_N N_Q_N_M1021_d N_Q_N_M1020_d N_Q_N_c_2304_n
+ N_Q_N_c_2305_n Q_N Q_N Q_N Q_N N_Q_N_c_2306_n PM_SKY130_FD_SC_LP__SDFBBN_1%Q_N
x_PM_SKY130_FD_SC_LP__SDFBBN_1%Q N_Q_M1023_d N_Q_M1004_d N_Q_c_2336_n
+ N_Q_c_2337_n N_Q_c_2333_n Q Q N_Q_c_2335_n Q PM_SKY130_FD_SC_LP__SDFBBN_1%Q
x_PM_SKY130_FD_SC_LP__SDFBBN_1%VGND N_VGND_M1032_s N_VGND_M1013_d N_VGND_M1015_s
+ N_VGND_M1039_d N_VGND_M1040_d N_VGND_M1027_s N_VGND_M1025_d N_VGND_M1006_d
+ N_VGND_M1041_d N_VGND_c_2358_n N_VGND_c_2359_n N_VGND_c_2360_n N_VGND_c_2361_n
+ N_VGND_c_2362_n N_VGND_c_2363_n N_VGND_c_2364_n N_VGND_c_2365_n
+ N_VGND_c_2366_n N_VGND_c_2367_n N_VGND_c_2368_n N_VGND_c_2369_n
+ N_VGND_c_2370_n N_VGND_c_2371_n N_VGND_c_2372_n VGND N_VGND_c_2373_n
+ N_VGND_c_2374_n N_VGND_c_2375_n N_VGND_c_2376_n N_VGND_c_2377_n
+ N_VGND_c_2378_n N_VGND_c_2379_n N_VGND_c_2380_n N_VGND_c_2381_n
+ N_VGND_c_2382_n N_VGND_c_2383_n N_VGND_c_2384_n N_VGND_c_2385_n
+ PM_SKY130_FD_SC_LP__SDFBBN_1%VGND
x_PM_SKY130_FD_SC_LP__SDFBBN_1%A_1752_60# N_A_1752_60#_M1035_d
+ N_A_1752_60#_M1008_d N_A_1752_60#_c_2540_n N_A_1752_60#_c_2537_n
+ N_A_1752_60#_c_2544_n PM_SKY130_FD_SC_LP__SDFBBN_1%A_1752_60#
x_PM_SKY130_FD_SC_LP__SDFBBN_1%A_2636_119# N_A_2636_119#_M1022_d
+ N_A_2636_119#_M1017_d N_A_2636_119#_c_2567_n N_A_2636_119#_c_2568_n
+ N_A_2636_119#_c_2569_n PM_SKY130_FD_SC_LP__SDFBBN_1%A_2636_119#
cc_1 VNB N_SCD_c_349_n 0.0214477f $X=-0.19 $Y=-0.245 $X2=0.415 $Y2=1.69
cc_2 VNB N_SCD_M1032_g 0.0281569f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=0.805
cc_3 VNB N_SCD_c_351_n 0.0233877f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.38
cc_4 VNB N_SCD_c_352_n 0.0187576f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.38
cc_5 VNB N_D_M1007_g 0.0164933f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=1.215
cc_6 VNB N_D_c_382_n 0.0244557f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB D 8.6426e-19 $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.38
cc_8 VNB N_D_c_384_n 0.0231976f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_328_429#_M1013_g 0.0206581f $X=-0.19 $Y=-0.245 $X2=0.415 $Y2=1.38
cc_10 VNB N_A_328_429#_c_431_n 0.00873642f $X=-0.19 $Y=-0.245 $X2=0.415
+ $Y2=1.215
cc_11 VNB N_A_328_429#_c_432_n 0.00907398f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_328_429#_c_433_n 0.0138383f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_328_429#_c_434_n 0.0462703f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_328_429#_c_435_n 0.00314773f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_328_429#_c_436_n 0.00595775f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_328_429#_c_437_n 0.0165665f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_328_429#_c_438_n 0.00466621f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_SCE_M1012_g 0.0364036f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=2.69
cc_19 VNB N_SCE_M1042_g 0.00562267f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=1.215
cc_20 VNB N_SCE_c_505_n 0.15002f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=0.805
cc_21 VNB N_SCE_c_506_n 0.0125534f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_SCE_M1010_g 0.0633162f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_SCE_c_508_n 0.0315617f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_SCE_c_509_n 0.00561632f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.55
cc_25 VNB N_CLK_N_M1015_g 0.0295765f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.885
cc_26 VNB N_CLK_N_c_569_n 0.00996808f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_CLK_N_c_570_n 0.0267776f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_28 VNB N_CLK_N_c_571_n 0.0181805f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_CLK_N_c_572_n 0.0176201f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.55
cc_30 VNB N_CLK_N_c_573_n 0.00944441f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_838_50#_M1039_g 0.0133978f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_838_50#_M1018_g 0.00645638f $X=-0.19 $Y=-0.245 $X2=0.415 $Y2=1.38
cc_33 VNB N_A_838_50#_c_619_n 0.135533f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.38
cc_34 VNB N_A_838_50#_c_620_n 0.012806f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.38
cc_35 VNB N_A_838_50#_M1028_g 0.0301209f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_A_838_50#_c_622_n 0.122956f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_838_50#_c_623_n 0.0354055f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_838_50#_c_624_n 0.00177279f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_838_50#_c_625_n 0.00215208f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_838_50#_c_626_n 0.00469123f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_838_50#_c_627_n 0.0383084f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_838_50#_c_628_n 0.0157956f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_838_50#_c_629_n 0.00165058f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_838_50#_c_630_n 0.0163544f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_838_50#_c_631_n 0.00729763f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_838_50#_c_632_n 2.33994e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_838_50#_c_633_n 0.00698745f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_838_50#_c_634_n 0.0154261f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_838_50#_c_635_n 0.00991418f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_838_50#_c_636_n 0.00406917f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_838_50#_c_637_n 0.00420583f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_838_50#_c_638_n 0.0223114f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_838_50#_c_639_n 0.01841f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_1445_324#_c_866_n 0.00394549f $X=-0.19 $Y=-0.245 $X2=0.415
+ $Y2=1.885
cc_55 VNB N_A_1445_324#_M1040_g 0.0420158f $X=-0.19 $Y=-0.245 $X2=0.415 $Y2=1.38
cc_56 VNB N_A_1445_324#_M1027_g 0.0193017f $X=-0.19 $Y=-0.245 $X2=0.24 $Y2=1.55
cc_57 VNB N_A_1445_324#_c_869_n 0.00189714f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_1445_324#_c_870_n 0.0353526f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_1445_324#_c_871_n 0.00504312f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_1445_324#_c_872_n 0.0037876f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_A_1445_324#_c_873_n 0.0235567f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_A_1445_324#_c_874_n 0.00599775f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_A_1445_324#_c_875_n 9.39767e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_64 VNB N_A_1445_324#_c_876_n 0.00982162f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_SET_B_M1035_g 0.0239598f $X=-0.19 $Y=-0.245 $X2=0.495 $Y2=1.885
cc_66 VNB N_SET_B_M1030_g 0.0143588f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=1.215
cc_67 VNB N_SET_B_c_1008_n 0.0290476f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_SET_B_c_1009_n 0.0026055f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_SET_B_c_1010_n 0.00533774f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_SET_B_c_1011_n 0.00155964f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_SET_B_c_1012_n 0.00185772f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_SET_B_c_1013_n 0.0322355f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_SET_B_c_1014_n 0.0260768f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_SET_B_c_1015_n 0.0163194f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_A_1295_379#_M1000_g 0.0387256f $X=-0.19 $Y=-0.245 $X2=0.535
+ $Y2=0.805
cc_76 VNB N_A_1295_379#_c_1147_n 0.0137914f $X=-0.19 $Y=-0.245 $X2=0.415
+ $Y2=1.885
cc_77 VNB N_A_1295_379#_c_1148_n 0.0312413f $X=-0.19 $Y=-0.245 $X2=0.155
+ $Y2=1.58
cc_78 VNB N_A_1295_379#_c_1149_n 0.0147531f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_A_1295_379#_c_1150_n 0.00365671f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_A_1295_379#_c_1151_n 0.0162949f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_A_1295_379#_c_1152_n 0.0022362f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_A_1295_379#_c_1153_n 0.00794818f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_A_1295_379#_c_1154_n 0.00770197f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_A_1295_379#_c_1155_n 8.06062e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_A_1295_379#_c_1156_n 0.00459633f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_A_995_66#_c_1275_n 0.0235022f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=1.215
cc_87 VNB N_A_995_66#_M1005_g 0.0333333f $X=-0.19 $Y=-0.245 $X2=0.415 $Y2=1.885
cc_88 VNB N_A_995_66#_c_1277_n 0.0168884f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_A_995_66#_c_1278_n 0.0289109f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.38
cc_90 VNB N_A_995_66#_c_1279_n 0.0142017f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_A_995_66#_c_1280_n 0.0133793f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_A_995_66#_c_1281_n 0.00538457f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_93 VNB N_A_995_66#_c_1282_n 0.0178097f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_94 VNB N_A_995_66#_c_1283_n 0.010339f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_95 VNB N_A_995_66#_c_1284_n 0.00622102f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_96 VNB N_A_995_66#_c_1285_n 0.00113286f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_97 VNB N_A_995_66#_c_1286_n 0.0328526f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_98 VNB N_A_2449_137#_c_1397_n 0.0159321f $X=-0.19 $Y=-0.245 $X2=0.535
+ $Y2=1.215
cc_99 VNB N_A_2449_137#_c_1398_n 0.0322275f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_100 VNB N_A_2449_137#_c_1399_n 0.00751986f $X=-0.19 $Y=-0.245 $X2=0.415
+ $Y2=1.885
cc_101 VNB N_A_2449_137#_M1021_g 0.026594f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_102 VNB N_A_2449_137#_c_1401_n 0.0586355f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_103 VNB N_A_2449_137#_c_1402_n 0.0231336f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_104 VNB N_A_2449_137#_M1002_g 0.00999973f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_105 VNB N_A_2449_137#_c_1404_n 0.017518f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_106 VNB N_A_2449_137#_c_1405_n 0.0116908f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_107 VNB N_A_2449_137#_c_1406_n 0.00391059f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_108 VNB N_A_2449_137#_c_1407_n 5.82258e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_109 VNB N_A_2449_137#_c_1408_n 0.00564451f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_110 VNB N_A_2449_137#_c_1409_n 0.00473438f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_111 VNB N_A_2449_137#_c_1410_n 0.00414001f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_112 VNB N_A_2449_137#_c_1411_n 0.0153729f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_113 VNB N_A_2449_137#_c_1412_n 0.0252773f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_114 VNB N_A_2299_119#_M1036_g 0.0225443f $X=-0.19 $Y=-0.245 $X2=0.535
+ $Y2=0.805
cc_115 VNB N_A_2299_119#_c_1584_n 0.00732847f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_116 VNB N_A_2299_119#_c_1585_n 0.002624f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_117 VNB N_A_2299_119#_c_1586_n 0.00369232f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_118 VNB N_A_2299_119#_c_1587_n 0.0267912f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_119 VNB N_A_2299_119#_c_1588_n 0.00113995f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_120 VNB N_A_1926_21#_M1008_g 0.00560268f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_121 VNB N_A_1926_21#_c_1682_n 0.342046f $X=-0.19 $Y=-0.245 $X2=0.415
+ $Y2=1.885
cc_122 VNB N_A_1926_21#_c_1683_n 0.0113948f $X=-0.19 $Y=-0.245 $X2=0.155
+ $Y2=1.58
cc_123 VNB N_A_1926_21#_c_1684_n 0.0373631f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_124 VNB N_A_1926_21#_c_1685_n 0.00781239f $X=-0.19 $Y=-0.245 $X2=0.415
+ $Y2=1.38
cc_125 VNB N_A_1926_21#_M1003_g 0.0265197f $X=-0.19 $Y=-0.245 $X2=0.415
+ $Y2=1.215
cc_126 VNB N_A_1926_21#_M1017_g 0.0137722f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_127 VNB N_A_1926_21#_c_1688_n 0.00727896f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_128 VNB N_A_1926_21#_c_1689_n 0.0289948f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_129 VNB N_A_1926_21#_c_1690_n 0.0264124f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_130 VNB N_A_1926_21#_c_1691_n 0.0183305f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_131 VNB N_A_1926_21#_c_1692_n 0.00589937f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_132 VNB N_A_1926_21#_c_1693_n 0.0111812f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_133 VNB N_RESET_B_M1006_g 0.0551382f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=1.215
cc_134 VNB N_RESET_B_c_1804_n 0.0255668f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_135 VNB N_RESET_B_c_1805_n 0.0043203f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_136 VNB N_A_3279_367#_M1023_g 0.0258656f $X=-0.19 $Y=-0.245 $X2=0.535
+ $Y2=0.805
cc_137 VNB N_A_3279_367#_M1004_g 0.00114141f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_138 VNB N_A_3279_367#_c_1843_n 0.0153531f $X=-0.19 $Y=-0.245 $X2=0.415
+ $Y2=1.215
cc_139 VNB N_A_3279_367#_c_1844_n 0.00670802f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_140 VNB N_A_3279_367#_c_1845_n 0.0360412f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_141 VNB N_A_3279_367#_c_1846_n 0.00223902f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_142 VNB N_VPWR_c_1940_n 0.740851f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_143 VNB N_A_200_119#_c_2126_n 0.00256999f $X=-0.19 $Y=-0.245 $X2=0.385
+ $Y2=1.38
cc_144 VNB N_A_200_119#_c_2127_n 0.00620164f $X=-0.19 $Y=-0.245 $X2=0.415
+ $Y2=1.215
cc_145 VNB N_A_200_119#_c_2128_n 0.00265362f $X=-0.19 $Y=-0.245 $X2=0.24
+ $Y2=1.55
cc_146 VNB N_A_200_119#_c_2129_n 0.00405027f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_147 VNB N_A_200_119#_c_2130_n 0.00995888f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_148 VNB N_A_200_119#_c_2131_n 0.0107839f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_149 VNB N_Q_N_c_2304_n 0.0102988f $X=-0.19 $Y=-0.245 $X2=0.535 $Y2=0.805
cc_150 VNB N_Q_N_c_2305_n 0.00637308f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_151 VNB N_Q_N_c_2306_n 0.00499313f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_152 VNB N_Q_c_2333_n 0.0250379f $X=-0.19 $Y=-0.245 $X2=0.385 $Y2=1.38
cc_153 VNB Q 0.0111388f $X=-0.19 $Y=-0.245 $X2=0.415 $Y2=1.215
cc_154 VNB N_Q_c_2335_n 0.0292706f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_155 VNB N_VGND_c_2358_n 0.0134927f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_156 VNB N_VGND_c_2359_n 0.0425682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_157 VNB N_VGND_c_2360_n 0.01451f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_158 VNB N_VGND_c_2361_n 0.0218982f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_159 VNB N_VGND_c_2362_n 0.0199414f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_160 VNB N_VGND_c_2363_n 0.0100818f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_161 VNB N_VGND_c_2364_n 0.0117815f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_162 VNB N_VGND_c_2365_n 0.0524399f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_163 VNB N_VGND_c_2366_n 0.0190236f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_164 VNB N_VGND_c_2367_n 0.0157811f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_165 VNB N_VGND_c_2368_n 0.00478154f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_166 VNB N_VGND_c_2369_n 0.0282712f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_167 VNB N_VGND_c_2370_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_168 VNB N_VGND_c_2371_n 0.0308597f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_169 VNB N_VGND_c_2372_n 0.00397464f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_170 VNB N_VGND_c_2373_n 0.0507567f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_171 VNB N_VGND_c_2374_n 0.0397277f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_172 VNB N_VGND_c_2375_n 0.058416f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_173 VNB N_VGND_c_2376_n 0.056007f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_174 VNB N_VGND_c_2377_n 0.0604952f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_175 VNB N_VGND_c_2378_n 0.0202074f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_176 VNB N_VGND_c_2379_n 0.88759f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_177 VNB N_VGND_c_2380_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_178 VNB N_VGND_c_2381_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_179 VNB N_VGND_c_2382_n 0.00631792f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_180 VNB N_VGND_c_2383_n 0.00332923f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_181 VNB N_VGND_c_2384_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_182 VNB N_VGND_c_2385_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_183 VNB N_A_1752_60#_c_2537_n 0.00292629f $X=-0.19 $Y=-0.245 $X2=0.415
+ $Y2=1.38
cc_184 VNB N_A_2636_119#_c_2567_n 0.0146285f $X=-0.19 $Y=-0.245 $X2=0.535
+ $Y2=1.215
cc_185 VNB N_A_2636_119#_c_2568_n 0.00357136f $X=-0.19 $Y=-0.245 $X2=0.415
+ $Y2=1.885
cc_186 VNB N_A_2636_119#_c_2569_n 0.00798634f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_187 VPB N_SCD_c_349_n 0.00298862f $X=-0.19 $Y=1.655 $X2=0.415 $Y2=1.69
cc_188 VPB N_SCD_M1024_g 0.0457368f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=2.69
cc_189 VPB N_SCD_c_355_n 0.0234049f $X=-0.19 $Y=1.655 $X2=0.415 $Y2=1.885
cc_190 VPB N_SCD_c_352_n 0.00971735f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.38
cc_191 VPB N_D_M1046_g 0.0328851f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=1.885
cc_192 VPB N_D_c_382_n 0.0436825f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_193 VPB N_A_328_429#_c_439_n 0.0177856f $X=-0.19 $Y=1.655 $X2=0.535 $Y2=1.215
cc_194 VPB N_A_328_429#_c_440_n 0.0313225f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_195 VPB N_A_328_429#_c_441_n 0.00667472f $X=-0.19 $Y=1.655 $X2=0.415
+ $Y2=1.885
cc_196 VPB N_A_328_429#_c_431_n 0.0296082f $X=-0.19 $Y=1.655 $X2=0.415 $Y2=1.215
cc_197 VPB N_A_328_429#_c_436_n 0.0120157f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_198 VPB N_SCE_M1042_g 0.0445552f $X=-0.19 $Y=1.655 $X2=0.535 $Y2=1.215
cc_199 VPB N_SCE_M1010_g 0.0373653f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_200 VPB N_SCE_c_509_n 0.00629667f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.55
cc_201 VPB N_CLK_N_c_569_n 0.0100207f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_202 VPB N_CLK_N_c_575_n 0.0216206f $X=-0.19 $Y=1.655 $X2=0.535 $Y2=1.215
cc_203 VPB N_CLK_N_c_576_n 0.0327792f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.38
cc_204 VPB N_A_838_50#_M1018_g 0.0569428f $X=-0.19 $Y=1.655 $X2=0.415 $Y2=1.38
cc_205 VPB N_A_838_50#_c_641_n 0.0744605f $X=-0.19 $Y=1.655 $X2=0.415 $Y2=1.215
cc_206 VPB N_A_838_50#_c_642_n 0.0129911f $X=-0.19 $Y=1.655 $X2=0.24 $Y2=1.55
cc_207 VPB N_A_838_50#_M1033_g 0.0641245f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.55
cc_208 VPB N_A_838_50#_c_644_n 0.0157934f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_209 VPB N_A_838_50#_c_645_n 0.0375757f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_210 VPB N_A_838_50#_c_625_n 0.0193585f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_211 VPB N_A_838_50#_c_633_n 0.00420577f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_212 VPB N_A_838_50#_c_648_n 0.00669695f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_213 VPB N_A_838_50#_c_649_n 0.00839291f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_214 VPB N_A_838_50#_c_650_n 0.00222326f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_215 VPB N_A_838_50#_c_651_n 0.0043737f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_216 VPB N_A_838_50#_c_652_n 0.0504076f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_217 VPB N_A_838_50#_c_638_n 0.00739466f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_218 VPB N_A_1445_324#_c_877_n 0.0219665f $X=-0.19 $Y=1.655 $X2=0.535
+ $Y2=1.215
cc_219 VPB N_A_1445_324#_c_866_n 0.00393767f $X=-0.19 $Y=1.655 $X2=0.415
+ $Y2=1.885
cc_220 VPB N_A_1445_324#_M1043_g 0.021346f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_221 VPB N_A_1445_324#_c_869_n 0.00274301f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_222 VPB N_A_1445_324#_c_870_n 0.0275686f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_223 VPB N_A_1445_324#_c_882_n 0.00493905f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_224 VPB N_A_1445_324#_c_872_n 0.0110683f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_225 VPB N_A_1445_324#_c_873_n 0.0151829f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_226 VPB N_A_1445_324#_c_885_n 0.00289127f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_227 VPB N_A_1445_324#_c_876_n 0.00889014f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_228 VPB N_SET_B_M1030_g 0.0318413f $X=-0.19 $Y=1.655 $X2=0.535 $Y2=1.215
cc_229 VPB N_SET_B_c_1017_n 0.0177884f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_230 VPB N_SET_B_M1011_g 0.0195077f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.38
cc_231 VPB N_SET_B_c_1019_n 0.0223113f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_232 VPB N_SET_B_c_1012_n 0.00274999f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_233 VPB N_SET_B_c_1014_n 0.00647704f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_234 VPB N_A_1295_379#_c_1147_n 0.0131126f $X=-0.19 $Y=1.655 $X2=0.415
+ $Y2=1.885
cc_235 VPB N_A_1295_379#_c_1148_n 0.0134813f $X=-0.19 $Y=1.655 $X2=0.155
+ $Y2=1.58
cc_236 VPB N_A_1295_379#_M1001_g 0.0224782f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.38
cc_237 VPB N_A_1295_379#_c_1149_n 0.00166945f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_238 VPB N_A_1295_379#_c_1161_n 0.00524413f $X=-0.19 $Y=1.655 $X2=0.385
+ $Y2=1.55
cc_239 VPB N_A_1295_379#_c_1150_n 0.00185252f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_240 VPB N_A_1295_379#_c_1154_n 0.00636682f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_241 VPB N_A_1295_379#_c_1155_n 0.00293096f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_242 VPB N_A_1295_379#_c_1165_n 0.0126991f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_243 VPB N_A_1295_379#_c_1156_n 0.00342769f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_244 VPB N_A_995_66#_c_1278_n 0.0130806f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.38
cc_245 VPB N_A_995_66#_M1034_g 0.0665799f $X=-0.19 $Y=1.655 $X2=0.24 $Y2=1.55
cc_246 VPB N_A_995_66#_c_1289_n 0.379496f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_247 VPB N_A_995_66#_c_1290_n 0.0103267f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_248 VPB N_A_995_66#_M1038_g 0.0103825f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_249 VPB N_A_995_66#_c_1292_n 0.02577f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_250 VPB N_A_995_66#_c_1293_n 0.00845077f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_251 VPB N_A_995_66#_c_1279_n 0.0167653f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_252 VPB N_A_995_66#_c_1295_n 0.00614339f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_253 VPB N_A_995_66#_c_1284_n 0.00435334f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_254 VPB N_A_995_66#_c_1286_n 0.0125101f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_255 VPB N_A_2449_137#_M1037_g 0.0291987f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.38
cc_256 VPB N_A_2449_137#_M1020_g 0.0253502f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_257 VPB N_A_2449_137#_M1002_g 0.0257445f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_258 VPB N_A_2449_137#_c_1416_n 0.0186682f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_259 VPB N_A_2449_137#_c_1417_n 0.0360965f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_260 VPB N_A_2449_137#_c_1408_n 0.00369291f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_261 VPB N_A_2449_137#_c_1419_n 0.0152241f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_262 VPB N_A_2449_137#_c_1420_n 0.00139956f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_263 VPB N_A_2449_137#_c_1411_n 0.0179972f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_264 VPB N_A_2449_137#_c_1412_n 0.00674696f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_265 VPB N_A_2299_119#_M1045_g 0.0352244f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_266 VPB N_A_2299_119#_c_1590_n 0.00345227f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_267 VPB N_A_2299_119#_c_1585_n 0.00372898f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_268 VPB N_A_2299_119#_c_1586_n 0.00286103f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_269 VPB N_A_2299_119#_c_1587_n 0.0171199f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_270 VPB N_A_1926_21#_M1003_g 0.0220021f $X=-0.19 $Y=1.655 $X2=0.415 $Y2=1.215
cc_271 VPB N_A_1926_21#_M1044_g 0.0350209f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.55
cc_272 VPB N_A_1926_21#_c_1688_n 0.0221989f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_273 VPB N_A_1926_21#_c_1697_n 0.00370839f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_274 VPB N_A_1926_21#_c_1698_n 0.00640151f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_275 VPB N_A_1926_21#_c_1699_n 0.0102441f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_276 VPB N_RESET_B_M1019_g 0.0211451f $X=-0.19 $Y=1.655 $X2=0.495 $Y2=1.885
cc_277 VPB N_RESET_B_c_1804_n 0.00652585f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_278 VPB N_RESET_B_c_1805_n 0.00449264f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_279 VPB N_A_3279_367#_M1004_g 0.0281049f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_280 VPB N_A_3279_367#_c_1848_n 0.00647595f $X=-0.19 $Y=1.655 $X2=0.385
+ $Y2=1.55
cc_281 VPB N_A_27_474#_c_1894_n 0.0330052f $X=-0.19 $Y=1.655 $X2=0.535 $Y2=0.805
cc_282 VPB N_A_27_474#_c_1895_n 0.0171528f $X=-0.19 $Y=1.655 $X2=0.415 $Y2=1.885
cc_283 VPB N_A_27_474#_c_1896_n 0.00993659f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_284 VPB N_A_27_474#_c_1897_n 8.03639e-19 $X=-0.19 $Y=1.655 $X2=0.415 $Y2=1.38
cc_285 VPB N_A_27_474#_c_1898_n 0.00709754f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.38
cc_286 VPB N_A_27_474#_c_1899_n 0.00107431f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.38
cc_287 VPB N_A_27_474#_c_1900_n 0.00866679f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_288 VPB N_VPWR_c_1941_n 0.00426277f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_289 VPB N_VPWR_c_1942_n 0.0166081f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_290 VPB N_VPWR_c_1943_n 0.0154267f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_291 VPB N_VPWR_c_1944_n 0.00978424f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_292 VPB N_VPWR_c_1945_n 0.0401468f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_293 VPB N_VPWR_c_1946_n 0.0125415f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_294 VPB N_VPWR_c_1947_n 0.00793993f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_295 VPB N_VPWR_c_1948_n 0.0132256f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_296 VPB N_VPWR_c_1949_n 0.0132256f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_297 VPB N_VPWR_c_1950_n 0.0176382f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_298 VPB N_VPWR_c_1951_n 0.04053f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_299 VPB N_VPWR_c_1952_n 0.00324402f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_300 VPB N_VPWR_c_1953_n 0.0310571f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_301 VPB N_VPWR_c_1954_n 0.00324402f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_302 VPB N_VPWR_c_1955_n 0.0507727f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_303 VPB N_VPWR_c_1956_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_304 VPB N_VPWR_c_1957_n 0.0248802f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_305 VPB N_VPWR_c_1958_n 0.00510392f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_306 VPB N_VPWR_c_1959_n 0.0168624f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_307 VPB N_VPWR_c_1960_n 0.036328f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_308 VPB N_VPWR_c_1961_n 0.0774965f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_309 VPB N_VPWR_c_1962_n 0.064146f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_310 VPB N_VPWR_c_1963_n 0.0204067f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_311 VPB N_VPWR_c_1964_n 0.0327055f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_312 VPB N_VPWR_c_1965_n 0.0187754f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_313 VPB N_VPWR_c_1940_n 0.183635f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_314 VPB N_VPWR_c_1967_n 0.00421413f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_315 VPB N_VPWR_c_1968_n 0.00455177f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_316 VPB N_VPWR_c_1969_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_317 VPB N_VPWR_c_1970_n 0.0047828f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_318 VPB N_VPWR_c_1971_n 0.00510392f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_319 VPB N_VPWR_c_1972_n 0.0047828f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_320 VPB N_A_200_119#_c_2132_n 0.00185133f $X=-0.19 $Y=1.655 $X2=0.385
+ $Y2=1.55
cc_321 VPB N_A_200_119#_c_2133_n 0.0093765f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_322 VPB N_A_200_119#_c_2134_n 0.00198304f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_323 VPB N_A_200_119#_c_2135_n 0.00168925f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_324 VPB N_A_200_119#_c_2136_n 0.0214991f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_325 VPB N_A_200_119#_c_2137_n 0.00475124f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_326 VPB N_A_200_119#_c_2138_n 0.0211538f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_327 VPB N_A_200_119#_c_2139_n 0.00326464f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_328 VPB N_A_200_119#_c_2140_n 0.0222658f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_329 VPB N_A_200_119#_c_2141_n 0.0268974f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_330 VPB N_A_200_119#_c_2142_n 0.00919848f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_331 VPB N_A_200_119#_c_2143_n 0.00586934f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_332 VPB N_A_200_119#_c_2144_n 0.0289016f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_333 VPB N_A_200_119#_c_2145_n 0.00326464f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_334 VPB N_A_200_119#_c_2146_n 0.0062406f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_335 VPB N_A_200_119#_c_2147_n 0.0121325f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_336 VPB N_A_200_119#_c_2148_n 2.08773e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_337 VPB N_A_200_119#_c_2149_n 0.004864f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_338 VPB N_A_200_119#_c_2150_n 0.00458171f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_339 VPB N_A_200_119#_c_2151_n 0.00124796f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_340 VPB N_A_200_119#_c_2130_n 0.0060442f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_341 VPB Q_N 0.00454816f $X=-0.19 $Y=1.655 $X2=0.415 $Y2=1.38
cc_342 VPB Q_N 0.0183979f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_343 VPB N_Q_N_c_2306_n 0.00347423f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_344 VPB N_Q_c_2336_n 0.0423813f $X=-0.19 $Y=1.655 $X2=0.535 $Y2=0.805
cc_345 VPB N_Q_c_2337_n 0.0126596f $X=-0.19 $Y=1.655 $X2=0.415 $Y2=1.38
cc_346 VPB N_Q_c_2333_n 0.00769959f $X=-0.19 $Y=1.655 $X2=0.385 $Y2=1.38
cc_347 N_SCD_M1032_g N_SCE_M1012_g 0.0244496f $X=0.535 $Y=0.805 $X2=0 $Y2=0
cc_348 N_SCD_c_349_n N_SCE_M1042_g 0.0244496f $X=0.415 $Y=1.69 $X2=0 $Y2=0
cc_349 N_SCD_M1024_g N_SCE_M1042_g 0.0380122f $X=0.495 $Y=2.69 $X2=0 $Y2=0
cc_350 N_SCD_c_351_n N_SCE_c_508_n 0.0244496f $X=0.385 $Y=1.38 $X2=0 $Y2=0
cc_351 N_SCD_c_352_n N_SCE_c_508_n 0.00237421f $X=0.385 $Y=1.38 $X2=0 $Y2=0
cc_352 N_SCD_c_351_n N_SCE_c_509_n 0.00221828f $X=0.385 $Y=1.38 $X2=0 $Y2=0
cc_353 N_SCD_c_352_n N_SCE_c_509_n 0.0281146f $X=0.385 $Y=1.38 $X2=0 $Y2=0
cc_354 N_SCD_M1024_g N_A_27_474#_c_1894_n 0.00422578f $X=0.495 $Y=2.69 $X2=0
+ $Y2=0
cc_355 N_SCD_M1024_g N_A_27_474#_c_1895_n 0.0163546f $X=0.495 $Y=2.69 $X2=0
+ $Y2=0
cc_356 N_SCD_c_355_n N_A_27_474#_c_1895_n 0.00305832f $X=0.415 $Y=1.885 $X2=0
+ $Y2=0
cc_357 N_SCD_c_352_n N_A_27_474#_c_1895_n 0.0135489f $X=0.385 $Y=1.38 $X2=0
+ $Y2=0
cc_358 N_SCD_c_355_n N_A_27_474#_c_1896_n 0.00387047f $X=0.415 $Y=1.885 $X2=0
+ $Y2=0
cc_359 N_SCD_c_352_n N_A_27_474#_c_1896_n 0.0208104f $X=0.385 $Y=1.38 $X2=0
+ $Y2=0
cc_360 N_SCD_M1024_g N_A_27_474#_c_1897_n 7.44326e-19 $X=0.495 $Y=2.69 $X2=0
+ $Y2=0
cc_361 N_SCD_M1024_g N_VPWR_c_1941_n 0.0140978f $X=0.495 $Y=2.69 $X2=0 $Y2=0
cc_362 N_SCD_M1024_g N_VPWR_c_1959_n 0.00418439f $X=0.495 $Y=2.69 $X2=0 $Y2=0
cc_363 N_SCD_M1024_g N_VPWR_c_1940_n 0.00830975f $X=0.495 $Y=2.69 $X2=0 $Y2=0
cc_364 N_SCD_M1032_g N_A_200_119#_c_2126_n 0.00113653f $X=0.535 $Y=0.805 $X2=0
+ $Y2=0
cc_365 N_SCD_M1032_g N_A_200_119#_c_2128_n 4.61477e-19 $X=0.535 $Y=0.805 $X2=0
+ $Y2=0
cc_366 N_SCD_M1032_g N_VGND_c_2359_n 0.0140549f $X=0.535 $Y=0.805 $X2=0 $Y2=0
cc_367 N_SCD_c_351_n N_VGND_c_2359_n 0.00642189f $X=0.385 $Y=1.38 $X2=0 $Y2=0
cc_368 N_SCD_c_352_n N_VGND_c_2359_n 0.0280299f $X=0.385 $Y=1.38 $X2=0 $Y2=0
cc_369 N_SCD_M1032_g N_VGND_c_2373_n 0.0035863f $X=0.535 $Y=0.805 $X2=0 $Y2=0
cc_370 N_SCD_M1032_g N_VGND_c_2379_n 0.00401353f $X=0.535 $Y=0.805 $X2=0 $Y2=0
cc_371 N_D_M1046_g N_A_328_429#_c_441_n 0.0280698f $X=1.285 $Y=2.69 $X2=0 $Y2=0
cc_372 N_D_c_382_n N_A_328_429#_c_441_n 0.0117795f $X=1.62 $Y=1.785 $X2=0 $Y2=0
cc_373 N_D_M1007_g N_A_328_429#_M1013_g 0.0135168f $X=1.495 $Y=0.805 $X2=0 $Y2=0
cc_374 D N_A_328_429#_M1013_g 0.00197155f $X=1.595 $Y=0.84 $X2=0 $Y2=0
cc_375 N_D_c_384_n N_A_328_429#_M1013_g 0.0140408f $X=1.655 $Y=1.315 $X2=0 $Y2=0
cc_376 N_D_M1046_g N_A_328_429#_c_431_n 0.0021027f $X=1.285 $Y=2.69 $X2=0 $Y2=0
cc_377 N_D_c_382_n N_A_328_429#_c_431_n 0.0140408f $X=1.62 $Y=1.785 $X2=0 $Y2=0
cc_378 N_D_c_382_n N_A_328_429#_c_432_n 0.0140408f $X=1.62 $Y=1.785 $X2=0 $Y2=0
cc_379 N_D_M1007_g N_SCE_M1012_g 0.0138415f $X=1.495 $Y=0.805 $X2=0 $Y2=0
cc_380 D N_SCE_M1012_g 9.68477e-19 $X=1.595 $Y=0.84 $X2=0 $Y2=0
cc_381 N_D_c_382_n N_SCE_M1042_g 0.0890219f $X=1.62 $Y=1.785 $X2=0 $Y2=0
cc_382 D N_SCE_M1042_g 3.33332e-19 $X=1.595 $Y=0.84 $X2=0 $Y2=0
cc_383 N_D_M1007_g N_SCE_c_505_n 0.00895556f $X=1.495 $Y=0.805 $X2=0 $Y2=0
cc_384 D N_SCE_c_508_n 2.96468e-19 $X=1.595 $Y=0.84 $X2=0 $Y2=0
cc_385 N_D_c_384_n N_SCE_c_508_n 0.0174492f $X=1.655 $Y=1.315 $X2=0 $Y2=0
cc_386 N_D_c_382_n N_SCE_c_509_n 0.00558444f $X=1.62 $Y=1.785 $X2=0 $Y2=0
cc_387 D N_SCE_c_509_n 0.0439567f $X=1.595 $Y=0.84 $X2=0 $Y2=0
cc_388 N_D_c_384_n N_SCE_c_509_n 0.00477122f $X=1.655 $Y=1.315 $X2=0 $Y2=0
cc_389 N_D_M1046_g N_A_27_474#_c_1895_n 0.00125192f $X=1.285 $Y=2.69 $X2=0 $Y2=0
cc_390 N_D_M1046_g N_A_27_474#_c_1897_n 0.00500666f $X=1.285 $Y=2.69 $X2=0 $Y2=0
cc_391 N_D_M1046_g N_A_27_474#_c_1898_n 0.0127943f $X=1.285 $Y=2.69 $X2=0 $Y2=0
cc_392 N_D_M1046_g N_A_27_474#_c_1900_n 6.44854e-19 $X=1.285 $Y=2.69 $X2=0 $Y2=0
cc_393 N_D_M1046_g N_VPWR_c_1951_n 0.00306988f $X=1.285 $Y=2.69 $X2=0 $Y2=0
cc_394 N_D_M1046_g N_VPWR_c_1940_n 0.00438306f $X=1.285 $Y=2.69 $X2=0 $Y2=0
cc_395 N_D_M1007_g N_A_200_119#_c_2126_n 0.00670476f $X=1.495 $Y=0.805 $X2=0
+ $Y2=0
cc_396 D N_A_200_119#_c_2126_n 0.0167425f $X=1.595 $Y=0.84 $X2=0 $Y2=0
cc_397 N_D_M1007_g N_A_200_119#_c_2127_n 0.0121885f $X=1.495 $Y=0.805 $X2=0
+ $Y2=0
cc_398 D N_A_200_119#_c_2127_n 0.0199759f $X=1.595 $Y=0.84 $X2=0 $Y2=0
cc_399 N_D_c_384_n N_A_200_119#_c_2127_n 7.69817e-19 $X=1.655 $Y=1.315 $X2=0
+ $Y2=0
cc_400 N_D_M1046_g N_A_200_119#_c_2132_n 0.00782017f $X=1.285 $Y=2.69 $X2=0
+ $Y2=0
cc_401 N_D_c_382_n N_A_200_119#_c_2133_n 0.00299411f $X=1.62 $Y=1.785 $X2=0
+ $Y2=0
cc_402 D N_A_200_119#_c_2133_n 0.0178656f $X=1.595 $Y=0.84 $X2=0 $Y2=0
cc_403 N_D_M1046_g N_A_200_119#_c_2134_n 0.0067262f $X=1.285 $Y=2.69 $X2=0 $Y2=0
cc_404 N_D_c_382_n N_A_200_119#_c_2134_n 0.0095336f $X=1.62 $Y=1.785 $X2=0 $Y2=0
cc_405 D N_A_200_119#_c_2134_n 0.00805447f $X=1.595 $Y=0.84 $X2=0 $Y2=0
cc_406 N_D_M1007_g N_A_200_119#_c_2129_n 0.00369033f $X=1.495 $Y=0.805 $X2=0
+ $Y2=0
cc_407 D N_A_200_119#_c_2129_n 0.0637353f $X=1.595 $Y=0.84 $X2=0 $Y2=0
cc_408 N_D_c_384_n N_A_200_119#_c_2129_n 0.00311411f $X=1.655 $Y=1.315 $X2=0
+ $Y2=0
cc_409 N_D_M1046_g N_A_200_119#_c_2135_n 8.91745e-19 $X=1.285 $Y=2.69 $X2=0
+ $Y2=0
cc_410 N_D_c_382_n N_A_200_119#_c_2135_n 0.0016691f $X=1.62 $Y=1.785 $X2=0 $Y2=0
cc_411 N_D_c_382_n N_A_200_119#_c_2151_n 0.00189173f $X=1.62 $Y=1.785 $X2=0
+ $Y2=0
cc_412 D N_A_200_119#_c_2151_n 0.0108693f $X=1.595 $Y=0.84 $X2=0 $Y2=0
cc_413 D A_314_119# 0.00438307f $X=1.595 $Y=0.84 $X2=-0.19 $Y2=-0.245
cc_414 N_A_328_429#_M1013_g N_SCE_c_505_n 0.00934409f $X=2.135 $Y=0.805 $X2=0
+ $Y2=0
cc_415 N_A_328_429#_M1013_g N_SCE_M1010_g 0.00876974f $X=2.135 $Y=0.805 $X2=0
+ $Y2=0
cc_416 N_A_328_429#_c_431_n N_SCE_M1010_g 0.0104365f $X=2.135 $Y=2.145 $X2=0
+ $Y2=0
cc_417 N_A_328_429#_c_433_n N_SCE_M1010_g 0.0272498f $X=3.095 $Y=1.34 $X2=0
+ $Y2=0
cc_418 N_A_328_429#_c_434_n N_SCE_M1010_g 0.0214137f $X=2.515 $Y=1.34 $X2=0
+ $Y2=0
cc_419 N_A_328_429#_c_436_n N_SCE_M1010_g 0.0155703f $X=3.18 $Y=2.2 $X2=0 $Y2=0
cc_420 N_A_328_429#_c_437_n N_SCE_M1010_g 0.0147751f $X=3.26 $Y=0.805 $X2=0
+ $Y2=0
cc_421 N_A_328_429#_c_437_n N_CLK_N_M1015_g 0.00437437f $X=3.26 $Y=0.805 $X2=0
+ $Y2=0
cc_422 N_A_328_429#_c_435_n N_CLK_N_c_570_n 0.00224269f $X=3.18 $Y=1.175 $X2=0
+ $Y2=0
cc_423 N_A_328_429#_c_438_n N_CLK_N_c_570_n 0.0057324f $X=3.18 $Y=1.34 $X2=0
+ $Y2=0
cc_424 N_A_328_429#_c_436_n N_CLK_N_c_571_n 5.6235e-19 $X=3.18 $Y=2.2 $X2=0
+ $Y2=0
cc_425 N_A_328_429#_c_437_n N_CLK_N_c_572_n 0.0031253f $X=3.26 $Y=0.805 $X2=0
+ $Y2=0
cc_426 N_A_328_429#_c_435_n N_CLK_N_c_573_n 0.00402969f $X=3.18 $Y=1.175 $X2=0
+ $Y2=0
cc_427 N_A_328_429#_c_436_n N_CLK_N_c_573_n 0.00100289f $X=3.18 $Y=2.2 $X2=0
+ $Y2=0
cc_428 N_A_328_429#_c_437_n N_CLK_N_c_573_n 0.00648875f $X=3.26 $Y=0.805 $X2=0
+ $Y2=0
cc_429 N_A_328_429#_c_438_n N_CLK_N_c_573_n 0.0108214f $X=3.18 $Y=1.34 $X2=0
+ $Y2=0
cc_430 N_A_328_429#_c_439_n N_A_27_474#_c_1898_n 0.0119176f $X=1.715 $Y=2.295
+ $X2=0 $Y2=0
cc_431 N_A_328_429#_c_439_n N_A_27_474#_c_1900_n 0.0078667f $X=1.715 $Y=2.295
+ $X2=0 $Y2=0
cc_432 N_A_328_429#_c_440_n N_A_27_474#_c_1900_n 0.00730447f $X=2.06 $Y=2.22
+ $X2=0 $Y2=0
cc_433 N_A_328_429#_c_439_n N_VPWR_c_1942_n 0.00367438f $X=1.715 $Y=2.295 $X2=0
+ $Y2=0
cc_434 N_A_328_429#_c_431_n N_VPWR_c_1942_n 0.00463056f $X=2.135 $Y=2.145 $X2=0
+ $Y2=0
cc_435 N_A_328_429#_c_439_n N_VPWR_c_1951_n 0.0030696f $X=1.715 $Y=2.295 $X2=0
+ $Y2=0
cc_436 N_A_328_429#_c_439_n N_VPWR_c_1940_n 0.00499887f $X=1.715 $Y=2.295 $X2=0
+ $Y2=0
cc_437 N_A_328_429#_M1013_g N_A_200_119#_c_2127_n 0.00574801f $X=2.135 $Y=0.805
+ $X2=0 $Y2=0
cc_438 N_A_328_429#_c_441_n N_A_200_119#_c_2132_n 0.00493105f $X=1.79 $Y=2.22
+ $X2=0 $Y2=0
cc_439 N_A_328_429#_c_440_n N_A_200_119#_c_2133_n 0.0117405f $X=2.06 $Y=2.22
+ $X2=0 $Y2=0
cc_440 N_A_328_429#_c_441_n N_A_200_119#_c_2133_n 0.00736166f $X=1.79 $Y=2.22
+ $X2=0 $Y2=0
cc_441 N_A_328_429#_c_431_n N_A_200_119#_c_2133_n 0.00583818f $X=2.135 $Y=2.145
+ $X2=0 $Y2=0
cc_442 N_A_328_429#_M1013_g N_A_200_119#_c_2129_n 0.0192016f $X=2.135 $Y=0.805
+ $X2=0 $Y2=0
cc_443 N_A_328_429#_c_431_n N_A_200_119#_c_2129_n 0.00910508f $X=2.135 $Y=2.145
+ $X2=0 $Y2=0
cc_444 N_A_328_429#_c_432_n N_A_200_119#_c_2129_n 0.00928273f $X=2.135 $Y=1.34
+ $X2=0 $Y2=0
cc_445 N_A_328_429#_c_433_n N_A_200_119#_c_2129_n 0.0238596f $X=3.095 $Y=1.34
+ $X2=0 $Y2=0
cc_446 N_A_328_429#_c_431_n N_A_200_119#_c_2135_n 0.00480634f $X=2.135 $Y=2.145
+ $X2=0 $Y2=0
cc_447 N_A_328_429#_c_431_n N_A_200_119#_c_2136_n 0.00738298f $X=2.135 $Y=2.145
+ $X2=0 $Y2=0
cc_448 N_A_328_429#_c_433_n N_A_200_119#_c_2136_n 0.0428932f $X=3.095 $Y=1.34
+ $X2=0 $Y2=0
cc_449 N_A_328_429#_c_434_n N_A_200_119#_c_2136_n 0.0125341f $X=2.515 $Y=1.34
+ $X2=0 $Y2=0
cc_450 N_A_328_429#_c_436_n N_A_200_119#_c_2136_n 0.0130055f $X=3.18 $Y=2.2
+ $X2=0 $Y2=0
cc_451 N_A_328_429#_c_431_n N_A_200_119#_c_2137_n 0.00158737f $X=2.135 $Y=2.145
+ $X2=0 $Y2=0
cc_452 N_A_328_429#_c_436_n N_A_200_119#_c_2137_n 0.0356849f $X=3.18 $Y=2.2
+ $X2=0 $Y2=0
cc_453 N_A_328_429#_c_436_n N_A_200_119#_c_2138_n 0.0126934f $X=3.18 $Y=2.2
+ $X2=0 $Y2=0
cc_454 N_A_328_429#_c_436_n N_A_200_119#_c_2140_n 0.0587633f $X=3.18 $Y=2.2
+ $X2=0 $Y2=0
cc_455 N_A_328_429#_c_436_n N_A_200_119#_c_2142_n 0.0137874f $X=3.18 $Y=2.2
+ $X2=0 $Y2=0
cc_456 N_A_328_429#_c_431_n N_A_200_119#_c_2151_n 0.00242835f $X=2.135 $Y=2.145
+ $X2=0 $Y2=0
cc_457 N_A_328_429#_M1013_g N_VGND_c_2360_n 0.00543267f $X=2.135 $Y=0.805 $X2=0
+ $Y2=0
cc_458 N_A_328_429#_c_433_n N_VGND_c_2360_n 0.025913f $X=3.095 $Y=1.34 $X2=0
+ $Y2=0
cc_459 N_A_328_429#_c_434_n N_VGND_c_2360_n 0.00760331f $X=2.515 $Y=1.34 $X2=0
+ $Y2=0
cc_460 N_A_328_429#_c_437_n N_VGND_c_2360_n 0.00917501f $X=3.26 $Y=0.805 $X2=0
+ $Y2=0
cc_461 N_A_328_429#_c_437_n N_VGND_c_2361_n 0.00775327f $X=3.26 $Y=0.805 $X2=0
+ $Y2=0
cc_462 N_A_328_429#_c_437_n N_VGND_c_2369_n 0.00745886f $X=3.26 $Y=0.805 $X2=0
+ $Y2=0
cc_463 N_A_328_429#_M1013_g N_VGND_c_2379_n 2.50464e-19 $X=2.135 $Y=0.805 $X2=0
+ $Y2=0
cc_464 N_A_328_429#_c_437_n N_VGND_c_2379_n 0.0103146f $X=3.26 $Y=0.805 $X2=0
+ $Y2=0
cc_465 N_SCE_M1042_g N_A_27_474#_c_1895_n 0.0134025f $X=0.925 $Y=2.69 $X2=0
+ $Y2=0
cc_466 N_SCE_c_508_n N_A_27_474#_c_1895_n 6.94062e-19 $X=1.015 $Y=1.38 $X2=0
+ $Y2=0
cc_467 N_SCE_c_509_n N_A_27_474#_c_1895_n 0.0168229f $X=1.015 $Y=1.38 $X2=0
+ $Y2=0
cc_468 N_SCE_M1042_g N_A_27_474#_c_1897_n 0.0119843f $X=0.925 $Y=2.69 $X2=0
+ $Y2=0
cc_469 N_SCE_M1042_g N_A_27_474#_c_1899_n 0.00347647f $X=0.925 $Y=2.69 $X2=0
+ $Y2=0
cc_470 N_SCE_M1042_g N_VPWR_c_1941_n 0.00294318f $X=0.925 $Y=2.69 $X2=0 $Y2=0
cc_471 N_SCE_M1010_g N_VPWR_c_1942_n 0.00340607f $X=2.965 $Y=0.805 $X2=0 $Y2=0
cc_472 N_SCE_M1042_g N_VPWR_c_1951_n 0.00471106f $X=0.925 $Y=2.69 $X2=0 $Y2=0
cc_473 N_SCE_M1010_g N_VPWR_c_1953_n 2.23678e-19 $X=2.965 $Y=0.805 $X2=0 $Y2=0
cc_474 N_SCE_M1042_g N_VPWR_c_1940_n 0.0089056f $X=0.925 $Y=2.69 $X2=0 $Y2=0
cc_475 N_SCE_M1012_g N_A_200_119#_c_2126_n 0.00734793f $X=0.925 $Y=0.805 $X2=0
+ $Y2=0
cc_476 N_SCE_c_508_n N_A_200_119#_c_2126_n 0.00138585f $X=1.015 $Y=1.38 $X2=0
+ $Y2=0
cc_477 N_SCE_c_509_n N_A_200_119#_c_2126_n 0.0277564f $X=1.015 $Y=1.38 $X2=0
+ $Y2=0
cc_478 N_SCE_c_505_n N_A_200_119#_c_2127_n 0.0142384f $X=2.89 $Y=0.18 $X2=0
+ $Y2=0
cc_479 N_SCE_M1012_g N_A_200_119#_c_2128_n 0.00554337f $X=0.925 $Y=0.805 $X2=0
+ $Y2=0
cc_480 N_SCE_c_505_n N_A_200_119#_c_2128_n 0.00479582f $X=2.89 $Y=0.18 $X2=0
+ $Y2=0
cc_481 N_SCE_M1042_g N_A_200_119#_c_2132_n 4.41958e-19 $X=0.925 $Y=2.69 $X2=0
+ $Y2=0
cc_482 N_SCE_M1042_g N_A_200_119#_c_2134_n 4.06466e-19 $X=0.925 $Y=2.69 $X2=0
+ $Y2=0
cc_483 N_SCE_M1010_g N_A_200_119#_c_2136_n 0.00572249f $X=2.965 $Y=0.805 $X2=0
+ $Y2=0
cc_484 N_SCE_M1010_g N_A_200_119#_c_2137_n 0.0272063f $X=2.965 $Y=0.805 $X2=0
+ $Y2=0
cc_485 N_SCE_M1010_g N_A_200_119#_c_2138_n 0.00576606f $X=2.965 $Y=0.805 $X2=0
+ $Y2=0
cc_486 N_SCE_M1010_g N_A_200_119#_c_2140_n 0.00310283f $X=2.965 $Y=0.805 $X2=0
+ $Y2=0
cc_487 N_SCE_M1012_g N_VGND_c_2359_n 0.00161717f $X=0.925 $Y=0.805 $X2=0 $Y2=0
cc_488 N_SCE_c_506_n N_VGND_c_2359_n 0.00971161f $X=1 $Y=0.18 $X2=0 $Y2=0
cc_489 N_SCE_c_505_n N_VGND_c_2360_n 0.0258591f $X=2.89 $Y=0.18 $X2=0 $Y2=0
cc_490 N_SCE_M1010_g N_VGND_c_2360_n 0.015224f $X=2.965 $Y=0.805 $X2=0 $Y2=0
cc_491 N_SCE_c_505_n N_VGND_c_2361_n 0.00991844f $X=2.89 $Y=0.18 $X2=0 $Y2=0
cc_492 N_SCE_c_505_n N_VGND_c_2369_n 0.013563f $X=2.89 $Y=0.18 $X2=0 $Y2=0
cc_493 N_SCE_c_506_n N_VGND_c_2373_n 0.0388559f $X=1 $Y=0.18 $X2=0 $Y2=0
cc_494 N_SCE_c_505_n N_VGND_c_2379_n 0.0609655f $X=2.89 $Y=0.18 $X2=0 $Y2=0
cc_495 N_SCE_c_506_n N_VGND_c_2379_n 0.010892f $X=1 $Y=0.18 $X2=0 $Y2=0
cc_496 N_CLK_N_c_576_n N_A_838_50#_c_622_n 5.6815e-19 $X=4.365 $Y=1.855 $X2=0
+ $Y2=0
cc_497 N_CLK_N_c_572_n N_A_838_50#_c_622_n 0.0369487f $X=4.025 $Y=1.035 $X2=0
+ $Y2=0
cc_498 N_CLK_N_c_573_n N_A_838_50#_c_622_n 0.00202757f $X=4.025 $Y=1.035 $X2=0
+ $Y2=0
cc_499 N_CLK_N_c_570_n N_A_838_50#_c_624_n 7.78245e-19 $X=4.025 $Y=1.375 $X2=0
+ $Y2=0
cc_500 N_CLK_N_c_569_n N_A_838_50#_c_625_n 0.00591454f $X=4.115 $Y=1.78 $X2=0
+ $Y2=0
cc_501 N_CLK_N_c_576_n N_A_838_50#_c_625_n 0.00730034f $X=4.365 $Y=1.855 $X2=0
+ $Y2=0
cc_502 N_CLK_N_M1015_g N_A_838_50#_c_634_n 0.00590992f $X=4.115 $Y=0.46 $X2=0
+ $Y2=0
cc_503 N_CLK_N_c_573_n N_A_838_50#_c_634_n 0.00221754f $X=4.025 $Y=1.035 $X2=0
+ $Y2=0
cc_504 N_CLK_N_c_572_n N_A_838_50#_c_635_n 7.78245e-19 $X=4.025 $Y=1.035 $X2=0
+ $Y2=0
cc_505 N_CLK_N_c_573_n N_A_838_50#_c_635_n 0.0541784f $X=4.025 $Y=1.035 $X2=0
+ $Y2=0
cc_506 N_CLK_N_M1015_g N_A_838_50#_c_636_n 0.0060129f $X=4.115 $Y=0.46 $X2=0
+ $Y2=0
cc_507 N_CLK_N_c_571_n N_A_838_50#_c_637_n 7.78245e-19 $X=4.025 $Y=1.54 $X2=0
+ $Y2=0
cc_508 N_CLK_N_c_576_n N_A_838_50#_c_637_n 0.00249866f $X=4.365 $Y=1.855 $X2=0
+ $Y2=0
cc_509 N_CLK_N_c_575_n N_VPWR_c_1943_n 0.00376577f $X=4.365 $Y=1.93 $X2=0 $Y2=0
cc_510 N_CLK_N_c_575_n N_VPWR_c_1960_n 2.23678e-19 $X=4.365 $Y=1.93 $X2=0 $Y2=0
cc_511 N_CLK_N_c_575_n N_A_200_119#_c_2140_n 0.00130692f $X=4.365 $Y=1.93 $X2=0
+ $Y2=0
cc_512 N_CLK_N_c_576_n N_A_200_119#_c_2140_n 7.92796e-19 $X=4.365 $Y=1.855 $X2=0
+ $Y2=0
cc_513 N_CLK_N_c_569_n N_A_200_119#_c_2141_n 0.00528978f $X=4.115 $Y=1.78 $X2=0
+ $Y2=0
cc_514 N_CLK_N_c_571_n N_A_200_119#_c_2141_n 0.00123144f $X=4.025 $Y=1.54 $X2=0
+ $Y2=0
cc_515 N_CLK_N_c_576_n N_A_200_119#_c_2141_n 0.0120747f $X=4.365 $Y=1.855 $X2=0
+ $Y2=0
cc_516 N_CLK_N_c_573_n N_A_200_119#_c_2141_n 0.0252679f $X=4.025 $Y=1.035 $X2=0
+ $Y2=0
cc_517 N_CLK_N_c_575_n N_A_200_119#_c_2143_n 0.028934f $X=4.365 $Y=1.93 $X2=0
+ $Y2=0
cc_518 N_CLK_N_c_576_n N_A_200_119#_c_2143_n 0.00512907f $X=4.365 $Y=1.855 $X2=0
+ $Y2=0
cc_519 N_CLK_N_c_575_n N_A_200_119#_c_2144_n 0.00576606f $X=4.365 $Y=1.93 $X2=0
+ $Y2=0
cc_520 N_CLK_N_c_575_n N_A_200_119#_c_2146_n 0.00261662f $X=4.365 $Y=1.93 $X2=0
+ $Y2=0
cc_521 N_CLK_N_M1015_g N_VGND_c_2361_n 0.0130079f $X=4.115 $Y=0.46 $X2=0 $Y2=0
cc_522 N_CLK_N_c_572_n N_VGND_c_2361_n 9.56064e-19 $X=4.025 $Y=1.035 $X2=0 $Y2=0
cc_523 N_CLK_N_c_573_n N_VGND_c_2361_n 0.0104884f $X=4.025 $Y=1.035 $X2=0 $Y2=0
cc_524 N_CLK_N_M1015_g N_VGND_c_2374_n 0.00534858f $X=4.115 $Y=0.46 $X2=0 $Y2=0
cc_525 N_CLK_N_M1015_g N_VGND_c_2379_n 0.0123058f $X=4.115 $Y=0.46 $X2=0 $Y2=0
cc_526 N_CLK_N_c_572_n N_VGND_c_2379_n 6.75321e-19 $X=4.025 $Y=1.035 $X2=0 $Y2=0
cc_527 N_A_838_50#_c_628_n N_A_1445_324#_M1000_d 0.00405136f $X=10.265 $Y=0.35
+ $X2=-0.19 $Y2=-0.245
cc_528 N_A_838_50#_c_626_n N_A_1445_324#_c_866_n 4.05318e-19 $X=7.21 $Y=1.215
+ $X2=0 $Y2=0
cc_529 N_A_838_50#_c_627_n N_A_1445_324#_c_866_n 0.0090932f $X=7.21 $Y=1.215
+ $X2=0 $Y2=0
cc_530 N_A_838_50#_M1028_g N_A_1445_324#_M1040_g 0.0190128f $X=7.12 $Y=0.73
+ $X2=0 $Y2=0
cc_531 N_A_838_50#_c_626_n N_A_1445_324#_M1040_g 0.00387156f $X=7.21 $Y=1.215
+ $X2=0 $Y2=0
cc_532 N_A_838_50#_c_627_n N_A_1445_324#_M1040_g 0.017189f $X=7.21 $Y=1.215
+ $X2=0 $Y2=0
cc_533 N_A_838_50#_c_673_p N_A_1445_324#_M1040_g 0.014479f $X=8.385 $Y=0.79
+ $X2=0 $Y2=0
cc_534 N_A_838_50#_c_674_p N_A_1445_324#_M1040_g 0.00394726f $X=8.47 $Y=0.705
+ $X2=0 $Y2=0
cc_535 N_A_838_50#_c_630_n N_A_1445_324#_M1027_g 0.00502057f $X=10.35 $Y=1.085
+ $X2=0 $Y2=0
cc_536 N_A_838_50#_c_631_n N_A_1445_324#_M1027_g 0.0149519f $X=11.12 $Y=1.17
+ $X2=0 $Y2=0
cc_537 N_A_838_50#_c_633_n N_A_1445_324#_M1027_g 0.00537674f $X=11.205 $Y=1.675
+ $X2=0 $Y2=0
cc_538 N_A_838_50#_c_638_n N_A_1445_324#_M1027_g 0.020664f $X=11.365 $Y=1.51
+ $X2=0 $Y2=0
cc_539 N_A_838_50#_c_639_n N_A_1445_324#_M1027_g 0.0290031f $X=11.365 $Y=1.345
+ $X2=0 $Y2=0
cc_540 N_A_838_50#_c_632_n N_A_1445_324#_c_871_n 7.47982e-19 $X=10.435 $Y=1.17
+ $X2=0 $Y2=0
cc_541 N_A_838_50#_c_631_n N_A_1445_324#_c_872_n 0.0305714f $X=11.12 $Y=1.17
+ $X2=0 $Y2=0
cc_542 N_A_838_50#_c_632_n N_A_1445_324#_c_872_n 0.010315f $X=10.435 $Y=1.17
+ $X2=0 $Y2=0
cc_543 N_A_838_50#_c_633_n N_A_1445_324#_c_872_n 0.0196132f $X=11.205 $Y=1.675
+ $X2=0 $Y2=0
cc_544 N_A_838_50#_c_648_n N_A_1445_324#_c_872_n 0.0037127f $X=11.205 $Y=2.895
+ $X2=0 $Y2=0
cc_545 N_A_838_50#_c_638_n N_A_1445_324#_c_872_n 2.33631e-19 $X=11.365 $Y=1.51
+ $X2=0 $Y2=0
cc_546 N_A_838_50#_c_631_n N_A_1445_324#_c_873_n 0.00525942f $X=11.12 $Y=1.17
+ $X2=0 $Y2=0
cc_547 N_A_838_50#_c_648_n N_A_1445_324#_c_873_n 0.0173763f $X=11.205 $Y=2.895
+ $X2=0 $Y2=0
cc_548 N_A_838_50#_c_630_n N_A_1445_324#_c_874_n 0.00109361f $X=10.35 $Y=1.085
+ $X2=0 $Y2=0
cc_549 N_A_838_50#_c_632_n N_A_1445_324#_c_874_n 0.00586392f $X=10.435 $Y=1.17
+ $X2=0 $Y2=0
cc_550 N_A_838_50#_c_628_n N_SET_B_M1035_g 0.0125497f $X=10.265 $Y=0.35 $X2=0
+ $Y2=0
cc_551 N_A_838_50#_c_631_n N_SET_B_c_1008_n 0.0315496f $X=11.12 $Y=1.17 $X2=0
+ $Y2=0
cc_552 N_A_838_50#_c_632_n N_SET_B_c_1008_n 0.0111681f $X=10.435 $Y=1.17 $X2=0
+ $Y2=0
cc_553 N_A_838_50#_c_633_n N_SET_B_c_1008_n 0.0365917f $X=11.205 $Y=1.675 $X2=0
+ $Y2=0
cc_554 N_A_838_50#_c_651_n N_SET_B_c_1008_n 0.0126936f $X=12.265 $Y=1.865 $X2=0
+ $Y2=0
cc_555 N_A_838_50#_c_638_n N_SET_B_c_1008_n 0.00100787f $X=11.365 $Y=1.51 $X2=0
+ $Y2=0
cc_556 N_A_838_50#_c_639_n N_SET_B_c_1008_n 0.007222f $X=11.365 $Y=1.345 $X2=0
+ $Y2=0
cc_557 N_A_838_50#_c_628_n N_SET_B_c_1010_n 0.00343517f $X=10.265 $Y=0.35 $X2=0
+ $Y2=0
cc_558 N_A_838_50#_c_651_n N_SET_B_c_1012_n 0.00253088f $X=12.265 $Y=1.865 $X2=0
+ $Y2=0
cc_559 N_A_838_50#_c_673_p N_SET_B_c_1013_n 0.00205173f $X=8.385 $Y=0.79 $X2=0
+ $Y2=0
cc_560 N_A_838_50#_c_628_n N_A_1295_379#_M1000_g 0.0103183f $X=10.265 $Y=0.35
+ $X2=0 $Y2=0
cc_561 N_A_838_50#_c_619_n N_A_1295_379#_c_1149_n 0.00704409f $X=7.045 $Y=0.18
+ $X2=0 $Y2=0
cc_562 N_A_838_50#_M1033_g N_A_1295_379#_c_1149_n 9.36938e-19 $X=6.4 $Y=2.105
+ $X2=0 $Y2=0
cc_563 N_A_838_50#_M1028_g N_A_1295_379#_c_1149_n 0.0106295f $X=7.12 $Y=0.73
+ $X2=0 $Y2=0
cc_564 N_A_838_50#_c_626_n N_A_1295_379#_c_1149_n 0.0375185f $X=7.21 $Y=1.215
+ $X2=0 $Y2=0
cc_565 N_A_838_50#_c_705_p N_A_1295_379#_c_1149_n 0.0133994f $X=7.31 $Y=0.79
+ $X2=0 $Y2=0
cc_566 N_A_838_50#_c_626_n N_A_1295_379#_c_1161_n 0.00902988f $X=7.21 $Y=1.215
+ $X2=0 $Y2=0
cc_567 N_A_838_50#_c_627_n N_A_1295_379#_c_1161_n 0.0013276f $X=7.21 $Y=1.215
+ $X2=0 $Y2=0
cc_568 N_A_838_50#_c_626_n N_A_1295_379#_c_1150_n 0.0109374f $X=7.21 $Y=1.215
+ $X2=0 $Y2=0
cc_569 N_A_838_50#_c_627_n N_A_1295_379#_c_1150_n 9.99763e-19 $X=7.21 $Y=1.215
+ $X2=0 $Y2=0
cc_570 N_A_838_50#_c_673_p N_A_1295_379#_c_1151_n 0.0506393f $X=8.385 $Y=0.79
+ $X2=0 $Y2=0
cc_571 N_A_838_50#_c_626_n N_A_1295_379#_c_1152_n 0.0135289f $X=7.21 $Y=1.215
+ $X2=0 $Y2=0
cc_572 N_A_838_50#_c_627_n N_A_1295_379#_c_1152_n 0.00127177f $X=7.21 $Y=1.215
+ $X2=0 $Y2=0
cc_573 N_A_838_50#_c_673_p N_A_1295_379#_c_1152_n 0.0112499f $X=8.385 $Y=0.79
+ $X2=0 $Y2=0
cc_574 N_A_838_50#_M1033_g N_A_1295_379#_c_1165_n 0.00253632f $X=6.4 $Y=2.105
+ $X2=0 $Y2=0
cc_575 N_A_838_50#_M1033_g N_A_995_66#_c_1275_n 0.00950983f $X=6.4 $Y=2.105
+ $X2=0 $Y2=0
cc_576 N_A_838_50#_c_619_n N_A_995_66#_M1005_g 0.00895007f $X=7.045 $Y=0.18
+ $X2=0 $Y2=0
cc_577 N_A_838_50#_M1028_g N_A_995_66#_M1005_g 0.0107685f $X=7.12 $Y=0.73 $X2=0
+ $Y2=0
cc_578 N_A_838_50#_M1033_g N_A_995_66#_c_1278_n 2.92137e-19 $X=6.4 $Y=2.105
+ $X2=0 $Y2=0
cc_579 N_A_838_50#_c_627_n N_A_995_66#_c_1278_n 0.00220046f $X=7.21 $Y=1.215
+ $X2=0 $Y2=0
cc_580 N_A_838_50#_M1033_g N_A_995_66#_M1034_g 0.0221327f $X=6.4 $Y=2.105 $X2=0
+ $Y2=0
cc_581 N_A_838_50#_c_644_n N_A_995_66#_c_1289_n 0.0100606f $X=11.93 $Y=2.455
+ $X2=0 $Y2=0
cc_582 N_A_838_50#_c_650_n N_A_995_66#_c_1289_n 0.00332551f $X=11.29 $Y=2.98
+ $X2=0 $Y2=0
cc_583 N_A_838_50#_c_641_n N_A_995_66#_c_1290_n 0.0221327f $X=6.325 $Y=3.135
+ $X2=0 $Y2=0
cc_584 N_A_838_50#_c_645_n N_A_995_66#_M1038_g 0.0100606f $X=12.265 $Y=2.305
+ $X2=0 $Y2=0
cc_585 N_A_838_50#_c_649_n N_A_995_66#_M1038_g 0.0151989f $X=12.1 $Y=2.98 $X2=0
+ $Y2=0
cc_586 N_A_838_50#_c_651_n N_A_995_66#_M1038_g 2.93889e-19 $X=12.265 $Y=1.865
+ $X2=0 $Y2=0
cc_587 N_A_838_50#_c_652_n N_A_995_66#_M1038_g 0.00258692f $X=12.265 $Y=1.865
+ $X2=0 $Y2=0
cc_588 N_A_838_50#_c_645_n N_A_995_66#_c_1292_n 0.00214523f $X=12.265 $Y=2.305
+ $X2=0 $Y2=0
cc_589 N_A_838_50#_c_633_n N_A_995_66#_c_1293_n 0.00119508f $X=11.205 $Y=1.675
+ $X2=0 $Y2=0
cc_590 N_A_838_50#_c_648_n N_A_995_66#_c_1293_n 0.0077349f $X=11.205 $Y=2.895
+ $X2=0 $Y2=0
cc_591 N_A_838_50#_c_638_n N_A_995_66#_c_1293_n 0.0102687f $X=11.365 $Y=1.51
+ $X2=0 $Y2=0
cc_592 N_A_838_50#_c_648_n N_A_995_66#_c_1279_n 0.00131551f $X=11.205 $Y=2.895
+ $X2=0 $Y2=0
cc_593 N_A_838_50#_c_651_n N_A_995_66#_c_1279_n 0.00122995f $X=12.265 $Y=1.865
+ $X2=0 $Y2=0
cc_594 N_A_838_50#_c_652_n N_A_995_66#_c_1279_n 0.0218791f $X=12.265 $Y=1.865
+ $X2=0 $Y2=0
cc_595 N_A_838_50#_c_639_n N_A_995_66#_c_1280_n 0.0144238f $X=11.365 $Y=1.345
+ $X2=0 $Y2=0
cc_596 N_A_838_50#_c_633_n N_A_995_66#_c_1282_n 4.04794e-19 $X=11.205 $Y=1.675
+ $X2=0 $Y2=0
cc_597 N_A_838_50#_c_638_n N_A_995_66#_c_1282_n 0.0213156f $X=11.365 $Y=1.51
+ $X2=0 $Y2=0
cc_598 N_A_838_50#_c_639_n N_A_995_66#_c_1282_n 0.00192706f $X=11.365 $Y=1.345
+ $X2=0 $Y2=0
cc_599 N_A_838_50#_M1039_g N_A_995_66#_c_1283_n 0.0127128f $X=5.345 $Y=0.54
+ $X2=0 $Y2=0
cc_600 N_A_838_50#_c_622_n N_A_995_66#_c_1283_n 0.0283427f $X=5.27 $Y=1.205
+ $X2=0 $Y2=0
cc_601 N_A_838_50#_c_623_n N_A_995_66#_c_1283_n 0.0202028f $X=5.345 $Y=1.205
+ $X2=0 $Y2=0
cc_602 N_A_838_50#_c_634_n N_A_995_66#_c_1283_n 0.0251394f $X=4.33 $Y=0.475
+ $X2=0 $Y2=0
cc_603 N_A_838_50#_c_635_n N_A_995_66#_c_1283_n 0.0322506f $X=4.595 $Y=1.035
+ $X2=0 $Y2=0
cc_604 N_A_838_50#_M1018_g N_A_995_66#_c_1295_n 0.0239057f $X=5.345 $Y=2.155
+ $X2=0 $Y2=0
cc_605 N_A_838_50#_c_625_n N_A_995_66#_c_1295_n 0.0350016f $X=4.58 $Y=2.2 $X2=0
+ $Y2=0
cc_606 N_A_838_50#_M1018_g N_A_995_66#_c_1284_n 0.00659585f $X=5.345 $Y=2.155
+ $X2=0 $Y2=0
cc_607 N_A_838_50#_c_623_n N_A_995_66#_c_1284_n 0.0102875f $X=5.345 $Y=1.205
+ $X2=0 $Y2=0
cc_608 N_A_838_50#_M1018_g N_A_995_66#_c_1285_n 0.00304296f $X=5.345 $Y=2.155
+ $X2=0 $Y2=0
cc_609 N_A_838_50#_c_622_n N_A_995_66#_c_1285_n 0.0160963f $X=5.27 $Y=1.205
+ $X2=0 $Y2=0
cc_610 N_A_838_50#_c_623_n N_A_995_66#_c_1285_n 9.78204e-19 $X=5.345 $Y=1.205
+ $X2=0 $Y2=0
cc_611 N_A_838_50#_c_624_n N_A_995_66#_c_1285_n 0.0246945f $X=4.567 $Y=1.348
+ $X2=0 $Y2=0
cc_612 N_A_838_50#_c_623_n N_A_995_66#_c_1286_n 0.017302f $X=5.345 $Y=1.205
+ $X2=0 $Y2=0
cc_613 N_A_838_50#_c_651_n N_A_2449_137#_c_1399_n 0.00134249f $X=12.265 $Y=1.865
+ $X2=0 $Y2=0
cc_614 N_A_838_50#_c_652_n N_A_2449_137#_c_1399_n 0.01029f $X=12.265 $Y=1.865
+ $X2=0 $Y2=0
cc_615 N_A_838_50#_c_644_n N_A_2449_137#_M1037_g 0.00621587f $X=11.93 $Y=2.455
+ $X2=0 $Y2=0
cc_616 N_A_838_50#_c_649_n N_A_2449_137#_M1037_g 0.00252975f $X=12.1 $Y=2.98
+ $X2=0 $Y2=0
cc_617 N_A_838_50#_c_651_n N_A_2449_137#_M1037_g 0.00713085f $X=12.265 $Y=1.865
+ $X2=0 $Y2=0
cc_618 N_A_838_50#_c_652_n N_A_2449_137#_M1037_g 0.00959621f $X=12.265 $Y=1.865
+ $X2=0 $Y2=0
cc_619 N_A_838_50#_c_651_n N_A_2449_137#_c_1416_n 0.02209f $X=12.265 $Y=1.865
+ $X2=0 $Y2=0
cc_620 N_A_838_50#_c_652_n N_A_2449_137#_c_1416_n 0.00114003f $X=12.265 $Y=1.865
+ $X2=0 $Y2=0
cc_621 N_A_838_50#_c_651_n N_A_2449_137#_c_1417_n 4.14293e-19 $X=12.265 $Y=1.865
+ $X2=0 $Y2=0
cc_622 N_A_838_50#_c_651_n N_A_2449_137#_c_1411_n 0.00151562f $X=12.265 $Y=1.865
+ $X2=0 $Y2=0
cc_623 N_A_838_50#_c_652_n N_A_2449_137#_c_1411_n 0.0372091f $X=12.265 $Y=1.865
+ $X2=0 $Y2=0
cc_624 N_A_838_50#_c_649_n N_A_2299_119#_M1038_d 0.00267852f $X=12.1 $Y=2.98
+ $X2=0 $Y2=0
cc_625 N_A_838_50#_c_633_n N_A_2299_119#_c_1584_n 0.00255382f $X=11.205 $Y=1.675
+ $X2=0 $Y2=0
cc_626 N_A_838_50#_c_639_n N_A_2299_119#_c_1584_n 0.0148976f $X=11.365 $Y=1.345
+ $X2=0 $Y2=0
cc_627 N_A_838_50#_c_644_n N_A_2299_119#_c_1590_n 0.00715527f $X=11.93 $Y=2.455
+ $X2=0 $Y2=0
cc_628 N_A_838_50#_c_645_n N_A_2299_119#_c_1590_n 0.00521228f $X=12.265 $Y=2.305
+ $X2=0 $Y2=0
cc_629 N_A_838_50#_c_633_n N_A_2299_119#_c_1590_n 0.00229002f $X=11.205 $Y=1.675
+ $X2=0 $Y2=0
cc_630 N_A_838_50#_c_648_n N_A_2299_119#_c_1590_n 0.0227323f $X=11.205 $Y=2.895
+ $X2=0 $Y2=0
cc_631 N_A_838_50#_c_649_n N_A_2299_119#_c_1590_n 0.0209848f $X=12.1 $Y=2.98
+ $X2=0 $Y2=0
cc_632 N_A_838_50#_c_633_n N_A_2299_119#_c_1585_n 0.0275506f $X=11.205 $Y=1.675
+ $X2=0 $Y2=0
cc_633 N_A_838_50#_c_648_n N_A_2299_119#_c_1585_n 0.0153054f $X=11.205 $Y=2.895
+ $X2=0 $Y2=0
cc_634 N_A_838_50#_c_651_n N_A_2299_119#_c_1585_n 0.0634032f $X=12.265 $Y=1.865
+ $X2=0 $Y2=0
cc_635 N_A_838_50#_c_652_n N_A_2299_119#_c_1585_n 0.00368182f $X=12.265 $Y=1.865
+ $X2=0 $Y2=0
cc_636 N_A_838_50#_c_638_n N_A_2299_119#_c_1585_n 9.68817e-19 $X=11.365 $Y=1.51
+ $X2=0 $Y2=0
cc_637 N_A_838_50#_c_639_n N_A_2299_119#_c_1585_n 8.16432e-19 $X=11.365 $Y=1.345
+ $X2=0 $Y2=0
cc_638 N_A_838_50#_c_628_n N_A_1926_21#_M1008_g 0.0106943f $X=10.265 $Y=0.35
+ $X2=0 $Y2=0
cc_639 N_A_838_50#_c_630_n N_A_1926_21#_M1008_g 0.00482903f $X=10.35 $Y=1.085
+ $X2=0 $Y2=0
cc_640 N_A_838_50#_c_628_n N_A_1926_21#_c_1682_n 0.0134096f $X=10.265 $Y=0.35
+ $X2=0 $Y2=0
cc_641 N_A_838_50#_c_639_n N_A_1926_21#_c_1682_n 0.0103003f $X=11.365 $Y=1.345
+ $X2=0 $Y2=0
cc_642 N_A_838_50#_c_628_n N_A_1926_21#_c_1684_n 0.00435005f $X=10.265 $Y=0.35
+ $X2=0 $Y2=0
cc_643 N_A_838_50#_c_630_n N_A_1926_21#_c_1684_n 0.00440571f $X=10.35 $Y=1.085
+ $X2=0 $Y2=0
cc_644 N_A_838_50#_c_632_n N_A_1926_21#_c_1684_n 0.00559162f $X=10.435 $Y=1.17
+ $X2=0 $Y2=0
cc_645 N_A_838_50#_c_632_n N_A_1926_21#_M1003_g 0.00296837f $X=10.435 $Y=1.17
+ $X2=0 $Y2=0
cc_646 N_A_838_50#_M1018_g N_VPWR_c_1944_n 0.00669734f $X=5.345 $Y=2.155 $X2=0
+ $Y2=0
cc_647 N_A_838_50#_c_641_n N_VPWR_c_1944_n 0.0244196f $X=6.325 $Y=3.135 $X2=0
+ $Y2=0
cc_648 N_A_838_50#_M1033_g N_VPWR_c_1944_n 0.00984036f $X=6.4 $Y=2.105 $X2=0
+ $Y2=0
cc_649 N_A_838_50#_c_648_n N_VPWR_c_1946_n 0.037359f $X=11.205 $Y=2.895 $X2=0
+ $Y2=0
cc_650 N_A_838_50#_c_650_n N_VPWR_c_1946_n 0.00755092f $X=11.29 $Y=2.98 $X2=0
+ $Y2=0
cc_651 N_A_838_50#_c_649_n N_VPWR_c_1947_n 0.00535867f $X=12.1 $Y=2.98 $X2=0
+ $Y2=0
cc_652 N_A_838_50#_c_651_n N_VPWR_c_1947_n 0.0119115f $X=12.265 $Y=1.865 $X2=0
+ $Y2=0
cc_653 N_A_838_50#_c_642_n N_VPWR_c_1960_n 0.00726972f $X=5.42 $Y=3.135 $X2=0
+ $Y2=0
cc_654 N_A_838_50#_c_641_n N_VPWR_c_1961_n 0.0240383f $X=6.325 $Y=3.135 $X2=0
+ $Y2=0
cc_655 N_A_838_50#_c_644_n N_VPWR_c_1962_n 0.00392127f $X=11.93 $Y=2.455 $X2=0
+ $Y2=0
cc_656 N_A_838_50#_c_649_n N_VPWR_c_1962_n 0.0704502f $X=12.1 $Y=2.98 $X2=0
+ $Y2=0
cc_657 N_A_838_50#_c_650_n N_VPWR_c_1962_n 0.0114583f $X=11.29 $Y=2.98 $X2=0
+ $Y2=0
cc_658 N_A_838_50#_c_641_n N_VPWR_c_1940_n 0.0264759f $X=6.325 $Y=3.135 $X2=0
+ $Y2=0
cc_659 N_A_838_50#_c_642_n N_VPWR_c_1940_n 0.00663227f $X=5.42 $Y=3.135 $X2=0
+ $Y2=0
cc_660 N_A_838_50#_c_644_n N_VPWR_c_1940_n 0.00542671f $X=11.93 $Y=2.455 $X2=0
+ $Y2=0
cc_661 N_A_838_50#_c_649_n N_VPWR_c_1940_n 0.0420089f $X=12.1 $Y=2.98 $X2=0
+ $Y2=0
cc_662 N_A_838_50#_c_650_n N_VPWR_c_1940_n 0.00589978f $X=11.29 $Y=2.98 $X2=0
+ $Y2=0
cc_663 N_A_838_50#_c_625_n N_A_200_119#_c_2141_n 0.0137113f $X=4.58 $Y=2.2 $X2=0
+ $Y2=0
cc_664 N_A_838_50#_c_625_n N_A_200_119#_c_2143_n 0.0337157f $X=4.58 $Y=2.2 $X2=0
+ $Y2=0
cc_665 N_A_838_50#_M1018_g N_A_200_119#_c_2144_n 0.00634342f $X=5.345 $Y=2.155
+ $X2=0 $Y2=0
cc_666 N_A_838_50#_c_642_n N_A_200_119#_c_2144_n 3.7398e-19 $X=5.42 $Y=3.135
+ $X2=0 $Y2=0
cc_667 N_A_838_50#_c_625_n N_A_200_119#_c_2144_n 0.0198711f $X=4.58 $Y=2.2 $X2=0
+ $Y2=0
cc_668 N_A_838_50#_M1018_g N_A_200_119#_c_2146_n 0.0163885f $X=5.345 $Y=2.155
+ $X2=0 $Y2=0
cc_669 N_A_838_50#_c_625_n N_A_200_119#_c_2146_n 0.0101821f $X=4.58 $Y=2.2 $X2=0
+ $Y2=0
cc_670 N_A_838_50#_M1018_g N_A_200_119#_c_2147_n 0.0127336f $X=5.345 $Y=2.155
+ $X2=0 $Y2=0
cc_671 N_A_838_50#_c_641_n N_A_200_119#_c_2147_n 0.0116989f $X=6.325 $Y=3.135
+ $X2=0 $Y2=0
cc_672 N_A_838_50#_M1033_g N_A_200_119#_c_2147_n 0.00825997f $X=6.4 $Y=2.105
+ $X2=0 $Y2=0
cc_673 N_A_838_50#_M1018_g N_A_200_119#_c_2148_n 0.00356962f $X=5.345 $Y=2.155
+ $X2=0 $Y2=0
cc_674 N_A_838_50#_c_625_n N_A_200_119#_c_2148_n 0.00850606f $X=4.58 $Y=2.2
+ $X2=0 $Y2=0
cc_675 N_A_838_50#_M1018_g N_A_200_119#_c_2149_n 0.010657f $X=5.345 $Y=2.155
+ $X2=0 $Y2=0
cc_676 N_A_838_50#_M1033_g N_A_200_119#_c_2149_n 0.0024289f $X=6.4 $Y=2.105
+ $X2=0 $Y2=0
cc_677 N_A_838_50#_M1033_g N_A_200_119#_c_2150_n 0.00342448f $X=6.4 $Y=2.105
+ $X2=0 $Y2=0
cc_678 N_A_838_50#_M1033_g N_A_200_119#_c_2130_n 0.00365546f $X=6.4 $Y=2.105
+ $X2=0 $Y2=0
cc_679 N_A_838_50#_M1039_g N_A_200_119#_c_2131_n 0.00811556f $X=5.345 $Y=0.54
+ $X2=0 $Y2=0
cc_680 N_A_838_50#_c_619_n N_A_200_119#_c_2131_n 0.00601704f $X=7.045 $Y=0.18
+ $X2=0 $Y2=0
cc_681 N_A_838_50#_c_648_n A_2198_379# 0.0198147f $X=11.205 $Y=2.895 $X2=-0.19
+ $Y2=-0.245
cc_682 N_A_838_50#_c_650_n A_2198_379# 0.00172167f $X=11.29 $Y=2.98 $X2=-0.19
+ $Y2=-0.245
cc_683 N_A_838_50#_c_649_n A_2401_506# 0.0021694f $X=12.1 $Y=2.98 $X2=-0.19
+ $Y2=-0.245
cc_684 N_A_838_50#_c_651_n A_2401_506# 0.0134456f $X=12.265 $Y=1.865 $X2=-0.19
+ $Y2=-0.245
cc_685 N_A_838_50#_c_673_p N_VGND_M1040_d 0.0251424f $X=8.385 $Y=0.79 $X2=0
+ $Y2=0
cc_686 N_A_838_50#_c_674_p N_VGND_M1040_d 0.00520668f $X=8.47 $Y=0.705 $X2=0
+ $Y2=0
cc_687 N_A_838_50#_c_629_n N_VGND_M1040_d 0.00182835f $X=8.555 $Y=0.35 $X2=0
+ $Y2=0
cc_688 N_A_838_50#_c_631_n N_VGND_M1027_s 0.00501179f $X=11.12 $Y=1.17 $X2=0
+ $Y2=0
cc_689 N_A_838_50#_c_634_n N_VGND_c_2361_n 0.0163242f $X=4.33 $Y=0.475 $X2=0
+ $Y2=0
cc_690 N_A_838_50#_M1039_g N_VGND_c_2362_n 0.00829723f $X=5.345 $Y=0.54 $X2=0
+ $Y2=0
cc_691 N_A_838_50#_c_619_n N_VGND_c_2362_n 0.0241326f $X=7.045 $Y=0.18 $X2=0
+ $Y2=0
cc_692 N_A_838_50#_c_619_n N_VGND_c_2363_n 0.00525646f $X=7.045 $Y=0.18 $X2=0
+ $Y2=0
cc_693 N_A_838_50#_c_673_p N_VGND_c_2363_n 0.0242832f $X=8.385 $Y=0.79 $X2=0
+ $Y2=0
cc_694 N_A_838_50#_c_674_p N_VGND_c_2363_n 0.00655701f $X=8.47 $Y=0.705 $X2=0
+ $Y2=0
cc_695 N_A_838_50#_c_629_n N_VGND_c_2363_n 0.013989f $X=8.555 $Y=0.35 $X2=0
+ $Y2=0
cc_696 N_A_838_50#_c_628_n N_VGND_c_2364_n 0.0141601f $X=10.265 $Y=0.35 $X2=0
+ $Y2=0
cc_697 N_A_838_50#_c_630_n N_VGND_c_2364_n 0.0345265f $X=10.35 $Y=1.085 $X2=0
+ $Y2=0
cc_698 N_A_838_50#_c_631_n N_VGND_c_2364_n 0.0135595f $X=11.12 $Y=1.17 $X2=0
+ $Y2=0
cc_699 N_A_838_50#_c_639_n N_VGND_c_2364_n 0.00153768f $X=11.365 $Y=1.345 $X2=0
+ $Y2=0
cc_700 N_A_838_50#_c_620_n N_VGND_c_2374_n 0.00736894f $X=5.42 $Y=0.18 $X2=0
+ $Y2=0
cc_701 N_A_838_50#_c_634_n N_VGND_c_2374_n 0.0228286f $X=4.33 $Y=0.475 $X2=0
+ $Y2=0
cc_702 N_A_838_50#_c_619_n N_VGND_c_2375_n 0.0411899f $X=7.045 $Y=0.18 $X2=0
+ $Y2=0
cc_703 N_A_838_50#_c_673_p N_VGND_c_2375_n 0.00753747f $X=8.385 $Y=0.79 $X2=0
+ $Y2=0
cc_704 N_A_838_50#_c_705_p N_VGND_c_2375_n 0.00373503f $X=7.31 $Y=0.79 $X2=0
+ $Y2=0
cc_705 N_A_838_50#_c_673_p N_VGND_c_2376_n 0.00269352f $X=8.385 $Y=0.79 $X2=0
+ $Y2=0
cc_706 N_A_838_50#_c_628_n N_VGND_c_2376_n 0.11379f $X=10.265 $Y=0.35 $X2=0
+ $Y2=0
cc_707 N_A_838_50#_c_629_n N_VGND_c_2376_n 0.0113687f $X=8.555 $Y=0.35 $X2=0
+ $Y2=0
cc_708 N_A_838_50#_c_619_n N_VGND_c_2379_n 0.0563018f $X=7.045 $Y=0.18 $X2=0
+ $Y2=0
cc_709 N_A_838_50#_c_620_n N_VGND_c_2379_n 0.0109396f $X=5.42 $Y=0.18 $X2=0
+ $Y2=0
cc_710 N_A_838_50#_c_622_n N_VGND_c_2379_n 0.0074388f $X=5.27 $Y=1.205 $X2=0
+ $Y2=0
cc_711 N_A_838_50#_c_673_p N_VGND_c_2379_n 0.0213925f $X=8.385 $Y=0.79 $X2=0
+ $Y2=0
cc_712 N_A_838_50#_c_705_p N_VGND_c_2379_n 0.00685961f $X=7.31 $Y=0.79 $X2=0
+ $Y2=0
cc_713 N_A_838_50#_c_628_n N_VGND_c_2379_n 0.0657755f $X=10.265 $Y=0.35 $X2=0
+ $Y2=0
cc_714 N_A_838_50#_c_629_n N_VGND_c_2379_n 0.00655847f $X=8.555 $Y=0.35 $X2=0
+ $Y2=0
cc_715 N_A_838_50#_c_634_n N_VGND_c_2379_n 0.0144161f $X=4.33 $Y=0.475 $X2=0
+ $Y2=0
cc_716 N_A_838_50#_c_639_n N_VGND_c_2379_n 9.39239e-19 $X=11.365 $Y=1.345 $X2=0
+ $Y2=0
cc_717 N_A_838_50#_c_626_n A_1439_104# 8.72273e-19 $X=7.21 $Y=1.215 $X2=-0.19
+ $Y2=-0.245
cc_718 N_A_838_50#_c_673_p A_1439_104# 0.0110593f $X=8.385 $Y=0.79 $X2=-0.19
+ $Y2=-0.245
cc_719 N_A_838_50#_c_705_p A_1439_104# 0.00112373f $X=7.31 $Y=0.79 $X2=-0.19
+ $Y2=-0.245
cc_720 N_A_838_50#_c_628_n N_A_1752_60#_M1035_d 0.00185121f $X=10.265 $Y=0.35
+ $X2=-0.19 $Y2=-0.245
cc_721 N_A_838_50#_c_628_n N_A_1752_60#_M1008_d 0.00288258f $X=10.265 $Y=0.35
+ $X2=0 $Y2=0
cc_722 N_A_838_50#_c_628_n N_A_1752_60#_c_2540_n 0.0689952f $X=10.265 $Y=0.35
+ $X2=0 $Y2=0
cc_723 N_A_838_50#_c_630_n N_A_1752_60#_c_2537_n 0.0205142f $X=10.35 $Y=1.085
+ $X2=0 $Y2=0
cc_724 N_A_838_50#_c_631_n A_2198_119# 0.0027472f $X=11.12 $Y=1.17 $X2=-0.19
+ $Y2=-0.245
cc_725 N_A_838_50#_c_633_n A_2198_119# 0.00810107f $X=11.205 $Y=1.675 $X2=-0.19
+ $Y2=-0.245
cc_726 N_A_1445_324#_c_869_n N_SET_B_M1030_g 0.00381373f $X=7.94 $Y=1.57 $X2=0
+ $Y2=0
cc_727 N_A_1445_324#_c_870_n N_SET_B_M1030_g 0.00507869f $X=7.94 $Y=1.57 $X2=0
+ $Y2=0
cc_728 N_A_1445_324#_c_912_p N_SET_B_M1030_g 0.0192094f $X=9.525 $Y=2.025 $X2=0
+ $Y2=0
cc_729 N_A_1445_324#_c_885_n N_SET_B_M1030_g 0.0145499f $X=9.69 $Y=2.08 $X2=0
+ $Y2=0
cc_730 N_A_1445_324#_M1000_d N_SET_B_c_1008_n 3.02582e-19 $X=9.195 $Y=0.3 $X2=0
+ $Y2=0
cc_731 N_A_1445_324#_M1027_g N_SET_B_c_1008_n 0.00477151f $X=10.915 $Y=0.915
+ $X2=0 $Y2=0
cc_732 N_A_1445_324#_c_912_p N_SET_B_c_1008_n 0.00137022f $X=9.525 $Y=2.025
+ $X2=0 $Y2=0
cc_733 N_A_1445_324#_c_871_n N_SET_B_c_1008_n 0.0160926f $X=9.77 $Y=1.435 $X2=0
+ $Y2=0
cc_734 N_A_1445_324#_c_872_n N_SET_B_c_1008_n 0.0358898f $X=10.775 $Y=1.56 $X2=0
+ $Y2=0
cc_735 N_A_1445_324#_c_873_n N_SET_B_c_1008_n 0.00603145f $X=10.775 $Y=1.56
+ $X2=0 $Y2=0
cc_736 N_A_1445_324#_c_874_n N_SET_B_c_1008_n 0.0157749f $X=9.41 $Y=1.13 $X2=0
+ $Y2=0
cc_737 N_A_1445_324#_c_885_n N_SET_B_c_1008_n 0.00587717f $X=9.69 $Y=2.08 $X2=0
+ $Y2=0
cc_738 N_A_1445_324#_c_874_n N_SET_B_c_1009_n 0.00131878f $X=9.41 $Y=1.13 $X2=0
+ $Y2=0
cc_739 N_A_1445_324#_c_874_n N_SET_B_c_1010_n 0.00900086f $X=9.41 $Y=1.13 $X2=0
+ $Y2=0
cc_740 N_A_1445_324#_c_871_n N_A_1295_379#_M1000_g 0.00311788f $X=9.77 $Y=1.435
+ $X2=0 $Y2=0
cc_741 N_A_1445_324#_c_874_n N_A_1295_379#_M1000_g 0.00553667f $X=9.41 $Y=1.13
+ $X2=0 $Y2=0
cc_742 N_A_1445_324#_c_912_p N_A_1295_379#_c_1147_n 6.26426e-19 $X=9.525
+ $Y=2.025 $X2=0 $Y2=0
cc_743 N_A_1445_324#_c_882_n N_A_1295_379#_c_1147_n 0.00382197f $X=9.77 $Y=1.915
+ $X2=0 $Y2=0
cc_744 N_A_1445_324#_c_872_n N_A_1295_379#_c_1147_n 0.0101093f $X=10.775 $Y=1.56
+ $X2=0 $Y2=0
cc_745 N_A_1445_324#_c_874_n N_A_1295_379#_c_1147_n 0.0036871f $X=9.41 $Y=1.13
+ $X2=0 $Y2=0
cc_746 N_A_1445_324#_c_885_n N_A_1295_379#_c_1147_n 0.00650665f $X=9.69 $Y=2.08
+ $X2=0 $Y2=0
cc_747 N_A_1445_324#_c_875_n N_A_1295_379#_c_1147_n 0.00686361f $X=9.77 $Y=1.58
+ $X2=0 $Y2=0
cc_748 N_A_1445_324#_c_912_p N_A_1295_379#_c_1148_n 0.00218686f $X=9.525
+ $Y=2.025 $X2=0 $Y2=0
cc_749 N_A_1445_324#_c_874_n N_A_1295_379#_c_1148_n 0.0017102f $X=9.41 $Y=1.13
+ $X2=0 $Y2=0
cc_750 N_A_1445_324#_c_875_n N_A_1295_379#_c_1148_n 7.70718e-19 $X=9.77 $Y=1.58
+ $X2=0 $Y2=0
cc_751 N_A_1445_324#_c_882_n N_A_1295_379#_M1001_g 0.00568271f $X=9.77 $Y=1.915
+ $X2=0 $Y2=0
cc_752 N_A_1445_324#_c_885_n N_A_1295_379#_M1001_g 0.0170541f $X=9.69 $Y=2.08
+ $X2=0 $Y2=0
cc_753 N_A_1445_324#_c_866_n N_A_1295_379#_c_1149_n 4.5415e-19 $X=7.375 $Y=1.695
+ $X2=0 $Y2=0
cc_754 N_A_1445_324#_c_877_n N_A_1295_379#_c_1161_n 0.0161515f $X=7.3 $Y=1.77
+ $X2=0 $Y2=0
cc_755 N_A_1445_324#_c_869_n N_A_1295_379#_c_1161_n 0.00515113f $X=7.94 $Y=1.57
+ $X2=0 $Y2=0
cc_756 N_A_1445_324#_c_940_p N_A_1295_379#_c_1161_n 0.00906837f $X=8.04 $Y=2.025
+ $X2=0 $Y2=0
cc_757 N_A_1445_324#_c_876_n N_A_1295_379#_c_1161_n 0.00418853f $X=7.615
+ $Y=1.587 $X2=0 $Y2=0
cc_758 N_A_1445_324#_c_877_n N_A_1295_379#_c_1150_n 0.00264287f $X=7.3 $Y=1.77
+ $X2=0 $Y2=0
cc_759 N_A_1445_324#_M1040_g N_A_1295_379#_c_1150_n 0.0051404f $X=7.69 $Y=0.73
+ $X2=0 $Y2=0
cc_760 N_A_1445_324#_c_869_n N_A_1295_379#_c_1150_n 0.0315837f $X=7.94 $Y=1.57
+ $X2=0 $Y2=0
cc_761 N_A_1445_324#_c_870_n N_A_1295_379#_c_1150_n 0.0111362f $X=7.94 $Y=1.57
+ $X2=0 $Y2=0
cc_762 N_A_1445_324#_c_876_n N_A_1295_379#_c_1150_n 0.0099726f $X=7.615 $Y=1.587
+ $X2=0 $Y2=0
cc_763 N_A_1445_324#_M1040_g N_A_1295_379#_c_1151_n 0.0114239f $X=7.69 $Y=0.73
+ $X2=0 $Y2=0
cc_764 N_A_1445_324#_c_869_n N_A_1295_379#_c_1151_n 0.0151939f $X=7.94 $Y=1.57
+ $X2=0 $Y2=0
cc_765 N_A_1445_324#_c_870_n N_A_1295_379#_c_1151_n 0.00671941f $X=7.94 $Y=1.57
+ $X2=0 $Y2=0
cc_766 N_A_1445_324#_M1040_g N_A_1295_379#_c_1152_n 0.00238028f $X=7.69 $Y=0.73
+ $X2=0 $Y2=0
cc_767 N_A_1445_324#_M1040_g N_A_1295_379#_c_1153_n 0.00291229f $X=7.69 $Y=0.73
+ $X2=0 $Y2=0
cc_768 N_A_1445_324#_c_869_n N_A_1295_379#_c_1153_n 0.0127902f $X=7.94 $Y=1.57
+ $X2=0 $Y2=0
cc_769 N_A_1445_324#_c_870_n N_A_1295_379#_c_1153_n 0.00212643f $X=7.94 $Y=1.57
+ $X2=0 $Y2=0
cc_770 N_A_1445_324#_c_912_p N_A_1295_379#_c_1154_n 0.0498275f $X=9.525 $Y=2.025
+ $X2=0 $Y2=0
cc_771 N_A_1445_324#_c_869_n N_A_1295_379#_c_1155_n 0.0132787f $X=7.94 $Y=1.57
+ $X2=0 $Y2=0
cc_772 N_A_1445_324#_c_870_n N_A_1295_379#_c_1155_n 0.00225681f $X=7.94 $Y=1.57
+ $X2=0 $Y2=0
cc_773 N_A_1445_324#_c_912_p N_A_1295_379#_c_1155_n 0.0135988f $X=9.525 $Y=2.025
+ $X2=0 $Y2=0
cc_774 N_A_1445_324#_c_877_n N_A_1295_379#_c_1165_n 0.00198585f $X=7.3 $Y=1.77
+ $X2=0 $Y2=0
cc_775 N_A_1445_324#_c_912_p N_A_1295_379#_c_1156_n 0.0223079f $X=9.525 $Y=2.025
+ $X2=0 $Y2=0
cc_776 N_A_1445_324#_c_871_n N_A_1295_379#_c_1156_n 0.00213344f $X=9.77 $Y=1.435
+ $X2=0 $Y2=0
cc_777 N_A_1445_324#_c_882_n N_A_1295_379#_c_1156_n 0.00199917f $X=9.77 $Y=1.915
+ $X2=0 $Y2=0
cc_778 N_A_1445_324#_c_874_n N_A_1295_379#_c_1156_n 0.0158213f $X=9.41 $Y=1.13
+ $X2=0 $Y2=0
cc_779 N_A_1445_324#_c_875_n N_A_1295_379#_c_1156_n 0.0234658f $X=9.77 $Y=1.58
+ $X2=0 $Y2=0
cc_780 N_A_1445_324#_c_866_n N_A_995_66#_c_1278_n 0.0226038f $X=7.375 $Y=1.695
+ $X2=0 $Y2=0
cc_781 N_A_1445_324#_c_877_n N_A_995_66#_M1034_g 0.0226038f $X=7.3 $Y=1.77 $X2=0
+ $Y2=0
cc_782 N_A_1445_324#_c_877_n N_A_995_66#_c_1289_n 0.00346109f $X=7.3 $Y=1.77
+ $X2=0 $Y2=0
cc_783 N_A_1445_324#_M1043_g N_A_995_66#_c_1289_n 0.0104164f $X=10.915 $Y=2.315
+ $X2=0 $Y2=0
cc_784 N_A_1445_324#_c_885_n N_A_995_66#_c_1289_n 0.00624358f $X=9.69 $Y=2.08
+ $X2=0 $Y2=0
cc_785 N_A_1445_324#_M1043_g N_A_995_66#_c_1293_n 0.024046f $X=10.915 $Y=2.315
+ $X2=0 $Y2=0
cc_786 N_A_1445_324#_M1027_g N_A_2299_119#_c_1584_n 0.00191906f $X=10.915
+ $Y=0.915 $X2=0 $Y2=0
cc_787 N_A_1445_324#_c_874_n N_A_1926_21#_M1008_g 0.00270963f $X=9.41 $Y=1.13
+ $X2=0 $Y2=0
cc_788 N_A_1445_324#_M1027_g N_A_1926_21#_c_1682_n 0.0103107f $X=10.915 $Y=0.915
+ $X2=0 $Y2=0
cc_789 N_A_1445_324#_M1027_g N_A_1926_21#_c_1684_n 0.00842571f $X=10.915
+ $Y=0.915 $X2=0 $Y2=0
cc_790 N_A_1445_324#_c_872_n N_A_1926_21#_c_1684_n 0.00810132f $X=10.775 $Y=1.56
+ $X2=0 $Y2=0
cc_791 N_A_1445_324#_c_874_n N_A_1926_21#_c_1684_n 0.00576447f $X=9.41 $Y=1.13
+ $X2=0 $Y2=0
cc_792 N_A_1445_324#_c_874_n N_A_1926_21#_c_1685_n 0.00848564f $X=9.41 $Y=1.13
+ $X2=0 $Y2=0
cc_793 N_A_1445_324#_M1043_g N_A_1926_21#_M1003_g 0.0162605f $X=10.915 $Y=2.315
+ $X2=0 $Y2=0
cc_794 N_A_1445_324#_c_871_n N_A_1926_21#_M1003_g 0.00414445f $X=9.77 $Y=1.435
+ $X2=0 $Y2=0
cc_795 N_A_1445_324#_c_882_n N_A_1926_21#_M1003_g 9.22822e-19 $X=9.77 $Y=1.915
+ $X2=0 $Y2=0
cc_796 N_A_1445_324#_c_872_n N_A_1926_21#_M1003_g 0.019681f $X=10.775 $Y=1.56
+ $X2=0 $Y2=0
cc_797 N_A_1445_324#_c_873_n N_A_1926_21#_M1003_g 0.018427f $X=10.775 $Y=1.56
+ $X2=0 $Y2=0
cc_798 N_A_1445_324#_c_874_n N_A_1926_21#_M1003_g 5.33645e-19 $X=9.41 $Y=1.13
+ $X2=0 $Y2=0
cc_799 N_A_1445_324#_c_885_n N_A_1926_21#_M1003_g 0.00237499f $X=9.69 $Y=2.08
+ $X2=0 $Y2=0
cc_800 N_A_1445_324#_c_869_n N_VPWR_M1009_d 0.00120223f $X=7.94 $Y=1.57 $X2=0
+ $Y2=0
cc_801 N_A_1445_324#_c_912_p N_VPWR_M1009_d 0.0271455f $X=9.525 $Y=2.025 $X2=0
+ $Y2=0
cc_802 N_A_1445_324#_c_940_p N_VPWR_M1009_d 0.0129227f $X=8.04 $Y=2.025 $X2=0
+ $Y2=0
cc_803 N_A_1445_324#_c_912_p N_VPWR_c_1945_n 0.0254908f $X=9.525 $Y=2.025 $X2=0
+ $Y2=0
cc_804 N_A_1445_324#_M1043_g N_VPWR_c_1946_n 0.0108626f $X=10.915 $Y=2.315 $X2=0
+ $Y2=0
cc_805 N_A_1445_324#_c_882_n N_VPWR_c_1946_n 2.87166e-19 $X=9.77 $Y=1.915 $X2=0
+ $Y2=0
cc_806 N_A_1445_324#_c_872_n N_VPWR_c_1946_n 0.0232879f $X=10.775 $Y=1.56 $X2=0
+ $Y2=0
cc_807 N_A_1445_324#_c_873_n N_VPWR_c_1946_n 0.00148357f $X=10.775 $Y=1.56 $X2=0
+ $Y2=0
cc_808 N_A_1445_324#_c_885_n N_VPWR_c_1946_n 0.0269238f $X=9.69 $Y=2.08 $X2=0
+ $Y2=0
cc_809 N_A_1445_324#_c_885_n N_VPWR_c_1955_n 0.00749462f $X=9.69 $Y=2.08 $X2=0
+ $Y2=0
cc_810 N_A_1445_324#_c_877_n N_VPWR_c_1940_n 9.4209e-19 $X=7.3 $Y=1.77 $X2=0
+ $Y2=0
cc_811 N_A_1445_324#_M1043_g N_VPWR_c_1940_n 9.39239e-19 $X=10.915 $Y=2.315
+ $X2=0 $Y2=0
cc_812 N_A_1445_324#_c_885_n N_VPWR_c_1940_n 0.00907254f $X=9.69 $Y=2.08 $X2=0
+ $Y2=0
cc_813 N_A_1445_324#_M1040_g N_VGND_c_2363_n 0.00534506f $X=7.69 $Y=0.73 $X2=0
+ $Y2=0
cc_814 N_A_1445_324#_M1027_g N_VGND_c_2364_n 0.0113526f $X=10.915 $Y=0.915 $X2=0
+ $Y2=0
cc_815 N_A_1445_324#_M1040_g N_VGND_c_2375_n 0.00370445f $X=7.69 $Y=0.73 $X2=0
+ $Y2=0
cc_816 N_A_1445_324#_M1040_g N_VGND_c_2379_n 0.00499434f $X=7.69 $Y=0.73 $X2=0
+ $Y2=0
cc_817 N_A_1445_324#_M1027_g N_VGND_c_2379_n 7.88961e-19 $X=10.915 $Y=0.915
+ $X2=0 $Y2=0
cc_818 N_A_1445_324#_c_872_n N_A_1752_60#_c_2537_n 0.00327398f $X=10.775 $Y=1.56
+ $X2=0 $Y2=0
cc_819 N_A_1445_324#_c_874_n N_A_1752_60#_c_2537_n 0.00529344f $X=9.41 $Y=1.13
+ $X2=0 $Y2=0
cc_820 N_A_1445_324#_M1000_d N_A_1752_60#_c_2544_n 0.00721354f $X=9.195 $Y=0.3
+ $X2=0 $Y2=0
cc_821 N_A_1445_324#_c_874_n N_A_1752_60#_c_2544_n 0.0295055f $X=9.41 $Y=1.13
+ $X2=0 $Y2=0
cc_822 N_SET_B_M1035_g N_A_1295_379#_M1000_g 0.0239466f $X=8.685 $Y=0.62 $X2=0
+ $Y2=0
cc_823 N_SET_B_c_1008_n N_A_1295_379#_M1000_g 0.00663051f $X=13.055 $Y=1.295
+ $X2=0 $Y2=0
cc_824 N_SET_B_c_1009_n N_A_1295_379#_M1000_g 0.00147849f $X=9.025 $Y=1.295
+ $X2=0 $Y2=0
cc_825 N_SET_B_c_1010_n N_A_1295_379#_M1000_g 0.00515477f $X=8.88 $Y=1.295 $X2=0
+ $Y2=0
cc_826 N_SET_B_c_1013_n N_A_1295_379#_M1000_g 0.0149533f $X=8.67 $Y=1.245 $X2=0
+ $Y2=0
cc_827 N_SET_B_c_1008_n N_A_1295_379#_c_1147_n 0.00329006f $X=13.055 $Y=1.295
+ $X2=0 $Y2=0
cc_828 N_SET_B_M1030_g N_A_1295_379#_c_1148_n 0.0212f $X=8.76 $Y=2.315 $X2=0
+ $Y2=0
cc_829 N_SET_B_M1035_g N_A_1295_379#_c_1151_n 9.57837e-19 $X=8.685 $Y=0.62 $X2=0
+ $Y2=0
cc_830 N_SET_B_c_1009_n N_A_1295_379#_c_1151_n 2.60497e-19 $X=9.025 $Y=1.295
+ $X2=0 $Y2=0
cc_831 N_SET_B_c_1010_n N_A_1295_379#_c_1151_n 0.0116223f $X=8.88 $Y=1.295 $X2=0
+ $Y2=0
cc_832 N_SET_B_c_1013_n N_A_1295_379#_c_1151_n 0.00365672f $X=8.67 $Y=1.245
+ $X2=0 $Y2=0
cc_833 N_SET_B_M1030_g N_A_1295_379#_c_1153_n 0.00359952f $X=8.76 $Y=2.315 $X2=0
+ $Y2=0
cc_834 N_SET_B_c_1009_n N_A_1295_379#_c_1153_n 9.1209e-19 $X=9.025 $Y=1.295
+ $X2=0 $Y2=0
cc_835 N_SET_B_c_1010_n N_A_1295_379#_c_1153_n 0.0126462f $X=8.88 $Y=1.295 $X2=0
+ $Y2=0
cc_836 N_SET_B_c_1013_n N_A_1295_379#_c_1153_n 0.004384f $X=8.67 $Y=1.245 $X2=0
+ $Y2=0
cc_837 N_SET_B_M1030_g N_A_1295_379#_c_1154_n 0.0120251f $X=8.76 $Y=2.315 $X2=0
+ $Y2=0
cc_838 N_SET_B_c_1008_n N_A_1295_379#_c_1154_n 0.00593081f $X=13.055 $Y=1.295
+ $X2=0 $Y2=0
cc_839 N_SET_B_c_1009_n N_A_1295_379#_c_1154_n 0.00809369f $X=9.025 $Y=1.295
+ $X2=0 $Y2=0
cc_840 N_SET_B_c_1010_n N_A_1295_379#_c_1154_n 0.0273813f $X=8.88 $Y=1.295 $X2=0
+ $Y2=0
cc_841 N_SET_B_c_1013_n N_A_1295_379#_c_1154_n 0.00526971f $X=8.67 $Y=1.245
+ $X2=0 $Y2=0
cc_842 N_SET_B_M1030_g N_A_1295_379#_c_1156_n 2.10119e-19 $X=8.76 $Y=2.315 $X2=0
+ $Y2=0
cc_843 N_SET_B_c_1008_n N_A_1295_379#_c_1156_n 0.0101711f $X=13.055 $Y=1.295
+ $X2=0 $Y2=0
cc_844 N_SET_B_c_1009_n N_A_1295_379#_c_1156_n 2.46208e-19 $X=9.025 $Y=1.295
+ $X2=0 $Y2=0
cc_845 N_SET_B_c_1013_n N_A_1295_379#_c_1156_n 7.24757e-19 $X=8.67 $Y=1.245
+ $X2=0 $Y2=0
cc_846 N_SET_B_M1030_g N_A_995_66#_c_1289_n 0.0104164f $X=8.76 $Y=2.315 $X2=0
+ $Y2=0
cc_847 N_SET_B_c_1008_n N_A_995_66#_c_1292_n 0.00306946f $X=13.055 $Y=1.295
+ $X2=0 $Y2=0
cc_848 N_SET_B_c_1008_n N_A_995_66#_c_1280_n 0.0016469f $X=13.055 $Y=1.295 $X2=0
+ $Y2=0
cc_849 N_SET_B_c_1008_n N_A_995_66#_c_1282_n 0.0049252f $X=13.055 $Y=1.295 $X2=0
+ $Y2=0
cc_850 N_SET_B_c_1008_n N_A_2449_137#_c_1397_n 0.00327119f $X=13.055 $Y=1.295
+ $X2=0 $Y2=0
cc_851 N_SET_B_c_1012_n N_A_2449_137#_c_1397_n 8.45641e-19 $X=13.2 $Y=1.295
+ $X2=0 $Y2=0
cc_852 N_SET_B_c_1015_n N_A_2449_137#_c_1397_n 0.0116588f $X=13.165 $Y=1.345
+ $X2=0 $Y2=0
cc_853 N_SET_B_c_1008_n N_A_2449_137#_c_1398_n 0.0149603f $X=13.055 $Y=1.295
+ $X2=0 $Y2=0
cc_854 N_SET_B_c_1012_n N_A_2449_137#_c_1398_n 0.00293444f $X=13.2 $Y=1.295
+ $X2=0 $Y2=0
cc_855 N_SET_B_c_1014_n N_A_2449_137#_c_1398_n 0.0218574f $X=13.165 $Y=1.51
+ $X2=0 $Y2=0
cc_856 N_SET_B_c_1015_n N_A_2449_137#_c_1398_n 0.00201317f $X=13.165 $Y=1.345
+ $X2=0 $Y2=0
cc_857 N_SET_B_c_1008_n N_A_2449_137#_c_1399_n 0.00209625f $X=13.055 $Y=1.295
+ $X2=0 $Y2=0
cc_858 N_SET_B_M1011_g N_A_2449_137#_M1037_g 0.00956465f $X=13.485 $Y=2.675
+ $X2=0 $Y2=0
cc_859 N_SET_B_c_1017_n N_A_2449_137#_c_1416_n 0.00267797f $X=13.255 $Y=1.975
+ $X2=0 $Y2=0
cc_860 N_SET_B_M1011_g N_A_2449_137#_c_1416_n 0.0123545f $X=13.485 $Y=2.675
+ $X2=0 $Y2=0
cc_861 N_SET_B_c_1019_n N_A_2449_137#_c_1416_n 0.0155305f $X=13.485 $Y=2.05
+ $X2=0 $Y2=0
cc_862 N_SET_B_c_1008_n N_A_2449_137#_c_1416_n 0.0102483f $X=13.055 $Y=1.295
+ $X2=0 $Y2=0
cc_863 N_SET_B_c_1011_n N_A_2449_137#_c_1416_n 0.00153029f $X=13.2 $Y=1.295
+ $X2=0 $Y2=0
cc_864 N_SET_B_c_1012_n N_A_2449_137#_c_1416_n 0.0254703f $X=13.2 $Y=1.295 $X2=0
+ $Y2=0
cc_865 N_SET_B_c_1014_n N_A_2449_137#_c_1416_n 0.0010031f $X=13.165 $Y=1.51
+ $X2=0 $Y2=0
cc_866 N_SET_B_c_1017_n N_A_2449_137#_c_1417_n 0.0106827f $X=13.255 $Y=1.975
+ $X2=0 $Y2=0
cc_867 N_SET_B_M1011_g N_A_2449_137#_c_1417_n 0.0039509f $X=13.485 $Y=2.675
+ $X2=0 $Y2=0
cc_868 N_SET_B_c_1008_n N_A_2449_137#_c_1417_n 0.0034753f $X=13.055 $Y=1.295
+ $X2=0 $Y2=0
cc_869 N_SET_B_M1011_g N_A_2449_137#_c_1453_n 0.00771458f $X=13.485 $Y=2.675
+ $X2=0 $Y2=0
cc_870 N_SET_B_M1011_g N_A_2449_137#_c_1454_n 0.0079779f $X=13.485 $Y=2.675
+ $X2=0 $Y2=0
cc_871 N_SET_B_c_1017_n N_A_2449_137#_c_1411_n 0.00944115f $X=13.255 $Y=1.975
+ $X2=0 $Y2=0
cc_872 N_SET_B_c_1012_n N_A_2449_137#_c_1411_n 0.00146194f $X=13.2 $Y=1.295
+ $X2=0 $Y2=0
cc_873 N_SET_B_c_1008_n N_A_2299_119#_M1016_d 0.00155613f $X=13.055 $Y=1.295
+ $X2=-0.19 $Y2=-0.245
cc_874 N_SET_B_c_1012_n N_A_2299_119#_M1036_g 5.69934e-19 $X=13.2 $Y=1.295 $X2=0
+ $Y2=0
cc_875 N_SET_B_c_1014_n N_A_2299_119#_M1036_g 0.00402075f $X=13.165 $Y=1.51
+ $X2=0 $Y2=0
cc_876 N_SET_B_c_1015_n N_A_2299_119#_M1036_g 0.0213423f $X=13.165 $Y=1.345
+ $X2=0 $Y2=0
cc_877 N_SET_B_c_1017_n N_A_2299_119#_M1045_g 0.00591636f $X=13.255 $Y=1.975
+ $X2=0 $Y2=0
cc_878 N_SET_B_c_1019_n N_A_2299_119#_M1045_g 0.0241099f $X=13.485 $Y=2.05 $X2=0
+ $Y2=0
cc_879 N_SET_B_c_1008_n N_A_2299_119#_c_1615_n 0.0464772f $X=13.055 $Y=1.295
+ $X2=0 $Y2=0
cc_880 N_SET_B_c_1011_n N_A_2299_119#_c_1615_n 0.00277178f $X=13.2 $Y=1.295
+ $X2=0 $Y2=0
cc_881 N_SET_B_c_1012_n N_A_2299_119#_c_1615_n 0.0153976f $X=13.2 $Y=1.295 $X2=0
+ $Y2=0
cc_882 N_SET_B_c_1014_n N_A_2299_119#_c_1615_n 6.00022e-19 $X=13.165 $Y=1.51
+ $X2=0 $Y2=0
cc_883 N_SET_B_c_1015_n N_A_2299_119#_c_1615_n 0.011959f $X=13.165 $Y=1.345
+ $X2=0 $Y2=0
cc_884 N_SET_B_c_1008_n N_A_2299_119#_c_1584_n 0.012104f $X=13.055 $Y=1.295
+ $X2=0 $Y2=0
cc_885 N_SET_B_c_1008_n N_A_2299_119#_c_1585_n 0.026166f $X=13.055 $Y=1.295
+ $X2=0 $Y2=0
cc_886 N_SET_B_c_1014_n N_A_2299_119#_c_1586_n 0.0011048f $X=13.165 $Y=1.51
+ $X2=0 $Y2=0
cc_887 N_SET_B_c_1019_n N_A_2299_119#_c_1587_n 0.00130767f $X=13.485 $Y=2.05
+ $X2=0 $Y2=0
cc_888 N_SET_B_c_1012_n N_A_2299_119#_c_1587_n 0.00118003f $X=13.2 $Y=1.295
+ $X2=0 $Y2=0
cc_889 N_SET_B_c_1014_n N_A_2299_119#_c_1587_n 0.0199946f $X=13.165 $Y=1.51
+ $X2=0 $Y2=0
cc_890 N_SET_B_c_1011_n N_A_2299_119#_c_1588_n 0.00717504f $X=13.2 $Y=1.295
+ $X2=0 $Y2=0
cc_891 N_SET_B_c_1012_n N_A_2299_119#_c_1588_n 0.0344418f $X=13.2 $Y=1.295 $X2=0
+ $Y2=0
cc_892 N_SET_B_c_1014_n N_A_2299_119#_c_1588_n 4.91579e-19 $X=13.165 $Y=1.51
+ $X2=0 $Y2=0
cc_893 N_SET_B_c_1015_n N_A_2299_119#_c_1588_n 0.00359807f $X=13.165 $Y=1.345
+ $X2=0 $Y2=0
cc_894 N_SET_B_c_1015_n N_A_1926_21#_c_1682_n 0.0100396f $X=13.165 $Y=1.345
+ $X2=0 $Y2=0
cc_895 N_SET_B_c_1008_n N_A_1926_21#_c_1684_n 0.00737091f $X=13.055 $Y=1.295
+ $X2=0 $Y2=0
cc_896 N_SET_B_c_1008_n N_A_1926_21#_M1003_g 0.0062067f $X=13.055 $Y=1.295 $X2=0
+ $Y2=0
cc_897 N_SET_B_M1030_g N_VPWR_c_1945_n 0.013968f $X=8.76 $Y=2.315 $X2=0 $Y2=0
cc_898 N_SET_B_M1011_g N_VPWR_c_1947_n 0.00647602f $X=13.485 $Y=2.675 $X2=0
+ $Y2=0
cc_899 N_SET_B_c_1019_n N_VPWR_c_1947_n 9.25689e-19 $X=13.485 $Y=2.05 $X2=0
+ $Y2=0
cc_900 N_SET_B_M1011_g N_VPWR_c_1957_n 0.00549284f $X=13.485 $Y=2.675 $X2=0
+ $Y2=0
cc_901 N_SET_B_M1030_g N_VPWR_c_1940_n 9.39239e-19 $X=8.76 $Y=2.315 $X2=0 $Y2=0
cc_902 N_SET_B_M1011_g N_VPWR_c_1940_n 0.0113256f $X=13.485 $Y=2.675 $X2=0 $Y2=0
cc_903 N_SET_B_c_1008_n N_VGND_M1025_d 0.00507456f $X=13.055 $Y=1.295 $X2=0
+ $Y2=0
cc_904 N_SET_B_M1035_g N_VGND_c_2363_n 0.0029201f $X=8.685 $Y=0.62 $X2=0 $Y2=0
cc_905 N_SET_B_c_1008_n N_VGND_c_2364_n 0.00153488f $X=13.055 $Y=1.295 $X2=0
+ $Y2=0
cc_906 N_SET_B_c_1015_n N_VGND_c_2366_n 0.00415562f $X=13.165 $Y=1.345 $X2=0
+ $Y2=0
cc_907 N_SET_B_M1035_g N_VGND_c_2376_n 0.00318662f $X=8.685 $Y=0.62 $X2=0 $Y2=0
cc_908 N_SET_B_M1035_g N_VGND_c_2379_n 0.00547455f $X=8.685 $Y=0.62 $X2=0 $Y2=0
cc_909 N_SET_B_c_1015_n N_VGND_c_2379_n 9.39239e-19 $X=13.165 $Y=1.345 $X2=0
+ $Y2=0
cc_910 N_SET_B_M1035_g N_A_1752_60#_c_2540_n 0.00455439f $X=8.685 $Y=0.62 $X2=0
+ $Y2=0
cc_911 N_SET_B_c_1008_n N_A_1752_60#_c_2540_n 0.00143785f $X=13.055 $Y=1.295
+ $X2=0 $Y2=0
cc_912 N_SET_B_c_1009_n N_A_1752_60#_c_2540_n 0.00293608f $X=9.025 $Y=1.295
+ $X2=0 $Y2=0
cc_913 N_SET_B_c_1010_n N_A_1752_60#_c_2540_n 0.0160798f $X=8.88 $Y=1.295 $X2=0
+ $Y2=0
cc_914 N_SET_B_c_1013_n N_A_1752_60#_c_2540_n 0.00183899f $X=8.67 $Y=1.245 $X2=0
+ $Y2=0
cc_915 N_SET_B_c_1008_n N_A_1752_60#_c_2537_n 0.00633611f $X=13.055 $Y=1.295
+ $X2=0 $Y2=0
cc_916 N_SET_B_c_1008_n N_A_1752_60#_c_2544_n 0.00691092f $X=13.055 $Y=1.295
+ $X2=0 $Y2=0
cc_917 N_SET_B_c_1008_n A_2198_119# 0.00205389f $X=13.055 $Y=1.295 $X2=-0.19
+ $Y2=-0.245
cc_918 N_SET_B_c_1008_n A_2401_163# 0.00201638f $X=13.055 $Y=1.295 $X2=-0.19
+ $Y2=-0.245
cc_919 N_SET_B_c_1011_n N_A_2636_119#_M1022_d 0.00138713f $X=13.2 $Y=1.295
+ $X2=-0.19 $Y2=-0.245
cc_920 N_SET_B_c_1012_n N_A_2636_119#_M1022_d 7.81362e-19 $X=13.2 $Y=1.295
+ $X2=-0.19 $Y2=-0.245
cc_921 N_SET_B_c_1015_n N_A_2636_119#_c_2569_n 0.00175602f $X=13.165 $Y=1.345
+ $X2=0 $Y2=0
cc_922 N_A_1295_379#_c_1149_n N_A_995_66#_M1005_g 0.00988007f $X=6.7 $Y=0.78
+ $X2=0 $Y2=0
cc_923 N_A_1295_379#_c_1149_n N_A_995_66#_c_1277_n 0.0114143f $X=6.7 $Y=0.78
+ $X2=0 $Y2=0
cc_924 N_A_1295_379#_c_1149_n N_A_995_66#_c_1278_n 0.0243902f $X=6.7 $Y=0.78
+ $X2=0 $Y2=0
cc_925 N_A_1295_379#_c_1150_n N_A_995_66#_c_1278_n 0.00152607f $X=7.575 $Y=1.875
+ $X2=0 $Y2=0
cc_926 N_A_1295_379#_c_1149_n N_A_995_66#_M1034_g 0.0032166f $X=6.7 $Y=0.78
+ $X2=0 $Y2=0
cc_927 N_A_1295_379#_c_1161_n N_A_995_66#_M1034_g 0.0141724f $X=7.49 $Y=1.96
+ $X2=0 $Y2=0
cc_928 N_A_1295_379#_c_1165_n N_A_995_66#_M1034_g 0.00858385f $X=6.697 $Y=1.96
+ $X2=0 $Y2=0
cc_929 N_A_1295_379#_M1001_g N_A_995_66#_c_1289_n 0.0103003f $X=9.905 $Y=2.315
+ $X2=0 $Y2=0
cc_930 N_A_1295_379#_M1000_g N_A_1926_21#_c_1683_n 0.0274866f $X=9.12 $Y=0.62
+ $X2=0 $Y2=0
cc_931 N_A_1295_379#_c_1147_n N_A_1926_21#_c_1685_n 0.0096417f $X=9.83 $Y=1.66
+ $X2=0 $Y2=0
cc_932 N_A_1295_379#_c_1147_n N_A_1926_21#_M1003_g 0.0644444f $X=9.83 $Y=1.66
+ $X2=0 $Y2=0
cc_933 N_A_1295_379#_c_1148_n N_A_1926_21#_M1003_g 0.00166896f $X=9.505 $Y=1.66
+ $X2=0 $Y2=0
cc_934 N_A_1295_379#_c_1161_n N_VPWR_M1009_d 0.0120976f $X=7.49 $Y=1.96 $X2=0
+ $Y2=0
cc_935 N_A_1295_379#_M1001_g N_VPWR_c_1946_n 0.00295094f $X=9.905 $Y=2.315 $X2=0
+ $Y2=0
cc_936 N_A_1295_379#_M1001_g N_VPWR_c_1940_n 9.39239e-19 $X=9.905 $Y=2.315 $X2=0
+ $Y2=0
cc_937 N_A_1295_379#_c_1165_n N_A_200_119#_c_2147_n 8.04338e-19 $X=6.697 $Y=1.96
+ $X2=0 $Y2=0
cc_938 N_A_1295_379#_c_1165_n N_A_200_119#_c_2149_n 0.0171783f $X=6.697 $Y=1.96
+ $X2=0 $Y2=0
cc_939 N_A_1295_379#_c_1149_n N_A_200_119#_c_2130_n 0.0584174f $X=6.7 $Y=0.78
+ $X2=0 $Y2=0
cc_940 N_A_1295_379#_c_1149_n N_A_200_119#_c_2131_n 0.0180055f $X=6.7 $Y=0.78
+ $X2=0 $Y2=0
cc_941 N_A_1295_379#_c_1161_n A_1397_379# 0.0048076f $X=7.49 $Y=1.96 $X2=-0.19
+ $Y2=-0.245
cc_942 N_A_1295_379#_c_1149_n N_VGND_c_2375_n 0.00905745f $X=6.7 $Y=0.78 $X2=0
+ $Y2=0
cc_943 N_A_1295_379#_M1000_g N_VGND_c_2376_n 0.00318662f $X=9.12 $Y=0.62 $X2=0
+ $Y2=0
cc_944 N_A_1295_379#_M1000_g N_VGND_c_2379_n 0.00492863f $X=9.12 $Y=0.62 $X2=0
+ $Y2=0
cc_945 N_A_1295_379#_c_1149_n N_VGND_c_2379_n 0.00966388f $X=6.7 $Y=0.78 $X2=0
+ $Y2=0
cc_946 N_A_1295_379#_M1000_g N_A_1752_60#_c_2540_n 0.00324578f $X=9.12 $Y=0.62
+ $X2=0 $Y2=0
cc_947 N_A_1295_379#_M1000_g N_A_1752_60#_c_2537_n 4.03553e-19 $X=9.12 $Y=0.62
+ $X2=0 $Y2=0
cc_948 N_A_1295_379#_M1000_g N_A_1752_60#_c_2544_n 0.00935256f $X=9.12 $Y=0.62
+ $X2=0 $Y2=0
cc_949 N_A_1295_379#_c_1148_n N_A_1752_60#_c_2544_n 3.5249e-19 $X=9.505 $Y=1.66
+ $X2=0 $Y2=0
cc_950 N_A_1295_379#_c_1156_n N_A_1752_60#_c_2544_n 4.22825e-19 $X=9.34 $Y=1.57
+ $X2=0 $Y2=0
cc_951 N_A_995_66#_c_1280_n N_A_2449_137#_c_1397_n 0.0216242f $X=11.93 $Y=1.31
+ $X2=0 $Y2=0
cc_952 N_A_995_66#_c_1282_n N_A_2449_137#_c_1399_n 0.0216242f $X=11.93 $Y=1.385
+ $X2=0 $Y2=0
cc_953 N_A_995_66#_c_1280_n N_A_2299_119#_c_1615_n 0.00730876f $X=11.93 $Y=1.31
+ $X2=0 $Y2=0
cc_954 N_A_995_66#_c_1280_n N_A_2299_119#_c_1584_n 0.0136083f $X=11.93 $Y=1.31
+ $X2=0 $Y2=0
cc_955 N_A_995_66#_M1038_g N_A_2299_119#_c_1590_n 0.0101675f $X=11.42 $Y=2.56
+ $X2=0 $Y2=0
cc_956 N_A_995_66#_c_1292_n N_A_2299_119#_c_1590_n 0.00913f $X=11.74 $Y=1.99
+ $X2=0 $Y2=0
cc_957 N_A_995_66#_c_1292_n N_A_2299_119#_c_1585_n 0.010404f $X=11.74 $Y=1.99
+ $X2=0 $Y2=0
cc_958 N_A_995_66#_c_1279_n N_A_2299_119#_c_1585_n 0.0197994f $X=11.815 $Y=1.915
+ $X2=0 $Y2=0
cc_959 N_A_995_66#_c_1280_n N_A_2299_119#_c_1585_n 0.00445645f $X=11.93 $Y=1.31
+ $X2=0 $Y2=0
cc_960 N_A_995_66#_c_1282_n N_A_2299_119#_c_1585_n 0.00762831f $X=11.93 $Y=1.385
+ $X2=0 $Y2=0
cc_961 N_A_995_66#_c_1280_n N_A_1926_21#_c_1682_n 0.00410485f $X=11.93 $Y=1.31
+ $X2=0 $Y2=0
cc_962 N_A_995_66#_c_1289_n N_A_1926_21#_M1003_g 0.0103107f $X=11.345 $Y=3.15
+ $X2=0 $Y2=0
cc_963 N_A_995_66#_c_1289_n N_VPWR_c_1945_n 0.0261591f $X=11.345 $Y=3.15 $X2=0
+ $Y2=0
cc_964 N_A_995_66#_c_1289_n N_VPWR_c_1946_n 0.025796f $X=11.345 $Y=3.15 $X2=0
+ $Y2=0
cc_965 N_A_995_66#_M1038_g N_VPWR_c_1946_n 0.0010345f $X=11.42 $Y=2.56 $X2=0
+ $Y2=0
cc_966 N_A_995_66#_c_1289_n N_VPWR_c_1955_n 0.0567941f $X=11.345 $Y=3.15 $X2=0
+ $Y2=0
cc_967 N_A_995_66#_c_1290_n N_VPWR_c_1961_n 0.0525681f $X=6.985 $Y=3.15 $X2=0
+ $Y2=0
cc_968 N_A_995_66#_c_1289_n N_VPWR_c_1962_n 0.0241625f $X=11.345 $Y=3.15 $X2=0
+ $Y2=0
cc_969 N_A_995_66#_c_1289_n N_VPWR_c_1940_n 0.176313f $X=11.345 $Y=3.15 $X2=0
+ $Y2=0
cc_970 N_A_995_66#_c_1290_n N_VPWR_c_1940_n 0.0104981f $X=6.985 $Y=3.15 $X2=0
+ $Y2=0
cc_971 N_A_995_66#_M1034_g N_A_200_119#_c_2147_n 7.53526e-19 $X=6.91 $Y=2.105
+ $X2=0 $Y2=0
cc_972 N_A_995_66#_c_1284_n N_A_200_119#_c_2147_n 0.0183115f $X=5.835 $Y=1.51
+ $X2=0 $Y2=0
cc_973 N_A_995_66#_c_1286_n N_A_200_119#_c_2147_n 0.0050931f $X=5.835 $Y=1.42
+ $X2=0 $Y2=0
cc_974 N_A_995_66#_M1018_s N_A_200_119#_c_2148_n 0.00322301f $X=4.99 $Y=1.835
+ $X2=0 $Y2=0
cc_975 N_A_995_66#_c_1295_n N_A_200_119#_c_2148_n 0.00960786f $X=5.13 $Y=1.98
+ $X2=0 $Y2=0
cc_976 N_A_995_66#_c_1275_n N_A_200_119#_c_2149_n 0.00512762f $X=6.33 $Y=1.42
+ $X2=0 $Y2=0
cc_977 N_A_995_66#_c_1275_n N_A_200_119#_c_2130_n 0.0112192f $X=6.33 $Y=1.42
+ $X2=0 $Y2=0
cc_978 N_A_995_66#_M1005_g N_A_200_119#_c_2130_n 0.00809257f $X=6.405 $Y=0.835
+ $X2=0 $Y2=0
cc_979 N_A_995_66#_c_1278_n N_A_200_119#_c_2130_n 9.66655e-19 $X=6.91 $Y=1.77
+ $X2=0 $Y2=0
cc_980 N_A_995_66#_M1034_g N_A_200_119#_c_2130_n 2.12666e-19 $X=6.91 $Y=2.105
+ $X2=0 $Y2=0
cc_981 N_A_995_66#_c_1281_n N_A_200_119#_c_2130_n 0.00262173f $X=6.405 $Y=1.42
+ $X2=0 $Y2=0
cc_982 N_A_995_66#_c_1284_n N_A_200_119#_c_2130_n 0.0245349f $X=5.835 $Y=1.51
+ $X2=0 $Y2=0
cc_983 N_A_995_66#_c_1286_n N_A_200_119#_c_2130_n 7.52082e-19 $X=5.835 $Y=1.42
+ $X2=0 $Y2=0
cc_984 N_A_995_66#_c_1275_n N_A_200_119#_c_2131_n 0.00530563f $X=6.33 $Y=1.42
+ $X2=0 $Y2=0
cc_985 N_A_995_66#_M1005_g N_A_200_119#_c_2131_n 0.00667446f $X=6.405 $Y=0.835
+ $X2=0 $Y2=0
cc_986 N_A_995_66#_M1005_g N_VGND_c_2362_n 0.00314964f $X=6.405 $Y=0.835 $X2=0
+ $Y2=0
cc_987 N_A_995_66#_c_1283_n N_VGND_c_2362_n 0.018006f $X=5.12 $Y=0.54 $X2=0
+ $Y2=0
cc_988 N_A_995_66#_c_1284_n N_VGND_c_2362_n 0.0119025f $X=5.835 $Y=1.51 $X2=0
+ $Y2=0
cc_989 N_A_995_66#_c_1286_n N_VGND_c_2362_n 0.00219291f $X=5.835 $Y=1.42 $X2=0
+ $Y2=0
cc_990 N_A_995_66#_c_1283_n N_VGND_c_2374_n 0.0173762f $X=5.12 $Y=0.54 $X2=0
+ $Y2=0
cc_991 N_A_995_66#_M1005_g N_VGND_c_2379_n 9.49986e-19 $X=6.405 $Y=0.835 $X2=0
+ $Y2=0
cc_992 N_A_995_66#_c_1280_n N_VGND_c_2379_n 8.16873e-19 $X=11.93 $Y=1.31 $X2=0
+ $Y2=0
cc_993 N_A_995_66#_c_1283_n N_VGND_c_2379_n 0.0123312f $X=5.12 $Y=0.54 $X2=0
+ $Y2=0
cc_994 N_A_2449_137#_c_1407_n N_A_2299_119#_M1036_g 0.00841591f $X=13.99
+ $Y=0.935 $X2=0 $Y2=0
cc_995 N_A_2449_137#_c_1408_n N_A_2299_119#_M1036_g 0.00238093f $X=14.135
+ $Y=2.47 $X2=0 $Y2=0
cc_996 N_A_2449_137#_c_1416_n N_A_2299_119#_M1045_g 0.00735586f $X=13.535
+ $Y=2.125 $X2=0 $Y2=0
cc_997 N_A_2449_137#_c_1453_n N_A_2299_119#_M1045_g 0.00183554f $X=13.7 $Y=2.4
+ $X2=0 $Y2=0
cc_998 N_A_2449_137#_c_1463_p N_A_2299_119#_M1045_g 0.0119774f $X=14.05 $Y=2.555
+ $X2=0 $Y2=0
cc_999 N_A_2449_137#_c_1454_n N_A_2299_119#_M1045_g 0.00886867f $X=13.7 $Y=2.555
+ $X2=0 $Y2=0
cc_1000 N_A_2449_137#_c_1397_n N_A_2299_119#_c_1615_n 0.0111405f $X=12.32
+ $Y=1.31 $X2=0 $Y2=0
cc_1001 N_A_2449_137#_c_1398_n N_A_2299_119#_c_1615_n 0.00951474f $X=12.64
+ $Y=1.385 $X2=0 $Y2=0
cc_1002 N_A_2449_137#_c_1407_n N_A_2299_119#_c_1615_n 0.0123421f $X=13.99
+ $Y=0.935 $X2=0 $Y2=0
cc_1003 N_A_2449_137#_c_1397_n N_A_2299_119#_c_1584_n 0.00217131f $X=12.32
+ $Y=1.31 $X2=0 $Y2=0
cc_1004 N_A_2449_137#_c_1399_n N_A_2299_119#_c_1585_n 0.00137569f $X=12.395
+ $Y=1.385 $X2=0 $Y2=0
cc_1005 N_A_2449_137#_c_1416_n N_A_2299_119#_c_1586_n 0.0253057f $X=13.535
+ $Y=2.125 $X2=0 $Y2=0
cc_1006 N_A_2449_137#_c_1408_n N_A_2299_119#_c_1586_n 0.0237544f $X=14.135
+ $Y=2.47 $X2=0 $Y2=0
cc_1007 N_A_2449_137#_c_1416_n N_A_2299_119#_c_1587_n 0.00223972f $X=13.535
+ $Y=2.125 $X2=0 $Y2=0
cc_1008 N_A_2449_137#_c_1408_n N_A_2299_119#_c_1587_n 0.0114928f $X=14.135
+ $Y=2.47 $X2=0 $Y2=0
cc_1009 N_A_2449_137#_c_1409_n N_A_2299_119#_c_1587_n 0.00327718f $X=14.062
+ $Y=1.255 $X2=0 $Y2=0
cc_1010 N_A_2449_137#_c_1407_n N_A_2299_119#_c_1588_n 0.0165547f $X=13.99
+ $Y=0.935 $X2=0 $Y2=0
cc_1011 N_A_2449_137#_c_1408_n N_A_2299_119#_c_1588_n 0.00764731f $X=14.135
+ $Y=2.47 $X2=0 $Y2=0
cc_1012 N_A_2449_137#_c_1419_n N_A_1926_21#_M1019_s 0.00245596f $X=15.55
+ $Y=2.555 $X2=0 $Y2=0
cc_1013 N_A_2449_137#_c_1397_n N_A_1926_21#_c_1682_n 0.0042225f $X=12.32 $Y=1.31
+ $X2=0 $Y2=0
cc_1014 N_A_2449_137#_c_1416_n N_A_1926_21#_M1044_g 2.6083e-19 $X=13.535
+ $Y=2.125 $X2=0 $Y2=0
cc_1015 N_A_2449_137#_c_1408_n N_A_1926_21#_M1044_g 0.016608f $X=14.135 $Y=2.47
+ $X2=0 $Y2=0
cc_1016 N_A_2449_137#_c_1419_n N_A_1926_21#_M1044_g 0.0146662f $X=15.55 $Y=2.555
+ $X2=0 $Y2=0
cc_1017 N_A_2449_137#_c_1454_n N_A_1926_21#_M1044_g 0.00156652f $X=13.7 $Y=2.555
+ $X2=0 $Y2=0
cc_1018 N_A_2449_137#_c_1483_p N_A_1926_21#_M1044_g 0.00230613f $X=14.135
+ $Y=2.555 $X2=0 $Y2=0
cc_1019 N_A_2449_137#_c_1407_n N_A_1926_21#_M1017_g 0.00336698f $X=13.99
+ $Y=0.935 $X2=0 $Y2=0
cc_1020 N_A_2449_137#_c_1409_n N_A_1926_21#_M1017_g 5.91445e-19 $X=14.062
+ $Y=1.255 $X2=0 $Y2=0
cc_1021 N_A_2449_137#_c_1408_n N_A_1926_21#_c_1688_n 0.00358982f $X=14.135
+ $Y=2.47 $X2=0 $Y2=0
cc_1022 N_A_2449_137#_c_1409_n N_A_1926_21#_c_1689_n 0.00447937f $X=14.062
+ $Y=1.255 $X2=0 $Y2=0
cc_1023 N_A_2449_137#_c_1409_n N_A_1926_21#_c_1697_n 0.0564867f $X=14.062
+ $Y=1.255 $X2=0 $Y2=0
cc_1024 N_A_2449_137#_c_1408_n N_A_1926_21#_c_1690_n 0.0018108f $X=14.135
+ $Y=2.47 $X2=0 $Y2=0
cc_1025 N_A_2449_137#_c_1407_n N_A_1926_21#_c_1692_n 0.00600185f $X=13.99
+ $Y=0.935 $X2=0 $Y2=0
cc_1026 N_A_2449_137#_c_1409_n N_A_1926_21#_c_1692_n 0.00611007f $X=14.062
+ $Y=1.255 $X2=0 $Y2=0
cc_1027 N_A_2449_137#_c_1408_n N_A_1926_21#_c_1698_n 0.023891f $X=14.135 $Y=2.47
+ $X2=0 $Y2=0
cc_1028 N_A_2449_137#_c_1419_n N_A_1926_21#_c_1698_n 0.0254784f $X=15.55
+ $Y=2.555 $X2=0 $Y2=0
cc_1029 N_A_2449_137#_M1020_g N_A_1926_21#_c_1699_n 2.92644e-19 $X=15.77
+ $Y=2.465 $X2=0 $Y2=0
cc_1030 N_A_2449_137#_c_1419_n N_A_1926_21#_c_1699_n 0.0312897f $X=15.55
+ $Y=2.555 $X2=0 $Y2=0
cc_1031 N_A_2449_137#_c_1420_n N_A_1926_21#_c_1699_n 0.0150776f $X=15.635
+ $Y=2.47 $X2=0 $Y2=0
cc_1032 N_A_2449_137#_M1020_g N_RESET_B_M1019_g 0.0277037f $X=15.77 $Y=2.465
+ $X2=0 $Y2=0
cc_1033 N_A_2449_137#_c_1419_n N_RESET_B_M1019_g 0.0150993f $X=15.55 $Y=2.555
+ $X2=0 $Y2=0
cc_1034 N_A_2449_137#_c_1420_n N_RESET_B_M1019_g 0.0101641f $X=15.635 $Y=2.47
+ $X2=0 $Y2=0
cc_1035 N_A_2449_137#_M1021_g N_RESET_B_M1006_g 0.0240812f $X=15.8 $Y=0.705
+ $X2=0 $Y2=0
cc_1036 N_A_2449_137#_c_1410_n N_RESET_B_M1006_g 0.00219674f $X=15.74 $Y=1.49
+ $X2=0 $Y2=0
cc_1037 N_A_2449_137#_c_1412_n N_RESET_B_M1006_g 0.0206453f $X=15.74 $Y=1.4
+ $X2=0 $Y2=0
cc_1038 N_A_2449_137#_M1020_g N_RESET_B_c_1804_n 6.69069e-19 $X=15.77 $Y=2.465
+ $X2=0 $Y2=0
cc_1039 N_A_2449_137#_M1020_g N_RESET_B_c_1805_n 3.11547e-19 $X=15.77 $Y=2.465
+ $X2=0 $Y2=0
cc_1040 N_A_2449_137#_c_1420_n N_RESET_B_c_1805_n 0.00931617f $X=15.635 $Y=2.47
+ $X2=0 $Y2=0
cc_1041 N_A_2449_137#_c_1410_n N_RESET_B_c_1805_n 0.0233352f $X=15.74 $Y=1.49
+ $X2=0 $Y2=0
cc_1042 N_A_2449_137#_c_1412_n N_RESET_B_c_1805_n 3.66753e-19 $X=15.74 $Y=1.4
+ $X2=0 $Y2=0
cc_1043 N_A_2449_137#_c_1402_n N_A_3279_367#_M1023_g 0.0118131f $X=16.755
+ $Y=1.325 $X2=0 $Y2=0
cc_1044 N_A_2449_137#_c_1404_n N_A_3279_367#_M1023_g 0.0136922f $X=16.772
+ $Y=0.78 $X2=0 $Y2=0
cc_1045 N_A_2449_137#_M1002_g N_A_3279_367#_M1004_g 0.0167472f $X=16.755
+ $Y=2.155 $X2=0 $Y2=0
cc_1046 N_A_2449_137#_M1021_g N_A_3279_367#_c_1843_n 0.00227445f $X=15.8
+ $Y=0.705 $X2=0 $Y2=0
cc_1047 N_A_2449_137#_c_1404_n N_A_3279_367#_c_1843_n 0.00298952f $X=16.772
+ $Y=0.78 $X2=0 $Y2=0
cc_1048 N_A_2449_137#_c_1405_n N_A_3279_367#_c_1843_n 0.0177398f $X=16.772
+ $Y=0.93 $X2=0 $Y2=0
cc_1049 N_A_2449_137#_M1020_g N_A_3279_367#_c_1848_n 0.00159595f $X=15.77
+ $Y=2.465 $X2=0 $Y2=0
cc_1050 N_A_2449_137#_M1002_g N_A_3279_367#_c_1848_n 0.0151894f $X=16.755
+ $Y=2.155 $X2=0 $Y2=0
cc_1051 N_A_2449_137#_c_1402_n N_A_3279_367#_c_1844_n 0.00626967f $X=16.755
+ $Y=1.325 $X2=0 $Y2=0
cc_1052 N_A_2449_137#_M1002_g N_A_3279_367#_c_1844_n 0.00918163f $X=16.755
+ $Y=2.155 $X2=0 $Y2=0
cc_1053 N_A_2449_137#_c_1405_n N_A_3279_367#_c_1844_n 9.82692e-19 $X=16.772
+ $Y=0.93 $X2=0 $Y2=0
cc_1054 N_A_2449_137#_c_1406_n N_A_3279_367#_c_1844_n 0.00312825f $X=16.755
+ $Y=1.4 $X2=0 $Y2=0
cc_1055 N_A_2449_137#_c_1402_n N_A_3279_367#_c_1845_n 0.0213474f $X=16.755
+ $Y=1.325 $X2=0 $Y2=0
cc_1056 N_A_2449_137#_c_1401_n N_A_3279_367#_c_1846_n 0.014258f $X=16.68 $Y=1.4
+ $X2=0 $Y2=0
cc_1057 N_A_2449_137#_c_1402_n N_A_3279_367#_c_1846_n 0.00162808f $X=16.755
+ $Y=1.325 $X2=0 $Y2=0
cc_1058 N_A_2449_137#_M1002_g N_A_3279_367#_c_1846_n 0.00337243f $X=16.755
+ $Y=2.155 $X2=0 $Y2=0
cc_1059 N_A_2449_137#_c_1406_n N_A_3279_367#_c_1846_n 3.53117e-19 $X=16.755
+ $Y=1.4 $X2=0 $Y2=0
cc_1060 N_A_2449_137#_c_1416_n N_VPWR_M1037_d 0.00247834f $X=13.535 $Y=2.125
+ $X2=0 $Y2=0
cc_1061 N_A_2449_137#_c_1419_n N_VPWR_M1044_d 0.0058655f $X=15.55 $Y=2.555 $X2=0
+ $Y2=0
cc_1062 N_A_2449_137#_c_1419_n N_VPWR_M1019_d 0.00841372f $X=15.55 $Y=2.555
+ $X2=0 $Y2=0
cc_1063 N_A_2449_137#_c_1420_n N_VPWR_M1019_d 0.00737561f $X=15.635 $Y=2.47
+ $X2=0 $Y2=0
cc_1064 N_A_2449_137#_M1037_g N_VPWR_c_1947_n 0.00715117f $X=12.745 $Y=2.74
+ $X2=0 $Y2=0
cc_1065 N_A_2449_137#_c_1416_n N_VPWR_c_1947_n 0.0202354f $X=13.535 $Y=2.125
+ $X2=0 $Y2=0
cc_1066 N_A_2449_137#_c_1419_n N_VPWR_c_1948_n 0.0198746f $X=15.55 $Y=2.555
+ $X2=0 $Y2=0
cc_1067 N_A_2449_137#_c_1454_n N_VPWR_c_1948_n 0.00819705f $X=13.7 $Y=2.555
+ $X2=0 $Y2=0
cc_1068 N_A_2449_137#_M1020_g N_VPWR_c_1949_n 0.00993676f $X=15.77 $Y=2.465
+ $X2=0 $Y2=0
cc_1069 N_A_2449_137#_c_1419_n N_VPWR_c_1949_n 0.0206531f $X=15.55 $Y=2.555
+ $X2=0 $Y2=0
cc_1070 N_A_2449_137#_M1002_g N_VPWR_c_1950_n 0.00526768f $X=16.755 $Y=2.155
+ $X2=0 $Y2=0
cc_1071 N_A_2449_137#_c_1463_p N_VPWR_c_1957_n 0.00230529f $X=14.05 $Y=2.555
+ $X2=0 $Y2=0
cc_1072 N_A_2449_137#_c_1419_n N_VPWR_c_1957_n 0.00149954f $X=15.55 $Y=2.555
+ $X2=0 $Y2=0
cc_1073 N_A_2449_137#_c_1454_n N_VPWR_c_1957_n 0.0177952f $X=13.7 $Y=2.555 $X2=0
+ $Y2=0
cc_1074 N_A_2449_137#_c_1483_p N_VPWR_c_1957_n 0.00238351f $X=14.135 $Y=2.555
+ $X2=0 $Y2=0
cc_1075 N_A_2449_137#_M1037_g N_VPWR_c_1962_n 0.00570944f $X=12.745 $Y=2.74
+ $X2=0 $Y2=0
cc_1076 N_A_2449_137#_c_1419_n N_VPWR_c_1963_n 0.011951f $X=15.55 $Y=2.555 $X2=0
+ $Y2=0
cc_1077 N_A_2449_137#_M1020_g N_VPWR_c_1964_n 0.00486043f $X=15.77 $Y=2.465
+ $X2=0 $Y2=0
cc_1078 N_A_2449_137#_M1002_g N_VPWR_c_1964_n 0.00312414f $X=16.755 $Y=2.155
+ $X2=0 $Y2=0
cc_1079 N_A_2449_137#_M1011_d N_VPWR_c_1940_n 0.00223819f $X=13.56 $Y=2.255
+ $X2=0 $Y2=0
cc_1080 N_A_2449_137#_M1037_g N_VPWR_c_1940_n 0.00542671f $X=12.745 $Y=2.74
+ $X2=0 $Y2=0
cc_1081 N_A_2449_137#_M1020_g N_VPWR_c_1940_n 0.00954696f $X=15.77 $Y=2.465
+ $X2=0 $Y2=0
cc_1082 N_A_2449_137#_M1002_g N_VPWR_c_1940_n 0.00410284f $X=16.755 $Y=2.155
+ $X2=0 $Y2=0
cc_1083 N_A_2449_137#_c_1463_p N_VPWR_c_1940_n 0.00441867f $X=14.05 $Y=2.555
+ $X2=0 $Y2=0
cc_1084 N_A_2449_137#_c_1419_n N_VPWR_c_1940_n 0.0253849f $X=15.55 $Y=2.555
+ $X2=0 $Y2=0
cc_1085 N_A_2449_137#_c_1454_n N_VPWR_c_1940_n 0.0123247f $X=13.7 $Y=2.555 $X2=0
+ $Y2=0
cc_1086 N_A_2449_137#_c_1483_p N_VPWR_c_1940_n 0.00483686f $X=14.135 $Y=2.555
+ $X2=0 $Y2=0
cc_1087 N_A_2449_137#_c_1408_n A_2798_451# 0.00143151f $X=14.135 $Y=2.47
+ $X2=-0.19 $Y2=-0.245
cc_1088 N_A_2449_137#_c_1483_p A_2798_451# 0.00178582f $X=14.135 $Y=2.555
+ $X2=-0.19 $Y2=-0.245
cc_1089 N_A_2449_137#_M1021_g N_Q_N_c_2304_n 0.0110933f $X=15.8 $Y=0.705 $X2=0
+ $Y2=0
cc_1090 N_A_2449_137#_M1021_g N_Q_N_c_2305_n 0.00287837f $X=15.8 $Y=0.705 $X2=0
+ $Y2=0
cc_1091 N_A_2449_137#_c_1401_n N_Q_N_c_2305_n 0.00487999f $X=16.68 $Y=1.4 $X2=0
+ $Y2=0
cc_1092 N_A_2449_137#_c_1410_n N_Q_N_c_2305_n 0.00425349f $X=15.74 $Y=1.49 $X2=0
+ $Y2=0
cc_1093 N_A_2449_137#_c_1401_n Q_N 0.00638348f $X=16.68 $Y=1.4 $X2=0 $Y2=0
cc_1094 N_A_2449_137#_M1002_g Q_N 0.00198641f $X=16.755 $Y=2.155 $X2=0 $Y2=0
cc_1095 N_A_2449_137#_M1020_g N_Q_N_c_2306_n 0.00251684f $X=15.77 $Y=2.465 $X2=0
+ $Y2=0
cc_1096 N_A_2449_137#_M1021_g N_Q_N_c_2306_n 0.00424694f $X=15.8 $Y=0.705 $X2=0
+ $Y2=0
cc_1097 N_A_2449_137#_c_1401_n N_Q_N_c_2306_n 0.0147906f $X=16.68 $Y=1.4 $X2=0
+ $Y2=0
cc_1098 N_A_2449_137#_M1002_g N_Q_N_c_2306_n 0.00285219f $X=16.755 $Y=2.155
+ $X2=0 $Y2=0
cc_1099 N_A_2449_137#_c_1420_n N_Q_N_c_2306_n 0.00524694f $X=15.635 $Y=2.47
+ $X2=0 $Y2=0
cc_1100 N_A_2449_137#_c_1410_n N_Q_N_c_2306_n 0.0232923f $X=15.74 $Y=1.49 $X2=0
+ $Y2=0
cc_1101 N_A_2449_137#_c_1412_n N_Q_N_c_2306_n 0.00124625f $X=15.74 $Y=1.4 $X2=0
+ $Y2=0
cc_1102 N_A_2449_137#_c_1402_n N_Q_c_2335_n 6.06302e-19 $X=16.755 $Y=1.325 $X2=0
+ $Y2=0
cc_1103 N_A_2449_137#_c_1404_n N_Q_c_2335_n 8.35721e-19 $X=16.772 $Y=0.78 $X2=0
+ $Y2=0
cc_1104 N_A_2449_137#_M1021_g N_VGND_c_2367_n 0.00368477f $X=15.8 $Y=0.705 $X2=0
+ $Y2=0
cc_1105 N_A_2449_137#_c_1410_n N_VGND_c_2367_n 0.00971705f $X=15.74 $Y=1.49
+ $X2=0 $Y2=0
cc_1106 N_A_2449_137#_c_1412_n N_VGND_c_2367_n 0.002179f $X=15.74 $Y=1.4 $X2=0
+ $Y2=0
cc_1107 N_A_2449_137#_c_1404_n N_VGND_c_2368_n 0.0105591f $X=16.772 $Y=0.78
+ $X2=0 $Y2=0
cc_1108 N_A_2449_137#_M1021_g N_VGND_c_2371_n 0.00502664f $X=15.8 $Y=0.705 $X2=0
+ $Y2=0
cc_1109 N_A_2449_137#_c_1404_n N_VGND_c_2371_n 0.00445056f $X=16.772 $Y=0.78
+ $X2=0 $Y2=0
cc_1110 N_A_2449_137#_c_1405_n N_VGND_c_2371_n 6.82495e-19 $X=16.772 $Y=0.93
+ $X2=0 $Y2=0
cc_1111 N_A_2449_137#_c_1397_n N_VGND_c_2379_n 9.72468e-19 $X=12.32 $Y=1.31
+ $X2=0 $Y2=0
cc_1112 N_A_2449_137#_M1021_g N_VGND_c_2379_n 0.0104609f $X=15.8 $Y=0.705 $X2=0
+ $Y2=0
cc_1113 N_A_2449_137#_c_1404_n N_VGND_c_2379_n 0.00899805f $X=16.772 $Y=0.78
+ $X2=0 $Y2=0
cc_1114 N_A_2449_137#_c_1405_n N_VGND_c_2379_n 9.27201e-19 $X=16.772 $Y=0.93
+ $X2=0 $Y2=0
cc_1115 N_A_2449_137#_M1036_d N_A_2636_119#_c_2567_n 0.00587704f $X=13.77
+ $Y=0.595 $X2=0 $Y2=0
cc_1116 N_A_2449_137#_c_1407_n N_A_2636_119#_c_2567_n 0.0178901f $X=13.99
+ $Y=0.935 $X2=0 $Y2=0
cc_1117 N_A_2449_137#_c_1409_n N_A_2636_119#_c_2567_n 0.00122727f $X=14.062
+ $Y=1.255 $X2=0 $Y2=0
cc_1118 N_A_2299_119#_M1036_g N_A_1926_21#_c_1682_n 0.00881852f $X=13.695
+ $Y=0.915 $X2=0 $Y2=0
cc_1119 N_A_2299_119#_c_1615_n N_A_1926_21#_c_1682_n 0.0128253f $X=13.54
+ $Y=0.915 $X2=0 $Y2=0
cc_1120 N_A_2299_119#_c_1584_n N_A_1926_21#_c_1682_n 0.00755492f $X=11.635
+ $Y=0.87 $X2=0 $Y2=0
cc_1121 N_A_2299_119#_M1045_g N_A_1926_21#_M1044_g 0.0484557f $X=13.915 $Y=2.675
+ $X2=0 $Y2=0
cc_1122 N_A_2299_119#_M1036_g N_A_1926_21#_M1017_g 0.0155126f $X=13.695 $Y=0.915
+ $X2=0 $Y2=0
cc_1123 N_A_2299_119#_c_1587_n N_A_1926_21#_c_1688_n 0.0484557f $X=13.705 $Y=1.6
+ $X2=0 $Y2=0
cc_1124 N_A_2299_119#_M1036_g N_A_1926_21#_c_1690_n 0.00106796f $X=13.695
+ $Y=0.915 $X2=0 $Y2=0
cc_1125 N_A_2299_119#_c_1587_n N_A_1926_21#_c_1690_n 0.00146988f $X=13.705
+ $Y=1.6 $X2=0 $Y2=0
cc_1126 N_A_2299_119#_M1045_g N_VPWR_c_1948_n 0.00194884f $X=13.915 $Y=2.675
+ $X2=0 $Y2=0
cc_1127 N_A_2299_119#_M1045_g N_VPWR_c_1957_n 0.0042231f $X=13.915 $Y=2.675
+ $X2=0 $Y2=0
cc_1128 N_A_2299_119#_M1045_g N_VPWR_c_1940_n 0.00581407f $X=13.915 $Y=2.675
+ $X2=0 $Y2=0
cc_1129 N_A_2299_119#_c_1615_n N_VGND_M1025_d 0.0114901f $X=13.54 $Y=0.915 $X2=0
+ $Y2=0
cc_1130 N_A_2299_119#_c_1584_n N_VGND_c_2364_n 0.00862234f $X=11.635 $Y=0.87
+ $X2=0 $Y2=0
cc_1131 N_A_2299_119#_c_1584_n N_VGND_c_2365_n 0.00927944f $X=11.635 $Y=0.87
+ $X2=0 $Y2=0
cc_1132 N_A_2299_119#_c_1615_n N_VGND_c_2366_n 0.0239631f $X=13.54 $Y=0.915
+ $X2=0 $Y2=0
cc_1133 N_A_2299_119#_c_1615_n N_VGND_c_2379_n 0.0326482f $X=13.54 $Y=0.915
+ $X2=0 $Y2=0
cc_1134 N_A_2299_119#_c_1584_n N_VGND_c_2379_n 0.0112444f $X=11.635 $Y=0.87
+ $X2=0 $Y2=0
cc_1135 N_A_2299_119#_c_1615_n A_2401_163# 0.002809f $X=13.54 $Y=0.915 $X2=-0.19
+ $Y2=-0.245
cc_1136 N_A_2299_119#_c_1615_n N_A_2636_119#_M1022_d 0.0122918f $X=13.54
+ $Y=0.915 $X2=-0.19 $Y2=-0.245
cc_1137 N_A_2299_119#_c_1588_n N_A_2636_119#_M1022_d 0.00291866f $X=13.705
+ $Y=1.435 $X2=-0.19 $Y2=-0.245
cc_1138 N_A_2299_119#_M1036_g N_A_2636_119#_c_2567_n 0.00249882f $X=13.695
+ $Y=0.915 $X2=0 $Y2=0
cc_1139 N_A_2299_119#_c_1615_n N_A_2636_119#_c_2567_n 0.00443108f $X=13.54
+ $Y=0.915 $X2=0 $Y2=0
cc_1140 N_A_2299_119#_M1036_g N_A_2636_119#_c_2568_n 7.17317e-19 $X=13.695
+ $Y=0.915 $X2=0 $Y2=0
cc_1141 N_A_2299_119#_M1036_g N_A_2636_119#_c_2569_n 0.0040979f $X=13.695
+ $Y=0.915 $X2=0 $Y2=0
cc_1142 N_A_2299_119#_c_1615_n N_A_2636_119#_c_2569_n 0.0234346f $X=13.54
+ $Y=0.915 $X2=0 $Y2=0
cc_1143 N_A_1926_21#_c_1688_n N_RESET_B_M1019_g 0.00213292f $X=14.565 $Y=1.62
+ $X2=0 $Y2=0
cc_1144 N_A_1926_21#_c_1697_n N_RESET_B_M1019_g 0.00469867f $X=14.565 $Y=1.265
+ $X2=0 $Y2=0
cc_1145 N_A_1926_21#_c_1699_n N_RESET_B_M1019_g 0.00534731f $X=15.045 $Y=2.125
+ $X2=0 $Y2=0
cc_1146 N_A_1926_21#_c_1689_n N_RESET_B_M1006_g 0.00648102f $X=14.565 $Y=1.25
+ $X2=0 $Y2=0
cc_1147 N_A_1926_21#_c_1697_n N_RESET_B_M1006_g 9.66234e-19 $X=14.565 $Y=1.265
+ $X2=0 $Y2=0
cc_1148 N_A_1926_21#_c_1691_n N_RESET_B_M1006_g 0.00603812f $X=14.91 $Y=1.08
+ $X2=0 $Y2=0
cc_1149 N_A_1926_21#_c_1693_n N_RESET_B_M1006_g 0.0146955f $X=15.075 $Y=0.495
+ $X2=0 $Y2=0
cc_1150 N_A_1926_21#_c_1697_n N_RESET_B_c_1804_n 4.04573e-19 $X=14.565 $Y=1.265
+ $X2=0 $Y2=0
cc_1151 N_A_1926_21#_c_1690_n N_RESET_B_c_1804_n 0.0132425f $X=14.565 $Y=1.265
+ $X2=0 $Y2=0
cc_1152 N_A_1926_21#_c_1691_n N_RESET_B_c_1804_n 0.00141132f $X=14.91 $Y=1.08
+ $X2=0 $Y2=0
cc_1153 N_A_1926_21#_c_1699_n N_RESET_B_c_1804_n 7.26845e-19 $X=15.045 $Y=2.125
+ $X2=0 $Y2=0
cc_1154 N_A_1926_21#_c_1697_n N_RESET_B_c_1805_n 0.0242595f $X=14.565 $Y=1.265
+ $X2=0 $Y2=0
cc_1155 N_A_1926_21#_c_1690_n N_RESET_B_c_1805_n 0.00317952f $X=14.565 $Y=1.265
+ $X2=0 $Y2=0
cc_1156 N_A_1926_21#_c_1691_n N_RESET_B_c_1805_n 0.0193651f $X=14.91 $Y=1.08
+ $X2=0 $Y2=0
cc_1157 N_A_1926_21#_c_1699_n N_RESET_B_c_1805_n 0.0140104f $X=15.045 $Y=2.125
+ $X2=0 $Y2=0
cc_1158 N_A_1926_21#_c_1698_n N_VPWR_M1044_d 0.0030328f $X=14.73 $Y=2.125 $X2=0
+ $Y2=0
cc_1159 N_A_1926_21#_M1003_g N_VPWR_c_1946_n 0.020285f $X=10.295 $Y=2.315 $X2=0
+ $Y2=0
cc_1160 N_A_1926_21#_M1044_g N_VPWR_c_1948_n 0.0106437f $X=14.275 $Y=2.675 $X2=0
+ $Y2=0
cc_1161 N_A_1926_21#_M1044_g N_VPWR_c_1957_n 0.00360067f $X=14.275 $Y=2.675
+ $X2=0 $Y2=0
cc_1162 N_A_1926_21#_M1003_g N_VPWR_c_1940_n 7.88961e-19 $X=10.295 $Y=2.315
+ $X2=0 $Y2=0
cc_1163 N_A_1926_21#_M1044_g N_VPWR_c_1940_n 0.00413657f $X=14.275 $Y=2.675
+ $X2=0 $Y2=0
cc_1164 N_A_1926_21#_c_1682_n N_VGND_c_2364_n 0.0211465f $X=14.21 $Y=0.18 $X2=0
+ $Y2=0
cc_1165 N_A_1926_21#_c_1682_n N_VGND_c_2365_n 0.0581842f $X=14.21 $Y=0.18 $X2=0
+ $Y2=0
cc_1166 N_A_1926_21#_c_1682_n N_VGND_c_2366_n 0.0252872f $X=14.21 $Y=0.18 $X2=0
+ $Y2=0
cc_1167 N_A_1926_21#_c_1691_n N_VGND_c_2367_n 0.0118036f $X=14.91 $Y=1.08 $X2=0
+ $Y2=0
cc_1168 N_A_1926_21#_c_1693_n N_VGND_c_2367_n 0.0379291f $X=15.075 $Y=0.495
+ $X2=0 $Y2=0
cc_1169 N_A_1926_21#_c_1683_n N_VGND_c_2376_n 0.0235248f $X=9.78 $Y=0.18 $X2=0
+ $Y2=0
cc_1170 N_A_1926_21#_c_1682_n N_VGND_c_2377_n 0.0328628f $X=14.21 $Y=0.18 $X2=0
+ $Y2=0
cc_1171 N_A_1926_21#_c_1693_n N_VGND_c_2377_n 0.0220321f $X=15.075 $Y=0.495
+ $X2=0 $Y2=0
cc_1172 N_A_1926_21#_c_1682_n N_VGND_c_2379_n 0.121388f $X=14.21 $Y=0.18 $X2=0
+ $Y2=0
cc_1173 N_A_1926_21#_c_1683_n N_VGND_c_2379_n 0.00547013f $X=9.78 $Y=0.18 $X2=0
+ $Y2=0
cc_1174 N_A_1926_21#_c_1693_n N_VGND_c_2379_n 0.0125808f $X=15.075 $Y=0.495
+ $X2=0 $Y2=0
cc_1175 N_A_1926_21#_M1008_g N_A_1752_60#_c_2540_n 5.12695e-19 $X=9.705 $Y=0.65
+ $X2=0 $Y2=0
cc_1176 N_A_1926_21#_M1008_g N_A_1752_60#_c_2537_n 0.0028996f $X=9.705 $Y=0.65
+ $X2=0 $Y2=0
cc_1177 N_A_1926_21#_c_1684_n N_A_1752_60#_c_2537_n 0.00675361f $X=10.22 $Y=1.12
+ $X2=0 $Y2=0
cc_1178 N_A_1926_21#_M1008_g N_A_1752_60#_c_2544_n 0.00854264f $X=9.705 $Y=0.65
+ $X2=0 $Y2=0
cc_1179 N_A_1926_21#_c_1682_n N_A_2636_119#_c_2567_n 0.0104791f $X=14.21 $Y=0.18
+ $X2=0 $Y2=0
cc_1180 N_A_1926_21#_M1017_g N_A_2636_119#_c_2567_n 0.0152145f $X=14.285 $Y=0.67
+ $X2=0 $Y2=0
cc_1181 N_A_1926_21#_c_1693_n N_A_2636_119#_c_2567_n 0.0116404f $X=15.075
+ $Y=0.495 $X2=0 $Y2=0
cc_1182 N_A_1926_21#_M1017_g N_A_2636_119#_c_2568_n 0.0086165f $X=14.285 $Y=0.67
+ $X2=0 $Y2=0
cc_1183 N_A_1926_21#_c_1689_n N_A_2636_119#_c_2568_n 0.00150824f $X=14.565
+ $Y=1.25 $X2=0 $Y2=0
cc_1184 N_A_1926_21#_c_1692_n N_A_2636_119#_c_2568_n 0.0222418f $X=14.73 $Y=1.08
+ $X2=0 $Y2=0
cc_1185 N_A_1926_21#_c_1693_n N_A_2636_119#_c_2568_n 0.0244934f $X=15.075
+ $Y=0.495 $X2=0 $Y2=0
cc_1186 N_A_1926_21#_c_1682_n N_A_2636_119#_c_2569_n 0.00788421f $X=14.21
+ $Y=0.18 $X2=0 $Y2=0
cc_1187 N_A_1926_21#_M1017_g N_A_2636_119#_c_2569_n 0.00133936f $X=14.285
+ $Y=0.67 $X2=0 $Y2=0
cc_1188 N_RESET_B_M1019_g N_VPWR_c_1963_n 5.15685e-19 $X=15.26 $Y=2.155 $X2=0
+ $Y2=0
cc_1189 N_RESET_B_M1006_g N_VGND_c_2367_n 0.00858349f $X=15.29 $Y=0.495 $X2=0
+ $Y2=0
cc_1190 N_RESET_B_M1006_g N_VGND_c_2377_n 0.00502664f $X=15.29 $Y=0.495 $X2=0
+ $Y2=0
cc_1191 N_RESET_B_M1006_g N_VGND_c_2379_n 0.0104609f $X=15.29 $Y=0.495 $X2=0
+ $Y2=0
cc_1192 N_RESET_B_M1006_g N_A_2636_119#_c_2567_n 4.39068e-19 $X=15.29 $Y=0.495
+ $X2=0 $Y2=0
cc_1193 N_RESET_B_M1006_g N_A_2636_119#_c_2568_n 9.46918e-19 $X=15.29 $Y=0.495
+ $X2=0 $Y2=0
cc_1194 N_A_3279_367#_M1004_g N_VPWR_c_1950_n 0.00698192f $X=17.265 $Y=2.465
+ $X2=0 $Y2=0
cc_1195 N_A_3279_367#_c_1848_n N_VPWR_c_1950_n 0.0248129f $X=16.54 $Y=1.98 $X2=0
+ $Y2=0
cc_1196 N_A_3279_367#_c_1844_n N_VPWR_c_1950_n 0.0206753f $X=17.205 $Y=1.47
+ $X2=0 $Y2=0
cc_1197 N_A_3279_367#_c_1845_n N_VPWR_c_1950_n 0.002179f $X=17.205 $Y=1.47 $X2=0
+ $Y2=0
cc_1198 N_A_3279_367#_M1004_g N_VPWR_c_1965_n 0.00549284f $X=17.265 $Y=2.465
+ $X2=0 $Y2=0
cc_1199 N_A_3279_367#_M1004_g N_VPWR_c_1940_n 0.0120439f $X=17.265 $Y=2.465
+ $X2=0 $Y2=0
cc_1200 N_A_3279_367#_c_1848_n N_VPWR_c_1940_n 0.00972751f $X=16.54 $Y=1.98
+ $X2=0 $Y2=0
cc_1201 N_A_3279_367#_c_1843_n N_Q_N_c_2304_n 0.0747023f $X=16.575 $Y=0.495
+ $X2=0 $Y2=0
cc_1202 N_A_3279_367#_c_1848_n N_Q_N_c_2306_n 0.0614497f $X=16.54 $Y=1.98 $X2=0
+ $Y2=0
cc_1203 N_A_3279_367#_c_1846_n N_Q_N_c_2306_n 0.0235793f $X=16.58 $Y=1.47 $X2=0
+ $Y2=0
cc_1204 N_A_3279_367#_M1004_g N_Q_c_2336_n 0.0145249f $X=17.265 $Y=2.465 $X2=0
+ $Y2=0
cc_1205 N_A_3279_367#_M1004_g N_Q_c_2337_n 0.00349143f $X=17.265 $Y=2.465 $X2=0
+ $Y2=0
cc_1206 N_A_3279_367#_c_1845_n N_Q_c_2337_n 0.00131892f $X=17.205 $Y=1.47 $X2=0
+ $Y2=0
cc_1207 N_A_3279_367#_M1023_g N_Q_c_2333_n 0.00448208f $X=17.265 $Y=0.705 $X2=0
+ $Y2=0
cc_1208 N_A_3279_367#_M1004_g N_Q_c_2333_n 0.00448208f $X=17.265 $Y=2.465 $X2=0
+ $Y2=0
cc_1209 N_A_3279_367#_c_1844_n N_Q_c_2333_n 0.0250952f $X=17.205 $Y=1.47 $X2=0
+ $Y2=0
cc_1210 N_A_3279_367#_c_1845_n N_Q_c_2333_n 0.00782465f $X=17.205 $Y=1.47 $X2=0
+ $Y2=0
cc_1211 N_A_3279_367#_M1023_g Q 0.00470167f $X=17.265 $Y=0.705 $X2=0 $Y2=0
cc_1212 N_A_3279_367#_M1023_g N_Q_c_2335_n 0.0131031f $X=17.265 $Y=0.705 $X2=0
+ $Y2=0
cc_1213 N_A_3279_367#_c_1843_n N_Q_c_2335_n 0.0108311f $X=16.575 $Y=0.495 $X2=0
+ $Y2=0
cc_1214 N_A_3279_367#_M1023_g N_VGND_c_2368_n 0.0042292f $X=17.265 $Y=0.705
+ $X2=0 $Y2=0
cc_1215 N_A_3279_367#_c_1843_n N_VGND_c_2368_n 0.017213f $X=16.575 $Y=0.495
+ $X2=0 $Y2=0
cc_1216 N_A_3279_367#_c_1844_n N_VGND_c_2368_n 0.00872859f $X=17.205 $Y=1.47
+ $X2=0 $Y2=0
cc_1217 N_A_3279_367#_c_1845_n N_VGND_c_2368_n 8.63177e-19 $X=17.205 $Y=1.47
+ $X2=0 $Y2=0
cc_1218 N_A_3279_367#_c_1843_n N_VGND_c_2371_n 0.0136872f $X=16.575 $Y=0.495
+ $X2=0 $Y2=0
cc_1219 N_A_3279_367#_M1023_g N_VGND_c_2378_n 0.00502664f $X=17.265 $Y=0.705
+ $X2=0 $Y2=0
cc_1220 N_A_3279_367#_M1023_g N_VGND_c_2379_n 0.0102873f $X=17.265 $Y=0.705
+ $X2=0 $Y2=0
cc_1221 N_A_3279_367#_c_1843_n N_VGND_c_2379_n 0.00785471f $X=16.575 $Y=0.495
+ $X2=0 $Y2=0
cc_1222 N_A_27_474#_c_1894_n N_VPWR_c_1941_n 0.0218522f $X=0.28 $Y=2.515 $X2=0
+ $Y2=0
cc_1223 N_A_27_474#_c_1895_n N_VPWR_c_1941_n 0.0170169f $X=0.975 $Y=2.15 $X2=0
+ $Y2=0
cc_1224 N_A_27_474#_c_1899_n N_VPWR_c_1941_n 0.00891552f $X=1.145 $Y=2.98 $X2=0
+ $Y2=0
cc_1225 N_A_27_474#_c_1898_n N_VPWR_c_1942_n 0.00966617f $X=1.765 $Y=2.98 $X2=0
+ $Y2=0
cc_1226 N_A_27_474#_c_1900_n N_VPWR_c_1942_n 0.0286078f $X=1.93 $Y=2.515 $X2=0
+ $Y2=0
cc_1227 N_A_27_474#_c_1898_n N_VPWR_c_1951_n 0.0590012f $X=1.765 $Y=2.98 $X2=0
+ $Y2=0
cc_1228 N_A_27_474#_c_1899_n N_VPWR_c_1951_n 0.0113756f $X=1.145 $Y=2.98 $X2=0
+ $Y2=0
cc_1229 N_A_27_474#_c_1894_n N_VPWR_c_1959_n 0.0138268f $X=0.28 $Y=2.515 $X2=0
+ $Y2=0
cc_1230 N_A_27_474#_c_1894_n N_VPWR_c_1940_n 0.00942507f $X=0.28 $Y=2.515 $X2=0
+ $Y2=0
cc_1231 N_A_27_474#_c_1898_n N_VPWR_c_1940_n 0.0345757f $X=1.765 $Y=2.98 $X2=0
+ $Y2=0
cc_1232 N_A_27_474#_c_1899_n N_VPWR_c_1940_n 0.00646268f $X=1.145 $Y=2.98 $X2=0
+ $Y2=0
cc_1233 N_A_27_474#_c_1897_n A_200_474# 0.00527525f $X=1.06 $Y=2.895 $X2=-0.19
+ $Y2=1.655
cc_1234 N_A_27_474#_c_1898_n A_200_474# 2.67089e-19 $X=1.765 $Y=2.98 $X2=-0.19
+ $Y2=1.655
cc_1235 N_A_27_474#_c_1898_n N_A_200_119#_M1046_d 0.00180746f $X=1.765 $Y=2.98
+ $X2=0 $Y2=0
cc_1236 N_A_27_474#_c_1895_n N_A_200_119#_c_2132_n 0.00491459f $X=0.975 $Y=2.15
+ $X2=0 $Y2=0
cc_1237 N_A_27_474#_c_1897_n N_A_200_119#_c_2132_n 0.0319857f $X=1.06 $Y=2.895
+ $X2=0 $Y2=0
cc_1238 N_A_27_474#_c_1898_n N_A_200_119#_c_2132_n 0.0136999f $X=1.765 $Y=2.98
+ $X2=0 $Y2=0
cc_1239 N_A_27_474#_c_1900_n N_A_200_119#_c_2132_n 0.01381f $X=1.93 $Y=2.515
+ $X2=0 $Y2=0
cc_1240 N_A_27_474#_c_1900_n N_A_200_119#_c_2133_n 0.0260027f $X=1.93 $Y=2.515
+ $X2=0 $Y2=0
cc_1241 N_A_27_474#_c_1895_n N_A_200_119#_c_2134_n 0.00860182f $X=0.975 $Y=2.15
+ $X2=0 $Y2=0
cc_1242 N_VPWR_c_1942_n N_A_200_119#_c_2133_n 0.00853273f $X=2.48 $Y=2.2 $X2=0
+ $Y2=0
cc_1243 N_VPWR_c_1942_n N_A_200_119#_c_2136_n 0.0136256f $X=2.48 $Y=2.2 $X2=0
+ $Y2=0
cc_1244 N_VPWR_M1047_s N_A_200_119#_c_2137_n 0.00671509f $X=2.34 $Y=2.055 $X2=0
+ $Y2=0
cc_1245 N_VPWR_c_1942_n N_A_200_119#_c_2137_n 0.0604263f $X=2.48 $Y=2.2 $X2=0
+ $Y2=0
cc_1246 N_VPWR_c_1943_n N_A_200_119#_c_2138_n 0.0137879f $X=3.88 $Y=2.39 $X2=0
+ $Y2=0
cc_1247 N_VPWR_c_1953_n N_A_200_119#_c_2138_n 0.0435439f $X=3.795 $Y=3.33 $X2=0
+ $Y2=0
cc_1248 N_VPWR_c_1940_n N_A_200_119#_c_2138_n 0.0263773f $X=17.52 $Y=3.33 $X2=0
+ $Y2=0
cc_1249 N_VPWR_c_1942_n N_A_200_119#_c_2139_n 0.0137879f $X=2.48 $Y=2.2 $X2=0
+ $Y2=0
cc_1250 N_VPWR_c_1953_n N_A_200_119#_c_2139_n 0.0114622f $X=3.795 $Y=3.33 $X2=0
+ $Y2=0
cc_1251 N_VPWR_c_1940_n N_A_200_119#_c_2139_n 0.00657784f $X=17.52 $Y=3.33 $X2=0
+ $Y2=0
cc_1252 N_VPWR_c_1943_n N_A_200_119#_c_2140_n 0.0587853f $X=3.88 $Y=2.39 $X2=0
+ $Y2=0
cc_1253 N_VPWR_c_1943_n N_A_200_119#_c_2141_n 0.013324f $X=3.88 $Y=2.39 $X2=0
+ $Y2=0
cc_1254 N_VPWR_M1029_s N_A_200_119#_c_2143_n 0.00708059f $X=3.735 $Y=2.055 $X2=0
+ $Y2=0
cc_1255 N_VPWR_c_1943_n N_A_200_119#_c_2143_n 0.0579357f $X=3.88 $Y=2.39 $X2=0
+ $Y2=0
cc_1256 N_VPWR_c_1944_n N_A_200_119#_c_2144_n 0.0136002f $X=5.635 $Y=2.84 $X2=0
+ $Y2=0
cc_1257 N_VPWR_c_1960_n N_A_200_119#_c_2144_n 0.0601491f $X=5.47 $Y=3.33 $X2=0
+ $Y2=0
cc_1258 N_VPWR_c_1940_n N_A_200_119#_c_2144_n 0.0365628f $X=17.52 $Y=3.33 $X2=0
+ $Y2=0
cc_1259 N_VPWR_c_1943_n N_A_200_119#_c_2145_n 0.0137879f $X=3.88 $Y=2.39 $X2=0
+ $Y2=0
cc_1260 N_VPWR_c_1960_n N_A_200_119#_c_2145_n 0.0114622f $X=5.47 $Y=3.33 $X2=0
+ $Y2=0
cc_1261 N_VPWR_c_1940_n N_A_200_119#_c_2145_n 0.00657784f $X=17.52 $Y=3.33 $X2=0
+ $Y2=0
cc_1262 N_VPWR_c_1944_n N_A_200_119#_c_2146_n 0.0158804f $X=5.635 $Y=2.84 $X2=0
+ $Y2=0
cc_1263 N_VPWR_M1018_d N_A_200_119#_c_2147_n 0.0102695f $X=5.42 $Y=1.835 $X2=0
+ $Y2=0
cc_1264 N_VPWR_c_1944_n N_A_200_119#_c_2147_n 0.0250423f $X=5.635 $Y=2.84 $X2=0
+ $Y2=0
cc_1265 N_VPWR_c_1940_n N_A_200_119#_c_2147_n 0.0246599f $X=17.52 $Y=3.33 $X2=0
+ $Y2=0
cc_1266 N_VPWR_c_1940_n A_2798_451# 0.00260855f $X=17.52 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_1267 N_VPWR_c_1940_n N_Q_N_M1020_d 0.00419266f $X=17.52 $Y=3.33 $X2=0 $Y2=0
cc_1268 N_VPWR_c_1950_n Q_N 0.0187326f $X=17.05 $Y=1.98 $X2=0 $Y2=0
cc_1269 N_VPWR_c_1964_n Q_N 0.0234637f $X=16.885 $Y=3.33 $X2=0 $Y2=0
cc_1270 N_VPWR_c_1940_n Q_N 0.0136532f $X=17.52 $Y=3.33 $X2=0 $Y2=0
cc_1271 N_VPWR_c_1940_n N_Q_M1004_d 0.0023218f $X=17.52 $Y=3.33 $X2=0 $Y2=0
cc_1272 N_VPWR_c_1965_n N_Q_c_2336_n 0.0214436f $X=17.52 $Y=3.33 $X2=0 $Y2=0
cc_1273 N_VPWR_c_1940_n N_Q_c_2336_n 0.0134754f $X=17.52 $Y=3.33 $X2=0 $Y2=0
cc_1274 N_VPWR_c_1950_n N_Q_c_2337_n 0.045997f $X=17.05 $Y=1.98 $X2=0 $Y2=0
cc_1275 N_A_200_119#_c_2126_n N_VGND_c_2359_n 0.0127019f $X=1.145 $Y=0.805 $X2=0
+ $Y2=0
cc_1276 N_A_200_119#_c_2128_n N_VGND_c_2359_n 0.00568209f $X=1.31 $Y=0.545 $X2=0
+ $Y2=0
cc_1277 N_A_200_119#_c_2127_n N_VGND_c_2360_n 0.013629f $X=2 $Y=0.545 $X2=0
+ $Y2=0
cc_1278 N_A_200_119#_c_2129_n N_VGND_c_2360_n 0.0258118f $X=2.085 $Y=1.685 $X2=0
+ $Y2=0
cc_1279 N_A_200_119#_c_2131_n N_VGND_c_2362_n 0.0111241f $X=6.19 $Y=0.835 $X2=0
+ $Y2=0
cc_1280 N_A_200_119#_c_2127_n N_VGND_c_2373_n 0.024463f $X=2 $Y=0.545 $X2=0
+ $Y2=0
cc_1281 N_A_200_119#_c_2128_n N_VGND_c_2373_n 0.00999549f $X=1.31 $Y=0.545 $X2=0
+ $Y2=0
cc_1282 N_A_200_119#_c_2131_n N_VGND_c_2375_n 0.00691436f $X=6.19 $Y=0.835 $X2=0
+ $Y2=0
cc_1283 N_A_200_119#_c_2127_n N_VGND_c_2379_n 0.024934f $X=2 $Y=0.545 $X2=0
+ $Y2=0
cc_1284 N_A_200_119#_c_2128_n N_VGND_c_2379_n 0.00991134f $X=1.31 $Y=0.545 $X2=0
+ $Y2=0
cc_1285 N_A_200_119#_c_2131_n N_VGND_c_2379_n 0.0087685f $X=6.19 $Y=0.835 $X2=0
+ $Y2=0
cc_1286 N_A_200_119#_c_2127_n A_314_119# 0.00897965f $X=2 $Y=0.545 $X2=-0.19
+ $Y2=-0.245
cc_1287 N_A_200_119#_c_2129_n A_314_119# 0.00452873f $X=2.085 $Y=1.685 $X2=-0.19
+ $Y2=-0.245
cc_1288 N_Q_N_c_2304_n N_VGND_c_2367_n 0.0339633f $X=16.015 $Y=0.43 $X2=0 $Y2=0
cc_1289 N_Q_N_c_2304_n N_VGND_c_2371_n 0.0270889f $X=16.015 $Y=0.43 $X2=0 $Y2=0
cc_1290 N_Q_N_c_2304_n N_VGND_c_2379_n 0.0154828f $X=16.015 $Y=0.43 $X2=0 $Y2=0
cc_1291 N_Q_c_2335_n N_VGND_c_2368_n 0.0283668f $X=17.48 $Y=0.43 $X2=0 $Y2=0
cc_1292 N_Q_c_2335_n N_VGND_c_2378_n 0.0237177f $X=17.48 $Y=0.43 $X2=0 $Y2=0
cc_1293 N_Q_c_2335_n N_VGND_c_2379_n 0.0135481f $X=17.48 $Y=0.43 $X2=0 $Y2=0
cc_1294 N_VGND_c_2377_n N_A_2636_119#_c_2567_n 0.0681098f $X=15.42 $Y=0 $X2=0
+ $Y2=0
cc_1295 N_VGND_c_2379_n N_A_2636_119#_c_2567_n 0.0381807f $X=17.52 $Y=0 $X2=0
+ $Y2=0
cc_1296 N_VGND_c_2366_n N_A_2636_119#_c_2569_n 0.0203686f $X=12.81 $Y=0.485
+ $X2=0 $Y2=0
cc_1297 N_VGND_c_2377_n N_A_2636_119#_c_2569_n 0.0211946f $X=15.42 $Y=0 $X2=0
+ $Y2=0
cc_1298 N_VGND_c_2379_n N_A_2636_119#_c_2569_n 0.0111959f $X=17.52 $Y=0 $X2=0
+ $Y2=0
