* NGSPICE file created from sky130_fd_sc_lp__nor4_2.ext - technology: sky130A

.subckt sky130_fd_sc_lp__nor4_2 A B C D VGND VNB VPB VPWR Y
M1000 VPWR A a_157_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=3.528e+11p pd=3.08e+06u as=7.056e+11p ps=6.16e+06u
M1001 a_74_367# C a_553_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=1.3482e+12p pd=9.7e+06u as=7.056e+11p ps=6.16e+06u
M1002 Y D VGND VNB nshort w=840000u l=150000u
+  ad=9.408e+11p pd=8.96e+06u as=1.3104e+12p ps=1.152e+07u
M1003 VGND B Y VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 Y B VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_157_367# A VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 Y D a_553_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=3.528e+11p pd=3.08e+06u as=0p ps=0u
M1007 a_157_367# B a_74_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_553_367# D Y VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_553_367# C a_74_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND A Y VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND C Y VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 Y C VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VGND D Y VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 Y A VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_74_367# B a_157_367# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

