* File: sky130_fd_sc_lp__and3b_1.pex.spice
* Created: Wed Sep  2 09:32:06 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__AND3B_1%A_N 2 5 9 11 12 13 14 15 21
c27 21 0 1.27661e-19 $X=0.27 $Y=1.005
r28 21 23 46.8028 $w=4.45e-07 $l=1.65e-07 $layer=POLY_cond $X=0.327 $Y=1.005
+ $X2=0.327 $Y2=0.84
r29 14 15 13.755 $w=3.08e-07 $l=3.7e-07 $layer=LI1_cond $X=0.24 $Y=1.665
+ $X2=0.24 $Y2=2.035
r30 13 14 13.755 $w=3.08e-07 $l=3.7e-07 $layer=LI1_cond $X=0.24 $Y=1.295
+ $X2=0.24 $Y2=1.665
r31 12 13 13.755 $w=3.08e-07 $l=3.7e-07 $layer=LI1_cond $X=0.24 $Y=0.925
+ $X2=0.24 $Y2=1.295
r32 12 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.27
+ $Y=1.005 $X2=0.27 $Y2=1.005
r33 9 11 646.085 $w=1.5e-07 $l=1.26e-06 $layer=POLY_cond $X=0.475 $Y=2.77
+ $X2=0.475 $Y2=1.51
r34 5 23 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=0.475 $Y=0.445
+ $X2=0.475 $Y2=0.84
r35 2 11 53.9265 $w=4.45e-07 $l=2.22e-07 $layer=POLY_cond $X=0.327 $Y=1.288
+ $X2=0.327 $Y2=1.51
r36 1 21 7.12377 $w=4.45e-07 $l=5.7e-08 $layer=POLY_cond $X=0.327 $Y=1.062
+ $X2=0.327 $Y2=1.005
r37 1 2 28.2451 $w=4.45e-07 $l=2.26e-07 $layer=POLY_cond $X=0.327 $Y=1.062
+ $X2=0.327 $Y2=1.288
.ends

.subckt PM_SKY130_FD_SC_LP__AND3B_1%A_110_47# 1 2 7 8 11 13 15 20 24 29 30 34 35
r58 34 35 7.92688 $w=2.88e-07 $l=1.65e-07 $layer=LI1_cond $X=0.71 $Y=2.77
+ $X2=0.71 $Y2=2.605
r59 32 35 68.2967 $w=1.88e-07 $l=1.17e-06 $layer=LI1_cond $X=0.66 $Y=1.435
+ $X2=0.66 $Y2=2.605
r60 29 32 17.0441 $w=4.83e-07 $l=5.05e-07 $layer=LI1_cond $X=0.807 $Y=0.93
+ $X2=0.807 $Y2=1.435
r61 29 31 5.98742 $w=4.83e-07 $l=1.65e-07 $layer=LI1_cond $X=0.807 $Y=0.93
+ $X2=0.807 $Y2=0.765
r62 29 30 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.955
+ $Y=0.93 $X2=0.955 $Y2=0.93
r63 24 31 12.7166 $w=2.88e-07 $l=3.2e-07 $layer=LI1_cond $X=0.71 $Y=0.445
+ $X2=0.71 $Y2=0.765
r64 18 30 62.0758 $w=3.3e-07 $l=3.55e-07 $layer=POLY_cond $X=0.955 $Y=1.285
+ $X2=0.955 $Y2=0.93
r65 18 20 158.957 $w=1.5e-07 $l=3.1e-07 $layer=POLY_cond $X=0.955 $Y=1.36
+ $X2=1.265 $Y2=1.36
r66 16 30 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=0.955 $Y=0.915
+ $X2=0.955 $Y2=0.93
r67 13 15 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.445 $Y=0.765
+ $X2=1.445 $Y2=0.445
r68 9 20 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.265 $Y=1.435
+ $X2=1.265 $Y2=1.36
r69 9 11 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.265 $Y=1.435
+ $X2=1.265 $Y2=2.045
r70 8 16 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=1.12 $Y=0.84
+ $X2=0.955 $Y2=0.915
r71 7 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.37 $Y=0.84
+ $X2=1.445 $Y2=0.765
r72 7 8 128.191 $w=1.5e-07 $l=2.5e-07 $layer=POLY_cond $X=1.37 $Y=0.84 $X2=1.12
+ $Y2=0.84
r73 2 34 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=2.56 $X2=0.69 $Y2=2.77
r74 1 24 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.235 $X2=0.69 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__AND3B_1%B 3 7 9 10 11 16
c37 9 0 1.91367e-19 $X=1.68 $Y=0.555
r38 16 19 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.715 $Y=1.32
+ $X2=1.715 $Y2=1.485
r39 16 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.715 $Y=1.32
+ $X2=1.715 $Y2=1.155
r40 11 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.715
+ $Y=1.32 $X2=1.715 $Y2=1.32
r41 10 11 14.4544 $w=2.93e-07 $l=3.7e-07 $layer=LI1_cond $X=1.712 $Y=0.925
+ $X2=1.712 $Y2=1.295
r42 9 10 14.4544 $w=2.93e-07 $l=3.7e-07 $layer=LI1_cond $X=1.712 $Y=0.555
+ $X2=1.712 $Y2=0.925
r43 7 18 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=1.805 $Y=0.445
+ $X2=1.805 $Y2=1.155
r44 3 19 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=1.78 $Y=2.045
+ $X2=1.78 $Y2=1.485
.ends

.subckt PM_SKY130_FD_SC_LP__AND3B_1%C 3 6 9 10 11 12 13 14 19
c40 12 0 8.69356e-20 $X=2.16 $Y=0.555
c41 6 0 1.91367e-19 $X=2.245 $Y=2.045
r42 19 20 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.255
+ $Y=0.93 $X2=2.255 $Y2=0.93
r43 14 20 13.5691 $w=3.08e-07 $l=3.65e-07 $layer=LI1_cond $X=2.185 $Y=1.295
+ $X2=2.185 $Y2=0.93
r44 13 20 0.185878 $w=3.08e-07 $l=5e-09 $layer=LI1_cond $X=2.185 $Y=0.925
+ $X2=2.185 $Y2=0.93
r45 12 13 13.755 $w=3.08e-07 $l=3.7e-07 $layer=LI1_cond $X=2.185 $Y=0.555
+ $X2=2.185 $Y2=0.925
r46 10 19 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.255 $Y=1.27
+ $X2=2.255 $Y2=0.93
r47 10 11 38.0424 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.255 $Y=1.27
+ $X2=2.255 $Y2=1.435
r48 9 19 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.255 $Y=0.765
+ $X2=2.255 $Y2=0.93
r49 6 11 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.245 $Y=2.045
+ $X2=2.245 $Y2=1.435
r50 3 9 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.165 $Y=0.445
+ $X2=2.165 $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_LP__AND3B_1%A_185_367# 1 2 3 12 16 20 23 24 25 30 38 40
+ 42 43
c79 43 0 1.93477e-19 $X=2.795 $Y=1.505
r80 43 47 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.795 $Y=1.505
+ $X2=2.795 $Y2=1.67
r81 43 46 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.795 $Y=1.505
+ $X2=2.795 $Y2=1.34
r82 42 43 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.795
+ $Y=1.505 $X2=2.795 $Y2=1.505
r83 36 38 2.90945 $w=3.03e-07 $l=7.7e-08 $layer=LI1_cond $X=1.23 $Y=0.432
+ $X2=1.307 $Y2=0.432
r84 31 40 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=2.125 $Y=1.76
+ $X2=1.99 $Y2=1.76
r85 30 42 10.5816 $w=2.94e-07 $l=3.33054e-07 $layer=LI1_cond $X=2.53 $Y=1.76
+ $X2=2.71 $Y2=1.505
r86 30 31 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=2.53 $Y=1.76
+ $X2=2.125 $Y2=1.76
r87 26 40 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.99 $Y=1.845
+ $X2=1.99 $Y2=1.76
r88 26 28 8.53661 $w=2.68e-07 $l=2e-07 $layer=LI1_cond $X=1.99 $Y=1.845 $X2=1.99
+ $Y2=2.045
r89 25 34 5.74118 $w=1.68e-07 $l=8.8e-08 $layer=LI1_cond $X=1.395 $Y=1.76
+ $X2=1.307 $Y2=1.76
r90 24 40 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=1.855 $Y=1.76
+ $X2=1.99 $Y2=1.76
r91 24 25 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=1.855 $Y=1.76
+ $X2=1.395 $Y2=1.76
r92 23 34 0.574824 $w=1.75e-07 $l=8.5e-08 $layer=LI1_cond $X=1.307 $Y=1.675
+ $X2=1.307 $Y2=1.76
r93 22 38 4.00781 $w=1.75e-07 $l=1.53e-07 $layer=LI1_cond $X=1.307 $Y=0.585
+ $X2=1.307 $Y2=0.432
r94 22 23 69.0805 $w=1.73e-07 $l=1.09e-06 $layer=LI1_cond $X=1.307 $Y=0.585
+ $X2=1.307 $Y2=1.675
r95 18 34 16.4406 $w=1.68e-07 $l=2.52e-07 $layer=LI1_cond $X=1.055 $Y=1.76
+ $X2=1.307 $Y2=1.76
r96 18 20 8.86495 $w=2.58e-07 $l=2e-07 $layer=LI1_cond $X=1.055 $Y=1.845
+ $X2=1.055 $Y2=2.045
r97 16 46 351.245 $w=1.5e-07 $l=6.85e-07 $layer=POLY_cond $X=2.87 $Y=0.655
+ $X2=2.87 $Y2=1.34
r98 12 47 407.649 $w=1.5e-07 $l=7.95e-07 $layer=POLY_cond $X=2.77 $Y=2.465
+ $X2=2.77 $Y2=1.67
r99 3 28 600 $w=1.7e-07 $l=2.78747e-07 $layer=licon1_PDIFF $count=1 $X=1.855
+ $Y=1.835 $X2=2.015 $Y2=2.045
r100 2 20 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=0.925
+ $Y=1.835 $X2=1.05 $Y2=2.045
r101 1 36 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=1.105
+ $Y=0.235 $X2=1.23 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__AND3B_1%VPWR 1 2 3 10 12 16 20 25 26 28 29 30 40 41
c35 20 0 1.06542e-19 $X=2.46 $Y=2.1
r36 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r37 40 41 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r38 38 41 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r39 37 38 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r40 35 45 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.24 $Y2=3.33
r41 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r42 32 44 4.49698 $w=1.7e-07 $l=1.98e-07 $layer=LI1_cond $X=0.395 $Y=3.33
+ $X2=0.197 $Y2=3.33
r43 32 34 52.5187 $w=1.68e-07 $l=8.05e-07 $layer=LI1_cond $X=0.395 $Y=3.33
+ $X2=1.2 $Y2=3.33
r44 30 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r45 30 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r46 28 37 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=2.295 $Y=3.33
+ $X2=2.16 $Y2=3.33
r47 28 29 9.23004 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=2.295 $Y=3.33
+ $X2=2.477 $Y2=3.33
r48 27 40 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=2.66 $Y=3.33
+ $X2=3.12 $Y2=3.33
r49 27 29 9.23004 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=2.66 $Y=3.33
+ $X2=2.477 $Y2=3.33
r50 25 34 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=1.355 $Y=3.33
+ $X2=1.2 $Y2=3.33
r51 25 26 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.355 $Y=3.33
+ $X2=1.52 $Y2=3.33
r52 24 37 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=1.685 $Y=3.33
+ $X2=2.16 $Y2=3.33
r53 24 26 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.685 $Y=3.33
+ $X2=1.52 $Y2=3.33
r54 20 23 14.5239 $w=3.63e-07 $l=4.6e-07 $layer=LI1_cond $X=2.477 $Y=2.1
+ $X2=2.477 $Y2=2.56
r55 18 29 1.2012 $w=3.65e-07 $l=8.5e-08 $layer=LI1_cond $X=2.477 $Y=3.245
+ $X2=2.477 $Y2=3.33
r56 18 23 21.628 $w=3.63e-07 $l=6.85e-07 $layer=LI1_cond $X=2.477 $Y=3.245
+ $X2=2.477 $Y2=2.56
r57 14 26 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.52 $Y=3.245
+ $X2=1.52 $Y2=3.33
r58 14 16 38.9386 $w=3.28e-07 $l=1.115e-06 $layer=LI1_cond $X=1.52 $Y=3.245
+ $X2=1.52 $Y2=2.13
r59 10 44 3.0207 $w=3e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.245 $Y=3.245
+ $X2=0.197 $Y2=3.33
r60 10 12 18.247 $w=2.98e-07 $l=4.75e-07 $layer=LI1_cond $X=0.245 $Y=3.245
+ $X2=0.245 $Y2=2.77
r61 3 23 300 $w=1.7e-07 $l=8.34266e-07 $layer=licon1_PDIFF $count=2 $X=2.32
+ $Y=1.835 $X2=2.555 $Y2=2.56
r62 3 20 600 $w=1.7e-07 $l=3.27605e-07 $layer=licon1_PDIFF $count=1 $X=2.32
+ $Y=1.835 $X2=2.46 $Y2=2.1
r63 2 16 600 $w=1.7e-07 $l=3.74333e-07 $layer=licon1_PDIFF $count=1 $X=1.34
+ $Y=1.835 $X2=1.52 $Y2=2.13
r64 1 12 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.56 $X2=0.26 $Y2=2.77
.ends

.subckt PM_SKY130_FD_SC_LP__AND3B_1%X 1 2 9 13 14 15 16 31 35
r18 33 35 0.583515 $w=3.93e-07 $l=2e-08 $layer=LI1_cond $X=3.077 $Y=2.015
+ $X2=3.077 $Y2=2.035
r19 21 35 0.350109 $w=3.93e-07 $l=1.2e-08 $layer=LI1_cond $X=3.077 $Y=2.047
+ $X2=3.077 $Y2=2.035
r20 16 28 3.93873 $w=3.93e-07 $l=1.35e-07 $layer=LI1_cond $X=3.077 $Y=2.775
+ $X2=3.077 $Y2=2.91
r21 15 16 10.795 $w=3.93e-07 $l=3.7e-07 $layer=LI1_cond $X=3.077 $Y=2.405
+ $X2=3.077 $Y2=2.775
r22 14 33 0.495988 $w=3.93e-07 $l=1.7e-08 $layer=LI1_cond $X=3.077 $Y=1.998
+ $X2=3.077 $Y2=2.015
r23 14 31 6.6945 $w=3.93e-07 $l=1.48e-07 $layer=LI1_cond $X=3.077 $Y=1.998
+ $X2=3.077 $Y2=1.85
r24 14 15 9.3946 $w=3.93e-07 $l=3.22e-07 $layer=LI1_cond $X=3.077 $Y=2.083
+ $X2=3.077 $Y2=2.405
r25 14 21 1.05033 $w=3.93e-07 $l=3.6e-08 $layer=LI1_cond $X=3.077 $Y=2.083
+ $X2=3.077 $Y2=2.047
r26 13 31 40.4695 $w=2.13e-07 $l=7.55e-07 $layer=LI1_cond $X=3.167 $Y=1.095
+ $X2=3.167 $Y2=1.85
r27 7 13 6.46398 $w=2.83e-07 $l=1.42e-07 $layer=LI1_cond $X=3.132 $Y=0.953
+ $X2=3.132 $Y2=1.095
r28 7 9 21.5527 $w=2.83e-07 $l=5.33e-07 $layer=LI1_cond $X=3.132 $Y=0.953
+ $X2=3.132 $Y2=0.42
r29 2 33 400 $w=1.7e-07 $l=2.4e-07 $layer=licon1_PDIFF $count=1 $X=2.845
+ $Y=1.835 $X2=2.985 $Y2=2.015
r30 2 28 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=2.845
+ $Y=1.835 $X2=2.985 $Y2=2.91
r31 1 9 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=2.945
+ $Y=0.235 $X2=3.085 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__AND3B_1%VGND 1 2 7 9 13 17 19 29 30 36
c50 30 0 1.27661e-19 $X=3.12 $Y=0
r51 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r52 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r53 30 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.64
+ $Y2=0
r54 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r55 27 36 8.23795 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=2.82 $Y=0 $X2=2.665
+ $Y2=0
r56 27 29 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=2.82 $Y=0 $X2=3.12
+ $Y2=0
r57 26 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r58 25 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r59 23 34 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r60 22 25 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=0.72 $Y=0 $X2=2.16
+ $Y2=0
r61 22 23 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r62 20 33 4.49698 $w=1.7e-07 $l=1.98e-07 $layer=LI1_cond $X=0.395 $Y=0 $X2=0.197
+ $Y2=0
r63 20 22 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.395 $Y=0 $X2=0.72
+ $Y2=0
r64 19 36 8.23795 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=2.51 $Y=0 $X2=2.665
+ $Y2=0
r65 19 25 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=2.51 $Y=0 $X2=2.16
+ $Y2=0
r66 17 26 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r67 17 23 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=0.72
+ $Y2=0
r68 13 15 20.4466 $w=3.08e-07 $l=5.5e-07 $layer=LI1_cond $X=2.665 $Y=0.38
+ $X2=2.665 $Y2=0.93
r69 11 36 0.701276 $w=3.1e-07 $l=8.5e-08 $layer=LI1_cond $X=2.665 $Y=0.085
+ $X2=2.665 $Y2=0
r70 11 13 10.9668 $w=3.08e-07 $l=2.95e-07 $layer=LI1_cond $X=2.665 $Y=0.085
+ $X2=2.665 $Y2=0.38
r71 7 33 3.0207 $w=3e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.245 $Y=0.085
+ $X2=0.197 $Y2=0
r72 7 9 13.8293 $w=2.98e-07 $l=3.6e-07 $layer=LI1_cond $X=0.245 $Y=0.085
+ $X2=0.245 $Y2=0.445
r73 2 15 182 $w=1.7e-07 $l=8.78322e-07 $layer=licon1_NDIFF $count=1 $X=2.24
+ $Y=0.235 $X2=2.655 $Y2=0.93
r74 2 13 182 $w=1.7e-07 $l=4.21307e-07 $layer=licon1_NDIFF $count=1 $X=2.24
+ $Y=0.235 $X2=2.595 $Y2=0.38
r75 1 9 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.445
.ends

