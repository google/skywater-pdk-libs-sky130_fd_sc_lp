* File: sky130_fd_sc_lp__a2111o_lp.pex.spice
* Created: Fri Aug 28 09:46:11 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A2111O_LP%D1 3 7 9 13 16 19 20 21 25 26
r47 25 26 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.365
+ $Y=1.02 $X2=0.365 $Y2=1.02
r48 20 21 10.5285 $w=4.03e-07 $l=3.7e-07 $layer=LI1_cond $X=0.327 $Y=1.295
+ $X2=0.327 $Y2=1.665
r49 20 26 7.82523 $w=4.03e-07 $l=2.75e-07 $layer=LI1_cond $X=0.327 $Y=1.295
+ $X2=0.327 $Y2=1.02
r50 18 25 55.3649 $w=3.7e-07 $l=3.55e-07 $layer=POLY_cond $X=0.385 $Y=1.375
+ $X2=0.385 $Y2=1.02
r51 18 19 29.492 $w=3.7e-07 $l=1.5e-07 $layer=POLY_cond $X=0.435 $Y=1.375
+ $X2=0.435 $Y2=1.525
r52 15 25 13.2564 $w=3.7e-07 $l=8.5e-08 $layer=POLY_cond $X=0.385 $Y=0.935
+ $X2=0.385 $Y2=1.02
r53 15 16 12.6443 $w=2.6e-07 $l=7.5e-08 $layer=POLY_cond $X=0.385 $Y=0.935
+ $X2=0.385 $Y2=0.86
r54 11 13 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=0.885 $Y=0.785
+ $X2=0.885 $Y2=0.445
r55 10 16 13.3547 $w=1.5e-07 $l=1.85e-07 $layer=POLY_cond $X=0.57 $Y=0.86
+ $X2=0.385 $Y2=0.86
r56 9 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.81 $Y=0.86
+ $X2=0.885 $Y2=0.785
r57 9 10 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=0.81 $Y=0.86 $X2=0.57
+ $Y2=0.86
r58 7 19 253.423 $w=2.5e-07 $l=1.02e-06 $layer=POLY_cond $X=0.545 $Y=2.545
+ $X2=0.545 $Y2=1.525
r59 1 16 12.6443 $w=2.6e-07 $l=1.42653e-07 $layer=POLY_cond $X=0.495 $Y=0.785
+ $X2=0.385 $Y2=0.86
r60 1 3 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=0.495 $Y=0.785
+ $X2=0.495 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__A2111O_LP%C1 3 5 7 10 12 14 15 16 17 21 23
r56 21 24 68.5216 $w=4.8e-07 $l=5.05e-07 $layer=POLY_cond $X=1.15 $Y=1.34
+ $X2=1.15 $Y2=1.845
r57 21 23 45.9721 $w=4.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.15 $Y=1.34
+ $X2=1.15 $Y2=1.175
r58 16 17 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.225 $Y=1.295
+ $X2=1.225 $Y2=1.665
r59 16 21 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.225
+ $Y=1.34 $X2=1.225 $Y2=1.34
r60 12 14 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=1.675 $Y=0.73
+ $X2=1.675 $Y2=0.445
r61 11 15 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.39 $Y=0.805
+ $X2=1.315 $Y2=0.805
r62 10 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.6 $Y=0.805
+ $X2=1.675 $Y2=0.73
r63 10 11 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=1.6 $Y=0.805
+ $X2=1.39 $Y2=0.805
r64 8 15 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.315 $Y=0.88
+ $X2=1.315 $Y2=0.805
r65 8 23 151.266 $w=1.5e-07 $l=2.95e-07 $layer=POLY_cond $X=1.315 $Y=0.88
+ $X2=1.315 $Y2=1.175
r66 5 15 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.315 $Y=0.73
+ $X2=1.315 $Y2=0.805
r67 5 7 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=1.315 $Y=0.73 $X2=1.315
+ $Y2=0.445
r68 3 24 173.918 $w=2.5e-07 $l=7e-07 $layer=POLY_cond $X=1.035 $Y=2.545
+ $X2=1.035 $Y2=1.845
.ends

.subckt PM_SKY130_FD_SC_LP__A2111O_LP%A_27_409# 1 2 3 4 15 19 23 25 27 29 33 36
+ 37 41 46 50 52 56 60 62 64 68
r136 67 68 14.3881 $w=6.7e-07 $l=2e-07 $layer=POLY_cond $X=2.265 $Y=1.307
+ $X2=2.465 $Y2=1.307
r137 63 68 20.503 $w=6.7e-07 $l=2.85e-07 $layer=POLY_cond $X=2.75 $Y=1.307
+ $X2=2.465 $Y2=1.307
r138 62 63 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.75
+ $Y=0.99 $X2=2.75 $Y2=0.99
r139 54 56 11.5244 $w=3.28e-07 $l=3.3e-07 $layer=LI1_cond $X=4.87 $Y=0.825
+ $X2=4.87 $Y2=0.495
r140 53 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.425 $Y=0.91
+ $X2=3.26 $Y2=0.91
r141 52 54 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.705 $Y=0.91
+ $X2=4.87 $Y2=0.825
r142 52 53 83.508 $w=1.68e-07 $l=1.28e-06 $layer=LI1_cond $X=4.705 $Y=0.91
+ $X2=3.425 $Y2=0.91
r143 48 64 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.26 $Y=0.825
+ $X2=3.26 $Y2=0.91
r144 48 50 11.5244 $w=3.28e-07 $l=3.3e-07 $layer=LI1_cond $X=3.26 $Y=0.825
+ $X2=3.26 $Y2=0.495
r145 47 62 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.915 $Y=0.91
+ $X2=2.75 $Y2=0.91
r146 46 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.095 $Y=0.91
+ $X2=3.26 $Y2=0.91
r147 46 47 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=3.095 $Y=0.91
+ $X2=2.915 $Y2=0.91
r148 41 42 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.89
+ $Y=1.285 $X2=1.89 $Y2=1.285
r149 39 41 10.1275 $w=3.28e-07 $l=2.9e-07 $layer=LI1_cond $X=1.89 $Y=0.995
+ $X2=1.89 $Y2=1.285
r150 38 60 4.16724 $w=1.7e-07 $l=2.78e-07 $layer=LI1_cond $X=1.265 $Y=0.91
+ $X2=0.987 $Y2=0.91
r151 37 39 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.725 $Y=0.91
+ $X2=1.89 $Y2=0.995
r152 37 38 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=1.725 $Y=0.91
+ $X2=1.265 $Y2=0.91
r153 35 60 2.64909 $w=3.62e-07 $l=2.30617e-07 $layer=LI1_cond $X=0.795 $Y=0.995
+ $X2=0.987 $Y2=0.91
r154 35 36 67.1979 $w=1.68e-07 $l=1.03e-06 $layer=LI1_cond $X=0.795 $Y=0.995
+ $X2=0.795 $Y2=2.025
r155 31 60 2.64909 $w=3.62e-07 $l=8.5e-08 $layer=LI1_cond $X=0.987 $Y=0.825
+ $X2=0.987 $Y2=0.91
r156 31 33 7.65059 $w=5.53e-07 $l=3.55e-07 $layer=LI1_cond $X=0.987 $Y=0.825
+ $X2=0.987 $Y2=0.47
r157 30 59 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.445 $Y=2.11
+ $X2=0.28 $Y2=2.11
r158 29 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.71 $Y=2.11
+ $X2=0.795 $Y2=2.025
r159 29 30 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.71 $Y=2.11
+ $X2=0.445 $Y2=2.11
r160 25 59 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.28 $Y=2.195
+ $X2=0.28 $Y2=2.11
r161 25 27 24.6204 $w=3.28e-07 $l=7.05e-07 $layer=LI1_cond $X=0.28 $Y=2.195
+ $X2=0.28 $Y2=2.9
r162 21 68 38.9565 $w=1.5e-07 $l=4.82e-07 $layer=POLY_cond $X=2.465 $Y=0.825
+ $X2=2.465 $Y2=1.307
r163 21 23 194.851 $w=1.5e-07 $l=3.8e-07 $layer=POLY_cond $X=2.465 $Y=0.825
+ $X2=2.465 $Y2=0.445
r164 17 67 25.9839 $w=2.5e-07 $l=4.83e-07 $layer=POLY_cond $X=2.265 $Y=1.79
+ $X2=2.265 $Y2=1.307
r165 17 19 163.979 $w=2.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.265 $Y=1.79
+ $X2=2.265 $Y2=2.45
r166 13 67 11.5104 $w=6.7e-07 $l=1.6e-07 $layer=POLY_cond $X=2.105 $Y=1.307
+ $X2=2.265 $Y2=1.307
r167 13 42 15.4672 $w=6.7e-07 $l=2.15e-07 $layer=POLY_cond $X=2.105 $Y=1.307
+ $X2=1.89 $Y2=1.307
r168 13 15 346.117 $w=1.5e-07 $l=6.75e-07 $layer=POLY_cond $X=2.105 $Y=1.12
+ $X2=2.105 $Y2=0.445
r169 4 59 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.045 $X2=0.28 $Y2=2.19
r170 4 27 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.045 $X2=0.28 $Y2=2.9
r171 3 56 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=4.73
+ $Y=0.285 $X2=4.87 $Y2=0.495
r172 2 50 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=3.115
+ $Y=0.285 $X2=3.26 $Y2=0.495
r173 1 33 182 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=1 $X=0.96
+ $Y=0.235 $X2=1.1 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_LP__A2111O_LP%B1 1 3 8 10 12 14 16 17 18 19 20 21 25
r60 20 21 12.183 $w=3.48e-07 $l=3.7e-07 $layer=LI1_cond $X=3.54 $Y=1.295
+ $X2=3.54 $Y2=1.665
r61 20 25 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.53
+ $Y=1.34 $X2=3.53 $Y2=1.34
r62 17 25 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=3.53 $Y=1.68
+ $X2=3.53 $Y2=1.34
r63 17 18 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.53 $Y=1.68
+ $X2=3.53 $Y2=1.845
r64 16 25 41.3509 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.53 $Y=1.175
+ $X2=3.53 $Y2=1.34
r65 12 14 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.835 $Y=0.78
+ $X2=3.835 $Y2=0.495
r66 11 19 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.55 $Y=0.855
+ $X2=3.475 $Y2=0.855
r67 10 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.76 $Y=0.855
+ $X2=3.835 $Y2=0.78
r68 10 11 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=3.76 $Y=0.855
+ $X2=3.55 $Y2=0.855
r69 8 18 173.918 $w=2.5e-07 $l=7e-07 $layer=POLY_cond $X=3.57 $Y=2.545 $X2=3.57
+ $Y2=1.845
r70 4 19 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.475 $Y=0.93
+ $X2=3.475 $Y2=0.855
r71 4 16 125.628 $w=1.5e-07 $l=2.45e-07 $layer=POLY_cond $X=3.475 $Y=0.93
+ $X2=3.475 $Y2=1.175
r72 1 19 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.475 $Y=0.78
+ $X2=3.475 $Y2=0.855
r73 1 3 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.475 $Y=0.78 $X2=3.475
+ $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__A2111O_LP%A2 2 5 9 11 12 13 17
c43 5 0 2.34935e-19 $X=4.1 $Y=2.545
r44 17 19 45.79 $w=4.05e-07 $l=1.65e-07 $layer=POLY_cond $X=4.137 $Y=1.34
+ $X2=4.137 $Y2=1.175
r45 12 13 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=4.1 $Y=1.295 $X2=4.1
+ $Y2=1.665
r46 12 17 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.1 $Y=1.34
+ $X2=4.1 $Y2=1.34
r47 9 19 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=4.265 $Y=0.495
+ $X2=4.265 $Y2=1.175
r48 5 11 173.918 $w=2.5e-07 $l=7e-07 $layer=POLY_cond $X=4.1 $Y=2.545 $X2=4.1
+ $Y2=1.845
r49 2 11 33.0779 $w=4.05e-07 $l=2.02e-07 $layer=POLY_cond $X=4.137 $Y=1.643
+ $X2=4.137 $Y2=1.845
r50 1 17 5.08091 $w=4.05e-07 $l=3.7e-08 $layer=POLY_cond $X=4.137 $Y=1.377
+ $X2=4.137 $Y2=1.34
r51 1 2 36.5276 $w=4.05e-07 $l=2.66e-07 $layer=POLY_cond $X=4.137 $Y=1.377
+ $X2=4.137 $Y2=1.643
.ends

.subckt PM_SKY130_FD_SC_LP__A2111O_LP%A1 3 7 11 12 13 15 22
r33 22 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.745
+ $Y=1.34 $X2=4.745 $Y2=1.34
r34 15 23 5.26632 $w=6.68e-07 $l=2.95e-07 $layer=LI1_cond $X=5.04 $Y=1.51
+ $X2=4.745 $Y2=1.51
r35 13 23 3.3026 $w=6.68e-07 $l=1.85e-07 $layer=LI1_cond $X=4.56 $Y=1.51
+ $X2=4.745 $Y2=1.51
r36 11 22 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=4.745 $Y=1.68
+ $X2=4.745 $Y2=1.34
r37 11 12 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.745 $Y=1.68
+ $X2=4.745 $Y2=1.845
r38 10 22 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.745 $Y=1.175
+ $X2=4.745 $Y2=1.34
r39 7 12 173.918 $w=2.5e-07 $l=7e-07 $layer=POLY_cond $X=4.705 $Y=2.545
+ $X2=4.705 $Y2=1.845
r40 3 10 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=4.655 $Y=0.495
+ $X2=4.655 $Y2=1.175
.ends

.subckt PM_SKY130_FD_SC_LP__A2111O_LP%A_232_409# 1 2 9 13 15 19 23 25 26
c40 26 0 1.25754e-19 $X=3.305 $Y=2.445
c41 25 0 1.25754e-19 $X=1.3 $Y=2.445
c42 23 0 1.43055e-19 $X=3.305 $Y=2.9
c43 19 0 9.18794e-20 $X=3.305 $Y=2.19
r44 21 26 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.305 $Y=2.53
+ $X2=3.305 $Y2=2.445
r45 21 23 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=3.305 $Y=2.53
+ $X2=3.305 $Y2=2.9
r46 17 26 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.305 $Y=2.36
+ $X2=3.305 $Y2=2.445
r47 17 19 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=3.305 $Y=2.36
+ $X2=3.305 $Y2=2.19
r48 16 25 3.80956 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.465 $Y=2.445
+ $X2=1.3 $Y2=2.445
r49 15 26 3.80956 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.14 $Y=2.445
+ $X2=3.305 $Y2=2.445
r50 15 16 109.278 $w=1.68e-07 $l=1.675e-06 $layer=LI1_cond $X=3.14 $Y=2.445
+ $X2=1.465 $Y2=2.445
r51 11 25 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.3 $Y=2.53 $X2=1.3
+ $Y2=2.445
r52 11 13 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=1.3 $Y=2.53 $X2=1.3
+ $Y2=2.9
r53 7 25 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.3 $Y=2.36 $X2=1.3
+ $Y2=2.445
r54 7 9 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=1.3 $Y=2.36 $X2=1.3
+ $Y2=2.19
r55 2 23 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=3.16
+ $Y=2.045 $X2=3.305 $Y2=2.9
r56 2 19 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=3.16
+ $Y=2.045 $X2=3.305 $Y2=2.19
r57 1 13 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=1.16
+ $Y=2.045 $X2=1.3 $Y2=2.9
r58 1 9 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.16
+ $Y=2.045 $X2=1.3 $Y2=2.19
.ends

.subckt PM_SKY130_FD_SC_LP__A2111O_LP%VPWR 1 2 9 13 16 17 18 20 33 34 37
r44 37 38 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r45 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r46 31 34 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=5.04 $Y2=3.33
r47 30 31 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r48 28 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.165 $Y=3.33 $X2=2
+ $Y2=3.33
r49 28 30 124.936 $w=1.68e-07 $l=1.915e-06 $layer=LI1_cond $X=2.165 $Y=3.33
+ $X2=4.08 $Y2=3.33
r50 27 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r51 26 27 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r52 23 27 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.68 $Y2=3.33
r53 22 26 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=0.24 $Y=3.33
+ $X2=1.68 $Y2=3.33
r54 22 23 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r55 20 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.835 $Y=3.33 $X2=2
+ $Y2=3.33
r56 20 26 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=1.835 $Y=3.33
+ $X2=1.68 $Y2=3.33
r57 18 31 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=4.08 $Y2=3.33
r58 18 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r59 16 30 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=4.2 $Y=3.33 $X2=4.08
+ $Y2=3.33
r60 16 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.2 $Y=3.33
+ $X2=4.365 $Y2=3.33
r61 15 33 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=4.53 $Y=3.33
+ $X2=5.04 $Y2=3.33
r62 15 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.53 $Y=3.33
+ $X2=4.365 $Y2=3.33
r63 11 17 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.365 $Y=3.245
+ $X2=4.365 $Y2=3.33
r64 11 13 24.6204 $w=3.28e-07 $l=7.05e-07 $layer=LI1_cond $X=4.365 $Y=3.245
+ $X2=4.365 $Y2=2.54
r65 7 37 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2 $Y=3.245 $X2=2
+ $Y2=3.33
r66 7 9 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=2 $Y=3.245 $X2=2
+ $Y2=2.8
r67 2 13 300 $w=1.7e-07 $l=5.60647e-07 $layer=licon1_PDIFF $count=2 $X=4.225
+ $Y=2.045 $X2=4.365 $Y2=2.54
r68 1 9 600 $w=1.7e-07 $l=9.19647e-07 $layer=licon1_PDIFF $count=1 $X=1.855
+ $Y=1.95 $X2=2 $Y2=2.8
.ends

.subckt PM_SKY130_FD_SC_LP__A2111O_LP%X 1 2 8 12 14 15
r29 15 18 4.87572 $w=2.58e-07 $l=1.1e-07 $layer=LI1_cond $X=2.64 $Y=2.05
+ $X2=2.53 $Y2=2.05
r30 14 18 5.54059 $w=2.58e-07 $l=1.25e-07 $layer=LI1_cond $X=2.405 $Y=2.05
+ $X2=2.53 $Y2=2.05
r31 9 12 10.9179 $w=3.78e-07 $l=3.6e-07 $layer=LI1_cond $X=2.32 $Y=0.455
+ $X2=2.68 $Y2=0.455
r32 8 14 7.21222 $w=2.6e-07 $l=1.67183e-07 $layer=LI1_cond $X=2.32 $Y=1.92
+ $X2=2.405 $Y2=2.05
r33 7 9 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.32 $Y=0.645 $X2=2.32
+ $Y2=0.455
r34 7 8 83.1818 $w=1.68e-07 $l=1.275e-06 $layer=LI1_cond $X=2.32 $Y=0.645
+ $X2=2.32 $Y2=1.92
r35 2 18 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.39
+ $Y=1.95 $X2=2.53 $Y2=2.095
r36 1 12 182 $w=1.7e-07 $l=2.81425e-07 $layer=licon1_NDIFF $count=1 $X=2.54
+ $Y=0.235 $X2=2.68 $Y2=0.455
.ends

.subckt PM_SKY130_FD_SC_LP__A2111O_LP%A_739_409# 1 2 7 9 11 13 15
r35 13 20 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.97 $Y=2.195 $X2=4.97
+ $Y2=2.11
r36 13 15 24.6204 $w=3.28e-07 $l=7.05e-07 $layer=LI1_cond $X=4.97 $Y=2.195
+ $X2=4.97 $Y2=2.9
r37 12 18 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4 $Y=2.11 $X2=3.835
+ $Y2=2.11
r38 11 20 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.805 $Y=2.11
+ $X2=4.97 $Y2=2.11
r39 11 12 52.5187 $w=1.68e-07 $l=8.05e-07 $layer=LI1_cond $X=4.805 $Y=2.11 $X2=4
+ $Y2=2.11
r40 7 18 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.835 $Y=2.195
+ $X2=3.835 $Y2=2.11
r41 7 9 24.6204 $w=3.28e-07 $l=7.05e-07 $layer=LI1_cond $X=3.835 $Y=2.195
+ $X2=3.835 $Y2=2.9
r42 2 20 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=4.83
+ $Y=2.045 $X2=4.97 $Y2=2.19
r43 2 15 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=4.83
+ $Y=2.045 $X2=4.97 $Y2=2.9
r44 1 18 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=3.695
+ $Y=2.045 $X2=3.835 $Y2=2.19
r45 1 9 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=3.695
+ $Y=2.045 $X2=3.835 $Y2=2.9
.ends

.subckt PM_SKY130_FD_SC_LP__A2111O_LP%VGND 1 2 3 10 12 16 20 23 24 25 34 43 44
+ 50
r72 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r73 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r74 44 51 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=4.08
+ $Y2=0
r75 43 44 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r76 41 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.215 $Y=0 $X2=4.05
+ $Y2=0
r77 41 43 53.8235 $w=1.68e-07 $l=8.25e-07 $layer=LI1_cond $X=4.215 $Y=0 $X2=5.04
+ $Y2=0
r78 40 51 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r79 39 40 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r80 36 39 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=2.16 $Y=0 $X2=3.6
+ $Y2=0
r81 36 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r82 34 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.885 $Y=0 $X2=4.05
+ $Y2=0
r83 34 39 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=3.885 $Y=0 $X2=3.6
+ $Y2=0
r84 33 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r85 32 33 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r86 30 33 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r87 30 48 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r88 29 32 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r89 29 30 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r90 27 47 4.73185 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=0 $X2=0.222
+ $Y2=0
r91 27 29 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.445 $Y=0 $X2=0.72
+ $Y2=0
r92 25 40 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r93 25 37 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=2.16
+ $Y2=0
r94 23 32 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=1.725 $Y=0 $X2=1.68
+ $Y2=0
r95 23 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.725 $Y=0 $X2=1.89
+ $Y2=0
r96 22 36 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=2.055 $Y=0 $X2=2.16
+ $Y2=0
r97 22 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.055 $Y=0 $X2=1.89
+ $Y2=0
r98 18 50 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.05 $Y=0.085
+ $X2=4.05 $Y2=0
r99 18 20 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=4.05 $Y=0.085
+ $X2=4.05 $Y2=0.455
r100 14 24 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.89 $Y=0.085
+ $X2=1.89 $Y2=0
r101 14 16 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=1.89 $Y=0.085
+ $X2=1.89 $Y2=0.43
r102 10 47 3.03433 $w=3.3e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.28 $Y=0.085
+ $X2=0.222 $Y2=0
r103 10 12 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=0.28 $Y=0.085
+ $X2=0.28 $Y2=0.445
r104 3 20 182 $w=1.7e-07 $l=2.29565e-07 $layer=licon1_NDIFF $count=1 $X=3.91
+ $Y=0.285 $X2=4.05 $Y2=0.455
r105 2 16 182 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_NDIFF $count=1 $X=1.75
+ $Y=0.235 $X2=1.89 $Y2=0.43
r106 1 12 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.28 $Y2=0.445
.ends

