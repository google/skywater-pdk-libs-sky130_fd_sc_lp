* File: sky130_fd_sc_lp__sdfrtp_4.spice
* Created: Fri Aug 28 11:28:36 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__sdfrtp_4.pex.spice"
.subckt sky130_fd_sc_lp__sdfrtp_4  VNB VPB SCE D SCD RESET_B CLK VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* CLK	CLK
* RESET_B	RESET_B
* SCD	SCD
* D	D
* SCE	SCE
* VPB	VPB
* VNB	VNB
MM1000 N_VGND_M1000_d N_SCE_M1000_g N_A_27_74#_M1000_s VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.1113 PD=1.37 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1021 noxref_25 N_A_27_74#_M1021_g N_noxref_24_M1021_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1113 PD=0.63 PS=1.37 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.5 A=0.063 P=1.14 MULT=1
MM1023 N_A_372_50#_M1023_d N_D_M1023_g noxref_25 VNB NSHORT L=0.15 W=0.42
+ AD=0.129575 AS=0.0441 PD=1.085 PS=0.63 NRD=34.284 NRS=14.28 M=1 R=2.8
+ SA=75000.6 SB=75001.2 A=0.063 P=1.14 MULT=1
MM1029 noxref_26 N_SCE_M1029_g N_A_372_50#_M1023_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.129575 PD=0.63 PS=1.085 NRD=14.28 NRS=32.856 M=1 R=2.8
+ SA=75000.9 SB=75001 A=0.063 P=1.14 MULT=1
MM1032 N_noxref_24_M1032_d N_SCD_M1032_g noxref_26 VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1001 N_VGND_M1001_d N_RESET_B_M1001_g N_noxref_24_M1032_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75001.7
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1030 N_A_881_463#_M1030_d N_A_975_255#_M1030_g N_A_372_50#_M1030_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.0588 AS=0.126 PD=0.7 PS=1.44 NRD=0 NRS=9.996 M=1 R=2.8
+ SA=75000.2 SB=75004.7 A=0.063 P=1.14 MULT=1
MM1024 A_1107_119# N_A_851_242#_M1024_g N_A_881_463#_M1030_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0672 AS=0.0588 PD=0.74 PS=0.7 NRD=30 NRS=0 M=1 R=2.8 SA=75000.7
+ SB=75004.3 A=0.063 P=1.14 MULT=1
MM1045 A_1201_119# N_A_1047_369#_M1045_g A_1107_119# VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0672 PD=0.63 PS=0.74 NRD=14.28 NRS=30 M=1 R=2.8 SA=75001.1
+ SB=75003.8 A=0.063 P=1.14 MULT=1
MM1036 N_VGND_M1036_d N_RESET_B_M1036_g A_1201_119# VNB NSHORT L=0.15 W=0.42
+ AD=0.112568 AS=0.0441 PD=0.903396 PS=0.63 NRD=27.132 NRS=14.28 M=1 R=2.8
+ SA=75001.5 SB=75003.5 A=0.063 P=1.14 MULT=1
MM1015 N_A_1047_369#_M1015_d N_A_881_463#_M1015_g N_VGND_M1036_d VNB NSHORT
+ L=0.15 W=0.64 AD=0.1552 AS=0.171532 PD=1.125 PS=1.3766 NRD=17.808 NRS=17.808
+ M=1 R=4.26667 SA=75001.4 SB=75002.3 A=0.096 P=1.58 MULT=1
MM1019 N_A_1524_69#_M1019_d N_A_851_242#_M1019_g N_A_1047_369#_M1015_d VNB
+ NSHORT L=0.15 W=0.64 AD=0.226657 AS=0.1552 PD=1.68453 PS=1.125 NRD=0
+ NRS=20.616 M=1 R=4.26667 SA=75002 SB=75001.6 A=0.096 P=1.58 MULT=1
MM1006 A_1705_113# N_A_975_255#_M1006_g N_A_1524_69#_M1019_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.148743 PD=0.63 PS=1.10547 NRD=14.28 NRS=137.136 M=1
+ R=2.8 SA=75003.5 SB=75001.5 A=0.063 P=1.14 MULT=1
MM1039 N_VGND_M1039_d N_A_1747_21#_M1039_g A_1705_113# VNB NSHORT L=0.15 W=0.42
+ AD=0.1035 AS=0.0441 PD=0.925 PS=0.63 NRD=27.132 NRS=14.28 M=1 R=2.8 SA=75003.9
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1026 A_1902_119# N_RESET_B_M1026_g N_VGND_M1039_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1035 PD=0.63 PS=0.925 NRD=14.28 NRS=28.56 M=1 R=2.8 SA=75004.3
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1016 N_A_1747_21#_M1016_d N_A_1524_69#_M1016_g A_1902_119# VNB NSHORT L=0.15
+ W=0.42 AD=0.1113 AS=0.0441 PD=1.37 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8
+ SA=75004.7 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1031 N_VGND_M1031_d N_A_975_255#_M1031_g N_A_851_242#_M1031_s VNB NSHORT
+ L=0.15 W=0.84 AD=0.24485 AS=0.2394 PD=1.495 PS=2.25 NRD=12.132 NRS=0 M=1 R=5.6
+ SA=75000.2 SB=75000.9 A=0.126 P=1.98 MULT=1
MM1011 N_A_975_255#_M1011_d N_CLK_M1011_g N_VGND_M1031_d VNB NSHORT L=0.15
+ W=0.84 AD=0.2394 AS=0.24485 PD=2.25 PS=1.495 NRD=0 NRS=27.132 M=1 R=5.6
+ SA=75000.9 SB=75000.2 A=0.126 P=1.98 MULT=1
MM1041 N_VGND_M1041_d N_A_1524_69#_M1041_g N_A_2555_47#_M1041_s VNB NSHORT
+ L=0.15 W=0.84 AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6
+ SA=75000.2 SB=75001.9 A=0.126 P=1.98 MULT=1
MM1014 N_VGND_M1041_d N_A_2555_47#_M1014_g N_Q_M1014_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75001.5 A=0.126 P=1.98 MULT=1
MM1027 N_VGND_M1027_d N_A_2555_47#_M1027_g N_Q_M1014_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.1
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1040 N_VGND_M1027_d N_A_2555_47#_M1040_g N_Q_M1040_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1344 PD=1.12 PS=1.16 NRD=0 NRS=0 M=1 R=5.6 SA=75001.5
+ SB=75000.7 A=0.126 P=1.98 MULT=1
MM1043 N_VGND_M1043_d N_A_2555_47#_M1043_g N_Q_M1040_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1344 PD=2.21 PS=1.16 NRD=0 NRS=5.712 M=1 R=5.6 SA=75001.9
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1002 N_VPWR_M1002_d N_SCE_M1002_g N_A_27_74#_M1002_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0896 AS=0.1696 PD=0.92 PS=1.81 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75003.8 A=0.096 P=1.58 MULT=1
MM1035 A_407_463# N_SCE_M1035_g N_VPWR_M1002_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0672 AS=0.0896 PD=0.85 PS=0.92 NRD=15.3857 NRS=0 M=1 R=4.26667 SA=75000.6
+ SB=75003.4 A=0.096 P=1.58 MULT=1
MM1038 N_A_372_50#_M1038_d N_D_M1038_g A_407_463# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0896 AS=0.0672 PD=0.92 PS=0.85 NRD=0 NRS=15.3857 M=1 R=4.26667 SA=75001
+ SB=75003.1 A=0.096 P=1.58 MULT=1
MM1020 A_565_463# N_A_27_74#_M1020_g N_A_372_50#_M1038_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1024 AS=0.0896 PD=0.96 PS=0.92 NRD=32.308 NRS=0 M=1 R=4.26667
+ SA=75001.4 SB=75002.6 A=0.096 P=1.58 MULT=1
MM1012 N_VPWR_M1012_d N_SCD_M1012_g A_565_463# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1392 AS=0.1024 PD=1.075 PS=0.96 NRD=26.1616 NRS=32.308 M=1 R=4.26667
+ SA=75001.9 SB=75002.2 A=0.096 P=1.58 MULT=1
MM1033 N_A_372_50#_M1033_d N_RESET_B_M1033_g N_VPWR_M1012_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.130294 AS=0.1392 PD=1.22566 PS=1.075 NRD=0 NRS=21.5321 M=1
+ R=4.26667 SA=75002.5 SB=75001.6 A=0.096 P=1.58 MULT=1
MM1017 N_A_881_463#_M1017_d N_A_851_242#_M1017_g N_A_372_50#_M1033_d VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.0987 AS=0.0855057 PD=0.89 PS=0.80434 NRD=44.5417
+ NRS=45.7237 M=1 R=2.8 SA=75003 SB=75001.8 A=0.063 P=1.14 MULT=1
MM1007 A_1005_463# N_A_975_255#_M1007_g N_A_881_463#_M1017_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0441 AS=0.0987 PD=0.63 PS=0.89 NRD=23.443 NRS=44.5417 M=1 R=2.8
+ SA=75003.6 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1003 N_VPWR_M1003_d N_A_1047_369#_M1003_g A_1005_463# VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0945 AS=0.0441 PD=0.87 PS=0.63 NRD=4.6886 NRS=23.443 M=1 R=2.8
+ SA=75004 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1009 N_A_881_463#_M1009_d N_RESET_B_M1009_g N_VPWR_M1003_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1113 AS=0.0945 PD=1.37 PS=0.87 NRD=0 NRS=75.0373 M=1 R=2.8
+ SA=75004.6 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1022 N_A_1047_369#_M1022_d N_A_881_463#_M1022_g N_VPWR_M1022_s VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.1176 AS=0.3679 PD=1.12 PS=2.7 NRD=0 NRS=28.1316 M=1 R=5.6
+ SA=75000.3 SB=75000.9 A=0.126 P=1.98 MULT=1
MM1010 N_A_1524_69#_M1010_d N_A_975_255#_M1010_g N_A_1047_369#_M1022_d VPB
+ PHIGHVT L=0.15 W=0.84 AD=0.290733 AS=0.1176 PD=2.21333 PS=1.12 NRD=16.4101
+ NRS=0 M=1 R=5.6 SA=75000.8 SB=75000.5 A=0.126 P=1.98 MULT=1
MM1013 A_1662_533# N_A_851_242#_M1013_g N_A_1524_69#_M1010_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0924 AS=0.145367 PD=0.86 PS=1.10667 NRD=77.3816 NRS=136.541 M=1
+ R=2.8 SA=75000.5 SB=75002 A=0.063 P=1.14 MULT=1
MM1028 N_VPWR_M1028_d N_A_1747_21#_M1028_g A_1662_533# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.1197 AS=0.0924 PD=0.99 PS=0.86 NRD=60.9715 NRS=77.3816 M=1 R=2.8
+ SA=75001.1 SB=75001.5 A=0.063 P=1.14 MULT=1
MM1018 N_A_1747_21#_M1018_d N_RESET_B_M1018_g N_VPWR_M1028_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0588 AS=0.1197 PD=0.7 PS=0.99 NRD=0 NRS=75.0373 M=1 R=2.8
+ SA=75001.8 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1042 N_VPWR_M1042_d N_A_1524_69#_M1042_g N_A_1747_21#_M1018_d VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.1596 AS=0.0588 PD=1.6 PS=0.7 NRD=53.9386 NRS=0 M=1 R=2.8
+ SA=75002.2 SB=75000.3 A=0.063 P=1.14 MULT=1
MM1004 N_VPWR_M1004_d N_A_975_255#_M1004_g N_A_851_242#_M1004_s VPB PHIGHVT
+ L=0.15 W=1.26 AD=0.34335 AS=0.3402 PD=1.805 PS=3.06 NRD=27.6194 NRS=0.7683 M=1
+ R=8.4 SA=75000.2 SB=75000.9 A=0.189 P=2.82 MULT=1
MM1037 N_A_975_255#_M1037_d N_CLK_M1037_g N_VPWR_M1004_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.34335 PD=3.05 PS=1.805 NRD=0 NRS=13.8097 M=1 R=8.4
+ SA=75000.9 SB=75000.2 A=0.189 P=2.82 MULT=1
MM1044 N_VPWR_M1044_d N_A_1524_69#_M1044_g N_A_2555_47#_M1044_s VPB PHIGHVT
+ L=0.15 W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.2 SB=75002 A=0.189 P=2.82 MULT=1
MM1005 N_Q_M1005_d N_A_2555_47#_M1005_g N_VPWR_M1044_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75001.5 A=0.189 P=2.82 MULT=1
MM1008 N_Q_M1005_d N_A_2555_47#_M1008_g N_VPWR_M1008_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.2016 PD=1.54 PS=1.58 NRD=0 NRS=3.1126 M=1 R=8.4 SA=75001.1
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1025 N_Q_M1025_d N_A_2555_47#_M1025_g N_VPWR_M1008_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.2016 PD=1.54 PS=1.58 NRD=0 NRS=3.1126 M=1 R=8.4 SA=75001.5
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1034 N_Q_M1025_d N_A_2555_47#_M1034_g N_VPWR_M1034_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75002 SB=75000.2
+ A=0.189 P=2.82 MULT=1
DX46_noxref VNB VPB NWDIODE A=29.3551 P=35.21
c_164 VNB 0 9.46857e-21 $X=0 $Y=0
c_308 VPB 0 1.28163e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_lp__sdfrtp_4.pxi.spice"
*
.ends
*
*
