* NGSPICE file created from sky130_fd_sc_lp__nand4_4.ext - technology: sky130A

.subckt sky130_fd_sc_lp__nand4_4 A B C D VGND VNB VPB VPWR Y
M1000 Y D VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=2.8224e+12p pd=2.464e+07u as=3.906e+12p ps=2.888e+07u
M1001 a_27_65# D VGND VNB nshort w=840000u l=150000u
+  ad=1.2348e+12p pd=1.134e+07u as=4.704e+11p ps=4.48e+06u
M1002 Y C VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 Y A VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_843_67# A Y VNB nshort w=840000u l=150000u
+  ad=1.1844e+12p pd=1.122e+07u as=4.704e+11p ps=4.48e+06u
M1005 a_843_67# A Y VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_27_65# C a_454_65# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=9.408e+11p ps=8.96e+06u
M1007 Y C VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPWR A Y VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_454_65# C a_27_65# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 Y B VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND D a_27_65# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VPWR D Y VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_454_65# B a_843_67# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_843_67# B a_454_65# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 Y B VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VPWR C Y VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VPWR A Y VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_27_65# C a_454_65# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VPWR D Y VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_843_67# B a_454_65# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 Y A VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VPWR B Y VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 VGND D a_27_65# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 Y A a_843_67# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 Y A a_843_67# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_454_65# B a_843_67# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 Y D VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 VPWR C Y VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 VPWR B Y VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 a_454_65# C a_27_65# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_27_65# D VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

