* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__o311a_lp A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
X0 X a_84_115# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X1 VPWR C1 a_84_115# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X2 a_84_115# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X3 VGND A3 a_273_141# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 VPWR A1 a_258_419# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X5 a_273_141# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 a_356_419# A3 a_84_115# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X7 a_563_141# C1 a_84_115# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 a_258_419# A2 a_356_419# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X9 a_114_141# a_84_115# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 a_273_141# B1 a_563_141# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X11 X a_84_115# a_114_141# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 VGND A1 a_273_141# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
