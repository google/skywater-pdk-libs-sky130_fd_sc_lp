* File: sky130_fd_sc_lp__busreceiver_1.pxi.spice
* Created: Wed Sep  2 09:37:54 2020
* 
x_PM_SKY130_FD_SC_LP__BUSRECEIVER_1%A_70_237# N_A_70_237#_M1002_d
+ N_A_70_237#_M1000_d N_A_70_237#_M1001_g N_A_70_237#_M1003_g N_A_70_237#_c_36_n
+ N_A_70_237#_c_37_n N_A_70_237#_c_38_n N_A_70_237#_c_47_p N_A_70_237#_c_79_p
+ N_A_70_237#_c_39_n N_A_70_237#_c_45_n N_A_70_237#_c_46_n N_A_70_237#_c_40_n
+ N_A_70_237#_c_41_n N_A_70_237#_c_42_n
+ PM_SKY130_FD_SC_LP__BUSRECEIVER_1%A_70_237#
x_PM_SKY130_FD_SC_LP__BUSRECEIVER_1%A N_A_c_91_n N_A_M1002_g N_A_M1000_g A
+ N_A_c_94_n PM_SKY130_FD_SC_LP__BUSRECEIVER_1%A
x_PM_SKY130_FD_SC_LP__BUSRECEIVER_1%X N_X_M1001_s N_X_M1003_s X X X X X
+ N_X_c_119_n X X N_X_c_121_n PM_SKY130_FD_SC_LP__BUSRECEIVER_1%X
x_PM_SKY130_FD_SC_LP__BUSRECEIVER_1%VPWR N_VPWR_M1003_d N_VPWR_c_138_n VPWR
+ N_VPWR_c_139_n N_VPWR_c_140_n N_VPWR_c_137_n N_VPWR_c_142_n
+ PM_SKY130_FD_SC_LP__BUSRECEIVER_1%VPWR
x_PM_SKY130_FD_SC_LP__BUSRECEIVER_1%VGND N_VGND_M1001_d N_VGND_c_157_n VGND
+ N_VGND_c_158_n N_VGND_c_159_n N_VGND_c_160_n N_VGND_c_161_n
+ PM_SKY130_FD_SC_LP__BUSRECEIVER_1%VGND
cc_1 VNB N_A_70_237#_M1003_g 0.00742137f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.465
cc_2 VNB N_A_70_237#_c_36_n 0.00100477f $X=-0.19 $Y=-0.245 $X2=0.562 $Y2=1.317
cc_3 VNB N_A_70_237#_c_37_n 0.00262171f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=1.35
cc_4 VNB N_A_70_237#_c_38_n 0.0351264f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=1.35
cc_5 VNB N_A_70_237#_c_39_n 0.00676608f $X=-0.19 $Y=-0.245 $X2=1.025 $Y2=1.69
cc_6 VNB N_A_70_237#_c_40_n 0.00106484f $X=-0.19 $Y=-0.245 $X2=0.562 $Y2=1.185
cc_7 VNB N_A_70_237#_c_41_n 0.0135215f $X=-0.19 $Y=-0.245 $X2=1.18 $Y2=0.855
cc_8 VNB N_A_70_237#_c_42_n 0.0209045f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=1.185
cc_9 VNB N_A_c_91_n 0.0248221f $X=-0.19 $Y=-0.245 $X2=1.04 $Y2=0.655
cc_10 VNB N_A_M1000_g 0.0104722f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB A 0.0100552f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.655
cc_12 VNB N_A_c_94_n 0.0465513f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_X_c_119_n 0.0247509f $X=-0.19 $Y=-0.245 $X2=1.025 $Y2=1.69
cc_14 VNB X 0.0051537f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_X_c_121_n 0.0286293f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_VPWR_c_137_n 0.0641695f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.185
cc_17 VNB N_VGND_c_157_n 0.0152379f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_VGND_c_158_n 0.0152818f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.515
cc_19 VNB N_VGND_c_159_n 0.0194904f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=1.35
cc_20 VNB N_VGND_c_160_n 0.114066f $X=-0.19 $Y=-0.245 $X2=0.515 $Y2=1.35
cc_21 VNB N_VGND_c_161_n 0.00513431f $X=-0.19 $Y=-0.245 $X2=1.025 $Y2=0.935
cc_22 VPB N_A_70_237#_M1003_g 0.0250607f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.465
cc_23 VPB N_A_70_237#_c_39_n 0.00812746f $X=-0.19 $Y=1.655 $X2=1.025 $Y2=1.69
cc_24 VPB N_A_70_237#_c_45_n 0.00135893f $X=-0.19 $Y=1.655 $X2=0.695 $Y2=1.69
cc_25 VPB N_A_70_237#_c_46_n 0.033797f $X=-0.19 $Y=1.655 $X2=1.18 $Y2=1.98
cc_26 VPB N_A_M1000_g 0.0272606f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_27 VPB X 0.0051537f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.465
cc_28 VPB X 0.0413572f $X=-0.19 $Y=1.655 $X2=1.18 $Y2=0.855
cc_29 VPB N_X_c_121_n 0.00967316f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_30 VPB N_VPWR_c_138_n 0.0229311f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_31 VPB N_VPWR_c_139_n 0.0152818f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.465
cc_32 VPB N_VPWR_c_140_n 0.0207592f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=1.02
cc_33 VPB N_VPWR_c_137_n 0.0521093f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=1.185
cc_34 VPB N_VPWR_c_142_n 0.00510842f $X=-0.19 $Y=1.655 $X2=1.025 $Y2=1.69
cc_35 N_A_70_237#_c_47_p N_A_c_91_n 0.0112496f $X=1.025 $Y=0.935 $X2=-0.19
+ $Y2=-0.245
cc_36 N_A_70_237#_c_40_n N_A_c_91_n 0.00298918f $X=0.562 $Y=1.185 $X2=-0.19
+ $Y2=-0.245
cc_37 N_A_70_237#_c_41_n N_A_c_91_n 0.00422733f $X=1.18 $Y=0.855 $X2=-0.19
+ $Y2=-0.245
cc_38 N_A_70_237#_c_42_n N_A_c_91_n 0.017543f $X=0.515 $Y=1.185 $X2=-0.19
+ $Y2=-0.245
cc_39 N_A_70_237#_M1003_g N_A_M1000_g 0.0225139f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_40 N_A_70_237#_c_37_n N_A_M1000_g 0.00298918f $X=0.515 $Y=1.35 $X2=0 $Y2=0
cc_41 N_A_70_237#_c_39_n N_A_M1000_g 0.017511f $X=1.025 $Y=1.69 $X2=0 $Y2=0
cc_42 N_A_70_237#_c_46_n N_A_M1000_g 0.0100119f $X=1.18 $Y=1.98 $X2=0 $Y2=0
cc_43 N_A_70_237#_c_36_n A 0.0122057f $X=0.562 $Y=1.317 $X2=0 $Y2=0
cc_44 N_A_70_237#_c_38_n A 2.57346e-19 $X=0.515 $Y=1.35 $X2=0 $Y2=0
cc_45 N_A_70_237#_c_47_p A 0.00133217f $X=1.025 $Y=0.935 $X2=0 $Y2=0
cc_46 N_A_70_237#_c_39_n A 0.0278482f $X=1.025 $Y=1.69 $X2=0 $Y2=0
cc_47 N_A_70_237#_c_41_n A 0.0221127f $X=1.18 $Y=0.855 $X2=0 $Y2=0
cc_48 N_A_70_237#_c_36_n N_A_c_94_n 0.00298918f $X=0.562 $Y=1.317 $X2=0 $Y2=0
cc_49 N_A_70_237#_c_38_n N_A_c_94_n 0.0211722f $X=0.515 $Y=1.35 $X2=0 $Y2=0
cc_50 N_A_70_237#_c_39_n N_A_c_94_n 0.00756864f $X=1.025 $Y=1.69 $X2=0 $Y2=0
cc_51 N_A_70_237#_c_41_n N_A_c_94_n 0.00661542f $X=1.18 $Y=0.855 $X2=0 $Y2=0
cc_52 N_A_70_237#_M1003_g N_X_c_121_n 0.00784563f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_53 N_A_70_237#_c_36_n N_X_c_121_n 0.0310031f $X=0.562 $Y=1.317 $X2=0 $Y2=0
cc_54 N_A_70_237#_c_38_n N_X_c_121_n 0.0081393f $X=0.515 $Y=1.35 $X2=0 $Y2=0
cc_55 N_A_70_237#_c_45_n N_X_c_121_n 0.0122619f $X=0.695 $Y=1.69 $X2=0 $Y2=0
cc_56 N_A_70_237#_c_40_n N_X_c_121_n 0.00786796f $X=0.562 $Y=1.185 $X2=0 $Y2=0
cc_57 N_A_70_237#_c_42_n N_X_c_121_n 0.00270466f $X=0.515 $Y=1.185 $X2=0 $Y2=0
cc_58 N_A_70_237#_M1003_g N_VPWR_c_138_n 0.0207725f $X=0.475 $Y=2.465 $X2=0
+ $Y2=0
cc_59 N_A_70_237#_c_38_n N_VPWR_c_138_n 4.72889e-19 $X=0.515 $Y=1.35 $X2=0 $Y2=0
cc_60 N_A_70_237#_c_39_n N_VPWR_c_138_n 0.0121673f $X=1.025 $Y=1.69 $X2=0 $Y2=0
cc_61 N_A_70_237#_c_45_n N_VPWR_c_138_n 0.0127495f $X=0.695 $Y=1.69 $X2=0 $Y2=0
cc_62 N_A_70_237#_c_46_n N_VPWR_c_138_n 0.0205413f $X=1.18 $Y=1.98 $X2=0 $Y2=0
cc_63 N_A_70_237#_M1003_g N_VPWR_c_139_n 0.00486043f $X=0.475 $Y=2.465 $X2=0
+ $Y2=0
cc_64 N_A_70_237#_M1003_g N_VPWR_c_137_n 0.00917987f $X=0.475 $Y=2.465 $X2=0
+ $Y2=0
cc_65 N_A_70_237#_c_46_n N_VPWR_c_137_n 0.0124293f $X=1.18 $Y=1.98 $X2=0 $Y2=0
cc_66 N_A_70_237#_c_47_p N_VGND_M1001_d 0.0039601f $X=1.025 $Y=0.935 $X2=-0.19
+ $Y2=-0.245
cc_67 N_A_70_237#_c_79_p N_VGND_M1001_d 9.61307e-19 $X=0.695 $Y=0.935 $X2=-0.19
+ $Y2=-0.245
cc_68 N_A_70_237#_c_40_n N_VGND_M1001_d 6.37289e-19 $X=0.562 $Y=1.185 $X2=-0.19
+ $Y2=-0.245
cc_69 N_A_70_237#_c_38_n N_VGND_c_157_n 4.13391e-19 $X=0.515 $Y=1.35 $X2=0 $Y2=0
cc_70 N_A_70_237#_c_47_p N_VGND_c_157_n 0.010956f $X=1.025 $Y=0.935 $X2=0 $Y2=0
cc_71 N_A_70_237#_c_79_p N_VGND_c_157_n 0.00969245f $X=0.695 $Y=0.935 $X2=0
+ $Y2=0
cc_72 N_A_70_237#_c_42_n N_VGND_c_157_n 0.0139049f $X=0.515 $Y=1.185 $X2=0 $Y2=0
cc_73 N_A_70_237#_c_42_n N_VGND_c_158_n 0.00486043f $X=0.515 $Y=1.185 $X2=0
+ $Y2=0
cc_74 N_A_70_237#_c_41_n N_VGND_c_159_n 0.004748f $X=1.18 $Y=0.855 $X2=0 $Y2=0
cc_75 N_A_70_237#_c_47_p N_VGND_c_160_n 0.00590405f $X=1.025 $Y=0.935 $X2=0
+ $Y2=0
cc_76 N_A_70_237#_c_79_p N_VGND_c_160_n 5.97684e-19 $X=0.695 $Y=0.935 $X2=0
+ $Y2=0
cc_77 N_A_70_237#_c_41_n N_VGND_c_160_n 0.00893333f $X=1.18 $Y=0.855 $X2=0 $Y2=0
cc_78 N_A_70_237#_c_42_n N_VGND_c_160_n 0.00917987f $X=0.515 $Y=1.185 $X2=0
+ $Y2=0
cc_79 N_A_M1000_g N_VPWR_c_138_n 0.00626576f $X=0.965 $Y=2.155 $X2=0 $Y2=0
cc_80 N_A_M1000_g N_VPWR_c_140_n 0.00312414f $X=0.965 $Y=2.155 $X2=0 $Y2=0
cc_81 N_A_M1000_g N_VPWR_c_137_n 0.00410284f $X=0.965 $Y=2.155 $X2=0 $Y2=0
cc_82 N_A_c_91_n N_VGND_c_157_n 0.00382433f $X=0.965 $Y=1.185 $X2=0 $Y2=0
cc_83 N_A_c_91_n N_VGND_c_159_n 0.00391716f $X=0.965 $Y=1.185 $X2=0 $Y2=0
cc_84 N_A_c_91_n N_VGND_c_160_n 0.0046122f $X=0.965 $Y=1.185 $X2=0 $Y2=0
cc_85 X N_VPWR_c_139_n 0.018528f $X=0.24 $Y=2.035 $X2=0 $Y2=0
cc_86 N_X_M1003_s N_VPWR_c_137_n 0.00371702f $X=0.135 $Y=1.835 $X2=0 $Y2=0
cc_87 X N_VPWR_c_137_n 0.0104192f $X=0.24 $Y=2.035 $X2=0 $Y2=0
cc_88 N_X_c_119_n N_VGND_c_158_n 0.018528f $X=0.26 $Y=0.42 $X2=0 $Y2=0
cc_89 N_X_M1001_s N_VGND_c_160_n 0.00371702f $X=0.135 $Y=0.235 $X2=0 $Y2=0
cc_90 N_X_c_119_n N_VGND_c_160_n 0.0104192f $X=0.26 $Y=0.42 $X2=0 $Y2=0
