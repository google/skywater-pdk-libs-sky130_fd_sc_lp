* File: sky130_fd_sc_lp__and3_4.pxi.spice
* Created: Fri Aug 28 10:06:14 2020
* 
x_PM_SKY130_FD_SC_LP__AND3_4%A N_A_M1003_g N_A_M1000_g A A N_A_c_76_n N_A_c_77_n
+ PM_SKY130_FD_SC_LP__AND3_4%A
x_PM_SKY130_FD_SC_LP__AND3_4%B N_B_M1004_g N_B_M1001_g B N_B_c_104_n
+ PM_SKY130_FD_SC_LP__AND3_4%B
x_PM_SKY130_FD_SC_LP__AND3_4%C N_C_M1007_g N_C_M1011_g C N_C_c_133_n
+ PM_SKY130_FD_SC_LP__AND3_4%C
x_PM_SKY130_FD_SC_LP__AND3_4%A_77_47# N_A_77_47#_M1003_s N_A_77_47#_M1000_s
+ N_A_77_47#_M1001_d N_A_77_47#_M1006_g N_A_77_47#_M1002_g N_A_77_47#_M1008_g
+ N_A_77_47#_M1005_g N_A_77_47#_M1009_g N_A_77_47#_M1010_g N_A_77_47#_M1013_g
+ N_A_77_47#_M1012_g N_A_77_47#_c_168_n N_A_77_47#_c_178_n N_A_77_47#_c_179_n
+ N_A_77_47#_c_180_n N_A_77_47#_c_191_n N_A_77_47#_c_169_n N_A_77_47#_c_209_n
+ N_A_77_47#_c_181_n N_A_77_47#_c_170_n N_A_77_47#_c_171_n N_A_77_47#_c_172_n
+ N_A_77_47#_c_183_n N_A_77_47#_c_173_n PM_SKY130_FD_SC_LP__AND3_4%A_77_47#
x_PM_SKY130_FD_SC_LP__AND3_4%VPWR N_VPWR_M1000_d N_VPWR_M1011_d N_VPWR_M1005_s
+ N_VPWR_M1012_s N_VPWR_c_302_n N_VPWR_c_303_n N_VPWR_c_304_n N_VPWR_c_305_n
+ N_VPWR_c_306_n N_VPWR_c_307_n N_VPWR_c_308_n N_VPWR_c_309_n N_VPWR_c_310_n
+ N_VPWR_c_311_n N_VPWR_c_312_n VPWR N_VPWR_c_313_n N_VPWR_c_301_n
+ N_VPWR_c_315_n PM_SKY130_FD_SC_LP__AND3_4%VPWR
x_PM_SKY130_FD_SC_LP__AND3_4%X N_X_M1006_d N_X_M1009_d N_X_M1002_d N_X_M1010_d
+ N_X_c_420_p N_X_c_406_n N_X_c_362_n N_X_c_363_n N_X_c_368_n N_X_c_369_n
+ N_X_c_417_p N_X_c_410_n N_X_c_370_n N_X_c_364_n N_X_c_371_n X X X X X
+ PM_SKY130_FD_SC_LP__AND3_4%X
x_PM_SKY130_FD_SC_LP__AND3_4%VGND N_VGND_M1007_d N_VGND_M1008_s N_VGND_M1013_s
+ N_VGND_c_431_n N_VGND_c_432_n N_VGND_c_433_n N_VGND_c_434_n N_VGND_c_435_n
+ N_VGND_c_436_n N_VGND_c_437_n N_VGND_c_438_n VGND N_VGND_c_439_n
+ N_VGND_c_440_n N_VGND_c_441_n PM_SKY130_FD_SC_LP__AND3_4%VGND
cc_1 VNB N_A_M1000_g 0.0116861f $X=-0.19 $Y=-0.245 $X2=0.725 $Y2=2.465
cc_2 VNB A 0.0370845f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_3 VNB N_A_c_76_n 0.0337675f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.35
cc_4 VNB N_A_c_77_n 0.0216251f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.185
cc_5 VNB N_B_M1004_g 0.0183128f $X=-0.19 $Y=-0.245 $X2=0.725 $Y2=0.655
cc_6 VNB N_B_M1001_g 0.00651524f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB B 0.00331121f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_8 VNB N_B_c_104_n 0.0326994f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.35
cc_9 VNB N_C_M1007_g 0.0203534f $X=-0.19 $Y=-0.245 $X2=0.725 $Y2=0.655
cc_10 VNB N_C_M1011_g 0.00656774f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB C 0.00165097f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_12 VNB N_C_c_133_n 0.032523f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.35
cc_13 VNB N_A_77_47#_M1006_g 0.0238878f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.35
cc_14 VNB N_A_77_47#_M1008_g 0.0222554f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.362
cc_15 VNB N_A_77_47#_M1009_g 0.0222627f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_77_47#_M1013_g 0.0275792f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_77_47#_c_168_n 0.0240525f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_77_47#_c_169_n 0.00753748f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_77_47#_c_170_n 0.0026076f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_77_47#_c_171_n 0.00160869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_77_47#_c_172_n 0.0834119f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_77_47#_c_173_n 0.00189527f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_VPWR_c_301_n 0.183584f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_X_c_362_n 0.00310505f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_X_c_363_n 0.00267635f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_X_c_364_n 0.00147023f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB X 0.037026f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB X 0.0197357f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB X 0.0222686f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_431_n 0.00501393f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.35
cc_31 VNB N_VGND_c_432_n 3.21684e-19 $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.515
cc_32 VNB N_VGND_c_433_n 0.0129398f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_434_n 0.00250565f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_435_n 0.0544595f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_436_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_437_n 0.0163732f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_438_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_439_n 0.0162485f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_440_n 0.247225f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_441_n 0.00426875f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VPB N_A_M1000_g 0.0260004f $X=-0.19 $Y=1.655 $X2=0.725 $Y2=2.465
cc_42 VPB N_B_M1001_g 0.0199624f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_43 VPB N_C_M1011_g 0.0201898f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_44 VPB N_A_77_47#_M1002_g 0.0197001f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.515
cc_45 VPB N_A_77_47#_M1005_g 0.018348f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_46 VPB N_A_77_47#_M1010_g 0.0183546f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_47 VPB N_A_77_47#_M1012_g 0.0223492f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_48 VPB N_A_77_47#_c_178_n 0.0437226f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_49 VPB N_A_77_47#_c_179_n 0.00462069f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_50 VPB N_A_77_47#_c_180_n 0.0116387f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_51 VPB N_A_77_47#_c_181_n 0.00291273f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_52 VPB N_A_77_47#_c_172_n 0.0150337f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_53 VPB N_A_77_47#_c_183_n 0.00339591f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_54 VPB N_A_77_47#_c_173_n 8.15258e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_55 VPB N_VPWR_c_302_n 0.00502942f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.185
cc_56 VPB N_VPWR_c_303_n 0.00435859f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_57 VPB N_VPWR_c_304_n 3.18512e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_58 VPB N_VPWR_c_305_n 0.0129398f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_59 VPB N_VPWR_c_306_n 0.0415892f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_60 VPB N_VPWR_c_307_n 0.025557f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_61 VPB N_VPWR_c_308_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_62 VPB N_VPWR_c_309_n 0.0172488f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_63 VPB N_VPWR_c_310_n 0.00631825f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_64 VPB N_VPWR_c_311_n 0.0157368f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_312_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_313_n 0.0164632f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_67 VPB N_VPWR_c_301_n 0.069365f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_315_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_69 VPB N_X_c_368_n 0.00304538f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_70 VPB N_X_c_369_n 0.00202885f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_71 VPB N_X_c_370_n 0.027677f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_72 VPB N_X_c_371_n 0.00144145f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_73 VPB X 0.00557628f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_74 N_A_c_77_n N_B_M1004_g 0.0454996f $X=0.635 $Y=1.185 $X2=0 $Y2=0
cc_75 N_A_M1000_g N_B_M1001_g 0.0211543f $X=0.725 $Y=2.465 $X2=0 $Y2=0
cc_76 A B 0.0222735f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_77 N_A_c_76_n B 5.49944e-19 $X=0.635 $Y=1.35 $X2=0 $Y2=0
cc_78 A N_B_c_104_n 0.00189238f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_79 N_A_c_76_n N_B_c_104_n 0.0454996f $X=0.635 $Y=1.35 $X2=0 $Y2=0
cc_80 N_A_c_77_n N_A_77_47#_c_168_n 0.013551f $X=0.635 $Y=1.185 $X2=0 $Y2=0
cc_81 N_A_M1000_g N_A_77_47#_c_179_n 0.0175125f $X=0.725 $Y=2.465 $X2=0 $Y2=0
cc_82 A N_A_77_47#_c_179_n 0.012435f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_83 N_A_c_76_n N_A_77_47#_c_179_n 7.74134e-19 $X=0.635 $Y=1.35 $X2=0 $Y2=0
cc_84 A N_A_77_47#_c_180_n 0.0209519f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_85 N_A_c_76_n N_A_77_47#_c_180_n 0.00333538f $X=0.635 $Y=1.35 $X2=0 $Y2=0
cc_86 A N_A_77_47#_c_191_n 0.00904214f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_87 N_A_c_77_n N_A_77_47#_c_191_n 0.0106483f $X=0.635 $Y=1.185 $X2=0 $Y2=0
cc_88 A N_A_77_47#_c_169_n 0.0250124f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_89 N_A_c_76_n N_A_77_47#_c_169_n 0.00413884f $X=0.635 $Y=1.35 $X2=0 $Y2=0
cc_90 N_A_c_77_n N_A_77_47#_c_169_n 7.32094e-19 $X=0.635 $Y=1.185 $X2=0 $Y2=0
cc_91 N_A_M1000_g N_VPWR_c_302_n 0.00332716f $X=0.725 $Y=2.465 $X2=0 $Y2=0
cc_92 N_A_M1000_g N_VPWR_c_307_n 0.00585385f $X=0.725 $Y=2.465 $X2=0 $Y2=0
cc_93 N_A_M1000_g N_VPWR_c_301_n 0.0118409f $X=0.725 $Y=2.465 $X2=0 $Y2=0
cc_94 N_A_c_77_n N_VGND_c_435_n 0.0054895f $X=0.635 $Y=1.185 $X2=0 $Y2=0
cc_95 N_A_c_77_n N_VGND_c_440_n 0.0109514f $X=0.635 $Y=1.185 $X2=0 $Y2=0
cc_96 N_B_M1004_g N_C_M1007_g 0.0375114f $X=1.085 $Y=0.655 $X2=0 $Y2=0
cc_97 N_B_M1001_g N_C_M1011_g 0.0262423f $X=1.235 $Y=2.465 $X2=0 $Y2=0
cc_98 B C 0.0173425f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_99 N_B_c_104_n C 0.00107695f $X=1.175 $Y=1.375 $X2=0 $Y2=0
cc_100 B N_C_c_133_n 0.00118972f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_101 N_B_c_104_n N_C_c_133_n 0.0202736f $X=1.175 $Y=1.375 $X2=0 $Y2=0
cc_102 N_B_M1004_g N_A_77_47#_c_168_n 0.00308147f $X=1.085 $Y=0.655 $X2=0 $Y2=0
cc_103 N_B_M1001_g N_A_77_47#_c_179_n 0.0163027f $X=1.235 $Y=2.465 $X2=0 $Y2=0
cc_104 B N_A_77_47#_c_179_n 0.024644f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_105 N_B_c_104_n N_A_77_47#_c_179_n 0.00126238f $X=1.175 $Y=1.375 $X2=0 $Y2=0
cc_106 N_B_M1004_g N_A_77_47#_c_191_n 0.0150723f $X=1.085 $Y=0.655 $X2=0 $Y2=0
cc_107 B N_A_77_47#_c_191_n 0.0219008f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_108 N_B_c_104_n N_A_77_47#_c_191_n 0.00112336f $X=1.175 $Y=1.375 $X2=0 $Y2=0
cc_109 N_B_M1001_g N_VPWR_c_302_n 0.0018561f $X=1.235 $Y=2.465 $X2=0 $Y2=0
cc_110 N_B_M1001_g N_VPWR_c_309_n 0.00585385f $X=1.235 $Y=2.465 $X2=0 $Y2=0
cc_111 N_B_M1001_g N_VPWR_c_301_n 0.0107676f $X=1.235 $Y=2.465 $X2=0 $Y2=0
cc_112 N_B_M1004_g N_VGND_c_435_n 0.00585385f $X=1.085 $Y=0.655 $X2=0 $Y2=0
cc_113 N_B_M1004_g N_VGND_c_440_n 0.011101f $X=1.085 $Y=0.655 $X2=0 $Y2=0
cc_114 N_C_M1007_g N_A_77_47#_M1006_g 0.0261484f $X=1.625 $Y=0.655 $X2=0 $Y2=0
cc_115 C N_A_77_47#_M1006_g 2.91659e-19 $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_116 N_C_c_133_n N_A_77_47#_M1006_g 0.0167507f $X=1.715 $Y=1.375 $X2=0 $Y2=0
cc_117 N_C_M1007_g N_A_77_47#_c_191_n 0.0168063f $X=1.625 $Y=0.655 $X2=0 $Y2=0
cc_118 C N_A_77_47#_c_191_n 0.0134757f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_119 N_C_c_133_n N_A_77_47#_c_191_n 0.00258174f $X=1.715 $Y=1.375 $X2=0 $Y2=0
cc_120 N_C_M1011_g N_A_77_47#_c_209_n 0.012727f $X=1.665 $Y=2.465 $X2=0 $Y2=0
cc_121 N_C_M1011_g N_A_77_47#_c_181_n 0.0125569f $X=1.665 $Y=2.465 $X2=0 $Y2=0
cc_122 C N_A_77_47#_c_181_n 0.0155486f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_123 N_C_c_133_n N_A_77_47#_c_181_n 0.0024279f $X=1.715 $Y=1.375 $X2=0 $Y2=0
cc_124 N_C_M1007_g N_A_77_47#_c_170_n 0.00326623f $X=1.625 $Y=0.655 $X2=0 $Y2=0
cc_125 C N_A_77_47#_c_170_n 0.0239745f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_126 N_C_c_133_n N_A_77_47#_c_170_n 0.00217772f $X=1.715 $Y=1.375 $X2=0 $Y2=0
cc_127 N_C_M1011_g N_A_77_47#_c_172_n 0.0164882f $X=1.665 $Y=2.465 $X2=0 $Y2=0
cc_128 N_C_M1011_g N_A_77_47#_c_183_n 0.00256592f $X=1.665 $Y=2.465 $X2=0 $Y2=0
cc_129 N_C_c_133_n N_A_77_47#_c_183_n 0.00136482f $X=1.715 $Y=1.375 $X2=0 $Y2=0
cc_130 N_C_M1011_g N_A_77_47#_c_173_n 0.0035765f $X=1.665 $Y=2.465 $X2=0 $Y2=0
cc_131 N_C_M1011_g N_VPWR_c_303_n 0.00199498f $X=1.665 $Y=2.465 $X2=0 $Y2=0
cc_132 N_C_M1011_g N_VPWR_c_309_n 0.00579312f $X=1.665 $Y=2.465 $X2=0 $Y2=0
cc_133 N_C_M1011_g N_VPWR_c_301_n 0.0107078f $X=1.665 $Y=2.465 $X2=0 $Y2=0
cc_134 N_C_M1007_g N_VGND_c_431_n 0.00601737f $X=1.625 $Y=0.655 $X2=0 $Y2=0
cc_135 N_C_M1007_g N_VGND_c_435_n 0.00585385f $X=1.625 $Y=0.655 $X2=0 $Y2=0
cc_136 N_C_M1007_g N_VGND_c_440_n 0.011482f $X=1.625 $Y=0.655 $X2=0 $Y2=0
cc_137 N_A_77_47#_c_179_n N_VPWR_M1000_d 0.00269806f $X=1.35 $Y=1.817 $X2=-0.19
+ $Y2=-0.245
cc_138 N_A_77_47#_c_181_n N_VPWR_M1011_d 0.00211177f $X=1.98 $Y=1.795 $X2=0
+ $Y2=0
cc_139 N_A_77_47#_c_173_n N_VPWR_M1011_d 0.00107162f $X=2.065 $Y=1.5 $X2=0 $Y2=0
cc_140 N_A_77_47#_c_179_n N_VPWR_c_302_n 0.0194846f $X=1.35 $Y=1.817 $X2=0 $Y2=0
cc_141 N_A_77_47#_M1002_g N_VPWR_c_303_n 0.0019225f $X=2.2 $Y=2.465 $X2=0 $Y2=0
cc_142 N_A_77_47#_c_181_n N_VPWR_c_303_n 0.0148886f $X=1.98 $Y=1.795 $X2=0 $Y2=0
cc_143 N_A_77_47#_c_173_n N_VPWR_c_303_n 0.00784407f $X=2.065 $Y=1.5 $X2=0 $Y2=0
cc_144 N_A_77_47#_M1002_g N_VPWR_c_304_n 7.49374e-19 $X=2.2 $Y=2.465 $X2=0 $Y2=0
cc_145 N_A_77_47#_M1005_g N_VPWR_c_304_n 0.0144646f $X=2.63 $Y=2.465 $X2=0 $Y2=0
cc_146 N_A_77_47#_M1010_g N_VPWR_c_304_n 0.0143393f $X=3.06 $Y=2.465 $X2=0 $Y2=0
cc_147 N_A_77_47#_M1012_g N_VPWR_c_304_n 7.27171e-19 $X=3.49 $Y=2.465 $X2=0
+ $Y2=0
cc_148 N_A_77_47#_M1010_g N_VPWR_c_305_n 0.00486043f $X=3.06 $Y=2.465 $X2=0
+ $Y2=0
cc_149 N_A_77_47#_M1012_g N_VPWR_c_305_n 0.00486043f $X=3.49 $Y=2.465 $X2=0
+ $Y2=0
cc_150 N_A_77_47#_M1010_g N_VPWR_c_306_n 7.27171e-19 $X=3.06 $Y=2.465 $X2=0
+ $Y2=0
cc_151 N_A_77_47#_M1012_g N_VPWR_c_306_n 0.0153838f $X=3.49 $Y=2.465 $X2=0 $Y2=0
cc_152 N_A_77_47#_c_178_n N_VPWR_c_307_n 0.0181659f $X=0.51 $Y=1.98 $X2=0 $Y2=0
cc_153 N_A_77_47#_c_209_n N_VPWR_c_309_n 0.014502f $X=1.45 $Y=1.98 $X2=0 $Y2=0
cc_154 N_A_77_47#_M1002_g N_VPWR_c_311_n 0.00585385f $X=2.2 $Y=2.465 $X2=0 $Y2=0
cc_155 N_A_77_47#_M1005_g N_VPWR_c_311_n 0.00486043f $X=2.63 $Y=2.465 $X2=0
+ $Y2=0
cc_156 N_A_77_47#_M1000_s N_VPWR_c_301_n 0.00336915f $X=0.385 $Y=1.835 $X2=0
+ $Y2=0
cc_157 N_A_77_47#_M1001_d N_VPWR_c_301_n 0.00362709f $X=1.31 $Y=1.835 $X2=0
+ $Y2=0
cc_158 N_A_77_47#_M1002_g N_VPWR_c_301_n 0.0108346f $X=2.2 $Y=2.465 $X2=0 $Y2=0
cc_159 N_A_77_47#_M1005_g N_VPWR_c_301_n 0.00824727f $X=2.63 $Y=2.465 $X2=0
+ $Y2=0
cc_160 N_A_77_47#_M1010_g N_VPWR_c_301_n 0.00824727f $X=3.06 $Y=2.465 $X2=0
+ $Y2=0
cc_161 N_A_77_47#_M1012_g N_VPWR_c_301_n 0.00824727f $X=3.49 $Y=2.465 $X2=0
+ $Y2=0
cc_162 N_A_77_47#_c_178_n N_VPWR_c_301_n 0.0104192f $X=0.51 $Y=1.98 $X2=0 $Y2=0
cc_163 N_A_77_47#_c_209_n N_VPWR_c_301_n 0.0093558f $X=1.45 $Y=1.98 $X2=0 $Y2=0
cc_164 N_A_77_47#_M1008_g N_X_c_362_n 0.0138138f $X=2.63 $Y=0.655 $X2=0 $Y2=0
cc_165 N_A_77_47#_M1009_g N_X_c_362_n 0.01419f $X=3.06 $Y=0.655 $X2=0 $Y2=0
cc_166 N_A_77_47#_c_171_n N_X_c_362_n 0.0447065f $X=3.65 $Y=1.5 $X2=0 $Y2=0
cc_167 N_A_77_47#_c_172_n N_X_c_362_n 0.00244902f $X=3.65 $Y=1.5 $X2=0 $Y2=0
cc_168 N_A_77_47#_M1006_g N_X_c_363_n 0.00131587f $X=2.2 $Y=0.655 $X2=0 $Y2=0
cc_169 N_A_77_47#_c_170_n N_X_c_363_n 0.0132012f $X=2.065 $Y=1.415 $X2=0 $Y2=0
cc_170 N_A_77_47#_c_171_n N_X_c_363_n 0.014687f $X=3.65 $Y=1.5 $X2=0 $Y2=0
cc_171 N_A_77_47#_c_172_n N_X_c_363_n 0.00255521f $X=3.65 $Y=1.5 $X2=0 $Y2=0
cc_172 N_A_77_47#_M1005_g N_X_c_368_n 0.0130035f $X=2.63 $Y=2.465 $X2=0 $Y2=0
cc_173 N_A_77_47#_M1010_g N_X_c_368_n 0.0131657f $X=3.06 $Y=2.465 $X2=0 $Y2=0
cc_174 N_A_77_47#_c_171_n N_X_c_368_n 0.0467265f $X=3.65 $Y=1.5 $X2=0 $Y2=0
cc_175 N_A_77_47#_c_172_n N_X_c_368_n 0.00246472f $X=3.65 $Y=1.5 $X2=0 $Y2=0
cc_176 N_A_77_47#_M1002_g N_X_c_369_n 6.55961e-19 $X=2.2 $Y=2.465 $X2=0 $Y2=0
cc_177 N_A_77_47#_c_171_n N_X_c_369_n 0.0153308f $X=3.65 $Y=1.5 $X2=0 $Y2=0
cc_178 N_A_77_47#_c_172_n N_X_c_369_n 0.00256759f $X=3.65 $Y=1.5 $X2=0 $Y2=0
cc_179 N_A_77_47#_c_173_n N_X_c_369_n 0.00793934f $X=2.065 $Y=1.5 $X2=0 $Y2=0
cc_180 N_A_77_47#_M1012_g N_X_c_370_n 0.0151718f $X=3.49 $Y=2.465 $X2=0 $Y2=0
cc_181 N_A_77_47#_c_171_n N_X_c_370_n 0.0312279f $X=3.65 $Y=1.5 $X2=0 $Y2=0
cc_182 N_A_77_47#_c_172_n N_X_c_370_n 0.0061618f $X=3.65 $Y=1.5 $X2=0 $Y2=0
cc_183 N_A_77_47#_c_171_n N_X_c_364_n 0.014687f $X=3.65 $Y=1.5 $X2=0 $Y2=0
cc_184 N_A_77_47#_c_172_n N_X_c_364_n 0.00255521f $X=3.65 $Y=1.5 $X2=0 $Y2=0
cc_185 N_A_77_47#_c_171_n N_X_c_371_n 0.0153308f $X=3.65 $Y=1.5 $X2=0 $Y2=0
cc_186 N_A_77_47#_c_172_n N_X_c_371_n 0.00256759f $X=3.65 $Y=1.5 $X2=0 $Y2=0
cc_187 N_A_77_47#_M1013_g X 0.00257405f $X=3.49 $Y=0.655 $X2=0 $Y2=0
cc_188 N_A_77_47#_M1013_g X 0.0161962f $X=3.49 $Y=0.655 $X2=0 $Y2=0
cc_189 N_A_77_47#_c_171_n X 0.0298871f $X=3.65 $Y=1.5 $X2=0 $Y2=0
cc_190 N_A_77_47#_c_172_n X 0.00612256f $X=3.65 $Y=1.5 $X2=0 $Y2=0
cc_191 N_A_77_47#_M1013_g X 0.00266999f $X=3.49 $Y=0.655 $X2=0 $Y2=0
cc_192 N_A_77_47#_M1012_g X 0.00240029f $X=3.49 $Y=2.465 $X2=0 $Y2=0
cc_193 N_A_77_47#_c_171_n X 0.013141f $X=3.65 $Y=1.5 $X2=0 $Y2=0
cc_194 N_A_77_47#_c_172_n X 0.00803399f $X=3.65 $Y=1.5 $X2=0 $Y2=0
cc_195 N_A_77_47#_c_191_n A_160_47# 0.00558659f $X=1.98 $Y=0.955 $X2=-0.19
+ $Y2=-0.245
cc_196 N_A_77_47#_c_191_n A_232_47# 0.014897f $X=1.98 $Y=0.955 $X2=-0.19
+ $Y2=-0.245
cc_197 N_A_77_47#_c_191_n N_VGND_M1007_d 0.00731953f $X=1.98 $Y=0.955 $X2=-0.19
+ $Y2=-0.245
cc_198 N_A_77_47#_c_170_n N_VGND_M1007_d 4.29653e-19 $X=2.065 $Y=1.415 $X2=-0.19
+ $Y2=-0.245
cc_199 N_A_77_47#_M1006_g N_VGND_c_431_n 0.0045244f $X=2.2 $Y=0.655 $X2=0 $Y2=0
cc_200 N_A_77_47#_c_191_n N_VGND_c_431_n 0.0260407f $X=1.98 $Y=0.955 $X2=0 $Y2=0
cc_201 N_A_77_47#_M1006_g N_VGND_c_432_n 6.61067e-19 $X=2.2 $Y=0.655 $X2=0 $Y2=0
cc_202 N_A_77_47#_M1008_g N_VGND_c_432_n 0.0111931f $X=2.63 $Y=0.655 $X2=0 $Y2=0
cc_203 N_A_77_47#_M1009_g N_VGND_c_432_n 0.0110241f $X=3.06 $Y=0.655 $X2=0 $Y2=0
cc_204 N_A_77_47#_M1013_g N_VGND_c_432_n 6.30983e-19 $X=3.49 $Y=0.655 $X2=0
+ $Y2=0
cc_205 N_A_77_47#_M1009_g N_VGND_c_433_n 0.00486043f $X=3.06 $Y=0.655 $X2=0
+ $Y2=0
cc_206 N_A_77_47#_M1013_g N_VGND_c_433_n 0.00486043f $X=3.49 $Y=0.655 $X2=0
+ $Y2=0
cc_207 N_A_77_47#_M1009_g N_VGND_c_434_n 6.28331e-19 $X=3.06 $Y=0.655 $X2=0
+ $Y2=0
cc_208 N_A_77_47#_M1013_g N_VGND_c_434_n 0.0117528f $X=3.49 $Y=0.655 $X2=0 $Y2=0
cc_209 N_A_77_47#_c_168_n N_VGND_c_435_n 0.0210467f $X=0.51 $Y=0.38 $X2=0 $Y2=0
cc_210 N_A_77_47#_M1006_g N_VGND_c_437_n 0.00585385f $X=2.2 $Y=0.655 $X2=0 $Y2=0
cc_211 N_A_77_47#_M1008_g N_VGND_c_437_n 0.00486043f $X=2.63 $Y=0.655 $X2=0
+ $Y2=0
cc_212 N_A_77_47#_M1003_s N_VGND_c_440_n 0.00215158f $X=0.385 $Y=0.235 $X2=0
+ $Y2=0
cc_213 N_A_77_47#_M1006_g N_VGND_c_440_n 0.0110998f $X=2.2 $Y=0.655 $X2=0 $Y2=0
cc_214 N_A_77_47#_M1008_g N_VGND_c_440_n 0.00824727f $X=2.63 $Y=0.655 $X2=0
+ $Y2=0
cc_215 N_A_77_47#_M1009_g N_VGND_c_440_n 0.00824727f $X=3.06 $Y=0.655 $X2=0
+ $Y2=0
cc_216 N_A_77_47#_M1013_g N_VGND_c_440_n 0.00824727f $X=3.49 $Y=0.655 $X2=0
+ $Y2=0
cc_217 N_A_77_47#_c_168_n N_VGND_c_440_n 0.0125689f $X=0.51 $Y=0.38 $X2=0 $Y2=0
cc_218 N_VPWR_c_301_n N_X_M1002_d 0.00536646f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_219 N_VPWR_c_301_n N_X_M1010_d 0.00536646f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_220 N_VPWR_c_311_n N_X_c_406_n 0.0124525f $X=2.68 $Y=3.33 $X2=0 $Y2=0
cc_221 N_VPWR_c_301_n N_X_c_406_n 0.00730901f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_222 N_VPWR_M1005_s N_X_c_368_n 0.00176461f $X=2.705 $Y=1.835 $X2=0 $Y2=0
cc_223 N_VPWR_c_304_n N_X_c_368_n 0.0170777f $X=2.845 $Y=2.18 $X2=0 $Y2=0
cc_224 N_VPWR_c_305_n N_X_c_410_n 0.0124525f $X=3.54 $Y=3.33 $X2=0 $Y2=0
cc_225 N_VPWR_c_301_n N_X_c_410_n 0.00730901f $X=4.08 $Y=3.33 $X2=0 $Y2=0
cc_226 N_VPWR_M1012_s N_X_c_370_n 0.00262981f $X=3.565 $Y=1.835 $X2=0 $Y2=0
cc_227 N_VPWR_c_306_n N_X_c_370_n 0.0220026f $X=3.705 $Y=2.18 $X2=0 $Y2=0
cc_228 N_X_c_362_n N_VGND_M1008_s 0.00176461f $X=3.18 $Y=1.15 $X2=0 $Y2=0
cc_229 X N_VGND_M1013_s 0.00241858f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_230 N_X_c_362_n N_VGND_c_432_n 0.0170777f $X=3.18 $Y=1.15 $X2=0 $Y2=0
cc_231 N_X_c_417_p N_VGND_c_433_n 0.0124525f $X=3.275 $Y=0.42 $X2=0 $Y2=0
cc_232 X N_VGND_c_434_n 0.0397208f $X=3.995 $Y=0.47 $X2=0 $Y2=0
cc_233 X N_VGND_c_434_n 0.0182205f $X=3.995 $Y=1.21 $X2=0 $Y2=0
cc_234 N_X_c_420_p N_VGND_c_437_n 0.0124525f $X=2.415 $Y=0.42 $X2=0 $Y2=0
cc_235 X N_VGND_c_439_n 0.00876216f $X=3.995 $Y=0.47 $X2=0 $Y2=0
cc_236 N_X_M1006_d N_VGND_c_440_n 0.00536646f $X=2.275 $Y=0.235 $X2=0 $Y2=0
cc_237 N_X_M1009_d N_VGND_c_440_n 0.00536646f $X=3.135 $Y=0.235 $X2=0 $Y2=0
cc_238 N_X_c_420_p N_VGND_c_440_n 0.00730901f $X=2.415 $Y=0.42 $X2=0 $Y2=0
cc_239 N_X_c_417_p N_VGND_c_440_n 0.00730901f $X=3.275 $Y=0.42 $X2=0 $Y2=0
cc_240 X N_VGND_c_440_n 0.00821462f $X=3.995 $Y=0.47 $X2=0 $Y2=0
cc_241 A_160_47# N_VGND_c_440_n 0.00899413f $X=0.8 $Y=0.235 $X2=0.51 $Y2=0.38
cc_242 A_232_47# N_VGND_c_440_n 0.0167135f $X=1.16 $Y=0.235 $X2=0.51 $Y2=0.38
