* File: sky130_fd_sc_lp__nand2b_4.spice
* Created: Wed Sep  2 10:03:40 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__nand2b_4.pex.spice"
.subckt sky130_fd_sc_lp__nand2b_4  VNB VPB A_N B VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B	B
* A_N	A_N
* VPB	VPB
* VNB	VNB
MM1011 N_VGND_M1011_d N_A_N_M1011_g N_A_27_51#_M1011_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.2226 PD=2.21 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1000 N_Y_M1000_d N_A_27_51#_M1000_g N_A_217_65#_M1000_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75003.3 A=0.126 P=1.98 MULT=1
MM1001 N_Y_M1000_d N_A_27_51#_M1001_g N_A_217_65#_M1001_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.147 PD=1.12 PS=1.19 NRD=0 NRS=9.996 M=1 R=5.6 SA=75000.6
+ SB=75002.9 A=0.126 P=1.98 MULT=1
MM1008 N_Y_M1008_d N_A_27_51#_M1008_g N_A_217_65#_M1001_s VNB NSHORT L=0.15
+ W=0.84 AD=0.147 AS=0.147 PD=1.19 PS=1.19 NRD=9.996 NRS=0 M=1 R=5.6 SA=75001.1
+ SB=75002.4 A=0.126 P=1.98 MULT=1
MM1015 N_Y_M1008_d N_A_27_51#_M1015_g N_A_217_65#_M1015_s VNB NSHORT L=0.15
+ W=0.84 AD=0.147 AS=0.1176 PD=1.19 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.6
+ SB=75001.9 A=0.126 P=1.98 MULT=1
MM1003 N_VGND_M1003_d N_B_M1003_g N_A_217_65#_M1015_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002.1
+ SB=75001.5 A=0.126 P=1.98 MULT=1
MM1005 N_VGND_M1003_d N_B_M1005_g N_A_217_65#_M1005_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002.5
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1010 N_VGND_M1010_d N_B_M1010_g N_A_217_65#_M1005_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002.9
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1014 N_VGND_M1010_d N_B_M1014_g N_A_217_65#_M1014_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75003.3
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1016 N_VPWR_M1016_d N_A_N_M1016_g N_A_27_51#_M1016_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.4536 AS=0.3339 PD=1.98 PS=3.05 NRD=34.3962 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75004.4 A=0.189 P=2.82 MULT=1
MM1002 N_VPWR_M1016_d N_A_27_51#_M1002_g N_Y_M1002_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.4536 AS=0.1764 PD=1.98 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75003.5 A=0.189 P=2.82 MULT=1
MM1006 N_VPWR_M1006_d N_A_27_51#_M1006_g N_Y_M1002_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.2268 AS=0.1764 PD=1.62 PS=1.54 NRD=6.2449 NRS=0 M=1 R=8.4 SA=75001.5
+ SB=75003.1 A=0.189 P=2.82 MULT=1
MM1007 N_VPWR_M1006_d N_A_27_51#_M1007_g N_Y_M1007_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.2268 AS=0.1764 PD=1.62 PS=1.54 NRD=6.2449 NRS=0 M=1 R=8.4 SA=75002
+ SB=75002.5 A=0.189 P=2.82 MULT=1
MM1012 N_VPWR_M1012_d N_A_27_51#_M1012_g N_Y_M1007_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.2646 AS=0.1764 PD=1.68 PS=1.54 NRD=10.9335 NRS=0 M=1 R=8.4 SA=75002.4
+ SB=75002.1 A=0.189 P=2.82 MULT=1
MM1004 N_VPWR_M1012_d N_B_M1004_g N_Y_M1004_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.2646 AS=0.2142 PD=1.68 PS=1.6 NRD=10.9335 NRS=3.9006 M=1 R=8.4 SA=75003
+ SB=75001.5 A=0.189 P=2.82 MULT=1
MM1009 N_VPWR_M1009_d N_B_M1009_g N_Y_M1004_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.2142 PD=1.54 PS=1.6 NRD=0 NRS=5.4569 M=1 R=8.4 SA=75003.5
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1013 N_VPWR_M1009_d N_B_M1013_g N_Y_M1013_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75003.9
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1017 N_VPWR_M1017_d N_B_M1017_g N_Y_M1013_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75004.4
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX18_noxref VNB VPB NWDIODE A=10.5559 P=15.05
*
.include "sky130_fd_sc_lp__nand2b_4.pxi.spice"
*
.ends
*
*
