* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__sdlclkp_1 CLK GATE SCE VGND VNB VPB VPWR GCLK
X0 a_1231_367# a_737_329# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X1 a_254_357# CLK VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 VGND CLK a_1194_52# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 a_721_133# a_737_329# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 a_110_468# GATE a_154_69# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X5 VPWR a_1231_367# GCLK VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X6 VGND a_254_357# a_334_69# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 a_254_357# CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X8 VPWR SCE a_110_468# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X9 a_736_463# a_737_329# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X10 a_623_133# a_334_69# a_721_133# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X11 VPWR a_623_133# a_737_329# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X12 VPWR CLK a_1231_367# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X13 VGND a_623_133# a_737_329# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X14 VGND SCE a_154_69# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X15 a_154_69# GATE VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X16 a_1194_52# a_737_329# a_1231_367# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X17 a_154_69# a_254_357# a_623_133# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X18 VPWR a_254_357# a_334_69# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X19 a_623_133# a_254_357# a_736_463# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X20 VGND a_1231_367# GCLK VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X21 a_154_69# a_334_69# a_623_133# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
.ends
