* File: sky130_fd_sc_lp__dfbbn_2.pxi.spice
* Created: Fri Aug 28 10:21:17 2020
* 
x_PM_SKY130_FD_SC_LP__DFBBN_2%CLK_N N_CLK_N_c_294_n N_CLK_N_M1025_g
+ N_CLK_N_c_301_n N_CLK_N_M1034_g N_CLK_N_c_296_n N_CLK_N_c_297_n
+ N_CLK_N_c_302_n CLK_N CLK_N CLK_N N_CLK_N_c_298_n N_CLK_N_c_299_n
+ PM_SKY130_FD_SC_LP__DFBBN_2%CLK_N
x_PM_SKY130_FD_SC_LP__DFBBN_2%D N_D_c_328_n N_D_c_329_n N_D_c_334_n N_D_M1042_g
+ N_D_c_330_n N_D_M1012_g N_D_c_335_n D N_D_c_331_n N_D_c_332_n
+ PM_SKY130_FD_SC_LP__DFBBN_2%D
x_PM_SKY130_FD_SC_LP__DFBBN_2%A_113_57# N_A_113_57#_M1025_d N_A_113_57#_M1034_d
+ N_A_113_57#_c_383_n N_A_113_57#_c_384_n N_A_113_57#_c_406_n
+ N_A_113_57#_c_407_n N_A_113_57#_M1002_g N_A_113_57#_M1035_g
+ N_A_113_57#_c_386_n N_A_113_57#_c_387_n N_A_113_57#_c_409_n
+ N_A_113_57#_c_410_n N_A_113_57#_M1023_g N_A_113_57#_M1041_g
+ N_A_113_57#_M1019_g N_A_113_57#_c_412_n N_A_113_57#_M1016_g
+ N_A_113_57#_c_413_n N_A_113_57#_c_389_n N_A_113_57#_c_415_n
+ N_A_113_57#_c_390_n N_A_113_57#_c_391_n N_A_113_57#_c_392_n
+ N_A_113_57#_c_393_n N_A_113_57#_c_394_n N_A_113_57#_c_395_n
+ N_A_113_57#_c_396_n N_A_113_57#_c_397_n N_A_113_57#_c_398_n
+ N_A_113_57#_c_417_n N_A_113_57#_c_418_n N_A_113_57#_c_419_n
+ N_A_113_57#_c_420_n N_A_113_57#_c_421_n N_A_113_57#_c_399_n
+ N_A_113_57#_c_400_n N_A_113_57#_c_401_n N_A_113_57#_c_402_n
+ N_A_113_57#_c_403_n N_A_113_57#_c_404_n N_A_113_57#_c_405_n
+ PM_SKY130_FD_SC_LP__DFBBN_2%A_113_57#
x_PM_SKY130_FD_SC_LP__DFBBN_2%A_789_78# N_A_789_78#_M1010_d N_A_789_78#_M1024_d
+ N_A_789_78#_M1037_g N_A_789_78#_M1039_g N_A_789_78#_M1043_g
+ N_A_789_78#_M1005_g N_A_789_78#_c_642_n N_A_789_78#_c_643_n
+ N_A_789_78#_c_687_p N_A_789_78#_c_671_p N_A_789_78#_c_633_n
+ N_A_789_78#_c_644_n N_A_789_78#_c_669_p N_A_789_78#_c_645_n
+ N_A_789_78#_c_634_n N_A_789_78#_c_635_n N_A_789_78#_c_636_n
+ N_A_789_78#_c_637_n N_A_789_78#_c_638_n PM_SKY130_FD_SC_LP__DFBBN_2%A_789_78#
x_PM_SKY130_FD_SC_LP__DFBBN_2%SET_B N_SET_B_M1017_g N_SET_B_M1024_g
+ N_SET_B_M1031_g N_SET_B_c_764_n N_SET_B_M1014_g SET_B N_SET_B_c_766_n
+ N_SET_B_c_767_n N_SET_B_c_768_n N_SET_B_c_769_n N_SET_B_c_770_n
+ PM_SKY130_FD_SC_LP__DFBBN_2%SET_B
x_PM_SKY130_FD_SC_LP__DFBBN_2%A_549_449# N_A_549_449#_M1013_d
+ N_A_549_449#_M1023_d N_A_549_449#_M1010_g N_A_549_449#_M1040_g
+ N_A_549_449#_c_890_n N_A_549_449#_c_891_n N_A_549_449#_c_899_n
+ N_A_549_449#_c_892_n N_A_549_449#_c_893_n N_A_549_449#_c_894_n
+ N_A_549_449#_c_895_n N_A_549_449#_c_944_n N_A_549_449#_c_902_n
+ N_A_549_449#_c_903_n N_A_549_449#_c_896_n N_A_549_449#_c_921_n
+ N_A_549_449#_c_905_n PM_SKY130_FD_SC_LP__DFBBN_2%A_549_449#
x_PM_SKY130_FD_SC_LP__DFBBN_2%A_223_119# N_A_223_119#_M1002_s
+ N_A_223_119#_M1035_s N_A_223_119#_M1013_g N_A_223_119#_c_1038_n
+ N_A_223_119#_c_1039_n N_A_223_119#_c_1040_n N_A_223_119#_M1030_g
+ N_A_223_119#_c_1042_n N_A_223_119#_c_1043_n N_A_223_119#_M1020_g
+ N_A_223_119#_c_1045_n N_A_223_119#_c_1046_n N_A_223_119#_c_1029_n
+ N_A_223_119#_c_1030_n N_A_223_119#_c_1031_n N_A_223_119#_c_1032_n
+ N_A_223_119#_M1015_g N_A_223_119#_c_1033_n N_A_223_119#_c_1034_n
+ N_A_223_119#_c_1035_n N_A_223_119#_c_1051_n N_A_223_119#_c_1052_n
+ N_A_223_119#_c_1036_n N_A_223_119#_c_1037_n N_A_223_119#_c_1054_n
+ PM_SKY130_FD_SC_LP__DFBBN_2%A_223_119#
x_PM_SKY130_FD_SC_LP__DFBBN_2%A_1746_137# N_A_1746_137#_M1004_d
+ N_A_1746_137#_M1014_d N_A_1746_137#_c_1197_n N_A_1746_137#_M1000_g
+ N_A_1746_137#_M1021_g N_A_1746_137#_M1011_g N_A_1746_137#_M1008_g
+ N_A_1746_137#_c_1199_n N_A_1746_137#_M1029_g N_A_1746_137#_c_1201_n
+ N_A_1746_137#_M1028_g N_A_1746_137#_c_1202_n N_A_1746_137#_c_1203_n
+ N_A_1746_137#_M1032_g N_A_1746_137#_M1006_g N_A_1746_137#_c_1205_n
+ N_A_1746_137#_c_1206_n N_A_1746_137#_c_1207_n N_A_1746_137#_c_1217_n
+ N_A_1746_137#_c_1253_p N_A_1746_137#_c_1251_p N_A_1746_137#_c_1208_n
+ N_A_1746_137#_c_1219_n N_A_1746_137#_c_1220_n N_A_1746_137#_c_1221_n
+ N_A_1746_137#_c_1222_n N_A_1746_137#_c_1223_n N_A_1746_137#_c_1262_p
+ N_A_1746_137#_c_1274_p N_A_1746_137#_c_1209_n N_A_1746_137#_c_1210_n
+ N_A_1746_137#_c_1211_n N_A_1746_137#_c_1212_n
+ PM_SKY130_FD_SC_LP__DFBBN_2%A_1746_137#
x_PM_SKY130_FD_SC_LP__DFBBN_2%A_1542_428# N_A_1542_428#_M1019_d
+ N_A_1542_428#_M1020_d N_A_1542_428#_c_1375_n N_A_1542_428#_M1004_g
+ N_A_1542_428#_M1022_g N_A_1542_428#_c_1382_n N_A_1542_428#_c_1383_n
+ N_A_1542_428#_c_1376_n N_A_1542_428#_c_1377_n N_A_1542_428#_c_1384_n
+ N_A_1542_428#_c_1378_n N_A_1542_428#_c_1379_n N_A_1542_428#_c_1380_n
+ N_A_1542_428#_c_1381_n PM_SKY130_FD_SC_LP__DFBBN_2%A_1542_428#
x_PM_SKY130_FD_SC_LP__DFBBN_2%A_1191_21# N_A_1191_21#_M1001_s
+ N_A_1191_21#_M1026_s N_A_1191_21#_M1003_g N_A_1191_21#_M1036_g
+ N_A_1191_21#_c_1472_n N_A_1191_21#_c_1473_n N_A_1191_21#_M1038_g
+ N_A_1191_21#_M1009_g N_A_1191_21#_c_1475_n N_A_1191_21#_c_1476_n
+ N_A_1191_21#_c_1477_n N_A_1191_21#_c_1478_n N_A_1191_21#_c_1483_n
+ N_A_1191_21#_c_1484_n N_A_1191_21#_c_1479_n
+ PM_SKY130_FD_SC_LP__DFBBN_2%A_1191_21#
x_PM_SKY130_FD_SC_LP__DFBBN_2%RESET_B N_RESET_B_c_1581_n N_RESET_B_M1026_g
+ N_RESET_B_M1001_g N_RESET_B_c_1584_n RESET_B N_RESET_B_c_1585_n
+ N_RESET_B_c_1586_n PM_SKY130_FD_SC_LP__DFBBN_2%RESET_B
x_PM_SKY130_FD_SC_LP__DFBBN_2%A_2618_131# N_A_2618_131#_M1032_s
+ N_A_2618_131#_M1006_s N_A_2618_131#_M1018_g N_A_2618_131#_M1007_g
+ N_A_2618_131#_c_1621_n N_A_2618_131#_M1033_g N_A_2618_131#_M1027_g
+ N_A_2618_131#_c_1624_n N_A_2618_131#_c_1625_n N_A_2618_131#_c_1626_n
+ N_A_2618_131#_c_1627_n N_A_2618_131#_c_1628_n N_A_2618_131#_c_1629_n
+ PM_SKY130_FD_SC_LP__DFBBN_2%A_2618_131#
x_PM_SKY130_FD_SC_LP__DFBBN_2%VPWR N_VPWR_M1034_s N_VPWR_M1035_d N_VPWR_M1039_d
+ N_VPWR_M1036_d N_VPWR_M1021_d N_VPWR_M1009_d N_VPWR_M1026_d N_VPWR_M1029_d
+ N_VPWR_M1006_d N_VPWR_M1027_s N_VPWR_c_1696_n N_VPWR_c_1697_n N_VPWR_c_1698_n
+ N_VPWR_c_1699_n N_VPWR_c_1700_n N_VPWR_c_1701_n N_VPWR_c_1702_n
+ N_VPWR_c_1703_n N_VPWR_c_1704_n N_VPWR_c_1705_n N_VPWR_c_1706_n
+ N_VPWR_c_1707_n N_VPWR_c_1708_n N_VPWR_c_1709_n N_VPWR_c_1710_n
+ N_VPWR_c_1711_n VPWR N_VPWR_c_1712_n N_VPWR_c_1713_n N_VPWR_c_1714_n
+ N_VPWR_c_1715_n N_VPWR_c_1716_n N_VPWR_c_1717_n N_VPWR_c_1718_n
+ N_VPWR_c_1719_n N_VPWR_c_1720_n N_VPWR_c_1721_n N_VPWR_c_1722_n
+ N_VPWR_c_1723_n N_VPWR_c_1724_n N_VPWR_c_1695_n
+ PM_SKY130_FD_SC_LP__DFBBN_2%VPWR
x_PM_SKY130_FD_SC_LP__DFBBN_2%A_463_449# N_A_463_449#_M1012_d
+ N_A_463_449#_M1042_d N_A_463_449#_c_1849_n N_A_463_449#_c_1850_n
+ N_A_463_449#_c_1853_n N_A_463_449#_c_1851_n
+ PM_SKY130_FD_SC_LP__DFBBN_2%A_463_449#
x_PM_SKY130_FD_SC_LP__DFBBN_2%Q_N N_Q_N_M1008_d N_Q_N_M1011_s N_Q_N_c_1907_n
+ N_Q_N_c_1908_n N_Q_N_c_1915_n N_Q_N_c_1906_n Q_N N_Q_N_c_1927_n
+ PM_SKY130_FD_SC_LP__DFBBN_2%Q_N
x_PM_SKY130_FD_SC_LP__DFBBN_2%Q N_Q_M1018_d N_Q_M1007_d N_Q_c_1945_n
+ N_Q_c_1940_n N_Q_c_1943_n Q Q N_Q_c_1965_n Q PM_SKY130_FD_SC_LP__DFBBN_2%Q
x_PM_SKY130_FD_SC_LP__DFBBN_2%VGND N_VGND_M1025_s N_VGND_M1002_d N_VGND_M1037_d
+ N_VGND_M1043_s N_VGND_M1000_d N_VGND_M1001_d N_VGND_M1028_s N_VGND_M1032_d
+ N_VGND_M1033_s N_VGND_c_1975_n N_VGND_c_1976_n N_VGND_c_1977_n N_VGND_c_1978_n
+ N_VGND_c_1979_n N_VGND_c_1980_n N_VGND_c_1981_n N_VGND_c_1982_n
+ N_VGND_c_1983_n N_VGND_c_1984_n N_VGND_c_1985_n N_VGND_c_1986_n
+ N_VGND_c_1987_n VGND N_VGND_c_1988_n N_VGND_c_1989_n N_VGND_c_1990_n
+ N_VGND_c_1991_n N_VGND_c_1992_n N_VGND_c_1993_n N_VGND_c_1994_n
+ N_VGND_c_1995_n N_VGND_c_1996_n N_VGND_c_1997_n N_VGND_c_1998_n
+ N_VGND_c_1999_n N_VGND_c_2000_n N_VGND_c_2001_n
+ PM_SKY130_FD_SC_LP__DFBBN_2%VGND
x_PM_SKY130_FD_SC_LP__DFBBN_2%A_1018_60# N_A_1018_60#_M1017_d
+ N_A_1018_60#_M1003_d N_A_1018_60#_c_2123_n N_A_1018_60#_c_2124_n
+ N_A_1018_60#_c_2125_n PM_SKY130_FD_SC_LP__DFBBN_2%A_1018_60#
x_PM_SKY130_FD_SC_LP__DFBBN_2%A_1911_119# N_A_1911_119#_M1031_d
+ N_A_1911_119#_M1038_d N_A_1911_119#_c_2148_n N_A_1911_119#_c_2149_n
+ N_A_1911_119#_c_2150_n N_A_1911_119#_c_2151_n
+ PM_SKY130_FD_SC_LP__DFBBN_2%A_1911_119#
cc_1 VNB N_CLK_N_c_294_n 0.0045875f $X=-0.19 $Y=-0.245 $X2=0.36 $Y2=2.18
cc_2 VNB N_CLK_N_M1025_g 0.0324132f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=0.495
cc_3 VNB N_CLK_N_c_296_n 0.034855f $X=-0.19 $Y=-0.245 $X2=0.335 $Y2=1.06
cc_4 VNB N_CLK_N_c_297_n 0.0222509f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.58
cc_5 VNB N_CLK_N_c_298_n 0.0383496f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.075
cc_6 VNB N_CLK_N_c_299_n 0.00767254f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.075
cc_7 VNB N_D_c_328_n 0.00894256f $X=-0.19 $Y=-0.245 $X2=0.36 $Y2=2.18
cc_8 VNB N_D_c_329_n 0.0284751f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=0.91
cc_9 VNB N_D_c_330_n 0.0160067f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=2.725
cc_10 VNB N_D_c_331_n 0.0442973f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=2.255
cc_11 VNB N_D_c_332_n 0.0104929f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.95
cc_12 VNB N_A_113_57#_c_383_n 0.0336595f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=2.33
cc_13 VNB N_A_113_57#_c_384_n 0.0163801f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=2.725
cc_14 VNB N_A_113_57#_M1002_g 0.039936f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.58
cc_15 VNB N_A_113_57#_c_386_n 0.153256f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_16 VNB N_A_113_57#_c_387_n 0.012806f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_17 VNB N_A_113_57#_M1041_g 0.032268f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.295
cc_18 VNB N_A_113_57#_c_389_n 0.00118519f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_113_57#_c_390_n 0.0484447f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_113_57#_c_391_n 0.044682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_113_57#_c_392_n 0.00466338f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_113_57#_c_393_n 0.00329926f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_113_57#_c_394_n 0.0215835f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_113_57#_c_395_n 0.00165293f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_113_57#_c_396_n 0.0153813f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_113_57#_c_397_n 0.00883394f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_113_57#_c_398_n 0.0042523f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_113_57#_c_399_n 0.0117145f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_113_57#_c_400_n 0.00664267f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_113_57#_c_401_n 0.0123356f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_113_57#_c_402_n 0.0117849f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_113_57#_c_403_n 0.00387779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_113_57#_c_404_n 0.0239236f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_113_57#_c_405_n 0.0186391f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_789_78#_M1037_g 0.0585965f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=2.725
cc_36 VNB N_A_789_78#_M1043_g 0.024468f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=2.255
cc_37 VNB N_A_789_78#_c_633_n 0.0015086f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_789_78#_c_634_n 0.00714372f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_789_78#_c_635_n 0.00124707f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_789_78#_c_636_n 6.43647e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_789_78#_c_637_n 0.0271889f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_789_78#_c_638_n 0.0213795f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_SET_B_M1017_g 0.0438126f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=0.91
cc_44 VNB N_SET_B_M1031_g 0.0220454f $X=-0.19 $Y=-0.245 $X2=0.335 $Y2=0.91
cc_45 VNB N_SET_B_c_764_n 0.0147187f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.415
cc_46 VNB SET_B 0.00580316f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_SET_B_c_766_n 0.0203228f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_SET_B_c_767_n 5.76378e-19 $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_49 VNB N_SET_B_c_768_n 0.00103874f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.075
cc_50 VNB N_SET_B_c_769_n 0.0234425f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_SET_B_c_770_n 0.00250627f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.295
cc_52 VNB N_A_549_449#_M1010_g 0.0388507f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=2.725
cc_53 VNB N_A_549_449#_c_890_n 0.00212616f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=2.255
cc_54 VNB N_A_549_449#_c_891_n 0.0109327f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_55 VNB N_A_549_449#_c_892_n 4.72401e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_549_449#_c_893_n 0.0161638f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.075
cc_57 VNB N_A_549_449#_c_894_n 0.0022362f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.075
cc_58 VNB N_A_549_449#_c_895_n 0.00163838f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.075
cc_59 VNB N_A_549_449#_c_896_n 0.0216532f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=2.035
cc_60 VNB N_A_223_119#_M1013_g 0.0358666f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=2.725
cc_61 VNB N_A_223_119#_c_1029_n 0.011445f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.075
cc_62 VNB N_A_223_119#_c_1030_n 0.0222083f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_A_223_119#_c_1031_n 0.00817729f $X=-0.19 $Y=-0.245 $X2=0.27
+ $Y2=1.295
cc_64 VNB N_A_223_119#_c_1032_n 0.0155813f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_65 VNB N_A_223_119#_c_1033_n 0.0207648f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=2.035
cc_66 VNB N_A_223_119#_c_1034_n 0.00621013f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_A_223_119#_c_1035_n 0.00954073f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_A_223_119#_c_1036_n 0.00276064f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_223_119#_c_1037_n 0.00782901f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_A_1746_137#_c_1197_n 0.015331f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=2.33
cc_71 VNB N_A_1746_137#_M1011_g 6.92337e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_A_1746_137#_c_1199_n 0.0141455f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_A_1746_137#_M1029_g 0.0110774f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.075
cc_74 VNB N_A_1746_137#_c_1201_n 0.0194771f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_A_1746_137#_c_1202_n 0.0577467f $X=-0.19 $Y=-0.245 $X2=0.27
+ $Y2=1.665
cc_76 VNB N_A_1746_137#_c_1203_n 0.0205703f $X=-0.19 $Y=-0.245 $X2=0.27
+ $Y2=2.035
cc_77 VNB N_A_1746_137#_M1006_g 0.0184049f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_A_1746_137#_c_1205_n 0.0195533f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_A_1746_137#_c_1206_n 0.0025471f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_A_1746_137#_c_1207_n 0.00515104f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_A_1746_137#_c_1208_n 0.00275509f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_A_1746_137#_c_1209_n 0.00327461f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_A_1746_137#_c_1210_n 0.0109072f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_A_1746_137#_c_1211_n 0.0304352f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_A_1746_137#_c_1212_n 0.0193752f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_A_1542_428#_c_1375_n 0.0153044f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=2.33
cc_87 VNB N_A_1542_428#_c_1376_n 0.00865175f $X=-0.19 $Y=-0.245 $X2=0.155
+ $Y2=1.21
cc_88 VNB N_A_1542_428#_c_1377_n 0.00928006f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_A_1542_428#_c_1378_n 0.00227559f $X=-0.19 $Y=-0.245 $X2=0.27
+ $Y2=1.075
cc_90 VNB N_A_1542_428#_c_1379_n 9.85316e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_A_1542_428#_c_1380_n 0.00779479f $X=-0.19 $Y=-0.245 $X2=0.27
+ $Y2=1.295
cc_92 VNB N_A_1542_428#_c_1381_n 0.0297039f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_93 VNB N_A_1191_21#_M1003_g 0.0485541f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=2.725
cc_94 VNB N_A_1191_21#_c_1472_n 0.34851f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.415
cc_95 VNB N_A_1191_21#_c_1473_n 0.011382f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.58
cc_96 VNB N_A_1191_21#_M1038_g 0.0293122f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_97 VNB N_A_1191_21#_c_1475_n 0.00707796f $X=-0.19 $Y=-0.245 $X2=0.27
+ $Y2=1.075
cc_98 VNB N_A_1191_21#_c_1476_n 0.0376552f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.075
cc_99 VNB N_A_1191_21#_c_1477_n 0.0121008f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.075
cc_100 VNB N_A_1191_21#_c_1478_n 0.00273074f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_101 VNB N_A_1191_21#_c_1479_n 0.00261783f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_102 VNB N_RESET_B_c_1581_n 0.011873f $X=-0.19 $Y=-0.245 $X2=0.36 $Y2=2.18
cc_103 VNB N_RESET_B_M1026_g 0.00109887f $X=-0.19 $Y=-0.245 $X2=0.49 $Y2=0.495
cc_104 VNB N_RESET_B_M1001_g 0.0228988f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=2.725
cc_105 VNB N_RESET_B_c_1584_n 0.022018f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.415
cc_106 VNB N_RESET_B_c_1585_n 0.00350543f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.95
cc_107 VNB N_RESET_B_c_1586_n 0.0321013f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_108 VNB N_A_2618_131#_M1018_g 0.0241958f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=2.725
cc_109 VNB N_A_2618_131#_M1007_g 0.00270422f $X=-0.19 $Y=-0.245 $X2=0.27
+ $Y2=1.415
cc_110 VNB N_A_2618_131#_c_1621_n 0.0117009f $X=-0.19 $Y=-0.245 $X2=0.36
+ $Y2=2.255
cc_111 VNB N_A_2618_131#_M1033_g 0.0284516f $X=-0.19 $Y=-0.245 $X2=0.155
+ $Y2=1.21
cc_112 VNB N_A_2618_131#_M1027_g 0.0169713f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_113 VNB N_A_2618_131#_c_1624_n 0.0106548f $X=-0.19 $Y=-0.245 $X2=0.27
+ $Y2=1.075
cc_114 VNB N_A_2618_131#_c_1625_n 0.00922808f $X=-0.19 $Y=-0.245 $X2=0.27
+ $Y2=1.075
cc_115 VNB N_A_2618_131#_c_1626_n 8.37508e-19 $X=-0.19 $Y=-0.245 $X2=0.27
+ $Y2=1.665
cc_116 VNB N_A_2618_131#_c_1627_n 0.00889868f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_117 VNB N_A_2618_131#_c_1628_n 0.00384711f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_118 VNB N_A_2618_131#_c_1629_n 0.0276806f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_119 VNB N_VPWR_c_1695_n 0.621437f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_120 VNB N_A_463_449#_c_1849_n 0.0022778f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=2.725
cc_121 VNB N_A_463_449#_c_1850_n 0.00422891f $X=-0.19 $Y=-0.245 $X2=0.335
+ $Y2=1.06
cc_122 VNB N_A_463_449#_c_1851_n 0.00491568f $X=-0.19 $Y=-0.245 $X2=0.6
+ $Y2=2.255
cc_123 VNB N_Q_N_c_1906_n 0.00221375f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=2.255
cc_124 VNB N_Q_c_1940_n 0.00291898f $X=-0.19 $Y=-0.245 $X2=0.36 $Y2=2.255
cc_125 VNB Q 0.00497765f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_126 VNB N_VGND_c_1975_n 0.0105185f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.075
cc_127 VNB N_VGND_c_1976_n 0.0257426f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.295
cc_128 VNB N_VGND_c_1977_n 0.015112f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=2.035
cc_129 VNB N_VGND_c_1978_n 0.0109935f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_130 VNB N_VGND_c_1979_n 0.0117815f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_131 VNB N_VGND_c_1980_n 0.0229811f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_132 VNB N_VGND_c_1981_n 0.00841408f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_133 VNB N_VGND_c_1982_n 0.0241118f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_134 VNB N_VGND_c_1983_n 0.0194232f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_135 VNB N_VGND_c_1984_n 0.0105185f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_136 VNB N_VGND_c_1985_n 0.0247507f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_137 VNB N_VGND_c_1986_n 0.0683427f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_138 VNB N_VGND_c_1987_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_139 VNB N_VGND_c_1988_n 0.033678f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_140 VNB N_VGND_c_1989_n 0.054773f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_141 VNB N_VGND_c_1990_n 0.0574553f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_142 VNB N_VGND_c_1991_n 0.0567805f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_143 VNB N_VGND_c_1992_n 0.0188675f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_144 VNB N_VGND_c_1993_n 0.0220244f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_145 VNB N_VGND_c_1994_n 0.0188675f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_146 VNB N_VGND_c_1995_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_147 VNB N_VGND_c_1996_n 0.00332923f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_148 VNB N_VGND_c_1997_n 0.00439458f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_149 VNB N_VGND_c_1998_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_150 VNB N_VGND_c_1999_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_151 VNB N_VGND_c_2000_n 0.00480869f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_152 VNB N_VGND_c_2001_n 0.747047f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_153 VNB N_A_1018_60#_c_2123_n 0.00113325f $X=-0.19 $Y=-0.245 $X2=0.6 $Y2=2.33
cc_154 VNB N_A_1018_60#_c_2124_n 0.00819986f $X=-0.19 $Y=-0.245 $X2=0.335
+ $Y2=1.06
cc_155 VNB N_A_1018_60#_c_2125_n 0.00135248f $X=-0.19 $Y=-0.245 $X2=0.36
+ $Y2=2.255
cc_156 VNB N_A_1911_119#_c_2148_n 7.02193e-19 $X=-0.19 $Y=-0.245 $X2=0.6
+ $Y2=2.725
cc_157 VNB N_A_1911_119#_c_2149_n 0.00794203f $X=-0.19 $Y=-0.245 $X2=0.335
+ $Y2=0.91
cc_158 VNB N_A_1911_119#_c_2150_n 0.00339258f $X=-0.19 $Y=-0.245 $X2=0.335
+ $Y2=1.06
cc_159 VNB N_A_1911_119#_c_2151_n 0.00621621f $X=-0.19 $Y=-0.245 $X2=0.27
+ $Y2=1.415
cc_160 VPB N_CLK_N_c_294_n 0.0341664f $X=-0.19 $Y=1.655 $X2=0.36 $Y2=2.18
cc_161 VPB N_CLK_N_c_301_n 0.0218224f $X=-0.19 $Y=1.655 $X2=0.6 $Y2=2.33
cc_162 VPB N_CLK_N_c_302_n 0.0372746f $X=-0.19 $Y=1.655 $X2=0.6 $Y2=2.255
cc_163 VPB N_CLK_N_c_299_n 0.0213933f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.075
cc_164 VPB N_D_c_328_n 0.0214798f $X=-0.19 $Y=1.655 $X2=0.36 $Y2=2.18
cc_165 VPB N_D_c_334_n 0.0148263f $X=-0.19 $Y=1.655 $X2=0.49 $Y2=0.495
cc_166 VPB N_D_c_335_n 0.0288009f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.415
cc_167 VPB N_A_113_57#_c_406_n 0.0454269f $X=-0.19 $Y=1.655 $X2=0.6 $Y2=2.725
cc_168 VPB N_A_113_57#_c_407_n 0.0163801f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.06
cc_169 VPB N_A_113_57#_M1035_g 0.0249616f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_170 VPB N_A_113_57#_c_409_n 0.0771781f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.95
cc_171 VPB N_A_113_57#_c_410_n 0.01298f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_172 VPB N_A_113_57#_M1023_g 0.0343117f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.075
cc_173 VPB N_A_113_57#_c_412_n 0.0158937f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=2.035
cc_174 VPB N_A_113_57#_c_413_n 0.0372569f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_175 VPB N_A_113_57#_c_389_n 0.018142f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_176 VPB N_A_113_57#_c_415_n 0.00230797f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_177 VPB N_A_113_57#_c_390_n 0.0146617f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_178 VPB N_A_113_57#_c_417_n 0.00615028f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_179 VPB N_A_113_57#_c_418_n 0.00826537f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_180 VPB N_A_113_57#_c_419_n 0.00448393f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_181 VPB N_A_113_57#_c_420_n 0.00320051f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_182 VPB N_A_113_57#_c_421_n 0.0511693f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_183 VPB N_A_113_57#_c_401_n 0.00949494f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_184 VPB N_A_113_57#_c_403_n 0.0030602f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_185 VPB N_A_113_57#_c_404_n 0.0068863f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_186 VPB N_A_789_78#_M1037_g 0.00543354f $X=-0.19 $Y=1.655 $X2=0.6 $Y2=2.725
cc_187 VPB N_A_789_78#_M1039_g 0.0205587f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.415
cc_188 VPB N_A_789_78#_M1005_g 0.0240798f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.95
cc_189 VPB N_A_789_78#_c_642_n 0.00488486f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.075
cc_190 VPB N_A_789_78#_c_643_n 0.055182f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.075
cc_191 VPB N_A_789_78#_c_644_n 0.0013286f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_192 VPB N_A_789_78#_c_645_n 0.00226117f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_193 VPB N_A_789_78#_c_636_n 0.00101696f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_194 VPB N_A_789_78#_c_637_n 0.0164463f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_195 VPB N_SET_B_M1024_g 0.0193697f $X=-0.19 $Y=1.655 $X2=0.6 $Y2=2.33
cc_196 VPB N_SET_B_c_764_n 0.0648922f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.415
cc_197 VPB SET_B 0.00780964f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_198 VPB N_SET_B_c_766_n 0.044356f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_199 VPB N_SET_B_c_767_n 0.00168997f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_200 VPB N_SET_B_c_768_n 0.00254874f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.075
cc_201 VPB N_SET_B_c_769_n 0.0105079f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_202 VPB N_SET_B_c_770_n 5.71498e-19 $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.295
cc_203 VPB N_A_549_449#_M1040_g 0.0170589f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.415
cc_204 VPB N_A_549_449#_c_891_n 0.00485084f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_205 VPB N_A_549_449#_c_899_n 0.00572233f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.95
cc_206 VPB N_A_549_449#_c_892_n 0.0051743f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_207 VPB N_A_549_449#_c_895_n 0.00563448f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.075
cc_208 VPB N_A_549_449#_c_902_n 0.00266878f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.295
cc_209 VPB N_A_549_449#_c_903_n 0.00231243f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_210 VPB N_A_549_449#_c_896_n 0.00975948f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=2.035
cc_211 VPB N_A_549_449#_c_905_n 0.00616579f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_212 VPB N_A_223_119#_c_1038_n 0.012397f $X=-0.19 $Y=1.655 $X2=0.335 $Y2=1.06
cc_213 VPB N_A_223_119#_c_1039_n 0.0285616f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.415
cc_214 VPB N_A_223_119#_c_1040_n 0.0132591f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.58
cc_215 VPB N_A_223_119#_M1030_g 0.0410009f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_216 VPB N_A_223_119#_c_1042_n 0.32504f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_217 VPB N_A_223_119#_c_1043_n 0.0118952f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_218 VPB N_A_223_119#_M1020_g 0.0105781f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_219 VPB N_A_223_119#_c_1045_n 0.0264454f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.075
cc_220 VPB N_A_223_119#_c_1046_n 0.00830324f $X=-0.19 $Y=1.655 $X2=0.27
+ $Y2=1.075
cc_221 VPB N_A_223_119#_c_1029_n 0.0159779f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.075
cc_222 VPB N_A_223_119#_c_1033_n 0.0215608f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=2.035
cc_223 VPB N_A_223_119#_c_1034_n 0.0277337f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_224 VPB N_A_223_119#_c_1035_n 0.00353284f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_225 VPB N_A_223_119#_c_1051_n 0.0109388f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_226 VPB N_A_223_119#_c_1052_n 0.0133734f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_227 VPB N_A_223_119#_c_1036_n 0.00113661f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_228 VPB N_A_223_119#_c_1054_n 7.52486e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_229 VPB N_A_1746_137#_M1021_g 0.0244725f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.58
cc_230 VPB N_A_1746_137#_M1011_g 0.0217807f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_231 VPB N_A_1746_137#_M1029_g 0.0225454f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.075
cc_232 VPB N_A_1746_137#_M1006_g 0.0259848f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_233 VPB N_A_1746_137#_c_1217_n 0.00661303f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_234 VPB N_A_1746_137#_c_1208_n 0.00438727f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_235 VPB N_A_1746_137#_c_1219_n 0.0245978f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_236 VPB N_A_1746_137#_c_1220_n 0.00173733f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_237 VPB N_A_1746_137#_c_1221_n 0.00852246f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_238 VPB N_A_1746_137#_c_1222_n 0.0342917f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_239 VPB N_A_1746_137#_c_1223_n 0.00232136f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_240 VPB N_A_1746_137#_c_1210_n 0.0193031f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_241 VPB N_A_1542_428#_c_1382_n 0.0141154f $X=-0.19 $Y=1.655 $X2=0.36
+ $Y2=2.255
cc_242 VPB N_A_1542_428#_c_1383_n 0.0265306f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_243 VPB N_A_1542_428#_c_1384_n 0.00249191f $X=-0.19 $Y=1.655 $X2=0.27
+ $Y2=1.075
cc_244 VPB N_A_1542_428#_c_1378_n 0.00382998f $X=-0.19 $Y=1.655 $X2=0.27
+ $Y2=1.075
cc_245 VPB N_A_1542_428#_c_1380_n 0.00400609f $X=-0.19 $Y=1.655 $X2=0.27
+ $Y2=1.295
cc_246 VPB N_A_1542_428#_c_1381_n 0.00845771f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_247 VPB N_A_1191_21#_M1003_g 0.0267835f $X=-0.19 $Y=1.655 $X2=0.6 $Y2=2.725
cc_248 VPB N_A_1191_21#_M1009_g 0.0387486f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.95
cc_249 VPB N_A_1191_21#_c_1476_n 0.0156993f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.075
cc_250 VPB N_A_1191_21#_c_1483_n 0.00990936f $X=-0.19 $Y=1.655 $X2=0.27
+ $Y2=1.295
cc_251 VPB N_A_1191_21#_c_1484_n 0.0112496f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.665
cc_252 VPB N_RESET_B_M1026_g 0.0282022f $X=-0.19 $Y=1.655 $X2=0.49 $Y2=0.495
cc_253 VPB N_A_2618_131#_M1007_g 0.0230272f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.415
cc_254 VPB N_A_2618_131#_M1027_g 0.027002f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_255 VPB N_A_2618_131#_c_1626_n 0.014571f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.665
cc_256 VPB N_VPWR_c_1696_n 0.0129883f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_257 VPB N_VPWR_c_1697_n 0.0365848f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_258 VPB N_VPWR_c_1698_n 0.0109716f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_259 VPB N_VPWR_c_1699_n 0.0220921f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_260 VPB N_VPWR_c_1700_n 0.024766f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_261 VPB N_VPWR_c_1701_n 0.00906969f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_262 VPB N_VPWR_c_1702_n 0.0254052f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_263 VPB N_VPWR_c_1703_n 0.0250032f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_264 VPB N_VPWR_c_1704_n 0.0362339f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_265 VPB N_VPWR_c_1705_n 0.0268954f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_266 VPB N_VPWR_c_1706_n 0.0104926f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_267 VPB N_VPWR_c_1707_n 0.0413598f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_268 VPB N_VPWR_c_1708_n 0.0336598f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_269 VPB N_VPWR_c_1709_n 0.00522307f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_270 VPB N_VPWR_c_1710_n 0.0775185f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_271 VPB N_VPWR_c_1711_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_272 VPB N_VPWR_c_1712_n 0.0367642f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_273 VPB N_VPWR_c_1713_n 0.0758757f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_274 VPB N_VPWR_c_1714_n 0.0278365f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_275 VPB N_VPWR_c_1715_n 0.0233255f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_276 VPB N_VPWR_c_1716_n 0.0173868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_277 VPB N_VPWR_c_1717_n 0.0234846f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_278 VPB N_VPWR_c_1718_n 0.0188675f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_279 VPB N_VPWR_c_1719_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_280 VPB N_VPWR_c_1720_n 0.0047828f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_281 VPB N_VPWR_c_1721_n 0.00598038f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_282 VPB N_VPWR_c_1722_n 0.0060562f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_283 VPB N_VPWR_c_1723_n 0.0047828f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_284 VPB N_VPWR_c_1724_n 0.0047828f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_285 VPB N_VPWR_c_1695_n 0.174711f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_286 VPB N_A_463_449#_c_1850_n 0.00538697f $X=-0.19 $Y=1.655 $X2=0.335
+ $Y2=1.06
cc_287 VPB N_A_463_449#_c_1853_n 0.0028426f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.58
cc_288 VPB N_Q_N_c_1907_n 0.00129605f $X=-0.19 $Y=1.655 $X2=0.6 $Y2=2.33
cc_289 VPB N_Q_N_c_1908_n 0.00203429f $X=-0.19 $Y=1.655 $X2=0.6 $Y2=2.725
cc_290 VPB N_Q_N_c_1906_n 0.00114162f $X=-0.19 $Y=1.655 $X2=0.6 $Y2=2.255
cc_291 VPB N_Q_c_1940_n 8.09705e-19 $X=-0.19 $Y=1.655 $X2=0.36 $Y2=2.255
cc_292 VPB N_Q_c_1943_n 0.00277912f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_293 N_CLK_N_c_298_n N_A_113_57#_c_384_n 0.011491f $X=0.27 $Y=1.075 $X2=0
+ $Y2=0
cc_294 N_CLK_N_c_299_n N_A_113_57#_c_384_n 8.1212e-19 $X=0.27 $Y=1.075 $X2=0
+ $Y2=0
cc_295 N_CLK_N_c_294_n N_A_113_57#_c_407_n 0.011491f $X=0.36 $Y=2.18 $X2=0 $Y2=0
cc_296 N_CLK_N_c_294_n N_A_113_57#_c_389_n 0.0045399f $X=0.36 $Y=2.18 $X2=0
+ $Y2=0
cc_297 N_CLK_N_c_301_n N_A_113_57#_c_389_n 0.0118675f $X=0.6 $Y=2.33 $X2=0 $Y2=0
cc_298 N_CLK_N_c_302_n N_A_113_57#_c_389_n 0.0106572f $X=0.6 $Y=2.255 $X2=0
+ $Y2=0
cc_299 N_CLK_N_M1025_g N_A_113_57#_c_399_n 0.00771309f $X=0.49 $Y=0.495 $X2=0
+ $Y2=0
cc_300 N_CLK_N_c_297_n N_A_113_57#_c_400_n 0.0045399f $X=0.27 $Y=1.58 $X2=0
+ $Y2=0
cc_301 N_CLK_N_c_297_n N_A_113_57#_c_401_n 0.011491f $X=0.27 $Y=1.58 $X2=0 $Y2=0
cc_302 N_CLK_N_M1025_g N_A_113_57#_c_402_n 0.0112284f $X=0.49 $Y=0.495 $X2=0
+ $Y2=0
cc_303 N_CLK_N_c_298_n N_A_113_57#_c_402_n 0.0045399f $X=0.27 $Y=1.075 $X2=0
+ $Y2=0
cc_304 N_CLK_N_c_299_n N_A_113_57#_c_402_n 0.0816843f $X=0.27 $Y=1.075 $X2=0
+ $Y2=0
cc_305 N_CLK_N_c_302_n N_A_223_119#_c_1051_n 0.00161331f $X=0.6 $Y=2.255 $X2=0
+ $Y2=0
cc_306 N_CLK_N_M1025_g N_A_223_119#_c_1037_n 3.32013e-19 $X=0.49 $Y=0.495 $X2=0
+ $Y2=0
cc_307 N_CLK_N_c_301_n N_VPWR_c_1697_n 0.0171119f $X=0.6 $Y=2.33 $X2=0 $Y2=0
cc_308 N_CLK_N_c_302_n N_VPWR_c_1697_n 0.00649475f $X=0.6 $Y=2.255 $X2=0 $Y2=0
cc_309 N_CLK_N_c_299_n N_VPWR_c_1697_n 0.0211391f $X=0.27 $Y=1.075 $X2=0 $Y2=0
cc_310 N_CLK_N_c_301_n N_VPWR_c_1708_n 0.00502664f $X=0.6 $Y=2.33 $X2=0 $Y2=0
cc_311 N_CLK_N_c_301_n N_VPWR_c_1695_n 0.0110321f $X=0.6 $Y=2.33 $X2=0 $Y2=0
cc_312 N_CLK_N_M1025_g N_VGND_c_1976_n 0.00533583f $X=0.49 $Y=0.495 $X2=0 $Y2=0
cc_313 N_CLK_N_c_296_n N_VGND_c_1976_n 0.00192064f $X=0.335 $Y=1.06 $X2=0 $Y2=0
cc_314 N_CLK_N_c_299_n N_VGND_c_1976_n 0.0207349f $X=0.27 $Y=1.075 $X2=0 $Y2=0
cc_315 N_CLK_N_M1025_g N_VGND_c_1988_n 0.00502664f $X=0.49 $Y=0.495 $X2=0 $Y2=0
cc_316 N_CLK_N_M1025_g N_VGND_c_2001_n 0.0109735f $X=0.49 $Y=0.495 $X2=0 $Y2=0
cc_317 N_D_c_328_n N_A_113_57#_c_406_n 0.00986581f $X=1.98 $Y=2.02 $X2=0 $Y2=0
cc_318 N_D_c_332_n N_A_113_57#_c_406_n 0.00247124f $X=1.92 $Y=1.345 $X2=0 $Y2=0
cc_319 N_D_c_331_n N_A_113_57#_M1002_g 0.0230397f $X=1.92 $Y=1.165 $X2=0 $Y2=0
cc_320 N_D_c_332_n N_A_113_57#_M1002_g 0.00229009f $X=1.92 $Y=1.345 $X2=0 $Y2=0
cc_321 N_D_c_334_n N_A_113_57#_M1035_g 0.00963216f $X=2.24 $Y=2.17 $X2=0 $Y2=0
cc_322 N_D_c_335_n N_A_113_57#_M1035_g 0.00986581f $X=2.24 $Y=2.095 $X2=0 $Y2=0
cc_323 N_D_c_330_n N_A_113_57#_c_386_n 0.0103003f $X=2.395 $Y=1.09 $X2=0 $Y2=0
cc_324 N_D_c_334_n N_A_113_57#_c_409_n 0.0104235f $X=2.24 $Y=2.17 $X2=0 $Y2=0
cc_325 N_D_c_335_n N_A_113_57#_M1023_g 0.0134253f $X=2.24 $Y=2.095 $X2=0 $Y2=0
cc_326 N_D_c_330_n N_A_223_119#_M1013_g 0.0177261f $X=2.395 $Y=1.09 $X2=0 $Y2=0
cc_327 N_D_c_331_n N_A_223_119#_M1013_g 0.00261043f $X=1.92 $Y=1.165 $X2=0 $Y2=0
cc_328 N_D_c_332_n N_A_223_119#_M1013_g 3.3113e-19 $X=1.92 $Y=1.345 $X2=0 $Y2=0
cc_329 N_D_c_335_n N_A_223_119#_c_1040_n 0.0010987f $X=2.24 $Y=2.095 $X2=0 $Y2=0
cc_330 N_D_c_328_n N_A_223_119#_c_1033_n 0.017832f $X=1.98 $Y=2.02 $X2=0 $Y2=0
cc_331 N_D_c_329_n N_A_223_119#_c_1033_n 0.0097091f $X=2.32 $Y=1.165 $X2=0 $Y2=0
cc_332 N_D_c_335_n N_A_223_119#_c_1033_n 0.00130767f $X=2.24 $Y=2.095 $X2=0
+ $Y2=0
cc_333 N_D_c_331_n N_A_223_119#_c_1033_n 0.00198685f $X=1.92 $Y=1.165 $X2=0
+ $Y2=0
cc_334 N_D_c_328_n N_A_223_119#_c_1035_n 0.00751343f $X=1.98 $Y=2.02 $X2=0 $Y2=0
cc_335 N_D_c_331_n N_A_223_119#_c_1035_n 3.70559e-19 $X=1.92 $Y=1.165 $X2=0
+ $Y2=0
cc_336 N_D_c_332_n N_A_223_119#_c_1035_n 0.0249384f $X=1.92 $Y=1.345 $X2=0 $Y2=0
cc_337 N_D_c_334_n N_A_223_119#_c_1051_n 3.37307e-19 $X=2.24 $Y=2.17 $X2=0 $Y2=0
cc_338 N_D_c_335_n N_A_223_119#_c_1051_n 6.81575e-19 $X=2.24 $Y=2.095 $X2=0
+ $Y2=0
cc_339 N_D_c_328_n N_A_223_119#_c_1052_n 0.00982076f $X=1.98 $Y=2.02 $X2=0 $Y2=0
cc_340 N_D_c_329_n N_A_223_119#_c_1052_n 0.00442355f $X=2.32 $Y=1.165 $X2=0
+ $Y2=0
cc_341 N_D_c_335_n N_A_223_119#_c_1052_n 0.0172458f $X=2.24 $Y=2.095 $X2=0 $Y2=0
cc_342 N_D_c_331_n N_A_223_119#_c_1052_n 0.00330121f $X=1.92 $Y=1.165 $X2=0
+ $Y2=0
cc_343 N_D_c_332_n N_A_223_119#_c_1052_n 0.0219435f $X=1.92 $Y=1.345 $X2=0 $Y2=0
cc_344 N_D_c_328_n N_A_223_119#_c_1036_n 0.00410683f $X=1.98 $Y=2.02 $X2=0 $Y2=0
cc_345 N_D_c_329_n N_A_223_119#_c_1036_n 0.00112825f $X=2.32 $Y=1.165 $X2=0
+ $Y2=0
cc_346 N_D_c_332_n N_A_223_119#_c_1036_n 0.00188136f $X=1.92 $Y=1.345 $X2=0
+ $Y2=0
cc_347 N_D_c_334_n N_VPWR_c_1698_n 0.0090293f $X=2.24 $Y=2.17 $X2=0 $Y2=0
cc_348 N_D_c_335_n N_VPWR_c_1698_n 0.00453517f $X=2.24 $Y=2.095 $X2=0 $Y2=0
cc_349 N_D_c_334_n N_VPWR_c_1695_n 8.60012e-19 $X=2.24 $Y=2.17 $X2=0 $Y2=0
cc_350 N_D_c_329_n N_A_463_449#_c_1849_n 0.00241686f $X=2.32 $Y=1.165 $X2=0
+ $Y2=0
cc_351 N_D_c_330_n N_A_463_449#_c_1849_n 0.0137714f $X=2.395 $Y=1.09 $X2=0 $Y2=0
cc_352 N_D_c_328_n N_A_463_449#_c_1850_n 4.50256e-19 $X=1.98 $Y=2.02 $X2=0 $Y2=0
cc_353 N_D_c_335_n N_A_463_449#_c_1850_n 0.00206788f $X=2.24 $Y=2.095 $X2=0
+ $Y2=0
cc_354 N_D_c_331_n N_A_463_449#_c_1850_n 4.72213e-19 $X=1.92 $Y=1.165 $X2=0
+ $Y2=0
cc_355 N_D_c_332_n N_A_463_449#_c_1850_n 0.00361125f $X=1.92 $Y=1.345 $X2=0
+ $Y2=0
cc_356 N_D_c_334_n N_A_463_449#_c_1853_n 0.00577737f $X=2.24 $Y=2.17 $X2=0 $Y2=0
cc_357 N_D_c_329_n N_A_463_449#_c_1851_n 0.00546286f $X=2.32 $Y=1.165 $X2=0
+ $Y2=0
cc_358 N_D_c_331_n N_A_463_449#_c_1851_n 2.91775e-19 $X=1.92 $Y=1.165 $X2=0
+ $Y2=0
cc_359 N_D_c_332_n N_A_463_449#_c_1851_n 0.00547679f $X=1.92 $Y=1.345 $X2=0
+ $Y2=0
cc_360 N_D_c_330_n N_VGND_c_1977_n 0.0108538f $X=2.395 $Y=1.09 $X2=0 $Y2=0
cc_361 N_D_c_331_n N_VGND_c_1977_n 0.00479201f $X=1.92 $Y=1.165 $X2=0 $Y2=0
cc_362 N_D_c_332_n N_VGND_c_1977_n 0.0265086f $X=1.92 $Y=1.345 $X2=0 $Y2=0
cc_363 N_D_c_330_n N_VGND_c_2001_n 9.39239e-19 $X=2.395 $Y=1.09 $X2=0 $Y2=0
cc_364 N_A_113_57#_c_394_n N_A_789_78#_M1010_d 0.00377155f $X=6.51 $Y=0.35
+ $X2=-0.19 $Y2=-0.245
cc_365 N_A_113_57#_M1041_g N_A_789_78#_M1037_g 0.0199736f $X=3.45 $Y=0.73 $X2=0
+ $Y2=0
cc_366 N_A_113_57#_c_415_n N_A_789_78#_M1037_g 0.00133964f $X=3.54 $Y=1.255
+ $X2=0 $Y2=0
cc_367 N_A_113_57#_c_390_n N_A_789_78#_M1037_g 0.0179917f $X=3.54 $Y=1.255 $X2=0
+ $Y2=0
cc_368 N_A_113_57#_c_391_n N_A_789_78#_M1037_g 0.0168632f $X=4.715 $Y=1.14 $X2=0
+ $Y2=0
cc_369 N_A_113_57#_c_393_n N_A_789_78#_M1037_g 0.0043076f $X=4.8 $Y=1.055 $X2=0
+ $Y2=0
cc_370 N_A_113_57#_c_396_n N_A_789_78#_M1043_g 0.0054108f $X=6.595 $Y=1.085
+ $X2=0 $Y2=0
cc_371 N_A_113_57#_c_397_n N_A_789_78#_M1043_g 0.0157419f $X=7.335 $Y=1.17 $X2=0
+ $Y2=0
cc_372 N_A_113_57#_c_403_n N_A_789_78#_M1043_g 0.0184148f $X=7.555 $Y=1.17 $X2=0
+ $Y2=0
cc_373 N_A_113_57#_c_404_n N_A_789_78#_M1043_g 0.0209026f $X=7.61 $Y=1.51 $X2=0
+ $Y2=0
cc_374 N_A_113_57#_c_405_n N_A_789_78#_M1043_g 0.030814f $X=7.61 $Y=1.345 $X2=0
+ $Y2=0
cc_375 N_A_113_57#_c_390_n N_A_789_78#_c_643_n 0.0179917f $X=3.54 $Y=1.255 $X2=0
+ $Y2=0
cc_376 N_A_113_57#_c_398_n N_A_789_78#_c_634_n 0.00539963f $X=6.68 $Y=1.17 $X2=0
+ $Y2=0
cc_377 N_A_113_57#_c_403_n N_A_789_78#_c_636_n 0.0220473f $X=7.555 $Y=1.17 $X2=0
+ $Y2=0
cc_378 N_A_113_57#_c_404_n N_A_789_78#_c_636_n 2.54383e-19 $X=7.61 $Y=1.51 $X2=0
+ $Y2=0
cc_379 N_A_113_57#_c_397_n N_A_789_78#_c_637_n 0.0059998f $X=7.335 $Y=1.17 $X2=0
+ $Y2=0
cc_380 N_A_113_57#_c_417_n N_A_789_78#_c_637_n 0.0181191f $X=7.42 $Y=2.895 $X2=0
+ $Y2=0
cc_381 N_A_113_57#_c_397_n N_A_789_78#_c_638_n 0.0314296f $X=7.335 $Y=1.17 $X2=0
+ $Y2=0
cc_382 N_A_113_57#_c_398_n N_A_789_78#_c_638_n 0.0127556f $X=6.68 $Y=1.17 $X2=0
+ $Y2=0
cc_383 N_A_113_57#_c_391_n N_SET_B_M1017_g 0.00792239f $X=4.715 $Y=1.14 $X2=0
+ $Y2=0
cc_384 N_A_113_57#_c_393_n N_SET_B_M1017_g 0.0137959f $X=4.8 $Y=1.055 $X2=0
+ $Y2=0
cc_385 N_A_113_57#_c_394_n N_SET_B_M1017_g 0.0145373f $X=6.51 $Y=0.35 $X2=0
+ $Y2=0
cc_386 N_A_113_57#_c_420_n SET_B 0.00661053f $X=8.51 $Y=1.865 $X2=0 $Y2=0
cc_387 N_A_113_57#_c_421_n SET_B 5.75095e-19 $X=8.51 $Y=1.865 $X2=0 $Y2=0
cc_388 N_A_113_57#_c_413_n N_SET_B_c_766_n 0.00401519f $X=8.51 $Y=2.305 $X2=0
+ $Y2=0
cc_389 N_A_113_57#_c_397_n N_SET_B_c_766_n 0.00883354f $X=7.335 $Y=1.17 $X2=0
+ $Y2=0
cc_390 N_A_113_57#_c_398_n N_SET_B_c_766_n 0.00102239f $X=6.68 $Y=1.17 $X2=0
+ $Y2=0
cc_391 N_A_113_57#_c_417_n N_SET_B_c_766_n 0.0119196f $X=7.42 $Y=2.895 $X2=0
+ $Y2=0
cc_392 N_A_113_57#_c_420_n N_SET_B_c_766_n 0.0189491f $X=8.51 $Y=1.865 $X2=0
+ $Y2=0
cc_393 N_A_113_57#_c_421_n N_SET_B_c_766_n 0.00477956f $X=8.51 $Y=1.865 $X2=0
+ $Y2=0
cc_394 N_A_113_57#_c_403_n N_SET_B_c_766_n 0.030562f $X=7.555 $Y=1.17 $X2=0
+ $Y2=0
cc_395 N_A_113_57#_c_404_n N_SET_B_c_766_n 9.29903e-19 $X=7.61 $Y=1.51 $X2=0
+ $Y2=0
cc_396 N_A_113_57#_c_420_n N_SET_B_c_768_n 0.00135882f $X=8.51 $Y=1.865 $X2=0
+ $Y2=0
cc_397 N_A_113_57#_c_421_n N_SET_B_c_768_n 7.41173e-19 $X=8.51 $Y=1.865 $X2=0
+ $Y2=0
cc_398 N_A_113_57#_c_391_n N_SET_B_c_769_n 0.0021982f $X=4.715 $Y=1.14 $X2=0
+ $Y2=0
cc_399 N_A_113_57#_c_394_n N_A_549_449#_M1010_g 0.0102984f $X=6.51 $Y=0.35 $X2=0
+ $Y2=0
cc_400 N_A_113_57#_c_386_n N_A_549_449#_c_890_n 0.0047569f $X=3.375 $Y=0.18
+ $X2=0 $Y2=0
cc_401 N_A_113_57#_M1041_g N_A_549_449#_c_890_n 0.00678963f $X=3.45 $Y=0.73
+ $X2=0 $Y2=0
cc_402 N_A_113_57#_M1023_g N_A_549_449#_c_891_n 2.36136e-19 $X=2.67 $Y=2.455
+ $X2=0 $Y2=0
cc_403 N_A_113_57#_c_415_n N_A_549_449#_c_891_n 0.037026f $X=3.54 $Y=1.255 $X2=0
+ $Y2=0
cc_404 N_A_113_57#_c_390_n N_A_549_449#_c_891_n 0.00678963f $X=3.54 $Y=1.255
+ $X2=0 $Y2=0
cc_405 N_A_113_57#_c_392_n N_A_549_449#_c_891_n 0.0129662f $X=3.64 $Y=1.14 $X2=0
+ $Y2=0
cc_406 N_A_113_57#_c_415_n N_A_549_449#_c_899_n 0.00702011f $X=3.54 $Y=1.255
+ $X2=0 $Y2=0
cc_407 N_A_113_57#_c_390_n N_A_549_449#_c_899_n 0.00260653f $X=3.54 $Y=1.255
+ $X2=0 $Y2=0
cc_408 N_A_113_57#_c_415_n N_A_549_449#_c_892_n 0.0127902f $X=3.54 $Y=1.255
+ $X2=0 $Y2=0
cc_409 N_A_113_57#_c_390_n N_A_549_449#_c_892_n 0.00119377f $X=3.54 $Y=1.255
+ $X2=0 $Y2=0
cc_410 N_A_113_57#_c_391_n N_A_549_449#_c_893_n 0.0534343f $X=4.715 $Y=1.14
+ $X2=0 $Y2=0
cc_411 N_A_113_57#_c_415_n N_A_549_449#_c_894_n 0.0132787f $X=3.54 $Y=1.255
+ $X2=0 $Y2=0
cc_412 N_A_113_57#_c_390_n N_A_549_449#_c_894_n 0.00127177f $X=3.54 $Y=1.255
+ $X2=0 $Y2=0
cc_413 N_A_113_57#_c_391_n N_A_549_449#_c_894_n 0.0134116f $X=4.715 $Y=1.14
+ $X2=0 $Y2=0
cc_414 N_A_113_57#_c_390_n N_A_549_449#_c_921_n 0.00678963f $X=3.54 $Y=1.255
+ $X2=0 $Y2=0
cc_415 N_A_113_57#_M1023_g N_A_549_449#_c_905_n 0.00281161f $X=2.67 $Y=2.455
+ $X2=0 $Y2=0
cc_416 N_A_113_57#_c_390_n N_A_549_449#_c_905_n 2.20559e-19 $X=3.54 $Y=1.255
+ $X2=0 $Y2=0
cc_417 N_A_113_57#_c_386_n N_A_223_119#_M1013_g 0.0103003f $X=3.375 $Y=0.18
+ $X2=0 $Y2=0
cc_418 N_A_113_57#_M1041_g N_A_223_119#_M1013_g 0.0107747f $X=3.45 $Y=0.73 $X2=0
+ $Y2=0
cc_419 N_A_113_57#_c_415_n N_A_223_119#_c_1039_n 4.95434e-19 $X=3.54 $Y=1.255
+ $X2=0 $Y2=0
cc_420 N_A_113_57#_c_390_n N_A_223_119#_c_1039_n 0.010277f $X=3.54 $Y=1.255
+ $X2=0 $Y2=0
cc_421 N_A_113_57#_M1023_g N_A_223_119#_c_1040_n 0.00188478f $X=2.67 $Y=2.455
+ $X2=0 $Y2=0
cc_422 N_A_113_57#_M1023_g N_A_223_119#_M1030_g 0.00730422f $X=2.67 $Y=2.455
+ $X2=0 $Y2=0
cc_423 N_A_113_57#_c_412_n N_A_223_119#_c_1042_n 0.0100806f $X=8.145 $Y=2.455
+ $X2=0 $Y2=0
cc_424 N_A_113_57#_c_419_n N_A_223_119#_c_1042_n 0.00332103f $X=7.505 $Y=2.98
+ $X2=0 $Y2=0
cc_425 N_A_113_57#_c_409_n N_A_223_119#_c_1043_n 0.00730422f $X=2.595 $Y=3.08
+ $X2=0 $Y2=0
cc_426 N_A_113_57#_c_413_n N_A_223_119#_M1020_g 0.0100806f $X=8.51 $Y=2.305
+ $X2=0 $Y2=0
cc_427 N_A_113_57#_c_418_n N_A_223_119#_M1020_g 0.0151989f $X=8.345 $Y=2.98
+ $X2=0 $Y2=0
cc_428 N_A_113_57#_c_421_n N_A_223_119#_M1020_g 0.00228806f $X=8.51 $Y=1.865
+ $X2=0 $Y2=0
cc_429 N_A_113_57#_c_413_n N_A_223_119#_c_1045_n 0.00379301f $X=8.51 $Y=2.305
+ $X2=0 $Y2=0
cc_430 N_A_113_57#_c_417_n N_A_223_119#_c_1046_n 0.00676641f $X=7.42 $Y=2.895
+ $X2=0 $Y2=0
cc_431 N_A_113_57#_c_403_n N_A_223_119#_c_1046_n 0.00206075f $X=7.555 $Y=1.17
+ $X2=0 $Y2=0
cc_432 N_A_113_57#_c_404_n N_A_223_119#_c_1046_n 0.0117925f $X=7.61 $Y=1.51
+ $X2=0 $Y2=0
cc_433 N_A_113_57#_c_417_n N_A_223_119#_c_1029_n 0.00122494f $X=7.42 $Y=2.895
+ $X2=0 $Y2=0
cc_434 N_A_113_57#_c_420_n N_A_223_119#_c_1029_n 0.00124311f $X=8.51 $Y=1.865
+ $X2=0 $Y2=0
cc_435 N_A_113_57#_c_421_n N_A_223_119#_c_1029_n 0.0223548f $X=8.51 $Y=1.865
+ $X2=0 $Y2=0
cc_436 N_A_113_57#_c_420_n N_A_223_119#_c_1030_n 8.68446e-19 $X=8.51 $Y=1.865
+ $X2=0 $Y2=0
cc_437 N_A_113_57#_c_421_n N_A_223_119#_c_1030_n 0.00825601f $X=8.51 $Y=1.865
+ $X2=0 $Y2=0
cc_438 N_A_113_57#_c_403_n N_A_223_119#_c_1031_n 5.59496e-19 $X=7.555 $Y=1.17
+ $X2=0 $Y2=0
cc_439 N_A_113_57#_c_404_n N_A_223_119#_c_1031_n 0.0210121f $X=7.61 $Y=1.51
+ $X2=0 $Y2=0
cc_440 N_A_113_57#_c_405_n N_A_223_119#_c_1031_n 0.0018943f $X=7.61 $Y=1.345
+ $X2=0 $Y2=0
cc_441 N_A_113_57#_c_403_n N_A_223_119#_c_1032_n 2.06829e-19 $X=7.555 $Y=1.17
+ $X2=0 $Y2=0
cc_442 N_A_113_57#_c_405_n N_A_223_119#_c_1032_n 0.00747575f $X=7.61 $Y=1.345
+ $X2=0 $Y2=0
cc_443 N_A_113_57#_M1023_g N_A_223_119#_c_1033_n 0.00762016f $X=2.67 $Y=2.455
+ $X2=0 $Y2=0
cc_444 N_A_113_57#_c_390_n N_A_223_119#_c_1034_n 0.0160225f $X=3.54 $Y=1.255
+ $X2=0 $Y2=0
cc_445 N_A_113_57#_c_383_n N_A_223_119#_c_1035_n 0.0125499f $X=1.395 $Y=1.375
+ $X2=0 $Y2=0
cc_446 N_A_113_57#_c_406_n N_A_223_119#_c_1035_n 0.00510473f $X=1.515 $Y=1.895
+ $X2=0 $Y2=0
cc_447 N_A_113_57#_M1002_g N_A_223_119#_c_1035_n 0.00976283f $X=1.47 $Y=0.805
+ $X2=0 $Y2=0
cc_448 N_A_113_57#_c_400_n N_A_223_119#_c_1035_n 0.0368496f $X=0.84 $Y=1.465
+ $X2=0 $Y2=0
cc_449 N_A_113_57#_c_401_n N_A_223_119#_c_1035_n 0.00416296f $X=0.84 $Y=1.465
+ $X2=0 $Y2=0
cc_450 N_A_113_57#_c_402_n N_A_223_119#_c_1035_n 0.0141955f $X=0.827 $Y=1.3
+ $X2=0 $Y2=0
cc_451 N_A_113_57#_M1035_g N_A_223_119#_c_1051_n 0.0154003f $X=1.59 $Y=2.565
+ $X2=0 $Y2=0
cc_452 N_A_113_57#_c_389_n N_A_223_119#_c_1051_n 0.0631119f $X=0.815 $Y=2.55
+ $X2=0 $Y2=0
cc_453 N_A_113_57#_c_406_n N_A_223_119#_c_1052_n 0.00398066f $X=1.515 $Y=1.895
+ $X2=0 $Y2=0
cc_454 N_A_113_57#_M1035_g N_A_223_119#_c_1052_n 0.00707993f $X=1.59 $Y=2.565
+ $X2=0 $Y2=0
cc_455 N_A_113_57#_c_383_n N_A_223_119#_c_1037_n 0.00397348f $X=1.395 $Y=1.375
+ $X2=0 $Y2=0
cc_456 N_A_113_57#_M1002_g N_A_223_119#_c_1037_n 0.00703355f $X=1.47 $Y=0.805
+ $X2=0 $Y2=0
cc_457 N_A_113_57#_c_399_n N_A_223_119#_c_1037_n 0.0289462f $X=0.705 $Y=0.495
+ $X2=0 $Y2=0
cc_458 N_A_113_57#_c_383_n N_A_223_119#_c_1054_n 0.00100297f $X=1.395 $Y=1.375
+ $X2=0 $Y2=0
cc_459 N_A_113_57#_c_406_n N_A_223_119#_c_1054_n 0.0145571f $X=1.515 $Y=1.895
+ $X2=0 $Y2=0
cc_460 N_A_113_57#_M1035_g N_A_223_119#_c_1054_n 0.00166926f $X=1.59 $Y=2.565
+ $X2=0 $Y2=0
cc_461 N_A_113_57#_c_389_n N_A_223_119#_c_1054_n 0.0124018f $X=0.815 $Y=2.55
+ $X2=0 $Y2=0
cc_462 N_A_113_57#_c_412_n N_A_1746_137#_M1021_g 0.00590258f $X=8.145 $Y=2.455
+ $X2=0 $Y2=0
cc_463 N_A_113_57#_c_413_n N_A_1746_137#_M1021_g 0.00504495f $X=8.51 $Y=2.305
+ $X2=0 $Y2=0
cc_464 N_A_113_57#_c_418_n N_A_1746_137#_M1021_g 0.00454173f $X=8.345 $Y=2.98
+ $X2=0 $Y2=0
cc_465 N_A_113_57#_c_420_n N_A_1746_137#_M1021_g 0.0103367f $X=8.51 $Y=1.865
+ $X2=0 $Y2=0
cc_466 N_A_113_57#_c_420_n N_A_1746_137#_c_1221_n 0.0168274f $X=8.51 $Y=1.865
+ $X2=0 $Y2=0
cc_467 N_A_113_57#_c_421_n N_A_1746_137#_c_1221_n 0.00122747f $X=8.51 $Y=1.865
+ $X2=0 $Y2=0
cc_468 N_A_113_57#_c_413_n N_A_1746_137#_c_1222_n 0.0212003f $X=8.51 $Y=2.305
+ $X2=0 $Y2=0
cc_469 N_A_113_57#_c_420_n N_A_1746_137#_c_1210_n 0.00255717f $X=8.51 $Y=1.865
+ $X2=0 $Y2=0
cc_470 N_A_113_57#_c_421_n N_A_1746_137#_c_1210_n 0.0212003f $X=8.51 $Y=1.865
+ $X2=0 $Y2=0
cc_471 N_A_113_57#_c_418_n N_A_1542_428#_M1020_d 0.00267852f $X=8.345 $Y=2.98
+ $X2=0 $Y2=0
cc_472 N_A_113_57#_c_405_n N_A_1542_428#_c_1376_n 0.0141349f $X=7.61 $Y=1.345
+ $X2=0 $Y2=0
cc_473 N_A_113_57#_c_420_n N_A_1542_428#_c_1377_n 0.00576025f $X=8.51 $Y=1.865
+ $X2=0 $Y2=0
cc_474 N_A_113_57#_c_421_n N_A_1542_428#_c_1377_n 0.00232851f $X=8.51 $Y=1.865
+ $X2=0 $Y2=0
cc_475 N_A_113_57#_c_412_n N_A_1542_428#_c_1384_n 0.00812282f $X=8.145 $Y=2.455
+ $X2=0 $Y2=0
cc_476 N_A_113_57#_c_413_n N_A_1542_428#_c_1384_n 0.0059583f $X=8.51 $Y=2.305
+ $X2=0 $Y2=0
cc_477 N_A_113_57#_c_417_n N_A_1542_428#_c_1384_n 0.0229716f $X=7.42 $Y=2.895
+ $X2=0 $Y2=0
cc_478 N_A_113_57#_c_418_n N_A_1542_428#_c_1384_n 0.0229954f $X=8.345 $Y=2.98
+ $X2=0 $Y2=0
cc_479 N_A_113_57#_c_403_n N_A_1542_428#_c_1384_n 0.00198059f $X=7.555 $Y=1.17
+ $X2=0 $Y2=0
cc_480 N_A_113_57#_c_417_n N_A_1542_428#_c_1378_n 0.0156917f $X=7.42 $Y=2.895
+ $X2=0 $Y2=0
cc_481 N_A_113_57#_c_420_n N_A_1542_428#_c_1378_n 0.0618901f $X=8.51 $Y=1.865
+ $X2=0 $Y2=0
cc_482 N_A_113_57#_c_421_n N_A_1542_428#_c_1378_n 0.0037009f $X=8.51 $Y=1.865
+ $X2=0 $Y2=0
cc_483 N_A_113_57#_c_403_n N_A_1542_428#_c_1378_n 0.0277695f $X=7.555 $Y=1.17
+ $X2=0 $Y2=0
cc_484 N_A_113_57#_c_404_n N_A_1542_428#_c_1378_n 0.00163913f $X=7.61 $Y=1.51
+ $X2=0 $Y2=0
cc_485 N_A_113_57#_c_403_n N_A_1542_428#_c_1379_n 0.00967259f $X=7.555 $Y=1.17
+ $X2=0 $Y2=0
cc_486 N_A_113_57#_c_405_n N_A_1542_428#_c_1379_n 7.75352e-19 $X=7.61 $Y=1.345
+ $X2=0 $Y2=0
cc_487 N_A_113_57#_c_394_n N_A_1191_21#_M1003_g 0.0124247f $X=6.51 $Y=0.35 $X2=0
+ $Y2=0
cc_488 N_A_113_57#_c_396_n N_A_1191_21#_M1003_g 0.00728312f $X=6.595 $Y=1.085
+ $X2=0 $Y2=0
cc_489 N_A_113_57#_c_398_n N_A_1191_21#_M1003_g 0.00310437f $X=6.68 $Y=1.17
+ $X2=0 $Y2=0
cc_490 N_A_113_57#_c_394_n N_A_1191_21#_c_1472_n 0.0115412f $X=6.51 $Y=0.35
+ $X2=0 $Y2=0
cc_491 N_A_113_57#_c_405_n N_A_1191_21#_c_1472_n 0.0104164f $X=7.61 $Y=1.345
+ $X2=0 $Y2=0
cc_492 N_A_113_57#_c_389_n N_VPWR_c_1697_n 0.0261645f $X=0.815 $Y=2.55 $X2=0
+ $Y2=0
cc_493 N_A_113_57#_M1035_g N_VPWR_c_1698_n 0.0103306f $X=1.59 $Y=2.565 $X2=0
+ $Y2=0
cc_494 N_A_113_57#_c_409_n N_VPWR_c_1698_n 0.0284081f $X=2.595 $Y=3.08 $X2=0
+ $Y2=0
cc_495 N_A_113_57#_M1023_g N_VPWR_c_1698_n 0.00544232f $X=2.67 $Y=2.455 $X2=0
+ $Y2=0
cc_496 N_A_113_57#_c_410_n N_VPWR_c_1708_n 0.00675559f $X=1.665 $Y=3.08 $X2=0
+ $Y2=0
cc_497 N_A_113_57#_c_389_n N_VPWR_c_1708_n 0.0237177f $X=0.815 $Y=2.55 $X2=0
+ $Y2=0
cc_498 N_A_113_57#_c_409_n N_VPWR_c_1710_n 0.0192298f $X=2.595 $Y=3.08 $X2=0
+ $Y2=0
cc_499 N_A_113_57#_c_412_n N_VPWR_c_1713_n 0.00392127f $X=8.145 $Y=2.455 $X2=0
+ $Y2=0
cc_500 N_A_113_57#_c_418_n N_VPWR_c_1713_n 0.0682237f $X=8.345 $Y=2.98 $X2=0
+ $Y2=0
cc_501 N_A_113_57#_c_419_n N_VPWR_c_1713_n 0.0114245f $X=7.505 $Y=2.98 $X2=0
+ $Y2=0
cc_502 N_A_113_57#_c_409_n N_VPWR_c_1695_n 0.0278029f $X=2.595 $Y=3.08 $X2=0
+ $Y2=0
cc_503 N_A_113_57#_c_410_n N_VPWR_c_1695_n 0.00953141f $X=1.665 $Y=3.08 $X2=0
+ $Y2=0
cc_504 N_A_113_57#_c_412_n N_VPWR_c_1695_n 0.00542671f $X=8.145 $Y=2.455 $X2=0
+ $Y2=0
cc_505 N_A_113_57#_c_413_n N_VPWR_c_1695_n 0.00153096f $X=8.51 $Y=2.305 $X2=0
+ $Y2=0
cc_506 N_A_113_57#_c_389_n N_VPWR_c_1695_n 0.0135481f $X=0.815 $Y=2.55 $X2=0
+ $Y2=0
cc_507 N_A_113_57#_c_418_n N_VPWR_c_1695_n 0.0408085f $X=8.345 $Y=2.98 $X2=0
+ $Y2=0
cc_508 N_A_113_57#_c_419_n N_VPWR_c_1695_n 0.00589433f $X=7.505 $Y=2.98 $X2=0
+ $Y2=0
cc_509 N_A_113_57#_c_386_n N_A_463_449#_c_1849_n 0.00582439f $X=3.375 $Y=0.18
+ $X2=0 $Y2=0
cc_510 N_A_113_57#_M1023_g N_A_463_449#_c_1850_n 0.0045615f $X=2.67 $Y=2.455
+ $X2=0 $Y2=0
cc_511 N_A_113_57#_c_409_n N_A_463_449#_c_1853_n 0.00389513f $X=2.595 $Y=3.08
+ $X2=0 $Y2=0
cc_512 N_A_113_57#_M1023_g N_A_463_449#_c_1853_n 0.014848f $X=2.67 $Y=2.455
+ $X2=0 $Y2=0
cc_513 N_A_113_57#_c_417_n A_1447_379# 0.0197069f $X=7.42 $Y=2.895 $X2=-0.19
+ $Y2=-0.245
cc_514 N_A_113_57#_c_419_n A_1447_379# 0.00404611f $X=7.505 $Y=2.98 $X2=-0.19
+ $Y2=-0.245
cc_515 N_A_113_57#_c_418_n A_1644_506# 0.00246829f $X=8.345 $Y=2.98 $X2=-0.19
+ $Y2=-0.245
cc_516 N_A_113_57#_c_420_n A_1644_506# 0.0121105f $X=8.51 $Y=1.865 $X2=-0.19
+ $Y2=-0.245
cc_517 N_A_113_57#_c_393_n N_VGND_M1037_d 0.00895164f $X=4.8 $Y=1.055 $X2=0
+ $Y2=0
cc_518 N_A_113_57#_c_395_n N_VGND_M1037_d 0.00182835f $X=4.885 $Y=0.35 $X2=0
+ $Y2=0
cc_519 N_A_113_57#_c_397_n N_VGND_M1043_s 0.00501179f $X=7.335 $Y=1.17 $X2=0
+ $Y2=0
cc_520 N_A_113_57#_c_399_n N_VGND_c_1976_n 0.0179429f $X=0.705 $Y=0.495 $X2=0
+ $Y2=0
cc_521 N_A_113_57#_M1002_g N_VGND_c_1977_n 0.0216434f $X=1.47 $Y=0.805 $X2=0
+ $Y2=0
cc_522 N_A_113_57#_c_386_n N_VGND_c_1977_n 0.0248025f $X=3.375 $Y=0.18 $X2=0
+ $Y2=0
cc_523 N_A_113_57#_c_386_n N_VGND_c_1978_n 0.00594862f $X=3.375 $Y=0.18 $X2=0
+ $Y2=0
cc_524 N_A_113_57#_c_391_n N_VGND_c_1978_n 0.0260135f $X=4.715 $Y=1.14 $X2=0
+ $Y2=0
cc_525 N_A_113_57#_c_393_n N_VGND_c_1978_n 0.0321918f $X=4.8 $Y=1.055 $X2=0
+ $Y2=0
cc_526 N_A_113_57#_c_395_n N_VGND_c_1978_n 0.013989f $X=4.885 $Y=0.35 $X2=0
+ $Y2=0
cc_527 N_A_113_57#_c_394_n N_VGND_c_1979_n 0.0141601f $X=6.51 $Y=0.35 $X2=0
+ $Y2=0
cc_528 N_A_113_57#_c_396_n N_VGND_c_1979_n 0.0345265f $X=6.595 $Y=1.085 $X2=0
+ $Y2=0
cc_529 N_A_113_57#_c_397_n N_VGND_c_1979_n 0.0147238f $X=7.335 $Y=1.17 $X2=0
+ $Y2=0
cc_530 N_A_113_57#_c_405_n N_VGND_c_1979_n 0.00207662f $X=7.61 $Y=1.345 $X2=0
+ $Y2=0
cc_531 N_A_113_57#_c_386_n N_VGND_c_1986_n 0.0507481f $X=3.375 $Y=0.18 $X2=0
+ $Y2=0
cc_532 N_A_113_57#_c_387_n N_VGND_c_1988_n 0.00768994f $X=1.545 $Y=0.18 $X2=0
+ $Y2=0
cc_533 N_A_113_57#_c_399_n N_VGND_c_1988_n 0.0218253f $X=0.705 $Y=0.495 $X2=0
+ $Y2=0
cc_534 N_A_113_57#_c_394_n N_VGND_c_1989_n 0.108638f $X=6.51 $Y=0.35 $X2=0 $Y2=0
cc_535 N_A_113_57#_c_395_n N_VGND_c_1989_n 0.0114622f $X=4.885 $Y=0.35 $X2=0
+ $Y2=0
cc_536 N_A_113_57#_c_386_n N_VGND_c_2001_n 0.0725353f $X=3.375 $Y=0.18 $X2=0
+ $Y2=0
cc_537 N_A_113_57#_c_387_n N_VGND_c_2001_n 0.0106678f $X=1.545 $Y=0.18 $X2=0
+ $Y2=0
cc_538 N_A_113_57#_c_394_n N_VGND_c_2001_n 0.0629179f $X=6.51 $Y=0.35 $X2=0
+ $Y2=0
cc_539 N_A_113_57#_c_395_n N_VGND_c_2001_n 0.00657784f $X=4.885 $Y=0.35 $X2=0
+ $Y2=0
cc_540 N_A_113_57#_c_399_n N_VGND_c_2001_n 0.0125375f $X=0.705 $Y=0.495 $X2=0
+ $Y2=0
cc_541 N_A_113_57#_c_405_n N_VGND_c_2001_n 9.39239e-19 $X=7.61 $Y=1.345 $X2=0
+ $Y2=0
cc_542 N_A_113_57#_c_394_n N_A_1018_60#_M1017_d 0.00186629f $X=6.51 $Y=0.35
+ $X2=-0.19 $Y2=-0.245
cc_543 N_A_113_57#_c_393_n N_A_1018_60#_c_2124_n 0.0137213f $X=4.8 $Y=1.055
+ $X2=0 $Y2=0
cc_544 N_A_113_57#_c_394_n N_A_1018_60#_c_2124_n 0.0597876f $X=6.51 $Y=0.35
+ $X2=0 $Y2=0
cc_545 N_A_113_57#_c_394_n N_A_1018_60#_c_2125_n 0.0120137f $X=6.51 $Y=0.35
+ $X2=0 $Y2=0
cc_546 N_A_113_57#_c_396_n N_A_1018_60#_c_2125_n 0.0234464f $X=6.595 $Y=1.085
+ $X2=0 $Y2=0
cc_547 N_A_113_57#_c_397_n A_1447_119# 0.00201179f $X=7.335 $Y=1.17 $X2=-0.19
+ $Y2=-0.245
cc_548 N_A_113_57#_c_403_n A_1447_119# 0.00944092f $X=7.555 $Y=1.17 $X2=-0.19
+ $Y2=-0.245
cc_549 N_A_789_78#_c_642_n N_SET_B_M1024_g 0.00408644f $X=4.27 $Y=1.92 $X2=0
+ $Y2=0
cc_550 N_A_789_78#_c_643_n N_SET_B_M1024_g 0.00449738f $X=4.27 $Y=1.92 $X2=0
+ $Y2=0
cc_551 N_A_789_78#_c_669_p N_SET_B_M1024_g 0.00902665f $X=5.14 $Y=2.532 $X2=0
+ $Y2=0
cc_552 N_A_789_78#_c_645_n N_SET_B_M1024_g 0.0105234f $X=5.47 $Y=2.532 $X2=0
+ $Y2=0
cc_553 N_A_789_78#_c_671_p N_SET_B_c_766_n 0.00556066f $X=5.885 $Y=2.395 $X2=0
+ $Y2=0
cc_554 N_A_789_78#_c_644_n N_SET_B_c_766_n 0.0162125f $X=5.97 $Y=2.31 $X2=0
+ $Y2=0
cc_555 N_A_789_78#_c_645_n N_SET_B_c_766_n 0.00114414f $X=5.47 $Y=2.532 $X2=0
+ $Y2=0
cc_556 N_A_789_78#_c_634_n N_SET_B_c_766_n 0.00851884f $X=5.74 $Y=1.13 $X2=0
+ $Y2=0
cc_557 N_A_789_78#_c_635_n N_SET_B_c_766_n 0.00868974f $X=5.97 $Y=1.52 $X2=0
+ $Y2=0
cc_558 N_A_789_78#_c_636_n N_SET_B_c_766_n 0.0190576f $X=6.99 $Y=1.57 $X2=0
+ $Y2=0
cc_559 N_A_789_78#_c_637_n N_SET_B_c_766_n 0.0122447f $X=6.99 $Y=1.57 $X2=0
+ $Y2=0
cc_560 N_A_789_78#_c_638_n N_SET_B_c_766_n 0.0388725f $X=6.825 $Y=1.585 $X2=0
+ $Y2=0
cc_561 N_A_789_78#_c_633_n N_A_549_449#_M1010_g 0.00191797f $X=5.97 $Y=1.435
+ $X2=0 $Y2=0
cc_562 N_A_789_78#_c_634_n N_A_549_449#_M1010_g 0.00999403f $X=5.74 $Y=1.13
+ $X2=0 $Y2=0
cc_563 N_A_789_78#_c_671_p N_A_549_449#_M1040_g 0.00736475f $X=5.885 $Y=2.395
+ $X2=0 $Y2=0
cc_564 N_A_789_78#_c_644_n N_A_549_449#_M1040_g 0.00436666f $X=5.97 $Y=2.31
+ $X2=0 $Y2=0
cc_565 N_A_789_78#_c_645_n N_A_549_449#_M1040_g 0.00705291f $X=5.47 $Y=2.532
+ $X2=0 $Y2=0
cc_566 N_A_789_78#_c_643_n N_A_549_449#_c_891_n 0.0011387f $X=4.27 $Y=1.92 $X2=0
+ $Y2=0
cc_567 N_A_789_78#_M1039_g N_A_549_449#_c_899_n 0.00574363f $X=4.02 $Y=2.455
+ $X2=0 $Y2=0
cc_568 N_A_789_78#_c_642_n N_A_549_449#_c_899_n 0.00645469f $X=4.27 $Y=1.92
+ $X2=0 $Y2=0
cc_569 N_A_789_78#_c_687_p N_A_549_449#_c_899_n 0.00710479f $X=4.37 $Y=2.395
+ $X2=0 $Y2=0
cc_570 N_A_789_78#_M1037_g N_A_549_449#_c_892_n 0.00487622f $X=4.02 $Y=0.73
+ $X2=0 $Y2=0
cc_571 N_A_789_78#_M1039_g N_A_549_449#_c_892_n 0.00298185f $X=4.02 $Y=2.455
+ $X2=0 $Y2=0
cc_572 N_A_789_78#_c_642_n N_A_549_449#_c_892_n 0.0312888f $X=4.27 $Y=1.92 $X2=0
+ $Y2=0
cc_573 N_A_789_78#_c_643_n N_A_549_449#_c_892_n 0.0108641f $X=4.27 $Y=1.92 $X2=0
+ $Y2=0
cc_574 N_A_789_78#_M1037_g N_A_549_449#_c_893_n 0.0116457f $X=4.02 $Y=0.73 $X2=0
+ $Y2=0
cc_575 N_A_789_78#_c_642_n N_A_549_449#_c_893_n 0.01515f $X=4.27 $Y=1.92 $X2=0
+ $Y2=0
cc_576 N_A_789_78#_c_643_n N_A_549_449#_c_893_n 0.00665566f $X=4.27 $Y=1.92
+ $X2=0 $Y2=0
cc_577 N_A_789_78#_M1037_g N_A_549_449#_c_894_n 0.00238028f $X=4.02 $Y=0.73
+ $X2=0 $Y2=0
cc_578 N_A_789_78#_M1037_g N_A_549_449#_c_895_n 0.00291229f $X=4.02 $Y=0.73
+ $X2=0 $Y2=0
cc_579 N_A_789_78#_c_642_n N_A_549_449#_c_895_n 0.0141145f $X=4.27 $Y=1.92 $X2=0
+ $Y2=0
cc_580 N_A_789_78#_c_643_n N_A_549_449#_c_895_n 0.00236957f $X=4.27 $Y=1.92
+ $X2=0 $Y2=0
cc_581 N_A_789_78#_M1024_d N_A_549_449#_c_944_n 0.00387952f $X=5.165 $Y=1.895
+ $X2=0 $Y2=0
cc_582 N_A_789_78#_c_644_n N_A_549_449#_c_944_n 0.0132518f $X=5.97 $Y=2.31 $X2=0
+ $Y2=0
cc_583 N_A_789_78#_c_669_p N_A_549_449#_c_944_n 0.0367981f $X=5.14 $Y=2.532
+ $X2=0 $Y2=0
cc_584 N_A_789_78#_c_645_n N_A_549_449#_c_944_n 0.0156317f $X=5.47 $Y=2.532
+ $X2=0 $Y2=0
cc_585 N_A_789_78#_c_642_n N_A_549_449#_c_902_n 0.0134543f $X=4.27 $Y=1.92 $X2=0
+ $Y2=0
cc_586 N_A_789_78#_c_643_n N_A_549_449#_c_902_n 0.00157436f $X=4.27 $Y=1.92
+ $X2=0 $Y2=0
cc_587 N_A_789_78#_c_669_p N_A_549_449#_c_902_n 0.0133439f $X=5.14 $Y=2.532
+ $X2=0 $Y2=0
cc_588 N_A_789_78#_M1024_d N_A_549_449#_c_903_n 9.03792e-19 $X=5.165 $Y=1.895
+ $X2=0 $Y2=0
cc_589 N_A_789_78#_c_644_n N_A_549_449#_c_903_n 0.0251821f $X=5.97 $Y=2.31 $X2=0
+ $Y2=0
cc_590 N_A_789_78#_c_634_n N_A_549_449#_c_903_n 0.009602f $X=5.74 $Y=1.13 $X2=0
+ $Y2=0
cc_591 N_A_789_78#_c_635_n N_A_549_449#_c_903_n 0.0103517f $X=5.97 $Y=1.52 $X2=0
+ $Y2=0
cc_592 N_A_789_78#_c_671_p N_A_549_449#_c_896_n 2.76184e-19 $X=5.885 $Y=2.395
+ $X2=0 $Y2=0
cc_593 N_A_789_78#_c_633_n N_A_549_449#_c_896_n 6.03658e-19 $X=5.97 $Y=1.435
+ $X2=0 $Y2=0
cc_594 N_A_789_78#_c_644_n N_A_549_449#_c_896_n 5.6361e-19 $X=5.97 $Y=2.31 $X2=0
+ $Y2=0
cc_595 N_A_789_78#_c_634_n N_A_549_449#_c_896_n 0.00330499f $X=5.74 $Y=1.13
+ $X2=0 $Y2=0
cc_596 N_A_789_78#_c_635_n N_A_549_449#_c_896_n 0.00194982f $X=5.97 $Y=1.52
+ $X2=0 $Y2=0
cc_597 N_A_789_78#_M1039_g N_A_549_449#_c_905_n 0.00133465f $X=4.02 $Y=2.455
+ $X2=0 $Y2=0
cc_598 N_A_789_78#_c_643_n N_A_223_119#_c_1039_n 0.0117935f $X=4.27 $Y=1.92
+ $X2=0 $Y2=0
cc_599 N_A_789_78#_M1039_g N_A_223_119#_M1030_g 0.0117935f $X=4.02 $Y=2.455
+ $X2=0 $Y2=0
cc_600 N_A_789_78#_M1039_g N_A_223_119#_c_1042_n 0.00760304f $X=4.02 $Y=2.455
+ $X2=0 $Y2=0
cc_601 N_A_789_78#_M1005_g N_A_223_119#_c_1042_n 0.0104164f $X=7.16 $Y=2.315
+ $X2=0 $Y2=0
cc_602 N_A_789_78#_c_687_p N_A_223_119#_c_1042_n 0.00525608f $X=4.37 $Y=2.395
+ $X2=0 $Y2=0
cc_603 N_A_789_78#_c_671_p N_A_223_119#_c_1042_n 0.00739236f $X=5.885 $Y=2.395
+ $X2=0 $Y2=0
cc_604 N_A_789_78#_c_669_p N_A_223_119#_c_1042_n 0.00712962f $X=5.14 $Y=2.532
+ $X2=0 $Y2=0
cc_605 N_A_789_78#_c_645_n N_A_223_119#_c_1042_n 0.00565192f $X=5.47 $Y=2.532
+ $X2=0 $Y2=0
cc_606 N_A_789_78#_M1005_g N_A_223_119#_c_1046_n 0.0273224f $X=7.16 $Y=2.315
+ $X2=0 $Y2=0
cc_607 N_A_789_78#_c_671_p N_A_1191_21#_M1003_g 0.00634225f $X=5.885 $Y=2.395
+ $X2=0 $Y2=0
cc_608 N_A_789_78#_c_633_n N_A_1191_21#_M1003_g 0.00743398f $X=5.97 $Y=1.435
+ $X2=0 $Y2=0
cc_609 N_A_789_78#_c_644_n N_A_1191_21#_M1003_g 0.0214666f $X=5.97 $Y=2.31 $X2=0
+ $Y2=0
cc_610 N_A_789_78#_c_645_n N_A_1191_21#_M1003_g 0.0012908f $X=5.47 $Y=2.532
+ $X2=0 $Y2=0
cc_611 N_A_789_78#_c_634_n N_A_1191_21#_M1003_g 0.00963959f $X=5.74 $Y=1.13
+ $X2=0 $Y2=0
cc_612 N_A_789_78#_c_635_n N_A_1191_21#_M1003_g 0.00236416f $X=5.97 $Y=1.52
+ $X2=0 $Y2=0
cc_613 N_A_789_78#_c_637_n N_A_1191_21#_M1003_g 0.00376099f $X=6.99 $Y=1.57
+ $X2=0 $Y2=0
cc_614 N_A_789_78#_c_638_n N_A_1191_21#_M1003_g 0.00685627f $X=6.825 $Y=1.585
+ $X2=0 $Y2=0
cc_615 N_A_789_78#_M1043_g N_A_1191_21#_c_1472_n 0.0103107f $X=7.16 $Y=0.915
+ $X2=0 $Y2=0
cc_616 N_A_789_78#_c_642_n N_VPWR_M1039_d 0.00215169f $X=4.27 $Y=1.92 $X2=0
+ $Y2=0
cc_617 N_A_789_78#_c_687_p N_VPWR_M1039_d 0.00579347f $X=4.37 $Y=2.395 $X2=0
+ $Y2=0
cc_618 N_A_789_78#_c_669_p N_VPWR_M1039_d 0.0192874f $X=5.14 $Y=2.532 $X2=0
+ $Y2=0
cc_619 N_A_789_78#_M1039_g N_VPWR_c_1699_n 0.00341996f $X=4.02 $Y=2.455 $X2=0
+ $Y2=0
cc_620 N_A_789_78#_c_669_p N_VPWR_c_1699_n 0.0248544f $X=5.14 $Y=2.532 $X2=0
+ $Y2=0
cc_621 N_A_789_78#_c_645_n N_VPWR_c_1699_n 0.00410938f $X=5.47 $Y=2.532 $X2=0
+ $Y2=0
cc_622 N_A_789_78#_M1005_g N_VPWR_c_1700_n 0.025462f $X=7.16 $Y=2.315 $X2=0
+ $Y2=0
cc_623 N_A_789_78#_c_671_p N_VPWR_c_1700_n 0.0133993f $X=5.885 $Y=2.395 $X2=0
+ $Y2=0
cc_624 N_A_789_78#_c_644_n N_VPWR_c_1700_n 0.0307988f $X=5.97 $Y=2.31 $X2=0
+ $Y2=0
cc_625 N_A_789_78#_c_638_n N_VPWR_c_1700_n 0.014464f $X=6.825 $Y=1.585 $X2=0
+ $Y2=0
cc_626 N_A_789_78#_c_645_n N_VPWR_c_1712_n 0.00722409f $X=5.47 $Y=2.532 $X2=0
+ $Y2=0
cc_627 N_A_789_78#_M1039_g N_VPWR_c_1695_n 9.6081e-19 $X=4.02 $Y=2.455 $X2=0
+ $Y2=0
cc_628 N_A_789_78#_M1005_g N_VPWR_c_1695_n 9.39239e-19 $X=7.16 $Y=2.315 $X2=0
+ $Y2=0
cc_629 N_A_789_78#_c_687_p N_VPWR_c_1695_n 0.00702095f $X=4.37 $Y=2.395 $X2=0
+ $Y2=0
cc_630 N_A_789_78#_c_671_p N_VPWR_c_1695_n 0.0177904f $X=5.885 $Y=2.395 $X2=0
+ $Y2=0
cc_631 N_A_789_78#_c_669_p N_VPWR_c_1695_n 0.0140835f $X=5.14 $Y=2.532 $X2=0
+ $Y2=0
cc_632 N_A_789_78#_c_645_n N_VPWR_c_1695_n 0.0088922f $X=5.47 $Y=2.532 $X2=0
+ $Y2=0
cc_633 N_A_789_78#_c_671_p A_1119_379# 0.0062271f $X=5.885 $Y=2.395 $X2=-0.19
+ $Y2=-0.245
cc_634 N_A_789_78#_c_644_n A_1119_379# 0.00438272f $X=5.97 $Y=2.31 $X2=-0.19
+ $Y2=-0.245
cc_635 N_A_789_78#_M1037_g N_VGND_c_1978_n 0.0192026f $X=4.02 $Y=0.73 $X2=0
+ $Y2=0
cc_636 N_A_789_78#_M1043_g N_VGND_c_1979_n 0.0113215f $X=7.16 $Y=0.915 $X2=0
+ $Y2=0
cc_637 N_A_789_78#_M1037_g N_VGND_c_1986_n 0.00475172f $X=4.02 $Y=0.73 $X2=0
+ $Y2=0
cc_638 N_A_789_78#_M1037_g N_VGND_c_2001_n 0.00499434f $X=4.02 $Y=0.73 $X2=0
+ $Y2=0
cc_639 N_A_789_78#_M1043_g N_VGND_c_2001_n 7.88961e-19 $X=7.16 $Y=0.915 $X2=0
+ $Y2=0
cc_640 N_A_789_78#_M1010_d N_A_1018_60#_c_2123_n 0.00709133f $X=5.525 $Y=0.3
+ $X2=0 $Y2=0
cc_641 N_A_789_78#_c_634_n N_A_1018_60#_c_2123_n 0.027978f $X=5.74 $Y=1.13 $X2=0
+ $Y2=0
cc_642 N_A_789_78#_c_638_n N_A_1018_60#_c_2123_n 0.00189874f $X=6.825 $Y=1.585
+ $X2=0 $Y2=0
cc_643 N_A_789_78#_c_638_n N_A_1018_60#_c_2125_n 0.00611341f $X=6.825 $Y=1.585
+ $X2=0 $Y2=0
cc_644 N_SET_B_M1017_g N_A_549_449#_M1010_g 0.0378368f $X=5.015 $Y=0.62 $X2=0
+ $Y2=0
cc_645 N_SET_B_M1024_g N_A_549_449#_M1040_g 0.0338471f $X=5.09 $Y=2.315 $X2=0
+ $Y2=0
cc_646 N_SET_B_c_767_n N_A_549_449#_c_893_n 6.42609e-19 $X=5.185 $Y=1.665 $X2=0
+ $Y2=0
cc_647 N_SET_B_c_769_n N_A_549_449#_c_893_n 0.0042644f $X=5 $Y=1.57 $X2=0 $Y2=0
cc_648 N_SET_B_c_770_n N_A_549_449#_c_893_n 0.013199f $X=5 $Y=1.57 $X2=0 $Y2=0
cc_649 N_SET_B_M1024_g N_A_549_449#_c_895_n 0.00206847f $X=5.09 $Y=2.315 $X2=0
+ $Y2=0
cc_650 N_SET_B_c_767_n N_A_549_449#_c_895_n 0.00586111f $X=5.185 $Y=1.665 $X2=0
+ $Y2=0
cc_651 N_SET_B_c_769_n N_A_549_449#_c_895_n 0.0038462f $X=5 $Y=1.57 $X2=0 $Y2=0
cc_652 N_SET_B_c_770_n N_A_549_449#_c_895_n 0.0122685f $X=5 $Y=1.57 $X2=0 $Y2=0
cc_653 N_SET_B_M1024_g N_A_549_449#_c_944_n 0.0116183f $X=5.09 $Y=2.315 $X2=0
+ $Y2=0
cc_654 N_SET_B_c_766_n N_A_549_449#_c_944_n 0.00812408f $X=8.735 $Y=1.665 $X2=0
+ $Y2=0
cc_655 N_SET_B_c_767_n N_A_549_449#_c_944_n 0.00314855f $X=5.185 $Y=1.665 $X2=0
+ $Y2=0
cc_656 N_SET_B_c_769_n N_A_549_449#_c_944_n 0.00288324f $X=5 $Y=1.57 $X2=0 $Y2=0
cc_657 N_SET_B_c_770_n N_A_549_449#_c_944_n 0.0139692f $X=5 $Y=1.57 $X2=0 $Y2=0
cc_658 N_SET_B_M1024_g N_A_549_449#_c_903_n 0.00214772f $X=5.09 $Y=2.315 $X2=0
+ $Y2=0
cc_659 N_SET_B_c_766_n N_A_549_449#_c_903_n 0.0247977f $X=8.735 $Y=1.665 $X2=0
+ $Y2=0
cc_660 N_SET_B_c_767_n N_A_549_449#_c_903_n 0.00259051f $X=5.185 $Y=1.665 $X2=0
+ $Y2=0
cc_661 N_SET_B_c_769_n N_A_549_449#_c_903_n 8.53228e-19 $X=5 $Y=1.57 $X2=0 $Y2=0
cc_662 N_SET_B_c_770_n N_A_549_449#_c_903_n 0.0164934f $X=5 $Y=1.57 $X2=0 $Y2=0
cc_663 N_SET_B_c_766_n N_A_549_449#_c_896_n 0.00150476f $X=8.735 $Y=1.665 $X2=0
+ $Y2=0
cc_664 N_SET_B_c_767_n N_A_549_449#_c_896_n 6.74491e-19 $X=5.185 $Y=1.665 $X2=0
+ $Y2=0
cc_665 N_SET_B_c_769_n N_A_549_449#_c_896_n 0.0221991f $X=5 $Y=1.57 $X2=0 $Y2=0
cc_666 N_SET_B_c_770_n N_A_549_449#_c_896_n 0.0014184f $X=5 $Y=1.57 $X2=0 $Y2=0
cc_667 N_SET_B_M1024_g N_A_223_119#_c_1042_n 0.00999935f $X=5.09 $Y=2.315 $X2=0
+ $Y2=0
cc_668 N_SET_B_c_766_n N_A_223_119#_c_1046_n 0.00661017f $X=8.735 $Y=1.665 $X2=0
+ $Y2=0
cc_669 SET_B N_A_223_119#_c_1029_n 0.00251875f $X=9.275 $Y=1.58 $X2=0 $Y2=0
cc_670 N_SET_B_c_766_n N_A_223_119#_c_1029_n 0.00215453f $X=8.735 $Y=1.665 $X2=0
+ $Y2=0
cc_671 N_SET_B_c_768_n N_A_223_119#_c_1029_n 8.33819e-19 $X=8.88 $Y=1.665 $X2=0
+ $Y2=0
cc_672 N_SET_B_c_766_n N_A_223_119#_c_1030_n 0.00656245f $X=8.735 $Y=1.665 $X2=0
+ $Y2=0
cc_673 N_SET_B_M1031_g N_A_1746_137#_c_1197_n 0.012159f $X=9.48 $Y=0.915 $X2=0
+ $Y2=0
cc_674 N_SET_B_c_764_n N_A_1746_137#_M1021_g 0.00855392f $X=9.735 $Y=2.065 $X2=0
+ $Y2=0
cc_675 N_SET_B_M1031_g N_A_1746_137#_c_1205_n 0.00661319f $X=9.48 $Y=0.915 $X2=0
+ $Y2=0
cc_676 SET_B N_A_1746_137#_c_1205_n 0.00288594f $X=9.275 $Y=1.58 $X2=0 $Y2=0
cc_677 N_SET_B_c_768_n N_A_1746_137#_c_1205_n 0.00186167f $X=8.88 $Y=1.665 $X2=0
+ $Y2=0
cc_678 N_SET_B_c_764_n N_A_1746_137#_c_1217_n 0.025114f $X=9.735 $Y=2.065 $X2=0
+ $Y2=0
cc_679 SET_B N_A_1746_137#_c_1217_n 0.0141034f $X=9.275 $Y=1.58 $X2=0 $Y2=0
cc_680 N_SET_B_c_764_n N_A_1746_137#_c_1221_n 0.00103892f $X=9.735 $Y=2.065
+ $X2=0 $Y2=0
cc_681 SET_B N_A_1746_137#_c_1221_n 0.0184689f $X=9.275 $Y=1.58 $X2=0 $Y2=0
cc_682 N_SET_B_c_768_n N_A_1746_137#_c_1221_n 9.47546e-19 $X=8.88 $Y=1.665 $X2=0
+ $Y2=0
cc_683 N_SET_B_c_764_n N_A_1746_137#_c_1222_n 0.00971149f $X=9.735 $Y=2.065
+ $X2=0 $Y2=0
cc_684 SET_B N_A_1746_137#_c_1222_n 0.0012483f $X=9.275 $Y=1.58 $X2=0 $Y2=0
cc_685 N_SET_B_c_764_n N_A_1746_137#_c_1223_n 0.0149063f $X=9.735 $Y=2.065 $X2=0
+ $Y2=0
cc_686 N_SET_B_c_764_n N_A_1746_137#_c_1210_n 0.0307118f $X=9.735 $Y=2.065 $X2=0
+ $Y2=0
cc_687 SET_B N_A_1746_137#_c_1210_n 0.0155957f $X=9.275 $Y=1.58 $X2=0 $Y2=0
cc_688 N_SET_B_M1031_g N_A_1542_428#_c_1375_n 0.02231f $X=9.48 $Y=0.915 $X2=0
+ $Y2=0
cc_689 N_SET_B_c_764_n N_A_1542_428#_c_1382_n 0.00617485f $X=9.735 $Y=2.065
+ $X2=0 $Y2=0
cc_690 SET_B N_A_1542_428#_c_1382_n 6.68025e-19 $X=9.275 $Y=1.58 $X2=0 $Y2=0
cc_691 N_SET_B_c_764_n N_A_1542_428#_c_1383_n 0.0234774f $X=9.735 $Y=2.065 $X2=0
+ $Y2=0
cc_692 N_SET_B_M1031_g N_A_1542_428#_c_1377_n 0.0157287f $X=9.48 $Y=0.915 $X2=0
+ $Y2=0
cc_693 N_SET_B_c_764_n N_A_1542_428#_c_1377_n 0.00911259f $X=9.735 $Y=2.065
+ $X2=0 $Y2=0
cc_694 SET_B N_A_1542_428#_c_1377_n 0.0551483f $X=9.275 $Y=1.58 $X2=0 $Y2=0
cc_695 N_SET_B_c_766_n N_A_1542_428#_c_1377_n 0.0136023f $X=8.735 $Y=1.665 $X2=0
+ $Y2=0
cc_696 N_SET_B_c_768_n N_A_1542_428#_c_1377_n 0.00377658f $X=8.88 $Y=1.665 $X2=0
+ $Y2=0
cc_697 N_SET_B_c_766_n N_A_1542_428#_c_1384_n 0.00971822f $X=8.735 $Y=1.665
+ $X2=0 $Y2=0
cc_698 SET_B N_A_1542_428#_c_1378_n 0.00409081f $X=9.275 $Y=1.58 $X2=0 $Y2=0
cc_699 N_SET_B_c_766_n N_A_1542_428#_c_1378_n 0.0234144f $X=8.735 $Y=1.665 $X2=0
+ $Y2=0
cc_700 N_SET_B_c_768_n N_A_1542_428#_c_1378_n 9.30425e-19 $X=8.88 $Y=1.665 $X2=0
+ $Y2=0
cc_701 N_SET_B_c_766_n N_A_1542_428#_c_1379_n 0.00738362f $X=8.735 $Y=1.665
+ $X2=0 $Y2=0
cc_702 N_SET_B_M1031_g N_A_1542_428#_c_1380_n 0.00377985f $X=9.48 $Y=0.915 $X2=0
+ $Y2=0
cc_703 N_SET_B_c_764_n N_A_1542_428#_c_1380_n 0.00108617f $X=9.735 $Y=2.065
+ $X2=0 $Y2=0
cc_704 SET_B N_A_1542_428#_c_1380_n 0.0146873f $X=9.275 $Y=1.58 $X2=0 $Y2=0
cc_705 N_SET_B_M1031_g N_A_1542_428#_c_1381_n 0.00628089f $X=9.48 $Y=0.915 $X2=0
+ $Y2=0
cc_706 N_SET_B_c_764_n N_A_1542_428#_c_1381_n 0.013423f $X=9.735 $Y=2.065 $X2=0
+ $Y2=0
cc_707 SET_B N_A_1542_428#_c_1381_n 2.50891e-19 $X=9.275 $Y=1.58 $X2=0 $Y2=0
cc_708 N_SET_B_c_766_n N_A_1191_21#_M1003_g 0.00366367f $X=8.735 $Y=1.665 $X2=0
+ $Y2=0
cc_709 N_SET_B_M1031_g N_A_1191_21#_c_1472_n 0.0103118f $X=9.48 $Y=0.915 $X2=0
+ $Y2=0
cc_710 N_SET_B_M1024_g N_VPWR_c_1699_n 0.00652951f $X=5.09 $Y=2.315 $X2=0 $Y2=0
cc_711 N_SET_B_c_766_n N_VPWR_c_1700_n 0.00957433f $X=8.735 $Y=1.665 $X2=0 $Y2=0
cc_712 N_SET_B_c_764_n N_VPWR_c_1701_n 0.00393161f $X=9.735 $Y=2.065 $X2=0 $Y2=0
cc_713 N_SET_B_c_764_n N_VPWR_c_1714_n 0.00449508f $X=9.735 $Y=2.065 $X2=0 $Y2=0
cc_714 N_SET_B_M1024_g N_VPWR_c_1695_n 9.39239e-19 $X=5.09 $Y=2.315 $X2=0 $Y2=0
cc_715 N_SET_B_c_764_n N_VPWR_c_1695_n 0.00877693f $X=9.735 $Y=2.065 $X2=0 $Y2=0
cc_716 N_SET_B_M1017_g N_VGND_c_1978_n 0.00352591f $X=5.015 $Y=0.62 $X2=0 $Y2=0
cc_717 N_SET_B_M1031_g N_VGND_c_1980_n 0.00660997f $X=9.48 $Y=0.915 $X2=0 $Y2=0
cc_718 N_SET_B_M1017_g N_VGND_c_1989_n 0.00318662f $X=5.015 $Y=0.62 $X2=0 $Y2=0
cc_719 N_SET_B_M1017_g N_VGND_c_2001_n 0.00547455f $X=5.015 $Y=0.62 $X2=0 $Y2=0
cc_720 N_SET_B_M1031_g N_VGND_c_2001_n 8.79083e-19 $X=9.48 $Y=0.915 $X2=0 $Y2=0
cc_721 N_SET_B_M1017_g N_A_1018_60#_c_2124_n 0.00490817f $X=5.015 $Y=0.62 $X2=0
+ $Y2=0
cc_722 N_SET_B_c_767_n N_A_1018_60#_c_2124_n 0.00126491f $X=5.185 $Y=1.665 $X2=0
+ $Y2=0
cc_723 N_SET_B_c_769_n N_A_1018_60#_c_2124_n 4.55546e-19 $X=5 $Y=1.57 $X2=0
+ $Y2=0
cc_724 N_SET_B_c_770_n N_A_1018_60#_c_2124_n 0.0031303f $X=5 $Y=1.57 $X2=0 $Y2=0
cc_725 N_SET_B_M1031_g N_A_1911_119#_c_2148_n 0.00639462f $X=9.48 $Y=0.915 $X2=0
+ $Y2=0
cc_726 N_A_549_449#_c_890_n N_A_223_119#_M1013_g 0.00535476f $X=3.12 $Y=0.725
+ $X2=0 $Y2=0
cc_727 N_A_549_449#_c_891_n N_A_223_119#_M1013_g 0.00349937f $X=3.175 $Y=2.225
+ $X2=0 $Y2=0
cc_728 N_A_549_449#_c_891_n N_A_223_119#_c_1038_n 0.00548166f $X=3.175 $Y=2.225
+ $X2=0 $Y2=0
cc_729 N_A_549_449#_c_891_n N_A_223_119#_c_1039_n 0.00962018f $X=3.175 $Y=2.225
+ $X2=0 $Y2=0
cc_730 N_A_549_449#_c_892_n N_A_223_119#_c_1039_n 0.00218303f $X=3.905 $Y=2.225
+ $X2=0 $Y2=0
cc_731 N_A_549_449#_c_905_n N_A_223_119#_c_1039_n 0.0058172f $X=3.42 $Y=2.455
+ $X2=0 $Y2=0
cc_732 N_A_549_449#_c_891_n N_A_223_119#_c_1040_n 0.00252046f $X=3.175 $Y=2.225
+ $X2=0 $Y2=0
cc_733 N_A_549_449#_c_905_n N_A_223_119#_c_1040_n 0.00127737f $X=3.42 $Y=2.455
+ $X2=0 $Y2=0
cc_734 N_A_549_449#_c_891_n N_A_223_119#_M1030_g 0.0010298f $X=3.175 $Y=2.225
+ $X2=0 $Y2=0
cc_735 N_A_549_449#_c_899_n N_A_223_119#_M1030_g 0.0120447f $X=3.82 $Y=2.31
+ $X2=0 $Y2=0
cc_736 N_A_549_449#_c_905_n N_A_223_119#_M1030_g 0.00836223f $X=3.42 $Y=2.455
+ $X2=0 $Y2=0
cc_737 N_A_549_449#_M1040_g N_A_223_119#_c_1042_n 0.00999935f $X=5.52 $Y=2.315
+ $X2=0 $Y2=0
cc_738 N_A_549_449#_c_899_n N_A_223_119#_c_1042_n 0.00609554f $X=3.82 $Y=2.31
+ $X2=0 $Y2=0
cc_739 N_A_549_449#_c_891_n N_A_223_119#_c_1034_n 0.00524877f $X=3.175 $Y=2.225
+ $X2=0 $Y2=0
cc_740 N_A_549_449#_c_892_n N_A_223_119#_c_1034_n 0.00103072f $X=3.905 $Y=2.225
+ $X2=0 $Y2=0
cc_741 N_A_549_449#_M1040_g N_A_1191_21#_M1003_g 0.0361146f $X=5.52 $Y=2.315
+ $X2=0 $Y2=0
cc_742 N_A_549_449#_c_944_n N_A_1191_21#_M1003_g 6.21434e-19 $X=5.375 $Y=2.045
+ $X2=0 $Y2=0
cc_743 N_A_549_449#_c_903_n N_A_1191_21#_M1003_g 0.0010935f $X=5.54 $Y=1.57
+ $X2=0 $Y2=0
cc_744 N_A_549_449#_c_896_n N_A_1191_21#_M1003_g 0.0171877f $X=5.54 $Y=1.57
+ $X2=0 $Y2=0
cc_745 N_A_549_449#_M1010_g N_A_1191_21#_c_1473_n 0.0314416f $X=5.45 $Y=0.62
+ $X2=0 $Y2=0
cc_746 N_A_549_449#_c_895_n N_VPWR_M1039_d 0.0011867f $X=4.635 $Y=1.96 $X2=0
+ $Y2=0
cc_747 N_A_549_449#_c_944_n N_VPWR_M1039_d 0.00919665f $X=5.375 $Y=2.045 $X2=0
+ $Y2=0
cc_748 N_A_549_449#_c_902_n N_VPWR_M1039_d 0.00144282f $X=4.72 $Y=2.045 $X2=0
+ $Y2=0
cc_749 N_A_549_449#_c_905_n N_VPWR_c_1710_n 0.00627379f $X=3.42 $Y=2.455 $X2=0
+ $Y2=0
cc_750 N_A_549_449#_M1040_g N_VPWR_c_1695_n 9.39239e-19 $X=5.52 $Y=2.315 $X2=0
+ $Y2=0
cc_751 N_A_549_449#_c_905_n N_VPWR_c_1695_n 0.00961952f $X=3.42 $Y=2.455 $X2=0
+ $Y2=0
cc_752 N_A_549_449#_c_890_n N_A_463_449#_c_1849_n 0.0203767f $X=3.12 $Y=0.725
+ $X2=0 $Y2=0
cc_753 N_A_549_449#_c_891_n N_A_463_449#_c_1849_n 0.0083955f $X=3.175 $Y=2.225
+ $X2=0 $Y2=0
cc_754 N_A_549_449#_M1023_d N_A_463_449#_c_1850_n 5.87996e-19 $X=2.745 $Y=2.245
+ $X2=0 $Y2=0
cc_755 N_A_549_449#_c_905_n N_A_463_449#_c_1850_n 0.00657775f $X=3.42 $Y=2.455
+ $X2=0 $Y2=0
cc_756 N_A_549_449#_M1023_d N_A_463_449#_c_1853_n 0.00427072f $X=2.745 $Y=2.245
+ $X2=0 $Y2=0
cc_757 N_A_549_449#_c_905_n N_A_463_449#_c_1853_n 0.0216786f $X=3.42 $Y=2.455
+ $X2=0 $Y2=0
cc_758 N_A_549_449#_c_891_n N_A_463_449#_c_1851_n 0.0780793f $X=3.175 $Y=2.225
+ $X2=0 $Y2=0
cc_759 N_A_549_449#_c_899_n A_709_449# 0.00630734f $X=3.82 $Y=2.31 $X2=-0.19
+ $Y2=-0.245
cc_760 N_A_549_449#_c_944_n A_1119_379# 0.00214968f $X=5.375 $Y=2.045 $X2=-0.19
+ $Y2=-0.245
cc_761 N_A_549_449#_c_903_n A_1119_379# 5.75572e-19 $X=5.54 $Y=1.57 $X2=-0.19
+ $Y2=-0.245
cc_762 N_A_549_449#_c_890_n N_VGND_c_1986_n 0.00611431f $X=3.12 $Y=0.725 $X2=0
+ $Y2=0
cc_763 N_A_549_449#_M1010_g N_VGND_c_1989_n 0.00318662f $X=5.45 $Y=0.62 $X2=0
+ $Y2=0
cc_764 N_A_549_449#_M1010_g N_VGND_c_2001_n 0.00492332f $X=5.45 $Y=0.62 $X2=0
+ $Y2=0
cc_765 N_A_549_449#_c_890_n N_VGND_c_2001_n 0.00653993f $X=3.12 $Y=0.725 $X2=0
+ $Y2=0
cc_766 N_A_549_449#_M1010_g N_A_1018_60#_c_2123_n 0.0122347f $X=5.45 $Y=0.62
+ $X2=0 $Y2=0
cc_767 N_A_549_449#_c_896_n N_A_1018_60#_c_2123_n 8.84098e-19 $X=5.54 $Y=1.57
+ $X2=0 $Y2=0
cc_768 N_A_549_449#_M1010_g N_A_1018_60#_c_2124_n 0.00480277f $X=5.45 $Y=0.62
+ $X2=0 $Y2=0
cc_769 N_A_549_449#_c_903_n N_A_1018_60#_c_2124_n 6.11501e-19 $X=5.54 $Y=1.57
+ $X2=0 $Y2=0
cc_770 N_A_223_119#_c_1032_n N_A_1746_137#_c_1197_n 0.0213733f $X=8.415 $Y=1.31
+ $X2=0 $Y2=0
cc_771 N_A_223_119#_c_1030_n N_A_1746_137#_c_1205_n 0.0213733f $X=8.34 $Y=1.385
+ $X2=0 $Y2=0
cc_772 N_A_223_119#_c_1032_n N_A_1542_428#_c_1376_n 0.006368f $X=8.415 $Y=1.31
+ $X2=0 $Y2=0
cc_773 N_A_223_119#_c_1030_n N_A_1542_428#_c_1377_n 0.00217836f $X=8.34 $Y=1.385
+ $X2=0 $Y2=0
cc_774 N_A_223_119#_c_1032_n N_A_1542_428#_c_1377_n 0.015156f $X=8.415 $Y=1.31
+ $X2=0 $Y2=0
cc_775 N_A_223_119#_M1020_g N_A_1542_428#_c_1384_n 0.0101949f $X=7.635 $Y=2.56
+ $X2=0 $Y2=0
cc_776 N_A_223_119#_c_1045_n N_A_1542_428#_c_1384_n 0.00997989f $X=7.985 $Y=1.99
+ $X2=0 $Y2=0
cc_777 N_A_223_119#_M1020_g N_A_1542_428#_c_1378_n 5.56793e-19 $X=7.635 $Y=2.56
+ $X2=0 $Y2=0
cc_778 N_A_223_119#_c_1045_n N_A_1542_428#_c_1378_n 0.0101706f $X=7.985 $Y=1.99
+ $X2=0 $Y2=0
cc_779 N_A_223_119#_c_1029_n N_A_1542_428#_c_1378_n 0.0144732f $X=8.06 $Y=1.915
+ $X2=0 $Y2=0
cc_780 N_A_223_119#_c_1031_n N_A_1542_428#_c_1378_n 0.00863083f $X=8.135
+ $Y=1.385 $X2=0 $Y2=0
cc_781 N_A_223_119#_c_1032_n N_A_1542_428#_c_1378_n 4.24368e-19 $X=8.415 $Y=1.31
+ $X2=0 $Y2=0
cc_782 N_A_223_119#_c_1031_n N_A_1542_428#_c_1379_n 0.00780864f $X=8.135
+ $Y=1.385 $X2=0 $Y2=0
cc_783 N_A_223_119#_c_1042_n N_A_1191_21#_M1003_g 0.0101786f $X=7.56 $Y=3.15
+ $X2=0 $Y2=0
cc_784 N_A_223_119#_c_1032_n N_A_1191_21#_c_1472_n 0.00495681f $X=8.415 $Y=1.31
+ $X2=0 $Y2=0
cc_785 N_A_223_119#_c_1051_n N_VPWR_c_1698_n 0.0258905f $X=1.375 $Y=2.39 $X2=0
+ $Y2=0
cc_786 N_A_223_119#_c_1052_n N_VPWR_c_1698_n 0.0260518f $X=2.295 $Y=1.96 $X2=0
+ $Y2=0
cc_787 N_A_223_119#_c_1042_n N_VPWR_c_1699_n 0.0253641f $X=7.56 $Y=3.15 $X2=0
+ $Y2=0
cc_788 N_A_223_119#_c_1042_n N_VPWR_c_1700_n 0.0261591f $X=7.56 $Y=3.15 $X2=0
+ $Y2=0
cc_789 N_A_223_119#_c_1051_n N_VPWR_c_1708_n 0.0111657f $X=1.375 $Y=2.39 $X2=0
+ $Y2=0
cc_790 N_A_223_119#_c_1043_n N_VPWR_c_1710_n 0.0441847f $X=3.545 $Y=3.15 $X2=0
+ $Y2=0
cc_791 N_A_223_119#_c_1042_n N_VPWR_c_1712_n 0.0412435f $X=7.56 $Y=3.15 $X2=0
+ $Y2=0
cc_792 N_A_223_119#_c_1042_n N_VPWR_c_1713_n 0.0356346f $X=7.56 $Y=3.15 $X2=0
+ $Y2=0
cc_793 N_A_223_119#_c_1042_n N_VPWR_c_1695_n 0.134269f $X=7.56 $Y=3.15 $X2=0
+ $Y2=0
cc_794 N_A_223_119#_c_1043_n N_VPWR_c_1695_n 0.0104239f $X=3.545 $Y=3.15 $X2=0
+ $Y2=0
cc_795 N_A_223_119#_c_1051_n N_VPWR_c_1695_n 0.0114323f $X=1.375 $Y=2.39 $X2=0
+ $Y2=0
cc_796 N_A_223_119#_M1013_g N_A_463_449#_c_1849_n 0.00943133f $X=2.825 $Y=0.805
+ $X2=0 $Y2=0
cc_797 N_A_223_119#_M1013_g N_A_463_449#_c_1850_n 0.00596599f $X=2.825 $Y=0.805
+ $X2=0 $Y2=0
cc_798 N_A_223_119#_c_1038_n N_A_463_449#_c_1850_n 0.006209f $X=3.06 $Y=2 $X2=0
+ $Y2=0
cc_799 N_A_223_119#_M1030_g N_A_463_449#_c_1850_n 2.64472e-19 $X=3.47 $Y=2.455
+ $X2=0 $Y2=0
cc_800 N_A_223_119#_c_1033_n N_A_463_449#_c_1850_n 0.00497011f $X=2.75 $Y=1.645
+ $X2=0 $Y2=0
cc_801 N_A_223_119#_c_1034_n N_A_463_449#_c_1850_n 0.0120367f $X=2.825 $Y=1.66
+ $X2=0 $Y2=0
cc_802 N_A_223_119#_c_1052_n N_A_463_449#_c_1850_n 0.0137875f $X=2.295 $Y=1.96
+ $X2=0 $Y2=0
cc_803 N_A_223_119#_c_1036_n N_A_463_449#_c_1850_n 0.0269458f $X=2.46 $Y=1.645
+ $X2=0 $Y2=0
cc_804 N_A_223_119#_c_1033_n N_A_463_449#_c_1853_n 0.00161187f $X=2.75 $Y=1.645
+ $X2=0 $Y2=0
cc_805 N_A_223_119#_c_1052_n N_A_463_449#_c_1853_n 0.0146267f $X=2.295 $Y=1.96
+ $X2=0 $Y2=0
cc_806 N_A_223_119#_M1013_g N_A_463_449#_c_1851_n 0.0121041f $X=2.825 $Y=0.805
+ $X2=0 $Y2=0
cc_807 N_A_223_119#_c_1033_n N_A_463_449#_c_1851_n 0.0087512f $X=2.75 $Y=1.645
+ $X2=0 $Y2=0
cc_808 N_A_223_119#_c_1036_n N_A_463_449#_c_1851_n 0.00951907f $X=2.46 $Y=1.645
+ $X2=0 $Y2=0
cc_809 N_A_223_119#_c_1037_n N_VGND_c_1977_n 0.0159918f $X=1.255 $Y=0.785 $X2=0
+ $Y2=0
cc_810 N_A_223_119#_c_1037_n N_VGND_c_1988_n 0.00738549f $X=1.255 $Y=0.785 $X2=0
+ $Y2=0
cc_811 N_A_223_119#_M1013_g N_VGND_c_2001_n 9.39239e-19 $X=2.825 $Y=0.805 $X2=0
+ $Y2=0
cc_812 N_A_223_119#_c_1032_n N_VGND_c_2001_n 9.72468e-19 $X=8.415 $Y=1.31 $X2=0
+ $Y2=0
cc_813 N_A_223_119#_c_1037_n N_VGND_c_2001_n 0.0101768f $X=1.255 $Y=0.785 $X2=0
+ $Y2=0
cc_814 N_A_1746_137#_c_1251_p N_A_1542_428#_c_1375_n 0.00813722f $X=10.22
+ $Y=0.89 $X2=0 $Y2=0
cc_815 N_A_1746_137#_c_1208_n N_A_1542_428#_c_1375_n 0.00127126f $X=10.39 $Y=2.2
+ $X2=0 $Y2=0
cc_816 N_A_1746_137#_c_1253_p N_A_1542_428#_c_1383_n 0.0140926f $X=10.305
+ $Y=2.285 $X2=0 $Y2=0
cc_817 N_A_1746_137#_c_1208_n N_A_1542_428#_c_1383_n 0.00645239f $X=10.39 $Y=2.2
+ $X2=0 $Y2=0
cc_818 N_A_1746_137#_c_1223_n N_A_1542_428#_c_1383_n 0.0126811f $X=9.95 $Y=2.365
+ $X2=0 $Y2=0
cc_819 N_A_1746_137#_c_1197_n N_A_1542_428#_c_1377_n 0.0150964f $X=8.805 $Y=1.31
+ $X2=0 $Y2=0
cc_820 N_A_1746_137#_c_1205_n N_A_1542_428#_c_1377_n 0.00485975f $X=8.96
+ $Y=1.385 $X2=0 $Y2=0
cc_821 N_A_1746_137#_c_1205_n N_A_1542_428#_c_1378_n 5.27174e-19 $X=8.96
+ $Y=1.385 $X2=0 $Y2=0
cc_822 N_A_1746_137#_c_1253_p N_A_1542_428#_c_1380_n 2.70995e-19 $X=10.305
+ $Y=2.285 $X2=0 $Y2=0
cc_823 N_A_1746_137#_c_1208_n N_A_1542_428#_c_1380_n 0.0318835f $X=10.39 $Y=2.2
+ $X2=0 $Y2=0
cc_824 N_A_1746_137#_c_1223_n N_A_1542_428#_c_1380_n 0.00921981f $X=9.95
+ $Y=2.365 $X2=0 $Y2=0
cc_825 N_A_1746_137#_c_1262_p N_A_1542_428#_c_1380_n 0.00355462f $X=10.305
+ $Y=1.165 $X2=0 $Y2=0
cc_826 N_A_1746_137#_c_1208_n N_A_1542_428#_c_1381_n 0.00751936f $X=10.39 $Y=2.2
+ $X2=0 $Y2=0
cc_827 N_A_1746_137#_c_1223_n N_A_1542_428#_c_1381_n 0.00126241f $X=9.95
+ $Y=2.365 $X2=0 $Y2=0
cc_828 N_A_1746_137#_c_1262_p N_A_1542_428#_c_1381_n 0.00297214f $X=10.305
+ $Y=1.165 $X2=0 $Y2=0
cc_829 N_A_1746_137#_c_1219_n N_A_1191_21#_M1026_s 0.0031491f $X=11.795 $Y=2.285
+ $X2=0 $Y2=0
cc_830 N_A_1746_137#_c_1197_n N_A_1191_21#_c_1472_n 0.00495681f $X=8.805 $Y=1.31
+ $X2=0 $Y2=0
cc_831 N_A_1746_137#_c_1251_p N_A_1191_21#_M1038_g 0.015989f $X=10.22 $Y=0.89
+ $X2=0 $Y2=0
cc_832 N_A_1746_137#_c_1208_n N_A_1191_21#_M1038_g 0.00389707f $X=10.39 $Y=2.2
+ $X2=0 $Y2=0
cc_833 N_A_1746_137#_c_1262_p N_A_1191_21#_M1038_g 0.00430892f $X=10.305
+ $Y=1.165 $X2=0 $Y2=0
cc_834 N_A_1746_137#_c_1208_n N_A_1191_21#_M1009_g 0.0154947f $X=10.39 $Y=2.2
+ $X2=0 $Y2=0
cc_835 N_A_1746_137#_c_1219_n N_A_1191_21#_M1009_g 0.0162535f $X=11.795 $Y=2.285
+ $X2=0 $Y2=0
cc_836 N_A_1746_137#_c_1223_n N_A_1191_21#_M1009_g 0.0021245f $X=9.95 $Y=2.365
+ $X2=0 $Y2=0
cc_837 N_A_1746_137#_c_1274_p N_A_1191_21#_M1009_g 0.00316892f $X=10.39 $Y=2.285
+ $X2=0 $Y2=0
cc_838 N_A_1746_137#_c_1262_p N_A_1191_21#_c_1475_n 0.0376918f $X=10.305
+ $Y=1.165 $X2=0 $Y2=0
cc_839 N_A_1746_137#_c_1208_n N_A_1191_21#_c_1476_n 0.00793511f $X=10.39 $Y=2.2
+ $X2=0 $Y2=0
cc_840 N_A_1746_137#_c_1219_n N_A_1191_21#_c_1476_n 0.00141173f $X=11.795
+ $Y=2.285 $X2=0 $Y2=0
cc_841 N_A_1746_137#_c_1251_p N_A_1191_21#_c_1478_n 0.0134574f $X=10.22 $Y=0.89
+ $X2=0 $Y2=0
cc_842 N_A_1746_137#_c_1208_n N_A_1191_21#_c_1483_n 0.027189f $X=10.39 $Y=2.2
+ $X2=0 $Y2=0
cc_843 N_A_1746_137#_c_1219_n N_A_1191_21#_c_1483_n 0.0197178f $X=11.795
+ $Y=2.285 $X2=0 $Y2=0
cc_844 N_A_1746_137#_M1011_g N_A_1191_21#_c_1484_n 2.91174e-19 $X=12.02 $Y=2.34
+ $X2=0 $Y2=0
cc_845 N_A_1746_137#_c_1219_n N_A_1191_21#_c_1484_n 0.0309089f $X=11.795
+ $Y=2.285 $X2=0 $Y2=0
cc_846 N_A_1746_137#_c_1220_n N_A_1191_21#_c_1484_n 0.0152162f $X=11.88 $Y=2.2
+ $X2=0 $Y2=0
cc_847 N_A_1746_137#_c_1212_n N_RESET_B_c_1581_n 0.00144422f $X=11.96 $Y=1.185
+ $X2=0 $Y2=0
cc_848 N_A_1746_137#_M1011_g N_RESET_B_M1026_g 0.0292262f $X=12.02 $Y=2.34 $X2=0
+ $Y2=0
cc_849 N_A_1746_137#_c_1219_n N_RESET_B_M1026_g 0.0203764f $X=11.795 $Y=2.285
+ $X2=0 $Y2=0
cc_850 N_A_1746_137#_c_1220_n N_RESET_B_M1026_g 0.00976358f $X=11.88 $Y=2.2
+ $X2=0 $Y2=0
cc_851 N_A_1746_137#_c_1212_n N_RESET_B_M1001_g 0.0145949f $X=11.96 $Y=1.185
+ $X2=0 $Y2=0
cc_852 N_A_1746_137#_c_1209_n N_RESET_B_c_1585_n 0.018794f $X=11.96 $Y=1.35
+ $X2=0 $Y2=0
cc_853 N_A_1746_137#_c_1211_n N_RESET_B_c_1585_n 0.00116723f $X=11.96 $Y=1.26
+ $X2=0 $Y2=0
cc_854 N_A_1746_137#_c_1209_n N_RESET_B_c_1586_n 0.0012048f $X=11.96 $Y=1.35
+ $X2=0 $Y2=0
cc_855 N_A_1746_137#_c_1211_n N_RESET_B_c_1586_n 0.0208775f $X=11.96 $Y=1.26
+ $X2=0 $Y2=0
cc_856 N_A_1746_137#_c_1203_n N_A_2618_131#_M1018_g 0.0158431f $X=13.45 $Y=1.185
+ $X2=0 $Y2=0
cc_857 N_A_1746_137#_M1006_g N_A_2618_131#_M1007_g 0.0181462f $X=13.45 $Y=2.155
+ $X2=0 $Y2=0
cc_858 N_A_1746_137#_c_1201_n N_A_2618_131#_c_1625_n 0.00222112f $X=12.46
+ $Y=1.185 $X2=0 $Y2=0
cc_859 N_A_1746_137#_c_1202_n N_A_2618_131#_c_1625_n 0.0100769f $X=13.375
+ $Y=1.26 $X2=0 $Y2=0
cc_860 N_A_1746_137#_c_1203_n N_A_2618_131#_c_1625_n 0.0101691f $X=13.45
+ $Y=1.185 $X2=0 $Y2=0
cc_861 N_A_1746_137#_c_1207_n N_A_2618_131#_c_1625_n 0.0017395f $X=13.45 $Y=1.26
+ $X2=0 $Y2=0
cc_862 N_A_1746_137#_M1029_g N_A_2618_131#_c_1626_n 0.00270855f $X=12.45 $Y=2.34
+ $X2=0 $Y2=0
cc_863 N_A_1746_137#_M1006_g N_A_2618_131#_c_1626_n 0.0167639f $X=13.45 $Y=2.155
+ $X2=0 $Y2=0
cc_864 N_A_1746_137#_M1006_g N_A_2618_131#_c_1627_n 0.0117789f $X=13.45 $Y=2.155
+ $X2=0 $Y2=0
cc_865 N_A_1746_137#_c_1207_n N_A_2618_131#_c_1627_n 0.00722589f $X=13.45
+ $Y=1.26 $X2=0 $Y2=0
cc_866 N_A_1746_137#_M1029_g N_A_2618_131#_c_1628_n 0.00447424f $X=12.45 $Y=2.34
+ $X2=0 $Y2=0
cc_867 N_A_1746_137#_c_1202_n N_A_2618_131#_c_1628_n 0.00873042f $X=13.375
+ $Y=1.26 $X2=0 $Y2=0
cc_868 N_A_1746_137#_M1006_g N_A_2618_131#_c_1628_n 0.00606798f $X=13.45
+ $Y=2.155 $X2=0 $Y2=0
cc_869 N_A_1746_137#_c_1207_n N_A_2618_131#_c_1629_n 0.0181351f $X=13.45 $Y=1.26
+ $X2=0 $Y2=0
cc_870 N_A_1746_137#_c_1217_n N_VPWR_M1021_d 0.00603025f $X=9.785 $Y=2.285 $X2=0
+ $Y2=0
cc_871 N_A_1746_137#_c_1219_n N_VPWR_M1009_d 0.00659114f $X=11.795 $Y=2.285
+ $X2=0 $Y2=0
cc_872 N_A_1746_137#_c_1219_n N_VPWR_M1026_d 0.00830173f $X=11.795 $Y=2.285
+ $X2=0 $Y2=0
cc_873 N_A_1746_137#_c_1220_n N_VPWR_M1026_d 0.00561339f $X=11.88 $Y=2.2 $X2=0
+ $Y2=0
cc_874 N_A_1746_137#_M1021_g N_VPWR_c_1701_n 0.0115296f $X=8.99 $Y=2.74 $X2=0
+ $Y2=0
cc_875 N_A_1746_137#_c_1217_n N_VPWR_c_1701_n 0.0192803f $X=9.785 $Y=2.285 $X2=0
+ $Y2=0
cc_876 N_A_1746_137#_c_1223_n N_VPWR_c_1701_n 0.0168566f $X=9.95 $Y=2.365 $X2=0
+ $Y2=0
cc_877 N_A_1746_137#_c_1219_n N_VPWR_c_1702_n 0.0210602f $X=11.795 $Y=2.285
+ $X2=0 $Y2=0
cc_878 N_A_1746_137#_c_1223_n N_VPWR_c_1702_n 0.0150558f $X=9.95 $Y=2.365 $X2=0
+ $Y2=0
cc_879 N_A_1746_137#_M1011_g N_VPWR_c_1703_n 0.0105837f $X=12.02 $Y=2.34 $X2=0
+ $Y2=0
cc_880 N_A_1746_137#_M1029_g N_VPWR_c_1703_n 5.19309e-19 $X=12.45 $Y=2.34 $X2=0
+ $Y2=0
cc_881 N_A_1746_137#_c_1219_n N_VPWR_c_1703_n 0.0216349f $X=11.795 $Y=2.285
+ $X2=0 $Y2=0
cc_882 N_A_1746_137#_M1029_g N_VPWR_c_1704_n 0.0114295f $X=12.45 $Y=2.34 $X2=0
+ $Y2=0
cc_883 N_A_1746_137#_c_1202_n N_VPWR_c_1704_n 0.0046297f $X=13.375 $Y=1.26 $X2=0
+ $Y2=0
cc_884 N_A_1746_137#_M1006_g N_VPWR_c_1704_n 0.00436498f $X=13.45 $Y=2.155 $X2=0
+ $Y2=0
cc_885 N_A_1746_137#_M1006_g N_VPWR_c_1705_n 0.00661754f $X=13.45 $Y=2.155 $X2=0
+ $Y2=0
cc_886 N_A_1746_137#_M1021_g N_VPWR_c_1713_n 0.00570944f $X=8.99 $Y=2.74 $X2=0
+ $Y2=0
cc_887 N_A_1746_137#_c_1223_n N_VPWR_c_1714_n 0.0157615f $X=9.95 $Y=2.365 $X2=0
+ $Y2=0
cc_888 N_A_1746_137#_M1011_g N_VPWR_c_1716_n 0.00389963f $X=12.02 $Y=2.34 $X2=0
+ $Y2=0
cc_889 N_A_1746_137#_M1029_g N_VPWR_c_1716_n 0.00430227f $X=12.45 $Y=2.34 $X2=0
+ $Y2=0
cc_890 N_A_1746_137#_M1006_g N_VPWR_c_1717_n 0.00312414f $X=13.45 $Y=2.155 $X2=0
+ $Y2=0
cc_891 N_A_1746_137#_M1021_g N_VPWR_c_1695_n 0.00542671f $X=8.99 $Y=2.74 $X2=0
+ $Y2=0
cc_892 N_A_1746_137#_M1011_g N_VPWR_c_1695_n 0.00764692f $X=12.02 $Y=2.34 $X2=0
+ $Y2=0
cc_893 N_A_1746_137#_M1029_g N_VPWR_c_1695_n 0.00815169f $X=12.45 $Y=2.34 $X2=0
+ $Y2=0
cc_894 N_A_1746_137#_M1006_g N_VPWR_c_1695_n 0.00410284f $X=13.45 $Y=2.155 $X2=0
+ $Y2=0
cc_895 N_A_1746_137#_c_1223_n N_VPWR_c_1695_n 0.0120285f $X=9.95 $Y=2.365 $X2=0
+ $Y2=0
cc_896 N_A_1746_137#_c_1253_p A_2048_428# 5.34178e-19 $X=10.305 $Y=2.285
+ $X2=-0.19 $Y2=-0.245
cc_897 N_A_1746_137#_c_1208_n A_2048_428# 6.49906e-19 $X=10.39 $Y=2.2 $X2=-0.19
+ $Y2=-0.245
cc_898 N_A_1746_137#_c_1274_p A_2048_428# 0.00392462f $X=10.39 $Y=2.285
+ $X2=-0.19 $Y2=-0.245
cc_899 N_A_1746_137#_M1011_g N_Q_N_c_1907_n 0.00103358f $X=12.02 $Y=2.34 $X2=0
+ $Y2=0
cc_900 N_A_1746_137#_c_1199_n N_Q_N_c_1907_n 0.00325129f $X=12.375 $Y=1.26 $X2=0
+ $Y2=0
cc_901 N_A_1746_137#_M1029_g N_Q_N_c_1907_n 0.00163541f $X=12.45 $Y=2.34 $X2=0
+ $Y2=0
cc_902 N_A_1746_137#_c_1220_n N_Q_N_c_1907_n 0.0164907f $X=11.88 $Y=2.2 $X2=0
+ $Y2=0
cc_903 N_A_1746_137#_M1029_g N_Q_N_c_1908_n 0.0156888f $X=12.45 $Y=2.34 $X2=0
+ $Y2=0
cc_904 N_A_1746_137#_c_1199_n N_Q_N_c_1915_n 0.00183f $X=12.375 $Y=1.26 $X2=0
+ $Y2=0
cc_905 N_A_1746_137#_c_1201_n N_Q_N_c_1915_n 0.00180034f $X=12.46 $Y=1.185 $X2=0
+ $Y2=0
cc_906 N_A_1746_137#_c_1212_n N_Q_N_c_1915_n 0.00308283f $X=11.96 $Y=1.185 $X2=0
+ $Y2=0
cc_907 N_A_1746_137#_M1011_g N_Q_N_c_1906_n 0.00126615f $X=12.02 $Y=2.34 $X2=0
+ $Y2=0
cc_908 N_A_1746_137#_c_1199_n N_Q_N_c_1906_n 0.00852334f $X=12.375 $Y=1.26 $X2=0
+ $Y2=0
cc_909 N_A_1746_137#_M1029_g N_Q_N_c_1906_n 0.0105158f $X=12.45 $Y=2.34 $X2=0
+ $Y2=0
cc_910 N_A_1746_137#_c_1201_n N_Q_N_c_1906_n 0.0040404f $X=12.46 $Y=1.185 $X2=0
+ $Y2=0
cc_911 N_A_1746_137#_c_1206_n N_Q_N_c_1906_n 0.00477804f $X=12.455 $Y=1.26 $X2=0
+ $Y2=0
cc_912 N_A_1746_137#_c_1220_n N_Q_N_c_1906_n 0.00894766f $X=11.88 $Y=2.2 $X2=0
+ $Y2=0
cc_913 N_A_1746_137#_c_1209_n N_Q_N_c_1906_n 0.0227977f $X=11.96 $Y=1.35 $X2=0
+ $Y2=0
cc_914 N_A_1746_137#_c_1211_n N_Q_N_c_1906_n 0.00119022f $X=11.96 $Y=1.26 $X2=0
+ $Y2=0
cc_915 N_A_1746_137#_c_1212_n N_Q_N_c_1906_n 0.00375693f $X=11.96 $Y=1.185 $X2=0
+ $Y2=0
cc_916 N_A_1746_137#_c_1201_n N_Q_N_c_1927_n 0.00671124f $X=12.46 $Y=1.185 $X2=0
+ $Y2=0
cc_917 N_A_1746_137#_c_1212_n N_Q_N_c_1927_n 0.00645722f $X=11.96 $Y=1.185 $X2=0
+ $Y2=0
cc_918 N_A_1746_137#_M1006_g N_Q_c_1943_n 2.83548e-19 $X=13.45 $Y=2.155 $X2=0
+ $Y2=0
cc_919 N_A_1746_137#_c_1197_n N_VGND_c_1980_n 0.00673404f $X=8.805 $Y=1.31 $X2=0
+ $Y2=0
cc_920 N_A_1746_137#_c_1209_n N_VGND_c_1981_n 0.0083854f $X=11.96 $Y=1.35 $X2=0
+ $Y2=0
cc_921 N_A_1746_137#_c_1211_n N_VGND_c_1981_n 8.03164e-19 $X=11.96 $Y=1.26 $X2=0
+ $Y2=0
cc_922 N_A_1746_137#_c_1212_n N_VGND_c_1981_n 0.00328271f $X=11.96 $Y=1.185
+ $X2=0 $Y2=0
cc_923 N_A_1746_137#_c_1201_n N_VGND_c_1982_n 0.00800849f $X=12.46 $Y=1.185
+ $X2=0 $Y2=0
cc_924 N_A_1746_137#_c_1202_n N_VGND_c_1982_n 0.00619922f $X=13.375 $Y=1.26
+ $X2=0 $Y2=0
cc_925 N_A_1746_137#_c_1203_n N_VGND_c_1982_n 0.00359522f $X=13.45 $Y=1.185
+ $X2=0 $Y2=0
cc_926 N_A_1746_137#_c_1203_n N_VGND_c_1983_n 0.00546662f $X=13.45 $Y=1.185
+ $X2=0 $Y2=0
cc_927 N_A_1746_137#_c_1201_n N_VGND_c_1992_n 0.00549284f $X=12.46 $Y=1.185
+ $X2=0 $Y2=0
cc_928 N_A_1746_137#_c_1212_n N_VGND_c_1992_n 0.00549284f $X=11.96 $Y=1.185
+ $X2=0 $Y2=0
cc_929 N_A_1746_137#_c_1203_n N_VGND_c_1993_n 0.00385415f $X=13.45 $Y=1.185
+ $X2=0 $Y2=0
cc_930 N_A_1746_137#_c_1197_n N_VGND_c_2001_n 9.72468e-19 $X=8.805 $Y=1.31 $X2=0
+ $Y2=0
cc_931 N_A_1746_137#_c_1201_n N_VGND_c_2001_n 0.0110929f $X=12.46 $Y=1.185 $X2=0
+ $Y2=0
cc_932 N_A_1746_137#_c_1203_n N_VGND_c_2001_n 0.0046122f $X=13.45 $Y=1.185 $X2=0
+ $Y2=0
cc_933 N_A_1746_137#_c_1212_n N_VGND_c_2001_n 0.00999943f $X=11.96 $Y=1.185
+ $X2=0 $Y2=0
cc_934 N_A_1746_137#_c_1251_p N_A_1911_119#_c_2148_n 0.0182563f $X=10.22 $Y=0.89
+ $X2=0 $Y2=0
cc_935 N_A_1746_137#_M1004_d N_A_1911_119#_c_2149_n 0.00597944f $X=10 $Y=0.595
+ $X2=0 $Y2=0
cc_936 N_A_1746_137#_c_1251_p N_A_1911_119#_c_2149_n 0.0200452f $X=10.22 $Y=0.89
+ $X2=0 $Y2=0
cc_937 N_A_1746_137#_c_1251_p N_A_1911_119#_c_2151_n 0.00255071f $X=10.22
+ $Y=0.89 $X2=0 $Y2=0
cc_938 N_A_1542_428#_c_1375_n N_A_1191_21#_c_1472_n 0.00881791f $X=9.925
+ $Y=1.345 $X2=0 $Y2=0
cc_939 N_A_1542_428#_c_1376_n N_A_1191_21#_c_1472_n 0.00666129f $X=8.12 $Y=0.74
+ $X2=0 $Y2=0
cc_940 N_A_1542_428#_c_1375_n N_A_1191_21#_M1038_g 0.0191168f $X=9.925 $Y=1.345
+ $X2=0 $Y2=0
cc_941 N_A_1542_428#_c_1380_n N_A_1191_21#_M1038_g 2.1676e-19 $X=9.955 $Y=1.205
+ $X2=0 $Y2=0
cc_942 N_A_1542_428#_c_1382_n N_A_1191_21#_M1009_g 0.0111297f $X=10.145 $Y=1.915
+ $X2=0 $Y2=0
cc_943 N_A_1542_428#_c_1383_n N_A_1191_21#_M1009_g 0.0710987f $X=10.145 $Y=2.065
+ $X2=0 $Y2=0
cc_944 N_A_1542_428#_c_1380_n N_A_1191_21#_c_1476_n 2.90401e-19 $X=9.955
+ $Y=1.205 $X2=0 $Y2=0
cc_945 N_A_1542_428#_c_1381_n N_A_1191_21#_c_1476_n 0.0175267f $X=10.125 $Y=1.51
+ $X2=0 $Y2=0
cc_946 N_A_1542_428#_c_1383_n N_VPWR_c_1702_n 0.00186217f $X=10.145 $Y=2.065
+ $X2=0 $Y2=0
cc_947 N_A_1542_428#_c_1383_n N_VPWR_c_1714_n 0.00449508f $X=10.145 $Y=2.065
+ $X2=0 $Y2=0
cc_948 N_A_1542_428#_c_1383_n N_VPWR_c_1695_n 0.00854629f $X=10.145 $Y=2.065
+ $X2=0 $Y2=0
cc_949 N_A_1542_428#_c_1377_n N_VGND_M1000_d 0.00821569f $X=9.785 $Y=1.205 $X2=0
+ $Y2=0
cc_950 N_A_1542_428#_c_1377_n N_VGND_c_1980_n 0.0243215f $X=9.785 $Y=1.205 $X2=0
+ $Y2=0
cc_951 N_A_1542_428#_c_1376_n N_VGND_c_1990_n 0.00756512f $X=8.12 $Y=0.74 $X2=0
+ $Y2=0
cc_952 N_A_1542_428#_c_1376_n N_VGND_c_2001_n 0.00911172f $X=8.12 $Y=0.74 $X2=0
+ $Y2=0
cc_953 N_A_1542_428#_c_1377_n A_1698_163# 0.0048076f $X=9.785 $Y=1.205 $X2=-0.19
+ $Y2=-0.245
cc_954 N_A_1542_428#_c_1377_n N_A_1911_119#_M1031_d 0.00187279f $X=9.785
+ $Y=1.205 $X2=-0.19 $Y2=-0.245
cc_955 N_A_1542_428#_c_1375_n N_A_1911_119#_c_2148_n 0.0092507f $X=9.925
+ $Y=1.345 $X2=0 $Y2=0
cc_956 N_A_1542_428#_c_1377_n N_A_1911_119#_c_2148_n 0.014057f $X=9.785 $Y=1.205
+ $X2=0 $Y2=0
cc_957 N_A_1542_428#_c_1380_n N_A_1911_119#_c_2148_n 0.00254886f $X=9.955
+ $Y=1.205 $X2=0 $Y2=0
cc_958 N_A_1542_428#_c_1375_n N_A_1911_119#_c_2149_n 0.00311859f $X=9.925
+ $Y=1.345 $X2=0 $Y2=0
cc_959 N_A_1191_21#_c_1475_n N_RESET_B_c_1581_n 0.0047176f $X=10.82 $Y=1.51
+ $X2=0 $Y2=0
cc_960 N_A_1191_21#_c_1477_n N_RESET_B_c_1581_n 0.00404524f $X=11.22 $Y=0.915
+ $X2=0 $Y2=0
cc_961 N_A_1191_21#_c_1476_n N_RESET_B_M1026_g 0.0037997f $X=10.82 $Y=1.51 $X2=0
+ $Y2=0
cc_962 N_A_1191_21#_c_1483_n N_RESET_B_M1026_g 0.00124824f $X=10.985 $Y=1.855
+ $X2=0 $Y2=0
cc_963 N_A_1191_21#_c_1484_n N_RESET_B_M1026_g 0.00575014f $X=11.295 $Y=1.855
+ $X2=0 $Y2=0
cc_964 N_A_1191_21#_c_1479_n N_RESET_B_M1001_g 0.0085564f $X=11.305 $Y=0.47
+ $X2=0 $Y2=0
cc_965 N_A_1191_21#_M1038_g N_RESET_B_c_1584_n 0.00600071f $X=10.515 $Y=0.66
+ $X2=0 $Y2=0
cc_966 N_A_1191_21#_c_1477_n N_RESET_B_c_1584_n 0.00609609f $X=11.22 $Y=0.915
+ $X2=0 $Y2=0
cc_967 N_A_1191_21#_c_1479_n N_RESET_B_c_1584_n 0.00625706f $X=11.305 $Y=0.47
+ $X2=0 $Y2=0
cc_968 N_A_1191_21#_c_1475_n N_RESET_B_c_1585_n 0.0260253f $X=10.82 $Y=1.51
+ $X2=0 $Y2=0
cc_969 N_A_1191_21#_c_1476_n N_RESET_B_c_1585_n 0.00109089f $X=10.82 $Y=1.51
+ $X2=0 $Y2=0
cc_970 N_A_1191_21#_c_1477_n N_RESET_B_c_1585_n 0.0237062f $X=11.22 $Y=0.915
+ $X2=0 $Y2=0
cc_971 N_A_1191_21#_c_1484_n N_RESET_B_c_1585_n 0.0225327f $X=11.295 $Y=1.855
+ $X2=0 $Y2=0
cc_972 N_A_1191_21#_c_1475_n N_RESET_B_c_1586_n 8.01768e-19 $X=10.82 $Y=1.51
+ $X2=0 $Y2=0
cc_973 N_A_1191_21#_c_1476_n N_RESET_B_c_1586_n 0.00881529f $X=10.82 $Y=1.51
+ $X2=0 $Y2=0
cc_974 N_A_1191_21#_c_1477_n N_RESET_B_c_1586_n 6.08141e-19 $X=11.22 $Y=0.915
+ $X2=0 $Y2=0
cc_975 N_A_1191_21#_c_1484_n N_RESET_B_c_1586_n 0.00522227f $X=11.295 $Y=1.855
+ $X2=0 $Y2=0
cc_976 N_A_1191_21#_M1003_g N_VPWR_c_1700_n 0.0273542f $X=6.03 $Y=0.955 $X2=0
+ $Y2=0
cc_977 N_A_1191_21#_M1009_g N_VPWR_c_1702_n 0.0134608f $X=10.525 $Y=2.56 $X2=0
+ $Y2=0
cc_978 N_A_1191_21#_M1009_g N_VPWR_c_1714_n 0.00396895f $X=10.525 $Y=2.56 $X2=0
+ $Y2=0
cc_979 N_A_1191_21#_M1003_g N_VPWR_c_1695_n 9.39239e-19 $X=6.03 $Y=0.955 $X2=0
+ $Y2=0
cc_980 N_A_1191_21#_M1009_g N_VPWR_c_1695_n 0.0076824f $X=10.525 $Y=2.56 $X2=0
+ $Y2=0
cc_981 N_A_1191_21#_c_1472_n N_VGND_c_1979_n 0.0211465f $X=10.44 $Y=0.18 $X2=0
+ $Y2=0
cc_982 N_A_1191_21#_c_1472_n N_VGND_c_1980_n 0.0260404f $X=10.44 $Y=0.18 $X2=0
+ $Y2=0
cc_983 N_A_1191_21#_c_1477_n N_VGND_c_1981_n 0.0136306f $X=11.22 $Y=0.915 $X2=0
+ $Y2=0
cc_984 N_A_1191_21#_c_1479_n N_VGND_c_1981_n 0.0260048f $X=11.305 $Y=0.47 $X2=0
+ $Y2=0
cc_985 N_A_1191_21#_c_1473_n N_VGND_c_1989_n 0.0219031f $X=6.105 $Y=0.18 $X2=0
+ $Y2=0
cc_986 N_A_1191_21#_c_1472_n N_VGND_c_1990_n 0.0642068f $X=10.44 $Y=0.18 $X2=0
+ $Y2=0
cc_987 N_A_1191_21#_c_1472_n N_VGND_c_1991_n 0.0283875f $X=10.44 $Y=0.18 $X2=0
+ $Y2=0
cc_988 N_A_1191_21#_c_1479_n N_VGND_c_1991_n 0.0144775f $X=11.305 $Y=0.47 $X2=0
+ $Y2=0
cc_989 N_A_1191_21#_M1001_s N_VGND_c_2001_n 0.00271024f $X=11.16 $Y=0.235 $X2=0
+ $Y2=0
cc_990 N_A_1191_21#_c_1472_n N_VGND_c_2001_n 0.139555f $X=10.44 $Y=0.18 $X2=0
+ $Y2=0
cc_991 N_A_1191_21#_c_1473_n N_VGND_c_2001_n 0.0054647f $X=6.105 $Y=0.18 $X2=0
+ $Y2=0
cc_992 N_A_1191_21#_c_1477_n N_VGND_c_2001_n 0.00816097f $X=11.22 $Y=0.915 $X2=0
+ $Y2=0
cc_993 N_A_1191_21#_c_1478_n N_VGND_c_2001_n 0.00372917f $X=10.985 $Y=0.915
+ $X2=0 $Y2=0
cc_994 N_A_1191_21#_c_1479_n N_VGND_c_2001_n 0.00948536f $X=11.305 $Y=0.47 $X2=0
+ $Y2=0
cc_995 N_A_1191_21#_M1003_g N_A_1018_60#_c_2123_n 0.0107997f $X=6.03 $Y=0.955
+ $X2=0 $Y2=0
cc_996 N_A_1191_21#_M1003_g N_A_1018_60#_c_2124_n 7.84604e-19 $X=6.03 $Y=0.955
+ $X2=0 $Y2=0
cc_997 N_A_1191_21#_c_1478_n N_A_1911_119#_M1038_d 0.00576772f $X=10.985
+ $Y=0.915 $X2=0 $Y2=0
cc_998 N_A_1191_21#_M1038_g N_A_1911_119#_c_2148_n 0.00164244f $X=10.515 $Y=0.66
+ $X2=0 $Y2=0
cc_999 N_A_1191_21#_c_1472_n N_A_1911_119#_c_2149_n 0.00902132f $X=10.44 $Y=0.18
+ $X2=0 $Y2=0
cc_1000 N_A_1191_21#_M1038_g N_A_1911_119#_c_2149_n 0.0144598f $X=10.515 $Y=0.66
+ $X2=0 $Y2=0
cc_1001 N_A_1191_21#_c_1472_n N_A_1911_119#_c_2150_n 0.00752773f $X=10.44
+ $Y=0.18 $X2=0 $Y2=0
cc_1002 N_A_1191_21#_M1038_g N_A_1911_119#_c_2151_n 6.13408e-19 $X=10.515
+ $Y=0.66 $X2=0 $Y2=0
cc_1003 N_A_1191_21#_c_1476_n N_A_1911_119#_c_2151_n 6.84168e-19 $X=10.82
+ $Y=1.51 $X2=0 $Y2=0
cc_1004 N_A_1191_21#_c_1478_n N_A_1911_119#_c_2151_n 0.0199813f $X=10.985
+ $Y=0.915 $X2=0 $Y2=0
cc_1005 N_A_1191_21#_c_1479_n N_A_1911_119#_c_2151_n 0.0194391f $X=11.305
+ $Y=0.47 $X2=0 $Y2=0
cc_1006 N_RESET_B_M1026_g N_VPWR_c_1695_n 0.00381575f $X=11.51 $Y=2.03 $X2=0
+ $Y2=0
cc_1007 N_RESET_B_M1001_g N_VGND_c_1981_n 0.0077437f $X=11.52 $Y=0.445 $X2=0
+ $Y2=0
cc_1008 N_RESET_B_M1001_g N_VGND_c_1991_n 0.00549284f $X=11.52 $Y=0.445 $X2=0
+ $Y2=0
cc_1009 N_RESET_B_M1001_g N_VGND_c_2001_n 0.011593f $X=11.52 $Y=0.445 $X2=0
+ $Y2=0
cc_1010 N_RESET_B_M1001_g N_A_1911_119#_c_2151_n 8.51193e-19 $X=11.52 $Y=0.445
+ $X2=0 $Y2=0
cc_1011 N_A_2618_131#_c_1626_n N_VPWR_c_1704_n 0.0531549f $X=13.235 $Y=1.98
+ $X2=0 $Y2=0
cc_1012 N_A_2618_131#_M1007_g N_VPWR_c_1705_n 0.00698192f $X=13.96 $Y=2.465
+ $X2=0 $Y2=0
cc_1013 N_A_2618_131#_c_1626_n N_VPWR_c_1705_n 0.025828f $X=13.235 $Y=1.98 $X2=0
+ $Y2=0
cc_1014 N_A_2618_131#_c_1627_n N_VPWR_c_1705_n 0.0186319f $X=13.93 $Y=1.44 $X2=0
+ $Y2=0
cc_1015 N_A_2618_131#_c_1629_n N_VPWR_c_1705_n 0.00146036f $X=13.93 $Y=1.35
+ $X2=0 $Y2=0
cc_1016 N_A_2618_131#_M1027_g N_VPWR_c_1707_n 0.0094801f $X=14.39 $Y=2.465 $X2=0
+ $Y2=0
cc_1017 N_A_2618_131#_M1007_g N_VPWR_c_1718_n 0.00549284f $X=13.96 $Y=2.465
+ $X2=0 $Y2=0
cc_1018 N_A_2618_131#_M1027_g N_VPWR_c_1718_n 0.00549284f $X=14.39 $Y=2.465
+ $X2=0 $Y2=0
cc_1019 N_A_2618_131#_M1007_g N_VPWR_c_1695_n 0.0110929f $X=13.96 $Y=2.465 $X2=0
+ $Y2=0
cc_1020 N_A_2618_131#_M1027_g N_VPWR_c_1695_n 0.0107398f $X=14.39 $Y=2.465 $X2=0
+ $Y2=0
cc_1021 N_A_2618_131#_c_1626_n N_VPWR_c_1695_n 0.0128958f $X=13.235 $Y=1.98
+ $X2=0 $Y2=0
cc_1022 N_A_2618_131#_c_1625_n N_Q_N_c_1906_n 0.0044826f $X=13.235 $Y=0.865
+ $X2=0 $Y2=0
cc_1023 N_A_2618_131#_c_1626_n N_Q_N_c_1906_n 0.00228272f $X=13.235 $Y=1.98
+ $X2=0 $Y2=0
cc_1024 N_A_2618_131#_c_1628_n N_Q_N_c_1906_n 0.00927367f $X=13.235 $Y=1.44
+ $X2=0 $Y2=0
cc_1025 N_A_2618_131#_M1007_g N_Q_c_1945_n 0.0137061f $X=13.96 $Y=2.465 $X2=0
+ $Y2=0
cc_1026 N_A_2618_131#_M1027_g N_Q_c_1945_n 0.0197981f $X=14.39 $Y=2.465 $X2=0
+ $Y2=0
cc_1027 N_A_2618_131#_M1018_g N_Q_c_1940_n 0.00246747f $X=13.96 $Y=0.655 $X2=0
+ $Y2=0
cc_1028 N_A_2618_131#_M1007_g N_Q_c_1940_n 0.00246747f $X=13.96 $Y=2.465 $X2=0
+ $Y2=0
cc_1029 N_A_2618_131#_c_1621_n N_Q_c_1940_n 0.00358637f $X=14.315 $Y=1.35 $X2=0
+ $Y2=0
cc_1030 N_A_2618_131#_M1033_g N_Q_c_1940_n 0.0101468f $X=14.39 $Y=0.655 $X2=0
+ $Y2=0
cc_1031 N_A_2618_131#_M1027_g N_Q_c_1940_n 0.0194308f $X=14.39 $Y=2.465 $X2=0
+ $Y2=0
cc_1032 N_A_2618_131#_c_1624_n N_Q_c_1940_n 0.0073295f $X=14.39 $Y=1.35 $X2=0
+ $Y2=0
cc_1033 N_A_2618_131#_c_1627_n N_Q_c_1940_n 0.0245348f $X=13.93 $Y=1.44 $X2=0
+ $Y2=0
cc_1034 N_A_2618_131#_c_1629_n N_Q_c_1940_n 5.36405e-19 $X=13.93 $Y=1.35 $X2=0
+ $Y2=0
cc_1035 N_A_2618_131#_M1007_g N_Q_c_1943_n 0.00298817f $X=13.96 $Y=2.465 $X2=0
+ $Y2=0
cc_1036 N_A_2618_131#_c_1621_n N_Q_c_1943_n 0.00650242f $X=14.315 $Y=1.35 $X2=0
+ $Y2=0
cc_1037 N_A_2618_131#_M1027_g N_Q_c_1943_n 0.0150137f $X=14.39 $Y=2.465 $X2=0
+ $Y2=0
cc_1038 N_A_2618_131#_c_1626_n N_Q_c_1943_n 7.97843e-19 $X=13.235 $Y=1.98 $X2=0
+ $Y2=0
cc_1039 N_A_2618_131#_c_1627_n N_Q_c_1943_n 0.00667629f $X=13.93 $Y=1.44 $X2=0
+ $Y2=0
cc_1040 N_A_2618_131#_c_1629_n N_Q_c_1943_n 0.00162496f $X=13.93 $Y=1.35 $X2=0
+ $Y2=0
cc_1041 N_A_2618_131#_M1018_g Q 0.00236686f $X=13.96 $Y=0.655 $X2=0 $Y2=0
cc_1042 N_A_2618_131#_c_1621_n Q 0.00406666f $X=14.315 $Y=1.35 $X2=0 $Y2=0
cc_1043 N_A_2618_131#_M1033_g Q 0.0146525f $X=14.39 $Y=0.655 $X2=0 $Y2=0
cc_1044 N_A_2618_131#_c_1627_n Q 0.00667752f $X=13.93 $Y=1.44 $X2=0 $Y2=0
cc_1045 N_A_2618_131#_M1018_g N_Q_c_1965_n 0.00854555f $X=13.96 $Y=0.655 $X2=0
+ $Y2=0
cc_1046 N_A_2618_131#_M1033_g N_Q_c_1965_n 0.0145269f $X=14.39 $Y=0.655 $X2=0
+ $Y2=0
cc_1047 N_A_2618_131#_c_1625_n N_VGND_c_1982_n 0.0303742f $X=13.235 $Y=0.865
+ $X2=0 $Y2=0
cc_1048 N_A_2618_131#_M1018_g N_VGND_c_1983_n 0.00550224f $X=13.96 $Y=0.655
+ $X2=0 $Y2=0
cc_1049 N_A_2618_131#_c_1625_n N_VGND_c_1983_n 0.0179429f $X=13.235 $Y=0.865
+ $X2=0 $Y2=0
cc_1050 N_A_2618_131#_c_1627_n N_VGND_c_1983_n 0.0208003f $X=13.93 $Y=1.44 $X2=0
+ $Y2=0
cc_1051 N_A_2618_131#_c_1629_n N_VGND_c_1983_n 0.00148357f $X=13.93 $Y=1.35
+ $X2=0 $Y2=0
cc_1052 N_A_2618_131#_M1033_g N_VGND_c_1985_n 0.00677163f $X=14.39 $Y=0.655
+ $X2=0 $Y2=0
cc_1053 N_A_2618_131#_c_1625_n N_VGND_c_1993_n 0.00658678f $X=13.235 $Y=0.865
+ $X2=0 $Y2=0
cc_1054 N_A_2618_131#_M1018_g N_VGND_c_1994_n 0.00549284f $X=13.96 $Y=0.655
+ $X2=0 $Y2=0
cc_1055 N_A_2618_131#_M1033_g N_VGND_c_1994_n 0.00549284f $X=14.39 $Y=0.655
+ $X2=0 $Y2=0
cc_1056 N_A_2618_131#_M1018_g N_VGND_c_2001_n 0.0110929f $X=13.96 $Y=0.655 $X2=0
+ $Y2=0
cc_1057 N_A_2618_131#_M1033_g N_VGND_c_2001_n 0.0109199f $X=14.39 $Y=0.655 $X2=0
+ $Y2=0
cc_1058 N_A_2618_131#_c_1625_n N_VGND_c_2001_n 0.00992454f $X=13.235 $Y=0.865
+ $X2=0 $Y2=0
cc_1059 N_VPWR_c_1698_n N_A_463_449#_c_1853_n 0.0232432f $X=1.885 $Y=2.39 $X2=0
+ $Y2=0
cc_1060 N_VPWR_c_1710_n N_A_463_449#_c_1853_n 0.006147f $X=4.63 $Y=3.33 $X2=0
+ $Y2=0
cc_1061 N_VPWR_c_1695_n N_A_463_449#_c_1853_n 0.018109f $X=14.64 $Y=3.33 $X2=0
+ $Y2=0
cc_1062 N_VPWR_c_1703_n N_Q_N_c_1908_n 0.0165025f $X=11.805 $Y=2.77 $X2=0 $Y2=0
cc_1063 N_VPWR_c_1716_n N_Q_N_c_1908_n 0.0118895f $X=12.59 $Y=3.33 $X2=0 $Y2=0
cc_1064 N_VPWR_c_1695_n N_Q_N_c_1908_n 0.00942244f $X=14.64 $Y=3.33 $X2=0 $Y2=0
cc_1065 N_VPWR_c_1704_n N_Q_N_c_1906_n 0.0928358f $X=12.675 $Y=1.855 $X2=0 $Y2=0
cc_1066 N_VPWR_c_1695_n N_Q_M1007_d 0.00223819f $X=14.64 $Y=3.33 $X2=0 $Y2=0
cc_1067 N_VPWR_c_1718_n N_Q_c_1945_n 0.0177952f $X=14.52 $Y=3.33 $X2=0 $Y2=0
cc_1068 N_VPWR_c_1695_n N_Q_c_1945_n 0.0123247f $X=14.64 $Y=3.33 $X2=0 $Y2=0
cc_1069 N_VPWR_c_1705_n N_Q_c_1943_n 0.0457104f $X=13.745 $Y=1.98 $X2=0 $Y2=0
cc_1070 N_VPWR_c_1704_n N_VGND_c_1982_n 0.00958683f $X=12.675 $Y=1.855 $X2=0
+ $Y2=0
cc_1071 N_A_463_449#_c_1849_n N_VGND_c_1977_n 0.0139674f $X=2.61 $Y=0.805 $X2=0
+ $Y2=0
cc_1072 N_A_463_449#_c_1849_n N_VGND_c_1986_n 0.00743798f $X=2.61 $Y=0.805 $X2=0
+ $Y2=0
cc_1073 N_A_463_449#_c_1849_n N_VGND_c_2001_n 0.00904485f $X=2.61 $Y=0.805 $X2=0
+ $Y2=0
cc_1074 N_Q_N_c_1927_n N_VGND_c_1982_n 0.0300958f $X=12.245 $Y=0.43 $X2=0 $Y2=0
cc_1075 N_Q_N_c_1927_n N_VGND_c_1992_n 0.0177952f $X=12.245 $Y=0.43 $X2=0 $Y2=0
cc_1076 N_Q_N_M1008_d N_VGND_c_2001_n 0.00223819f $X=12.105 $Y=0.235 $X2=0 $Y2=0
cc_1077 N_Q_N_c_1927_n N_VGND_c_2001_n 0.0123247f $X=12.245 $Y=0.43 $X2=0 $Y2=0
cc_1078 N_Q_c_1965_n N_VGND_c_1983_n 0.0307034f $X=14.175 $Y=0.43 $X2=0 $Y2=0
cc_1079 N_Q_c_1965_n N_VGND_c_1994_n 0.0177952f $X=14.175 $Y=0.43 $X2=0 $Y2=0
cc_1080 N_Q_M1018_d N_VGND_c_2001_n 0.00223819f $X=14.035 $Y=0.235 $X2=0 $Y2=0
cc_1081 N_Q_c_1965_n N_VGND_c_2001_n 0.0123247f $X=14.175 $Y=0.43 $X2=0 $Y2=0
cc_1082 N_VGND_c_1980_n N_A_1911_119#_c_2148_n 0.0245387f $X=9.2 $Y=0.755 $X2=0
+ $Y2=0
cc_1083 N_VGND_c_1991_n N_A_1911_119#_c_2149_n 0.0468271f $X=11.65 $Y=0 $X2=0
+ $Y2=0
cc_1084 N_VGND_c_2001_n N_A_1911_119#_c_2149_n 0.0261772f $X=14.64 $Y=0 $X2=0
+ $Y2=0
cc_1085 N_VGND_c_1980_n N_A_1911_119#_c_2150_n 0.0144411f $X=9.2 $Y=0.755 $X2=0
+ $Y2=0
cc_1086 N_VGND_c_1991_n N_A_1911_119#_c_2150_n 0.0222284f $X=11.65 $Y=0 $X2=0
+ $Y2=0
cc_1087 N_VGND_c_2001_n N_A_1911_119#_c_2150_n 0.0114499f $X=14.64 $Y=0 $X2=0
+ $Y2=0
cc_1088 N_VGND_c_1991_n N_A_1911_119#_c_2151_n 0.0160316f $X=11.65 $Y=0 $X2=0
+ $Y2=0
cc_1089 N_VGND_c_2001_n N_A_1911_119#_c_2151_n 0.00945436f $X=14.64 $Y=0 $X2=0
+ $Y2=0
