* File: sky130_fd_sc_lp__fahcin_1.pxi.spice
* Created: Fri Aug 28 10:35:37 2020
* 
x_PM_SKY130_FD_SC_LP__FAHCIN_1%A N_A_M1016_g N_A_M1012_g A N_A_c_250_n
+ N_A_c_251_n PM_SKY130_FD_SC_LP__FAHCIN_1%A
x_PM_SKY130_FD_SC_LP__FAHCIN_1%A_29_47# N_A_29_47#_M1016_s N_A_29_47#_M1026_d
+ N_A_29_47#_M1012_s N_A_29_47#_M1002_d N_A_29_47#_M1005_g N_A_29_47#_M1007_g
+ N_A_29_47#_c_285_n N_A_29_47#_c_286_n N_A_29_47#_c_287_n N_A_29_47#_c_300_n
+ N_A_29_47#_c_301_n N_A_29_47#_c_288_n N_A_29_47#_c_316_n N_A_29_47#_c_289_n
+ N_A_29_47#_c_290_n N_A_29_47#_c_303_n N_A_29_47#_c_291_n N_A_29_47#_c_292_n
+ N_A_29_47#_c_304_n N_A_29_47#_c_305_n N_A_29_47#_c_306_n N_A_29_47#_c_293_n
+ N_A_29_47#_c_294_n N_A_29_47#_c_295_n N_A_29_47#_c_308_n N_A_29_47#_c_296_n
+ PM_SKY130_FD_SC_LP__FAHCIN_1%A_29_47#
x_PM_SKY130_FD_SC_LP__FAHCIN_1%A_439_47# N_A_439_47#_M1004_s N_A_439_47#_M1013_s
+ N_A_439_47#_M1026_g N_A_439_47#_M1021_g N_A_439_47#_M1002_g
+ N_A_439_47#_c_397_n N_A_439_47#_M1009_g N_A_439_47#_c_398_n
+ N_A_439_47#_M1019_g N_A_439_47#_c_400_n N_A_439_47#_M1015_g
+ N_A_439_47#_c_401_n N_A_439_47#_c_402_n N_A_439_47#_c_403_n
+ N_A_439_47#_c_404_n N_A_439_47#_c_405_n N_A_439_47#_c_406_n
+ N_A_439_47#_c_407_n N_A_439_47#_c_408_n N_A_439_47#_c_409_n
+ N_A_439_47#_c_454_p N_A_439_47#_c_410_n N_A_439_47#_c_411_n
+ N_A_439_47#_c_419_n N_A_439_47#_c_412_n PM_SKY130_FD_SC_LP__FAHCIN_1%A_439_47#
x_PM_SKY130_FD_SC_LP__FAHCIN_1%B N_B_c_575_n N_B_M1006_g N_B_M1010_g N_B_c_576_n
+ N_B_c_577_n N_B_c_588_n N_B_c_589_n N_B_c_590_n N_B_M1014_g N_B_M1000_g
+ N_B_c_591_n N_B_c_579_n N_B_c_592_n N_B_c_580_n N_B_M1004_g N_B_M1013_g
+ N_B_c_594_n N_B_c_582_n N_B_c_583_n N_B_c_584_n N_B_c_585_n B
+ PM_SKY130_FD_SC_LP__FAHCIN_1%B
x_PM_SKY130_FD_SC_LP__FAHCIN_1%A_555_73# N_A_555_73#_M1006_d N_A_555_73#_M1010_d
+ N_A_555_73#_M1030_g N_A_555_73#_M1008_g N_A_555_73#_M1031_g
+ N_A_555_73#_M1020_g N_A_555_73#_c_710_n N_A_555_73#_c_742_n
+ N_A_555_73#_c_711_n N_A_555_73#_c_743_n N_A_555_73#_c_726_n
+ N_A_555_73#_c_727_n N_A_555_73#_c_728_n N_A_555_73#_c_761_n
+ N_A_555_73#_c_762_n N_A_555_73#_c_765_n N_A_555_73#_c_712_n
+ N_A_555_73#_c_713_n N_A_555_73#_c_731_n N_A_555_73#_c_732_n
+ N_A_555_73#_c_733_n N_A_555_73#_c_734_n N_A_555_73#_c_714_n
+ N_A_555_73#_c_715_n N_A_555_73#_c_735_n N_A_555_73#_c_736_n
+ N_A_555_73#_c_716_n N_A_555_73#_c_717_n N_A_555_73#_c_718_n
+ N_A_555_73#_c_719_n N_A_555_73#_c_720_n N_A_555_73#_c_721_n
+ N_A_555_73#_c_739_n N_A_555_73#_c_722_n N_A_555_73#_c_741_n
+ PM_SKY130_FD_SC_LP__FAHCIN_1%A_555_73#
x_PM_SKY130_FD_SC_LP__FAHCIN_1%A_364_73# N_A_364_73#_M1026_s N_A_364_73#_M1000_d
+ N_A_364_73#_M1021_s N_A_364_73#_M1014_d N_A_364_73#_c_959_n
+ N_A_364_73#_M1027_g N_A_364_73#_c_960_n N_A_364_73#_c_961_n
+ N_A_364_73#_c_962_n N_A_364_73#_c_981_n N_A_364_73#_c_982_n
+ N_A_364_73#_c_983_n N_A_364_73#_M1029_g N_A_364_73#_M1024_g
+ N_A_364_73#_M1028_g N_A_364_73#_c_964_n N_A_364_73#_c_986_n
+ N_A_364_73#_c_965_n N_A_364_73#_c_966_n N_A_364_73#_c_967_n
+ N_A_364_73#_c_968_n N_A_364_73#_c_969_n N_A_364_73#_c_970_n
+ N_A_364_73#_c_971_n N_A_364_73#_c_972_n N_A_364_73#_c_973_n
+ N_A_364_73#_c_974_n N_A_364_73#_c_975_n N_A_364_73#_c_976_n
+ N_A_364_73#_c_977_n N_A_364_73#_c_978_n N_A_364_73#_c_979_n
+ PM_SKY130_FD_SC_LP__FAHCIN_1%A_364_73#
x_PM_SKY130_FD_SC_LP__FAHCIN_1%CIN N_CIN_M1003_g N_CIN_c_1202_n N_CIN_M1011_g
+ N_CIN_c_1203_n N_CIN_M1023_g N_CIN_c_1205_n N_CIN_M1022_g CIN
+ PM_SKY130_FD_SC_LP__FAHCIN_1%CIN
x_PM_SKY130_FD_SC_LP__FAHCIN_1%A_1774_367# N_A_1774_367#_M1022_d
+ N_A_1774_367#_M1023_d N_A_1774_367#_M1024_d N_A_1774_367#_M1017_g
+ N_A_1774_367#_M1025_g N_A_1774_367#_c_1271_n N_A_1774_367#_c_1282_n
+ N_A_1774_367#_c_1272_n N_A_1774_367#_c_1273_n N_A_1774_367#_c_1274_n
+ N_A_1774_367#_c_1266_n N_A_1774_367#_c_1267_n N_A_1774_367#_c_1276_n
+ N_A_1774_367#_c_1277_n N_A_1774_367#_c_1268_n N_A_1774_367#_c_1269_n
+ PM_SKY130_FD_SC_LP__FAHCIN_1%A_1774_367#
x_PM_SKY130_FD_SC_LP__FAHCIN_1%A_1926_135# N_A_1926_135#_M1031_d
+ N_A_1926_135#_M1020_d N_A_1926_135#_c_1363_n N_A_1926_135#_M1001_g
+ N_A_1926_135#_M1018_g N_A_1926_135#_c_1364_n N_A_1926_135#_c_1380_n
+ N_A_1926_135#_c_1365_n N_A_1926_135#_c_1366_n N_A_1926_135#_c_1367_n
+ N_A_1926_135#_c_1368_n N_A_1926_135#_c_1369_n N_A_1926_135#_c_1370_n
+ N_A_1926_135#_c_1389_n N_A_1926_135#_c_1371_n N_A_1926_135#_c_1372_n
+ PM_SKY130_FD_SC_LP__FAHCIN_1%A_1926_135#
x_PM_SKY130_FD_SC_LP__FAHCIN_1%VPWR N_VPWR_M1012_d N_VPWR_M1013_d N_VPWR_M1003_d
+ N_VPWR_M1025_d N_VPWR_c_1461_n N_VPWR_c_1462_n N_VPWR_c_1463_n N_VPWR_c_1464_n
+ N_VPWR_c_1465_n N_VPWR_c_1466_n N_VPWR_c_1467_n N_VPWR_c_1468_n VPWR
+ N_VPWR_c_1469_n N_VPWR_c_1470_n N_VPWR_c_1471_n N_VPWR_c_1460_n
+ N_VPWR_c_1473_n N_VPWR_c_1474_n PM_SKY130_FD_SC_LP__FAHCIN_1%VPWR
x_PM_SKY130_FD_SC_LP__FAHCIN_1%A_256_87# N_A_256_87#_M1005_d N_A_256_87#_M1009_d
+ N_A_256_87#_M1007_d N_A_256_87#_M1021_d N_A_256_87#_c_1575_n
+ N_A_256_87#_c_1568_n N_A_256_87#_c_1576_n N_A_256_87#_c_1577_n
+ N_A_256_87#_c_1569_n N_A_256_87#_c_1598_n N_A_256_87#_c_1570_n
+ N_A_256_87#_c_1571_n N_A_256_87#_c_1572_n N_A_256_87#_c_1573_n
+ N_A_256_87#_c_1574_n PM_SKY130_FD_SC_LP__FAHCIN_1%A_256_87#
x_PM_SKY130_FD_SC_LP__FAHCIN_1%A_1152_389# N_A_1152_389#_M1015_d
+ N_A_1152_389#_M1019_d N_A_1152_389#_c_1651_n N_A_1152_389#_c_1652_n
+ N_A_1152_389#_c_1653_n PM_SKY130_FD_SC_LP__FAHCIN_1%A_1152_389#
x_PM_SKY130_FD_SC_LP__FAHCIN_1%COUT N_COUT_M1027_d N_COUT_M1030_d
+ N_COUT_c_1685_n N_COUT_c_1681_n COUT COUT COUT N_COUT_c_1682_n
+ PM_SKY130_FD_SC_LP__FAHCIN_1%COUT
x_PM_SKY130_FD_SC_LP__FAHCIN_1%A_1500_63# N_A_1500_63#_M1008_d
+ N_A_1500_63#_M1029_d N_A_1500_63#_c_1719_n N_A_1500_63#_c_1721_n
+ N_A_1500_63#_c_1720_n N_A_1500_63#_c_1734_n
+ PM_SKY130_FD_SC_LP__FAHCIN_1%A_1500_63#
x_PM_SKY130_FD_SC_LP__FAHCIN_1%A_1883_395# N_A_1883_395#_M1028_d
+ N_A_1883_395#_M1020_s N_A_1883_395#_M1025_s N_A_1883_395#_c_1757_n
+ N_A_1883_395#_c_1752_n N_A_1883_395#_c_1753_n N_A_1883_395#_c_1758_n
+ N_A_1883_395#_c_1754_n N_A_1883_395#_c_1756_n
+ PM_SKY130_FD_SC_LP__FAHCIN_1%A_1883_395#
x_PM_SKY130_FD_SC_LP__FAHCIN_1%SUM N_SUM_M1001_d N_SUM_M1018_d SUM SUM SUM SUM
+ SUM SUM SUM N_SUM_c_1802_n PM_SKY130_FD_SC_LP__FAHCIN_1%SUM
x_PM_SKY130_FD_SC_LP__FAHCIN_1%VGND N_VGND_M1016_d N_VGND_M1004_d N_VGND_M1011_d
+ N_VGND_M1017_d N_VGND_c_1816_n N_VGND_c_1817_n N_VGND_c_1818_n N_VGND_c_1819_n
+ N_VGND_c_1820_n N_VGND_c_1821_n VGND N_VGND_c_1822_n N_VGND_c_1823_n
+ N_VGND_c_1824_n N_VGND_c_1825_n N_VGND_c_1826_n N_VGND_c_1827_n
+ N_VGND_c_1828_n N_VGND_c_1829_n PM_SKY130_FD_SC_LP__FAHCIN_1%VGND
cc_1 VNB N_A_M1016_g 0.03313f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=0.655
cc_2 VNB N_A_c_250_n 0.0289188f $X=-0.19 $Y=-0.245 $X2=0.625 $Y2=1.51
cc_3 VNB N_A_c_251_n 0.00409837f $X=-0.19 $Y=-0.245 $X2=0.625 $Y2=1.51
cc_4 VNB N_A_29_47#_M1005_g 0.023613f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.675
cc_5 VNB N_A_29_47#_c_285_n 0.0235029f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_6 VNB N_A_29_47#_c_286_n 0.00724895f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_A_29_47#_c_287_n 0.0284857f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_A_29_47#_c_288_n 0.00789792f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A_29_47#_c_289_n 0.00759958f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A_29_47#_c_290_n 0.00164259f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_29_47#_c_291_n 0.0178496f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_12 VNB N_A_29_47#_c_292_n 0.00246543f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_29_47#_c_293_n 0.0136024f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_29_47#_c_294_n 0.0232197f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_29_47#_c_295_n 0.0185776f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_29_47#_c_296_n 0.00239374f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_439_47#_M1026_g 0.04017f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_18 VNB N_A_439_47#_M1021_g 0.0234105f $X=-0.19 $Y=-0.245 $X2=0.625 $Y2=1.51
cc_19 VNB N_A_439_47#_c_397_n 0.0171371f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_439_47#_c_398_n 0.0612879f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_439_47#_M1019_g 0.00297236f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_439_47#_c_400_n 0.0185112f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_439_47#_c_401_n 0.00694327f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_439_47#_c_402_n 9.12604e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_439_47#_c_403_n 0.0351046f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_439_47#_c_404_n 0.00145481f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_A_439_47#_c_405_n 0.0119871f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_A_439_47#_c_406_n 0.00252335f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_439_47#_c_407_n 0.00314884f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_439_47#_c_408_n 2.73397e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_439_47#_c_409_n 0.00157591f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_439_47#_c_410_n 0.00148026f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_439_47#_c_411_n 0.00307484f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_439_47#_c_412_n 0.0591339f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_B_c_575_n 0.0166057f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.345
cc_36 VNB N_B_c_576_n 0.0884473f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_B_c_577_n 0.0122516f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_38 VNB N_B_M1000_g 0.032822f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_B_c_579_n 0.032317f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_B_c_580_n 0.0582273f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_B_M1004_g 0.0223703f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_B_c_582_n 0.00749069f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_B_c_583_n 0.0139121f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_B_c_584_n 0.016494f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_B_c_585_n 0.0104886f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB B 0.00466408f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_555_73#_M1008_g 0.0264657f $X=-0.19 $Y=-0.245 $X2=0.625 $Y2=1.51
cc_48 VNB N_A_555_73#_M1031_g 0.0142722f $X=-0.19 $Y=-0.245 $X2=0.632 $Y2=1.665
cc_49 VNB N_A_555_73#_M1020_g 0.00477426f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_555_73#_c_710_n 0.0291121f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_555_73#_c_711_n 0.00534596f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_A_555_73#_c_712_n 0.00208537f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_555_73#_c_713_n 0.0217963f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_A_555_73#_c_714_n 0.00471236f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_555_73#_c_715_n 0.0373059f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_555_73#_c_716_n 0.00377482f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_555_73#_c_717_n 0.00214925f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_58 VNB N_A_555_73#_c_718_n 0.00269376f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_555_73#_c_719_n 0.00164384f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_555_73#_c_720_n 0.00654172f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_A_555_73#_c_721_n 0.0458556f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VNB N_A_555_73#_c_722_n 0.00409703f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_63 VNB N_A_364_73#_c_959_n 0.0202112f $X=-0.19 $Y=-0.245 $X2=0.625 $Y2=1.51
cc_64 VNB N_A_364_73#_c_960_n 0.0358121f $X=-0.19 $Y=-0.245 $X2=0.632 $Y2=1.51
cc_65 VNB N_A_364_73#_c_961_n 0.00809269f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_66 VNB N_A_364_73#_c_962_n 0.0163806f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_A_364_73#_M1028_g 0.0233088f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_A_364_73#_c_964_n 0.0019663f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_364_73#_c_965_n 0.0146077f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_A_364_73#_c_966_n 0.00250285f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_A_364_73#_c_967_n 0.0104907f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_A_364_73#_c_968_n 0.0115723f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_73 VNB N_A_364_73#_c_969_n 0.00881423f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_74 VNB N_A_364_73#_c_970_n 0.0049567f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_A_364_73#_c_971_n 0.0201566f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_A_364_73#_c_972_n 0.00120757f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_A_364_73#_c_973_n 0.00161117f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_A_364_73#_c_974_n 0.00102098f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_A_364_73#_c_975_n 0.0359038f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_A_364_73#_c_976_n 0.0179748f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_A_364_73#_c_977_n 0.00174443f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_A_364_73#_c_978_n 0.0226464f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_A_364_73#_c_979_n 0.00539282f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_CIN_M1003_g 0.00626498f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=0.655
cc_85 VNB N_CIN_c_1202_n 0.022684f $X=-0.19 $Y=-0.245 $X2=0.505 $Y2=1.675
cc_86 VNB N_CIN_c_1203_n 0.103285f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_CIN_M1023_g 0.0147491f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_CIN_c_1205_n 0.0205785f $X=-0.19 $Y=-0.245 $X2=0.625 $Y2=1.51
cc_89 VNB CIN 0.00309594f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.675
cc_90 VNB N_A_1774_367#_M1017_g 0.037341f $X=-0.19 $Y=-0.245 $X2=0.625 $Y2=1.51
cc_91 VNB N_A_1774_367#_c_1266_n 0.00658655f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VNB N_A_1774_367#_c_1267_n 0.00434256f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_93 VNB N_A_1774_367#_c_1268_n 0.00348854f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_94 VNB N_A_1774_367#_c_1269_n 0.0149982f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_95 VNB N_A_1926_135#_c_1363_n 0.0219979f $X=-0.19 $Y=-0.245 $X2=0.505
+ $Y2=2.465
cc_96 VNB N_A_1926_135#_c_1364_n 0.00347379f $X=-0.19 $Y=-0.245 $X2=0.61
+ $Y2=1.675
cc_97 VNB N_A_1926_135#_c_1365_n 0.00469021f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_98 VNB N_A_1926_135#_c_1366_n 0.0221716f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_99 VNB N_A_1926_135#_c_1367_n 0.00395223f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_100 VNB N_A_1926_135#_c_1368_n 0.00245002f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_101 VNB N_A_1926_135#_c_1369_n 0.0175105f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_102 VNB N_A_1926_135#_c_1370_n 0.00114172f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_103 VNB N_A_1926_135#_c_1371_n 0.00437414f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_104 VNB N_A_1926_135#_c_1372_n 0.0392166f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_105 VNB N_VPWR_c_1460_n 0.521925f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_106 VNB N_A_256_87#_c_1568_n 0.00898735f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_107 VNB N_A_256_87#_c_1569_n 0.0046576f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_108 VNB N_A_256_87#_c_1570_n 0.0147027f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_109 VNB N_A_256_87#_c_1571_n 9.14949e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_110 VNB N_A_256_87#_c_1572_n 0.00218483f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_111 VNB N_A_256_87#_c_1573_n 0.00529985f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_112 VNB N_A_256_87#_c_1574_n 0.00153512f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_113 VNB N_A_1152_389#_c_1651_n 0.00218577f $X=-0.19 $Y=-0.245 $X2=0.635
+ $Y2=1.58
cc_114 VNB N_A_1152_389#_c_1652_n 0.0109166f $X=-0.19 $Y=-0.245 $X2=0.625
+ $Y2=1.51
cc_115 VNB N_A_1152_389#_c_1653_n 0.0027253f $X=-0.19 $Y=-0.245 $X2=0.61
+ $Y2=1.675
cc_116 VNB N_COUT_c_1681_n 0.011422f $X=-0.19 $Y=-0.245 $X2=0.625 $Y2=1.51
cc_117 VNB N_COUT_c_1682_n 0.00321455f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_118 VNB N_A_1500_63#_c_1719_n 0.00268243f $X=-0.19 $Y=-0.245 $X2=0.61
+ $Y2=1.51
cc_119 VNB N_A_1500_63#_c_1720_n 0.00962662f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_120 VNB N_A_1883_395#_c_1752_n 5.85565e-19 $X=-0.19 $Y=-0.245 $X2=0.61
+ $Y2=1.345
cc_121 VNB N_A_1883_395#_c_1753_n 0.00748944f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_122 VNB N_A_1883_395#_c_1754_n 5.50952e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_123 VNB SUM 0.0287167f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_124 VNB N_SUM_c_1802_n 0.038521f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_125 VNB N_VGND_c_1816_n 0.00472864f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.675
cc_126 VNB N_VGND_c_1817_n 0.00801633f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_127 VNB N_VGND_c_1818_n 0.00805673f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_128 VNB N_VGND_c_1819_n 0.0134347f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_129 VNB N_VGND_c_1820_n 0.066854f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_130 VNB N_VGND_c_1821_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_131 VNB N_VGND_c_1822_n 0.0191859f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_132 VNB N_VGND_c_1823_n 0.106499f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_133 VNB N_VGND_c_1824_n 0.070998f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_134 VNB N_VGND_c_1825_n 0.0246757f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_135 VNB N_VGND_c_1826_n 0.664336f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_136 VNB N_VGND_c_1827_n 0.00326991f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_137 VNB N_VGND_c_1828_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_138 VNB N_VGND_c_1829_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_139 VPB N_A_M1012_g 0.0240586f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=2.465
cc_140 VPB N_A_c_250_n 0.00748205f $X=-0.19 $Y=1.655 $X2=0.625 $Y2=1.51
cc_141 VPB N_A_c_251_n 0.00329586f $X=-0.19 $Y=1.655 $X2=0.625 $Y2=1.51
cc_142 VPB N_A_29_47#_M1007_g 0.0255606f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_143 VPB N_A_29_47#_c_285_n 0.00157399f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_144 VPB N_A_29_47#_c_286_n 0.011521f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_145 VPB N_A_29_47#_c_300_n 0.00495495f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_146 VPB N_A_29_47#_c_301_n 0.0367383f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_147 VPB N_A_29_47#_c_290_n 2.09827e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_148 VPB N_A_29_47#_c_303_n 0.0020123f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_149 VPB N_A_29_47#_c_304_n 0.0405163f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_150 VPB N_A_29_47#_c_305_n 0.00129628f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_151 VPB N_A_29_47#_c_306_n 0.00420487f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_152 VPB N_A_29_47#_c_294_n 0.0129964f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_153 VPB N_A_29_47#_c_308_n 0.00509527f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_154 VPB N_A_439_47#_M1021_g 0.0221672f $X=-0.19 $Y=1.655 $X2=0.625 $Y2=1.51
cc_155 VPB N_A_439_47#_M1002_g 0.0242732f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_156 VPB N_A_439_47#_M1019_g 0.028643f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_157 VPB N_A_439_47#_c_402_n 0.00159168f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_158 VPB N_A_439_47#_c_403_n 0.0153189f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_159 VPB N_A_439_47#_c_410_n 0.00205621f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_160 VPB N_A_439_47#_c_419_n 0.00337416f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_161 VPB N_B_M1010_g 0.0239916f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=2.465
cc_162 VPB N_B_c_588_n 0.0850613f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_163 VPB N_B_c_589_n 0.012806f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=1.51
cc_164 VPB N_B_c_590_n 0.0172775f $X=-0.19 $Y=1.655 $X2=0.625 $Y2=1.51
cc_165 VPB N_B_c_591_n 0.029817f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_166 VPB N_B_c_592_n 0.0670172f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_167 VPB N_B_M1013_g 0.0244373f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_168 VPB N_B_c_594_n 0.0255399f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_169 VPB N_B_c_583_n 7.64796e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_170 VPB N_B_c_584_n 0.00665786f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_171 VPB N_B_c_585_n 5.28154e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_172 VPB N_A_555_73#_M1030_g 0.0234321f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_173 VPB N_A_555_73#_M1020_g 0.0302715f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_174 VPB N_A_555_73#_c_711_n 0.00481766f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_175 VPB N_A_555_73#_c_726_n 0.00117385f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_176 VPB N_A_555_73#_c_727_n 0.00654621f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_177 VPB N_A_555_73#_c_728_n 0.00250017f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_178 VPB N_A_555_73#_c_712_n 0.00141099f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_179 VPB N_A_555_73#_c_713_n 0.0172482f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_180 VPB N_A_555_73#_c_731_n 0.00373639f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_181 VPB N_A_555_73#_c_732_n 0.0343975f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_182 VPB N_A_555_73#_c_733_n 0.00342181f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_183 VPB N_A_555_73#_c_734_n 0.0054467f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_184 VPB N_A_555_73#_c_735_n 0.00983119f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_185 VPB N_A_555_73#_c_736_n 0.00436967f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_186 VPB N_A_555_73#_c_716_n 0.0116209f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_187 VPB N_A_555_73#_c_717_n 0.00109931f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_188 VPB N_A_555_73#_c_739_n 0.00244613f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_189 VPB N_A_555_73#_c_722_n 0.00405985f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_190 VPB N_A_555_73#_c_741_n 0.00125213f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_191 VPB N_A_364_73#_c_962_n 0.00207067f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_192 VPB N_A_364_73#_c_981_n 0.0269016f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_193 VPB N_A_364_73#_c_982_n 0.0144397f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_194 VPB N_A_364_73#_c_983_n 0.0201752f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_195 VPB N_A_364_73#_M1024_g 0.0212061f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_196 VPB N_A_364_73#_c_964_n 0.00816794f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_197 VPB N_A_364_73#_c_986_n 0.0110745f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_198 VPB N_A_364_73#_c_967_n 0.0106566f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_199 VPB N_A_364_73#_c_969_n 0.0168232f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_200 VPB N_A_364_73#_c_970_n 0.0035927f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_201 VPB N_A_364_73#_c_971_n 0.0217056f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_202 VPB N_A_364_73#_c_972_n 0.00566058f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_203 VPB N_A_364_73#_c_973_n 0.00192642f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_204 VPB N_A_364_73#_c_974_n 0.00130179f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_205 VPB N_A_364_73#_c_976_n 0.01645f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_206 VPB N_A_364_73#_c_977_n 0.00150793f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_207 VPB N_A_364_73#_c_979_n 0.00488142f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_208 VPB N_CIN_M1003_g 0.0306565f $X=-0.19 $Y=1.655 $X2=0.505 $Y2=0.655
cc_209 VPB N_CIN_M1023_g 0.0281566f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_210 VPB N_A_1774_367#_M1025_g 0.024752f $X=-0.19 $Y=1.655 $X2=0.632 $Y2=1.51
cc_211 VPB N_A_1774_367#_c_1271_n 0.013367f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_212 VPB N_A_1774_367#_c_1272_n 0.00615719f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_213 VPB N_A_1774_367#_c_1273_n 4.78886e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_214 VPB N_A_1774_367#_c_1274_n 0.00340278f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_215 VPB N_A_1774_367#_c_1266_n 0.00552121f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_216 VPB N_A_1774_367#_c_1276_n 0.0218002f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_217 VPB N_A_1774_367#_c_1277_n 0.00563461f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_218 VPB N_A_1774_367#_c_1268_n 0.012028f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_219 VPB N_A_1774_367#_c_1269_n 0.0359174f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_220 VPB N_A_1926_135#_M1018_g 0.0244567f $X=-0.19 $Y=1.655 $X2=0.625 $Y2=1.51
cc_221 VPB N_A_1926_135#_c_1364_n 0.00229576f $X=-0.19 $Y=1.655 $X2=0.61
+ $Y2=1.675
cc_222 VPB N_A_1926_135#_c_1371_n 0.00519569f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_223 VPB N_A_1926_135#_c_1372_n 0.0104902f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_224 VPB N_VPWR_c_1461_n 0.00345454f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=1.675
cc_225 VPB N_VPWR_c_1462_n 0.00477712f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_226 VPB N_VPWR_c_1463_n 0.00472864f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_227 VPB N_VPWR_c_1464_n 0.00240024f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_228 VPB N_VPWR_c_1465_n 0.0995147f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_229 VPB N_VPWR_c_1466_n 0.00510584f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_230 VPB N_VPWR_c_1467_n 0.0736639f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_231 VPB N_VPWR_c_1468_n 0.00324402f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_232 VPB N_VPWR_c_1469_n 0.0163313f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_233 VPB N_VPWR_c_1470_n 0.0716449f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_234 VPB N_VPWR_c_1471_n 0.0159924f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_235 VPB N_VPWR_c_1460_n 0.1187f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_236 VPB N_VPWR_c_1473_n 0.00510842f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_237 VPB N_VPWR_c_1474_n 0.00356964f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_238 VPB N_A_256_87#_c_1575_n 0.00509192f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=1.675
cc_239 VPB N_A_256_87#_c_1576_n 0.0121872f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_240 VPB N_A_256_87#_c_1577_n 2.87297e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_241 VPB N_A_256_87#_c_1569_n 0.00245378f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_242 VPB N_A_1152_389#_c_1652_n 0.00487698f $X=-0.19 $Y=1.655 $X2=0.625
+ $Y2=1.51
cc_243 VPB N_COUT_c_1681_n 0.00581862f $X=-0.19 $Y=1.655 $X2=0.625 $Y2=1.51
cc_244 VPB N_A_1500_63#_c_1721_n 0.00205339f $X=-0.19 $Y=1.655 $X2=0.632
+ $Y2=1.51
cc_245 VPB N_A_1500_63#_c_1720_n 0.00182107f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_246 VPB N_A_1883_395#_c_1753_n 0.0101469f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_247 VPB N_A_1883_395#_c_1756_n 0.0123253f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_248 VPB SUM 0.0553437f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_249 N_A_M1016_g N_A_29_47#_M1005_g 0.0110323f $X=0.505 $Y=0.655 $X2=0 $Y2=0
cc_250 N_A_M1012_g N_A_29_47#_M1007_g 0.00949565f $X=0.505 $Y=2.465 $X2=0 $Y2=0
cc_251 N_A_M1012_g N_A_29_47#_c_285_n 0.00448581f $X=0.505 $Y=2.465 $X2=0 $Y2=0
cc_252 N_A_M1016_g N_A_29_47#_c_287_n 0.0116694f $X=0.505 $Y=0.655 $X2=0 $Y2=0
cc_253 N_A_M1016_g N_A_29_47#_c_288_n 0.0124479f $X=0.505 $Y=0.655 $X2=0 $Y2=0
cc_254 N_A_c_250_n N_A_29_47#_c_288_n 0.00146208f $X=0.625 $Y=1.51 $X2=0 $Y2=0
cc_255 N_A_c_251_n N_A_29_47#_c_288_n 0.0249495f $X=0.625 $Y=1.51 $X2=0 $Y2=0
cc_256 N_A_M1016_g N_A_29_47#_c_316_n 0.00196465f $X=0.505 $Y=0.655 $X2=0 $Y2=0
cc_257 N_A_M1016_g N_A_29_47#_c_289_n 0.00343434f $X=0.505 $Y=0.655 $X2=0 $Y2=0
cc_258 N_A_c_251_n N_A_29_47#_c_289_n 0.00382359f $X=0.625 $Y=1.51 $X2=0 $Y2=0
cc_259 N_A_M1012_g N_A_29_47#_c_290_n 2.57404e-19 $X=0.505 $Y=2.465 $X2=0 $Y2=0
cc_260 N_A_c_250_n N_A_29_47#_c_290_n 9.57737e-19 $X=0.625 $Y=1.51 $X2=0 $Y2=0
cc_261 N_A_c_251_n N_A_29_47#_c_290_n 0.0313487f $X=0.625 $Y=1.51 $X2=0 $Y2=0
cc_262 N_A_M1012_g N_A_29_47#_c_303_n 0.00280383f $X=0.505 $Y=2.465 $X2=0 $Y2=0
cc_263 N_A_M1016_g N_A_29_47#_c_293_n 0.0035087f $X=0.505 $Y=0.655 $X2=0 $Y2=0
cc_264 N_A_M1016_g N_A_29_47#_c_294_n 0.0218245f $X=0.505 $Y=0.655 $X2=0 $Y2=0
cc_265 N_A_c_251_n N_A_29_47#_c_294_n 0.0313839f $X=0.625 $Y=1.51 $X2=0 $Y2=0
cc_266 N_A_M1016_g N_A_29_47#_c_295_n 0.00306263f $X=0.505 $Y=0.655 $X2=0 $Y2=0
cc_267 N_A_c_250_n N_A_29_47#_c_295_n 0.0181301f $X=0.625 $Y=1.51 $X2=0 $Y2=0
cc_268 N_A_c_251_n N_A_29_47#_c_295_n 0.00141225f $X=0.625 $Y=1.51 $X2=0 $Y2=0
cc_269 N_A_M1012_g N_A_29_47#_c_308_n 0.00185402f $X=0.505 $Y=2.465 $X2=0 $Y2=0
cc_270 N_A_M1012_g N_VPWR_c_1461_n 0.018103f $X=0.505 $Y=2.465 $X2=0 $Y2=0
cc_271 N_A_c_250_n N_VPWR_c_1461_n 0.00108746f $X=0.625 $Y=1.51 $X2=0 $Y2=0
cc_272 N_A_c_251_n N_VPWR_c_1461_n 0.0135716f $X=0.625 $Y=1.51 $X2=0 $Y2=0
cc_273 N_A_M1012_g N_VPWR_c_1469_n 0.00486043f $X=0.505 $Y=2.465 $X2=0 $Y2=0
cc_274 N_A_M1012_g N_VPWR_c_1460_n 0.00920706f $X=0.505 $Y=2.465 $X2=0 $Y2=0
cc_275 N_A_M1016_g N_VGND_c_1816_n 0.00659033f $X=0.505 $Y=0.655 $X2=0 $Y2=0
cc_276 N_A_M1016_g N_VGND_c_1822_n 0.00549284f $X=0.505 $Y=0.655 $X2=0 $Y2=0
cc_277 N_A_M1016_g N_VGND_c_1826_n 0.0122601f $X=0.505 $Y=0.655 $X2=0 $Y2=0
cc_278 N_A_29_47#_c_291_n N_A_439_47#_M1026_g 0.0100446f $X=2.32 $Y=0.35 $X2=0
+ $Y2=0
cc_279 N_A_29_47#_c_296_n N_A_439_47#_M1026_g 0.0124007f $X=2.445 $Y=0.35 $X2=0
+ $Y2=0
cc_280 N_A_29_47#_c_304_n N_A_439_47#_M1021_g 0.00982453f $X=3.505 $Y=2.98 $X2=0
+ $Y2=0
cc_281 N_A_29_47#_c_304_n N_A_439_47#_M1002_g 0.00376655f $X=3.505 $Y=2.98 $X2=0
+ $Y2=0
cc_282 N_A_29_47#_c_306_n N_A_439_47#_M1002_g 0.00373758f $X=3.59 $Y=2.53 $X2=0
+ $Y2=0
cc_283 N_A_29_47#_c_296_n N_B_c_575_n 7.36008e-19 $X=2.445 $Y=0.35 $X2=-0.19
+ $Y2=-0.245
cc_284 N_A_29_47#_c_304_n N_B_M1010_g 0.016339f $X=3.505 $Y=2.98 $X2=0 $Y2=0
cc_285 N_A_29_47#_c_304_n N_B_c_588_n 0.0162984f $X=3.505 $Y=2.98 $X2=0 $Y2=0
cc_286 N_A_29_47#_c_306_n N_B_c_590_n 0.00171059f $X=3.59 $Y=2.53 $X2=0 $Y2=0
cc_287 N_A_29_47#_c_304_n N_B_c_594_n 9.68559e-19 $X=3.505 $Y=2.98 $X2=0 $Y2=0
cc_288 N_A_29_47#_c_304_n N_A_555_73#_c_742_n 0.0277254f $X=3.505 $Y=2.98 $X2=0
+ $Y2=0
cc_289 N_A_29_47#_M1002_d N_A_555_73#_c_743_n 0.0155031f $X=3.45 $Y=1.895 $X2=0
+ $Y2=0
cc_290 N_A_29_47#_c_306_n N_A_555_73#_c_743_n 0.0125711f $X=3.59 $Y=2.53 $X2=0
+ $Y2=0
cc_291 N_A_29_47#_M1002_d N_A_555_73#_c_726_n 0.0066111f $X=3.45 $Y=1.895 $X2=0
+ $Y2=0
cc_292 N_A_29_47#_c_306_n N_A_555_73#_c_726_n 0.0410836f $X=3.59 $Y=2.53 $X2=0
+ $Y2=0
cc_293 N_A_29_47#_c_304_n N_A_555_73#_c_728_n 0.0152908f $X=3.505 $Y=2.98 $X2=0
+ $Y2=0
cc_294 N_A_29_47#_c_291_n N_A_364_73#_M1026_s 0.00597963f $X=2.32 $Y=0.35
+ $X2=-0.19 $Y2=-0.245
cc_295 N_A_29_47#_c_286_n N_A_364_73#_c_964_n 0.00492535f $X=1.195 $Y=1.875
+ $X2=0 $Y2=0
cc_296 N_A_29_47#_c_303_n N_A_364_73#_c_964_n 0.00467862f $X=1.15 $Y=2.895 $X2=0
+ $Y2=0
cc_297 N_A_29_47#_c_308_n N_A_364_73#_c_964_n 0.00306968f $X=1.172 $Y=1.875
+ $X2=0 $Y2=0
cc_298 N_A_29_47#_c_285_n N_A_364_73#_c_968_n 0.00672135f $X=1.195 $Y=1.71 $X2=0
+ $Y2=0
cc_299 N_A_29_47#_c_290_n N_A_364_73#_c_968_n 0.00730371f $X=1.172 $Y=1.688
+ $X2=0 $Y2=0
cc_300 N_A_29_47#_c_285_n N_A_364_73#_c_978_n 0.00800017f $X=1.195 $Y=1.71 $X2=0
+ $Y2=0
cc_301 N_A_29_47#_c_289_n N_A_364_73#_c_978_n 0.00763099f $X=1.172 $Y=1.392
+ $X2=0 $Y2=0
cc_302 N_A_29_47#_c_290_n N_A_364_73#_c_978_n 0.0191559f $X=1.172 $Y=1.688 $X2=0
+ $Y2=0
cc_303 N_A_29_47#_c_295_n N_A_364_73#_c_978_n 0.00118432f $X=1.195 $Y=1.37 $X2=0
+ $Y2=0
cc_304 N_A_29_47#_c_303_n N_VPWR_M1012_d 0.00839025f $X=1.15 $Y=2.895 $X2=-0.19
+ $Y2=-0.245
cc_305 N_A_29_47#_c_305_n N_VPWR_M1012_d 0.00140476f $X=1.235 $Y=2.98 $X2=-0.19
+ $Y2=-0.245
cc_306 N_A_29_47#_M1007_g N_VPWR_c_1461_n 0.00480937f $X=1.285 $Y=2.535 $X2=0
+ $Y2=0
cc_307 N_A_29_47#_c_303_n N_VPWR_c_1461_n 0.0614885f $X=1.15 $Y=2.895 $X2=0
+ $Y2=0
cc_308 N_A_29_47#_c_305_n N_VPWR_c_1461_n 0.0139721f $X=1.235 $Y=2.98 $X2=0
+ $Y2=0
cc_309 N_A_29_47#_M1007_g N_VPWR_c_1465_n 0.00321624f $X=1.285 $Y=2.535 $X2=0
+ $Y2=0
cc_310 N_A_29_47#_c_304_n N_VPWR_c_1465_n 0.148244f $X=3.505 $Y=2.98 $X2=0 $Y2=0
cc_311 N_A_29_47#_c_305_n N_VPWR_c_1465_n 0.0113756f $X=1.235 $Y=2.98 $X2=0
+ $Y2=0
cc_312 N_A_29_47#_c_301_n N_VPWR_c_1469_n 0.0173887f $X=0.29 $Y=2.125 $X2=0
+ $Y2=0
cc_313 N_A_29_47#_M1012_s N_VPWR_c_1460_n 0.0042346f $X=0.145 $Y=1.835 $X2=0
+ $Y2=0
cc_314 N_A_29_47#_M1007_g N_VPWR_c_1460_n 0.00596139f $X=1.285 $Y=2.535 $X2=0
+ $Y2=0
cc_315 N_A_29_47#_c_301_n N_VPWR_c_1460_n 0.0101709f $X=0.29 $Y=2.125 $X2=0
+ $Y2=0
cc_316 N_A_29_47#_c_304_n N_VPWR_c_1460_n 0.0865887f $X=3.505 $Y=2.98 $X2=0
+ $Y2=0
cc_317 N_A_29_47#_c_305_n N_VPWR_c_1460_n 0.00646268f $X=1.235 $Y=2.98 $X2=0
+ $Y2=0
cc_318 N_A_29_47#_c_304_n N_A_256_87#_M1007_d 0.00329037f $X=3.505 $Y=2.98 $X2=0
+ $Y2=0
cc_319 N_A_29_47#_c_291_n N_A_256_87#_c_1568_n 0.0217648f $X=2.32 $Y=0.35 $X2=0
+ $Y2=0
cc_320 N_A_29_47#_c_296_n N_A_256_87#_c_1568_n 0.0136706f $X=2.445 $Y=0.35 $X2=0
+ $Y2=0
cc_321 N_A_29_47#_c_304_n N_A_256_87#_c_1576_n 0.0620761f $X=3.505 $Y=2.98 $X2=0
+ $Y2=0
cc_322 N_A_29_47#_c_304_n N_A_256_87#_c_1577_n 0.0180286f $X=3.505 $Y=2.98 $X2=0
+ $Y2=0
cc_323 N_A_29_47#_c_296_n N_A_256_87#_c_1571_n 0.0106464f $X=2.445 $Y=0.35 $X2=0
+ $Y2=0
cc_324 N_A_29_47#_c_289_n N_A_256_87#_c_1573_n 0.00188903f $X=1.172 $Y=1.392
+ $X2=0 $Y2=0
cc_325 N_A_29_47#_c_291_n N_A_256_87#_c_1573_n 0.0176855f $X=2.32 $Y=0.35 $X2=0
+ $Y2=0
cc_326 N_A_29_47#_M1026_d N_A_256_87#_c_1574_n 0.00178407f $X=2.345 $Y=0.365
+ $X2=0 $Y2=0
cc_327 N_A_29_47#_c_288_n N_VGND_M1016_d 0.0092404f $X=0.985 $Y=1.08 $X2=-0.19
+ $Y2=-0.245
cc_328 N_A_29_47#_c_316_n N_VGND_M1016_d 0.0060449f $X=1.07 $Y=0.995 $X2=-0.19
+ $Y2=-0.245
cc_329 N_A_29_47#_M1005_g N_VGND_c_1816_n 0.00140078f $X=1.205 $Y=0.755 $X2=0
+ $Y2=0
cc_330 N_A_29_47#_c_288_n N_VGND_c_1816_n 0.0130182f $X=0.985 $Y=1.08 $X2=0
+ $Y2=0
cc_331 N_A_29_47#_c_316_n N_VGND_c_1816_n 0.0264174f $X=1.07 $Y=0.995 $X2=0
+ $Y2=0
cc_332 N_A_29_47#_c_292_n N_VGND_c_1816_n 0.0135569f $X=1.155 $Y=0.35 $X2=0
+ $Y2=0
cc_333 N_A_29_47#_c_287_n N_VGND_c_1822_n 0.0207694f $X=0.29 $Y=0.43 $X2=0 $Y2=0
cc_334 N_A_29_47#_M1005_g N_VGND_c_1823_n 8.70381e-19 $X=1.205 $Y=0.755 $X2=0
+ $Y2=0
cc_335 N_A_29_47#_c_291_n N_VGND_c_1823_n 0.0702539f $X=2.32 $Y=0.35 $X2=0 $Y2=0
cc_336 N_A_29_47#_c_292_n N_VGND_c_1823_n 0.0114622f $X=1.155 $Y=0.35 $X2=0
+ $Y2=0
cc_337 N_A_29_47#_c_296_n N_VGND_c_1823_n 0.0160274f $X=2.445 $Y=0.35 $X2=0
+ $Y2=0
cc_338 N_A_29_47#_M1016_s N_VGND_c_1826_n 0.0023218f $X=0.145 $Y=0.235 $X2=0
+ $Y2=0
cc_339 N_A_29_47#_c_287_n N_VGND_c_1826_n 0.0130884f $X=0.29 $Y=0.43 $X2=0 $Y2=0
cc_340 N_A_29_47#_c_291_n N_VGND_c_1826_n 0.0429633f $X=2.32 $Y=0.35 $X2=0 $Y2=0
cc_341 N_A_29_47#_c_292_n N_VGND_c_1826_n 0.00657784f $X=1.155 $Y=0.35 $X2=0
+ $Y2=0
cc_342 N_A_29_47#_c_296_n N_VGND_c_1826_n 0.00935889f $X=2.445 $Y=0.35 $X2=0
+ $Y2=0
cc_343 N_A_439_47#_c_397_n N_B_c_575_n 0.00603486f $X=3.4 $Y=1.375 $X2=-0.19
+ $Y2=-0.245
cc_344 N_A_439_47#_c_412_n N_B_c_575_n 0.00873921f $X=3.3 $Y=1.54 $X2=-0.19
+ $Y2=-0.245
cc_345 N_A_439_47#_M1021_g N_B_M1010_g 0.0184304f $X=2.285 $Y=2.455 $X2=0 $Y2=0
cc_346 N_A_439_47#_M1002_g N_B_M1010_g 0.0160947f $X=3.375 $Y=2.315 $X2=0 $Y2=0
cc_347 N_A_439_47#_c_412_n N_B_M1010_g 0.00526391f $X=3.3 $Y=1.54 $X2=0 $Y2=0
cc_348 N_A_439_47#_c_397_n N_B_c_576_n 0.00738071f $X=3.4 $Y=1.375 $X2=0 $Y2=0
cc_349 N_A_439_47#_c_406_n N_B_c_576_n 0.00123167f $X=4.05 $Y=0.35 $X2=0 $Y2=0
cc_350 N_A_439_47#_M1026_g N_B_c_577_n 0.0250317f $X=2.27 $Y=0.685 $X2=0 $Y2=0
cc_351 N_A_439_47#_M1002_g N_B_c_588_n 0.00881852f $X=3.375 $Y=2.315 $X2=0 $Y2=0
cc_352 N_A_439_47#_M1002_g N_B_c_590_n 0.0167083f $X=3.375 $Y=2.315 $X2=0 $Y2=0
cc_353 N_A_439_47#_c_397_n N_B_M1000_g 0.0112356f $X=3.4 $Y=1.375 $X2=0 $Y2=0
cc_354 N_A_439_47#_c_403_n N_B_M1000_g 0.00109491f $X=3.615 $Y=1.54 $X2=0 $Y2=0
cc_355 N_A_439_47#_c_404_n N_B_M1000_g 0.0196054f $X=3.965 $Y=1.2 $X2=0 $Y2=0
cc_356 N_A_439_47#_c_405_n N_B_M1000_g 0.0106246f $X=4.715 $Y=0.35 $X2=0 $Y2=0
cc_357 N_A_439_47#_c_406_n N_B_M1000_g 0.00366581f $X=4.05 $Y=0.35 $X2=0 $Y2=0
cc_358 N_A_439_47#_c_411_n N_B_M1000_g 0.00517851f $X=3.965 $Y=1.285 $X2=0 $Y2=0
cc_359 N_A_439_47#_c_405_n N_B_c_579_n 0.00397031f $X=4.715 $Y=0.35 $X2=0 $Y2=0
cc_360 N_A_439_47#_c_419_n N_B_c_592_n 0.00387526f $X=4.88 $Y=1.935 $X2=0 $Y2=0
cc_361 N_A_439_47#_c_404_n N_B_c_580_n 7.21138e-19 $X=3.965 $Y=1.2 $X2=0 $Y2=0
cc_362 N_A_439_47#_c_405_n N_B_c_580_n 0.0151063f $X=4.715 $Y=0.35 $X2=0 $Y2=0
cc_363 N_A_439_47#_c_407_n N_B_c_580_n 0.00487119f $X=4.88 $Y=0.46 $X2=0 $Y2=0
cc_364 N_A_439_47#_c_409_n N_B_c_580_n 0.00178734f $X=5.045 $Y=0.915 $X2=0 $Y2=0
cc_365 N_A_439_47#_c_398_n N_B_M1004_g 0.0252325f $X=5.685 $Y=1.595 $X2=0 $Y2=0
cc_366 N_A_439_47#_c_400_n N_B_M1004_g 0.0125433f $X=5.805 $Y=1.065 $X2=0 $Y2=0
cc_367 N_A_439_47#_c_405_n N_B_M1004_g 0.00270755f $X=4.715 $Y=0.35 $X2=0 $Y2=0
cc_368 N_A_439_47#_c_407_n N_B_M1004_g 0.00631089f $X=4.88 $Y=0.46 $X2=0 $Y2=0
cc_369 N_A_439_47#_c_408_n N_B_M1004_g 0.00964494f $X=5.38 $Y=0.915 $X2=0 $Y2=0
cc_370 N_A_439_47#_c_409_n N_B_M1004_g 7.4149e-19 $X=5.045 $Y=0.915 $X2=0 $Y2=0
cc_371 N_A_439_47#_c_410_n N_B_M1004_g 0.00605372f $X=5.545 $Y=1.43 $X2=0 $Y2=0
cc_372 N_A_439_47#_c_454_p N_B_M1013_g 0.0101898f $X=5.38 $Y=1.935 $X2=0 $Y2=0
cc_373 N_A_439_47#_c_419_n N_B_M1013_g 0.00660964f $X=4.88 $Y=1.935 $X2=0 $Y2=0
cc_374 N_A_439_47#_c_409_n N_B_c_584_n 9.23198e-19 $X=5.045 $Y=0.915 $X2=0 $Y2=0
cc_375 N_A_439_47#_c_419_n N_B_c_584_n 0.00313846f $X=4.88 $Y=1.935 $X2=0 $Y2=0
cc_376 N_A_439_47#_M1019_g N_B_c_585_n 0.033513f $X=5.685 $Y=2.445 $X2=0 $Y2=0
cc_377 N_A_439_47#_c_410_n N_B_c_585_n 0.00419105f $X=5.545 $Y=1.43 $X2=0 $Y2=0
cc_378 N_A_439_47#_c_398_n B 0.00122947f $X=5.685 $Y=1.595 $X2=0 $Y2=0
cc_379 N_A_439_47#_c_408_n B 0.00750985f $X=5.38 $Y=0.915 $X2=0 $Y2=0
cc_380 N_A_439_47#_c_409_n B 0.0249621f $X=5.045 $Y=0.915 $X2=0 $Y2=0
cc_381 N_A_439_47#_c_454_p B 0.00613307f $X=5.38 $Y=1.935 $X2=0 $Y2=0
cc_382 N_A_439_47#_c_410_n B 0.0293512f $X=5.545 $Y=1.43 $X2=0 $Y2=0
cc_383 N_A_439_47#_c_419_n B 0.0184794f $X=4.88 $Y=1.935 $X2=0 $Y2=0
cc_384 N_A_439_47#_M1019_g N_A_555_73#_M1030_g 0.0259674f $X=5.685 $Y=2.445
+ $X2=0 $Y2=0
cc_385 N_A_439_47#_c_397_n N_A_555_73#_c_711_n 0.00252243f $X=3.4 $Y=1.375 $X2=0
+ $Y2=0
cc_386 N_A_439_47#_c_402_n N_A_555_73#_c_711_n 0.0226269f $X=3.615 $Y=1.54 $X2=0
+ $Y2=0
cc_387 N_A_439_47#_c_403_n N_A_555_73#_c_711_n 0.0110807f $X=3.615 $Y=1.54 $X2=0
+ $Y2=0
cc_388 N_A_439_47#_c_411_n N_A_555_73#_c_711_n 0.010367f $X=3.965 $Y=1.285 $X2=0
+ $Y2=0
cc_389 N_A_439_47#_c_412_n N_A_555_73#_c_711_n 0.013808f $X=3.3 $Y=1.54 $X2=0
+ $Y2=0
cc_390 N_A_439_47#_M1002_g N_A_555_73#_c_743_n 0.0173005f $X=3.375 $Y=2.315
+ $X2=0 $Y2=0
cc_391 N_A_439_47#_c_402_n N_A_555_73#_c_743_n 0.0119497f $X=3.615 $Y=1.54 $X2=0
+ $Y2=0
cc_392 N_A_439_47#_c_403_n N_A_555_73#_c_743_n 0.00197112f $X=3.615 $Y=1.54
+ $X2=0 $Y2=0
cc_393 N_A_439_47#_c_411_n N_A_555_73#_c_743_n 0.00218066f $X=3.965 $Y=1.285
+ $X2=0 $Y2=0
cc_394 N_A_439_47#_M1002_g N_A_555_73#_c_726_n 0.002275f $X=3.375 $Y=2.315 $X2=0
+ $Y2=0
cc_395 N_A_439_47#_M1013_s N_A_555_73#_c_727_n 0.00461378f $X=4.735 $Y=1.835
+ $X2=0 $Y2=0
cc_396 N_A_439_47#_c_419_n N_A_555_73#_c_727_n 0.00232075f $X=4.88 $Y=1.935
+ $X2=0 $Y2=0
cc_397 N_A_439_47#_M1013_s N_A_555_73#_c_761_n 0.00420864f $X=4.735 $Y=1.835
+ $X2=0 $Y2=0
cc_398 N_A_439_47#_M1019_g N_A_555_73#_c_762_n 0.0173467f $X=5.685 $Y=2.445
+ $X2=0 $Y2=0
cc_399 N_A_439_47#_c_454_p N_A_555_73#_c_762_n 0.0180195f $X=5.38 $Y=1.935 $X2=0
+ $Y2=0
cc_400 N_A_439_47#_c_419_n N_A_555_73#_c_762_n 0.00167262f $X=4.88 $Y=1.935
+ $X2=0 $Y2=0
cc_401 N_A_439_47#_M1013_s N_A_555_73#_c_765_n 0.00421212f $X=4.735 $Y=1.835
+ $X2=0 $Y2=0
cc_402 N_A_439_47#_c_419_n N_A_555_73#_c_765_n 0.013891f $X=4.88 $Y=1.935 $X2=0
+ $Y2=0
cc_403 N_A_439_47#_M1019_g N_A_555_73#_c_712_n 0.00122564f $X=5.685 $Y=2.445
+ $X2=0 $Y2=0
cc_404 N_A_439_47#_c_398_n N_A_555_73#_c_713_n 0.0118f $X=5.685 $Y=1.595 $X2=0
+ $Y2=0
cc_405 N_A_439_47#_M1019_g N_A_555_73#_c_731_n 0.0016473f $X=5.685 $Y=2.445
+ $X2=0 $Y2=0
cc_406 N_A_439_47#_M1019_g N_A_555_73#_c_733_n 0.00492071f $X=5.685 $Y=2.445
+ $X2=0 $Y2=0
cc_407 N_A_439_47#_M1002_g N_A_555_73#_c_739_n 0.00146042f $X=3.375 $Y=2.315
+ $X2=0 $Y2=0
cc_408 N_A_439_47#_c_412_n N_A_555_73#_c_739_n 0.00746776f $X=3.3 $Y=1.54 $X2=0
+ $Y2=0
cc_409 N_A_439_47#_c_400_n N_A_364_73#_c_959_n 0.00882135f $X=5.805 $Y=1.065
+ $X2=0 $Y2=0
cc_410 N_A_439_47#_c_398_n N_A_364_73#_c_961_n 0.00882135f $X=5.685 $Y=1.595
+ $X2=0 $Y2=0
cc_411 N_A_439_47#_M1021_g N_A_364_73#_c_964_n 0.005694f $X=2.285 $Y=2.455 $X2=0
+ $Y2=0
cc_412 N_A_439_47#_c_419_n N_A_364_73#_c_986_n 0.0264961f $X=4.88 $Y=1.935 $X2=0
+ $Y2=0
cc_413 N_A_439_47#_c_402_n N_A_364_73#_c_965_n 0.00675009f $X=3.615 $Y=1.54
+ $X2=0 $Y2=0
cc_414 N_A_439_47#_c_403_n N_A_364_73#_c_965_n 0.00333125f $X=3.615 $Y=1.54
+ $X2=0 $Y2=0
cc_415 N_A_439_47#_c_404_n N_A_364_73#_c_965_n 0.040522f $X=3.965 $Y=1.2 $X2=0
+ $Y2=0
cc_416 N_A_439_47#_c_405_n N_A_364_73#_c_965_n 0.0187372f $X=4.715 $Y=0.35 $X2=0
+ $Y2=0
cc_417 N_A_439_47#_c_407_n N_A_364_73#_c_965_n 0.0139332f $X=4.88 $Y=0.46 $X2=0
+ $Y2=0
cc_418 N_A_439_47#_c_409_n N_A_364_73#_c_965_n 0.011731f $X=5.045 $Y=0.915 $X2=0
+ $Y2=0
cc_419 N_A_439_47#_c_411_n N_A_364_73#_c_965_n 0.0130004f $X=3.965 $Y=1.285
+ $X2=0 $Y2=0
cc_420 N_A_439_47#_M1021_g N_A_364_73#_c_967_n 0.00903287f $X=2.285 $Y=2.455
+ $X2=0 $Y2=0
cc_421 N_A_439_47#_M1002_g N_A_364_73#_c_967_n 0.00236133f $X=3.375 $Y=2.315
+ $X2=0 $Y2=0
cc_422 N_A_439_47#_c_401_n N_A_364_73#_c_967_n 4.43336e-19 $X=2.277 $Y=1.45
+ $X2=0 $Y2=0
cc_423 N_A_439_47#_c_402_n N_A_364_73#_c_967_n 0.0116206f $X=3.615 $Y=1.54 $X2=0
+ $Y2=0
cc_424 N_A_439_47#_c_403_n N_A_364_73#_c_967_n 0.0125858f $X=3.615 $Y=1.54 $X2=0
+ $Y2=0
cc_425 N_A_439_47#_c_411_n N_A_364_73#_c_967_n 0.00581316f $X=3.965 $Y=1.285
+ $X2=0 $Y2=0
cc_426 N_A_439_47#_c_412_n N_A_364_73#_c_967_n 0.00879517f $X=3.3 $Y=1.54 $X2=0
+ $Y2=0
cc_427 N_A_439_47#_c_398_n N_A_364_73#_c_969_n 0.00620379f $X=5.685 $Y=1.595
+ $X2=0 $Y2=0
cc_428 N_A_439_47#_M1019_g N_A_364_73#_c_969_n 0.00617891f $X=5.685 $Y=2.445
+ $X2=0 $Y2=0
cc_429 N_A_439_47#_c_408_n N_A_364_73#_c_969_n 0.00707507f $X=5.38 $Y=0.915
+ $X2=0 $Y2=0
cc_430 N_A_439_47#_c_409_n N_A_364_73#_c_969_n 0.0012805f $X=5.045 $Y=0.915
+ $X2=0 $Y2=0
cc_431 N_A_439_47#_c_454_p N_A_364_73#_c_969_n 0.0131719f $X=5.38 $Y=1.935 $X2=0
+ $Y2=0
cc_432 N_A_439_47#_c_410_n N_A_364_73#_c_969_n 0.0338548f $X=5.545 $Y=1.43 $X2=0
+ $Y2=0
cc_433 N_A_439_47#_c_419_n N_A_364_73#_c_969_n 0.00897219f $X=4.88 $Y=1.935
+ $X2=0 $Y2=0
cc_434 N_A_439_47#_M1002_g N_A_364_73#_c_970_n 7.94915e-19 $X=3.375 $Y=2.315
+ $X2=0 $Y2=0
cc_435 N_A_439_47#_c_402_n N_A_364_73#_c_970_n 0.00133525f $X=3.615 $Y=1.54
+ $X2=0 $Y2=0
cc_436 N_A_439_47#_c_403_n N_A_364_73#_c_970_n 0.00129186f $X=3.615 $Y=1.54
+ $X2=0 $Y2=0
cc_437 N_A_439_47#_c_411_n N_A_364_73#_c_970_n 0.00329208f $X=3.965 $Y=1.285
+ $X2=0 $Y2=0
cc_438 N_A_439_47#_M1026_g N_A_364_73#_c_978_n 0.00863186f $X=2.27 $Y=0.685
+ $X2=0 $Y2=0
cc_439 N_A_439_47#_M1021_g N_A_364_73#_c_978_n 0.00533997f $X=2.285 $Y=2.455
+ $X2=0 $Y2=0
cc_440 N_A_439_47#_M1002_g N_A_364_73#_c_979_n 0.00124343f $X=3.375 $Y=2.315
+ $X2=0 $Y2=0
cc_441 N_A_439_47#_c_402_n N_A_364_73#_c_979_n 0.00969407f $X=3.615 $Y=1.54
+ $X2=0 $Y2=0
cc_442 N_A_439_47#_c_403_n N_A_364_73#_c_979_n 0.00293704f $X=3.615 $Y=1.54
+ $X2=0 $Y2=0
cc_443 N_A_439_47#_c_411_n N_A_364_73#_c_979_n 0.00521681f $X=3.965 $Y=1.285
+ $X2=0 $Y2=0
cc_444 N_A_439_47#_c_454_p N_VPWR_M1013_d 0.00804985f $X=5.38 $Y=1.935 $X2=0
+ $Y2=0
cc_445 N_A_439_47#_c_410_n N_VPWR_M1013_d 2.13439e-19 $X=5.545 $Y=1.43 $X2=0
+ $Y2=0
cc_446 N_A_439_47#_M1019_g N_VPWR_c_1462_n 0.00761672f $X=5.685 $Y=2.445 $X2=0
+ $Y2=0
cc_447 N_A_439_47#_M1021_g N_VPWR_c_1465_n 8.06546e-19 $X=2.285 $Y=2.455 $X2=0
+ $Y2=0
cc_448 N_A_439_47#_M1019_g N_VPWR_c_1467_n 0.00443639f $X=5.685 $Y=2.445 $X2=0
+ $Y2=0
cc_449 N_A_439_47#_M1013_s N_VPWR_c_1460_n 0.00259949f $X=4.735 $Y=1.835 $X2=0
+ $Y2=0
cc_450 N_A_439_47#_M1019_g N_VPWR_c_1460_n 0.0054106f $X=5.685 $Y=2.445 $X2=0
+ $Y2=0
cc_451 N_A_439_47#_c_404_n N_A_256_87#_M1009_d 0.00680793f $X=3.965 $Y=1.2 $X2=0
+ $Y2=0
cc_452 N_A_439_47#_c_411_n N_A_256_87#_M1009_d 0.00900512f $X=3.965 $Y=1.285
+ $X2=0 $Y2=0
cc_453 N_A_439_47#_M1021_g N_A_256_87#_c_1575_n 0.00307981f $X=2.285 $Y=2.455
+ $X2=0 $Y2=0
cc_454 N_A_439_47#_M1026_g N_A_256_87#_c_1568_n 0.0123409f $X=2.27 $Y=0.685
+ $X2=0 $Y2=0
cc_455 N_A_439_47#_M1021_g N_A_256_87#_c_1576_n 0.0139394f $X=2.285 $Y=2.455
+ $X2=0 $Y2=0
cc_456 N_A_439_47#_M1026_g N_A_256_87#_c_1569_n 0.0154698f $X=2.27 $Y=0.685
+ $X2=0 $Y2=0
cc_457 N_A_439_47#_M1021_g N_A_256_87#_c_1569_n 0.0218068f $X=2.285 $Y=2.455
+ $X2=0 $Y2=0
cc_458 N_A_439_47#_M1002_g N_A_256_87#_c_1569_n 2.09225e-19 $X=3.375 $Y=2.315
+ $X2=0 $Y2=0
cc_459 N_A_439_47#_c_401_n N_A_256_87#_c_1569_n 0.00170337f $X=2.277 $Y=1.45
+ $X2=0 $Y2=0
cc_460 N_A_439_47#_c_412_n N_A_256_87#_c_1569_n 0.0171161f $X=3.3 $Y=1.54 $X2=0
+ $Y2=0
cc_461 N_A_439_47#_M1026_g N_A_256_87#_c_1598_n 8.21167e-19 $X=2.27 $Y=0.685
+ $X2=0 $Y2=0
cc_462 N_A_439_47#_c_397_n N_A_256_87#_c_1598_n 0.00129355f $X=3.4 $Y=1.375
+ $X2=0 $Y2=0
cc_463 N_A_439_47#_c_397_n N_A_256_87#_c_1570_n 0.00307326f $X=3.4 $Y=1.375
+ $X2=0 $Y2=0
cc_464 N_A_439_47#_c_406_n N_A_256_87#_c_1570_n 0.0152909f $X=4.05 $Y=0.35 $X2=0
+ $Y2=0
cc_465 N_A_439_47#_c_397_n N_A_256_87#_c_1572_n 0.00910135f $X=3.4 $Y=1.375
+ $X2=0 $Y2=0
cc_466 N_A_439_47#_c_404_n N_A_256_87#_c_1572_n 0.0423947f $X=3.965 $Y=1.2 $X2=0
+ $Y2=0
cc_467 N_A_439_47#_c_411_n N_A_256_87#_c_1572_n 0.0142567f $X=3.965 $Y=1.285
+ $X2=0 $Y2=0
cc_468 N_A_439_47#_M1026_g N_A_256_87#_c_1573_n 0.00580048f $X=2.27 $Y=0.685
+ $X2=0 $Y2=0
cc_469 N_A_439_47#_M1026_g N_A_256_87#_c_1574_n 0.00228676f $X=2.27 $Y=0.685
+ $X2=0 $Y2=0
cc_470 N_A_439_47#_c_412_n N_A_256_87#_c_1574_n 0.0052783f $X=3.3 $Y=1.54 $X2=0
+ $Y2=0
cc_471 N_A_439_47#_c_400_n N_A_1152_389#_c_1651_n 0.00977465f $X=5.805 $Y=1.065
+ $X2=0 $Y2=0
cc_472 N_A_439_47#_c_398_n N_A_1152_389#_c_1652_n 0.015597f $X=5.685 $Y=1.595
+ $X2=0 $Y2=0
cc_473 N_A_439_47#_c_400_n N_A_1152_389#_c_1652_n 0.00172526f $X=5.805 $Y=1.065
+ $X2=0 $Y2=0
cc_474 N_A_439_47#_c_454_p N_A_1152_389#_c_1652_n 0.010104f $X=5.38 $Y=1.935
+ $X2=0 $Y2=0
cc_475 N_A_439_47#_c_410_n N_A_1152_389#_c_1652_n 0.0584065f $X=5.545 $Y=1.43
+ $X2=0 $Y2=0
cc_476 N_A_439_47#_c_400_n N_A_1152_389#_c_1653_n 0.00317954f $X=5.805 $Y=1.065
+ $X2=0 $Y2=0
cc_477 N_A_439_47#_c_408_n N_A_1152_389#_c_1653_n 0.0134824f $X=5.38 $Y=0.915
+ $X2=0 $Y2=0
cc_478 N_A_439_47#_c_408_n N_VGND_M1004_d 0.0109911f $X=5.38 $Y=0.915 $X2=0
+ $Y2=0
cc_479 N_A_439_47#_c_410_n N_VGND_M1004_d 0.00215798f $X=5.545 $Y=1.43 $X2=0
+ $Y2=0
cc_480 N_A_439_47#_c_398_n N_VGND_c_1817_n 5.74223e-19 $X=5.685 $Y=1.595 $X2=0
+ $Y2=0
cc_481 N_A_439_47#_c_400_n N_VGND_c_1817_n 0.0059071f $X=5.805 $Y=1.065 $X2=0
+ $Y2=0
cc_482 N_A_439_47#_c_405_n N_VGND_c_1817_n 0.00880411f $X=4.715 $Y=0.35 $X2=0
+ $Y2=0
cc_483 N_A_439_47#_c_408_n N_VGND_c_1817_n 0.0261572f $X=5.38 $Y=0.915 $X2=0
+ $Y2=0
cc_484 N_A_439_47#_M1026_g N_VGND_c_1823_n 0.00283533f $X=2.27 $Y=0.685 $X2=0
+ $Y2=0
cc_485 N_A_439_47#_c_405_n N_VGND_c_1823_n 0.0616564f $X=4.715 $Y=0.35 $X2=0
+ $Y2=0
cc_486 N_A_439_47#_c_406_n N_VGND_c_1823_n 0.0113569f $X=4.05 $Y=0.35 $X2=0
+ $Y2=0
cc_487 N_A_439_47#_c_400_n N_VGND_c_1824_n 0.00425753f $X=5.805 $Y=1.065 $X2=0
+ $Y2=0
cc_488 N_A_439_47#_M1026_g N_VGND_c_1826_n 0.0037193f $X=2.27 $Y=0.685 $X2=0
+ $Y2=0
cc_489 N_A_439_47#_c_400_n N_VGND_c_1826_n 0.00798825f $X=5.805 $Y=1.065 $X2=0
+ $Y2=0
cc_490 N_A_439_47#_c_405_n N_VGND_c_1826_n 0.0348083f $X=4.715 $Y=0.35 $X2=0
+ $Y2=0
cc_491 N_A_439_47#_c_406_n N_VGND_c_1826_n 0.005852f $X=4.05 $Y=0.35 $X2=0 $Y2=0
cc_492 N_A_439_47#_c_408_n N_VGND_c_1826_n 0.00979413f $X=5.38 $Y=0.915 $X2=0
+ $Y2=0
cc_493 N_B_M1010_g N_A_555_73#_c_742_n 0.00606163f $X=2.715 $Y=2.455 $X2=0 $Y2=0
cc_494 N_B_c_575_n N_A_555_73#_c_711_n 0.00204713f $X=2.7 $Y=0.255 $X2=0 $Y2=0
cc_495 N_B_c_590_n N_A_555_73#_c_743_n 0.00553632f $X=4.065 $Y=2.845 $X2=0 $Y2=0
cc_496 N_B_c_590_n N_A_555_73#_c_726_n 0.0174127f $X=4.065 $Y=2.845 $X2=0 $Y2=0
cc_497 N_B_c_592_n N_A_555_73#_c_726_n 7.63452e-19 $X=4.585 $Y=2.845 $X2=0 $Y2=0
cc_498 N_B_c_594_n N_A_555_73#_c_726_n 0.00297649f $X=4.065 $Y=2.92 $X2=0 $Y2=0
cc_499 N_B_c_591_n N_A_555_73#_c_727_n 0.0273287f $X=4.51 $Y=2.92 $X2=0 $Y2=0
cc_500 N_B_c_594_n N_A_555_73#_c_727_n 0.00954135f $X=4.065 $Y=2.92 $X2=0 $Y2=0
cc_501 N_B_c_588_n N_A_555_73#_c_728_n 0.0011085f $X=3.99 $Y=3.15 $X2=0 $Y2=0
cc_502 N_B_c_594_n N_A_555_73#_c_728_n 0.00376332f $X=4.065 $Y=2.92 $X2=0 $Y2=0
cc_503 N_B_c_592_n N_A_555_73#_c_761_n 0.00504992f $X=4.585 $Y=2.845 $X2=0 $Y2=0
cc_504 N_B_M1013_g N_A_555_73#_c_762_n 0.0135537f $X=5.095 $Y=2.465 $X2=0 $Y2=0
cc_505 N_B_c_592_n N_A_555_73#_c_765_n 0.00172966f $X=4.585 $Y=2.845 $X2=0 $Y2=0
cc_506 N_B_M1010_g N_A_555_73#_c_739_n 0.0024346f $X=2.715 $Y=2.455 $X2=0 $Y2=0
cc_507 N_B_c_590_n N_A_364_73#_c_986_n 0.00755721f $X=4.065 $Y=2.845 $X2=0 $Y2=0
cc_508 N_B_c_591_n N_A_364_73#_c_986_n 0.00401797f $X=4.51 $Y=2.92 $X2=0 $Y2=0
cc_509 N_B_c_592_n N_A_364_73#_c_986_n 0.0142702f $X=4.585 $Y=2.845 $X2=0 $Y2=0
cc_510 N_B_M1000_g N_A_364_73#_c_965_n 0.00330041f $X=4.095 $Y=0.945 $X2=0 $Y2=0
cc_511 N_B_c_580_n N_A_364_73#_c_965_n 0.00990292f $X=4.595 $Y=1.34 $X2=0 $Y2=0
cc_512 N_B_c_583_n N_A_364_73#_c_965_n 0.00538885f $X=4.59 $Y=1.505 $X2=0 $Y2=0
cc_513 B N_A_364_73#_c_965_n 0.0282981f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_514 N_B_M1010_g N_A_364_73#_c_967_n 0.00188655f $X=2.715 $Y=2.455 $X2=0 $Y2=0
cc_515 N_B_c_592_n N_A_364_73#_c_969_n 0.00768171f $X=4.585 $Y=2.845 $X2=0 $Y2=0
cc_516 N_B_M1013_g N_A_364_73#_c_969_n 0.00232294f $X=5.095 $Y=2.465 $X2=0 $Y2=0
cc_517 N_B_c_583_n N_A_364_73#_c_969_n 0.00736514f $X=4.59 $Y=1.505 $X2=0 $Y2=0
cc_518 N_B_c_584_n N_A_364_73#_c_969_n 0.00163641f $X=5.02 $Y=1.505 $X2=0 $Y2=0
cc_519 N_B_c_585_n N_A_364_73#_c_969_n 9.00145e-19 $X=5.095 $Y=1.505 $X2=0 $Y2=0
cc_520 B N_A_364_73#_c_969_n 0.0195401f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_521 N_B_c_590_n N_A_364_73#_c_970_n 0.00527853f $X=4.065 $Y=2.845 $X2=0 $Y2=0
cc_522 N_B_M1000_g N_A_364_73#_c_970_n 0.0029131f $X=4.095 $Y=0.945 $X2=0 $Y2=0
cc_523 N_B_c_590_n N_A_364_73#_c_979_n 0.00537865f $X=4.065 $Y=2.845 $X2=0 $Y2=0
cc_524 N_B_M1000_g N_A_364_73#_c_979_n 0.00329507f $X=4.095 $Y=0.945 $X2=0 $Y2=0
cc_525 N_B_c_583_n N_A_364_73#_c_979_n 0.00741589f $X=4.59 $Y=1.505 $X2=0 $Y2=0
cc_526 B N_A_364_73#_c_979_n 0.00830519f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_527 N_B_M1013_g N_VPWR_c_1462_n 0.0102151f $X=5.095 $Y=2.465 $X2=0 $Y2=0
cc_528 N_B_c_589_n N_VPWR_c_1465_n 0.0348528f $X=2.79 $Y=3.15 $X2=0 $Y2=0
cc_529 N_B_c_591_n N_VPWR_c_1465_n 0.00274426f $X=4.51 $Y=2.92 $X2=0 $Y2=0
cc_530 N_B_M1013_g N_VPWR_c_1465_n 0.00364083f $X=5.095 $Y=2.465 $X2=0 $Y2=0
cc_531 N_B_c_588_n N_VPWR_c_1460_n 0.0337988f $X=3.99 $Y=3.15 $X2=0 $Y2=0
cc_532 N_B_c_589_n N_VPWR_c_1460_n 0.00604685f $X=2.79 $Y=3.15 $X2=0 $Y2=0
cc_533 N_B_M1013_g N_VPWR_c_1460_n 0.00577754f $X=5.095 $Y=2.465 $X2=0 $Y2=0
cc_534 N_B_c_594_n N_VPWR_c_1460_n 0.0060468f $X=4.065 $Y=2.92 $X2=0 $Y2=0
cc_535 N_B_M1010_g N_A_256_87#_c_1576_n 0.00230329f $X=2.715 $Y=2.455 $X2=0
+ $Y2=0
cc_536 N_B_c_575_n N_A_256_87#_c_1569_n 0.0037661f $X=2.7 $Y=0.255 $X2=0 $Y2=0
cc_537 N_B_M1010_g N_A_256_87#_c_1569_n 0.00922294f $X=2.715 $Y=2.455 $X2=0
+ $Y2=0
cc_538 N_B_c_575_n N_A_256_87#_c_1598_n 0.0111059f $X=2.7 $Y=0.255 $X2=0 $Y2=0
cc_539 N_B_c_576_n N_A_256_87#_c_1570_n 0.0161153f $X=4.02 $Y=0.18 $X2=0 $Y2=0
cc_540 N_B_M1000_g N_A_256_87#_c_1570_n 9.70705e-19 $X=4.095 $Y=0.945 $X2=0
+ $Y2=0
cc_541 N_B_c_575_n N_A_256_87#_c_1571_n 0.00607618f $X=2.7 $Y=0.255 $X2=0 $Y2=0
cc_542 N_B_c_576_n N_A_256_87#_c_1571_n 0.00134409f $X=4.02 $Y=0.18 $X2=0 $Y2=0
cc_543 N_B_c_575_n N_A_256_87#_c_1572_n 4.16909e-19 $X=2.7 $Y=0.255 $X2=0 $Y2=0
cc_544 N_B_M1000_g N_A_256_87#_c_1572_n 0.0018577f $X=4.095 $Y=0.945 $X2=0 $Y2=0
cc_545 N_B_c_575_n N_A_256_87#_c_1574_n 0.0104208f $X=2.7 $Y=0.255 $X2=0 $Y2=0
cc_546 N_B_M1004_g N_A_1152_389#_c_1651_n 8.90528e-19 $X=5.095 $Y=0.735 $X2=0
+ $Y2=0
cc_547 N_B_c_579_n N_VGND_c_1817_n 0.0014037f $X=4.52 $Y=0.18 $X2=0 $Y2=0
cc_548 N_B_M1004_g N_VGND_c_1817_n 0.00513393f $X=5.095 $Y=0.735 $X2=0 $Y2=0
cc_549 N_B_c_577_n N_VGND_c_1823_n 0.0489628f $X=2.775 $Y=0.18 $X2=0 $Y2=0
cc_550 N_B_M1004_g N_VGND_c_1823_n 0.00475301f $X=5.095 $Y=0.735 $X2=0 $Y2=0
cc_551 N_B_c_576_n N_VGND_c_1826_n 0.0348552f $X=4.02 $Y=0.18 $X2=0 $Y2=0
cc_552 N_B_c_577_n N_VGND_c_1826_n 0.00690017f $X=2.775 $Y=0.18 $X2=0 $Y2=0
cc_553 N_B_c_579_n N_VGND_c_1826_n 0.0138572f $X=4.52 $Y=0.18 $X2=0 $Y2=0
cc_554 N_B_M1004_g N_VGND_c_1826_n 0.00565064f $X=5.095 $Y=0.735 $X2=0 $Y2=0
cc_555 N_B_c_582_n N_VGND_c_1826_n 0.0037101f $X=4.095 $Y=0.18 $X2=0 $Y2=0
cc_556 N_A_555_73#_c_712_n N_A_364_73#_c_961_n 0.00124844f $X=6.255 $Y=1.62
+ $X2=0 $Y2=0
cc_557 N_A_555_73#_c_713_n N_A_364_73#_c_961_n 0.014694f $X=6.255 $Y=1.62 $X2=0
+ $Y2=0
cc_558 N_A_555_73#_c_713_n N_A_364_73#_c_962_n 0.00523248f $X=6.255 $Y=1.62
+ $X2=0 $Y2=0
cc_559 N_A_555_73#_c_714_n N_A_364_73#_c_962_n 0.00255287f $X=7.515 $Y=1.28
+ $X2=0 $Y2=0
cc_560 N_A_555_73#_c_715_n N_A_364_73#_c_962_n 0.0118097f $X=7.515 $Y=1.28 $X2=0
+ $Y2=0
cc_561 N_A_555_73#_c_722_n N_A_364_73#_c_962_n 0.00192647f $X=7.44 $Y=1.745
+ $X2=0 $Y2=0
cc_562 N_A_555_73#_c_734_n N_A_364_73#_c_981_n 0.00666662f $X=7.35 $Y=2.895
+ $X2=0 $Y2=0
cc_563 N_A_555_73#_c_715_n N_A_364_73#_c_981_n 0.00966628f $X=7.515 $Y=1.28
+ $X2=0 $Y2=0
cc_564 N_A_555_73#_c_722_n N_A_364_73#_c_981_n 0.0103386f $X=7.44 $Y=1.745 $X2=0
+ $Y2=0
cc_565 N_A_555_73#_M1030_g N_A_364_73#_c_982_n 5.41349e-19 $X=6.23 $Y=2.365
+ $X2=0 $Y2=0
cc_566 N_A_555_73#_c_734_n N_A_364_73#_c_983_n 0.0330011f $X=7.35 $Y=2.895 $X2=0
+ $Y2=0
cc_567 N_A_555_73#_c_735_n N_A_364_73#_c_983_n 0.00592729f $X=8.145 $Y=2.98
+ $X2=0 $Y2=0
cc_568 N_A_555_73#_c_741_n N_A_364_73#_c_983_n 0.00163657f $X=7.35 $Y=2.98 $X2=0
+ $Y2=0
cc_569 N_A_555_73#_M1020_g N_A_364_73#_M1024_g 0.0357608f $X=9.77 $Y=2.395 $X2=0
+ $Y2=0
cc_570 N_A_555_73#_M1031_g N_A_364_73#_M1028_g 0.00953054f $X=9.555 $Y=0.995
+ $X2=0 $Y2=0
cc_571 N_A_555_73#_c_710_n N_A_364_73#_M1028_g 0.00193838f $X=9.77 $Y=1.5 $X2=0
+ $Y2=0
cc_572 N_A_555_73#_c_721_n N_A_364_73#_M1028_g 5.51888e-19 $X=9.61 $Y=0.4 $X2=0
+ $Y2=0
cc_573 N_A_555_73#_c_743_n N_A_364_73#_c_986_n 0.0132229f $X=3.855 $Y=2.045
+ $X2=0 $Y2=0
cc_574 N_A_555_73#_c_726_n N_A_364_73#_c_986_n 0.0407847f $X=3.94 $Y=2.895 $X2=0
+ $Y2=0
cc_575 N_A_555_73#_c_727_n N_A_364_73#_c_986_n 0.0192314f $X=4.795 $Y=2.98 $X2=0
+ $Y2=0
cc_576 N_A_555_73#_c_761_n N_A_364_73#_c_986_n 0.00541095f $X=4.88 $Y=2.895
+ $X2=0 $Y2=0
cc_577 N_A_555_73#_c_765_n N_A_364_73#_c_986_n 0.00932269f $X=4.965 $Y=2.52
+ $X2=0 $Y2=0
cc_578 N_A_555_73#_M1008_g N_A_364_73#_c_966_n 0.00117722f $X=7.425 $Y=0.635
+ $X2=0 $Y2=0
cc_579 N_A_555_73#_c_714_n N_A_364_73#_c_966_n 0.0171581f $X=7.515 $Y=1.28 $X2=0
+ $Y2=0
cc_580 N_A_555_73#_c_711_n N_A_364_73#_c_967_n 0.0226056f $X=3.185 $Y=0.78 $X2=0
+ $Y2=0
cc_581 N_A_555_73#_c_743_n N_A_364_73#_c_967_n 0.019495f $X=3.855 $Y=2.045 $X2=0
+ $Y2=0
cc_582 N_A_555_73#_c_739_n N_A_364_73#_c_967_n 0.0119485f $X=3.045 $Y=2.04 $X2=0
+ $Y2=0
cc_583 N_A_555_73#_c_712_n N_A_364_73#_c_969_n 0.0190027f $X=6.255 $Y=1.62 $X2=0
+ $Y2=0
cc_584 N_A_555_73#_c_713_n N_A_364_73#_c_969_n 0.0102068f $X=6.255 $Y=1.62 $X2=0
+ $Y2=0
cc_585 N_A_555_73#_c_743_n N_A_364_73#_c_970_n 0.00260866f $X=3.855 $Y=2.045
+ $X2=0 $Y2=0
cc_586 N_A_555_73#_M1020_g N_A_364_73#_c_971_n 0.00695833f $X=9.77 $Y=2.395
+ $X2=0 $Y2=0
cc_587 N_A_555_73#_c_710_n N_A_364_73#_c_971_n 0.00607197f $X=9.77 $Y=1.5 $X2=0
+ $Y2=0
cc_588 N_A_555_73#_c_715_n N_A_364_73#_c_971_n 0.00161502f $X=7.515 $Y=1.28
+ $X2=0 $Y2=0
cc_589 N_A_555_73#_c_716_n N_A_364_73#_c_971_n 0.0439705f $X=8.755 $Y=1.675
+ $X2=0 $Y2=0
cc_590 N_A_555_73#_c_717_n N_A_364_73#_c_971_n 0.0160454f $X=8.315 $Y=1.675
+ $X2=0 $Y2=0
cc_591 N_A_555_73#_c_722_n N_A_364_73#_c_971_n 0.0348702f $X=7.44 $Y=1.745 $X2=0
+ $Y2=0
cc_592 N_A_555_73#_c_714_n N_A_364_73#_c_972_n 6.03099e-19 $X=7.515 $Y=1.28
+ $X2=0 $Y2=0
cc_593 N_A_555_73#_c_722_n N_A_364_73#_c_972_n 0.00163729f $X=7.44 $Y=1.745
+ $X2=0 $Y2=0
cc_594 N_A_555_73#_c_714_n N_A_364_73#_c_973_n 0.00884353f $X=7.515 $Y=1.28
+ $X2=0 $Y2=0
cc_595 N_A_555_73#_c_722_n N_A_364_73#_c_973_n 0.0119189f $X=7.44 $Y=1.745 $X2=0
+ $Y2=0
cc_596 N_A_555_73#_M1008_g N_A_364_73#_c_975_n 0.0118097f $X=7.425 $Y=0.635
+ $X2=0 $Y2=0
cc_597 N_A_555_73#_c_714_n N_A_364_73#_c_975_n 0.00118899f $X=7.515 $Y=1.28
+ $X2=0 $Y2=0
cc_598 N_A_555_73#_c_710_n N_A_364_73#_c_976_n 0.0163774f $X=9.77 $Y=1.5 $X2=0
+ $Y2=0
cc_599 N_A_555_73#_c_710_n N_A_364_73#_c_977_n 4.40797e-19 $X=9.77 $Y=1.5 $X2=0
+ $Y2=0
cc_600 N_A_555_73#_c_743_n N_A_364_73#_c_979_n 0.0030439f $X=3.855 $Y=2.045
+ $X2=0 $Y2=0
cc_601 N_A_555_73#_c_734_n N_CIN_M1003_g 0.00122704f $X=7.35 $Y=2.895 $X2=0
+ $Y2=0
cc_602 N_A_555_73#_c_735_n N_CIN_M1003_g 0.0149171f $X=8.145 $Y=2.98 $X2=0 $Y2=0
cc_603 N_A_555_73#_c_736_n N_CIN_M1003_g 0.0152823f $X=8.23 $Y=2.895 $X2=0 $Y2=0
cc_604 N_A_555_73#_c_717_n N_CIN_M1003_g 0.00171484f $X=8.315 $Y=1.675 $X2=0
+ $Y2=0
cc_605 N_A_555_73#_c_722_n N_CIN_M1003_g 6.84362e-19 $X=7.44 $Y=1.745 $X2=0
+ $Y2=0
cc_606 N_A_555_73#_M1008_g N_CIN_c_1202_n 0.012361f $X=7.425 $Y=0.635 $X2=0
+ $Y2=0
cc_607 N_A_555_73#_c_718_n N_CIN_c_1202_n 0.00444907f $X=8.84 $Y=1.59 $X2=0
+ $Y2=0
cc_608 N_A_555_73#_c_714_n N_CIN_c_1203_n 7.11696e-19 $X=7.515 $Y=1.28 $X2=0
+ $Y2=0
cc_609 N_A_555_73#_c_715_n N_CIN_c_1203_n 0.0102179f $X=7.515 $Y=1.28 $X2=0
+ $Y2=0
cc_610 N_A_555_73#_c_716_n N_CIN_c_1203_n 0.0119624f $X=8.755 $Y=1.675 $X2=0
+ $Y2=0
cc_611 N_A_555_73#_c_717_n N_CIN_c_1203_n 0.00767492f $X=8.315 $Y=1.675 $X2=0
+ $Y2=0
cc_612 N_A_555_73#_c_718_n N_CIN_c_1203_n 0.0118384f $X=8.84 $Y=1.59 $X2=0 $Y2=0
cc_613 N_A_555_73#_M1031_g N_CIN_M1023_g 0.0020273f $X=9.555 $Y=0.995 $X2=0
+ $Y2=0
cc_614 N_A_555_73#_c_736_n N_CIN_M1023_g 0.00451029f $X=8.23 $Y=2.895 $X2=0
+ $Y2=0
cc_615 N_A_555_73#_c_716_n N_CIN_M1023_g 0.0161188f $X=8.755 $Y=1.675 $X2=0
+ $Y2=0
cc_616 N_A_555_73#_c_718_n N_CIN_M1023_g 0.00622329f $X=8.84 $Y=1.59 $X2=0 $Y2=0
cc_617 N_A_555_73#_M1031_g N_CIN_c_1205_n 0.0168951f $X=9.555 $Y=0.995 $X2=0
+ $Y2=0
cc_618 N_A_555_73#_c_718_n N_CIN_c_1205_n 0.0118012f $X=8.84 $Y=1.59 $X2=0 $Y2=0
cc_619 N_A_555_73#_c_720_n N_CIN_c_1205_n 0.0219563f $X=9.61 $Y=0.4 $X2=0 $Y2=0
cc_620 N_A_555_73#_c_721_n N_CIN_c_1205_n 0.0109782f $X=9.61 $Y=0.4 $X2=0 $Y2=0
cc_621 N_A_555_73#_c_716_n CIN 0.0168267f $X=8.755 $Y=1.675 $X2=0 $Y2=0
cc_622 N_A_555_73#_c_717_n CIN 0.00510303f $X=8.315 $Y=1.675 $X2=0 $Y2=0
cc_623 N_A_555_73#_c_718_n CIN 0.023108f $X=8.84 $Y=1.59 $X2=0 $Y2=0
cc_624 N_A_555_73#_c_720_n N_A_1774_367#_M1022_d 0.00213864f $X=9.61 $Y=0.4
+ $X2=-0.19 $Y2=-0.245
cc_625 N_A_555_73#_M1020_g N_A_1774_367#_c_1271_n 0.00499618f $X=9.77 $Y=2.395
+ $X2=0 $Y2=0
cc_626 N_A_555_73#_M1031_g N_A_1774_367#_c_1282_n 0.00841983f $X=9.555 $Y=0.995
+ $X2=0 $Y2=0
cc_627 N_A_555_73#_c_720_n N_A_1774_367#_c_1282_n 0.0256538f $X=9.61 $Y=0.4
+ $X2=0 $Y2=0
cc_628 N_A_555_73#_c_716_n N_A_1774_367#_c_1274_n 0.00419599f $X=8.755 $Y=1.675
+ $X2=0 $Y2=0
cc_629 N_A_555_73#_M1031_g N_A_1774_367#_c_1266_n 0.00277058f $X=9.555 $Y=0.995
+ $X2=0 $Y2=0
cc_630 N_A_555_73#_M1020_g N_A_1774_367#_c_1266_n 0.0149835f $X=9.77 $Y=2.395
+ $X2=0 $Y2=0
cc_631 N_A_555_73#_c_716_n N_A_1774_367#_c_1266_n 0.011158f $X=8.755 $Y=1.675
+ $X2=0 $Y2=0
cc_632 N_A_555_73#_M1031_g N_A_1774_367#_c_1267_n 0.0041705f $X=9.555 $Y=0.995
+ $X2=0 $Y2=0
cc_633 N_A_555_73#_c_718_n N_A_1774_367#_c_1267_n 0.0298268f $X=8.84 $Y=1.59
+ $X2=0 $Y2=0
cc_634 N_A_555_73#_M1020_g N_A_1774_367#_c_1276_n 0.00778052f $X=9.77 $Y=2.395
+ $X2=0 $Y2=0
cc_635 N_A_555_73#_M1031_g N_A_1926_135#_c_1364_n 0.00139336f $X=9.555 $Y=0.995
+ $X2=0 $Y2=0
cc_636 N_A_555_73#_M1020_g N_A_1926_135#_c_1364_n 0.0118197f $X=9.77 $Y=2.395
+ $X2=0 $Y2=0
cc_637 N_A_555_73#_c_710_n N_A_1926_135#_c_1364_n 0.00643673f $X=9.77 $Y=1.5
+ $X2=0 $Y2=0
cc_638 N_A_555_73#_M1031_g N_A_1926_135#_c_1380_n 0.00180275f $X=9.555 $Y=0.995
+ $X2=0 $Y2=0
cc_639 N_A_555_73#_c_710_n N_A_1926_135#_c_1380_n 5.17548e-19 $X=9.77 $Y=1.5
+ $X2=0 $Y2=0
cc_640 N_A_555_73#_c_720_n N_A_1926_135#_c_1380_n 5.67848e-19 $X=9.61 $Y=0.4
+ $X2=0 $Y2=0
cc_641 N_A_555_73#_c_721_n N_A_1926_135#_c_1380_n 3.2992e-19 $X=9.61 $Y=0.4
+ $X2=0 $Y2=0
cc_642 N_A_555_73#_M1031_g N_A_1926_135#_c_1365_n 0.00710803f $X=9.555 $Y=0.995
+ $X2=0 $Y2=0
cc_643 N_A_555_73#_c_720_n N_A_1926_135#_c_1365_n 0.0101143f $X=9.61 $Y=0.4
+ $X2=0 $Y2=0
cc_644 N_A_555_73#_c_721_n N_A_1926_135#_c_1365_n 8.57466e-19 $X=9.61 $Y=0.4
+ $X2=0 $Y2=0
cc_645 N_A_555_73#_c_720_n N_A_1926_135#_c_1367_n 0.0144263f $X=9.61 $Y=0.4
+ $X2=0 $Y2=0
cc_646 N_A_555_73#_c_721_n N_A_1926_135#_c_1367_n 0.00132764f $X=9.61 $Y=0.4
+ $X2=0 $Y2=0
cc_647 N_A_555_73#_M1020_g N_A_1926_135#_c_1389_n 0.00529063f $X=9.77 $Y=2.395
+ $X2=0 $Y2=0
cc_648 N_A_555_73#_c_762_n N_VPWR_M1013_d 0.0101725f $X=6.165 $Y=2.52 $X2=0
+ $Y2=0
cc_649 N_A_555_73#_c_735_n N_VPWR_M1003_d 0.0013163f $X=8.145 $Y=2.98 $X2=0
+ $Y2=0
cc_650 N_A_555_73#_c_736_n N_VPWR_M1003_d 0.0250912f $X=8.23 $Y=2.895 $X2=0
+ $Y2=0
cc_651 N_A_555_73#_c_762_n N_VPWR_c_1462_n 0.020016f $X=6.165 $Y=2.52 $X2=0
+ $Y2=0
cc_652 N_A_555_73#_c_735_n N_VPWR_c_1463_n 0.0134673f $X=8.145 $Y=2.98 $X2=0
+ $Y2=0
cc_653 N_A_555_73#_c_736_n N_VPWR_c_1463_n 0.0664508f $X=8.23 $Y=2.895 $X2=0
+ $Y2=0
cc_654 N_A_555_73#_c_716_n N_VPWR_c_1463_n 0.0119019f $X=8.755 $Y=1.675 $X2=0
+ $Y2=0
cc_655 N_A_555_73#_c_727_n N_VPWR_c_1465_n 0.0573512f $X=4.795 $Y=2.98 $X2=0
+ $Y2=0
cc_656 N_A_555_73#_c_728_n N_VPWR_c_1465_n 0.0113092f $X=4.025 $Y=2.98 $X2=0
+ $Y2=0
cc_657 N_A_555_73#_c_762_n N_VPWR_c_1465_n 0.00208901f $X=6.165 $Y=2.52 $X2=0
+ $Y2=0
cc_658 N_A_555_73#_M1030_g N_VPWR_c_1467_n 8.42392e-19 $X=6.23 $Y=2.365 $X2=0
+ $Y2=0
cc_659 N_A_555_73#_c_762_n N_VPWR_c_1467_n 0.00863735f $X=6.165 $Y=2.52 $X2=0
+ $Y2=0
cc_660 N_A_555_73#_c_732_n N_VPWR_c_1467_n 0.0557292f $X=7.265 $Y=2.98 $X2=0
+ $Y2=0
cc_661 N_A_555_73#_c_733_n N_VPWR_c_1467_n 0.0121364f $X=6.345 $Y=2.98 $X2=0
+ $Y2=0
cc_662 N_A_555_73#_c_735_n N_VPWR_c_1467_n 0.0540284f $X=8.145 $Y=2.98 $X2=0
+ $Y2=0
cc_663 N_A_555_73#_c_741_n N_VPWR_c_1467_n 0.0114282f $X=7.35 $Y=2.98 $X2=0
+ $Y2=0
cc_664 N_A_555_73#_M1020_g N_VPWR_c_1470_n 6.93234e-19 $X=9.77 $Y=2.395 $X2=0
+ $Y2=0
cc_665 N_A_555_73#_M1030_g N_VPWR_c_1460_n 3.28073e-19 $X=6.23 $Y=2.365 $X2=0
+ $Y2=0
cc_666 N_A_555_73#_c_727_n N_VPWR_c_1460_n 0.0347965f $X=4.795 $Y=2.98 $X2=0
+ $Y2=0
cc_667 N_A_555_73#_c_728_n N_VPWR_c_1460_n 0.00584408f $X=4.025 $Y=2.98 $X2=0
+ $Y2=0
cc_668 N_A_555_73#_c_762_n N_VPWR_c_1460_n 0.0237164f $X=6.165 $Y=2.52 $X2=0
+ $Y2=0
cc_669 N_A_555_73#_c_732_n N_VPWR_c_1460_n 0.034375f $X=7.265 $Y=2.98 $X2=0
+ $Y2=0
cc_670 N_A_555_73#_c_733_n N_VPWR_c_1460_n 0.00696477f $X=6.345 $Y=2.98 $X2=0
+ $Y2=0
cc_671 N_A_555_73#_c_735_n N_VPWR_c_1460_n 0.0330161f $X=8.145 $Y=2.98 $X2=0
+ $Y2=0
cc_672 N_A_555_73#_c_741_n N_VPWR_c_1460_n 0.00657239f $X=7.35 $Y=2.98 $X2=0
+ $Y2=0
cc_673 N_A_555_73#_c_742_n N_A_256_87#_c_1576_n 0.0118236f $X=3.045 $Y=2.55
+ $X2=0 $Y2=0
cc_674 N_A_555_73#_c_742_n N_A_256_87#_c_1569_n 0.0271806f $X=3.045 $Y=2.55
+ $X2=0 $Y2=0
cc_675 N_A_555_73#_c_711_n N_A_256_87#_c_1569_n 0.0311445f $X=3.185 $Y=0.78
+ $X2=0 $Y2=0
cc_676 N_A_555_73#_c_739_n N_A_256_87#_c_1569_n 0.017718f $X=3.045 $Y=2.04 $X2=0
+ $Y2=0
cc_677 N_A_555_73#_M1006_d N_A_256_87#_c_1598_n 0.00517636f $X=2.775 $Y=0.365
+ $X2=0 $Y2=0
cc_678 N_A_555_73#_c_711_n N_A_256_87#_c_1598_n 0.0167202f $X=3.185 $Y=0.78
+ $X2=0 $Y2=0
cc_679 N_A_555_73#_M1006_d N_A_256_87#_c_1570_n 0.00423552f $X=2.775 $Y=0.365
+ $X2=0 $Y2=0
cc_680 N_A_555_73#_c_711_n N_A_256_87#_c_1570_n 0.0126927f $X=3.185 $Y=0.78
+ $X2=0 $Y2=0
cc_681 N_A_555_73#_c_711_n N_A_256_87#_c_1572_n 0.0142363f $X=3.185 $Y=0.78
+ $X2=0 $Y2=0
cc_682 N_A_555_73#_M1006_d N_A_256_87#_c_1574_n 0.00169871f $X=2.775 $Y=0.365
+ $X2=0 $Y2=0
cc_683 N_A_555_73#_c_711_n N_A_256_87#_c_1574_n 0.0131302f $X=3.185 $Y=0.78
+ $X2=0 $Y2=0
cc_684 N_A_555_73#_c_762_n N_A_1152_389#_M1019_d 0.0117153f $X=6.165 $Y=2.52
+ $X2=0 $Y2=0
cc_685 N_A_555_73#_M1030_g N_A_1152_389#_c_1652_n 0.00320307f $X=6.23 $Y=2.365
+ $X2=0 $Y2=0
cc_686 N_A_555_73#_c_762_n N_A_1152_389#_c_1652_n 0.0130182f $X=6.165 $Y=2.52
+ $X2=0 $Y2=0
cc_687 N_A_555_73#_c_712_n N_A_1152_389#_c_1652_n 0.0538898f $X=6.255 $Y=1.62
+ $X2=0 $Y2=0
cc_688 N_A_555_73#_c_713_n N_A_1152_389#_c_1652_n 0.00236638f $X=6.255 $Y=1.62
+ $X2=0 $Y2=0
cc_689 N_A_555_73#_c_712_n N_A_1152_389#_c_1653_n 5.43431e-19 $X=6.255 $Y=1.62
+ $X2=0 $Y2=0
cc_690 N_A_555_73#_c_713_n N_A_1152_389#_c_1653_n 0.00228866f $X=6.255 $Y=1.62
+ $X2=0 $Y2=0
cc_691 N_A_555_73#_c_734_n N_COUT_M1030_d 0.015233f $X=7.35 $Y=2.895 $X2=0 $Y2=0
cc_692 N_A_555_73#_c_732_n N_COUT_c_1685_n 0.0242662f $X=7.265 $Y=2.98 $X2=0
+ $Y2=0
cc_693 N_A_555_73#_c_734_n N_COUT_c_1685_n 0.0301521f $X=7.35 $Y=2.895 $X2=0
+ $Y2=0
cc_694 N_A_555_73#_M1030_g N_COUT_c_1681_n 0.00604926f $X=6.23 $Y=2.365 $X2=0
+ $Y2=0
cc_695 N_A_555_73#_M1008_g N_COUT_c_1681_n 0.0037357f $X=7.425 $Y=0.635 $X2=0
+ $Y2=0
cc_696 N_A_555_73#_c_712_n N_COUT_c_1681_n 0.0520243f $X=6.255 $Y=1.62 $X2=0
+ $Y2=0
cc_697 N_A_555_73#_c_713_n N_COUT_c_1681_n 0.00325901f $X=6.255 $Y=1.62 $X2=0
+ $Y2=0
cc_698 N_A_555_73#_c_734_n N_COUT_c_1681_n 0.00558113f $X=7.35 $Y=2.895 $X2=0
+ $Y2=0
cc_699 N_A_555_73#_M1008_g COUT 0.0258832f $X=7.425 $Y=0.635 $X2=0 $Y2=0
cc_700 N_A_555_73#_c_714_n COUT 0.0113072f $X=7.515 $Y=1.28 $X2=0 $Y2=0
cc_701 N_A_555_73#_M1008_g N_COUT_c_1682_n 0.00324375f $X=7.425 $Y=0.635 $X2=0
+ $Y2=0
cc_702 N_A_555_73#_c_735_n N_A_1500_63#_M1029_d 0.00257746f $X=8.145 $Y=2.98
+ $X2=0 $Y2=0
cc_703 N_A_555_73#_M1008_g N_A_1500_63#_c_1719_n 0.0051447f $X=7.425 $Y=0.635
+ $X2=0 $Y2=0
cc_704 N_A_555_73#_c_734_n N_A_1500_63#_c_1721_n 0.056196f $X=7.35 $Y=2.895
+ $X2=0 $Y2=0
cc_705 N_A_555_73#_c_715_n N_A_1500_63#_c_1721_n 0.0020535f $X=7.515 $Y=1.28
+ $X2=0 $Y2=0
cc_706 N_A_555_73#_c_735_n N_A_1500_63#_c_1721_n 0.0209107f $X=8.145 $Y=2.98
+ $X2=0 $Y2=0
cc_707 N_A_555_73#_M1008_g N_A_1500_63#_c_1720_n 0.00307078f $X=7.425 $Y=0.635
+ $X2=0 $Y2=0
cc_708 N_A_555_73#_c_734_n N_A_1500_63#_c_1720_n 0.00730823f $X=7.35 $Y=2.895
+ $X2=0 $Y2=0
cc_709 N_A_555_73#_c_714_n N_A_1500_63#_c_1720_n 0.0447849f $X=7.515 $Y=1.28
+ $X2=0 $Y2=0
cc_710 N_A_555_73#_c_715_n N_A_1500_63#_c_1720_n 0.0026349f $X=7.515 $Y=1.28
+ $X2=0 $Y2=0
cc_711 N_A_555_73#_c_736_n N_A_1500_63#_c_1720_n 0.0672907f $X=8.23 $Y=2.895
+ $X2=0 $Y2=0
cc_712 N_A_555_73#_c_717_n N_A_1500_63#_c_1720_n 0.0115071f $X=8.315 $Y=1.675
+ $X2=0 $Y2=0
cc_713 N_A_555_73#_M1008_g N_A_1500_63#_c_1734_n 0.00122521f $X=7.425 $Y=0.635
+ $X2=0 $Y2=0
cc_714 N_A_555_73#_M1020_g N_A_1883_395#_c_1757_n 0.00974008f $X=9.77 $Y=2.395
+ $X2=0 $Y2=0
cc_715 N_A_555_73#_M1020_g N_A_1883_395#_c_1758_n 0.005159f $X=9.77 $Y=2.395
+ $X2=0 $Y2=0
cc_716 N_A_555_73#_c_718_n N_VGND_M1011_d 0.00917614f $X=8.84 $Y=1.59 $X2=0
+ $Y2=0
cc_717 N_A_555_73#_c_719_n N_VGND_M1011_d 0.00257008f $X=8.925 $Y=0.415 $X2=0
+ $Y2=0
cc_718 N_A_555_73#_c_718_n N_VGND_c_1818_n 0.0245013f $X=8.84 $Y=1.59 $X2=0
+ $Y2=0
cc_719 N_A_555_73#_c_719_n N_VGND_c_1818_n 0.024647f $X=8.925 $Y=0.415 $X2=0
+ $Y2=0
cc_720 N_A_555_73#_c_719_n N_VGND_c_1820_n 0.0114622f $X=8.925 $Y=0.415 $X2=0
+ $Y2=0
cc_721 N_A_555_73#_c_720_n N_VGND_c_1820_n 0.052114f $X=9.61 $Y=0.4 $X2=0 $Y2=0
cc_722 N_A_555_73#_c_721_n N_VGND_c_1820_n 0.00593319f $X=9.61 $Y=0.4 $X2=0
+ $Y2=0
cc_723 N_A_555_73#_M1008_g N_VGND_c_1824_n 0.00337135f $X=7.425 $Y=0.635 $X2=0
+ $Y2=0
cc_724 N_A_555_73#_M1008_g N_VGND_c_1826_n 0.00555452f $X=7.425 $Y=0.635 $X2=0
+ $Y2=0
cc_725 N_A_555_73#_c_719_n N_VGND_c_1826_n 0.00657784f $X=8.925 $Y=0.415 $X2=0
+ $Y2=0
cc_726 N_A_555_73#_c_720_n N_VGND_c_1826_n 0.0299744f $X=9.61 $Y=0.4 $X2=0 $Y2=0
cc_727 N_A_555_73#_c_721_n N_VGND_c_1826_n 0.00774851f $X=9.61 $Y=0.4 $X2=0
+ $Y2=0
cc_728 N_A_364_73#_c_981_n N_CIN_M1003_g 0.0212287f $X=7.375 $Y=1.76 $X2=0 $Y2=0
cc_729 N_A_364_73#_c_971_n N_CIN_M1003_g 0.00992847f $X=10.175 $Y=1.665 $X2=0
+ $Y2=0
cc_730 N_A_364_73#_c_971_n N_CIN_c_1203_n 0.00671808f $X=10.175 $Y=1.665 $X2=0
+ $Y2=0
cc_731 N_A_364_73#_c_971_n CIN 0.00247476f $X=10.175 $Y=1.665 $X2=0 $Y2=0
cc_732 N_A_364_73#_M1028_g N_A_1774_367#_M1017_g 0.013679f $X=10.255 $Y=0.995
+ $X2=0 $Y2=0
cc_733 N_A_364_73#_c_976_n N_A_1774_367#_M1017_g 0.00672066f $X=10.27 $Y=1.65
+ $X2=0 $Y2=0
cc_734 N_A_364_73#_M1028_g N_A_1774_367#_c_1282_n 2.50761e-19 $X=10.255 $Y=0.995
+ $X2=0 $Y2=0
cc_735 N_A_364_73#_c_971_n N_A_1774_367#_c_1274_n 0.0105413f $X=10.175 $Y=1.665
+ $X2=0 $Y2=0
cc_736 N_A_364_73#_c_971_n N_A_1774_367#_c_1266_n 0.0251205f $X=10.175 $Y=1.665
+ $X2=0 $Y2=0
cc_737 N_A_364_73#_c_971_n N_A_1774_367#_c_1267_n 0.0100513f $X=10.175 $Y=1.665
+ $X2=0 $Y2=0
cc_738 N_A_364_73#_M1024_g N_A_1774_367#_c_1276_n 0.00794256f $X=10.2 $Y=2.395
+ $X2=0 $Y2=0
cc_739 N_A_364_73#_M1024_g N_A_1774_367#_c_1277_n 0.00648172f $X=10.2 $Y=2.395
+ $X2=0 $Y2=0
cc_740 N_A_364_73#_c_976_n N_A_1774_367#_c_1269_n 8.27185e-19 $X=10.27 $Y=1.65
+ $X2=0 $Y2=0
cc_741 N_A_364_73#_M1024_g N_A_1926_135#_c_1364_n 0.00419434f $X=10.2 $Y=2.395
+ $X2=0 $Y2=0
cc_742 N_A_364_73#_M1028_g N_A_1926_135#_c_1364_n 0.00365511f $X=10.255 $Y=0.995
+ $X2=0 $Y2=0
cc_743 N_A_364_73#_c_971_n N_A_1926_135#_c_1364_n 0.0114068f $X=10.175 $Y=1.665
+ $X2=0 $Y2=0
cc_744 N_A_364_73#_c_974_n N_A_1926_135#_c_1364_n 5.62211e-19 $X=10.32 $Y=1.665
+ $X2=0 $Y2=0
cc_745 N_A_364_73#_c_976_n N_A_1926_135#_c_1364_n 9.53831e-19 $X=10.27 $Y=1.65
+ $X2=0 $Y2=0
cc_746 N_A_364_73#_c_977_n N_A_1926_135#_c_1364_n 0.0220364f $X=10.27 $Y=1.65
+ $X2=0 $Y2=0
cc_747 N_A_364_73#_M1028_g N_A_1926_135#_c_1380_n 0.00453443f $X=10.255 $Y=0.995
+ $X2=0 $Y2=0
cc_748 N_A_364_73#_c_971_n N_A_1926_135#_c_1380_n 0.00828603f $X=10.175 $Y=1.665
+ $X2=0 $Y2=0
cc_749 N_A_364_73#_c_976_n N_A_1926_135#_c_1380_n 0.00175589f $X=10.27 $Y=1.65
+ $X2=0 $Y2=0
cc_750 N_A_364_73#_c_977_n N_A_1926_135#_c_1380_n 0.00475191f $X=10.27 $Y=1.65
+ $X2=0 $Y2=0
cc_751 N_A_364_73#_M1028_g N_A_1926_135#_c_1365_n 0.0113081f $X=10.255 $Y=0.995
+ $X2=0 $Y2=0
cc_752 N_A_364_73#_M1028_g N_A_1926_135#_c_1366_n 0.00551905f $X=10.255 $Y=0.995
+ $X2=0 $Y2=0
cc_753 N_A_364_73#_M1028_g N_A_1926_135#_c_1368_n 4.17189e-19 $X=10.255 $Y=0.995
+ $X2=0 $Y2=0
cc_754 N_A_364_73#_M1024_g N_A_1926_135#_c_1389_n 0.0037427f $X=10.2 $Y=2.395
+ $X2=0 $Y2=0
cc_755 N_A_364_73#_c_971_n N_A_1926_135#_c_1389_n 0.00805591f $X=10.175 $Y=1.665
+ $X2=0 $Y2=0
cc_756 N_A_364_73#_c_977_n N_A_1926_135#_c_1389_n 0.00189377f $X=10.27 $Y=1.65
+ $X2=0 $Y2=0
cc_757 N_A_364_73#_c_971_n N_VPWR_c_1463_n 0.00136271f $X=10.175 $Y=1.665 $X2=0
+ $Y2=0
cc_758 N_A_364_73#_c_983_n N_VPWR_c_1467_n 6.63031e-19 $X=7.45 $Y=1.835 $X2=0
+ $Y2=0
cc_759 N_A_364_73#_M1024_g N_VPWR_c_1470_n 6.93234e-19 $X=10.2 $Y=2.395 $X2=0
+ $Y2=0
cc_760 N_A_364_73#_c_964_n N_A_256_87#_c_1575_n 0.0194589f $X=2.07 $Y=2.19 $X2=0
+ $Y2=0
cc_761 N_A_364_73#_c_968_n N_A_256_87#_c_1575_n 0.00230128f $X=1.825 $Y=1.665
+ $X2=0 $Y2=0
cc_762 N_A_364_73#_c_978_n N_A_256_87#_c_1575_n 0.0044098f $X=1.95 $Y=1.37 $X2=0
+ $Y2=0
cc_763 N_A_364_73#_M1026_s N_A_256_87#_c_1568_n 0.00974948f $X=1.82 $Y=0.365
+ $X2=0 $Y2=0
cc_764 N_A_364_73#_c_967_n N_A_256_87#_c_1568_n 0.00589823f $X=3.935 $Y=1.665
+ $X2=0 $Y2=0
cc_765 N_A_364_73#_c_968_n N_A_256_87#_c_1568_n 0.00144373f $X=1.825 $Y=1.665
+ $X2=0 $Y2=0
cc_766 N_A_364_73#_c_978_n N_A_256_87#_c_1568_n 0.0323636f $X=1.95 $Y=1.37 $X2=0
+ $Y2=0
cc_767 N_A_364_73#_M1021_s N_A_256_87#_c_1576_n 0.00583812f $X=1.925 $Y=2.035
+ $X2=0 $Y2=0
cc_768 N_A_364_73#_c_964_n N_A_256_87#_c_1576_n 0.0193144f $X=2.07 $Y=2.19 $X2=0
+ $Y2=0
cc_769 N_A_364_73#_c_964_n N_A_256_87#_c_1569_n 0.0306607f $X=2.07 $Y=2.19 $X2=0
+ $Y2=0
cc_770 N_A_364_73#_c_967_n N_A_256_87#_c_1569_n 0.0332146f $X=3.935 $Y=1.665
+ $X2=0 $Y2=0
cc_771 N_A_364_73#_c_968_n N_A_256_87#_c_1569_n 3.30859e-19 $X=1.825 $Y=1.665
+ $X2=0 $Y2=0
cc_772 N_A_364_73#_c_978_n N_A_256_87#_c_1569_n 0.0425632f $X=1.95 $Y=1.37 $X2=0
+ $Y2=0
cc_773 N_A_364_73#_c_968_n N_A_256_87#_c_1573_n 0.00125301f $X=1.825 $Y=1.665
+ $X2=0 $Y2=0
cc_774 N_A_364_73#_c_978_n N_A_256_87#_c_1573_n 4.24005e-19 $X=1.95 $Y=1.37
+ $X2=0 $Y2=0
cc_775 N_A_364_73#_c_967_n N_A_256_87#_c_1574_n 0.00825847f $X=3.935 $Y=1.665
+ $X2=0 $Y2=0
cc_776 N_A_364_73#_c_959_n N_A_1152_389#_c_1651_n 0.00579716f $X=6.235 $Y=1.065
+ $X2=0 $Y2=0
cc_777 N_A_364_73#_c_959_n N_A_1152_389#_c_1652_n 0.00242883f $X=6.235 $Y=1.065
+ $X2=0 $Y2=0
cc_778 N_A_364_73#_c_969_n N_A_1152_389#_c_1652_n 0.0211983f $X=6.815 $Y=1.665
+ $X2=0 $Y2=0
cc_779 N_A_364_73#_c_959_n N_A_1152_389#_c_1653_n 0.0029684f $X=6.235 $Y=1.065
+ $X2=0 $Y2=0
cc_780 N_A_364_73#_c_969_n N_A_1152_389#_c_1653_n 0.00607991f $X=6.815 $Y=1.665
+ $X2=0 $Y2=0
cc_781 N_A_364_73#_c_983_n N_COUT_c_1685_n 0.00396013f $X=7.45 $Y=1.835 $X2=0
+ $Y2=0
cc_782 N_A_364_73#_c_969_n N_COUT_c_1685_n 0.00596316f $X=6.815 $Y=1.665 $X2=0
+ $Y2=0
cc_783 N_A_364_73#_c_972_n N_COUT_c_1685_n 0.00212161f $X=7.105 $Y=1.665 $X2=0
+ $Y2=0
cc_784 N_A_364_73#_c_975_n N_COUT_c_1685_n 0.00129567f $X=6.975 $Y=1.14 $X2=0
+ $Y2=0
cc_785 N_A_364_73#_c_959_n N_COUT_c_1681_n 0.00371767f $X=6.235 $Y=1.065 $X2=0
+ $Y2=0
cc_786 N_A_364_73#_c_960_n N_COUT_c_1681_n 0.014588f $X=6.81 $Y=1.14 $X2=0 $Y2=0
cc_787 N_A_364_73#_c_962_n N_COUT_c_1681_n 0.00120542f $X=7.065 $Y=1.685 $X2=0
+ $Y2=0
cc_788 N_A_364_73#_c_982_n N_COUT_c_1681_n 6.84802e-19 $X=7.14 $Y=1.76 $X2=0
+ $Y2=0
cc_789 N_A_364_73#_c_983_n N_COUT_c_1681_n 5.45099e-19 $X=7.45 $Y=1.835 $X2=0
+ $Y2=0
cc_790 N_A_364_73#_c_966_n N_COUT_c_1681_n 0.0489993f $X=6.975 $Y=1.23 $X2=0
+ $Y2=0
cc_791 N_A_364_73#_c_969_n N_COUT_c_1681_n 0.0191804f $X=6.815 $Y=1.665 $X2=0
+ $Y2=0
cc_792 N_A_364_73#_c_972_n N_COUT_c_1681_n 0.00273887f $X=7.105 $Y=1.665 $X2=0
+ $Y2=0
cc_793 N_A_364_73#_c_975_n N_COUT_c_1681_n 0.00432988f $X=6.975 $Y=1.14 $X2=0
+ $Y2=0
cc_794 N_A_364_73#_c_966_n COUT 0.0209852f $X=6.975 $Y=1.23 $X2=0 $Y2=0
cc_795 N_A_364_73#_c_975_n COUT 0.00552322f $X=6.975 $Y=1.14 $X2=0 $Y2=0
cc_796 N_A_364_73#_c_959_n N_COUT_c_1682_n 0.0113369f $X=6.235 $Y=1.065 $X2=0
+ $Y2=0
cc_797 N_A_364_73#_c_960_n N_COUT_c_1682_n 0.0106892f $X=6.81 $Y=1.14 $X2=0
+ $Y2=0
cc_798 N_A_364_73#_c_983_n N_A_1500_63#_c_1721_n 0.00670059f $X=7.45 $Y=1.835
+ $X2=0 $Y2=0
cc_799 N_A_364_73#_c_971_n N_A_1500_63#_c_1721_n 0.00924338f $X=10.175 $Y=1.665
+ $X2=0 $Y2=0
cc_800 N_A_364_73#_c_981_n N_A_1500_63#_c_1720_n 0.0015624f $X=7.375 $Y=1.76
+ $X2=0 $Y2=0
cc_801 N_A_364_73#_c_966_n N_A_1500_63#_c_1720_n 0.00131404f $X=6.975 $Y=1.23
+ $X2=0 $Y2=0
cc_802 N_A_364_73#_c_971_n N_A_1500_63#_c_1720_n 0.023427f $X=10.175 $Y=1.665
+ $X2=0 $Y2=0
cc_803 N_A_364_73#_c_975_n N_A_1500_63#_c_1720_n 2.71911e-19 $X=6.975 $Y=1.14
+ $X2=0 $Y2=0
cc_804 N_A_364_73#_M1024_g N_A_1883_395#_c_1757_n 0.0149746f $X=10.2 $Y=2.395
+ $X2=0 $Y2=0
cc_805 N_A_364_73#_c_974_n N_A_1883_395#_c_1757_n 0.0024267f $X=10.32 $Y=1.665
+ $X2=0 $Y2=0
cc_806 N_A_364_73#_c_976_n N_A_1883_395#_c_1757_n 0.00260215f $X=10.27 $Y=1.65
+ $X2=0 $Y2=0
cc_807 N_A_364_73#_c_977_n N_A_1883_395#_c_1757_n 0.00592096f $X=10.27 $Y=1.65
+ $X2=0 $Y2=0
cc_808 N_A_364_73#_M1028_g N_A_1883_395#_c_1752_n 0.00714816f $X=10.255 $Y=0.995
+ $X2=0 $Y2=0
cc_809 N_A_364_73#_M1024_g N_A_1883_395#_c_1753_n 0.00933807f $X=10.2 $Y=2.395
+ $X2=0 $Y2=0
cc_810 N_A_364_73#_M1028_g N_A_1883_395#_c_1753_n 0.00355411f $X=10.255 $Y=0.995
+ $X2=0 $Y2=0
cc_811 N_A_364_73#_c_974_n N_A_1883_395#_c_1753_n 0.00742586f $X=10.32 $Y=1.665
+ $X2=0 $Y2=0
cc_812 N_A_364_73#_c_976_n N_A_1883_395#_c_1753_n 0.001186f $X=10.27 $Y=1.65
+ $X2=0 $Y2=0
cc_813 N_A_364_73#_c_977_n N_A_1883_395#_c_1753_n 0.0207418f $X=10.27 $Y=1.65
+ $X2=0 $Y2=0
cc_814 N_A_364_73#_M1024_g N_A_1883_395#_c_1758_n 8.64731e-19 $X=10.2 $Y=2.395
+ $X2=0 $Y2=0
cc_815 N_A_364_73#_c_974_n N_A_1883_395#_c_1754_n 0.00163359f $X=10.32 $Y=1.665
+ $X2=0 $Y2=0
cc_816 N_A_364_73#_c_976_n N_A_1883_395#_c_1754_n 3.24106e-19 $X=10.27 $Y=1.65
+ $X2=0 $Y2=0
cc_817 N_A_364_73#_c_977_n N_A_1883_395#_c_1754_n 0.00100164f $X=10.27 $Y=1.65
+ $X2=0 $Y2=0
cc_818 N_A_364_73#_M1024_g N_A_1883_395#_c_1756_n 0.0095034f $X=10.2 $Y=2.395
+ $X2=0 $Y2=0
cc_819 N_A_364_73#_M1028_g N_VGND_c_1820_n 2.04887e-19 $X=10.255 $Y=0.995 $X2=0
+ $Y2=0
cc_820 N_A_364_73#_c_959_n N_VGND_c_1824_n 0.00477421f $X=6.235 $Y=1.065 $X2=0
+ $Y2=0
cc_821 N_A_364_73#_c_959_n N_VGND_c_1826_n 0.00980949f $X=6.235 $Y=1.065 $X2=0
+ $Y2=0
cc_822 N_CIN_M1023_g N_A_1774_367#_c_1271_n 0.0103818f $X=8.795 $Y=2.465 $X2=0
+ $Y2=0
cc_823 N_CIN_c_1203_n N_A_1774_367#_c_1274_n 0.00532335f $X=8.795 $Y=1.415 $X2=0
+ $Y2=0
cc_824 N_CIN_M1023_g N_A_1774_367#_c_1274_n 0.00275293f $X=8.795 $Y=2.465 $X2=0
+ $Y2=0
cc_825 N_CIN_c_1203_n N_A_1774_367#_c_1266_n 0.00264515f $X=8.795 $Y=1.415 $X2=0
+ $Y2=0
cc_826 N_CIN_M1023_g N_A_1774_367#_c_1266_n 0.00679111f $X=8.795 $Y=2.465 $X2=0
+ $Y2=0
cc_827 N_CIN_c_1205_n N_A_1774_367#_c_1267_n 0.00264515f $X=9.01 $Y=1.265 $X2=0
+ $Y2=0
cc_828 N_CIN_M1003_g N_VPWR_c_1463_n 0.00194683f $X=7.995 $Y=2.445 $X2=0 $Y2=0
cc_829 N_CIN_M1023_g N_VPWR_c_1463_n 0.00493471f $X=8.795 $Y=2.465 $X2=0 $Y2=0
cc_830 N_CIN_M1003_g N_VPWR_c_1467_n 0.00389795f $X=7.995 $Y=2.445 $X2=0 $Y2=0
cc_831 N_CIN_M1023_g N_VPWR_c_1470_n 0.0054778f $X=8.795 $Y=2.465 $X2=0 $Y2=0
cc_832 N_CIN_M1003_g N_VPWR_c_1460_n 0.0054106f $X=7.995 $Y=2.445 $X2=0 $Y2=0
cc_833 N_CIN_M1023_g N_VPWR_c_1460_n 0.0123556f $X=8.795 $Y=2.465 $X2=0 $Y2=0
cc_834 N_CIN_c_1202_n N_A_1500_63#_c_1719_n 0.00728242f $X=8.115 $Y=1.08 $X2=0
+ $Y2=0
cc_835 N_CIN_M1003_g N_A_1500_63#_c_1721_n 0.0114689f $X=7.995 $Y=2.445 $X2=0
+ $Y2=0
cc_836 N_CIN_M1003_g N_A_1500_63#_c_1720_n 0.00875953f $X=7.995 $Y=2.445 $X2=0
+ $Y2=0
cc_837 N_CIN_c_1202_n N_A_1500_63#_c_1720_n 0.00766293f $X=8.115 $Y=1.08 $X2=0
+ $Y2=0
cc_838 N_CIN_c_1203_n N_A_1500_63#_c_1720_n 0.0100996f $X=8.795 $Y=1.415 $X2=0
+ $Y2=0
cc_839 CIN N_A_1500_63#_c_1720_n 0.017077f $X=8.315 $Y=1.21 $X2=0 $Y2=0
cc_840 N_CIN_c_1202_n N_A_1500_63#_c_1734_n 0.00607821f $X=8.115 $Y=1.08 $X2=0
+ $Y2=0
cc_841 N_CIN_c_1203_n N_A_1500_63#_c_1734_n 0.00161608f $X=8.795 $Y=1.415 $X2=0
+ $Y2=0
cc_842 N_CIN_M1023_g N_A_1883_395#_c_1758_n 4.03363e-19 $X=8.795 $Y=2.465 $X2=0
+ $Y2=0
cc_843 N_CIN_c_1202_n N_VGND_c_1818_n 0.0158334f $X=8.115 $Y=1.08 $X2=0 $Y2=0
cc_844 N_CIN_c_1203_n N_VGND_c_1818_n 0.00256652f $X=8.795 $Y=1.415 $X2=0 $Y2=0
cc_845 N_CIN_c_1205_n N_VGND_c_1818_n 0.00394027f $X=9.01 $Y=1.265 $X2=0 $Y2=0
cc_846 CIN N_VGND_c_1818_n 0.0259927f $X=8.315 $Y=1.21 $X2=0 $Y2=0
cc_847 N_CIN_c_1205_n N_VGND_c_1820_n 0.00309864f $X=9.01 $Y=1.265 $X2=0 $Y2=0
cc_848 N_CIN_c_1202_n N_VGND_c_1824_n 0.00477421f $X=8.115 $Y=1.08 $X2=0 $Y2=0
cc_849 N_CIN_c_1202_n N_VGND_c_1826_n 0.00992346f $X=8.115 $Y=1.08 $X2=0 $Y2=0
cc_850 N_CIN_c_1205_n N_VGND_c_1826_n 0.00564376f $X=9.01 $Y=1.265 $X2=0 $Y2=0
cc_851 N_A_1774_367#_M1017_g N_A_1926_135#_c_1363_n 0.00794016f $X=10.915
+ $Y=0.915 $X2=0 $Y2=0
cc_852 N_A_1774_367#_c_1273_n N_A_1926_135#_M1018_g 0.00141295f $X=11.425
+ $Y=2.895 $X2=0 $Y2=0
cc_853 N_A_1774_367#_c_1268_n N_A_1926_135#_M1018_g 8.66941e-19 $X=11.2 $Y=1.77
+ $X2=0 $Y2=0
cc_854 N_A_1774_367#_c_1269_n N_A_1926_135#_M1018_g 0.0164881f $X=11.2 $Y=1.77
+ $X2=0 $Y2=0
cc_855 N_A_1774_367#_c_1266_n N_A_1926_135#_c_1364_n 0.0223803f $X=9.067 $Y=1.94
+ $X2=0 $Y2=0
cc_856 N_A_1774_367#_c_1267_n N_A_1926_135#_c_1364_n 0.00169496f $X=9.312
+ $Y=1.335 $X2=0 $Y2=0
cc_857 N_A_1774_367#_c_1282_n N_A_1926_135#_c_1380_n 0.010058f $X=9.312 $Y=1.143
+ $X2=0 $Y2=0
cc_858 N_A_1774_367#_M1017_g N_A_1926_135#_c_1365_n 0.00218349f $X=10.915
+ $Y=0.915 $X2=0 $Y2=0
cc_859 N_A_1774_367#_c_1282_n N_A_1926_135#_c_1365_n 0.014119f $X=9.312 $Y=1.143
+ $X2=0 $Y2=0
cc_860 N_A_1774_367#_M1017_g N_A_1926_135#_c_1366_n 0.00602577f $X=10.915
+ $Y=0.915 $X2=0 $Y2=0
cc_861 N_A_1774_367#_M1017_g N_A_1926_135#_c_1368_n 0.0230022f $X=10.915
+ $Y=0.915 $X2=0 $Y2=0
cc_862 N_A_1774_367#_c_1268_n N_A_1926_135#_c_1369_n 0.0234136f $X=11.2 $Y=1.77
+ $X2=0 $Y2=0
cc_863 N_A_1774_367#_c_1269_n N_A_1926_135#_c_1369_n 0.00158541f $X=11.2 $Y=1.77
+ $X2=0 $Y2=0
cc_864 N_A_1774_367#_M1017_g N_A_1926_135#_c_1370_n 0.00630602f $X=10.915
+ $Y=0.915 $X2=0 $Y2=0
cc_865 N_A_1774_367#_c_1268_n N_A_1926_135#_c_1370_n 0.00825061f $X=11.2 $Y=1.77
+ $X2=0 $Y2=0
cc_866 N_A_1774_367#_c_1269_n N_A_1926_135#_c_1370_n 0.00261558f $X=11.2 $Y=1.77
+ $X2=0 $Y2=0
cc_867 N_A_1774_367#_c_1274_n N_A_1926_135#_c_1389_n 0.00649939f $X=9.01
+ $Y=2.105 $X2=0 $Y2=0
cc_868 N_A_1774_367#_M1017_g N_A_1926_135#_c_1371_n 9.95492e-19 $X=10.915
+ $Y=0.915 $X2=0 $Y2=0
cc_869 N_A_1774_367#_c_1268_n N_A_1926_135#_c_1371_n 0.00393751f $X=11.2 $Y=1.77
+ $X2=0 $Y2=0
cc_870 N_A_1774_367#_M1017_g N_A_1926_135#_c_1372_n 0.0049382f $X=10.915
+ $Y=0.915 $X2=0 $Y2=0
cc_871 N_A_1774_367#_c_1268_n N_A_1926_135#_c_1372_n 2.76493e-19 $X=11.2 $Y=1.77
+ $X2=0 $Y2=0
cc_872 N_A_1774_367#_c_1269_n N_A_1926_135#_c_1372_n 0.00373936f $X=11.2 $Y=1.77
+ $X2=0 $Y2=0
cc_873 N_A_1774_367#_c_1272_n N_VPWR_M1025_d 0.00252815f $X=11.34 $Y=2.98 $X2=0
+ $Y2=0
cc_874 N_A_1774_367#_c_1273_n N_VPWR_M1025_d 0.00748694f $X=11.425 $Y=2.895
+ $X2=0 $Y2=0
cc_875 N_A_1774_367#_M1025_g N_VPWR_c_1464_n 0.00238497f $X=11.29 $Y=2.595 $X2=0
+ $Y2=0
cc_876 N_A_1774_367#_c_1272_n N_VPWR_c_1464_n 0.0136053f $X=11.34 $Y=2.98 $X2=0
+ $Y2=0
cc_877 N_A_1774_367#_c_1273_n N_VPWR_c_1464_n 0.0623862f $X=11.425 $Y=2.895
+ $X2=0 $Y2=0
cc_878 N_A_1774_367#_c_1268_n N_VPWR_c_1464_n 0.0135103f $X=11.2 $Y=1.77 $X2=0
+ $Y2=0
cc_879 N_A_1774_367#_c_1269_n N_VPWR_c_1464_n 0.00351211f $X=11.2 $Y=1.77 $X2=0
+ $Y2=0
cc_880 N_A_1774_367#_M1025_g N_VPWR_c_1470_n 0.0035993f $X=11.29 $Y=2.595 $X2=0
+ $Y2=0
cc_881 N_A_1774_367#_c_1271_n N_VPWR_c_1470_n 0.0276229f $X=9.067 $Y=2.895 $X2=0
+ $Y2=0
cc_882 N_A_1774_367#_c_1272_n N_VPWR_c_1470_n 0.00928977f $X=11.34 $Y=2.98 $X2=0
+ $Y2=0
cc_883 N_A_1774_367#_c_1276_n N_VPWR_c_1470_n 0.123005f $X=10.36 $Y=2.9 $X2=0
+ $Y2=0
cc_884 N_A_1774_367#_M1023_d N_VPWR_c_1460_n 0.00223793f $X=8.87 $Y=1.835 $X2=0
+ $Y2=0
cc_885 N_A_1774_367#_M1025_g N_VPWR_c_1460_n 0.0074086f $X=11.29 $Y=2.595 $X2=0
+ $Y2=0
cc_886 N_A_1774_367#_c_1271_n N_VPWR_c_1460_n 0.0170251f $X=9.067 $Y=2.895 $X2=0
+ $Y2=0
cc_887 N_A_1774_367#_c_1272_n N_VPWR_c_1460_n 0.00645723f $X=11.34 $Y=2.98 $X2=0
+ $Y2=0
cc_888 N_A_1774_367#_c_1276_n N_VPWR_c_1460_n 0.0762176f $X=10.36 $Y=2.9 $X2=0
+ $Y2=0
cc_889 N_A_1774_367#_c_1272_n N_A_1883_395#_M1025_s 0.00549859f $X=11.34 $Y=2.98
+ $X2=0 $Y2=0
cc_890 N_A_1774_367#_M1024_d N_A_1883_395#_c_1757_n 0.0125345f $X=10.275
+ $Y=1.975 $X2=0 $Y2=0
cc_891 N_A_1774_367#_c_1276_n N_A_1883_395#_c_1757_n 0.0210188f $X=10.36 $Y=2.9
+ $X2=0 $Y2=0
cc_892 N_A_1774_367#_c_1277_n N_A_1883_395#_c_1757_n 0.0179895f $X=10.69 $Y=2.9
+ $X2=0 $Y2=0
cc_893 N_A_1774_367#_M1024_d N_A_1883_395#_c_1753_n 0.00374237f $X=10.275
+ $Y=1.975 $X2=0 $Y2=0
cc_894 N_A_1774_367#_M1025_g N_A_1883_395#_c_1753_n 0.00341452f $X=11.29
+ $Y=2.595 $X2=0 $Y2=0
cc_895 N_A_1774_367#_c_1273_n N_A_1883_395#_c_1753_n 0.00525457f $X=11.425
+ $Y=2.895 $X2=0 $Y2=0
cc_896 N_A_1774_367#_c_1268_n N_A_1883_395#_c_1753_n 0.0237464f $X=11.2 $Y=1.77
+ $X2=0 $Y2=0
cc_897 N_A_1774_367#_c_1269_n N_A_1883_395#_c_1753_n 0.0073273f $X=11.2 $Y=1.77
+ $X2=0 $Y2=0
cc_898 N_A_1774_367#_c_1271_n N_A_1883_395#_c_1758_n 0.0259752f $X=9.067
+ $Y=2.895 $X2=0 $Y2=0
cc_899 N_A_1774_367#_c_1276_n N_A_1883_395#_c_1758_n 0.0152912f $X=10.36 $Y=2.9
+ $X2=0 $Y2=0
cc_900 N_A_1774_367#_M1017_g N_A_1883_395#_c_1754_n 0.00630592f $X=10.915
+ $Y=0.915 $X2=0 $Y2=0
cc_901 N_A_1774_367#_M1024_d N_A_1883_395#_c_1756_n 0.00427433f $X=10.275
+ $Y=1.975 $X2=0 $Y2=0
cc_902 N_A_1774_367#_c_1272_n N_A_1883_395#_c_1756_n 0.0273101f $X=11.34 $Y=2.98
+ $X2=0 $Y2=0
cc_903 N_A_1774_367#_c_1277_n N_A_1883_395#_c_1756_n 0.00592503f $X=10.69 $Y=2.9
+ $X2=0 $Y2=0
cc_904 N_A_1774_367#_c_1268_n N_A_1883_395#_c_1756_n 0.0103187f $X=11.2 $Y=1.77
+ $X2=0 $Y2=0
cc_905 N_A_1774_367#_c_1269_n N_A_1883_395#_c_1756_n 0.00717505f $X=11.2 $Y=1.77
+ $X2=0 $Y2=0
cc_906 N_A_1774_367#_M1017_g N_VGND_c_1819_n 0.00198731f $X=10.915 $Y=0.915
+ $X2=0 $Y2=0
cc_907 N_A_1774_367#_M1017_g N_VGND_c_1820_n 2.4468e-19 $X=10.915 $Y=0.915 $X2=0
+ $Y2=0
cc_908 N_A_1926_135#_M1018_g N_VPWR_c_1464_n 0.0217229f $X=11.99 $Y=2.465 $X2=0
+ $Y2=0
cc_909 N_A_1926_135#_c_1371_n N_VPWR_c_1464_n 0.017453f $X=11.775 $Y=1.34 $X2=0
+ $Y2=0
cc_910 N_A_1926_135#_c_1372_n N_VPWR_c_1464_n 0.0015674f $X=11.99 $Y=1.51 $X2=0
+ $Y2=0
cc_911 N_A_1926_135#_M1018_g N_VPWR_c_1471_n 0.00486043f $X=11.99 $Y=2.465 $X2=0
+ $Y2=0
cc_912 N_A_1926_135#_M1018_g N_VPWR_c_1460_n 0.00919377f $X=11.99 $Y=2.465 $X2=0
+ $Y2=0
cc_913 N_A_1926_135#_M1020_d N_A_1883_395#_c_1757_n 0.00418283f $X=9.845
+ $Y=1.975 $X2=0 $Y2=0
cc_914 N_A_1926_135#_c_1389_n N_A_1883_395#_c_1757_n 0.0189039f $X=9.985 $Y=2.12
+ $X2=0 $Y2=0
cc_915 N_A_1926_135#_c_1365_n N_A_1883_395#_c_1752_n 0.0333521f $X=10.04 $Y=0.98
+ $X2=0 $Y2=0
cc_916 N_A_1926_135#_c_1366_n N_A_1883_395#_c_1752_n 0.0268637f $X=10.965
+ $Y=0.35 $X2=0 $Y2=0
cc_917 N_A_1926_135#_c_1389_n N_A_1883_395#_c_1753_n 0.00577441f $X=9.985
+ $Y=2.12 $X2=0 $Y2=0
cc_918 N_A_1926_135#_c_1380_n N_A_1883_395#_c_1754_n 0.0112705f $X=10.08
+ $Y=1.135 $X2=0 $Y2=0
cc_919 N_A_1926_135#_c_1368_n N_A_1883_395#_c_1754_n 0.0214565f $X=11.05
+ $Y=1.255 $X2=0 $Y2=0
cc_920 N_A_1926_135#_c_1370_n N_A_1883_395#_c_1754_n 0.0131379f $X=11.135
+ $Y=1.34 $X2=0 $Y2=0
cc_921 N_A_1926_135#_c_1363_n SUM 0.005843f $X=11.775 $Y=1.345 $X2=0 $Y2=0
cc_922 N_A_1926_135#_c_1371_n SUM 0.0315208f $X=11.775 $Y=1.34 $X2=0 $Y2=0
cc_923 N_A_1926_135#_c_1372_n SUM 0.018341f $X=11.99 $Y=1.51 $X2=0 $Y2=0
cc_924 N_A_1926_135#_c_1363_n N_SUM_c_1802_n 0.00866446f $X=11.775 $Y=1.345
+ $X2=0 $Y2=0
cc_925 N_A_1926_135#_c_1371_n N_SUM_c_1802_n 0.0069456f $X=11.775 $Y=1.34 $X2=0
+ $Y2=0
cc_926 N_A_1926_135#_c_1372_n N_SUM_c_1802_n 0.00586694f $X=11.99 $Y=1.51 $X2=0
+ $Y2=0
cc_927 N_A_1926_135#_c_1368_n N_VGND_M1017_d 0.00734574f $X=11.05 $Y=1.255 $X2=0
+ $Y2=0
cc_928 N_A_1926_135#_c_1363_n N_VGND_c_1819_n 0.0118704f $X=11.775 $Y=1.345
+ $X2=0 $Y2=0
cc_929 N_A_1926_135#_c_1366_n N_VGND_c_1819_n 0.014441f $X=10.965 $Y=0.35 $X2=0
+ $Y2=0
cc_930 N_A_1926_135#_c_1368_n N_VGND_c_1819_n 0.0473041f $X=11.05 $Y=1.255 $X2=0
+ $Y2=0
cc_931 N_A_1926_135#_c_1369_n N_VGND_c_1819_n 0.0233169f $X=11.61 $Y=1.34 $X2=0
+ $Y2=0
cc_932 N_A_1926_135#_c_1371_n N_VGND_c_1819_n 0.00276232f $X=11.775 $Y=1.34
+ $X2=0 $Y2=0
cc_933 N_A_1926_135#_c_1372_n N_VGND_c_1819_n 2.04868e-19 $X=11.99 $Y=1.51 $X2=0
+ $Y2=0
cc_934 N_A_1926_135#_c_1366_n N_VGND_c_1820_n 0.0574898f $X=10.965 $Y=0.35 $X2=0
+ $Y2=0
cc_935 N_A_1926_135#_c_1367_n N_VGND_c_1820_n 0.0168561f $X=10.205 $Y=0.35 $X2=0
+ $Y2=0
cc_936 N_A_1926_135#_c_1363_n N_VGND_c_1825_n 0.00534051f $X=11.775 $Y=1.345
+ $X2=0 $Y2=0
cc_937 N_A_1926_135#_c_1363_n N_VGND_c_1826_n 0.00537853f $X=11.775 $Y=1.345
+ $X2=0 $Y2=0
cc_938 N_A_1926_135#_c_1366_n N_VGND_c_1826_n 0.0349731f $X=10.965 $Y=0.35 $X2=0
+ $Y2=0
cc_939 N_A_1926_135#_c_1367_n N_VGND_c_1826_n 0.00967329f $X=10.205 $Y=0.35
+ $X2=0 $Y2=0
cc_940 N_VPWR_c_1460_n N_A_1883_395#_M1025_s 0.00228827f $X=12.24 $Y=3.33 $X2=0
+ $Y2=0
cc_941 N_VPWR_c_1460_n N_SUM_M1018_d 0.00419266f $X=12.24 $Y=3.33 $X2=0 $Y2=0
cc_942 N_VPWR_c_1471_n SUM 0.0163841f $X=12.24 $Y=3.33 $X2=0 $Y2=0
cc_943 N_VPWR_c_1460_n SUM 0.00959046f $X=12.24 $Y=3.33 $X2=0 $Y2=0
cc_944 N_A_256_87#_c_1570_n N_VGND_c_1823_n 0.0489186f $X=3.45 $Y=0.35 $X2=0
+ $Y2=0
cc_945 N_A_256_87#_c_1571_n N_VGND_c_1823_n 0.0112553f $X=2.92 $Y=0.35 $X2=0
+ $Y2=0
cc_946 N_A_256_87#_c_1568_n N_VGND_c_1826_n 0.0079269f $X=2.335 $Y=0.94 $X2=0
+ $Y2=0
cc_947 N_A_256_87#_c_1570_n N_VGND_c_1826_n 0.0263614f $X=3.45 $Y=0.35 $X2=0
+ $Y2=0
cc_948 N_A_256_87#_c_1571_n N_VGND_c_1826_n 0.00583019f $X=2.92 $Y=0.35 $X2=0
+ $Y2=0
cc_949 N_A_1152_389#_c_1652_n N_COUT_c_1681_n 0.0155954f $X=5.9 $Y=2.09 $X2=0
+ $Y2=0
cc_950 N_A_1152_389#_c_1653_n N_COUT_c_1681_n 0.00396362f $X=6 $Y=0.975 $X2=0
+ $Y2=0
cc_951 N_A_1152_389#_c_1651_n N_COUT_c_1682_n 0.022229f $X=6.02 $Y=0.46 $X2=0
+ $Y2=0
cc_952 N_A_1152_389#_c_1651_n N_VGND_c_1817_n 0.0200957f $X=6.02 $Y=0.46 $X2=0
+ $Y2=0
cc_953 N_A_1152_389#_c_1651_n N_VGND_c_1824_n 0.0207498f $X=6.02 $Y=0.46 $X2=0
+ $Y2=0
cc_954 N_A_1152_389#_c_1651_n N_VGND_c_1826_n 0.0136103f $X=6.02 $Y=0.46 $X2=0
+ $Y2=0
cc_955 COUT N_VGND_c_1824_n 0.0245596f $X=7.355 $Y=0.47 $X2=0 $Y2=0
cc_956 N_COUT_c_1682_n N_VGND_c_1824_n 0.0185698f $X=6.695 $Y=0.59 $X2=0 $Y2=0
cc_957 COUT N_VGND_c_1826_n 0.0287268f $X=7.355 $Y=0.47 $X2=0 $Y2=0
cc_958 N_COUT_c_1682_n N_VGND_c_1826_n 0.0125141f $X=6.695 $Y=0.59 $X2=0 $Y2=0
cc_959 N_A_1500_63#_c_1719_n N_VGND_c_1818_n 0.0224074f $X=7.9 $Y=0.615 $X2=0
+ $Y2=0
cc_960 N_A_1500_63#_c_1719_n N_VGND_c_1824_n 0.0186334f $X=7.9 $Y=0.615 $X2=0
+ $Y2=0
cc_961 N_A_1500_63#_c_1719_n N_VGND_c_1826_n 0.0123754f $X=7.9 $Y=0.615 $X2=0
+ $Y2=0
cc_962 N_SUM_c_1802_n N_VGND_c_1819_n 0.0278485f $X=11.99 $Y=0.54 $X2=0 $Y2=0
cc_963 N_SUM_c_1802_n N_VGND_c_1825_n 0.0219719f $X=11.99 $Y=0.54 $X2=0 $Y2=0
cc_964 N_SUM_c_1802_n N_VGND_c_1826_n 0.0197403f $X=11.99 $Y=0.54 $X2=0 $Y2=0
