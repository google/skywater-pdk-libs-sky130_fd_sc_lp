* File: sky130_fd_sc_lp__or3_4.spice
* Created: Fri Aug 28 11:23:26 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__or3_4.pex.spice"
.subckt sky130_fd_sc_lp__or3_4  VNB VPB C B A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* B	B
* C	C
* VPB	VPB
* VNB	VNB
MM1001 N_VGND_M1001_d N_C_M1001_g N_A_77_49#_M1001_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1512 AS=0.2226 PD=1.2 PS=2.21 NRD=4.992 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75003 A=0.126 P=1.98 MULT=1
MM1006 N_A_77_49#_M1006_d N_B_M1006_g N_VGND_M1001_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1512 PD=1.12 PS=1.2 NRD=0 NRS=6.42 M=1 R=5.6 SA=75000.7
+ SB=75002.4 A=0.126 P=1.98 MULT=1
MM1013 N_VGND_M1013_d N_A_M1013_g N_A_77_49#_M1006_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1617 AS=0.1176 PD=1.225 PS=1.12 NRD=7.14 NRS=0 M=1 R=5.6 SA=75001.1
+ SB=75002 A=0.126 P=1.98 MULT=1
MM1004 N_X_M1004_d N_A_77_49#_M1004_g N_VGND_M1013_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1617 PD=1.12 PS=1.225 NRD=0 NRS=7.848 M=1 R=5.6 SA=75001.7
+ SB=75001.5 A=0.126 P=1.98 MULT=1
MM1008 N_X_M1004_d N_A_77_49#_M1008_g N_VGND_M1008_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002.1
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1009 N_X_M1009_d N_A_77_49#_M1009_g N_VGND_M1008_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002.5
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1012 N_X_M1009_d N_A_77_49#_M1012_g N_VGND_M1012_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75003 SB=75000.2
+ A=0.126 P=1.98 MULT=1
MM1000 A_160_367# N_C_M1000_g N_A_77_49#_M1000_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1323 AS=0.3339 PD=1.47 PS=3.05 NRD=7.8012 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75003 A=0.189 P=2.82 MULT=1
MM1003 A_232_367# N_B_M1003_g A_160_367# VPB PHIGHVT L=0.15 W=1.26 AD=0.2457
+ AS=0.1323 PD=1.65 PS=1.47 NRD=21.8867 NRS=7.8012 M=1 R=8.4 SA=75000.6
+ SB=75002.6 A=0.189 P=2.82 MULT=1
MM1007 N_VPWR_M1007_d N_A_M1007_g A_232_367# VPB PHIGHVT L=0.15 W=1.26
+ AD=0.26775 AS=0.2457 PD=1.685 PS=1.65 NRD=10.9335 NRS=21.8867 M=1 R=8.4
+ SA=75001.1 SB=75002.1 A=0.189 P=2.82 MULT=1
MM1002 N_X_M1002_d N_A_77_49#_M1002_g N_VPWR_M1007_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.26775 PD=1.54 PS=1.685 NRD=0 NRS=11.7215 M=1 R=8.4 SA=75001.7
+ SB=75001.5 A=0.189 P=2.82 MULT=1
MM1005 N_X_M1002_d N_A_77_49#_M1005_g N_VPWR_M1005_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.1
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1010 N_X_M1010_d N_A_77_49#_M1010_g N_VPWR_M1005_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.5
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1011 N_X_M1010_d N_A_77_49#_M1011_g N_VPWR_M1011_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75003 SB=75000.2
+ A=0.189 P=2.82 MULT=1
DX14_noxref VNB VPB NWDIODE A=8.7655 P=13.13
*
.include "sky130_fd_sc_lp__or3_4.pxi.spice"
*
.ends
*
*
