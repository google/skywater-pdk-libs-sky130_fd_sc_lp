* File: sky130_fd_sc_lp__and3b_lp.pex.spice
* Created: Fri Aug 28 10:06:59 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__AND3B_LP%A_N 1 3 6 8 10 12 14 17 18 19 23 24
r42 23 24 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.29
+ $Y=1.07 $X2=0.29 $Y2=1.07
r43 18 19 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.29 $Y=1.295
+ $X2=0.29 $Y2=1.665
r44 18 24 7.85757 $w=3.28e-07 $l=2.25e-07 $layer=LI1_cond $X=0.29 $Y=1.295
+ $X2=0.29 $Y2=1.07
r45 16 23 42.9206 $w=4.6e-07 $l=3.55e-07 $layer=POLY_cond $X=0.355 $Y=1.425
+ $X2=0.355 $Y2=1.07
r46 16 17 29.6465 $w=4.6e-07 $l=1.5e-07 $layer=POLY_cond $X=0.405 $Y=1.425
+ $X2=0.405 $Y2=1.575
r47 13 23 16.9264 $w=4.6e-07 $l=1.4e-07 $layer=POLY_cond $X=0.355 $Y=0.93
+ $X2=0.355 $Y2=1.07
r48 13 14 10.9339 $w=3.05e-07 $l=7.5e-08 $layer=POLY_cond $X=0.355 $Y=0.93
+ $X2=0.355 $Y2=0.855
r49 10 12 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.885 $Y=0.78
+ $X2=0.885 $Y2=0.495
r50 9 14 15.748 $w=1.5e-07 $l=2.3e-07 $layer=POLY_cond $X=0.585 $Y=0.855
+ $X2=0.355 $Y2=0.855
r51 8 10 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.81 $Y=0.855
+ $X2=0.885 $Y2=0.78
r52 8 9 115.372 $w=1.5e-07 $l=2.25e-07 $layer=POLY_cond $X=0.81 $Y=0.855
+ $X2=0.585 $Y2=0.855
r53 6 17 239.758 $w=2.5e-07 $l=9.65e-07 $layer=POLY_cond $X=0.56 $Y=2.54
+ $X2=0.56 $Y2=1.575
r54 1 14 10.9339 $w=3.05e-07 $l=1.73494e-07 $layer=POLY_cond $X=0.495 $Y=0.78
+ $X2=0.355 $Y2=0.855
r55 1 3 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.495 $Y=0.78 $X2=0.495
+ $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__AND3B_LP%A_137_408# 1 2 9 13 15 18 22 24 28 32 34 35
+ 39
r61 35 40 59.3755 $w=7.2e-07 $l=5.05e-07 $layer=POLY_cond $X=1.415 $Y=1.335
+ $X2=1.415 $Y2=1.84
r62 35 39 50.9599 $w=7.2e-07 $l=1.65e-07 $layer=POLY_cond $X=1.415 $Y=1.335
+ $X2=1.415 $Y2=1.17
r63 34 37 17.1263 $w=5.63e-07 $l=5.05e-07 $layer=LI1_cond $X=1.102 $Y=1.335
+ $X2=1.102 $Y2=1.84
r64 34 36 4.06573 $w=5.63e-07 $l=1.65e-07 $layer=LI1_cond $X=1.102 $Y=1.335
+ $X2=1.102 $Y2=1.17
r65 34 35 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.22
+ $Y=1.335 $X2=1.22 $Y2=1.335
r66 32 37 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=0.905 $Y=2.02
+ $X2=0.905 $Y2=1.84
r67 28 36 17.4809 $w=4.43e-07 $l=6.75e-07 $layer=LI1_cond $X=1.042 $Y=0.495
+ $X2=1.042 $Y2=1.17
r68 22 32 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.825 $Y=2.185
+ $X2=0.825 $Y2=2.02
r69 22 24 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=0.825 $Y=2.185
+ $X2=0.825 $Y2=2.895
r70 16 18 92.2979 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=1.7 $Y=0.855
+ $X2=1.88 $Y2=0.855
r71 13 18 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.88 $Y=0.78
+ $X2=1.88 $Y2=0.855
r72 13 15 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=1.88 $Y=0.78 $X2=1.88
+ $Y2=0.495
r73 11 16 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.7 $Y=0.93 $X2=1.7
+ $Y2=0.855
r74 11 39 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=1.7 $Y=0.93 $X2=1.7
+ $Y2=1.17
r75 9 40 175.16 $w=2.5e-07 $l=7.05e-07 $layer=POLY_cond $X=1.65 $Y=2.545
+ $X2=1.65 $Y2=1.84
r76 2 24 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=0.685
+ $Y=2.04 $X2=0.825 $Y2=2.895
r77 2 22 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.685
+ $Y=2.04 $X2=0.825 $Y2=2.185
r78 1 28 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.96
+ $Y=0.285 $X2=1.1 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__AND3B_LP%B 1 3 7 11 12 14 21 22
r44 21 22 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.18
+ $Y=1.335 $X2=2.18 $Y2=1.335
r45 14 22 0.357038 $w=6.68e-07 $l=2e-08 $layer=LI1_cond $X=2.16 $Y=1.505
+ $X2=2.18 $Y2=1.505
r46 12 14 8.56892 $w=6.68e-07 $l=4.8e-07 $layer=LI1_cond $X=1.68 $Y=1.505
+ $X2=2.16 $Y2=1.505
r47 11 21 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.18 $Y=1.675
+ $X2=2.18 $Y2=1.335
r48 10 21 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.18 $Y=1.17
+ $X2=2.18 $Y2=1.335
r49 7 10 346.117 $w=1.5e-07 $l=6.75e-07 $layer=POLY_cond $X=2.27 $Y=0.495
+ $X2=2.27 $Y2=1.17
r50 1 11 30.6163 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.18 $Y=1.84
+ $X2=2.18 $Y2=1.675
r51 1 3 175.16 $w=2.5e-07 $l=7.05e-07 $layer=POLY_cond $X=2.18 $Y=1.84 $X2=2.18
+ $Y2=2.545
.ends

.subckt PM_SKY130_FD_SC_LP__AND3B_LP%C 3 7 11 12 13 14 18
r46 18 19 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.75
+ $Y=1.335 $X2=2.75 $Y2=1.335
r47 14 19 9.75144 $w=3.88e-07 $l=3.3e-07 $layer=LI1_cond $X=2.72 $Y=1.665
+ $X2=2.72 $Y2=1.335
r48 13 19 1.18199 $w=3.88e-07 $l=4e-08 $layer=LI1_cond $X=2.72 $Y=1.295 $X2=2.72
+ $Y2=1.335
r49 11 18 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.75 $Y=1.675
+ $X2=2.75 $Y2=1.335
r50 11 12 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.75 $Y=1.675
+ $X2=2.75 $Y2=1.84
r51 10 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.75 $Y=1.17
+ $X2=2.75 $Y2=1.335
r52 7 12 175.16 $w=2.5e-07 $l=7.05e-07 $layer=POLY_cond $X=2.71 $Y=2.545
+ $X2=2.71 $Y2=1.84
r53 3 10 346.117 $w=1.5e-07 $l=6.75e-07 $layer=POLY_cond $X=2.66 $Y=0.495
+ $X2=2.66 $Y2=1.17
.ends

.subckt PM_SKY130_FD_SC_LP__AND3B_LP%A_248_409# 1 2 3 10 12 15 17 19 24 28 30 31
+ 32 33 38 40 42 43 45 46 49 50
r113 49 52 65.7961 $w=5.35e-07 $l=5.05e-07 $layer=POLY_cond $X=3.422 $Y=0.985
+ $X2=3.422 $Y2=1.49
r114 48 49 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.32
+ $Y=0.985 $X2=3.32 $Y2=0.985
r115 45 50 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=3.18 $Y=2.02
+ $X2=3.18 $Y2=1.49
r116 43 50 9.49412 $w=3.88e-07 $l=1.95e-07 $layer=LI1_cond $X=3.29 $Y=1.295
+ $X2=3.29 $Y2=1.49
r117 42 48 2.51472 $w=3.9e-07 $l=8.5e-08 $layer=LI1_cond $X=3.29 $Y=0.99
+ $X2=3.29 $Y2=0.905
r118 42 43 9.0127 $w=3.88e-07 $l=3.05e-07 $layer=LI1_cond $X=3.29 $Y=0.99
+ $X2=3.29 $Y2=1.295
r119 41 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.61 $Y=2.105
+ $X2=2.445 $Y2=2.105
r120 40 45 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.095 $Y=2.105
+ $X2=3.18 $Y2=2.02
r121 40 41 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=3.095 $Y=2.105
+ $X2=2.61 $Y2=2.105
r122 36 46 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.445 $Y=2.19
+ $X2=2.445 $Y2=2.105
r123 36 38 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=2.445 $Y=2.19
+ $X2=2.445 $Y2=2.9
r124 32 48 5.76906 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=3.095 $Y=0.905
+ $X2=3.29 $Y2=0.905
r125 32 33 82.5294 $w=1.68e-07 $l=1.265e-06 $layer=LI1_cond $X=3.095 $Y=0.905
+ $X2=1.83 $Y2=0.905
r126 30 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.28 $Y=2.105
+ $X2=2.445 $Y2=2.105
r127 30 31 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=2.28 $Y=2.105
+ $X2=1.55 $Y2=2.105
r128 26 33 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.665 $Y=0.82
+ $X2=1.83 $Y2=0.905
r129 26 28 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=1.665 $Y=0.82
+ $X2=1.665 $Y2=0.495
r130 22 31 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.385 $Y=2.19
+ $X2=1.55 $Y2=2.105
r131 22 24 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=1.385 $Y=2.19
+ $X2=1.385 $Y2=2.9
r132 17 49 31.8222 $w=2.67e-07 $l=2.62857e-07 $layer=POLY_cond $X=3.615 $Y=0.82
+ $X2=3.422 $Y2=0.985
r133 17 19 104.433 $w=1.5e-07 $l=3.25e-07 $layer=POLY_cond $X=3.615 $Y=0.82
+ $X2=3.615 $Y2=0.495
r134 15 52 262.119 $w=2.5e-07 $l=1.055e-06 $layer=POLY_cond $X=3.345 $Y=2.545
+ $X2=3.345 $Y2=1.49
r135 10 49 31.8222 $w=2.67e-07 $l=2.35465e-07 $layer=POLY_cond $X=3.255 $Y=0.82
+ $X2=3.422 $Y2=0.985
r136 10 12 104.433 $w=1.5e-07 $l=3.25e-07 $layer=POLY_cond $X=3.255 $Y=0.82
+ $X2=3.255 $Y2=0.495
r137 3 38 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=2.305
+ $Y=2.045 $X2=2.445 $Y2=2.9
r138 3 36 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.305
+ $Y=2.045 $X2=2.445 $Y2=2.19
r139 2 24 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=1.24
+ $Y=2.045 $X2=1.385 $Y2=2.9
r140 2 22 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=1.24
+ $Y=2.045 $X2=1.385 $Y2=2.19
r141 1 28 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=1.52
+ $Y=0.285 $X2=1.665 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__AND3B_LP%VPWR 1 2 3 10 12 18 22 25 26 27 36 42 43 49
r47 49 50 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r48 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r49 43 50 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.12 $Y2=3.33
r50 42 43 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r51 40 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.14 $Y=3.33
+ $X2=2.975 $Y2=3.33
r52 40 42 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=3.14 $Y=3.33
+ $X2=4.08 $Y2=3.33
r53 39 50 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r54 38 39 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r55 36 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.81 $Y=3.33
+ $X2=2.975 $Y2=3.33
r56 36 38 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=2.81 $Y=3.33
+ $X2=2.64 $Y2=3.33
r57 34 35 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r58 32 35 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r59 32 47 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r60 31 34 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.72 $Y=3.33 $X2=1.68
+ $Y2=3.33
r61 31 32 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r62 29 46 4.70058 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=0.46 $Y=3.33 $X2=0.23
+ $Y2=3.33
r63 29 31 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=0.46 $Y=3.33
+ $X2=0.72 $Y2=3.33
r64 27 39 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r65 27 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r66 25 34 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=1.75 $Y=3.33 $X2=1.68
+ $Y2=3.33
r67 25 26 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.75 $Y=3.33
+ $X2=1.915 $Y2=3.33
r68 24 38 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=2.08 $Y=3.33
+ $X2=2.64 $Y2=3.33
r69 24 26 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.08 $Y=3.33
+ $X2=1.915 $Y2=3.33
r70 20 49 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.975 $Y=3.245
+ $X2=2.975 $Y2=3.33
r71 20 22 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=2.975 $Y=3.245
+ $X2=2.975 $Y2=2.535
r72 16 26 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.915 $Y=3.245
+ $X2=1.915 $Y2=3.33
r73 16 18 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=1.915 $Y=3.245
+ $X2=1.915 $Y2=2.535
r74 12 15 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=0.295 $Y=2.185
+ $X2=0.295 $Y2=2.895
r75 10 46 3.0656 $w=3.3e-07 $l=1.12916e-07 $layer=LI1_cond $X=0.295 $Y=3.245
+ $X2=0.23 $Y2=3.33
r76 10 15 12.2229 $w=3.28e-07 $l=3.5e-07 $layer=LI1_cond $X=0.295 $Y=3.245
+ $X2=0.295 $Y2=2.895
r77 3 22 300 $w=1.7e-07 $l=5.55608e-07 $layer=licon1_PDIFF $count=2 $X=2.835
+ $Y=2.045 $X2=2.975 $Y2=2.535
r78 2 18 300 $w=1.7e-07 $l=5.55608e-07 $layer=licon1_PDIFF $count=2 $X=1.775
+ $Y=2.045 $X2=1.915 $Y2=2.535
r79 1 15 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.15
+ $Y=2.04 $X2=0.295 $Y2=2.895
r80 1 12 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.15
+ $Y=2.04 $X2=0.295 $Y2=2.185
.ends

.subckt PM_SKY130_FD_SC_LP__AND3B_LP%X 1 2 9 11 12 13 14 15 31
r27 31 32 1.20415 $w=7.48e-07 $l=1e-08 $layer=LI1_cond $X=3.82 $Y=2.035 $X2=3.82
+ $Y2=2.025
r28 15 41 1.99346 $w=7.48e-07 $l=1.25e-07 $layer=LI1_cond $X=3.82 $Y=2.775
+ $X2=3.82 $Y2=2.9
r29 14 15 5.90065 $w=7.48e-07 $l=3.7e-07 $layer=LI1_cond $X=3.82 $Y=2.405
+ $X2=3.82 $Y2=2.775
r30 14 35 3.42876 $w=7.48e-07 $l=2.15e-07 $layer=LI1_cond $X=3.82 $Y=2.405
+ $X2=3.82 $Y2=2.19
r31 13 35 1.88183 $w=7.48e-07 $l=1.18e-07 $layer=LI1_cond $X=3.82 $Y=2.072
+ $X2=3.82 $Y2=2.19
r32 13 31 0.590065 $w=7.48e-07 $l=3.7e-08 $layer=LI1_cond $X=3.82 $Y=2.072
+ $X2=3.82 $Y2=2.035
r33 13 32 0.857566 $w=5.28e-07 $l=3.8e-08 $layer=LI1_cond $X=3.93 $Y=1.987
+ $X2=3.93 $Y2=2.025
r34 12 13 7.26674 $w=5.28e-07 $l=3.22e-07 $layer=LI1_cond $X=3.93 $Y=1.665
+ $X2=3.93 $Y2=1.987
r35 12 22 4.96485 $w=5.28e-07 $l=2.2e-07 $layer=LI1_cond $X=3.93 $Y=1.665
+ $X2=3.93 $Y2=1.445
r36 11 22 3.38513 $w=5.28e-07 $l=1.5e-07 $layer=LI1_cond $X=3.93 $Y=1.295
+ $X2=3.93 $Y2=1.445
r37 11 28 4.28868 $w=5.28e-07 $l=1.15e-07 $layer=LI1_cond $X=3.93 $Y=1.295
+ $X2=3.93 $Y2=1.18
r38 9 28 23.9219 $w=3.28e-07 $l=6.85e-07 $layer=LI1_cond $X=3.83 $Y=0.495
+ $X2=3.83 $Y2=1.18
r39 2 41 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=3.47
+ $Y=2.045 $X2=3.61 $Y2=2.9
r40 2 35 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=3.47
+ $Y=2.045 $X2=3.61 $Y2=2.19
r41 1 9 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=3.69
+ $Y=0.285 $X2=3.83 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__AND3B_LP%VGND 1 2 7 9 13 16 17 18 31 32
r42 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r43 31 32 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r44 29 32 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=4.08
+ $Y2=0
r45 28 31 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=3.12 $Y=0 $X2=4.08
+ $Y2=0
r46 28 29 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r47 26 29 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r48 25 26 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r49 23 36 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r50 22 25 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=0.72 $Y=0 $X2=2.64
+ $Y2=0
r51 22 23 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r52 20 35 4.73185 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=0 $X2=0.222
+ $Y2=0
r53 20 22 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.445 $Y=0 $X2=0.72
+ $Y2=0
r54 18 26 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r55 18 23 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=2.16 $Y=0 $X2=0.72
+ $Y2=0
r56 16 25 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=2.71 $Y=0 $X2=2.64
+ $Y2=0
r57 16 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.71 $Y=0 $X2=2.875
+ $Y2=0
r58 15 28 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=3.04 $Y=0 $X2=3.12
+ $Y2=0
r59 15 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.04 $Y=0 $X2=2.875
+ $Y2=0
r60 11 17 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.875 $Y=0.085
+ $X2=2.875 $Y2=0
r61 11 13 12.7467 $w=3.28e-07 $l=3.65e-07 $layer=LI1_cond $X=2.875 $Y=0.085
+ $X2=2.875 $Y2=0.45
r62 7 35 3.03433 $w=3.3e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.28 $Y=0.085
+ $X2=0.222 $Y2=0
r63 7 9 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=0.28 $Y=0.085 $X2=0.28
+ $Y2=0.495
r64 2 13 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=2.735
+ $Y=0.285 $X2=2.875 $Y2=0.45
r65 1 9 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.285 $X2=0.28 $Y2=0.495
.ends

