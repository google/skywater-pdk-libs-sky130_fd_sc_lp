* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__sdfbbn_1 CLK_N D RESET_B SCD SCE SET_B VGND VNB VPB VPWR
+ Q Q_N
X0 a_27_474# SCD VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X1 a_1295_379# a_995_66# a_1397_379# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X2 a_2198_379# a_995_66# a_2299_119# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X3 VGND a_1445_324# a_2198_119# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X4 a_2198_119# a_838_50# a_2299_119# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X5 a_1439_104# a_1445_324# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 VPWR CLK_N a_838_50# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X7 a_995_66# a_838_50# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X8 a_200_119# a_328_429# a_27_474# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X9 VPWR SCE a_200_474# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X10 a_200_474# D a_200_119# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X11 VGND SET_B a_1752_60# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X12 a_1752_60# a_1295_379# a_1445_324# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X13 a_995_66# a_838_50# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X14 VPWR a_2449_137# Q_N VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X15 a_2299_119# a_995_66# a_2401_163# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X16 a_1445_324# a_1926_21# a_1752_60# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X17 VGND a_3279_367# Q VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X18 a_1445_324# a_1295_379# a_1996_379# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X19 VGND SCD a_122_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X20 a_2636_119# a_2299_119# a_2449_137# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X21 a_2401_506# a_2449_137# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X22 a_1295_379# a_838_50# a_1439_104# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X23 VGND SET_B a_2636_119# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X24 a_2449_137# a_2299_119# a_2798_451# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X25 VGND CLK_N a_838_50# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X26 VPWR SET_B a_2449_137# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X27 a_2449_137# a_1926_21# a_2636_119# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X28 a_200_119# a_995_66# a_1295_379# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X29 a_3279_367# a_2449_137# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X30 a_1397_379# a_1445_324# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X31 VPWR SET_B a_1445_324# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X32 a_200_119# a_838_50# a_1295_379# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X33 a_122_119# SCE a_200_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X34 VPWR a_1445_324# a_2198_379# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X35 a_1996_379# a_1926_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X36 a_2798_451# a_1926_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X37 a_200_119# D a_314_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X38 a_2299_119# a_838_50# a_2401_506# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X39 a_314_119# a_328_429# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X40 VPWR a_3279_367# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X41 a_1926_21# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X42 a_1926_21# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X43 a_2401_163# a_2449_137# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X44 a_3279_367# a_2449_137# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X45 VPWR SCE a_328_429# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X46 VGND SCE a_328_429# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X47 VGND a_2449_137# Q_N VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
.ends
