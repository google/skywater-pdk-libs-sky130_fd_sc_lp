* File: sky130_fd_sc_lp__maj3_lp.spice
* Created: Wed Sep  2 09:59:44 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__maj3_lp.pex.spice"
.subckt sky130_fd_sc_lp__maj3_lp  VNB VPB A B C VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* C	C
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1000 A_154_125# N_B_M1000_g N_A_29_419#_M1000_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.1197 PD=0.66 PS=1.41 NRD=18.564 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.1 A=0.063 P=1.14 MULT=1
MM1010 N_VGND_M1010_d N_A_M1010_g A_154_125# VNB NSHORT L=0.15 W=0.42
+ AD=0.133725 AS=0.0504 PD=1.145 PS=0.66 NRD=75.252 NRS=18.564 M=1 R=2.8
+ SA=75000.6 SB=75001.7 A=0.063 P=1.14 MULT=1
MM1014 A_350_125# N_A_M1014_g N_VGND_M1010_d VNB NSHORT L=0.15 W=0.42 AD=0.0504
+ AS=0.133725 PD=0.66 PS=1.145 NRD=18.564 NRS=75.252 M=1 R=2.8 SA=75001.2
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1006 N_A_29_419#_M1006_d N_C_M1006_g A_350_125# VNB NSHORT L=0.15 W=0.42
+ AD=0.100537 AS=0.0504 PD=1.065 PS=0.66 NRD=24.276 NRS=18.564 M=1 R=2.8
+ SA=75001.6 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1011 A_530_68# N_B_M1011_g N_A_29_419#_M1006_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0651 AS=0.100537 PD=0.73 PS=1.065 NRD=28.56 NRS=0 M=1 R=2.8 SA=75000.8
+ SB=75001.5 A=0.063 P=1.14 MULT=1
MM1001 N_VGND_M1001_d N_C_M1001_g A_530_68# VNB NSHORT L=0.15 W=0.42 AD=0.0588
+ AS=0.0651 PD=0.7 PS=0.73 NRD=0 NRS=28.56 M=1 R=2.8 SA=75001.3 SB=75001 A=0.063
+ P=1.14 MULT=1
MM1009 A_708_68# N_A_29_419#_M1009_g N_VGND_M1001_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75001.7
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1007 N_X_M1007_d N_A_29_419#_M1007_g A_708_68# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75002.1
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1004 A_152_419# N_B_M1004_g N_A_29_419#_M1004_s VPB PHIGHVT L=0.25 W=1
+ AD=0.105 AS=0.365 PD=1.21 PS=2.73 NRD=9.8303 NRS=15.7403 M=1 R=4 SA=125000
+ SB=125003 A=0.25 P=2.5 MULT=1
MM1013 N_VPWR_M1013_d N_A_M1013_g A_152_419# VPB PHIGHVT L=0.25 W=1 AD=0.14
+ AS=0.105 PD=1.28 PS=1.21 NRD=0 NRS=9.8303 M=1 R=4 SA=125001 SB=125003 A=0.25
+ P=2.5 MULT=1
MM1012 A_350_419# N_A_M1012_g N_VPWR_M1013_d VPB PHIGHVT L=0.25 W=1 AD=0.105
+ AS=0.14 PD=1.21 PS=1.28 NRD=9.8303 NRS=0 M=1 R=4 SA=125001 SB=125002 A=0.25
+ P=2.5 MULT=1
MM1008 N_A_29_419#_M1008_d N_C_M1008_g A_350_419# VPB PHIGHVT L=0.25 W=1 AD=0.14
+ AS=0.105 PD=1.28 PS=1.21 NRD=0 NRS=9.8303 M=1 R=4 SA=125002 SB=125002 A=0.25
+ P=2.5 MULT=1
MM1002 A_548_419# N_B_M1002_g N_A_29_419#_M1008_d VPB PHIGHVT L=0.25 W=1
+ AD=0.125 AS=0.14 PD=1.25 PS=1.28 NRD=13.7703 NRS=0 M=1 R=4 SA=125002 SB=125001
+ A=0.25 P=2.5 MULT=1
MM1005 N_VPWR_M1005_d N_C_M1005_g A_548_419# VPB PHIGHVT L=0.25 W=1 AD=0.145
+ AS=0.125 PD=1.29 PS=1.25 NRD=0 NRS=13.7703 M=1 R=4 SA=125003 SB=125001 A=0.25
+ P=2.5 MULT=1
MM1003 N_X_M1003_d N_A_29_419#_M1003_g N_VPWR_M1005_d VPB PHIGHVT L=0.25 W=1
+ AD=0.285 AS=0.145 PD=2.57 PS=1.29 NRD=0 NRS=1.9503 M=1 R=4 SA=125003 SB=125000
+ A=0.25 P=2.5 MULT=1
DX15_noxref VNB VPB NWDIODE A=8.7655 P=13.13
*
.include "sky130_fd_sc_lp__maj3_lp.pxi.spice"
*
.ends
*
*
