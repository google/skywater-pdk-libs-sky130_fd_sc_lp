* File: sky130_fd_sc_lp__o21ai_lp.pxi.spice
* Created: Fri Aug 28 11:05:08 2020
* 
x_PM_SKY130_FD_SC_LP__O21AI_LP%A1 N_A1_M1000_g N_A1_M1001_g N_A1_c_47_n
+ N_A1_c_48_n A1 A1 N_A1_c_50_n PM_SKY130_FD_SC_LP__O21AI_LP%A1
x_PM_SKY130_FD_SC_LP__O21AI_LP%A2 N_A2_M1004_g N_A2_M1003_g N_A2_c_80_n
+ N_A2_c_81_n A2 A2 N_A2_c_83_n PM_SKY130_FD_SC_LP__O21AI_LP%A2
x_PM_SKY130_FD_SC_LP__O21AI_LP%B1 N_B1_M1002_g N_B1_M1005_g N_B1_c_119_n
+ N_B1_c_120_n B1 B1 N_B1_c_122_n PM_SKY130_FD_SC_LP__O21AI_LP%B1
x_PM_SKY130_FD_SC_LP__O21AI_LP%VPWR N_VPWR_M1000_s N_VPWR_M1002_d N_VPWR_c_155_n
+ N_VPWR_c_156_n N_VPWR_c_157_n N_VPWR_c_158_n VPWR N_VPWR_c_159_n
+ N_VPWR_c_154_n PM_SKY130_FD_SC_LP__O21AI_LP%VPWR
x_PM_SKY130_FD_SC_LP__O21AI_LP%Y N_Y_M1005_d N_Y_M1004_d N_Y_c_181_n N_Y_c_179_n
+ N_Y_c_180_n Y Y PM_SKY130_FD_SC_LP__O21AI_LP%Y
x_PM_SKY130_FD_SC_LP__O21AI_LP%A_64_57# N_A_64_57#_M1001_s N_A_64_57#_M1003_d
+ N_A_64_57#_c_210_n N_A_64_57#_c_211_n N_A_64_57#_c_212_n N_A_64_57#_c_213_n
+ PM_SKY130_FD_SC_LP__O21AI_LP%A_64_57#
x_PM_SKY130_FD_SC_LP__O21AI_LP%VGND N_VGND_M1001_d N_VGND_c_242_n N_VGND_c_243_n
+ N_VGND_c_244_n VGND N_VGND_c_245_n N_VGND_c_246_n
+ PM_SKY130_FD_SC_LP__O21AI_LP%VGND
cc_1 VNB N_A1_M1001_g 0.0456132f $X=-0.19 $Y=-0.245 $X2=0.68 $Y2=0.495
cc_2 VNB N_A1_c_47_n 0.025421f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.63
cc_3 VNB N_A1_c_48_n 0.00188025f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.795
cc_4 VNB A1 0.0367954f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_5 VNB N_A1_c_50_n 0.01709f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.29
cc_6 VNB N_A2_M1003_g 0.0343212f $X=-0.19 $Y=-0.245 $X2=0.68 $Y2=0.495
cc_7 VNB N_A2_c_80_n 0.0238826f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.63
cc_8 VNB N_A2_c_81_n 0.00176646f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.795
cc_9 VNB A2 0.00171359f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_10 VNB N_A2_c_83_n 0.0167493f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_B1_M1005_g 0.037026f $X=-0.19 $Y=-0.245 $X2=0.68 $Y2=0.495
cc_12 VNB N_B1_c_119_n 0.023974f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.63
cc_13 VNB N_B1_c_120_n 0.00177322f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.795
cc_14 VNB B1 0.00750659f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_15 VNB N_B1_c_122_n 0.0168121f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_VPWR_c_154_n 0.103974f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_Y_c_179_n 0.0454093f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.125
cc_18 VNB N_Y_c_180_n 0.0319758f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_64_57#_c_210_n 0.0219254f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.29
cc_20 VNB N_A_64_57#_c_211_n 0.0226191f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.63
cc_21 VNB N_A_64_57#_c_212_n 0.0100927f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.795
cc_22 VNB N_A_64_57#_c_213_n 0.00207453f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_23 VNB N_VGND_c_242_n 0.00712794f $X=-0.19 $Y=-0.245 $X2=0.68 $Y2=0.495
cc_24 VNB N_VGND_c_243_n 0.0248931f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.29
cc_25 VNB N_VGND_c_244_n 0.00632158f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.125
cc_26 VNB N_VGND_c_245_n 0.0352041f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.29
cc_27 VNB N_VGND_c_246_n 0.169132f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.29
cc_28 VPB N_A1_M1000_g 0.0402348f $X=-0.19 $Y=1.655 $X2=0.65 $Y2=2.545
cc_29 VPB N_A1_c_48_n 0.0126461f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=1.795
cc_30 VPB A1 0.015971f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_31 VPB N_A2_M1004_g 0.0316723f $X=-0.19 $Y=1.655 $X2=0.65 $Y2=2.545
cc_32 VPB N_A2_c_81_n 0.012129f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=1.795
cc_33 VPB A2 7.54819e-19 $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_34 VPB N_B1_M1002_g 0.0354587f $X=-0.19 $Y=1.655 $X2=0.65 $Y2=2.545
cc_35 VPB N_B1_c_120_n 0.012185f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=1.795
cc_36 VPB B1 0.00184675f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_37 VPB N_VPWR_c_155_n 0.0147062f $X=-0.19 $Y=1.655 $X2=0.68 $Y2=0.495
cc_38 VPB N_VPWR_c_156_n 0.0470528f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=1.29
cc_39 VPB N_VPWR_c_157_n 0.0159821f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_40 VPB N_VPWR_c_158_n 0.0328593f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_41 VPB N_VPWR_c_159_n 0.0345234f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_42 VPB N_VPWR_c_154_n 0.0677165f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_43 VPB N_Y_c_181_n 0.020173f $X=-0.19 $Y=1.655 $X2=0.68 $Y2=0.495
cc_44 VPB N_Y_c_179_n 0.0156431f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=1.125
cc_45 VPB Y 0.011981f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_46 N_A1_M1000_g N_A2_M1004_g 0.0279407f $X=0.65 $Y=2.545 $X2=0 $Y2=0
cc_47 N_A1_M1001_g N_A2_M1003_g 0.0232293f $X=0.68 $Y=0.495 $X2=0 $Y2=0
cc_48 N_A1_c_47_n N_A2_c_80_n 0.0279407f $X=0.61 $Y=1.63 $X2=0 $Y2=0
cc_49 N_A1_c_48_n N_A2_c_81_n 0.0279407f $X=0.61 $Y=1.795 $X2=0 $Y2=0
cc_50 A1 A2 0.0540841f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_51 N_A1_c_50_n A2 7.5249e-19 $X=0.61 $Y=1.29 $X2=0 $Y2=0
cc_52 A1 N_A2_c_83_n 0.00437388f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_53 N_A1_c_50_n N_A2_c_83_n 0.0279407f $X=0.61 $Y=1.29 $X2=0 $Y2=0
cc_54 N_A1_M1000_g N_VPWR_c_156_n 0.0268199f $X=0.65 $Y=2.545 $X2=0 $Y2=0
cc_55 N_A1_c_48_n N_VPWR_c_156_n 0.00207134f $X=0.61 $Y=1.795 $X2=0 $Y2=0
cc_56 A1 N_VPWR_c_156_n 0.0241167f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_57 N_A1_M1000_g N_VPWR_c_159_n 0.00802402f $X=0.65 $Y=2.545 $X2=0 $Y2=0
cc_58 N_A1_M1000_g N_VPWR_c_154_n 0.0142664f $X=0.65 $Y=2.545 $X2=0 $Y2=0
cc_59 N_A1_M1000_g Y 0.00422969f $X=0.65 $Y=2.545 $X2=0 $Y2=0
cc_60 N_A1_M1001_g N_A_64_57#_c_210_n 0.00979067f $X=0.68 $Y=0.495 $X2=0 $Y2=0
cc_61 N_A1_M1001_g N_A_64_57#_c_211_n 0.00915924f $X=0.68 $Y=0.495 $X2=0 $Y2=0
cc_62 A1 N_A_64_57#_c_211_n 0.0153682f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_63 N_A1_c_50_n N_A_64_57#_c_211_n 5.23484e-19 $X=0.61 $Y=1.29 $X2=0 $Y2=0
cc_64 N_A1_M1001_g N_A_64_57#_c_212_n 0.00419316f $X=0.68 $Y=0.495 $X2=0 $Y2=0
cc_65 A1 N_A_64_57#_c_212_n 0.0285664f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_66 N_A1_c_50_n N_A_64_57#_c_212_n 0.00429552f $X=0.61 $Y=1.29 $X2=0 $Y2=0
cc_67 N_A1_M1001_g N_A_64_57#_c_213_n 8.76764e-19 $X=0.68 $Y=0.495 $X2=0 $Y2=0
cc_68 N_A1_M1001_g N_VGND_c_242_n 0.00479877f $X=0.68 $Y=0.495 $X2=0 $Y2=0
cc_69 N_A1_M1001_g N_VGND_c_243_n 0.00502664f $X=0.68 $Y=0.495 $X2=0 $Y2=0
cc_70 N_A1_M1001_g N_VGND_c_246_n 0.00652763f $X=0.68 $Y=0.495 $X2=0 $Y2=0
cc_71 N_A2_M1004_g N_B1_M1002_g 0.0169128f $X=1.14 $Y=2.545 $X2=0 $Y2=0
cc_72 N_A2_M1003_g N_B1_M1005_g 0.0276106f $X=1.27 $Y=0.495 $X2=0 $Y2=0
cc_73 N_A2_c_80_n N_B1_c_119_n 0.01184f $X=1.18 $Y=1.63 $X2=0 $Y2=0
cc_74 N_A2_c_81_n N_B1_c_120_n 0.01184f $X=1.18 $Y=1.795 $X2=0 $Y2=0
cc_75 A2 B1 0.0438819f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_76 N_A2_c_83_n B1 0.00410205f $X=1.18 $Y=1.29 $X2=0 $Y2=0
cc_77 A2 N_B1_c_122_n 8.23261e-19 $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_78 N_A2_c_83_n N_B1_c_122_n 0.01184f $X=1.18 $Y=1.29 $X2=0 $Y2=0
cc_79 N_A2_M1004_g N_VPWR_c_156_n 0.00414308f $X=1.14 $Y=2.545 $X2=0 $Y2=0
cc_80 N_A2_M1004_g N_VPWR_c_158_n 8.46069e-19 $X=1.14 $Y=2.545 $X2=0 $Y2=0
cc_81 N_A2_M1004_g N_VPWR_c_159_n 0.00673673f $X=1.14 $Y=2.545 $X2=0 $Y2=0
cc_82 N_A2_M1004_g N_VPWR_c_154_n 0.0102002f $X=1.14 $Y=2.545 $X2=0 $Y2=0
cc_83 N_A2_M1004_g Y 0.0363457f $X=1.14 $Y=2.545 $X2=0 $Y2=0
cc_84 N_A2_c_81_n Y 6.13398e-19 $X=1.18 $Y=1.795 $X2=0 $Y2=0
cc_85 A2 Y 0.0141565f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_86 N_A2_M1003_g N_A_64_57#_c_210_n 8.76764e-19 $X=1.27 $Y=0.495 $X2=0 $Y2=0
cc_87 N_A2_M1003_g N_A_64_57#_c_211_n 0.0118802f $X=1.27 $Y=0.495 $X2=0 $Y2=0
cc_88 A2 N_A_64_57#_c_211_n 0.0246663f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_89 N_A2_c_83_n N_A_64_57#_c_211_n 0.00122995f $X=1.18 $Y=1.29 $X2=0 $Y2=0
cc_90 N_A2_M1003_g N_A_64_57#_c_213_n 0.00876498f $X=1.27 $Y=0.495 $X2=0 $Y2=0
cc_91 N_A2_M1003_g N_VGND_c_242_n 0.00479877f $X=1.27 $Y=0.495 $X2=0 $Y2=0
cc_92 N_A2_M1003_g N_VGND_c_245_n 0.00502664f $X=1.27 $Y=0.495 $X2=0 $Y2=0
cc_93 N_A2_M1003_g N_VGND_c_246_n 0.00579934f $X=1.27 $Y=0.495 $X2=0 $Y2=0
cc_94 N_B1_M1002_g N_VPWR_c_158_n 0.0167591f $X=1.71 $Y=2.545 $X2=0 $Y2=0
cc_95 N_B1_M1002_g N_VPWR_c_159_n 0.00802402f $X=1.71 $Y=2.545 $X2=0 $Y2=0
cc_96 N_B1_M1002_g N_VPWR_c_154_n 0.0144019f $X=1.71 $Y=2.545 $X2=0 $Y2=0
cc_97 N_B1_M1002_g N_Y_c_181_n 0.0223083f $X=1.71 $Y=2.545 $X2=0 $Y2=0
cc_98 N_B1_c_120_n N_Y_c_181_n 5.43485e-19 $X=1.75 $Y=1.795 $X2=0 $Y2=0
cc_99 B1 N_Y_c_181_n 0.0253793f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_100 N_B1_M1002_g N_Y_c_179_n 0.00590404f $X=1.71 $Y=2.545 $X2=0 $Y2=0
cc_101 N_B1_M1005_g N_Y_c_179_n 0.00926209f $X=1.7 $Y=0.495 $X2=0 $Y2=0
cc_102 B1 N_Y_c_179_n 0.0483772f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_103 N_B1_c_122_n N_Y_c_179_n 0.0148853f $X=1.75 $Y=1.29 $X2=0 $Y2=0
cc_104 N_B1_M1005_g N_Y_c_180_n 0.00891322f $X=1.7 $Y=0.495 $X2=0 $Y2=0
cc_105 B1 N_Y_c_180_n 0.00380507f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_106 N_B1_c_122_n N_Y_c_180_n 5.52087e-19 $X=1.75 $Y=1.29 $X2=0 $Y2=0
cc_107 N_B1_M1002_g Y 2.07053e-19 $X=1.71 $Y=2.545 $X2=0 $Y2=0
cc_108 N_B1_M1005_g N_A_64_57#_c_211_n 0.00535193f $X=1.7 $Y=0.495 $X2=0 $Y2=0
cc_109 B1 N_A_64_57#_c_211_n 0.00713614f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_110 N_B1_c_122_n N_A_64_57#_c_211_n 3.08957e-19 $X=1.75 $Y=1.29 $X2=0 $Y2=0
cc_111 N_B1_M1005_g N_A_64_57#_c_213_n 0.00743855f $X=1.7 $Y=0.495 $X2=0 $Y2=0
cc_112 N_B1_M1005_g N_VGND_c_245_n 0.00502664f $X=1.7 $Y=0.495 $X2=0 $Y2=0
cc_113 N_B1_M1005_g N_VGND_c_246_n 0.0103089f $X=1.7 $Y=0.495 $X2=0 $Y2=0
cc_114 N_VPWR_M1002_d N_Y_c_181_n 0.00305415f $X=1.835 $Y=2.045 $X2=0 $Y2=0
cc_115 N_VPWR_c_158_n N_Y_c_181_n 0.0213634f $X=1.975 $Y=2.49 $X2=0 $Y2=0
cc_116 N_VPWR_c_156_n Y 0.0181604f $X=0.385 $Y=2.19 $X2=0 $Y2=0
cc_117 N_VPWR_c_158_n Y 0.0217731f $X=1.975 $Y=2.49 $X2=0 $Y2=0
cc_118 N_VPWR_c_159_n Y 0.026783f $X=1.81 $Y=3.33 $X2=0 $Y2=0
cc_119 N_VPWR_c_154_n Y 0.0172601f $X=2.16 $Y=3.33 $X2=0 $Y2=0
cc_120 N_Y_c_179_n N_A_64_57#_c_211_n 0.00656559f $X=2.18 $Y=1.975 $X2=0 $Y2=0
cc_121 N_Y_c_179_n N_A_64_57#_c_213_n 0.00180948f $X=2.18 $Y=1.975 $X2=0 $Y2=0
cc_122 N_Y_c_180_n N_A_64_57#_c_213_n 0.0179956f $X=2.18 $Y=0.495 $X2=0 $Y2=0
cc_123 N_Y_c_180_n N_VGND_c_245_n 0.0283101f $X=2.18 $Y=0.495 $X2=0 $Y2=0
cc_124 N_Y_c_180_n N_VGND_c_246_n 0.0166475f $X=2.18 $Y=0.495 $X2=0 $Y2=0
cc_125 N_A_64_57#_c_210_n N_VGND_c_242_n 0.0125869f $X=0.465 $Y=0.495 $X2=0
+ $Y2=0
cc_126 N_A_64_57#_c_211_n N_VGND_c_242_n 0.025061f $X=1.32 $Y=0.86 $X2=0 $Y2=0
cc_127 N_A_64_57#_c_213_n N_VGND_c_242_n 0.0125869f $X=1.485 $Y=0.495 $X2=0
+ $Y2=0
cc_128 N_A_64_57#_c_210_n N_VGND_c_243_n 0.0220321f $X=0.465 $Y=0.495 $X2=0
+ $Y2=0
cc_129 N_A_64_57#_c_213_n N_VGND_c_245_n 0.021949f $X=1.485 $Y=0.495 $X2=0 $Y2=0
cc_130 N_A_64_57#_c_210_n N_VGND_c_246_n 0.0125808f $X=0.465 $Y=0.495 $X2=0
+ $Y2=0
cc_131 N_A_64_57#_c_211_n N_VGND_c_246_n 0.0125928f $X=1.32 $Y=0.86 $X2=0 $Y2=0
cc_132 N_A_64_57#_c_213_n N_VGND_c_246_n 0.0124703f $X=1.485 $Y=0.495 $X2=0
+ $Y2=0
