* File: sky130_fd_sc_lp__nor4_4.pex.spice
* Created: Fri Aug 28 10:57:42 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__NOR4_4%A 3 5 7 10 12 14 17 19 21 24 26 28 29 30 31
+ 32 37 53 55
c78 55 0 1.15464e-19 $X=2.06 $Y=1.405
c79 24 0 1.83481e-20 $X=1.99 $Y=2.465
r80 54 55 8.8479 $w=4.4e-07 $l=7e-08 $layer=POLY_cond $X=1.99 $Y=1.405 $X2=2.06
+ $Y2=1.405
r81 52 54 2.52797 $w=4.4e-07 $l=2e-08 $layer=POLY_cond $X=1.97 $Y=1.405 $X2=1.99
+ $Y2=1.405
r82 52 53 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.97
+ $Y=1.46 $X2=1.97 $Y2=1.46
r83 50 52 42.9755 $w=4.4e-07 $l=3.4e-07 $layer=POLY_cond $X=1.63 $Y=1.405
+ $X2=1.97 $Y2=1.405
r84 49 50 8.8479 $w=4.4e-07 $l=7e-08 $layer=POLY_cond $X=1.56 $Y=1.405 $X2=1.63
+ $Y2=1.405
r85 48 49 45.5035 $w=4.4e-07 $l=3.6e-07 $layer=POLY_cond $X=1.2 $Y=1.405
+ $X2=1.56 $Y2=1.405
r86 47 48 8.8479 $w=4.4e-07 $l=7e-08 $layer=POLY_cond $X=1.13 $Y=1.405 $X2=1.2
+ $Y2=1.405
r87 45 47 22.7517 $w=4.4e-07 $l=1.8e-07 $layer=POLY_cond $X=0.95 $Y=1.405
+ $X2=1.13 $Y2=1.405
r88 45 46 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.95
+ $Y=1.46 $X2=0.95 $Y2=1.46
r89 43 45 22.7517 $w=4.4e-07 $l=1.8e-07 $layer=POLY_cond $X=0.77 $Y=1.405
+ $X2=0.95 $Y2=1.405
r90 42 43 8.8479 $w=4.4e-07 $l=7e-08 $layer=POLY_cond $X=0.7 $Y=1.405 $X2=0.77
+ $Y2=1.405
r91 39 40 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.61
+ $Y=1.46 $X2=0.61 $Y2=1.46
r92 37 42 9.4799 $w=4.4e-07 $l=7.5e-08 $layer=POLY_cond $X=0.625 $Y=1.405
+ $X2=0.7 $Y2=1.405
r93 37 39 1.89598 $w=4.4e-07 $l=1.5e-08 $layer=POLY_cond $X=0.625 $Y=1.405
+ $X2=0.61 $Y2=1.405
r94 32 53 8.25206 $w=4.03e-07 $l=2.9e-07 $layer=LI1_cond $X=1.68 $Y=1.547
+ $X2=1.97 $Y2=1.547
r95 31 32 13.6586 $w=4.03e-07 $l=4.8e-07 $layer=LI1_cond $X=1.2 $Y=1.547
+ $X2=1.68 $Y2=1.547
r96 31 46 7.11385 $w=4.03e-07 $l=2.5e-07 $layer=LI1_cond $X=1.2 $Y=1.547
+ $X2=0.95 $Y2=1.547
r97 30 46 6.54474 $w=4.03e-07 $l=2.3e-07 $layer=LI1_cond $X=0.72 $Y=1.547
+ $X2=0.95 $Y2=1.547
r98 30 40 3.13009 $w=4.03e-07 $l=1.1e-07 $layer=LI1_cond $X=0.72 $Y=1.547
+ $X2=0.61 $Y2=1.547
r99 29 40 10.5285 $w=4.03e-07 $l=3.7e-07 $layer=LI1_cond $X=0.24 $Y=1.547
+ $X2=0.61 $Y2=1.547
r100 26 55 28.2085 $w=1.5e-07 $l=2.2e-07 $layer=POLY_cond $X=2.06 $Y=1.185
+ $X2=2.06 $Y2=1.405
r101 26 28 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.06 $Y=1.185
+ $X2=2.06 $Y2=0.655
r102 22 54 28.2085 $w=1.5e-07 $l=2.2e-07 $layer=POLY_cond $X=1.99 $Y=1.625
+ $X2=1.99 $Y2=1.405
r103 22 24 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=1.99 $Y=1.625
+ $X2=1.99 $Y2=2.465
r104 19 50 28.2085 $w=1.5e-07 $l=2.2e-07 $layer=POLY_cond $X=1.63 $Y=1.185
+ $X2=1.63 $Y2=1.405
r105 19 21 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.63 $Y=1.185
+ $X2=1.63 $Y2=0.655
r106 15 49 28.2085 $w=1.5e-07 $l=2.2e-07 $layer=POLY_cond $X=1.56 $Y=1.625
+ $X2=1.56 $Y2=1.405
r107 15 17 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=1.56 $Y=1.625
+ $X2=1.56 $Y2=2.465
r108 12 48 28.2085 $w=1.5e-07 $l=2.2e-07 $layer=POLY_cond $X=1.2 $Y=1.185
+ $X2=1.2 $Y2=1.405
r109 12 14 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.2 $Y=1.185
+ $X2=1.2 $Y2=0.655
r110 8 47 28.2085 $w=1.5e-07 $l=2.2e-07 $layer=POLY_cond $X=1.13 $Y=1.625
+ $X2=1.13 $Y2=1.405
r111 8 10 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=1.13 $Y=1.625
+ $X2=1.13 $Y2=2.465
r112 5 43 28.2085 $w=1.5e-07 $l=2.2e-07 $layer=POLY_cond $X=0.77 $Y=1.185
+ $X2=0.77 $Y2=1.405
r113 5 7 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.77 $Y=1.185
+ $X2=0.77 $Y2=0.655
r114 1 42 28.2085 $w=1.5e-07 $l=2.2e-07 $layer=POLY_cond $X=0.7 $Y=1.625 $X2=0.7
+ $Y2=1.405
r115 1 3 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=0.7 $Y=1.625 $X2=0.7
+ $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4_4%B 1 3 4 6 7 9 10 12 13 15 16 18 19 21 22 24
+ 25 26 40 41
r83 40 42 1.94355 $w=4.96e-07 $l=2e-08 $layer=POLY_cond $X=4.21 $Y=1.455
+ $X2=4.23 $Y2=1.455
r84 40 41 48.4267 $w=1.7e-07 $l=5.1e-07 $layer=licon1_POLY $count=3 $X=4.21
+ $Y=1.35 $X2=4.21 $Y2=1.35
r85 38 40 39.8427 $w=4.96e-07 $l=4.1e-07 $layer=POLY_cond $X=3.8 $Y=1.455
+ $X2=4.21 $Y2=1.455
r86 37 38 8.74597 $w=4.96e-07 $l=9e-08 $layer=POLY_cond $X=3.71 $Y=1.455 $X2=3.8
+ $Y2=1.455
r87 36 37 33.0403 $w=4.96e-07 $l=3.4e-07 $layer=POLY_cond $X=3.37 $Y=1.455
+ $X2=3.71 $Y2=1.455
r88 35 36 8.74597 $w=4.96e-07 $l=9e-08 $layer=POLY_cond $X=3.28 $Y=1.455
+ $X2=3.37 $Y2=1.455
r89 34 35 33.0403 $w=4.96e-07 $l=3.4e-07 $layer=POLY_cond $X=2.94 $Y=1.455
+ $X2=3.28 $Y2=1.455
r90 33 34 8.74597 $w=4.96e-07 $l=9e-08 $layer=POLY_cond $X=2.85 $Y=1.455
+ $X2=2.94 $Y2=1.455
r91 31 33 33.0403 $w=4.96e-07 $l=3.4e-07 $layer=POLY_cond $X=2.51 $Y=1.455
+ $X2=2.85 $Y2=1.455
r92 31 32 48.4267 $w=1.7e-07 $l=5.1e-07 $layer=licon1_POLY $count=3 $X=2.51
+ $Y=1.35 $X2=2.51 $Y2=1.35
r93 29 31 8.74597 $w=4.96e-07 $l=9e-08 $layer=POLY_cond $X=2.42 $Y=1.455
+ $X2=2.51 $Y2=1.455
r94 26 41 38.6512 $w=3.23e-07 $l=1.09e-06 $layer=LI1_cond $X=3.12 $Y=1.372
+ $X2=4.21 $Y2=1.372
r95 25 26 17.0207 $w=3.23e-07 $l=4.8e-07 $layer=LI1_cond $X=2.64 $Y=1.372
+ $X2=3.12 $Y2=1.372
r96 25 32 4.60977 $w=3.23e-07 $l=1.3e-07 $layer=LI1_cond $X=2.64 $Y=1.372
+ $X2=2.51 $Y2=1.372
r97 22 42 31.2052 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=4.23 $Y=1.185
+ $X2=4.23 $Y2=1.455
r98 22 24 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=4.23 $Y=1.185
+ $X2=4.23 $Y2=0.655
r99 19 38 31.2052 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=3.8 $Y=1.185 $X2=3.8
+ $Y2=1.455
r100 19 21 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=3.8 $Y=1.185
+ $X2=3.8 $Y2=0.655
r101 16 37 31.2052 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=3.71 $Y=1.725
+ $X2=3.71 $Y2=1.455
r102 16 18 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=3.71 $Y=1.725
+ $X2=3.71 $Y2=2.465
r103 13 36 31.2052 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=3.37 $Y=1.185
+ $X2=3.37 $Y2=1.455
r104 13 15 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=3.37 $Y=1.185
+ $X2=3.37 $Y2=0.655
r105 10 35 31.2052 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=3.28 $Y=1.725
+ $X2=3.28 $Y2=1.455
r106 10 12 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=3.28 $Y=1.725
+ $X2=3.28 $Y2=2.465
r107 7 34 31.2052 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=2.94 $Y=1.185
+ $X2=2.94 $Y2=1.455
r108 7 9 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.94 $Y=1.185
+ $X2=2.94 $Y2=0.655
r109 4 33 31.2052 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=2.85 $Y=1.725
+ $X2=2.85 $Y2=1.455
r110 4 6 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=2.85 $Y=1.725
+ $X2=2.85 $Y2=2.465
r111 1 29 31.2052 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=2.42 $Y=1.725
+ $X2=2.42 $Y2=1.455
r112 1 3 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=2.42 $Y=1.725
+ $X2=2.42 $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4_4%C 1 3 6 8 10 13 15 17 20 22 24 27 29 30 31 45
r89 43 45 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=5.86 $Y=1.35 $X2=5.95
+ $Y2=1.35
r90 43 44 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.86
+ $Y=1.35 $X2=5.86 $Y2=1.35
r91 41 43 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=5.52 $Y=1.35
+ $X2=5.86 $Y2=1.35
r92 40 41 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=5.09 $Y=1.35
+ $X2=5.52 $Y2=1.35
r93 38 40 43.7153 $w=3.3e-07 $l=2.5e-07 $layer=POLY_cond $X=4.84 $Y=1.35
+ $X2=5.09 $Y2=1.35
r94 38 39 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.84
+ $Y=1.35 $X2=4.84 $Y2=1.35
r95 35 38 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=4.66 $Y=1.35 $X2=4.84
+ $Y2=1.35
r96 31 44 4.96437 $w=3.23e-07 $l=1.4e-07 $layer=LI1_cond $X=6 $Y=1.372 $X2=5.86
+ $Y2=1.372
r97 30 44 12.0563 $w=3.23e-07 $l=3.4e-07 $layer=LI1_cond $X=5.52 $Y=1.372
+ $X2=5.86 $Y2=1.372
r98 29 30 17.0207 $w=3.23e-07 $l=4.8e-07 $layer=LI1_cond $X=5.04 $Y=1.372
+ $X2=5.52 $Y2=1.372
r99 29 39 7.09196 $w=3.23e-07 $l=2e-07 $layer=LI1_cond $X=5.04 $Y=1.372 $X2=4.84
+ $Y2=1.372
r100 25 45 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.95 $Y=1.515
+ $X2=5.95 $Y2=1.35
r101 25 27 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=5.95 $Y=1.515
+ $X2=5.95 $Y2=2.465
r102 22 45 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.95 $Y=1.185
+ $X2=5.95 $Y2=1.35
r103 22 24 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=5.95 $Y=1.185
+ $X2=5.95 $Y2=0.655
r104 18 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.52 $Y=1.515
+ $X2=5.52 $Y2=1.35
r105 18 20 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=5.52 $Y=1.515
+ $X2=5.52 $Y2=2.465
r106 15 41 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.52 $Y=1.185
+ $X2=5.52 $Y2=1.35
r107 15 17 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=5.52 $Y=1.185
+ $X2=5.52 $Y2=0.655
r108 11 40 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.09 $Y=1.515
+ $X2=5.09 $Y2=1.35
r109 11 13 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=5.09 $Y=1.515
+ $X2=5.09 $Y2=2.465
r110 8 40 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.09 $Y=1.185
+ $X2=5.09 $Y2=1.35
r111 8 10 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=5.09 $Y=1.185
+ $X2=5.09 $Y2=0.655
r112 4 35 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.66 $Y=1.515
+ $X2=4.66 $Y2=1.35
r113 4 6 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=4.66 $Y=1.515
+ $X2=4.66 $Y2=2.465
r114 1 35 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.66 $Y=1.185
+ $X2=4.66 $Y2=1.35
r115 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=4.66 $Y=1.185
+ $X2=4.66 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4_4%D 3 7 11 15 19 23 27 31 35 38 39 50 52 59 61
r88 52 59 1.02439 $w=3.13e-07 $l=2.8e-08 $layer=LI1_cond $X=6.988 $Y=1.367
+ $X2=6.96 $Y2=1.367
r89 46 48 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=6.81 $Y=1.44
+ $X2=7.24 $Y2=1.44
r90 46 47 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.81
+ $Y=1.44 $X2=6.81 $Y2=1.44
r91 43 46 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=6.38 $Y=1.44
+ $X2=6.81 $Y2=1.44
r92 39 61 7.14549 $w=3.13e-07 $l=1.29e-07 $layer=LI1_cond $X=7.016 $Y=1.367
+ $X2=7.145 $Y2=1.367
r93 39 52 1.02439 $w=3.13e-07 $l=2.8e-08 $layer=LI1_cond $X=7.016 $Y=1.367
+ $X2=6.988 $Y2=1.367
r94 39 59 1.06098 $w=3.13e-07 $l=2.9e-08 $layer=LI1_cond $X=6.931 $Y=1.367
+ $X2=6.96 $Y2=1.367
r95 39 47 4.42684 $w=3.13e-07 $l=1.21e-07 $layer=LI1_cond $X=6.931 $Y=1.367
+ $X2=6.81 $Y2=1.367
r96 38 47 12.0732 $w=3.13e-07 $l=3.3e-07 $layer=LI1_cond $X=6.48 $Y=1.367
+ $X2=6.81 $Y2=1.367
r97 36 50 31.475 $w=3.3e-07 $l=1.8e-07 $layer=POLY_cond $X=7.49 $Y=1.44 $X2=7.67
+ $Y2=1.44
r98 36 48 43.7153 $w=3.3e-07 $l=2.5e-07 $layer=POLY_cond $X=7.49 $Y=1.44
+ $X2=7.24 $Y2=1.44
r99 35 61 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=7.49 $Y=1.44
+ $X2=7.145 $Y2=1.44
r100 35 36 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.49
+ $Y=1.44 $X2=7.49 $Y2=1.44
r101 29 50 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.67 $Y=1.605
+ $X2=7.67 $Y2=1.44
r102 29 31 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=7.67 $Y=1.605
+ $X2=7.67 $Y2=2.465
r103 25 50 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.67 $Y=1.275
+ $X2=7.67 $Y2=1.44
r104 25 27 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=7.67 $Y=1.275
+ $X2=7.67 $Y2=0.655
r105 21 48 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.24 $Y=1.605
+ $X2=7.24 $Y2=1.44
r106 21 23 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=7.24 $Y=1.605
+ $X2=7.24 $Y2=2.465
r107 17 48 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.24 $Y=1.275
+ $X2=7.24 $Y2=1.44
r108 17 19 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=7.24 $Y=1.275
+ $X2=7.24 $Y2=0.655
r109 13 46 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.81 $Y=1.605
+ $X2=6.81 $Y2=1.44
r110 13 15 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=6.81 $Y=1.605
+ $X2=6.81 $Y2=2.465
r111 9 46 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.81 $Y=1.275
+ $X2=6.81 $Y2=1.44
r112 9 11 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=6.81 $Y=1.275
+ $X2=6.81 $Y2=0.655
r113 5 43 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.38 $Y=1.605
+ $X2=6.38 $Y2=1.44
r114 5 7 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=6.38 $Y=1.605
+ $X2=6.38 $Y2=2.465
r115 1 43 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.38 $Y=1.275
+ $X2=6.38 $Y2=1.44
r116 1 3 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=6.38 $Y=1.275
+ $X2=6.38 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4_4%A_72_367# 1 2 3 4 5 16 18 20 24 26 28 29 30
+ 34 36 38 40 45 51
c63 28 0 1.15464e-19 $X=2.227 $Y=2.09
r64 38 53 2.71076 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=3.937 $Y=2.895
+ $X2=3.937 $Y2=2.98
r65 38 40 25.5049 $w=3.03e-07 $l=6.75e-07 $layer=LI1_cond $X=3.937 $Y=2.895
+ $X2=3.937 $Y2=2.22
r66 37 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.23 $Y=2.98
+ $X2=3.065 $Y2=2.98
r67 36 53 4.84748 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=3.785 $Y=2.98
+ $X2=3.937 $Y2=2.98
r68 36 37 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=3.785 $Y=2.98
+ $X2=3.23 $Y2=2.98
r69 32 51 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.065 $Y=2.895
+ $X2=3.065 $Y2=2.98
r70 32 34 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=3.065 $Y=2.895
+ $X2=3.065 $Y2=2.22
r71 31 49 4.0965 $w=1.7e-07 $l=1.18e-07 $layer=LI1_cond $X=2.345 $Y=2.98
+ $X2=2.227 $Y2=2.98
r72 30 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.9 $Y=2.98
+ $X2=3.065 $Y2=2.98
r73 30 31 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=2.9 $Y=2.98
+ $X2=2.345 $Y2=2.98
r74 29 49 2.95087 $w=2.35e-07 $l=8.5e-08 $layer=LI1_cond $X=2.227 $Y=2.895
+ $X2=2.227 $Y2=2.98
r75 28 47 2.96548 $w=2.35e-07 $l=8.5e-08 $layer=LI1_cond $X=2.227 $Y=2.09
+ $X2=2.227 $Y2=2.005
r76 28 29 39.4773 $w=2.33e-07 $l=8.05e-07 $layer=LI1_cond $X=2.227 $Y=2.09
+ $X2=2.227 $Y2=2.895
r77 27 45 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.44 $Y=2.005
+ $X2=1.345 $Y2=2.005
r78 26 47 4.08189 $w=1.7e-07 $l=1.17e-07 $layer=LI1_cond $X=2.11 $Y=2.005
+ $X2=2.227 $Y2=2.005
r79 26 27 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.11 $Y=2.005
+ $X2=1.44 $Y2=2.005
r80 22 45 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.345 $Y=2.09
+ $X2=1.345 $Y2=2.005
r81 22 24 47.2823 $w=1.88e-07 $l=8.1e-07 $layer=LI1_cond $X=1.345 $Y=2.09
+ $X2=1.345 $Y2=2.9
r82 21 43 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.58 $Y=2.005
+ $X2=0.45 $Y2=2.005
r83 20 45 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.25 $Y=2.005
+ $X2=1.345 $Y2=2.005
r84 20 21 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.25 $Y=2.005
+ $X2=0.58 $Y2=2.005
r85 16 43 2.85134 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=0.45 $Y=2.09 $X2=0.45
+ $Y2=2.005
r86 16 18 35.903 $w=2.58e-07 $l=8.1e-07 $layer=LI1_cond $X=0.45 $Y=2.09 $X2=0.45
+ $Y2=2.9
r87 5 53 400 $w=1.7e-07 $l=1.13284e-06 $layer=licon1_PDIFF $count=1 $X=3.785
+ $Y=1.835 $X2=3.925 $Y2=2.9
r88 5 40 400 $w=1.7e-07 $l=4.49583e-07 $layer=licon1_PDIFF $count=1 $X=3.785
+ $Y=1.835 $X2=3.925 $Y2=2.22
r89 4 51 400 $w=1.7e-07 $l=1.13284e-06 $layer=licon1_PDIFF $count=1 $X=2.925
+ $Y=1.835 $X2=3.065 $Y2=2.9
r90 4 34 400 $w=1.7e-07 $l=4.49583e-07 $layer=licon1_PDIFF $count=1 $X=2.925
+ $Y=1.835 $X2=3.065 $Y2=2.22
r91 3 49 400 $w=1.7e-07 $l=1.13284e-06 $layer=licon1_PDIFF $count=1 $X=2.065
+ $Y=1.835 $X2=2.205 $Y2=2.9
r92 3 47 400 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_PDIFF $count=1 $X=2.065
+ $Y=1.835 $X2=2.205 $Y2=2.085
r93 2 45 400 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_PDIFF $count=1 $X=1.205
+ $Y=1.835 $X2=1.345 $Y2=2.085
r94 2 24 400 $w=1.7e-07 $l=1.13284e-06 $layer=licon1_PDIFF $count=1 $X=1.205
+ $Y=1.835 $X2=1.345 $Y2=2.9
r95 1 43 400 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_PDIFF $count=1 $X=0.36
+ $Y=1.835 $X2=0.485 $Y2=2.085
r96 1 18 400 $w=1.7e-07 $l=1.12577e-06 $layer=licon1_PDIFF $count=1 $X=0.36
+ $Y=1.835 $X2=0.485 $Y2=2.9
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4_4%VPWR 1 2 9 11 15 17 18 19 30 31 34
r100 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r101 30 31 1.43077 $w=1.7e-07 $l=1.105e-06 $layer=mcon $count=6 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r102 28 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=1.68 $Y2=3.33
r103 27 30 375.786 $w=1.68e-07 $l=5.76e-06 $layer=LI1_cond $X=2.16 $Y=3.33
+ $X2=7.92 $Y2=3.33
r104 27 28 1.43077 $w=1.7e-07 $l=1.105e-06 $layer=mcon $count=6 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r105 25 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.94 $Y=3.33
+ $X2=1.775 $Y2=3.33
r106 25 27 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=1.94 $Y=3.33
+ $X2=2.16 $Y2=3.33
r107 23 35 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r108 22 23 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r109 19 31 1.07034 $w=4.9e-07 $l=3.84e-06 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=7.92 $Y2=3.33
r110 19 28 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=2.16 $Y2=3.33
r111 17 22 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=0.75 $Y=3.33 $X2=0.72
+ $Y2=3.33
r112 17 18 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.75 $Y=3.33
+ $X2=0.915 $Y2=3.33
r113 13 34 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.775 $Y=3.245
+ $X2=1.775 $Y2=3.33
r114 13 15 30.208 $w=3.28e-07 $l=8.65e-07 $layer=LI1_cond $X=1.775 $Y=3.245
+ $X2=1.775 $Y2=2.38
r115 12 18 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.08 $Y=3.33
+ $X2=0.915 $Y2=3.33
r116 11 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.61 $Y=3.33
+ $X2=1.775 $Y2=3.33
r117 11 12 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=1.61 $Y=3.33
+ $X2=1.08 $Y2=3.33
r118 7 18 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.915 $Y=3.245
+ $X2=0.915 $Y2=3.33
r119 7 9 28.6365 $w=3.28e-07 $l=8.2e-07 $layer=LI1_cond $X=0.915 $Y=3.245
+ $X2=0.915 $Y2=2.425
r120 2 15 300 $w=1.7e-07 $l=6.11003e-07 $layer=licon1_PDIFF $count=2 $X=1.635
+ $Y=1.835 $X2=1.775 $Y2=2.38
r121 1 9 300 $w=1.7e-07 $l=6.56277e-07 $layer=licon1_PDIFF $count=2 $X=0.775
+ $Y=1.835 $X2=0.915 $Y2=2.425
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4_4%A_499_367# 1 2 3 4 15 17 18 21 23 27 29 33 35
+ 36
c48 18 0 1.83481e-20 $X=2.73 $Y=1.79
r49 31 33 6.4697 $w=1.78e-07 $l=1.05e-07 $layer=LI1_cond $X=5.73 $Y=1.875
+ $X2=5.73 $Y2=1.98
r50 30 36 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=4.97 $Y=1.79
+ $X2=4.875 $Y2=1.79
r51 29 31 6.82373 $w=1.7e-07 $l=1.25499e-07 $layer=LI1_cond $X=5.64 $Y=1.79
+ $X2=5.73 $Y2=1.875
r52 29 30 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.64 $Y=1.79
+ $X2=4.97 $Y2=1.79
r53 25 36 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=4.875 $Y=1.875
+ $X2=4.875 $Y2=1.79
r54 25 27 6.12919 $w=1.88e-07 $l=1.05e-07 $layer=LI1_cond $X=4.875 $Y=1.875
+ $X2=4.875 $Y2=1.98
r55 24 35 6.25164 $w=1.7e-07 $l=1.08e-07 $layer=LI1_cond $X=3.615 $Y=1.79
+ $X2=3.507 $Y2=1.79
r56 23 36 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=4.78 $Y=1.79
+ $X2=4.875 $Y2=1.79
r57 23 24 76.0053 $w=1.68e-07 $l=1.165e-06 $layer=LI1_cond $X=4.78 $Y=1.79
+ $X2=3.615 $Y2=1.79
r58 19 35 0.512231 $w=2.15e-07 $l=8.5e-08 $layer=LI1_cond $X=3.507 $Y=1.875
+ $X2=3.507 $Y2=1.79
r59 19 21 5.62821 $w=2.13e-07 $l=1.05e-07 $layer=LI1_cond $X=3.507 $Y=1.875
+ $X2=3.507 $Y2=1.98
r60 17 35 6.25164 $w=1.7e-07 $l=1.07e-07 $layer=LI1_cond $X=3.4 $Y=1.79
+ $X2=3.507 $Y2=1.79
r61 17 18 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.4 $Y=1.79 $X2=2.73
+ $Y2=1.79
r62 13 18 6.93832 $w=1.7e-07 $l=1.44375e-07 $layer=LI1_cond $X=2.622 $Y=1.875
+ $X2=2.73 $Y2=1.79
r63 13 15 5.62821 $w=2.13e-07 $l=1.05e-07 $layer=LI1_cond $X=2.622 $Y=1.875
+ $X2=2.622 $Y2=1.98
r64 4 33 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=5.595
+ $Y=1.835 $X2=5.735 $Y2=1.98
r65 3 27 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=4.735
+ $Y=1.835 $X2=4.875 $Y2=1.98
r66 2 21 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=3.355
+ $Y=1.835 $X2=3.495 $Y2=1.98
r67 1 15 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=2.495
+ $Y=1.835 $X2=2.635 $Y2=1.98
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4_4%A_864_367# 1 2 3 4 5 16 18 20 24 26 30 32 36
+ 38 40 42 47 49 51
r80 40 53 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.885 $Y=2.905
+ $X2=7.885 $Y2=2.99
r81 40 42 26.7157 $w=3.28e-07 $l=7.65e-07 $layer=LI1_cond $X=7.885 $Y=2.905
+ $X2=7.885 $Y2=2.14
r82 39 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.19 $Y=2.99
+ $X2=7.025 $Y2=2.99
r83 38 53 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.72 $Y=2.99
+ $X2=7.885 $Y2=2.99
r84 38 39 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=7.72 $Y=2.99
+ $X2=7.19 $Y2=2.99
r85 34 51 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.025 $Y=2.905
+ $X2=7.025 $Y2=2.99
r86 34 36 26.7157 $w=3.28e-07 $l=7.65e-07 $layer=LI1_cond $X=7.025 $Y=2.905
+ $X2=7.025 $Y2=2.14
r87 33 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.33 $Y=2.99
+ $X2=6.165 $Y2=2.99
r88 32 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.86 $Y=2.99
+ $X2=7.025 $Y2=2.99
r89 32 33 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=6.86 $Y=2.99
+ $X2=6.33 $Y2=2.99
r90 28 49 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.165 $Y=2.905
+ $X2=6.165 $Y2=2.99
r91 28 30 26.7157 $w=3.28e-07 $l=7.65e-07 $layer=LI1_cond $X=6.165 $Y=2.905
+ $X2=6.165 $Y2=2.14
r92 27 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.47 $Y=2.99
+ $X2=5.305 $Y2=2.99
r93 26 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6 $Y=2.99 $X2=6.165
+ $Y2=2.99
r94 26 27 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=6 $Y=2.99 $X2=5.47
+ $Y2=2.99
r95 22 47 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.305 $Y=2.905
+ $X2=5.305 $Y2=2.99
r96 22 24 26.7157 $w=3.28e-07 $l=7.65e-07 $layer=LI1_cond $X=5.305 $Y=2.905
+ $X2=5.305 $Y2=2.14
r97 21 45 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.61 $Y=2.99
+ $X2=4.445 $Y2=2.99
r98 20 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.14 $Y=2.99
+ $X2=5.305 $Y2=2.99
r99 20 21 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=5.14 $Y=2.99
+ $X2=4.61 $Y2=2.99
r100 16 45 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.445 $Y=2.905
+ $X2=4.445 $Y2=2.99
r101 16 18 26.7157 $w=3.28e-07 $l=7.65e-07 $layer=LI1_cond $X=4.445 $Y=2.905
+ $X2=4.445 $Y2=2.14
r102 5 53 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=7.745
+ $Y=1.835 $X2=7.885 $Y2=2.91
r103 5 42 400 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_PDIFF $count=1 $X=7.745
+ $Y=1.835 $X2=7.885 $Y2=2.14
r104 4 51 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=6.885
+ $Y=1.835 $X2=7.025 $Y2=2.91
r105 4 36 400 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_PDIFF $count=1 $X=6.885
+ $Y=1.835 $X2=7.025 $Y2=2.14
r106 3 49 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=6.025
+ $Y=1.835 $X2=6.165 $Y2=2.91
r107 3 30 400 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_PDIFF $count=1 $X=6.025
+ $Y=1.835 $X2=6.165 $Y2=2.14
r108 2 47 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=5.165
+ $Y=1.835 $X2=5.305 $Y2=2.91
r109 2 24 400 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_PDIFF $count=1 $X=5.165
+ $Y=1.835 $X2=5.305 $Y2=2.14
r110 1 45 400 $w=1.7e-07 $l=1.13578e-06 $layer=licon1_PDIFF $count=1 $X=4.32
+ $Y=1.835 $X2=4.445 $Y2=2.91
r111 1 18 400 $w=1.7e-07 $l=3.62146e-07 $layer=licon1_PDIFF $count=1 $X=4.32
+ $Y=1.835 $X2=4.445 $Y2=2.14
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4_4%Y 1 2 3 4 5 6 7 8 9 10 33 35 36 39 41 45 47
+ 51 53 57 59 63 65 69 73 75 77 78 81 85 87 89 91 93 94 95 96 97 102 105
r127 104 105 18.8154 $w=2.43e-07 $l=4e-07 $layer=LI1_cond $X=7.947 $Y=1.695
+ $X2=7.947 $Y2=1.295
r128 103 105 5.17423 $w=2.43e-07 $l=1.1e-07 $layer=LI1_cond $X=7.947 $Y=1.185
+ $X2=7.947 $Y2=1.295
r129 91 92 8.9027 $w=1.85e-07 $l=1.35e-07 $layer=LI1_cond $X=1.845 $Y=0.955
+ $X2=1.845 $Y2=1.09
r130 90 102 5.40251 $w=1.8e-07 $l=9.5e-08 $layer=LI1_cond $X=7.55 $Y=1.785
+ $X2=7.455 $Y2=1.785
r131 89 104 7.02594 $w=1.8e-07 $l=1.60823e-07 $layer=LI1_cond $X=7.825 $Y=1.785
+ $X2=7.947 $Y2=1.695
r132 89 90 16.9444 $w=1.78e-07 $l=2.75e-07 $layer=LI1_cond $X=7.825 $Y=1.785
+ $X2=7.55 $Y2=1.785
r133 88 100 2.30104 $w=1.8e-07 $l=1.18e-07 $layer=LI1_cond $X=7.55 $Y=1.095
+ $X2=7.432 $Y2=1.095
r134 87 103 7.02594 $w=1.8e-07 $l=1.60823e-07 $layer=LI1_cond $X=7.825 $Y=1.095
+ $X2=7.947 $Y2=1.185
r135 87 88 16.9444 $w=1.78e-07 $l=2.75e-07 $layer=LI1_cond $X=7.825 $Y=1.095
+ $X2=7.55 $Y2=1.095
r136 83 102 1.14861 $w=1.9e-07 $l=9e-08 $layer=LI1_cond $X=7.455 $Y=1.875
+ $X2=7.455 $Y2=1.785
r137 83 85 6.12919 $w=1.88e-07 $l=1.05e-07 $layer=LI1_cond $X=7.455 $Y=1.875
+ $X2=7.455 $Y2=1.98
r138 81 99 26.2679 $w=1.88e-07 $l=4.5e-07 $layer=LI1_cond $X=7.455 $Y=0.42
+ $X2=7.455 $Y2=0.87
r139 77 102 5.40251 $w=1.8e-07 $l=9.5e-08 $layer=LI1_cond $X=7.36 $Y=1.785
+ $X2=7.455 $Y2=1.785
r140 77 78 41.2828 $w=1.78e-07 $l=6.7e-07 $layer=LI1_cond $X=7.36 $Y=1.785
+ $X2=6.69 $Y2=1.785
r141 76 97 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=6.69 $Y=0.955
+ $X2=6.595 $Y2=0.955
r142 75 100 6.86562 $w=2.33e-07 $l=1.4e-07 $layer=LI1_cond $X=7.432 $Y=0.955
+ $X2=7.432 $Y2=1.095
r143 75 99 4.6247 $w=2.33e-07 $l=8.5e-08 $layer=LI1_cond $X=7.432 $Y=0.955
+ $X2=7.432 $Y2=0.87
r144 75 76 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=7.315 $Y=0.955
+ $X2=6.69 $Y2=0.955
r145 71 78 6.82297 $w=1.8e-07 $l=1.32571e-07 $layer=LI1_cond $X=6.595 $Y=1.875
+ $X2=6.69 $Y2=1.785
r146 71 73 6.12919 $w=1.88e-07 $l=1.05e-07 $layer=LI1_cond $X=6.595 $Y=1.875
+ $X2=6.595 $Y2=1.98
r147 67 97 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=6.595 $Y=0.87
+ $X2=6.595 $Y2=0.955
r148 67 69 25.6842 $w=1.88e-07 $l=4.4e-07 $layer=LI1_cond $X=6.595 $Y=0.87
+ $X2=6.595 $Y2=0.43
r149 66 96 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=5.83 $Y=0.955
+ $X2=5.735 $Y2=0.955
r150 65 97 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=6.5 $Y=0.955
+ $X2=6.595 $Y2=0.955
r151 65 66 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=6.5 $Y=0.955
+ $X2=5.83 $Y2=0.955
r152 61 96 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=5.735 $Y=0.87
+ $X2=5.735 $Y2=0.955
r153 61 63 25.6842 $w=1.88e-07 $l=4.4e-07 $layer=LI1_cond $X=5.735 $Y=0.87
+ $X2=5.735 $Y2=0.43
r154 60 95 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=4.97 $Y=0.955
+ $X2=4.875 $Y2=0.955
r155 59 96 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=5.64 $Y=0.955
+ $X2=5.735 $Y2=0.955
r156 59 60 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.64 $Y=0.955
+ $X2=4.97 $Y2=0.955
r157 55 95 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=4.875 $Y=0.87
+ $X2=4.875 $Y2=0.955
r158 55 57 25.6842 $w=1.88e-07 $l=4.4e-07 $layer=LI1_cond $X=4.875 $Y=0.87
+ $X2=4.875 $Y2=0.43
r159 54 94 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=4.11 $Y=0.955
+ $X2=4.015 $Y2=0.955
r160 53 95 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=4.78 $Y=0.955
+ $X2=4.875 $Y2=0.955
r161 53 54 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.78 $Y=0.955
+ $X2=4.11 $Y2=0.955
r162 49 94 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=4.015 $Y=0.87
+ $X2=4.015 $Y2=0.955
r163 49 51 25.6842 $w=1.88e-07 $l=4.4e-07 $layer=LI1_cond $X=4.015 $Y=0.87
+ $X2=4.015 $Y2=0.43
r164 48 93 5.78184 $w=1.7e-07 $l=9.8e-08 $layer=LI1_cond $X=3.25 $Y=0.955
+ $X2=3.152 $Y2=0.955
r165 47 94 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=3.92 $Y=0.955
+ $X2=4.015 $Y2=0.955
r166 47 48 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.92 $Y=0.955
+ $X2=3.25 $Y2=0.955
r167 43 93 0.85348 $w=1.95e-07 $l=8.5e-08 $layer=LI1_cond $X=3.152 $Y=0.87
+ $X2=3.152 $Y2=0.955
r168 43 45 25.0256 $w=1.93e-07 $l=4.4e-07 $layer=LI1_cond $X=3.152 $Y=0.87
+ $X2=3.152 $Y2=0.43
r169 42 91 1.22693 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.94 $Y=0.955
+ $X2=1.845 $Y2=0.955
r170 41 93 5.78184 $w=1.7e-07 $l=9.7e-08 $layer=LI1_cond $X=3.055 $Y=0.955
+ $X2=3.152 $Y2=0.955
r171 41 42 72.7433 $w=1.68e-07 $l=1.115e-06 $layer=LI1_cond $X=3.055 $Y=0.955
+ $X2=1.94 $Y2=0.955
r172 37 91 5.45789 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.845 $Y=0.87
+ $X2=1.845 $Y2=0.955
r173 37 39 26.2679 $w=1.88e-07 $l=4.5e-07 $layer=LI1_cond $X=1.845 $Y=0.87
+ $X2=1.845 $Y2=0.42
r174 35 92 1.22693 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.75 $Y=1.09
+ $X2=1.845 $Y2=1.09
r175 35 36 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.75 $Y=1.09
+ $X2=1.08 $Y2=1.09
r176 31 36 6.93832 $w=1.7e-07 $l=1.44375e-07 $layer=LI1_cond $X=0.972 $Y=1.005
+ $X2=1.08 $Y2=1.09
r177 31 33 31.3572 $w=2.13e-07 $l=5.85e-07 $layer=LI1_cond $X=0.972 $Y=1.005
+ $X2=0.972 $Y2=0.42
r178 10 85 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=7.315
+ $Y=1.835 $X2=7.455 $Y2=1.98
r179 9 73 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=6.455
+ $Y=1.835 $X2=6.595 $Y2=1.98
r180 8 81 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=7.315
+ $Y=0.235 $X2=7.455 $Y2=0.42
r181 7 69 91 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_NDIFF $count=2 $X=6.455
+ $Y=0.235 $X2=6.595 $Y2=0.43
r182 6 63 91 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_NDIFF $count=2 $X=5.595
+ $Y=0.235 $X2=5.735 $Y2=0.43
r183 5 57 91 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_NDIFF $count=2 $X=4.735
+ $Y=0.235 $X2=4.875 $Y2=0.43
r184 4 51 91 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_NDIFF $count=2 $X=3.875
+ $Y=0.235 $X2=4.015 $Y2=0.43
r185 3 45 91 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_NDIFF $count=2 $X=3.015
+ $Y=0.235 $X2=3.155 $Y2=0.43
r186 2 39 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=1.705
+ $Y=0.235 $X2=1.845 $Y2=0.42
r187 1 33 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=0.845
+ $Y=0.235 $X2=0.985 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__NOR4_4%VGND 1 2 3 4 5 6 7 8 9 30 34 40 44 48 50 54
+ 58 60 62 65 66 67 68 70 71 72 73 74 83 95 100 108 114 116 119 122 126
r133 125 126 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=0
+ $X2=7.92 $Y2=0
r134 122 123 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.96 $Y=0
+ $X2=6.96 $Y2=0
r135 119 120 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=0 $X2=6
+ $Y2=0
r136 116 117 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r137 113 114 11.2653 $w=7.83e-07 $l=1.6e-07 $layer=LI1_cond $X=2.725 $Y=0.307
+ $X2=2.885 $Y2=0.307
r138 110 113 1.29512 $w=7.83e-07 $l=8.5e-08 $layer=LI1_cond $X=2.64 $Y=0.307
+ $X2=2.725 $Y2=0.307
r139 110 111 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0
+ $X2=2.64 $Y2=0
r140 107 111 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0
+ $X2=2.64 $Y2=0
r141 106 110 7.3136 $w=7.83e-07 $l=4.8e-07 $layer=LI1_cond $X=2.16 $Y=0.307
+ $X2=2.64 $Y2=0.307
r142 106 108 9.58928 $w=7.83e-07 $l=5e-08 $layer=LI1_cond $X=2.16 $Y=0.307
+ $X2=2.11 $Y2=0.307
r143 106 107 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0
+ $X2=2.16 $Y2=0
r144 104 126 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0
+ $X2=7.92 $Y2=0
r145 104 123 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=0
+ $X2=6.96 $Y2=0
r146 103 104 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=0
+ $X2=7.44 $Y2=0
r147 101 122 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.19 $Y=0
+ $X2=7.025 $Y2=0
r148 101 103 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=7.19 $Y=0
+ $X2=7.44 $Y2=0
r149 100 125 4.746 $w=1.7e-07 $l=2.2e-07 $layer=LI1_cond $X=7.72 $Y=0 $X2=7.94
+ $Y2=0
r150 100 103 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=7.72 $Y=0
+ $X2=7.44 $Y2=0
r151 99 123 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0
+ $X2=6.96 $Y2=0
r152 99 120 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6
+ $Y2=0
r153 98 99 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r154 96 119 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.33 $Y=0
+ $X2=6.165 $Y2=0
r155 96 98 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=6.33 $Y=0 $X2=6.48
+ $Y2=0
r156 95 122 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.86 $Y=0
+ $X2=7.025 $Y2=0
r157 95 98 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=6.86 $Y=0 $X2=6.48
+ $Y2=0
r158 94 120 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=6
+ $Y2=0
r159 93 94 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r160 88 116 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.75 $Y=0
+ $X2=3.585 $Y2=0
r161 88 90 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=3.75 $Y=0 $X2=4.08
+ $Y2=0
r162 87 117 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r163 87 111 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0
+ $X2=2.64 $Y2=0
r164 86 114 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=3.12 $Y=0
+ $X2=2.885 $Y2=0
r165 86 87 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r166 83 116 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.42 $Y=0
+ $X2=3.585 $Y2=0
r167 83 86 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=3.42 $Y=0 $X2=3.12
+ $Y2=0
r168 82 107 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r169 81 82 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r170 78 82 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r171 77 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r172 74 94 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=5.04
+ $Y2=0
r173 74 117 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.6
+ $Y2=0
r174 74 90 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r175 72 93 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=5.14 $Y=0 $X2=5.04
+ $Y2=0
r176 72 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.14 $Y=0 $X2=5.305
+ $Y2=0
r177 70 90 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=4.28 $Y=0 $X2=4.08
+ $Y2=0
r178 70 71 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.28 $Y=0 $X2=4.445
+ $Y2=0
r179 69 93 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=4.61 $Y=0 $X2=5.04
+ $Y2=0
r180 69 71 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.61 $Y=0 $X2=4.445
+ $Y2=0
r181 67 81 3.26203 $w=1.68e-07 $l=5e-08 $layer=LI1_cond $X=1.25 $Y=0 $X2=1.2
+ $Y2=0
r182 67 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.25 $Y=0 $X2=1.415
+ $Y2=0
r183 65 77 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=0.39 $Y=0 $X2=0.24
+ $Y2=0
r184 65 66 8.14251 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=0.39 $Y=0 $X2=0.542
+ $Y2=0
r185 64 81 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=0.695 $Y=0 $X2=1.2
+ $Y2=0
r186 64 66 8.14251 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=0.695 $Y=0
+ $X2=0.542 $Y2=0
r187 60 125 3.02018 $w=3.3e-07 $l=1.09087e-07 $layer=LI1_cond $X=7.885 $Y=0.085
+ $X2=7.94 $Y2=0
r188 60 62 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=7.885 $Y=0.085
+ $X2=7.885 $Y2=0.38
r189 56 122 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.025 $Y=0.085
+ $X2=7.025 $Y2=0
r190 56 58 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=7.025 $Y=0.085
+ $X2=7.025 $Y2=0.535
r191 52 119 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.165 $Y=0.085
+ $X2=6.165 $Y2=0
r192 52 54 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=6.165 $Y=0.085
+ $X2=6.165 $Y2=0.535
r193 51 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.47 $Y=0 $X2=5.305
+ $Y2=0
r194 50 119 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6 $Y=0 $X2=6.165
+ $Y2=0
r195 50 51 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=6 $Y=0 $X2=5.47
+ $Y2=0
r196 46 73 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.305 $Y=0.085
+ $X2=5.305 $Y2=0
r197 46 48 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=5.305 $Y=0.085
+ $X2=5.305 $Y2=0.535
r198 42 71 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.445 $Y=0.085
+ $X2=4.445 $Y2=0
r199 42 44 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=4.445 $Y=0.085
+ $X2=4.445 $Y2=0.535
r200 38 116 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.585 $Y=0.085
+ $X2=3.585 $Y2=0
r201 38 40 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=3.585 $Y=0.085
+ $X2=3.585 $Y2=0.535
r202 37 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.58 $Y=0 $X2=1.415
+ $Y2=0
r203 37 108 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=1.58 $Y=0 $X2=2.11
+ $Y2=0
r204 32 68 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.415 $Y=0.085
+ $X2=1.415 $Y2=0
r205 32 34 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.415 $Y=0.085
+ $X2=1.415 $Y2=0.38
r206 28 66 0.649941 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.542 $Y=0.085
+ $X2=0.542 $Y2=0
r207 28 30 11.1466 $w=3.03e-07 $l=2.95e-07 $layer=LI1_cond $X=0.542 $Y=0.085
+ $X2=0.542 $Y2=0.38
r208 9 62 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=7.745
+ $Y=0.235 $X2=7.885 $Y2=0.38
r209 8 58 182 $w=1.7e-07 $l=3.63318e-07 $layer=licon1_NDIFF $count=1 $X=6.885
+ $Y=0.235 $X2=7.025 $Y2=0.535
r210 7 54 182 $w=1.7e-07 $l=3.63318e-07 $layer=licon1_NDIFF $count=1 $X=6.025
+ $Y=0.235 $X2=6.165 $Y2=0.535
r211 6 48 182 $w=1.7e-07 $l=3.63318e-07 $layer=licon1_NDIFF $count=1 $X=5.165
+ $Y=0.235 $X2=5.305 $Y2=0.535
r212 5 44 182 $w=1.7e-07 $l=3.63318e-07 $layer=licon1_NDIFF $count=1 $X=4.305
+ $Y=0.235 $X2=4.445 $Y2=0.535
r213 4 40 182 $w=1.7e-07 $l=3.63318e-07 $layer=licon1_NDIFF $count=1 $X=3.445
+ $Y=0.235 $X2=3.585 $Y2=0.535
r214 3 113 91 $w=1.7e-07 $l=7.24638e-07 $layer=licon1_NDIFF $count=2 $X=2.135
+ $Y=0.235 $X2=2.725 $Y2=0.535
r215 2 34 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.275
+ $Y=0.235 $X2=1.415 $Y2=0.38
r216 1 30 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.43
+ $Y=0.235 $X2=0.555 $Y2=0.38
.ends

