* File: sky130_fd_sc_lp__o32a_lp.pex.spice
* Created: Wed Sep  2 10:26:19 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O32A_LP%B1 1 3 5 6 8 10 11 12 13
c33 12 0 5.0416e-20 $X=0.24 $Y=1.295
r34 12 13 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.27 $Y=1.295
+ $X2=0.27 $Y2=1.665
r35 12 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=1.345 $X2=0.27 $Y2=1.345
r36 10 17 41.0924 $w=3.3e-07 $l=2.35e-07 $layer=POLY_cond $X=0.505 $Y=1.345
+ $X2=0.27 $Y2=1.345
r37 6 10 107.981 $w=1.54e-07 $l=3.48977e-07 $layer=POLY_cond $X=0.595 $Y=1
+ $X2=0.587 $Y2=1.345
r38 6 8 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.595 $Y=1 $X2=0.595
+ $Y2=0.715
r39 3 11 40.9178 $w=2.5e-07 $l=1.25e-07 $layer=POLY_cond $X=0.63 $Y=2.09
+ $X2=0.63 $Y2=1.965
r40 3 5 97.364 $w=2.5e-07 $l=5.05e-07 $layer=POLY_cond $X=0.63 $Y=2.09 $X2=0.63
+ $Y2=2.595
r41 1 10 51.6429 $w=1.54e-07 $l=1.68464e-07 $layer=POLY_cond $X=0.58 $Y=1.51
+ $X2=0.587 $Y2=1.345
r42 1 11 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=0.58 $Y=1.51
+ $X2=0.58 $Y2=1.965
.ends

.subckt PM_SKY130_FD_SC_LP__O32A_LP%B2 3 5 8 10 11 12 13 14 20 21
c48 21 0 6.35613e-20 $X=1.06 $Y=1.59
c49 20 0 5.0416e-20 $X=1.06 $Y=1.59
c50 10 0 1.04659e-19 $X=1.12 $Y=1.965
c51 8 0 1.89026e-19 $X=1.105 $Y=0.655
r52 20 23 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.06 $Y=1.59
+ $X2=1.06 $Y2=1.755
r53 20 22 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.06 $Y=1.59
+ $X2=1.06 $Y2=1.425
r54 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.06
+ $Y=1.59 $X2=1.06 $Y2=1.59
r55 13 14 7.2549 $w=6.08e-07 $l=3.7e-07 $layer=LI1_cond $X=0.92 $Y=2.405
+ $X2=0.92 $Y2=2.775
r56 12 13 7.2549 $w=6.08e-07 $l=3.7e-07 $layer=LI1_cond $X=0.92 $Y=2.035
+ $X2=0.92 $Y2=2.405
r57 11 12 7.2549 $w=6.08e-07 $l=3.7e-07 $layer=LI1_cond $X=0.92 $Y=1.665
+ $X2=0.92 $Y2=2.035
r58 11 21 1.47059 $w=6.08e-07 $l=7.5e-08 $layer=LI1_cond $X=0.92 $Y=1.665
+ $X2=0.92 $Y2=1.59
r59 10 23 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=1.07 $Y=1.965
+ $X2=1.07 $Y2=1.755
r60 8 22 394.83 $w=1.5e-07 $l=7.7e-07 $layer=POLY_cond $X=1.105 $Y=0.655
+ $X2=1.105 $Y2=1.425
r61 3 10 40.9178 $w=2.5e-07 $l=1.25e-07 $layer=POLY_cond $X=1.12 $Y=2.09
+ $X2=1.12 $Y2=1.965
r62 3 5 97.364 $w=2.5e-07 $l=5.05e-07 $layer=POLY_cond $X=1.12 $Y=2.09 $X2=1.12
+ $Y2=2.595
.ends

.subckt PM_SKY130_FD_SC_LP__O32A_LP%A3 3 9 10 11 12 15 16
c48 16 0 2.75793e-19 $X=1.6 $Y=1.56
c49 11 0 6.35613e-20 $X=1.747 $Y=2.02
r50 15 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.6 $Y=1.56 $X2=1.6
+ $Y2=1.725
r51 15 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.6 $Y=1.56 $X2=1.6
+ $Y2=1.395
r52 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.6
+ $Y=1.56 $X2=1.6 $Y2=1.56
r53 12 16 3.36129 $w=3.58e-07 $l=1.05e-07 $layer=LI1_cond $X=1.615 $Y=1.665
+ $X2=1.615 $Y2=1.56
r54 10 11 47.1291 $w=2.5e-07 $l=1.5e-07 $layer=POLY_cond $X=1.747 $Y=1.87
+ $X2=1.747 $Y2=2.02
r55 10 18 74.3511 $w=1.5e-07 $l=1.45e-07 $layer=POLY_cond $X=1.69 $Y=1.87
+ $X2=1.69 $Y2=1.725
r56 9 11 110.86 $w=2.5e-07 $l=5.75e-07 $layer=POLY_cond $X=1.755 $Y=2.595
+ $X2=1.755 $Y2=2.02
r57 3 17 379.447 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=1.535 $Y=0.655
+ $X2=1.535 $Y2=1.395
.ends

.subckt PM_SKY130_FD_SC_LP__O32A_LP%A2 3 7 9 10 11 14 15
c48 15 0 1.70596e-19 $X=2.14 $Y=1.495
r49 14 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.14 $Y=1.495
+ $X2=2.14 $Y2=1.66
r50 14 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.14 $Y=1.495
+ $X2=2.14 $Y2=1.33
r51 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.14
+ $Y=1.495 $X2=2.14 $Y2=1.495
r52 11 15 5.93683 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=2.14 $Y=1.665
+ $X2=2.14 $Y2=1.495
r53 10 17 156.394 $w=1.5e-07 $l=3.05e-07 $layer=POLY_cond $X=2.195 $Y=1.965
+ $X2=2.195 $Y2=1.66
r54 7 10 40.9178 $w=2.5e-07 $l=1.25e-07 $layer=POLY_cond $X=2.245 $Y=2.09
+ $X2=2.245 $Y2=1.965
r55 7 9 97.364 $w=2.5e-07 $l=5.05e-07 $layer=POLY_cond $X=2.245 $Y=2.09
+ $X2=2.245 $Y2=2.595
r56 3 16 346.117 $w=1.5e-07 $l=6.75e-07 $layer=POLY_cond $X=2.125 $Y=0.655
+ $X2=2.125 $Y2=1.33
.ends

.subckt PM_SKY130_FD_SC_LP__O32A_LP%A1 3 8 10 11 12 13 14 17 18 19
c48 18 0 1.64536e-19 $X=2.68 $Y=1.56
c49 13 0 3.26804e-19 $X=2.735 $Y=1.95
c50 11 0 1.44963e-19 $X=2.587 $Y=0.94
c51 8 0 2.9647e-19 $X=2.735 $Y=2.075
r52 17 20 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.68 $Y=1.56
+ $X2=2.68 $Y2=1.725
r53 17 19 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.68 $Y=1.56
+ $X2=2.68 $Y2=1.395
r54 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.68
+ $Y=1.56 $X2=2.68 $Y2=1.56
r55 14 18 3.66686 $w=3.28e-07 $l=1.05e-07 $layer=LI1_cond $X=2.68 $Y=1.665
+ $X2=2.68 $Y2=1.56
r56 13 20 115.372 $w=1.5e-07 $l=2.25e-07 $layer=POLY_cond $X=2.685 $Y=1.95
+ $X2=2.685 $Y2=1.725
r57 12 19 156.394 $w=1.5e-07 $l=3.05e-07 $layer=POLY_cond $X=2.62 $Y=1.09
+ $X2=2.62 $Y2=1.395
r58 11 12 44.7709 $w=2.15e-07 $l=1.5e-07 $layer=POLY_cond $X=2.587 $Y=0.94
+ $X2=2.587 $Y2=1.09
r59 8 13 40.9178 $w=2.5e-07 $l=1.25e-07 $layer=POLY_cond $X=2.735 $Y=2.075
+ $X2=2.735 $Y2=1.95
r60 8 10 100.256 $w=2.5e-07 $l=5.2e-07 $layer=POLY_cond $X=2.735 $Y=2.075
+ $X2=2.735 $Y2=2.595
r61 3 11 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.555 $Y=0.655
+ $X2=2.555 $Y2=0.94
.ends

.subckt PM_SKY130_FD_SC_LP__O32A_LP%A_134_101# 1 2 7 9 12 16 19 21 24 26 27 30
+ 32 33 37 38 40 41
c96 41 0 1.56208e-19 $X=3.205 $Y=1.74
c97 40 0 1.96001e-19 $X=3.11 $Y=1.96
c98 33 0 1.78918e-20 $X=1.655 $Y=2.045
c99 21 0 5.01836e-20 $X=3.237 $Y=1.74
c100 12 0 1.14352e-19 $X=3.275 $Y=2.595
r101 40 41 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=3.11 $Y=1.96
+ $X2=3.11 $Y2=1.74
r102 37 38 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.22
+ $Y=1.235 $X2=3.22 $Y2=1.235
r103 35 41 8.99121 $w=3.58e-07 $l=1.8e-07 $layer=LI1_cond $X=3.205 $Y=1.56
+ $X2=3.205 $Y2=1.74
r104 35 37 10.404 $w=3.58e-07 $l=3.25e-07 $layer=LI1_cond $X=3.205 $Y=1.56
+ $X2=3.205 $Y2=1.235
r105 34 37 2.72105 $w=3.58e-07 $l=8.5e-08 $layer=LI1_cond $X=3.205 $Y=1.15
+ $X2=3.205 $Y2=1.235
r106 32 40 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.025 $Y=2.045
+ $X2=3.11 $Y2=1.96
r107 32 33 89.3797 $w=1.68e-07 $l=1.37e-06 $layer=LI1_cond $X=3.025 $Y=2.045
+ $X2=1.655 $Y2=2.045
r108 28 33 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.53 $Y=2.13
+ $X2=1.655 $Y2=2.045
r109 28 30 5.07075 $w=2.48e-07 $l=1.1e-07 $layer=LI1_cond $X=1.53 $Y=2.13
+ $X2=1.53 $Y2=2.24
r110 26 34 23.5781 $w=9e-08 $l=2.18403e-07 $layer=LI1_cond $X=3.025 $Y=1.065
+ $X2=3.205 $Y2=1.15
r111 26 27 133.743 $w=1.68e-07 $l=2.05e-06 $layer=LI1_cond $X=3.025 $Y=1.065
+ $X2=0.975 $Y2=1.065
r112 22 27 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.81 $Y=0.98
+ $X2=0.975 $Y2=1.065
r113 22 24 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=0.81 $Y=0.98 $X2=0.81
+ $Y2=0.78
r114 20 38 51.0643 $w=3.65e-07 $l=3.23e-07 $layer=POLY_cond $X=3.237 $Y=1.558
+ $X2=3.237 $Y2=1.235
r115 20 21 33.1107 $w=3.65e-07 $l=1.82e-07 $layer=POLY_cond $X=3.237 $Y=1.558
+ $X2=3.237 $Y2=1.74
r116 19 38 22.9236 $w=3.65e-07 $l=1.45e-07 $layer=POLY_cond $X=3.237 $Y=1.09
+ $X2=3.237 $Y2=1.235
r117 12 21 212.428 $w=2.5e-07 $l=8.55e-07 $layer=POLY_cond $X=3.275 $Y=2.595
+ $X2=3.275 $Y2=1.74
r118 7 19 25.7148 $w=3.65e-07 $l=1.5e-07 $layer=POLY_cond $X=3.165 $Y=0.94
+ $X2=3.165 $Y2=1.09
r119 7 16 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.345 $Y=0.94
+ $X2=3.345 $Y2=0.655
r120 7 9 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.985 $Y=0.94
+ $X2=2.985 $Y2=0.655
r121 2 30 300 $w=1.7e-07 $l=3.09112e-07 $layer=licon1_PDIFF $count=2 $X=1.245
+ $Y=2.095 $X2=1.49 $Y2=2.24
r122 1 24 182 $w=1.7e-07 $l=3.37824e-07 $layer=licon1_NDIFF $count=1 $X=0.67
+ $Y=0.505 $X2=0.81 $Y2=0.78
.ends

.subckt PM_SKY130_FD_SC_LP__O32A_LP%VPWR 1 2 7 9 15 18 19 20 30 31
r42 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r43 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r44 28 31 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r45 27 28 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r46 25 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r47 24 27 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=0.72 $Y=3.33
+ $X2=2.64 $Y2=3.33
r48 24 25 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r49 22 34 3.93235 $w=1.7e-07 $l=2.18e-07 $layer=LI1_cond $X=0.435 $Y=3.33
+ $X2=0.217 $Y2=3.33
r50 22 24 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.435 $Y=3.33
+ $X2=0.72 $Y2=3.33
r51 20 28 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=2.64 $Y2=3.33
r52 20 25 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=0.72 $Y2=3.33
r53 18 27 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=2.835 $Y=3.33
+ $X2=2.64 $Y2=3.33
r54 18 19 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.835 $Y=3.33 $X2=3
+ $Y2=3.33
r55 17 30 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=3.165 $Y=3.33
+ $X2=3.6 $Y2=3.33
r56 17 19 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.165 $Y=3.33 $X2=3
+ $Y2=3.33
r57 13 19 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3 $Y=3.245 $X2=3
+ $Y2=3.33
r58 13 15 26.8903 $w=3.28e-07 $l=7.7e-07 $layer=LI1_cond $X=3 $Y=3.245 $X2=3
+ $Y2=2.475
r59 9 12 32.7294 $w=2.48e-07 $l=7.1e-07 $layer=LI1_cond $X=0.31 $Y=2.24 $X2=0.31
+ $Y2=2.95
r60 7 34 3.21082 $w=2.5e-07 $l=1.28662e-07 $layer=LI1_cond $X=0.31 $Y=3.245
+ $X2=0.217 $Y2=3.33
r61 7 12 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=0.31 $Y=3.245
+ $X2=0.31 $Y2=2.95
r62 2 15 300 $w=1.7e-07 $l=4.44522e-07 $layer=licon1_PDIFF $count=2 $X=2.86
+ $Y=2.095 $X2=3 $Y2=2.475
r63 1 12 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.205
+ $Y=2.095 $X2=0.35 $Y2=2.95
r64 1 9 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.205
+ $Y=2.095 $X2=0.35 $Y2=2.24
.ends

.subckt PM_SKY130_FD_SC_LP__O32A_LP%X 1 2 10 13 14 15 30 32
c23 13 0 1.00469e-19 $X=3.515 $Y=1.95
r24 20 32 2.0808 $w=3.58e-07 $l=6.5e-08 $layer=LI1_cond $X=3.555 $Y=2.1
+ $X2=3.555 $Y2=2.035
r25 14 15 11.8446 $w=3.58e-07 $l=3.7e-07 $layer=LI1_cond $X=3.555 $Y=2.405
+ $X2=3.555 $Y2=2.775
r26 14 23 5.28203 $w=3.58e-07 $l=1.65e-07 $layer=LI1_cond $X=3.555 $Y=2.405
+ $X2=3.555 $Y2=2.24
r27 13 32 0.320123 $w=3.58e-07 $l=1e-08 $layer=LI1_cond $X=3.555 $Y=2.025
+ $X2=3.555 $Y2=2.035
r28 13 30 6.59029 $w=3.58e-07 $l=1.05e-07 $layer=LI1_cond $X=3.555 $Y=2.025
+ $X2=3.555 $Y2=1.92
r29 13 23 4.1616 $w=3.58e-07 $l=1.3e-07 $layer=LI1_cond $X=3.555 $Y=2.11
+ $X2=3.555 $Y2=2.24
r30 13 20 0.320123 $w=3.58e-07 $l=1e-08 $layer=LI1_cond $X=3.555 $Y=2.11
+ $X2=3.555 $Y2=2.1
r31 12 30 67.5241 $w=1.68e-07 $l=1.035e-06 $layer=LI1_cond $X=3.65 $Y=0.885
+ $X2=3.65 $Y2=1.92
r32 10 12 10.6751 $w=3.38e-07 $l=2.3e-07 $layer=LI1_cond $X=3.565 $Y=0.655
+ $X2=3.565 $Y2=0.885
r33 2 23 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=3.4
+ $Y=2.095 $X2=3.54 $Y2=2.24
r34 1 10 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=3.42
+ $Y=0.445 $X2=3.56 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__O32A_LP%A_31_101# 1 2 3 12 14 15 19 20 21 23
c42 23 0 1.44963e-19 $X=2.34 $Y=0.61
r43 23 25 4.84026 $w=2.48e-07 $l=1.05e-07 $layer=LI1_cond $X=2.3 $Y=0.61 $X2=2.3
+ $Y2=0.715
r44 20 25 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.175 $Y=0.715
+ $X2=2.3 $Y2=0.715
r45 20 21 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.175 $Y=0.715
+ $X2=1.485 $Y2=0.715
r46 17 21 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.32 $Y=0.63
+ $X2=1.485 $Y2=0.715
r47 17 19 0.69845 $w=3.28e-07 $l=2e-08 $layer=LI1_cond $X=1.32 $Y=0.63 $X2=1.32
+ $Y2=0.61
r48 16 19 6.11144 $w=3.28e-07 $l=1.75e-07 $layer=LI1_cond $X=1.32 $Y=0.435
+ $X2=1.32 $Y2=0.61
r49 14 16 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.155 $Y=0.35
+ $X2=1.32 $Y2=0.435
r50 14 15 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.155 $Y=0.35
+ $X2=0.465 $Y2=0.35
r51 10 15 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.3 $Y=0.435
+ $X2=0.465 $Y2=0.35
r52 10 12 9.7783 $w=3.28e-07 $l=2.8e-07 $layer=LI1_cond $X=0.3 $Y=0.435 $X2=0.3
+ $Y2=0.715
r53 3 23 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=2.2
+ $Y=0.445 $X2=2.34 $Y2=0.61
r54 2 19 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=1.18
+ $Y=0.445 $X2=1.32 $Y2=0.61
r55 1 12 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.155
+ $Y=0.505 $X2=0.3 $Y2=0.715
.ends

.subckt PM_SKY130_FD_SC_LP__O32A_LP%VGND 1 2 9 11 15 17 19 26 27 30 33
r43 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r44 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r45 27 34 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=2.64
+ $Y2=0
r46 26 27 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r47 24 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.935 $Y=0 $X2=2.77
+ $Y2=0
r48 24 26 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=2.935 $Y=0 $X2=3.6
+ $Y2=0
r49 22 31 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=0.24 $Y=0 $X2=1.68
+ $Y2=0
r50 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r51 19 30 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.665 $Y=0 $X2=1.83
+ $Y2=0
r52 19 21 92.9679 $w=1.68e-07 $l=1.425e-06 $layer=LI1_cond $X=1.665 $Y=0
+ $X2=0.24 $Y2=0
r53 17 34 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=2.64
+ $Y2=0
r54 17 31 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=1.68
+ $Y2=0
r55 13 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.77 $Y=0.085
+ $X2=2.77 $Y2=0
r56 13 15 18.3343 $w=3.28e-07 $l=5.25e-07 $layer=LI1_cond $X=2.77 $Y=0.085
+ $X2=2.77 $Y2=0.61
r57 12 30 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.995 $Y=0 $X2=1.83
+ $Y2=0
r58 11 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.605 $Y=0 $X2=2.77
+ $Y2=0
r59 11 12 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=2.605 $Y=0 $X2=1.995
+ $Y2=0
r60 7 30 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.83 $Y=0.085 $X2=1.83
+ $Y2=0
r61 7 9 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=1.83 $Y=0.085 $X2=1.83
+ $Y2=0.285
r62 2 15 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=2.63
+ $Y=0.445 $X2=2.77 $Y2=0.61
r63 1 9 182 $w=1.7e-07 $l=2.89137e-07 $layer=licon1_NDIFF $count=1 $X=1.61
+ $Y=0.445 $X2=1.83 $Y2=0.285
.ends

