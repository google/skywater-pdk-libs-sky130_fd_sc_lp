* File: sky130_fd_sc_lp__inv_2.pex.spice
* Created: Fri Aug 28 10:38:13 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__INV_2%A 1 3 6 8 10 13 15 16 24
r33 23 24 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=0.485 $Y=1.46
+ $X2=0.915 $Y2=1.46
r34 20 23 27.1035 $w=3.3e-07 $l=1.55e-07 $layer=POLY_cond $X=0.33 $Y=1.46
+ $X2=0.485 $Y2=1.46
r35 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.33
+ $Y=1.46 $X2=0.33 $Y2=1.46
r36 16 21 6.75002 $w=3.48e-07 $l=2.05e-07 $layer=LI1_cond $X=0.26 $Y=1.665
+ $X2=0.26 $Y2=1.46
r37 15 21 5.43295 $w=3.48e-07 $l=1.65e-07 $layer=LI1_cond $X=0.26 $Y=1.295
+ $X2=0.26 $Y2=1.46
r38 11 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.915 $Y=1.625
+ $X2=0.915 $Y2=1.46
r39 11 13 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=0.915 $Y=1.625
+ $X2=0.915 $Y2=2.465
r40 8 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.915 $Y=1.295
+ $X2=0.915 $Y2=1.46
r41 8 10 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.915 $Y=1.295
+ $X2=0.915 $Y2=0.765
r42 4 23 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.485 $Y=1.625
+ $X2=0.485 $Y2=1.46
r43 4 6 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=0.485 $Y=1.625
+ $X2=0.485 $Y2=2.465
r44 1 23 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.485 $Y=1.295
+ $X2=0.485 $Y2=1.46
r45 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.485 $Y=1.295
+ $X2=0.485 $Y2=0.765
.ends

.subckt PM_SKY130_FD_SC_LP__INV_2%VPWR 1 2 7 9 13 15 19 21 31
r21 30 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r22 27 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r23 22 27 4.75569 $w=1.7e-07 $l=2.18e-07 $layer=LI1_cond $X=0.435 $Y=3.33
+ $X2=0.217 $Y2=3.33
r24 22 24 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.435 $Y=3.33
+ $X2=0.72 $Y2=3.33
r25 21 30 4.31554 $w=1.7e-07 $l=2.17e-07 $layer=LI1_cond $X=1.005 $Y=3.33
+ $X2=1.222 $Y2=3.33
r26 21 24 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.005 $Y=3.33
+ $X2=0.72 $Y2=3.33
r27 19 31 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r28 19 28 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r29 19 24 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r30 15 18 38.5472 $w=2.88e-07 $l=9.7e-07 $layer=LI1_cond $X=1.15 $Y=1.98
+ $X2=1.15 $Y2=2.95
r31 13 30 3.1223 $w=2.9e-07 $l=1.15521e-07 $layer=LI1_cond $X=1.15 $Y=3.245
+ $X2=1.222 $Y2=3.33
r32 13 18 11.7231 $w=2.88e-07 $l=2.95e-07 $layer=LI1_cond $X=1.15 $Y=3.245
+ $X2=1.15 $Y2=2.95
r33 9 12 30.208 $w=3.28e-07 $l=8.65e-07 $layer=LI1_cond $X=0.27 $Y=2.085
+ $X2=0.27 $Y2=2.95
r34 7 27 3.01048 $w=3.3e-07 $l=1.08305e-07 $layer=LI1_cond $X=0.27 $Y=3.245
+ $X2=0.217 $Y2=3.33
r35 7 12 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.27 $Y=3.245
+ $X2=0.27 $Y2=2.95
r36 2 18 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=0.99
+ $Y=1.835 $X2=1.13 $Y2=2.95
r37 2 15 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.99
+ $Y=1.835 $X2=1.13 $Y2=1.98
r38 1 12 400 $w=1.7e-07 $l=1.17584e-06 $layer=licon1_PDIFF $count=1 $X=0.145
+ $Y=1.835 $X2=0.27 $Y2=2.95
r39 1 9 400 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_PDIFF $count=1 $X=0.145
+ $Y=1.835 $X2=0.27 $Y2=2.085
.ends

.subckt PM_SKY130_FD_SC_LP__INV_2%Y 1 2 7 8 9 10 11 12 13
r16 13 39 6.76434 $w=2.28e-07 $l=1.35e-07 $layer=LI1_cond $X=0.72 $Y=2.775
+ $X2=0.72 $Y2=2.91
r17 12 13 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.72 $Y=2.405
+ $X2=0.72 $Y2=2.775
r18 11 12 19.5414 $w=2.28e-07 $l=3.9e-07 $layer=LI1_cond $X=0.72 $Y=2.015
+ $X2=0.72 $Y2=2.405
r19 10 11 17.5372 $w=2.28e-07 $l=3.5e-07 $layer=LI1_cond $X=0.72 $Y=1.665
+ $X2=0.72 $Y2=2.015
r20 9 10 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.72 $Y=1.295
+ $X2=0.72 $Y2=1.665
r21 8 9 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.72 $Y=0.925 $X2=0.72
+ $Y2=1.295
r22 7 8 22.7983 $w=2.28e-07 $l=4.55e-07 $layer=LI1_cond $X=0.72 $Y=0.47 $X2=0.72
+ $Y2=0.925
r23 2 39 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=0.56
+ $Y=1.835 $X2=0.7 $Y2=2.91
r24 2 11 400 $w=1.7e-07 $l=2.4e-07 $layer=licon1_PDIFF $count=1 $X=0.56 $Y=1.835
+ $X2=0.7 $Y2=2.015
r25 1 7 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=0.56
+ $Y=0.345 $X2=0.7 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_LP__INV_2%VGND 1 2 7 9 11 13 15 17 27
r20 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r21 23 24 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r22 18 23 4.75569 $w=1.7e-07 $l=2.18e-07 $layer=LI1_cond $X=0.435 $Y=0 $X2=0.217
+ $Y2=0
r23 18 20 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.435 $Y=0 $X2=0.72
+ $Y2=0
r24 17 26 4.31554 $w=1.7e-07 $l=2.17e-07 $layer=LI1_cond $X=1.005 $Y=0 $X2=1.222
+ $Y2=0
r25 17 20 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.005 $Y=0 $X2=0.72
+ $Y2=0
r26 15 27 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r27 15 24 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r28 15 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r29 11 26 3.1223 $w=2.9e-07 $l=1.15521e-07 $layer=LI1_cond $X=1.15 $Y=0.085
+ $X2=1.222 $Y2=0
r30 11 13 16.0945 $w=2.88e-07 $l=4.05e-07 $layer=LI1_cond $X=1.15 $Y=0.085
+ $X2=1.15 $Y2=0.49
r31 7 23 3.01048 $w=3.3e-07 $l=1.08305e-07 $layer=LI1_cond $X=0.27 $Y=0.085
+ $X2=0.217 $Y2=0
r32 7 9 14.1436 $w=3.28e-07 $l=4.05e-07 $layer=LI1_cond $X=0.27 $Y=0.085
+ $X2=0.27 $Y2=0.49
r33 2 13 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=0.99
+ $Y=0.345 $X2=1.13 $Y2=0.49
r34 1 9 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.145
+ $Y=0.345 $X2=0.27 $Y2=0.49
.ends

