* NGSPICE file created from sky130_fd_sc_lp__a2111oi_0.ext - technology: sky130A

.subckt sky130_fd_sc_lp__a2111oi_0 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
M1000 a_432_47# A1 Y VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=2.352e+11p ps=2.8e+06u
M1001 a_318_483# A2 VPWR VPB phighvt w=640000u l=150000u
+  ad=3.488e+11p pd=3.65e+06u as=2.432e+11p ps=2.04e+06u
M1002 Y D1 VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=3.696e+11p ps=4.28e+06u
M1003 a_174_483# D1 Y VPB phighvt w=640000u l=150000u
+  ad=1.344e+11p pd=1.7e+06u as=1.888e+11p ps=1.87e+06u
M1004 a_246_483# C1 a_174_483# VPB phighvt w=640000u l=150000u
+  ad=1.344e+11p pd=1.7e+06u as=0p ps=0u
M1005 VPWR A1 a_318_483# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 Y B1 VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND A2 a_432_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND C1 Y VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_318_483# B1 a_246_483# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

