* File: sky130_fd_sc_lp__sdfstp_lp.pex.spice
* Created: Fri Aug 28 11:30:03 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__SDFSTP_LP%SCE 3 7 11 15 19 23 24 30 31 32 36 37 39
+ 40 48 51 55
r96 44 46 17.4861 $w=3.3e-07 $l=1e-07 $layer=POLY_cond $X=0.545 $Y=1.02
+ $X2=0.645 $Y2=1.02
r97 40 55 8.06514 $w=4.68e-07 $l=1.15e-07 $layer=LI1_cond $X=2.16 $Y=1.045
+ $X2=2.275 $Y2=1.045
r98 39 51 4.00199 $w=4.68e-07 $l=1.15e-07 $layer=LI1_cond $X=1.68 $Y=1.045
+ $X2=1.565 $Y2=1.045
r99 36 37 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.675
+ $Y=1.285 $X2=2.675 $Y2=1.285
r100 34 36 0.177299 $w=3.23e-07 $l=5e-09 $layer=LI1_cond $X=2.672 $Y=1.28
+ $X2=2.672 $Y2=1.285
r101 32 34 7.72402 $w=1.7e-07 $l=2.00035e-07 $layer=LI1_cond $X=2.51 $Y=1.195
+ $X2=2.672 $Y2=1.28
r102 32 55 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=2.51 $Y=1.195
+ $X2=2.275 $Y2=1.195
r103 31 39 3.05382 $w=4.68e-07 $l=1.2e-07 $layer=LI1_cond $X=1.8 $Y=1.045
+ $X2=1.68 $Y2=1.045
r104 30 40 3.05382 $w=4.68e-07 $l=1.2e-07 $layer=LI1_cond $X=2.04 $Y=1.045
+ $X2=2.16 $Y2=1.045
r105 30 31 6.10763 $w=4.68e-07 $l=2.4e-07 $layer=LI1_cond $X=2.04 $Y=1.045
+ $X2=1.8 $Y2=1.045
r106 28 48 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=0.915 $Y=1.02
+ $X2=1.005 $Y2=1.02
r107 28 46 47.2125 $w=3.3e-07 $l=2.7e-07 $layer=POLY_cond $X=0.915 $Y=1.02
+ $X2=0.645 $Y2=1.02
r108 27 51 22.6996 $w=3.28e-07 $l=6.5e-07 $layer=LI1_cond $X=0.915 $Y=1.02
+ $X2=1.565 $Y2=1.02
r109 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.915
+ $Y=1.02 $X2=0.915 $Y2=1.02
r110 23 37 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.675 $Y=1.625
+ $X2=2.675 $Y2=1.285
r111 23 24 31.2043 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.675 $Y=1.625
+ $X2=2.675 $Y2=1.79
r112 22 37 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.675 $Y=1.12
+ $X2=2.675 $Y2=1.285
r113 19 24 183.856 $w=2.5e-07 $l=7.4e-07 $layer=POLY_cond $X=2.655 $Y=2.53
+ $X2=2.655 $Y2=1.79
r114 15 22 346.117 $w=1.5e-07 $l=6.75e-07 $layer=POLY_cond $X=2.585 $Y=0.445
+ $X2=2.585 $Y2=1.12
r115 9 48 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.005 $Y=0.855
+ $X2=1.005 $Y2=1.02
r116 9 11 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=1.005 $Y=0.855
+ $X2=1.005 $Y2=0.445
r117 5 46 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.645 $Y=0.855
+ $X2=0.645 $Y2=1.02
r118 5 7 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=0.645 $Y=0.855
+ $X2=0.645 $Y2=0.445
r119 1 44 9.34494 $w=2.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.545 $Y=1.185
+ $X2=0.545 $Y2=1.02
r120 1 3 337.897 $w=2.5e-07 $l=1.36e-06 $layer=POLY_cond $X=0.545 $Y=1.185
+ $X2=0.545 $Y2=2.545
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSTP_LP%A_27_409# 1 2 9 12 13 15 16 17 20 23 26 32
+ 36 39
c69 32 0 1.32997e-19 $X=1.22 $Y=1.625
r70 36 38 6.28597 $w=4.78e-07 $l=2.05e-07 $layer=LI1_cond $X=0.355 $Y=0.47
+ $X2=0.355 $Y2=0.675
r71 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.22
+ $Y=1.625 $X2=1.22 $Y2=1.625
r72 30 39 1.34256 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=0.445 $Y=1.625
+ $X2=0.28 $Y2=1.625
r73 30 32 27.0649 $w=3.28e-07 $l=7.75e-07 $layer=LI1_cond $X=0.445 $Y=1.625
+ $X2=1.22 $Y2=1.625
r74 26 28 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=0.28 $Y=2.19 $X2=0.28
+ $Y2=2.9
r75 24 39 5.16603 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=0.28 $Y=1.79
+ $X2=0.28 $Y2=1.625
r76 24 26 13.969 $w=3.28e-07 $l=4e-07 $layer=LI1_cond $X=0.28 $Y=1.79 $X2=0.28
+ $Y2=2.19
r77 23 39 5.16603 $w=3.3e-07 $l=1.65e-07 $layer=LI1_cond $X=0.28 $Y=1.46
+ $X2=0.28 $Y2=1.625
r78 23 38 27.4142 $w=3.28e-07 $l=7.85e-07 $layer=LI1_cond $X=0.28 $Y=1.46
+ $X2=0.28 $Y2=0.675
r79 18 20 41.0213 $w=1.5e-07 $l=8e-08 $layer=POLY_cond $X=1.685 $Y=0.805
+ $X2=1.765 $Y2=0.805
r80 16 33 50.7098 $w=3.3e-07 $l=2.9e-07 $layer=POLY_cond $X=1.51 $Y=1.625
+ $X2=1.22 $Y2=1.625
r81 16 17 1.50692 $w=3.3e-07 $l=1.25e-07 $layer=POLY_cond $X=1.51 $Y=1.625
+ $X2=1.635 $Y2=1.625
r82 13 20 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.765 $Y=0.73
+ $X2=1.765 $Y2=0.805
r83 13 15 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=1.765 $Y=0.73
+ $X2=1.765 $Y2=0.445
r84 12 17 30.2679 $w=2e-07 $l=1.88348e-07 $layer=POLY_cond $X=1.685 $Y=1.46
+ $X2=1.635 $Y2=1.625
r85 11 18 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.685 $Y=0.88
+ $X2=1.685 $Y2=0.805
r86 11 12 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=1.685 $Y=0.88
+ $X2=1.685 $Y2=1.46
r87 7 17 30.2679 $w=2e-07 $l=1.65e-07 $layer=POLY_cond $X=1.635 $Y=1.79
+ $X2=1.635 $Y2=1.625
r88 7 9 183.856 $w=2.5e-07 $l=7.4e-07 $layer=POLY_cond $X=1.635 $Y=1.79
+ $X2=1.635 $Y2=2.53
r89 2 28 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.045 $X2=0.28 $Y2=2.9
r90 2 26 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.045 $X2=0.28 $Y2=2.19
r91 1 36 182 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_NDIFF $count=1 $X=0.285
+ $Y=0.235 $X2=0.43 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSTP_LP%D 3 7 9 10 14
c41 14 0 1.32997e-19 $X=2.135 $Y=1.625
r42 14 17 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.135 $Y=1.625
+ $X2=2.135 $Y2=1.79
r43 14 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.135 $Y=1.625
+ $X2=2.135 $Y2=1.46
r44 10 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.135
+ $Y=1.625 $X2=2.135 $Y2=1.625
r45 9 10 15.8897 $w=3.28e-07 $l=4.55e-07 $layer=LI1_cond $X=1.68 $Y=1.625
+ $X2=2.135 $Y2=1.625
r46 7 16 520.457 $w=1.5e-07 $l=1.015e-06 $layer=POLY_cond $X=2.155 $Y=0.445
+ $X2=2.155 $Y2=1.46
r47 3 17 183.856 $w=2.5e-07 $l=7.4e-07 $layer=POLY_cond $X=2.165 $Y=2.53
+ $X2=2.165 $Y2=1.79
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSTP_LP%SCD 1 3 8 12 14 15 19 21
r50 19 22 63.0283 $w=6.3e-07 $l=5.05e-07 $layer=POLY_cond $X=3.375 $Y=1.325
+ $X2=3.375 $Y2=1.83
r51 19 21 50.3829 $w=6.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.375 $Y=1.325
+ $X2=3.375 $Y2=1.16
r52 14 15 13.3251 $w=3.18e-07 $l=3.7e-07 $layer=LI1_cond $X=3.525 $Y=1.295
+ $X2=3.525 $Y2=1.665
r53 14 19 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.525
+ $Y=1.325 $X2=3.525 $Y2=1.325
r54 10 12 82.0426 $w=1.5e-07 $l=1.6e-07 $layer=POLY_cond $X=2.975 $Y=0.805
+ $X2=3.135 $Y2=0.805
r55 8 22 173.918 $w=2.5e-07 $l=7e-07 $layer=POLY_cond $X=3.185 $Y=2.53 $X2=3.185
+ $Y2=1.83
r56 4 12 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.135 $Y=0.88
+ $X2=3.135 $Y2=0.805
r57 4 21 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=3.135 $Y=0.88
+ $X2=3.135 $Y2=1.16
r58 1 10 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.975 $Y=0.73
+ $X2=2.975 $Y2=0.805
r59 1 3 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.975 $Y=0.73 $X2=2.975
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSTP_LP%CLK 3 6 9 13 16 17 20
c53 9 0 4.93603e-20 $X=4.275 $Y=2.545
c54 3 0 3.76099e-20 $X=4.11 $Y=0.75
r55 20 22 31.0702 $w=4.35e-07 $l=1.65e-07 $layer=POLY_cond $X=4.252 $Y=1.675
+ $X2=4.252 $Y2=1.84
r56 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.305
+ $Y=1.675 $X2=4.305 $Y2=1.675
r57 17 21 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=4.56 $Y=1.675
+ $X2=4.305 $Y2=1.675
r58 9 22 175.16 $w=2.5e-07 $l=7.05e-07 $layer=POLY_cond $X=4.275 $Y=2.545
+ $X2=4.275 $Y2=1.84
r59 6 20 6.64828 $w=4.35e-07 $l=5.2e-08 $layer=POLY_cond $X=4.252 $Y=1.623
+ $X2=4.252 $Y2=1.675
r60 6 16 39.3783 $w=4.35e-07 $l=3.08e-07 $layer=POLY_cond $X=4.252 $Y=1.623
+ $X2=4.252 $Y2=1.315
r61 1 16 24.5823 $w=4.35e-07 $l=1.5e-07 $layer=POLY_cond $X=4.305 $Y=1.165
+ $X2=4.305 $Y2=1.315
r62 1 13 212.798 $w=1.5e-07 $l=4.15e-07 $layer=POLY_cond $X=4.5 $Y=1.165 $X2=4.5
+ $Y2=0.75
r63 1 3 212.798 $w=1.5e-07 $l=4.15e-07 $layer=POLY_cond $X=4.11 $Y=1.165
+ $X2=4.11 $Y2=0.75
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSTP_LP%A_986_409# 1 2 9 13 17 21 25 27 28 32 35
+ 36 38 41 42 43 45 46 51 53 54 57 59 64 65 70
c206 65 0 1.43583e-19 $X=10.18 $Y=1.465
c207 64 0 1.422e-19 $X=10.015 $Y=1.465
c208 54 0 1.76636e-19 $X=5.875 $Y=1.3
c209 36 0 6.73817e-20 $X=6.73 $Y=1.465
c210 28 0 4.93603e-20 $X=5.235 $Y=2.98
r211 70 82 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=10.915 $Y=1.77
+ $X2=10.915 $Y2=1.935
r212 69 70 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.915
+ $Y=1.77 $X2=10.915 $Y2=1.77
r213 64 78 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=10.015 $Y=1.465
+ $X2=10.015 $Y2=1.3
r214 63 65 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=10.015 $Y=1.465
+ $X2=10.18 $Y2=1.465
r215 63 64 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.015
+ $Y=1.465 $X2=10.015 $Y2=1.465
r216 60 63 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=9.935 $Y=1.465
+ $X2=10.015 $Y2=1.465
r217 57 74 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.83 $Y=1.675
+ $X2=5.83 $Y2=1.84
r218 56 58 9.45624 $w=4.88e-07 $l=1.65e-07 $layer=LI1_cond $X=5.875 $Y=1.675
+ $X2=5.875 $Y2=1.84
r219 56 57 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.83
+ $Y=1.675 $X2=5.83 $Y2=1.675
r220 53 56 5.12605 $w=4.88e-07 $l=2.1e-07 $layer=LI1_cond $X=5.875 $Y=1.465
+ $X2=5.875 $Y2=1.675
r221 53 54 9.45624 $w=4.88e-07 $l=1.65e-07 $layer=LI1_cond $X=5.875 $Y=1.465
+ $X2=5.875 $Y2=1.3
r222 49 51 6.63049 $w=3.63e-07 $l=2.1e-07 $layer=LI1_cond $X=5.505 $Y=0.797
+ $X2=5.715 $Y2=0.797
r223 46 69 8.50163 $w=3.03e-07 $l=2.25e-07 $layer=LI1_cond $X=10.902 $Y=1.545
+ $X2=10.902 $Y2=1.77
r224 46 65 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=10.75 $Y=1.545
+ $X2=10.18 $Y2=1.545
r225 44 60 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.935 $Y=1.63
+ $X2=9.935 $Y2=1.465
r226 44 45 57.0856 $w=1.68e-07 $l=8.75e-07 $layer=LI1_cond $X=9.935 $Y=1.63
+ $X2=9.935 $Y2=2.505
r227 42 45 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=9.85 $Y=2.59
+ $X2=9.935 $Y2=2.505
r228 42 43 187.241 $w=1.68e-07 $l=2.87e-06 $layer=LI1_cond $X=9.85 $Y=2.59
+ $X2=6.98 $Y2=2.59
r229 40 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.895 $Y=2.675
+ $X2=6.98 $Y2=2.59
r230 40 41 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=6.895 $Y=2.675
+ $X2=6.895 $Y2=2.895
r231 39 59 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.12 $Y=2.98
+ $X2=6.035 $Y2=2.98
r232 38 41 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.81 $Y=2.98
+ $X2=6.895 $Y2=2.895
r233 38 39 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=6.81 $Y=2.98
+ $X2=6.12 $Y2=2.98
r234 36 76 16.6207 $w=3.19e-07 $l=1.1e-07 $layer=POLY_cond $X=6.73 $Y=1.465
+ $X2=6.84 $Y2=1.465
r235 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.73
+ $Y=1.465 $X2=6.73 $Y2=1.465
r236 33 53 3.05139 $w=3.3e-07 $l=2.45e-07 $layer=LI1_cond $X=6.12 $Y=1.465
+ $X2=5.875 $Y2=1.465
r237 33 35 21.3027 $w=3.28e-07 $l=6.1e-07 $layer=LI1_cond $X=6.12 $Y=1.465
+ $X2=6.73 $Y2=1.465
r238 32 59 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.035 $Y=2.895
+ $X2=6.035 $Y2=2.98
r239 32 58 68.8289 $w=1.68e-07 $l=1.055e-06 $layer=LI1_cond $X=6.035 $Y=2.895
+ $X2=6.035 $Y2=1.84
r240 29 51 5.2253 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=5.715 $Y=0.98
+ $X2=5.715 $Y2=0.797
r241 29 54 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=5.715 $Y=0.98
+ $X2=5.715 $Y2=1.3
r242 27 59 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.95 $Y=2.98
+ $X2=6.035 $Y2=2.98
r243 27 28 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=5.95 $Y=2.98
+ $X2=5.235 $Y2=2.98
r244 23 28 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.07 $Y=2.895
+ $X2=5.235 $Y2=2.98
r245 23 25 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=5.07 $Y=2.895
+ $X2=5.07 $Y2=2.535
r246 21 82 163.979 $w=2.5e-07 $l=6.6e-07 $layer=POLY_cond $X=10.905 $Y=2.595
+ $X2=10.905 $Y2=1.935
r247 17 78 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=9.955 $Y=0.835
+ $X2=9.955 $Y2=1.3
r248 11 76 20.418 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.84 $Y=1.3
+ $X2=6.84 $Y2=1.465
r249 11 13 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=6.84 $Y=1.3
+ $X2=6.84 $Y2=0.835
r250 9 74 187.582 $w=2.5e-07 $l=7.55e-07 $layer=POLY_cond $X=5.87 $Y=2.595
+ $X2=5.87 $Y2=1.84
r251 2 25 300 $w=1.7e-07 $l=5.55608e-07 $layer=licon1_PDIFF $count=2 $X=4.93
+ $Y=2.045 $X2=5.07 $Y2=2.535
r252 1 49 182 $w=1.7e-07 $l=3.17372e-07 $layer=licon1_NDIFF $count=1 $X=5.365
+ $Y=0.54 $X2=5.505 $Y2=0.795
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSTP_LP%A_1425_99# 1 2 9 11 13 15 16 17 19 21 24
+ 31
c76 17 0 7.21954e-20 $X=8.095 $Y=1.3
c77 13 0 1.23194e-19 $X=7.26 $Y=2.595
c78 11 0 5.62448e-20 $X=7.26 $Y=1.885
c79 9 0 8.63956e-20 $X=7.2 $Y=0.835
r80 28 31 5.5817 $w=4.48e-07 $l=2.1e-07 $layer=LI1_cond $X=8.18 $Y=0.84 $X2=8.39
+ $Y2=0.84
r81 26 27 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.59
+ $Y=1.38 $X2=7.59 $Y2=1.38
r82 23 28 6.50032 $w=1.7e-07 $l=2.25e-07 $layer=LI1_cond $X=8.18 $Y=1.065
+ $X2=8.18 $Y2=0.84
r83 23 24 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=8.18 $Y=1.065
+ $X2=8.18 $Y2=1.215
r84 19 21 30.8855 $w=2.48e-07 $l=6.7e-07 $layer=LI1_cond $X=7.755 $Y=2.2
+ $X2=8.425 $Y2=2.2
r85 18 26 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.755 $Y=1.3
+ $X2=7.59 $Y2=1.3
r86 17 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.095 $Y=1.3
+ $X2=8.18 $Y2=1.215
r87 17 18 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=8.095 $Y=1.3
+ $X2=7.755 $Y2=1.3
r88 16 19 6.98653 $w=2.5e-07 $l=2.18746e-07 $layer=LI1_cond $X=7.59 $Y=2.075
+ $X2=7.755 $Y2=2.2
r89 15 26 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.59 $Y=1.385 $X2=7.59
+ $Y2=1.3
r90 15 16 24.0965 $w=3.28e-07 $l=6.9e-07 $layer=LI1_cond $X=7.59 $Y=1.385
+ $X2=7.59 $Y2=2.075
r91 11 27 56.9292 $w=6.22e-07 $l=5.88154e-07 $layer=POLY_cond $X=7.26 $Y=1.885
+ $X2=7.44 $Y2=1.38
r92 11 13 176.402 $w=2.5e-07 $l=7.1e-07 $layer=POLY_cond $X=7.26 $Y=1.885
+ $X2=7.26 $Y2=2.595
r93 7 27 45.1746 $w=6.22e-07 $l=3.11769e-07 $layer=POLY_cond $X=7.2 $Y=1.215
+ $X2=7.44 $Y2=1.38
r94 7 9 194.851 $w=1.5e-07 $l=3.8e-07 $layer=POLY_cond $X=7.2 $Y=1.215 $X2=7.2
+ $Y2=0.835
r95 2 21 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=8.285
+ $Y=2.095 $X2=8.425 $Y2=2.24
r96 1 31 182 $w=1.7e-07 $l=2.78209e-07 $layer=licon1_NDIFF $count=1 $X=8.245
+ $Y=0.625 $X2=8.39 $Y2=0.84
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSTP_LP%A_1199_419# 1 2 9 13 14 17 21 25 29 30 33
+ 35 36 37 40 41 44 45 46 47 50 53 55 56 57 61 65 70 71 74
c186 71 0 1.43583e-19 $X=9.475 $Y=1.41
c187 70 0 1.96053e-19 $X=9.475 $Y=1.41
c188 61 0 8.63956e-20 $X=6.56 $Y=0.835
c189 57 0 5.62448e-20 $X=8.905 $Y=1.33
c190 56 0 1.99585e-19 $X=9.31 $Y=1.33
c191 50 0 2.901e-19 $X=8.16 $Y=1.73
c192 36 0 6.73817e-20 $X=6.63 $Y=2.16
c193 30 0 2.94985e-20 $X=9.475 $Y=1.915
r194 70 71 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=9.475
+ $Y=1.41 $X2=9.475 $Y2=1.41
r195 66 68 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=8.53 $Y=1.33
+ $X2=8.82 $Y2=1.33
r196 61 63 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=6.56 $Y=0.835
+ $X2=6.56 $Y2=0.965
r197 57 68 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=8.905 $Y=1.33
+ $X2=8.82 $Y2=1.33
r198 56 70 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.31 $Y=1.33
+ $X2=9.475 $Y2=1.33
r199 56 57 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=9.31 $Y=1.33
+ $X2=8.905 $Y2=1.33
r200 55 68 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.82 $Y=1.245
+ $X2=8.82 $Y2=1.33
r201 54 55 52.8449 $w=1.68e-07 $l=8.1e-07 $layer=LI1_cond $X=8.82 $Y=0.435
+ $X2=8.82 $Y2=1.245
r202 52 66 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.53 $Y=1.415
+ $X2=8.53 $Y2=1.33
r203 52 53 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=8.53 $Y=1.415
+ $X2=8.53 $Y2=1.565
r204 50 74 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.16 $Y=1.73
+ $X2=8.16 $Y2=1.565
r205 49 50 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.16
+ $Y=1.73 $X2=8.16 $Y2=1.73
r206 47 53 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=8.445 $Y=1.73
+ $X2=8.53 $Y2=1.565
r207 47 49 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=8.445 $Y=1.73
+ $X2=8.16 $Y2=1.73
r208 45 54 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.735 $Y=0.35
+ $X2=8.82 $Y2=0.435
r209 45 46 53.4973 $w=1.68e-07 $l=8.2e-07 $layer=LI1_cond $X=8.735 $Y=0.35
+ $X2=7.915 $Y2=0.35
r210 43 46 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.83 $Y=0.435
+ $X2=7.915 $Y2=0.35
r211 43 44 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=7.83 $Y=0.435
+ $X2=7.83 $Y2=0.865
r212 42 65 4.81226 $w=1.85e-07 $l=9.21954e-08 $layer=LI1_cond $X=7.245 $Y=0.95
+ $X2=7.16 $Y2=0.965
r213 41 44 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.745 $Y=0.95
+ $X2=7.83 $Y2=0.865
r214 41 42 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=7.745 $Y=0.95
+ $X2=7.245 $Y2=0.95
r215 39 65 1.64875 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=7.16 $Y=1.065 $X2=7.16
+ $Y2=0.965
r216 39 40 65.8931 $w=1.68e-07 $l=1.01e-06 $layer=LI1_cond $X=7.16 $Y=1.065
+ $X2=7.16 $Y2=2.075
r217 38 63 3.66692 $w=2e-07 $l=1.65e-07 $layer=LI1_cond $X=6.725 $Y=0.965
+ $X2=6.56 $Y2=0.965
r218 37 65 4.81226 $w=1.85e-07 $l=8.5e-08 $layer=LI1_cond $X=7.075 $Y=0.965
+ $X2=7.16 $Y2=0.965
r219 37 38 19.4091 $w=1.98e-07 $l=3.5e-07 $layer=LI1_cond $X=7.075 $Y=0.965
+ $X2=6.725 $Y2=0.965
r220 35 40 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.075 $Y=2.16
+ $X2=7.16 $Y2=2.075
r221 35 36 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=7.075 $Y=2.16
+ $X2=6.63 $Y2=2.16
r222 31 36 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.465 $Y=2.245
+ $X2=6.63 $Y2=2.16
r223 31 33 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=6.465 $Y=2.245
+ $X2=6.465 $Y2=2.395
r224 29 71 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=9.475 $Y=1.75
+ $X2=9.475 $Y2=1.41
r225 29 30 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=9.475 $Y=1.75
+ $X2=9.475 $Y2=1.915
r226 28 71 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=9.475 $Y=1.245
+ $X2=9.475 $Y2=1.41
r227 25 28 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=9.565 $Y=0.835
+ $X2=9.565 $Y2=1.245
r228 21 30 168.948 $w=2.5e-07 $l=6.8e-07 $layer=POLY_cond $X=9.515 $Y=2.595
+ $X2=9.515 $Y2=1.915
r229 15 17 194.851 $w=1.5e-07 $l=3.8e-07 $layer=POLY_cond $X=8.605 $Y=1.215
+ $X2=8.605 $Y2=0.835
r230 13 15 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.53 $Y=1.29
+ $X2=8.605 $Y2=1.215
r231 13 14 105.117 $w=1.5e-07 $l=2.05e-07 $layer=POLY_cond $X=8.53 $Y=1.29
+ $X2=8.325 $Y2=1.29
r232 11 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.25 $Y=1.365
+ $X2=8.325 $Y2=1.29
r233 11 74 102.553 $w=1.5e-07 $l=2e-07 $layer=POLY_cond $X=8.25 $Y=1.365
+ $X2=8.25 $Y2=1.565
r234 7 50 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.16 $Y=1.895
+ $X2=8.16 $Y2=1.73
r235 7 9 173.918 $w=2.5e-07 $l=7e-07 $layer=POLY_cond $X=8.16 $Y=1.895 $X2=8.16
+ $Y2=2.595
r236 2 33 600 $w=1.7e-07 $l=6.01581e-07 $layer=licon1_PDIFF $count=1 $X=5.995
+ $Y=2.095 $X2=6.465 $Y2=2.395
r237 1 61 182 $w=1.7e-07 $l=2.95212e-07 $layer=licon1_NDIFF $count=1 $X=6.355
+ $Y=0.625 $X2=6.56 $Y2=0.835
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSTP_LP%SET_B 3 7 9 11 12 13 16 20 21 22 27 30 31
+ 36 37
c126 37 0 1.99585e-19 $X=8.995 $Y=1.77
c127 36 0 1.66906e-19 $X=8.935 $Y=1.77
c128 21 0 2.94985e-20 $X=12.095 $Y=2.035
c129 7 0 7.21954e-20 $X=8.995 $Y=0.835
r130 35 37 10.4917 $w=3.3e-07 $l=6e-08 $layer=POLY_cond $X=8.935 $Y=1.77
+ $X2=8.995 $Y2=1.77
r131 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.935
+ $Y=1.77 $X2=8.935 $Y2=1.77
r132 32 35 42.841 $w=3.3e-07 $l=2.45e-07 $layer=POLY_cond $X=8.69 $Y=1.77
+ $X2=8.935 $Y2=1.77
r133 31 46 21.1281 $w=3.28e-07 $l=6.05e-07 $layer=LI1_cond $X=12.265 $Y=1.43
+ $X2=12.265 $Y2=2.035
r134 30 31 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=12.265
+ $Y=1.43 $X2=12.265 $Y2=1.43
r135 27 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.24 $Y=2.035
+ $X2=12.24 $Y2=2.035
r136 25 36 10.013 $w=3.03e-07 $l=2.65e-07 $layer=LI1_cond $X=8.947 $Y=2.035
+ $X2=8.947 $Y2=1.77
r137 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=2.035
+ $X2=8.88 $Y2=2.035
r138 22 24 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=9.025 $Y=2.035
+ $X2=8.88 $Y2=2.035
r139 21 27 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=12.095 $Y=2.035
+ $X2=12.24 $Y2=2.035
r140 21 22 3.7995 $w=1.4e-07 $l=3.07e-06 $layer=MET1_cond $X=12.095 $Y=2.035
+ $X2=9.025 $Y2=2.035
r141 19 30 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=12.265 $Y=1.77
+ $X2=12.265 $Y2=1.43
r142 19 20 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=12.265 $Y=1.77
+ $X2=12.265 $Y2=1.935
r143 18 30 79.5619 $w=3.3e-07 $l=4.55e-07 $layer=POLY_cond $X=12.265 $Y=0.975
+ $X2=12.265 $Y2=1.43
r144 16 20 163.979 $w=2.5e-07 $l=6.6e-07 $layer=POLY_cond $X=12.225 $Y=2.595
+ $X2=12.225 $Y2=1.935
r145 12 18 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=12.1 $Y=0.9
+ $X2=12.265 $Y2=0.975
r146 12 13 358.936 $w=1.5e-07 $l=7e-07 $layer=POLY_cond $X=12.1 $Y=0.9 $X2=11.4
+ $Y2=0.9
r147 9 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=11.325 $Y=0.825
+ $X2=11.4 $Y2=0.9
r148 9 11 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=11.325 $Y=0.825
+ $X2=11.325 $Y2=0.54
r149 5 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.995 $Y=1.605
+ $X2=8.995 $Y2=1.77
r150 5 7 394.83 $w=1.5e-07 $l=7.7e-07 $layer=POLY_cond $X=8.995 $Y=1.605
+ $X2=8.995 $Y2=0.835
r151 1 32 9.34494 $w=2.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.69 $Y=1.935
+ $X2=8.69 $Y2=1.77
r152 1 3 163.979 $w=2.5e-07 $l=6.6e-07 $layer=POLY_cond $X=8.69 $Y=1.935
+ $X2=8.69 $Y2=2.595
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSTP_LP%A_750_108# 1 2 9 13 16 17 21 23 28 30 31
+ 32 33 34 35 37 38 40 41 42 44 48 49 50 51 54 60 63 64 68 69 72 75
c208 54 0 1.84917e-19 $X=10.545 $Y=1.195
c209 49 0 1.98095e-19 $X=4.93 $Y=1.195
c210 42 0 5.38522e-20 $X=10.13 $Y=1.945
c211 16 0 1.76636e-19 $X=4.93 $Y=1.555
r212 76 78 21.8577 $w=3.3e-07 $l=1.25e-07 $layer=POLY_cond $X=4.805 $Y=1.72
+ $X2=4.93 $Y2=1.72
r213 72 74 9.71523 $w=2.48e-07 $l=1.85e-07 $layer=LI1_cond $X=3.935 $Y=0.795
+ $X2=3.935 $Y2=0.98
r214 69 78 5.24584 $w=3.3e-07 $l=3e-08 $layer=POLY_cond $X=4.96 $Y=1.72 $X2=4.93
+ $Y2=1.72
r215 68 69 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.96
+ $Y=1.72 $X2=4.96 $Y2=1.72
r216 66 68 12.5721 $w=2.73e-07 $l=3e-07 $layer=LI1_cond $X=4.962 $Y=2.02
+ $X2=4.962 $Y2=1.72
r217 65 75 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.175 $Y=2.105
+ $X2=4.01 $Y2=2.105
r218 64 66 7.32204 $w=1.7e-07 $l=1.74396e-07 $layer=LI1_cond $X=4.825 $Y=2.105
+ $X2=4.962 $Y2=2.02
r219 64 65 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=4.825 $Y=2.105
+ $X2=4.175 $Y2=2.105
r220 63 75 3.70735 $w=2.5e-07 $l=1.11018e-07 $layer=LI1_cond $X=3.95 $Y=2.02
+ $X2=4.01 $Y2=2.105
r221 63 74 67.8503 $w=1.68e-07 $l=1.04e-06 $layer=LI1_cond $X=3.95 $Y=2.02
+ $X2=3.95 $Y2=0.98
r222 58 75 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.01 $Y=2.19
+ $X2=4.01 $Y2=2.105
r223 58 60 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=4.01 $Y=2.19
+ $X2=4.01 $Y2=2.9
r224 52 54 41.0213 $w=1.5e-07 $l=8e-08 $layer=POLY_cond $X=10.465 $Y=1.195
+ $X2=10.545 $Y2=1.195
r225 46 54 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=10.545 $Y=1.12
+ $X2=10.545 $Y2=1.195
r226 46 48 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=10.545 $Y=1.12
+ $X2=10.545 $Y2=0.54
r227 45 48 146.138 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=10.545 $Y=0.255
+ $X2=10.545 $Y2=0.54
r228 43 52 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=10.465 $Y=1.27
+ $X2=10.465 $Y2=1.195
r229 43 44 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=10.465 $Y=1.27
+ $X2=10.465 $Y2=1.87
r230 41 44 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=10.39 $Y=1.945
+ $X2=10.465 $Y2=1.87
r231 41 42 133.319 $w=1.5e-07 $l=2.6e-07 $layer=POLY_cond $X=10.39 $Y=1.945
+ $X2=10.13 $Y2=1.945
r232 38 42 29.1797 $w=1.5e-07 $l=1.58114e-07 $layer=POLY_cond $X=10.005 $Y=2.02
+ $X2=10.13 $Y2=1.945
r233 38 40 110.86 $w=2.5e-07 $l=5.75e-07 $layer=POLY_cond $X=10.005 $Y=2.02
+ $X2=10.005 $Y2=2.595
r234 35 37 110.86 $w=2.5e-07 $l=5.75e-07 $layer=POLY_cond $X=6.73 $Y=2.02
+ $X2=6.73 $Y2=2.595
r235 33 35 29.1797 $w=1.5e-07 $l=1.58114e-07 $layer=POLY_cond $X=6.605 $Y=1.945
+ $X2=6.73 $Y2=2.02
r236 33 34 128.191 $w=1.5e-07 $l=2.5e-07 $layer=POLY_cond $X=6.605 $Y=1.945
+ $X2=6.355 $Y2=1.945
r237 31 45 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=10.47 $Y=0.18
+ $X2=10.545 $Y2=0.255
r238 31 32 2110.03 $w=1.5e-07 $l=4.115e-06 $layer=POLY_cond $X=10.47 $Y=0.18
+ $X2=6.355 $Y2=0.18
r239 30 34 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.28 $Y=1.87
+ $X2=6.355 $Y2=1.945
r240 29 51 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.28 $Y=1.27
+ $X2=6.28 $Y2=1.195
r241 29 30 307.66 $w=1.5e-07 $l=6e-07 $layer=POLY_cond $X=6.28 $Y=1.27 $X2=6.28
+ $Y2=1.87
r242 26 51 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.28 $Y=1.12
+ $X2=6.28 $Y2=1.195
r243 26 28 146.138 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=6.28 $Y=1.12
+ $X2=6.28 $Y2=0.835
r244 25 32 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=6.28 $Y=0.255
+ $X2=6.355 $Y2=0.18
r245 25 28 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=6.28 $Y=0.255
+ $X2=6.28 $Y2=0.835
r246 24 50 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.365 $Y=1.195
+ $X2=5.29 $Y2=1.195
r247 23 51 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.205 $Y=1.195
+ $X2=6.28 $Y2=1.195
r248 23 24 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=6.205 $Y=1.195
+ $X2=5.365 $Y2=1.195
r249 19 50 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.29 $Y=1.12
+ $X2=5.29 $Y2=1.195
r250 19 21 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=5.29 $Y=1.12
+ $X2=5.29 $Y2=0.75
r251 18 49 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.005 $Y=1.195
+ $X2=4.93 $Y2=1.195
r252 17 50 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.215 $Y=1.195
+ $X2=5.29 $Y2=1.195
r253 17 18 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=5.215 $Y=1.195
+ $X2=5.005 $Y2=1.195
r254 16 78 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.93 $Y=1.555
+ $X2=4.93 $Y2=1.72
r255 15 49 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.93 $Y=1.27
+ $X2=4.93 $Y2=1.195
r256 15 16 146.138 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=4.93 $Y=1.27
+ $X2=4.93 $Y2=1.555
r257 11 49 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.93 $Y=1.12
+ $X2=4.93 $Y2=1.195
r258 11 13 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=4.93 $Y=1.12
+ $X2=4.93 $Y2=0.75
r259 7 76 9.34494 $w=2.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.805 $Y=1.885
+ $X2=4.805 $Y2=1.72
r260 7 9 163.979 $w=2.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.805 $Y=1.885
+ $X2=4.805 $Y2=2.545
r261 2 60 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=3.865
+ $Y=2.045 $X2=4.01 $Y2=2.9
r262 2 58 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=3.865
+ $Y=2.045 $X2=4.01 $Y2=2.19
r263 1 72 182 $w=1.7e-07 $l=3.19374e-07 $layer=licon1_NDIFF $count=1 $X=3.75
+ $Y=0.54 $X2=3.895 $Y2=0.795
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSTP_LP%A_2172_40# 1 2 9 11 12 15 19 22 23 26 28
+ 30 35
c83 35 0 1.32475e-20 $X=11.605 $Y=1.29
r84 28 30 36.6477 $w=2.48e-07 $l=7.95e-07 $layer=LI1_cond $X=13.01 $Y=1.085
+ $X2=13.01 $Y2=1.88
r85 24 28 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=12.63 $Y=1 $X2=13.01
+ $Y2=1
r86 24 26 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=12.63 $Y=0.915
+ $X2=12.63 $Y2=0.495
r87 22 24 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=12.465 $Y=1
+ $X2=12.63 $Y2=1
r88 22 23 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=12.465 $Y=1
+ $X2=11.89 $Y2=1
r89 20 38 64.545 $w=5.7e-07 $l=5.05e-07 $layer=POLY_cond $X=11.605 $Y=1.38
+ $X2=11.605 $Y2=1.885
r90 20 35 8.44783 $w=5.7e-07 $l=9e-08 $layer=POLY_cond $X=11.605 $Y=1.38
+ $X2=11.605 $Y2=1.29
r91 19 20 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=11.725
+ $Y=1.38 $X2=11.725 $Y2=1.38
r92 17 23 7.55824 $w=1.7e-07 $l=1.90825e-07 $layer=LI1_cond $X=11.737 $Y=1.085
+ $X2=11.89 $Y2=1
r93 17 19 11.1466 $w=3.03e-07 $l=2.95e-07 $layer=LI1_cond $X=11.737 $Y=1.085
+ $X2=11.737 $Y2=1.38
r94 15 38 176.402 $w=2.5e-07 $l=7.1e-07 $layer=POLY_cond $X=11.445 $Y=2.595
+ $X2=11.445 $Y2=1.885
r95 11 35 34.7497 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=11.32 $Y=1.29
+ $X2=11.605 $Y2=1.29
r96 11 12 158.957 $w=1.5e-07 $l=3.1e-07 $layer=POLY_cond $X=11.32 $Y=1.29
+ $X2=11.01 $Y2=1.29
r97 7 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=10.935 $Y=1.215
+ $X2=11.01 $Y2=1.29
r98 7 9 346.117 $w=1.5e-07 $l=6.75e-07 $layer=POLY_cond $X=10.935 $Y=1.215
+ $X2=10.935 $Y2=0.54
r99 2 30 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=12.905
+ $Y=1.735 $X2=13.05 $Y2=1.88
r100 1 26 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=12.485
+ $Y=0.285 $X2=12.63 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSTP_LP%A_2006_125# 1 2 3 10 12 13 14 15 17 20 22
+ 26 28 32 36 39 41 42 43 46 50 52 53 54 57 58 60 61 62 63 66 67 70 72 75 78
c181 57 0 1.84917e-19 $X=11.32 $Y=2.33
r182 72 74 6.11144 $w=3.28e-07 $l=1.75e-07 $layer=LI1_cond $X=10.405 $Y=2.24
+ $X2=10.405 $Y2=2.415
r183 70 78 86.1176 $w=1.68e-07 $l=1.32e-06 $layer=LI1_cond $X=13.4 $Y=2.895
+ $X2=13.4 $Y2=1.575
r184 66 67 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=13.48
+ $Y=1.07 $X2=13.48 $Y2=1.07
r185 64 78 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=13.48 $Y=1.41
+ $X2=13.48 $Y2=1.575
r186 64 66 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=13.48 $Y=1.41
+ $X2=13.48 $Y2=1.07
r187 62 70 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=13.315 $Y=2.98
+ $X2=13.4 $Y2=2.895
r188 62 63 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=13.315 $Y=2.98
+ $X2=12.655 $Y2=2.98
r189 61 63 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=12.49 $Y=2.895
+ $X2=12.655 $Y2=2.98
r190 60 77 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=12.49 $Y=2.5
+ $X2=12.49 $Y2=2.415
r191 60 61 13.7944 $w=3.28e-07 $l=3.95e-07 $layer=LI1_cond $X=12.49 $Y=2.5
+ $X2=12.49 $Y2=2.895
r192 59 75 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.405 $Y=2.415
+ $X2=11.32 $Y2=2.415
r193 58 77 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.325 $Y=2.415
+ $X2=12.49 $Y2=2.415
r194 58 59 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=12.325 $Y=2.415
+ $X2=11.405 $Y2=2.415
r195 57 75 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.32 $Y=2.33
+ $X2=11.32 $Y2=2.415
r196 56 57 81.2246 $w=1.68e-07 $l=1.245e-06 $layer=LI1_cond $X=11.32 $Y=1.085
+ $X2=11.32 $Y2=2.33
r197 55 74 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.57 $Y=2.415
+ $X2=10.405 $Y2=2.415
r198 54 75 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.235 $Y=2.415
+ $X2=11.32 $Y2=2.415
r199 54 55 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=11.235 $Y=2.415
+ $X2=10.57 $Y2=2.415
r200 52 56 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=11.235 $Y=1
+ $X2=11.32 $Y2=1.085
r201 52 53 45.9947 $w=1.68e-07 $l=7.05e-07 $layer=LI1_cond $X=11.235 $Y=1
+ $X2=10.53 $Y2=1
r202 48 74 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=10.405 $Y=2.5
+ $X2=10.405 $Y2=2.415
r203 48 50 13.969 $w=3.28e-07 $l=4e-07 $layer=LI1_cond $X=10.405 $Y=2.5
+ $X2=10.405 $Y2=2.9
r204 44 53 8.76165 $w=1.7e-07 $l=2.62076e-07 $layer=LI1_cond $X=10.307 $Y=0.915
+ $X2=10.53 $Y2=1
r205 44 46 11.3949 $w=4.43e-07 $l=4.4e-07 $layer=LI1_cond $X=10.307 $Y=0.915
+ $X2=10.307 $Y2=0.475
r206 40 67 43.3922 $w=4.55e-07 $l=3.55e-07 $layer=POLY_cond $X=13.417 $Y=1.425
+ $X2=13.417 $Y2=1.07
r207 40 41 9.56592 $w=3.52e-07 $l=7.5e-08 $layer=POLY_cond $X=13.417 $Y=1.425
+ $X2=13.417 $Y2=1.5
r208 38 67 11.612 $w=4.55e-07 $l=9.5e-08 $layer=POLY_cond $X=13.417 $Y=0.975
+ $X2=13.417 $Y2=1.07
r209 38 39 11.0167 $w=3.02e-07 $l=8.87412e-08 $layer=POLY_cond $X=13.417
+ $Y=0.975 $X2=13.387 $Y2=0.9
r210 34 43 15.9654 $w=2e-07 $l=8.44097e-08 $layer=POLY_cond $X=14.555 $Y=1.425
+ $X2=14.575 $Y2=1.5
r211 34 36 476.872 $w=1.5e-07 $l=9.3e-07 $layer=POLY_cond $X=14.555 $Y=1.425
+ $X2=14.555 $Y2=0.495
r212 30 43 15.9654 $w=2e-07 $l=7.5e-08 $layer=POLY_cond $X=14.575 $Y=1.575
+ $X2=14.575 $Y2=1.5
r213 30 32 197.521 $w=2.5e-07 $l=7.95e-07 $layer=POLY_cond $X=14.575 $Y=1.575
+ $X2=14.575 $Y2=2.37
r214 29 42 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=14.27 $Y=1.5
+ $X2=14.195 $Y2=1.5
r215 28 43 9.46703 $w=1.5e-07 $l=1.25e-07 $layer=POLY_cond $X=14.45 $Y=1.5
+ $X2=14.575 $Y2=1.5
r216 28 29 92.2979 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=14.45 $Y=1.5
+ $X2=14.27 $Y2=1.5
r217 24 42 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=14.195 $Y=1.425
+ $X2=14.195 $Y2=1.5
r218 24 26 476.872 $w=1.5e-07 $l=9.3e-07 $layer=POLY_cond $X=14.195 $Y=1.425
+ $X2=14.195 $Y2=0.495
r219 23 41 17.931 $w=1.5e-07 $l=2.28e-07 $layer=POLY_cond $X=13.645 $Y=1.5
+ $X2=13.417 $Y2=1.5
r220 22 42 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=14.12 $Y=1.5
+ $X2=14.195 $Y2=1.5
r221 22 23 243.564 $w=1.5e-07 $l=4.75e-07 $layer=POLY_cond $X=14.12 $Y=1.5
+ $X2=13.645 $Y2=1.5
r222 18 41 9.56592 $w=3.52e-07 $l=1.34365e-07 $layer=POLY_cond $X=13.315
+ $Y=1.575 $X2=13.417 $Y2=1.5
r223 18 20 163.979 $w=2.5e-07 $l=6.6e-07 $layer=POLY_cond $X=13.315 $Y=1.575
+ $X2=13.315 $Y2=2.235
r224 15 39 11.0167 $w=3.02e-07 $l=2.16273e-07 $layer=POLY_cond $X=13.205
+ $Y=0.825 $X2=13.387 $Y2=0.9
r225 15 17 106.04 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=13.205 $Y=0.825
+ $X2=13.205 $Y2=0.495
r226 13 39 15.6242 $w=1.5e-07 $l=2.57e-07 $layer=POLY_cond $X=13.13 $Y=0.9
+ $X2=13.387 $Y2=0.9
r227 13 14 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=13.13 $Y=0.9
+ $X2=12.92 $Y2=0.9
r228 10 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=12.845 $Y=0.825
+ $X2=12.92 $Y2=0.9
r229 10 12 106.04 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=12.845 $Y=0.825
+ $X2=12.845 $Y2=0.495
r230 3 77 300 $w=1.7e-07 $l=4.64758e-07 $layer=licon1_PDIFF $count=2 $X=12.35
+ $Y=2.095 $X2=12.49 $Y2=2.495
r231 2 72 600 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=1 $X=10.13
+ $Y=2.095 $X2=10.405 $Y2=2.24
r232 2 50 600 $w=1.7e-07 $l=9.32416e-07 $layer=licon1_PDIFF $count=1 $X=10.13
+ $Y=2.095 $X2=10.405 $Y2=2.9
r233 1 46 91 $w=1.7e-07 $l=2.85307e-07 $layer=licon1_NDIFF $count=2 $X=10.03
+ $Y=0.625 $X2=10.25 $Y2=0.475
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSTP_LP%A_2767_57# 1 2 9 13 17 23 26 28 31 35 42
+ 44 46 47
c74 26 0 6.94276e-20 $X=15.075 $Y=1.66
r75 46 47 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=15.075
+ $Y=1.155 $X2=15.075 $Y2=1.155
r76 40 42 5.20034 $w=4.58e-07 $l=2e-07 $layer=LI1_cond $X=13.98 $Y=0.495
+ $X2=14.18 $Y2=0.495
r77 36 44 3.11956 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=14.475 $Y=1.075
+ $X2=14.285 $Y2=1.075
r78 35 46 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=14.91 $Y=1.075
+ $X2=15.075 $Y2=1.075
r79 35 36 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=14.91 $Y=1.075
+ $X2=14.475 $Y2=1.075
r80 31 33 21.5325 $w=3.78e-07 $l=7.1e-07 $layer=LI1_cond $X=14.285 $Y=2.015
+ $X2=14.285 $Y2=2.725
r81 29 44 3.40559 $w=2.75e-07 $l=8.5e-08 $layer=LI1_cond $X=14.285 $Y=1.16
+ $X2=14.285 $Y2=1.075
r82 29 31 25.93 $w=3.78e-07 $l=8.55e-07 $layer=LI1_cond $X=14.285 $Y=1.16
+ $X2=14.285 $Y2=2.015
r83 28 44 3.40559 $w=2.75e-07 $l=1.41244e-07 $layer=LI1_cond $X=14.18 $Y=0.99
+ $X2=14.285 $Y2=1.075
r84 27 42 6.6364 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=14.18 $Y=0.725
+ $X2=14.18 $Y2=0.495
r85 27 28 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=14.18 $Y=0.725
+ $X2=14.18 $Y2=0.99
r86 25 47 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=15.075 $Y=1.495
+ $X2=15.075 $Y2=1.155
r87 25 26 31.6748 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=15.075 $Y=1.495
+ $X2=15.075 $Y2=1.66
r88 22 47 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=15.075 $Y=1.14
+ $X2=15.075 $Y2=1.155
r89 22 23 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=15.075 $Y=1.065
+ $X2=15.345 $Y2=1.065
r90 19 22 46.1489 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=14.985 $Y=1.065
+ $X2=15.075 $Y2=1.065
r91 15 23 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=15.345 $Y=0.99
+ $X2=15.345 $Y2=1.065
r92 15 17 253.819 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=15.345 $Y=0.99
+ $X2=15.345 $Y2=0.495
r93 13 26 176.402 $w=2.5e-07 $l=7.1e-07 $layer=POLY_cond $X=15.105 $Y=2.37
+ $X2=15.105 $Y2=1.66
r94 7 19 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=14.985 $Y=0.99
+ $X2=14.985 $Y2=1.065
r95 7 9 253.819 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=14.985 $Y=0.99
+ $X2=14.985 $Y2=0.495
r96 2 33 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=14.165
+ $Y=1.87 $X2=14.31 $Y2=2.725
r97 2 31 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=14.165
+ $Y=1.87 $X2=14.31 $Y2=2.015
r98 1 40 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=13.835
+ $Y=0.285 $X2=13.98 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSTP_LP%VPWR 1 2 3 4 5 6 7 8 29 35 39 43 47 51 55
+ 59 64 65 67 68 69 78 85 90 95 103 113 114 117 120 123 126 129 132
r166 132 133 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=13.68 $Y=3.33
+ $X2=13.68 $Y2=3.33
r167 129 130 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.76 $Y=3.33
+ $X2=11.76 $Y2=3.33
r168 126 127 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r169 123 124 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r170 120 121 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r171 117 118 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r172 113 114 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=15.6 $Y=3.33
+ $X2=15.6 $Y2=3.33
r173 111 114 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=14.64 $Y=3.33
+ $X2=15.6 $Y2=3.33
r174 111 133 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=14.64 $Y=3.33
+ $X2=13.68 $Y2=3.33
r175 110 111 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=14.64 $Y=3.33
+ $X2=14.64 $Y2=3.33
r176 108 132 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=13.915 $Y=3.33
+ $X2=13.79 $Y2=3.33
r177 108 110 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=13.915 $Y=3.33
+ $X2=14.64 $Y2=3.33
r178 107 133 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=12.24 $Y=3.33
+ $X2=13.68 $Y2=3.33
r179 107 130 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=12.24 $Y=3.33
+ $X2=11.76 $Y2=3.33
r180 106 107 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=12.24 $Y=3.33
+ $X2=12.24 $Y2=3.33
r181 104 129 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.875 $Y=3.33
+ $X2=11.71 $Y2=3.33
r182 104 106 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=11.875 $Y=3.33
+ $X2=12.24 $Y2=3.33
r183 103 132 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=13.665 $Y=3.33
+ $X2=13.79 $Y2=3.33
r184 103 106 92.9679 $w=1.68e-07 $l=1.425e-06 $layer=LI1_cond $X=13.665 $Y=3.33
+ $X2=12.24 $Y2=3.33
r185 102 130 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=3.33
+ $X2=11.76 $Y2=3.33
r186 101 102 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=11.28 $Y=3.33
+ $X2=11.28 $Y2=3.33
r187 99 102 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=11.28 $Y2=3.33
r188 99 127 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=8.88 $Y2=3.33
r189 98 101 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=9.36 $Y=3.33
+ $X2=11.28 $Y2=3.33
r190 98 99 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r191 96 126 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.12 $Y=3.33
+ $X2=8.955 $Y2=3.33
r192 96 98 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=9.12 $Y=3.33
+ $X2=9.36 $Y2=3.33
r193 95 129 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.545 $Y=3.33
+ $X2=11.71 $Y2=3.33
r194 95 101 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=11.545 $Y=3.33
+ $X2=11.28 $Y2=3.33
r195 94 127 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=8.88 $Y2=3.33
r196 93 94 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r197 91 123 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.77 $Y=3.33
+ $X2=7.605 $Y2=3.33
r198 91 93 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=7.77 $Y=3.33
+ $X2=8.4 $Y2=3.33
r199 90 126 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.79 $Y=3.33
+ $X2=8.955 $Y2=3.33
r200 90 93 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=8.79 $Y=3.33
+ $X2=8.4 $Y2=3.33
r201 89 124 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=7.44 $Y2=3.33
r202 89 121 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=3.33
+ $X2=4.56 $Y2=3.33
r203 88 89 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r204 86 120 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.705 $Y=3.33
+ $X2=4.54 $Y2=3.33
r205 86 88 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=4.705 $Y=3.33
+ $X2=5.04 $Y2=3.33
r206 85 123 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.44 $Y=3.33
+ $X2=7.605 $Y2=3.33
r207 85 88 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=7.44 $Y=3.33
+ $X2=5.04 $Y2=3.33
r208 84 121 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r209 83 84 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r210 81 84 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=4.08 $Y2=3.33
r211 80 83 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=3.12 $Y=3.33
+ $X2=4.08 $Y2=3.33
r212 80 81 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r213 78 120 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.375 $Y=3.33
+ $X2=4.54 $Y2=3.33
r214 78 83 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=4.375 $Y=3.33
+ $X2=4.08 $Y2=3.33
r215 77 81 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r216 76 77 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r217 74 77 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r218 74 118 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r219 73 76 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r220 73 74 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r221 71 117 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.975 $Y=3.33
+ $X2=0.81 $Y2=3.33
r222 71 73 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=0.975 $Y=3.33
+ $X2=1.2 $Y2=3.33
r223 69 94 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=8.4 $Y2=3.33
r224 69 124 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=3.33
+ $X2=7.44 $Y2=3.33
r225 67 110 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=14.675 $Y=3.33
+ $X2=14.64 $Y2=3.33
r226 67 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=14.675 $Y=3.33
+ $X2=14.84 $Y2=3.33
r227 66 113 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=15.005 $Y=3.33
+ $X2=15.6 $Y2=3.33
r228 66 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=15.005 $Y=3.33
+ $X2=14.84 $Y2=3.33
r229 64 76 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=2.755 $Y=3.33
+ $X2=2.64 $Y2=3.33
r230 64 65 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.755 $Y=3.33
+ $X2=2.92 $Y2=3.33
r231 63 80 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=3.085 $Y=3.33
+ $X2=3.12 $Y2=3.33
r232 63 65 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.085 $Y=3.33
+ $X2=2.92 $Y2=3.33
r233 59 62 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=14.84 $Y=2.015
+ $X2=14.84 $Y2=2.725
r234 57 68 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=14.84 $Y=3.245
+ $X2=14.84 $Y2=3.33
r235 57 62 18.1597 $w=3.28e-07 $l=5.2e-07 $layer=LI1_cond $X=14.84 $Y=3.245
+ $X2=14.84 $Y2=2.725
r236 53 132 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=13.79 $Y=3.245
+ $X2=13.79 $Y2=3.33
r237 53 55 61.0795 $w=2.48e-07 $l=1.325e-06 $layer=LI1_cond $X=13.79 $Y=3.245
+ $X2=13.79 $Y2=1.92
r238 49 129 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=11.71 $Y=3.245
+ $X2=11.71 $Y2=3.33
r239 49 51 12.2229 $w=3.28e-07 $l=3.5e-07 $layer=LI1_cond $X=11.71 $Y=3.245
+ $X2=11.71 $Y2=2.895
r240 45 126 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.955 $Y=3.245
+ $X2=8.955 $Y2=3.33
r241 45 47 10.4768 $w=3.28e-07 $l=3e-07 $layer=LI1_cond $X=8.955 $Y=3.245
+ $X2=8.955 $Y2=2.945
r242 41 123 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.605 $Y=3.245
+ $X2=7.605 $Y2=3.33
r243 41 43 7.85757 $w=3.28e-07 $l=2.25e-07 $layer=LI1_cond $X=7.605 $Y=3.245
+ $X2=7.605 $Y2=3.02
r244 37 120 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.54 $Y=3.245
+ $X2=4.54 $Y2=3.33
r245 37 39 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=4.54 $Y=3.245
+ $X2=4.54 $Y2=2.535
r246 33 65 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.92 $Y=3.245
+ $X2=2.92 $Y2=3.33
r247 33 35 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=2.92 $Y=3.245
+ $X2=2.92 $Y2=2.86
r248 29 32 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=0.81 $Y=2.19
+ $X2=0.81 $Y2=2.9
r249 27 117 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.81 $Y=3.245
+ $X2=0.81 $Y2=3.33
r250 27 32 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=0.81 $Y=3.245
+ $X2=0.81 $Y2=2.9
r251 8 62 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=14.7
+ $Y=1.87 $X2=14.84 $Y2=2.725
r252 8 59 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=14.7
+ $Y=1.87 $X2=14.84 $Y2=2.015
r253 7 55 300 $w=1.7e-07 $l=3.91727e-07 $layer=licon1_PDIFF $count=2 $X=13.44
+ $Y=1.735 $X2=13.75 $Y2=1.92
r254 6 51 600 $w=1.7e-07 $l=8.67179e-07 $layer=licon1_PDIFF $count=1 $X=11.57
+ $Y=2.095 $X2=11.71 $Y2=2.895
r255 5 47 600 $w=1.7e-07 $l=9.17333e-07 $layer=licon1_PDIFF $count=1 $X=8.815
+ $Y=2.095 $X2=8.955 $Y2=2.945
r256 4 43 600 $w=1.7e-07 $l=1.02914e-06 $layer=licon1_PDIFF $count=1 $X=7.385
+ $Y=2.095 $X2=7.605 $Y2=3.02
r257 3 39 300 $w=1.7e-07 $l=5.55608e-07 $layer=licon1_PDIFF $count=2 $X=4.4
+ $Y=2.045 $X2=4.54 $Y2=2.535
r258 2 35 600 $w=1.7e-07 $l=8.97274e-07 $layer=licon1_PDIFF $count=1 $X=2.78
+ $Y=2.03 $X2=2.92 $Y2=2.86
r259 1 32 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=0.67
+ $Y=2.045 $X2=0.81 $Y2=2.9
r260 1 29 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.67
+ $Y=2.045 $X2=0.81 $Y2=2.19
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSTP_LP%A_245_406# 1 2 9 13 14 16 17 18 21 25 27
r60 23 27 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.49 $Y=2.49 $X2=3.49
+ $Y2=2.405
r61 23 25 1.84391 $w=2.48e-07 $l=4e-08 $layer=LI1_cond $X=3.49 $Y=2.49 $X2=3.49
+ $Y2=2.53
r62 19 27 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.49 $Y=2.32 $X2=3.49
+ $Y2=2.405
r63 19 21 6.68417 $w=2.48e-07 $l=1.45e-07 $layer=LI1_cond $X=3.49 $Y=2.32
+ $X2=3.49 $Y2=2.175
r64 17 27 2.76166 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.365 $Y=2.405
+ $X2=3.49 $Y2=2.405
r65 17 18 61.9786 $w=1.68e-07 $l=9.5e-07 $layer=LI1_cond $X=3.365 $Y=2.405
+ $X2=2.415 $Y2=2.405
r66 15 18 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.33 $Y=2.49
+ $X2=2.415 $Y2=2.405
r67 15 16 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=2.33 $Y=2.49
+ $X2=2.33 $Y2=2.895
r68 13 16 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.245 $Y=2.98
+ $X2=2.33 $Y2=2.895
r69 13 14 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=2.245 $Y=2.98
+ $X2=1.535 $Y2=2.98
r70 9 12 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=1.37 $Y=2.175 $X2=1.37
+ $Y2=2.885
r71 7 14 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.37 $Y=2.895
+ $X2=1.535 $Y2=2.98
r72 7 12 0.349225 $w=3.28e-07 $l=1e-08 $layer=LI1_cond $X=1.37 $Y=2.895 $X2=1.37
+ $Y2=2.885
r73 2 25 300 $w=1.7e-07 $l=5.65685e-07 $layer=licon1_PDIFF $count=2 $X=3.31
+ $Y=2.03 $X2=3.45 $Y2=2.53
r74 2 21 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=3.31
+ $Y=2.03 $X2=3.45 $Y2=2.175
r75 1 12 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=1.225
+ $Y=2.03 $X2=1.37 $Y2=2.885
r76 1 9 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=1.225
+ $Y=2.03 $X2=1.37 $Y2=2.175
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSTP_LP%A_352_406# 1 2 3 4 15 17 18 19 22 23 26 27
+ 28 30 31 32 34 35 36 41 45 48 50 52 54 55
c171 52 0 1.98095e-19 $X=5.365 $Y=1.245
c172 50 0 1.29843e-19 $X=3.1 $Y=0.845
c173 32 0 6.89731e-20 $X=4.41 $Y=1.245
r174 54 55 8.63679 $w=3.28e-07 $l=1.7e-07 $layer=LI1_cond $X=5.525 $Y=2.02
+ $X2=5.525 $Y2=2.19
r175 51 52 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=5.075 $Y=1.245
+ $X2=5.365 $Y2=1.245
r176 43 45 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=6.065 $Y=0.435
+ $X2=6.065 $Y2=0.835
r177 41 55 7.15912 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=5.605 $Y=2.395
+ $X2=5.605 $Y2=2.19
r178 37 52 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.365 $Y=1.33
+ $X2=5.365 $Y2=1.245
r179 37 54 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=5.365 $Y=1.33
+ $X2=5.365 $Y2=2.02
r180 35 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.98 $Y=0.35
+ $X2=6.065 $Y2=0.435
r181 35 36 53.4973 $w=1.68e-07 $l=8.2e-07 $layer=LI1_cond $X=5.98 $Y=0.35
+ $X2=5.16 $Y2=0.35
r182 34 51 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.075 $Y=1.16
+ $X2=5.075 $Y2=1.245
r183 33 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.075 $Y=0.435
+ $X2=5.16 $Y2=0.35
r184 33 34 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=5.075 $Y=0.435
+ $X2=5.075 $Y2=1.16
r185 31 51 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=4.99 $Y=1.245
+ $X2=5.075 $Y2=1.245
r186 31 32 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=4.99 $Y=1.245
+ $X2=4.41 $Y2=1.245
r187 30 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.325 $Y=1.16
+ $X2=4.41 $Y2=1.245
r188 29 30 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=4.325 $Y=0.435
+ $X2=4.325 $Y2=1.16
r189 27 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.24 $Y=0.35
+ $X2=4.325 $Y2=0.435
r190 27 28 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=4.24 $Y=0.35
+ $X2=3.625 $Y2=0.35
r191 25 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.54 $Y=0.435
+ $X2=3.625 $Y2=0.35
r192 25 26 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=3.54 $Y=0.435
+ $X2=3.54 $Y2=0.76
r193 24 50 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.185 $Y=0.845
+ $X2=3.1 $Y2=0.845
r194 23 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.455 $Y=0.845
+ $X2=3.54 $Y2=0.76
r195 23 24 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=3.455 $Y=0.845
+ $X2=3.185 $Y2=0.845
r196 21 50 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.1 $Y=0.93 $X2=3.1
+ $Y2=0.845
r197 21 22 67.8503 $w=1.68e-07 $l=1.04e-06 $layer=LI1_cond $X=3.1 $Y=0.93
+ $X2=3.1 $Y2=1.97
r198 20 48 15.8958 $w=3.07e-07 $l=4.93964e-07 $layer=LI1_cond $X=2.625 $Y=0.845
+ $X2=2.415 $Y2=0.445
r199 19 50 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.015 $Y=0.845
+ $X2=3.1 $Y2=0.845
r200 19 20 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=3.015 $Y=0.845
+ $X2=2.625 $Y2=0.845
r201 17 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.015 $Y=2.055
+ $X2=3.1 $Y2=1.97
r202 17 18 61.9786 $w=1.68e-07 $l=9.5e-07 $layer=LI1_cond $X=3.015 $Y=2.055
+ $X2=2.065 $Y2=2.055
r203 13 18 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.9 $Y=2.14
+ $X2=2.065 $Y2=2.055
r204 13 15 1.22229 $w=3.28e-07 $l=3.5e-08 $layer=LI1_cond $X=1.9 $Y=2.14 $X2=1.9
+ $Y2=2.175
r205 4 41 600 $w=1.7e-07 $l=3.61248e-07 $layer=licon1_PDIFF $count=1 $X=5.47
+ $Y=2.095 $X2=5.605 $Y2=2.395
r206 3 15 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=1.76
+ $Y=2.03 $X2=1.9 $Y2=2.175
r207 2 45 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=5.92
+ $Y=0.625 $X2=6.065 $Y2=0.835
r208 1 48 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.23
+ $Y=0.235 $X2=2.37 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSTP_LP%Q 1 2 9 12 13 14 15 16 38 42
c21 38 0 6.94276e-20 $X=15.37 $Y=2.015
r22 38 39 7.29421 $w=5.18e-07 $l=1.65e-07 $layer=LI1_cond $X=15.465 $Y=2.015
+ $X2=15.465 $Y2=1.85
r23 28 42 1.72511 $w=5.18e-07 $l=7.5e-08 $layer=LI1_cond $X=15.465 $Y=2.11
+ $X2=15.465 $Y2=2.035
r24 16 33 1.15008 $w=5.18e-07 $l=5e-08 $layer=LI1_cond $X=15.465 $Y=2.775
+ $X2=15.465 $Y2=2.725
r25 15 33 7.36048 $w=5.18e-07 $l=3.2e-07 $layer=LI1_cond $X=15.465 $Y=2.405
+ $X2=15.465 $Y2=2.725
r26 14 42 0.115008 $w=5.18e-07 $l=5e-09 $layer=LI1_cond $X=15.465 $Y=2.03
+ $X2=15.465 $Y2=2.035
r27 14 38 0.345023 $w=5.18e-07 $l=1.5e-08 $layer=LI1_cond $X=15.465 $Y=2.03
+ $X2=15.465 $Y2=2.015
r28 14 15 6.67044 $w=5.18e-07 $l=2.9e-07 $layer=LI1_cond $X=15.465 $Y=2.115
+ $X2=15.465 $Y2=2.405
r29 14 28 0.115008 $w=5.18e-07 $l=5e-09 $layer=LI1_cond $X=15.465 $Y=2.115
+ $X2=15.465 $Y2=2.11
r30 13 39 8.88342 $w=2.38e-07 $l=1.85e-07 $layer=LI1_cond $X=15.605 $Y=1.665
+ $X2=15.605 $Y2=1.85
r31 12 13 17.7668 $w=2.38e-07 $l=3.7e-07 $layer=LI1_cond $X=15.605 $Y=1.295
+ $X2=15.605 $Y2=1.665
r32 11 12 27.3705 $w=2.38e-07 $l=5.7e-07 $layer=LI1_cond $X=15.605 $Y=0.725
+ $X2=15.605 $Y2=1.295
r33 9 11 8.90991 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=15.56 $Y=0.495
+ $X2=15.56 $Y2=0.725
r34 2 38 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=15.23
+ $Y=1.87 $X2=15.37 $Y2=2.015
r35 2 33 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=15.23
+ $Y=1.87 $X2=15.37 $Y2=2.725
r36 1 9 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=15.42
+ $Y=0.285 $X2=15.56 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__SDFSTP_LP%VGND 1 2 3 4 5 6 7 8 27 31 35 39 43 47 51
+ 55 58 59 61 62 64 65 66 68 73 88 95 113 119 120 123 126 129 132 135
c172 73 0 1.29843e-19 $X=3.025 $Y=0
c173 47 0 1.32475e-20 $X=11.54 $Y=0.52
r174 135 136 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=14.64 $Y=0
+ $X2=14.64 $Y2=0
r175 132 133 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=9.36 $Y=0
+ $X2=9.36 $Y2=0
r176 129 130 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.44 $Y=0
+ $X2=7.44 $Y2=0
r177 126 127 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0
+ $X2=3.12 $Y2=0
r178 123 124 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r179 120 136 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=15.6 $Y=0
+ $X2=14.64 $Y2=0
r180 119 120 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=15.6 $Y=0
+ $X2=15.6 $Y2=0
r181 117 135 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=14.935 $Y=0
+ $X2=14.77 $Y2=0
r182 117 119 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=14.935 $Y=0
+ $X2=15.6 $Y2=0
r183 116 136 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=13.68 $Y=0
+ $X2=14.64 $Y2=0
r184 115 116 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=13.68 $Y=0
+ $X2=13.68 $Y2=0
r185 113 135 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=14.605 $Y=0
+ $X2=14.77 $Y2=0
r186 113 115 60.3476 $w=1.68e-07 $l=9.25e-07 $layer=LI1_cond $X=14.605 $Y=0
+ $X2=13.68 $Y2=0
r187 112 116 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=13.2 $Y=0
+ $X2=13.68 $Y2=0
r188 111 112 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=13.2 $Y=0
+ $X2=13.2 $Y2=0
r189 109 112 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=11.76 $Y=0
+ $X2=13.2 $Y2=0
r190 108 111 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=11.76 $Y=0
+ $X2=13.2 $Y2=0
r191 108 109 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.76 $Y=0
+ $X2=11.76 $Y2=0
r192 106 109 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=11.28 $Y=0
+ $X2=11.76 $Y2=0
r193 106 133 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=11.28 $Y=0
+ $X2=9.36 $Y2=0
r194 105 106 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=11.28 $Y=0
+ $X2=11.28 $Y2=0
r195 103 132 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.415 $Y=0
+ $X2=9.25 $Y2=0
r196 103 105 121.674 $w=1.68e-07 $l=1.865e-06 $layer=LI1_cond $X=9.415 $Y=0
+ $X2=11.28 $Y2=0
r197 102 133 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=0
+ $X2=9.36 $Y2=0
r198 101 102 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.88 $Y=0
+ $X2=8.88 $Y2=0
r199 98 101 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=7.92 $Y=0 $X2=8.88
+ $Y2=0
r200 96 129 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.565 $Y=0
+ $X2=7.44 $Y2=0
r201 96 98 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=7.565 $Y=0
+ $X2=7.92 $Y2=0
r202 95 132 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.085 $Y=0
+ $X2=9.25 $Y2=0
r203 95 101 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=9.085 $Y=0
+ $X2=8.88 $Y2=0
r204 94 130 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.96 $Y=0
+ $X2=7.44 $Y2=0
r205 93 94 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.96 $Y=0
+ $X2=6.96 $Y2=0
r206 91 94 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=5.04 $Y=0
+ $X2=6.96 $Y2=0
r207 90 93 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=5.04 $Y=0 $X2=6.96
+ $Y2=0
r208 90 91 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.04 $Y=0
+ $X2=5.04 $Y2=0
r209 88 129 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.315 $Y=0
+ $X2=7.44 $Y2=0
r210 88 93 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=7.315 $Y=0
+ $X2=6.96 $Y2=0
r211 87 91 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.04
+ $Y2=0
r212 86 87 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r213 84 87 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.56
+ $Y2=0
r214 84 127 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=3.12
+ $Y2=0
r215 83 86 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=3.6 $Y=0 $X2=4.56
+ $Y2=0
r216 83 84 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r217 81 126 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.275 $Y=0
+ $X2=3.15 $Y2=0
r218 81 83 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=3.275 $Y=0 $X2=3.6
+ $Y2=0
r219 80 127 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0
+ $X2=3.12 $Y2=0
r220 79 80 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r221 77 80 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r222 77 124 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r223 76 79 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r224 76 77 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r225 74 123 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.385 $Y=0
+ $X2=1.22 $Y2=0
r226 74 76 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.385 $Y=0 $X2=1.68
+ $Y2=0
r227 73 126 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.025 $Y=0
+ $X2=3.15 $Y2=0
r228 73 79 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=3.025 $Y=0
+ $X2=2.64 $Y2=0
r229 71 124 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r230 70 71 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r231 68 123 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.055 $Y=0
+ $X2=1.22 $Y2=0
r232 68 70 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.055 $Y=0
+ $X2=0.72 $Y2=0
r233 66 102 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.92 $Y=0
+ $X2=8.88 $Y2=0
r234 66 130 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.92 $Y=0
+ $X2=7.44 $Y2=0
r235 66 98 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r236 64 111 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=13.255 $Y=0
+ $X2=13.2 $Y2=0
r237 64 65 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.255 $Y=0
+ $X2=13.42 $Y2=0
r238 63 115 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=13.585 $Y=0
+ $X2=13.68 $Y2=0
r239 63 65 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.585 $Y=0
+ $X2=13.42 $Y2=0
r240 61 105 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=11.375 $Y=0
+ $X2=11.28 $Y2=0
r241 61 62 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.375 $Y=0
+ $X2=11.54 $Y2=0
r242 60 108 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=11.705 $Y=0
+ $X2=11.76 $Y2=0
r243 60 62 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.705 $Y=0
+ $X2=11.54 $Y2=0
r244 58 86 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=4.63 $Y=0 $X2=4.56
+ $Y2=0
r245 58 59 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.63 $Y=0 $X2=4.715
+ $Y2=0
r246 57 90 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=4.8 $Y=0 $X2=5.04
+ $Y2=0
r247 57 59 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.8 $Y=0 $X2=4.715
+ $Y2=0
r248 53 135 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=14.77 $Y=0.085
+ $X2=14.77 $Y2=0
r249 53 55 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=14.77 $Y=0.085
+ $X2=14.77 $Y2=0.495
r250 49 65 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=13.42 $Y=0.085
+ $X2=13.42 $Y2=0
r251 49 51 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=13.42 $Y=0.085
+ $X2=13.42 $Y2=0.495
r252 45 62 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=11.54 $Y=0.085
+ $X2=11.54 $Y2=0
r253 45 47 15.1913 $w=3.28e-07 $l=4.35e-07 $layer=LI1_cond $X=11.54 $Y=0.085
+ $X2=11.54 $Y2=0.52
r254 41 132 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.25 $Y=0.085
+ $X2=9.25 $Y2=0
r255 41 43 26.1919 $w=3.28e-07 $l=7.5e-07 $layer=LI1_cond $X=9.25 $Y=0.085
+ $X2=9.25 $Y2=0.835
r256 37 129 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.44 $Y=0.085
+ $X2=7.44 $Y2=0
r257 37 39 20.0525 $w=2.48e-07 $l=4.35e-07 $layer=LI1_cond $X=7.44 $Y=0.085
+ $X2=7.44 $Y2=0.52
r258 33 59 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.715 $Y=0.085
+ $X2=4.715 $Y2=0
r259 33 35 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=4.715 $Y=0.085
+ $X2=4.715 $Y2=0.75
r260 29 126 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.15 $Y=0.085
+ $X2=3.15 $Y2=0
r261 29 31 14.2903 $w=2.48e-07 $l=3.1e-07 $layer=LI1_cond $X=3.15 $Y=0.085
+ $X2=3.15 $Y2=0.395
r262 25 123 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.22 $Y=0.085
+ $X2=1.22 $Y2=0
r263 25 27 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=1.22 $Y=0.085
+ $X2=1.22 $Y2=0.445
r264 8 55 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=14.63
+ $Y=0.285 $X2=14.77 $Y2=0.495
r265 7 51 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=13.28
+ $Y=0.285 $X2=13.42 $Y2=0.495
r266 6 47 182 $w=1.7e-07 $l=2.504e-07 $layer=licon1_NDIFF $count=1 $X=11.4
+ $Y=0.33 $X2=11.54 $Y2=0.52
r267 5 43 182 $w=1.7e-07 $l=2.86182e-07 $layer=licon1_NDIFF $count=1 $X=9.07
+ $Y=0.625 $X2=9.25 $Y2=0.835
r268 4 39 182 $w=1.7e-07 $l=2.52091e-07 $layer=licon1_NDIFF $count=1 $X=7.275
+ $Y=0.625 $X2=7.48 $Y2=0.52
r269 3 35 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=4.575
+ $Y=0.54 $X2=4.715 $Y2=0.75
r270 2 31 182 $w=1.7e-07 $l=2.19089e-07 $layer=licon1_NDIFF $count=1 $X=3.05
+ $Y=0.235 $X2=3.19 $Y2=0.395
r271 1 27 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.08
+ $Y=0.235 $X2=1.22 $Y2=0.445
.ends

