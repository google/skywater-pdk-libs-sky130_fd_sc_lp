# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_sc_lp__sdfsbp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_lp__sdfsbp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  15.36000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.105000 0.765000 1.915000 1.775000 ;
        RECT 1.105000 1.775000 1.555000 1.945000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.573300 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 13.915000 1.020000 14.250000 3.075000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.556500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 14.835000 1.840000 15.275000 3.075000 ;
        RECT 15.005000 0.380000 15.275000 1.840000 ;
    END
  END Q_N
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.545000 1.080000 2.735000 2.205000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.560000 1.915000 0.935000 2.125000 ;
        RECT 0.560000 2.125000 2.375000 2.295000 ;
        RECT 2.125000 0.995000 2.375000 2.125000 ;
    END
  END SCE
  PIN SET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT  7.295000 1.920000  7.585000 1.965000 ;
        RECT  7.295000 1.965000 10.945000 2.105000 ;
        RECT  7.295000 2.105000  7.585000 2.150000 ;
        RECT 10.655000 1.920000 10.945000 1.965000 ;
        RECT 10.655000 2.105000 10.945000 2.150000 ;
    END
  END SET_B
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 3.275000 0.830000 3.755000 1.885000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 15.360000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.000000 0.000000 15.360000 0.245000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.655000 15.550000 3.520000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 15.360000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 15.360000 0.085000 ;
      RECT  0.000000  3.245000 15.360000 3.415000 ;
      RECT  0.130000  0.280000  0.635000 0.610000 ;
      RECT  0.130000  0.610000  0.380000 1.125000 ;
      RECT  0.130000  1.125000  0.935000 1.455000 ;
      RECT  0.130000  1.455000  0.390000 3.065000 ;
      RECT  0.560000  2.465000  0.890000 3.245000 ;
      RECT  0.805000  0.085000  1.135000 0.595000 ;
      RECT  1.460000  2.475000  3.075000 2.645000 ;
      RECT  1.460000  2.645000  1.790000 3.025000 ;
      RECT  1.595000  0.280000  2.540000 0.595000 ;
      RECT  2.370000  0.595000  2.540000 0.655000 ;
      RECT  2.370000  0.655000  3.075000 0.825000 ;
      RECT  2.405000  2.815000  2.735000 3.245000 ;
      RECT  2.790000  0.085000  3.120000 0.485000 ;
      RECT  2.905000  0.825000  3.075000 2.475000 ;
      RECT  2.905000  2.645000  3.075000 2.895000 ;
      RECT  2.905000  2.895000  3.775000 3.065000 ;
      RECT  3.245000  2.230000  4.125000 2.435000 ;
      RECT  3.245000  2.435000  3.435000 2.725000 ;
      RECT  3.290000  0.330000  4.125000 0.660000 ;
      RECT  3.605000  2.615000  5.575000 2.785000 ;
      RECT  3.605000  2.785000  3.775000 2.895000 ;
      RECT  3.925000  0.660000  4.125000 2.230000 ;
      RECT  3.955000  2.955000  4.285000 3.245000 ;
      RECT  4.295000  0.085000  4.535000 0.730000 ;
      RECT  4.480000  1.375000  5.105000 2.435000 ;
      RECT  4.705000  0.400000  5.005000 1.375000 ;
      RECT  5.255000  0.585000  5.670000 0.865000 ;
      RECT  5.255000  0.865000  5.455000 1.035000 ;
      RECT  5.275000  1.035000  5.455000 2.360000 ;
      RECT  5.275000  2.360000  5.575000 2.615000 ;
      RECT  5.625000  1.035000  8.335000 1.205000 ;
      RECT  5.625000  1.205000  5.795000 1.885000 ;
      RECT  5.625000  1.885000  6.035000 2.055000 ;
      RECT  5.745000  2.055000  6.035000 2.690000 ;
      RECT  5.840000  0.640000  6.100000 1.025000 ;
      RECT  5.840000  1.025000  8.335000 1.035000 ;
      RECT  5.965000  1.375000  7.985000 1.545000 ;
      RECT  5.965000  1.545000  6.225000 1.705000 ;
      RECT  6.455000  1.905000  7.175000 2.190000 ;
      RECT  6.505000  2.360000  6.835000 3.245000 ;
      RECT  6.560000  0.085000  6.890000 0.855000 ;
      RECT  7.005000  2.190000  7.175000 2.300000 ;
      RECT  7.005000  2.300000  9.475000 2.470000 ;
      RECT  7.005000  2.470000  7.480000 2.690000 ;
      RECT  7.060000  0.525000  7.250000 1.025000 ;
      RECT  7.345000  1.790000  7.645000 2.130000 ;
      RECT  7.420000  0.635000  8.685000 0.855000 ;
      RECT  7.650000  2.640000  8.885000 3.245000 ;
      RECT  7.815000  1.545000  7.985000 1.780000 ;
      RECT  7.815000  1.780000  9.125000 1.950000 ;
      RECT  8.165000  1.205000  8.335000 1.420000 ;
      RECT  8.165000  1.420000  8.775000 1.610000 ;
      RECT  8.515000  0.855000  8.685000 1.080000 ;
      RECT  8.515000  1.080000 10.130000 1.250000 ;
      RECT  8.855000  0.085000  9.055000 0.910000 ;
      RECT  8.955000  1.420000  9.790000 1.610000 ;
      RECT  8.955000  1.610000  9.125000 1.780000 ;
      RECT  9.305000  1.780000 10.130000 1.950000 ;
      RECT  9.305000  1.950000  9.475000 2.300000 ;
      RECT  9.575000  0.640000 10.480000 0.910000 ;
      RECT  9.645000  2.120000 10.480000 2.300000 ;
      RECT  9.645000  2.300000 11.655000 2.470000 ;
      RECT  9.645000  2.470000 10.150000 2.880000 ;
      RECT  9.960000  1.250000 10.130000 1.780000 ;
      RECT 10.310000  0.910000 10.480000 2.120000 ;
      RECT 10.460000  2.640000 11.225000 3.245000 ;
      RECT 10.650000  1.920000 11.530000 2.130000 ;
      RECT 10.660000  1.495000 12.150000 1.750000 ;
      RECT 10.820000  0.085000 11.150000 0.960000 ;
      RECT 11.375000  0.795000 11.730000 1.495000 ;
      RECT 11.395000  2.470000 11.655000 2.905000 ;
      RECT 11.395000  2.905000 12.685000 3.075000 ;
      RECT 11.900000  0.085000 12.455000 1.080000 ;
      RECT 11.975000  1.750000 12.150000 2.465000 ;
      RECT 11.975000  2.465000 12.345000 2.735000 ;
      RECT 12.320000  1.590000 12.795000 2.010000 ;
      RECT 12.320000  2.010000 12.685000 2.260000 ;
      RECT 12.515000  2.260000 12.685000 2.905000 ;
      RECT 12.625000  0.450000 13.735000 0.620000 ;
      RECT 12.625000  0.620000 12.795000 1.590000 ;
      RECT 12.855000  2.180000 13.115000 3.245000 ;
      RECT 12.965000  0.790000 13.235000 1.160000 ;
      RECT 12.965000  1.160000 13.665000 1.330000 ;
      RECT 13.285000  1.330000 13.665000 1.830000 ;
      RECT 13.285000  1.830000 13.545000 2.860000 ;
      RECT 13.405000  0.330000 13.735000 0.450000 ;
      RECT 13.405000  0.620000 13.735000 0.680000 ;
      RECT 13.405000  0.680000 14.835000 0.850000 ;
      RECT 14.425000  0.085000 14.755000 0.510000 ;
      RECT 14.425000  1.840000 14.615000 3.245000 ;
      RECT 14.665000  0.850000 14.835000 1.670000 ;
    LAYER mcon ;
      RECT  0.155000 -0.085000  0.325000 0.085000 ;
      RECT  0.155000  3.245000  0.325000 3.415000 ;
      RECT  0.635000 -0.085000  0.805000 0.085000 ;
      RECT  0.635000  3.245000  0.805000 3.415000 ;
      RECT  1.115000 -0.085000  1.285000 0.085000 ;
      RECT  1.115000  3.245000  1.285000 3.415000 ;
      RECT  1.595000 -0.085000  1.765000 0.085000 ;
      RECT  1.595000  3.245000  1.765000 3.415000 ;
      RECT  2.075000 -0.085000  2.245000 0.085000 ;
      RECT  2.075000  3.245000  2.245000 3.415000 ;
      RECT  2.555000 -0.085000  2.725000 0.085000 ;
      RECT  2.555000  3.245000  2.725000 3.415000 ;
      RECT  3.035000 -0.085000  3.205000 0.085000 ;
      RECT  3.035000  3.245000  3.205000 3.415000 ;
      RECT  3.515000 -0.085000  3.685000 0.085000 ;
      RECT  3.515000  3.245000  3.685000 3.415000 ;
      RECT  3.995000 -0.085000  4.165000 0.085000 ;
      RECT  3.995000  3.245000  4.165000 3.415000 ;
      RECT  4.475000 -0.085000  4.645000 0.085000 ;
      RECT  4.475000  3.245000  4.645000 3.415000 ;
      RECT  4.955000 -0.085000  5.125000 0.085000 ;
      RECT  4.955000  3.245000  5.125000 3.415000 ;
      RECT  5.435000 -0.085000  5.605000 0.085000 ;
      RECT  5.435000  3.245000  5.605000 3.415000 ;
      RECT  5.915000 -0.085000  6.085000 0.085000 ;
      RECT  5.915000  3.245000  6.085000 3.415000 ;
      RECT  6.395000 -0.085000  6.565000 0.085000 ;
      RECT  6.395000  3.245000  6.565000 3.415000 ;
      RECT  6.875000 -0.085000  7.045000 0.085000 ;
      RECT  6.875000  3.245000  7.045000 3.415000 ;
      RECT  7.355000 -0.085000  7.525000 0.085000 ;
      RECT  7.355000  1.950000  7.525000 2.120000 ;
      RECT  7.355000  3.245000  7.525000 3.415000 ;
      RECT  7.835000 -0.085000  8.005000 0.085000 ;
      RECT  7.835000  3.245000  8.005000 3.415000 ;
      RECT  8.315000 -0.085000  8.485000 0.085000 ;
      RECT  8.315000  3.245000  8.485000 3.415000 ;
      RECT  8.795000 -0.085000  8.965000 0.085000 ;
      RECT  8.795000  3.245000  8.965000 3.415000 ;
      RECT  9.275000 -0.085000  9.445000 0.085000 ;
      RECT  9.275000  3.245000  9.445000 3.415000 ;
      RECT  9.755000 -0.085000  9.925000 0.085000 ;
      RECT  9.755000  3.245000  9.925000 3.415000 ;
      RECT 10.235000 -0.085000 10.405000 0.085000 ;
      RECT 10.235000  3.245000 10.405000 3.415000 ;
      RECT 10.715000 -0.085000 10.885000 0.085000 ;
      RECT 10.715000  1.950000 10.885000 2.120000 ;
      RECT 10.715000  3.245000 10.885000 3.415000 ;
      RECT 11.195000 -0.085000 11.365000 0.085000 ;
      RECT 11.195000  3.245000 11.365000 3.415000 ;
      RECT 11.675000 -0.085000 11.845000 0.085000 ;
      RECT 11.675000  3.245000 11.845000 3.415000 ;
      RECT 12.155000 -0.085000 12.325000 0.085000 ;
      RECT 12.155000  3.245000 12.325000 3.415000 ;
      RECT 12.635000 -0.085000 12.805000 0.085000 ;
      RECT 12.635000  3.245000 12.805000 3.415000 ;
      RECT 13.115000 -0.085000 13.285000 0.085000 ;
      RECT 13.115000  3.245000 13.285000 3.415000 ;
      RECT 13.595000 -0.085000 13.765000 0.085000 ;
      RECT 13.595000  3.245000 13.765000 3.415000 ;
      RECT 14.075000 -0.085000 14.245000 0.085000 ;
      RECT 14.075000  3.245000 14.245000 3.415000 ;
      RECT 14.555000 -0.085000 14.725000 0.085000 ;
      RECT 14.555000  3.245000 14.725000 3.415000 ;
      RECT 15.035000 -0.085000 15.205000 0.085000 ;
      RECT 15.035000  3.245000 15.205000 3.415000 ;
  END
END sky130_fd_sc_lp__sdfsbp_1
END LIBRARY
