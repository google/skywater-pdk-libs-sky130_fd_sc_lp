* File: sky130_fd_sc_lp__o2bb2a_m.spice
* Created: Fri Aug 28 11:12:17 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__o2bb2a_m.pex.spice"
.subckt sky130_fd_sc_lp__o2bb2a_m  VNB VPB A1_N A2_N B2 B1 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* B1	B1
* B2	B2
* A2_N	A2_N
* A1_N	A1_N
* VPB	VPB
* VNB	VNB
MM1006 N_VGND_M1006_d N_A_85_187#_M1006_g N_X_M1006_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75001.2
+ A=0.063 P=1.14 MULT=1
MM1007 A_223_47# N_A1_N_M1007_g N_VGND_M1006_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.8 A=0.063 P=1.14 MULT=1
MM1008 N_A_209_535#_M1008_d N_A2_N_M1008_g A_223_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.2172 AS=0.0441 PD=2.02 PS=0.63 NRD=87.132 NRS=14.28 M=1 R=2.8 SA=75001
+ SB=75000.4 A=0.063 P=1.14 MULT=1
MM1003 N_A_487_167#_M1003_d N_A_209_535#_M1003_g N_A_85_187#_M1003_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1004 N_VGND_M1004_d N_B2_M1004_g N_A_487_167#_M1003_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0672 AS=0.0588 PD=0.74 PS=0.7 NRD=5.712 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1005 N_A_487_167#_M1005_d N_B1_M1005_g N_VGND_M1004_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.0672 PD=1.37 PS=0.74 NRD=0 NRS=5.712 M=1 R=2.8 SA=75001.1
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1001 N_VPWR_M1001_d N_A_85_187#_M1001_g N_X_M1001_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0672 AS=0.1113 PD=0.74 PS=1.37 NRD=9.3772 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.8 A=0.063 P=1.14 MULT=1
MM1011 N_A_209_535#_M1011_d N_A1_N_M1011_g N_VPWR_M1001_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0588 AS=0.0672 PD=0.7 PS=0.74 NRD=0 NRS=9.3772 M=1 R=2.8
+ SA=75000.7 SB=75002.3 A=0.063 P=1.14 MULT=1
MM1002 N_VPWR_M1002_d N_A2_N_M1002_g N_A_209_535#_M1011_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1554 AS=0.0588 PD=1.16 PS=0.7 NRD=114.91 NRS=0 M=1 R=2.8
+ SA=75001.1 SB=75001.9 A=0.063 P=1.14 MULT=1
MM1000 N_A_85_187#_M1000_d N_A_209_535#_M1000_g N_VPWR_M1002_d VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.0588 AS=0.1554 PD=0.7 PS=1.16 NRD=0 NRS=100.844 M=1 R=2.8
+ SA=75002 SB=75001 A=0.063 P=1.14 MULT=1
MM1009 A_559_535# N_B2_M1009_g N_A_85_187#_M1000_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=23.443 NRS=0 M=1 R=2.8 SA=75002.4
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1010 N_VPWR_M1010_d N_B1_M1010_g A_559_535# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.1113 AS=0.0441 PD=1.37 PS=0.63 NRD=0 NRS=23.443 M=1 R=2.8 SA=75002.8
+ SB=75000.2 A=0.063 P=1.14 MULT=1
DX12_noxref VNB VPB NWDIODE A=7.8703 P=12.17
*
.include "sky130_fd_sc_lp__o2bb2a_m.pxi.spice"
*
.ends
*
*
