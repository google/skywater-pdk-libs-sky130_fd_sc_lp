* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__a31o_lp A1 A2 A3 B1 VGND VNB VPB VPWR X
X0 a_352_56# A3 VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 a_155_409# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X2 a_48_409# B1 a_155_409# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X3 a_274_56# A2 a_352_56# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 a_516_56# a_48_409# X VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 a_155_409# A3 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X6 VPWR A2 a_155_409# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
X7 a_116_56# B1 a_48_409# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 VGND B1 a_116_56# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 a_48_409# A1 a_274_56# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 VGND a_48_409# a_516_56# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X11 VPWR a_48_409# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=250000u
.ends
