# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__sdfxtp_2
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__sdfxtp_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  11.04000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.115000 0.385000 1.765000 1.455000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.588000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.225000 0.375000 10.465000 3.075000 ;
    END
  END Q
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.035000 1.455000 2.725000 1.775000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.450000 1.140000 0.830000 2.130000 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 3.255000 1.200000 3.735000 2.120000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT  0.000000 -0.085000 11.040000 0.085000 ;
        RECT  0.725000  0.085000  0.945000 0.970000 ;
        RECT  2.695000  0.085000  3.025000 0.945000 ;
        RECT  3.695000  0.085000  4.025000 0.530000 ;
        RECT  6.205000  0.085000  6.545000 0.555000 ;
        RECT  8.830000  0.085000  9.040000 0.885000 ;
        RECT  9.745000  0.085000 10.055000 1.175000 ;
        RECT 10.635000  0.085000 10.935000 1.255000 ;
      LAYER mcon ;
        RECT  0.155000 -0.085000  0.325000 0.085000 ;
        RECT  0.635000 -0.085000  0.805000 0.085000 ;
        RECT  1.115000 -0.085000  1.285000 0.085000 ;
        RECT  1.595000 -0.085000  1.765000 0.085000 ;
        RECT  2.075000 -0.085000  2.245000 0.085000 ;
        RECT  2.555000 -0.085000  2.725000 0.085000 ;
        RECT  3.035000 -0.085000  3.205000 0.085000 ;
        RECT  3.515000 -0.085000  3.685000 0.085000 ;
        RECT  3.995000 -0.085000  4.165000 0.085000 ;
        RECT  4.475000 -0.085000  4.645000 0.085000 ;
        RECT  4.955000 -0.085000  5.125000 0.085000 ;
        RECT  5.435000 -0.085000  5.605000 0.085000 ;
        RECT  5.915000 -0.085000  6.085000 0.085000 ;
        RECT  6.395000 -0.085000  6.565000 0.085000 ;
        RECT  6.875000 -0.085000  7.045000 0.085000 ;
        RECT  7.355000 -0.085000  7.525000 0.085000 ;
        RECT  7.835000 -0.085000  8.005000 0.085000 ;
        RECT  8.315000 -0.085000  8.485000 0.085000 ;
        RECT  8.795000 -0.085000  8.965000 0.085000 ;
        RECT  9.275000 -0.085000  9.445000 0.085000 ;
        RECT  9.755000 -0.085000  9.925000 0.085000 ;
        RECT 10.235000 -0.085000 10.405000 0.085000 ;
        RECT 10.715000 -0.085000 10.885000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.245000 11.040000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT  0.000000 3.245000 11.040000 3.415000 ;
        RECT  0.780000 2.640000  1.110000 3.245000 ;
        RECT  2.625000 2.690000  2.845000 3.245000 ;
        RECT  3.555000 2.640000  3.805000 3.245000 ;
        RECT  6.095000 2.455000  6.375000 3.245000 ;
        RECT  8.450000 2.325000  9.125000 3.245000 ;
        RECT  9.745000 1.845000 10.055000 3.245000 ;
        RECT 10.635000 1.815000 10.935000 3.245000 ;
      LAYER mcon ;
        RECT  0.155000 3.245000  0.325000 3.415000 ;
        RECT  0.635000 3.245000  0.805000 3.415000 ;
        RECT  1.115000 3.245000  1.285000 3.415000 ;
        RECT  1.595000 3.245000  1.765000 3.415000 ;
        RECT  2.075000 3.245000  2.245000 3.415000 ;
        RECT  2.555000 3.245000  2.725000 3.415000 ;
        RECT  3.035000 3.245000  3.205000 3.415000 ;
        RECT  3.515000 3.245000  3.685000 3.415000 ;
        RECT  3.995000 3.245000  4.165000 3.415000 ;
        RECT  4.475000 3.245000  4.645000 3.415000 ;
        RECT  4.955000 3.245000  5.125000 3.415000 ;
        RECT  5.435000 3.245000  5.605000 3.415000 ;
        RECT  5.915000 3.245000  6.085000 3.415000 ;
        RECT  6.395000 3.245000  6.565000 3.415000 ;
        RECT  6.875000 3.245000  7.045000 3.415000 ;
        RECT  7.355000 3.245000  7.525000 3.415000 ;
        RECT  7.835000 3.245000  8.005000 3.415000 ;
        RECT  8.315000 3.245000  8.485000 3.415000 ;
        RECT  8.795000 3.245000  8.965000 3.415000 ;
        RECT  9.275000 3.245000  9.445000 3.415000 ;
        RECT  9.755000 3.245000  9.925000 3.415000 ;
        RECT 10.235000 3.245000 10.405000 3.415000 ;
        RECT 10.715000 3.245000 10.885000 3.415000 ;
      LAYER met1 ;
        RECT 0.000000 3.085000 11.040000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.110000 0.640000  0.555000 0.970000 ;
      RECT 0.110000 0.970000  0.280000 2.300000 ;
      RECT 0.110000 2.300000  1.170000 2.470000 ;
      RECT 0.315000 2.470000  0.610000 3.075000 ;
      RECT 1.000000 1.635000  1.250000 1.945000 ;
      RECT 1.000000 1.945000  2.115000 2.275000 ;
      RECT 1.000000 2.275000  1.170000 2.300000 ;
      RECT 1.615000 2.445000  2.725000 2.520000 ;
      RECT 1.615000 2.520000  2.455000 2.645000 ;
      RECT 1.615000 2.645000  1.945000 3.075000 ;
      RECT 1.935000 0.635000  2.135000 1.115000 ;
      RECT 1.935000 1.115000  3.075000 1.285000 ;
      RECT 2.285000 1.950000  3.075000 2.120000 ;
      RECT 2.285000 2.120000  2.725000 2.445000 ;
      RECT 2.905000 1.285000  3.075000 1.950000 ;
      RECT 3.025000 2.300000  4.145000 2.470000 ;
      RECT 3.025000 2.470000  3.355000 3.025000 ;
      RECT 3.225000 0.700000  3.905000 0.860000 ;
      RECT 3.225000 0.860000  4.145000 1.030000 ;
      RECT 3.905000 1.030000  4.145000 2.300000 ;
      RECT 3.975000 2.470000  4.145000 2.835000 ;
      RECT 3.975000 2.835000  5.845000 3.005000 ;
      RECT 4.195000 0.265000  5.965000 0.485000 ;
      RECT 4.195000 0.485000  4.535000 0.610000 ;
      RECT 4.315000 0.610000  4.535000 1.175000 ;
      RECT 4.315000 1.175000  4.625000 2.665000 ;
      RECT 4.760000 0.655000  5.090000 0.905000 ;
      RECT 4.760000 0.905000  4.965000 0.955000 ;
      RECT 4.795000 0.955000  4.965000 2.275000 ;
      RECT 4.795000 2.275000  5.135000 2.590000 ;
      RECT 5.145000 1.075000  6.935000 1.245000 ;
      RECT 5.145000 1.245000  5.315000 1.935000 ;
      RECT 5.145000 1.935000  5.495000 2.105000 ;
      RECT 5.270000 0.670000  5.490000 1.075000 ;
      RECT 5.305000 2.105000  5.495000 2.630000 ;
      RECT 5.485000 1.425000  5.845000 1.755000 ;
      RECT 5.660000 0.485000  5.965000 0.725000 ;
      RECT 5.660000 0.725000  6.935000 0.895000 ;
      RECT 5.675000 1.755000  5.845000 2.115000 ;
      RECT 5.675000 2.115000  6.715000 2.285000 ;
      RECT 5.675000 2.285000  5.845000 2.835000 ;
      RECT 6.025000 1.425000  6.355000 1.495000 ;
      RECT 6.025000 1.495000  7.295000 1.665000 ;
      RECT 6.025000 1.665000  7.125000 1.945000 ;
      RECT 6.545000 2.285000  6.715000 2.745000 ;
      RECT 6.545000 2.745000  7.465000 2.915000 ;
      RECT 6.605000 1.245000  6.935000 1.325000 ;
      RECT 6.715000 0.255000  7.795000 0.425000 ;
      RECT 6.715000 0.425000  6.935000 0.725000 ;
      RECT 6.885000 1.945000  7.125000 2.575000 ;
      RECT 7.105000 0.595000  7.295000 1.495000 ;
      RECT 7.295000 1.835000  7.635000 2.065000 ;
      RECT 7.295000 2.065000  7.465000 2.745000 ;
      RECT 7.465000 0.425000  7.795000 1.095000 ;
      RECT 7.465000 1.275000  8.320000 1.445000 ;
      RECT 7.465000 1.445000  7.635000 1.835000 ;
      RECT 7.635000 2.235000  7.985000 3.075000 ;
      RECT 7.815000 1.635000  9.210000 1.805000 ;
      RECT 7.815000 1.805000  7.985000 2.235000 ;
      RECT 7.975000 0.335000  8.660000 0.665000 ;
      RECT 8.020000 0.845000  8.320000 1.275000 ;
      RECT 8.325000 1.975000  9.550000 2.155000 ;
      RECT 8.490000 0.665000  8.660000 1.135000 ;
      RECT 8.490000 1.135000  9.210000 1.635000 ;
      RECT 9.210000 0.255000  9.550000 0.895000 ;
      RECT 9.295000 2.155000  9.550000 2.905000 ;
      RECT 9.380000 0.895000  9.550000 1.345000 ;
      RECT 9.380000 1.345000 10.055000 1.675000 ;
      RECT 9.380000 1.675000  9.550000 1.975000 ;
    LAYER mcon ;
      RECT 2.555000 2.320000 2.725000 2.490000 ;
      RECT 4.955000 2.320000 5.125000 2.490000 ;
    LAYER met1 ;
      RECT 2.495000 2.290000 2.785000 2.335000 ;
      RECT 2.495000 2.335000 5.185000 2.475000 ;
      RECT 2.495000 2.475000 2.785000 2.520000 ;
      RECT 4.895000 2.290000 5.185000 2.335000 ;
      RECT 4.895000 2.475000 5.185000 2.520000 ;
  END
END sky130_fd_sc_lp__sdfxtp_2
