* File: sky130_fd_sc_lp__dfxbp_lp.pex.spice
* Created: Wed Sep  2 09:45:00 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__DFXBP_LP%CLK 3 5 7 8 10 11 12 18
c36 3 0 8.71038e-20 $X=0.54 $Y=2.515
r37 18 20 19.9686 $w=3.5e-07 $l=1.45e-07 $layer=POLY_cond $X=0.765 $Y=1.182
+ $X2=0.91 $Y2=1.182
r38 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.765
+ $Y=1.12 $X2=0.765 $Y2=1.12
r39 16 18 29.6086 $w=3.5e-07 $l=2.15e-07 $layer=POLY_cond $X=0.55 $Y=1.182
+ $X2=0.765 $Y2=1.182
r40 15 16 1.37714 $w=3.5e-07 $l=1e-08 $layer=POLY_cond $X=0.54 $Y=1.182 $X2=0.55
+ $Y2=1.182
r41 12 19 6.80989 $w=3.28e-07 $l=1.95e-07 $layer=LI1_cond $X=0.765 $Y=0.925
+ $X2=0.765 $Y2=1.12
r42 11 12 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.765 $Y=0.555
+ $X2=0.765 $Y2=0.925
r43 8 20 22.6286 $w=1.5e-07 $l=2.27e-07 $layer=POLY_cond $X=0.91 $Y=0.955
+ $X2=0.91 $Y2=1.182
r44 8 10 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.91 $Y=0.955
+ $X2=0.91 $Y2=0.635
r45 5 16 22.6286 $w=1.5e-07 $l=2.27e-07 $layer=POLY_cond $X=0.55 $Y=0.955
+ $X2=0.55 $Y2=1.182
r46 5 7 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.55 $Y=0.955 $X2=0.55
+ $Y2=0.635
r47 1 15 10.701 $w=2.5e-07 $l=2.28e-07 $layer=POLY_cond $X=0.54 $Y=1.41 $X2=0.54
+ $Y2=1.182
r48 1 3 274.541 $w=2.5e-07 $l=1.105e-06 $layer=POLY_cond $X=0.54 $Y=1.41
+ $X2=0.54 $Y2=2.515
.ends

.subckt PM_SKY130_FD_SC_LP__DFXBP_LP%D 3 7 10 11 15 17 18 25
r49 23 25 45.4639 $w=3.3e-07 $l=2.6e-07 $layer=POLY_cond $X=1.15 $Y=1.69
+ $X2=1.41 $Y2=1.69
r50 20 23 13.9889 $w=3.3e-07 $l=8e-08 $layer=POLY_cond $X=1.07 $Y=1.69 $X2=1.15
+ $Y2=1.69
r51 18 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.15
+ $Y=1.69 $X2=1.15 $Y2=1.69
r52 13 15 235.872 $w=1.5e-07 $l=4.6e-07 $layer=POLY_cond $X=1.77 $Y=1.095
+ $X2=1.77 $Y2=0.635
r53 12 17 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.485 $Y=1.17
+ $X2=1.41 $Y2=1.17
r54 11 13 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.695 $Y=1.17
+ $X2=1.77 $Y2=1.095
r55 11 12 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=1.695 $Y=1.17
+ $X2=1.485 $Y2=1.17
r56 10 25 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.41 $Y=1.525
+ $X2=1.41 $Y2=1.69
r57 9 17 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.41 $Y=1.245
+ $X2=1.41 $Y2=1.17
r58 9 10 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=1.41 $Y=1.245
+ $X2=1.41 $Y2=1.525
r59 5 17 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.41 $Y=1.095
+ $X2=1.41 $Y2=1.17
r60 5 7 235.872 $w=1.5e-07 $l=4.6e-07 $layer=POLY_cond $X=1.41 $Y=1.095 $X2=1.41
+ $Y2=0.635
r61 1 20 9.34494 $w=2.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.07 $Y=1.855
+ $X2=1.07 $Y2=1.69
r62 1 3 163.979 $w=2.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.07 $Y=1.855 $X2=1.07
+ $Y2=2.515
.ends

.subckt PM_SKY130_FD_SC_LP__DFXBP_LP%A_615_93# 1 2 3 4 13 15 16 18 20 21 26 29
+ 30 33 36 37 38 42 43 44 45 49 52 55 56 57 59 60
c177 59 0 1.31451e-19 $X=6.305 $Y=2.24
c178 45 0 1.66108e-19 $X=3.24 $Y=1.05
r179 60 63 10.4768 $w=3.28e-07 $l=3e-07 $layer=LI1_cond $X=7.435 $Y=0.7
+ $X2=7.435 $Y2=1
r180 55 57 8.3814 $w=3.83e-07 $l=2.8e-07 $layer=LI1_cond $X=4.587 $Y=1.92
+ $X2=4.587 $Y2=2.2
r181 55 56 8.58894 $w=3.83e-07 $l=1.65e-07 $layer=LI1_cond $X=4.587 $Y=1.92
+ $X2=4.587 $Y2=1.755
r182 48 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.24
+ $Y=1.29 $X2=3.24 $Y2=1.29
r183 45 48 8.3814 $w=3.28e-07 $l=2.4e-07 $layer=LI1_cond $X=3.24 $Y=1.05
+ $X2=3.24 $Y2=1.29
r184 43 60 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.27 $Y=0.7
+ $X2=7.435 $Y2=0.7
r185 43 44 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=7.27 $Y=0.7
+ $X2=6.74 $Y2=0.7
r186 41 44 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.655 $Y=0.785
+ $X2=6.74 $Y2=0.7
r187 41 42 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=6.655 $Y=0.785
+ $X2=6.655 $Y2=1.335
r188 37 42 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.57 $Y=1.42
+ $X2=6.655 $Y2=1.335
r189 37 38 71.1123 $w=1.68e-07 $l=1.09e-06 $layer=LI1_cond $X=6.57 $Y=1.42
+ $X2=5.48 $Y2=1.42
r190 36 38 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.395 $Y=1.335
+ $X2=5.48 $Y2=1.42
r191 35 36 58.7166 $w=1.68e-07 $l=9e-07 $layer=LI1_cond $X=5.395 $Y=0.435
+ $X2=5.395 $Y2=1.335
r192 34 57 5.54671 $w=1.7e-07 $l=1.93e-07 $layer=LI1_cond $X=4.78 $Y=2.2
+ $X2=4.587 $Y2=2.2
r193 33 59 4.95428 $w=1.7e-07 $l=1.74714e-07 $layer=LI1_cond $X=6.14 $Y=2.2
+ $X2=6.305 $Y2=2.18
r194 33 34 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=6.14 $Y=2.2
+ $X2=4.78 $Y2=2.2
r195 31 52 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.695 $Y=1.135
+ $X2=4.695 $Y2=1.05
r196 31 56 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=4.695 $Y=1.135
+ $X2=4.695 $Y2=1.755
r197 29 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.31 $Y=0.35
+ $X2=5.395 $Y2=0.435
r198 29 30 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=5.31 $Y=0.35
+ $X2=4.48 $Y2=0.35
r199 24 52 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=4.315 $Y=1.05
+ $X2=4.695 $Y2=1.05
r200 24 26 5.5876 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=4.315 $Y=0.965
+ $X2=4.315 $Y2=0.805
r201 23 30 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.315 $Y=0.435
+ $X2=4.48 $Y2=0.35
r202 23 26 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=4.315 $Y=0.435
+ $X2=4.315 $Y2=0.805
r203 22 45 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.405 $Y=1.05
+ $X2=3.24 $Y2=1.05
r204 21 24 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=4.15 $Y=1.05
+ $X2=4.315 $Y2=1.05
r205 21 22 48.6043 $w=1.68e-07 $l=7.45e-07 $layer=LI1_cond $X=4.15 $Y=1.05
+ $X2=3.405 $Y2=1.05
r206 18 20 110.86 $w=2.5e-07 $l=5.75e-07 $layer=POLY_cond $X=3.765 $Y=1.66
+ $X2=3.765 $Y2=2.235
r207 17 49 54.4789 $w=2.61e-07 $l=3.68375e-07 $layer=POLY_cond $X=3.405 $Y=1.585
+ $X2=3.24 $Y2=1.29
r208 16 18 29.1797 $w=1.5e-07 $l=1.58114e-07 $layer=POLY_cond $X=3.64 $Y=1.585
+ $X2=3.765 $Y2=1.66
r209 16 17 120.5 $w=1.5e-07 $l=2.35e-07 $layer=POLY_cond $X=3.64 $Y=1.585
+ $X2=3.405 $Y2=1.585
r210 13 49 39.116 $w=2.61e-07 $l=2.05122e-07 $layer=POLY_cond $X=3.15 $Y=1.125
+ $X2=3.24 $Y2=1.29
r211 13 15 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=3.15 $Y=1.125
+ $X2=3.15 $Y2=0.805
r212 4 59 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=6.16
+ $Y=2.095 $X2=6.305 $Y2=2.24
r213 3 55 300 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_PDIFF $count=2 $X=4.42
+ $Y=1.735 $X2=4.56 $Y2=1.92
r214 2 63 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=7.295
+ $Y=0.855 $X2=7.435 $Y2=1
r215 1 26 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=4.175
+ $Y=0.595 $X2=4.315 $Y2=0.805
.ends

.subckt PM_SKY130_FD_SC_LP__DFXBP_LP%A_455_85# 1 2 7 9 10 11 12 14 15 17 19 21
+ 23 28
c90 17 0 2.19317e-19 $X=4.295 $Y=2.235
c91 7 0 1.66108e-19 $X=3.74 $Y=1.12
r92 29 31 29.274 $w=3.54e-07 $l=2.15e-07 $layer=POLY_cond $X=4.227 $Y=1.41
+ $X2=4.227 $Y2=1.195
r93 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.265
+ $Y=1.41 $X2=4.265 $Y2=1.41
r94 24 26 4.29183 $w=1.7e-07 $l=2.07485e-07 $layer=LI1_cond $X=2.66 $Y=1.72
+ $X2=2.455 $Y2=1.725
r95 23 28 13.3169 $w=2.84e-07 $l=3.94487e-07 $layer=LI1_cond $X=4.045 $Y=1.72
+ $X2=4.237 $Y2=1.41
r96 23 24 90.3583 $w=1.68e-07 $l=1.385e-06 $layer=LI1_cond $X=4.045 $Y=1.72
+ $X2=2.66 $Y2=1.72
r97 19 26 3.47434 $w=3.3e-07 $l=1.48661e-07 $layer=LI1_cond $X=2.495 $Y=1.595
+ $X2=2.455 $Y2=1.725
r98 19 21 30.5572 $w=3.28e-07 $l=8.75e-07 $layer=LI1_cond $X=2.495 $Y=1.595
+ $X2=2.495 $Y2=0.72
r99 15 29 26.6882 $w=3.54e-07 $l=1.96074e-07 $layer=POLY_cond $X=4.295 $Y=1.575
+ $X2=4.227 $Y2=1.41
r100 15 17 163.979 $w=2.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.295 $Y=1.575
+ $X2=4.295 $Y2=2.235
r101 12 31 26.5778 $w=3.54e-07 $l=1.60169e-07 $layer=POLY_cond $X=4.1 $Y=1.12
+ $X2=4.227 $Y2=1.195
r102 12 14 101.22 $w=1.5e-07 $l=3.15e-07 $layer=POLY_cond $X=4.1 $Y=1.12 $X2=4.1
+ $Y2=0.805
r103 10 31 22.9014 $w=1.5e-07 $l=2.02e-07 $layer=POLY_cond $X=4.025 $Y=1.195
+ $X2=4.227 $Y2=1.195
r104 10 11 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=4.025 $Y=1.195
+ $X2=3.815 $Y2=1.195
r105 7 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.74 $Y=1.12
+ $X2=3.815 $Y2=1.195
r106 7 9 101.22 $w=1.5e-07 $l=3.15e-07 $layer=POLY_cond $X=3.74 $Y=1.12 $X2=3.74
+ $Y2=0.805
r107 2 26 600 $w=1.7e-07 $l=2.08567e-07 $layer=licon1_PDIFF $count=1 $X=2.275
+ $Y=1.615 $X2=2.415 $Y2=1.765
r108 1 21 182 $w=1.7e-07 $l=3.89776e-07 $layer=licon1_NDIFF $count=1 $X=2.275
+ $Y=0.425 $X2=2.495 $Y2=0.72
.ends

.subckt PM_SKY130_FD_SC_LP__DFXBP_LP%A_27_403# 1 2 7 10 13 15 17 19 20 21 22 24
+ 25 27 29 30 33 34 38 42 45 46 47 48 51 54 56 59 61 64 65 67 68 71
c174 65 0 8.71038e-20 $X=1.32 $Y=2.92
c175 33 0 9.24756e-20 $X=5.95 $Y=3.075
c176 29 0 1.49367e-19 $X=5.53 $Y=1.48
c177 25 0 1.36058e-19 $X=5.53 $Y=1.12
c178 20 0 8.93026e-20 $X=5.455 $Y=1.195
r179 68 73 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=2.15 $Y=2.94
+ $X2=2.15 $Y2=3.15
r180 67 68 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.15
+ $Y=2.94 $X2=2.15 $Y2=2.94
r181 65 67 32.9837 $w=2.88e-07 $l=8.3e-07 $layer=LI1_cond $X=1.32 $Y=2.92
+ $X2=2.15 $Y2=2.92
r182 64 65 7.43784 $w=2.9e-07 $l=1.8262e-07 $layer=LI1_cond $X=1.235 $Y=2.775
+ $X2=1.32 $Y2=2.92
r183 63 64 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=1.235 $Y=2.595
+ $X2=1.235 $Y2=2.775
r184 62 71 3.80956 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.44 $Y=2.51
+ $X2=0.275 $Y2=2.51
r185 61 63 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.15 $Y=2.51
+ $X2=1.235 $Y2=2.595
r186 61 62 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=1.15 $Y=2.51
+ $X2=0.44 $Y2=2.51
r187 57 71 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.275 $Y=2.595
+ $X2=0.275 $Y2=2.51
r188 57 59 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=0.275 $Y=2.595
+ $X2=0.275 $Y2=2.87
r189 56 70 5.81909 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.275 $Y=2.16
+ $X2=0.275 $Y2=1.995
r190 54 71 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.275 $Y=2.425
+ $X2=0.275 $Y2=2.51
r191 54 56 9.25447 $w=3.28e-07 $l=2.65e-07 $layer=LI1_cond $X=0.275 $Y=2.425
+ $X2=0.275 $Y2=2.16
r192 51 70 50.5588 $w=3.08e-07 $l=1.36e-06 $layer=LI1_cond $X=0.265 $Y=0.635
+ $X2=0.265 $Y2=1.995
r193 40 48 15.9654 $w=2e-07 $l=9.68246e-08 $layer=POLY_cond $X=6.62 $Y=1.48
+ $X2=6.57 $Y2=1.555
r194 40 42 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=6.62 $Y=1.48
+ $X2=6.62 $Y2=0.975
r195 36 48 15.9654 $w=2e-07 $l=7.5e-08 $layer=POLY_cond $X=6.57 $Y=1.63 $X2=6.57
+ $Y2=1.555
r196 36 38 239.758 $w=2.5e-07 $l=9.65e-07 $layer=POLY_cond $X=6.57 $Y=1.63
+ $X2=6.57 $Y2=2.595
r197 35 47 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=6.025 $Y=1.555
+ $X2=5.95 $Y2=1.555
r198 34 48 9.46703 $w=1.5e-07 $l=1.25e-07 $layer=POLY_cond $X=6.445 $Y=1.555
+ $X2=6.57 $Y2=1.555
r199 34 35 215.362 $w=1.5e-07 $l=4.2e-07 $layer=POLY_cond $X=6.445 $Y=1.555
+ $X2=6.025 $Y2=1.555
r200 32 47 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.95 $Y=1.63
+ $X2=5.95 $Y2=1.555
r201 32 33 740.947 $w=1.5e-07 $l=1.445e-06 $layer=POLY_cond $X=5.95 $Y=1.63
+ $X2=5.95 $Y2=3.075
r202 31 45 9.46703 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=5.605 $Y=1.555
+ $X2=5.435 $Y2=1.555
r203 30 47 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.875 $Y=1.555
+ $X2=5.95 $Y2=1.555
r204 30 31 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=5.875 $Y=1.555
+ $X2=5.605 $Y2=1.555
r205 29 45 15.9654 $w=2e-07 $l=1.27083e-07 $layer=POLY_cond $X=5.53 $Y=1.48
+ $X2=5.435 $Y2=1.555
r206 28 46 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.53 $Y=1.27
+ $X2=5.53 $Y2=1.195
r207 28 29 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=5.53 $Y=1.27
+ $X2=5.53 $Y2=1.48
r208 25 46 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.53 $Y=1.12
+ $X2=5.53 $Y2=1.195
r209 25 27 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=5.53 $Y=1.12
+ $X2=5.53 $Y2=0.835
r210 22 45 15.9654 $w=2e-07 $l=9.48683e-08 $layer=POLY_cond $X=5.39 $Y=1.63
+ $X2=5.435 $Y2=1.555
r211 22 24 110.86 $w=2.5e-07 $l=5.75e-07 $layer=POLY_cond $X=5.39 $Y=1.63
+ $X2=5.39 $Y2=2.205
r212 20 46 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=5.455 $Y=1.195
+ $X2=5.53 $Y2=1.195
r213 20 21 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=5.455 $Y=1.195
+ $X2=5.245 $Y2=1.195
r214 17 21 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.17 $Y=1.12
+ $X2=5.245 $Y2=1.195
r215 17 19 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=5.17 $Y=1.12
+ $X2=5.17 $Y2=0.835
r216 16 73 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.315 $Y=3.15
+ $X2=2.15 $Y2=3.15
r217 15 33 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.875 $Y=3.15
+ $X2=5.95 $Y2=3.075
r218 15 16 1825.45 $w=1.5e-07 $l=3.56e-06 $layer=POLY_cond $X=5.875 $Y=3.15
+ $X2=2.315 $Y2=3.15
r219 13 44 435.851 $w=1.5e-07 $l=8.5e-07 $layer=POLY_cond $X=2.2 $Y=0.635
+ $X2=2.2 $Y2=1.485
r220 8 68 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.15 $Y=2.775
+ $X2=2.15 $Y2=2.94
r221 8 10 163.979 $w=2.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.15 $Y=2.775
+ $X2=2.15 $Y2=2.115
r222 7 44 40.9178 $w=2.5e-07 $l=1.25e-07 $layer=POLY_cond $X=2.15 $Y=1.61
+ $X2=2.15 $Y2=1.485
r223 7 10 125.469 $w=2.5e-07 $l=5.05e-07 $layer=POLY_cond $X=2.15 $Y=1.61
+ $X2=2.15 $Y2=2.115
r224 2 59 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.015 $X2=0.275 $Y2=2.87
r225 2 56 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.015 $X2=0.275 $Y2=2.16
r226 1 51 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.19
+ $Y=0.425 $X2=0.335 $Y2=0.635
.ends

.subckt PM_SKY130_FD_SC_LP__DFXBP_LP%A_511_218# 1 2 9 14 15 16 19 24 26 28 34 40
+ 42 43 44
c121 44 0 8.93026e-20 $X=6.935 $Y=1.775
c122 34 0 1.36058e-19 $X=5.045 $Y=0.7
c123 28 0 1.49367e-19 $X=5.045 $Y=1.685
c124 19 0 1.31451e-19 $X=7.1 $Y=2.595
c125 9 0 1.6807e-19 $X=2.68 $Y=2.115
r126 43 48 31.8923 $w=3.6e-07 $l=1.65e-07 $layer=POLY_cond $X=7.115 $Y=1.77
+ $X2=7.115 $Y2=1.935
r127 43 47 46.5827 $w=3.6e-07 $l=1.65e-07 $layer=POLY_cond $X=7.115 $Y=1.77
+ $X2=7.115 $Y2=1.605
r128 42 44 8.46025 $w=3.18e-07 $l=1.65e-07 $layer=LI1_cond $X=7.1 $Y=1.775
+ $X2=6.935 $Y2=1.775
r129 42 43 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.1
+ $Y=1.77 $X2=7.1 $Y2=1.77
r130 40 44 107.321 $w=1.68e-07 $l=1.645e-06 $layer=LI1_cond $X=5.29 $Y=1.77
+ $X2=6.935 $Y2=1.77
r131 39 40 8.79328 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=5.125 $Y=1.81
+ $X2=5.29 $Y2=1.81
r132 36 39 3.68782 $w=2.48e-07 $l=8e-08 $layer=LI1_cond $X=5.045 $Y=1.81
+ $X2=5.125 $Y2=1.81
r133 32 34 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=4.875 $Y=0.7
+ $X2=5.045 $Y2=0.7
r134 28 36 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.045 $Y=1.685
+ $X2=5.045 $Y2=1.81
r135 27 34 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.045 $Y=0.785
+ $X2=5.045 $Y2=0.7
r136 27 28 58.7166 $w=1.68e-07 $l=9e-07 $layer=LI1_cond $X=5.045 $Y=0.785
+ $X2=5.045 $Y2=1.685
r137 25 26 47.1291 $w=2.5e-07 $l=1.5e-07 $layer=POLY_cond $X=2.71 $Y=1.09
+ $X2=2.71 $Y2=1.24
r138 24 47 276.894 $w=1.5e-07 $l=5.4e-07 $layer=POLY_cond $X=7.22 $Y=1.065
+ $X2=7.22 $Y2=1.605
r139 21 24 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=7.22 $Y=0.255
+ $X2=7.22 $Y2=1.065
r140 19 48 163.979 $w=2.5e-07 $l=6.6e-07 $layer=POLY_cond $X=7.1 $Y=2.595
+ $X2=7.1 $Y2=1.935
r141 15 21 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.145 $Y=0.18
+ $X2=7.22 $Y2=0.255
r142 15 16 2194.64 $w=1.5e-07 $l=4.28e-06 $layer=POLY_cond $X=7.145 $Y=0.18
+ $X2=2.865 $Y2=0.18
r143 14 25 146.138 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.79 $Y=0.805
+ $X2=2.79 $Y2=1.09
r144 11 16 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.79 $Y=0.255
+ $X2=2.865 $Y2=0.18
r145 11 14 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=2.79 $Y=0.255
+ $X2=2.79 $Y2=0.805
r146 9 26 217.397 $w=2.5e-07 $l=8.75e-07 $layer=POLY_cond $X=2.68 $Y=2.115
+ $X2=2.68 $Y2=1.24
r147 2 39 600 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=4.98
+ $Y=1.705 $X2=5.125 $Y2=1.85
r148 1 32 182 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=1 $X=4.73
+ $Y=0.555 $X2=4.875 $Y2=0.7
.ends

.subckt PM_SKY130_FD_SC_LP__DFXBP_LP%A_1507_321# 1 2 9 12 13 15 18 22 26 30 34
+ 38 42 46 49 50 53 56 57 62 68 69 71 76 78 80 86
c149 38 0 1.1898e-19 $X=11.125 $Y=0.845
c150 13 0 1.1902e-19 $X=8.205 $Y=0.78
r151 95 96 62.9501 $w=3.3e-07 $l=3.6e-07 $layer=POLY_cond $X=10.765 $Y=1.42
+ $X2=11.125 $Y2=1.42
r152 90 91 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=9.975 $Y=1.42
+ $X2=10.185 $Y2=1.42
r153 88 90 55.9556 $w=3.3e-07 $l=3.2e-07 $layer=POLY_cond $X=9.655 $Y=1.42
+ $X2=9.975 $Y2=1.42
r154 80 96 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=11.2 $Y=1.42
+ $X2=11.125 $Y2=1.42
r155 79 93 16.6118 $w=3.3e-07 $l=9.5e-08 $layer=POLY_cond $X=10.24 $Y=1.42
+ $X2=10.335 $Y2=1.42
r156 79 91 9.61737 $w=3.3e-07 $l=5.5e-08 $layer=POLY_cond $X=10.24 $Y=1.42
+ $X2=10.185 $Y2=1.42
r157 78 79 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=10.24
+ $Y=1.42 $X2=10.24 $Y2=1.42
r158 75 76 9.2801 $w=4.58e-07 $l=1.65e-07 $layer=LI1_cond $X=9.21 $Y=0.495
+ $X2=9.375 $Y2=0.495
r159 72 75 6.50043 $w=4.58e-07 $l=2.5e-07 $layer=LI1_cond $X=8.96 $Y=0.495
+ $X2=9.21 $Y2=0.495
r160 69 80 69.9445 $w=3.3e-07 $l=4e-07 $layer=POLY_cond $X=11.6 $Y=1.42 $X2=11.2
+ $Y2=1.42
r161 68 69 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=11.6
+ $Y=1.42 $X2=11.6 $Y2=1.42
r162 66 95 32.3493 $w=3.3e-07 $l=1.85e-07 $layer=POLY_cond $X=10.58 $Y=1.42
+ $X2=10.765 $Y2=1.42
r163 66 93 42.841 $w=3.3e-07 $l=2.45e-07 $layer=POLY_cond $X=10.58 $Y=1.42
+ $X2=10.335 $Y2=1.42
r164 65 68 35.621 $w=3.28e-07 $l=1.02e-06 $layer=LI1_cond $X=10.58 $Y=1.42
+ $X2=11.6 $Y2=1.42
r165 65 66 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=10.58
+ $Y=1.42 $X2=10.58 $Y2=1.42
r166 63 78 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.275 $Y=1.42
+ $X2=10.19 $Y2=1.42
r167 63 65 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=10.275 $Y=1.42
+ $X2=10.58 $Y2=1.42
r168 62 78 3.80956 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.19 $Y=1.255
+ $X2=10.19 $Y2=1.42
r169 61 62 53.4973 $w=1.68e-07 $l=8.2e-07 $layer=LI1_cond $X=10.19 $Y=0.435
+ $X2=10.19 $Y2=1.255
r170 57 61 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.105 $Y=0.35
+ $X2=10.19 $Y2=0.435
r171 57 76 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=10.105 $Y=0.35
+ $X2=9.375 $Y2=0.35
r172 56 71 3.03453 $w=3.12e-07 $l=1.80566e-07 $layer=LI1_cond $X=8.96 $Y=2.02
+ $X2=8.817 $Y2=2.105
r173 55 72 6.6364 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=8.96 $Y=0.725
+ $X2=8.96 $Y2=0.495
r174 55 56 84.4866 $w=1.68e-07 $l=1.295e-06 $layer=LI1_cond $X=8.96 $Y=0.725
+ $X2=8.96 $Y2=2.02
r175 51 71 3.03453 $w=3.12e-07 $l=8.5e-08 $layer=LI1_cond $X=8.817 $Y=2.19
+ $X2=8.817 $Y2=2.105
r176 51 53 1.31437 $w=4.53e-07 $l=5e-08 $layer=LI1_cond $X=8.817 $Y=2.19
+ $X2=8.817 $Y2=2.24
r177 49 71 3.60271 $w=1.7e-07 $l=2.27e-07 $layer=LI1_cond $X=8.59 $Y=2.105
+ $X2=8.817 $Y2=2.105
r178 49 50 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=8.59 $Y=2.105
+ $X2=8.125 $Y2=2.105
r179 47 86 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=7.96 $Y=1.77 $X2=8.05
+ $Y2=1.77
r180 47 83 52.4584 $w=3.3e-07 $l=3e-07 $layer=POLY_cond $X=7.96 $Y=1.77 $X2=7.66
+ $Y2=1.77
r181 46 47 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.96
+ $Y=1.77 $X2=7.96 $Y2=1.77
r182 44 50 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=7.96 $Y=2.02
+ $X2=8.125 $Y2=2.105
r183 44 46 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=7.96 $Y=2.02
+ $X2=7.96 $Y2=1.77
r184 40 42 79.4787 $w=1.5e-07 $l=1.55e-07 $layer=POLY_cond $X=8.05 $Y=0.855
+ $X2=8.205 $Y2=0.855
r185 36 96 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=11.125 $Y=1.255
+ $X2=11.125 $Y2=1.42
r186 36 38 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=11.125 $Y=1.255
+ $X2=11.125 $Y2=0.845
r187 32 95 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.765 $Y=1.255
+ $X2=10.765 $Y2=1.42
r188 32 34 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=10.765 $Y=1.255
+ $X2=10.765 $Y2=0.845
r189 28 93 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.335 $Y=1.255
+ $X2=10.335 $Y2=1.42
r190 28 30 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=10.335 $Y=1.255
+ $X2=10.335 $Y2=0.845
r191 24 91 9.34494 $w=2.5e-07 $l=1.65e-07 $layer=POLY_cond $X=10.185 $Y=1.585
+ $X2=10.185 $Y2=1.42
r192 24 26 186.34 $w=2.5e-07 $l=7.5e-07 $layer=POLY_cond $X=10.185 $Y=1.585
+ $X2=10.185 $Y2=2.335
r193 20 90 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.975 $Y=1.255
+ $X2=9.975 $Y2=1.42
r194 20 22 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=9.975 $Y=1.255
+ $X2=9.975 $Y2=0.845
r195 16 88 9.34494 $w=2.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.655 $Y=1.585
+ $X2=9.655 $Y2=1.42
r196 16 18 186.34 $w=2.5e-07 $l=7.5e-07 $layer=POLY_cond $X=9.655 $Y=1.585
+ $X2=9.655 $Y2=2.335
r197 13 42 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.205 $Y=0.78
+ $X2=8.205 $Y2=0.855
r198 13 15 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=8.205 $Y=0.78
+ $X2=8.205 $Y2=0.495
r199 12 86 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.05 $Y=1.605
+ $X2=8.05 $Y2=1.77
r200 11 40 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.05 $Y=0.93
+ $X2=8.05 $Y2=0.855
r201 11 12 346.117 $w=1.5e-07 $l=6.75e-07 $layer=POLY_cond $X=8.05 $Y=0.93
+ $X2=8.05 $Y2=1.605
r202 7 83 9.34494 $w=2.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.66 $Y=1.935
+ $X2=7.66 $Y2=1.77
r203 7 9 163.979 $w=2.5e-07 $l=6.6e-07 $layer=POLY_cond $X=7.66 $Y=1.935
+ $X2=7.66 $Y2=2.595
r204 2 53 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=8.615
+ $Y=2.095 $X2=8.755 $Y2=2.24
r205 1 75 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=9.07
+ $Y=0.285 $X2=9.21 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__DFXBP_LP%A_1339_153# 1 2 9 13 15 19 22 24 29 31 33
+ 34 36 37 42 43 45 46
c103 42 0 9.24756e-20 $X=6.835 $Y=2.28
c104 13 0 1.69058e-19 $X=8.635 $Y=0.495
r105 45 46 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=8.53
+ $Y=1.335 $X2=8.53 $Y2=1.335
r106 38 43 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.615 $Y=1.35
+ $X2=7.53 $Y2=1.35
r107 37 45 4.78091 $w=1.7e-07 $l=1.8747e-07 $layer=LI1_cond $X=8.365 $Y=1.35
+ $X2=8.53 $Y2=1.302
r108 37 38 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=8.365 $Y=1.35
+ $X2=7.615 $Y2=1.35
r109 35 43 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.53 $Y=1.435
+ $X2=7.53 $Y2=1.35
r110 35 36 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=7.53 $Y=1.435
+ $X2=7.53 $Y2=2.115
r111 33 43 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.445 $Y=1.35
+ $X2=7.53 $Y2=1.35
r112 33 34 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=7.445 $Y=1.35
+ $X2=7.09 $Y2=1.35
r113 32 42 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7 $Y=2.2 $X2=6.835
+ $Y2=2.2
r114 31 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.445 $Y=2.2
+ $X2=7.53 $Y2=2.115
r115 31 32 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=7.445 $Y=2.2 $X2=7
+ $Y2=2.2
r116 27 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.005 $Y=1.265
+ $X2=7.09 $Y2=1.35
r117 27 29 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=7.005 $Y=1.265
+ $X2=7.005 $Y2=1.13
r118 23 46 55.6971 $w=3.45e-07 $l=3.33e-07 $layer=POLY_cond $X=8.537 $Y=1.668
+ $X2=8.537 $Y2=1.335
r119 23 24 33.2433 $w=3.45e-07 $l=1.72e-07 $layer=POLY_cond $X=8.537 $Y=1.668
+ $X2=8.537 $Y2=1.84
r120 21 46 2.50888 $w=3.45e-07 $l=1.5e-08 $layer=POLY_cond $X=8.537 $Y=1.32
+ $X2=8.537 $Y2=1.335
r121 21 22 13.218 $w=2.47e-07 $l=7.5e-08 $layer=POLY_cond $X=8.537 $Y=1.32
+ $X2=8.537 $Y2=1.245
r122 17 19 346.117 $w=1.5e-07 $l=6.75e-07 $layer=POLY_cond $X=8.995 $Y=1.17
+ $X2=8.995 $Y2=0.495
r123 16 22 12.6197 $w=1.5e-07 $l=1.73e-07 $layer=POLY_cond $X=8.71 $Y=1.245
+ $X2=8.537 $Y2=1.245
r124 15 17 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.92 $Y=1.245
+ $X2=8.995 $Y2=1.17
r125 15 16 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=8.92 $Y=1.245
+ $X2=8.71 $Y2=1.245
r126 11 22 13.218 $w=2.47e-07 $l=1.30208e-07 $layer=POLY_cond $X=8.635 $Y=1.17
+ $X2=8.537 $Y2=1.245
r127 11 13 346.117 $w=1.5e-07 $l=6.75e-07 $layer=POLY_cond $X=8.635 $Y=1.17
+ $X2=8.635 $Y2=0.495
r128 9 24 187.582 $w=2.5e-07 $l=7.55e-07 $layer=POLY_cond $X=8.49 $Y=2.595
+ $X2=8.49 $Y2=1.84
r129 2 42 300 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_PDIFF $count=2 $X=6.695
+ $Y=2.095 $X2=6.835 $Y2=2.28
r130 1 29 182 $w=1.7e-07 $l=4.96362e-07 $layer=licon1_NDIFF $count=1 $X=6.695
+ $Y=0.765 $X2=7.005 $Y2=1.13
.ends

.subckt PM_SKY130_FD_SC_LP__DFXBP_LP%A_2062_367# 1 2 9 11 13 16 20 21 24 28 29
+ 30 37 38 40 44
c62 30 0 1.1898e-19 $X=12.005 $Y=0.99
c63 20 0 9.72338e-20 $X=12.272 $Y=1.365
r64 40 42 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=11.34 $Y=0.845
+ $X2=11.34 $Y2=0.99
r65 37 44 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=12.17 $Y=1.38
+ $X2=12.17 $Y2=1.215
r66 37 38 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=12.17
+ $Y=1.38 $X2=12.17 $Y2=1.38
r67 35 37 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=12.17 $Y=1.765
+ $X2=12.17 $Y2=1.38
r68 32 44 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=12.09 $Y=1.075
+ $X2=12.09 $Y2=1.215
r69 31 42 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.505 $Y=0.99
+ $X2=11.34 $Y2=0.99
r70 30 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=12.005 $Y=0.99
+ $X2=12.09 $Y2=1.075
r71 30 31 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=12.005 $Y=0.99
+ $X2=11.505 $Y2=0.99
r72 28 35 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=12.005 $Y=1.85
+ $X2=12.17 $Y2=1.765
r73 28 29 90.6845 $w=1.68e-07 $l=1.39e-06 $layer=LI1_cond $X=12.005 $Y=1.85
+ $X2=10.615 $Y2=1.85
r74 24 26 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=10.45 $Y=1.98
+ $X2=10.45 $Y2=2.69
r75 22 29 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=10.45 $Y=1.935
+ $X2=10.615 $Y2=1.85
r76 22 24 1.57151 $w=3.28e-07 $l=4.5e-08 $layer=LI1_cond $X=10.45 $Y=1.935
+ $X2=10.45 $Y2=1.98
r77 21 38 36.8212 $w=4.35e-07 $l=2.88e-07 $layer=POLY_cond $X=12.222 $Y=1.668
+ $X2=12.222 $Y2=1.38
r78 20 38 1.91777 $w=4.35e-07 $l=1.5e-08 $layer=POLY_cond $X=12.222 $Y=1.365
+ $X2=12.222 $Y2=1.38
r79 11 21 44.9166 $w=3.67e-07 $l=4.2775e-07 $layer=POLY_cond $X=12.415 $Y=2.01
+ $X2=12.222 $Y2=1.668
r80 11 13 103.148 $w=2.5e-07 $l=5.35e-07 $layer=POLY_cond $X=12.415 $Y=2.01
+ $X2=12.415 $Y2=2.545
r81 7 20 24.5823 $w=4.35e-07 $l=1.5e-07 $layer=POLY_cond $X=12.272 $Y=1.215
+ $X2=12.272 $Y2=1.365
r82 7 16 369.191 $w=1.5e-07 $l=7.2e-07 $layer=POLY_cond $X=12.465 $Y=1.215
+ $X2=12.465 $Y2=0.495
r83 7 9 369.191 $w=1.5e-07 $l=7.2e-07 $layer=POLY_cond $X=12.105 $Y=1.215
+ $X2=12.105 $Y2=0.495
r84 2 26 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=10.31
+ $Y=1.835 $X2=10.45 $Y2=2.69
r85 2 24 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=10.31
+ $Y=1.835 $X2=10.45 $Y2=1.98
r86 1 40 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=11.2
+ $Y=0.635 $X2=11.34 $Y2=0.845
.ends

.subckt PM_SKY130_FD_SC_LP__DFXBP_LP%VPWR 1 2 3 4 5 6 23 27 31 35 39 45 48 49 50
+ 52 60 65 73 89 90 93 96 99 102 105
r120 105 106 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.84 $Y=3.33
+ $X2=9.84 $Y2=3.33
r121 102 103 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r122 99 100 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r123 96 97 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r124 93 94 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r125 89 90 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=12.72 $Y=3.33
+ $X2=12.72 $Y2=3.33
r126 87 90 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=11.76 $Y=3.33
+ $X2=12.72 $Y2=3.33
r127 86 87 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.76 $Y=3.33
+ $X2=11.76 $Y2=3.33
r128 84 87 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=10.32 $Y=3.33
+ $X2=11.76 $Y2=3.33
r129 84 106 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=3.33
+ $X2=9.84 $Y2=3.33
r130 83 86 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=10.32 $Y=3.33
+ $X2=11.76 $Y2=3.33
r131 83 84 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.32 $Y=3.33
+ $X2=10.32 $Y2=3.33
r132 81 105 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.085 $Y=3.33
+ $X2=9.92 $Y2=3.33
r133 81 83 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=10.085 $Y=3.33
+ $X2=10.32 $Y2=3.33
r134 80 106 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=9.36 $Y=3.33
+ $X2=9.84 $Y2=3.33
r135 79 80 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=9.36 $Y=3.33
+ $X2=9.36 $Y2=3.33
r136 77 80 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=9.36 $Y2=3.33
r137 77 103 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=7.92 $Y2=3.33
r138 76 79 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=8.4 $Y=3.33 $X2=9.36
+ $Y2=3.33
r139 76 77 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.4 $Y=3.33
+ $X2=8.4 $Y2=3.33
r140 74 102 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.125 $Y=3.33
+ $X2=7.96 $Y2=3.33
r141 74 76 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=8.125 $Y=3.33
+ $X2=8.4 $Y2=3.33
r142 73 105 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.755 $Y=3.33
+ $X2=9.92 $Y2=3.33
r143 73 79 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=9.755 $Y=3.33
+ $X2=9.36 $Y2=3.33
r144 72 103 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=7.92 $Y2=3.33
r145 71 72 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r146 69 100 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33
+ $X2=5.52 $Y2=3.33
r147 68 71 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=6 $Y=3.33 $X2=7.44
+ $Y2=3.33
r148 68 69 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r149 66 99 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.82 $Y=3.33
+ $X2=5.655 $Y2=3.33
r150 66 68 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=5.82 $Y=3.33 $X2=6
+ $Y2=3.33
r151 65 102 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.795 $Y=3.33
+ $X2=7.96 $Y2=3.33
r152 65 71 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=7.795 $Y=3.33
+ $X2=7.44 $Y2=3.33
r153 64 100 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.52 $Y2=3.33
r154 64 97 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=4.08 $Y2=3.33
r155 63 64 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r156 61 96 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.195 $Y=3.33
+ $X2=4.03 $Y2=3.33
r157 61 63 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=4.195 $Y=3.33
+ $X2=4.56 $Y2=3.33
r158 60 99 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.49 $Y=3.33
+ $X2=5.655 $Y2=3.33
r159 60 63 60.6738 $w=1.68e-07 $l=9.3e-07 $layer=LI1_cond $X=5.49 $Y=3.33
+ $X2=4.56 $Y2=3.33
r160 59 97 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r161 58 59 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r162 56 59 0.668963 $w=4.9e-07 $l=2.4e-06 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=3.6 $Y2=3.33
r163 56 94 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r164 55 58 156.578 $w=1.68e-07 $l=2.4e-06 $layer=LI1_cond $X=1.2 $Y=3.33 $X2=3.6
+ $Y2=3.33
r165 55 56 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r166 53 93 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.97 $Y=3.33
+ $X2=0.805 $Y2=3.33
r167 53 55 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=0.97 $Y=3.33
+ $X2=1.2 $Y2=3.33
r168 52 96 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.865 $Y=3.33
+ $X2=4.03 $Y2=3.33
r169 52 58 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=3.865 $Y=3.33
+ $X2=3.6 $Y2=3.33
r170 50 72 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6.48 $Y=3.33
+ $X2=7.44 $Y2=3.33
r171 50 69 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33 $X2=6
+ $Y2=3.33
r172 48 86 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=11.985 $Y=3.33
+ $X2=11.76 $Y2=3.33
r173 48 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.985 $Y=3.33
+ $X2=12.15 $Y2=3.33
r174 47 89 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=12.315 $Y=3.33
+ $X2=12.72 $Y2=3.33
r175 47 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.315 $Y=3.33
+ $X2=12.15 $Y2=3.33
r176 43 49 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=12.15 $Y=3.245
+ $X2=12.15 $Y2=3.33
r177 43 45 33.7002 $w=3.28e-07 $l=9.65e-07 $layer=LI1_cond $X=12.15 $Y=3.245
+ $X2=12.15 $Y2=2.28
r178 39 42 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=9.92 $Y=1.98
+ $X2=9.92 $Y2=2.69
r179 37 105 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.92 $Y=3.245
+ $X2=9.92 $Y2=3.33
r180 37 42 19.382 $w=3.28e-07 $l=5.55e-07 $layer=LI1_cond $X=9.92 $Y=3.245
+ $X2=9.92 $Y2=2.69
r181 33 102 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.96 $Y=3.245
+ $X2=7.96 $Y2=3.33
r182 33 35 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=7.96 $Y=3.245
+ $X2=7.96 $Y2=2.535
r183 29 99 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.655 $Y=3.245
+ $X2=5.655 $Y2=3.33
r184 29 31 24.0965 $w=3.28e-07 $l=6.9e-07 $layer=LI1_cond $X=5.655 $Y=3.245
+ $X2=5.655 $Y2=2.555
r185 25 96 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.03 $Y=3.245
+ $X2=4.03 $Y2=3.33
r186 25 27 38.2402 $w=3.28e-07 $l=1.095e-06 $layer=LI1_cond $X=4.03 $Y=3.245
+ $X2=4.03 $Y2=2.15
r187 21 93 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.805 $Y=3.245
+ $X2=0.805 $Y2=3.33
r188 21 23 13.2706 $w=3.28e-07 $l=3.8e-07 $layer=LI1_cond $X=0.805 $Y=3.245
+ $X2=0.805 $Y2=2.865
r189 6 45 300 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_PDIFF $count=2 $X=12.005
+ $Y=2.045 $X2=12.15 $Y2=2.28
r190 5 42 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=9.78
+ $Y=1.835 $X2=9.92 $Y2=2.69
r191 5 39 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=9.78
+ $Y=1.835 $X2=9.92 $Y2=1.98
r192 4 35 300 $w=1.7e-07 $l=5.20192e-07 $layer=licon1_PDIFF $count=2 $X=7.785
+ $Y=2.095 $X2=7.96 $Y2=2.535
r193 3 31 600 $w=1.7e-07 $l=9.17333e-07 $layer=licon1_PDIFF $count=1 $X=5.515
+ $Y=1.705 $X2=5.655 $Y2=2.555
r194 2 27 300 $w=1.7e-07 $l=4.79922e-07 $layer=licon1_PDIFF $count=2 $X=3.89
+ $Y=1.735 $X2=4.03 $Y2=2.15
r195 1 23 600 $w=1.7e-07 $l=9.17333e-07 $layer=licon1_PDIFF $count=1 $X=0.665
+ $Y=2.015 $X2=0.805 $Y2=2.865
.ends

.subckt PM_SKY130_FD_SC_LP__DFXBP_LP%A_239_403# 1 2 3 10 13 19 21 24 26 27
r53 26 27 8.69362 $w=2.58e-07 $l=1.65e-07 $layer=LI1_cond $X=2.945 $Y=2.115
+ $X2=2.78 $Y2=2.115
r54 21 23 10.7321 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=1.985 $Y=0.635
+ $X2=1.985 $Y2=0.865
r55 17 19 9.14916 $w=2.08e-07 $l=1.65e-07 $layer=LI1_cond $X=1.335 $Y=2.14
+ $X2=1.5 $Y2=2.14
r56 15 24 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.99 $Y=2.12
+ $X2=1.905 $Y2=2.12
r57 15 27 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=1.99 $Y=2.12
+ $X2=2.78 $Y2=2.12
r58 13 24 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.905 $Y=2.035
+ $X2=1.905 $Y2=2.12
r59 13 23 76.3316 $w=1.68e-07 $l=1.17e-06 $layer=LI1_cond $X=1.905 $Y=2.035
+ $X2=1.905 $Y2=0.865
r60 10 24 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.82 $Y=2.12
+ $X2=1.905 $Y2=2.12
r61 10 19 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=1.82 $Y=2.12 $X2=1.5
+ $Y2=2.12
r62 3 26 600 $w=1.7e-07 $l=5.25357e-07 $layer=licon1_PDIFF $count=1 $X=2.805
+ $Y=1.615 $X2=2.945 $Y2=2.075
r63 2 17 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.195
+ $Y=2.015 $X2=1.335 $Y2=2.16
r64 1 21 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.845
+ $Y=0.425 $X2=1.985 $Y2=0.635
.ends

.subckt PM_SKY130_FD_SC_LP__DFXBP_LP%A_349_323# 1 2 7 11 16
c33 16 0 1.6807e-19 $X=2.05 $Y=2.49
c34 11 0 1.29275e-19 $X=3.5 $Y=2.15
c35 7 0 9.0042e-20 $X=3.335 $Y=2.51
r36 14 16 9.14916 $w=2.08e-07 $l=1.65e-07 $layer=LI1_cond $X=1.885 $Y=2.49
+ $X2=2.05 $Y2=2.49
r37 9 11 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=3.5 $Y=2.425 $X2=3.5
+ $Y2=2.15
r38 7 9 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.335 $Y=2.51
+ $X2=3.5 $Y2=2.425
r39 7 16 83.8342 $w=1.68e-07 $l=1.285e-06 $layer=LI1_cond $X=3.335 $Y=2.51
+ $X2=2.05 $Y2=2.51
r40 2 11 300 $w=1.7e-07 $l=4.79922e-07 $layer=licon1_PDIFF $count=2 $X=3.36
+ $Y=1.735 $X2=3.5 $Y2=2.15
r41 1 14 600 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=1.745
+ $Y=1.615 $X2=1.885 $Y2=2.47
.ends

.subckt PM_SKY130_FD_SC_LP__DFXBP_LP%Q 1 2 8 11 12 13 14 15
r26 14 15 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=9.39 $Y=2.405
+ $X2=9.39 $Y2=2.69
r27 13 14 14.8421 $w=3.28e-07 $l=4.25e-07 $layer=LI1_cond $X=9.39 $Y=1.98
+ $X2=9.39 $Y2=2.405
r28 12 13 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=9.39 $Y=1.665
+ $X2=9.39 $Y2=1.98
r29 11 12 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=9.39 $Y=1.295
+ $X2=9.39 $Y2=1.665
r30 8 11 7.68295 $w=3.28e-07 $l=2.2e-07 $layer=LI1_cond $X=9.39 $Y=1.075
+ $X2=9.39 $Y2=1.295
r31 8 10 14.7516 $w=3.06e-07 $l=5.03438e-07 $layer=LI1_cond $X=9.39 $Y=1.075
+ $X2=9.76 $Y2=0.76
r32 2 15 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=9.245
+ $Y=1.835 $X2=9.39 $Y2=2.69
r33 2 13 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=9.245
+ $Y=1.835 $X2=9.39 $Y2=1.98
r34 1 10 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=9.62
+ $Y=0.635 $X2=9.76 $Y2=0.845
.ends

.subckt PM_SKY130_FD_SC_LP__DFXBP_LP%Q_N 1 2 7 8 9 10 11 12 13
r18 13 40 4.36531 $w=3.28e-07 $l=1.25e-07 $layer=LI1_cond $X=12.68 $Y=2.775
+ $X2=12.68 $Y2=2.9
r19 12 13 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=12.68 $Y=2.405
+ $X2=12.68 $Y2=2.775
r20 12 34 7.50834 $w=3.28e-07 $l=2.15e-07 $layer=LI1_cond $X=12.68 $Y=2.405
+ $X2=12.68 $Y2=2.19
r21 11 34 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=12.68 $Y=2.035
+ $X2=12.68 $Y2=2.19
r22 10 11 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=12.68 $Y=1.665
+ $X2=12.68 $Y2=2.035
r23 9 10 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=12.68 $Y=1.295
+ $X2=12.68 $Y2=1.665
r24 8 9 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=12.68 $Y=0.925
+ $X2=12.68 $Y2=1.295
r25 7 8 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=12.68 $Y=0.495
+ $X2=12.68 $Y2=0.925
r26 2 40 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=12.54
+ $Y=2.045 $X2=12.68 $Y2=2.9
r27 2 34 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=12.54
+ $Y=2.045 $X2=12.68 $Y2=2.19
r28 1 7 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=12.54
+ $Y=0.285 $X2=12.68 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__DFXBP_LP%VGND 1 2 3 4 5 6 21 25 29 33 37 41 44 45 47
+ 48 49 51 56 68 79 85 86 89 92 95 98
c130 41 0 9.72338e-20 $X=11.89 $Y=0.495
r131 98 99 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=11.76 $Y=0
+ $X2=11.76 $Y2=0
r132 95 96 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r133 92 93 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r134 89 90 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r135 86 99 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=12.72 $Y=0
+ $X2=11.76 $Y2=0
r136 85 86 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=12.72 $Y=0
+ $X2=12.72 $Y2=0
r137 83 98 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.055 $Y=0
+ $X2=11.89 $Y2=0
r138 83 85 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=12.055 $Y=0
+ $X2=12.72 $Y2=0
r139 82 99 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=10.8 $Y=0
+ $X2=11.76 $Y2=0
r140 81 82 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=10.8 $Y=0 $X2=10.8
+ $Y2=0
r141 79 98 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.725 $Y=0
+ $X2=11.89 $Y2=0
r142 79 81 60.3476 $w=1.68e-07 $l=9.25e-07 $layer=LI1_cond $X=11.725 $Y=0
+ $X2=10.8 $Y2=0
r143 78 82 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=10.32 $Y=0
+ $X2=10.8 $Y2=0
r144 77 78 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.32 $Y=0
+ $X2=10.32 $Y2=0
r145 75 78 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=8.88 $Y=0
+ $X2=10.32 $Y2=0
r146 75 96 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.88 $Y=0 $X2=8.4
+ $Y2=0
r147 74 77 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=8.88 $Y=0
+ $X2=10.32 $Y2=0
r148 74 75 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.88 $Y=0 $X2=8.88
+ $Y2=0
r149 72 95 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.585 $Y=0 $X2=8.46
+ $Y2=0
r150 72 74 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=8.585 $Y=0 $X2=8.88
+ $Y2=0
r151 70 71 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=6 $Y=0 $X2=6 $Y2=0
r152 68 95 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.335 $Y=0 $X2=8.46
+ $Y2=0
r153 68 70 152.337 $w=1.68e-07 $l=2.335e-06 $layer=LI1_cond $X=8.335 $Y=0 $X2=6
+ $Y2=0
r154 67 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=6
+ $Y2=0
r155 67 93 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=5.52 $Y=0 $X2=3.6
+ $Y2=0
r156 66 67 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.52 $Y=0
+ $X2=5.52 $Y2=0
r157 64 92 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.61 $Y=0 $X2=3.445
+ $Y2=0
r158 64 66 124.61 $w=1.68e-07 $l=1.91e-06 $layer=LI1_cond $X=3.61 $Y=0 $X2=5.52
+ $Y2=0
r159 63 93 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r160 62 63 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r161 60 63 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.68 $Y=0
+ $X2=3.12 $Y2=0
r162 60 90 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r163 59 62 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.68 $Y=0 $X2=3.12
+ $Y2=0
r164 59 60 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r165 57 89 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.36 $Y=0 $X2=1.235
+ $Y2=0
r166 57 59 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=1.36 $Y=0 $X2=1.68
+ $Y2=0
r167 56 92 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.28 $Y=0 $X2=3.445
+ $Y2=0
r168 56 62 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=3.28 $Y=0 $X2=3.12
+ $Y2=0
r169 54 90 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r170 53 54 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r171 51 89 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.11 $Y=0 $X2=1.235
+ $Y2=0
r172 51 53 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=1.11 $Y=0 $X2=0.72
+ $Y2=0
r173 49 96 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=6.48 $Y=0 $X2=8.4
+ $Y2=0
r174 49 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=0 $X2=6
+ $Y2=0
r175 47 77 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=10.465 $Y=0
+ $X2=10.32 $Y2=0
r176 47 48 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.465 $Y=0
+ $X2=10.59 $Y2=0
r177 46 81 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=10.715 $Y=0
+ $X2=10.8 $Y2=0
r178 46 48 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.715 $Y=0
+ $X2=10.59 $Y2=0
r179 44 66 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=5.66 $Y=0 $X2=5.52
+ $Y2=0
r180 44 45 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.66 $Y=0 $X2=5.785
+ $Y2=0
r181 43 70 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=5.91 $Y=0 $X2=6 $Y2=0
r182 43 45 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.91 $Y=0 $X2=5.785
+ $Y2=0
r183 39 98 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=11.89 $Y=0.085
+ $X2=11.89 $Y2=0
r184 39 41 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=11.89 $Y=0.085
+ $X2=11.89 $Y2=0.495
r185 35 48 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=10.59 $Y=0.085
+ $X2=10.59 $Y2=0
r186 35 37 35.0343 $w=2.48e-07 $l=7.6e-07 $layer=LI1_cond $X=10.59 $Y=0.085
+ $X2=10.59 $Y2=0.845
r187 31 95 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=8.46 $Y=0.085
+ $X2=8.46 $Y2=0
r188 31 33 18.9001 $w=2.48e-07 $l=4.1e-07 $layer=LI1_cond $X=8.46 $Y=0.085
+ $X2=8.46 $Y2=0.495
r189 27 45 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.785 $Y=0.085
+ $X2=5.785 $Y2=0
r190 27 29 34.5733 $w=2.48e-07 $l=7.5e-07 $layer=LI1_cond $X=5.785 $Y=0.085
+ $X2=5.785 $Y2=0.835
r191 23 92 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.445 $Y=0.085
+ $X2=3.445 $Y2=0
r192 23 25 18.6835 $w=3.28e-07 $l=5.35e-07 $layer=LI1_cond $X=3.445 $Y=0.085
+ $X2=3.445 $Y2=0.62
r193 19 89 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.235 $Y=0.085
+ $X2=1.235 $Y2=0
r194 19 21 25.3537 $w=2.48e-07 $l=5.5e-07 $layer=LI1_cond $X=1.235 $Y=0.085
+ $X2=1.235 $Y2=0.635
r195 6 41 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=11.75
+ $Y=0.285 $X2=11.89 $Y2=0.495
r196 5 37 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=10.41
+ $Y=0.635 $X2=10.55 $Y2=0.845
r197 4 33 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=8.28
+ $Y=0.285 $X2=8.42 $Y2=0.495
r198 3 29 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=5.605
+ $Y=0.625 $X2=5.745 $Y2=0.835
r199 2 25 182 $w=1.7e-07 $l=2.32164e-07 $layer=licon1_NDIFF $count=1 $X=3.225
+ $Y=0.595 $X2=3.445 $Y2=0.62
r200 1 21 182 $w=1.7e-07 $l=2.96985e-07 $layer=licon1_NDIFF $count=1 $X=0.985
+ $Y=0.425 $X2=1.195 $Y2=0.635
.ends

.subckt PM_SKY130_FD_SC_LP__DFXBP_LP%A_1232_153# 1 2 9 11 12 13
c32 13 0 1.69058e-19 $X=7.99 $Y=0.35
c33 11 0 1.1902e-19 $X=7.825 $Y=0.35
r34 13 16 5.06376 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=7.99 $Y=0.35
+ $X2=7.99 $Y2=0.495
r35 11 13 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.825 $Y=0.35
+ $X2=7.99 $Y2=0.35
r36 11 12 93.6203 $w=1.68e-07 $l=1.435e-06 $layer=LI1_cond $X=7.825 $Y=0.35
+ $X2=6.39 $Y2=0.35
r37 7 12 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=6.265 $Y=0.435
+ $X2=6.39 $Y2=0.35
r38 7 9 23.7403 $w=2.48e-07 $l=5.15e-07 $layer=LI1_cond $X=6.265 $Y=0.435
+ $X2=6.265 $Y2=0.95
r39 2 16 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=7.845
+ $Y=0.285 $X2=7.99 $Y2=0.495
r40 1 9 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=6.16
+ $Y=0.765 $X2=6.305 $Y2=0.95
.ends

