# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__einvn_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_lp__einvn_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.360000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.905000 1.195000 3.275000 1.525000 ;
    END
  END A
  PIN TE_B
    ANTENNAGATEAREA  0.537000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.550000 0.840000 0.945000 1.510000 ;
    END
  END TE_B
  PIN Z
    ANTENNADIFFAREA  0.903000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.110000 1.705000 3.265000 1.875000 ;
        RECT 2.110000 1.875000 2.370000 2.155000 ;
        RECT 2.495000 0.595000 2.835000 0.885000 ;
        RECT 2.495000 0.885000 2.735000 1.705000 ;
        RECT 2.975000 1.875000 3.265000 3.075000 ;
    END
  END Z
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.360000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.360000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.360000 0.085000 ;
      RECT 0.000000  3.245000 3.360000 3.415000 ;
      RECT 0.100000  0.355000 0.370000 1.680000 ;
      RECT 0.100000  1.680000 1.940000 1.850000 ;
      RECT 0.100000  1.850000 0.430000 2.485000 ;
      RECT 0.550000  0.085000 0.880000 0.560000 ;
      RECT 0.600000  2.020000 0.930000 3.245000 ;
      RECT 1.100000  2.020000 1.405000 2.325000 ;
      RECT 1.100000  2.325000 2.805000 2.495000 ;
      RECT 1.100000  2.495000 1.335000 3.075000 ;
      RECT 1.215000  0.255000 1.475000 1.005000 ;
      RECT 1.215000  1.005000 2.325000 1.175000 ;
      RECT 1.505000  2.665000 1.835000 3.245000 ;
      RECT 1.645000  0.085000 1.975000 0.835000 ;
      RECT 1.770000  1.345000 2.100000 1.535000 ;
      RECT 1.770000  1.535000 1.940000 1.680000 ;
      RECT 2.145000  0.255000 3.265000 0.425000 ;
      RECT 2.145000  0.425000 2.325000 1.005000 ;
      RECT 2.505000  2.495000 2.805000 3.075000 ;
      RECT 2.540000  2.045000 2.805000 2.325000 ;
      RECT 3.005000  0.425000 3.265000 1.025000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
  END
END sky130_fd_sc_lp__einvn_2
END LIBRARY
