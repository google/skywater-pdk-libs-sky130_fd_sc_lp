* File: sky130_fd_sc_lp__or2b_1.spice
* Created: Wed Sep  2 10:29:42 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__or2b_1.pex.spice"
.subckt sky130_fd_sc_lp__or2b_1  VNB VPB B_N A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* B_N	B_N
* VPB	VPB
* VNB	VNB
MM1000 N_VGND_M1000_d N_B_N_M1000_g N_A_27_535#_M1000_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75001.6
+ A=0.063 P=1.14 MULT=1
MM1003 N_A_224_382#_M1003_d N_A_27_535#_M1003_g N_VGND_M1000_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1007 N_VGND_M1007_d N_A_M1007_g N_A_224_382#_M1003_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0896 AS=0.0588 PD=0.81 PS=0.7 NRD=12.852 NRS=0 M=1 R=2.8 SA=75001.1
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1002 N_X_M1002_d N_A_224_382#_M1002_g N_VGND_M1007_d VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1792 PD=2.21 PS=1.62 NRD=0 NRS=3.564 M=1 R=5.6 SA=75000.9
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1006 N_VPWR_M1006_d N_B_N_M1006_g N_A_27_535#_M1006_s VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1113 AS=0.1113 PD=1.37 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1004 A_307_367# N_A_27_535#_M1004_g N_A_224_382#_M1004_s VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0441 AS=0.110175 PD=0.63 PS=1.37 NRD=23.443 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1005 N_VPWR_M1005_d N_A_M1005_g A_307_367# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.095025 AS=0.0441 PD=0.8175 PS=0.63 NRD=18.7544 NRS=23.443 M=1 R=2.8
+ SA=75000.5 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1001 N_X_M1001_d N_A_224_382#_M1001_g N_VPWR_M1005_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.285075 PD=3.05 PS=2.4525 NRD=0 NRS=2.8565 M=1 R=8.4 SA=75000.5
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX8_noxref VNB VPB NWDIODE A=6.0799 P=10.25
*
.include "sky130_fd_sc_lp__or2b_1.pxi.spice"
*
.ends
*
*
