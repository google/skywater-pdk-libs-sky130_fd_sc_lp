* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__busdrivernovlp2_20 A TE_B VGND VNB VPB VPWR Z
X0 VPWR A a_217_367# VPB sky130_fd_pr__pfet_01v8 w=1.26e+06u l=150000u
X1 VPWR a_217_367# Z VPB sky130_fd_pr__pfet_01v8 w=1.26e+06u l=150000u
X2 a_1238_47# a_726_47# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 a_217_367# a_1238_47# a_1451_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X4 a_726_47# A VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X5 a_27_367# TE_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 a_381_85# a_217_367# VPWR VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X7 VPWR a_217_367# Z VPB sky130_fd_pr__pfet_01v8 w=1.26e+06u l=150000u
X8 Z a_726_47# VGND VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X9 a_658_367# a_381_85# a_726_47# VPB sky130_fd_pr__pfet_01v8 w=1.26e+06u l=150000u
X10 VGND a_27_367# a_303_85# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X11 VGND A a_726_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X12 Z a_726_47# VGND VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X13 Z a_217_367# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.26e+06u l=150000u
X14 VPWR TE_B a_1260_373# VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X15 a_217_367# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.26e+06u l=150000u
X16 Z a_217_367# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.26e+06u l=150000u
X17 VGND a_726_47# Z VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X18 Z a_217_367# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.26e+06u l=150000u
X19 Z a_217_367# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.26e+06u l=150000u
X20 Z a_217_367# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.26e+06u l=150000u
X21 VGND TE_B a_1238_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X22 a_1451_47# A VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X23 Z a_217_367# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.26e+06u l=150000u
X24 VGND a_726_47# Z VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X25 VPWR a_217_367# Z VPB sky130_fd_pr__pfet_01v8 w=1.26e+06u l=150000u
X26 a_27_367# TE_B VPWR VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X27 VPWR a_217_367# Z VPB sky130_fd_pr__pfet_01v8 w=1.26e+06u l=150000u
X28 Z a_726_47# VGND VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X29 VGND a_726_47# Z VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X30 VPWR a_217_367# Z VPB sky130_fd_pr__pfet_01v8 w=1.26e+06u l=150000u
X31 Z a_726_47# VGND VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X32 VPWR A a_658_367# VPB sky130_fd_pr__pfet_01v8 w=1.26e+06u l=150000u
X33 VPWR a_217_367# Z VPB sky130_fd_pr__pfet_01v8 w=1.26e+06u l=150000u
X34 VPWR a_217_367# Z VPB sky130_fd_pr__pfet_01v8 w=1.26e+06u l=150000u
X35 VGND a_726_47# Z VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X36 VPWR a_27_367# a_217_367# VPB sky130_fd_pr__pfet_01v8 w=1.26e+06u l=150000u
X37 VGND TE_B a_726_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X38 VPWR a_217_367# Z VPB sky130_fd_pr__pfet_01v8 w=1.26e+06u l=150000u
X39 a_726_47# TE_B VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X40 VPWR a_217_367# Z VPB sky130_fd_pr__pfet_01v8 w=1.26e+06u l=150000u
X41 VPWR a_217_367# Z VPB sky130_fd_pr__pfet_01v8 w=1.26e+06u l=150000u
X42 VGND a_726_47# Z VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X43 a_658_367# A VPWR VPB sky130_fd_pr__pfet_01v8 w=1.26e+06u l=150000u
X44 Z a_217_367# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.26e+06u l=150000u
X45 Z a_217_367# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.26e+06u l=150000u
X46 VGND a_726_47# Z VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X47 Z a_217_367# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.26e+06u l=150000u
X48 Z a_726_47# VGND VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X49 VPWR a_27_367# a_381_85# VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X50 a_303_85# a_217_367# a_381_85# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X51 VGND A a_1451_47# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X52 Z a_726_47# VGND VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X53 a_726_47# a_381_85# a_658_367# VPB sky130_fd_pr__pfet_01v8 w=1.26e+06u l=150000u
X54 VGND a_726_47# Z VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X55 a_217_367# a_27_367# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.26e+06u l=150000u
X56 a_1260_373# a_726_47# a_1238_47# VPB sky130_fd_pr__pfet_01v8 w=840000u l=150000u
X57 Z a_217_367# VPWR VPB sky130_fd_pr__pfet_01v8 w=1.26e+06u l=150000u
X58 a_1451_47# a_1238_47# a_217_367# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X59 Z a_726_47# VGND VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
.ends
