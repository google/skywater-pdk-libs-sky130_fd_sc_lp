# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__xor2_0
  CLASS CORE ;
  FOREIGN sky130_fd_sc_lp__xor2_0 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.360000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.625000 1.210000 1.350000 1.395000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.205000 1.185000 0.455000 1.565000 ;
        RECT 0.205000 1.565000 1.940000 1.855000 ;
        RECT 1.520000 1.210000 1.940000 1.565000 ;
    END
  END B
  PIN X
    ANTENNADIFFAREA  0.516100 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.970000 0.410000 2.815000 0.700000 ;
        RECT 2.545000 1.815000 2.815000 2.495000 ;
        RECT 2.645000 0.700000 2.815000 1.815000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 3.360000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 3.360000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.360000 0.085000 ;
      RECT 0.000000  3.245000 3.360000 3.415000 ;
      RECT 0.095000  2.025000 2.375000 2.195000 ;
      RECT 0.095000  2.195000 0.425000 3.065000 ;
      RECT 0.270000  0.085000 0.560000 0.800000 ;
      RECT 0.730000  0.395000 0.960000 0.870000 ;
      RECT 0.730000  0.870000 2.475000 1.040000 ;
      RECT 0.915000  2.385000 1.210000 3.245000 ;
      RECT 1.130000  0.085000 1.460000 0.700000 ;
      RECT 1.380000  2.365000 2.375000 2.535000 ;
      RECT 1.380000  2.535000 1.640000 3.065000 ;
      RECT 1.810000  2.705000 2.035000 3.245000 ;
      RECT 2.205000  1.040000 2.475000 1.625000 ;
      RECT 2.205000  1.625000 2.375000 2.025000 ;
      RECT 2.205000  2.535000 2.375000 2.665000 ;
      RECT 2.205000  2.665000 3.255000 2.835000 ;
      RECT 2.985000  0.085000 3.255000 0.800000 ;
      RECT 2.985000  1.815000 3.255000 2.665000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
  END
END sky130_fd_sc_lp__xor2_0
END LIBRARY
