* File: sky130_fd_sc_lp__a32o_2.pex.spice
* Created: Wed Sep  2 09:27:41 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A32O_2%A_108_267# 1 2 9 13 17 21 24 25 26 27 29 35
+ 43
c78 29 0 2.42403e-19 $X=2.28 $Y=1.98
c79 24 0 6.64853e-20 $X=1.33 $Y=1.405
r80 42 43 30 $w=2.41e-07 $l=1.5e-07 $layer=POLY_cond $X=1.045 $Y=1.5 $X2=1.195
+ $Y2=1.5
r81 33 43 11 $w=2.41e-07 $l=5.5e-08 $layer=POLY_cond $X=1.25 $Y=1.5 $X2=1.195
+ $Y2=1.5
r82 32 35 4.43636 $w=1.98e-07 $l=8e-08 $layer=LI1_cond $X=1.25 $Y=1.505 $X2=1.33
+ $Y2=1.505
r83 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.25
+ $Y=1.5 $X2=1.25 $Y2=1.5
r84 27 29 46.9904 $w=1.88e-07 $l=8.05e-07 $layer=LI1_cond $X=2.28 $Y=1.175
+ $X2=2.28 $Y2=1.98
r85 25 27 7.67083 $w=5.73e-07 $l=1.30767e-07 $layer=LI1_cond $X=2.185 $Y=1.09
+ $X2=2.28 $Y2=1.175
r86 25 38 14.2653 $w=5.73e-07 $l=8.22618e-07 $layer=LI1_cond $X=2.185 $Y=1.09
+ $X2=2.525 $Y2=0.42
r87 25 26 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=2.185 $Y=1.09
+ $X2=1.415 $Y2=1.09
r88 24 35 1.68994 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=1.33 $Y=1.405 $X2=1.33
+ $Y2=1.505
r89 23 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.33 $Y=1.175
+ $X2=1.415 $Y2=1.09
r90 23 24 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=1.33 $Y=1.175
+ $X2=1.33 $Y2=1.405
r91 19 43 13.8727 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.195 $Y=1.335
+ $X2=1.195 $Y2=1.5
r92 19 21 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=1.195 $Y=1.335
+ $X2=1.195 $Y2=0.655
r93 15 42 13.8727 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.045 $Y=1.665
+ $X2=1.045 $Y2=1.5
r94 15 17 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=1.045 $Y=1.665
+ $X2=1.045 $Y2=2.465
r95 11 42 56 $w=2.41e-07 $l=3.52987e-07 $layer=POLY_cond $X=0.765 $Y=1.335
+ $X2=1.045 $Y2=1.5
r96 11 13 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=0.765 $Y=1.335
+ $X2=0.765 $Y2=0.655
r97 7 11 30 $w=2.41e-07 $l=2.12132e-07 $layer=POLY_cond $X=0.615 $Y=1.485
+ $X2=0.765 $Y2=1.335
r98 7 9 502.511 $w=1.5e-07 $l=9.8e-07 $layer=POLY_cond $X=0.615 $Y=1.485
+ $X2=0.615 $Y2=2.465
r99 2 29 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=2.14
+ $Y=1.835 $X2=2.28 $Y2=1.98
r100 1 38 91 $w=1.7e-07 $l=2.93258e-07 $layer=licon1_NDIFF $count=2 $X=2.52
+ $Y=0.235 $X2=2.735 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__A32O_2%B2 1 3 6 8 12 13
c38 13 0 6.64853e-20 $X=2.065 $Y=1.535
r39 13 14 2.60541 $w=3.7e-07 $l=2e-08 $layer=POLY_cond $X=2.065 $Y=1.535
+ $X2=2.085 $Y2=1.535
r40 11 13 31.9162 $w=3.7e-07 $l=2.45e-07 $layer=POLY_cond $X=1.82 $Y=1.535
+ $X2=2.065 $Y2=1.535
r41 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.82
+ $Y=1.51 $X2=1.82 $Y2=1.51
r42 8 12 4.15415 $w=4.28e-07 $l=1.55e-07 $layer=LI1_cond $X=1.8 $Y=1.665 $X2=1.8
+ $Y2=1.51
r43 4 14 23.9667 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=2.085 $Y=1.345
+ $X2=2.085 $Y2=1.535
r44 4 6 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.085 $Y=1.345
+ $X2=2.085 $Y2=0.655
r45 1 13 23.9667 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=2.065 $Y=1.725
+ $X2=2.065 $Y2=1.535
r46 1 3 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=2.065 $Y=1.725
+ $X2=2.065 $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__A32O_2%B1 1 3 6 8 9 10 11 17
r39 17 19 21.1266 $w=3.08e-07 $l=1.35e-07 $layer=POLY_cond $X=2.495 $Y=1.35
+ $X2=2.63 $Y2=1.35
r40 16 17 7.82468 $w=3.08e-07 $l=5e-08 $layer=POLY_cond $X=2.445 $Y=1.35
+ $X2=2.495 $Y2=1.35
r41 10 11 21.5981 $w=1.88e-07 $l=3.7e-07 $layer=LI1_cond $X=2.64 $Y=2.035
+ $X2=2.64 $Y2=2.405
r42 9 10 21.5981 $w=1.88e-07 $l=3.7e-07 $layer=LI1_cond $X=2.64 $Y=1.665
+ $X2=2.64 $Y2=2.035
r43 8 9 21.5981 $w=1.88e-07 $l=3.7e-07 $layer=LI1_cond $X=2.64 $Y=1.295 $X2=2.64
+ $Y2=1.665
r44 8 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.63
+ $Y=1.35 $X2=2.63 $Y2=1.35
r45 4 17 19.5884 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.495 $Y=1.515
+ $X2=2.495 $Y2=1.35
r46 4 6 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=2.495 $Y=1.515
+ $X2=2.495 $Y2=2.465
r47 1 16 19.5884 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.445 $Y=1.185
+ $X2=2.445 $Y2=1.35
r48 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.445 $Y=1.185
+ $X2=2.445 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__A32O_2%A1 3 6 8 9 10 15 17
c39 17 0 5.12769e-20 $X=3.17 $Y=1.185
c40 8 0 1.91126e-19 $X=3.12 $Y=0.555
r41 15 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.17 $Y=1.35
+ $X2=3.17 $Y2=1.515
r42 15 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.17 $Y=1.35
+ $X2=3.17 $Y2=1.185
r43 10 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.17
+ $Y=1.35 $X2=3.17 $Y2=1.35
r44 9 10 19.382 $w=2.18e-07 $l=3.7e-07 $layer=LI1_cond $X=3.145 $Y=0.925
+ $X2=3.145 $Y2=1.295
r45 8 9 19.382 $w=2.18e-07 $l=3.7e-07 $layer=LI1_cond $X=3.145 $Y=0.555
+ $X2=3.145 $Y2=0.925
r46 6 18 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=3.205 $Y=2.465
+ $X2=3.205 $Y2=1.515
r47 3 17 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=3.08 $Y=0.655
+ $X2=3.08 $Y2=1.185
.ends

.subckt PM_SKY130_FD_SC_LP__A32O_2%A2 3 6 8 9 10 21 23
c34 21 0 1.64508e-19 $X=3.71 $Y=1.35
c35 6 0 9.4196e-20 $X=3.73 $Y=2.465
r36 21 24 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.71 $Y=1.35
+ $X2=3.71 $Y2=1.515
r37 21 23 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.71 $Y=1.35
+ $X2=3.71 $Y2=1.185
r38 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.71
+ $Y=1.35 $X2=3.71 $Y2=1.35
r39 10 22 0.888977 $w=7.38e-07 $l=5.5e-08 $layer=LI1_cond $X=3.795 $Y=1.295
+ $X2=3.795 $Y2=1.35
r40 9 10 5.98039 $w=7.38e-07 $l=3.7e-07 $layer=LI1_cond $X=3.795 $Y=0.925
+ $X2=3.795 $Y2=1.295
r41 8 9 5.98039 $w=7.38e-07 $l=3.7e-07 $layer=LI1_cond $X=3.795 $Y=0.555
+ $X2=3.795 $Y2=0.925
r42 6 24 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=3.73 $Y=2.465
+ $X2=3.73 $Y2=1.515
r43 3 23 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=3.62 $Y=0.655
+ $X2=3.62 $Y2=1.185
.ends

.subckt PM_SKY130_FD_SC_LP__A32O_2%A3 3 7 9 10 16
c23 9 0 2.58704e-19 $X=4.56 $Y=1.295
r24 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.43
+ $Y=1.375 $X2=4.43 $Y2=1.375
r25 13 16 47.2125 $w=3.3e-07 $l=2.7e-07 $layer=POLY_cond $X=4.16 $Y=1.375
+ $X2=4.43 $Y2=1.375
r26 10 17 9.03266 $w=3.68e-07 $l=2.9e-07 $layer=LI1_cond $X=4.53 $Y=1.665
+ $X2=4.53 $Y2=1.375
r27 9 17 2.49177 $w=3.68e-07 $l=8e-08 $layer=LI1_cond $X=4.53 $Y=1.295 $X2=4.53
+ $Y2=1.375
r28 5 13 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.16 $Y=1.54
+ $X2=4.16 $Y2=1.375
r29 5 7 474.309 $w=1.5e-07 $l=9.25e-07 $layer=POLY_cond $X=4.16 $Y=1.54 $X2=4.16
+ $Y2=2.465
r30 1 13 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.16 $Y=1.21
+ $X2=4.16 $Y2=1.375
r31 1 3 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=4.16 $Y=1.21 $X2=4.16
+ $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__A32O_2%X 1 2 3 12 16 20 24 30 32 33
r42 31 33 1.82734 $w=7.18e-07 $l=1.1e-07 $layer=LI1_cond $X=0.515 $Y=1.775
+ $X2=0.515 $Y2=1.665
r43 31 32 1.85714 $w=5.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.515 $Y=1.775
+ $X2=0.515 $Y2=1.86
r44 30 33 7.14325 $w=7.18e-07 $l=4.3e-07 $layer=LI1_cond $X=0.515 $Y=1.235
+ $X2=0.515 $Y2=1.665
r45 29 30 10.2049 $w=7.18e-07 $l=1.7e-07 $layer=LI1_cond $X=0.615 $Y=1.065
+ $X2=0.615 $Y2=1.235
r46 24 26 42.8709 $w=2.48e-07 $l=9.3e-07 $layer=LI1_cond $X=1.29 $Y=1.98
+ $X2=1.29 $Y2=2.91
r47 22 24 1.61342 $w=2.48e-07 $l=3.5e-08 $layer=LI1_cond $X=1.29 $Y=1.945
+ $X2=1.29 $Y2=1.98
r48 20 29 37.6507 $w=1.88e-07 $l=6.45e-07 $layer=LI1_cond $X=0.98 $Y=0.42
+ $X2=0.98 $Y2=1.065
r49 17 32 5.62386 $w=1.7e-07 $l=3.6e-07 $layer=LI1_cond $X=0.875 $Y=1.86
+ $X2=0.515 $Y2=1.86
r50 16 22 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.165 $Y=1.86
+ $X2=1.29 $Y2=1.945
r51 16 17 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=1.165 $Y=1.86
+ $X2=0.875 $Y2=1.86
r52 12 14 31.5227 $w=3.38e-07 $l=9.3e-07 $layer=LI1_cond $X=0.325 $Y=1.98
+ $X2=0.325 $Y2=2.91
r53 10 32 1.85714 $w=5.3e-07 $l=2.28583e-07 $layer=LI1_cond $X=0.325 $Y=1.945
+ $X2=0.515 $Y2=1.86
r54 10 12 1.18634 $w=3.38e-07 $l=3.5e-08 $layer=LI1_cond $X=0.325 $Y=1.945
+ $X2=0.325 $Y2=1.98
r55 3 26 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=1.12
+ $Y=1.835 $X2=1.26 $Y2=2.91
r56 3 24 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.12
+ $Y=1.835 $X2=1.26 $Y2=1.98
r57 2 14 400 $w=1.7e-07 $l=1.13578e-06 $layer=licon1_PDIFF $count=1 $X=0.275
+ $Y=1.835 $X2=0.4 $Y2=2.91
r58 2 12 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.275
+ $Y=1.835 $X2=0.4 $Y2=1.98
r59 1 20 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=0.84
+ $Y=0.235 $X2=0.98 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__A32O_2%VPWR 1 2 3 14 20 24 26 31 32 33 42 47 51
r55 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r56 47 48 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r57 45 51 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r58 44 45 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r59 42 50 4.4922 $w=1.7e-07 $l=2.95e-07 $layer=LI1_cond $X=4.21 $Y=3.33
+ $X2=4.505 $Y2=3.33
r60 42 44 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=4.21 $Y=3.33
+ $X2=4.08 $Y2=3.33
r61 41 45 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=4.08 $Y2=3.33
r62 40 41 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r63 38 48 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r64 37 40 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=3.12 $Y2=3.33
r65 37 38 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r66 35 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.995 $Y=3.33
+ $X2=0.83 $Y2=3.33
r67 35 37 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=0.995 $Y=3.33
+ $X2=1.2 $Y2=3.33
r68 33 41 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.4 $Y=3.33
+ $X2=3.12 $Y2=3.33
r69 33 38 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=2.4 $Y=3.33 $X2=1.2
+ $Y2=3.33
r70 31 40 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=3.3 $Y=3.33 $X2=3.12
+ $Y2=3.33
r71 31 32 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.3 $Y=3.33
+ $X2=3.465 $Y2=3.33
r72 30 44 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=3.63 $Y=3.33
+ $X2=4.08 $Y2=3.33
r73 30 32 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.63 $Y=3.33
+ $X2=3.465 $Y2=3.33
r74 26 29 33.0018 $w=3.28e-07 $l=9.45e-07 $layer=LI1_cond $X=4.375 $Y=2.005
+ $X2=4.375 $Y2=2.95
r75 24 50 3.27398 $w=3.3e-07 $l=1.67183e-07 $layer=LI1_cond $X=4.375 $Y=3.245
+ $X2=4.505 $Y2=3.33
r76 24 29 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=4.375 $Y=3.245
+ $X2=4.375 $Y2=2.95
r77 20 23 26.5411 $w=3.28e-07 $l=7.6e-07 $layer=LI1_cond $X=3.465 $Y=2.19
+ $X2=3.465 $Y2=2.95
r78 18 32 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.465 $Y=3.245
+ $X2=3.465 $Y2=3.33
r79 18 23 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=3.465 $Y=3.245
+ $X2=3.465 $Y2=2.95
r80 14 17 26.8903 $w=3.28e-07 $l=7.7e-07 $layer=LI1_cond $X=0.83 $Y=2.2 $X2=0.83
+ $Y2=2.97
r81 12 47 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.83 $Y=3.245
+ $X2=0.83 $Y2=3.33
r82 12 17 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=0.83 $Y=3.245
+ $X2=0.83 $Y2=2.97
r83 3 29 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=4.235
+ $Y=1.835 $X2=4.375 $Y2=2.95
r84 3 26 400 $w=1.7e-07 $l=2.29565e-07 $layer=licon1_PDIFF $count=1 $X=4.235
+ $Y=1.835 $X2=4.375 $Y2=2.005
r85 2 23 400 $w=1.7e-07 $l=1.20395e-06 $layer=licon1_PDIFF $count=1 $X=3.28
+ $Y=1.835 $X2=3.465 $Y2=2.95
r86 2 20 400 $w=1.7e-07 $l=4.37836e-07 $layer=licon1_PDIFF $count=1 $X=3.28
+ $Y=1.835 $X2=3.465 $Y2=2.19
r87 1 17 400 $w=1.7e-07 $l=1.20297e-06 $layer=licon1_PDIFF $count=1 $X=0.69
+ $Y=1.835 $X2=0.83 $Y2=2.97
r88 1 14 400 $w=1.7e-07 $l=4.29331e-07 $layer=licon1_PDIFF $count=1 $X=0.69
+ $Y=1.835 $X2=0.83 $Y2=2.2
.ends

.subckt PM_SKY130_FD_SC_LP__A32O_2%A_345_367# 1 2 3 10 12 19 20 21 24 32 33
r49 31 33 10.7212 $w=3.28e-07 $l=3.07e-07 $layer=LI1_cond $X=2.71 $Y=2.91
+ $X2=3.017 $Y2=2.91
r50 31 32 7.76373 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=2.71 $Y=2.91
+ $X2=2.565 $Y2=2.91
r51 24 26 44.6572 $w=2.38e-07 $l=9.3e-07 $layer=LI1_cond $X=3.92 $Y=1.98
+ $X2=3.92 $Y2=2.91
r52 22 24 2.64102 $w=2.38e-07 $l=5.5e-08 $layer=LI1_cond $X=3.92 $Y=1.925
+ $X2=3.92 $Y2=1.98
r53 20 22 7.07814 $w=1.7e-07 $l=1.56844e-07 $layer=LI1_cond $X=3.8 $Y=1.84
+ $X2=3.92 $Y2=1.925
r54 20 21 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.8 $Y=1.84 $X2=3.13
+ $Y2=1.84
r55 17 33 2.99809 $w=2.25e-07 $l=1.65e-07 $layer=LI1_cond $X=3.017 $Y=2.745
+ $X2=3.017 $Y2=2.91
r56 17 19 39.1831 $w=2.23e-07 $l=7.65e-07 $layer=LI1_cond $X=3.017 $Y=2.745
+ $X2=3.017 $Y2=1.98
r57 16 21 6.9898 $w=1.7e-07 $l=1.49579e-07 $layer=LI1_cond $X=3.017 $Y=1.925
+ $X2=3.13 $Y2=1.84
r58 16 19 2.81708 $w=2.23e-07 $l=5.5e-08 $layer=LI1_cond $X=3.017 $Y=1.925
+ $X2=3.017 $Y2=1.98
r59 15 29 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.015 $Y=2.99
+ $X2=1.85 $Y2=2.99
r60 15 32 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=2.015 $Y=2.99
+ $X2=2.565 $Y2=2.99
r61 10 29 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.85 $Y=2.905 $X2=1.85
+ $Y2=2.99
r62 10 12 31.081 $w=3.28e-07 $l=8.9e-07 $layer=LI1_cond $X=1.85 $Y=2.905
+ $X2=1.85 $Y2=2.015
r63 3 26 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=3.805
+ $Y=1.835 $X2=3.945 $Y2=2.91
r64 3 24 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=3.805
+ $Y=1.835 $X2=3.945 $Y2=1.98
r65 2 31 600 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=2.57
+ $Y=1.835 $X2=2.71 $Y2=2.91
r66 2 19 300 $w=1.7e-07 $l=4.87134e-07 $layer=licon1_PDIFF $count=2 $X=2.57
+ $Y=1.835 $X2=2.99 $Y2=1.98
r67 1 29 400 $w=1.7e-07 $l=1.17083e-06 $layer=licon1_PDIFF $count=1 $X=1.725
+ $Y=1.835 $X2=1.85 $Y2=2.945
r68 1 12 400 $w=1.7e-07 $l=2.34307e-07 $layer=licon1_PDIFF $count=1 $X=1.725
+ $Y=1.835 $X2=1.85 $Y2=2.015
.ends

.subckt PM_SKY130_FD_SC_LP__A32O_2%VGND 1 2 3 12 14 16 19 20 21 27 31 41 48
r54 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r55 41 44 5.75329 $w=7.88e-07 $l=3.8e-07 $layer=LI1_cond $X=1.64 $Y=0 $X2=1.64
+ $Y2=0.38
r56 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r57 38 48 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=4.56
+ $Y2=0
r58 37 38 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r59 35 42 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.68
+ $Y2=0
r60 34 37 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=2.16 $Y=0 $X2=4.08
+ $Y2=0
r61 34 35 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r62 32 41 10.1246 $w=1.7e-07 $l=3.95e-07 $layer=LI1_cond $X=2.035 $Y=0 $X2=1.64
+ $Y2=0
r63 32 34 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=2.035 $Y=0 $X2=2.16
+ $Y2=0
r64 31 47 3.94577 $w=1.7e-07 $l=2.32e-07 $layer=LI1_cond $X=4.335 $Y=0 $X2=4.567
+ $Y2=0
r65 31 37 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=4.335 $Y=0 $X2=4.08
+ $Y2=0
r66 30 42 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r67 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r68 27 41 10.1246 $w=1.7e-07 $l=3.95e-07 $layer=LI1_cond $X=1.245 $Y=0 $X2=1.64
+ $Y2=0
r69 27 29 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=1.245 $Y=0 $X2=1.2
+ $Y2=0
r70 25 30 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=1.2
+ $Y2=0
r71 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r72 21 38 0.468274 $w=4.9e-07 $l=1.68e-06 $layer=MET1_cond $X=2.4 $Y=0 $X2=4.08
+ $Y2=0
r73 21 35 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.4 $Y=0 $X2=2.16
+ $Y2=0
r74 19 24 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=0.385 $Y=0 $X2=0.24
+ $Y2=0
r75 19 20 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.385 $Y=0 $X2=0.55
+ $Y2=0
r76 18 29 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=0.715 $Y=0 $X2=1.2
+ $Y2=0
r77 18 20 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.715 $Y=0 $X2=0.55
+ $Y2=0
r78 14 47 3.23145 $w=2.55e-07 $l=1.41244e-07 $layer=LI1_cond $X=4.462 $Y=0.085
+ $X2=4.567 $Y2=0
r79 14 16 13.3322 $w=2.53e-07 $l=2.95e-07 $layer=LI1_cond $X=4.462 $Y=0.085
+ $X2=4.462 $Y2=0.38
r80 10 20 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.55 $Y=0.085
+ $X2=0.55 $Y2=0
r81 10 12 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.55 $Y=0.085
+ $X2=0.55 $Y2=0.38
r82 3 16 91 $w=1.7e-07 $l=2.5229e-07 $layer=licon1_NDIFF $count=2 $X=4.235
+ $Y=0.235 $X2=4.425 $Y2=0.38
r83 2 44 45.5 $w=1.7e-07 $l=6.68581e-07 $layer=licon1_NDIFF $count=4 $X=1.27
+ $Y=0.235 $X2=1.87 $Y2=0.38
r84 1 12 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.425
+ $Y=0.235 $X2=0.55 $Y2=0.38
.ends

