* File: sky130_fd_sc_lp__iso0n_lp2.spice
* Created: Wed Sep  2 09:57:34 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__iso0n_lp2.pex.spice"
.subckt sky130_fd_sc_lp__iso0n_lp2  VNB VPB A SLEEP_B VPWR X KAGND VGND
* 
* KAGND	KAGND
* X	X
* VPWR	VPWR
* SLEEP_B	SLEEP_B
* A	A
* VPB	VPB
* VNB	VNB
MM1001 A_152_65# N_A_M1001_g N_A_65_65#_M1001_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.1197 PD=0.66 PS=1.41 NRD=18.564 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1002 N_KAGND_M1002_d N_SLEEP_B_M1002_g A_152_65# VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0504 PD=0.7 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75000.6
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1004 A_316_65# N_A_65_65#_M1004_g N_KAGND_M1002_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.0588 PD=0.66 PS=0.7 NRD=18.564 NRS=0 M=1 R=2.8 SA=75001
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1003 N_X_M1003_d N_A_65_65#_M1003_g A_316_65# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0504 PD=1.41 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75001.4
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1005 N_A_65_65#_M1005_d N_A_M1005_g N_VPWR_M1005_s VPB PHIGHVT L=0.25 W=1
+ AD=0.14 AS=0.35 PD=1.28 PS=2.7 NRD=0 NRS=12.7853 M=1 R=4 SA=125000 SB=125001
+ A=0.25 P=2.5 MULT=1
MM1000 N_VPWR_M1000_d N_SLEEP_B_M1000_g N_A_65_65#_M1005_d VPB PHIGHVT L=0.25
+ W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125001 SB=125001
+ A=0.25 P=2.5 MULT=1
MM1006 N_X_M1006_d N_A_65_65#_M1006_g N_VPWR_M1000_d VPB PHIGHVT L=0.25 W=1
+ AD=0.285 AS=0.14 PD=2.57 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125001 SB=125000
+ A=0.25 P=2.5 MULT=1
DX7_noxref VNB VPB NWDIODE A=5.1847 P=9.29
*
.include "sky130_fd_sc_lp__iso0n_lp2.pxi.spice"
*
.ends
*
*
