* File: sky130_fd_sc_lp__maj3_1.pex.spice
* Created: Wed Sep  2 09:59:24 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__MAJ3_1%A 3 7 11 15 17 18 26
c40 3 0 4.15925e-20 $X=0.87 $Y=2.165
r41 24 26 17.4217 $w=2.49e-07 $l=9e-08 $layer=POLY_cond $X=1.21 $Y=1.29 $X2=1.3
+ $Y2=1.29
r42 22 24 36.7791 $w=2.49e-07 $l=1.9e-07 $layer=POLY_cond $X=1.02 $Y=1.29
+ $X2=1.21 $Y2=1.29
r43 18 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.21
+ $Y=1.29 $X2=1.21 $Y2=1.29
r44 17 18 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=0.72 $Y=1.29 $X2=1.2
+ $Y2=1.29
r45 13 26 38.7149 $w=2.49e-07 $l=2.70185e-07 $layer=POLY_cond $X=1.5 $Y=1.125
+ $X2=1.3 $Y2=1.29
r46 13 15 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=1.5 $Y=1.125 $X2=1.5
+ $Y2=0.495
r47 9 26 14.627 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.3 $Y=1.455 $X2=1.3
+ $Y2=1.29
r48 9 11 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=1.3 $Y=1.455 $X2=1.3
+ $Y2=2.165
r49 5 22 14.627 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.02 $Y=1.125
+ $X2=1.02 $Y2=1.29
r50 5 7 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=1.02 $Y=1.125 $X2=1.02
+ $Y2=0.495
r51 1 22 29.0361 $w=2.49e-07 $l=2.2798e-07 $layer=POLY_cond $X=0.87 $Y=1.455
+ $X2=1.02 $Y2=1.29
r52 1 3 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=0.87 $Y=1.455 $X2=0.87
+ $Y2=2.165
.ends

.subckt PM_SKY130_FD_SC_LP__MAJ3_1%B 1 3 6 9 12 16 20 22 23 31
r47 29 31 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.98 $Y=1.345
+ $X2=2.32 $Y2=1.345
r48 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.98
+ $Y=1.345 $X2=1.98 $Y2=1.345
r49 26 29 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=1.89 $Y=1.345 $X2=1.98
+ $Y2=1.345
r50 23 30 6.28605 $w=3.28e-07 $l=1.8e-07 $layer=LI1_cond $X=2.16 $Y=1.345
+ $X2=1.98 $Y2=1.345
r51 22 30 10.4768 $w=3.28e-07 $l=3e-07 $layer=LI1_cond $X=1.68 $Y=1.345 $X2=1.98
+ $Y2=1.345
r52 18 20 117.936 $w=1.5e-07 $l=2.3e-07 $layer=POLY_cond $X=1.66 $Y=1.77
+ $X2=1.89 $Y2=1.77
r53 14 31 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.32 $Y=1.51
+ $X2=2.32 $Y2=1.345
r54 14 16 330.734 $w=1.5e-07 $l=6.45e-07 $layer=POLY_cond $X=2.32 $Y=1.51
+ $X2=2.32 $Y2=2.155
r55 10 31 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.32 $Y=1.18
+ $X2=2.32 $Y2=1.345
r56 10 12 351.245 $w=1.5e-07 $l=6.85e-07 $layer=POLY_cond $X=2.32 $Y=1.18
+ $X2=2.32 $Y2=0.495
r57 9 20 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.89 $Y=1.695
+ $X2=1.89 $Y2=1.77
r58 8 26 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.89 $Y=1.51
+ $X2=1.89 $Y2=1.345
r59 8 9 94.8617 $w=1.5e-07 $l=1.85e-07 $layer=POLY_cond $X=1.89 $Y=1.51 $X2=1.89
+ $Y2=1.695
r60 4 26 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.89 $Y=1.18
+ $X2=1.89 $Y2=1.345
r61 4 6 351.245 $w=1.5e-07 $l=6.85e-07 $layer=POLY_cond $X=1.89 $Y=1.18 $X2=1.89
+ $Y2=0.495
r62 1 18 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.66 $Y=1.845
+ $X2=1.66 $Y2=1.77
r63 1 3 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.66 $Y=1.845 $X2=1.66
+ $Y2=2.165
.ends

.subckt PM_SKY130_FD_SC_LP__MAJ3_1%C 3 6 7 8 11 14 15 16 17 22
c53 17 0 1.87895e-19 $X=2.64 $Y=2.775
c54 11 0 6.76105e-20 $X=2.68 $Y=0.495
r55 22 25 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=2.59 $Y=2.9 $X2=2.59
+ $Y2=2.99
r56 22 24 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.59 $Y=2.9
+ $X2=2.59 $Y2=2.735
r57 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.59
+ $Y=2.9 $X2=2.59 $Y2=2.9
r58 17 23 1.42277 $w=4.03e-07 $l=5e-08 $layer=LI1_cond $X=2.64 $Y=2.862 $X2=2.59
+ $Y2=2.862
r59 16 23 12.2358 $w=4.03e-07 $l=4.3e-07 $layer=LI1_cond $X=2.16 $Y=2.862
+ $X2=2.59 $Y2=2.862
r60 15 16 13.6586 $w=4.03e-07 $l=4.8e-07 $layer=LI1_cond $X=1.68 $Y=2.862
+ $X2=2.16 $Y2=2.862
r61 14 24 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=2.68 $Y=2.155
+ $X2=2.68 $Y2=2.735
r62 11 14 851.191 $w=1.5e-07 $l=1.66e-06 $layer=POLY_cond $X=2.68 $Y=0.495
+ $X2=2.68 $Y2=2.155
r63 7 25 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.425 $Y=2.99
+ $X2=2.59 $Y2=2.99
r64 7 8 943.489 $w=1.5e-07 $l=1.84e-06 $layer=POLY_cond $X=2.425 $Y=2.99
+ $X2=0.585 $Y2=2.99
r65 3 6 856.319 $w=1.5e-07 $l=1.67e-06 $layer=POLY_cond $X=0.51 $Y=0.495
+ $X2=0.51 $Y2=2.165
r66 1 8 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.51 $Y=2.915
+ $X2=0.585 $Y2=2.99
r67 1 6 384.574 $w=1.5e-07 $l=7.5e-07 $layer=POLY_cond $X=0.51 $Y=2.915 $X2=0.51
+ $Y2=2.165
.ends

.subckt PM_SKY130_FD_SC_LP__MAJ3_1%A_30_57# 1 2 3 4 15 19 23 29 32 34 37 40 42
+ 43 45 52 53 55 59
c90 45 0 6.76105e-20 $X=1.99 $Y=2.01
c91 19 0 1.46302e-19 $X=3.345 $Y=2.465
r92 58 59 6.99445 $w=3.3e-07 $l=4e-08 $layer=POLY_cond $X=3.305 $Y=1.49
+ $X2=3.345 $Y2=1.49
r93 51 53 7.65138 $w=6.78e-07 $l=4.35e-07 $layer=LI1_cond $X=2.105 $Y=0.605
+ $X2=2.54 $Y2=0.605
r94 51 52 10.6764 $w=6.78e-07 $l=1.65e-07 $layer=LI1_cond $X=2.105 $Y=0.605
+ $X2=1.94 $Y2=0.605
r95 45 48 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=1.99 $Y=2.01
+ $X2=1.99 $Y2=2.16
r96 42 43 10.7321 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=0.295 $Y=2.165
+ $X2=0.295 $Y2=1.935
r97 38 58 30.6007 $w=3.3e-07 $l=1.75e-07 $layer=POLY_cond $X=3.13 $Y=1.49
+ $X2=3.305 $Y2=1.49
r98 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.13
+ $Y=1.49 $X2=3.13 $Y2=1.49
r99 35 55 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.625 $Y=1.49
+ $X2=2.54 $Y2=1.49
r100 35 37 17.6359 $w=3.28e-07 $l=5.05e-07 $layer=LI1_cond $X=2.625 $Y=1.49
+ $X2=3.13 $Y2=1.49
r101 33 55 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.54 $Y=1.655
+ $X2=2.54 $Y2=1.49
r102 33 34 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=2.54 $Y=1.655
+ $X2=2.54 $Y2=1.925
r103 32 55 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.54 $Y=1.325
+ $X2=2.54 $Y2=1.49
r104 31 53 9.13095 $w=1.7e-07 $l=3.4e-07 $layer=LI1_cond $X=2.54 $Y=0.945
+ $X2=2.54 $Y2=0.605
r105 31 32 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=2.54 $Y=0.945
+ $X2=2.54 $Y2=1.325
r106 30 45 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.155 $Y=2.01
+ $X2=1.99 $Y2=2.01
r107 29 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.455 $Y=2.01
+ $X2=2.54 $Y2=1.925
r108 29 30 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=2.455 $Y=2.01
+ $X2=2.155 $Y2=2.01
r109 28 40 2.11342 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.38 $Y=0.86
+ $X2=0.255 $Y2=0.86
r110 28 52 101.775 $w=1.68e-07 $l=1.56e-06 $layer=LI1_cond $X=0.38 $Y=0.86
+ $X2=1.94 $Y2=0.86
r111 25 40 4.3182 $w=2.1e-07 $l=1.03078e-07 $layer=LI1_cond $X=0.215 $Y=0.945
+ $X2=0.255 $Y2=0.86
r112 25 43 64.5882 $w=1.68e-07 $l=9.9e-07 $layer=LI1_cond $X=0.215 $Y=0.945
+ $X2=0.215 $Y2=1.935
r113 21 40 4.3182 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=0.255 $Y=0.775
+ $X2=0.255 $Y2=0.86
r114 21 23 12.9074 $w=2.48e-07 $l=2.8e-07 $layer=LI1_cond $X=0.255 $Y=0.775
+ $X2=0.255 $Y2=0.495
r115 17 59 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.345 $Y=1.655
+ $X2=3.345 $Y2=1.49
r116 17 19 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=3.345 $Y=1.655
+ $X2=3.345 $Y2=2.465
r117 13 58 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.305 $Y=1.325
+ $X2=3.305 $Y2=1.49
r118 13 15 317.915 $w=1.5e-07 $l=6.2e-07 $layer=POLY_cond $X=3.305 $Y=1.325
+ $X2=3.305 $Y2=0.705
r119 4 48 600 $w=1.7e-07 $l=3.42491e-07 $layer=licon1_PDIFF $count=1 $X=1.735
+ $Y=1.955 $X2=1.99 $Y2=2.16
r120 3 42 600 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=1 $X=0.15
+ $Y=1.955 $X2=0.295 $Y2=2.165
r121 2 51 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.965
+ $Y=0.285 $X2=2.105 $Y2=0.495
r122 1 23 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.15
+ $Y=0.285 $X2=0.295 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__MAJ3_1%VPWR 1 2 9 13 17 19 24 31 32 35 38
r36 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r37 35 36 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r38 32 39 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=3.12 $Y2=3.33
r39 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r40 29 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.295 $Y=3.33
+ $X2=3.13 $Y2=3.33
r41 29 31 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3.295 $Y=3.33
+ $X2=3.6 $Y2=3.33
r42 28 39 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r43 27 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r44 25 35 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.25 $Y=3.33
+ $X2=1.085 $Y2=3.33
r45 25 27 90.6845 $w=1.68e-07 $l=1.39e-06 $layer=LI1_cond $X=1.25 $Y=3.33
+ $X2=2.64 $Y2=3.33
r46 24 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.965 $Y=3.33
+ $X2=3.13 $Y2=3.33
r47 24 27 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=2.965 $Y=3.33
+ $X2=2.64 $Y2=3.33
r48 22 36 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r49 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r50 19 35 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.92 $Y=3.33
+ $X2=1.085 $Y2=3.33
r51 19 21 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=0.92 $Y=3.33 $X2=0.72
+ $Y2=3.33
r52 17 28 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=2.64 $Y2=3.33
r53 17 36 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=3.33
+ $X2=1.2 $Y2=3.33
r54 13 16 16.239 $w=3.28e-07 $l=4.65e-07 $layer=LI1_cond $X=3.13 $Y=2 $X2=3.13
+ $Y2=2.465
r55 11 38 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.13 $Y=3.245
+ $X2=3.13 $Y2=3.33
r56 11 16 27.2396 $w=3.28e-07 $l=7.8e-07 $layer=LI1_cond $X=3.13 $Y=3.245
+ $X2=3.13 $Y2=2.465
r57 7 35 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.085 $Y=3.245
+ $X2=1.085 $Y2=3.33
r58 7 9 37.7163 $w=3.28e-07 $l=1.08e-06 $layer=LI1_cond $X=1.085 $Y=3.245
+ $X2=1.085 $Y2=2.165
r59 2 16 300 $w=1.7e-07 $l=6.82202e-07 $layer=licon1_PDIFF $count=2 $X=2.755
+ $Y=1.945 $X2=3.13 $Y2=2.465
r60 2 13 600 $w=1.7e-07 $l=4.01559e-07 $layer=licon1_PDIFF $count=1 $X=2.755
+ $Y=1.945 $X2=3.13 $Y2=2
r61 1 9 600 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_PDIFF $count=1 $X=0.945
+ $Y=1.955 $X2=1.085 $Y2=2.165
.ends

.subckt PM_SKY130_FD_SC_LP__MAJ3_1%X 1 2 7 8 9 10 11 12 13 24 30
r16 22 30 1.09015 $w=3.68e-07 $l=3.5e-08 $layer=LI1_cond $X=3.54 $Y=0.96
+ $X2=3.54 $Y2=0.925
r17 13 44 5.76222 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=3.6 $Y=2.775
+ $X2=3.6 $Y2=2.9
r18 12 13 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=3.6 $Y=2.405 $X2=3.6
+ $Y2=2.775
r19 11 12 20.5135 $w=2.48e-07 $l=4.45e-07 $layer=LI1_cond $X=3.6 $Y=1.96 $X2=3.6
+ $Y2=2.405
r20 10 11 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=3.6 $Y=1.665
+ $X2=3.6 $Y2=1.96
r21 9 10 17.0562 $w=2.48e-07 $l=3.7e-07 $layer=LI1_cond $X=3.6 $Y=1.295 $X2=3.6
+ $Y2=1.665
r22 9 47 6.91466 $w=2.48e-07 $l=1.5e-07 $layer=LI1_cond $X=3.6 $Y=1.295 $X2=3.6
+ $Y2=1.145
r23 8 47 6.20149 $w=3.68e-07 $l=1.6e-07 $layer=LI1_cond $X=3.54 $Y=0.985
+ $X2=3.54 $Y2=1.145
r24 8 22 0.778678 $w=3.68e-07 $l=2.5e-08 $layer=LI1_cond $X=3.54 $Y=0.985
+ $X2=3.54 $Y2=0.96
r25 8 30 0.778678 $w=3.68e-07 $l=2.5e-08 $layer=LI1_cond $X=3.54 $Y=0.9 $X2=3.54
+ $Y2=0.925
r26 7 8 10.7458 $w=3.68e-07 $l=3.45e-07 $layer=LI1_cond $X=3.54 $Y=0.555
+ $X2=3.54 $Y2=0.9
r27 7 24 3.89339 $w=3.68e-07 $l=1.25e-07 $layer=LI1_cond $X=3.54 $Y=0.555
+ $X2=3.54 $Y2=0.43
r28 2 44 400 $w=1.7e-07 $l=1.13284e-06 $layer=licon1_PDIFF $count=1 $X=3.42
+ $Y=1.835 $X2=3.56 $Y2=2.9
r29 2 11 400 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=3.42
+ $Y=1.835 $X2=3.56 $Y2=1.96
r30 1 24 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.38
+ $Y=0.285 $X2=3.52 $Y2=0.43
.ends

.subckt PM_SKY130_FD_SC_LP__MAJ3_1%VGND 1 2 9 13 18 19 20 22 35 36 39
r44 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r45 35 36 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r46 33 36 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r47 32 33 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r48 30 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r49 29 32 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r50 29 30 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r51 27 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.4 $Y=0 $X2=1.235
+ $Y2=0
r52 27 29 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=1.4 $Y=0 $X2=1.68
+ $Y2=0
r53 25 40 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r54 24 25 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r55 22 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.07 $Y=0 $X2=1.235
+ $Y2=0
r56 22 24 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=1.07 $Y=0 $X2=0.72
+ $Y2=0
r57 20 33 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=2.64
+ $Y2=0
r58 20 30 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=1.92 $Y=0 $X2=1.68
+ $Y2=0
r59 18 32 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=2.845 $Y=0 $X2=2.64
+ $Y2=0
r60 18 19 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.845 $Y=0 $X2=3.01
+ $Y2=0
r61 17 35 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=3.175 $Y=0 $X2=3.6
+ $Y2=0
r62 17 19 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.175 $Y=0 $X2=3.01
+ $Y2=0
r63 13 15 19.2074 $w=3.28e-07 $l=5.5e-07 $layer=LI1_cond $X=3.01 $Y=0.43
+ $X2=3.01 $Y2=0.98
r64 11 19 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.01 $Y=0.085
+ $X2=3.01 $Y2=0
r65 11 13 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=3.01 $Y=0.085
+ $X2=3.01 $Y2=0.43
r66 7 39 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.235 $Y=0.085
+ $X2=1.235 $Y2=0
r67 7 9 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=1.235 $Y=0.085
+ $X2=1.235 $Y2=0.43
r68 2 15 182 $w=1.7e-07 $l=8.12558e-07 $layer=licon1_NDIFF $count=1 $X=2.755
+ $Y=0.285 $X2=3.01 $Y2=0.98
r69 2 13 182 $w=1.7e-07 $l=3.19374e-07 $layer=licon1_NDIFF $count=1 $X=2.755
+ $Y=0.285 $X2=3.01 $Y2=0.43
r70 1 9 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=1.095
+ $Y=0.285 $X2=1.235 $Y2=0.43
.ends

