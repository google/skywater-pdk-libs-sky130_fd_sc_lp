* File: sky130_fd_sc_lp__a2bb2oi_0.pxi.spice
* Created: Wed Sep  2 09:24:16 2020
* 
x_PM_SKY130_FD_SC_LP__A2BB2OI_0%A1_N N_A1_N_c_64_n N_A1_N_M1003_g N_A1_N_M1007_g
+ N_A1_N_c_67_n A1_N A1_N A1_N N_A1_N_c_69_n PM_SKY130_FD_SC_LP__A2BB2OI_0%A1_N
x_PM_SKY130_FD_SC_LP__A2BB2OI_0%A2_N N_A2_N_M1005_g N_A2_N_M1006_g A2_N A2_N
+ N_A2_N_c_94_n N_A2_N_c_95_n PM_SKY130_FD_SC_LP__A2BB2OI_0%A2_N
x_PM_SKY130_FD_SC_LP__A2BB2OI_0%A_110_47# N_A_110_47#_M1003_d
+ N_A_110_47#_M1005_d N_A_110_47#_c_132_n N_A_110_47#_M1008_g
+ N_A_110_47#_c_134_n N_A_110_47#_M1009_g N_A_110_47#_c_135_n
+ N_A_110_47#_c_129_n N_A_110_47#_c_136_n N_A_110_47#_c_185_p
+ N_A_110_47#_c_130_n N_A_110_47#_c_131_n
+ PM_SKY130_FD_SC_LP__A2BB2OI_0%A_110_47#
x_PM_SKY130_FD_SC_LP__A2BB2OI_0%B2 N_B2_M1000_g N_B2_M1004_g N_B2_c_192_n
+ N_B2_c_193_n B2 B2 N_B2_c_195_n PM_SKY130_FD_SC_LP__A2BB2OI_0%B2
x_PM_SKY130_FD_SC_LP__A2BB2OI_0%B1 N_B1_M1002_g N_B1_M1001_g N_B1_c_233_n
+ N_B1_c_234_n B1 B1 N_B1_c_236_n PM_SKY130_FD_SC_LP__A2BB2OI_0%B1
x_PM_SKY130_FD_SC_LP__A2BB2OI_0%VPWR N_VPWR_M1007_s N_VPWR_M1004_d
+ N_VPWR_c_261_n N_VPWR_c_262_n N_VPWR_c_263_n VPWR N_VPWR_c_264_n
+ N_VPWR_c_265_n N_VPWR_c_260_n N_VPWR_c_267_n
+ PM_SKY130_FD_SC_LP__A2BB2OI_0%VPWR
x_PM_SKY130_FD_SC_LP__A2BB2OI_0%Y N_Y_M1008_d N_Y_M1009_s N_Y_c_309_n Y Y Y Y Y
+ Y N_Y_c_301_n Y Y PM_SKY130_FD_SC_LP__A2BB2OI_0%Y
x_PM_SKY130_FD_SC_LP__A2BB2OI_0%A_420_387# N_A_420_387#_M1009_d
+ N_A_420_387#_M1001_d N_A_420_387#_c_344_n N_A_420_387#_c_342_n
+ N_A_420_387#_c_343_n N_A_420_387#_c_347_n
+ PM_SKY130_FD_SC_LP__A2BB2OI_0%A_420_387#
x_PM_SKY130_FD_SC_LP__A2BB2OI_0%VGND N_VGND_M1003_s N_VGND_M1006_d
+ N_VGND_M1002_d N_VGND_c_370_n N_VGND_c_371_n N_VGND_c_372_n N_VGND_c_373_n
+ VGND N_VGND_c_374_n N_VGND_c_375_n N_VGND_c_376_n
+ PM_SKY130_FD_SC_LP__A2BB2OI_0%VGND
cc_1 VNB N_A1_N_c_64_n 0.0207126f $X=-0.19 $Y=-0.245 $X2=0.327 $Y2=1.288
cc_2 VNB N_A1_N_M1003_g 0.0282237f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.445
cc_3 VNB N_A1_N_M1007_g 0.00872834f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.455
cc_4 VNB N_A1_N_c_67_n 0.028948f $X=-0.19 $Y=-0.245 $X2=0.327 $Y2=1.51
cc_5 VNB A1_N 0.034183f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_6 VNB N_A1_N_c_69_n 0.028948f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.005
cc_7 VNB N_A2_N_M1005_g 0.0123577f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.84
cc_8 VNB A2_N 0.00293821f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.455
cc_9 VNB N_A2_N_c_94_n 0.0879857f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_10 VNB N_A2_N_c_95_n 0.0222618f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_110_47#_M1008_g 0.0701433f $X=-0.19 $Y=-0.245 $X2=0.327 $Y2=1.51
cc_12 VNB N_A_110_47#_c_129_n 0.00781153f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.005
cc_13 VNB N_A_110_47#_c_130_n 0.00245708f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_14 VNB N_A_110_47#_c_131_n 0.0100721f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_B2_M1000_g 0.0195676f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.84
cc_16 VNB N_B2_M1004_g 0.0103766f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.51
cc_17 VNB N_B2_c_192_n 0.0196784f $X=-0.19 $Y=-0.245 $X2=0.327 $Y2=1.51
cc_18 VNB N_B2_c_193_n 0.0147436f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_19 VNB B2 0.0175203f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_20 VNB N_B2_c_195_n 0.0147436f $X=-0.19 $Y=-0.245 $X2=0.327 $Y2=1.005
cc_21 VNB N_B1_M1002_g 0.025294f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.84
cc_22 VNB N_B1_M1001_g 0.0144909f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.51
cc_23 VNB N_B1_c_233_n 0.0275318f $X=-0.19 $Y=-0.245 $X2=0.327 $Y2=1.51
cc_24 VNB N_B1_c_234_n 0.0185186f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_25 VNB B1 0.0331792f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_26 VNB N_B1_c_236_n 0.0185778f $X=-0.19 $Y=-0.245 $X2=0.327 $Y2=1.005
cc_27 VNB N_VPWR_c_260_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB Y 0.0123665f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_29 VNB N_Y_c_301_n 0.0039352f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A_420_387#_c_342_n 0.0114511f $X=-0.19 $Y=-0.245 $X2=0.327 $Y2=1.51
cc_31 VNB N_A_420_387#_c_343_n 0.00183194f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_32 VNB N_VGND_c_370_n 0.0107842f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_371_n 0.0191775f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_34 VNB N_VGND_c_372_n 0.011138f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_35 VNB N_VGND_c_373_n 0.0174842f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_374_n 0.0338112f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.005
cc_37 VNB N_VGND_c_375_n 0.037253f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.295
cc_38 VNB N_VGND_c_376_n 0.187043f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VPB N_A1_N_M1007_g 0.0464428f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.455
cc_40 VPB A1_N 0.0115654f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_41 VPB N_A2_N_M1005_g 0.0333749f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.84
cc_42 VPB N_A_110_47#_c_132_n 0.0284274f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=1.51
cc_43 VPB N_A_110_47#_M1008_g 4.91864e-19 $X=-0.19 $Y=1.655 $X2=0.327 $Y2=1.51
cc_44 VPB N_A_110_47#_c_134_n 0.0193339f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_45 VPB N_A_110_47#_c_135_n 0.0167788f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_46 VPB N_A_110_47#_c_136_n 0.0125478f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_47 VPB N_A_110_47#_c_130_n 0.0129662f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_48 VPB N_A_110_47#_c_131_n 0.0301047f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_49 VPB N_B2_M1004_g 0.0245145f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=1.51
cc_50 VPB N_B1_M1001_g 0.0303213f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=1.51
cc_51 VPB N_VPWR_c_261_n 0.0115529f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=1.51
cc_52 VPB N_VPWR_c_262_n 0.0540948f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.455
cc_53 VPB N_VPWR_c_263_n 0.0314903f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_54 VPB N_VPWR_c_264_n 0.0608278f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_55 VPB N_VPWR_c_265_n 0.0179326f $X=-0.19 $Y=1.655 $X2=0.27 $Y2=1.665
cc_56 VPB N_VPWR_c_260_n 0.096528f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_57 VPB N_VPWR_c_267_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_58 VPB Y 0.00127078f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_59 VPB Y 0.0280374f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_60 VPB N_A_420_387#_c_344_n 0.00602862f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.455
cc_61 VPB N_A_420_387#_c_342_n 0.01319f $X=-0.19 $Y=1.655 $X2=0.327 $Y2=1.51
cc_62 VPB N_A_420_387#_c_343_n 0.00158627f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_63 VPB N_A_420_387#_c_347_n 0.0346418f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_64 N_A1_N_c_64_n N_A2_N_M1005_g 0.0636233f $X=0.327 $Y=1.288 $X2=0 $Y2=0
cc_65 N_A1_N_M1003_g N_A2_N_c_94_n 0.0636233f $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_66 A1_N N_A2_N_c_94_n 6.66073e-19 $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_67 N_A1_N_M1003_g N_A2_N_c_95_n 0.0116011f $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_68 N_A1_N_M1003_g N_A_110_47#_c_129_n 0.0106606f $X=0.475 $Y=0.445 $X2=0
+ $Y2=0
cc_69 A1_N N_A_110_47#_c_129_n 0.0617871f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_70 N_A1_N_M1007_g N_A_110_47#_c_136_n 0.00174197f $X=0.475 $Y=2.455 $X2=0
+ $Y2=0
cc_71 N_A1_N_M1007_g N_A_110_47#_c_130_n 0.0098514f $X=0.475 $Y=2.455 $X2=0
+ $Y2=0
cc_72 A1_N N_A_110_47#_c_130_n 0.0164878f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_73 N_A1_N_M1007_g N_VPWR_c_262_n 0.0165019f $X=0.475 $Y=2.455 $X2=0 $Y2=0
cc_74 N_A1_N_c_67_n N_VPWR_c_262_n 0.00119546f $X=0.327 $Y=1.51 $X2=0 $Y2=0
cc_75 A1_N N_VPWR_c_262_n 0.0217025f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_76 N_A1_N_M1007_g N_VPWR_c_264_n 0.00377474f $X=0.475 $Y=2.455 $X2=0 $Y2=0
cc_77 N_A1_N_M1007_g N_VPWR_c_260_n 0.00410937f $X=0.475 $Y=2.455 $X2=0 $Y2=0
cc_78 N_A1_N_M1003_g N_VGND_c_371_n 0.00369776f $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_79 A1_N N_VGND_c_371_n 0.0175586f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_80 N_A1_N_c_69_n N_VGND_c_371_n 0.00195491f $X=0.27 $Y=1.005 $X2=0 $Y2=0
cc_81 N_A1_N_M1003_g N_VGND_c_374_n 0.00585385f $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_82 N_A1_N_M1003_g N_VGND_c_376_n 0.0101809f $X=0.475 $Y=0.445 $X2=0 $Y2=0
cc_83 A1_N N_VGND_c_376_n 0.00372952f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_84 A2_N N_A_110_47#_M1008_g 5.94669e-19 $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_85 N_A2_N_c_94_n N_A_110_47#_M1008_g 0.0146965f $X=1.2 $Y=0.93 $X2=0 $Y2=0
cc_86 N_A2_N_M1005_g N_A_110_47#_c_129_n 0.0106927f $X=0.835 $Y=2.455 $X2=0
+ $Y2=0
cc_87 A2_N N_A_110_47#_c_129_n 0.0478059f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_88 N_A2_N_c_94_n N_A_110_47#_c_129_n 0.0191038f $X=1.2 $Y=0.93 $X2=0 $Y2=0
cc_89 N_A2_N_c_95_n N_A_110_47#_c_129_n 0.00296311f $X=1.062 $Y=0.765 $X2=0
+ $Y2=0
cc_90 N_A2_N_M1005_g N_A_110_47#_c_136_n 0.010989f $X=0.835 $Y=2.455 $X2=0 $Y2=0
cc_91 N_A2_N_M1005_g N_A_110_47#_c_130_n 0.0274567f $X=0.835 $Y=2.455 $X2=0
+ $Y2=0
cc_92 A2_N N_A_110_47#_c_130_n 0.0258325f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_93 N_A2_N_c_94_n N_A_110_47#_c_130_n 0.00540812f $X=1.2 $Y=0.93 $X2=0 $Y2=0
cc_94 N_A2_N_M1005_g N_A_110_47#_c_131_n 0.018116f $X=0.835 $Y=2.455 $X2=0 $Y2=0
cc_95 A2_N N_A_110_47#_c_131_n 7.44118e-19 $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_96 N_A2_N_c_94_n N_A_110_47#_c_131_n 0.0135905f $X=1.2 $Y=0.93 $X2=0 $Y2=0
cc_97 N_A2_N_M1005_g N_VPWR_c_262_n 0.00233081f $X=0.835 $Y=2.455 $X2=0 $Y2=0
cc_98 N_A2_N_M1005_g N_VPWR_c_264_n 0.00436277f $X=0.835 $Y=2.455 $X2=0 $Y2=0
cc_99 N_A2_N_M1005_g N_VPWR_c_260_n 0.00489211f $X=0.835 $Y=2.455 $X2=0 $Y2=0
cc_100 N_A2_N_M1005_g Y 0.00471814f $X=0.835 $Y=2.455 $X2=0 $Y2=0
cc_101 A2_N Y 0.0451856f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_102 N_A2_N_c_94_n Y 0.00615761f $X=1.2 $Y=0.93 $X2=0 $Y2=0
cc_103 N_A2_N_M1005_g Y 0.00442224f $X=0.835 $Y=2.455 $X2=0 $Y2=0
cc_104 N_A2_N_c_94_n N_Y_c_301_n 2.76648e-19 $X=1.2 $Y=0.93 $X2=0 $Y2=0
cc_105 A2_N N_VGND_c_374_n 0.0291411f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_106 N_A2_N_c_94_n N_VGND_c_374_n 0.0103869f $X=1.2 $Y=0.93 $X2=0 $Y2=0
cc_107 N_A2_N_c_95_n N_VGND_c_374_n 0.00960456f $X=1.062 $Y=0.765 $X2=0 $Y2=0
cc_108 A2_N N_VGND_c_376_n 0.00130731f $X=1.115 $Y=0.84 $X2=0 $Y2=0
cc_109 N_A2_N_c_94_n N_VGND_c_376_n 5.56241e-19 $X=1.2 $Y=0.93 $X2=0 $Y2=0
cc_110 N_A2_N_c_95_n N_VGND_c_376_n 0.0121919f $X=1.062 $Y=0.765 $X2=0 $Y2=0
cc_111 N_A_110_47#_M1008_g N_B2_M1000_g 0.0146171f $X=1.9 $Y=0.445 $X2=0 $Y2=0
cc_112 N_A_110_47#_M1008_g N_B2_M1004_g 0.00572225f $X=1.9 $Y=0.445 $X2=0 $Y2=0
cc_113 N_A_110_47#_c_135_n N_B2_M1004_g 0.0160381f $X=2.025 $Y=1.74 $X2=0 $Y2=0
cc_114 N_A_110_47#_M1008_g B2 0.00477631f $X=1.9 $Y=0.445 $X2=0 $Y2=0
cc_115 N_A_110_47#_c_135_n B2 0.00207515f $X=2.025 $Y=1.74 $X2=0 $Y2=0
cc_116 N_A_110_47#_M1008_g N_B2_c_195_n 0.0329726f $X=1.9 $Y=0.445 $X2=0 $Y2=0
cc_117 N_A_110_47#_c_136_n N_VPWR_c_262_n 0.0214127f $X=1.05 $Y=2.29 $X2=0 $Y2=0
cc_118 N_A_110_47#_c_130_n N_VPWR_c_262_n 0.00287649f $X=1.315 $Y=1.81 $X2=0
+ $Y2=0
cc_119 N_A_110_47#_c_134_n N_VPWR_c_263_n 5.01764e-19 $X=2.025 $Y=1.815 $X2=0
+ $Y2=0
cc_120 N_A_110_47#_c_134_n N_VPWR_c_264_n 0.00352953f $X=2.025 $Y=1.815 $X2=0
+ $Y2=0
cc_121 N_A_110_47#_c_136_n N_VPWR_c_264_n 0.0082118f $X=1.05 $Y=2.29 $X2=0 $Y2=0
cc_122 N_A_110_47#_c_134_n N_VPWR_c_260_n 0.00434946f $X=2.025 $Y=1.815 $X2=0
+ $Y2=0
cc_123 N_A_110_47#_c_136_n N_VPWR_c_260_n 0.0106498f $X=1.05 $Y=2.29 $X2=0 $Y2=0
cc_124 N_A_110_47#_c_130_n A_110_427# 0.00356976f $X=1.315 $Y=1.81 $X2=-0.19
+ $Y2=-0.245
cc_125 N_A_110_47#_M1008_g N_Y_c_309_n 0.0160675f $X=1.9 $Y=0.445 $X2=0 $Y2=0
cc_126 N_A_110_47#_c_132_n Y 0.0178116f $X=1.825 $Y=1.74 $X2=0 $Y2=0
cc_127 N_A_110_47#_M1008_g Y 0.0256479f $X=1.9 $Y=0.445 $X2=0 $Y2=0
cc_128 N_A_110_47#_c_134_n Y 0.00102544f $X=2.025 $Y=1.815 $X2=0 $Y2=0
cc_129 N_A_110_47#_c_135_n Y 0.00398468f $X=2.025 $Y=1.74 $X2=0 $Y2=0
cc_130 N_A_110_47#_c_130_n Y 0.0428221f $X=1.315 $Y=1.81 $X2=0 $Y2=0
cc_131 N_A_110_47#_c_131_n Y 0.00183349f $X=1.48 $Y=1.81 $X2=0 $Y2=0
cc_132 N_A_110_47#_c_134_n Y 0.00398971f $X=2.025 $Y=1.815 $X2=0 $Y2=0
cc_133 N_A_110_47#_c_135_n Y 0.00255832f $X=2.025 $Y=1.74 $X2=0 $Y2=0
cc_134 N_A_110_47#_c_136_n Y 0.0322772f $X=1.05 $Y=2.29 $X2=0 $Y2=0
cc_135 N_A_110_47#_M1008_g N_Y_c_301_n 0.00640185f $X=1.9 $Y=0.445 $X2=0 $Y2=0
cc_136 N_A_110_47#_c_134_n N_A_420_387#_c_344_n 0.00119014f $X=2.025 $Y=1.815
+ $X2=0 $Y2=0
cc_137 N_A_110_47#_c_135_n N_A_420_387#_c_343_n 0.00181949f $X=2.025 $Y=1.74
+ $X2=0 $Y2=0
cc_138 N_A_110_47#_M1008_g N_VGND_c_374_n 0.00643531f $X=1.9 $Y=0.445 $X2=0
+ $Y2=0
cc_139 N_A_110_47#_c_185_p N_VGND_c_374_n 0.0133089f $X=0.69 $Y=0.445 $X2=0
+ $Y2=0
cc_140 N_A_110_47#_M1008_g N_VGND_c_375_n 0.00362032f $X=1.9 $Y=0.445 $X2=0
+ $Y2=0
cc_141 N_A_110_47#_M1003_d N_VGND_c_376_n 0.00246193f $X=0.55 $Y=0.235 $X2=0
+ $Y2=0
cc_142 N_A_110_47#_M1008_g N_VGND_c_376_n 0.0068533f $X=1.9 $Y=0.445 $X2=0 $Y2=0
cc_143 N_A_110_47#_c_185_p N_VGND_c_376_n 0.0104333f $X=0.69 $Y=0.445 $X2=0
+ $Y2=0
cc_144 N_B2_M1000_g N_B1_M1002_g 0.0226329f $X=2.33 $Y=0.445 $X2=0 $Y2=0
cc_145 B2 N_B1_M1002_g 0.00514384f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_146 N_B2_M1004_g N_B1_M1001_g 0.0271215f $X=2.455 $Y=2.255 $X2=0 $Y2=0
cc_147 N_B2_c_192_n N_B1_c_233_n 0.0118752f $X=2.38 $Y=1.31 $X2=0 $Y2=0
cc_148 N_B2_c_193_n N_B1_c_234_n 0.0118752f $X=2.38 $Y=1.475 $X2=0 $Y2=0
cc_149 B2 B1 0.0364245f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_150 N_B2_c_195_n B1 7.496e-19 $X=2.38 $Y=0.97 $X2=0 $Y2=0
cc_151 N_B2_c_195_n N_B1_c_236_n 0.0118752f $X=2.38 $Y=0.97 $X2=0 $Y2=0
cc_152 N_B2_M1004_g N_VPWR_c_263_n 0.0105766f $X=2.455 $Y=2.255 $X2=0 $Y2=0
cc_153 N_B2_M1004_g N_VPWR_c_264_n 0.00293417f $X=2.455 $Y=2.255 $X2=0 $Y2=0
cc_154 N_B2_M1004_g N_VPWR_c_260_n 0.00365355f $X=2.455 $Y=2.255 $X2=0 $Y2=0
cc_155 N_B2_M1000_g N_Y_c_309_n 0.00709441f $X=2.33 $Y=0.445 $X2=0 $Y2=0
cc_156 B2 N_Y_c_309_n 0.0163729f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_157 N_B2_M1004_g Y 9.41121e-19 $X=2.455 $Y=2.255 $X2=0 $Y2=0
cc_158 N_B2_c_192_n Y 2.76722e-19 $X=2.38 $Y=1.31 $X2=0 $Y2=0
cc_159 B2 Y 0.0566001f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_160 N_B2_c_195_n Y 2.76722e-19 $X=2.38 $Y=0.97 $X2=0 $Y2=0
cc_161 N_B2_M1000_g N_Y_c_301_n 8.22435e-19 $X=2.33 $Y=0.445 $X2=0 $Y2=0
cc_162 N_B2_M1004_g N_A_420_387#_c_344_n 0.00317376f $X=2.455 $Y=2.255 $X2=0
+ $Y2=0
cc_163 N_B2_M1004_g N_A_420_387#_c_342_n 0.0140077f $X=2.455 $Y=2.255 $X2=0
+ $Y2=0
cc_164 N_B2_c_193_n N_A_420_387#_c_342_n 4.15267e-19 $X=2.38 $Y=1.475 $X2=0
+ $Y2=0
cc_165 B2 N_A_420_387#_c_342_n 0.0165513f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_166 N_B2_c_193_n N_A_420_387#_c_343_n 9.38777e-19 $X=2.38 $Y=1.475 $X2=0
+ $Y2=0
cc_167 B2 N_A_420_387#_c_343_n 0.0210391f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_168 N_B2_M1000_g N_VGND_c_373_n 0.00212557f $X=2.33 $Y=0.445 $X2=0 $Y2=0
cc_169 N_B2_M1000_g N_VGND_c_375_n 0.00548159f $X=2.33 $Y=0.445 $X2=0 $Y2=0
cc_170 N_B2_M1000_g N_VGND_c_376_n 0.00651572f $X=2.33 $Y=0.445 $X2=0 $Y2=0
cc_171 B2 N_VGND_c_376_n 0.0106805f $X=2.075 $Y=0.84 $X2=0 $Y2=0
cc_172 N_B1_M1001_g N_VPWR_c_263_n 0.013846f $X=2.885 $Y=2.255 $X2=0 $Y2=0
cc_173 N_B1_M1001_g N_VPWR_c_265_n 0.00293417f $X=2.885 $Y=2.255 $X2=0 $Y2=0
cc_174 N_B1_M1001_g N_VPWR_c_260_n 0.00365355f $X=2.885 $Y=2.255 $X2=0 $Y2=0
cc_175 N_B1_M1002_g N_Y_c_309_n 0.00103192f $X=2.86 $Y=0.445 $X2=0 $Y2=0
cc_176 N_B1_M1001_g N_A_420_387#_c_342_n 0.0173873f $X=2.885 $Y=2.255 $X2=0
+ $Y2=0
cc_177 N_B1_c_234_n N_A_420_387#_c_342_n 0.00220138f $X=2.95 $Y=1.475 $X2=0
+ $Y2=0
cc_178 B1 N_A_420_387#_c_342_n 0.0345462f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_179 N_B1_M1001_g N_A_420_387#_c_347_n 0.00527749f $X=2.885 $Y=2.255 $X2=0
+ $Y2=0
cc_180 N_B1_M1002_g N_VGND_c_373_n 0.013834f $X=2.86 $Y=0.445 $X2=0 $Y2=0
cc_181 B1 N_VGND_c_373_n 0.0265987f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_182 N_B1_c_236_n N_VGND_c_373_n 0.00114754f $X=2.95 $Y=0.97 $X2=0 $Y2=0
cc_183 N_B1_M1002_g N_VGND_c_375_n 0.00486043f $X=2.86 $Y=0.445 $X2=0 $Y2=0
cc_184 N_B1_M1002_g N_VGND_c_376_n 0.0072416f $X=2.86 $Y=0.445 $X2=0 $Y2=0
cc_185 B1 N_VGND_c_376_n 0.00428397f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_186 N_VPWR_c_263_n Y 0.0123797f $X=2.67 $Y=2.07 $X2=0 $Y2=0
cc_187 N_VPWR_c_264_n Y 0.0144531f $X=2.505 $Y=3.33 $X2=0 $Y2=0
cc_188 N_VPWR_c_260_n Y 0.0131616f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_189 N_VPWR_c_263_n N_A_420_387#_c_344_n 0.0236371f $X=2.67 $Y=2.07 $X2=0
+ $Y2=0
cc_190 N_VPWR_c_264_n N_A_420_387#_c_344_n 0.00380048f $X=2.505 $Y=3.33 $X2=0
+ $Y2=0
cc_191 N_VPWR_c_260_n N_A_420_387#_c_344_n 0.00642502f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_192 N_VPWR_c_263_n N_A_420_387#_c_342_n 0.0216087f $X=2.67 $Y=2.07 $X2=0
+ $Y2=0
cc_193 N_VPWR_c_263_n N_A_420_387#_c_347_n 0.0225912f $X=2.67 $Y=2.07 $X2=0
+ $Y2=0
cc_194 N_VPWR_c_265_n N_A_420_387#_c_347_n 0.00413386f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_195 N_VPWR_c_260_n N_A_420_387#_c_347_n 0.00698862f $X=3.12 $Y=3.33 $X2=0
+ $Y2=0
cc_196 Y N_A_420_387#_c_344_n 0.00666735f $X=1.595 $Y=0.84 $X2=0 $Y2=0
cc_197 Y N_A_420_387#_c_344_n 0.00310207f $X=1.595 $Y=1.95 $X2=0 $Y2=0
cc_198 Y N_A_420_387#_c_343_n 0.011749f $X=1.595 $Y=0.84 $X2=0 $Y2=0
cc_199 N_Y_c_309_n N_VGND_M1006_d 0.0043579f $X=2.115 $Y=0.445 $X2=0 $Y2=0
cc_200 N_Y_c_301_n N_VGND_M1006_d 0.00186668f $X=1.727 $Y=0.78 $X2=0 $Y2=0
cc_201 N_Y_c_309_n N_VGND_c_373_n 0.00878856f $X=2.115 $Y=0.445 $X2=0 $Y2=0
cc_202 N_Y_c_309_n N_VGND_c_374_n 0.0289956f $X=2.115 $Y=0.445 $X2=0 $Y2=0
cc_203 N_Y_c_309_n N_VGND_c_375_n 0.0282143f $X=2.115 $Y=0.445 $X2=0 $Y2=0
cc_204 N_Y_M1008_d N_VGND_c_376_n 0.00225919f $X=1.975 $Y=0.235 $X2=0 $Y2=0
cc_205 N_Y_c_309_n N_VGND_c_376_n 0.0205037f $X=2.115 $Y=0.445 $X2=0 $Y2=0
cc_206 Y N_VGND_c_376_n 0.00598742f $X=1.595 $Y=0.84 $X2=0 $Y2=0
cc_207 N_VGND_c_376_n A_481_47# 0.0120342f $X=3.12 $Y=0 $X2=-0.19 $Y2=-0.245
