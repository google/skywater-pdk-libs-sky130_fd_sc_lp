* File: sky130_fd_sc_lp__o21ai_lp.pex.spice
* Created: Fri Aug 28 11:05:08 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O21AI_LP%A1 3 7 11 12 13 15 22
r33 22 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.61
+ $Y=1.29 $X2=0.61 $Y2=1.29
r34 15 23 1.96371 $w=6.68e-07 $l=1.1e-07 $layer=LI1_cond $X=0.72 $Y=1.46
+ $X2=0.61 $Y2=1.46
r35 13 23 6.60521 $w=6.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.24 $Y=1.46
+ $X2=0.61 $Y2=1.46
r36 11 22 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.61 $Y=1.63
+ $X2=0.61 $Y2=1.29
r37 11 12 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.61 $Y=1.63
+ $X2=0.61 $Y2=1.795
r38 10 22 43.0552 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.61 $Y=1.125
+ $X2=0.61 $Y2=1.29
r39 7 10 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=0.68 $Y=0.495
+ $X2=0.68 $Y2=1.125
r40 3 12 186.34 $w=2.5e-07 $l=7.5e-07 $layer=POLY_cond $X=0.65 $Y=2.545 $X2=0.65
+ $Y2=1.795
.ends

.subckt PM_SKY130_FD_SC_LP__O21AI_LP%A2 3 7 11 12 13 14 18
r39 13 14 13.0959 $w=3.28e-07 $l=3.75e-07 $layer=LI1_cond $X=1.18 $Y=1.29
+ $X2=1.18 $Y2=1.665
r40 13 18 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.18
+ $Y=1.29 $X2=1.18 $Y2=1.29
r41 11 18 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.18 $Y=1.63
+ $X2=1.18 $Y2=1.29
r42 11 12 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.18 $Y=1.63
+ $X2=1.18 $Y2=1.795
r43 10 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.18 $Y=1.125
+ $X2=1.18 $Y2=1.29
r44 7 10 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=1.27 $Y=0.495
+ $X2=1.27 $Y2=1.125
r45 3 12 186.34 $w=2.5e-07 $l=7.5e-07 $layer=POLY_cond $X=1.14 $Y=2.545 $X2=1.14
+ $Y2=1.795
.ends

.subckt PM_SKY130_FD_SC_LP__O21AI_LP%B1 3 7 11 12 13 14 18
r36 13 14 12.3476 $w=3.48e-07 $l=3.75e-07 $layer=LI1_cond $X=1.74 $Y=1.29
+ $X2=1.74 $Y2=1.665
r37 13 18 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.75
+ $Y=1.29 $X2=1.75 $Y2=1.29
r38 11 18 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.75 $Y=1.63
+ $X2=1.75 $Y2=1.29
r39 11 12 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.75 $Y=1.63
+ $X2=1.75 $Y2=1.795
r40 10 18 40.8701 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.75 $Y=1.125
+ $X2=1.75 $Y2=1.29
r41 7 10 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=1.7 $Y=0.495 $X2=1.7
+ $Y2=1.125
r42 3 12 186.34 $w=2.5e-07 $l=7.5e-07 $layer=POLY_cond $X=1.71 $Y=2.545 $X2=1.71
+ $Y2=1.795
.ends

.subckt PM_SKY130_FD_SC_LP__O21AI_LP%VPWR 1 2 7 9 13 15 17 19 32
r25 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r26 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r27 26 32 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r28 25 26 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r29 23 29 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r30 22 25 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.72 $Y=3.33 $X2=1.68
+ $Y2=3.33
r31 22 23 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r32 20 28 4.54404 $w=1.7e-07 $l=2.75e-07 $layer=LI1_cond $X=0.55 $Y=3.33
+ $X2=0.275 $Y2=3.33
r33 20 22 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=0.55 $Y=3.33
+ $X2=0.72 $Y2=3.33
r34 19 31 4.4922 $w=1.7e-07 $l=2.95e-07 $layer=LI1_cond $X=1.81 $Y=3.33
+ $X2=2.105 $Y2=3.33
r35 19 25 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=1.81 $Y=3.33
+ $X2=1.68 $Y2=3.33
r36 17 26 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=1.68 $Y2=3.33
r37 17 23 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r38 13 31 3.27398 $w=3.3e-07 $l=1.67183e-07 $layer=LI1_cond $X=1.975 $Y=3.245
+ $X2=2.105 $Y2=3.33
r39 13 15 26.3665 $w=3.28e-07 $l=7.55e-07 $layer=LI1_cond $X=1.975 $Y=3.245
+ $X2=1.975 $Y2=2.49
r40 9 12 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=0.385 $Y=2.19
+ $X2=0.385 $Y2=2.9
r41 7 28 3.22214 $w=3.3e-07 $l=1.46458e-07 $layer=LI1_cond $X=0.385 $Y=3.245
+ $X2=0.275 $Y2=3.33
r42 7 12 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=0.385 $Y=3.245
+ $X2=0.385 $Y2=2.9
r43 2 15 300 $w=1.7e-07 $l=5.10221e-07 $layer=licon1_PDIFF $count=2 $X=1.835
+ $Y=2.045 $X2=1.975 $Y2=2.49
r44 1 12 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.24
+ $Y=2.045 $X2=0.385 $Y2=2.9
r45 1 9 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.24
+ $Y=2.045 $X2=0.385 $Y2=2.19
.ends

.subckt PM_SKY130_FD_SC_LP__O21AI_LP%Y 1 2 7 10 14 16 17
r31 20 22 3.82169 $w=4.15e-07 $l=1.3e-07 $layer=LI1_cond $X=1.327 $Y=2.06
+ $X2=1.327 $Y2=2.19
r32 17 28 3.6747 $w=4.15e-07 $l=1.25e-07 $layer=LI1_cond $X=1.327 $Y=2.775
+ $X2=1.327 $Y2=2.9
r33 16 17 10.8771 $w=4.15e-07 $l=3.7e-07 $layer=LI1_cond $X=1.327 $Y=2.405
+ $X2=1.327 $Y2=2.775
r34 16 22 6.32048 $w=4.15e-07 $l=2.15e-07 $layer=LI1_cond $X=1.327 $Y=2.405
+ $X2=1.327 $Y2=2.19
r35 12 14 4.81032 $w=4.58e-07 $l=1.85e-07 $layer=LI1_cond $X=1.995 $Y=0.495
+ $X2=2.18 $Y2=0.495
r36 9 14 6.6364 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=2.18 $Y=0.725 $X2=2.18
+ $Y2=0.495
r37 9 10 81.5508 $w=1.68e-07 $l=1.25e-06 $layer=LI1_cond $X=2.18 $Y=0.725
+ $X2=2.18 $Y2=1.975
r38 8 20 6.00275 $w=1.7e-07 $l=2.43e-07 $layer=LI1_cond $X=1.57 $Y=2.06
+ $X2=1.327 $Y2=2.06
r39 7 10 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.095 $Y=2.06
+ $X2=2.18 $Y2=1.975
r40 7 8 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=2.095 $Y=2.06
+ $X2=1.57 $Y2=2.06
r41 2 28 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=1.265
+ $Y=2.045 $X2=1.405 $Y2=2.9
r42 2 22 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.265
+ $Y=2.045 $X2=1.405 $Y2=2.19
r43 1 12 182 $w=1.7e-07 $l=3.07571e-07 $layer=licon1_NDIFF $count=1 $X=1.775
+ $Y=0.285 $X2=1.995 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__O21AI_LP%A_64_57# 1 2 9 11 12 15
r32 13 15 9.7783 $w=3.28e-07 $l=2.8e-07 $layer=LI1_cond $X=1.485 $Y=0.775
+ $X2=1.485 $Y2=0.495
r33 11 13 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.32 $Y=0.86
+ $X2=1.485 $Y2=0.775
r34 11 12 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.32 $Y=0.86 $X2=0.63
+ $Y2=0.86
r35 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.465 $Y=0.775
+ $X2=0.63 $Y2=0.86
r36 7 9 9.7783 $w=3.28e-07 $l=2.8e-07 $layer=LI1_cond $X=0.465 $Y=0.775
+ $X2=0.465 $Y2=0.495
r37 2 15 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.345
+ $Y=0.285 $X2=1.485 $Y2=0.495
r38 1 9 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=0.32
+ $Y=0.285 $X2=0.465 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_LP__O21AI_LP%VGND 1 6 9 10 11 21 22
r23 21 22 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r24 18 21 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r25 14 15 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r26 11 22 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r27 11 15 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r28 11 18 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r29 9 14 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=0.81 $Y=0 $X2=0.72
+ $Y2=0
r30 9 10 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.81 $Y=0 $X2=0.975
+ $Y2=0
r31 8 18 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=1.14 $Y=0 $X2=1.2 $Y2=0
r32 8 10 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.14 $Y=0 $X2=0.975
+ $Y2=0
r33 4 10 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.975 $Y=0.085
+ $X2=0.975 $Y2=0
r34 4 6 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=0.975 $Y=0.085
+ $X2=0.975 $Y2=0.43
r35 1 6 182 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_NDIFF $count=1 $X=0.755
+ $Y=0.285 $X2=0.975 $Y2=0.43
.ends

