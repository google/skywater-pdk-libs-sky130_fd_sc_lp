* File: sky130_fd_sc_lp__o211a_0.pex.spice
* Created: Wed Sep  2 10:13:37 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O211A_0%A_80_21# 1 2 3 12 14 15 16 18 20 25 29 31 34
+ 35 37 39 40 42 45 47 48 49
c103 40 0 1.65825e-19 $X=2.745 $Y=1.275
c104 37 0 1.99675e-19 $X=3.1 $Y=0.445
c105 34 0 1.01278e-19 $X=2.66 $Y=1.19
c106 25 0 3.08377e-20 $X=2.065 $Y=2.142
r107 43 49 3.11846 $w=3.3e-07 $l=9.3e-08 $layer=LI1_cond $X=3.1 $Y=2.235 $X2=3.1
+ $Y2=2.142
r108 43 45 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=3.1 $Y=2.235
+ $X2=3.1 $Y2=2.57
r109 42 49 3.11846 $w=3.3e-07 $l=9.2e-08 $layer=LI1_cond $X=3.1 $Y=2.05 $X2=3.1
+ $Y2=2.142
r110 41 42 24.0965 $w=3.28e-07 $l=6.9e-07 $layer=LI1_cond $X=3.1 $Y=1.36 $X2=3.1
+ $Y2=2.05
r111 39 41 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.935 $Y=1.275
+ $X2=3.1 $Y2=1.36
r112 39 40 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=2.935 $Y=1.275
+ $X2=2.745 $Y2=1.275
r113 35 37 12.5882 $w=3.23e-07 $l=3.55e-07 $layer=LI1_cond $X=2.745 $Y=0.442
+ $X2=3.1 $Y2=0.442
r114 34 40 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.66 $Y=1.19
+ $X2=2.745 $Y2=1.275
r115 33 35 7.72402 $w=3.25e-07 $l=2.01057e-07 $layer=LI1_cond $X=2.66 $Y=0.605
+ $X2=2.745 $Y2=0.442
r116 33 34 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=2.66 $Y=0.605
+ $X2=2.66 $Y2=1.19
r117 32 48 6.98765 $w=1.85e-07 $l=1.35e-07 $layer=LI1_cond $X=2.335 $Y=2.142
+ $X2=2.2 $Y2=2.142
r118 31 49 3.48878 $w=1.85e-07 $l=1.65e-07 $layer=LI1_cond $X=2.935 $Y=2.142
+ $X2=3.1 $Y2=2.142
r119 31 32 35.9705 $w=1.83e-07 $l=6e-07 $layer=LI1_cond $X=2.935 $Y=2.142
+ $X2=2.335 $Y2=2.142
r120 27 48 0.0237744 $w=2.7e-07 $l=9.3e-08 $layer=LI1_cond $X=2.2 $Y=2.235
+ $X2=2.2 $Y2=2.142
r121 27 29 13.4452 $w=2.68e-07 $l=3.15e-07 $layer=LI1_cond $X=2.2 $Y=2.235
+ $X2=2.2 $Y2=2.55
r122 25 48 6.98765 $w=1.85e-07 $l=1.35e-07 $layer=LI1_cond $X=2.065 $Y=2.142
+ $X2=2.2 $Y2=2.142
r123 25 47 16.4865 $w=1.83e-07 $l=2.75e-07 $layer=LI1_cond $X=2.065 $Y=2.142
+ $X2=1.79 $Y2=2.142
r124 22 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.05
+ $Y=2.1 $X2=1.05 $Y2=2.1
r125 20 47 7.4448 $w=2.98e-07 $l=1.5e-07 $layer=LI1_cond $X=1.64 $Y=2.085
+ $X2=1.79 $Y2=2.085
r126 20 22 22.6647 $w=2.98e-07 $l=5.9e-07 $layer=LI1_cond $X=1.64 $Y=2.085
+ $X2=1.05 $Y2=2.085
r127 16 23 21.5735 $w=1.5e-07 $l=1.70895e-07 $layer=POLY_cond $X=1.115 $Y=2.265
+ $X2=1.127 $Y2=2.1
r128 16 18 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.115 $Y=2.265
+ $X2=1.115 $Y2=2.745
r129 14 23 10.6039 $w=3.3e-07 $l=8.7e-08 $layer=POLY_cond $X=1.04 $Y=2.1
+ $X2=1.127 $Y2=2.1
r130 14 15 85.682 $w=3.3e-07 $l=4.9e-07 $layer=POLY_cond $X=1.04 $Y=2.1 $X2=0.55
+ $Y2=2.1
r131 10 15 32.1775 $w=3.3e-07 $l=1.98997e-07 $layer=POLY_cond $X=0.475 $Y=1.935
+ $X2=0.55 $Y2=2.1
r132 10 12 764.021 $w=1.5e-07 $l=1.49e-06 $layer=POLY_cond $X=0.475 $Y=1.935
+ $X2=0.475 $Y2=0.445
r133 3 45 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=2.96
+ $Y=2.425 $X2=3.1 $Y2=2.57
r134 2 29 300 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=2 $X=2.06
+ $Y=2.425 $X2=2.2 $Y2=2.55
r135 1 37 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.96
+ $Y=0.235 $X2=3.1 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__O211A_0%A1 3 7 9 10 11 15
c39 7 0 1.7152e-19 $X=1.625 $Y=2.745
r40 14 15 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.535
+ $Y=1.4 $X2=1.535 $Y2=1.4
r41 11 15 8.67569 $w=4.43e-07 $l=3.35e-07 $layer=LI1_cond $X=1.2 $Y=1.342
+ $X2=1.535 $Y2=1.342
r42 9 14 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=1.55 $Y=1.4 $X2=1.535
+ $Y2=1.4
r43 9 10 5.03009 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=1.55 $Y=1.4 $X2=1.625
+ $Y2=1.4
r44 5 10 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.625 $Y=1.565
+ $X2=1.625 $Y2=1.4
r45 5 7 605.064 $w=1.5e-07 $l=1.18e-06 $layer=POLY_cond $X=1.625 $Y=1.565
+ $X2=1.625 $Y2=2.745
r46 1 10 37.0704 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.625 $Y=1.235
+ $X2=1.625 $Y2=1.4
r47 1 3 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.625 $Y=1.235
+ $X2=1.625 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__O211A_0%A2 3 7 11 12 13 14 18
c47 18 0 1.90167e-19 $X=2.075 $Y=1.33
c48 12 0 3.08377e-20 $X=2.075 $Y=1.835
c49 3 0 1.41676e-19 $X=1.985 $Y=2.745
r50 13 14 13.3251 $w=3.18e-07 $l=3.7e-07 $layer=LI1_cond $X=2.12 $Y=1.295
+ $X2=2.12 $Y2=1.665
r51 13 18 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.075
+ $Y=1.33 $X2=2.075 $Y2=1.33
r52 11 18 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.075 $Y=1.67
+ $X2=2.075 $Y2=1.33
r53 11 12 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.075 $Y=1.67
+ $X2=2.075 $Y2=1.835
r54 10 18 38.0424 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.075 $Y=1.165
+ $X2=2.075 $Y2=1.33
r55 7 10 369.191 $w=1.5e-07 $l=7.2e-07 $layer=POLY_cond $X=2.065 $Y=0.445
+ $X2=2.065 $Y2=1.165
r56 3 12 466.617 $w=1.5e-07 $l=9.1e-07 $layer=POLY_cond $X=1.985 $Y=2.745
+ $X2=1.985 $Y2=1.835
.ends

.subckt PM_SKY130_FD_SC_LP__O211A_0%B1 3 7 11 12 13 16
c52 13 0 1.41676e-19 $X=2.64 $Y=1.665
c53 7 0 1.98559e-19 $X=2.525 $Y=0.445
r54 16 19 46.536 $w=4.35e-07 $l=1.65e-07 $layer=POLY_cond $X=2.667 $Y=1.695
+ $X2=2.667 $Y2=1.86
r55 16 18 50.3716 $w=4.35e-07 $l=1.95e-07 $layer=POLY_cond $X=2.667 $Y=1.695
+ $X2=2.667 $Y2=1.5
r56 13 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.615
+ $Y=1.695 $X2=2.615 $Y2=1.695
r57 11 12 43.7534 $w=2.2e-07 $l=1.5e-07 $layer=POLY_cond $X=2.49 $Y=2.075
+ $X2=2.49 $Y2=2.225
r58 11 19 110.245 $w=1.5e-07 $l=2.15e-07 $layer=POLY_cond $X=2.525 $Y=2.075
+ $X2=2.525 $Y2=1.86
r59 7 18 540.968 $w=1.5e-07 $l=1.055e-06 $layer=POLY_cond $X=2.525 $Y=0.445
+ $X2=2.525 $Y2=1.5
r60 3 12 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=2.455 $Y=2.745
+ $X2=2.455 $Y2=2.225
.ends

.subckt PM_SKY130_FD_SC_LP__O211A_0%C1 1 3 6 9 12 14 21
c37 14 0 1.98559e-19 $X=3.12 $Y=0.925
c38 9 0 7.69365e-20 $X=3.17 $Y=2.07
r39 19 21 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=3.08 $Y=0.93 $X2=3.17
+ $Y2=0.93
r40 16 19 34.0979 $w=3.3e-07 $l=1.95e-07 $layer=POLY_cond $X=2.885 $Y=0.93
+ $X2=3.08 $Y2=0.93
r41 14 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.08
+ $Y=0.93 $X2=3.08 $Y2=0.93
r42 10 12 146.138 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.885 $Y=2.145
+ $X2=3.17 $Y2=2.145
r43 9 12 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.17 $Y=2.07 $X2=3.17
+ $Y2=2.145
r44 8 21 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.17 $Y=1.095
+ $X2=3.17 $Y2=0.93
r45 8 9 499.947 $w=1.5e-07 $l=9.75e-07 $layer=POLY_cond $X=3.17 $Y=1.095
+ $X2=3.17 $Y2=2.07
r46 4 10 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.885 $Y=2.22
+ $X2=2.885 $Y2=2.145
r47 4 6 269.202 $w=1.5e-07 $l=5.25e-07 $layer=POLY_cond $X=2.885 $Y=2.22
+ $X2=2.885 $Y2=2.745
r48 1 16 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.885 $Y=0.765
+ $X2=2.885 $Y2=0.93
r49 1 3 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.885 $Y=0.765
+ $X2=2.885 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__O211A_0%X 1 2 9 11 12 13 14 15 16 28
c19 9 0 1.7152e-19 $X=0.9 $Y=2.57
r20 15 16 13.4589 $w=2.78e-07 $l=3.27e-07 $layer=LI1_cond $X=0.225 $Y=2.035
+ $X2=0.225 $Y2=2.362
r21 14 15 15.2287 $w=2.78e-07 $l=3.7e-07 $layer=LI1_cond $X=0.225 $Y=1.665
+ $X2=0.225 $Y2=2.035
r22 13 14 15.2287 $w=2.78e-07 $l=3.7e-07 $layer=LI1_cond $X=0.225 $Y=1.295
+ $X2=0.225 $Y2=1.665
r23 12 13 15.2287 $w=2.78e-07 $l=3.7e-07 $layer=LI1_cond $X=0.225 $Y=0.925
+ $X2=0.225 $Y2=1.295
r24 11 12 15.2287 $w=2.78e-07 $l=3.7e-07 $layer=LI1_cond $X=0.225 $Y=0.555
+ $X2=0.225 $Y2=0.925
r25 11 28 4.52745 $w=2.78e-07 $l=1.1e-07 $layer=LI1_cond $X=0.225 $Y=0.555
+ $X2=0.225 $Y2=0.445
r26 7 16 2.48464 $w=6.7e-07 $l=1.4e-07 $layer=LI1_cond $X=0.365 $Y=2.74
+ $X2=0.225 $Y2=2.74
r27 7 9 9.55078 $w=6.68e-07 $l=5.35e-07 $layer=LI1_cond $X=0.365 $Y=2.74 $X2=0.9
+ $Y2=2.74
r28 2 9 150 $w=1.7e-07 $l=5.32588e-07 $layer=licon1_PDIFF $count=4 $X=0.435
+ $Y=2.425 $X2=0.9 $Y2=2.57
r29 1 28 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__O211A_0%VPWR 1 2 9 13 16 17 18 27 33 34 37
r40 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r41 34 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.64 $Y2=3.33
r42 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r43 31 37 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.765 $Y=3.33
+ $X2=2.635 $Y2=3.33
r44 31 33 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=2.765 $Y=3.33
+ $X2=3.12 $Y2=3.33
r45 30 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=2.64 $Y2=3.33
r46 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r47 27 37 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.505 $Y=3.33
+ $X2=2.635 $Y2=3.33
r48 27 29 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=2.505 $Y=3.33
+ $X2=2.16 $Y2=3.33
r49 25 26 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r50 22 26 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.2 $Y2=3.33
r51 21 25 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.24 $Y=3.33 $X2=1.2
+ $Y2=3.33
r52 21 22 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r53 18 30 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r54 18 26 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r55 16 25 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=1.245 $Y=3.33
+ $X2=1.2 $Y2=3.33
r56 16 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.245 $Y=3.33
+ $X2=1.41 $Y2=3.33
r57 15 29 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=1.575 $Y=3.33
+ $X2=2.16 $Y2=3.33
r58 15 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.575 $Y=3.33
+ $X2=1.41 $Y2=3.33
r59 11 37 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=2.635 $Y=3.245
+ $X2=2.635 $Y2=3.33
r60 11 13 29.9192 $w=2.58e-07 $l=6.75e-07 $layer=LI1_cond $X=2.635 $Y=3.245
+ $X2=2.635 $Y2=2.57
r61 7 17 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.41 $Y=3.245 $X2=1.41
+ $Y2=3.33
r62 7 9 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=1.41 $Y=3.245
+ $X2=1.41 $Y2=2.57
r63 2 13 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=2.53
+ $Y=2.425 $X2=2.67 $Y2=2.57
r64 1 9 300 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_PDIFF $count=2 $X=1.19
+ $Y=2.425 $X2=1.41 $Y2=2.57
.ends

.subckt PM_SKY130_FD_SC_LP__O211A_0%VGND 1 2 9 13 16 17 18 20 33 34 37
r41 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r42 33 34 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r43 31 34 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r44 30 33 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r45 30 31 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r46 25 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.875 $Y=0 $X2=0.71
+ $Y2=0
r47 25 27 52.5187 $w=1.68e-07 $l=8.05e-07 $layer=LI1_cond $X=0.875 $Y=0 $X2=1.68
+ $Y2=0
r48 23 38 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r49 22 23 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r50 20 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.545 $Y=0 $X2=0.71
+ $Y2=0
r51 20 22 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.545 $Y=0 $X2=0.24
+ $Y2=0
r52 18 31 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.16
+ $Y2=0
r53 18 38 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=0.72
+ $Y2=0
r54 18 27 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r55 16 27 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=1.745 $Y=0 $X2=1.68
+ $Y2=0
r56 16 17 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.745 $Y=0 $X2=1.875
+ $Y2=0
r57 15 30 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=2.005 $Y=0 $X2=2.16
+ $Y2=0
r58 15 17 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.005 $Y=0 $X2=1.875
+ $Y2=0
r59 11 17 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=1.875 $Y=0.085
+ $X2=1.875 $Y2=0
r60 11 13 15.9569 $w=2.58e-07 $l=3.6e-07 $layer=LI1_cond $X=1.875 $Y=0.085
+ $X2=1.875 $Y2=0.445
r61 7 37 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.71 $Y=0.085 $X2=0.71
+ $Y2=0
r62 7 9 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=0.71 $Y=0.085 $X2=0.71
+ $Y2=0.445
r63 2 13 182 $w=1.7e-07 $l=2.74955e-07 $layer=licon1_NDIFF $count=1 $X=1.7
+ $Y=0.235 $X2=1.85 $Y2=0.445
r64 1 9 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.235 $X2=0.69 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__O211A_0%A_257_47# 1 2 9 11 12 15
r28 13 15 16.7856 $w=2.28e-07 $l=3.35e-07 $layer=LI1_cond $X=2.29 $Y=0.78
+ $X2=2.29 $Y2=0.445
r29 11 13 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=2.175 $Y=0.865
+ $X2=2.29 $Y2=0.78
r30 11 12 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=2.175 $Y=0.865
+ $X2=1.575 $Y2=0.865
r31 7 12 7.68211 $w=1.7e-07 $l=1.9799e-07 $layer=LI1_cond $X=1.415 $Y=0.78
+ $X2=1.575 $Y2=0.865
r32 7 9 12.0646 $w=3.18e-07 $l=3.35e-07 $layer=LI1_cond $X=1.415 $Y=0.78
+ $X2=1.415 $Y2=0.445
r33 2 15 182 $w=1.7e-07 $l=2.82489e-07 $layer=licon1_NDIFF $count=1 $X=2.14
+ $Y=0.235 $X2=2.31 $Y2=0.445
r34 1 9 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=1.285
+ $Y=0.235 $X2=1.41 $Y2=0.445
.ends

