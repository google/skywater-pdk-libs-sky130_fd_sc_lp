* File: sky130_fd_sc_lp__and4_0.spice
* Created: Wed Sep  2 09:32:39 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__and4_0.pex.spice"
.subckt sky130_fd_sc_lp__and4_0  VNB VPB A B C D VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* D	D
* C	C
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1002 A_167_58# N_A_M1002_g N_A_84_58#_M1002_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1113 PD=0.63 PS=1.37 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002 A=0.063 P=1.14 MULT=1
MM1003 A_239_58# N_B_M1003_g A_167_58# VNB NSHORT L=0.15 W=0.42 AD=0.0441
+ AS=0.0441 PD=0.63 PS=0.63 NRD=14.28 NRS=14.28 M=1 R=2.8 SA=75000.6 SB=75001.7
+ A=0.063 P=1.14 MULT=1
MM1006 A_311_58# N_C_M1006_g A_239_58# VNB NSHORT L=0.15 W=0.42 AD=0.0441
+ AS=0.0441 PD=0.63 PS=0.63 NRD=14.28 NRS=14.28 M=1 R=2.8 SA=75000.9 SB=75001.3
+ A=0.063 P=1.14 MULT=1
MM1008 N_VGND_M1008_d N_D_M1008_g A_311_58# VNB NSHORT L=0.15 W=0.42 AD=0.1302
+ AS=0.0441 PD=1.04 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.3 SB=75001
+ A=0.063 P=1.14 MULT=1
MM1005 N_X_M1005_d N_A_84_58#_M1005_g N_VGND_M1008_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.1302 PD=1.37 PS=1.04 NRD=0 NRS=0 M=1 R=2.8 SA=75002 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1009 N_A_84_58#_M1009_d N_A_M1009_g N_VPWR_M1009_s VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2 SB=75002.4
+ A=0.063 P=1.14 MULT=1
MM1000 N_VPWR_M1000_d N_B_M1000_g N_A_84_58#_M1009_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0693 AS=0.0588 PD=0.75 PS=0.7 NRD=7.0329 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75001.9 A=0.063 P=1.14 MULT=1
MM1007 N_A_84_58#_M1007_d N_C_M1007_g N_VPWR_M1000_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0588 AS=0.0693 PD=0.7 PS=0.75 NRD=0 NRS=16.4101 M=1 R=2.8 SA=75001.1
+ SB=75001.5 A=0.063 P=1.14 MULT=1
MM1004 N_VPWR_M1004_d N_D_M1004_g N_A_84_58#_M1007_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.137094 AS=0.0588 PD=1.05 PS=0.7 NRD=127.301 NRS=0 M=1 R=2.8 SA=75001.5
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1001 N_X_M1001_d N_A_84_58#_M1001_g N_VPWR_M1004_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1696 AS=0.208906 PD=1.81 PS=1.6 NRD=0 NRS=0 M=1 R=4.26667 SA=75001.6
+ SB=75000.2 A=0.096 P=1.58 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9751 P=11.21
*
.include "sky130_fd_sc_lp__and4_0.pxi.spice"
*
.ends
*
*
