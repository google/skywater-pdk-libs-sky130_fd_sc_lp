* File: sky130_fd_sc_lp__a21o_4.pex.spice
* Created: Fri Aug 28 09:51:10 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A21O_4%A_134_269# 1 2 3 12 16 20 24 28 32 36 40 42
+ 49 51 52 53 56 60 64 67 68 69 71
c138 69 0 4.75122e-20 $X=3.215 $Y=0.95
c139 42 0 1.58172e-19 $X=2.205 $Y=1.512
r140 83 84 20.9834 $w=3.3e-07 $l=1.2e-07 $layer=POLY_cond $X=2.035 $Y=1.51
+ $X2=2.155 $Y2=1.51
r141 82 83 54.207 $w=3.3e-07 $l=3.1e-07 $layer=POLY_cond $X=1.725 $Y=1.51
+ $X2=2.035 $Y2=1.51
r142 81 82 20.9834 $w=3.3e-07 $l=1.2e-07 $layer=POLY_cond $X=1.605 $Y=1.51
+ $X2=1.725 $Y2=1.51
r143 80 81 54.207 $w=3.3e-07 $l=3.1e-07 $layer=POLY_cond $X=1.295 $Y=1.51
+ $X2=1.605 $Y2=1.51
r144 79 80 20.9834 $w=3.3e-07 $l=1.2e-07 $layer=POLY_cond $X=1.175 $Y=1.51
+ $X2=1.295 $Y2=1.51
r145 75 77 20.9834 $w=3.3e-07 $l=1.2e-07 $layer=POLY_cond $X=0.745 $Y=1.51
+ $X2=0.865 $Y2=1.51
r146 71 73 9.16716 $w=2.18e-07 $l=1.75e-07 $layer=LI1_cond $X=4.515 $Y=0.77
+ $X2=4.515 $Y2=0.945
r147 67 68 2.64593 $w=3.28e-07 $l=6e-08 $layer=LI1_cond $X=3.2 $Y=1.97 $X2=3.2
+ $Y2=1.91
r148 65 69 4.30018 $w=1.7e-07 $l=1.5248e-07 $layer=LI1_cond $X=3.365 $Y=0.945
+ $X2=3.215 $Y2=0.95
r149 64 73 2.2496 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=4.405 $Y=0.945
+ $X2=4.515 $Y2=0.945
r150 64 65 67.8503 $w=1.68e-07 $l=1.04e-06 $layer=LI1_cond $X=4.405 $Y=0.945
+ $X2=3.365 $Y2=0.945
r151 62 69 1.96316 $w=2.6e-07 $l=9.94987e-08 $layer=LI1_cond $X=3.235 $Y=1.04
+ $X2=3.215 $Y2=0.95
r152 62 68 38.5625 $w=2.58e-07 $l=8.7e-07 $layer=LI1_cond $X=3.235 $Y=1.04
+ $X2=3.235 $Y2=1.91
r153 58 69 1.96316 $w=2.4e-07 $l=1.03923e-07 $layer=LI1_cond $X=3.185 $Y=0.86
+ $X2=3.215 $Y2=0.95
r154 58 60 21.1281 $w=2.38e-07 $l=4.4e-07 $layer=LI1_cond $X=3.185 $Y=0.86
+ $X2=3.185 $Y2=0.42
r155 54 67 3.66686 $w=3.28e-07 $l=1.05e-07 $layer=LI1_cond $X=3.2 $Y=2.075
+ $X2=3.2 $Y2=1.97
r156 54 56 20.0804 $w=3.28e-07 $l=5.75e-07 $layer=LI1_cond $X=3.2 $Y=2.075
+ $X2=3.2 $Y2=2.65
r157 52 69 4.30018 $w=1.7e-07 $l=1.5248e-07 $layer=LI1_cond $X=3.065 $Y=0.955
+ $X2=3.215 $Y2=0.95
r158 52 53 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.065 $Y=0.955
+ $X2=2.375 $Y2=0.955
r159 50 53 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.29 $Y=1.04
+ $X2=2.375 $Y2=0.955
r160 50 51 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=2.29 $Y=1.04
+ $X2=2.29 $Y2=1.415
r161 49 84 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=2.17 $Y=1.51
+ $X2=2.155 $Y2=1.51
r162 48 49 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.17
+ $Y=1.51 $X2=2.17 $Y2=1.51
r163 45 79 4.37153 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=1.15 $Y=1.51
+ $X2=1.175 $Y2=1.51
r164 45 77 49.8355 $w=3.3e-07 $l=2.85e-07 $layer=POLY_cond $X=1.15 $Y=1.51
+ $X2=0.865 $Y2=1.51
r165 44 48 58.014 $w=1.93e-07 $l=1.02e-06 $layer=LI1_cond $X=1.15 $Y=1.512
+ $X2=2.17 $Y2=1.512
r166 44 45 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.15
+ $Y=1.51 $X2=1.15 $Y2=1.51
r167 42 51 6.85817 $w=1.95e-07 $l=1.32868e-07 $layer=LI1_cond $X=2.205 $Y=1.512
+ $X2=2.29 $Y2=1.415
r168 42 48 1.99068 $w=1.93e-07 $l=3.5e-08 $layer=LI1_cond $X=2.205 $Y=1.512
+ $X2=2.17 $Y2=1.512
r169 38 84 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.155 $Y=1.345
+ $X2=2.155 $Y2=1.51
r170 38 40 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=2.155 $Y=1.345
+ $X2=2.155 $Y2=0.665
r171 34 83 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.035 $Y=1.675
+ $X2=2.035 $Y2=1.51
r172 34 36 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.035 $Y=1.675
+ $X2=2.035 $Y2=2.465
r173 30 82 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.725 $Y=1.345
+ $X2=1.725 $Y2=1.51
r174 30 32 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=1.725 $Y=1.345
+ $X2=1.725 $Y2=0.665
r175 26 81 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.605 $Y=1.675
+ $X2=1.605 $Y2=1.51
r176 26 28 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.605 $Y=1.675
+ $X2=1.605 $Y2=2.465
r177 22 80 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.295 $Y=1.345
+ $X2=1.295 $Y2=1.51
r178 22 24 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=1.295 $Y=1.345
+ $X2=1.295 $Y2=0.665
r179 18 79 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.175 $Y=1.675
+ $X2=1.175 $Y2=1.51
r180 18 20 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=1.175 $Y=1.675
+ $X2=1.175 $Y2=2.465
r181 14 77 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.865 $Y=1.345
+ $X2=0.865 $Y2=1.51
r182 14 16 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=0.865 $Y=1.345
+ $X2=0.865 $Y2=0.665
r183 10 75 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.745 $Y=1.675
+ $X2=0.745 $Y2=1.51
r184 10 12 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=0.745 $Y=1.675
+ $X2=0.745 $Y2=2.465
r185 3 67 400 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_PDIFF $count=1 $X=3.06
+ $Y=1.835 $X2=3.2 $Y2=1.97
r186 3 56 400 $w=1.7e-07 $l=8.82227e-07 $layer=licon1_PDIFF $count=1 $X=3.06
+ $Y=1.835 $X2=3.2 $Y2=2.65
r187 2 71 182 $w=1.7e-07 $l=5.90868e-07 $layer=licon1_NDIFF $count=1 $X=4.39
+ $Y=0.245 $X2=4.53 $Y2=0.77
r188 1 60 91 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=2 $X=3.06
+ $Y=0.245 $X2=3.2 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__A21O_4%B1 3 6 8 10 12 15 17 18 19 22 23
c62 6 0 1.58172e-19 $X=2.985 $Y=2.465
r63 25 27 45.1558 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=2.872 $Y=1.375
+ $X2=2.872 $Y2=1.54
r64 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.85
+ $Y=1.375 $X2=2.85 $Y2=1.375
r65 22 25 13.3477 $w=3.75e-07 $l=9e-08 $layer=POLY_cond $X=2.872 $Y=1.285
+ $X2=2.872 $Y2=1.375
r66 22 23 31.8081 $w=3.75e-07 $l=7.5e-08 $layer=POLY_cond $X=2.872 $Y=1.285
+ $X2=2.872 $Y2=1.21
r67 19 26 8.79496 $w=3.78e-07 $l=2.9e-07 $layer=LI1_cond $X=2.745 $Y=1.665
+ $X2=2.745 $Y2=1.375
r68 18 26 2.4262 $w=3.78e-07 $l=8e-08 $layer=LI1_cond $X=2.745 $Y=1.295
+ $X2=2.745 $Y2=1.375
r69 13 17 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.415 $Y=1.36
+ $X2=3.415 $Y2=1.285
r70 13 15 566.606 $w=1.5e-07 $l=1.105e-06 $layer=POLY_cond $X=3.415 $Y=1.36
+ $X2=3.415 $Y2=2.465
r71 10 17 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.415 $Y=1.21
+ $X2=3.415 $Y2=1.285
r72 10 12 175.127 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=3.415 $Y=1.21
+ $X2=3.415 $Y2=0.665
r73 9 22 24.2915 $w=1.5e-07 $l=1.88e-07 $layer=POLY_cond $X=3.06 $Y=1.285
+ $X2=2.872 $Y2=1.285
r74 8 17 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.34 $Y=1.285
+ $X2=3.415 $Y2=1.285
r75 8 9 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=3.34 $Y=1.285 $X2=3.06
+ $Y2=1.285
r76 6 27 474.309 $w=1.5e-07 $l=9.25e-07 $layer=POLY_cond $X=2.985 $Y=2.465
+ $X2=2.985 $Y2=1.54
r77 3 23 175.127 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=2.985 $Y=0.665
+ $X2=2.985 $Y2=1.21
.ends

.subckt PM_SKY130_FD_SC_LP__A21O_4%A2 3 7 11 15 19 21 28 29 31 32 33
c83 29 0 1.46692e-19 $X=5.265 $Y=1.51
c84 7 0 4.75122e-20 $X=3.885 $Y=0.665
c85 3 0 1.19057e-19 $X=3.845 $Y=2.465
r86 32 33 16.2679 $w=3.38e-07 $l=3.95e-07 $layer=LI1_cond $X=4.56 $Y=2.035
+ $X2=4.955 $Y2=2.035
r87 31 48 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4 $Y=2.035 $X2=4.085
+ $Y2=2.035
r88 31 32 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=4.125 $Y=2.035
+ $X2=4.56 $Y2=2.035
r89 31 48 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=4.125 $Y=2.035
+ $X2=4.085 $Y2=2.035
r90 29 46 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.265 $Y=1.51
+ $X2=5.265 $Y2=1.675
r91 29 45 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.265 $Y=1.51
+ $X2=5.265 $Y2=1.345
r92 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.265
+ $Y=1.51 $X2=5.265 $Y2=1.51
r93 25 33 11.7777 $w=3.38e-07 $l=3.05e-07 $layer=LI1_cond $X=5.04 $Y=1.645
+ $X2=5.04 $Y2=1.95
r94 24 28 8.64332 $w=2.98e-07 $l=2.25e-07 $layer=LI1_cond $X=5.04 $Y=1.495
+ $X2=5.265 $Y2=1.495
r95 24 25 4.061 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=5.04 $Y=1.495 $X2=5.04
+ $Y2=1.645
r96 22 31 15.6476 $w=2.58e-07 $l=3.25e-07 $layer=LI1_cond $X=4 $Y=1.625 $X2=4
+ $Y2=1.95
r97 21 22 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4 $Y=1.46 $X2=4
+ $Y2=1.625
r98 19 43 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.865 $Y=1.46
+ $X2=3.865 $Y2=1.625
r99 19 42 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.865 $Y=1.46
+ $X2=3.865 $Y2=1.295
r100 18 21 4.71454 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=3.865 $Y=1.46
+ $X2=4 $Y2=1.46
r101 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.865
+ $Y=1.46 $X2=3.865 $Y2=1.46
r102 15 46 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=5.175 $Y=2.465
+ $X2=5.175 $Y2=1.675
r103 11 45 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=5.175 $Y=0.665
+ $X2=5.175 $Y2=1.345
r104 7 42 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=3.885 $Y=0.665
+ $X2=3.885 $Y2=1.295
r105 3 43 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=3.845 $Y=2.465
+ $X2=3.845 $Y2=1.625
.ends

.subckt PM_SKY130_FD_SC_LP__A21O_4%A1 1 3 6 8 10 13 15 16 24
c51 15 0 2.65748e-19 $X=4.56 $Y=1.295
r52 22 24 55.0813 $w=3.3e-07 $l=3.15e-07 $layer=POLY_cond $X=4.43 $Y=1.36
+ $X2=4.745 $Y2=1.36
r53 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.43
+ $Y=1.36 $X2=4.43 $Y2=1.36
r54 19 22 20.109 $w=3.3e-07 $l=1.15e-07 $layer=POLY_cond $X=4.315 $Y=1.36
+ $X2=4.43 $Y2=1.36
r55 16 23 9.24987 $w=3.78e-07 $l=3.05e-07 $layer=LI1_cond $X=4.455 $Y=1.665
+ $X2=4.455 $Y2=1.36
r56 15 23 1.97128 $w=3.78e-07 $l=6.5e-08 $layer=LI1_cond $X=4.455 $Y=1.295
+ $X2=4.455 $Y2=1.36
r57 11 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.745 $Y=1.525
+ $X2=4.745 $Y2=1.36
r58 11 13 482 $w=1.5e-07 $l=9.4e-07 $layer=POLY_cond $X=4.745 $Y=1.525 $X2=4.745
+ $Y2=2.465
r59 8 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.745 $Y=1.195
+ $X2=4.745 $Y2=1.36
r60 8 10 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=4.745 $Y=1.195
+ $X2=4.745 $Y2=0.665
r61 4 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.315 $Y=1.525
+ $X2=4.315 $Y2=1.36
r62 4 6 482 $w=1.5e-07 $l=9.4e-07 $layer=POLY_cond $X=4.315 $Y=1.525 $X2=4.315
+ $Y2=2.465
r63 1 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.315 $Y=1.195
+ $X2=4.315 $Y2=1.36
r64 1 3 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=4.315 $Y=1.195
+ $X2=4.315 $Y2=0.665
.ends

.subckt PM_SKY130_FD_SC_LP__A21O_4%VPWR 1 2 3 4 5 18 24 28 32 38 42 45 46 47 48
+ 49 58 66 73 74 77 80 83
r93 83 84 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r94 80 81 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r95 77 78 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r96 74 84 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=5.04 $Y2=3.33
r97 73 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r98 71 83 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.125 $Y=3.33
+ $X2=4.96 $Y2=3.33
r99 71 73 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=5.125 $Y=3.33
+ $X2=5.52 $Y2=3.33
r100 70 84 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.04 $Y2=3.33
r101 70 81 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=4.08 $Y2=3.33
r102 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r103 67 80 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.245 $Y=3.33
+ $X2=4.08 $Y2=3.33
r104 67 69 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=4.245 $Y=3.33
+ $X2=4.56 $Y2=3.33
r105 66 83 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.795 $Y=3.33
+ $X2=4.96 $Y2=3.33
r106 66 69 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=4.795 $Y=3.33
+ $X2=4.56 $Y2=3.33
r107 65 81 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r108 64 65 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r109 62 78 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r110 61 64 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.64 $Y=3.33 $X2=3.6
+ $Y2=3.33
r111 61 62 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r112 59 77 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=2.385 $Y=3.33
+ $X2=2.235 $Y2=3.33
r113 59 61 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=2.385 $Y=3.33
+ $X2=2.64 $Y2=3.33
r114 58 80 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.915 $Y=3.33
+ $X2=4.08 $Y2=3.33
r115 58 64 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=3.915 $Y=3.33
+ $X2=3.6 $Y2=3.33
r116 57 78 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=2.16 $Y2=3.33
r117 56 57 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r118 53 57 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=1.2 $Y2=3.33
r119 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r120 49 65 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.88 $Y=3.33
+ $X2=3.6 $Y2=3.33
r121 49 62 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.88 $Y=3.33
+ $X2=2.64 $Y2=3.33
r122 47 56 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=1.225 $Y=3.33
+ $X2=1.2 $Y2=3.33
r123 47 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.225 $Y=3.33
+ $X2=1.39 $Y2=3.33
r124 45 52 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=0.365 $Y=3.33
+ $X2=0.24 $Y2=3.33
r125 45 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.365 $Y=3.33
+ $X2=0.53 $Y2=3.33
r126 44 56 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=0.695 $Y=3.33
+ $X2=1.2 $Y2=3.33
r127 44 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.695 $Y=3.33
+ $X2=0.53 $Y2=3.33
r128 40 83 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.96 $Y=3.245
+ $X2=4.96 $Y2=3.33
r129 40 42 15.3659 $w=3.28e-07 $l=4.4e-07 $layer=LI1_cond $X=4.96 $Y=3.245
+ $X2=4.96 $Y2=2.805
r130 36 80 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.08 $Y=3.245
+ $X2=4.08 $Y2=3.33
r131 36 38 15.3659 $w=3.28e-07 $l=4.4e-07 $layer=LI1_cond $X=4.08 $Y=3.245
+ $X2=4.08 $Y2=2.805
r132 32 35 37.2623 $w=2.98e-07 $l=9.7e-07 $layer=LI1_cond $X=2.235 $Y=1.98
+ $X2=2.235 $Y2=2.95
r133 30 77 0.597483 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.235 $Y=3.245
+ $X2=2.235 $Y2=3.33
r134 30 35 11.3324 $w=2.98e-07 $l=2.95e-07 $layer=LI1_cond $X=2.235 $Y=3.245
+ $X2=2.235 $Y2=2.95
r135 29 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.555 $Y=3.33
+ $X2=1.39 $Y2=3.33
r136 28 77 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=2.085 $Y=3.33
+ $X2=2.235 $Y2=3.33
r137 28 29 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=2.085 $Y=3.33
+ $X2=1.555 $Y2=3.33
r138 24 27 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=1.39 $Y=2.24
+ $X2=1.39 $Y2=2.95
r139 22 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.39 $Y=3.245
+ $X2=1.39 $Y2=3.33
r140 22 27 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.39 $Y=3.245
+ $X2=1.39 $Y2=2.95
r141 18 21 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=0.53 $Y=2.24
+ $X2=0.53 $Y2=2.95
r142 16 46 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.53 $Y=3.245
+ $X2=0.53 $Y2=3.33
r143 16 21 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.53 $Y=3.245
+ $X2=0.53 $Y2=2.95
r144 5 42 600 $w=1.7e-07 $l=1.03764e-06 $layer=licon1_PDIFF $count=1 $X=4.82
+ $Y=1.835 $X2=4.96 $Y2=2.805
r145 4 38 600 $w=1.7e-07 $l=1.04695e-06 $layer=licon1_PDIFF $count=1 $X=3.92
+ $Y=1.835 $X2=4.08 $Y2=2.805
r146 3 35 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=2.11
+ $Y=1.835 $X2=2.25 $Y2=2.95
r147 3 32 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.11
+ $Y=1.835 $X2=2.25 $Y2=1.98
r148 2 27 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=1.25
+ $Y=1.835 $X2=1.39 $Y2=2.95
r149 2 24 400 $w=1.7e-07 $l=4.69814e-07 $layer=licon1_PDIFF $count=1 $X=1.25
+ $Y=1.835 $X2=1.39 $Y2=2.24
r150 1 21 400 $w=1.7e-07 $l=1.17584e-06 $layer=licon1_PDIFF $count=1 $X=0.405
+ $Y=1.835 $X2=0.53 $Y2=2.95
r151 1 18 400 $w=1.7e-07 $l=4.63303e-07 $layer=licon1_PDIFF $count=1 $X=0.405
+ $Y=1.835 $X2=0.53 $Y2=2.24
.ends

.subckt PM_SKY130_FD_SC_LP__A21O_4%X 1 2 3 4 15 19 21 23 25 27 31 35 36 37 40 47
+ 49
r57 47 49 0.92006 $w=6.48e-07 $l=5e-08 $layer=LI1_cond $X=0.48 $Y=1.245 $X2=0.48
+ $Y2=1.295
r58 40 47 2.16256 $w=6.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.48 $Y=1.16 $X2=0.48
+ $Y2=1.245
r59 40 49 0.31282 $w=6.48e-07 $l=1.7e-08 $layer=LI1_cond $X=0.48 $Y=1.312
+ $X2=0.48 $Y2=1.295
r60 36 40 10.0944 $w=2.03e-07 $l=1.8e-07 $layer=LI1_cond $X=0.985 $Y=1.16
+ $X2=0.805 $Y2=1.16
r61 36 37 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=0.985 $Y=1.16
+ $X2=1.08 $Y2=1.16
r62 33 40 8.61176 $w=6.48e-07 $l=4.68e-07 $layer=LI1_cond $X=0.48 $Y=1.78
+ $X2=0.48 $Y2=1.312
r63 33 35 2.74833 $w=4.2e-07 $l=1.68449e-07 $layer=LI1_cond $X=0.48 $Y=1.78
+ $X2=0.605 $Y2=1.882
r64 29 31 38.2345 $w=1.88e-07 $l=6.55e-07 $layer=LI1_cond $X=1.94 $Y=1.075
+ $X2=1.94 $Y2=0.42
r65 25 39 3.55261 $w=1.9e-07 $l=1.03e-07 $layer=LI1_cond $X=1.82 $Y=1.985
+ $X2=1.82 $Y2=1.882
r66 25 27 53.9952 $w=1.88e-07 $l=9.25e-07 $layer=LI1_cond $X=1.82 $Y=1.985
+ $X2=1.82 $Y2=2.91
r67 24 37 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.175 $Y=1.16
+ $X2=1.08 $Y2=1.16
r68 23 29 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=1.845 $Y=1.16
+ $X2=1.94 $Y2=1.075
r69 23 24 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.845 $Y=1.16
+ $X2=1.175 $Y2=1.16
r70 22 35 4.01484 $w=2.05e-07 $l=4.5e-07 $layer=LI1_cond $X=1.055 $Y=1.882
+ $X2=0.605 $Y2=1.882
r71 21 39 3.27668 $w=2.05e-07 $l=9.5e-08 $layer=LI1_cond $X=1.725 $Y=1.882
+ $X2=1.82 $Y2=1.882
r72 21 22 36.2483 $w=2.03e-07 $l=6.7e-07 $layer=LI1_cond $X=1.725 $Y=1.882
+ $X2=1.055 $Y2=1.882
r73 17 37 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.08 $Y=1.075
+ $X2=1.08 $Y2=1.16
r74 17 19 38.2345 $w=1.88e-07 $l=6.55e-07 $layer=LI1_cond $X=1.08 $Y=1.075
+ $X2=1.08 $Y2=0.42
r75 13 35 2.74833 $w=4.2e-07 $l=4.03225e-07 $layer=LI1_cond $X=0.96 $Y=1.985
+ $X2=0.605 $Y2=1.882
r76 13 15 53.9952 $w=1.88e-07 $l=9.25e-07 $layer=LI1_cond $X=0.96 $Y=1.985
+ $X2=0.96 $Y2=2.91
r77 4 39 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.68
+ $Y=1.835 $X2=1.82 $Y2=1.98
r78 4 27 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=1.68
+ $Y=1.835 $X2=1.82 $Y2=2.91
r79 3 35 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.82
+ $Y=1.835 $X2=0.96 $Y2=1.98
r80 3 15 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=0.82
+ $Y=1.835 $X2=0.96 $Y2=2.91
r81 2 31 91 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=2 $X=1.8
+ $Y=0.245 $X2=1.94 $Y2=0.42
r82 1 19 91 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=2 $X=0.94
+ $Y=0.245 $X2=1.08 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__A21O_4%A_529_367# 1 2 3 4 13 15 17 21 25 29 33 40 42
+ 44
r54 31 44 4.50329 $w=2e-07 $l=8.5e-08 $layer=LI1_cond $X=5.395 $Y=2.3 $X2=5.395
+ $Y2=2.385
r55 31 33 17.7455 $w=1.98e-07 $l=3.2e-07 $layer=LI1_cond $X=5.395 $Y=2.3
+ $X2=5.395 $Y2=1.98
r56 30 42 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=4.625 $Y=2.385
+ $X2=4.52 $Y2=2.385
r57 29 44 1.93381 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=5.295 $Y=2.385
+ $X2=5.395 $Y2=2.385
r58 29 30 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.295 $Y=2.385
+ $X2=4.625 $Y2=2.385
r59 26 40 2.0246 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=3.745 $Y=2.385
+ $X2=3.64 $Y2=2.385
r60 25 42 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=4.415 $Y=2.385
+ $X2=4.52 $Y2=2.385
r61 25 26 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.415 $Y=2.385
+ $X2=3.745 $Y2=2.385
r62 23 40 4.40882 $w=2.05e-07 $l=8.74643e-08 $layer=LI1_cond $X=3.635 $Y=2.47
+ $X2=3.64 $Y2=2.385
r63 23 24 24.1227 $w=1.98e-07 $l=4.35e-07 $layer=LI1_cond $X=3.635 $Y=2.47
+ $X2=3.635 $Y2=2.905
r64 19 40 4.40882 $w=2.05e-07 $l=8.5e-08 $layer=LI1_cond $X=3.64 $Y=2.3 $X2=3.64
+ $Y2=2.385
r65 19 21 16.9004 $w=2.08e-07 $l=3.2e-07 $layer=LI1_cond $X=3.64 $Y=2.3 $X2=3.64
+ $Y2=1.98
r66 18 38 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.865 $Y=2.99
+ $X2=2.735 $Y2=2.99
r67 17 24 6.87494 $w=1.7e-07 $l=1.36015e-07 $layer=LI1_cond $X=3.535 $Y=2.99
+ $X2=3.635 $Y2=2.905
r68 17 18 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.535 $Y=2.99
+ $X2=2.865 $Y2=2.99
r69 13 38 2.85134 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=2.735 $Y=2.905
+ $X2=2.735 $Y2=2.99
r70 13 15 35.903 $w=2.58e-07 $l=8.1e-07 $layer=LI1_cond $X=2.735 $Y=2.905
+ $X2=2.735 $Y2=2.095
r71 4 44 300 $w=1.7e-07 $l=6.81414e-07 $layer=licon1_PDIFF $count=2 $X=5.25
+ $Y=1.835 $X2=5.39 $Y2=2.45
r72 4 33 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=5.25
+ $Y=1.835 $X2=5.39 $Y2=1.98
r73 3 42 300 $w=1.7e-07 $l=6.96491e-07 $layer=licon1_PDIFF $count=2 $X=4.39
+ $Y=1.835 $X2=4.53 $Y2=2.465
r74 2 40 300 $w=1.7e-07 $l=6.81414e-07 $layer=licon1_PDIFF $count=2 $X=3.49
+ $Y=1.835 $X2=3.63 $Y2=2.45
r75 2 21 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=3.49
+ $Y=1.835 $X2=3.63 $Y2=1.98
r76 1 38 400 $w=1.7e-07 $l=1.17584e-06 $layer=licon1_PDIFF $count=1 $X=2.645
+ $Y=1.835 $X2=2.77 $Y2=2.95
r77 1 15 400 $w=1.7e-07 $l=3.16386e-07 $layer=licon1_PDIFF $count=1 $X=2.645
+ $Y=1.835 $X2=2.77 $Y2=2.095
.ends

.subckt PM_SKY130_FD_SC_LP__A21O_4%VGND 1 2 3 4 5 18 22 26 28 30 33 34 35 37 46
+ 50 55 64 74 78
r83 77 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r84 74 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r85 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r86 62 78 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=5.52
+ $Y2=0
r87 61 62 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r88 59 62 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=5.04
+ $Y2=0
r89 59 75 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.6
+ $Y2=0
r90 58 61 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=4.08 $Y=0 $X2=5.04
+ $Y2=0
r91 58 59 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r92 56 74 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=3.815 $Y=0 $X2=3.645
+ $Y2=0
r93 56 58 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=3.815 $Y=0 $X2=4.08
+ $Y2=0
r94 55 77 4.26799 $w=1.7e-07 $l=2.5e-07 $layer=LI1_cond $X=5.26 $Y=0 $X2=5.51
+ $Y2=0
r95 55 61 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=5.26 $Y=0 $X2=5.04
+ $Y2=0
r96 54 75 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r97 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r98 51 53 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=2.895 $Y=0 $X2=3.12
+ $Y2=0
r99 50 74 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=3.475 $Y=0 $X2=3.645
+ $Y2=0
r100 50 53 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=3.475 $Y=0
+ $X2=3.12 $Y2=0
r101 49 69 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r102 48 49 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r103 46 71 9.7695 $w=6.53e-07 $l=5.35e-07 $layer=LI1_cond $X=2.567 $Y=0
+ $X2=2.567 $Y2=0.535
r104 46 51 8.8858 $w=1.7e-07 $l=3.28e-07 $layer=LI1_cond $X=2.567 $Y=0 $X2=2.895
+ $Y2=0
r105 46 69 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r106 46 48 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=2.24 $Y=0 $X2=2.16
+ $Y2=0
r107 45 49 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r108 45 65 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r109 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r110 42 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.815 $Y=0 $X2=0.65
+ $Y2=0
r111 42 44 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=0.815 $Y=0 $X2=1.2
+ $Y2=0
r112 40 65 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r113 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r114 37 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.485 $Y=0 $X2=0.65
+ $Y2=0
r115 37 39 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=0.485 $Y=0 $X2=0.24
+ $Y2=0
r116 35 54 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.88 $Y=0
+ $X2=3.12 $Y2=0
r117 35 69 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.88 $Y=0
+ $X2=2.64 $Y2=0
r118 33 44 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=1.345 $Y=0 $X2=1.2
+ $Y2=0
r119 33 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.345 $Y=0 $X2=1.51
+ $Y2=0
r120 32 48 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=1.675 $Y=0
+ $X2=2.16 $Y2=0
r121 32 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.675 $Y=0 $X2=1.51
+ $Y2=0
r122 28 77 3.20953 $w=2.95e-07 $l=1.39155e-07 $layer=LI1_cond $X=5.407 $Y=0.085
+ $X2=5.51 $Y2=0
r123 28 30 11.9151 $w=2.93e-07 $l=3.05e-07 $layer=LI1_cond $X=5.407 $Y=0.085
+ $X2=5.407 $Y2=0.39
r124 24 74 0.987631 $w=3.4e-07 $l=8.5e-08 $layer=LI1_cond $X=3.645 $Y=0.085
+ $X2=3.645 $Y2=0
r125 24 26 14.914 $w=3.38e-07 $l=4.4e-07 $layer=LI1_cond $X=3.645 $Y=0.085
+ $X2=3.645 $Y2=0.525
r126 20 34 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.51 $Y=0.085
+ $X2=1.51 $Y2=0
r127 20 22 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=1.51 $Y=0.085
+ $X2=1.51 $Y2=0.39
r128 16 64 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.65 $Y=0.085
+ $X2=0.65 $Y2=0
r129 16 18 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=0.65 $Y=0.085
+ $X2=0.65 $Y2=0.39
r130 5 30 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.25
+ $Y=0.245 $X2=5.39 $Y2=0.39
r131 4 26 182 $w=1.7e-07 $l=3.50999e-07 $layer=licon1_NDIFF $count=1 $X=3.49
+ $Y=0.245 $X2=3.65 $Y2=0.525
r132 3 71 91 $w=1.7e-07 $l=6.69477e-07 $layer=licon1_NDIFF $count=2 $X=2.23
+ $Y=0.245 $X2=2.77 $Y2=0.535
r133 2 22 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.37
+ $Y=0.245 $X2=1.51 $Y2=0.39
r134 1 18 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.525
+ $Y=0.245 $X2=0.65 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_LP__A21O_4%A_792_49# 1 2 7 11 17
r21 11 14 8.29759 $w=2.48e-07 $l=1.8e-07 $layer=LI1_cond $X=4.11 $Y=0.345
+ $X2=4.11 $Y2=0.525
r22 8 11 2.6621 $w=1.8e-07 $l=1.25e-07 $layer=LI1_cond $X=4.235 $Y=0.345
+ $X2=4.11 $Y2=0.345
r23 7 17 4.55851 $w=1.8e-07 $l=1.47e-07 $layer=LI1_cond $X=4.795 $Y=0.345
+ $X2=4.942 $Y2=0.345
r24 7 8 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=4.795 $Y=0.345
+ $X2=4.235 $Y2=0.345
r25 2 17 91 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_NDIFF $count=2 $X=4.82
+ $Y=0.245 $X2=4.96 $Y2=0.42
r26 1 14 182 $w=1.7e-07 $l=3.42929e-07 $layer=licon1_NDIFF $count=1 $X=3.96
+ $Y=0.245 $X2=4.1 $Y2=0.525
.ends

