* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__o221a_m A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
X0 VPWR a_27_179# X VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X1 a_110_179# B1 a_196_179# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 a_396_535# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X3 VGND A2 a_196_179# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 a_27_179# A2 a_396_535# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X5 a_238_535# B2 a_27_179# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X6 a_27_179# C1 a_110_179# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 a_196_179# B2 a_110_179# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 a_27_179# C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X9 a_196_179# A1 VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 VPWR B1 a_238_535# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X11 VGND a_27_179# X VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
