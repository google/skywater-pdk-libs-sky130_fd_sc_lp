* File: sky130_fd_sc_lp__or3b_1.spice
* Created: Fri Aug 28 11:23:55 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__or3b_1.pex.spice"
.subckt sky130_fd_sc_lp__or3b_1  VNB VPB C_N B A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* B	B
* C_N	C_N
* VPB	VPB
* VNB	VNB
MM1003 N_A_110_70#_M1003_d N_C_N_M1003_g N_VGND_M1003_s VNB NSHORT L=0.15 W=0.42
+ AD=0.1113 AS=0.1113 PD=1.37 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1008 N_VGND_M1008_d N_A_110_70#_M1008_g N_A_220_74#_M1008_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0672 AS=0.1113 PD=0.74 PS=1.37 NRD=5.712 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.6 A=0.063 P=1.14 MULT=1
MM1007 N_A_220_74#_M1007_d N_B_M1007_g N_VGND_M1008_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0672 PD=0.7 PS=0.74 NRD=0 NRS=5.712 M=1 R=2.8 SA=75000.7
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1002 N_VGND_M1002_d N_A_M1002_g N_A_220_74#_M1007_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0896 AS=0.0588 PD=0.81 PS=0.7 NRD=12.852 NRS=0 M=1 R=2.8 SA=75001.1
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1005 N_X_M1005_d N_A_220_74#_M1005_g N_VGND_M1002_d VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1792 PD=2.21 PS=1.62 NRD=0 NRS=3.564 M=1 R=5.6 SA=75000.9
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1006 N_A_110_70#_M1006_d N_C_N_M1006_g N_VPWR_M1006_s VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1113 AS=0.1113 PD=1.37 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1009 A_303_367# N_A_110_70#_M1009_g N_A_220_74#_M1009_s VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0441 AS=0.1113 PD=0.63 PS=1.37 NRD=23.443 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.6 A=0.063 P=1.14 MULT=1
MM1000 A_375_367# N_B_M1000_g A_303_367# VPB PHIGHVT L=0.15 W=0.42 AD=0.0819
+ AS=0.0441 PD=0.81 PS=0.63 NRD=65.6601 NRS=23.443 M=1 R=2.8 SA=75000.6
+ SB=75001.3 A=0.063 P=1.14 MULT=1
MM1004 N_VPWR_M1004_d N_A_M1004_g A_375_367# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.095025 AS=0.0819 PD=0.8175 PS=0.81 NRD=23.443 NRS=65.6601 M=1 R=2.8
+ SA=75001.1 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1001 N_X_M1001_d N_A_220_74#_M1001_g N_VPWR_M1004_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.285075 PD=3.05 PS=2.4525 NRD=0 NRS=2.3443 M=1 R=8.4 SA=75000.7
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9751 P=11.21
c_39 VNB 0 6.36774e-20 $X=0 $Y=0
*
.include "sky130_fd_sc_lp__or3b_1.pxi.spice"
*
.ends
*
*
