* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__dfxbp_1 CLK D VGND VNB VPB VPWR Q Q_N
X0 VGND a_526_463# a_697_93# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X1 a_1401_22# a_1149_93# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X2 a_440_463# a_110_82# a_526_463# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 a_997_119# a_110_82# a_1105_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 a_440_463# a_217_463# a_526_463# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X5 a_1401_22# a_1149_93# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 a_650_499# a_697_93# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X7 VPWR a_997_119# a_1149_93# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X8 a_697_93# a_217_463# a_997_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 VGND D a_440_463# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 VGND a_997_119# a_1149_93# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X11 VPWR CLK a_110_82# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X12 a_1137_379# a_1149_93# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X13 a_526_463# a_217_463# a_655_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X14 a_697_93# a_110_82# a_997_119# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X15 VPWR a_1401_22# Q_N VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X16 a_1105_119# a_1149_93# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X17 VPWR a_1149_93# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X18 a_217_463# a_110_82# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X19 VGND a_1401_22# Q_N VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X20 VPWR D a_440_463# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X21 a_655_119# a_697_93# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X22 VGND a_1149_93# Q VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X23 VGND CLK a_110_82# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X24 a_526_463# a_110_82# a_650_499# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X25 a_217_463# a_110_82# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X26 VPWR a_526_463# a_697_93# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X27 a_997_119# a_217_463# a_1137_379# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
.ends
