* File: sky130_fd_sc_lp__o211a_2.pxi.spice
* Created: Fri Aug 28 11:02:02 2020
* 
x_PM_SKY130_FD_SC_LP__O211A_2%C1 N_C1_M1006_g N_C1_c_70_n N_C1_M1010_g C1
+ N_C1_c_69_n PM_SKY130_FD_SC_LP__O211A_2%C1
x_PM_SKY130_FD_SC_LP__O211A_2%B1 N_B1_c_93_n N_B1_M1000_g N_B1_M1007_g B1
+ N_B1_c_96_n PM_SKY130_FD_SC_LP__O211A_2%B1
x_PM_SKY130_FD_SC_LP__O211A_2%A2 N_A2_c_129_n N_A2_M1004_g N_A2_c_130_n
+ N_A2_M1003_g A2 A2 A2 PM_SKY130_FD_SC_LP__O211A_2%A2
x_PM_SKY130_FD_SC_LP__O211A_2%A1 N_A1_M1005_g N_A1_M1011_g A1 A1 A1 N_A1_c_174_n
+ N_A1_c_175_n PM_SKY130_FD_SC_LP__O211A_2%A1
x_PM_SKY130_FD_SC_LP__O211A_2%A_27_47# N_A_27_47#_M1006_s N_A_27_47#_M1010_s
+ N_A_27_47#_M1007_d N_A_27_47#_M1002_g N_A_27_47#_M1001_g N_A_27_47#_M1008_g
+ N_A_27_47#_M1009_g N_A_27_47#_c_214_n N_A_27_47#_c_223_n N_A_27_47#_c_215_n
+ N_A_27_47#_c_216_n N_A_27_47#_c_250_n N_A_27_47#_c_252_n N_A_27_47#_c_217_n
+ N_A_27_47#_c_218_n N_A_27_47#_c_226_n N_A_27_47#_c_255_n N_A_27_47#_c_219_n
+ N_A_27_47#_c_220_n PM_SKY130_FD_SC_LP__O211A_2%A_27_47#
x_PM_SKY130_FD_SC_LP__O211A_2%VPWR N_VPWR_M1010_d N_VPWR_M1005_d N_VPWR_M1009_s
+ N_VPWR_c_320_n N_VPWR_c_321_n N_VPWR_c_322_n VPWR N_VPWR_c_323_n
+ N_VPWR_c_324_n N_VPWR_c_325_n N_VPWR_c_326_n N_VPWR_c_319_n
+ PM_SKY130_FD_SC_LP__O211A_2%VPWR
x_PM_SKY130_FD_SC_LP__O211A_2%X N_X_M1002_s N_X_M1001_d N_X_c_371_n N_X_c_388_n
+ X X X PM_SKY130_FD_SC_LP__O211A_2%X
x_PM_SKY130_FD_SC_LP__O211A_2%A_182_47# N_A_182_47#_M1000_d N_A_182_47#_M1004_d
+ N_A_182_47#_c_401_n N_A_182_47#_c_402_n N_A_182_47#_c_403_n
+ N_A_182_47#_c_417_n N_A_182_47#_c_404_n PM_SKY130_FD_SC_LP__O211A_2%A_182_47#
x_PM_SKY130_FD_SC_LP__O211A_2%VGND N_VGND_M1004_s N_VGND_M1011_d N_VGND_M1008_d
+ N_VGND_c_434_n N_VGND_c_435_n N_VGND_c_436_n N_VGND_c_437_n N_VGND_c_438_n
+ N_VGND_c_439_n N_VGND_c_440_n N_VGND_c_441_n VGND N_VGND_c_442_n
+ N_VGND_c_443_n PM_SKY130_FD_SC_LP__O211A_2%VGND
cc_1 VNB N_C1_M1006_g 0.0244531f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.655
cc_2 VNB C1 0.00326334f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_3 VNB N_C1_c_69_n 0.0627346f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.485
cc_4 VNB N_B1_c_93_n 0.0216028f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.245
cc_5 VNB N_B1_M1007_g 0.00793938f $X=-0.19 $Y=-0.245 $X2=0.645 $Y2=2.465
cc_6 VNB B1 0.00341502f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_7 VNB N_B1_c_96_n 0.0419665f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.41
cc_8 VNB N_A2_c_129_n 0.0205256f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.245
cc_9 VNB N_A2_c_130_n 0.0449888f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_10 VNB N_A2_M1003_g 7.39226e-19 $X=-0.19 $Y=-0.245 $X2=0.645 $Y2=2.465
cc_11 VNB A2 0.00131981f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_12 VNB N_A1_M1005_g 0.00420322f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.655
cc_13 VNB A1 0.00598061f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_14 VNB N_A1_c_174_n 0.032587f $X=-0.19 $Y=-0.245 $X2=0.255 $Y2=1.295
cc_15 VNB N_A1_c_175_n 0.0171045f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_27_47#_M1002_g 0.0201075f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.41
cc_17 VNB N_A_27_47#_M1001_g 0.00147254f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_27_47#_M1008_g 0.0228451f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_27_47#_M1009_g 0.00156298f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_27_47#_c_214_n 0.0237941f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_27_47#_c_215_n 0.0040499f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_27_47#_c_216_n 0.00704914f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_27_47#_c_217_n 7.64562e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_27_47#_c_218_n 0.00816863f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB N_A_27_47#_c_219_n 0.00481921f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_A_27_47#_c_220_n 0.0653565f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_VPWR_c_319_n 0.163682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_X_c_371_n 0.00203831f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB X 0.024651f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB X 0.00709178f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_182_47#_c_401_n 0.00671676f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_182_47#_c_402_n 0.0116411f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.41
cc_33 VNB N_A_182_47#_c_403_n 4.81195e-19 $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.41
cc_34 VNB N_A_182_47#_c_404_n 0.00181827f $X=-0.19 $Y=-0.245 $X2=0.255 $Y2=1.295
cc_35 VNB N_VGND_c_434_n 0.00803496f $X=-0.19 $Y=-0.245 $X2=0.27 $Y2=1.41
cc_36 VNB N_VGND_c_435_n 0.0048727f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_436_n 0.0166207f $X=-0.19 $Y=-0.245 $X2=0.255 $Y2=1.41
cc_38 VNB N_VGND_c_437_n 0.0394174f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_438_n 0.0406434f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_439_n 0.00547551f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_440_n 0.0159219f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_441_n 0.00442067f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_442_n 0.017949f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_443_n 0.232213f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VPB N_C1_c_70_n 0.0197428f $X=-0.19 $Y=1.655 $X2=0.645 $Y2=1.725
cc_46 VPB N_C1_c_69_n 0.0255096f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=1.485
cc_47 VPB N_B1_M1007_g 0.0209392f $X=-0.19 $Y=1.655 $X2=0.645 $Y2=2.465
cc_48 VPB N_A2_M1003_g 0.0208455f $X=-0.19 $Y=1.655 $X2=0.645 $Y2=2.465
cc_49 VPB A2 0.00123092f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_50 VPB N_A1_M1005_g 0.0200456f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.655
cc_51 VPB A1 0.00247198f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_52 VPB N_A_27_47#_M1001_g 0.022707f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_53 VPB N_A_27_47#_M1009_g 0.0227978f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_54 VPB N_A_27_47#_c_223_n 0.0442891f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_55 VPB N_A_27_47#_c_216_n 0.001484f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_56 VPB N_A_27_47#_c_217_n 0.00275268f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_57 VPB N_A_27_47#_c_226_n 0.0104464f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_58 VPB N_VPWR_c_320_n 4.89148e-19 $X=-0.19 $Y=1.655 $X2=0.645 $Y2=1.725
cc_59 VPB N_VPWR_c_321_n 0.0109777f $X=-0.19 $Y=1.655 $X2=0.255 $Y2=1.41
cc_60 VPB N_VPWR_c_322_n 0.0352627f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_61 VPB N_VPWR_c_323_n 0.0307198f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_62 VPB N_VPWR_c_324_n 0.0129657f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_63 VPB N_VPWR_c_325_n 0.0256026f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_64 VPB N_VPWR_c_326_n 0.0123114f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_319_n 0.0522338f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_66 VPB X 0.00841928f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_67 N_C1_M1006_g N_B1_c_93_n 0.0365354f $X=0.475 $Y=0.655 $X2=-0.19 $Y2=-0.245
cc_68 N_C1_c_69_n N_B1_M1007_g 0.0216603f $X=0.475 $Y=1.485 $X2=0 $Y2=0
cc_69 N_C1_c_69_n N_B1_c_96_n 0.0418835f $X=0.475 $Y=1.485 $X2=0 $Y2=0
cc_70 N_C1_M1006_g N_A_27_47#_c_214_n 0.0131664f $X=0.475 $Y=0.655 $X2=0 $Y2=0
cc_71 N_C1_M1006_g N_A_27_47#_c_215_n 0.0085199f $X=0.475 $Y=0.655 $X2=0 $Y2=0
cc_72 C1 N_A_27_47#_c_215_n 0.0252617f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_73 N_C1_c_69_n N_A_27_47#_c_215_n 0.0163186f $X=0.475 $Y=1.485 $X2=0 $Y2=0
cc_74 N_C1_c_70_n N_A_27_47#_c_216_n 0.00316071f $X=0.645 $Y=1.725 $X2=0 $Y2=0
cc_75 N_C1_c_69_n N_A_27_47#_c_216_n 0.00178105f $X=0.475 $Y=1.485 $X2=0 $Y2=0
cc_76 N_C1_M1006_g N_A_27_47#_c_218_n 0.0123416f $X=0.475 $Y=0.655 $X2=0 $Y2=0
cc_77 C1 N_A_27_47#_c_218_n 0.0152919f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_78 N_C1_c_69_n N_A_27_47#_c_218_n 0.00351078f $X=0.475 $Y=1.485 $X2=0 $Y2=0
cc_79 N_C1_c_70_n N_A_27_47#_c_226_n 0.0114329f $X=0.645 $Y=1.725 $X2=0 $Y2=0
cc_80 C1 N_A_27_47#_c_226_n 0.00759321f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_81 N_C1_c_69_n N_A_27_47#_c_226_n 0.0188041f $X=0.475 $Y=1.485 $X2=0 $Y2=0
cc_82 N_C1_c_70_n N_VPWR_c_320_n 0.0141348f $X=0.645 $Y=1.725 $X2=0 $Y2=0
cc_83 N_C1_c_70_n N_VPWR_c_325_n 0.00564095f $X=0.645 $Y=1.725 $X2=0 $Y2=0
cc_84 N_C1_c_70_n N_VPWR_c_319_n 0.0105414f $X=0.645 $Y=1.725 $X2=0 $Y2=0
cc_85 N_C1_M1006_g N_A_182_47#_c_401_n 0.00161761f $X=0.475 $Y=0.655 $X2=0 $Y2=0
cc_86 N_C1_M1006_g N_VGND_c_438_n 0.0054895f $X=0.475 $Y=0.655 $X2=0 $Y2=0
cc_87 N_C1_M1006_g N_VGND_c_443_n 0.00709137f $X=0.475 $Y=0.655 $X2=0 $Y2=0
cc_88 N_B1_c_96_n N_A2_c_129_n 0.00136734f $X=1.095 $Y=1.35 $X2=-0.19 $Y2=-0.245
cc_89 N_B1_M1007_g N_A2_c_130_n 0.00611892f $X=1.115 $Y=2.465 $X2=0 $Y2=0
cc_90 B1 N_A2_c_130_n 0.00178173f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_91 N_B1_c_96_n N_A2_c_130_n 0.0183919f $X=1.095 $Y=1.35 $X2=0 $Y2=0
cc_92 N_B1_M1007_g N_A2_M1003_g 0.0226384f $X=1.115 $Y=2.465 $X2=0 $Y2=0
cc_93 N_B1_M1007_g A2 0.00117084f $X=1.115 $Y=2.465 $X2=0 $Y2=0
cc_94 B1 A2 0.0128887f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_95 N_B1_c_96_n A2 5.63182e-19 $X=1.095 $Y=1.35 $X2=0 $Y2=0
cc_96 N_B1_c_93_n N_A_27_47#_c_214_n 0.00168111f $X=0.835 $Y=1.185 $X2=0 $Y2=0
cc_97 N_B1_c_93_n N_A_27_47#_c_215_n 0.00424744f $X=0.835 $Y=1.185 $X2=0 $Y2=0
cc_98 N_B1_M1007_g N_A_27_47#_c_215_n 0.00150382f $X=1.115 $Y=2.465 $X2=0 $Y2=0
cc_99 B1 N_A_27_47#_c_215_n 0.0159315f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_100 N_B1_c_96_n N_A_27_47#_c_215_n 0.0014587f $X=1.095 $Y=1.35 $X2=0 $Y2=0
cc_101 N_B1_M1007_g N_A_27_47#_c_216_n 0.0189167f $X=1.115 $Y=2.465 $X2=0 $Y2=0
cc_102 B1 N_A_27_47#_c_216_n 0.0271162f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_103 N_B1_c_96_n N_A_27_47#_c_216_n 0.0101184f $X=1.095 $Y=1.35 $X2=0 $Y2=0
cc_104 N_B1_M1007_g N_VPWR_c_320_n 0.0136743f $X=1.115 $Y=2.465 $X2=0 $Y2=0
cc_105 N_B1_M1007_g N_VPWR_c_323_n 0.00564095f $X=1.115 $Y=2.465 $X2=0 $Y2=0
cc_106 N_B1_M1007_g N_VPWR_c_319_n 0.0101267f $X=1.115 $Y=2.465 $X2=0 $Y2=0
cc_107 N_B1_c_93_n N_A_182_47#_c_401_n 0.0118182f $X=0.835 $Y=1.185 $X2=0 $Y2=0
cc_108 B1 N_A_182_47#_c_402_n 0.00522897f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_109 N_B1_c_96_n N_A_182_47#_c_402_n 0.00103667f $X=1.095 $Y=1.35 $X2=0 $Y2=0
cc_110 N_B1_c_93_n N_A_182_47#_c_403_n 0.00225996f $X=0.835 $Y=1.185 $X2=0 $Y2=0
cc_111 B1 N_A_182_47#_c_403_n 0.0215594f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_112 N_B1_c_96_n N_A_182_47#_c_403_n 0.00767923f $X=1.095 $Y=1.35 $X2=0 $Y2=0
cc_113 N_B1_c_93_n N_VGND_c_434_n 0.00338638f $X=0.835 $Y=1.185 $X2=0 $Y2=0
cc_114 N_B1_c_93_n N_VGND_c_438_n 0.0054945f $X=0.835 $Y=1.185 $X2=0 $Y2=0
cc_115 N_B1_c_93_n N_VGND_c_443_n 0.0112336f $X=0.835 $Y=1.185 $X2=0 $Y2=0
cc_116 N_A2_M1003_g N_A1_M1005_g 0.061083f $X=1.785 $Y=2.465 $X2=0 $Y2=0
cc_117 N_A2_c_129_n A1 0.00453785f $X=1.785 $Y=1.23 $X2=0 $Y2=0
cc_118 A2 A1 0.049049f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_119 N_A2_c_130_n N_A1_c_174_n 0.061083f $X=1.785 $Y=1.64 $X2=0 $Y2=0
cc_120 A2 N_A1_c_174_n 9.67795e-19 $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_121 N_A2_c_129_n N_A1_c_175_n 0.0167445f $X=1.785 $Y=1.23 $X2=0 $Y2=0
cc_122 A2 N_A_27_47#_M1007_d 0.00325389f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_123 N_A2_M1003_g N_A_27_47#_c_216_n 9.73652e-19 $X=1.785 $Y=2.465 $X2=0 $Y2=0
cc_124 A2 N_A_27_47#_c_216_n 0.023386f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_125 N_A2_M1003_g N_A_27_47#_c_250_n 0.00410407f $X=1.785 $Y=2.465 $X2=0 $Y2=0
cc_126 A2 N_A_27_47#_c_250_n 0.0153851f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_127 N_A2_c_130_n N_A_27_47#_c_252_n 2.02544e-19 $X=1.785 $Y=1.64 $X2=0 $Y2=0
cc_128 N_A2_M1003_g N_A_27_47#_c_252_n 0.0168584f $X=1.785 $Y=2.465 $X2=0 $Y2=0
cc_129 A2 N_A_27_47#_c_252_n 0.0109774f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_130 N_A2_c_130_n N_A_27_47#_c_255_n 0.00353749f $X=1.785 $Y=1.64 $X2=0 $Y2=0
cc_131 N_A2_M1003_g N_A_27_47#_c_255_n 0.0118661f $X=1.785 $Y=2.465 $X2=0 $Y2=0
cc_132 A2 N_A_27_47#_c_255_n 0.00171307f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_133 N_A2_M1003_g N_VPWR_c_320_n 0.0010085f $X=1.785 $Y=2.465 $X2=0 $Y2=0
cc_134 N_A2_M1003_g N_VPWR_c_323_n 0.00585385f $X=1.785 $Y=2.465 $X2=0 $Y2=0
cc_135 N_A2_M1003_g N_VPWR_c_326_n 0.00258111f $X=1.785 $Y=2.465 $X2=0 $Y2=0
cc_136 N_A2_M1003_g N_VPWR_c_319_n 0.0113489f $X=1.785 $Y=2.465 $X2=0 $Y2=0
cc_137 N_A2_c_129_n N_A_182_47#_c_401_n 0.00455563f $X=1.785 $Y=1.23 $X2=0 $Y2=0
cc_138 N_A2_c_129_n N_A_182_47#_c_402_n 0.0156701f $X=1.785 $Y=1.23 $X2=0 $Y2=0
cc_139 N_A2_c_130_n N_A_182_47#_c_402_n 0.00539168f $X=1.785 $Y=1.64 $X2=0 $Y2=0
cc_140 A2 N_A_182_47#_c_402_n 0.0153197f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_141 N_A2_c_129_n N_A_182_47#_c_404_n 6.2974e-19 $X=1.785 $Y=1.23 $X2=0 $Y2=0
cc_142 N_A2_c_129_n N_VGND_c_434_n 0.0115981f $X=1.785 $Y=1.23 $X2=0 $Y2=0
cc_143 N_A2_c_129_n N_VGND_c_440_n 0.00448994f $X=1.785 $Y=1.23 $X2=0 $Y2=0
cc_144 N_A2_c_129_n N_VGND_c_443_n 0.00814279f $X=1.785 $Y=1.23 $X2=0 $Y2=0
cc_145 A1 N_A_27_47#_M1002_g 7.6982e-19 $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_146 N_A1_c_174_n N_A_27_47#_M1002_g 0.0205185f $X=2.235 $Y=1.395 $X2=0 $Y2=0
cc_147 N_A1_c_175_n N_A_27_47#_M1002_g 0.0135438f $X=2.235 $Y=1.23 $X2=0 $Y2=0
cc_148 N_A1_M1005_g N_A_27_47#_M1001_g 0.0154407f $X=2.145 $Y=2.465 $X2=0 $Y2=0
cc_149 N_A1_M1005_g N_A_27_47#_c_252_n 0.0148306f $X=2.145 $Y=2.465 $X2=0 $Y2=0
cc_150 A1 N_A_27_47#_c_252_n 0.0148434f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_151 N_A1_M1005_g N_A_27_47#_c_217_n 0.00511112f $X=2.145 $Y=2.465 $X2=0 $Y2=0
cc_152 A1 N_A_27_47#_c_217_n 0.0380915f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_153 A1 N_A_27_47#_c_219_n 0.0263702f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_154 N_A1_c_174_n N_A_27_47#_c_219_n 0.0017709f $X=2.235 $Y=1.395 $X2=0 $Y2=0
cc_155 N_A1_M1005_g N_A_27_47#_c_220_n 0.00198404f $X=2.145 $Y=2.465 $X2=0 $Y2=0
cc_156 A1 N_A_27_47#_c_220_n 4.05909e-19 $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_157 A1 N_VPWR_M1005_d 0.00322827f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_158 N_A1_M1005_g N_VPWR_c_323_n 0.00487821f $X=2.145 $Y=2.465 $X2=0 $Y2=0
cc_159 N_A1_M1005_g N_VPWR_c_326_n 0.0173219f $X=2.145 $Y=2.465 $X2=0 $Y2=0
cc_160 N_A1_M1005_g N_VPWR_c_319_n 0.00818716f $X=2.145 $Y=2.465 $X2=0 $Y2=0
cc_161 N_A1_c_175_n X 3.59176e-19 $X=2.235 $Y=1.23 $X2=0 $Y2=0
cc_162 A1 N_A_182_47#_c_417_n 0.0099843f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_163 N_A1_c_174_n N_A_182_47#_c_417_n 3.51706e-19 $X=2.235 $Y=1.395 $X2=0
+ $Y2=0
cc_164 N_A1_c_175_n N_A_182_47#_c_417_n 0.00208374f $X=2.235 $Y=1.23 $X2=0 $Y2=0
cc_165 N_A1_c_175_n N_A_182_47#_c_404_n 0.00758856f $X=2.235 $Y=1.23 $X2=0 $Y2=0
cc_166 N_A1_c_175_n N_VGND_c_434_n 5.62083e-19 $X=2.235 $Y=1.23 $X2=0 $Y2=0
cc_167 N_A1_c_174_n N_VGND_c_435_n 0.00252309f $X=2.235 $Y=1.395 $X2=0 $Y2=0
cc_168 N_A1_c_175_n N_VGND_c_435_n 0.00180445f $X=2.235 $Y=1.23 $X2=0 $Y2=0
cc_169 N_A1_c_175_n N_VGND_c_440_n 0.00507287f $X=2.235 $Y=1.23 $X2=0 $Y2=0
cc_170 N_A1_c_175_n N_VGND_c_443_n 0.00955246f $X=2.235 $Y=1.23 $X2=0 $Y2=0
cc_171 N_A_27_47#_c_216_n N_VPWR_M1010_d 0.0022225f $X=1.215 $Y=1.777 $X2=-0.19
+ $Y2=-0.245
cc_172 N_A_27_47#_c_252_n N_VPWR_M1005_d 0.0155316f $X=2.49 $Y=2.375 $X2=0 $Y2=0
cc_173 N_A_27_47#_c_217_n N_VPWR_M1005_d 0.014077f $X=2.575 $Y=2.29 $X2=0 $Y2=0
cc_174 N_A_27_47#_c_216_n N_VPWR_c_320_n 0.0178669f $X=1.215 $Y=1.777 $X2=0
+ $Y2=0
cc_175 N_A_27_47#_M1001_g N_VPWR_c_322_n 6.72004e-19 $X=2.915 $Y=2.465 $X2=0
+ $Y2=0
cc_176 N_A_27_47#_M1009_g N_VPWR_c_322_n 0.0166575f $X=3.345 $Y=2.465 $X2=0
+ $Y2=0
cc_177 N_A_27_47#_c_255_n N_VPWR_c_323_n 0.0269046f $X=1.45 $Y=2.43 $X2=0 $Y2=0
cc_178 N_A_27_47#_M1001_g N_VPWR_c_324_n 0.00487821f $X=2.915 $Y=2.465 $X2=0
+ $Y2=0
cc_179 N_A_27_47#_M1009_g N_VPWR_c_324_n 0.00486043f $X=3.345 $Y=2.465 $X2=0
+ $Y2=0
cc_180 N_A_27_47#_c_223_n N_VPWR_c_325_n 0.0185207f $X=0.43 $Y=1.98 $X2=0 $Y2=0
cc_181 N_A_27_47#_M1001_g N_VPWR_c_326_n 0.01354f $X=2.915 $Y=2.465 $X2=0 $Y2=0
cc_182 N_A_27_47#_M1009_g N_VPWR_c_326_n 5.90548e-19 $X=3.345 $Y=2.465 $X2=0
+ $Y2=0
cc_183 N_A_27_47#_c_252_n N_VPWR_c_326_n 0.0343163f $X=2.49 $Y=2.375 $X2=0 $Y2=0
cc_184 N_A_27_47#_c_255_n N_VPWR_c_326_n 0.0140538f $X=1.45 $Y=2.43 $X2=0 $Y2=0
cc_185 N_A_27_47#_M1010_s N_VPWR_c_319_n 0.00302127f $X=0.305 $Y=1.835 $X2=0
+ $Y2=0
cc_186 N_A_27_47#_M1007_d N_VPWR_c_319_n 0.00847955f $X=1.19 $Y=1.835 $X2=0
+ $Y2=0
cc_187 N_A_27_47#_M1001_g N_VPWR_c_319_n 0.00824731f $X=2.915 $Y=2.465 $X2=0
+ $Y2=0
cc_188 N_A_27_47#_M1009_g N_VPWR_c_319_n 0.00824727f $X=3.345 $Y=2.465 $X2=0
+ $Y2=0
cc_189 N_A_27_47#_c_223_n N_VPWR_c_319_n 0.010808f $X=0.43 $Y=1.98 $X2=0 $Y2=0
cc_190 N_A_27_47#_c_255_n N_VPWR_c_319_n 0.0154733f $X=1.45 $Y=2.43 $X2=0 $Y2=0
cc_191 N_A_27_47#_c_252_n A_372_367# 0.00732587f $X=2.49 $Y=2.375 $X2=-0.19
+ $Y2=-0.245
cc_192 N_A_27_47#_M1002_g N_X_c_371_n 0.00938439f $X=2.685 $Y=0.7 $X2=0 $Y2=0
cc_193 N_A_27_47#_M1008_g N_X_c_371_n 0.0103034f $X=3.115 $Y=0.7 $X2=0 $Y2=0
cc_194 N_A_27_47#_M1002_g X 0.00622575f $X=2.685 $Y=0.7 $X2=0 $Y2=0
cc_195 N_A_27_47#_M1008_g X 0.0168397f $X=3.115 $Y=0.7 $X2=0 $Y2=0
cc_196 N_A_27_47#_c_219_n X 0.0246205f $X=2.775 $Y=1.46 $X2=0 $Y2=0
cc_197 N_A_27_47#_c_220_n X 0.0201247f $X=3.115 $Y=1.462 $X2=0 $Y2=0
cc_198 N_A_27_47#_M1009_g X 0.00972414f $X=3.345 $Y=2.465 $X2=0 $Y2=0
cc_199 N_A_27_47#_c_217_n X 0.0192136f $X=2.575 $Y=2.29 $X2=0 $Y2=0
cc_200 N_A_27_47#_c_219_n X 0.011426f $X=2.775 $Y=1.46 $X2=0 $Y2=0
cc_201 N_A_27_47#_c_220_n X 0.0147379f $X=3.115 $Y=1.462 $X2=0 $Y2=0
cc_202 N_A_27_47#_M1009_g X 0.0135118f $X=3.345 $Y=2.465 $X2=0 $Y2=0
cc_203 N_A_27_47#_c_215_n A_110_47# 2.83863e-19 $X=0.615 $Y=1.64 $X2=-0.19
+ $Y2=-0.245
cc_204 N_A_27_47#_c_218_n A_110_47# 0.00223753f $X=0.615 $Y=0.95 $X2=-0.19
+ $Y2=-0.245
cc_205 N_A_27_47#_c_214_n N_A_182_47#_c_401_n 0.0197398f $X=0.26 $Y=0.38 $X2=0
+ $Y2=0
cc_206 N_A_27_47#_c_216_n N_A_182_47#_c_402_n 0.00490595f $X=1.215 $Y=1.777
+ $X2=0 $Y2=0
cc_207 N_A_27_47#_c_216_n N_A_182_47#_c_403_n 0.00110939f $X=1.215 $Y=1.777
+ $X2=0 $Y2=0
cc_208 N_A_27_47#_M1002_g N_VGND_c_435_n 0.00178387f $X=2.685 $Y=0.7 $X2=0 $Y2=0
cc_209 N_A_27_47#_c_219_n N_VGND_c_435_n 0.0044237f $X=2.775 $Y=1.46 $X2=0 $Y2=0
cc_210 N_A_27_47#_M1008_g N_VGND_c_437_n 0.00750862f $X=3.115 $Y=0.7 $X2=0 $Y2=0
cc_211 N_A_27_47#_c_220_n N_VGND_c_437_n 0.00114149f $X=3.115 $Y=1.462 $X2=0
+ $Y2=0
cc_212 N_A_27_47#_c_214_n N_VGND_c_438_n 0.0208843f $X=0.26 $Y=0.38 $X2=0 $Y2=0
cc_213 N_A_27_47#_M1002_g N_VGND_c_442_n 0.00506844f $X=2.685 $Y=0.7 $X2=0 $Y2=0
cc_214 N_A_27_47#_M1008_g N_VGND_c_442_n 0.00506844f $X=3.115 $Y=0.7 $X2=0 $Y2=0
cc_215 N_A_27_47#_M1006_s N_VGND_c_443_n 0.00215158f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_216 N_A_27_47#_M1002_g N_VGND_c_443_n 0.0095335f $X=2.685 $Y=0.7 $X2=0 $Y2=0
cc_217 N_A_27_47#_M1008_g N_VGND_c_443_n 0.0102494f $X=3.115 $Y=0.7 $X2=0 $Y2=0
cc_218 N_A_27_47#_c_214_n N_VGND_c_443_n 0.0125302f $X=0.26 $Y=0.38 $X2=0 $Y2=0
cc_219 N_A_27_47#_c_218_n N_VGND_c_443_n 0.00869588f $X=0.615 $Y=0.95 $X2=0
+ $Y2=0
cc_220 N_VPWR_c_319_n A_372_367# 0.00899413f $X=3.6 $Y=3.33 $X2=-0.19 $Y2=-0.245
cc_221 N_VPWR_c_319_n N_X_M1001_d 0.00536646f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_222 N_VPWR_c_324_n N_X_c_388_n 0.0124525f $X=3.395 $Y=3.33 $X2=0 $Y2=0
cc_223 N_VPWR_c_319_n N_X_c_388_n 0.00730901f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_224 N_VPWR_M1009_s X 0.00244921f $X=3.42 $Y=1.835 $X2=0 $Y2=0
cc_225 N_VPWR_M1009_s X 0.00983132f $X=3.42 $Y=1.835 $X2=0 $Y2=0
cc_226 N_VPWR_c_322_n X 0.00262043f $X=3.56 $Y=2.395 $X2=0 $Y2=0
cc_227 N_X_c_371_n N_VGND_c_435_n 0.0271735f $X=2.9 $Y=0.42 $X2=0 $Y2=0
cc_228 N_X_c_371_n N_VGND_c_437_n 0.021958f $X=2.9 $Y=0.42 $X2=0 $Y2=0
cc_229 X N_VGND_c_437_n 0.0153239f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_230 N_X_c_371_n N_VGND_c_442_n 0.0233446f $X=2.9 $Y=0.42 $X2=0 $Y2=0
cc_231 N_X_c_371_n N_VGND_c_443_n 0.0125323f $X=2.9 $Y=0.42 $X2=0 $Y2=0
cc_232 A_110_47# N_VGND_c_443_n 0.00467646f $X=0.55 $Y=0.235 $X2=1.615 $Y2=2.375
cc_233 N_A_182_47#_c_402_n N_VGND_M1004_s 0.00591634f $X=1.905 $Y=0.955
+ $X2=-0.19 $Y2=-0.245
cc_234 N_A_182_47#_c_401_n N_VGND_c_434_n 0.033111f $X=1.05 $Y=0.435 $X2=0 $Y2=0
cc_235 N_A_182_47#_c_402_n N_VGND_c_434_n 0.0220026f $X=1.905 $Y=0.955 $X2=0
+ $Y2=0
cc_236 N_A_182_47#_c_404_n N_VGND_c_434_n 0.0164958f $X=2 $Y=0.435 $X2=0 $Y2=0
cc_237 N_A_182_47#_c_404_n N_VGND_c_435_n 0.0220242f $X=2 $Y=0.435 $X2=0 $Y2=0
cc_238 N_A_182_47#_c_401_n N_VGND_c_438_n 0.0192086f $X=1.05 $Y=0.435 $X2=0
+ $Y2=0
cc_239 N_A_182_47#_c_404_n N_VGND_c_440_n 0.0168098f $X=2 $Y=0.435 $X2=0 $Y2=0
cc_240 N_A_182_47#_M1000_d N_VGND_c_443_n 0.00215591f $X=0.91 $Y=0.235 $X2=0
+ $Y2=0
cc_241 N_A_182_47#_c_401_n N_VGND_c_443_n 0.0124769f $X=1.05 $Y=0.435 $X2=0
+ $Y2=0
cc_242 N_A_182_47#_c_404_n N_VGND_c_443_n 0.00984755f $X=2 $Y=0.435 $X2=0 $Y2=0
