* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
X0 VGND A2 a_792_49# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X1 VPWR a_134_269# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X2 X a_134_269# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X3 VGND B1 a_134_269# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X4 a_792_49# A1 a_134_269# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X5 a_134_269# A1 a_792_49# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X6 VPWR A1 a_529_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X7 VGND a_134_269# X VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X8 a_134_269# B1 a_529_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X9 X a_134_269# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X10 a_529_367# B1 a_134_269# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X11 VGND a_134_269# X VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X12 a_134_269# B1 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X13 VPWR A2 a_529_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X14 a_529_367# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X15 a_529_367# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X16 X a_134_269# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X17 X a_134_269# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X18 VPWR a_134_269# X VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X19 a_792_49# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
.ends
