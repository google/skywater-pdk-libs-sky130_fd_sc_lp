* File: sky130_fd_sc_lp__mux2_8.pex.spice
* Created: Fri Aug 28 10:44:13 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__MUX2_8%A_84_21# 1 2 3 4 15 19 23 27 31 35 39 43 47
+ 51 55 59 63 67 71 75 77 84 86 87 90 92 96 103 104 105 108 109 112 113 114 115
+ 117 118 121 122
c288 117 0 1.88674e-19 $X=6.785 $Y=0.725
c289 108 0 1.4579e-20 $X=4.67 $Y=0.725
c290 86 0 1.83364e-19 $X=3.71 $Y=2.32
c291 71 0 3.40629e-19 $X=3.505 $Y=2.465
r292 134 135 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=3.505 $Y=1.43
+ $X2=3.575 $Y2=1.43
r293 133 134 62.9501 $w=3.3e-07 $l=3.6e-07 $layer=POLY_cond $X=3.145 $Y=1.43
+ $X2=3.505 $Y2=1.43
r294 132 133 12.2403 $w=3.3e-07 $l=7e-08 $layer=POLY_cond $X=3.075 $Y=1.43
+ $X2=3.145 $Y2=1.43
r295 131 132 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=2.645 $Y=1.43
+ $X2=3.075 $Y2=1.43
r296 130 131 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=2.215 $Y=1.43
+ $X2=2.645 $Y2=1.43
r297 129 130 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=1.785 $Y=1.43
+ $X2=2.215 $Y2=1.43
r298 128 129 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=1.355 $Y=1.43
+ $X2=1.785 $Y2=1.43
r299 124 126 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=0.495 $Y=1.43
+ $X2=0.925 $Y2=1.43
r300 121 122 8.48463 $w=2.98e-07 $l=1.65e-07 $layer=LI1_cond $X=6.855 $Y=2.585
+ $X2=6.69 $Y2=2.585
r301 117 118 9.26861 $w=2.18e-07 $l=1.65e-07 $layer=LI1_cond $X=6.785 $Y=0.745
+ $X2=6.62 $Y2=0.745
r302 115 122 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=5.86 $Y=2.52
+ $X2=6.69 $Y2=2.52
r303 114 115 9.42727 $w=1.98e-07 $l=1.7e-07 $layer=LI1_cond $X=5.69 $Y=2.505
+ $X2=5.86 $Y2=2.505
r304 113 114 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.02 $Y=2.49
+ $X2=5.69 $Y2=2.49
r305 111 113 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=4.855 $Y=2.57
+ $X2=5.02 $Y2=2.57
r306 111 112 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=4.855 $Y=2.57
+ $X2=4.69 $Y2=2.57
r307 109 118 105.69 $w=1.68e-07 $l=1.62e-06 $layer=LI1_cond $X=5 $Y=0.77
+ $X2=6.62 $Y2=0.77
r308 107 109 8.69362 $w=2.58e-07 $l=1.65e-07 $layer=LI1_cond $X=4.835 $Y=0.725
+ $X2=5 $Y2=0.725
r309 107 108 8.69362 $w=2.58e-07 $l=1.65e-07 $layer=LI1_cond $X=4.835 $Y=0.725
+ $X2=4.67 $Y2=0.725
r310 105 112 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=4.225 $Y=2.49
+ $X2=4.69 $Y2=2.49
r311 104 105 7.68295 $w=2.53e-07 $l=1.7e-07 $layer=LI1_cond $X=4.055 $Y=2.447
+ $X2=4.225 $Y2=2.447
r312 96 108 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=4.305 $Y=0.77
+ $X2=4.67 $Y2=0.77
r313 91 96 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.22 $Y=0.855
+ $X2=4.305 $Y2=0.77
r314 91 92 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=4.22 $Y=0.855
+ $X2=4.22 $Y2=1.265
r315 90 104 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=3.795 $Y=2.405
+ $X2=4.055 $Y2=2.405
r316 88 103 3.70735 $w=2.5e-07 $l=1.18427e-07 $layer=LI1_cond $X=3.795 $Y=1.35
+ $X2=3.71 $Y2=1.43
r317 87 92 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.135 $Y=1.35
+ $X2=4.22 $Y2=1.265
r318 87 88 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=4.135 $Y=1.35
+ $X2=3.795 $Y2=1.35
r319 86 90 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.71 $Y=2.32
+ $X2=3.795 $Y2=2.405
r320 85 103 2.76166 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.71 $Y=1.595
+ $X2=3.71 $Y2=1.43
r321 85 86 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=3.71 $Y=1.595
+ $X2=3.71 $Y2=2.32
r322 84 135 1.74861 $w=3.3e-07 $l=1e-08 $layer=POLY_cond $X=3.585 $Y=1.43
+ $X2=3.575 $Y2=1.43
r323 83 84 36.32 $w=1.7e-07 $l=6.8e-07 $layer=licon1_POLY $count=4 $X=3.585
+ $Y=1.43 $X2=3.585 $Y2=1.43
r324 80 128 26.2292 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=1.205 $Y=1.43
+ $X2=1.355 $Y2=1.43
r325 80 126 48.9612 $w=3.3e-07 $l=2.8e-07 $layer=POLY_cond $X=1.205 $Y=1.43
+ $X2=0.925 $Y2=1.43
r326 79 83 83.1156 $w=3.28e-07 $l=2.38e-06 $layer=LI1_cond $X=1.205 $Y=1.43
+ $X2=3.585 $Y2=1.43
r327 79 80 36.32 $w=1.7e-07 $l=6.8e-07 $layer=licon1_POLY $count=4 $X=1.205
+ $Y=1.43 $X2=1.205 $Y2=1.43
r328 77 103 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.625 $Y=1.43
+ $X2=3.71 $Y2=1.43
r329 77 83 1.3969 $w=3.28e-07 $l=4e-08 $layer=LI1_cond $X=3.625 $Y=1.43
+ $X2=3.585 $Y2=1.43
r330 73 135 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.575 $Y=1.265
+ $X2=3.575 $Y2=1.43
r331 73 75 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.575 $Y=1.265
+ $X2=3.575 $Y2=0.655
r332 69 134 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.505 $Y=1.595
+ $X2=3.505 $Y2=1.43
r333 69 71 446.106 $w=1.5e-07 $l=8.7e-07 $layer=POLY_cond $X=3.505 $Y=1.595
+ $X2=3.505 $Y2=2.465
r334 65 133 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.145 $Y=1.265
+ $X2=3.145 $Y2=1.43
r335 65 67 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=3.145 $Y=1.265
+ $X2=3.145 $Y2=0.655
r336 61 132 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.075 $Y=1.595
+ $X2=3.075 $Y2=1.43
r337 61 63 446.106 $w=1.5e-07 $l=8.7e-07 $layer=POLY_cond $X=3.075 $Y=1.595
+ $X2=3.075 $Y2=2.465
r338 57 131 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.645 $Y=1.595
+ $X2=2.645 $Y2=1.43
r339 57 59 446.106 $w=1.5e-07 $l=8.7e-07 $layer=POLY_cond $X=2.645 $Y=1.595
+ $X2=2.645 $Y2=2.465
r340 53 131 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.645 $Y=1.265
+ $X2=2.645 $Y2=1.43
r341 53 55 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.645 $Y=1.265
+ $X2=2.645 $Y2=0.655
r342 49 130 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.215 $Y=1.595
+ $X2=2.215 $Y2=1.43
r343 49 51 446.106 $w=1.5e-07 $l=8.7e-07 $layer=POLY_cond $X=2.215 $Y=1.595
+ $X2=2.215 $Y2=2.465
r344 45 130 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.215 $Y=1.265
+ $X2=2.215 $Y2=1.43
r345 45 47 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.215 $Y=1.265
+ $X2=2.215 $Y2=0.655
r346 41 129 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.785 $Y=1.595
+ $X2=1.785 $Y2=1.43
r347 41 43 446.106 $w=1.5e-07 $l=8.7e-07 $layer=POLY_cond $X=1.785 $Y=1.595
+ $X2=1.785 $Y2=2.465
r348 37 129 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.785 $Y=1.265
+ $X2=1.785 $Y2=1.43
r349 37 39 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.785 $Y=1.265
+ $X2=1.785 $Y2=0.655
r350 33 128 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.355 $Y=1.595
+ $X2=1.355 $Y2=1.43
r351 33 35 446.106 $w=1.5e-07 $l=8.7e-07 $layer=POLY_cond $X=1.355 $Y=1.595
+ $X2=1.355 $Y2=2.465
r352 29 128 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.355 $Y=1.265
+ $X2=1.355 $Y2=1.43
r353 29 31 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=1.355 $Y=1.265
+ $X2=1.355 $Y2=0.655
r354 25 126 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.925 $Y=1.595
+ $X2=0.925 $Y2=1.43
r355 25 27 446.106 $w=1.5e-07 $l=8.7e-07 $layer=POLY_cond $X=0.925 $Y=1.595
+ $X2=0.925 $Y2=2.465
r356 21 126 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.925 $Y=1.265
+ $X2=0.925 $Y2=1.43
r357 21 23 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=0.925 $Y=1.265
+ $X2=0.925 $Y2=0.655
r358 17 124 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=1.595
+ $X2=0.495 $Y2=1.43
r359 17 19 446.106 $w=1.5e-07 $l=8.7e-07 $layer=POLY_cond $X=0.495 $Y=1.595
+ $X2=0.495 $Y2=2.465
r360 13 124 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=1.265
+ $X2=0.495 $Y2=1.43
r361 13 15 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=0.495 $Y=1.265
+ $X2=0.495 $Y2=0.655
r362 4 121 600 $w=1.7e-07 $l=5.85662e-07 $layer=licon1_PDIFF $count=1 $X=6.645
+ $Y=2.095 $X2=6.855 $Y2=2.585
r363 3 111 600 $w=1.7e-07 $l=5.40486e-07 $layer=licon1_PDIFF $count=1 $X=4.715
+ $Y=2.095 $X2=4.855 $Y2=2.57
r364 2 117 182 $w=1.7e-07 $l=5.55608e-07 $layer=licon1_NDIFF $count=1 $X=6.645
+ $Y=0.235 $X2=6.785 $Y2=0.725
r365 1 107 182 $w=1.7e-07 $l=5.44977e-07 $layer=licon1_NDIFF $count=1 $X=4.625
+ $Y=0.235 $X2=4.835 $Y2=0.685
.ends

.subckt PM_SKY130_FD_SC_LP__MUX2_8%S 3 7 11 15 19 23 27 28 30 31 39 40 42 43 45
+ 46 48 54 55 67
c181 42 0 2.21293e-19 $X=7.775 $Y=2.035
c182 40 0 3.01138e-19 $X=8.205 $Y=1.51
c183 30 0 1.71596e-19 $X=5.355 $Y=2.15
c184 23 0 2.03815e-19 $X=8.125 $Y=2.465
c185 15 0 9.83241e-21 $X=5.57 $Y=2.595
c186 11 0 1.06565e-19 $X=5.55 $Y=0.555
c187 3 0 3.35634e-19 $X=4.12 $Y=0.555
r188 55 64 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=5.52 $Y=1.72
+ $X2=5.52 $Y2=2.035
r189 54 57 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.52 $Y=1.72
+ $X2=5.52 $Y2=1.885
r190 54 56 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.52 $Y=1.72
+ $X2=5.52 $Y2=1.555
r191 54 55 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.52
+ $Y=1.72 $X2=5.52 $Y2=1.72
r192 48 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=2.035
+ $X2=5.52 $Y2=2.035
r193 46 67 6.56993 $w=2.28e-07 $l=1.15e-07 $layer=LI1_cond $X=7.92 $Y=2.035
+ $X2=7.92 $Y2=1.92
r194 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=2.035
+ $X2=7.92 $Y2=2.035
r195 43 48 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.665 $Y=2.035
+ $X2=5.52 $Y2=2.035
r196 42 45 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.775 $Y=2.035
+ $X2=7.92 $Y2=2.035
r197 42 43 2.61138 $w=1.4e-07 $l=2.11e-06 $layer=MET1_cond $X=7.775 $Y=2.035
+ $X2=5.665 $Y2=2.035
r198 40 60 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.205 $Y=1.51
+ $X2=8.205 $Y2=1.675
r199 40 59 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=8.205 $Y=1.51
+ $X2=8.205 $Y2=1.345
r200 39 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.205
+ $Y=1.51 $X2=8.205 $Y2=1.51
r201 36 39 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=7.95 $Y=1.51
+ $X2=8.205 $Y2=1.51
r202 35 64 1.04768 $w=3.28e-07 $l=3e-08 $layer=LI1_cond $X=5.52 $Y=2.065
+ $X2=5.52 $Y2=2.035
r203 32 36 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.95 $Y=1.675
+ $X2=7.95 $Y2=1.51
r204 32 67 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=7.95 $Y=1.675
+ $X2=7.95 $Y2=1.92
r205 30 35 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.355 $Y=2.15
+ $X2=5.52 $Y2=2.065
r206 30 31 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=5.355 $Y=2.15
+ $X2=4.565 $Y2=2.15
r207 28 52 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.19 $Y=1.77
+ $X2=4.19 $Y2=1.935
r208 28 51 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.19 $Y=1.77
+ $X2=4.19 $Y2=1.605
r209 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.19
+ $Y=1.77 $X2=4.19 $Y2=1.77
r210 25 31 27.2595 $w=1.94e-07 $l=4.50988e-07 $layer=LI1_cond $X=4.135 $Y=2.107
+ $X2=4.565 $Y2=2.15
r211 25 27 7.11803 $w=3.38e-07 $l=2.1e-07 $layer=LI1_cond $X=4.135 $Y=1.98
+ $X2=4.135 $Y2=1.77
r212 23 60 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=8.125 $Y=2.465
+ $X2=8.125 $Y2=1.675
r213 19 59 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=8.115 $Y=0.655
+ $X2=8.115 $Y2=1.345
r214 15 57 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=5.57 $Y=2.595
+ $X2=5.57 $Y2=1.885
r215 11 56 512.766 $w=1.5e-07 $l=1e-06 $layer=POLY_cond $X=5.55 $Y=0.555
+ $X2=5.55 $Y2=1.555
r216 7 52 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=4.14 $Y=2.595
+ $X2=4.14 $Y2=1.935
r217 3 51 538.404 $w=1.5e-07 $l=1.05e-06 $layer=POLY_cond $X=4.12 $Y=0.555
+ $X2=4.12 $Y2=1.605
.ends

.subckt PM_SKY130_FD_SC_LP__MUX2_8%A1 3 5 9 13 17 21 22 26 30 31 34 36 41 51
c121 36 0 1.11688e-19 $X=6.48 $Y=1.665
c122 26 0 1.06565e-19 $X=4.64 $Y=1.19
r123 48 51 3.53416 $w=3.73e-07 $l=1.15e-07 $layer=LI1_cond $X=6.48 $Y=1.737
+ $X2=6.595 $Y2=1.737
r124 36 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=1.665
+ $X2=6.48 $Y2=1.665
r125 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=1.665
+ $X2=4.56 $Y2=1.665
r126 31 33 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.705 $Y=1.665
+ $X2=4.56 $Y2=1.665
r127 30 36 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.335 $Y=1.665
+ $X2=6.48 $Y2=1.665
r128 30 31 2.01732 $w=1.4e-07 $l=1.63e-06 $layer=MET1_cond $X=6.335 $Y=1.665
+ $X2=4.705 $Y2=1.665
r129 29 34 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=4.56 $Y=1.355
+ $X2=4.56 $Y2=1.665
r130 27 41 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.64 $Y=1.19
+ $X2=4.805 $Y2=1.19
r131 27 38 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=4.64 $Y=1.19 $X2=4.55
+ $Y2=1.19
r132 26 29 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=4.64 $Y=1.19
+ $X2=4.64 $Y2=1.355
r133 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.64
+ $Y=1.19 $X2=4.64 $Y2=1.19
r134 22 44 26.4627 $w=2.55e-07 $l=1.4e-07 $layer=POLY_cond $X=6.93 $Y=1.76
+ $X2=7.07 $Y2=1.76
r135 21 51 10.7241 $w=3.58e-07 $l=3.35e-07 $layer=LI1_cond $X=6.93 $Y=1.745
+ $X2=6.595 $Y2=1.745
r136 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.93
+ $Y=1.76 $X2=6.93 $Y2=1.76
r137 15 44 15.178 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.07 $Y=1.925
+ $X2=7.07 $Y2=1.76
r138 15 17 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=7.07 $Y=1.925
+ $X2=7.07 $Y2=2.595
r139 11 22 68.0471 $w=2.55e-07 $l=4.34741e-07 $layer=POLY_cond $X=6.57 $Y=1.925
+ $X2=6.93 $Y2=1.76
r140 11 13 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=6.57 $Y=1.925
+ $X2=6.57 $Y2=2.595
r141 7 9 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=5.05 $Y=1.025 $X2=5.05
+ $Y2=0.555
r142 5 7 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.975 $Y=1.1
+ $X2=5.05 $Y2=1.025
r143 5 41 87.1702 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=4.975 $Y=1.1
+ $X2=4.805 $Y2=1.1
r144 1 38 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.55 $Y=1.025
+ $X2=4.55 $Y2=1.19
r145 1 3 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=4.55 $Y=1.025 $X2=4.55
+ $Y2=0.555
.ends

.subckt PM_SKY130_FD_SC_LP__MUX2_8%A0 3 7 11 15 19 20 22 23 24 26 33 36
c102 36 0 1.91001e-19 $X=6.93 $Y=1.11
c103 22 0 9.83241e-21 $X=4.98 $Y=1.73
r104 34 36 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=6.93 $Y=1.19 $X2=6.93
+ $Y2=1.11
r105 33 35 13.5502 $w=2.49e-07 $l=7e-08 $layer=POLY_cond $X=6.93 $Y=1.19 $X2=7
+ $Y2=1.19
r106 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.93
+ $Y=1.19 $X2=6.93 $Y2=1.19
r107 26 34 3.66686 $w=3.28e-07 $l=1.05e-07 $layer=LI1_cond $X=6.93 $Y=1.295
+ $X2=6.93 $Y2=1.19
r108 23 30 17.2143 $w=2.52e-07 $l=9e-08 $layer=POLY_cond $X=4.98 $Y=1.73
+ $X2=5.07 $Y2=1.73
r109 22 24 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=4.98 $Y=1.73
+ $X2=4.98 $Y2=1.565
r110 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.98
+ $Y=1.73 $X2=4.98 $Y2=1.73
r111 19 36 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.765 $Y=1.11
+ $X2=6.93 $Y2=1.11
r112 19 20 105.69 $w=1.68e-07 $l=1.62e-06 $layer=LI1_cond $X=6.765 $Y=1.11
+ $X2=5.145 $Y2=1.11
r113 17 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.06 $Y=1.195
+ $X2=5.145 $Y2=1.11
r114 17 24 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=5.06 $Y=1.195
+ $X2=5.06 $Y2=1.565
r115 13 35 14.627 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7 $Y=1.025 $X2=7
+ $Y2=1.19
r116 13 15 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=7 $Y=1.025 $X2=7
+ $Y2=0.555
r117 9 33 69.6867 $w=2.49e-07 $l=4.34741e-07 $layer=POLY_cond $X=6.57 $Y=1.025
+ $X2=6.93 $Y2=1.19
r118 9 11 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=6.57 $Y=1.025 $X2=6.57
+ $Y2=0.555
r119 5 30 14.904 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.07 $Y=1.895
+ $X2=5.07 $Y2=1.73
r120 5 7 358.936 $w=1.5e-07 $l=7e-07 $layer=POLY_cond $X=5.07 $Y=1.895 $X2=5.07
+ $Y2=2.595
r121 1 23 65.0317 $w=2.52e-07 $l=4.14367e-07 $layer=POLY_cond $X=4.64 $Y=1.895
+ $X2=4.98 $Y2=1.73
r122 1 3 358.936 $w=1.5e-07 $l=7e-07 $layer=POLY_cond $X=4.64 $Y=1.895 $X2=4.64
+ $Y2=2.595
.ends

.subckt PM_SKY130_FD_SC_LP__MUX2_8%A_1179_311# 1 2 9 13 17 21 25 26 28 29 33 34
+ 36 37 40 44 49 50 51 52 56
c152 52 0 7.90956e-20 $X=7.45 $Y=2.18
c153 50 0 3.69886e-19 $X=7.53 $Y=1.35
c154 49 0 3.38857e-19 $X=7.53 $Y=1.35
c155 37 0 9.87261e-20 $X=7.695 $Y=1.09
c156 33 0 1.37914e-19 $X=7.45 $Y=2.095
c157 26 0 1.80337e-19 $X=6.06 $Y=1.72
c158 17 0 3.79675e-19 $X=7.5 $Y=0.555
c159 13 0 3.68162e-19 $X=6.14 $Y=2.595
c160 9 0 1.11688e-19 $X=6.14 $Y=0.555
r161 52 53 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=7.45 $Y=2.18
+ $X2=7.45 $Y2=2.405
r162 50 62 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.53 $Y=1.35
+ $X2=7.53 $Y2=1.515
r163 50 61 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=7.53 $Y=1.35
+ $X2=7.53 $Y2=1.185
r164 49 51 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=7.53 $Y=1.35
+ $X2=7.53 $Y2=1.515
r165 49 50 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.53
+ $Y=1.35 $X2=7.53 $Y2=1.35
r166 42 56 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=8.38 $Y=2.32
+ $X2=8.38 $Y2=2.405
r167 42 44 14.2903 $w=2.48e-07 $l=3.1e-07 $layer=LI1_cond $X=8.38 $Y=2.32
+ $X2=8.38 $Y2=2.01
r168 38 40 20.4297 $w=3.28e-07 $l=5.85e-07 $layer=LI1_cond $X=8.33 $Y=1.005
+ $X2=8.33 $Y2=0.42
r169 36 38 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=8.165 $Y=1.09
+ $X2=8.33 $Y2=1.005
r170 36 37 30.6631 $w=1.68e-07 $l=4.7e-07 $layer=LI1_cond $X=8.165 $Y=1.09
+ $X2=7.695 $Y2=1.09
r171 35 53 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.535 $Y=2.405
+ $X2=7.45 $Y2=2.405
r172 34 56 2.76166 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.255 $Y=2.405
+ $X2=8.38 $Y2=2.405
r173 34 35 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=8.255 $Y=2.405
+ $X2=7.535 $Y2=2.405
r174 33 52 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=7.45 $Y=2.095
+ $X2=7.45 $Y2=2.18
r175 33 51 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=7.45 $Y=2.095
+ $X2=7.45 $Y2=1.515
r176 30 37 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=7.53 $Y=1.175
+ $X2=7.695 $Y2=1.09
r177 30 49 6.11144 $w=3.28e-07 $l=1.75e-07 $layer=LI1_cond $X=7.53 $Y=1.175
+ $X2=7.53 $Y2=1.35
r178 28 52 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.365 $Y=2.18
+ $X2=7.45 $Y2=2.18
r179 28 29 76.984 $w=1.68e-07 $l=1.18e-06 $layer=LI1_cond $X=7.365 $Y=2.18
+ $X2=6.185 $Y2=2.18
r180 26 59 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.06 $Y=1.72
+ $X2=6.06 $Y2=1.885
r181 26 58 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.06 $Y=1.72
+ $X2=6.06 $Y2=1.555
r182 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.06
+ $Y=1.72 $X2=6.06 $Y2=1.72
r183 23 29 13.8237 $w=1.23e-07 $l=1.8262e-07 $layer=LI1_cond $X=6.04 $Y=2.095
+ $X2=6.185 $Y2=2.18
r184 23 25 14.9023 $w=2.88e-07 $l=3.75e-07 $layer=LI1_cond $X=6.04 $Y=2.095
+ $X2=6.04 $Y2=1.72
r185 21 62 553.787 $w=1.5e-07 $l=1.08e-06 $layer=POLY_cond $X=7.58 $Y=2.595
+ $X2=7.58 $Y2=1.515
r186 17 61 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=7.5 $Y=0.555
+ $X2=7.5 $Y2=1.185
r187 13 59 364.064 $w=1.5e-07 $l=7.1e-07 $layer=POLY_cond $X=6.14 $Y=2.595
+ $X2=6.14 $Y2=1.885
r188 9 58 512.766 $w=1.5e-07 $l=1e-06 $layer=POLY_cond $X=6.14 $Y=0.555 $X2=6.14
+ $Y2=1.555
r189 2 56 300 $w=1.7e-07 $l=6.91466e-07 $layer=licon1_PDIFF $count=2 $X=8.2
+ $Y=1.835 $X2=8.34 $Y2=2.46
r190 2 44 600 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_PDIFF $count=1 $X=8.2
+ $Y=1.835 $X2=8.34 $Y2=2.01
r191 1 40 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=8.19
+ $Y=0.235 $X2=8.33 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__MUX2_8%VPWR 1 2 3 4 5 6 7 22 24 30 34 38 40 44 48 52
+ 55 56 58 59 60 61 62 74 82 89 90 96 99 102
r143 102 103 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r144 99 100 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r145 96 97 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r146 93 94 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r147 90 103 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=8.4 $Y=3.33
+ $X2=7.92 $Y2=3.33
r148 89 90 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.4 $Y=3.33 $X2=8.4
+ $Y2=3.33
r149 87 102 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.075 $Y=3.33
+ $X2=7.91 $Y2=3.33
r150 87 89 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=8.075 $Y=3.33
+ $X2=8.4 $Y2=3.33
r151 86 103 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=7.92 $Y2=3.33
r152 86 100 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=6 $Y2=3.33
r153 85 86 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r154 83 99 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.02 $Y=3.33
+ $X2=5.855 $Y2=3.33
r155 83 85 92.6417 $w=1.68e-07 $l=1.42e-06 $layer=LI1_cond $X=6.02 $Y=3.33
+ $X2=7.44 $Y2=3.33
r156 82 102 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.745 $Y=3.33
+ $X2=7.91 $Y2=3.33
r157 82 85 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=7.745 $Y=3.33
+ $X2=7.44 $Y2=3.33
r158 81 100 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=6 $Y2=3.33
r159 80 81 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r160 78 97 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.6 $Y2=3.33
r161 77 80 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=4.08 $Y=3.33
+ $X2=5.52 $Y2=3.33
r162 77 78 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r163 75 96 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.885 $Y=3.33
+ $X2=3.72 $Y2=3.33
r164 75 77 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=3.885 $Y=3.33
+ $X2=4.08 $Y2=3.33
r165 74 99 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.69 $Y=3.33
+ $X2=5.855 $Y2=3.33
r166 74 80 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=5.69 $Y=3.33
+ $X2=5.52 $Y2=3.33
r167 73 97 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.6 $Y2=3.33
r168 72 73 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r169 70 73 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r170 69 70 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r171 67 70 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.68 $Y2=3.33
r172 67 94 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r173 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r174 64 93 4.00981 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=0.365 $Y=3.33
+ $X2=0.182 $Y2=3.33
r175 64 66 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=0.365 $Y=3.33
+ $X2=0.72 $Y2=3.33
r176 62 81 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=4.32 $Y=3.33
+ $X2=5.52 $Y2=3.33
r177 62 78 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.32 $Y=3.33
+ $X2=4.08 $Y2=3.33
r178 60 72 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=2.775 $Y=3.33
+ $X2=2.64 $Y2=3.33
r179 60 61 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.775 $Y=3.33
+ $X2=2.86 $Y2=3.33
r180 58 69 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=1.915 $Y=3.33
+ $X2=1.68 $Y2=3.33
r181 58 59 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.915 $Y=3.33 $X2=2
+ $Y2=3.33
r182 57 72 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=2.085 $Y=3.33
+ $X2=2.64 $Y2=3.33
r183 57 59 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.085 $Y=3.33 $X2=2
+ $Y2=3.33
r184 55 66 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.055 $Y=3.33
+ $X2=0.72 $Y2=3.33
r185 55 56 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.055 $Y=3.33
+ $X2=1.14 $Y2=3.33
r186 54 69 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=1.225 $Y=3.33
+ $X2=1.68 $Y2=3.33
r187 54 56 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.225 $Y=3.33
+ $X2=1.14 $Y2=3.33
r188 50 102 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.91 $Y=3.245
+ $X2=7.91 $Y2=3.33
r189 50 52 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=7.91 $Y=3.245
+ $X2=7.91 $Y2=2.885
r190 46 99 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.855 $Y=3.245
+ $X2=5.855 $Y2=3.33
r191 46 48 10.4768 $w=3.28e-07 $l=3e-07 $layer=LI1_cond $X=5.855 $Y=3.245
+ $X2=5.855 $Y2=2.945
r192 42 96 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.72 $Y=3.245
+ $X2=3.72 $Y2=3.33
r193 42 44 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=3.72 $Y=3.245
+ $X2=3.72 $Y2=2.885
r194 41 61 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.945 $Y=3.33
+ $X2=2.86 $Y2=3.33
r195 40 96 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.555 $Y=3.33
+ $X2=3.72 $Y2=3.33
r196 40 41 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=3.555 $Y=3.33
+ $X2=2.945 $Y2=3.33
r197 36 61 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.86 $Y=3.245
+ $X2=2.86 $Y2=3.33
r198 36 38 60.3476 $w=1.68e-07 $l=9.25e-07 $layer=LI1_cond $X=2.86 $Y=3.245
+ $X2=2.86 $Y2=2.32
r199 32 59 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2 $Y=3.245 $X2=2
+ $Y2=3.33
r200 32 34 60.3476 $w=1.68e-07 $l=9.25e-07 $layer=LI1_cond $X=2 $Y=3.245 $X2=2
+ $Y2=2.32
r201 28 56 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.14 $Y=3.245
+ $X2=1.14 $Y2=3.33
r202 28 30 60.3476 $w=1.68e-07 $l=9.25e-07 $layer=LI1_cond $X=1.14 $Y=3.245
+ $X2=1.14 $Y2=2.32
r203 24 27 45.6367 $w=2.48e-07 $l=9.9e-07 $layer=LI1_cond $X=0.24 $Y=1.96
+ $X2=0.24 $Y2=2.95
r204 22 93 3.13335 $w=2.5e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.24 $Y=3.245
+ $X2=0.182 $Y2=3.33
r205 22 27 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=0.24 $Y=3.245
+ $X2=0.24 $Y2=2.95
r206 7 52 600 $w=1.7e-07 $l=9.08598e-07 $layer=licon1_PDIFF $count=1 $X=7.655
+ $Y=2.095 $X2=7.91 $Y2=2.885
r207 6 48 600 $w=1.7e-07 $l=9.4921e-07 $layer=licon1_PDIFF $count=1 $X=5.645
+ $Y=2.095 $X2=5.855 $Y2=2.945
r208 5 44 600 $w=1.7e-07 $l=1.11781e-06 $layer=licon1_PDIFF $count=1 $X=3.58
+ $Y=1.835 $X2=3.72 $Y2=2.885
r209 4 38 300 $w=1.7e-07 $l=5.50568e-07 $layer=licon1_PDIFF $count=2 $X=2.72
+ $Y=1.835 $X2=2.86 $Y2=2.32
r210 3 34 300 $w=1.7e-07 $l=5.50568e-07 $layer=licon1_PDIFF $count=2 $X=1.86
+ $Y=1.835 $X2=2 $Y2=2.32
r211 2 30 300 $w=1.7e-07 $l=5.50568e-07 $layer=licon1_PDIFF $count=2 $X=1
+ $Y=1.835 $X2=1.14 $Y2=2.32
r212 1 27 400 $w=1.7e-07 $l=1.18528e-06 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.835 $X2=0.28 $Y2=2.95
r213 1 24 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.835 $X2=0.28 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_LP__MUX2_8%X 1 2 3 4 5 6 7 8 27 31 33 35 39 43 45 47 51
+ 55 57 59 61 63 67 70 73 74 76 77 79 82 83
c136 61 0 1.88359e-19 $X=3.25 $Y=1.985
r137 82 83 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.71 $Y=1.295
+ $X2=0.71 $Y2=1.665
r138 71 83 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=0.71 $Y=1.815
+ $X2=0.71 $Y2=1.665
r139 71 73 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.71 $Y=1.815
+ $X2=0.71 $Y2=1.9
r140 69 82 6.9845 $w=3.28e-07 $l=2e-07 $layer=LI1_cond $X=0.71 $Y=1.095 $X2=0.71
+ $Y2=1.295
r141 69 70 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.71 $Y=1.095
+ $X2=0.71 $Y2=1.01
r142 65 67 19.0328 $w=3.28e-07 $l=5.45e-07 $layer=LI1_cond $X=3.36 $Y=0.925
+ $X2=3.36 $Y2=0.38
r143 61 81 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.25 $Y=1.985
+ $X2=3.25 $Y2=1.9
r144 61 63 42.6404 $w=2.48e-07 $l=9.25e-07 $layer=LI1_cond $X=3.25 $Y=1.985
+ $X2=3.25 $Y2=2.91
r145 60 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.595 $Y=1.9
+ $X2=2.43 $Y2=1.9
r146 59 81 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.125 $Y=1.9
+ $X2=3.25 $Y2=1.9
r147 59 60 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=3.125 $Y=1.9
+ $X2=2.595 $Y2=1.9
r148 58 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.595 $Y=1.01
+ $X2=2.43 $Y2=1.01
r149 57 65 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.195 $Y=1.01
+ $X2=3.36 $Y2=0.925
r150 57 58 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=3.195 $Y=1.01
+ $X2=2.595 $Y2=1.01
r151 53 79 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.43 $Y=1.985
+ $X2=2.43 $Y2=1.9
r152 53 55 32.3033 $w=3.28e-07 $l=9.25e-07 $layer=LI1_cond $X=2.43 $Y=1.985
+ $X2=2.43 $Y2=2.91
r153 49 77 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.43 $Y=0.925
+ $X2=2.43 $Y2=1.01
r154 49 51 19.0328 $w=3.28e-07 $l=5.45e-07 $layer=LI1_cond $X=2.43 $Y=0.925
+ $X2=2.43 $Y2=0.38
r155 48 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.735 $Y=1.9
+ $X2=1.57 $Y2=1.9
r156 47 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.265 $Y=1.9
+ $X2=2.43 $Y2=1.9
r157 47 48 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=2.265 $Y=1.9
+ $X2=1.735 $Y2=1.9
r158 46 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.735 $Y=1.01
+ $X2=1.57 $Y2=1.01
r159 45 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.265 $Y=1.01
+ $X2=2.43 $Y2=1.01
r160 45 46 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=2.265 $Y=1.01
+ $X2=1.735 $Y2=1.01
r161 41 76 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.57 $Y=1.985
+ $X2=1.57 $Y2=1.9
r162 41 43 32.3033 $w=3.28e-07 $l=9.25e-07 $layer=LI1_cond $X=1.57 $Y=1.985
+ $X2=1.57 $Y2=2.91
r163 37 74 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.57 $Y=0.925
+ $X2=1.57 $Y2=1.01
r164 37 39 19.0328 $w=3.28e-07 $l=5.45e-07 $layer=LI1_cond $X=1.57 $Y=0.925
+ $X2=1.57 $Y2=0.38
r165 36 73 3.80956 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.875 $Y=1.9
+ $X2=0.71 $Y2=1.9
r166 35 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.405 $Y=1.9
+ $X2=1.57 $Y2=1.9
r167 35 36 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=1.405 $Y=1.9
+ $X2=0.875 $Y2=1.9
r168 34 70 3.80956 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.875 $Y=1.01
+ $X2=0.71 $Y2=1.01
r169 33 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.405 $Y=1.01
+ $X2=1.57 $Y2=1.01
r170 33 34 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=1.405 $Y=1.01
+ $X2=0.875 $Y2=1.01
r171 29 73 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.71 $Y=1.985
+ $X2=0.71 $Y2=1.9
r172 29 31 32.3033 $w=3.28e-07 $l=9.25e-07 $layer=LI1_cond $X=0.71 $Y=1.985
+ $X2=0.71 $Y2=2.91
r173 25 70 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.71 $Y=0.925
+ $X2=0.71 $Y2=1.01
r174 25 27 19.0328 $w=3.28e-07 $l=5.45e-07 $layer=LI1_cond $X=0.71 $Y=0.925
+ $X2=0.71 $Y2=0.38
r175 8 81 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=3.15
+ $Y=1.835 $X2=3.29 $Y2=1.98
r176 8 63 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=3.15
+ $Y=1.835 $X2=3.29 $Y2=2.91
r177 7 79 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.29
+ $Y=1.835 $X2=2.43 $Y2=1.98
r178 7 55 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=2.29
+ $Y=1.835 $X2=2.43 $Y2=2.91
r179 6 76 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.43
+ $Y=1.835 $X2=1.57 $Y2=1.98
r180 6 43 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=1.43
+ $Y=1.835 $X2=1.57 $Y2=2.91
r181 5 73 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.57
+ $Y=1.835 $X2=0.71 $Y2=1.98
r182 5 31 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=0.57
+ $Y=1.835 $X2=0.71 $Y2=2.91
r183 4 67 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.22
+ $Y=0.235 $X2=3.36 $Y2=0.38
r184 3 51 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.29
+ $Y=0.235 $X2=2.43 $Y2=0.38
r185 2 39 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.43
+ $Y=0.235 $X2=1.57 $Y2=0.38
r186 1 27 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=0.57
+ $Y=0.235 $X2=0.71 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_LP__MUX2_8%A_843_419# 1 2 7 10 15
c23 15 0 1.96566e-19 $X=5.355 $Y=2.91
r24 15 17 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=5.355 $Y=2.91 $X2=5.355
+ $Y2=2.99
r25 10 12 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=4.355 $Y=2.91 $X2=4.355
+ $Y2=2.99
r26 8 12 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.52 $Y=2.99
+ $X2=4.355 $Y2=2.99
r27 7 17 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.19 $Y=2.99
+ $X2=5.355 $Y2=2.99
r28 7 8 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.19 $Y=2.99 $X2=4.52
+ $Y2=2.99
r29 2 15 600 $w=1.7e-07 $l=9.13989e-07 $layer=licon1_PDIFF $count=1 $X=5.145
+ $Y=2.095 $X2=5.355 $Y2=2.91
r30 1 10 600 $w=1.7e-07 $l=8.82227e-07 $layer=licon1_PDIFF $count=1 $X=4.215
+ $Y=2.095 $X2=4.355 $Y2=2.91
.ends

.subckt PM_SKY130_FD_SC_LP__MUX2_8%A_1243_419# 1 2 7 10 15
c27 15 0 1.24719e-19 $X=7.355 $Y=2.865
r28 15 17 4.36531 $w=3.28e-07 $l=1.25e-07 $layer=LI1_cond $X=7.355 $Y=2.865
+ $X2=7.355 $Y2=2.99
r29 10 12 3.66686 $w=3.28e-07 $l=1.05e-07 $layer=LI1_cond $X=6.355 $Y=2.885
+ $X2=6.355 $Y2=2.99
r30 8 12 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.52 $Y=2.99
+ $X2=6.355 $Y2=2.99
r31 7 17 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.19 $Y=2.99
+ $X2=7.355 $Y2=2.99
r32 7 8 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=7.19 $Y=2.99 $X2=6.52
+ $Y2=2.99
r33 2 15 600 $w=1.7e-07 $l=8.68677e-07 $layer=licon1_PDIFF $count=1 $X=7.145
+ $Y=2.095 $X2=7.355 $Y2=2.865
r34 1 10 600 $w=1.7e-07 $l=8.57146e-07 $layer=licon1_PDIFF $count=1 $X=6.215
+ $Y=2.095 $X2=6.355 $Y2=2.885
.ends

.subckt PM_SKY130_FD_SC_LP__MUX2_8%VGND 1 2 3 4 5 6 7 22 24 28 32 36 40 46 50 53
+ 54 56 57 59 60 62 63 65 66 67 82 94 95 101
c127 82 0 1.4579e-20 $X=5.68 $Y=0
c128 50 0 1.45368e-19 $X=7.83 $Y=0.525
c129 7 0 9.87261e-20 $X=7.575 $Y=0.235
r130 101 102 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6 $Y=0 $X2=6
+ $Y2=0
r131 98 99 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r132 94 95 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.4 $Y=0 $X2=8.4
+ $Y2=0
r133 92 95 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.44 $Y=0 $X2=8.4
+ $Y2=0
r134 92 102 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=7.44 $Y=0 $X2=6
+ $Y2=0
r135 91 92 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=0 $X2=7.44
+ $Y2=0
r136 89 101 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.01 $Y=0
+ $X2=5.845 $Y2=0
r137 89 91 93.2941 $w=1.68e-07 $l=1.43e-06 $layer=LI1_cond $X=6.01 $Y=0 $X2=7.44
+ $Y2=0
r138 88 102 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=0 $X2=6
+ $Y2=0
r139 87 88 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r140 84 87 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=4.08 $Y=0 $X2=5.52
+ $Y2=0
r141 84 85 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r142 82 101 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.68 $Y=0
+ $X2=5.845 $Y2=0
r143 82 87 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=5.68 $Y=0 $X2=5.52
+ $Y2=0
r144 81 85 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r145 80 81 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r146 78 81 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.6
+ $Y2=0
r147 77 78 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r148 75 78 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r149 74 75 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r150 72 75 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r151 72 99 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=0.24
+ $Y2=0
r152 71 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r153 69 98 4.09637 $w=1.7e-07 $l=1.88e-07 $layer=LI1_cond $X=0.375 $Y=0
+ $X2=0.187 $Y2=0
r154 69 71 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.375 $Y=0 $X2=0.72
+ $Y2=0
r155 67 88 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=4.32 $Y=0 $X2=5.52
+ $Y2=0
r156 67 85 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=4.32 $Y=0
+ $X2=4.08 $Y2=0
r157 65 91 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=7.665 $Y=0
+ $X2=7.44 $Y2=0
r158 65 66 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.665 $Y=0 $X2=7.83
+ $Y2=0
r159 64 94 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=7.995 $Y=0 $X2=8.4
+ $Y2=0
r160 64 66 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.995 $Y=0 $X2=7.83
+ $Y2=0
r161 62 80 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=3.705 $Y=0 $X2=3.6
+ $Y2=0
r162 62 63 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.705 $Y=0 $X2=3.83
+ $Y2=0
r163 61 84 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=3.955 $Y=0
+ $X2=4.08 $Y2=0
r164 61 63 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.955 $Y=0 $X2=3.83
+ $Y2=0
r165 59 77 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=2.775 $Y=0
+ $X2=2.64 $Y2=0
r166 59 60 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.775 $Y=0 $X2=2.9
+ $Y2=0
r167 58 80 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=3.025 $Y=0 $X2=3.6
+ $Y2=0
r168 58 60 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.025 $Y=0 $X2=2.9
+ $Y2=0
r169 56 74 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=1.915 $Y=0
+ $X2=1.68 $Y2=0
r170 56 57 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.915 $Y=0 $X2=2
+ $Y2=0
r171 55 77 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=2.085 $Y=0
+ $X2=2.64 $Y2=0
r172 55 57 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.085 $Y=0 $X2=2
+ $Y2=0
r173 53 71 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.055 $Y=0
+ $X2=0.72 $Y2=0
r174 53 54 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.055 $Y=0 $X2=1.14
+ $Y2=0
r175 52 74 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=1.225 $Y=0
+ $X2=1.68 $Y2=0
r176 52 54 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.225 $Y=0 $X2=1.14
+ $Y2=0
r177 48 66 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.83 $Y=0.085
+ $X2=7.83 $Y2=0
r178 48 50 15.3659 $w=3.28e-07 $l=4.4e-07 $layer=LI1_cond $X=7.83 $Y=0.085
+ $X2=7.83 $Y2=0.525
r179 44 101 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.845 $Y=0.085
+ $X2=5.845 $Y2=0
r180 44 46 9.25447 $w=3.28e-07 $l=2.65e-07 $layer=LI1_cond $X=5.845 $Y=0.085
+ $X2=5.845 $Y2=0.35
r181 40 42 25.3537 $w=2.48e-07 $l=5.5e-07 $layer=LI1_cond $X=3.83 $Y=0.38
+ $X2=3.83 $Y2=0.93
r182 38 63 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.83 $Y=0.085
+ $X2=3.83 $Y2=0
r183 38 40 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=3.83 $Y=0.085
+ $X2=3.83 $Y2=0.38
r184 34 60 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.9 $Y=0.085
+ $X2=2.9 $Y2=0
r185 34 36 18.4391 $w=2.48e-07 $l=4e-07 $layer=LI1_cond $X=2.9 $Y=0.085 $X2=2.9
+ $Y2=0.485
r186 30 57 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2 $Y=0.085 $X2=2
+ $Y2=0
r187 30 32 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=2 $Y=0.085 $X2=2
+ $Y2=0.485
r188 26 54 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.14 $Y=0.085
+ $X2=1.14 $Y2=0
r189 26 28 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=1.14 $Y=0.085
+ $X2=1.14 $Y2=0.485
r190 22 98 3.11585 $w=2.6e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.245 $Y=0.085
+ $X2=0.187 $Y2=0
r191 22 24 12.1893 $w=2.58e-07 $l=2.75e-07 $layer=LI1_cond $X=0.245 $Y=0.085
+ $X2=0.245 $Y2=0.36
r192 7 50 182 $w=1.7e-07 $l=3.97555e-07 $layer=licon1_NDIFF $count=1 $X=7.575
+ $Y=0.235 $X2=7.83 $Y2=0.525
r193 6 46 182 $w=1.7e-07 $l=2.71477e-07 $layer=licon1_NDIFF $count=1 $X=5.625
+ $Y=0.235 $X2=5.845 $Y2=0.35
r194 5 42 182 $w=1.7e-07 $l=7.61791e-07 $layer=licon1_NDIFF $count=1 $X=3.65
+ $Y=0.235 $X2=3.79 $Y2=0.93
r195 5 40 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=3.65
+ $Y=0.235 $X2=3.79 $Y2=0.38
r196 4 36 182 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=1 $X=2.72
+ $Y=0.235 $X2=2.86 $Y2=0.485
r197 3 32 182 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=1 $X=1.86
+ $Y=0.235 $X2=2 $Y2=0.485
r198 2 28 182 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_NDIFF $count=1 $X=1
+ $Y=0.235 $X2=1.14 $Y2=0.485
r199 1 24 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.28 $Y2=0.36
.ends

.subckt PM_SKY130_FD_SC_LP__MUX2_8%A_839_47# 1 2 7 9 14
r26 14 17 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=5.335 $Y=0.34
+ $X2=5.335 $Y2=0.425
r27 9 12 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=4.335 $Y=0.34
+ $X2=4.335 $Y2=0.425
r28 8 9 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.5 $Y=0.34 $X2=4.335
+ $Y2=0.34
r29 7 14 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.17 $Y=0.34
+ $X2=5.335 $Y2=0.34
r30 7 8 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.17 $Y=0.34 $X2=4.5
+ $Y2=0.34
r31 2 17 182 $w=1.7e-07 $l=2.89828e-07 $layer=licon1_NDIFF $count=1 $X=5.125
+ $Y=0.235 $X2=5.335 $Y2=0.425
r32 1 12 182 $w=1.7e-07 $l=2.504e-07 $layer=licon1_NDIFF $count=1 $X=4.195
+ $Y=0.235 $X2=4.335 $Y2=0.425
.ends

.subckt PM_SKY130_FD_SC_LP__MUX2_8%A_1243_47# 1 2 7 11
c17 11 0 1.83562e-19 $X=7.285 $Y=0.465
r18 11 13 2.21818 $w=3.3e-07 $l=6e-08 $layer=LI1_cond $X=7.285 $Y=0.465
+ $X2=7.285 $Y2=0.525
r19 7 11 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=7.12 $Y=0.38
+ $X2=7.285 $Y2=0.465
r20 7 9 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=7.12 $Y=0.38
+ $X2=6.355 $Y2=0.38
r21 2 13 182 $w=1.7e-07 $l=3.80789e-07 $layer=licon1_NDIFF $count=1 $X=7.075
+ $Y=0.235 $X2=7.285 $Y2=0.525
r22 1 9 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=6.215
+ $Y=0.235 $X2=6.355 $Y2=0.38
.ends

