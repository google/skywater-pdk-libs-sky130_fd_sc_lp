* File: sky130_fd_sc_lp__o21a_m.pxi.spice
* Created: Fri Aug 28 11:04:22 2020
* 
x_PM_SKY130_FD_SC_LP__O21A_M%A_80_23# N_A_80_23#_M1006_s N_A_80_23#_M1005_d
+ N_A_80_23#_M1002_g N_A_80_23#_c_67_n N_A_80_23#_c_68_n N_A_80_23#_M1000_g
+ N_A_80_23#_c_69_n N_A_80_23#_c_77_n N_A_80_23#_c_70_n N_A_80_23#_c_71_n
+ N_A_80_23#_c_72_n N_A_80_23#_c_79_n N_A_80_23#_c_80_n N_A_80_23#_c_130_p
+ N_A_80_23#_c_81_n N_A_80_23#_c_73_n N_A_80_23#_c_87_p N_A_80_23#_c_74_n
+ PM_SKY130_FD_SC_LP__O21A_M%A_80_23#
x_PM_SKY130_FD_SC_LP__O21A_M%B1 N_B1_M1005_g N_B1_M1006_g N_B1_c_143_n
+ N_B1_c_148_n B1 B1 B1 N_B1_c_145_n PM_SKY130_FD_SC_LP__O21A_M%B1
x_PM_SKY130_FD_SC_LP__O21A_M%A2 N_A2_c_191_n N_A2_M1001_g N_A2_M1003_g
+ N_A2_c_197_n A2 A2 A2 A2 N_A2_c_194_n PM_SKY130_FD_SC_LP__O21A_M%A2
x_PM_SKY130_FD_SC_LP__O21A_M%A1 N_A1_M1007_g N_A1_c_246_n N_A1_M1004_g
+ N_A1_c_247_n N_A1_c_242_n N_A1_c_249_n A1 A1 A1 A1 N_A1_c_244_n
+ PM_SKY130_FD_SC_LP__O21A_M%A1
x_PM_SKY130_FD_SC_LP__O21A_M%X N_X_M1002_s N_X_M1000_s N_X_c_297_p X X X X X
+ N_X_c_280_n N_X_c_281_n PM_SKY130_FD_SC_LP__O21A_M%X
x_PM_SKY130_FD_SC_LP__O21A_M%VPWR N_VPWR_M1000_d N_VPWR_M1007_d N_VPWR_c_301_n
+ N_VPWR_c_302_n N_VPWR_c_303_n N_VPWR_c_304_n VPWR N_VPWR_c_305_n
+ N_VPWR_c_306_n N_VPWR_c_300_n N_VPWR_c_308_n PM_SKY130_FD_SC_LP__O21A_M%VPWR
x_PM_SKY130_FD_SC_LP__O21A_M%VGND N_VGND_M1002_d N_VGND_M1003_d N_VGND_c_338_n
+ N_VGND_c_339_n N_VGND_c_340_n N_VGND_c_341_n VGND N_VGND_c_342_n
+ N_VGND_c_343_n N_VGND_c_344_n N_VGND_c_345_n PM_SKY130_FD_SC_LP__O21A_M%VGND
x_PM_SKY130_FD_SC_LP__O21A_M%A_300_74# N_A_300_74#_M1006_d N_A_300_74#_M1004_d
+ N_A_300_74#_c_376_n N_A_300_74#_c_377_n N_A_300_74#_c_378_n
+ N_A_300_74#_c_379_n PM_SKY130_FD_SC_LP__O21A_M%A_300_74#
cc_1 VNB N_A_80_23#_c_67_n 0.0268581f $X=-0.19 $Y=-0.245 $X2=0.577 $Y2=1.268
cc_2 VNB N_A_80_23#_c_68_n 0.0103415f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.12
cc_3 VNB N_A_80_23#_c_69_n 0.0192174f $X=-0.19 $Y=-0.245 $X2=0.577 $Y2=1.445
cc_4 VNB N_A_80_23#_c_70_n 0.00154569f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=0.945
cc_5 VNB N_A_80_23#_c_71_n 0.00180608f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=2.3
cc_6 VNB N_A_80_23#_c_72_n 0.0187567f $X=-0.19 $Y=-0.245 $X2=1.105 $Y2=0.86
cc_7 VNB N_A_80_23#_c_73_n 0.0204383f $X=-0.19 $Y=-0.245 $X2=0.59 $Y2=0.94
cc_8 VNB N_A_80_23#_c_74_n 0.0232189f $X=-0.19 $Y=-0.245 $X2=0.577 $Y2=0.775
cc_9 VNB N_B1_M1006_g 0.0290885f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.775
cc_10 VNB N_B1_c_143_n 0.0217044f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.445
cc_11 VNB B1 0.00109817f $X=-0.19 $Y=-0.245 $X2=0.765 $Y2=2.27
cc_12 VNB N_B1_c_145_n 0.0469119f $X=-0.19 $Y=-0.245 $X2=0.765 $Y2=2.195
cc_13 VNB N_A2_c_191_n 0.00258793f $X=-0.19 $Y=-0.245 $X2=1.27 $Y2=2.675
cc_14 VNB N_A2_M1003_g 0.0448499f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.455
cc_15 VNB A2 0.00348555f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.445
cc_16 VNB N_A2_c_194_n 0.0211297f $X=-0.19 $Y=-0.245 $X2=0.765 $Y2=2.195
cc_17 VNB N_A1_M1004_g 0.0568884f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.455
cc_18 VNB N_A1_c_242_n 0.00576183f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB A1 0.0132304f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.195
cc_20 VNB N_A1_c_244_n 0.0214147f $X=-0.19 $Y=-0.245 $X2=0.675 $Y2=2.385
cc_21 VNB X 0.0463672f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.445
cc_22 VNB N_VPWR_c_300_n 0.123877f $X=-0.19 $Y=-0.245 $X2=1.21 $Y2=0.645
cc_23 VNB N_VGND_c_338_n 0.00528824f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.455
cc_24 VNB N_VGND_c_339_n 0.00856386f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.12
cc_25 VNB N_VGND_c_340_n 0.0346511f $X=-0.19 $Y=-0.245 $X2=0.765 $Y2=2.885
cc_26 VNB N_VGND_c_341_n 0.0040393f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_342_n 0.0188402f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_343_n 0.0233193f $X=-0.19 $Y=-0.245 $X2=1.21 $Y2=0.645
cc_29 VNB N_VGND_c_344_n 0.190795f $X=-0.19 $Y=-0.245 $X2=1.21 $Y2=0.645
cc_30 VNB N_VGND_c_345_n 0.00401211f $X=-0.19 $Y=-0.245 $X2=1.33 $Y2=2.715
cc_31 VNB N_A_300_74#_c_376_n 0.00116323f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.455
cc_32 VNB N_A_300_74#_c_377_n 0.0236651f $X=-0.19 $Y=-0.245 $X2=0.577 $Y2=1.268
cc_33 VNB N_A_300_74#_c_378_n 0.00408137f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.445
cc_34 VNB N_A_300_74#_c_379_n 0.00317049f $X=-0.19 $Y=-0.245 $X2=0.765 $Y2=2.885
cc_35 VPB N_A_80_23#_c_68_n 0.0250455f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.12
cc_36 VPB N_A_80_23#_M1000_g 0.0372179f $X=-0.19 $Y=1.655 $X2=0.765 $Y2=2.885
cc_37 VPB N_A_80_23#_c_77_n 0.0321014f $X=-0.19 $Y=1.655 $X2=0.765 $Y2=2.195
cc_38 VPB N_A_80_23#_c_71_n 0.00470958f $X=-0.19 $Y=1.655 $X2=0.59 $Y2=2.3
cc_39 VPB N_A_80_23#_c_79_n 0.015741f $X=-0.19 $Y=1.655 $X2=1.245 $Y2=2.385
cc_40 VPB N_A_80_23#_c_80_n 0.00335026f $X=-0.19 $Y=1.655 $X2=0.675 $Y2=2.385
cc_41 VPB N_A_80_23#_c_81_n 0.00185172f $X=-0.19 $Y=1.655 $X2=1.33 $Y2=2.715
cc_42 VPB N_B1_M1005_g 0.0504512f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_43 VPB N_B1_c_143_n 0.00457043f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=1.445
cc_44 VPB N_B1_c_148_n 0.0181926f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.12
cc_45 VPB B1 0.00517954f $X=-0.19 $Y=1.655 $X2=0.765 $Y2=2.27
cc_46 VPB N_A2_c_191_n 0.0193788f $X=-0.19 $Y=1.655 $X2=1.27 $Y2=2.675
cc_47 VPB N_A2_M1001_g 0.0396247f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_48 VPB N_A2_c_197_n 0.0240888f $X=-0.19 $Y=1.655 $X2=0.577 $Y2=1.268
cc_49 VPB A2 0.00494808f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=1.445
cc_50 VPB N_A1_M1007_g 0.0267076f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_51 VPB N_A1_c_246_n 0.0152473f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_52 VPB N_A1_c_247_n 0.0316874f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.12
cc_53 VPB N_A1_c_242_n 0.0272466f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_54 VPB N_A1_c_249_n 0.0233834f $X=-0.19 $Y=1.655 $X2=0.577 $Y2=1.445
cc_55 VPB A1 0.0241868f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.195
cc_56 VPB X 0.050701f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=1.445
cc_57 VPB N_X_c_280_n 0.0111747f $X=-0.19 $Y=1.655 $X2=0.59 $Y2=2.3
cc_58 VPB N_X_c_281_n 0.00459604f $X=-0.19 $Y=1.655 $X2=0.59 $Y2=0.94
cc_59 VPB N_VPWR_c_301_n 0.0047158f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=0.455
cc_60 VPB N_VPWR_c_302_n 0.01277f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.12
cc_61 VPB N_VPWR_c_303_n 0.0266906f $X=-0.19 $Y=1.655 $X2=0.765 $Y2=2.885
cc_62 VPB N_VPWR_c_304_n 0.0032427f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_63 VPB N_VPWR_c_305_n 0.0274415f $X=-0.19 $Y=1.655 $X2=0.59 $Y2=2.3
cc_64 VPB N_VPWR_c_306_n 0.0185316f $X=-0.19 $Y=1.655 $X2=1.21 $Y2=0.645
cc_65 VPB N_VPWR_c_300_n 0.0645924f $X=-0.19 $Y=1.655 $X2=1.21 $Y2=0.645
cc_66 VPB N_VPWR_c_308_n 0.00510247f $X=-0.19 $Y=1.655 $X2=1.33 $Y2=2.715
cc_67 N_A_80_23#_c_68_n N_B1_M1005_g 0.00224765f $X=0.475 $Y=2.12 $X2=0 $Y2=0
cc_68 N_A_80_23#_c_77_n N_B1_M1005_g 0.0359356f $X=0.765 $Y=2.195 $X2=0 $Y2=0
cc_69 N_A_80_23#_c_71_n N_B1_M1005_g 0.00169512f $X=0.59 $Y=2.3 $X2=0 $Y2=0
cc_70 N_A_80_23#_c_79_n N_B1_M1005_g 0.0106882f $X=1.245 $Y=2.385 $X2=0 $Y2=0
cc_71 N_A_80_23#_c_81_n N_B1_M1005_g 0.00579869f $X=1.33 $Y=2.715 $X2=0 $Y2=0
cc_72 N_A_80_23#_c_87_p N_B1_M1005_g 0.00308082f $X=1.41 $Y=2.82 $X2=0 $Y2=0
cc_73 N_A_80_23#_c_71_n N_B1_M1006_g 4.16161e-19 $X=0.59 $Y=2.3 $X2=0 $Y2=0
cc_74 N_A_80_23#_c_72_n N_B1_M1006_g 0.00204979f $X=1.105 $Y=0.86 $X2=0 $Y2=0
cc_75 N_A_80_23#_c_73_n N_B1_M1006_g 0.00414685f $X=0.59 $Y=0.94 $X2=0 $Y2=0
cc_76 N_A_80_23#_c_68_n N_B1_c_143_n 0.00828856f $X=0.475 $Y=2.12 $X2=0 $Y2=0
cc_77 N_A_80_23#_c_69_n N_B1_c_143_n 0.00680319f $X=0.577 $Y=1.445 $X2=0 $Y2=0
cc_78 N_A_80_23#_c_71_n N_B1_c_143_n 0.00467137f $X=0.59 $Y=2.3 $X2=0 $Y2=0
cc_79 N_A_80_23#_c_79_n N_B1_c_148_n 0.00376465f $X=1.245 $Y=2.385 $X2=0 $Y2=0
cc_80 N_A_80_23#_c_67_n B1 7.89849e-19 $X=0.577 $Y=1.268 $X2=0 $Y2=0
cc_81 N_A_80_23#_c_68_n B1 8.3035e-19 $X=0.475 $Y=2.12 $X2=0 $Y2=0
cc_82 N_A_80_23#_c_71_n B1 0.0361407f $X=0.59 $Y=2.3 $X2=0 $Y2=0
cc_83 N_A_80_23#_c_72_n B1 0.0135762f $X=1.105 $Y=0.86 $X2=0 $Y2=0
cc_84 N_A_80_23#_c_79_n B1 0.0170098f $X=1.245 $Y=2.385 $X2=0 $Y2=0
cc_85 N_A_80_23#_c_67_n N_B1_c_145_n 0.0127409f $X=0.577 $Y=1.268 $X2=0 $Y2=0
cc_86 N_A_80_23#_c_71_n N_B1_c_145_n 0.00171261f $X=0.59 $Y=2.3 $X2=0 $Y2=0
cc_87 N_A_80_23#_c_72_n N_B1_c_145_n 0.00903569f $X=1.105 $Y=0.86 $X2=0 $Y2=0
cc_88 N_A_80_23#_c_79_n N_A2_M1001_g 0.00119549f $X=1.245 $Y=2.385 $X2=0 $Y2=0
cc_89 N_A_80_23#_c_81_n N_A2_M1001_g 0.0048329f $X=1.33 $Y=2.715 $X2=0 $Y2=0
cc_90 N_A_80_23#_c_87_p N_A2_M1001_g 0.00495015f $X=1.41 $Y=2.82 $X2=0 $Y2=0
cc_91 N_A_80_23#_c_79_n A2 0.0133007f $X=1.245 $Y=2.385 $X2=0 $Y2=0
cc_92 N_A_80_23#_c_81_n A2 0.00135305f $X=1.33 $Y=2.715 $X2=0 $Y2=0
cc_93 N_A_80_23#_c_87_p N_A1_M1007_g 8.63638e-19 $X=1.41 $Y=2.82 $X2=0 $Y2=0
cc_94 N_A_80_23#_M1000_g X 0.0071049f $X=0.765 $Y=2.885 $X2=0 $Y2=0
cc_95 N_A_80_23#_c_70_n X 0.0130058f $X=0.59 $Y=0.945 $X2=0 $Y2=0
cc_96 N_A_80_23#_c_71_n X 0.0927453f $X=0.59 $Y=2.3 $X2=0 $Y2=0
cc_97 N_A_80_23#_c_80_n X 0.0137873f $X=0.675 $Y=2.385 $X2=0 $Y2=0
cc_98 N_A_80_23#_c_74_n X 0.0433027f $X=0.577 $Y=0.775 $X2=0 $Y2=0
cc_99 N_A_80_23#_M1000_g N_X_c_281_n 0.0034112f $X=0.765 $Y=2.885 $X2=0 $Y2=0
cc_100 N_A_80_23#_c_77_n N_X_c_281_n 0.00402094f $X=0.765 $Y=2.195 $X2=0 $Y2=0
cc_101 N_A_80_23#_c_79_n N_X_c_281_n 0.0015466f $X=1.245 $Y=2.385 $X2=0 $Y2=0
cc_102 N_A_80_23#_c_80_n N_X_c_281_n 0.00906707f $X=0.675 $Y=2.385 $X2=0 $Y2=0
cc_103 N_A_80_23#_c_87_p N_X_c_281_n 0.00213492f $X=1.41 $Y=2.82 $X2=0 $Y2=0
cc_104 N_A_80_23#_M1000_g N_VPWR_c_301_n 0.00271808f $X=0.765 $Y=2.885 $X2=0
+ $Y2=0
cc_105 N_A_80_23#_c_79_n N_VPWR_c_301_n 0.00803245f $X=1.245 $Y=2.385 $X2=0
+ $Y2=0
cc_106 N_A_80_23#_c_87_p N_VPWR_c_302_n 0.0026493f $X=1.41 $Y=2.82 $X2=0 $Y2=0
cc_107 N_A_80_23#_M1000_g N_VPWR_c_303_n 0.00552362f $X=0.765 $Y=2.885 $X2=0
+ $Y2=0
cc_108 N_A_80_23#_c_87_p N_VPWR_c_305_n 0.00910408f $X=1.41 $Y=2.82 $X2=0 $Y2=0
cc_109 N_A_80_23#_M1005_d N_VPWR_c_300_n 0.00246398f $X=1.27 $Y=2.675 $X2=0
+ $Y2=0
cc_110 N_A_80_23#_M1000_g N_VPWR_c_300_n 0.00743912f $X=0.765 $Y=2.885 $X2=0
+ $Y2=0
cc_111 N_A_80_23#_c_79_n N_VPWR_c_300_n 0.0111221f $X=1.245 $Y=2.385 $X2=0 $Y2=0
cc_112 N_A_80_23#_c_87_p N_VPWR_c_300_n 0.0110346f $X=1.41 $Y=2.82 $X2=0 $Y2=0
cc_113 N_A_80_23#_c_70_n N_VGND_c_338_n 0.00520877f $X=0.59 $Y=0.945 $X2=0 $Y2=0
cc_114 N_A_80_23#_c_72_n N_VGND_c_338_n 0.00738693f $X=1.105 $Y=0.86 $X2=0 $Y2=0
cc_115 N_A_80_23#_c_130_p N_VGND_c_338_n 0.00361546f $X=1.21 $Y=0.645 $X2=0
+ $Y2=0
cc_116 N_A_80_23#_c_73_n N_VGND_c_338_n 0.00267327f $X=0.59 $Y=0.94 $X2=0 $Y2=0
cc_117 N_A_80_23#_c_74_n N_VGND_c_338_n 0.00452011f $X=0.577 $Y=0.775 $X2=0
+ $Y2=0
cc_118 N_A_80_23#_c_130_p N_VGND_c_340_n 0.0054404f $X=1.21 $Y=0.645 $X2=0 $Y2=0
cc_119 N_A_80_23#_c_73_n N_VGND_c_342_n 2.43213e-19 $X=0.59 $Y=0.94 $X2=0 $Y2=0
cc_120 N_A_80_23#_c_74_n N_VGND_c_342_n 0.00575161f $X=0.577 $Y=0.775 $X2=0
+ $Y2=0
cc_121 N_A_80_23#_c_70_n N_VGND_c_344_n 0.00317739f $X=0.59 $Y=0.945 $X2=0 $Y2=0
cc_122 N_A_80_23#_c_72_n N_VGND_c_344_n 0.0118038f $X=1.105 $Y=0.86 $X2=0 $Y2=0
cc_123 N_A_80_23#_c_130_p N_VGND_c_344_n 0.00694949f $X=1.21 $Y=0.645 $X2=0
+ $Y2=0
cc_124 N_A_80_23#_c_74_n N_VGND_c_344_n 0.0114831f $X=0.577 $Y=0.775 $X2=0 $Y2=0
cc_125 N_A_80_23#_c_72_n N_A_300_74#_c_376_n 0.00489317f $X=1.105 $Y=0.86 $X2=0
+ $Y2=0
cc_126 N_A_80_23#_c_72_n N_A_300_74#_c_378_n 0.00662791f $X=1.105 $Y=0.86 $X2=0
+ $Y2=0
cc_127 N_B1_M1005_g N_A2_c_191_n 0.0439817f $X=1.195 $Y=2.885 $X2=0 $Y2=0
cc_128 N_B1_c_148_n N_A2_c_191_n 0.0119216f $X=1.145 $Y=1.88 $X2=0 $Y2=0
cc_129 B1 N_A2_c_191_n 0.00161332f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_130 N_B1_M1006_g N_A2_M1003_g 0.0275538f $X=1.425 $Y=0.58 $X2=0 $Y2=0
cc_131 B1 N_A2_M1003_g 2.12013e-19 $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_132 N_B1_c_145_n N_A2_M1003_g 0.00517758f $X=1.145 $Y=1.375 $X2=0 $Y2=0
cc_133 N_B1_M1005_g A2 0.00149892f $X=1.195 $Y=2.885 $X2=0 $Y2=0
cc_134 N_B1_c_143_n A2 0.00156959f $X=1.145 $Y=1.715 $X2=0 $Y2=0
cc_135 B1 A2 0.0412593f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_136 N_B1_c_145_n A2 0.00180458f $X=1.145 $Y=1.375 $X2=0 $Y2=0
cc_137 N_B1_c_143_n N_A2_c_194_n 0.0119216f $X=1.145 $Y=1.715 $X2=0 $Y2=0
cc_138 B1 N_A2_c_194_n 0.00168046f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_139 N_B1_M1005_g N_VPWR_c_301_n 0.00271808f $X=1.195 $Y=2.885 $X2=0 $Y2=0
cc_140 N_B1_M1005_g N_VPWR_c_305_n 0.00552362f $X=1.195 $Y=2.885 $X2=0 $Y2=0
cc_141 N_B1_M1005_g N_VPWR_c_300_n 0.00625534f $X=1.195 $Y=2.885 $X2=0 $Y2=0
cc_142 N_B1_M1006_g N_VGND_c_338_n 0.00540096f $X=1.425 $Y=0.58 $X2=0 $Y2=0
cc_143 N_B1_M1006_g N_VGND_c_340_n 0.00461464f $X=1.425 $Y=0.58 $X2=0 $Y2=0
cc_144 N_B1_M1006_g N_VGND_c_344_n 0.00914415f $X=1.425 $Y=0.58 $X2=0 $Y2=0
cc_145 N_B1_M1006_g N_A_300_74#_c_376_n 5.67457e-19 $X=1.425 $Y=0.58 $X2=0 $Y2=0
cc_146 N_B1_M1006_g N_A_300_74#_c_378_n 0.00356175f $X=1.425 $Y=0.58 $X2=0 $Y2=0
cc_147 N_A2_M1001_g N_A1_c_246_n 0.00510169f $X=1.625 $Y=2.885 $X2=0 $Y2=0
cc_148 A2 N_A1_c_246_n 7.73432e-19 $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_149 N_A2_M1003_g N_A1_M1004_g 0.036501f $X=1.855 $Y=0.58 $X2=0 $Y2=0
cc_150 N_A2_M1001_g N_A1_c_247_n 0.0555149f $X=1.625 $Y=2.885 $X2=0 $Y2=0
cc_151 N_A2_c_197_n N_A1_c_247_n 0.00148092f $X=1.74 $Y=2.1 $X2=0 $Y2=0
cc_152 A2 N_A1_c_247_n 0.00114637f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_153 N_A2_c_191_n N_A1_c_242_n 0.0118047f $X=1.74 $Y=1.91 $X2=0 $Y2=0
cc_154 N_A2_c_197_n N_A1_c_249_n 0.0118047f $X=1.74 $Y=2.1 $X2=0 $Y2=0
cc_155 N_A2_M1001_g A1 9.68589e-19 $X=1.625 $Y=2.885 $X2=0 $Y2=0
cc_156 N_A2_M1003_g A1 0.00702457f $X=1.855 $Y=0.58 $X2=0 $Y2=0
cc_157 A2 A1 0.0695948f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_158 A2 N_A1_c_244_n 6.12233e-19 $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_159 N_A2_c_194_n N_A1_c_244_n 0.0118047f $X=1.715 $Y=1.595 $X2=0 $Y2=0
cc_160 N_A2_M1001_g N_VPWR_c_302_n 0.0022041f $X=1.625 $Y=2.885 $X2=0 $Y2=0
cc_161 N_A2_M1001_g N_VPWR_c_305_n 0.00552362f $X=1.625 $Y=2.885 $X2=0 $Y2=0
cc_162 N_A2_M1001_g N_VPWR_c_300_n 0.00684977f $X=1.625 $Y=2.885 $X2=0 $Y2=0
cc_163 A2 N_VPWR_c_300_n 0.00720306f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_164 N_A2_M1003_g N_VGND_c_339_n 0.00327258f $X=1.855 $Y=0.58 $X2=0 $Y2=0
cc_165 N_A2_M1003_g N_VGND_c_340_n 0.00461464f $X=1.855 $Y=0.58 $X2=0 $Y2=0
cc_166 N_A2_M1003_g N_VGND_c_344_n 0.00468324f $X=1.855 $Y=0.58 $X2=0 $Y2=0
cc_167 N_A2_M1003_g N_A_300_74#_c_376_n 9.4709e-19 $X=1.855 $Y=0.58 $X2=0 $Y2=0
cc_168 N_A2_M1003_g N_A_300_74#_c_377_n 0.0155156f $X=1.855 $Y=0.58 $X2=0 $Y2=0
cc_169 A2 N_A_300_74#_c_377_n 0.00418441f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_170 A2 N_A_300_74#_c_378_n 0.0131935f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_171 N_A2_c_194_n N_A_300_74#_c_378_n 0.00238471f $X=1.715 $Y=1.595 $X2=0
+ $Y2=0
cc_172 N_A1_M1007_g N_VPWR_c_302_n 0.0111975f $X=1.985 $Y=2.885 $X2=0 $Y2=0
cc_173 N_A1_c_247_n N_VPWR_c_302_n 0.00153758f $X=2.245 $Y=2.415 $X2=0 $Y2=0
cc_174 A1 N_VPWR_c_302_n 0.0116602f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_175 N_A1_M1007_g N_VPWR_c_305_n 0.00486043f $X=1.985 $Y=2.885 $X2=0 $Y2=0
cc_176 N_A1_M1007_g N_VPWR_c_300_n 0.00818711f $X=1.985 $Y=2.885 $X2=0 $Y2=0
cc_177 A1 N_VPWR_c_300_n 0.00356679f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_178 N_A1_M1004_g N_VGND_c_339_n 0.00327258f $X=2.285 $Y=0.58 $X2=0 $Y2=0
cc_179 N_A1_M1004_g N_VGND_c_343_n 0.00461464f $X=2.285 $Y=0.58 $X2=0 $Y2=0
cc_180 N_A1_M1004_g N_VGND_c_344_n 0.0047218f $X=2.285 $Y=0.58 $X2=0 $Y2=0
cc_181 N_A1_M1004_g N_A_300_74#_c_377_n 0.0132026f $X=2.285 $Y=0.58 $X2=0 $Y2=0
cc_182 A1 N_A_300_74#_c_377_n 0.026708f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_183 N_A1_c_244_n N_A_300_74#_c_377_n 0.00337939f $X=2.335 $Y=1.595 $X2=0
+ $Y2=0
cc_184 N_A1_M1004_g N_A_300_74#_c_379_n 0.0020107f $X=2.285 $Y=0.58 $X2=0 $Y2=0
cc_185 N_X_c_280_n N_VPWR_c_303_n 0.00617311f $X=0.24 $Y=2.715 $X2=0 $Y2=0
cc_186 N_X_c_281_n N_VPWR_c_303_n 0.0119708f $X=0.55 $Y=2.82 $X2=0 $Y2=0
cc_187 N_X_M1000_s N_VPWR_c_300_n 0.00236056f $X=0.425 $Y=2.675 $X2=0 $Y2=0
cc_188 N_X_c_280_n N_VPWR_c_300_n 0.00605229f $X=0.24 $Y=2.715 $X2=0 $Y2=0
cc_189 N_X_c_281_n N_VPWR_c_300_n 0.0132152f $X=0.55 $Y=2.82 $X2=0 $Y2=0
cc_190 N_X_c_297_p N_VGND_c_342_n 0.012998f $X=0.26 $Y=0.43 $X2=0 $Y2=0
cc_191 N_X_M1002_s N_VGND_c_344_n 0.00407306f $X=0.135 $Y=0.245 $X2=0 $Y2=0
cc_192 N_X_c_297_p N_VGND_c_344_n 0.0080203f $X=0.26 $Y=0.43 $X2=0 $Y2=0
cc_193 N_VPWR_c_300_n A_340_535# 0.00620535f $X=2.64 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_194 N_VGND_c_340_n N_A_300_74#_c_376_n 0.00523228f $X=1.965 $Y=0 $X2=0 $Y2=0
cc_195 N_VGND_c_344_n N_A_300_74#_c_376_n 0.00699584f $X=2.64 $Y=0 $X2=0 $Y2=0
cc_196 N_VGND_c_339_n N_A_300_74#_c_377_n 0.0142847f $X=2.07 $Y=0.515 $X2=0
+ $Y2=0
cc_197 N_VGND_c_344_n N_A_300_74#_c_377_n 0.0135041f $X=2.64 $Y=0 $X2=0 $Y2=0
cc_198 N_VGND_c_343_n N_A_300_74#_c_379_n 0.00549876f $X=2.64 $Y=0 $X2=0 $Y2=0
cc_199 N_VGND_c_344_n N_A_300_74#_c_379_n 0.00699584f $X=2.64 $Y=0 $X2=0 $Y2=0
