* File: sky130_fd_sc_lp__a211o_4.pex.spice
* Created: Wed Sep  2 09:17:39 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__A211O_4%A_103_263# 1 2 3 4 15 19 23 27 31 35 39 43
+ 45 54 56 57 58 60 63 65 69 71 75 77 79 83 84 87 99
c166 79 0 1.81713e-19 $X=3.095 $Y=0.93
c167 60 0 1.93692e-19 $X=2.645 $Y=2.12
r168 96 97 21.8577 $w=3.3e-07 $l=1.25e-07 $layer=POLY_cond $X=1.88 $Y=1.48
+ $X2=2.005 $Y2=1.48
r169 95 96 53.3327 $w=3.3e-07 $l=3.05e-07 $layer=POLY_cond $X=1.575 $Y=1.48
+ $X2=1.88 $Y2=1.48
r170 94 95 21.8577 $w=3.3e-07 $l=1.25e-07 $layer=POLY_cond $X=1.45 $Y=1.48
+ $X2=1.575 $Y2=1.48
r171 93 94 53.3327 $w=3.3e-07 $l=3.05e-07 $layer=POLY_cond $X=1.145 $Y=1.48
+ $X2=1.45 $Y2=1.48
r172 92 93 21.8577 $w=3.3e-07 $l=1.25e-07 $layer=POLY_cond $X=1.02 $Y=1.48
+ $X2=1.145 $Y2=1.48
r173 87 88 11.7205 $w=2.29e-07 $l=2.2e-07 $layer=LI1_cond $X=3.992 $Y=0.93
+ $X2=3.992 $Y2=1.15
r174 83 84 9.26861 $w=2.18e-07 $l=1.65e-07 $layer=LI1_cond $X=3.62 $Y=2.145
+ $X2=3.455 $Y2=2.145
r175 73 75 17.8038 $w=1.88e-07 $l=3.05e-07 $layer=LI1_cond $X=5.6 $Y=1.065
+ $X2=5.6 $Y2=0.76
r176 72 88 2.48377 $w=1.7e-07 $l=1.18e-07 $layer=LI1_cond $X=4.11 $Y=1.15
+ $X2=3.992 $Y2=1.15
r177 71 73 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=5.505 $Y=1.15
+ $X2=5.6 $Y2=1.065
r178 71 72 91.0107 $w=1.68e-07 $l=1.395e-06 $layer=LI1_cond $X=5.505 $Y=1.15
+ $X2=4.11 $Y2=1.15
r179 67 87 4.41277 $w=2.35e-07 $l=8.5e-08 $layer=LI1_cond $X=3.992 $Y=0.845
+ $X2=3.992 $Y2=0.93
r180 67 69 20.8421 $w=2.33e-07 $l=4.25e-07 $layer=LI1_cond $X=3.992 $Y=0.845
+ $X2=3.992 $Y2=0.42
r181 66 79 1.83547 $w=1.7e-07 $l=1.03e-07 $layer=LI1_cond $X=3.205 $Y=0.93
+ $X2=3.102 $Y2=0.93
r182 65 87 2.48377 $w=1.7e-07 $l=1.17e-07 $layer=LI1_cond $X=3.875 $Y=0.93
+ $X2=3.992 $Y2=0.93
r183 65 66 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.875 $Y=0.93
+ $X2=3.205 $Y2=0.93
r184 61 79 4.59867 $w=2.03e-07 $l=8.5e-08 $layer=LI1_cond $X=3.102 $Y=0.845
+ $X2=3.102 $Y2=0.93
r185 61 63 22.9933 $w=2.03e-07 $l=4.25e-07 $layer=LI1_cond $X=3.102 $Y=0.845
+ $X2=3.102 $Y2=0.42
r186 60 84 52.8449 $w=1.68e-07 $l=8.1e-07 $layer=LI1_cond $X=2.645 $Y=2.12
+ $X2=3.455 $Y2=2.12
r187 57 79 7.57428 $w=2.03e-07 $l=1.4e-07 $layer=LI1_cond $X=3.102 $Y=1.07
+ $X2=3.102 $Y2=0.93
r188 57 58 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=3 $Y=1.07
+ $X2=2.645 $Y2=1.07
r189 56 60 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.56 $Y=2.035
+ $X2=2.645 $Y2=2.12
r190 55 77 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.56 $Y=1.585
+ $X2=2.56 $Y2=1.49
r191 55 56 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=2.56 $Y=1.585
+ $X2=2.56 $Y2=2.035
r192 54 77 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.56 $Y=1.395
+ $X2=2.56 $Y2=1.49
r193 53 58 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.56 $Y=1.155
+ $X2=2.645 $Y2=1.07
r194 53 54 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=2.56 $Y=1.155
+ $X2=2.56 $Y2=1.395
r195 52 99 71.6931 $w=3.3e-07 $l=4.1e-07 $layer=POLY_cond $X=2.04 $Y=1.48
+ $X2=2.45 $Y2=1.48
r196 52 97 6.12014 $w=3.3e-07 $l=3.5e-08 $layer=POLY_cond $X=2.04 $Y=1.48
+ $X2=2.005 $Y2=1.48
r197 51 52 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=2.04
+ $Y=1.48 $X2=2.04 $Y2=1.48
r198 48 92 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.68 $Y=1.48
+ $X2=1.02 $Y2=1.48
r199 48 89 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=0.68 $Y=1.48 $X2=0.59
+ $Y2=1.48
r200 47 51 79.3876 $w=1.88e-07 $l=1.36e-06 $layer=LI1_cond $X=0.68 $Y=1.49
+ $X2=2.04 $Y2=1.49
r201 47 48 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=0.68
+ $Y=1.48 $X2=0.68 $Y2=1.48
r202 45 77 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=2.475 $Y=1.49
+ $X2=2.56 $Y2=1.49
r203 45 51 25.3923 $w=1.88e-07 $l=4.35e-07 $layer=LI1_cond $X=2.475 $Y=1.49
+ $X2=2.04 $Y2=1.49
r204 41 99 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.45 $Y=1.315
+ $X2=2.45 $Y2=1.48
r205 41 43 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.45 $Y=1.315
+ $X2=2.45 $Y2=0.655
r206 37 97 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.005 $Y=1.315
+ $X2=2.005 $Y2=1.48
r207 37 39 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=2.005 $Y=1.315
+ $X2=2.005 $Y2=0.655
r208 33 96 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.88 $Y=1.645
+ $X2=1.88 $Y2=1.48
r209 33 35 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=1.88 $Y=1.645
+ $X2=1.88 $Y2=2.465
r210 29 95 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.575 $Y=1.315
+ $X2=1.575 $Y2=1.48
r211 29 31 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.575 $Y=1.315
+ $X2=1.575 $Y2=0.655
r212 25 94 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.45 $Y=1.645
+ $X2=1.45 $Y2=1.48
r213 25 27 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=1.45 $Y=1.645
+ $X2=1.45 $Y2=2.465
r214 21 93 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.145 $Y=1.315
+ $X2=1.145 $Y2=1.48
r215 21 23 338.426 $w=1.5e-07 $l=6.6e-07 $layer=POLY_cond $X=1.145 $Y=1.315
+ $X2=1.145 $Y2=0.655
r216 17 92 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.02 $Y=1.645
+ $X2=1.02 $Y2=1.48
r217 17 19 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=1.02 $Y=1.645
+ $X2=1.02 $Y2=2.465
r218 13 89 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.59 $Y=1.645
+ $X2=0.59 $Y2=1.48
r219 13 15 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=0.59 $Y=1.645
+ $X2=0.59 $Y2=2.465
r220 4 83 600 $w=1.7e-07 $l=3.78583e-07 $layer=licon1_PDIFF $count=1 $X=3.48
+ $Y=1.835 $X2=3.62 $Y2=2.15
r221 3 75 182 $w=1.7e-07 $l=5.90868e-07 $layer=licon1_NDIFF $count=1 $X=5.46
+ $Y=0.235 $X2=5.6 $Y2=0.76
r222 2 87 182 $w=1.7e-07 $l=7.61791e-07 $layer=licon1_NDIFF $count=1 $X=3.83
+ $Y=0.235 $X2=3.97 $Y2=0.93
r223 2 69 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=3.83
+ $Y=0.235 $X2=3.97 $Y2=0.42
r224 1 79 182 $w=1.7e-07 $l=7.61791e-07 $layer=licon1_NDIFF $count=1 $X=2.955
+ $Y=0.235 $X2=3.095 $Y2=0.93
r225 1 63 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=2.955
+ $Y=0.235 $X2=3.095 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__A211O_4%B1 3 7 11 13 15 18 22 24 28 29
c100 28 0 1.39441e-19 $X=2.9 $Y=1.51
c101 3 0 1.81713e-19 $X=2.88 $Y=0.655
r102 28 31 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.9 $Y=1.51
+ $X2=2.9 $Y2=1.675
r103 28 30 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.9 $Y=1.51
+ $X2=2.9 $Y2=1.345
r104 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.9
+ $Y=1.51 $X2=2.9 $Y2=1.51
r105 24 39 3.39823 $w=3.88e-07 $l=1.15e-07 $layer=LI1_cond $X=3.01 $Y=1.665
+ $X2=3.01 $Y2=1.78
r106 24 39 5.6248 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=3.205 $Y=1.78
+ $X2=3.01 $Y2=1.78
r107 24 29 4.58022 $w=3.88e-07 $l=1.55e-07 $layer=LI1_cond $X=3.01 $Y=1.665
+ $X2=3.01 $Y2=1.51
r108 22 24 47.5816 $w=2.23e-07 $l=9.15e-07 $layer=LI1_cond $X=4.12 $Y=1.78
+ $X2=3.205 $Y2=1.78
r109 21 22 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.285 $Y=1.78
+ $X2=4.12 $Y2=1.78
r110 18 21 9.7783 $w=3.28e-07 $l=2.8e-07 $layer=LI1_cond $X=4.285 $Y=1.5
+ $X2=4.285 $Y2=1.78
r111 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.285
+ $Y=1.5 $X2=4.285 $Y2=1.5
r112 13 19 38.6069 $w=3.31e-07 $l=1.77059e-07 $layer=POLY_cond $X=4.305 $Y=1.665
+ $X2=4.28 $Y2=1.5
r113 13 15 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=4.305 $Y=1.665
+ $X2=4.305 $Y2=2.465
r114 9 19 38.6069 $w=3.31e-07 $l=2.07123e-07 $layer=POLY_cond $X=4.185 $Y=1.335
+ $X2=4.28 $Y2=1.5
r115 9 11 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=4.185 $Y=1.335
+ $X2=4.185 $Y2=0.655
r116 7 31 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.975 $Y=2.465
+ $X2=2.975 $Y2=1.675
r117 3 30 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.88 $Y=0.655
+ $X2=2.88 $Y2=1.345
.ends

.subckt PM_SKY130_FD_SC_LP__A211O_4%C1 1 3 6 8 10 13 15 22
c57 15 0 1.39441e-19 $X=3.6 $Y=1.295
r58 20 22 20.0833 $w=3.24e-07 $l=1.35e-07 $layer=POLY_cond $X=3.62 $Y=1.332
+ $X2=3.755 $Y2=1.332
r59 18 20 31.9846 $w=3.24e-07 $l=2.15e-07 $layer=POLY_cond $X=3.405 $Y=1.332
+ $X2=3.62 $Y2=1.332
r60 17 18 11.9012 $w=3.24e-07 $l=8e-08 $layer=POLY_cond $X=3.325 $Y=1.332
+ $X2=3.405 $Y2=1.332
r61 15 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.62
+ $Y=1.35 $X2=3.62 $Y2=1.35
r62 11 22 11.9012 $w=3.24e-07 $l=2.19383e-07 $layer=POLY_cond $X=3.835 $Y=1.515
+ $X2=3.755 $Y2=1.332
r63 11 13 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=3.835 $Y=1.515
+ $X2=3.835 $Y2=2.465
r64 8 22 20.7868 $w=1.5e-07 $l=1.82e-07 $layer=POLY_cond $X=3.755 $Y=1.15
+ $X2=3.755 $Y2=1.332
r65 8 10 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=3.755 $Y=1.15
+ $X2=3.755 $Y2=0.655
r66 4 18 20.7868 $w=1.5e-07 $l=1.83e-07 $layer=POLY_cond $X=3.405 $Y=1.515
+ $X2=3.405 $Y2=1.332
r67 4 6 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=3.405 $Y=1.515
+ $X2=3.405 $Y2=2.465
r68 1 17 20.7868 $w=1.5e-07 $l=1.82e-07 $layer=POLY_cond $X=3.325 $Y=1.15
+ $X2=3.325 $Y2=1.332
r69 1 3 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=3.325 $Y=1.15
+ $X2=3.325 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__A211O_4%A2 3 6 10 14 20 21 23 24 25 33 36
c76 36 0 5.4009e-20 $X=4.935 $Y=1.725
c77 21 0 1.55473e-19 $X=6.335 $Y=1.51
r78 33 36 54.9546 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=4.935 $Y=1.51
+ $X2=4.935 $Y2=1.725
r79 33 35 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.935 $Y=1.51
+ $X2=4.935 $Y2=1.345
r80 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.935
+ $Y=1.51 $X2=4.935 $Y2=1.51
r81 24 25 16.2679 $w=3.38e-07 $l=3.95e-07 $layer=LI1_cond $X=5.52 $Y=2.035
+ $X2=5.915 $Y2=2.035
r82 23 41 3.50848 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.935 $Y=2.035
+ $X2=5.1 $Y2=2.035
r83 23 34 23.4615 $w=2.73e-07 $l=5.25e-07 $layer=LI1_cond $X=4.935 $Y=2.035
+ $X2=4.935 $Y2=1.51
r84 23 24 26.6182 $w=1.68e-07 $l=4.08e-07 $layer=LI1_cond $X=5.112 $Y=2.035
+ $X2=5.52 $Y2=2.035
r85 23 41 0.782888 $w=1.68e-07 $l=1.2e-08 $layer=LI1_cond $X=5.112 $Y=2.035
+ $X2=5.1 $Y2=2.035
r86 21 39 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.335 $Y=1.51
+ $X2=6.335 $Y2=1.675
r87 21 38 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=6.335 $Y=1.51
+ $X2=6.335 $Y2=1.345
r88 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.335
+ $Y=1.51 $X2=6.335 $Y2=1.51
r89 17 25 10.547 $w=3.78e-07 $l=3.05e-07 $layer=LI1_cond $X=6.02 $Y=1.645
+ $X2=6.02 $Y2=1.95
r90 16 20 12.1007 $w=2.98e-07 $l=3.15e-07 $layer=LI1_cond $X=6.02 $Y=1.495
+ $X2=6.335 $Y2=1.495
r91 16 17 2.82627 $w=2.1e-07 $l=1.5e-07 $layer=LI1_cond $X=6.02 $Y=1.495
+ $X2=6.02 $Y2=1.645
r92 14 39 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=6.245 $Y=2.465
+ $X2=6.245 $Y2=1.675
r93 10 38 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=6.245 $Y=0.655
+ $X2=6.245 $Y2=1.345
r94 6 35 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=4.955 $Y=0.655
+ $X2=4.955 $Y2=1.345
r95 3 36 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=4.845 $Y=2.465
+ $X2=4.845 $Y2=1.725
.ends

.subckt PM_SKY130_FD_SC_LP__A211O_4%A1 3 7 11 15 17 23 24
c49 23 0 2.09482e-19 $X=5.475 $Y=1.51
r50 22 24 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=5.475 $Y=1.51
+ $X2=5.815 $Y2=1.51
r51 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.475
+ $Y=1.51 $X2=5.475 $Y2=1.51
r52 19 22 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=5.385 $Y=1.51
+ $X2=5.475 $Y2=1.51
r53 17 23 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=5.475 $Y=1.665
+ $X2=5.475 $Y2=1.51
r54 13 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.815 $Y=1.675
+ $X2=5.815 $Y2=1.51
r55 13 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=5.815 $Y=1.675
+ $X2=5.815 $Y2=2.465
r56 9 24 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.815 $Y=1.345
+ $X2=5.815 $Y2=1.51
r57 9 11 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=5.815 $Y=1.345
+ $X2=5.815 $Y2=0.655
r58 5 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.385 $Y=1.675
+ $X2=5.385 $Y2=1.51
r59 5 7 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=5.385 $Y=1.675
+ $X2=5.385 $Y2=2.465
r60 1 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.385 $Y=1.345
+ $X2=5.385 $Y2=1.51
r61 1 3 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=5.385 $Y=1.345
+ $X2=5.385 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__A211O_4%VPWR 1 2 3 4 5 16 18 24 30 36 40 42 44 49 54
+ 62 69 70 76 79 82 85
r103 85 86 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r104 82 83 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r105 79 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r106 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r107 73 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r108 70 86 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6.48 $Y=3.33 $X2=6
+ $Y2=3.33
r109 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r110 67 85 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.195 $Y=3.33
+ $X2=6.03 $Y2=3.33
r111 67 69 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=6.195 $Y=3.33
+ $X2=6.48 $Y2=3.33
r112 66 86 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33 $X2=6
+ $Y2=3.33
r113 66 83 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.52 $Y=3.33
+ $X2=5.04 $Y2=3.33
r114 65 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r115 63 82 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.225 $Y=3.33
+ $X2=5.06 $Y2=3.33
r116 63 65 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=5.225 $Y=3.33
+ $X2=5.52 $Y2=3.33
r117 62 85 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.865 $Y=3.33
+ $X2=6.03 $Y2=3.33
r118 62 65 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=5.865 $Y=3.33
+ $X2=5.52 $Y2=3.33
r119 61 83 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.04 $Y2=3.33
r120 60 61 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r121 58 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=2.16 $Y2=3.33
r122 57 60 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=2.64 $Y=3.33
+ $X2=4.56 $Y2=3.33
r123 57 58 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r124 55 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.26 $Y=3.33
+ $X2=2.095 $Y2=3.33
r125 55 57 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=2.26 $Y=3.33
+ $X2=2.64 $Y2=3.33
r126 54 82 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.895 $Y=3.33
+ $X2=5.06 $Y2=3.33
r127 54 60 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=4.895 $Y=3.33
+ $X2=4.56 $Y2=3.33
r128 53 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.16 $Y2=3.33
r129 53 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r130 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r131 50 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.4 $Y=3.33
+ $X2=1.235 $Y2=3.33
r132 50 52 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=1.4 $Y=3.33
+ $X2=1.68 $Y2=3.33
r133 49 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.93 $Y=3.33
+ $X2=2.095 $Y2=3.33
r134 49 52 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=1.93 $Y=3.33
+ $X2=1.68 $Y2=3.33
r135 48 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r136 48 74 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r137 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r138 45 73 4.55841 $w=1.7e-07 $l=2.7e-07 $layer=LI1_cond $X=0.54 $Y=3.33
+ $X2=0.27 $Y2=3.33
r139 45 47 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=0.54 $Y=3.33
+ $X2=0.72 $Y2=3.33
r140 44 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.07 $Y=3.33
+ $X2=1.235 $Y2=3.33
r141 44 47 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=1.07 $Y=3.33
+ $X2=0.72 $Y2=3.33
r142 42 61 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=3.36 $Y=3.33
+ $X2=4.56 $Y2=3.33
r143 42 58 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=3.36 $Y=3.33
+ $X2=2.64 $Y2=3.33
r144 38 85 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.03 $Y=3.245
+ $X2=6.03 $Y2=3.33
r145 38 40 16.0644 $w=3.28e-07 $l=4.6e-07 $layer=LI1_cond $X=6.03 $Y=3.245
+ $X2=6.03 $Y2=2.785
r146 34 82 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.06 $Y=3.245
+ $X2=5.06 $Y2=3.33
r147 34 36 16.5882 $w=3.28e-07 $l=4.75e-07 $layer=LI1_cond $X=5.06 $Y=3.245
+ $X2=5.06 $Y2=2.77
r148 30 33 33.8748 $w=3.28e-07 $l=9.7e-07 $layer=LI1_cond $X=2.095 $Y=1.98
+ $X2=2.095 $Y2=2.95
r149 28 79 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.095 $Y=3.245
+ $X2=2.095 $Y2=3.33
r150 28 33 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.095 $Y=3.245
+ $X2=2.095 $Y2=2.95
r151 24 27 26.5411 $w=3.28e-07 $l=7.6e-07 $layer=LI1_cond $X=1.235 $Y=2.19
+ $X2=1.235 $Y2=2.95
r152 22 76 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.235 $Y=3.245
+ $X2=1.235 $Y2=3.33
r153 22 27 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.235 $Y=3.245
+ $X2=1.235 $Y2=2.95
r154 18 21 26.8903 $w=3.28e-07 $l=7.7e-07 $layer=LI1_cond $X=0.375 $Y=2.18
+ $X2=0.375 $Y2=2.95
r155 16 73 3.20777 $w=3.3e-07 $l=1.41244e-07 $layer=LI1_cond $X=0.375 $Y=3.245
+ $X2=0.27 $Y2=3.33
r156 16 21 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.375 $Y=3.245
+ $X2=0.375 $Y2=2.95
r157 5 40 600 $w=1.7e-07 $l=1.0176e-06 $layer=licon1_PDIFF $count=1 $X=5.89
+ $Y=1.835 $X2=6.03 $Y2=2.785
r158 4 36 600 $w=1.7e-07 $l=1.00256e-06 $layer=licon1_PDIFF $count=1 $X=4.92
+ $Y=1.835 $X2=5.06 $Y2=2.77
r159 3 33 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=1.955
+ $Y=1.835 $X2=2.095 $Y2=2.95
r160 3 30 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.955
+ $Y=1.835 $X2=2.095 $Y2=1.98
r161 2 27 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=1.095
+ $Y=1.835 $X2=1.235 $Y2=2.95
r162 2 24 400 $w=1.7e-07 $l=4.19196e-07 $layer=licon1_PDIFF $count=1 $X=1.095
+ $Y=1.835 $X2=1.235 $Y2=2.19
r163 1 21 400 $w=1.7e-07 $l=1.17584e-06 $layer=licon1_PDIFF $count=1 $X=0.25
+ $Y=1.835 $X2=0.375 $Y2=2.95
r164 1 18 400 $w=1.7e-07 $l=4.02679e-07 $layer=licon1_PDIFF $count=1 $X=0.25
+ $Y=1.835 $X2=0.375 $Y2=2.18
.ends

.subckt PM_SKY130_FD_SC_LP__A211O_4%X 1 2 3 4 13 14 15 19 23 27 29 33 39 42 43
+ 44 45 46 47 61
r64 59 61 3.16357 $w=2.53e-07 $l=7e-08 $layer=LI1_cond $X=0.217 $Y=1.225
+ $X2=0.217 $Y2=1.295
r65 46 53 3.29812 $w=2.85e-07 $l=8.5e-08 $layer=LI1_cond $X=0.247 $Y=1.14
+ $X2=0.247 $Y2=1.055
r66 46 59 3.29812 $w=2.85e-07 $l=9.88686e-08 $layer=LI1_cond $X=0.247 $Y=1.14
+ $X2=0.217 $Y2=1.225
r67 46 47 16.4054 $w=2.53e-07 $l=3.63e-07 $layer=LI1_cond $X=0.217 $Y=1.302
+ $X2=0.217 $Y2=1.665
r68 46 61 0.316357 $w=2.53e-07 $l=7e-09 $layer=LI1_cond $X=0.217 $Y=1.302
+ $X2=0.217 $Y2=1.295
r69 45 53 4.75611 $w=3.13e-07 $l=1.3e-07 $layer=LI1_cond $X=0.247 $Y=0.925
+ $X2=0.247 $Y2=1.055
r70 44 45 13.5366 $w=3.13e-07 $l=3.7e-07 $layer=LI1_cond $X=0.247 $Y=0.555
+ $X2=0.247 $Y2=0.925
r71 41 47 4.06745 $w=2.53e-07 $l=9e-08 $layer=LI1_cond $X=0.217 $Y=1.755
+ $X2=0.217 $Y2=1.665
r72 37 39 38.5101 $w=1.78e-07 $l=6.25e-07 $layer=LI1_cond $X=2.215 $Y=1.045
+ $X2=2.215 $Y2=0.42
r73 33 35 54.2871 $w=1.88e-07 $l=9.3e-07 $layer=LI1_cond $X=1.665 $Y=1.98
+ $X2=1.665 $Y2=2.91
r74 31 33 3.21053 $w=1.88e-07 $l=5.5e-08 $layer=LI1_cond $X=1.665 $Y=1.925
+ $X2=1.665 $Y2=1.98
r75 30 43 5.52892 $w=1.75e-07 $l=9.5e-08 $layer=LI1_cond $X=1.455 $Y=1.135
+ $X2=1.36 $Y2=1.135
r76 29 37 6.81649 $w=1.8e-07 $l=1.27279e-07 $layer=LI1_cond $X=2.125 $Y=1.135
+ $X2=2.215 $Y2=1.045
r77 29 30 41.2828 $w=1.78e-07 $l=6.7e-07 $layer=LI1_cond $X=2.125 $Y=1.135
+ $X2=1.455 $Y2=1.135
r78 25 43 1.04816 $w=1.9e-07 $l=9e-08 $layer=LI1_cond $X=1.36 $Y=1.045 $X2=1.36
+ $Y2=1.135
r79 25 27 36.4833 $w=1.88e-07 $l=6.25e-07 $layer=LI1_cond $X=1.36 $Y=1.045
+ $X2=1.36 $Y2=0.42
r80 24 42 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=0.9 $Y=1.84 $X2=0.805
+ $Y2=1.84
r81 23 31 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=1.57 $Y=1.84
+ $X2=1.665 $Y2=1.925
r82 23 24 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.57 $Y=1.84 $X2=0.9
+ $Y2=1.84
r83 19 21 54.2871 $w=1.88e-07 $l=9.3e-07 $layer=LI1_cond $X=0.805 $Y=1.98
+ $X2=0.805 $Y2=2.91
r84 17 42 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=0.805 $Y=1.925
+ $X2=0.805 $Y2=1.84
r85 17 19 3.21053 $w=1.88e-07 $l=5.5e-08 $layer=LI1_cond $X=0.805 $Y=1.925
+ $X2=0.805 $Y2=1.98
r86 16 46 3.25423 $w=1.7e-07 $l=1.58e-07 $layer=LI1_cond $X=0.405 $Y=1.14
+ $X2=0.247 $Y2=1.14
r87 15 43 5.52892 $w=1.75e-07 $l=9.74679e-08 $layer=LI1_cond $X=1.265 $Y=1.14
+ $X2=1.36 $Y2=1.135
r88 15 16 56.107 $w=1.68e-07 $l=8.6e-07 $layer=LI1_cond $X=1.265 $Y=1.14
+ $X2=0.405 $Y2=1.14
r89 14 41 7.17723 $w=1.7e-07 $l=1.65118e-07 $layer=LI1_cond $X=0.345 $Y=1.84
+ $X2=0.217 $Y2=1.755
r90 13 42 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=0.71 $Y=1.84
+ $X2=0.805 $Y2=1.84
r91 13 14 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.71 $Y=1.84
+ $X2=0.345 $Y2=1.84
r92 4 35 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=1.525
+ $Y=1.835 $X2=1.665 $Y2=2.91
r93 4 33 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.525
+ $Y=1.835 $X2=1.665 $Y2=1.98
r94 3 21 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=0.665
+ $Y=1.835 $X2=0.805 $Y2=2.91
r95 3 19 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.665
+ $Y=1.835 $X2=0.805 $Y2=1.98
r96 2 39 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=2.08
+ $Y=0.235 $X2=2.22 $Y2=0.42
r97 1 27 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=1.22
+ $Y=0.235 $X2=1.36 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__A211O_4%A_527_367# 1 2 3 4 15 17 19 21 25 27 31 36
+ 41 43
c71 1 0 1.93692e-19 $X=2.635 $Y=1.835
r72 39 40 4.41555 $w=3.73e-07 $l=1.35e-07 $layer=LI1_cond $X=4.542 $Y=2.375
+ $X2=4.542 $Y2=2.51
r73 38 39 8.34048 $w=3.73e-07 $l=2.55e-07 $layer=LI1_cond $X=4.542 $Y=2.12
+ $X2=4.542 $Y2=2.375
r74 29 43 3.19717 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=6.46 $Y=2.29
+ $X2=6.46 $Y2=2.375
r75 29 31 10.826 $w=3.28e-07 $l=3.1e-07 $layer=LI1_cond $X=6.46 $Y=2.29 $X2=6.46
+ $Y2=1.98
r76 28 41 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=5.695 $Y=2.375
+ $X2=5.565 $Y2=2.375
r77 27 43 3.3845 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.295 $Y=2.375
+ $X2=6.46 $Y2=2.375
r78 27 28 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=6.295 $Y=2.375
+ $X2=5.695 $Y2=2.375
r79 23 41 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=5.565 $Y=2.46
+ $X2=5.565 $Y2=2.375
r80 23 25 0.221624 $w=2.58e-07 $l=5e-09 $layer=LI1_cond $X=5.565 $Y=2.46
+ $X2=5.565 $Y2=2.465
r81 22 39 5.35566 $w=1.7e-07 $l=1.88e-07 $layer=LI1_cond $X=4.73 $Y=2.375
+ $X2=4.542 $Y2=2.375
r82 21 41 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=5.435 $Y=2.375
+ $X2=5.565 $Y2=2.375
r83 21 22 45.9947 $w=1.68e-07 $l=7.05e-07 $layer=LI1_cond $X=5.435 $Y=2.375
+ $X2=4.73 $Y2=2.375
r84 17 40 2.89929 $w=3.73e-07 $l=9.12688e-08 $layer=LI1_cond $X=4.555 $Y=2.595
+ $X2=4.542 $Y2=2.51
r85 17 19 10.677 $w=3.38e-07 $l=3.15e-07 $layer=LI1_cond $X=4.555 $Y=2.595
+ $X2=4.555 $Y2=2.91
r86 16 36 4.09051 $w=1.7e-07 $l=1.77059e-07 $layer=LI1_cond $X=2.925 $Y=2.51
+ $X2=2.76 $Y2=2.485
r87 15 40 5.35566 $w=1.7e-07 $l=1.87e-07 $layer=LI1_cond $X=4.355 $Y=2.51
+ $X2=4.542 $Y2=2.51
r88 15 16 93.2941 $w=1.68e-07 $l=1.43e-06 $layer=LI1_cond $X=4.355 $Y=2.51
+ $X2=2.925 $Y2=2.51
r89 4 43 300 $w=1.7e-07 $l=6.56277e-07 $layer=licon1_PDIFF $count=2 $X=6.32
+ $Y=1.835 $X2=6.46 $Y2=2.425
r90 4 31 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=6.32
+ $Y=1.835 $X2=6.46 $Y2=1.98
r91 3 25 300 $w=1.7e-07 $l=6.96491e-07 $layer=licon1_PDIFF $count=2 $X=5.46
+ $Y=1.835 $X2=5.6 $Y2=2.465
r92 2 38 300 $w=1.7e-07 $l=3.65992e-07 $layer=licon1_PDIFF $count=2 $X=4.38
+ $Y=1.835 $X2=4.565 $Y2=2.12
r93 2 19 600 $w=1.7e-07 $l=1.16383e-06 $layer=licon1_PDIFF $count=1 $X=4.38
+ $Y=1.835 $X2=4.565 $Y2=2.91
r94 1 36 300 $w=1.7e-07 $l=7.64951e-07 $layer=licon1_PDIFF $count=2 $X=2.635
+ $Y=1.835 $X2=2.76 $Y2=2.54
.ends

.subckt PM_SKY130_FD_SC_LP__A211O_4%A_610_367# 1 2 11
r16 8 11 34.1759 $w=2.88e-07 $l=8.6e-07 $layer=LI1_cond $X=3.19 $Y=2.91 $X2=4.05
+ $Y2=2.91
r17 2 11 600 $w=1.7e-07 $l=1.12282e-06 $layer=licon1_PDIFF $count=1 $X=3.91
+ $Y=1.835 $X2=4.05 $Y2=2.89
r18 1 8 600 $w=1.7e-07 $l=1.12282e-06 $layer=licon1_PDIFF $count=1 $X=3.05
+ $Y=1.835 $X2=3.19 $Y2=2.89
.ends

.subckt PM_SKY130_FD_SC_LP__A211O_4%VGND 1 2 3 4 5 6 21 23 27 31 35 39 41 43 45
+ 46 47 53 58 63 68 77 80 83 86 90
r101 89 90 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=0 $X2=6.48
+ $Y2=0
r102 86 87 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r103 83 84 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r104 80 81 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r105 77 78 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r106 75 90 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=6.48
+ $Y2=0
r107 74 75 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6 $Y2=0
r108 72 75 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=6
+ $Y2=0
r109 72 87 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=4.56
+ $Y2=0
r110 71 74 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=5.04 $Y=0 $X2=6
+ $Y2=0
r111 71 72 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r112 69 86 12.0118 $w=1.7e-07 $l=2.78e-07 $layer=LI1_cond $X=4.835 $Y=0
+ $X2=4.557 $Y2=0
r113 69 71 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=4.835 $Y=0
+ $X2=5.04 $Y2=0
r114 68 89 4.13127 $w=1.7e-07 $l=1.77e-07 $layer=LI1_cond $X=6.365 $Y=0
+ $X2=6.542 $Y2=0
r115 68 74 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=6.365 $Y=0 $X2=6
+ $Y2=0
r116 67 87 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=4.56
+ $Y2=0
r117 67 84 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.6
+ $Y2=0
r118 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r119 64 83 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.705 $Y=0 $X2=3.54
+ $Y2=0
r120 64 66 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=3.705 $Y=0
+ $X2=4.08 $Y2=0
r121 63 86 12.0118 $w=1.7e-07 $l=2.77e-07 $layer=LI1_cond $X=4.28 $Y=0 $X2=4.557
+ $Y2=0
r122 63 66 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=4.28 $Y=0 $X2=4.08
+ $Y2=0
r123 62 81 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.64
+ $Y2=0
r124 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r125 59 80 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.83 $Y=0 $X2=2.665
+ $Y2=0
r126 59 61 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=2.83 $Y=0 $X2=3.12
+ $Y2=0
r127 58 83 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.375 $Y=0 $X2=3.54
+ $Y2=0
r128 58 61 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=3.375 $Y=0
+ $X2=3.12 $Y2=0
r129 57 81 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r130 57 78 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.68
+ $Y2=0
r131 56 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r132 54 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.955 $Y=0 $X2=1.79
+ $Y2=0
r133 54 56 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=1.955 $Y=0
+ $X2=2.16 $Y2=0
r134 53 80 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.5 $Y=0 $X2=2.665
+ $Y2=0
r135 53 56 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=2.5 $Y=0 $X2=2.16
+ $Y2=0
r136 51 78 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r137 50 51 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r138 47 84 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.36 $Y=0 $X2=3.6
+ $Y2=0
r139 47 62 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=3.36 $Y=0
+ $X2=3.12 $Y2=0
r140 45 50 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=0.765 $Y=0 $X2=0.72
+ $Y2=0
r141 45 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.765 $Y=0 $X2=0.93
+ $Y2=0
r142 41 89 3.08095 $w=2.6e-07 $l=1.05924e-07 $layer=LI1_cond $X=6.495 $Y=0.085
+ $X2=6.542 $Y2=0
r143 41 43 13.0758 $w=2.58e-07 $l=2.95e-07 $layer=LI1_cond $X=6.495 $Y=0.085
+ $X2=6.495 $Y2=0.38
r144 37 86 2.33542 $w=5.55e-07 $l=8.5e-08 $layer=LI1_cond $X=4.557 $Y=0.085
+ $X2=4.557 $Y2=0
r145 37 39 6.35753 $w=5.53e-07 $l=2.95e-07 $layer=LI1_cond $X=4.557 $Y=0.085
+ $X2=4.557 $Y2=0.38
r146 33 83 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.54 $Y=0.085
+ $X2=3.54 $Y2=0
r147 33 35 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=3.54 $Y=0.085
+ $X2=3.54 $Y2=0.53
r148 29 80 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.665 $Y=0.085
+ $X2=2.665 $Y2=0
r149 29 31 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.665 $Y=0.085
+ $X2=2.665 $Y2=0.36
r150 25 77 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.79 $Y=0.085
+ $X2=1.79 $Y2=0
r151 25 27 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=1.79 $Y=0.085
+ $X2=1.79 $Y2=0.36
r152 24 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.095 $Y=0 $X2=0.93
+ $Y2=0
r153 23 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.625 $Y=0 $X2=1.79
+ $Y2=0
r154 23 24 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=1.625 $Y=0
+ $X2=1.095 $Y2=0
r155 19 46 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.93 $Y=0.085
+ $X2=0.93 $Y2=0
r156 19 21 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.93 $Y=0.085
+ $X2=0.93 $Y2=0.38
r157 6 43 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=6.32
+ $Y=0.235 $X2=6.46 $Y2=0.38
r158 5 39 45.5 $w=1.7e-07 $l=5.47723e-07 $layer=licon1_NDIFF $count=4 $X=4.26
+ $Y=0.235 $X2=4.74 $Y2=0.38
r159 4 35 182 $w=1.7e-07 $l=3.58225e-07 $layer=licon1_NDIFF $count=1 $X=3.4
+ $Y=0.235 $X2=3.54 $Y2=0.53
r160 3 31 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=2.525
+ $Y=0.235 $X2=2.665 $Y2=0.36
r161 2 27 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=1.65
+ $Y=0.235 $X2=1.79 $Y2=0.36
r162 1 21 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.805
+ $Y=0.235 $X2=0.93 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_LP__A211O_4%A_1006_47# 1 2 9 14 16
r25 10 14 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.335 $Y=0.34
+ $X2=5.17 $Y2=0.34
r26 9 16 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.865 $Y=0.34
+ $X2=6.03 $Y2=0.34
r27 9 10 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=5.865 $Y=0.34
+ $X2=5.335 $Y2=0.34
r28 2 16 91 $w=1.7e-07 $l=1.9799e-07 $layer=licon1_NDIFF $count=2 $X=5.89
+ $Y=0.235 $X2=6.03 $Y2=0.375
r29 1 14 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.03
+ $Y=0.235 $X2=5.17 $Y2=0.38
.ends

