* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__einvn_4 A TE_B VGND VNB VPB VPWR Z
X0 a_87_367# TE_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X1 VPWR TE_B a_555_201# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X2 VPWR TE_B a_87_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X3 Z A a_87_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X4 a_87_367# TE_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X5 a_87_367# A Z VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X6 a_83_69# A Z VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X7 Z A a_83_69# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X8 VPWR TE_B a_87_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X9 VGND TE_B a_555_201# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X10 Z A a_83_69# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X11 VGND a_555_201# a_83_69# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X12 a_83_69# a_555_201# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X13 a_87_367# A Z VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X14 Z A a_87_367# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X15 a_83_69# A Z VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X16 VGND a_555_201# a_83_69# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X17 a_83_69# a_555_201# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
.ends
