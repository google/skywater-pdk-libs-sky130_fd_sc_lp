* File: sky130_fd_sc_lp__and4bb_4.pex.spice
* Created: Fri Aug 28 10:09:28 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__AND4BB_4%B_N 3 6 8 9 10 11 12 19 21
r31 19 22 46.504 $w=3.55e-07 $l=1.65e-07 $layer=POLY_cond $X=0.707 $Y=1.35
+ $X2=0.707 $Y2=1.515
r32 19 21 46.504 $w=3.55e-07 $l=1.65e-07 $layer=POLY_cond $X=0.707 $Y=1.35
+ $X2=0.707 $Y2=1.185
r33 11 12 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.74 $Y=1.665
+ $X2=0.74 $Y2=2.035
r34 10 11 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.74 $Y=1.295
+ $X2=0.74 $Y2=1.665
r35 10 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.72
+ $Y=1.35 $X2=0.72 $Y2=1.35
r36 9 10 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.74 $Y=0.925
+ $X2=0.74 $Y2=1.295
r37 8 9 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.74 $Y=0.555 $X2=0.74
+ $Y2=0.925
r38 6 22 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=0.605 $Y=2.045
+ $X2=0.605 $Y2=1.515
r39 3 21 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.605 $Y=0.865
+ $X2=0.605 $Y2=1.185
.ends

.subckt PM_SKY130_FD_SC_LP__AND4BB_4%A_254_21# 1 2 3 12 16 20 24 28 32 36 40 42
+ 49 51 53 55 56 60 64 66 67 68
c142 64 0 1.99703e-19 $X=4.935 $Y=0.42
c143 53 0 5.82218e-20 $X=2.77 $Y=1.965
c144 49 0 7.53854e-20 $X=2.65 $Y=1.5
c145 40 0 1.53355e-19 $X=2.635 $Y=2.465
c146 36 0 1.25546e-19 $X=2.635 $Y=0.655
r147 73 74 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=2.205 $Y=1.5
+ $X2=2.635 $Y2=1.5
r148 72 73 75.1904 $w=3.3e-07 $l=4.3e-07 $layer=POLY_cond $X=1.775 $Y=1.5
+ $X2=2.205 $Y2=1.5
r149 67 68 24.8349 $w=6.48e-07 $l=9.45e-07 $layer=LI1_cond $X=3.46 $Y=0.647
+ $X2=4.405 $Y2=0.647
r150 64 68 9.75264 $w=6.48e-07 $l=5.3e-07 $layer=LI1_cond $X=4.935 $Y=0.58
+ $X2=4.405 $Y2=0.58
r151 58 60 35.7956 $w=3.28e-07 $l=1.025e-06 $layer=LI1_cond $X=3.425 $Y=2.13
+ $X2=4.45 $Y2=2.13
r152 56 58 19.9058 $w=3.28e-07 $l=5.7e-07 $layer=LI1_cond $X=2.855 $Y=2.13
+ $X2=3.425 $Y2=2.13
r153 55 67 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=2.855 $Y=0.955
+ $X2=3.46 $Y2=0.955
r154 53 56 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.77 $Y=1.965
+ $X2=2.855 $Y2=2.13
r155 52 66 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=2.77 $Y=1.645
+ $X2=2.77 $Y2=1.53
r156 52 53 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=2.77 $Y=1.645
+ $X2=2.77 $Y2=1.965
r157 51 66 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=2.77 $Y=1.415
+ $X2=2.77 $Y2=1.53
r158 50 55 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.77 $Y=1.04
+ $X2=2.855 $Y2=0.955
r159 50 51 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=2.77 $Y=1.04
+ $X2=2.77 $Y2=1.415
r160 49 74 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=2.65 $Y=1.5
+ $X2=2.635 $Y2=1.5
r161 48 49 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.65
+ $Y=1.5 $X2=2.65 $Y2=1.5
r162 45 72 25.3549 $w=3.3e-07 $l=1.45e-07 $layer=POLY_cond $X=1.63 $Y=1.5
+ $X2=1.775 $Y2=1.5
r163 45 69 49.8355 $w=3.3e-07 $l=2.85e-07 $layer=POLY_cond $X=1.63 $Y=1.5
+ $X2=1.345 $Y2=1.5
r164 44 48 51.1083 $w=2.28e-07 $l=1.02e-06 $layer=LI1_cond $X=1.63 $Y=1.53
+ $X2=2.65 $Y2=1.53
r165 44 45 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.63
+ $Y=1.5 $X2=1.63 $Y2=1.5
r166 42 66 0.280307 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.685 $Y=1.53
+ $X2=2.77 $Y2=1.53
r167 42 48 1.75372 $w=2.28e-07 $l=3.5e-08 $layer=LI1_cond $X=2.685 $Y=1.53
+ $X2=2.65 $Y2=1.53
r168 38 74 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.635 $Y=1.665
+ $X2=2.635 $Y2=1.5
r169 38 40 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=2.635 $Y=1.665
+ $X2=2.635 $Y2=2.465
r170 34 74 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.635 $Y=1.335
+ $X2=2.635 $Y2=1.5
r171 34 36 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=2.635 $Y=1.335
+ $X2=2.635 $Y2=0.655
r172 30 73 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.205 $Y=1.665
+ $X2=2.205 $Y2=1.5
r173 30 32 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=2.205 $Y=1.665
+ $X2=2.205 $Y2=2.465
r174 26 73 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.205 $Y=1.335
+ $X2=2.205 $Y2=1.5
r175 26 28 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=2.205 $Y=1.335
+ $X2=2.205 $Y2=0.655
r176 22 72 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.775 $Y=1.665
+ $X2=1.775 $Y2=1.5
r177 22 24 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=1.775 $Y=1.665
+ $X2=1.775 $Y2=2.465
r178 18 72 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.775 $Y=1.335
+ $X2=1.775 $Y2=1.5
r179 18 20 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=1.775 $Y=1.335
+ $X2=1.775 $Y2=0.655
r180 14 69 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.345 $Y=1.665
+ $X2=1.345 $Y2=1.5
r181 14 16 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=1.345 $Y=1.665
+ $X2=1.345 $Y2=2.465
r182 10 69 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.345 $Y=1.335
+ $X2=1.345 $Y2=1.5
r183 10 12 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=1.345 $Y=1.335
+ $X2=1.345 $Y2=0.655
r184 3 60 600 $w=1.7e-07 $l=3.80197e-07 $layer=licon1_PDIFF $count=1 $X=4.255
+ $Y=1.835 $X2=4.45 $Y2=2.13
r185 2 58 600 $w=1.7e-07 $l=3.58225e-07 $layer=licon1_PDIFF $count=1 $X=3.285
+ $Y=1.835 $X2=3.425 $Y2=2.13
r186 1 64 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=4.795
+ $Y=0.235 $X2=4.935 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__AND4BB_4%D 3 7 9 10 14
c43 9 0 1.25546e-19 $X=3.12 $Y=1.295
r44 14 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.19 $Y=1.375
+ $X2=3.19 $Y2=1.54
r45 14 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.19 $Y=1.375
+ $X2=3.19 $Y2=1.21
r46 9 10 15.5056 $w=2.73e-07 $l=3.7e-07 $layer=LI1_cond $X=3.172 $Y=1.295
+ $X2=3.172 $Y2=1.665
r47 9 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.19
+ $Y=1.375 $X2=3.19 $Y2=1.375
r48 7 16 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=3.28 $Y=0.655
+ $X2=3.28 $Y2=1.21
r49 3 17 474.309 $w=1.5e-07 $l=9.25e-07 $layer=POLY_cond $X=3.21 $Y=2.465
+ $X2=3.21 $Y2=1.54
.ends

.subckt PM_SKY130_FD_SC_LP__AND4BB_4%C 3 7 9 10 14
r33 14 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.73 $Y=1.375
+ $X2=3.73 $Y2=1.54
r34 14 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.73 $Y=1.375
+ $X2=3.73 $Y2=1.21
r35 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.73
+ $Y=1.375 $X2=3.73 $Y2=1.375
r36 10 15 7.95734 $w=4.18e-07 $l=2.9e-07 $layer=LI1_cond $X=3.69 $Y=1.665
+ $X2=3.69 $Y2=1.375
r37 9 15 2.19513 $w=4.18e-07 $l=8e-08 $layer=LI1_cond $X=3.69 $Y=1.295 $X2=3.69
+ $Y2=1.375
r38 7 17 474.309 $w=1.5e-07 $l=9.25e-07 $layer=POLY_cond $X=3.64 $Y=2.465
+ $X2=3.64 $Y2=1.54
r39 3 16 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=3.64 $Y=0.655
+ $X2=3.64 $Y2=1.21
.ends

.subckt PM_SKY130_FD_SC_LP__AND4BB_4%A_49_131# 1 2 9 13 17 21 22 23 26 28 29
c89 29 0 3.23513e-19 $X=4.27 $Y=1.51
c90 28 0 1.68512e-19 $X=4.27 $Y=1.51
r91 29 35 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.27 $Y=1.51
+ $X2=4.27 $Y2=1.675
r92 29 34 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.27 $Y=1.51
+ $X2=4.27 $Y2=1.345
r93 28 31 6.44012 $w=3.38e-07 $l=1.9e-07 $layer=LI1_cond $X=4.275 $Y=1.51
+ $X2=4.275 $Y2=1.7
r94 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.27
+ $Y=1.51 $X2=4.27 $Y2=1.51
r95 25 26 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=4.875 $Y=1.785
+ $X2=4.875 $Y2=2.465
r96 24 31 4.80115 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=4.445 $Y=1.7
+ $X2=4.275 $Y2=1.7
r97 23 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.79 $Y=1.7
+ $X2=4.875 $Y2=1.785
r98 23 24 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=4.79 $Y=1.7
+ $X2=4.445 $Y2=1.7
r99 21 26 6.82373 $w=1.8e-07 $l=1.25499e-07 $layer=LI1_cond $X=4.79 $Y=2.555
+ $X2=4.875 $Y2=2.465
r100 21 22 267.106 $w=1.78e-07 $l=4.335e-06 $layer=LI1_cond $X=4.79 $Y=2.555
+ $X2=0.455 $Y2=2.555
r101 17 20 54.3953 $w=2.48e-07 $l=1.18e-06 $layer=LI1_cond $X=0.33 $Y=0.865
+ $X2=0.33 $Y2=2.045
r102 15 22 7.0541 $w=1.8e-07 $l=1.63936e-07 $layer=LI1_cond $X=0.33 $Y=2.465
+ $X2=0.455 $Y2=2.555
r103 15 20 19.361 $w=2.48e-07 $l=4.2e-07 $layer=LI1_cond $X=0.33 $Y=2.465
+ $X2=0.33 $Y2=2.045
r104 13 35 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=4.18 $Y=2.465
+ $X2=4.18 $Y2=1.675
r105 9 34 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=4.18 $Y=0.655
+ $X2=4.18 $Y2=1.345
r106 2 20 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=0.245
+ $Y=1.835 $X2=0.37 $Y2=2.045
r107 1 17 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.245
+ $Y=0.655 $X2=0.37 $Y2=0.865
.ends

.subckt PM_SKY130_FD_SC_LP__AND4BB_4%A_929_21# 1 2 9 12 14 18 22 24 28 30 32 33
+ 36
c54 24 0 1.2381e-19 $X=4.81 $Y=1.16
c55 12 0 1.68512e-19 $X=4.72 $Y=2.465
r56 32 33 8.48463 $w=2.98e-07 $l=1.65e-07 $layer=LI1_cond $X=5.49 $Y=2.095
+ $X2=5.49 $Y2=1.93
r57 28 37 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.81 $Y=1.35
+ $X2=4.81 $Y2=1.515
r58 28 36 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.81 $Y=1.35
+ $X2=4.81 $Y2=1.185
r59 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.81
+ $Y=1.35 $X2=4.81 $Y2=1.35
r60 24 27 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=4.81 $Y=1.16
+ $X2=4.81 $Y2=1.35
r61 20 22 9.52982 $w=2.58e-07 $l=2.15e-07 $layer=LI1_cond $X=6.015 $Y=1.075
+ $X2=6.015 $Y2=0.86
r62 19 30 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.51 $Y=1.16
+ $X2=5.425 $Y2=1.16
r63 18 20 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=5.885 $Y=1.16
+ $X2=6.015 $Y2=1.075
r64 18 19 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=5.885 $Y=1.16
+ $X2=5.51 $Y2=1.16
r65 16 30 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.425 $Y=1.245
+ $X2=5.425 $Y2=1.16
r66 16 33 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=5.425 $Y=1.245
+ $X2=5.425 $Y2=1.93
r67 15 24 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.975 $Y=1.16
+ $X2=4.81 $Y2=1.16
r68 14 30 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.34 $Y=1.16
+ $X2=5.425 $Y2=1.16
r69 14 15 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=5.34 $Y=1.16
+ $X2=4.975 $Y2=1.16
r70 12 37 487.128 $w=1.5e-07 $l=9.5e-07 $layer=POLY_cond $X=4.72 $Y=2.465
+ $X2=4.72 $Y2=1.515
r71 9 36 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=4.72 $Y=0.655
+ $X2=4.72 $Y2=1.185
r72 2 32 600 $w=1.7e-07 $l=3.2249e-07 $layer=licon1_PDIFF $count=1 $X=5.335
+ $Y=1.835 $X2=5.475 $Y2=2.095
r73 1 22 182 $w=1.7e-07 $l=2.7627e-07 $layer=licon1_NDIFF $count=1 $X=5.84
+ $Y=0.645 $X2=5.98 $Y2=0.86
.ends

.subckt PM_SKY130_FD_SC_LP__AND4BB_4%A_N 3 5 6 9 11 14 15
r30 14 17 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=5.855 $Y=1.51
+ $X2=5.855 $Y2=1.6
r31 14 16 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=5.855 $Y=1.51
+ $X2=5.855 $Y2=1.345
r32 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.855
+ $Y=1.51 $X2=5.855 $Y2=1.51
r33 11 15 4.11983 $w=4.48e-07 $l=1.55e-07 $layer=LI1_cond $X=5.915 $Y=1.665
+ $X2=5.915 $Y2=1.51
r34 9 16 251.255 $w=1.5e-07 $l=4.9e-07 $layer=POLY_cond $X=5.765 $Y=0.855
+ $X2=5.765 $Y2=1.345
r35 5 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.69 $Y=1.6
+ $X2=5.855 $Y2=1.6
r36 5 6 182.032 $w=1.5e-07 $l=3.55e-07 $layer=POLY_cond $X=5.69 $Y=1.6 $X2=5.335
+ $Y2=1.6
r37 1 6 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.26 $Y=1.675
+ $X2=5.335 $Y2=1.6
r38 1 3 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=5.26 $Y=1.675 $X2=5.26
+ $Y2=2.045
.ends

.subckt PM_SKY130_FD_SC_LP__AND4BB_4%VPWR 1 2 3 4 5 18 22 26 30 34 37 38 40 41
+ 43 44 45 47 62 68 69 72 75
r76 75 76 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r77 72 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r78 69 76 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=5.04
+ $Y2=3.33
r79 68 69 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r80 66 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.1 $Y=3.33
+ $X2=4.935 $Y2=3.33
r81 66 68 58.7166 $w=1.68e-07 $l=9e-07 $layer=LI1_cond $X=5.1 $Y=3.33 $X2=6
+ $Y2=3.33
r82 65 76 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.04 $Y2=3.33
r83 64 65 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r84 62 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.77 $Y=3.33
+ $X2=4.935 $Y2=3.33
r85 62 64 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=4.77 $Y=3.33
+ $X2=4.56 $Y2=3.33
r86 61 65 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.56 $Y2=3.33
r87 60 61 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r88 57 58 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r89 55 58 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r90 55 73 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r91 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r92 52 72 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.295 $Y=3.33
+ $X2=1.13 $Y2=3.33
r93 52 54 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=1.295 $Y=3.33
+ $X2=1.68 $Y2=3.33
r94 50 73 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r95 49 50 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r96 47 72 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.965 $Y=3.33
+ $X2=1.13 $Y2=3.33
r97 47 49 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=0.965 $Y=3.33
+ $X2=0.72 $Y2=3.33
r98 45 61 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r99 45 58 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=2.64 $Y2=3.33
r100 43 60 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=3.75 $Y=3.33 $X2=3.6
+ $Y2=3.33
r101 43 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.75 $Y=3.33
+ $X2=3.915 $Y2=3.33
r102 42 64 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r103 42 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.08 $Y=3.33
+ $X2=3.915 $Y2=3.33
r104 40 57 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=2.765 $Y=3.33
+ $X2=2.64 $Y2=3.33
r105 40 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.765 $Y=3.33
+ $X2=2.93 $Y2=3.33
r106 39 60 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=3.095 $Y=3.33
+ $X2=3.6 $Y2=3.33
r107 39 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.095 $Y=3.33
+ $X2=2.93 $Y2=3.33
r108 37 54 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=1.825 $Y=3.33
+ $X2=1.68 $Y2=3.33
r109 37 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.825 $Y=3.33
+ $X2=1.99 $Y2=3.33
r110 36 57 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=2.155 $Y=3.33
+ $X2=2.64 $Y2=3.33
r111 36 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.155 $Y=3.33
+ $X2=1.99 $Y2=3.33
r112 32 75 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.935 $Y=3.245
+ $X2=4.935 $Y2=3.33
r113 32 34 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=4.935 $Y=3.245
+ $X2=4.935 $Y2=2.95
r114 28 44 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.915 $Y=3.245
+ $X2=3.915 $Y2=3.33
r115 28 30 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=3.915 $Y=3.245
+ $X2=3.915 $Y2=2.95
r116 24 41 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.93 $Y=3.245
+ $X2=2.93 $Y2=3.33
r117 24 26 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.93 $Y=3.245
+ $X2=2.93 $Y2=2.95
r118 20 38 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.99 $Y=3.245
+ $X2=1.99 $Y2=3.33
r119 20 22 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.99 $Y=3.245
+ $X2=1.99 $Y2=2.95
r120 16 72 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.13 $Y=3.245
+ $X2=1.13 $Y2=3.33
r121 16 18 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.13 $Y=3.245
+ $X2=1.13 $Y2=2.95
r122 5 34 600 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=4.795
+ $Y=1.835 $X2=4.935 $Y2=2.95
r123 4 30 600 $w=1.7e-07 $l=1.21088e-06 $layer=licon1_PDIFF $count=1 $X=3.715
+ $Y=1.835 $X2=3.915 $Y2=2.95
r124 3 26 600 $w=1.7e-07 $l=1.22005e-06 $layer=licon1_PDIFF $count=1 $X=2.71
+ $Y=1.835 $X2=2.93 $Y2=2.95
r125 2 22 600 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=1.85
+ $Y=1.835 $X2=1.99 $Y2=2.95
r126 1 18 600 $w=1.7e-07 $l=1.32097e-06 $layer=licon1_PDIFF $count=1 $X=0.68
+ $Y=1.835 $X2=1.13 $Y2=2.95
.ends

.subckt PM_SKY130_FD_SC_LP__AND4BB_4%X 1 2 3 4 13 17 21 23 24 27 34
c53 17 0 1.53355e-19 $X=2.42 $Y=1.98
c54 13 0 1.63555e-19 $X=1.295 $Y=1.98
r55 33 34 9.24242 $w=1.78e-07 $l=1.5e-07 $layer=LI1_cond $X=1.205 $Y=1.815
+ $X2=1.205 $Y2=1.665
r56 30 34 25.8788 $w=1.78e-07 $l=4.2e-07 $layer=LI1_cond $X=1.205 $Y=1.245
+ $X2=1.205 $Y2=1.665
r57 29 30 0.364908 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=1.205 $Y=1.16
+ $X2=1.205 $Y2=1.245
r58 25 27 38.2345 $w=1.88e-07 $l=6.55e-07 $layer=LI1_cond $X=2.42 $Y=1.075
+ $X2=2.42 $Y2=0.42
r59 23 25 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=2.325 $Y=1.16
+ $X2=2.42 $Y2=1.075
r60 23 24 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.325 $Y=1.16
+ $X2=1.655 $Y2=1.16
r61 19 24 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=1.54 $Y=1.16
+ $X2=1.655 $Y2=1.16
r62 19 29 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.54 $Y=1.16
+ $X2=1.205 $Y2=1.16
r63 19 21 32.8196 $w=2.28e-07 $l=6.55e-07 $layer=LI1_cond $X=1.54 $Y=1.075
+ $X2=1.54 $Y2=0.42
r64 15 17 30.0334 $w=3.28e-07 $l=8.6e-07 $layer=LI1_cond $X=1.56 $Y=1.98
+ $X2=2.42 $Y2=1.98
r65 13 33 7.61292 $w=3.3e-07 $l=2.05122e-07 $layer=LI1_cond $X=1.295 $Y=1.98
+ $X2=1.205 $Y2=1.815
r66 13 15 9.25447 $w=3.28e-07 $l=2.65e-07 $layer=LI1_cond $X=1.295 $Y=1.98
+ $X2=1.56 $Y2=1.98
r67 4 17 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.28
+ $Y=1.835 $X2=2.42 $Y2=1.98
r68 3 15 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.42
+ $Y=1.835 $X2=1.56 $Y2=1.98
r69 2 27 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=2.28
+ $Y=0.235 $X2=2.42 $Y2=0.42
r70 1 21 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=1.42
+ $Y=0.235 $X2=1.56 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__AND4BB_4%VGND 1 2 3 4 15 19 23 27 30 31 33 34 36 37
+ 38 50 59 60 63
c76 23 0 7.53854e-20 $X=2.955 $Y=0.535
r77 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.52 $Y=0 $X2=5.52
+ $Y2=0
r78 60 64 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=0 $X2=5.52
+ $Y2=0
r79 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=0 $X2=6 $Y2=0
r80 57 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.715 $Y=0 $X2=5.55
+ $Y2=0
r81 57 59 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=5.715 $Y=0 $X2=6
+ $Y2=0
r82 56 64 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=5.04 $Y=0 $X2=5.52
+ $Y2=0
r83 55 56 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.04 $Y=0 $X2=5.04
+ $Y2=0
r84 52 55 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=3.12 $Y=0 $X2=5.04
+ $Y2=0
r85 50 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.385 $Y=0 $X2=5.55
+ $Y2=0
r86 50 55 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=5.385 $Y=0 $X2=5.04
+ $Y2=0
r87 48 49 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r88 46 49 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r89 45 46 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r90 42 46 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.68
+ $Y2=0
r91 41 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r92 38 56 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=3.12 $Y=0 $X2=5.04
+ $Y2=0
r93 38 49 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.64
+ $Y2=0
r94 38 52 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r95 37 52 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.955 $Y=0 $X2=3.12
+ $Y2=0
r96 36 48 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=2.79 $Y=0 $X2=2.64
+ $Y2=0
r97 36 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.79 $Y=0 $X2=2.955
+ $Y2=0
r98 33 45 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=1.825 $Y=0 $X2=1.68
+ $Y2=0
r99 33 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.825 $Y=0 $X2=1.99
+ $Y2=0
r100 32 48 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=2.155 $Y=0
+ $X2=2.64 $Y2=0
r101 32 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.155 $Y=0 $X2=1.99
+ $Y2=0
r102 30 41 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.025 $Y=0
+ $X2=0.72 $Y2=0
r103 30 31 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=1.025 $Y=0 $X2=1.14
+ $Y2=0
r104 29 45 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=1.255 $Y=0
+ $X2=1.68 $Y2=0
r105 29 31 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=1.255 $Y=0 $X2=1.14
+ $Y2=0
r106 25 63 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.55 $Y=0.085
+ $X2=5.55 $Y2=0
r107 25 27 24.9696 $w=3.28e-07 $l=7.15e-07 $layer=LI1_cond $X=5.55 $Y=0.085
+ $X2=5.55 $Y2=0.8
r108 21 37 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.955 $Y=0.085
+ $X2=2.955 $Y2=0
r109 21 23 15.7151 $w=3.28e-07 $l=4.5e-07 $layer=LI1_cond $X=2.955 $Y=0.085
+ $X2=2.955 $Y2=0.535
r110 17 34 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.99 $Y=0.085
+ $X2=1.99 $Y2=0
r111 17 19 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.99 $Y=0.085
+ $X2=1.99 $Y2=0.38
r112 13 31 0.280307 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.14 $Y=0.085
+ $X2=1.14 $Y2=0
r113 13 15 14.7813 $w=2.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.14 $Y=0.085
+ $X2=1.14 $Y2=0.38
r114 4 27 182 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=1 $X=5.425
+ $Y=0.645 $X2=5.55 $Y2=0.8
r115 3 23 182 $w=1.7e-07 $l=4.04351e-07 $layer=licon1_NDIFF $count=1 $X=2.71
+ $Y=0.235 $X2=2.955 $Y2=0.535
r116 2 19 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.85
+ $Y=0.235 $X2=1.99 $Y2=0.38
r117 1 15 91 $w=1.7e-07 $l=5.71183e-07 $layer=licon1_NDIFF $count=2 $X=0.68
+ $Y=0.655 $X2=1.13 $Y2=0.38
.ends

