* File: sky130_fd_sc_lp__o41a_1.spice
* Created: Wed Sep  2 10:27:26 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__o41a_1.pex.spice"
.subckt sky130_fd_sc_lp__o41a_1  VNB VPB B1 A4 A3 A2 A1 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* A1	A1
* A2	A2
* A3	A3
* A4	A4
* B1	B1
* VPB	VPB
* VNB	VNB
MM1001 N_VGND_M1001_d N_A_155_23#_M1001_g N_X_M1001_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.5082 PD=2.21 PS=2.89 NRD=0 NRS=24.276 M=1 R=5.6 SA=75000.5
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1002 N_A_375_49#_M1002_d N_B1_M1002_g N_A_155_23#_M1002_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75002.2 A=0.126 P=1.98 MULT=1
MM1005 N_VGND_M1005_d N_A4_M1005_g N_A_375_49#_M1002_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1806 AS=0.1176 PD=1.27 PS=1.12 NRD=9.996 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75001.7 A=0.126 P=1.98 MULT=1
MM1004 N_A_375_49#_M1004_d N_A3_M1004_g N_VGND_M1005_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1806 PD=1.12 PS=1.27 NRD=0 NRS=11.424 M=1 R=5.6 SA=75001.2
+ SB=75001.2 A=0.126 P=1.98 MULT=1
MM1007 N_VGND_M1007_d N_A2_M1007_g N_A_375_49#_M1004_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1638 AS=0.1176 PD=1.23 PS=1.12 NRD=9.996 NRS=0 M=1 R=5.6 SA=75001.6
+ SB=75000.7 A=0.126 P=1.98 MULT=1
MM1011 N_A_375_49#_M1011_d N_A1_M1011_g N_VGND_M1007_d VNB NSHORT L=0.15 W=0.84
+ AD=0.2226 AS=0.1638 PD=2.21 PS=1.23 NRD=0 NRS=5.712 M=1 R=5.6 SA=75002.2
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1008 N_VPWR_M1008_d N_A_155_23#_M1008_g N_X_M1008_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.2646 AS=0.7623 PD=1.68 PS=3.73 NRD=10.9335 NRS=0 M=1 R=8.4 SA=75000.5
+ SB=75002.9 A=0.189 P=2.82 MULT=1
MM1010 N_A_155_23#_M1010_d N_B1_M1010_g N_VPWR_M1008_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.25515 AS=0.2646 PD=1.665 PS=1.68 NRD=0 NRS=10.9335 M=1 R=8.4 SA=75001.1
+ SB=75002.4 A=0.189 P=2.82 MULT=1
MM1000 A_447_367# N_A4_M1000_g N_A_155_23#_M1010_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3024 AS=0.25515 PD=1.74 PS=1.665 NRD=28.9196 NRS=19.5424 M=1 R=8.4
+ SA=75001.7 SB=75001.8 A=0.189 P=2.82 MULT=1
MM1006 A_573_367# N_A3_M1006_g A_447_367# VPB PHIGHVT L=0.15 W=1.26 AD=0.189
+ AS=0.3024 PD=1.56 PS=1.74 NRD=14.8341 NRS=28.9196 M=1 R=8.4 SA=75002.3
+ SB=75001.2 A=0.189 P=2.82 MULT=1
MM1009 A_663_367# N_A2_M1009_g A_573_367# VPB PHIGHVT L=0.15 W=1.26 AD=0.2457
+ AS=0.189 PD=1.65 PS=1.56 NRD=21.8867 NRS=14.8341 M=1 R=8.4 SA=75002.7
+ SB=75000.7 A=0.189 P=2.82 MULT=1
MM1003 N_VPWR_M1003_d N_A1_M1003_g A_663_367# VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.2457 PD=3.05 PS=1.65 NRD=0 NRS=21.8867 M=1 R=8.4 SA=75003.3
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX12_noxref VNB VPB NWDIODE A=8.7655 P=13.13
c_67 VPB 0 1.17498e-19 $X=0 $Y=3.085
*
.include "sky130_fd_sc_lp__o41a_1.pxi.spice"
*
.ends
*
*
