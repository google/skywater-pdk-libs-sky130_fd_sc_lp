* NGSPICE file created from sky130_fd_sc_lp__a21boi_0.ext - technology: sky130A

.subckt sky130_fd_sc_lp__a21boi_0 A1 A2 B1_N VGND VNB VPB VPWR Y
M1000 a_350_47# A1 Y VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=1.176e+11p ps=1.4e+06u
M1001 a_324_483# a_27_47# Y VPB phighvt w=640000u l=150000u
+  ad=3.488e+11p pd=3.65e+06u as=1.696e+11p ps=1.81e+06u
M1002 VGND B1_N a_27_47# VNB nshort w=420000u l=150000u
+  ad=3.717e+11p pd=3.45e+06u as=1.113e+11p ps=1.37e+06u
M1003 a_324_483# A2 VPWR VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=2.905e+11p ps=3.21e+06u
M1004 VPWR B1_N a_27_47# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1005 VPWR A1 a_324_483# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 Y a_27_47# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND A2 a_350_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

