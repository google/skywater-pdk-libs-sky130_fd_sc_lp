* NGSPICE file created from sky130_fd_sc_lp__buflp_0.ext - technology: sky130A

.subckt sky130_fd_sc_lp__buflp_0 A VGND VNB VPB VPWR X
M1000 VPWR A a_128_490# VPB phighvt w=420000u l=150000u
+  ad=2.286e+11p pd=2.07e+06u as=1.008e+11p ps=1.32e+06u
M1001 X a_36_120# a_315_446# VPB phighvt w=640000u l=150000u
+  ad=1.824e+11p pd=1.85e+06u as=1.536e+11p ps=1.76e+06u
M1002 a_287_120# a_36_120# VGND VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=1.176e+11p ps=1.4e+06u
M1003 VGND A a_123_120# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1004 a_315_446# a_36_120# VPWR VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 X a_36_120# a_287_120# VNB nshort w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=0p ps=0u
M1006 a_128_490# A a_36_120# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1007 a_123_120# A a_36_120# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
.ends

