* File: sky130_fd_sc_lp__sdfxbp_lp.spice
* Created: Fri Aug 28 11:30:31 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__sdfxbp_lp.pex.spice"
.subckt sky130_fd_sc_lp__sdfxbp_lp  VNB VPB D SCE SCD CLK VPWR Q Q_N VGND
* 
* VGND	VGND
* Q_N	Q_N
* Q	Q
* VPWR	VPWR
* CLK	CLK
* SCD	SCD
* SCE	SCE
* D	D
* VPB	VPB
* VNB	VNB
MM1037 A_141_125# N_SCE_M1037_g N_A_27_409#_M1037_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.1197 PD=0.66 PS=1.41 NRD=18.564 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.5 A=0.063 P=1.14 MULT=1
MM1008 N_VGND_M1008_d N_SCE_M1008_g A_141_125# VNB NSHORT L=0.15 W=0.42
+ AD=0.0924 AS=0.0504 PD=0.86 PS=0.66 NRD=22.848 NRS=18.564 M=1 R=2.8 SA=75000.6
+ SB=75002.1 A=0.063 P=1.14 MULT=1
MM1015 A_337_125# N_A_27_409#_M1015_g N_VGND_M1008_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0504 AS=0.0924 PD=0.66 PS=0.86 NRD=18.564 NRS=22.848 M=1 R=2.8 SA=75001.2
+ SB=75001.5 A=0.063 P=1.14 MULT=1
MM1003 N_A_343_417#_M1003_d N_D_M1003_g A_337_125# VNB NSHORT L=0.15 W=0.42
+ AD=0.0819 AS=0.0504 PD=0.81 PS=0.66 NRD=31.428 NRS=18.564 M=1 R=2.8 SA=75001.6
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1020 A_523_125# N_SCE_M1020_g N_A_343_417#_M1003_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0819 PD=0.63 PS=0.81 NRD=14.28 NRS=0 M=1 R=2.8 SA=75002.1
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1012 N_VGND_M1012_d N_SCD_M1012_g A_523_125# VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75002.5
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1035 A_789_66# N_CLK_M1035_g N_A_706_66#_M1035_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1113 PD=0.63 PS=1.37 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.3 A=0.063 P=1.14 MULT=1
MM1021 N_VGND_M1021_d N_CLK_M1021_g A_789_66# VNB NSHORT L=0.15 W=0.42 AD=0.0588
+ AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6 SB=75001 A=0.063
+ P=1.14 MULT=1
MM1004 A_947_66# N_A_706_66#_M1004_g N_VGND_M1021_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75001
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1039 N_A_975_347#_M1039_d N_A_706_66#_M1039_g A_947_66# VNB NSHORT L=0.15
+ W=0.42 AD=0.1134 AS=0.0441 PD=1.38 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8
+ SA=75001.3 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1014 N_A_1278_155#_M1014_d N_A_975_347#_M1014_g N_A_1127_155#_M1014_s VNB
+ NSHORT L=0.15 W=0.42 AD=0.0609 AS=0.2541 PD=0.71 PS=2.05 NRD=2.856 NRS=97.14
+ M=1 R=2.8 SA=75000.5 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1041 N_A_343_417#_M1041_d N_A_706_66#_M1041_g N_A_1278_155#_M1014_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.1113 AS=0.0609 PD=1.37 PS=0.71 NRD=0 NRS=0 M=1 R=2.8
+ SA=75001 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1009 N_VGND_M1009_d N_A_1530_231#_M1009_g N_A_1127_155#_M1009_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.1147 AS=0.1113 PD=1.05 PS=1.37 NRD=62.304 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1028 A_1674_125# N_A_1278_155#_M1028_g N_VGND_M1009_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1147 PD=0.63 PS=1.05 NRD=14.28 NRS=19.992 M=1 R=2.8 SA=75000.7
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1018 N_A_1530_231#_M1018_d N_A_1278_155#_M1018_g A_1674_125# VNB NSHORT L=0.15
+ W=0.42 AD=0.1113 AS=0.0441 PD=1.37 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8
+ SA=75001.1 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1042 N_A_1902_347#_M1042_d N_A_706_66#_M1042_g N_A_1859_155#_M1042_s VNB
+ NSHORT L=0.15 W=0.42 AD=0.07245 AS=0.1113 PD=0.765 PS=1.37 NRD=18.564 NRS=0
+ M=1 R=2.8 SA=75000.2 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1022 N_A_1530_231#_M1022_d N_A_975_347#_M1022_g N_A_1902_347#_M1042_d VNB
+ NSHORT L=0.15 W=0.42 AD=0.28115 AS=0.07245 PD=2.64 PS=0.765 NRD=175.536 NRS=0
+ M=1 R=2.8 SA=75000.7 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1001 N_VGND_M1001_d N_A_2089_254#_M1001_g N_A_1859_155#_M1001_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.0588 AS=0.1134 PD=0.7 PS=1.38 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001 A=0.063 P=1.14 MULT=1
MM1016 A_2331_57# N_A_1902_347#_M1016_g N_VGND_M1001_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1002 N_A_2089_254#_M1002_d N_A_1902_347#_M1002_g A_2331_57# VNB NSHORT L=0.15
+ W=0.42 AD=0.1113 AS=0.0441 PD=1.37 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1043 A_2593_127# N_A_2089_254#_M1043_g N_Q_M1043_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1113 PD=0.63 PS=1.37 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.3 A=0.063 P=1.14 MULT=1
MM1025 N_VGND_M1025_d N_A_2089_254#_M1025_g A_2593_127# VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1029 A_2751_127# N_A_2089_254#_M1029_g N_VGND_M1025_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0588 PD=0.63 PS=0.7 NRD=14.28 NRS=0 M=1 R=2.8 SA=75001
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1023 N_A_2714_401#_M1023_d N_A_2089_254#_M1023_g A_2751_127# VNB NSHORT L=0.15
+ W=0.42 AD=0.1134 AS=0.0441 PD=1.38 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8
+ SA=75001.3 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1031 A_3015_57# N_A_2714_401#_M1031_g N_VGND_M1031_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1134 PD=0.63 PS=1.38 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1026 N_Q_N_M1026_d N_A_2714_401#_M1026_g A_3015_57# VNB NSHORT L=0.15 W=0.42
+ AD=0.1134 AS=0.0441 PD=1.38 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1017 N_VPWR_M1017_d N_SCE_M1017_g N_A_27_409#_M1017_s VPB PHIGHVT L=0.25 W=1
+ AD=0.27 AS=0.27 PD=2.54 PS=2.54 NRD=0 NRS=0 M=1 R=4 SA=125000 SB=125000 A=0.25
+ P=2.5 MULT=1
MM1036 N_A_343_417#_M1036_d N_A_27_409#_M1036_g N_A_239_417#_M1036_s VPB PHIGHVT
+ L=0.25 W=1 AD=0.14 AS=0.27 PD=1.28 PS=2.54 NRD=0 NRS=0 M=1 R=4 SA=125000
+ SB=125002 A=0.25 P=2.5 MULT=1
MM1019 A_449_417# N_D_M1019_g N_A_343_417#_M1036_d VPB PHIGHVT L=0.25 W=1
+ AD=0.11 AS=0.14 PD=1.22 PS=1.28 NRD=10.8153 NRS=0 M=1 R=4 SA=125001 SB=125001
+ A=0.25 P=2.5 MULT=1
MM1006 N_VPWR_M1006_d N_SCE_M1006_g A_449_417# VPB PHIGHVT L=0.25 W=1 AD=0.14
+ AS=0.11 PD=1.28 PS=1.22 NRD=0 NRS=10.8153 M=1 R=4 SA=125001 SB=125001 A=0.25
+ P=2.5 MULT=1
MM1040 N_A_239_417#_M1040_d N_SCD_M1040_g N_VPWR_M1006_d VPB PHIGHVT L=0.25 W=1
+ AD=0.285 AS=0.14 PD=2.57 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125002 SB=125000
+ A=0.25 P=2.5 MULT=1
MM1005 N_VPWR_M1005_d N_CLK_M1005_g N_A_706_66#_M1005_s VPB PHIGHVT L=0.25 W=1
+ AD=0.14 AS=0.285 PD=1.28 PS=2.57 NRD=0 NRS=0 M=1 R=4 SA=125000 SB=125001
+ A=0.25 P=2.5 MULT=1
MM1030 N_A_975_347#_M1030_d N_A_706_66#_M1030_g N_VPWR_M1005_d VPB PHIGHVT
+ L=0.25 W=1 AD=0.285 AS=0.14 PD=2.57 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125001
+ SB=125000 A=0.25 P=2.5 MULT=1
MM1010 N_A_1278_155#_M1010_d N_A_975_347#_M1010_g N_A_343_417#_M1010_s VPB
+ PHIGHVT L=0.25 W=1 AD=0.14 AS=0.285 PD=1.28 PS=2.57 NRD=0 NRS=0 M=1 R=4
+ SA=125000 SB=125005 A=0.25 P=2.5 MULT=1
MM1038 A_1482_347# N_A_706_66#_M1038_g N_A_1278_155#_M1010_d VPB PHIGHVT L=0.25
+ W=1 AD=0.12 AS=0.14 PD=1.24 PS=1.28 NRD=12.7853 NRS=0 M=1 R=4 SA=125001
+ SB=125004 A=0.25 P=2.5 MULT=1
MM1007 N_VPWR_M1007_d N_A_1530_231#_M1007_g A_1482_347# VPB PHIGHVT L=0.25 W=1
+ AD=0.31 AS=0.12 PD=1.62 PS=1.24 NRD=0 NRS=12.7853 M=1 R=4 SA=125001 SB=125004
+ A=0.25 P=2.5 MULT=1
MM1013 N_A_1530_231#_M1013_d N_A_1278_155#_M1013_g N_VPWR_M1007_d VPB PHIGHVT
+ L=0.25 W=1 AD=0.245 AS=0.31 PD=1.49 PS=1.62 NRD=0 NRS=66.98 M=1 R=4 SA=125002
+ SB=125003 A=0.25 P=2.5 MULT=1
MM1024 N_A_1902_347#_M1024_d N_A_706_66#_M1024_g N_A_1530_231#_M1013_d VPB
+ PHIGHVT L=0.25 W=1 AD=0.223625 AS=0.245 PD=1.465 PS=1.49 NRD=15.7403
+ NRS=41.3503 M=1 R=4 SA=125003 SB=125002 A=0.25 P=2.5 MULT=1
MM1033 A_2040_352# N_A_975_347#_M1033_g N_A_1902_347#_M1024_d VPB PHIGHVT L=0.25
+ W=1 AD=0.1225 AS=0.223625 PD=1.245 PS=1.465 NRD=13.2778 NRS=15.7403 M=1 R=4
+ SA=125003 SB=125001 A=0.25 P=2.5 MULT=1
MM1034 N_VPWR_M1034_d N_A_2089_254#_M1034_g A_2040_352# VPB PHIGHVT L=0.25 W=1
+ AD=0.226525 AS=0.1225 PD=1.485 PS=1.245 NRD=15.7403 NRS=13.2778 M=1 R=4
+ SA=125004 SB=125001 A=0.25 P=2.5 MULT=1
MM1000 N_A_2089_254#_M1000_d N_A_1902_347#_M1000_g N_VPWR_M1034_d VPB PHIGHVT
+ L=0.25 W=1 AD=0.285 AS=0.226525 PD=2.57 PS=1.485 NRD=0 NRS=15.7403 M=1 R=4
+ SA=125004 SB=125000 A=0.25 P=2.5 MULT=1
MM1032 N_VPWR_M1032_d N_A_2089_254#_M1032_g N_Q_M1032_s VPB PHIGHVT L=0.25 W=1
+ AD=0.14 AS=0.285 PD=1.28 PS=2.57 NRD=0 NRS=0 M=1 R=4 SA=125000 SB=125001
+ A=0.25 P=2.5 MULT=1
MM1011 N_A_2714_401#_M1011_d N_A_2089_254#_M1011_g N_VPWR_M1032_d VPB PHIGHVT
+ L=0.25 W=1 AD=0.285 AS=0.14 PD=2.57 PS=1.28 NRD=0 NRS=0 M=1 R=4 SA=125001
+ SB=125000 A=0.25 P=2.5 MULT=1
MM1027 N_Q_N_M1027_d N_A_2714_401#_M1027_g N_VPWR_M1027_s VPB PHIGHVT L=0.25 W=1
+ AD=0.285 AS=0.285 PD=2.57 PS=2.57 NRD=0 NRS=0 M=1 R=4 SA=125000 SB=125000
+ A=0.25 P=2.5 MULT=1
DX44_noxref VNB VPB NWDIODE A=31.0274 P=36.37
c_157 VNB 0 1.71737e-19 $X=0 $Y=0
*
.include "sky130_fd_sc_lp__sdfxbp_lp.pxi.spice"
*
.ends
*
*
