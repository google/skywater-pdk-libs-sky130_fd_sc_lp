* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__sdfsbp_2 CLK D SCD SCE SET_B VGND VNB VPB VPWR Q Q_N
X0 VGND a_2624_49# Q VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X1 VGND a_629_47# a_920_73# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 VGND a_1799_408# a_2624_49# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 VGND CLK a_629_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 a_268_467# a_629_47# a_1163_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 Q_N a_1799_408# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X6 Q a_2624_49# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X7 VPWR SET_B a_1799_408# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X8 Q a_2624_49# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X9 a_27_467# SCE VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 a_1735_119# a_920_73# a_1799_408# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X11 VPWR a_1799_408# a_2624_49# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X12 a_268_467# a_27_467# a_376_467# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X13 a_471_47# SCD VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X14 VGND a_1799_408# Q_N VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X15 a_2001_119# SET_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X16 VPWR SCE a_196_467# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X17 a_196_467# D a_268_467# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X18 a_1291_93# a_1163_119# a_1530_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X19 a_1799_408# a_629_47# a_1929_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X20 VPWR a_1163_119# a_1291_93# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X21 VGND a_27_467# a_268_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X22 Q_N a_1799_408# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X23 a_268_467# a_920_73# a_1163_119# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X24 VPWR a_1799_408# Q_N VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X25 a_27_467# SCE VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X26 a_1799_408# a_920_73# a_1904_492# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X27 a_1904_492# a_1946_369# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X28 a_376_467# SCD VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X29 VPWR a_1163_119# a_1697_379# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X30 a_1697_379# a_629_47# a_1799_408# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X31 a_268_467# SCE a_471_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X32 a_1249_119# a_1291_93# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X33 a_1946_369# a_1799_408# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X34 a_1291_93# SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X35 a_1946_369# a_1799_408# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X36 VPWR CLK a_629_47# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X37 a_1163_119# a_629_47# a_1275_463# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X38 a_1163_119# a_920_73# a_1249_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X39 a_1530_119# SET_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X40 VPWR a_629_47# a_920_73# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X41 a_1275_463# a_1291_93# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X42 a_1929_119# a_1946_369# a_2001_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X43 VPWR a_2624_49# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X44 a_268_47# D a_268_467# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X45 VGND a_1163_119# a_1735_119# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
.ends
