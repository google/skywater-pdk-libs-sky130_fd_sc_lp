* File: sky130_fd_sc_lp__o211ai_4.pex.spice
* Created: Fri Aug 28 11:03:09 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__O211AI_4%A1 3 7 11 15 19 23 27 31 33 41 42 43 45 46
+ 51 52 53 54 55 56 63 70 75
r122 63 66 13.1146 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=0.55 $Y=1.46
+ $X2=0.625 $Y2=1.46
r123 56 75 4.19663 $w=1.95e-07 $l=1.4e-07 $layer=LI1_cond $X=3.64 $Y=2.022
+ $X2=3.5 $Y2=2.022
r124 55 75 21.6131 $w=1.93e-07 $l=3.8e-07 $layer=LI1_cond $X=3.12 $Y=2.022
+ $X2=3.5 $Y2=2.022
r125 54 55 27.3007 $w=1.93e-07 $l=4.8e-07 $layer=LI1_cond $X=2.64 $Y=2.022
+ $X2=3.12 $Y2=2.022
r126 53 54 27.3007 $w=1.93e-07 $l=4.8e-07 $layer=LI1_cond $X=2.16 $Y=2.022
+ $X2=2.64 $Y2=2.022
r127 52 53 27.3007 $w=1.93e-07 $l=4.8e-07 $layer=LI1_cond $X=1.68 $Y=2.022
+ $X2=2.16 $Y2=2.022
r128 52 76 6.82517 $w=1.93e-07 $l=1.2e-07 $layer=LI1_cond $X=1.68 $Y=2.022
+ $X2=1.56 $Y2=2.022
r129 51 76 5.7603 $w=1.95e-07 $l=2.23e-07 $layer=LI1_cond $X=1.337 $Y=2.022
+ $X2=1.56 $Y2=2.022
r130 50 70 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=1.395 $Y=1.46
+ $X2=1.485 $Y2=1.46
r131 50 68 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.395 $Y=1.46
+ $X2=1.055 $Y2=1.46
r132 49 50 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.395
+ $Y=1.46 $X2=1.395 $Y2=1.46
r133 46 74 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.655 $Y=1.51
+ $X2=3.655 $Y2=1.675
r134 46 73 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.655 $Y=1.51
+ $X2=3.655 $Y2=1.345
r135 45 46 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.655
+ $Y=1.51 $X2=3.655 $Y2=1.51
r136 43 56 2.90766 $w=2.8e-07 $l=9.7e-08 $layer=LI1_cond $X=3.64 $Y=1.925
+ $X2=3.64 $Y2=2.022
r137 43 45 17.0809 $w=2.78e-07 $l=4.15e-07 $layer=LI1_cond $X=3.64 $Y=1.925
+ $X2=3.64 $Y2=1.51
r138 42 51 2.5056 $w=4.45e-07 $l=9.7e-08 $layer=LI1_cond $X=1.337 $Y=1.925
+ $X2=1.337 $Y2=2.022
r139 41 49 2.8409 $w=4.45e-07 $l=1.43e-07 $layer=LI1_cond $X=1.337 $Y=1.63
+ $X2=1.337 $Y2=1.487
r140 41 42 7.63979 $w=4.43e-07 $l=2.95e-07 $layer=LI1_cond $X=1.337 $Y=1.63
+ $X2=1.337 $Y2=1.925
r141 40 68 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.715 $Y=1.46
+ $X2=1.055 $Y2=1.46
r142 40 66 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=0.715 $Y=1.46
+ $X2=0.625 $Y2=1.46
r143 39 40 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.715
+ $Y=1.46 $X2=0.715 $Y2=1.46
r144 36 63 30.6007 $w=3.3e-07 $l=1.75e-07 $layer=POLY_cond $X=0.375 $Y=1.46
+ $X2=0.55 $Y2=1.46
r145 35 39 13.7484 $w=2.83e-07 $l=3.4e-07 $layer=LI1_cond $X=0.375 $Y=1.487
+ $X2=0.715 $Y2=1.487
r146 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.375
+ $Y=1.46 $X2=0.375 $Y2=1.46
r147 33 49 4.41035 $w=2.85e-07 $l=2.22e-07 $layer=LI1_cond $X=1.115 $Y=1.487
+ $X2=1.337 $Y2=1.487
r148 33 39 16.1746 $w=2.83e-07 $l=4e-07 $layer=LI1_cond $X=1.115 $Y=1.487
+ $X2=0.715 $Y2=1.487
r149 31 73 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.645 $Y=0.655
+ $X2=3.645 $Y2=1.345
r150 27 74 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.635 $Y=2.465
+ $X2=3.635 $Y2=1.675
r151 21 70 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.485 $Y=1.625
+ $X2=1.485 $Y2=1.46
r152 21 23 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=1.485 $Y=1.625
+ $X2=1.485 $Y2=2.465
r153 17 70 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.485 $Y=1.295
+ $X2=1.485 $Y2=1.46
r154 17 19 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=1.485 $Y=1.295
+ $X2=1.485 $Y2=0.655
r155 13 68 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.055 $Y=1.625
+ $X2=1.055 $Y2=1.46
r156 13 15 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=1.055 $Y=1.625
+ $X2=1.055 $Y2=2.465
r157 9 68 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.055 $Y=1.295
+ $X2=1.055 $Y2=1.46
r158 9 11 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=1.055 $Y=1.295
+ $X2=1.055 $Y2=0.655
r159 5 66 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.625 $Y=1.625
+ $X2=0.625 $Y2=1.46
r160 5 7 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=0.625 $Y=1.625
+ $X2=0.625 $Y2=2.465
r161 1 66 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.625 $Y=1.295
+ $X2=0.625 $Y2=1.46
r162 1 3 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=0.625 $Y=1.295
+ $X2=0.625 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__O211AI_4%A2 3 5 7 10 12 14 17 19 21 24 26 28 29 30
+ 31 45
r80 43 45 24.1488 $w=3.8e-07 $l=1.65e-07 $layer=POLY_cond $X=3.04 $Y=1.535
+ $X2=3.205 $Y2=1.535
r81 43 44 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.04
+ $Y=1.51 $X2=3.04 $Y2=1.51
r82 41 43 38.7844 $w=3.8e-07 $l=2.65e-07 $layer=POLY_cond $X=2.775 $Y=1.535
+ $X2=3.04 $Y2=1.535
r83 40 41 62.9332 $w=3.8e-07 $l=4.3e-07 $layer=POLY_cond $X=2.345 $Y=1.535
+ $X2=2.775 $Y2=1.535
r84 38 40 47.5658 $w=3.8e-07 $l=3.25e-07 $layer=POLY_cond $X=2.02 $Y=1.535
+ $X2=2.345 $Y2=1.535
r85 38 39 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.02
+ $Y=1.51 $X2=2.02 $Y2=1.51
r86 35 38 15.3674 $w=3.8e-07 $l=1.05e-07 $layer=POLY_cond $X=1.915 $Y=1.535
+ $X2=2.02 $Y2=1.535
r87 31 44 2.83678 $w=3.23e-07 $l=8e-08 $layer=LI1_cond $X=3.12 $Y=1.587 $X2=3.04
+ $Y2=1.587
r88 30 44 14.1839 $w=3.23e-07 $l=4e-07 $layer=LI1_cond $X=2.64 $Y=1.587 $X2=3.04
+ $Y2=1.587
r89 29 30 17.0207 $w=3.23e-07 $l=4.8e-07 $layer=LI1_cond $X=2.16 $Y=1.587
+ $X2=2.64 $Y2=1.587
r90 29 39 4.96437 $w=3.23e-07 $l=1.4e-07 $layer=LI1_cond $X=2.16 $Y=1.587
+ $X2=2.02 $Y2=1.587
r91 26 45 24.6126 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=3.205 $Y=1.725
+ $X2=3.205 $Y2=1.535
r92 26 28 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=3.205 $Y=1.725
+ $X2=3.205 $Y2=2.465
r93 22 45 24.6126 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=3.205 $Y=1.345
+ $X2=3.205 $Y2=1.535
r94 22 24 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.205 $Y=1.345
+ $X2=3.205 $Y2=0.655
r95 19 41 24.6126 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=2.775 $Y=1.725
+ $X2=2.775 $Y2=1.535
r96 19 21 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=2.775 $Y=1.725
+ $X2=2.775 $Y2=2.465
r97 15 41 24.6126 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=2.775 $Y=1.345
+ $X2=2.775 $Y2=1.535
r98 15 17 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.775 $Y=1.345
+ $X2=2.775 $Y2=0.655
r99 12 40 24.6126 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=2.345 $Y=1.725
+ $X2=2.345 $Y2=1.535
r100 12 14 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=2.345 $Y=1.725
+ $X2=2.345 $Y2=2.465
r101 8 40 24.6126 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=2.345 $Y=1.345
+ $X2=2.345 $Y2=1.535
r102 8 10 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=2.345 $Y=1.345
+ $X2=2.345 $Y2=0.655
r103 5 35 24.6126 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=1.915 $Y=1.725
+ $X2=1.915 $Y2=1.535
r104 5 7 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=1.915 $Y=1.725
+ $X2=1.915 $Y2=2.465
r105 1 35 24.6126 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=1.915 $Y=1.345
+ $X2=1.915 $Y2=1.535
r106 1 3 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.915 $Y=1.345
+ $X2=1.915 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__O211AI_4%B1 3 7 11 15 19 23 27 31 33 34 35 36 39 40
+ 42 43 44 58
r126 56 58 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=4.875 $Y=1.51
+ $X2=4.965 $Y2=1.51
r127 56 57 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=4.875
+ $Y=1.51 $X2=4.875 $Y2=1.51
r128 54 56 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=4.535 $Y=1.51
+ $X2=4.875 $Y2=1.51
r129 52 54 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=4.195 $Y=1.51
+ $X2=4.535 $Y2=1.51
r130 52 53 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=4.195
+ $Y=1.51 $X2=4.195 $Y2=1.51
r131 49 52 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=4.105 $Y=1.51
+ $X2=4.195 $Y2=1.51
r132 44 57 2.66204 $w=5.83e-07 $l=8e-08 $layer=LI1_cond $X=4.955 $Y=1.552
+ $X2=4.875 $Y2=1.552
r133 43 57 8.74746 $w=4.13e-07 $l=3.15e-07 $layer=LI1_cond $X=4.56 $Y=1.552
+ $X2=4.875 $Y2=1.552
r134 43 53 10.1359 $w=4.13e-07 $l=3.65e-07 $layer=LI1_cond $X=4.56 $Y=1.552
+ $X2=4.195 $Y2=1.552
r135 42 53 3.19352 $w=4.13e-07 $l=1.15e-07 $layer=LI1_cond $X=4.08 $Y=1.552
+ $X2=4.195 $Y2=1.552
r136 40 62 16.3138 $w=3.25e-07 $l=1.1e-07 $layer=POLY_cond $X=7.555 $Y=1.51
+ $X2=7.665 $Y2=1.51
r137 40 60 14.8308 $w=3.25e-07 $l=1e-07 $layer=POLY_cond $X=7.555 $Y=1.51
+ $X2=7.455 $Y2=1.51
r138 39 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.555
+ $Y=1.51 $X2=7.555 $Y2=1.51
r139 37 39 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=7.555 $Y=1.93
+ $X2=7.555 $Y2=1.51
r140 35 37 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=7.39 $Y=2.015
+ $X2=7.555 $Y2=1.93
r141 35 36 147.77 $w=1.68e-07 $l=2.265e-06 $layer=LI1_cond $X=7.39 $Y=2.015
+ $X2=5.125 $Y2=2.015
r142 34 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.04 $Y=1.93
+ $X2=5.125 $Y2=2.015
r143 33 44 6.03523 $w=1.7e-07 $l=2.08e-07 $layer=LI1_cond $X=5.04 $Y=1.76
+ $X2=5.04 $Y2=1.552
r144 33 34 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=5.04 $Y=1.76
+ $X2=5.04 $Y2=1.93
r145 29 62 20.86 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.665 $Y=1.345
+ $X2=7.665 $Y2=1.51
r146 29 31 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=7.665 $Y=1.345
+ $X2=7.665 $Y2=0.765
r147 25 60 20.86 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.455 $Y=1.675
+ $X2=7.455 $Y2=1.51
r148 25 27 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=7.455 $Y=1.675
+ $X2=7.455 $Y2=2.465
r149 21 58 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.965 $Y=1.675
+ $X2=4.965 $Y2=1.51
r150 21 23 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=4.965 $Y=1.675
+ $X2=4.965 $Y2=2.465
r151 17 58 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.965 $Y=1.345
+ $X2=4.965 $Y2=1.51
r152 17 19 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=4.965 $Y=1.345
+ $X2=4.965 $Y2=0.655
r153 13 54 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.535 $Y=1.675
+ $X2=4.535 $Y2=1.51
r154 13 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=4.535 $Y=1.675
+ $X2=4.535 $Y2=2.465
r155 9 54 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.535 $Y=1.345
+ $X2=4.535 $Y2=1.51
r156 9 11 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=4.535 $Y=1.345
+ $X2=4.535 $Y2=0.655
r157 5 49 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.105 $Y=1.675
+ $X2=4.105 $Y2=1.51
r158 5 7 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=4.105 $Y=1.675
+ $X2=4.105 $Y2=2.465
r159 1 49 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.105 $Y=1.345
+ $X2=4.105 $Y2=1.51
r160 1 3 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=4.105 $Y=1.345
+ $X2=4.105 $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__O211AI_4%C1 3 7 11 15 19 23 27 31 33 34 35 36 56
r77 56 57 7.41538 $w=3.25e-07 $l=5e-08 $layer=POLY_cond $X=7.025 $Y=1.51
+ $X2=7.075 $Y2=1.51
r78 54 56 21.5046 $w=3.25e-07 $l=1.45e-07 $layer=POLY_cond $X=6.88 $Y=1.51
+ $X2=7.025 $Y2=1.51
r79 54 55 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.88
+ $Y=1.51 $X2=6.88 $Y2=1.51
r80 52 54 34.8523 $w=3.25e-07 $l=2.35e-07 $layer=POLY_cond $X=6.645 $Y=1.51
+ $X2=6.88 $Y2=1.51
r81 51 52 57.84 $w=3.25e-07 $l=3.9e-07 $layer=POLY_cond $X=6.255 $Y=1.51
+ $X2=6.645 $Y2=1.51
r82 49 51 8.15692 $w=3.25e-07 $l=5.5e-08 $layer=POLY_cond $X=6.2 $Y=1.51
+ $X2=6.255 $Y2=1.51
r83 49 50 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.2 $Y=1.51
+ $X2=6.2 $Y2=1.51
r84 47 49 21.5046 $w=3.25e-07 $l=1.45e-07 $layer=POLY_cond $X=6.055 $Y=1.51
+ $X2=6.2 $Y2=1.51
r85 46 47 34.1108 $w=3.25e-07 $l=2.3e-07 $layer=POLY_cond $X=5.825 $Y=1.51
+ $X2=6.055 $Y2=1.51
r86 45 46 29.6615 $w=3.25e-07 $l=2e-07 $layer=POLY_cond $X=5.625 $Y=1.51
+ $X2=5.825 $Y2=1.51
r87 43 45 15.5723 $w=3.25e-07 $l=1.05e-07 $layer=POLY_cond $X=5.52 $Y=1.51
+ $X2=5.625 $Y2=1.51
r88 41 43 18.5385 $w=3.25e-07 $l=1.25e-07 $layer=POLY_cond $X=5.395 $Y=1.51
+ $X2=5.52 $Y2=1.51
r89 36 55 2.7521 $w=3.33e-07 $l=8e-08 $layer=LI1_cond $X=6.96 $Y=1.592 $X2=6.88
+ $Y2=1.592
r90 35 55 13.7605 $w=3.33e-07 $l=4e-07 $layer=LI1_cond $X=6.48 $Y=1.592 $X2=6.88
+ $Y2=1.592
r91 35 50 9.63236 $w=3.33e-07 $l=2.8e-07 $layer=LI1_cond $X=6.48 $Y=1.592
+ $X2=6.2 $Y2=1.592
r92 34 50 6.88026 $w=3.33e-07 $l=2e-07 $layer=LI1_cond $X=6 $Y=1.592 $X2=6.2
+ $Y2=1.592
r93 33 34 16.5126 $w=3.33e-07 $l=4.8e-07 $layer=LI1_cond $X=5.52 $Y=1.592 $X2=6
+ $Y2=1.592
r94 33 43 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.52
+ $Y=1.51 $X2=5.52 $Y2=1.51
r95 29 57 20.86 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.075 $Y=1.345
+ $X2=7.075 $Y2=1.51
r96 29 31 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=7.075 $Y=1.345
+ $X2=7.075 $Y2=0.765
r97 25 56 20.86 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.025 $Y=1.675
+ $X2=7.025 $Y2=1.51
r98 25 27 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=7.025 $Y=1.675
+ $X2=7.025 $Y2=2.465
r99 21 52 20.86 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.645 $Y=1.345
+ $X2=6.645 $Y2=1.51
r100 21 23 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=6.645 $Y=1.345
+ $X2=6.645 $Y2=0.765
r101 17 51 20.86 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.255 $Y=1.675
+ $X2=6.255 $Y2=1.51
r102 17 19 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=6.255 $Y=1.675
+ $X2=6.255 $Y2=2.465
r103 13 47 20.86 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.055 $Y=1.345
+ $X2=6.055 $Y2=1.51
r104 13 15 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=6.055 $Y=1.345
+ $X2=6.055 $Y2=0.765
r105 9 46 20.86 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.825 $Y=1.675
+ $X2=5.825 $Y2=1.51
r106 9 11 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=5.825 $Y=1.675
+ $X2=5.825 $Y2=2.465
r107 5 45 20.86 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.625 $Y=1.345
+ $X2=5.625 $Y2=1.51
r108 5 7 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=5.625 $Y=1.345
+ $X2=5.625 $Y2=0.765
r109 1 41 20.86 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.395 $Y=1.675
+ $X2=5.395 $Y2=1.51
r110 1 3 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=5.395 $Y=1.675
+ $X2=5.395 $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__O211AI_4%VPWR 1 2 3 4 5 6 7 22 24 30 34 38 40 44 48
+ 51 52 53 54 56 57 58 60 75 85 86 92 95 98
r125 101 102 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.48 $Y=3.33
+ $X2=6.48 $Y2=3.33
r126 98 101 9.37226 $w=6.68e-07 $l=5.25e-07 $layer=LI1_cond $X=6.64 $Y=2.805
+ $X2=6.64 $Y2=3.33
r127 95 96 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.52 $Y=3.33
+ $X2=5.52 $Y2=3.33
r128 92 93 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r129 89 90 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r130 85 86 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.92 $Y=3.33
+ $X2=7.92 $Y2=3.33
r131 83 86 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=7.92 $Y2=3.33
r132 83 102 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=7.44 $Y=3.33
+ $X2=6.48 $Y2=3.33
r133 82 83 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.44 $Y=3.33
+ $X2=7.44 $Y2=3.33
r134 80 101 9.03384 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=6.975 $Y=3.33
+ $X2=6.64 $Y2=3.33
r135 80 82 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=6.975 $Y=3.33
+ $X2=7.44 $Y2=3.33
r136 79 102 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33
+ $X2=6.48 $Y2=3.33
r137 79 96 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=6 $Y=3.33 $X2=5.52
+ $Y2=3.33
r138 78 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6 $Y=3.33 $X2=6
+ $Y2=3.33
r139 76 95 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.73 $Y=3.33
+ $X2=5.605 $Y2=3.33
r140 76 78 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=5.73 $Y=3.33 $X2=6
+ $Y2=3.33
r141 75 101 9.03384 $w=1.7e-07 $l=3.35e-07 $layer=LI1_cond $X=6.305 $Y=3.33
+ $X2=6.64 $Y2=3.33
r142 75 78 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=6.305 $Y=3.33
+ $X2=6 $Y2=3.33
r143 74 96 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.52 $Y2=3.33
r144 73 74 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r145 70 71 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.6 $Y=3.33
+ $X2=3.6 $Y2=3.33
r146 68 71 0.535171 $w=4.9e-07 $l=1.92e-06 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=3.6 $Y2=3.33
r147 68 93 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r148 67 70 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=1.68 $Y=3.33
+ $X2=3.6 $Y2=3.33
r149 67 68 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r150 65 92 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.435 $Y=3.33
+ $X2=1.27 $Y2=3.33
r151 65 67 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=1.435 $Y=3.33
+ $X2=1.68 $Y2=3.33
r152 64 93 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r153 64 90 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=0.24 $Y2=3.33
r154 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r155 61 89 4.18769 $w=1.7e-07 $l=2.68e-07 $layer=LI1_cond $X=0.535 $Y=3.33
+ $X2=0.267 $Y2=3.33
r156 61 63 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=0.535 $Y=3.33
+ $X2=0.72 $Y2=3.33
r157 60 92 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.105 $Y=3.33
+ $X2=1.27 $Y2=3.33
r158 60 63 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=1.105 $Y=3.33
+ $X2=0.72 $Y2=3.33
r159 58 74 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r160 58 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.6 $Y2=3.33
r161 56 82 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=7.505 $Y=3.33
+ $X2=7.44 $Y2=3.33
r162 56 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.505 $Y=3.33
+ $X2=7.67 $Y2=3.33
r163 55 85 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=7.835 $Y=3.33
+ $X2=7.92 $Y2=3.33
r164 55 57 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.835 $Y=3.33
+ $X2=7.67 $Y2=3.33
r165 53 73 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=4.585 $Y=3.33
+ $X2=4.56 $Y2=3.33
r166 53 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.585 $Y=3.33
+ $X2=4.75 $Y2=3.33
r167 51 70 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=3.705 $Y=3.33
+ $X2=3.6 $Y2=3.33
r168 51 52 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.705 $Y=3.33
+ $X2=3.87 $Y2=3.33
r169 50 73 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=4.035 $Y=3.33
+ $X2=4.56 $Y2=3.33
r170 50 52 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.035 $Y=3.33
+ $X2=3.87 $Y2=3.33
r171 46 57 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.67 $Y=3.245
+ $X2=7.67 $Y2=3.33
r172 46 48 14.6675 $w=3.28e-07 $l=4.2e-07 $layer=LI1_cond $X=7.67 $Y=3.245
+ $X2=7.67 $Y2=2.825
r173 42 95 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.605 $Y=3.245
+ $X2=5.605 $Y2=3.33
r174 42 44 21.6659 $w=2.48e-07 $l=4.7e-07 $layer=LI1_cond $X=5.605 $Y=3.245
+ $X2=5.605 $Y2=2.775
r175 41 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.915 $Y=3.33
+ $X2=4.75 $Y2=3.33
r176 40 95 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.48 $Y=3.33
+ $X2=5.605 $Y2=3.33
r177 40 41 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=5.48 $Y=3.33
+ $X2=4.915 $Y2=3.33
r178 36 54 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.75 $Y=3.245
+ $X2=4.75 $Y2=3.33
r179 36 38 17.4613 $w=3.28e-07 $l=5e-07 $layer=LI1_cond $X=4.75 $Y=3.245
+ $X2=4.75 $Y2=2.745
r180 32 52 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.87 $Y=3.245
+ $X2=3.87 $Y2=3.33
r181 32 34 15.3659 $w=3.28e-07 $l=4.4e-07 $layer=LI1_cond $X=3.87 $Y=3.245
+ $X2=3.87 $Y2=2.805
r182 28 92 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.27 $Y=3.245
+ $X2=1.27 $Y2=3.33
r183 28 30 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=1.27 $Y=3.245
+ $X2=1.27 $Y2=2.815
r184 24 27 38.5472 $w=2.88e-07 $l=9.7e-07 $layer=LI1_cond $X=0.39 $Y=1.98
+ $X2=0.39 $Y2=2.95
r185 22 89 3.25015 $w=2.9e-07 $l=1.5995e-07 $layer=LI1_cond $X=0.39 $Y=3.245
+ $X2=0.267 $Y2=3.33
r186 22 27 11.7231 $w=2.88e-07 $l=2.95e-07 $layer=LI1_cond $X=0.39 $Y=3.245
+ $X2=0.39 $Y2=2.95
r187 7 48 600 $w=1.7e-07 $l=1.05769e-06 $layer=licon1_PDIFF $count=1 $X=7.53
+ $Y=1.835 $X2=7.67 $Y2=2.825
r188 6 98 300 $w=1.7e-07 $l=1.18596e-06 $layer=licon1_PDIFF $count=2 $X=6.33
+ $Y=1.835 $X2=6.81 $Y2=2.805
r189 5 44 600 $w=1.7e-07 $l=1.00757e-06 $layer=licon1_PDIFF $count=1 $X=5.47
+ $Y=1.835 $X2=5.61 $Y2=2.775
r190 4 38 600 $w=1.7e-07 $l=9.77497e-07 $layer=licon1_PDIFF $count=1 $X=4.61
+ $Y=1.835 $X2=4.75 $Y2=2.745
r191 3 34 600 $w=1.7e-07 $l=1.04695e-06 $layer=licon1_PDIFF $count=1 $X=3.71
+ $Y=1.835 $X2=3.87 $Y2=2.805
r192 2 30 600 $w=1.7e-07 $l=1.04766e-06 $layer=licon1_PDIFF $count=1 $X=1.13
+ $Y=1.835 $X2=1.27 $Y2=2.815
r193 1 27 400 $w=1.7e-07 $l=1.17584e-06 $layer=licon1_PDIFF $count=1 $X=0.285
+ $Y=1.835 $X2=0.41 $Y2=2.95
r194 1 24 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.285
+ $Y=1.835 $X2=0.41 $Y2=1.98
.ends

.subckt PM_SKY130_FD_SC_LP__O211AI_4%A_140_367# 1 2 3 4 15 19 21 22 28 34 35
r41 34 35 4.31602 $w=3.93e-07 $l=1.05e-07 $layer=LI1_cond $X=3.42 $Y=2.877
+ $X2=3.315 $Y2=2.877
r42 26 35 32.8338 $w=2.63e-07 $l=7.55e-07 $layer=LI1_cond $X=2.56 $Y=2.942
+ $X2=3.315 $Y2=2.942
r43 24 32 3.01344 $w=2.65e-07 $l=1e-07 $layer=LI1_cond $X=1.805 $Y=2.942
+ $X2=1.705 $Y2=2.942
r44 24 26 32.8338 $w=2.63e-07 $l=7.55e-07 $layer=LI1_cond $X=1.805 $Y=2.942
+ $X2=2.56 $Y2=2.942
r45 22 32 3.97773 $w=2e-07 $l=1.32e-07 $layer=LI1_cond $X=1.705 $Y=2.81
+ $X2=1.705 $Y2=2.942
r46 21 30 3.66916 $w=2e-07 $l=1.15e-07 $layer=LI1_cond $X=1.705 $Y=2.52
+ $X2=1.705 $Y2=2.405
r47 21 22 16.0818 $w=1.98e-07 $l=2.9e-07 $layer=LI1_cond $X=1.705 $Y=2.52
+ $X2=1.705 $Y2=2.81
r48 20 28 1.18299 $w=2.3e-07 $l=1.1e-07 $layer=LI1_cond $X=0.925 $Y=2.405
+ $X2=0.815 $Y2=2.405
r49 19 30 3.19058 $w=2.3e-07 $l=1e-07 $layer=LI1_cond $X=1.605 $Y=2.405
+ $X2=1.705 $Y2=2.405
r50 19 20 34.0722 $w=2.28e-07 $l=6.8e-07 $layer=LI1_cond $X=1.605 $Y=2.405
+ $X2=0.925 $Y2=2.405
r51 13 28 5.35987 $w=2.2e-07 $l=1.15e-07 $layer=LI1_cond $X=0.815 $Y=2.29
+ $X2=0.815 $Y2=2.405
r52 13 15 16.239 $w=2.18e-07 $l=3.1e-07 $layer=LI1_cond $X=0.815 $Y=2.29
+ $X2=0.815 $Y2=1.98
r53 4 34 600 $w=1.7e-07 $l=1.07773e-06 $layer=licon1_PDIFF $count=1 $X=3.28
+ $Y=1.835 $X2=3.42 $Y2=2.845
r54 3 26 600 $w=1.7e-07 $l=1.14787e-06 $layer=licon1_PDIFF $count=1 $X=2.42
+ $Y=1.835 $X2=2.56 $Y2=2.915
r55 2 32 600 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=1.56
+ $Y=1.835 $X2=1.7 $Y2=2.91
r56 2 30 600 $w=1.7e-07 $l=6.8644e-07 $layer=licon1_PDIFF $count=1 $X=1.56
+ $Y=1.835 $X2=1.7 $Y2=2.455
r57 1 28 300 $w=1.7e-07 $l=6.71361e-07 $layer=licon1_PDIFF $count=2 $X=0.7
+ $Y=1.835 $X2=0.84 $Y2=2.44
r58 1 15 600 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=0.7
+ $Y=1.835 $X2=0.84 $Y2=1.98
.ends

.subckt PM_SKY130_FD_SC_LP__O211AI_4%Y 1 2 3 4 5 6 7 8 25 33 35 39 41 49 51 55
+ 58 59 65 67 68 70 72 73 74 75 76 77
r104 75 76 23.5393 $w=2.33e-07 $l=4.8e-07 $layer=LI1_cond $X=6.48 $Y=2.387
+ $X2=6.96 $Y2=2.387
r105 75 82 16.9188 $w=2.33e-07 $l=3.45e-07 $layer=LI1_cond $X=6.48 $Y=2.387
+ $X2=6.135 $Y2=2.387
r106 74 82 5.8365 $w=2.02e-07 $l=1.18e-07 $layer=LI1_cond $X=6.017 $Y=2.387
+ $X2=6.135 $Y2=2.387
r107 73 77 22.0681 $w=2.33e-07 $l=4.5e-07 $layer=LI1_cond $X=7.89 $Y=2.387
+ $X2=7.44 $Y2=2.387
r108 70 76 9.07242 $w=2.33e-07 $l=1.85e-07 $layer=LI1_cond $X=7.145 $Y=2.387
+ $X2=6.96 $Y2=2.387
r109 70 72 4.31353 $w=2.35e-07 $l=9.5e-08 $layer=LI1_cond $X=7.145 $Y=2.387
+ $X2=7.24 $Y2=2.387
r110 69 77 5.14921 $w=2.33e-07 $l=1.05e-07 $layer=LI1_cond $X=7.335 $Y=2.387
+ $X2=7.44 $Y2=2.387
r111 69 72 4.31353 $w=2.35e-07 $l=9.5e-08 $layer=LI1_cond $X=7.335 $Y=2.387
+ $X2=7.24 $Y2=2.387
r112 59 62 3.4329 $w=2.08e-07 $l=6.5e-08 $layer=LI1_cond $X=2.13 $Y=2.4 $X2=2.13
+ $Y2=2.465
r113 58 73 6.97338 $w=2.35e-07 $l=1.55625e-07 $layer=LI1_cond $X=7.98 $Y=2.27
+ $X2=7.89 $Y2=2.387
r114 57 58 62.5404 $w=1.78e-07 $l=1.015e-06 $layer=LI1_cond $X=7.98 $Y=1.255
+ $X2=7.98 $Y2=2.27
r115 53 72 2.11804 $w=1.9e-07 $l=1.18e-07 $layer=LI1_cond $X=7.24 $Y=2.505
+ $X2=7.24 $Y2=2.387
r116 53 55 23.6411 $w=1.88e-07 $l=4.05e-07 $layer=LI1_cond $X=7.24 $Y=2.505
+ $X2=7.24 $Y2=2.91
r117 51 57 6.81649 $w=1.8e-07 $l=1.27279e-07 $layer=LI1_cond $X=7.89 $Y=1.165
+ $X2=7.98 $Y2=1.255
r118 51 68 53.298 $w=1.78e-07 $l=8.65e-07 $layer=LI1_cond $X=7.89 $Y=1.165
+ $X2=7.025 $Y2=1.165
r119 47 74 0.812465 $w=2.35e-07 $l=1.18e-07 $layer=LI1_cond $X=6.017 $Y=2.505
+ $X2=6.017 $Y2=2.387
r120 47 49 19.8613 $w=2.33e-07 $l=4.05e-07 $layer=LI1_cond $X=6.017 $Y=2.505
+ $X2=6.017 $Y2=2.91
r121 43 46 40.5342 $w=2.88e-07 $l=1.02e-06 $layer=LI1_cond $X=5.84 $Y=1.11
+ $X2=6.86 $Y2=1.11
r122 41 68 7.4104 $w=2.88e-07 $l=1.45e-07 $layer=LI1_cond $X=6.88 $Y=1.11
+ $X2=7.025 $Y2=1.11
r123 41 46 0.794788 $w=2.88e-07 $l=2e-08 $layer=LI1_cond $X=6.88 $Y=1.11
+ $X2=6.86 $Y2=1.11
r124 40 67 6.47928 $w=1.7e-07 $l=1.13e-07 $layer=LI1_cond $X=5.31 $Y=2.355
+ $X2=5.197 $Y2=2.355
r125 39 74 5.8365 $w=2.02e-07 $l=1.32034e-07 $layer=LI1_cond $X=5.9 $Y=2.355
+ $X2=6.017 $Y2=2.387
r126 39 40 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=5.9 $Y=2.355
+ $X2=5.31 $Y2=2.355
r127 36 65 3.27902 $w=1.7e-07 $l=2.504e-07 $layer=LI1_cond $X=4.425 $Y=2.355
+ $X2=4.205 $Y2=2.29
r128 35 67 6.47928 $w=1.7e-07 $l=1.12e-07 $layer=LI1_cond $X=5.085 $Y=2.355
+ $X2=5.197 $Y2=2.355
r129 35 36 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=5.085 $Y=2.355
+ $X2=4.425 $Y2=2.355
r130 31 65 2.82707 $w=2.1e-07 $l=1.24599e-07 $layer=LI1_cond $X=4.32 $Y=2.27
+ $X2=4.205 $Y2=2.29
r131 31 33 9.24242 $w=2.08e-07 $l=1.75e-07 $layer=LI1_cond $X=4.32 $Y=2.27
+ $X2=4.32 $Y2=2.095
r132 26 59 0.430812 $w=2.2e-07 $l=1.05e-07 $layer=LI1_cond $X=2.235 $Y=2.4
+ $X2=2.13 $Y2=2.4
r133 26 28 39.5497 $w=2.18e-07 $l=7.55e-07 $layer=LI1_cond $X=2.235 $Y=2.4
+ $X2=2.99 $Y2=2.4
r134 25 65 3.27902 $w=2.2e-07 $l=1.1e-07 $layer=LI1_cond $X=4.205 $Y=2.4
+ $X2=4.205 $Y2=2.29
r135 25 28 63.6463 $w=2.18e-07 $l=1.215e-06 $layer=LI1_cond $X=4.205 $Y=2.4
+ $X2=2.99 $Y2=2.4
r136 8 72 600 $w=1.7e-07 $l=6.0597e-07 $layer=licon1_PDIFF $count=1 $X=7.1
+ $Y=1.835 $X2=7.24 $Y2=2.375
r137 8 55 600 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=7.1
+ $Y=1.835 $X2=7.24 $Y2=2.91
r138 7 74 600 $w=1.7e-07 $l=5.85833e-07 $layer=licon1_PDIFF $count=1 $X=5.9
+ $Y=1.835 $X2=6.04 $Y2=2.355
r139 7 49 600 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=5.9
+ $Y=1.835 $X2=6.04 $Y2=2.91
r140 6 67 300 $w=1.7e-07 $l=5.90868e-07 $layer=licon1_PDIFF $count=2 $X=5.04
+ $Y=1.835 $X2=5.18 $Y2=2.36
r141 5 65 300 $w=1.7e-07 $l=7.36682e-07 $layer=licon1_PDIFF $count=2 $X=4.18
+ $Y=1.835 $X2=4.32 $Y2=2.505
r142 5 33 600 $w=1.7e-07 $l=3.2249e-07 $layer=licon1_PDIFF $count=1 $X=4.18
+ $Y=1.835 $X2=4.32 $Y2=2.095
r143 4 28 600 $w=1.7e-07 $l=6.3616e-07 $layer=licon1_PDIFF $count=1 $X=2.85
+ $Y=1.835 $X2=2.99 $Y2=2.405
r144 3 62 600 $w=1.7e-07 $l=6.96491e-07 $layer=licon1_PDIFF $count=1 $X=1.99
+ $Y=1.835 $X2=2.13 $Y2=2.465
r145 2 46 182 $w=1.7e-07 $l=7.81873e-07 $layer=licon1_NDIFF $count=1 $X=6.72
+ $Y=0.345 $X2=6.86 $Y2=1.06
r146 1 43 182 $w=1.7e-07 $l=7.81873e-07 $layer=licon1_NDIFF $count=1 $X=5.7
+ $Y=0.345 $X2=5.84 $Y2=1.06
.ends

.subckt PM_SKY130_FD_SC_LP__O211AI_4%A_57_47# 1 2 3 4 5 6 7 24 26 27 30 32 36 38
+ 42 44 48 50 52 53 54 56 57 58 59 63
r105 63 65 8.3814 $w=3.28e-07 $l=2.4e-07 $layer=LI1_cond $X=7.88 $Y=0.47
+ $X2=7.88 $Y2=0.71
r106 55 61 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=4.915 $Y=0.71
+ $X2=4.785 $Y2=0.71
r107 54 65 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.715 $Y=0.71
+ $X2=7.88 $Y2=0.71
r108 54 55 182.674 $w=1.68e-07 $l=2.8e-06 $layer=LI1_cond $X=7.715 $Y=0.71
+ $X2=4.915 $Y2=0.71
r109 52 61 2.85134 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=4.785 $Y=0.795
+ $X2=4.785 $Y2=0.71
r110 52 53 8.86495 $w=2.58e-07 $l=2e-07 $layer=LI1_cond $X=4.785 $Y=0.795
+ $X2=4.785 $Y2=0.995
r111 51 59 6.30264 $w=1.8e-07 $l=1.15e-07 $layer=LI1_cond $X=3.985 $Y=1.085
+ $X2=3.87 $Y2=1.085
r112 50 53 7.11373 $w=1.8e-07 $l=1.69115e-07 $layer=LI1_cond $X=4.655 $Y=1.085
+ $X2=4.785 $Y2=0.995
r113 50 51 41.2828 $w=1.78e-07 $l=6.7e-07 $layer=LI1_cond $X=4.655 $Y=1.085
+ $X2=3.985 $Y2=1.085
r114 46 59 0.47666 $w=2.3e-07 $l=9e-08 $layer=LI1_cond $X=3.87 $Y=0.995 $X2=3.87
+ $Y2=1.085
r115 46 48 28.8111 $w=2.28e-07 $l=5.75e-07 $layer=LI1_cond $X=3.87 $Y=0.995
+ $X2=3.87 $Y2=0.42
r116 45 58 5.40251 $w=1.8e-07 $l=9.5e-08 $layer=LI1_cond $X=3.085 $Y=1.085
+ $X2=2.99 $Y2=1.085
r117 44 59 6.30264 $w=1.8e-07 $l=1.15e-07 $layer=LI1_cond $X=3.755 $Y=1.085
+ $X2=3.87 $Y2=1.085
r118 44 45 41.2828 $w=1.78e-07 $l=6.7e-07 $layer=LI1_cond $X=3.755 $Y=1.085
+ $X2=3.085 $Y2=1.085
r119 40 58 1.14861 $w=1.9e-07 $l=9e-08 $layer=LI1_cond $X=2.99 $Y=0.995 $X2=2.99
+ $Y2=1.085
r120 40 42 33.5646 $w=1.88e-07 $l=5.75e-07 $layer=LI1_cond $X=2.99 $Y=0.995
+ $X2=2.99 $Y2=0.42
r121 39 57 5.40251 $w=1.8e-07 $l=9.5e-08 $layer=LI1_cond $X=2.225 $Y=1.085
+ $X2=2.13 $Y2=1.085
r122 38 58 5.40251 $w=1.8e-07 $l=9.5e-08 $layer=LI1_cond $X=2.895 $Y=1.085
+ $X2=2.99 $Y2=1.085
r123 38 39 41.2828 $w=1.78e-07 $l=6.7e-07 $layer=LI1_cond $X=2.895 $Y=1.085
+ $X2=2.225 $Y2=1.085
r124 34 57 1.14861 $w=1.9e-07 $l=9e-08 $layer=LI1_cond $X=2.13 $Y=0.995 $X2=2.13
+ $Y2=1.085
r125 34 36 33.5646 $w=1.88e-07 $l=5.75e-07 $layer=LI1_cond $X=2.13 $Y=0.995
+ $X2=2.13 $Y2=0.42
r126 33 56 5.40251 $w=1.8e-07 $l=9.5e-08 $layer=LI1_cond $X=1.365 $Y=1.085
+ $X2=1.27 $Y2=1.085
r127 32 57 5.40251 $w=1.8e-07 $l=9.5e-08 $layer=LI1_cond $X=2.035 $Y=1.085
+ $X2=2.13 $Y2=1.085
r128 32 33 41.2828 $w=1.78e-07 $l=6.7e-07 $layer=LI1_cond $X=2.035 $Y=1.085
+ $X2=1.365 $Y2=1.085
r129 28 56 1.14861 $w=1.9e-07 $l=9e-08 $layer=LI1_cond $X=1.27 $Y=0.995 $X2=1.27
+ $Y2=1.085
r130 28 30 33.5646 $w=1.88e-07 $l=5.75e-07 $layer=LI1_cond $X=1.27 $Y=0.995
+ $X2=1.27 $Y2=0.42
r131 26 56 5.40251 $w=1.8e-07 $l=9.5e-08 $layer=LI1_cond $X=1.175 $Y=1.085
+ $X2=1.27 $Y2=1.085
r132 26 27 41.2828 $w=1.78e-07 $l=6.7e-07 $layer=LI1_cond $X=1.175 $Y=1.085
+ $X2=0.505 $Y2=1.085
r133 22 27 6.84108 $w=1.8e-07 $l=1.3784e-07 $layer=LI1_cond $X=0.405 $Y=0.995
+ $X2=0.505 $Y2=1.085
r134 22 24 31.8864 $w=1.98e-07 $l=5.75e-07 $layer=LI1_cond $X=0.405 $Y=0.995
+ $X2=0.405 $Y2=0.42
r135 7 63 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=7.74
+ $Y=0.345 $X2=7.88 $Y2=0.47
r136 6 61 182 $w=1.7e-07 $l=6.21068e-07 $layer=licon1_NDIFF $count=1 $X=4.61
+ $Y=0.235 $X2=4.75 $Y2=0.79
r137 5 48 91 $w=1.7e-07 $l=2.48948e-07 $layer=licon1_NDIFF $count=2 $X=3.72
+ $Y=0.235 $X2=3.87 $Y2=0.42
r138 4 42 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=2.85
+ $Y=0.235 $X2=2.99 $Y2=0.42
r139 3 36 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=1.99
+ $Y=0.235 $X2=2.13 $Y2=0.42
r140 2 30 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=1.13
+ $Y=0.235 $X2=1.27 $Y2=0.42
r141 1 24 91 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=2 $X=0.285
+ $Y=0.235 $X2=0.41 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__O211AI_4%VGND 1 2 3 4 17 21 25 29 32 33 34 36 41 54
+ 55 58 61 64
r96 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r97 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.68 $Y=0 $X2=1.68
+ $Y2=0
r98 58 59 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r99 54 55 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=7.92 $Y=0 $X2=7.92
+ $Y2=0
r100 51 54 281.84 $w=1.68e-07 $l=4.32e-06 $layer=LI1_cond $X=3.6 $Y=0 $X2=7.92
+ $Y2=0
r101 51 52 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r102 49 52 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=3.6
+ $Y2=0
r103 49 65 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.64
+ $Y2=0
r104 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r105 46 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.725 $Y=0 $X2=2.56
+ $Y2=0
r106 46 48 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=2.725 $Y=0
+ $X2=3.12 $Y2=0
r107 45 65 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=2.64
+ $Y2=0
r108 45 62 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=1.68
+ $Y2=0
r109 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r110 42 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.865 $Y=0 $X2=1.7
+ $Y2=0
r111 42 44 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.865 $Y=0 $X2=2.16
+ $Y2=0
r112 41 64 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.395 $Y=0 $X2=2.56
+ $Y2=0
r113 41 44 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=2.395 $Y=0
+ $X2=2.16 $Y2=0
r114 40 62 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=1.68
+ $Y2=0
r115 40 59 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r116 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r117 37 58 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.005 $Y=0 $X2=0.84
+ $Y2=0
r118 37 39 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=1.005 $Y=0 $X2=1.2
+ $Y2=0
r119 36 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.535 $Y=0 $X2=1.7
+ $Y2=0
r120 36 39 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.535 $Y=0 $X2=1.2
+ $Y2=0
r121 34 55 1.07034 $w=4.9e-07 $l=3.84e-06 $layer=MET1_cond $X=4.08 $Y=0 $X2=7.92
+ $Y2=0
r122 34 52 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=0 $X2=3.6
+ $Y2=0
r123 32 48 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=3.255 $Y=0
+ $X2=3.12 $Y2=0
r124 32 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.255 $Y=0 $X2=3.42
+ $Y2=0
r125 31 51 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=3.585 $Y=0 $X2=3.6
+ $Y2=0
r126 31 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.585 $Y=0 $X2=3.42
+ $Y2=0
r127 27 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.42 $Y=0.085
+ $X2=3.42 $Y2=0
r128 27 29 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=3.42 $Y=0.085
+ $X2=3.42 $Y2=0.36
r129 23 64 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.56 $Y=0.085
+ $X2=2.56 $Y2=0
r130 23 25 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.56 $Y=0.085
+ $X2=2.56 $Y2=0.36
r131 19 61 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.7 $Y=0.085 $X2=1.7
+ $Y2=0
r132 19 21 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=1.7 $Y=0.085
+ $X2=1.7 $Y2=0.36
r133 15 58 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.84 $Y=0.085
+ $X2=0.84 $Y2=0
r134 15 17 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=0.84 $Y=0.085
+ $X2=0.84 $Y2=0.36
r135 4 29 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=3.28
+ $Y=0.235 $X2=3.42 $Y2=0.36
r136 3 25 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=2.42
+ $Y=0.235 $X2=2.56 $Y2=0.36
r137 2 21 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=1.56
+ $Y=0.235 $X2=1.7 $Y2=0.36
r138 1 17 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=0.7
+ $Y=0.235 $X2=0.84 $Y2=0.36
.ends

.subckt PM_SKY130_FD_SC_LP__O211AI_4%A_836_47# 1 2 3 4 21 24
r32 19 21 59.5407 $w=1.88e-07 $l=1.02e-06 $layer=LI1_cond $X=6.35 $Y=0.36
+ $X2=7.37 $Y2=0.36
r33 17 19 61.5837 $w=1.88e-07 $l=1.055e-06 $layer=LI1_cond $X=5.295 $Y=0.36
+ $X2=6.35 $Y2=0.36
r34 15 24 4.74669 $w=1.9e-07 $l=1.65e-07 $layer=LI1_cond $X=4.485 $Y=0.36
+ $X2=4.32 $Y2=0.36
r35 15 17 47.2823 $w=1.88e-07 $l=8.1e-07 $layer=LI1_cond $X=4.485 $Y=0.36
+ $X2=5.295 $Y2=0.36
r36 4 21 182 $w=1.7e-07 $l=2.27376e-07 $layer=licon1_NDIFF $count=1 $X=7.15
+ $Y=0.345 $X2=7.37 $Y2=0.36
r37 3 19 182 $w=1.7e-07 $l=2.27376e-07 $layer=licon1_NDIFF $count=1 $X=6.13
+ $Y=0.345 $X2=6.35 $Y2=0.36
r38 2 17 182 $w=1.7e-07 $l=3.11288e-07 $layer=licon1_NDIFF $count=1 $X=5.04
+ $Y=0.235 $X2=5.295 $Y2=0.36
r39 1 24 91 $w=1.7e-07 $l=1.96214e-07 $layer=licon1_NDIFF $count=2 $X=4.18
+ $Y=0.235 $X2=4.32 $Y2=0.37
.ends

