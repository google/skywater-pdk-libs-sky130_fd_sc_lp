# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__a31oi_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_lp__a31oi_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.800000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.960000 1.425000 3.335000 1.750000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.625000 1.210000 1.635000 1.545000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 1.210000 0.455000 1.545000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.505000 1.425000 4.715000 1.750000 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  1.037400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.335000 0.605000 2.675000 1.085000 ;
        RECT 2.335000 1.085000 4.465000 1.255000 ;
        RECT 2.335000 1.255000 2.790000 1.950000 ;
        RECT 2.335000 1.950000 4.035000 2.130000 ;
        RECT 3.345000 0.325000 3.535000 1.085000 ;
        RECT 3.705000 2.130000 4.035000 2.735000 ;
        RECT 4.205000 0.325000 4.465000 1.085000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 4.800000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 4.800000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.800000 0.085000 ;
      RECT 0.000000  3.245000 4.800000 3.415000 ;
      RECT 0.095000  0.335000 0.345000 0.870000 ;
      RECT 0.095000  0.870000 2.145000 1.040000 ;
      RECT 0.095000  1.715000 2.165000 1.885000 ;
      RECT 0.095000  1.885000 0.355000 3.075000 ;
      RECT 0.525000  0.085000 0.855000 0.700000 ;
      RECT 0.525000  2.055000 0.855000 3.245000 ;
      RECT 1.025000  0.335000 1.255000 0.870000 ;
      RECT 1.025000  1.885000 1.260000 3.075000 ;
      RECT 1.425000  0.255000 3.175000 0.435000 ;
      RECT 1.425000  0.435000 1.645000 0.700000 ;
      RECT 1.430000  2.055000 1.760000 3.245000 ;
      RECT 1.815000  0.605000 2.145000 0.870000 ;
      RECT 1.815000  1.040000 2.145000 1.205000 ;
      RECT 1.930000  1.885000 2.165000 2.300000 ;
      RECT 1.930000  2.300000 3.535000 2.470000 ;
      RECT 1.930000  2.470000 2.155000 3.075000 ;
      RECT 2.325000  2.640000 3.175000 3.245000 ;
      RECT 2.845000  0.435000 3.175000 0.915000 ;
      RECT 3.345000  2.470000 3.535000 2.905000 ;
      RECT 3.345000  2.905000 4.465000 3.075000 ;
      RECT 3.705000  0.085000 4.035000 0.915000 ;
      RECT 4.205000  1.920000 4.465000 2.905000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
  END
END sky130_fd_sc_lp__a31oi_2
END LIBRARY
