# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__ebufn_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_lp__ebufn_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.240000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.315000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.405000 1.345000 5.805000 1.780000 ;
    END
  END A
  PIN TE_B
    ANTENNAGATEAREA  1.071000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.485000 1.180000 4.770000 1.410000 ;
        RECT 4.440000 1.410000 4.770000 1.595000 ;
    END
  END TE_B
  PIN Z
    ANTENNADIFFAREA  1.323000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 1.180000 0.705000 1.410000 ;
        RECT 0.535000 0.595000 0.875000 0.975000 ;
        RECT 0.535000 0.975000 1.875000 1.145000 ;
        RECT 0.535000 1.145000 0.705000 1.180000 ;
        RECT 0.535000 1.410000 0.705000 1.815000 ;
        RECT 0.535000 1.815000 1.875000 1.985000 ;
        RECT 0.535000 1.985000 0.875000 2.735000 ;
        RECT 1.545000 0.595000 1.875000 0.975000 ;
        RECT 1.545000 1.985000 1.875000 2.735000 ;
    END
  END Z
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 6.240000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 6.240000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.240000 0.085000 ;
      RECT 0.000000  3.245000 6.240000 3.415000 ;
      RECT 0.115000  0.255000 2.225000 0.425000 ;
      RECT 0.115000  0.425000 0.365000 1.010000 ;
      RECT 0.115000  1.815000 0.365000 2.905000 ;
      RECT 0.115000  2.905000 2.375000 3.075000 ;
      RECT 0.875000  1.315000 1.885000 1.475000 ;
      RECT 0.875000  1.475000 2.215000 1.645000 ;
      RECT 1.045000  0.425000 1.375000 0.805000 ;
      RECT 1.045000  2.155000 1.375000 2.905000 ;
      RECT 2.045000  1.645000 2.215000 2.015000 ;
      RECT 2.045000  2.015000 4.495000 2.185000 ;
      RECT 2.045000  2.355000 3.375000 2.525000 ;
      RECT 2.045000  2.525000 2.375000 2.905000 ;
      RECT 2.055000  0.425000 2.225000 1.135000 ;
      RECT 2.055000  1.135000 3.085000 1.305000 ;
      RECT 2.405000  0.085000 2.735000 0.965000 ;
      RECT 2.545000  2.695000 2.875000 3.245000 ;
      RECT 2.915000  0.255000 3.085000 0.840000 ;
      RECT 2.915000  0.840000 4.025000 1.010000 ;
      RECT 2.915000  1.010000 3.085000 1.135000 ;
      RECT 3.045000  2.525000 4.415000 2.695000 ;
      RECT 3.045000  2.695000 3.375000 3.075000 ;
      RECT 3.265000  0.085000 3.515000 0.670000 ;
      RECT 3.545000  2.865000 3.875000 3.245000 ;
      RECT 3.695000  0.255000 4.025000 0.840000 ;
      RECT 4.085000  2.695000 4.415000 3.075000 ;
      RECT 4.195000  0.340000 5.110000 1.010000 ;
      RECT 4.325000  2.185000 6.145000 2.355000 ;
      RECT 4.665000  1.765000 5.110000 2.015000 ;
      RECT 4.780000  0.255000 5.110000 0.340000 ;
      RECT 4.940000  1.010000 5.110000 1.765000 ;
      RECT 5.210000  2.525000 5.540000 3.245000 ;
      RECT 5.280000  0.085000 5.610000 1.135000 ;
      RECT 5.710000  1.950000 6.145000 2.185000 ;
      RECT 5.710000  2.355000 6.145000 3.075000 ;
      RECT 5.780000  0.255000 6.145000 1.135000 ;
      RECT 5.975000  1.135000 6.145000 1.950000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
  END
END sky130_fd_sc_lp__ebufn_4
END LIBRARY
