* File: sky130_fd_sc_lp__a2111o_0.pxi.spice
* Created: Fri Aug 28 09:45:42 2020
* 
x_PM_SKY130_FD_SC_LP__A2111O_0%A_80_159# N_A_80_159#_M1001_d N_A_80_159#_M1004_d
+ N_A_80_159#_M1002_s N_A_80_159#_c_91_n N_A_80_159#_M1005_g N_A_80_159#_M1008_g
+ N_A_80_159#_c_94_n N_A_80_159#_c_95_n N_A_80_159#_c_96_n N_A_80_159#_c_97_n
+ N_A_80_159#_c_105_n N_A_80_159#_c_106_n N_A_80_159#_c_107_n N_A_80_159#_c_98_n
+ N_A_80_159#_c_99_n N_A_80_159#_c_100_n N_A_80_159#_c_101_n N_A_80_159#_c_102_n
+ PM_SKY130_FD_SC_LP__A2111O_0%A_80_159#
x_PM_SKY130_FD_SC_LP__A2111O_0%D1 N_D1_M1001_g N_D1_c_181_n N_D1_c_182_n
+ N_D1_M1002_g N_D1_c_178_n N_D1_c_184_n N_D1_c_185_n D1 D1 N_D1_c_180_n
+ PM_SKY130_FD_SC_LP__A2111O_0%D1
x_PM_SKY130_FD_SC_LP__A2111O_0%C1 N_C1_M1007_g N_C1_c_232_n N_C1_M1009_g
+ N_C1_c_233_n N_C1_c_239_n C1 C1 C1 C1 C1 N_C1_c_235_n N_C1_c_236_n
+ PM_SKY130_FD_SC_LP__A2111O_0%C1
x_PM_SKY130_FD_SC_LP__A2111O_0%B1 N_B1_M1003_g N_B1_M1004_g N_B1_c_287_n
+ N_B1_c_292_n B1 B1 B1 B1 N_B1_c_289_n B1 PM_SKY130_FD_SC_LP__A2111O_0%B1
x_PM_SKY130_FD_SC_LP__A2111O_0%A1 N_A1_c_338_n N_A1_c_339_n N_A1_M1010_g
+ N_A1_M1006_g N_A1_c_341_n A1 A1 A1 PM_SKY130_FD_SC_LP__A2111O_0%A1
x_PM_SKY130_FD_SC_LP__A2111O_0%A2 N_A2_c_389_n N_A2_M1011_g N_A2_M1000_g
+ N_A2_c_390_n N_A2_c_391_n N_A2_c_397_n N_A2_c_392_n A2 A2 A2 N_A2_c_394_n
+ PM_SKY130_FD_SC_LP__A2111O_0%A2
x_PM_SKY130_FD_SC_LP__A2111O_0%X N_X_M1008_s N_X_M1005_s X X X X X X X
+ N_X_c_428_n PM_SKY130_FD_SC_LP__A2111O_0%X
x_PM_SKY130_FD_SC_LP__A2111O_0%VPWR N_VPWR_M1005_d N_VPWR_M1006_d N_VPWR_c_444_n
+ N_VPWR_c_445_n VPWR N_VPWR_c_446_n N_VPWR_c_447_n N_VPWR_c_448_n
+ N_VPWR_c_443_n N_VPWR_c_450_n N_VPWR_c_451_n PM_SKY130_FD_SC_LP__A2111O_0%VPWR
x_PM_SKY130_FD_SC_LP__A2111O_0%A_468_476# N_A_468_476#_M1003_d
+ N_A_468_476#_M1000_d N_A_468_476#_c_489_n N_A_468_476#_c_490_n
+ N_A_468_476#_c_491_n N_A_468_476#_c_492_n N_A_468_476#_c_493_n
+ PM_SKY130_FD_SC_LP__A2111O_0%A_468_476#
x_PM_SKY130_FD_SC_LP__A2111O_0%VGND N_VGND_M1008_d N_VGND_M1007_d N_VGND_M1011_d
+ N_VGND_c_523_n N_VGND_c_524_n N_VGND_c_525_n N_VGND_c_526_n N_VGND_c_527_n
+ VGND N_VGND_c_528_n N_VGND_c_529_n N_VGND_c_530_n N_VGND_c_531_n
+ PM_SKY130_FD_SC_LP__A2111O_0%VGND
cc_1 VNB N_A_80_159#_c_91_n 0.0222601f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.26
cc_2 VNB N_A_80_159#_M1005_g 0.0108375f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.735
cc_3 VNB N_A_80_159#_M1008_g 0.0216019f $X=-0.19 $Y=-0.245 $X2=0.735 $Y2=0.445
cc_4 VNB N_A_80_159#_c_94_n 0.0247989f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.465
cc_5 VNB N_A_80_159#_c_95_n 0.00129366f $X=-0.19 $Y=-0.245 $X2=0.672 $Y2=0.965
cc_6 VNB N_A_80_159#_c_96_n 0.00122097f $X=-0.19 $Y=-0.245 $X2=0.672 $Y2=2.055
cc_7 VNB N_A_80_159#_c_97_n 0.00935776f $X=-0.19 $Y=-0.245 $X2=1.245 $Y2=0.88
cc_8 VNB N_A_80_159#_c_98_n 0.00262864f $X=-0.19 $Y=-0.245 $X2=1.38 $Y2=0.445
cc_9 VNB N_A_80_159#_c_99_n 0.0259308f $X=-0.19 $Y=-0.245 $X2=2.49 $Y2=0.88
cc_10 VNB N_A_80_159#_c_100_n 0.00299574f $X=-0.19 $Y=-0.245 $X2=2.62 $Y2=0.445
cc_11 VNB N_A_80_159#_c_101_n 0.0238237f $X=-0.19 $Y=-0.245 $X2=0.645 $Y2=0.96
cc_12 VNB N_A_80_159#_c_102_n 0.00614282f $X=-0.19 $Y=-0.245 $X2=1.377 $Y2=0.88
cc_13 VNB N_D1_M1001_g 0.0385388f $X=-0.19 $Y=-0.245 $X2=1.145 $Y2=2.38
cc_14 VNB N_D1_c_178_n 0.0195796f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.465
cc_15 VNB D1 0.00607047f $X=-0.19 $Y=-0.245 $X2=0.735 $Y2=0.445
cc_16 VNB N_D1_c_180_n 0.0155663f $X=-0.19 $Y=-0.245 $X2=1.245 $Y2=0.88
cc_17 VNB N_C1_M1007_g 0.0238768f $X=-0.19 $Y=-0.245 $X2=1.145 $Y2=2.38
cc_18 VNB N_C1_c_232_n 0.0171481f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_C1_c_233_n 0.0163094f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB C1 0.00504539f $X=-0.19 $Y=-0.245 $X2=0.735 $Y2=0.445
cc_21 VNB N_C1_c_235_n 0.0167772f $X=-0.19 $Y=-0.245 $X2=1.27 $Y2=2.525
cc_22 VNB N_C1_c_236_n 0.0132687f $X=-0.19 $Y=-0.245 $X2=1.377 $Y2=0.795
cc_23 VNB N_B1_M1004_g 0.0447783f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_B1_c_287_n 0.0176172f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.26
cc_25 VNB B1 0.00582167f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.735
cc_26 VNB N_B1_c_289_n 0.0155431f $X=-0.19 $Y=-0.245 $X2=1.245 $Y2=0.88
cc_27 VNB N_A1_c_338_n 0.0246717f $X=-0.19 $Y=-0.245 $X2=1.24 $Y2=0.235
cc_28 VNB N_A1_c_339_n 0.0177361f $X=-0.19 $Y=-0.245 $X2=2.48 $Y2=0.235
cc_29 VNB N_A1_M1010_g 0.0384964f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_A1_c_341_n 0.00242546f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.26
cc_31 VNB A1 0.0115398f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.465
cc_32 VNB N_A2_c_389_n 0.0217754f $X=-0.19 $Y=-0.245 $X2=1.24 $Y2=0.235
cc_33 VNB N_A2_c_390_n 0.0089209f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A2_c_391_n 0.038391f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.735
cc_35 VNB N_A2_c_392_n 0.0185675f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.465
cc_36 VNB A2 0.0372835f $X=-0.19 $Y=-0.245 $X2=0.672 $Y2=0.965
cc_37 VNB N_A2_c_394_n 0.0355915f $X=-0.19 $Y=-0.245 $X2=1.24 $Y2=2.525
cc_38 VNB X 0.0564033f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_X_c_428_n 0.0210885f $X=-0.19 $Y=-0.245 $X2=1.377 $Y2=0.88
cc_40 VNB N_VPWR_c_443_n 0.163682f $X=-0.19 $Y=-0.245 $X2=1.38 $Y2=0.445
cc_41 VNB N_VGND_c_523_n 0.00462055f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.465
cc_42 VNB N_VGND_c_524_n 0.0159096f $X=-0.19 $Y=-0.245 $X2=0.735 $Y2=0.795
cc_43 VNB N_VGND_c_525_n 0.0180857f $X=-0.19 $Y=-0.245 $X2=0.735 $Y2=0.445
cc_44 VNB N_VGND_c_526_n 0.0230158f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=1.465
cc_45 VNB N_VGND_c_527_n 0.00497572f $X=-0.19 $Y=-0.245 $X2=0.672 $Y2=0.965
cc_46 VNB N_VGND_c_528_n 0.0251036f $X=-0.19 $Y=-0.245 $X2=1.24 $Y2=2.525
cc_47 VNB N_VGND_c_529_n 0.0168324f $X=-0.19 $Y=-0.245 $X2=1.51 $Y2=0.88
cc_48 VNB N_VGND_c_530_n 0.0190727f $X=-0.19 $Y=-0.245 $X2=0.645 $Y2=0.96
cc_49 VNB N_VGND_c_531_n 0.211479f $X=-0.19 $Y=-0.245 $X2=0.605 $Y2=0.96
cc_50 VPB N_A_80_159#_M1005_g 0.0614904f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.735
cc_51 VPB N_A_80_159#_c_96_n 0.00480924f $X=-0.19 $Y=1.655 $X2=0.672 $Y2=2.055
cc_52 VPB N_A_80_159#_c_105_n 0.0180746f $X=-0.19 $Y=1.655 $X2=1.105 $Y2=2.14
cc_53 VPB N_A_80_159#_c_106_n 0.00297831f $X=-0.19 $Y=1.655 $X2=0.81 $Y2=2.14
cc_54 VPB N_A_80_159#_c_107_n 0.0118159f $X=-0.19 $Y=1.655 $X2=1.27 $Y2=2.525
cc_55 VPB N_D1_c_181_n 0.0164111f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_56 VPB N_D1_c_182_n 0.0183464f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_57 VPB N_D1_c_178_n 0.00387641f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=1.465
cc_58 VPB N_D1_c_184_n 0.0169818f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.735
cc_59 VPB N_D1_c_185_n 0.0256757f $X=-0.19 $Y=1.655 $X2=0.735 $Y2=0.795
cc_60 VPB D1 0.00392514f $X=-0.19 $Y=1.655 $X2=0.735 $Y2=0.445
cc_61 VPB N_C1_c_232_n 0.00285802f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_62 VPB N_C1_M1009_g 0.0349895f $X=-0.19 $Y=1.655 $X2=0.605 $Y2=1.26
cc_63 VPB N_C1_c_239_n 0.0176853f $X=-0.19 $Y=1.655 $X2=0.735 $Y2=0.445
cc_64 VPB C1 0.00359142f $X=-0.19 $Y=1.655 $X2=0.735 $Y2=0.445
cc_65 VPB N_B1_M1003_g 0.0363665f $X=-0.19 $Y=1.655 $X2=1.145 $Y2=2.38
cc_66 VPB N_B1_c_287_n 0.00372549f $X=-0.19 $Y=1.655 $X2=0.605 $Y2=1.26
cc_67 VPB N_B1_c_292_n 0.0178816f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=1.465
cc_68 VPB B1 0.00482038f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.735
cc_69 VPB B1 0.00399581f $X=-0.19 $Y=1.655 $X2=0.735 $Y2=0.795
cc_70 VPB N_A1_M1006_g 0.0439891f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_71 VPB N_A1_c_341_n 0.0219175f $X=-0.19 $Y=1.655 $X2=0.605 $Y2=1.26
cc_72 VPB A1 0.00364517f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=1.465
cc_73 VPB N_A2_M1000_g 0.0223993f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_74 VPB N_A2_c_390_n 0.0307484f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_75 VPB N_A2_c_397_n 0.019395f $X=-0.19 $Y=1.655 $X2=0.735 $Y2=0.445
cc_76 VPB A2 0.0101494f $X=-0.19 $Y=1.655 $X2=0.672 $Y2=0.965
cc_77 VPB X 0.0680294f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_78 VPB N_VPWR_c_444_n 0.0135694f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_79 VPB N_VPWR_c_445_n 0.00970664f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.735
cc_80 VPB N_VPWR_c_446_n 0.0157693f $X=-0.19 $Y=1.655 $X2=0.735 $Y2=0.445
cc_81 VPB N_VPWR_c_447_n 0.0587056f $X=-0.19 $Y=1.655 $X2=0.672 $Y2=2.055
cc_82 VPB N_VPWR_c_448_n 0.018185f $X=-0.19 $Y=1.655 $X2=1.377 $Y2=0.445
cc_83 VPB N_VPWR_c_443_n 0.0767466f $X=-0.19 $Y=1.655 $X2=1.38 $Y2=0.445
cc_84 VPB N_VPWR_c_450_n 0.00526374f $X=-0.19 $Y=1.655 $X2=1.51 $Y2=0.88
cc_85 VPB N_VPWR_c_451_n 0.00507132f $X=-0.19 $Y=1.655 $X2=2.62 $Y2=0.445
cc_86 VPB N_A_468_476#_c_489_n 0.00345128f $X=-0.19 $Y=1.655 $X2=0.605 $Y2=1
cc_87 VPB N_A_468_476#_c_490_n 0.0190529f $X=-0.19 $Y=1.655 $X2=0.605 $Y2=1.26
cc_88 VPB N_A_468_476#_c_491_n 0.00863766f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=1.465
cc_89 VPB N_A_468_476#_c_492_n 0.0358666f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_90 VPB N_A_468_476#_c_493_n 0.00398857f $X=-0.19 $Y=1.655 $X2=0.605 $Y2=1.465
cc_91 N_A_80_159#_M1008_g N_D1_M1001_g 0.0332669f $X=0.735 $Y=0.445 $X2=0 $Y2=0
cc_92 N_A_80_159#_c_96_n N_D1_M1001_g 0.00113499f $X=0.672 $Y=2.055 $X2=0 $Y2=0
cc_93 N_A_80_159#_c_97_n N_D1_M1001_g 0.011812f $X=1.245 $Y=0.88 $X2=0 $Y2=0
cc_94 N_A_80_159#_c_98_n N_D1_M1001_g 0.00389978f $X=1.38 $Y=0.445 $X2=0 $Y2=0
cc_95 N_A_80_159#_M1005_g N_D1_c_181_n 0.00416986f $X=0.475 $Y=2.735 $X2=0 $Y2=0
cc_96 N_A_80_159#_c_96_n N_D1_c_181_n 0.0034737f $X=0.672 $Y=2.055 $X2=0 $Y2=0
cc_97 N_A_80_159#_c_105_n N_D1_c_181_n 0.00461789f $X=1.105 $Y=2.14 $X2=0 $Y2=0
cc_98 N_A_80_159#_c_107_n N_D1_c_182_n 0.00330239f $X=1.27 $Y=2.525 $X2=0 $Y2=0
cc_99 N_A_80_159#_M1005_g N_D1_c_178_n 0.00789186f $X=0.475 $Y=2.735 $X2=0 $Y2=0
cc_100 N_A_80_159#_c_94_n N_D1_c_178_n 0.00693201f $X=0.605 $Y=1.465 $X2=0 $Y2=0
cc_101 N_A_80_159#_c_96_n N_D1_c_178_n 0.0013724f $X=0.672 $Y=2.055 $X2=0 $Y2=0
cc_102 N_A_80_159#_c_105_n N_D1_c_184_n 0.00134656f $X=1.105 $Y=2.14 $X2=0 $Y2=0
cc_103 N_A_80_159#_c_105_n N_D1_c_185_n 0.00503575f $X=1.105 $Y=2.14 $X2=0 $Y2=0
cc_104 N_A_80_159#_c_107_n N_D1_c_185_n 0.00537398f $X=1.27 $Y=2.525 $X2=0 $Y2=0
cc_105 N_A_80_159#_c_91_n D1 0.00211977f $X=0.605 $Y=1.26 $X2=0 $Y2=0
cc_106 N_A_80_159#_M1005_g D1 9.61223e-19 $X=0.475 $Y=2.735 $X2=0 $Y2=0
cc_107 N_A_80_159#_c_96_n D1 0.0602584f $X=0.672 $Y=2.055 $X2=0 $Y2=0
cc_108 N_A_80_159#_c_97_n D1 0.0210165f $X=1.245 $Y=0.88 $X2=0 $Y2=0
cc_109 N_A_80_159#_c_105_n D1 0.0320758f $X=1.105 $Y=2.14 $X2=0 $Y2=0
cc_110 N_A_80_159#_c_102_n D1 0.0120921f $X=1.377 $Y=0.88 $X2=0 $Y2=0
cc_111 N_A_80_159#_c_91_n N_D1_c_180_n 0.00693201f $X=0.605 $Y=1.26 $X2=0 $Y2=0
cc_112 N_A_80_159#_c_96_n N_D1_c_180_n 2.87255e-19 $X=0.672 $Y=2.055 $X2=0 $Y2=0
cc_113 N_A_80_159#_c_97_n N_D1_c_180_n 2.57889e-19 $X=1.245 $Y=0.88 $X2=0 $Y2=0
cc_114 N_A_80_159#_c_102_n N_D1_c_180_n 0.00110462f $X=1.377 $Y=0.88 $X2=0 $Y2=0
cc_115 N_A_80_159#_c_98_n N_C1_M1007_g 0.00387458f $X=1.38 $Y=0.445 $X2=0 $Y2=0
cc_116 N_A_80_159#_c_99_n N_C1_M1007_g 0.00567779f $X=2.49 $Y=0.88 $X2=0 $Y2=0
cc_117 N_A_80_159#_c_99_n N_C1_c_233_n 0.011797f $X=2.49 $Y=0.88 $X2=0 $Y2=0
cc_118 N_A_80_159#_c_105_n C1 0.0137784f $X=1.105 $Y=2.14 $X2=0 $Y2=0
cc_119 N_A_80_159#_c_107_n C1 0.0327287f $X=1.27 $Y=2.525 $X2=0 $Y2=0
cc_120 N_A_80_159#_c_99_n C1 0.0257007f $X=2.49 $Y=0.88 $X2=0 $Y2=0
cc_121 N_A_80_159#_c_99_n N_C1_c_235_n 0.00362661f $X=2.49 $Y=0.88 $X2=0 $Y2=0
cc_122 N_A_80_159#_c_99_n N_B1_M1004_g 0.0148915f $X=2.49 $Y=0.88 $X2=0 $Y2=0
cc_123 N_A_80_159#_c_100_n N_B1_M1004_g 0.00384678f $X=2.62 $Y=0.445 $X2=0 $Y2=0
cc_124 N_A_80_159#_c_99_n B1 0.0304253f $X=2.49 $Y=0.88 $X2=0 $Y2=0
cc_125 N_A_80_159#_c_99_n N_B1_c_289_n 0.0013321f $X=2.49 $Y=0.88 $X2=0 $Y2=0
cc_126 N_A_80_159#_c_99_n N_A1_c_338_n 6.93845e-19 $X=2.49 $Y=0.88 $X2=-0.19
+ $Y2=-0.245
cc_127 N_A_80_159#_c_99_n N_A1_M1010_g 0.0014946f $X=2.49 $Y=0.88 $X2=0 $Y2=0
cc_128 N_A_80_159#_c_100_n N_A1_M1010_g 0.0035527f $X=2.62 $Y=0.445 $X2=0 $Y2=0
cc_129 N_A_80_159#_c_99_n A1 0.0150436f $X=2.49 $Y=0.88 $X2=0 $Y2=0
cc_130 N_A_80_159#_c_100_n A1 0.00118564f $X=2.62 $Y=0.445 $X2=0 $Y2=0
cc_131 N_A_80_159#_M1008_g X 0.00542503f $X=0.735 $Y=0.445 $X2=0 $Y2=0
cc_132 N_A_80_159#_c_95_n X 0.0140891f $X=0.672 $Y=0.965 $X2=0 $Y2=0
cc_133 N_A_80_159#_c_96_n X 0.0838258f $X=0.672 $Y=2.055 $X2=0 $Y2=0
cc_134 N_A_80_159#_c_106_n X 0.0140891f $X=0.81 $Y=2.14 $X2=0 $Y2=0
cc_135 N_A_80_159#_c_101_n X 0.0442221f $X=0.645 $Y=0.96 $X2=0 $Y2=0
cc_136 N_A_80_159#_c_95_n N_X_c_428_n 0.00658299f $X=0.672 $Y=0.965 $X2=0 $Y2=0
cc_137 N_A_80_159#_c_101_n N_X_c_428_n 0.0065749f $X=0.645 $Y=0.96 $X2=0 $Y2=0
cc_138 N_A_80_159#_M1005_g N_VPWR_c_444_n 0.0124402f $X=0.475 $Y=2.735 $X2=0
+ $Y2=0
cc_139 N_A_80_159#_c_105_n N_VPWR_c_444_n 0.00353232f $X=1.105 $Y=2.14 $X2=0
+ $Y2=0
cc_140 N_A_80_159#_c_106_n N_VPWR_c_444_n 0.0244741f $X=0.81 $Y=2.14 $X2=0 $Y2=0
cc_141 N_A_80_159#_c_107_n N_VPWR_c_444_n 0.0397188f $X=1.27 $Y=2.525 $X2=0
+ $Y2=0
cc_142 N_A_80_159#_M1005_g N_VPWR_c_446_n 0.00489337f $X=0.475 $Y=2.735 $X2=0
+ $Y2=0
cc_143 N_A_80_159#_c_107_n N_VPWR_c_447_n 0.0157217f $X=1.27 $Y=2.525 $X2=0
+ $Y2=0
cc_144 N_A_80_159#_M1005_g N_VPWR_c_443_n 0.00948861f $X=0.475 $Y=2.735 $X2=0
+ $Y2=0
cc_145 N_A_80_159#_c_107_n N_VPWR_c_443_n 0.0102395f $X=1.27 $Y=2.525 $X2=0
+ $Y2=0
cc_146 N_A_80_159#_M1008_g N_VGND_c_523_n 0.00319241f $X=0.735 $Y=0.445 $X2=0
+ $Y2=0
cc_147 N_A_80_159#_c_97_n N_VGND_c_523_n 0.0155344f $X=1.245 $Y=0.88 $X2=0 $Y2=0
cc_148 N_A_80_159#_M1008_g N_VGND_c_526_n 0.00585385f $X=0.735 $Y=0.445 $X2=0
+ $Y2=0
cc_149 N_A_80_159#_c_100_n N_VGND_c_528_n 0.0127495f $X=2.62 $Y=0.445 $X2=0
+ $Y2=0
cc_150 N_A_80_159#_c_98_n N_VGND_c_529_n 0.013059f $X=1.38 $Y=0.445 $X2=0 $Y2=0
cc_151 N_A_80_159#_c_99_n N_VGND_c_530_n 0.0440024f $X=2.49 $Y=0.88 $X2=0 $Y2=0
cc_152 N_A_80_159#_M1001_d N_VGND_c_531_n 0.00233419f $X=1.24 $Y=0.235 $X2=0
+ $Y2=0
cc_153 N_A_80_159#_M1004_d N_VGND_c_531_n 0.00286869f $X=2.48 $Y=0.235 $X2=0
+ $Y2=0
cc_154 N_A_80_159#_M1008_g N_VGND_c_531_n 0.00737685f $X=0.735 $Y=0.445 $X2=0
+ $Y2=0
cc_155 N_A_80_159#_c_95_n N_VGND_c_531_n 0.00573616f $X=0.672 $Y=0.965 $X2=0
+ $Y2=0
cc_156 N_A_80_159#_c_97_n N_VGND_c_531_n 0.00608283f $X=1.245 $Y=0.88 $X2=0
+ $Y2=0
cc_157 N_A_80_159#_c_98_n N_VGND_c_531_n 0.0101028f $X=1.38 $Y=0.445 $X2=0 $Y2=0
cc_158 N_A_80_159#_c_99_n N_VGND_c_531_n 0.0122597f $X=2.49 $Y=0.88 $X2=0 $Y2=0
cc_159 N_A_80_159#_c_100_n N_VGND_c_531_n 0.00971865f $X=2.62 $Y=0.445 $X2=0
+ $Y2=0
cc_160 N_D1_M1001_g N_C1_M1007_g 0.0218974f $X=1.165 $Y=0.445 $X2=0 $Y2=0
cc_161 N_D1_c_178_n N_C1_c_232_n 0.0139013f $X=1.215 $Y=1.71 $X2=0 $Y2=0
cc_162 N_D1_c_181_n N_C1_M1009_g 0.00542971f $X=1.305 $Y=2.12 $X2=0 $Y2=0
cc_163 N_D1_c_185_n N_C1_M1009_g 0.056652f $X=1.485 $Y=2.195 $X2=0 $Y2=0
cc_164 N_D1_c_184_n N_C1_c_239_n 0.0139013f $X=1.215 $Y=1.875 $X2=0 $Y2=0
cc_165 N_D1_c_182_n C1 0.0137207f $X=1.485 $Y=2.27 $X2=0 $Y2=0
cc_166 N_D1_c_185_n C1 0.00420305f $X=1.485 $Y=2.195 $X2=0 $Y2=0
cc_167 D1 C1 0.0594842f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_168 N_D1_c_180_n C1 0.00877015f $X=1.215 $Y=1.37 $X2=0 $Y2=0
cc_169 D1 N_C1_c_235_n 7.48023e-19 $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_170 N_D1_c_180_n N_C1_c_235_n 0.0139013f $X=1.215 $Y=1.37 $X2=0 $Y2=0
cc_171 N_D1_M1001_g N_C1_c_236_n 0.00714881f $X=1.165 $Y=0.445 $X2=0 $Y2=0
cc_172 D1 N_C1_c_236_n 2.27495e-19 $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_173 N_D1_c_180_n N_C1_c_236_n 2.16961e-19 $X=1.215 $Y=1.37 $X2=0 $Y2=0
cc_174 N_D1_c_182_n N_VPWR_c_444_n 0.00318696f $X=1.485 $Y=2.27 $X2=0 $Y2=0
cc_175 N_D1_c_182_n N_VPWR_c_447_n 0.00496106f $X=1.485 $Y=2.27 $X2=0 $Y2=0
cc_176 N_D1_c_182_n N_VPWR_c_443_n 0.0102513f $X=1.485 $Y=2.27 $X2=0 $Y2=0
cc_177 N_D1_M1001_g N_VGND_c_523_n 0.00168119f $X=1.165 $Y=0.445 $X2=0 $Y2=0
cc_178 N_D1_M1001_g N_VGND_c_529_n 0.00585385f $X=1.165 $Y=0.445 $X2=0 $Y2=0
cc_179 N_D1_M1001_g N_VGND_c_531_n 0.00624609f $X=1.165 $Y=0.445 $X2=0 $Y2=0
cc_180 N_C1_M1009_g N_B1_M1003_g 0.0638103f $X=1.875 $Y=2.7 $X2=0 $Y2=0
cc_181 C1 N_B1_M1003_g 0.00219395f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_182 N_C1_M1007_g N_B1_M1004_g 0.00647587f $X=1.595 $Y=0.445 $X2=0 $Y2=0
cc_183 N_C1_c_233_n N_B1_M1004_g 0.00792008f $X=1.71 $Y=0.92 $X2=0 $Y2=0
cc_184 N_C1_c_232_n N_B1_c_287_n 0.0138696f $X=1.77 $Y=1.7 $X2=0 $Y2=0
cc_185 N_C1_c_239_n N_B1_c_292_n 0.0138696f $X=1.77 $Y=1.88 $X2=0 $Y2=0
cc_186 C1 B1 0.0759353f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_187 N_C1_c_235_n B1 0.005861f $X=1.785 $Y=1.375 $X2=0 $Y2=0
cc_188 N_C1_c_236_n B1 2.60133e-19 $X=1.77 $Y=1.21 $X2=0 $Y2=0
cc_189 N_C1_M1009_g B1 0.00285315f $X=1.875 $Y=2.7 $X2=0 $Y2=0
cc_190 C1 B1 0.035278f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_191 C1 N_B1_c_289_n 5.83619e-19 $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_192 N_C1_c_235_n N_B1_c_289_n 0.0138696f $X=1.785 $Y=1.375 $X2=0 $Y2=0
cc_193 N_C1_M1009_g N_VPWR_c_447_n 0.00430047f $X=1.875 $Y=2.7 $X2=0 $Y2=0
cc_194 C1 N_VPWR_c_447_n 0.00992281f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_195 N_C1_M1009_g N_VPWR_c_443_n 0.00756384f $X=1.875 $Y=2.7 $X2=0 $Y2=0
cc_196 C1 N_VPWR_c_443_n 0.0112305f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_197 C1 A_312_476# 0.00160751f $X=1.595 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_198 N_C1_M1009_g N_A_468_476#_c_493_n 0.00112119f $X=1.875 $Y=2.7 $X2=0 $Y2=0
cc_199 C1 N_A_468_476#_c_493_n 0.0081562f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_200 N_C1_M1007_g N_VGND_c_529_n 0.00585385f $X=1.595 $Y=0.445 $X2=0 $Y2=0
cc_201 N_C1_M1007_g N_VGND_c_530_n 0.00243778f $X=1.595 $Y=0.445 $X2=0 $Y2=0
cc_202 N_C1_c_233_n N_VGND_c_530_n 5.78666e-19 $X=1.71 $Y=0.92 $X2=0 $Y2=0
cc_203 N_C1_M1007_g N_VGND_c_531_n 0.00694727f $X=1.595 $Y=0.445 $X2=0 $Y2=0
cc_204 N_B1_M1004_g N_A1_c_338_n 0.00221728f $X=2.405 $Y=0.445 $X2=-0.19
+ $Y2=-0.245
cc_205 B1 N_A1_c_338_n 0.00251555f $X=2.075 $Y=1.21 $X2=-0.19 $Y2=-0.245
cc_206 N_B1_c_289_n N_A1_c_338_n 0.0116999f $X=2.325 $Y=1.375 $X2=-0.19
+ $Y2=-0.245
cc_207 N_B1_c_287_n N_A1_c_339_n 0.0116999f $X=2.325 $Y=1.715 $X2=0 $Y2=0
cc_208 N_B1_M1004_g N_A1_M1010_g 0.0284396f $X=2.405 $Y=0.445 $X2=0 $Y2=0
cc_209 N_B1_M1003_g N_A1_M1006_g 0.0167171f $X=2.265 $Y=2.7 $X2=0 $Y2=0
cc_210 N_B1_c_292_n N_A1_M1006_g 0.00154898f $X=2.325 $Y=1.88 $X2=0 $Y2=0
cc_211 B1 N_A1_M1006_g 0.00305655f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_212 B1 N_A1_M1006_g 3.76911e-19 $X=2.075 $Y=2.32 $X2=0 $Y2=0
cc_213 N_B1_c_292_n N_A1_c_341_n 0.0116999f $X=2.325 $Y=1.88 $X2=0 $Y2=0
cc_214 B1 A1 0.0220309f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_215 N_B1_c_289_n A1 0.00180903f $X=2.325 $Y=1.375 $X2=0 $Y2=0
cc_216 N_B1_M1003_g N_VPWR_c_447_n 0.00480263f $X=2.265 $Y=2.7 $X2=0 $Y2=0
cc_217 N_B1_M1003_g N_VPWR_c_443_n 0.0077372f $X=2.265 $Y=2.7 $X2=0 $Y2=0
cc_218 B1 N_VPWR_c_443_n 0.00802014f $X=2.075 $Y=2.32 $X2=0 $Y2=0
cc_219 B1 A_390_476# 0.00342793f $X=2.075 $Y=2.32 $X2=-0.19 $Y2=-0.245
cc_220 N_B1_M1003_g N_A_468_476#_c_489_n 0.00621384f $X=2.265 $Y=2.7 $X2=0 $Y2=0
cc_221 B1 N_A_468_476#_c_489_n 0.0184965f $X=2.075 $Y=2.32 $X2=0 $Y2=0
cc_222 N_B1_M1003_g N_A_468_476#_c_491_n 6.63008e-19 $X=2.265 $Y=2.7 $X2=0 $Y2=0
cc_223 B1 N_A_468_476#_c_491_n 0.005754f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_224 B1 N_A_468_476#_c_491_n 0.00940668f $X=2.075 $Y=2.32 $X2=0 $Y2=0
cc_225 N_B1_M1003_g N_A_468_476#_c_493_n 0.00655094f $X=2.265 $Y=2.7 $X2=0 $Y2=0
cc_226 B1 N_A_468_476#_c_493_n 0.00285197f $X=2.075 $Y=2.32 $X2=0 $Y2=0
cc_227 N_B1_M1004_g N_VGND_c_528_n 0.00585385f $X=2.405 $Y=0.445 $X2=0 $Y2=0
cc_228 N_B1_M1004_g N_VGND_c_530_n 0.0040695f $X=2.405 $Y=0.445 $X2=0 $Y2=0
cc_229 N_B1_M1004_g N_VGND_c_531_n 0.00694727f $X=2.405 $Y=0.445 $X2=0 $Y2=0
cc_230 N_A1_M1010_g N_A2_c_389_n 0.0497825f $X=2.835 $Y=0.445 $X2=-0.19
+ $Y2=-0.245
cc_231 N_A1_M1006_g N_A2_c_390_n 0.00782772f $X=2.91 $Y=2.7 $X2=0 $Y2=0
cc_232 N_A1_c_341_n N_A2_c_390_n 0.0114116f $X=2.947 $Y=1.84 $X2=0 $Y2=0
cc_233 N_A1_c_338_n N_A2_c_391_n 0.00249419f $X=2.947 $Y=1.387 $X2=0 $Y2=0
cc_234 A1 N_A2_c_391_n 0.0104998f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_235 N_A1_M1006_g N_A2_c_397_n 0.0183286f $X=2.91 $Y=2.7 $X2=0 $Y2=0
cc_236 N_A1_c_339_n N_A2_c_392_n 0.0114116f $X=2.947 $Y=1.623 $X2=0 $Y2=0
cc_237 N_A1_c_338_n A2 6.98976e-19 $X=2.947 $Y=1.387 $X2=0 $Y2=0
cc_238 A1 A2 0.0833501f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_239 N_A1_c_338_n N_A2_c_394_n 0.0114116f $X=2.947 $Y=1.387 $X2=0 $Y2=0
cc_240 N_A1_M1010_g N_A2_c_394_n 0.00377314f $X=2.835 $Y=0.445 $X2=0 $Y2=0
cc_241 A1 N_A2_c_394_n 0.00620828f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_242 N_A1_M1006_g N_VPWR_c_445_n 0.00302461f $X=2.91 $Y=2.7 $X2=0 $Y2=0
cc_243 N_A1_M1006_g N_VPWR_c_447_n 0.00512921f $X=2.91 $Y=2.7 $X2=0 $Y2=0
cc_244 N_A1_M1006_g N_VPWR_c_443_n 0.0101328f $X=2.91 $Y=2.7 $X2=0 $Y2=0
cc_245 N_A1_M1006_g N_A_468_476#_c_489_n 0.00314229f $X=2.91 $Y=2.7 $X2=0 $Y2=0
cc_246 N_A1_M1006_g N_A_468_476#_c_490_n 0.0180639f $X=2.91 $Y=2.7 $X2=0 $Y2=0
cc_247 N_A1_c_341_n N_A_468_476#_c_490_n 0.00183707f $X=2.947 $Y=1.84 $X2=0
+ $Y2=0
cc_248 A1 N_A_468_476#_c_490_n 0.0256048f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_249 N_A1_c_341_n N_A_468_476#_c_491_n 0.00427685f $X=2.947 $Y=1.84 $X2=0
+ $Y2=0
cc_250 N_A1_M1006_g N_A_468_476#_c_493_n 0.00242446f $X=2.91 $Y=2.7 $X2=0 $Y2=0
cc_251 N_A1_M1010_g N_VGND_c_525_n 0.00241774f $X=2.835 $Y=0.445 $X2=0 $Y2=0
cc_252 A1 N_VGND_c_525_n 0.00271362f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_253 N_A1_M1010_g N_VGND_c_528_n 0.00585385f $X=2.835 $Y=0.445 $X2=0 $Y2=0
cc_254 N_A1_M1010_g N_VGND_c_531_n 0.0108402f $X=2.835 $Y=0.445 $X2=0 $Y2=0
cc_255 A1 N_VGND_c_531_n 0.0118449f $X=3.035 $Y=0.84 $X2=0 $Y2=0
cc_256 N_A2_M1000_g N_VPWR_c_445_n 0.00298017f $X=3.34 $Y=2.7 $X2=0 $Y2=0
cc_257 N_A2_M1000_g N_VPWR_c_448_n 0.00512921f $X=3.34 $Y=2.7 $X2=0 $Y2=0
cc_258 N_A2_M1000_g N_VPWR_c_443_n 0.0103953f $X=3.34 $Y=2.7 $X2=0 $Y2=0
cc_259 N_A2_c_390_n N_A_468_476#_c_490_n 0.00540061f $X=3.48 $Y=2.08 $X2=0 $Y2=0
cc_260 N_A2_c_397_n N_A_468_476#_c_490_n 0.015311f $X=3.48 $Y=2.155 $X2=0 $Y2=0
cc_261 N_A2_c_392_n N_A_468_476#_c_490_n 6.37586e-19 $X=3.57 $Y=1.51 $X2=0 $Y2=0
cc_262 A2 N_A_468_476#_c_490_n 0.0258916f $X=3.515 $Y=0.84 $X2=0 $Y2=0
cc_263 N_A2_M1000_g N_A_468_476#_c_492_n 0.00491829f $X=3.34 $Y=2.7 $X2=0 $Y2=0
cc_264 N_A2_c_397_n N_A_468_476#_c_492_n 0.00508223f $X=3.48 $Y=2.155 $X2=0
+ $Y2=0
cc_265 N_A2_c_391_n N_VGND_c_524_n 9.88622e-19 $X=3.57 $Y=0.93 $X2=0 $Y2=0
cc_266 N_A2_c_389_n N_VGND_c_525_n 0.0153833f $X=3.195 $Y=0.78 $X2=0 $Y2=0
cc_267 N_A2_c_391_n N_VGND_c_525_n 0.00627521f $X=3.57 $Y=0.93 $X2=0 $Y2=0
cc_268 A2 N_VGND_c_525_n 0.014807f $X=3.515 $Y=0.84 $X2=0 $Y2=0
cc_269 N_A2_c_389_n N_VGND_c_528_n 0.00368966f $X=3.195 $Y=0.78 $X2=0 $Y2=0
cc_270 N_A2_c_389_n N_VGND_c_531_n 0.00340079f $X=3.195 $Y=0.78 $X2=0 $Y2=0
cc_271 A2 N_VGND_c_531_n 0.00672002f $X=3.515 $Y=0.84 $X2=0 $Y2=0
cc_272 X N_VPWR_c_444_n 0.0261581f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_273 X N_VPWR_c_446_n 0.0199289f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_274 X N_VPWR_c_443_n 0.010808f $X=0.155 $Y=0.47 $X2=0 $Y2=0
cc_275 N_X_c_428_n N_VGND_c_526_n 0.0312811f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_276 N_X_M1008_s N_VGND_c_531_n 0.0022581f $X=0.395 $Y=0.235 $X2=0 $Y2=0
cc_277 N_X_c_428_n N_VGND_c_531_n 0.0210745f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_278 N_VPWR_c_445_n N_A_468_476#_c_489_n 7.19015e-19 $X=3.125 $Y=2.535 $X2=0
+ $Y2=0
cc_279 N_VPWR_c_445_n N_A_468_476#_c_490_n 0.0213306f $X=3.125 $Y=2.535 $X2=0
+ $Y2=0
cc_280 N_VPWR_c_445_n N_A_468_476#_c_492_n 0.00227218f $X=3.125 $Y=2.535 $X2=0
+ $Y2=0
cc_281 N_VPWR_c_448_n N_A_468_476#_c_492_n 0.0171883f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_282 N_VPWR_c_443_n N_A_468_476#_c_492_n 0.0111947f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_283 N_VPWR_c_445_n N_A_468_476#_c_493_n 0.00152987f $X=3.125 $Y=2.535 $X2=0
+ $Y2=0
cc_284 N_VPWR_c_447_n N_A_468_476#_c_493_n 0.027874f $X=2.99 $Y=3.33 $X2=0 $Y2=0
cc_285 N_VPWR_c_443_n N_A_468_476#_c_493_n 0.0187782f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_286 N_VGND_c_531_n A_582_47# 0.00307285f $X=3.6 $Y=0 $X2=-0.19 $Y2=-0.245
