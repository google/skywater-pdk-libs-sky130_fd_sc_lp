* File: sky130_fd_sc_lp__nor3b_2.pex.spice
* Created: Fri Aug 28 10:56:25 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__NOR3B_2%C_N 3 7 11 12 13 14 18 19
c33 19 0 6.87565e-20 $X=0.385 $Y=1.615
r34 18 19 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.385
+ $Y=1.615 $X2=0.385 $Y2=1.615
r35 13 14 11.0754 $w=3.83e-07 $l=3.7e-07 $layer=LI1_cond $X=0.277 $Y=1.665
+ $X2=0.277 $Y2=2.035
r36 13 19 1.49668 $w=3.83e-07 $l=5e-08 $layer=LI1_cond $X=0.277 $Y=1.665
+ $X2=0.277 $Y2=1.615
r37 11 18 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=0.385 $Y=1.955
+ $X2=0.385 $Y2=1.615
r38 11 12 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.385 $Y=1.955
+ $X2=0.385 $Y2=2.12
r39 10 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.385 $Y=1.45
+ $X2=0.385 $Y2=1.615
r40 7 12 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=0.475 $Y=2.75
+ $X2=0.475 $Y2=2.12
r41 3 10 299.968 $w=1.5e-07 $l=5.85e-07 $layer=POLY_cond $X=0.475 $Y=0.865
+ $X2=0.475 $Y2=1.45
.ends

.subckt PM_SKY130_FD_SC_LP__NOR3B_2%A_27_131# 1 2 9 11 13 16 18 20 21 24 28 32
+ 34 35 36 37 39 42 45
c87 21 0 6.87565e-20 $X=1.35 $Y=1.35
r88 42 43 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.34
+ $Y=1.35 $X2=1.34 $Y2=1.35
r89 40 45 3.70735 $w=2.5e-07 $l=1.0225e-07 $layer=LI1_cond $X=0.925 $Y=1.35
+ $X2=0.84 $Y2=1.312
r90 40 42 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=0.925 $Y=1.35
+ $X2=1.34 $Y2=1.35
r91 38 45 2.76166 $w=1.7e-07 $l=2.03e-07 $layer=LI1_cond $X=0.84 $Y=1.515
+ $X2=0.84 $Y2=1.312
r92 38 39 51.2139 $w=1.68e-07 $l=7.85e-07 $layer=LI1_cond $X=0.84 $Y=1.515
+ $X2=0.84 $Y2=2.3
r93 36 39 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.755 $Y=2.385
+ $X2=0.84 $Y2=2.3
r94 36 37 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=0.755 $Y=2.385
+ $X2=0.355 $Y2=2.385
r95 34 45 3.70735 $w=2.5e-07 $l=1.53734e-07 $layer=LI1_cond $X=0.755 $Y=1.195
+ $X2=0.84 $Y2=1.312
r96 34 35 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=0.755 $Y=1.195
+ $X2=0.355 $Y2=1.195
r97 30 37 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=0.225 $Y=2.47
+ $X2=0.355 $Y2=2.385
r98 30 32 12.4109 $w=2.58e-07 $l=2.8e-07 $layer=LI1_cond $X=0.225 $Y=2.47
+ $X2=0.225 $Y2=2.75
r99 26 35 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=0.225 $Y=1.11
+ $X2=0.355 $Y2=1.195
r100 26 28 10.8596 $w=2.58e-07 $l=2.45e-07 $layer=LI1_cond $X=0.225 $Y=1.11
+ $X2=0.225 $Y2=0.865
r101 23 24 61.4966 $w=2.9e-07 $l=3.7e-07 $layer=POLY_cond $X=1.485 $Y=1.35
+ $X2=1.855 $Y2=1.35
r102 22 23 9.97241 $w=2.9e-07 $l=6e-08 $layer=POLY_cond $X=1.425 $Y=1.35
+ $X2=1.485 $Y2=1.35
r103 21 43 1.74861 $w=3.3e-07 $l=1e-08 $layer=POLY_cond $X=1.35 $Y=1.35 $X2=1.34
+ $Y2=1.35
r104 21 22 11.7856 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=1.35 $Y=1.35
+ $X2=1.425 $Y2=1.35
r105 18 24 27.4241 $w=2.9e-07 $l=2.33345e-07 $layer=POLY_cond $X=2.02 $Y=1.185
+ $X2=1.855 $Y2=1.35
r106 18 20 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.02 $Y=1.185
+ $X2=2.02 $Y2=0.655
r107 14 24 18.1727 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.855 $Y=1.515
+ $X2=1.855 $Y2=1.35
r108 14 16 482 $w=1.5e-07 $l=9.4e-07 $layer=POLY_cond $X=1.855 $Y=1.515
+ $X2=1.855 $Y2=2.455
r109 11 23 18.1727 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.485 $Y=1.185
+ $X2=1.485 $Y2=1.35
r110 11 13 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.485 $Y=1.185
+ $X2=1.485 $Y2=0.655
r111 7 22 18.1727 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.425 $Y=1.515
+ $X2=1.425 $Y2=1.35
r112 7 9 482 $w=1.5e-07 $l=9.4e-07 $layer=POLY_cond $X=1.425 $Y=1.515 $X2=1.425
+ $Y2=2.455
r113 2 32 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.54 $X2=0.26 $Y2=2.75
r114 1 28 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.655 $X2=0.26 $Y2=0.865
.ends

.subckt PM_SKY130_FD_SC_LP__NOR3B_2%B 3 7 11 15 19 25 26
c56 11 0 1.40652e-19 $X=2.715 $Y=2.455
r57 25 27 4.24296 $w=2.84e-07 $l=2.5e-08 $layer=POLY_cond $X=2.945 $Y=1.5
+ $X2=2.97 $Y2=1.5
r58 25 26 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.945
+ $Y=1.5 $X2=2.945 $Y2=1.5
r59 23 25 39.0352 $w=2.84e-07 $l=2.3e-07 $layer=POLY_cond $X=2.715 $Y=1.5
+ $X2=2.945 $Y2=1.5
r60 22 23 29.7007 $w=2.84e-07 $l=1.75e-07 $layer=POLY_cond $X=2.54 $Y=1.5
+ $X2=2.715 $Y2=1.5
r61 19 26 4.8597 $w=4.13e-07 $l=1.75e-07 $layer=LI1_cond $X=3.12 $Y=1.542
+ $X2=2.945 $Y2=1.542
r62 13 27 17.6835 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.97 $Y=1.335
+ $X2=2.97 $Y2=1.5
r63 13 15 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=2.97 $Y=1.335
+ $X2=2.97 $Y2=0.655
r64 9 23 17.6835 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.715 $Y=1.665
+ $X2=2.715 $Y2=1.5
r65 9 11 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.715 $Y=1.665
+ $X2=2.715 $Y2=2.455
r66 5 22 17.6835 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.54 $Y=1.335
+ $X2=2.54 $Y2=1.5
r67 5 7 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=2.54 $Y=1.335 $X2=2.54
+ $Y2=0.655
r68 1 22 43.2782 $w=2.84e-07 $l=3.27261e-07 $layer=POLY_cond $X=2.285 $Y=1.665
+ $X2=2.54 $Y2=1.5
r69 1 3 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=2.285 $Y=1.665
+ $X2=2.285 $Y2=2.455
.ends

.subckt PM_SKY130_FD_SC_LP__NOR3B_2%A 3 7 11 15 17 18 19 33
c41 33 0 1.40652e-19 $X=4.32 $Y=1.51
r42 31 33 15.7375 $w=3.3e-07 $l=9e-08 $layer=POLY_cond $X=4.23 $Y=1.51 $X2=4.32
+ $Y2=1.51
r43 31 32 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=4.23
+ $Y=1.51 $X2=4.23 $Y2=1.51
r44 29 31 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=3.89 $Y=1.51
+ $X2=4.23 $Y2=1.51
r45 28 29 10.4917 $w=3.3e-07 $l=6e-08 $layer=POLY_cond $X=3.83 $Y=1.51 $X2=3.89
+ $Y2=1.51
r46 26 28 48.9612 $w=3.3e-07 $l=2.8e-07 $layer=POLY_cond $X=3.55 $Y=1.51
+ $X2=3.83 $Y2=1.51
r47 26 27 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=3.55
+ $Y=1.51 $X2=3.55 $Y2=1.51
r48 23 26 26.2292 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=3.4 $Y=1.51 $X2=3.55
+ $Y2=1.51
r49 19 32 9.164 $w=4.13e-07 $l=3.3e-07 $layer=LI1_cond $X=4.56 $Y=1.542 $X2=4.23
+ $Y2=1.542
r50 18 32 4.16546 $w=4.13e-07 $l=1.5e-07 $layer=LI1_cond $X=4.08 $Y=1.542
+ $X2=4.23 $Y2=1.542
r51 17 18 13.3295 $w=4.13e-07 $l=4.8e-07 $layer=LI1_cond $X=3.6 $Y=1.542
+ $X2=4.08 $Y2=1.542
r52 17 27 1.38849 $w=4.13e-07 $l=5e-08 $layer=LI1_cond $X=3.6 $Y=1.542 $X2=3.55
+ $Y2=1.542
r53 13 33 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.32 $Y=1.675
+ $X2=4.32 $Y2=1.51
r54 13 15 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=4.32 $Y=1.675
+ $X2=4.32 $Y2=2.465
r55 9 29 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.89 $Y=1.675
+ $X2=3.89 $Y2=1.51
r56 9 11 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=3.89 $Y=1.675
+ $X2=3.89 $Y2=2.465
r57 5 28 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.83 $Y=1.345
+ $X2=3.83 $Y2=1.51
r58 5 7 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.83 $Y=1.345 $X2=3.83
+ $Y2=0.655
r59 1 23 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.4 $Y=1.345 $X2=3.4
+ $Y2=1.51
r60 1 3 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=3.4 $Y=1.345 $X2=3.4
+ $Y2=0.655
.ends

.subckt PM_SKY130_FD_SC_LP__NOR3B_2%VPWR 1 2 3 12 16 18 20 24 26 31 39 45 48 52
r58 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r59 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r60 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r61 43 52 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=4.56 $Y2=3.33
r62 43 49 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.08 $Y=3.33
+ $X2=3.6 $Y2=3.33
r63 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r64 40 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.84 $Y=3.33
+ $X2=3.675 $Y2=3.33
r65 40 42 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=3.84 $Y=3.33
+ $X2=4.08 $Y2=3.33
r66 39 51 4.77065 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=4.37 $Y=3.33
+ $X2=4.585 $Y2=3.33
r67 39 42 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=4.37 $Y=3.33
+ $X2=4.08 $Y2=3.33
r68 38 49 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=3.33
+ $X2=3.6 $Y2=3.33
r69 37 38 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r70 35 46 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=3.33
+ $X2=0.72 $Y2=3.33
r71 34 37 125.262 $w=1.68e-07 $l=1.92e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=3.12 $Y2=3.33
r72 34 35 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33
+ $X2=1.2 $Y2=3.33
r73 32 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.855 $Y=3.33
+ $X2=0.69 $Y2=3.33
r74 32 34 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.855 $Y=3.33
+ $X2=1.2 $Y2=3.33
r75 31 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.51 $Y=3.33
+ $X2=3.675 $Y2=3.33
r76 31 37 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=3.51 $Y=3.33
+ $X2=3.12 $Y2=3.33
r77 29 46 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r78 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r79 26 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.525 $Y=3.33
+ $X2=0.69 $Y2=3.33
r80 26 28 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.525 $Y=3.33
+ $X2=0.24 $Y2=3.33
r81 24 38 0.200689 $w=4.9e-07 $l=7.2e-07 $layer=MET1_cond $X=2.4 $Y=3.33
+ $X2=3.12 $Y2=3.33
r82 24 35 0.334482 $w=4.9e-07 $l=1.2e-06 $layer=MET1_cond $X=2.4 $Y=3.33 $X2=1.2
+ $Y2=3.33
r83 20 23 33.0018 $w=3.28e-07 $l=9.45e-07 $layer=LI1_cond $X=4.535 $Y=2.005
+ $X2=4.535 $Y2=2.95
r84 18 51 2.99552 $w=3.3e-07 $l=1.07121e-07 $layer=LI1_cond $X=4.535 $Y=3.245
+ $X2=4.585 $Y2=3.33
r85 18 23 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=4.535 $Y=3.245
+ $X2=4.535 $Y2=2.95
r86 14 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.675 $Y=3.245
+ $X2=3.675 $Y2=3.33
r87 14 16 30.7318 $w=3.28e-07 $l=8.8e-07 $layer=LI1_cond $X=3.675 $Y=3.245
+ $X2=3.675 $Y2=2.365
r88 10 45 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=3.245
+ $X2=0.69 $Y2=3.33
r89 10 12 16.7628 $w=3.28e-07 $l=4.8e-07 $layer=LI1_cond $X=0.69 $Y=3.245
+ $X2=0.69 $Y2=2.765
r90 3 23 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=4.395
+ $Y=1.835 $X2=4.535 $Y2=2.95
r91 3 20 400 $w=1.7e-07 $l=2.29565e-07 $layer=licon1_PDIFF $count=1 $X=4.395
+ $Y=1.835 $X2=4.535 $Y2=2.005
r92 2 16 300 $w=1.7e-07 $l=5.89194e-07 $layer=licon1_PDIFF $count=2 $X=3.55
+ $Y=1.835 $X2=3.675 $Y2=2.365
r93 1 12 600 $w=1.7e-07 $l=2.86575e-07 $layer=licon1_PDIFF $count=1 $X=0.55
+ $Y=2.54 $X2=0.69 $Y2=2.765
.ends

.subckt PM_SKY130_FD_SC_LP__NOR3B_2%A_217_365# 1 2 3 10 12 14 18 20 24 29
r42 22 24 21.2759 $w=2.58e-07 $l=4.8e-07 $layer=LI1_cond $X=2.965 $Y=2.905
+ $X2=2.965 $Y2=2.425
r43 21 29 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.165 $Y=2.99
+ $X2=2.07 $Y2=2.99
r44 20 22 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=2.835 $Y=2.99
+ $X2=2.965 $Y2=2.905
r45 20 21 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.835 $Y=2.99
+ $X2=2.165 $Y2=2.99
r46 16 29 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=2.07 $Y=2.905
+ $X2=2.07 $Y2=2.99
r47 16 18 54.5789 $w=1.88e-07 $l=9.35e-07 $layer=LI1_cond $X=2.07 $Y=2.905
+ $X2=2.07 $Y2=1.97
r48 15 27 3.82155 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.305 $Y=2.99
+ $X2=1.2 $Y2=2.99
r49 14 29 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.975 $Y=2.99
+ $X2=2.07 $Y2=2.99
r50 14 15 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.975 $Y=2.99
+ $X2=1.305 $Y2=2.99
r51 10 27 3.09364 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=1.2 $Y=2.905 $X2=1.2
+ $Y2=2.99
r52 10 12 49.381 $w=2.08e-07 $l=9.35e-07 $layer=LI1_cond $X=1.2 $Y=2.905 $X2=1.2
+ $Y2=1.97
r53 3 24 300 $w=1.7e-07 $l=6.66333e-07 $layer=licon1_PDIFF $count=2 $X=2.79
+ $Y=1.825 $X2=2.93 $Y2=2.425
r54 2 29 400 $w=1.7e-07 $l=1.15288e-06 $layer=licon1_PDIFF $count=1 $X=1.93
+ $Y=1.825 $X2=2.07 $Y2=2.91
r55 2 18 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.93
+ $Y=1.825 $X2=2.07 $Y2=1.97
r56 1 27 400 $w=1.7e-07 $l=1.1458e-06 $layer=licon1_PDIFF $count=1 $X=1.085
+ $Y=1.825 $X2=1.21 $Y2=2.91
r57 1 12 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=1.085
+ $Y=1.825 $X2=1.21 $Y2=1.97
.ends

.subckt PM_SKY130_FD_SC_LP__NOR3B_2%Y 1 2 3 4 13 17 19 23 25 26 27 28 29 30 31
+ 42 48 57
r59 55 57 0.873063 $w=3.28e-07 $l=2.5e-08 $layer=LI1_cond $X=1.64 $Y=2.01
+ $X2=1.64 $Y2=2.035
r60 40 48 2.09535 $w=3.28e-07 $l=6e-08 $layer=LI1_cond $X=1.76 $Y=0.985 $X2=1.76
+ $Y2=0.925
r61 31 62 8.55602 $w=3.28e-07 $l=2.45e-07 $layer=LI1_cond $X=1.64 $Y=2.405
+ $X2=1.64 $Y2=2.65
r62 30 55 2.09535 $w=3.28e-07 $l=6e-08 $layer=LI1_cond $X=1.64 $Y=1.95 $X2=1.64
+ $Y2=2.01
r63 30 67 5.18491 $w=3.28e-07 $l=1.05e-07 $layer=LI1_cond $X=1.64 $Y=1.95
+ $X2=1.64 $Y2=1.845
r64 30 31 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=1.64 $Y=2.065
+ $X2=1.64 $Y2=2.405
r65 30 57 1.04768 $w=3.28e-07 $l=3e-08 $layer=LI1_cond $X=1.64 $Y=2.065 $X2=1.64
+ $Y2=2.035
r66 29 67 9.50649 $w=2.08e-07 $l=1.8e-07 $layer=LI1_cond $X=1.7 $Y=1.665 $X2=1.7
+ $Y2=1.845
r67 28 29 19.5411 $w=2.08e-07 $l=3.7e-07 $layer=LI1_cond $X=1.7 $Y=1.295 $X2=1.7
+ $Y2=1.665
r68 28 49 6.8658 $w=2.08e-07 $l=1.3e-07 $layer=LI1_cond $X=1.7 $Y=1.295 $X2=1.7
+ $Y2=1.165
r69 27 40 3.64284 $w=2.7e-07 $l=9e-08 $layer=LI1_cond $X=1.76 $Y=1.075 $X2=1.76
+ $Y2=0.985
r70 27 49 3.64284 $w=2.7e-07 $l=1.16189e-07 $layer=LI1_cond $X=1.76 $Y=1.075
+ $X2=1.7 $Y2=1.165
r71 27 48 0.453993 $w=3.28e-07 $l=1.3e-08 $layer=LI1_cond $X=1.76 $Y=0.912
+ $X2=1.76 $Y2=0.925
r72 26 27 12.4673 $w=3.28e-07 $l=3.57e-07 $layer=LI1_cond $X=1.76 $Y=0.555
+ $X2=1.76 $Y2=0.912
r73 26 42 4.71454 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=1.76 $Y=0.555
+ $X2=1.76 $Y2=0.42
r74 21 23 28.8111 $w=2.28e-07 $l=5.75e-07 $layer=LI1_cond $X=3.635 $Y=0.995
+ $X2=3.635 $Y2=0.42
r75 20 25 6.44382 $w=1.75e-07 $l=1.17473e-07 $layer=LI1_cond $X=2.85 $Y=1.08
+ $X2=2.735 $Y2=1.075
r76 19 21 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=3.52 $Y=1.08
+ $X2=3.635 $Y2=0.995
r77 19 20 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.52 $Y=1.08
+ $X2=2.85 $Y2=1.08
r78 15 25 0.379591 $w=2.3e-07 $l=9e-08 $layer=LI1_cond $X=2.735 $Y=0.985
+ $X2=2.735 $Y2=1.075
r79 15 17 28.31 $w=2.28e-07 $l=5.65e-07 $layer=LI1_cond $X=2.735 $Y=0.985
+ $X2=2.735 $Y2=0.42
r80 14 27 2.83584 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=1.925 $Y=1.075
+ $X2=1.76 $Y2=1.075
r81 13 25 6.44382 $w=1.75e-07 $l=1.15e-07 $layer=LI1_cond $X=2.62 $Y=1.075
+ $X2=2.735 $Y2=1.075
r82 13 14 42.8232 $w=1.78e-07 $l=6.95e-07 $layer=LI1_cond $X=2.62 $Y=1.075
+ $X2=1.925 $Y2=1.075
r83 4 30 400 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=1.5
+ $Y=1.825 $X2=1.64 $Y2=1.95
r84 4 62 400 $w=1.7e-07 $l=8.92258e-07 $layer=licon1_PDIFF $count=1 $X=1.5
+ $Y=1.825 $X2=1.64 $Y2=2.65
r85 3 23 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=3.475
+ $Y=0.235 $X2=3.615 $Y2=0.42
r86 2 17 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=2.615
+ $Y=0.235 $X2=2.755 $Y2=0.42
r87 1 42 91 $w=1.7e-07 $l=2.77489e-07 $layer=licon1_NDIFF $count=2 $X=1.56
+ $Y=0.235 $X2=1.76 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_LP__NOR3B_2%A_472_365# 1 2 7 9 11 13 15
r26 13 20 3.31438 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=4.1 $Y=2.09 $X2=4.1
+ $Y2=2.005
r27 13 15 50.5253 $w=1.78e-07 $l=8.2e-07 $layer=LI1_cond $X=4.1 $Y=2.09 $X2=4.1
+ $Y2=2.91
r28 12 18 4.83599 $w=1.7e-07 $l=1.83016e-07 $layer=LI1_cond $X=2.665 $Y=2.005
+ $X2=2.5 $Y2=1.967
r29 11 20 3.50935 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=4.01 $Y=2.005 $X2=4.1
+ $Y2=2.005
r30 11 12 87.7487 $w=1.68e-07 $l=1.345e-06 $layer=LI1_cond $X=4.01 $Y=2.005
+ $X2=2.665 $Y2=2.005
r31 7 18 2.93018 $w=3.3e-07 $l=1.23e-07 $layer=LI1_cond $X=2.5 $Y=2.09 $X2=2.5
+ $Y2=1.967
r32 7 9 19.5566 $w=3.28e-07 $l=5.6e-07 $layer=LI1_cond $X=2.5 $Y=2.09 $X2=2.5
+ $Y2=2.65
r33 2 20 400 $w=1.7e-07 $l=3.1225e-07 $layer=licon1_PDIFF $count=1 $X=3.965
+ $Y=1.835 $X2=4.105 $Y2=2.085
r34 2 15 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=3.965
+ $Y=1.835 $X2=4.105 $Y2=2.91
r35 1 18 400 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_PDIFF $count=1 $X=2.36
+ $Y=1.825 $X2=2.5 $Y2=1.95
r36 1 9 400 $w=1.7e-07 $l=8.92258e-07 $layer=licon1_PDIFF $count=1 $X=2.36
+ $Y=1.825 $X2=2.5 $Y2=2.65
.ends

.subckt PM_SKY130_FD_SC_LP__NOR3B_2%VGND 1 2 3 4 13 17 21 25 27 29 34 39 46 47
+ 51 63 66 69
r59 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r60 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r61 63 64 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r62 58 60 0.813333 $w=8.98e-07 $l=6e-08 $layer=LI1_cond $X=0.975 $Y=0.775
+ $X2=0.975 $Y2=0.835
r63 56 58 5.35444 $w=8.98e-07 $l=3.95e-07 $layer=LI1_cond $X=0.975 $Y=0.38
+ $X2=0.975 $Y2=0.775
r64 54 64 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r65 52 54 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r66 51 56 5.15111 $w=8.98e-07 $l=3.8e-07 $layer=LI1_cond $X=0.975 $Y=0 $X2=0.975
+ $Y2=0.38
r67 51 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r68 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r69 47 70 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=4.08
+ $Y2=0
r70 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r71 44 69 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=4.21 $Y=0 $X2=4.065
+ $Y2=0
r72 44 46 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=4.21 $Y=0 $X2=4.56
+ $Y2=0
r73 43 70 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r74 43 67 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=3.12
+ $Y2=0
r75 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r76 40 66 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.35 $Y=0 $X2=3.185
+ $Y2=0
r77 40 42 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=3.35 $Y=0 $X2=3.6
+ $Y2=0
r78 39 69 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=3.92 $Y=0 $X2=4.065
+ $Y2=0
r79 39 42 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=3.92 $Y=0 $X2=3.6
+ $Y2=0
r80 38 67 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=0 $X2=3.12
+ $Y2=0
r81 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r82 35 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.45 $Y=0 $X2=2.285
+ $Y2=0
r83 35 37 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=2.45 $Y=0 $X2=2.64
+ $Y2=0
r84 34 66 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.02 $Y=0 $X2=3.185
+ $Y2=0
r85 34 37 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=3.02 $Y=0 $X2=2.64
+ $Y2=0
r86 32 52 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r87 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r88 29 51 11.004 $w=1.7e-07 $l=4.5e-07 $layer=LI1_cond $X=0.525 $Y=0 $X2=0.975
+ $Y2=0
r89 29 31 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.525 $Y=0 $X2=0.24
+ $Y2=0
r90 27 38 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.4 $Y=0 $X2=2.64
+ $Y2=0
r91 27 64 0.0668963 $w=4.9e-07 $l=2.4e-07 $layer=MET1_cond $X=2.4 $Y=0 $X2=2.16
+ $Y2=0
r92 23 69 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=4.065 $Y=0.085
+ $X2=4.065 $Y2=0
r93 23 25 11.7231 $w=2.88e-07 $l=2.95e-07 $layer=LI1_cond $X=4.065 $Y=0.085
+ $X2=4.065 $Y2=0.38
r94 19 66 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.185 $Y=0.085
+ $X2=3.185 $Y2=0
r95 19 21 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=3.185 $Y=0.085
+ $X2=3.185 $Y2=0.36
r96 15 63 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.285 $Y=0.085
+ $X2=2.285 $Y2=0
r97 15 17 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.285 $Y=0.085
+ $X2=2.285 $Y2=0.36
r98 14 51 11.004 $w=1.7e-07 $l=4.5e-07 $layer=LI1_cond $X=1.425 $Y=0 $X2=0.975
+ $Y2=0
r99 13 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.12 $Y=0 $X2=2.285
+ $Y2=0
r100 13 14 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=2.12 $Y=0
+ $X2=1.425 $Y2=0
r101 4 25 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.905
+ $Y=0.235 $X2=4.045 $Y2=0.38
r102 3 21 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=3.045
+ $Y=0.235 $X2=3.185 $Y2=0.36
r103 2 17 91 $w=1.7e-07 $l=2.44643e-07 $layer=licon1_NDIFF $count=2 $X=2.095
+ $Y=0.235 $X2=2.285 $Y2=0.36
r104 1 60 182 $w=1.7e-07 $l=2.4e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.655 $X2=0.69 $Y2=0.835
r105 1 58 182 $w=1.7e-07 $l=7.77689e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.655 $X2=1.27 $Y2=0.775
r106 1 56 182 $w=1.7e-07 $l=8.46404e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.655 $X2=1.27 $Y2=0.38
.ends

