# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_lp__ha_lp
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_lp__ha_lp ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.280000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  0.626000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.785000 1.450000 3.205000 1.780000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.626000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.215000 1.605000 2.545000 1.960000 ;
        RECT 2.215000 1.960000 3.685000 2.130000 ;
        RECT 2.215000 2.130000 2.755000 2.890000 ;
        RECT 3.385000 1.605000 3.685000 1.960000 ;
    END
  END B
  PIN COUT
    ANTENNADIFFAREA  0.402600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.745000 2.075000 5.170000 3.065000 ;
        RECT 4.840000 0.440000 5.170000 1.045000 ;
        RECT 4.925000 1.045000 5.170000 2.075000 ;
    END
  END COUT
  PIN SUM
    ANTENNADIFFAREA  0.402600 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.110000 0.440000 0.440000 2.865000 ;
        RECT 0.110000 2.865000 0.975000 3.035000 ;
        RECT 0.645000 2.155000 0.975000 2.865000 ;
    END
  END SUM
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 5.280000 0.245000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 5.280000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.280000 0.085000 ;
      RECT 0.000000  3.245000 5.280000 3.415000 ;
      RECT 0.870000  1.565000 1.500000 1.725000 ;
      RECT 0.870000  1.725000 2.035000 1.895000 ;
      RECT 0.900000  0.085000 1.150000 1.335000 ;
      RECT 1.175000  2.075000 1.505000 3.245000 ;
      RECT 1.330000  0.265000 1.640000 0.645000 ;
      RECT 1.330000  0.645000 1.500000 1.565000 ;
      RECT 1.680000  1.100000 3.590000 1.225000 ;
      RECT 1.680000  1.225000 4.685000 1.270000 ;
      RECT 1.680000  1.270000 1.985000 1.430000 ;
      RECT 1.705000  1.895000 2.035000 3.065000 ;
      RECT 1.820000  0.265000 2.070000 0.750000 ;
      RECT 1.820000  0.750000 3.010000 0.920000 ;
      RECT 2.250000  0.085000 2.580000 0.570000 ;
      RECT 2.760000  0.265000 3.010000 0.750000 ;
      RECT 3.010000  2.310000 3.340000 3.245000 ;
      RECT 3.260000  0.605000 3.590000 1.100000 ;
      RECT 3.420000  1.270000 4.685000 1.395000 ;
      RECT 3.590000  2.310000 4.035000 3.065000 ;
      RECT 3.865000  1.395000 4.035000 2.310000 ;
      RECT 4.050000  0.085000 4.380000 1.045000 ;
      RECT 4.215000  2.075000 4.545000 3.245000 ;
      RECT 4.355000  1.395000 4.685000 1.895000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
  END
END sky130_fd_sc_lp__ha_lp
