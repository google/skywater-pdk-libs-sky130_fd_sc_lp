* File: sky130_fd_sc_lp__and4_lp2.pex.spice
* Created: Fri Aug 28 10:07:53 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__AND4_LP2%A_84_21# 1 2 3 10 12 15 19 22 24 25 26 28
+ 29 31 32 35 39 43 49 54 55 56
c109 31 0 6.1916e-20 $X=1.225 $Y=2.055
c110 15 0 1.86771e-19 $X=0.56 $Y=2.545
r111 53 54 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.615
+ $Y=1.105 $X2=0.615 $Y2=1.105
r112 47 49 10.4768 $w=3.28e-07 $l=3e-07 $layer=LI1_cond $X=2.78 $Y=0.77 $X2=2.78
+ $Y2=0.47
r113 43 45 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=2.53 $Y=2.19
+ $X2=2.53 $Y2=2.9
r114 41 43 1.74613 $w=3.28e-07 $l=5e-08 $layer=LI1_cond $X=2.53 $Y=2.14 $X2=2.53
+ $Y2=2.19
r115 40 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.555 $Y=2.055
+ $X2=1.39 $Y2=2.055
r116 39 41 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.365 $Y=2.055
+ $X2=2.53 $Y2=2.14
r117 39 40 52.8449 $w=1.68e-07 $l=8.1e-07 $layer=LI1_cond $X=2.365 $Y=2.055
+ $X2=1.555 $Y2=2.055
r118 35 37 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=1.39 $Y=2.19
+ $X2=1.39 $Y2=2.9
r119 33 56 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.39 $Y=2.14
+ $X2=1.39 $Y2=2.055
r120 33 35 1.74613 $w=3.28e-07 $l=5e-08 $layer=LI1_cond $X=1.39 $Y=2.14 $X2=1.39
+ $Y2=2.19
r121 31 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.225 $Y=2.055
+ $X2=1.39 $Y2=2.055
r122 31 32 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=1.225 $Y=2.055
+ $X2=0.81 $Y2=2.055
r123 30 53 11.4232 $w=2.67e-07 $l=3.27872e-07 $layer=LI1_cond $X=0.81 $Y=0.855
+ $X2=0.63 $Y2=1.105
r124 29 47 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.615 $Y=0.855
+ $X2=2.78 $Y2=0.77
r125 29 30 117.759 $w=1.68e-07 $l=1.805e-06 $layer=LI1_cond $X=2.615 $Y=0.855
+ $X2=0.81 $Y2=0.855
r126 28 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.725 $Y=1.97
+ $X2=0.81 $Y2=2.055
r127 28 55 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=0.725 $Y=1.97
+ $X2=0.725 $Y2=1.61
r128 26 55 8.99121 $w=3.58e-07 $l=1.8e-07 $layer=LI1_cond $X=0.63 $Y=1.43
+ $X2=0.63 $Y2=1.61
r129 25 53 1.34795 $w=3.6e-07 $l=1.5e-08 $layer=LI1_cond $X=0.63 $Y=1.12
+ $X2=0.63 $Y2=1.105
r130 25 26 9.92381 $w=3.58e-07 $l=3.1e-07 $layer=LI1_cond $X=0.63 $Y=1.12
+ $X2=0.63 $Y2=1.43
r131 23 54 55.6971 $w=3.45e-07 $l=3.33e-07 $layer=POLY_cond $X=0.607 $Y=1.438
+ $X2=0.607 $Y2=1.105
r132 23 24 33.2433 $w=3.45e-07 $l=1.72e-07 $layer=POLY_cond $X=0.607 $Y=1.438
+ $X2=0.607 $Y2=1.61
r133 22 54 37.6332 $w=3.45e-07 $l=2.25e-07 $layer=POLY_cond $X=0.607 $Y=0.88
+ $X2=0.607 $Y2=1.105
r134 15 24 232.304 $w=2.5e-07 $l=9.35e-07 $layer=POLY_cond $X=0.56 $Y=2.545
+ $X2=0.56 $Y2=1.61
r135 10 22 26.2249 $w=3.45e-07 $l=1.5e-07 $layer=POLY_cond $X=0.675 $Y=0.73
+ $X2=0.675 $Y2=0.88
r136 10 19 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.855 $Y=0.73
+ $X2=0.855 $Y2=0.445
r137 10 12 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.495 $Y=0.73
+ $X2=0.495 $Y2=0.445
r138 3 45 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=2.39
+ $Y=2.045 $X2=2.53 $Y2=2.9
r139 3 43 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.39
+ $Y=2.045 $X2=2.53 $Y2=2.19
r140 2 37 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=1.25
+ $Y=2.045 $X2=1.39 $Y2=2.9
r141 2 35 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=1.25
+ $Y=2.045 $X2=1.39 $Y2=2.19
r142 1 49 182 $w=1.7e-07 $l=2.96859e-07 $layer=licon1_NDIFF $count=1 $X=2.64
+ $Y=0.235 $X2=2.78 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_LP__AND4_LP2%D 3 7 9 11 12 13 16 18 19 23
c54 18 0 1.86771e-19 $X=1.2 $Y=1.295
c55 13 0 6.1916e-20 $X=1.155 $Y=1.79
c56 3 0 1.08032e-19 $X=1.125 $Y=2.545
r57 18 19 13.2706 $w=3.28e-07 $l=3.8e-07 $layer=LI1_cond $X=1.155 $Y=1.285
+ $X2=1.155 $Y2=1.665
r58 18 23 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.155
+ $Y=1.285 $X2=1.155 $Y2=1.285
r59 14 16 76.9149 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=1.245 $Y=0.805
+ $X2=1.395 $Y2=0.805
r60 12 23 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.155 $Y=1.625
+ $X2=1.155 $Y2=1.285
r61 12 13 31.6748 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.155 $Y=1.625
+ $X2=1.155 $Y2=1.79
r62 11 23 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.155 $Y=1.12
+ $X2=1.155 $Y2=1.285
r63 7 16 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.395 $Y=0.73
+ $X2=1.395 $Y2=0.805
r64 7 9 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=1.395 $Y=0.73 $X2=1.395
+ $Y2=0.445
r65 5 14 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.245 $Y=0.88
+ $X2=1.245 $Y2=0.805
r66 5 11 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=1.245 $Y=0.88
+ $X2=1.245 $Y2=1.12
r67 3 13 187.582 $w=2.5e-07 $l=7.55e-07 $layer=POLY_cond $X=1.125 $Y=2.545
+ $X2=1.125 $Y2=1.79
.ends

.subckt PM_SKY130_FD_SC_LP__AND4_LP2%C 3 7 11 12 13 14 18
r40 13 14 13.2706 $w=3.28e-07 $l=3.8e-07 $layer=LI1_cond $X=1.695 $Y=1.285
+ $X2=1.695 $Y2=1.665
r41 13 18 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.695
+ $Y=1.285 $X2=1.695 $Y2=1.285
r42 11 18 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=1.695 $Y=1.625
+ $X2=1.695 $Y2=1.285
r43 11 12 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.695 $Y=1.625
+ $X2=1.695 $Y2=1.79
r44 10 18 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.695 $Y=1.12
+ $X2=1.695 $Y2=1.285
r45 7 10 346.117 $w=1.5e-07 $l=6.75e-07 $layer=POLY_cond $X=1.785 $Y=0.445
+ $X2=1.785 $Y2=1.12
r46 3 12 187.582 $w=2.5e-07 $l=7.55e-07 $layer=POLY_cond $X=1.655 $Y=2.545
+ $X2=1.655 $Y2=1.79
.ends

.subckt PM_SKY130_FD_SC_LP__AND4_LP2%B 3 5 7 11 12 13 17 18
r40 17 18 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.265
+ $Y=1.285 $X2=2.265 $Y2=1.285
r41 12 13 11.0754 $w=3.83e-07 $l=3.7e-07 $layer=LI1_cond $X=2.237 $Y=1.295
+ $X2=2.237 $Y2=1.665
r42 12 18 0.299336 $w=3.83e-07 $l=1e-08 $layer=LI1_cond $X=2.237 $Y=1.295
+ $X2=2.237 $Y2=1.285
r43 11 17 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.265 $Y=1.625
+ $X2=2.265 $Y2=1.285
r44 10 17 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.265 $Y=1.12
+ $X2=2.265 $Y2=1.285
r45 5 11 30.6163 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.265 $Y=1.79
+ $X2=2.265 $Y2=1.625
r46 5 7 187.582 $w=2.5e-07 $l=7.55e-07 $layer=POLY_cond $X=2.265 $Y=1.79
+ $X2=2.265 $Y2=2.545
r47 3 10 346.117 $w=1.5e-07 $l=6.75e-07 $layer=POLY_cond $X=2.175 $Y=0.445
+ $X2=2.175 $Y2=1.12
.ends

.subckt PM_SKY130_FD_SC_LP__AND4_LP2%A 1 3 8 12 15 16 17 18 19 23 24
r36 23 24 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.835
+ $Y=1.285 $X2=2.835 $Y2=1.285
r37 18 19 7.83273 $w=5.63e-07 $l=3.7e-07 $layer=LI1_cond $X=2.952 $Y=1.295
+ $X2=2.952 $Y2=1.665
r38 18 24 0.211695 $w=5.63e-07 $l=1e-08 $layer=LI1_cond $X=2.952 $Y=1.295
+ $X2=2.952 $Y2=1.285
r39 16 23 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.835 $Y=1.625
+ $X2=2.835 $Y2=1.285
r40 16 17 32.3805 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.835 $Y=1.625
+ $X2=2.835 $Y2=1.79
r41 15 23 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.835 $Y=1.12
+ $X2=2.835 $Y2=1.285
r42 10 12 92.2979 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=2.565 $Y=0.805
+ $X2=2.745 $Y2=0.805
r43 8 17 187.582 $w=2.5e-07 $l=7.55e-07 $layer=POLY_cond $X=2.795 $Y=2.545
+ $X2=2.795 $Y2=1.79
r44 4 12 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.745 $Y=0.88
+ $X2=2.745 $Y2=0.805
r45 4 15 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=2.745 $Y=0.88
+ $X2=2.745 $Y2=1.12
r46 1 10 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.565 $Y=0.73
+ $X2=2.565 $Y2=0.805
r47 1 3 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.565 $Y=0.73 $X2=2.565
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_LP__AND4_LP2%X 1 2 10 13 14 15 31 33
c22 13 0 1.08032e-19 $X=0.155 $Y=1.95
r23 20 33 2.0808 $w=3.58e-07 $l=6.5e-08 $layer=LI1_cond $X=0.28 $Y=2.1 $X2=0.28
+ $Y2=2.035
r24 15 28 4.00154 $w=3.58e-07 $l=1.25e-07 $layer=LI1_cond $X=0.28 $Y=2.775
+ $X2=0.28 $Y2=2.9
r25 14 15 11.8446 $w=3.58e-07 $l=3.7e-07 $layer=LI1_cond $X=0.28 $Y=2.405
+ $X2=0.28 $Y2=2.775
r26 13 33 0.320123 $w=3.58e-07 $l=1e-08 $layer=LI1_cond $X=0.28 $Y=2.025
+ $X2=0.28 $Y2=2.035
r27 13 31 6.59029 $w=3.58e-07 $l=1.05e-07 $layer=LI1_cond $X=0.28 $Y=2.025
+ $X2=0.28 $Y2=1.92
r28 13 14 9.44363 $w=3.58e-07 $l=2.95e-07 $layer=LI1_cond $X=0.28 $Y=2.11
+ $X2=0.28 $Y2=2.405
r29 13 20 0.320123 $w=3.58e-07 $l=1e-08 $layer=LI1_cond $X=0.28 $Y=2.11 $X2=0.28
+ $Y2=2.1
r30 12 31 81.2246 $w=1.68e-07 $l=1.245e-06 $layer=LI1_cond $X=0.185 $Y=0.675
+ $X2=0.185 $Y2=1.92
r31 10 12 9.81557 $w=3.43e-07 $l=2.05e-07 $layer=LI1_cond $X=0.272 $Y=0.47
+ $X2=0.272 $Y2=0.675
r32 2 28 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.15
+ $Y=2.045 $X2=0.295 $Y2=2.9
r33 2 13 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.15
+ $Y=2.045 $X2=0.295 $Y2=2.19
r34 1 10 182 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.28 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_LP__AND4_LP2%VPWR 1 2 3 14 18 20 22 27 28 29 35 40 44
r47 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r48 40 41 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r49 38 44 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r50 37 38 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r51 35 43 4.69206 $w=1.7e-07 $l=2.32e-07 $layer=LI1_cond $X=2.895 $Y=3.33
+ $X2=3.127 $Y2=3.33
r52 35 37 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=2.895 $Y=3.33
+ $X2=2.64 $Y2=3.33
r53 31 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.99 $Y=3.33
+ $X2=0.825 $Y2=3.33
r54 31 33 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=0.99 $Y=3.33 $X2=1.68
+ $Y2=3.33
r55 29 38 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r56 29 41 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=0.72 $Y2=3.33
r57 29 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.68 $Y=3.33
+ $X2=1.68 $Y2=3.33
r58 27 33 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=1.755 $Y=3.33
+ $X2=1.68 $Y2=3.33
r59 27 28 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.755 $Y=3.33
+ $X2=1.92 $Y2=3.33
r60 26 37 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=2.085 $Y=3.33
+ $X2=2.64 $Y2=3.33
r61 26 28 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.085 $Y=3.33
+ $X2=1.92 $Y2=3.33
r62 22 25 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=3.06 $Y=2.19 $X2=3.06
+ $Y2=2.9
r63 20 43 3.07411 $w=3.3e-07 $l=1.13666e-07 $layer=LI1_cond $X=3.06 $Y=3.245
+ $X2=3.127 $Y2=3.33
r64 20 25 12.0483 $w=3.28e-07 $l=3.45e-07 $layer=LI1_cond $X=3.06 $Y=3.245
+ $X2=3.06 $Y2=2.9
r65 16 28 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.92 $Y=3.245
+ $X2=1.92 $Y2=3.33
r66 16 18 26.5411 $w=3.28e-07 $l=7.6e-07 $layer=LI1_cond $X=1.92 $Y=3.245
+ $X2=1.92 $Y2=2.485
r67 12 40 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.825 $Y=3.245
+ $X2=0.825 $Y2=3.33
r68 12 14 26.5411 $w=3.28e-07 $l=7.6e-07 $layer=LI1_cond $X=0.825 $Y=3.245
+ $X2=0.825 $Y2=2.485
r69 3 25 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=2.92
+ $Y=2.045 $X2=3.06 $Y2=2.9
r70 3 22 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.92
+ $Y=2.045 $X2=3.06 $Y2=2.19
r71 2 18 300 $w=1.7e-07 $l=5.05173e-07 $layer=licon1_PDIFF $count=2 $X=1.78
+ $Y=2.045 $X2=1.92 $Y2=2.485
r72 1 14 300 $w=1.7e-07 $l=5.05173e-07 $layer=licon1_PDIFF $count=2 $X=0.685
+ $Y=2.045 $X2=0.825 $Y2=2.485
.ends

.subckt PM_SKY130_FD_SC_LP__AND4_LP2%VGND 1 6 8 10 17 18 21
r37 21 22 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r38 17 18 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r39 15 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.235 $Y=0 $X2=1.07
+ $Y2=0
r40 15 17 122.979 $w=1.68e-07 $l=1.885e-06 $layer=LI1_cond $X=1.235 $Y=0
+ $X2=3.12 $Y2=0
r41 13 22 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r42 12 13 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r43 10 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.905 $Y=0 $X2=1.07
+ $Y2=0
r44 10 12 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=0.905 $Y=0 $X2=0.72
+ $Y2=0
r45 8 18 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=1.68 $Y=0 $X2=3.12
+ $Y2=0
r46 8 22 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r47 4 21 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.07 $Y=0.085 $X2=1.07
+ $Y2=0
r48 4 6 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=1.07 $Y=0.085
+ $X2=1.07 $Y2=0.4
r49 1 6 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=0.93
+ $Y=0.235 $X2=1.07 $Y2=0.4
.ends

