# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO sky130_fd_sc_lp__nand3_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_lp__nand3_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.760000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.395000 1.310000 1.750000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.170000 1.425000 3.180000 1.605000 ;
        RECT 2.795000 1.605000 3.180000 1.920000 ;
        RECT 2.795000 1.920000 5.430000 2.120000 ;
        RECT 5.200000 1.425000 5.540000 1.705000 ;
        RECT 5.200000 1.705000 5.430000 1.920000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  1.260000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.390000 1.425000 4.930000 1.750000 ;
    END
  END C
  PIN Y
    ANTENNADIFFAREA  2.587200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.595000 0.595000 0.815000 1.055000 ;
        RECT 0.595000 1.055000 1.710000 1.225000 ;
        RECT 0.645000 1.920000 2.625000 1.945000 ;
        RECT 0.645000 1.945000 1.695000 2.100000 ;
        RECT 0.645000 2.100000 0.835000 3.075000 ;
        RECT 1.485000 0.595000 1.710000 1.055000 ;
        RECT 1.495000 1.225000 1.710000 1.425000 ;
        RECT 1.495000 1.425000 2.000000 1.775000 ;
        RECT 1.495000 1.775000 2.625000 1.920000 ;
        RECT 1.505000 2.100000 1.695000 3.075000 ;
        RECT 2.365000 1.945000 2.625000 2.290000 ;
        RECT 2.365000 2.290000 5.165000 2.460000 ;
        RECT 2.365000 2.460000 2.545000 3.075000 ;
        RECT 3.225000 2.460000 3.415000 3.075000 ;
        RECT 4.105000 2.460000 4.305000 3.075000 ;
        RECT 4.975000 2.460000 5.165000 3.075000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 5.760000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.000000 0.000000 5.760000 0.245000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.655000 5.950000 3.520000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 5.760000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.760000 0.085000 ;
      RECT 0.000000  3.245000 5.760000 3.415000 ;
      RECT 0.125000  0.255000 2.105000 0.425000 ;
      RECT 0.125000  0.425000 0.425000 1.145000 ;
      RECT 0.145000  1.920000 0.475000 3.245000 ;
      RECT 0.985000  0.425000 1.315000 0.885000 ;
      RECT 1.005000  2.270000 1.335000 3.245000 ;
      RECT 1.865000  2.115000 2.195000 3.245000 ;
      RECT 1.880000  0.425000 2.105000 1.085000 ;
      RECT 1.880000  1.085000 5.665000 1.255000 ;
      RECT 2.275000  0.255000 3.505000 0.425000 ;
      RECT 2.275000  0.425000 2.605000 0.915000 ;
      RECT 2.725000  2.630000 3.055000 3.245000 ;
      RECT 2.775000  0.645000 3.005000 1.085000 ;
      RECT 3.175000  0.425000 3.505000 0.745000 ;
      RECT 3.175000  0.745000 5.235000 0.915000 ;
      RECT 3.585000  2.630000 3.915000 3.245000 ;
      RECT 3.675000  0.085000 3.945000 0.575000 ;
      RECT 4.065000  0.700000 4.355000 0.745000 ;
      RECT 4.475000  0.085000 4.805000 0.575000 ;
      RECT 4.475000  2.630000 4.805000 3.245000 ;
      RECT 4.930000  0.700000 5.235000 0.745000 ;
      RECT 5.335000  2.290000 5.665000 3.245000 ;
      RECT 5.405000  0.265000 5.665000 1.085000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
  END
END sky130_fd_sc_lp__nand3_4
END LIBRARY
