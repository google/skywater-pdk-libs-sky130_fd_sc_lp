* File: sky130_fd_sc_lp__nor4b_4.spice
* Created: Wed Sep  2 10:11:09 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__nor4b_4.pex.spice"
.subckt sky130_fd_sc_lp__nor4b_4  VNB VPB D_N C B A VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A	A
* B	B
* C	C
* D_N	D_N
* VPB	VPB
* VNB	VNB
MM1027 N_VGND_M1027_d N_D_N_M1027_g N_A_27_367#_M1027_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1386 AS=0.2226 PD=1.17 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75008.1 A=0.126 P=1.98 MULT=1
MM1004 N_VGND_M1027_d N_A_27_367#_M1004_g N_Y_M1004_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1386 AS=0.1176 PD=1.17 PS=1.12 NRD=7.14 NRS=0 M=1 R=5.6 SA=75000.7
+ SB=75007.6 A=0.126 P=1.98 MULT=1
MM1009 N_VGND_M1009_d N_A_27_367#_M1009_g N_Y_M1004_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1386 AS=0.1176 PD=1.17 PS=1.12 NRD=2.856 NRS=0 M=1 R=5.6 SA=75001.1
+ SB=75007.1 A=0.126 P=1.98 MULT=1
MM1024 N_VGND_M1009_d N_A_27_367#_M1024_g N_Y_M1024_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1386 AS=0.1176 PD=1.17 PS=1.12 NRD=4.284 NRS=0 M=1 R=5.6 SA=75001.6
+ SB=75006.7 A=0.126 P=1.98 MULT=1
MM1029 N_VGND_M1029_d N_A_27_367#_M1029_g N_Y_M1024_s VNB NSHORT L=0.15 W=0.84
+ AD=0.2646 AS=0.1176 PD=1.47 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002 SB=75006.2
+ A=0.126 P=1.98 MULT=1
MM1001 N_VGND_M1029_d N_C_M1001_g N_Y_M1001_s VNB NSHORT L=0.15 W=0.84 AD=0.2646
+ AS=0.1176 PD=1.47 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75002.8 SB=75005.5 A=0.126
+ P=1.98 MULT=1
MM1016 N_VGND_M1016_d N_C_M1016_g N_Y_M1001_s VNB NSHORT L=0.15 W=0.84 AD=0.1176
+ AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75003.2 SB=75005 A=0.126
+ P=1.98 MULT=1
MM1025 N_VGND_M1016_d N_C_M1025_g N_Y_M1025_s VNB NSHORT L=0.15 W=0.84 AD=0.1176
+ AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75003.6 SB=75004.6 A=0.126
+ P=1.98 MULT=1
MM1030 N_VGND_M1030_d N_C_M1030_g N_Y_M1025_s VNB NSHORT L=0.15 W=0.84 AD=0.3276
+ AS=0.1176 PD=1.62 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75004.1 SB=75004.2 A=0.126
+ P=1.98 MULT=1
MM1000 N_Y_M1000_d N_B_M1000_g N_VGND_M1030_d VNB NSHORT L=0.15 W=0.84 AD=0.1176
+ AS=0.3276 PD=1.12 PS=1.62 NRD=0 NRS=0 M=1 R=5.6 SA=75005 SB=75003.2 A=0.126
+ P=1.98 MULT=1
MM1003 N_Y_M1000_d N_B_M1003_g N_VGND_M1003_s VNB NSHORT L=0.15 W=0.84 AD=0.1176
+ AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75005.4 SB=75002.8 A=0.126
+ P=1.98 MULT=1
MM1015 N_Y_M1015_d N_B_M1015_g N_VGND_M1003_s VNB NSHORT L=0.15 W=0.84 AD=0.1176
+ AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75005.9 SB=75002.4 A=0.126
+ P=1.98 MULT=1
MM1017 N_Y_M1015_d N_B_M1017_g N_VGND_M1017_s VNB NSHORT L=0.15 W=0.84 AD=0.1176
+ AS=0.1218 PD=1.12 PS=1.13 NRD=0 NRS=0 M=1 R=5.6 SA=75006.3 SB=75001.9 A=0.126
+ P=1.98 MULT=1
MM1011 N_VGND_M1017_s N_A_M1011_g N_Y_M1011_s VNB NSHORT L=0.15 W=0.84 AD=0.1218
+ AS=0.1302 PD=1.13 PS=1.15 NRD=1.428 NRS=1.428 M=1 R=5.6 SA=75006.7 SB=75001.5
+ A=0.126 P=1.98 MULT=1
MM1013 N_VGND_M1013_d N_A_M1013_g N_Y_M1011_s VNB NSHORT L=0.15 W=0.84 AD=0.1176
+ AS=0.1302 PD=1.12 PS=1.15 NRD=0 NRS=2.856 M=1 R=5.6 SA=75007.2 SB=75001.1
+ A=0.126 P=1.98 MULT=1
MM1022 N_VGND_M1013_d N_A_M1022_g N_Y_M1022_s VNB NSHORT L=0.15 W=0.84 AD=0.1176
+ AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75007.6 SB=75000.6 A=0.126
+ P=1.98 MULT=1
MM1028 N_VGND_M1028_d N_A_M1028_g N_Y_M1022_s VNB NSHORT L=0.15 W=0.84 AD=0.2226
+ AS=0.1176 PD=2.21 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75008.1 SB=75000.2 A=0.126
+ P=1.98 MULT=1
MM1033 N_VPWR_M1033_d N_D_N_M1033_g N_A_27_367#_M1033_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.3339 PD=3.05 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75000.2 A=0.189 P=2.82 MULT=1
MM1005 N_Y_M1005_d N_A_27_367#_M1005_g N_A_217_367#_M1005_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75003.2 A=0.189 P=2.82 MULT=1
MM1006 N_Y_M1005_d N_A_27_367#_M1006_g N_A_217_367#_M1006_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75002.8 A=0.189 P=2.82 MULT=1
MM1018 N_Y_M1018_d N_A_27_367#_M1018_g N_A_217_367#_M1006_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75002.3 A=0.189 P=2.82 MULT=1
MM1031 N_Y_M1018_d N_A_27_367#_M1031_g N_A_217_367#_M1031_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.5
+ SB=75001.9 A=0.189 P=2.82 MULT=1
MM1008 N_A_217_367#_M1031_s N_C_M1008_g N_A_644_367#_M1008_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.9
+ SB=75001.5 A=0.189 P=2.82 MULT=1
MM1012 N_A_217_367#_M1012_d N_C_M1012_g N_A_644_367#_M1008_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.3
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1021 N_A_217_367#_M1012_d N_C_M1021_g N_A_644_367#_M1021_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.8
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1023 N_A_217_367#_M1023_d N_C_M1023_g N_A_644_367#_M1021_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75003.2
+ SB=75000.2 A=0.189 P=2.82 MULT=1
MM1007 N_A_1009_367#_M1007_d N_B_M1007_g N_A_644_367#_M1007_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75003.2 A=0.189 P=2.82 MULT=1
MM1014 N_A_1009_367#_M1014_d N_B_M1014_g N_A_644_367#_M1007_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75002.8 A=0.189 P=2.82 MULT=1
MM1019 N_A_1009_367#_M1014_d N_B_M1019_g N_A_644_367#_M1019_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75002.3 A=0.189 P=2.82 MULT=1
MM1026 N_A_1009_367#_M1026_d N_B_M1026_g N_A_644_367#_M1019_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.5
+ SB=75001.9 A=0.189 P=2.82 MULT=1
MM1002 N_VPWR_M1002_d N_A_M1002_g N_A_1009_367#_M1026_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.9
+ SB=75001.5 A=0.189 P=2.82 MULT=1
MM1010 N_VPWR_M1002_d N_A_M1010_g N_A_1009_367#_M1010_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.3
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1020 N_VPWR_M1020_d N_A_M1020_g N_A_1009_367#_M1010_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.8
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1032 N_VPWR_M1020_d N_A_M1032_g N_A_1009_367#_M1032_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4 SA=75003.2
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX34_noxref VNB VPB NWDIODE A=17.7175 P=22.73
*
.include "sky130_fd_sc_lp__nor4b_4.pxi.spice"
*
.ends
*
*
