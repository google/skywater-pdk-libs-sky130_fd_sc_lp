# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
MACRO sky130_fd_sc_lp__o211a_4
  CLASS CORE ;
  SOURCE USER ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.720000 BY  3.330000 ;
  SYMMETRY X Y R90 ;
  SITE unit ;
  PIN A1
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.670000 1.195000 6.635000 1.255000 ;
        RECT 4.670000 1.255000 5.000000 1.525000 ;
        RECT 4.830000 1.085000 6.635000 1.195000 ;
        RECT 6.315000 1.255000 6.635000 1.760000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.210000 1.425000 6.145000 1.760000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.545000 1.405000 3.275000 1.930000 ;
        RECT 2.545000 1.930000 4.460000 2.100000 ;
        RECT 4.130000 1.345000 4.460000 1.930000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  0.630000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.445000 1.405000 3.920000 1.760000 ;
    END
  END C1
  PIN X
    ANTENNADIFFAREA  1.176000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.045000 1.655000 1.215000 ;
        RECT 0.085000 1.215000 0.370000 1.755000 ;
        RECT 0.085000 1.755000 2.035000 1.925000 ;
        RECT 0.595000 0.255000 0.785000 1.045000 ;
        RECT 0.985000 1.925000 1.165000 3.075000 ;
        RECT 1.455000 0.255000 1.655000 1.045000 ;
        RECT 1.845000 1.925000 2.035000 3.075000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.245000 6.720000 0.245000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 0.000000 0.500000 0.500000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.800000 0.500000 3.300000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 3.085000 6.720000 3.575000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.720000 0.085000 ;
      RECT 0.000000  3.245000 6.720000 3.415000 ;
      RECT 0.095000  0.085000 0.425000 0.875000 ;
      RECT 0.485000  2.095000 0.815000 3.245000 ;
      RECT 0.540000  1.385000 2.375000 1.585000 ;
      RECT 0.955000  0.085000 1.285000 0.875000 ;
      RECT 1.345000  2.095000 1.675000 3.245000 ;
      RECT 1.850000  0.085000 2.085000 0.940000 ;
      RECT 2.205000  1.065000 3.700000 1.235000 ;
      RECT 2.205000  1.235000 2.375000 1.385000 ;
      RECT 2.205000  1.585000 2.375000 2.270000 ;
      RECT 2.205000  2.270000 5.665000 2.440000 ;
      RECT 2.205000  2.610000 2.535000 3.245000 ;
      RECT 2.335000  0.255000 2.665000 0.635000 ;
      RECT 2.335000  0.635000 4.665000 0.745000 ;
      RECT 2.335000  0.745000 6.525000 0.805000 ;
      RECT 2.335000  0.805000 2.665000 0.895000 ;
      RECT 2.705000  2.440000 3.295000 3.075000 ;
      RECT 2.845000  0.255000 4.225000 0.465000 ;
      RECT 3.370000  0.975000 3.700000 1.065000 ;
      RECT 3.465000  2.610000 3.795000 3.245000 ;
      RECT 3.965000  2.440000 4.300000 3.075000 ;
      RECT 4.365000  0.805000 6.525000 0.915000 ;
      RECT 4.365000  0.915000 4.660000 1.025000 ;
      RECT 4.395000  0.255000 4.665000 0.635000 ;
      RECT 4.470000  2.610000 4.735000 3.245000 ;
      RECT 4.835000  0.085000 5.165000 0.575000 ;
      RECT 4.905000  2.780000 6.025000 3.075000 ;
      RECT 5.335000  0.255000 5.665000 0.745000 ;
      RECT 5.335000  1.930000 5.665000 2.270000 ;
      RECT 5.335000  2.440000 5.665000 2.610000 ;
      RECT 5.835000  0.085000 6.025000 0.575000 ;
      RECT 5.835000  1.930000 6.025000 2.780000 ;
      RECT 6.195000  0.255000 6.525000 0.745000 ;
      RECT 6.195000  1.930000 6.525000 3.245000 ;
    LAYER mcon ;
      RECT 0.155000 -0.085000 0.325000 0.085000 ;
      RECT 0.155000  3.245000 0.325000 3.415000 ;
      RECT 0.635000 -0.085000 0.805000 0.085000 ;
      RECT 0.635000  3.245000 0.805000 3.415000 ;
      RECT 1.115000 -0.085000 1.285000 0.085000 ;
      RECT 1.115000  3.245000 1.285000 3.415000 ;
      RECT 1.595000 -0.085000 1.765000 0.085000 ;
      RECT 1.595000  3.245000 1.765000 3.415000 ;
      RECT 2.075000 -0.085000 2.245000 0.085000 ;
      RECT 2.075000  3.245000 2.245000 3.415000 ;
      RECT 2.555000 -0.085000 2.725000 0.085000 ;
      RECT 2.555000  3.245000 2.725000 3.415000 ;
      RECT 3.035000 -0.085000 3.205000 0.085000 ;
      RECT 3.035000  3.245000 3.205000 3.415000 ;
      RECT 3.515000 -0.085000 3.685000 0.085000 ;
      RECT 3.515000  3.245000 3.685000 3.415000 ;
      RECT 3.995000 -0.085000 4.165000 0.085000 ;
      RECT 3.995000  3.245000 4.165000 3.415000 ;
      RECT 4.475000 -0.085000 4.645000 0.085000 ;
      RECT 4.475000  3.245000 4.645000 3.415000 ;
      RECT 4.955000 -0.085000 5.125000 0.085000 ;
      RECT 4.955000  3.245000 5.125000 3.415000 ;
      RECT 5.435000 -0.085000 5.605000 0.085000 ;
      RECT 5.435000  3.245000 5.605000 3.415000 ;
      RECT 5.915000 -0.085000 6.085000 0.085000 ;
      RECT 5.915000  3.245000 6.085000 3.415000 ;
      RECT 6.395000 -0.085000 6.565000 0.085000 ;
      RECT 6.395000  3.245000 6.565000 3.415000 ;
  END
END sky130_fd_sc_lp__o211a_4
END LIBRARY
