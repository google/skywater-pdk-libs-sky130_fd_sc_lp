* File: sky130_fd_sc_lp__o221ai_2.spice
* Created: Fri Aug 28 11:08:37 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__o221ai_2.pex.spice"
.subckt sky130_fd_sc_lp__o221ai_2  VNB VPB C1 B1 B2 A1 A2 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A2	A2
* A1	A1
* B2	B2
* B1	B1
* C1	C1
* VPB	VPB
* VNB	VNB
MM1002 N_Y_M1002_d N_C1_M1002_g N_A_29_69#_M1002_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1005 N_Y_M1002_d N_C1_M1005_g N_A_29_69#_M1005_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1003 N_A_305_65#_M1003_d N_B1_M1003_g N_A_29_69#_M1003_s VNB NSHORT L=0.15
+ W=0.84 AD=0.2226 AS=0.147 PD=2.21 PS=1.19 NRD=0 NRS=9.996 M=1 R=5.6 SA=75000.2
+ SB=75003.5 A=0.126 P=1.98 MULT=1
MM1006 N_A_305_65#_M1006_d N_B2_M1006_g N_A_29_69#_M1003_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.147 PD=1.12 PS=1.19 NRD=0 NRS=0 M=1 R=5.6 SA=75000.7
+ SB=75003 A=0.126 P=1.98 MULT=1
MM1014 N_A_305_65#_M1006_d N_B2_M1014_g N_A_29_69#_M1014_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.189 PD=1.12 PS=1.29 NRD=0 NRS=13.56 M=1 R=5.6 SA=75001.1
+ SB=75002.6 A=0.126 P=1.98 MULT=1
MM1010 N_A_305_65#_M1010_d N_B1_M1010_g N_A_29_69#_M1014_s VNB NSHORT L=0.15
+ W=0.84 AD=0.1176 AS=0.189 PD=1.12 PS=1.29 NRD=0 NRS=10.704 M=1 R=5.6
+ SA=75001.7 SB=75002 A=0.126 P=1.98 MULT=1
MM1011 N_VGND_M1011_d N_A1_M1011_g N_A_305_65#_M1010_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1344 AS=0.1176 PD=1.16 PS=1.12 NRD=2.856 NRS=0 M=1 R=5.6 SA=75002.1
+ SB=75001.6 A=0.126 P=1.98 MULT=1
MM1009 N_A_305_65#_M1009_d N_A2_M1009_g N_VGND_M1011_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1344 PD=1.12 PS=1.16 NRD=0 NRS=2.856 M=1 R=5.6 SA=75002.6
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1017 N_A_305_65#_M1009_d N_A2_M1017_g N_VGND_M1017_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1344 PD=1.12 PS=1.16 NRD=0 NRS=2.856 M=1 R=5.6 SA=75003.1
+ SB=75000.7 A=0.126 P=1.98 MULT=1
MM1012 N_VGND_M1017_s N_A1_M1012_g N_A_305_65#_M1012_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1344 AS=0.2226 PD=1.16 PS=2.21 NRD=2.856 NRS=0 M=1 R=5.6 SA=75003.5
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1004 N_VPWR_M1004_d N_C1_M1004_g N_Y_M1004_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.2 SB=75005
+ A=0.189 P=2.82 MULT=1
MM1015 N_VPWR_M1015_d N_C1_M1015_g N_Y_M1004_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.504 AS=0.1764 PD=2.06 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6 SB=75004.5
+ A=0.189 P=2.82 MULT=1
MM1001 N_VPWR_M1015_d N_B1_M1001_g N_A_388_367#_M1001_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.504 AS=0.2205 PD=2.06 PS=1.61 NRD=0 NRS=5.4569 M=1 R=8.4
+ SA=75001.6 SB=75003.6 A=0.189 P=2.82 MULT=1
MM1007 N_A_388_367#_M1001_s N_B2_M1007_g N_Y_M1007_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.2205 AS=0.1764 PD=1.61 PS=1.54 NRD=5.4569 NRS=0 M=1 R=8.4 SA=75002.1
+ SB=75003.1 A=0.189 P=2.82 MULT=1
MM1019 N_A_388_367#_M1019_d N_B2_M1019_g N_Y_M1007_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75002.5
+ SB=75002.7 A=0.189 P=2.82 MULT=1
MM1013 N_VPWR_M1013_d N_B1_M1013_g N_A_388_367#_M1019_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3276 AS=0.1764 PD=1.78 PS=1.54 NRD=18.7544 NRS=0 M=1 R=8.4
+ SA=75002.9 SB=75002.2 A=0.189 P=2.82 MULT=1
MM1000 N_VPWR_M1013_d N_A1_M1000_g N_A_794_367#_M1000_s VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3276 AS=0.2268 PD=1.78 PS=1.62 NRD=18.7544 NRS=12.4898 M=1 R=8.4
+ SA=75003.6 SB=75001.6 A=0.189 P=2.82 MULT=1
MM1008 N_A_794_367#_M1000_s N_A2_M1008_g N_Y_M1008_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.2268 AS=0.1764 PD=1.62 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75004.1
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1018 N_A_794_367#_M1018_d N_A2_M1018_g N_Y_M1008_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75004.5
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1016 N_VPWR_M1016_d N_A1_M1016_g N_A_794_367#_M1018_d VPB PHIGHVT L=0.15
+ W=1.26 AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75005
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX20_noxref VNB VPB NWDIODE A=11.4511 P=16.01
*
.include "sky130_fd_sc_lp__o221ai_2.pxi.spice"
*
.ends
*
*
