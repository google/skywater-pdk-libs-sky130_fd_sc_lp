* NGSPICE file created from sky130_fd_sc_lp__dlrtn_4.ext - technology: sky130A

.subckt sky130_fd_sc_lp__dlrtn_4 D GATE_N RESET_B VGND VNB VPB VPWR Q
M1000 a_725_125# a_357_365# a_639_125# VNB nshort w=420000u l=150000u
+  ad=1.344e+11p pd=1.48e+06u as=1.176e+11p ps=1.4e+06u
M1001 a_250_70# GATE_N VGND VNB nshort w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=1.2075e+12p ps=1.137e+07u
M1002 VPWR a_250_70# a_357_365# VPB phighvt w=640000u l=150000u
+  ad=2.2795e+12p pd=1.789e+07u as=3.329e+11p ps=2.82e+06u
M1003 a_567_125# a_27_468# VGND VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1004 VGND a_789_99# a_725_125# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_250_70# GATE_N VPWR VPB phighvt w=640000u l=150000u
+  ad=1.696e+11p pd=1.81e+06u as=0p ps=0u
M1006 VPWR RESET_B a_789_99# VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=3.528e+11p ps=3.08e+06u
M1007 VPWR a_789_99# Q VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=7.182e+11p ps=6.18e+06u
M1008 VPWR a_789_99# a_748_447# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1009 VGND RESET_B a_1009_47# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=1.764e+11p ps=2.1e+06u
M1010 a_567_447# a_27_468# VPWR VPB phighvt w=640000u l=150000u
+  ad=1.344e+11p pd=1.7e+06u as=0p ps=0u
M1011 Q a_789_99# VGND VNB nshort w=840000u l=150000u
+  ad=4.704e+11p pd=4.48e+06u as=0p ps=0u
M1012 Q a_789_99# VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_639_125# a_357_365# a_567_447# VPB phighvt w=640000u l=150000u
+  ad=2.286e+11p pd=2.07e+06u as=0p ps=0u
M1014 Q a_789_99# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 Q a_789_99# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VGND D a_27_468# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.197e+11p ps=1.41e+06u
M1017 VGND a_250_70# a_357_365# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1018 a_1009_47# a_639_125# a_789_99# VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=2.226e+11p ps=2.21e+06u
M1019 a_789_99# a_639_125# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_748_447# a_250_70# a_639_125# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VGND a_789_99# Q VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VPWR D a_27_468# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.696e+11p ps=1.81e+06u
M1023 VGND a_789_99# Q VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_639_125# a_250_70# a_567_125# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 VPWR a_789_99# Q VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

