* NGSPICE file created from sky130_fd_sc_lp__and3b_1.ext - technology: sky130A

.subckt sky130_fd_sc_lp__and3b_1 A_N B C VGND VNB VPB VPWR X
M1000 X a_185_367# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=3.339e+11p pd=3.05e+06u as=6.447e+11p ps=6.21e+06u
M1001 VPWR C a_185_367# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=2.436e+11p ps=2.84e+06u
M1002 a_185_367# B VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_110_47# A_N VGND VNB nshort w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=4.557e+11p ps=4.16e+06u
M1004 VPWR a_110_47# a_185_367# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 X a_185_367# VGND VNB nshort w=840000u l=150000u
+  ad=2.226e+11p pd=2.21e+06u as=0p ps=0u
M1006 a_110_47# A_N VPWR VPB phighvt w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1007 a_304_47# a_110_47# a_185_367# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=1.113e+11p ps=1.37e+06u
M1008 a_376_47# B a_304_47# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1009 VGND C a_376_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

