* File: sky130_fd_sc_lp__dfrtp_4.spice
* Created: Fri Aug 28 10:22:30 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__dfrtp_4.pex.spice"
.subckt sky130_fd_sc_lp__dfrtp_4  VNB VPB CLK D RESET_B VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* RESET_B	RESET_B
* D	D
* CLK	CLK
* VPB	VPB
* VNB	VNB
MM1020 N_VGND_M1020_d N_CLK_M1020_g N_A_27_90#_M1020_s VNB NSHORT L=0.15 W=0.42
+ AD=0.1449 AS=0.1113 PD=1.11 PS=1.37 NRD=2.856 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.1 A=0.063 P=1.14 MULT=1
MM1021 N_A_216_462#_M1021_d N_A_27_90#_M1021_g N_VGND_M1020_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1197 AS=0.1449 PD=1.41 PS=1.11 NRD=5.712 NRS=114.276 M=1 R=2.8
+ SA=75001 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1022 A_531_119# N_RESET_B_M1022_g N_VGND_M1022_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1113 PD=0.63 PS=1.37 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75005.3 A=0.063 P=1.14 MULT=1
MM1018 N_A_340_535#_M1018_d N_D_M1018_g A_531_119# VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.6
+ SB=75005 A=0.063 P=1.14 MULT=1
MM1008 N_A_595_535#_M1008_d N_A_27_90#_M1008_g N_A_340_535#_M1018_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.1155 AS=0.0588 PD=0.97 PS=0.7 NRD=77.136 NRS=0 M=1 R=2.8
+ SA=75001 SB=75004.5 A=0.063 P=1.14 MULT=1
MM1031 A_829_119# N_A_216_462#_M1031_g N_A_595_535#_M1008_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0483 AS=0.1155 PD=0.65 PS=0.97 NRD=17.136 NRS=0 M=1 R=2.8
+ SA=75001.7 SB=75003.8 A=0.063 P=1.14 MULT=1
MM1033 A_905_119# N_A_731_405#_M1033_g A_829_119# VNB NSHORT L=0.15 W=0.42
+ AD=0.08575 AS=0.0483 PD=0.88 PS=0.65 NRD=42.612 NRS=17.136 M=1 R=2.8
+ SA=75002.1 SB=75003.4 A=0.063 P=1.14 MULT=1
MM1010 N_VGND_M1010_d N_RESET_B_M1010_g A_905_119# VNB NSHORT L=0.15 W=0.42
+ AD=0.139274 AS=0.08575 PD=1.04604 PS=0.88 NRD=79.02 NRS=42.612 M=1 R=2.8
+ SA=75002.2 SB=75003.3 A=0.063 P=1.14 MULT=1
MM1025 N_A_731_405#_M1025_d N_A_595_535#_M1025_g N_VGND_M1010_d VNB NSHORT
+ L=0.15 W=0.64 AD=0.1835 AS=0.212226 PD=1.29 PS=1.59396 NRD=22.488 NRS=22.5 M=1
+ R=4.26667 SA=75002 SB=75002.1 A=0.096 P=1.58 MULT=1
MM1012 N_A_1255_449#_M1012_d N_A_216_462#_M1012_g N_A_731_405#_M1025_d VNB
+ NSHORT L=0.15 W=0.64 AD=0.301162 AS=0.1835 PD=1.79925 PS=1.29 NRD=56.244
+ NRS=22.488 M=1 R=4.26667 SA=75002.6 SB=75001.5 A=0.096 P=1.58 MULT=1
MM1002 A_1449_133# N_A_27_90#_M1002_g N_A_1255_449#_M1012_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0819 AS=0.197638 PD=0.81 PS=1.18075 NRD=39.996 NRS=38.568 M=1
+ R=2.8 SA=75003.4 SB=75001.8 A=0.063 P=1.14 MULT=1
MM1019 N_VGND_M1019_d N_A_1475_426#_M1019_g A_1449_133# VNB NSHORT L=0.15 W=0.42
+ AD=0.1155 AS=0.0819 PD=0.97 PS=0.81 NRD=38.568 NRS=39.996 M=1 R=2.8 SA=75003.9
+ SB=75001.3 A=0.063 P=1.14 MULT=1
MM1003 A_1697_133# N_RESET_B_M1003_g N_VGND_M1019_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1155 PD=0.63 PS=0.97 NRD=14.28 NRS=38.568 M=1 R=2.8 SA=75004.6
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1032 N_A_1475_426#_M1032_d N_A_1255_449#_M1032_g A_1697_133# VNB NSHORT L=0.15
+ W=0.42 AD=0.1197 AS=0.0441 PD=1.41 PS=0.63 NRD=5.712 NRS=14.28 M=1 R=2.8
+ SA=75005 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1035 N_VGND_M1035_d N_A_1255_449#_M1035_g N_A_1891_47#_M1035_s VNB NSHORT
+ L=0.15 W=0.84 AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6
+ SA=75000.2 SB=75001.9 A=0.126 P=1.98 MULT=1
MM1004 N_Q_M1004_d N_A_1891_47#_M1004_g N_VGND_M1035_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75000.6
+ SB=75001.5 A=0.126 P=1.98 MULT=1
MM1006 N_Q_M1004_d N_A_1891_47#_M1006_g N_VGND_M1006_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.1
+ SB=75001.1 A=0.126 P=1.98 MULT=1
MM1015 N_Q_M1015_d N_A_1891_47#_M1015_g N_VGND_M1006_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.1176 PD=1.12 PS=1.12 NRD=0 NRS=0 M=1 R=5.6 SA=75001.5
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1029 N_Q_M1015_d N_A_1891_47#_M1029_g N_VGND_M1029_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2226 PD=1.12 PS=2.21 NRD=0 NRS=0 M=1 R=5.6 SA=75001.9
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1036 N_VPWR_M1036_d N_CLK_M1036_g N_A_27_90#_M1036_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0896 AS=0.1696 PD=0.92 PS=1.81 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75000.6 A=0.096 P=1.58 MULT=1
MM1013 N_A_216_462#_M1013_d N_A_27_90#_M1013_g N_VPWR_M1036_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1696 AS=0.0896 PD=1.81 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.6 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1034 N_VPWR_M1034_d N_RESET_B_M1034_g N_A_340_535#_M1034_s VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.4 A=0.063 P=1.14 MULT=1
MM1023 N_A_340_535#_M1023_d N_D_M1023_g N_VPWR_M1034_d VPB PHIGHVT L=0.15 W=0.42
+ AD=0.0588 AS=0.0588 PD=0.7 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6 SB=75002
+ A=0.063 P=1.14 MULT=1
MM1009 N_A_595_535#_M1009_d N_A_216_462#_M1009_g N_A_340_535#_M1023_d VPB
+ PHIGHVT L=0.15 W=0.42 AD=0.0672 AS=0.0588 PD=0.74 PS=0.7 NRD=18.7544 NRS=0 M=1
+ R=2.8 SA=75001.1 SB=75001.5 A=0.063 P=1.14 MULT=1
MM1001 A_689_535# N_A_27_90#_M1001_g N_A_595_535#_M1009_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.0441 AS=0.0672 PD=0.63 PS=0.74 NRD=23.443 NRS=0 M=1 R=2.8
+ SA=75001.5 SB=75001.1 A=0.063 P=1.14 MULT=1
MM1000 N_VPWR_M1000_d N_A_731_405#_M1000_g A_689_535# VPB PHIGHVT L=0.15 W=0.42
+ AD=0.07455 AS=0.0441 PD=0.775 PS=0.63 NRD=35.1645 NRS=23.443 M=1 R=2.8
+ SA=75001.9 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1007 N_A_595_535#_M1007_d N_RESET_B_M1007_g N_VPWR_M1000_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.1113 AS=0.07455 PD=1.37 PS=0.775 NRD=0 NRS=0 M=1 R=2.8 SA=75002.4
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1027 N_A_731_405#_M1027_d N_A_595_535#_M1027_g N_VPWR_M1027_s VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.1176 AS=0.3679 PD=1.12 PS=2.7 NRD=0 NRS=28.1316 M=1 R=5.6
+ SA=75000.3 SB=75002 A=0.126 P=1.98 MULT=1
MM1014 N_A_1255_449#_M1014_d N_A_27_90#_M1014_g N_A_731_405#_M1027_d VPB PHIGHVT
+ L=0.15 W=0.84 AD=0.222633 AS=0.1176 PD=1.75333 PS=1.12 NRD=18.7544 NRS=0 M=1
+ R=5.6 SA=75000.8 SB=75001.5 A=0.126 P=1.98 MULT=1
MM1028 A_1380_488# N_A_216_462#_M1028_g N_A_1255_449#_M1014_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.09975 AS=0.111317 PD=0.895 PS=0.876667 NRD=85.5965 NRS=56.2829 M=1
+ R=2.8 SA=75001.4 SB=75002.2 A=0.063 P=1.14 MULT=1
MM1016 N_VPWR_M1016_d N_A_1475_426#_M1016_g A_1380_488# VPB PHIGHVT L=0.15
+ W=0.42 AD=0.15015 AS=0.09975 PD=1.135 PS=0.895 NRD=100.844 NRS=85.5965 M=1
+ R=2.8 SA=75002 SB=75001.6 A=0.063 P=1.14 MULT=1
MM1024 N_A_1475_426#_M1024_d N_RESET_B_M1024_g N_VPWR_M1016_d VPB PHIGHVT L=0.15
+ W=0.42 AD=0.06405 AS=0.15015 PD=0.725 PS=1.135 NRD=0 NRS=103.189 M=1 R=2.8
+ SA=75002.9 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1030 N_VPWR_M1030_d N_A_1255_449#_M1030_g N_A_1475_426#_M1024_d VPB PHIGHVT
+ L=0.15 W=0.42 AD=0.1428 AS=0.06405 PD=1.52 PS=0.725 NRD=25.7873 NRS=11.7215
+ M=1 R=2.8 SA=75003.3 SB=75000.3 A=0.063 P=1.14 MULT=1
MM1011 N_VPWR_M1011_d N_A_1255_449#_M1011_g N_A_1891_47#_M1011_s VPB PHIGHVT
+ L=0.15 W=1.26 AD=0.1764 AS=0.3339 PD=1.54 PS=3.05 NRD=0 NRS=0 M=1 R=8.4
+ SA=75000.2 SB=75001.9 A=0.189 P=2.82 MULT=1
MM1005 N_VPWR_M1011_d N_A_1891_47#_M1005_g N_Q_M1005_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75000.6
+ SB=75001.5 A=0.189 P=2.82 MULT=1
MM1017 N_VPWR_M1017_d N_A_1891_47#_M1017_g N_Q_M1005_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75001.1 A=0.189 P=2.82 MULT=1
MM1026 N_VPWR_M1017_d N_A_1891_47#_M1026_g N_Q_M1026_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.1764 PD=1.54 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.5
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1037 N_VPWR_M1037_d N_A_1891_47#_M1037_g N_Q_M1026_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3339 AS=0.1764 PD=3.05 PS=1.54 NRD=0 NRS=0 M=1 R=8.4 SA=75001.9
+ SB=75000.2 A=0.189 P=2.82 MULT=1
DX38_noxref VNB VPB NWDIODE A=23.0887 P=28.49
c_131 VNB 0 6.36774e-20 $X=0 $Y=0
*
.include "sky130_fd_sc_lp__dfrtp_4.pxi.spice"
*
.ends
*
*
