* NGSPICE file created from sky130_fd_sc_lp__and3_lp.ext - technology: sky130A

.subckt sky130_fd_sc_lp__and3_lp A B C VGND VNB VPB VPWR X
M1000 a_38_416# B VPWR VPB phighvt w=1e+06u l=250000u
+  ad=5.65e+11p pd=5.13e+06u as=6e+11p ps=5.2e+06u
M1001 VGND C a_234_47# VNB nshort w=420000u l=150000u
+  ad=1.533e+11p pd=1.57e+06u as=1.008e+11p ps=1.32e+06u
M1002 a_415_47# a_38_416# VGND VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1003 VPWR A a_38_416# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1004 X a_38_416# a_415_47# VNB nshort w=420000u l=150000u
+  ad=1.197e+11p pd=1.41e+06u as=0p ps=0u
M1005 X a_38_416# VPWR VPB phighvt w=1e+06u l=250000u
+  ad=2.85e+11p pd=2.57e+06u as=0p ps=0u
M1006 a_156_47# A a_38_416# VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=1.197e+11p ps=1.41e+06u
M1007 a_234_47# B a_156_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPWR C a_38_416# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
.ends

