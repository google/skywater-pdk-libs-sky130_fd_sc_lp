* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__sregrbp_1 ASYNC CLK D SCD SCE VGND VNB VPB VPWR Q Q_N
X0 a_1225_463# a_1273_393# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X1 a_1831_373# a_761_357# a_1903_125# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X2 a_342_531# SCE a_486_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 a_1825_125# a_934_357# a_1903_125# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X4 a_264_531# D a_342_531# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X5 VGND a_761_357# a_934_357# VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X6 Q a_2083_65# VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X7 a_75_531# SCE VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X8 VPWR a_342_531# a_636_531# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X9 VPWR a_1903_125# a_2083_65# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X10 a_761_357# CLK VGND VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X11 VGND a_2083_65# a_2456_451# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 VGND a_2456_451# Q_N VNB sky130_fd_pr__nfet_01v8 w=840000u l=150000u
X13 VGND a_75_531# a_312_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X14 VGND SCE a_75_531# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X15 VPWR a_1273_393# a_1831_373# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X16 a_761_357# CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X17 a_1139_463# a_761_357# a_1225_463# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X18 a_1501_119# ASYNC a_1273_393# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X19 a_1139_463# a_934_357# a_1319_119# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X20 a_2083_65# ASYNC VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X21 VPWR SCE a_264_531# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X22 VPWR a_2083_65# a_2456_451# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=150000u
X23 Q a_2083_65# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X24 a_2222_47# ASYNC a_2083_65# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X25 a_342_531# a_75_531# a_428_531# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X26 VPWR a_761_357# a_934_357# VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X27 a_486_47# SCD VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X28 a_636_531# a_934_357# a_1139_463# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X29 a_1903_125# a_934_357# a_2042_451# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X30 VGND a_342_531# a_636_531# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X31 a_2042_451# a_2083_65# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X32 VGND a_1139_463# a_1501_119# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X33 VGND a_1273_393# a_1825_125# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X34 a_1273_393# a_1139_463# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X35 a_1319_119# a_1273_393# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X36 VPWR a_2456_451# Q_N VPB sky130_fd_pr__pfet_01v8_hvt w=1.26e+06u l=150000u
X37 a_1903_125# a_761_357# a_2035_91# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X38 a_428_531# SCD VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X39 a_312_47# D a_342_531# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X40 a_636_531# a_761_357# a_1139_463# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X41 VGND a_1903_125# a_2222_47# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X42 VPWR ASYNC a_1273_393# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=150000u
X43 a_2035_91# a_2083_65# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
