* File: sky130_fd_sc_lp__dlrbp_1.pxi.spice
* Created: Wed Sep  2 09:46:29 2020
* 
x_PM_SKY130_FD_SC_LP__DLRBP_1%GATE N_GATE_M1004_g N_GATE_c_172_n N_GATE_M1011_g
+ N_GATE_c_173_n GATE GATE N_GATE_c_174_n N_GATE_c_175_n N_GATE_c_176_n
+ PM_SKY130_FD_SC_LP__DLRBP_1%GATE
x_PM_SKY130_FD_SC_LP__DLRBP_1%D N_D_c_204_n N_D_M1003_g N_D_M1017_g N_D_c_210_n
+ D D N_D_c_207_n PM_SKY130_FD_SC_LP__DLRBP_1%D
x_PM_SKY130_FD_SC_LP__DLRBP_1%A_373_481# N_A_373_481#_M1017_s
+ N_A_373_481#_M1003_s N_A_373_481#_c_252_n N_A_373_481#_c_253_n
+ N_A_373_481#_M1018_g N_A_373_481#_M1009_g N_A_373_481#_c_255_n
+ N_A_373_481#_c_256_n N_A_373_481#_c_257_n N_A_373_481#_c_258_n
+ N_A_373_481#_c_264_n N_A_373_481#_c_259_n N_A_373_481#_c_265_n
+ PM_SKY130_FD_SC_LP__DLRBP_1%A_373_481#
x_PM_SKY130_FD_SC_LP__DLRBP_1%A_218_483# N_A_218_483#_M1023_d
+ N_A_218_483#_M1020_d N_A_218_483#_M1015_g N_A_218_483#_M1001_g
+ N_A_218_483#_c_339_n N_A_218_483#_c_352_n N_A_218_483#_c_340_n
+ N_A_218_483#_c_341_n N_A_218_483#_c_332_n N_A_218_483#_c_393_p
+ N_A_218_483#_c_343_n N_A_218_483#_c_344_n N_A_218_483#_c_345_n
+ N_A_218_483#_c_346_n N_A_218_483#_c_347_n N_A_218_483#_c_333_n
+ N_A_218_483#_c_334_n N_A_218_483#_c_335_n N_A_218_483#_c_336_n
+ N_A_218_483#_c_398_p N_A_218_483#_c_337_n
+ PM_SKY130_FD_SC_LP__DLRBP_1%A_218_483#
x_PM_SKY130_FD_SC_LP__DLRBP_1%A_49_93# N_A_49_93#_M1004_s N_A_49_93#_M1011_s
+ N_A_49_93#_M1020_g N_A_49_93#_c_461_n N_A_49_93#_M1023_g N_A_49_93#_c_462_n
+ N_A_49_93#_c_463_n N_A_49_93#_c_464_n N_A_49_93#_c_465_n N_A_49_93#_c_466_n
+ N_A_49_93#_M1014_g N_A_49_93#_c_474_n N_A_49_93#_c_475_n N_A_49_93#_M1021_g
+ N_A_49_93#_c_468_n N_A_49_93#_c_469_n N_A_49_93#_c_478_n N_A_49_93#_c_479_n
+ N_A_49_93#_c_470_n N_A_49_93#_c_480_n N_A_49_93#_c_481_n
+ PM_SKY130_FD_SC_LP__DLRBP_1%A_49_93#
x_PM_SKY130_FD_SC_LP__DLRBP_1%A_776_93# N_A_776_93#_M1013_s N_A_776_93#_M1006_d
+ N_A_776_93#_M1019_g N_A_776_93#_M1010_g N_A_776_93#_M1007_g
+ N_A_776_93#_M1016_g N_A_776_93#_M1000_g N_A_776_93#_M1008_g
+ N_A_776_93#_c_577_n N_A_776_93#_c_593_n N_A_776_93#_c_578_n
+ N_A_776_93#_c_579_n N_A_776_93#_c_596_n N_A_776_93#_c_597_n
+ N_A_776_93#_c_598_n N_A_776_93#_c_580_n N_A_776_93#_c_581_n
+ N_A_776_93#_c_582_n N_A_776_93#_c_657_p N_A_776_93#_c_583_n
+ N_A_776_93#_c_599_n N_A_776_93#_c_600_n N_A_776_93#_c_584_n
+ N_A_776_93#_c_602_n N_A_776_93#_c_603_n N_A_776_93#_c_585_n
+ N_A_776_93#_c_586_n N_A_776_93#_c_606_n N_A_776_93#_c_587_n
+ N_A_776_93#_c_588_n N_A_776_93#_c_589_n PM_SKY130_FD_SC_LP__DLRBP_1%A_776_93#
x_PM_SKY130_FD_SC_LP__DLRBP_1%A_626_119# N_A_626_119#_M1015_d
+ N_A_626_119#_M1014_d N_A_626_119#_M1006_g N_A_626_119#_c_774_n
+ N_A_626_119#_M1013_g N_A_626_119#_c_775_n N_A_626_119#_c_776_n
+ N_A_626_119#_c_777_n N_A_626_119#_c_781_n N_A_626_119#_c_778_n
+ N_A_626_119#_c_779_n PM_SKY130_FD_SC_LP__DLRBP_1%A_626_119#
x_PM_SKY130_FD_SC_LP__DLRBP_1%RESET_B N_RESET_B_M1005_g N_RESET_B_M1022_g
+ RESET_B RESET_B RESET_B N_RESET_B_c_855_n PM_SKY130_FD_SC_LP__DLRBP_1%RESET_B
x_PM_SKY130_FD_SC_LP__DLRBP_1%A_1187_131# N_A_1187_131#_M1007_d
+ N_A_1187_131#_M1016_d N_A_1187_131#_c_899_n N_A_1187_131#_c_900_n
+ N_A_1187_131#_M1012_g N_A_1187_131#_M1002_g N_A_1187_131#_c_903_n
+ N_A_1187_131#_c_904_n N_A_1187_131#_c_905_n N_A_1187_131#_c_906_n
+ N_A_1187_131#_c_907_n N_A_1187_131#_c_911_n N_A_1187_131#_c_908_n
+ PM_SKY130_FD_SC_LP__DLRBP_1%A_1187_131#
x_PM_SKY130_FD_SC_LP__DLRBP_1%VPWR N_VPWR_M1011_d N_VPWR_M1003_d N_VPWR_M1010_d
+ N_VPWR_M1022_d N_VPWR_M1012_d N_VPWR_c_955_n N_VPWR_c_956_n N_VPWR_c_957_n
+ N_VPWR_c_958_n N_VPWR_c_959_n N_VPWR_c_960_n N_VPWR_c_961_n VPWR
+ N_VPWR_c_962_n N_VPWR_c_963_n N_VPWR_c_964_n N_VPWR_c_965_n N_VPWR_c_954_n
+ N_VPWR_c_967_n N_VPWR_c_968_n N_VPWR_c_969_n N_VPWR_c_970_n
+ PM_SKY130_FD_SC_LP__DLRBP_1%VPWR
x_PM_SKY130_FD_SC_LP__DLRBP_1%Q_N N_Q_N_M1002_s N_Q_N_M1012_s Q_N Q_N Q_N Q_N
+ Q_N N_Q_N_c_1055_n PM_SKY130_FD_SC_LP__DLRBP_1%Q_N
x_PM_SKY130_FD_SC_LP__DLRBP_1%Q N_Q_M1008_d N_Q_M1000_d Q Q Q Q Q Q Q
+ N_Q_c_1079_n Q N_Q_c_1082_n Q PM_SKY130_FD_SC_LP__DLRBP_1%Q
x_PM_SKY130_FD_SC_LP__DLRBP_1%VGND N_VGND_M1004_d N_VGND_M1017_d N_VGND_M1019_d
+ N_VGND_M1005_d N_VGND_M1002_d N_VGND_c_1102_n N_VGND_c_1103_n N_VGND_c_1104_n
+ N_VGND_c_1105_n N_VGND_c_1106_n N_VGND_c_1107_n N_VGND_c_1108_n
+ N_VGND_c_1109_n VGND N_VGND_c_1110_n N_VGND_c_1111_n N_VGND_c_1112_n
+ N_VGND_c_1113_n N_VGND_c_1114_n N_VGND_c_1115_n N_VGND_c_1116_n
+ N_VGND_c_1117_n PM_SKY130_FD_SC_LP__DLRBP_1%VGND
cc_1 VNB N_GATE_c_172_n 0.0234998f $X=-0.19 $Y=-0.245 $X2=0.697 $Y2=1.478
cc_2 VNB N_GATE_c_173_n 0.0141478f $X=-0.19 $Y=-0.245 $X2=0.697 $Y2=1.665
cc_3 VNB N_GATE_c_174_n 0.0213409f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.16
cc_4 VNB N_GATE_c_175_n 0.00385522f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.16
cc_5 VNB N_GATE_c_176_n 0.0221345f $X=-0.19 $Y=-0.245 $X2=0.697 $Y2=0.995
cc_6 VNB N_D_c_204_n 0.00248774f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=0.675
cc_7 VNB N_D_M1017_g 0.0343727f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB D 0.00261626f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_9 VNB N_D_c_207_n 0.0187553f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.16
cc_10 VNB N_A_373_481#_c_252_n 0.00509211f $X=-0.19 $Y=-0.245 $X2=0.585
+ $Y2=2.735
cc_11 VNB N_A_373_481#_c_253_n 0.0134868f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=2.735
cc_12 VNB N_A_373_481#_M1018_g 0.0227644f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_13 VNB N_A_373_481#_c_255_n 0.00786487f $X=-0.19 $Y=-0.245 $X2=0.755 $Y2=1.16
cc_14 VNB N_A_373_481#_c_256_n 0.00554549f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_373_481#_c_257_n 0.0155785f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_373_481#_c_258_n 0.00345831f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_373_481#_c_259_n 0.00865517f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_218_483#_c_332_n 0.00268914f $X=-0.19 $Y=-0.245 $X2=0.755
+ $Y2=1.665
cc_19 VNB N_A_218_483#_c_333_n 0.0123067f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_218_483#_c_334_n 0.00372986f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_218_483#_c_335_n 0.00256512f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_218_483#_c_336_n 0.0366218f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_218_483#_c_337_n 0.0157443f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_A_49_93#_c_461_n 0.0193257f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_25 VNB N_A_49_93#_c_462_n 0.0353911f $X=-0.19 $Y=-0.245 $X2=0.697 $Y2=1.16
cc_26 VNB N_A_49_93#_c_463_n 0.0373469f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.16
cc_27 VNB N_A_49_93#_c_464_n 0.046633f $X=-0.19 $Y=-0.245 $X2=0.755 $Y2=1.16
cc_28 VNB N_A_49_93#_c_465_n 0.134355f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_A_49_93#_c_466_n 0.0126197f $X=-0.19 $Y=-0.245 $X2=0.755 $Y2=1.295
cc_30 VNB N_A_49_93#_M1021_g 0.0534401f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_A_49_93#_c_468_n 0.00741257f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_A_49_93#_c_469_n 0.0411554f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A_49_93#_c_470_n 0.0126278f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_A_776_93#_M1019_g 0.0257191f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VNB N_A_776_93#_M1007_g 0.0279521f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.16
cc_36 VNB N_A_776_93#_M1000_g 0.00494362f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A_776_93#_c_577_n 0.0244318f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VNB N_A_776_93#_c_578_n 0.00307401f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_A_776_93#_c_579_n 0.0178921f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_40 VNB N_A_776_93#_c_580_n 0.00443849f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_41 VNB N_A_776_93#_c_581_n 0.00101471f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_42 VNB N_A_776_93#_c_582_n 0.00185848f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_A_776_93#_c_583_n 0.00230825f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_A_776_93#_c_584_n 0.00100943f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_45 VNB N_A_776_93#_c_585_n 0.00224927f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_46 VNB N_A_776_93#_c_586_n 0.0268271f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_A_776_93#_c_587_n 0.00385621f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_A_776_93#_c_588_n 0.0379359f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_A_776_93#_c_589_n 0.020022f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_A_626_119#_M1006_g 0.0049249f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_A_626_119#_c_774_n 0.0188221f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_52 VNB N_A_626_119#_c_775_n 0.00157741f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_A_626_119#_c_776_n 0.0225685f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.16
cc_54 VNB N_A_626_119#_c_777_n 0.0102123f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_A_626_119#_c_778_n 0.00335596f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_A_626_119#_c_779_n 0.0459632f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_RESET_B_M1005_g 0.0196181f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=0.675
cc_58 VNB N_RESET_B_M1022_g 0.00293979f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=2.735
cc_59 VNB RESET_B 0.00461394f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_RESET_B_c_855_n 0.0328172f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.16
cc_61 VNB N_A_1187_131#_c_899_n 0.0236385f $X=-0.19 $Y=-0.245 $X2=0.585
+ $Y2=2.735
cc_62 VNB N_A_1187_131#_c_900_n 0.0180948f $X=-0.19 $Y=-0.245 $X2=0.585
+ $Y2=2.735
cc_63 VNB N_A_1187_131#_M1012_g 0.0136814f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_64 VNB N_A_1187_131#_M1002_g 0.0220478f $X=-0.19 $Y=-0.245 $X2=0.697 $Y2=1.16
cc_65 VNB N_A_1187_131#_c_903_n 0.00705697f $X=-0.19 $Y=-0.245 $X2=0.697
+ $Y2=0.995
cc_66 VNB N_A_1187_131#_c_904_n 0.00217584f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_67 VNB N_A_1187_131#_c_905_n 0.002696f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_68 VNB N_A_1187_131#_c_906_n 0.00652769f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_69 VNB N_A_1187_131#_c_907_n 0.0477231f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_70 VNB N_A_1187_131#_c_908_n 0.00882696f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_71 VNB N_VPWR_c_954_n 0.342803f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_72 VNB N_Q_N_c_1055_n 0.0246772f $X=-0.19 $Y=-0.245 $X2=0.697 $Y2=0.995
cc_73 VNB Q 0.0107012f $X=-0.19 $Y=-0.245 $X2=0.585 $Y2=2.735
cc_74 VNB Q 0.0308583f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_75 VNB N_Q_c_1079_n 0.0290875f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_76 VNB N_VGND_c_1102_n 0.0160002f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_77 VNB N_VGND_c_1103_n 0.0128611f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_78 VNB N_VGND_c_1104_n 0.0402755f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_79 VNB N_VGND_c_1105_n 0.0154915f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_80 VNB N_VGND_c_1106_n 0.0122653f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_81 VNB N_VGND_c_1107_n 0.00595504f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_82 VNB N_VGND_c_1108_n 0.043765f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_83 VNB N_VGND_c_1109_n 0.00403597f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_84 VNB N_VGND_c_1110_n 0.0372553f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_85 VNB N_VGND_c_1111_n 0.0255258f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_86 VNB N_VGND_c_1112_n 0.0208004f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_87 VNB N_VGND_c_1113_n 0.460194f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_88 VNB N_VGND_c_1114_n 0.029373f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_89 VNB N_VGND_c_1115_n 0.00392849f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_90 VNB N_VGND_c_1116_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_91 VNB N_VGND_c_1117_n 0.00510247f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_92 VPB N_GATE_M1011_g 0.056898f $X=-0.19 $Y=1.655 $X2=0.585 $Y2=2.735
cc_93 VPB N_GATE_c_173_n 0.00719306f $X=-0.19 $Y=1.655 $X2=0.697 $Y2=1.665
cc_94 VPB N_GATE_c_175_n 0.00291679f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=1.16
cc_95 VPB N_D_c_204_n 0.0227006f $X=-0.19 $Y=1.655 $X2=0.585 $Y2=0.675
cc_96 VPB N_D_M1003_g 0.0325997f $X=-0.19 $Y=1.655 $X2=0.697 $Y2=1.478
cc_97 VPB N_D_c_210_n 0.0196248f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_98 VPB D 0.00650176f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_99 VPB N_A_373_481#_c_253_n 0.00256103f $X=-0.19 $Y=1.655 $X2=0.585 $Y2=2.735
cc_100 VPB N_A_373_481#_M1009_g 0.0324273f $X=-0.19 $Y=1.655 $X2=0.697 $Y2=1.16
cc_101 VPB N_A_373_481#_c_255_n 0.015095f $X=-0.19 $Y=1.655 $X2=0.755 $Y2=1.16
cc_102 VPB N_A_373_481#_c_258_n 0.00303419f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_103 VPB N_A_373_481#_c_264_n 0.041256f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_104 VPB N_A_373_481#_c_265_n 0.0111341f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_105 VPB N_A_218_483#_M1001_g 0.0208687f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_106 VPB N_A_218_483#_c_339_n 0.0153465f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=1.16
cc_107 VPB N_A_218_483#_c_340_n 0.00970277f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_108 VPB N_A_218_483#_c_341_n 0.00366666f $X=-0.19 $Y=1.655 $X2=0.755
+ $Y2=1.295
cc_109 VPB N_A_218_483#_c_332_n 0.00552658f $X=-0.19 $Y=1.655 $X2=0.755
+ $Y2=1.665
cc_110 VPB N_A_218_483#_c_343_n 0.00407236f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_111 VPB N_A_218_483#_c_344_n 0.00136519f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_112 VPB N_A_218_483#_c_345_n 0.0113124f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_113 VPB N_A_218_483#_c_346_n 0.0441554f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_114 VPB N_A_218_483#_c_347_n 0.0140384f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_115 VPB N_A_218_483#_c_333_n 0.0156969f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_116 VPB N_A_49_93#_M1020_g 0.0231185f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_117 VPB N_A_49_93#_c_462_n 0.0218528f $X=-0.19 $Y=1.655 $X2=0.697 $Y2=1.16
cc_118 VPB N_A_49_93#_M1014_g 0.0353901f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_119 VPB N_A_49_93#_c_474_n 0.0269317f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_120 VPB N_A_49_93#_c_475_n 0.00826968f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_121 VPB N_A_49_93#_M1021_g 0.00330743f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_122 VPB N_A_49_93#_c_469_n 0.013506f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_123 VPB N_A_49_93#_c_478_n 0.0357423f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_124 VPB N_A_49_93#_c_479_n 0.00837261f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_125 VPB N_A_49_93#_c_480_n 0.0167985f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_126 VPB N_A_49_93#_c_481_n 0.0435295f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_127 VPB N_A_776_93#_M1010_g 0.0514079f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_128 VPB N_A_776_93#_M1016_g 0.023979f $X=-0.19 $Y=1.655 $X2=0.755 $Y2=1.295
cc_129 VPB N_A_776_93#_M1000_g 0.0235615f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_130 VPB N_A_776_93#_c_593_n 0.0262037f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_131 VPB N_A_776_93#_c_578_n 9.67053e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_132 VPB N_A_776_93#_c_579_n 0.00906961f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_133 VPB N_A_776_93#_c_596_n 0.00427573f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_134 VPB N_A_776_93#_c_597_n 0.00536519f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_135 VPB N_A_776_93#_c_598_n 0.0035097f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_136 VPB N_A_776_93#_c_599_n 0.00138687f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_137 VPB N_A_776_93#_c_600_n 0.0308669f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_138 VPB N_A_776_93#_c_584_n 0.00109152f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_139 VPB N_A_776_93#_c_602_n 0.00512402f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_140 VPB N_A_776_93#_c_603_n 0.00190656f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_141 VPB N_A_776_93#_c_585_n 5.15864e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_142 VPB N_A_776_93#_c_586_n 0.00735055f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_143 VPB N_A_776_93#_c_606_n 0.00179023f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_144 VPB N_A_626_119#_M1006_g 0.0216056f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_145 VPB N_A_626_119#_c_781_n 0.00105702f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_146 VPB N_A_626_119#_c_778_n 0.0107066f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_147 VPB N_RESET_B_M1022_g 0.0209342f $X=-0.19 $Y=1.655 $X2=0.585 $Y2=2.735
cc_148 VPB RESET_B 0.001183f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_149 VPB N_A_1187_131#_M1012_g 0.024467f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_150 VPB N_A_1187_131#_c_905_n 0.00531925f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_151 VPB N_A_1187_131#_c_911_n 0.00809333f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_152 VPB N_VPWR_c_955_n 0.00598367f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_153 VPB N_VPWR_c_956_n 0.00363629f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_154 VPB N_VPWR_c_957_n 0.00620907f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_155 VPB N_VPWR_c_958_n 0.0200918f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_156 VPB N_VPWR_c_959_n 4.89148e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_157 VPB N_VPWR_c_960_n 0.0435739f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_158 VPB N_VPWR_c_961_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_159 VPB N_VPWR_c_962_n 0.0409653f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_160 VPB N_VPWR_c_963_n 0.0427131f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_161 VPB N_VPWR_c_964_n 0.0149962f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_162 VPB N_VPWR_c_965_n 0.0194284f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_163 VPB N_VPWR_c_954_n 0.103264f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_164 VPB N_VPWR_c_967_n 0.0250062f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_165 VPB N_VPWR_c_968_n 0.0041411f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_166 VPB N_VPWR_c_969_n 0.00574453f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_167 VPB N_VPWR_c_970_n 0.00548753f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_168 VPB N_Q_N_c_1055_n 0.00269723f $X=-0.19 $Y=1.655 $X2=0.697 $Y2=0.995
cc_169 VPB Q 0.00432237f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_170 VPB Q 0.0140922f $X=-0.19 $Y=1.655 $X2=0.697 $Y2=1.665
cc_171 VPB N_Q_c_1082_n 0.0541945f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_172 N_GATE_c_174_n N_A_218_483#_c_333_n 3.54279e-19 $X=0.72 $Y=1.16 $X2=0
+ $Y2=0
cc_173 N_GATE_c_175_n N_A_218_483#_c_333_n 0.0249989f $X=0.72 $Y=1.16 $X2=0
+ $Y2=0
cc_174 N_GATE_c_176_n N_A_49_93#_c_461_n 0.0137249f $X=0.697 $Y=0.995 $X2=0
+ $Y2=0
cc_175 N_GATE_c_172_n N_A_49_93#_c_462_n 0.0216505f $X=0.697 $Y=1.478 $X2=0
+ $Y2=0
cc_176 N_GATE_M1011_g N_A_49_93#_c_462_n 0.00722859f $X=0.585 $Y=2.735 $X2=0
+ $Y2=0
cc_177 N_GATE_c_175_n N_A_49_93#_c_462_n 9.77808e-19 $X=0.72 $Y=1.16 $X2=0 $Y2=0
cc_178 N_GATE_c_174_n N_A_49_93#_c_468_n 0.0216505f $X=0.72 $Y=1.16 $X2=0 $Y2=0
cc_179 N_GATE_c_175_n N_A_49_93#_c_468_n 0.00281184f $X=0.72 $Y=1.16 $X2=0 $Y2=0
cc_180 N_GATE_c_175_n N_A_49_93#_c_469_n 0.0577043f $X=0.72 $Y=1.16 $X2=0 $Y2=0
cc_181 N_GATE_c_176_n N_A_49_93#_c_469_n 0.0313868f $X=0.697 $Y=0.995 $X2=0
+ $Y2=0
cc_182 N_GATE_M1011_g N_A_49_93#_c_478_n 0.00739514f $X=0.585 $Y=2.735 $X2=0
+ $Y2=0
cc_183 N_GATE_M1011_g N_A_49_93#_c_479_n 0.0282665f $X=0.585 $Y=2.735 $X2=0
+ $Y2=0
cc_184 N_GATE_c_173_n N_A_49_93#_c_479_n 0.00130072f $X=0.697 $Y=1.665 $X2=0
+ $Y2=0
cc_185 N_GATE_c_175_n N_A_49_93#_c_479_n 0.0225274f $X=0.72 $Y=1.16 $X2=0 $Y2=0
cc_186 N_GATE_c_176_n N_A_49_93#_c_470_n 0.00477214f $X=0.697 $Y=0.995 $X2=0
+ $Y2=0
cc_187 N_GATE_M1011_g N_A_49_93#_c_481_n 0.0283632f $X=0.585 $Y=2.735 $X2=0
+ $Y2=0
cc_188 N_GATE_M1011_g N_VPWR_c_955_n 0.00270385f $X=0.585 $Y=2.735 $X2=0 $Y2=0
cc_189 N_GATE_M1011_g N_VPWR_c_954_n 0.011101f $X=0.585 $Y=2.735 $X2=0 $Y2=0
cc_190 N_GATE_M1011_g N_VPWR_c_967_n 0.00545548f $X=0.585 $Y=2.735 $X2=0 $Y2=0
cc_191 N_GATE_c_174_n N_VGND_c_1102_n 0.00131222f $X=0.72 $Y=1.16 $X2=0 $Y2=0
cc_192 N_GATE_c_175_n N_VGND_c_1102_n 0.0146389f $X=0.72 $Y=1.16 $X2=0 $Y2=0
cc_193 N_GATE_c_176_n N_VGND_c_1102_n 0.00595587f $X=0.697 $Y=0.995 $X2=0 $Y2=0
cc_194 N_GATE_c_176_n N_VGND_c_1113_n 0.00515964f $X=0.697 $Y=0.995 $X2=0 $Y2=0
cc_195 N_GATE_c_176_n N_VGND_c_1114_n 0.00489592f $X=0.697 $Y=0.995 $X2=0 $Y2=0
cc_196 N_D_M1017_g N_A_373_481#_c_252_n 0.0110668f $X=2.265 $Y=0.805 $X2=0 $Y2=0
cc_197 D N_A_373_481#_c_253_n 0.00342126f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_198 N_D_c_207_n N_A_373_481#_c_253_n 0.0110668f $X=2.16 $Y=1.615 $X2=0 $Y2=0
cc_199 N_D_M1017_g N_A_373_481#_M1018_g 0.022355f $X=2.265 $Y=0.805 $X2=0 $Y2=0
cc_200 N_D_M1003_g N_A_373_481#_M1009_g 0.015968f $X=2.205 $Y=2.725 $X2=0 $Y2=0
cc_201 N_D_c_210_n N_A_373_481#_M1009_g 0.0018587f $X=2.167 $Y=2.12 $X2=0 $Y2=0
cc_202 D N_A_373_481#_M1009_g 0.00161862f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_203 N_D_M1003_g N_A_373_481#_c_255_n 0.00726867f $X=2.205 $Y=2.725 $X2=0
+ $Y2=0
cc_204 N_D_M1017_g N_A_373_481#_c_255_n 0.00507751f $X=2.265 $Y=0.805 $X2=0
+ $Y2=0
cc_205 D N_A_373_481#_c_255_n 0.0496524f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_206 N_D_c_207_n N_A_373_481#_c_255_n 0.0078059f $X=2.16 $Y=1.615 $X2=0 $Y2=0
cc_207 N_D_M1017_g N_A_373_481#_c_256_n 0.00208306f $X=2.265 $Y=0.805 $X2=0
+ $Y2=0
cc_208 N_D_M1017_g N_A_373_481#_c_257_n 0.016229f $X=2.265 $Y=0.805 $X2=0 $Y2=0
cc_209 N_D_M1017_g N_A_373_481#_c_258_n 0.00210816f $X=2.265 $Y=0.805 $X2=0
+ $Y2=0
cc_210 D N_A_373_481#_c_258_n 0.0335023f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_211 N_D_c_207_n N_A_373_481#_c_258_n 7.3197e-19 $X=2.16 $Y=1.615 $X2=0 $Y2=0
cc_212 N_D_c_204_n N_A_373_481#_c_264_n 0.0110668f $X=2.167 $Y=1.948 $X2=0 $Y2=0
cc_213 N_D_M1017_g N_A_373_481#_c_259_n 7.54522e-19 $X=2.265 $Y=0.805 $X2=0
+ $Y2=0
cc_214 D N_A_373_481#_c_259_n 0.0217003f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_215 N_D_c_207_n N_A_373_481#_c_259_n 0.00382741f $X=2.16 $Y=1.615 $X2=0 $Y2=0
cc_216 N_D_M1003_g N_A_373_481#_c_265_n 4.28647e-19 $X=2.205 $Y=2.725 $X2=0
+ $Y2=0
cc_217 N_D_c_210_n N_A_373_481#_c_265_n 0.00296752f $X=2.167 $Y=2.12 $X2=0 $Y2=0
cc_218 D N_A_373_481#_c_265_n 0.00114639f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_219 N_D_M1003_g N_A_218_483#_c_339_n 0.0149062f $X=2.205 $Y=2.725 $X2=0 $Y2=0
cc_220 N_D_M1003_g N_A_218_483#_c_352_n 0.0151588f $X=2.205 $Y=2.725 $X2=0 $Y2=0
cc_221 N_D_M1003_g N_A_218_483#_c_341_n 0.00579424f $X=2.205 $Y=2.725 $X2=0
+ $Y2=0
cc_222 N_D_c_210_n N_A_218_483#_c_341_n 4.69216e-19 $X=2.167 $Y=2.12 $X2=0 $Y2=0
cc_223 D N_A_218_483#_c_341_n 0.00783181f $X=2.075 $Y=1.58 $X2=0 $Y2=0
cc_224 N_D_M1003_g N_A_218_483#_c_347_n 3.39781e-19 $X=2.205 $Y=2.725 $X2=0
+ $Y2=0
cc_225 N_D_M1003_g N_A_218_483#_c_333_n 0.00480968f $X=2.205 $Y=2.725 $X2=0
+ $Y2=0
cc_226 N_D_M1017_g N_A_218_483#_c_333_n 6.19452e-19 $X=2.265 $Y=0.805 $X2=0
+ $Y2=0
cc_227 N_D_c_207_n N_A_49_93#_c_462_n 0.00361558f $X=2.16 $Y=1.615 $X2=0 $Y2=0
cc_228 N_D_M1017_g N_A_49_93#_c_464_n 0.0148316f $X=2.265 $Y=0.805 $X2=0 $Y2=0
cc_229 N_D_M1017_g N_A_49_93#_c_465_n 0.0104164f $X=2.265 $Y=0.805 $X2=0 $Y2=0
cc_230 N_D_c_204_n N_A_49_93#_c_481_n 0.00361558f $X=2.167 $Y=1.948 $X2=0 $Y2=0
cc_231 N_D_M1003_g N_VPWR_c_956_n 0.00279348f $X=2.205 $Y=2.725 $X2=0 $Y2=0
cc_232 N_D_M1003_g N_VPWR_c_962_n 0.00325872f $X=2.205 $Y=2.725 $X2=0 $Y2=0
cc_233 N_D_M1003_g N_VPWR_c_954_n 0.00614507f $X=2.205 $Y=2.725 $X2=0 $Y2=0
cc_234 N_D_M1017_g N_VGND_c_1103_n 0.00362665f $X=2.265 $Y=0.805 $X2=0 $Y2=0
cc_235 N_D_M1017_g N_VGND_c_1113_n 9.39239e-19 $X=2.265 $Y=0.805 $X2=0 $Y2=0
cc_236 N_A_373_481#_M1003_s N_A_218_483#_c_339_n 0.00287043f $X=1.865 $Y=2.405
+ $X2=0 $Y2=0
cc_237 N_A_373_481#_M1009_g N_A_218_483#_c_339_n 4.02509e-19 $X=2.905 $Y=2.725
+ $X2=0 $Y2=0
cc_238 N_A_373_481#_c_265_n N_A_218_483#_c_339_n 0.0253978f $X=1.99 $Y=2.57
+ $X2=0 $Y2=0
cc_239 N_A_373_481#_M1009_g N_A_218_483#_c_352_n 0.00127739f $X=2.905 $Y=2.725
+ $X2=0 $Y2=0
cc_240 N_A_373_481#_M1009_g N_A_218_483#_c_340_n 0.018945f $X=2.905 $Y=2.725
+ $X2=0 $Y2=0
cc_241 N_A_373_481#_c_258_n N_A_218_483#_c_340_n 0.0141502f $X=2.755 $Y=1.86
+ $X2=0 $Y2=0
cc_242 N_A_373_481#_c_264_n N_A_218_483#_c_340_n 0.00152209f $X=2.755 $Y=1.86
+ $X2=0 $Y2=0
cc_243 N_A_373_481#_c_255_n N_A_218_483#_c_341_n 0.00431466f $X=1.81 $Y=2.385
+ $X2=0 $Y2=0
cc_244 N_A_373_481#_c_265_n N_A_218_483#_c_341_n 0.00389792f $X=1.99 $Y=2.57
+ $X2=0 $Y2=0
cc_245 N_A_373_481#_c_253_n N_A_218_483#_c_332_n 0.00139956f $X=2.68 $Y=1.695
+ $X2=0 $Y2=0
cc_246 N_A_373_481#_c_264_n N_A_218_483#_c_332_n 0.00934779f $X=2.755 $Y=1.86
+ $X2=0 $Y2=0
cc_247 N_A_373_481#_M1009_g N_A_218_483#_c_344_n 6.80202e-19 $X=2.905 $Y=2.725
+ $X2=0 $Y2=0
cc_248 N_A_373_481#_c_255_n N_A_218_483#_c_333_n 0.0800025f $X=1.81 $Y=2.385
+ $X2=0 $Y2=0
cc_249 N_A_373_481#_c_256_n N_A_218_483#_c_333_n 0.0117808f $X=2.05 $Y=0.805
+ $X2=0 $Y2=0
cc_250 N_A_373_481#_c_259_n N_A_218_483#_c_333_n 0.0151021f $X=2.18 $Y=1.182
+ $X2=0 $Y2=0
cc_251 N_A_373_481#_c_265_n N_A_218_483#_c_333_n 0.0289991f $X=1.99 $Y=2.57
+ $X2=0 $Y2=0
cc_252 N_A_373_481#_c_256_n N_A_218_483#_c_334_n 0.0102945f $X=2.05 $Y=0.805
+ $X2=0 $Y2=0
cc_253 N_A_373_481#_M1018_g N_A_218_483#_c_335_n 3.40638e-19 $X=2.695 $Y=0.805
+ $X2=0 $Y2=0
cc_254 N_A_373_481#_c_257_n N_A_218_483#_c_335_n 0.011936f $X=2.59 $Y=1.195
+ $X2=0 $Y2=0
cc_255 N_A_373_481#_c_258_n N_A_218_483#_c_335_n 0.0525967f $X=2.755 $Y=1.86
+ $X2=0 $Y2=0
cc_256 N_A_373_481#_c_252_n N_A_218_483#_c_336_n 0.0299647f $X=2.68 $Y=1.445
+ $X2=0 $Y2=0
cc_257 N_A_373_481#_c_258_n N_A_218_483#_c_336_n 0.00105102f $X=2.755 $Y=1.86
+ $X2=0 $Y2=0
cc_258 N_A_373_481#_M1018_g N_A_218_483#_c_337_n 0.0299647f $X=2.695 $Y=0.805
+ $X2=0 $Y2=0
cc_259 N_A_373_481#_c_257_n N_A_218_483#_c_337_n 0.00122821f $X=2.59 $Y=1.195
+ $X2=0 $Y2=0
cc_260 N_A_373_481#_c_255_n N_A_49_93#_M1020_g 2.35073e-19 $X=1.81 $Y=2.385
+ $X2=0 $Y2=0
cc_261 N_A_373_481#_c_265_n N_A_49_93#_M1020_g 3.49685e-19 $X=1.99 $Y=2.57 $X2=0
+ $Y2=0
cc_262 N_A_373_481#_c_255_n N_A_49_93#_c_463_n 6.79817e-19 $X=1.81 $Y=2.385
+ $X2=0 $Y2=0
cc_263 N_A_373_481#_c_259_n N_A_49_93#_c_463_n 0.010078f $X=2.18 $Y=1.182 $X2=0
+ $Y2=0
cc_264 N_A_373_481#_c_256_n N_A_49_93#_c_464_n 0.00519577f $X=2.05 $Y=0.805
+ $X2=0 $Y2=0
cc_265 N_A_373_481#_M1018_g N_A_49_93#_c_465_n 0.0103107f $X=2.695 $Y=0.805
+ $X2=0 $Y2=0
cc_266 N_A_373_481#_c_256_n N_A_49_93#_c_465_n 0.00422946f $X=2.05 $Y=0.805
+ $X2=0 $Y2=0
cc_267 N_A_373_481#_M1009_g N_A_49_93#_M1014_g 0.0391128f $X=2.905 $Y=2.725
+ $X2=0 $Y2=0
cc_268 N_A_373_481#_c_258_n N_A_49_93#_c_475_n 2.25523e-19 $X=2.755 $Y=1.86
+ $X2=0 $Y2=0
cc_269 N_A_373_481#_c_264_n N_A_49_93#_c_475_n 0.044938f $X=2.755 $Y=1.86 $X2=0
+ $Y2=0
cc_270 N_A_373_481#_c_257_n N_A_626_119#_c_775_n 5.94015e-19 $X=2.59 $Y=1.195
+ $X2=0 $Y2=0
cc_271 N_A_373_481#_M1009_g N_VPWR_c_956_n 0.00994744f $X=2.905 $Y=2.725 $X2=0
+ $Y2=0
cc_272 N_A_373_481#_M1009_g N_VPWR_c_963_n 0.00445056f $X=2.905 $Y=2.725 $X2=0
+ $Y2=0
cc_273 N_A_373_481#_M1009_g N_VPWR_c_954_n 0.0079903f $X=2.905 $Y=2.725 $X2=0
+ $Y2=0
cc_274 N_A_373_481#_M1018_g N_VGND_c_1103_n 0.00987797f $X=2.695 $Y=0.805 $X2=0
+ $Y2=0
cc_275 N_A_373_481#_c_257_n N_VGND_c_1103_n 0.0198434f $X=2.59 $Y=1.195 $X2=0
+ $Y2=0
cc_276 N_A_373_481#_c_256_n N_VGND_c_1110_n 0.0050474f $X=2.05 $Y=0.805 $X2=0
+ $Y2=0
cc_277 N_A_373_481#_M1018_g N_VGND_c_1113_n 7.88961e-19 $X=2.695 $Y=0.805 $X2=0
+ $Y2=0
cc_278 N_A_373_481#_c_256_n N_VGND_c_1113_n 0.00753675f $X=2.05 $Y=0.805 $X2=0
+ $Y2=0
cc_279 N_A_218_483#_c_347_n N_A_49_93#_M1020_g 0.00748291f $X=1.23 $Y=2.56 $X2=0
+ $Y2=0
cc_280 N_A_218_483#_c_333_n N_A_49_93#_M1020_g 0.00361785f $X=1.305 $Y=2.425
+ $X2=0 $Y2=0
cc_281 N_A_218_483#_c_333_n N_A_49_93#_c_461_n 0.00247195f $X=1.305 $Y=2.425
+ $X2=0 $Y2=0
cc_282 N_A_218_483#_c_334_n N_A_49_93#_c_461_n 0.00504886f $X=1.385 $Y=0.675
+ $X2=0 $Y2=0
cc_283 N_A_218_483#_c_333_n N_A_49_93#_c_462_n 0.0264617f $X=1.305 $Y=2.425
+ $X2=0 $Y2=0
cc_284 N_A_218_483#_c_333_n N_A_49_93#_c_463_n 0.0150938f $X=1.305 $Y=2.425
+ $X2=0 $Y2=0
cc_285 N_A_218_483#_c_333_n N_A_49_93#_c_464_n 0.00153497f $X=1.305 $Y=2.425
+ $X2=0 $Y2=0
cc_286 N_A_218_483#_c_334_n N_A_49_93#_c_464_n 0.00540352f $X=1.385 $Y=0.675
+ $X2=0 $Y2=0
cc_287 N_A_218_483#_c_337_n N_A_49_93#_c_465_n 0.0104164f $X=3.145 $Y=1.125
+ $X2=0 $Y2=0
cc_288 N_A_218_483#_c_332_n N_A_49_93#_M1014_g 0.00646739f $X=3.11 $Y=2.29 $X2=0
+ $Y2=0
cc_289 N_A_218_483#_c_393_p N_A_49_93#_M1014_g 0.00800767f $X=3.11 $Y=2.905
+ $X2=0 $Y2=0
cc_290 N_A_218_483#_c_343_n N_A_49_93#_M1014_g 0.0121718f $X=3.755 $Y=2.99 $X2=0
+ $Y2=0
cc_291 N_A_218_483#_c_344_n N_A_49_93#_M1014_g 0.00110234f $X=3.195 $Y=2.99
+ $X2=0 $Y2=0
cc_292 N_A_218_483#_c_345_n N_A_49_93#_M1014_g 6.88433e-19 $X=3.93 $Y=2.3 $X2=0
+ $Y2=0
cc_293 N_A_218_483#_c_346_n N_A_49_93#_M1014_g 0.023789f $X=3.93 $Y=2.3 $X2=0
+ $Y2=0
cc_294 N_A_218_483#_c_398_p N_A_49_93#_M1014_g 0.00316831f $X=3.11 $Y=2.375
+ $X2=0 $Y2=0
cc_295 N_A_218_483#_c_332_n N_A_49_93#_c_475_n 0.00350633f $X=3.11 $Y=2.29 $X2=0
+ $Y2=0
cc_296 N_A_218_483#_c_335_n N_A_49_93#_c_475_n 3.63297e-19 $X=3.145 $Y=1.29
+ $X2=0 $Y2=0
cc_297 N_A_218_483#_c_336_n N_A_49_93#_c_475_n 0.0063097f $X=3.145 $Y=1.29 $X2=0
+ $Y2=0
cc_298 N_A_218_483#_c_332_n N_A_49_93#_M1021_g 0.00106545f $X=3.11 $Y=2.29 $X2=0
+ $Y2=0
cc_299 N_A_218_483#_c_335_n N_A_49_93#_M1021_g 3.08823e-19 $X=3.145 $Y=1.29
+ $X2=0 $Y2=0
cc_300 N_A_218_483#_c_336_n N_A_49_93#_M1021_g 0.0203656f $X=3.145 $Y=1.29 $X2=0
+ $Y2=0
cc_301 N_A_218_483#_c_337_n N_A_49_93#_M1021_g 0.00866639f $X=3.145 $Y=1.125
+ $X2=0 $Y2=0
cc_302 N_A_218_483#_c_334_n N_A_49_93#_c_468_n 0.0016786f $X=1.385 $Y=0.675
+ $X2=0 $Y2=0
cc_303 N_A_218_483#_c_347_n N_A_49_93#_c_479_n 0.00878828f $X=1.23 $Y=2.56 $X2=0
+ $Y2=0
cc_304 N_A_218_483#_c_333_n N_A_49_93#_c_479_n 0.0262086f $X=1.305 $Y=2.425
+ $X2=0 $Y2=0
cc_305 N_A_218_483#_c_347_n N_A_49_93#_c_481_n 0.0103484f $X=1.23 $Y=2.56 $X2=0
+ $Y2=0
cc_306 N_A_218_483#_M1001_g N_A_776_93#_M1010_g 0.0162912f $X=3.79 $Y=2.835
+ $X2=0 $Y2=0
cc_307 N_A_218_483#_c_343_n N_A_776_93#_M1010_g 0.00176785f $X=3.755 $Y=2.99
+ $X2=0 $Y2=0
cc_308 N_A_218_483#_c_345_n N_A_776_93#_M1010_g 0.0062326f $X=3.93 $Y=2.3 $X2=0
+ $Y2=0
cc_309 N_A_218_483#_c_346_n N_A_776_93#_M1010_g 0.0205444f $X=3.93 $Y=2.3 $X2=0
+ $Y2=0
cc_310 N_A_218_483#_c_346_n N_A_776_93#_c_593_n 0.00701312f $X=3.93 $Y=2.3 $X2=0
+ $Y2=0
cc_311 N_A_218_483#_c_345_n N_A_776_93#_c_596_n 0.0121399f $X=3.93 $Y=2.3 $X2=0
+ $Y2=0
cc_312 N_A_218_483#_c_346_n N_A_776_93#_c_596_n 0.00104016f $X=3.93 $Y=2.3 $X2=0
+ $Y2=0
cc_313 N_A_218_483#_c_345_n N_A_776_93#_c_598_n 0.0141251f $X=3.93 $Y=2.3 $X2=0
+ $Y2=0
cc_314 N_A_218_483#_c_346_n N_A_776_93#_c_598_n 0.00120976f $X=3.93 $Y=2.3 $X2=0
+ $Y2=0
cc_315 N_A_218_483#_c_345_n N_A_776_93#_c_602_n 0.00197651f $X=3.93 $Y=2.3 $X2=0
+ $Y2=0
cc_316 N_A_218_483#_c_346_n N_A_776_93#_c_602_n 6.09533e-19 $X=3.93 $Y=2.3 $X2=0
+ $Y2=0
cc_317 N_A_218_483#_c_343_n N_A_626_119#_M1014_d 0.00492676f $X=3.755 $Y=2.99
+ $X2=0 $Y2=0
cc_318 N_A_218_483#_c_335_n N_A_626_119#_c_775_n 0.00891911f $X=3.145 $Y=1.29
+ $X2=0 $Y2=0
cc_319 N_A_218_483#_c_336_n N_A_626_119#_c_775_n 0.00349704f $X=3.145 $Y=1.29
+ $X2=0 $Y2=0
cc_320 N_A_218_483#_c_337_n N_A_626_119#_c_775_n 0.00364822f $X=3.145 $Y=1.125
+ $X2=0 $Y2=0
cc_321 N_A_218_483#_M1001_g N_A_626_119#_c_781_n 0.00231621f $X=3.79 $Y=2.835
+ $X2=0 $Y2=0
cc_322 N_A_218_483#_c_343_n N_A_626_119#_c_781_n 0.0141662f $X=3.755 $Y=2.99
+ $X2=0 $Y2=0
cc_323 N_A_218_483#_c_398_p N_A_626_119#_c_781_n 0.00390582f $X=3.11 $Y=2.375
+ $X2=0 $Y2=0
cc_324 N_A_218_483#_c_332_n N_A_626_119#_c_778_n 0.0497139f $X=3.11 $Y=2.29
+ $X2=0 $Y2=0
cc_325 N_A_218_483#_c_345_n N_A_626_119#_c_778_n 0.0442782f $X=3.93 $Y=2.3 $X2=0
+ $Y2=0
cc_326 N_A_218_483#_c_346_n N_A_626_119#_c_778_n 0.00231621f $X=3.93 $Y=2.3
+ $X2=0 $Y2=0
cc_327 N_A_218_483#_c_335_n N_A_626_119#_c_778_n 0.0211001f $X=3.145 $Y=1.29
+ $X2=0 $Y2=0
cc_328 N_A_218_483#_c_336_n N_A_626_119#_c_778_n 0.00174112f $X=3.145 $Y=1.29
+ $X2=0 $Y2=0
cc_329 N_A_218_483#_c_398_p N_A_626_119#_c_778_n 0.00621363f $X=3.11 $Y=2.375
+ $X2=0 $Y2=0
cc_330 N_A_218_483#_c_339_n N_VPWR_M1003_d 0.00133555f $X=2.255 $Y=2.99 $X2=0
+ $Y2=0
cc_331 N_A_218_483#_c_352_n N_VPWR_M1003_d 0.00502614f $X=2.34 $Y=2.905 $X2=0
+ $Y2=0
cc_332 N_A_218_483#_c_340_n N_VPWR_M1003_d 0.00893588f $X=3.025 $Y=2.375 $X2=0
+ $Y2=0
cc_333 N_A_218_483#_c_347_n N_VPWR_c_955_n 0.026574f $X=1.23 $Y=2.56 $X2=0 $Y2=0
cc_334 N_A_218_483#_c_339_n N_VPWR_c_956_n 0.0143348f $X=2.255 $Y=2.99 $X2=0
+ $Y2=0
cc_335 N_A_218_483#_c_352_n N_VPWR_c_956_n 0.0205938f $X=2.34 $Y=2.905 $X2=0
+ $Y2=0
cc_336 N_A_218_483#_c_340_n N_VPWR_c_956_n 0.0161865f $X=3.025 $Y=2.375 $X2=0
+ $Y2=0
cc_337 N_A_218_483#_c_344_n N_VPWR_c_956_n 0.00753116f $X=3.195 $Y=2.99 $X2=0
+ $Y2=0
cc_338 N_A_218_483#_c_343_n N_VPWR_c_957_n 0.00643368f $X=3.755 $Y=2.99 $X2=0
+ $Y2=0
cc_339 N_A_218_483#_c_345_n N_VPWR_c_957_n 0.00913572f $X=3.93 $Y=2.3 $X2=0
+ $Y2=0
cc_340 N_A_218_483#_c_339_n N_VPWR_c_962_n 0.0574458f $X=2.255 $Y=2.99 $X2=0
+ $Y2=0
cc_341 N_A_218_483#_c_347_n N_VPWR_c_962_n 0.0341068f $X=1.23 $Y=2.56 $X2=0
+ $Y2=0
cc_342 N_A_218_483#_M1001_g N_VPWR_c_963_n 0.00325768f $X=3.79 $Y=2.835 $X2=0
+ $Y2=0
cc_343 N_A_218_483#_c_343_n N_VPWR_c_963_n 0.0537025f $X=3.755 $Y=2.99 $X2=0
+ $Y2=0
cc_344 N_A_218_483#_c_344_n N_VPWR_c_963_n 0.0121003f $X=3.195 $Y=2.99 $X2=0
+ $Y2=0
cc_345 N_A_218_483#_M1001_g N_VPWR_c_954_n 0.00528417f $X=3.79 $Y=2.835 $X2=0
+ $Y2=0
cc_346 N_A_218_483#_c_339_n N_VPWR_c_954_n 0.032617f $X=2.255 $Y=2.99 $X2=0
+ $Y2=0
cc_347 N_A_218_483#_c_343_n N_VPWR_c_954_n 0.0298062f $X=3.755 $Y=2.99 $X2=0
+ $Y2=0
cc_348 N_A_218_483#_c_344_n N_VPWR_c_954_n 0.00657636f $X=3.195 $Y=2.99 $X2=0
+ $Y2=0
cc_349 N_A_218_483#_c_346_n N_VPWR_c_954_n 0.0017992f $X=3.93 $Y=2.3 $X2=0 $Y2=0
cc_350 N_A_218_483#_c_347_n N_VPWR_c_954_n 0.0184595f $X=1.23 $Y=2.56 $X2=0
+ $Y2=0
cc_351 N_A_218_483#_c_343_n A_773_525# 0.00204994f $X=3.755 $Y=2.99 $X2=-0.19
+ $Y2=-0.245
cc_352 N_A_218_483#_c_345_n A_773_525# 0.00394633f $X=3.93 $Y=2.3 $X2=-0.19
+ $Y2=-0.245
cc_353 N_A_218_483#_c_337_n N_VGND_c_1103_n 0.00171025f $X=3.145 $Y=1.125 $X2=0
+ $Y2=0
cc_354 N_A_218_483#_c_334_n N_VGND_c_1110_n 0.00769038f $X=1.385 $Y=0.675 $X2=0
+ $Y2=0
cc_355 N_A_218_483#_c_334_n N_VGND_c_1113_n 0.0107127f $X=1.385 $Y=0.675 $X2=0
+ $Y2=0
cc_356 N_A_218_483#_c_337_n N_VGND_c_1113_n 9.39239e-19 $X=3.145 $Y=1.125 $X2=0
+ $Y2=0
cc_357 N_A_49_93#_M1021_g N_A_776_93#_M1019_g 0.0573542f $X=3.595 $Y=0.805 $X2=0
+ $Y2=0
cc_358 N_A_49_93#_M1014_g N_A_776_93#_c_593_n 3.44006e-19 $X=3.265 $Y=2.725
+ $X2=0 $Y2=0
cc_359 N_A_49_93#_c_474_n N_A_776_93#_c_593_n 0.00925517f $X=3.52 $Y=1.82 $X2=0
+ $Y2=0
cc_360 N_A_49_93#_M1021_g N_A_776_93#_c_578_n 0.00109724f $X=3.595 $Y=0.805
+ $X2=0 $Y2=0
cc_361 N_A_49_93#_M1021_g N_A_776_93#_c_579_n 0.00925517f $X=3.595 $Y=0.805
+ $X2=0 $Y2=0
cc_362 N_A_49_93#_c_474_n N_A_776_93#_c_602_n 0.00109724f $X=3.52 $Y=1.82 $X2=0
+ $Y2=0
cc_363 N_A_49_93#_c_465_n N_A_626_119#_c_775_n 0.00485162f $X=3.52 $Y=0.18 $X2=0
+ $Y2=0
cc_364 N_A_49_93#_M1021_g N_A_626_119#_c_775_n 0.0106873f $X=3.595 $Y=0.805
+ $X2=0 $Y2=0
cc_365 N_A_49_93#_M1021_g N_A_626_119#_c_776_n 0.0102642f $X=3.595 $Y=0.805
+ $X2=0 $Y2=0
cc_366 N_A_49_93#_c_474_n N_A_626_119#_c_781_n 0.00131103f $X=3.52 $Y=1.82 $X2=0
+ $Y2=0
cc_367 N_A_49_93#_M1014_g N_A_626_119#_c_778_n 0.00711312f $X=3.265 $Y=2.725
+ $X2=0 $Y2=0
cc_368 N_A_49_93#_c_474_n N_A_626_119#_c_778_n 0.0129501f $X=3.52 $Y=1.82 $X2=0
+ $Y2=0
cc_369 N_A_49_93#_M1021_g N_A_626_119#_c_778_n 0.0151649f $X=3.595 $Y=0.805
+ $X2=0 $Y2=0
cc_370 N_A_49_93#_M1020_g N_VPWR_c_955_n 0.00253142f $X=1.015 $Y=2.735 $X2=0
+ $Y2=0
cc_371 N_A_49_93#_c_478_n N_VPWR_c_955_n 0.0015231f $X=0.37 $Y=2.56 $X2=0 $Y2=0
cc_372 N_A_49_93#_c_479_n N_VPWR_c_955_n 0.0167738f $X=1.105 $Y=2.09 $X2=0 $Y2=0
cc_373 N_A_49_93#_M1014_g N_VPWR_c_956_n 0.00114059f $X=3.265 $Y=2.725 $X2=0
+ $Y2=0
cc_374 N_A_49_93#_M1020_g N_VPWR_c_962_n 0.00511358f $X=1.015 $Y=2.735 $X2=0
+ $Y2=0
cc_375 N_A_49_93#_M1014_g N_VPWR_c_963_n 0.00325896f $X=3.265 $Y=2.725 $X2=0
+ $Y2=0
cc_376 N_A_49_93#_M1020_g N_VPWR_c_954_n 0.0105214f $X=1.015 $Y=2.735 $X2=0
+ $Y2=0
cc_377 N_A_49_93#_M1014_g N_VPWR_c_954_n 0.00492529f $X=3.265 $Y=2.725 $X2=0
+ $Y2=0
cc_378 N_A_49_93#_c_478_n N_VPWR_c_954_n 0.0113912f $X=0.37 $Y=2.56 $X2=0 $Y2=0
cc_379 N_A_49_93#_c_478_n N_VPWR_c_967_n 0.0210042f $X=0.37 $Y=2.56 $X2=0 $Y2=0
cc_380 N_A_49_93#_c_461_n N_VGND_c_1102_n 0.00600242f $X=1.17 $Y=0.995 $X2=0
+ $Y2=0
cc_381 N_A_49_93#_c_466_n N_VGND_c_1102_n 0.00429842f $X=1.85 $Y=0.18 $X2=0
+ $Y2=0
cc_382 N_A_49_93#_c_464_n N_VGND_c_1103_n 0.00580625f $X=1.775 $Y=0.995 $X2=0
+ $Y2=0
cc_383 N_A_49_93#_c_465_n N_VGND_c_1103_n 0.0236334f $X=3.52 $Y=0.18 $X2=0 $Y2=0
cc_384 N_A_49_93#_c_465_n N_VGND_c_1104_n 0.0324909f $X=3.52 $Y=0.18 $X2=0 $Y2=0
cc_385 N_A_49_93#_c_465_n N_VGND_c_1105_n 0.0106942f $X=3.52 $Y=0.18 $X2=0 $Y2=0
cc_386 N_A_49_93#_M1021_g N_VGND_c_1105_n 0.00135753f $X=3.595 $Y=0.805 $X2=0
+ $Y2=0
cc_387 N_A_49_93#_c_461_n N_VGND_c_1110_n 0.00489592f $X=1.17 $Y=0.995 $X2=0
+ $Y2=0
cc_388 N_A_49_93#_c_466_n N_VGND_c_1110_n 0.0206801f $X=1.85 $Y=0.18 $X2=0 $Y2=0
cc_389 N_A_49_93#_c_461_n N_VGND_c_1113_n 0.00515964f $X=1.17 $Y=0.995 $X2=0
+ $Y2=0
cc_390 N_A_49_93#_c_465_n N_VGND_c_1113_n 0.0569965f $X=3.52 $Y=0.18 $X2=0 $Y2=0
cc_391 N_A_49_93#_c_466_n N_VGND_c_1113_n 0.0116041f $X=1.85 $Y=0.18 $X2=0 $Y2=0
cc_392 N_A_49_93#_c_470_n N_VGND_c_1113_n 0.0107802f $X=0.37 $Y=0.675 $X2=0
+ $Y2=0
cc_393 N_A_49_93#_c_470_n N_VGND_c_1114_n 0.00777897f $X=0.37 $Y=0.675 $X2=0
+ $Y2=0
cc_394 N_A_776_93#_c_593_n N_A_626_119#_M1006_g 0.0358966f $X=4.22 $Y=1.925
+ $X2=0 $Y2=0
cc_395 N_A_776_93#_c_578_n N_A_626_119#_M1006_g 0.00202605f $X=4.15 $Y=1.42
+ $X2=0 $Y2=0
cc_396 N_A_776_93#_c_579_n N_A_626_119#_M1006_g 0.0046757f $X=4.15 $Y=1.42 $X2=0
+ $Y2=0
cc_397 N_A_776_93#_c_597_n N_A_626_119#_M1006_g 0.0140545f $X=4.995 $Y=2.385
+ $X2=0 $Y2=0
cc_398 N_A_776_93#_c_602_n N_A_626_119#_M1006_g 0.0019912f $X=4.17 $Y=1.925
+ $X2=0 $Y2=0
cc_399 N_A_776_93#_c_603_n N_A_626_119#_M1006_g 2.96668e-19 $X=5.12 $Y=2.465
+ $X2=0 $Y2=0
cc_400 N_A_776_93#_c_580_n N_A_626_119#_c_774_n 0.00678038f $X=4.71 $Y=0.38
+ $X2=0 $Y2=0
cc_401 N_A_776_93#_c_581_n N_A_626_119#_c_774_n 0.0106239f $X=5.64 $Y=0.74 $X2=0
+ $Y2=0
cc_402 N_A_776_93#_c_582_n N_A_626_119#_c_774_n 0.00155434f $X=4.875 $Y=0.74
+ $X2=0 $Y2=0
cc_403 N_A_776_93#_M1019_g N_A_626_119#_c_775_n 0.00148033f $X=3.955 $Y=0.805
+ $X2=0 $Y2=0
cc_404 N_A_776_93#_M1013_s N_A_626_119#_c_776_n 0.00316686f $X=4.585 $Y=0.235
+ $X2=0 $Y2=0
cc_405 N_A_776_93#_M1019_g N_A_626_119#_c_776_n 0.0182838f $X=3.955 $Y=0.805
+ $X2=0 $Y2=0
cc_406 N_A_776_93#_c_577_n N_A_626_119#_c_776_n 0.00812738f $X=4.097 $Y=1.405
+ $X2=0 $Y2=0
cc_407 N_A_776_93#_c_593_n N_A_626_119#_c_776_n 0.00276736f $X=4.22 $Y=1.925
+ $X2=0 $Y2=0
cc_408 N_A_776_93#_c_578_n N_A_626_119#_c_776_n 0.0292404f $X=4.15 $Y=1.42 $X2=0
+ $Y2=0
cc_409 N_A_776_93#_c_582_n N_A_626_119#_c_776_n 0.0202029f $X=4.875 $Y=0.74
+ $X2=0 $Y2=0
cc_410 N_A_776_93#_M1019_g N_A_626_119#_c_777_n 8.7052e-19 $X=3.955 $Y=0.805
+ $X2=0 $Y2=0
cc_411 N_A_776_93#_c_577_n N_A_626_119#_c_777_n 7.95438e-19 $X=4.097 $Y=1.405
+ $X2=0 $Y2=0
cc_412 N_A_776_93#_c_578_n N_A_626_119#_c_777_n 0.0140945f $X=4.15 $Y=1.42 $X2=0
+ $Y2=0
cc_413 N_A_776_93#_M1019_g N_A_626_119#_c_778_n 0.00121707f $X=3.955 $Y=0.805
+ $X2=0 $Y2=0
cc_414 N_A_776_93#_c_593_n N_A_626_119#_c_778_n 2.67632e-19 $X=4.22 $Y=1.925
+ $X2=0 $Y2=0
cc_415 N_A_776_93#_c_578_n N_A_626_119#_c_778_n 0.0213791f $X=4.15 $Y=1.42 $X2=0
+ $Y2=0
cc_416 N_A_776_93#_c_579_n N_A_626_119#_c_778_n 0.00175649f $X=4.15 $Y=1.42
+ $X2=0 $Y2=0
cc_417 N_A_776_93#_c_596_n N_A_626_119#_c_778_n 0.00656462f $X=4.27 $Y=2.3 $X2=0
+ $Y2=0
cc_418 N_A_776_93#_M1019_g N_A_626_119#_c_779_n 0.001918f $X=3.955 $Y=0.805
+ $X2=0 $Y2=0
cc_419 N_A_776_93#_c_577_n N_A_626_119#_c_779_n 0.017178f $X=4.097 $Y=1.405
+ $X2=0 $Y2=0
cc_420 N_A_776_93#_c_578_n N_A_626_119#_c_779_n 0.00106867f $X=4.15 $Y=1.42
+ $X2=0 $Y2=0
cc_421 N_A_776_93#_c_582_n N_A_626_119#_c_779_n 0.00280183f $X=4.875 $Y=0.74
+ $X2=0 $Y2=0
cc_422 N_A_776_93#_M1007_g N_RESET_B_M1005_g 0.0164397f $X=5.86 $Y=0.865 $X2=0
+ $Y2=0
cc_423 N_A_776_93#_c_580_n N_RESET_B_M1005_g 0.00147554f $X=4.71 $Y=0.38 $X2=0
+ $Y2=0
cc_424 N_A_776_93#_c_581_n N_RESET_B_M1005_g 0.0130157f $X=5.64 $Y=0.74 $X2=0
+ $Y2=0
cc_425 N_A_776_93#_c_583_n N_RESET_B_M1005_g 0.0074215f $X=5.725 $Y=1.295 $X2=0
+ $Y2=0
cc_426 N_A_776_93#_M1016_g N_RESET_B_M1022_g 0.0279766f $X=5.86 $Y=2.105 $X2=0
+ $Y2=0
cc_427 N_A_776_93#_c_657_p N_RESET_B_M1022_g 0.0110108f $X=5.64 $Y=2.397 $X2=0
+ $Y2=0
cc_428 N_A_776_93#_c_599_n N_RESET_B_M1022_g 0.00506569f $X=5.725 $Y=2.3 $X2=0
+ $Y2=0
cc_429 N_A_776_93#_c_603_n N_RESET_B_M1022_g 2.785e-19 $X=5.12 $Y=2.465 $X2=0
+ $Y2=0
cc_430 N_A_776_93#_c_585_n N_RESET_B_M1022_g 2.8049e-19 $X=5.945 $Y=1.46 $X2=0
+ $Y2=0
cc_431 N_A_776_93#_c_586_n N_RESET_B_M1022_g 0.00263776f $X=5.945 $Y=1.46 $X2=0
+ $Y2=0
cc_432 N_A_776_93#_M1006_d RESET_B 0.00188202f $X=4.98 $Y=1.785 $X2=0 $Y2=0
cc_433 N_A_776_93#_M1016_g RESET_B 0.00144053f $X=5.86 $Y=2.105 $X2=0 $Y2=0
cc_434 N_A_776_93#_c_593_n RESET_B 0.00118063f $X=4.22 $Y=1.925 $X2=0 $Y2=0
cc_435 N_A_776_93#_c_578_n RESET_B 0.0177179f $X=4.15 $Y=1.42 $X2=0 $Y2=0
cc_436 N_A_776_93#_c_579_n RESET_B 2.77126e-19 $X=4.15 $Y=1.42 $X2=0 $Y2=0
cc_437 N_A_776_93#_c_597_n RESET_B 0.00244073f $X=4.995 $Y=2.385 $X2=0 $Y2=0
cc_438 N_A_776_93#_c_581_n RESET_B 0.0189102f $X=5.64 $Y=0.74 $X2=0 $Y2=0
cc_439 N_A_776_93#_c_657_p RESET_B 0.0109822f $X=5.64 $Y=2.397 $X2=0 $Y2=0
cc_440 N_A_776_93#_c_583_n RESET_B 0.00662241f $X=5.725 $Y=1.295 $X2=0 $Y2=0
cc_441 N_A_776_93#_c_599_n RESET_B 0.0397307f $X=5.725 $Y=2.3 $X2=0 $Y2=0
cc_442 N_A_776_93#_c_603_n RESET_B 0.0143367f $X=5.12 $Y=2.465 $X2=0 $Y2=0
cc_443 N_A_776_93#_c_585_n RESET_B 0.0277101f $X=5.945 $Y=1.46 $X2=0 $Y2=0
cc_444 N_A_776_93#_c_586_n RESET_B 4.57232e-19 $X=5.945 $Y=1.46 $X2=0 $Y2=0
cc_445 N_A_776_93#_M1007_g N_RESET_B_c_855_n 0.00427141f $X=5.86 $Y=0.865 $X2=0
+ $Y2=0
cc_446 N_A_776_93#_c_581_n N_RESET_B_c_855_n 0.00258804f $X=5.64 $Y=0.74 $X2=0
+ $Y2=0
cc_447 N_A_776_93#_c_583_n N_RESET_B_c_855_n 5.61579e-19 $X=5.725 $Y=1.295 $X2=0
+ $Y2=0
cc_448 N_A_776_93#_c_585_n N_RESET_B_c_855_n 0.00172393f $X=5.945 $Y=1.46 $X2=0
+ $Y2=0
cc_449 N_A_776_93#_c_586_n N_RESET_B_c_855_n 0.0127892f $X=5.945 $Y=1.46 $X2=0
+ $Y2=0
cc_450 N_A_776_93#_c_600_n N_A_1187_131#_M1016_d 0.00278905f $X=7.225 $Y=2.41
+ $X2=0 $Y2=0
cc_451 N_A_776_93#_c_586_n N_A_1187_131#_c_900_n 0.0087108f $X=5.945 $Y=1.46
+ $X2=0 $Y2=0
cc_452 N_A_776_93#_M1000_g N_A_1187_131#_M1012_g 0.0537136f $X=7.5 $Y=2.465
+ $X2=0 $Y2=0
cc_453 N_A_776_93#_c_600_n N_A_1187_131#_M1012_g 0.0165556f $X=7.225 $Y=2.41
+ $X2=0 $Y2=0
cc_454 N_A_776_93#_c_584_n N_A_1187_131#_M1012_g 0.00817911f $X=7.337 $Y=2.325
+ $X2=0 $Y2=0
cc_455 N_A_776_93#_c_587_n N_A_1187_131#_M1012_g 8.3095e-19 $X=7.55 $Y=1.395
+ $X2=0 $Y2=0
cc_456 N_A_776_93#_c_588_n N_A_1187_131#_M1012_g 0.00615509f $X=7.55 $Y=1.395
+ $X2=0 $Y2=0
cc_457 N_A_776_93#_c_587_n N_A_1187_131#_M1002_g 0.00158491f $X=7.55 $Y=1.395
+ $X2=0 $Y2=0
cc_458 N_A_776_93#_c_588_n N_A_1187_131#_M1002_g 0.0130132f $X=7.55 $Y=1.395
+ $X2=0 $Y2=0
cc_459 N_A_776_93#_c_589_n N_A_1187_131#_M1002_g 0.0138565f $X=7.572 $Y=1.23
+ $X2=0 $Y2=0
cc_460 N_A_776_93#_M1007_g N_A_1187_131#_c_904_n 0.00202686f $X=5.86 $Y=0.865
+ $X2=0 $Y2=0
cc_461 N_A_776_93#_c_583_n N_A_1187_131#_c_904_n 0.0104664f $X=5.725 $Y=1.295
+ $X2=0 $Y2=0
cc_462 N_A_776_93#_M1016_g N_A_1187_131#_c_905_n 0.00309626f $X=5.86 $Y=2.105
+ $X2=0 $Y2=0
cc_463 N_A_776_93#_c_599_n N_A_1187_131#_c_905_n 0.00678853f $X=5.725 $Y=2.3
+ $X2=0 $Y2=0
cc_464 N_A_776_93#_c_585_n N_A_1187_131#_c_906_n 0.00245048f $X=5.945 $Y=1.46
+ $X2=0 $Y2=0
cc_465 N_A_776_93#_c_586_n N_A_1187_131#_c_906_n 0.00397509f $X=5.945 $Y=1.46
+ $X2=0 $Y2=0
cc_466 N_A_776_93#_M1007_g N_A_1187_131#_c_907_n 0.0105684f $X=5.86 $Y=0.865
+ $X2=0 $Y2=0
cc_467 N_A_776_93#_c_583_n N_A_1187_131#_c_907_n 3.8554e-19 $X=5.725 $Y=1.295
+ $X2=0 $Y2=0
cc_468 N_A_776_93#_c_600_n N_A_1187_131#_c_911_n 0.0277605f $X=7.225 $Y=2.41
+ $X2=0 $Y2=0
cc_469 N_A_776_93#_c_585_n N_A_1187_131#_c_911_n 0.00289418f $X=5.945 $Y=1.46
+ $X2=0 $Y2=0
cc_470 N_A_776_93#_c_586_n N_A_1187_131#_c_911_n 0.00410003f $X=5.945 $Y=1.46
+ $X2=0 $Y2=0
cc_471 N_A_776_93#_c_585_n N_A_1187_131#_c_908_n 0.0246186f $X=5.945 $Y=1.46
+ $X2=0 $Y2=0
cc_472 N_A_776_93#_c_586_n N_A_1187_131#_c_908_n 0.00562348f $X=5.945 $Y=1.46
+ $X2=0 $Y2=0
cc_473 N_A_776_93#_c_597_n N_VPWR_M1010_d 0.0102601f $X=4.995 $Y=2.385 $X2=0
+ $Y2=0
cc_474 N_A_776_93#_c_657_p N_VPWR_M1022_d 0.00854487f $X=5.64 $Y=2.397 $X2=0
+ $Y2=0
cc_475 N_A_776_93#_c_599_n N_VPWR_M1022_d 0.00503529f $X=5.725 $Y=2.3 $X2=0
+ $Y2=0
cc_476 N_A_776_93#_c_606_n N_VPWR_M1022_d 3.71002e-19 $X=5.725 $Y=2.397 $X2=0
+ $Y2=0
cc_477 N_A_776_93#_c_600_n N_VPWR_M1012_d 0.00261951f $X=7.225 $Y=2.41 $X2=0
+ $Y2=0
cc_478 N_A_776_93#_c_584_n N_VPWR_M1012_d 0.0047614f $X=7.337 $Y=2.325 $X2=0
+ $Y2=0
cc_479 N_A_776_93#_M1010_g N_VPWR_c_957_n 0.00798116f $X=4.38 $Y=2.835 $X2=0
+ $Y2=0
cc_480 N_A_776_93#_c_597_n N_VPWR_c_957_n 0.0197374f $X=4.995 $Y=2.385 $X2=0
+ $Y2=0
cc_481 N_A_776_93#_c_603_n N_VPWR_c_957_n 0.00112187f $X=5.12 $Y=2.465 $X2=0
+ $Y2=0
cc_482 N_A_776_93#_c_657_p N_VPWR_c_958_n 0.0154514f $X=5.64 $Y=2.397 $X2=0
+ $Y2=0
cc_483 N_A_776_93#_c_603_n N_VPWR_c_958_n 0.0153691f $X=5.12 $Y=2.465 $X2=0
+ $Y2=0
cc_484 N_A_776_93#_c_606_n N_VPWR_c_958_n 0.00659973f $X=5.725 $Y=2.397 $X2=0
+ $Y2=0
cc_485 N_A_776_93#_M1000_g N_VPWR_c_959_n 0.0113958f $X=7.5 $Y=2.465 $X2=0 $Y2=0
cc_486 N_A_776_93#_c_600_n N_VPWR_c_959_n 0.0180131f $X=7.225 $Y=2.41 $X2=0
+ $Y2=0
cc_487 N_A_776_93#_M1016_g N_VPWR_c_960_n 0.00294244f $X=5.86 $Y=2.105 $X2=0
+ $Y2=0
cc_488 N_A_776_93#_M1010_g N_VPWR_c_963_n 0.0053602f $X=4.38 $Y=2.835 $X2=0
+ $Y2=0
cc_489 N_A_776_93#_c_603_n N_VPWR_c_964_n 0.0142733f $X=5.12 $Y=2.465 $X2=0
+ $Y2=0
cc_490 N_A_776_93#_M1000_g N_VPWR_c_965_n 0.00486043f $X=7.5 $Y=2.465 $X2=0
+ $Y2=0
cc_491 N_A_776_93#_M1010_g N_VPWR_c_954_n 0.00636546f $X=4.38 $Y=2.835 $X2=0
+ $Y2=0
cc_492 N_A_776_93#_M1016_g N_VPWR_c_954_n 0.00398527f $X=5.86 $Y=2.105 $X2=0
+ $Y2=0
cc_493 N_A_776_93#_M1000_g N_VPWR_c_954_n 0.00931409f $X=7.5 $Y=2.465 $X2=0
+ $Y2=0
cc_494 N_A_776_93#_c_597_n N_VPWR_c_954_n 0.0107054f $X=4.995 $Y=2.385 $X2=0
+ $Y2=0
cc_495 N_A_776_93#_c_598_n N_VPWR_c_954_n 0.00618754f $X=4.355 $Y=2.385 $X2=0
+ $Y2=0
cc_496 N_A_776_93#_c_657_p N_VPWR_c_954_n 0.00587091f $X=5.64 $Y=2.397 $X2=0
+ $Y2=0
cc_497 N_A_776_93#_c_600_n N_VPWR_c_954_n 0.0452856f $X=7.225 $Y=2.41 $X2=0
+ $Y2=0
cc_498 N_A_776_93#_c_603_n N_VPWR_c_954_n 0.00841451f $X=5.12 $Y=2.465 $X2=0
+ $Y2=0
cc_499 N_A_776_93#_c_606_n N_VPWR_c_954_n 0.00395689f $X=5.725 $Y=2.397 $X2=0
+ $Y2=0
cc_500 N_A_776_93#_c_600_n N_Q_N_M1012_s 0.00774352f $X=7.225 $Y=2.41 $X2=0
+ $Y2=0
cc_501 N_A_776_93#_M1000_g N_Q_N_c_1055_n 4.82647e-19 $X=7.5 $Y=2.465 $X2=0
+ $Y2=0
cc_502 N_A_776_93#_c_600_n N_Q_N_c_1055_n 0.0196663f $X=7.225 $Y=2.41 $X2=0
+ $Y2=0
cc_503 N_A_776_93#_c_584_n N_Q_N_c_1055_n 0.0449743f $X=7.337 $Y=2.325 $X2=0
+ $Y2=0
cc_504 N_A_776_93#_c_587_n N_Q_N_c_1055_n 0.026366f $X=7.55 $Y=1.395 $X2=0 $Y2=0
cc_505 N_A_776_93#_c_588_n N_Q_N_c_1055_n 2.58555e-19 $X=7.55 $Y=1.395 $X2=0
+ $Y2=0
cc_506 N_A_776_93#_c_589_n N_Q_N_c_1055_n 9.83921e-19 $X=7.572 $Y=1.23 $X2=0
+ $Y2=0
cc_507 N_A_776_93#_c_587_n Q 0.00201794f $X=7.55 $Y=1.395 $X2=0 $Y2=0
cc_508 N_A_776_93#_c_588_n Q 0.00366716f $X=7.55 $Y=1.395 $X2=0 $Y2=0
cc_509 N_A_776_93#_c_589_n Q 0.00240756f $X=7.572 $Y=1.23 $X2=0 $Y2=0
cc_510 N_A_776_93#_M1000_g Q 0.00256773f $X=7.5 $Y=2.465 $X2=0 $Y2=0
cc_511 N_A_776_93#_c_584_n Q 0.00554306f $X=7.337 $Y=2.325 $X2=0 $Y2=0
cc_512 N_A_776_93#_c_587_n Q 0.0260579f $X=7.55 $Y=1.395 $X2=0 $Y2=0
cc_513 N_A_776_93#_c_588_n Q 0.00883369f $X=7.55 $Y=1.395 $X2=0 $Y2=0
cc_514 N_A_776_93#_c_589_n Q 0.00402644f $X=7.572 $Y=1.23 $X2=0 $Y2=0
cc_515 N_A_776_93#_M1000_g Q 0.00507951f $X=7.5 $Y=2.465 $X2=0 $Y2=0
cc_516 N_A_776_93#_c_584_n Q 0.0247689f $X=7.337 $Y=2.325 $X2=0 $Y2=0
cc_517 N_A_776_93#_c_587_n Q 0.00193873f $X=7.55 $Y=1.395 $X2=0 $Y2=0
cc_518 N_A_776_93#_c_588_n Q 0.00399242f $X=7.55 $Y=1.395 $X2=0 $Y2=0
cc_519 N_A_776_93#_c_589_n N_Q_c_1079_n 0.00940433f $X=7.572 $Y=1.23 $X2=0 $Y2=0
cc_520 N_A_776_93#_c_581_n N_VGND_M1005_d 0.00969104f $X=5.64 $Y=0.74 $X2=0
+ $Y2=0
cc_521 N_A_776_93#_c_583_n N_VGND_M1005_d 0.00314657f $X=5.725 $Y=1.295 $X2=0
+ $Y2=0
cc_522 N_A_776_93#_M1019_g N_VGND_c_1104_n 0.0035863f $X=3.955 $Y=0.805 $X2=0
+ $Y2=0
cc_523 N_A_776_93#_M1019_g N_VGND_c_1105_n 0.00932459f $X=3.955 $Y=0.805 $X2=0
+ $Y2=0
cc_524 N_A_776_93#_c_580_n N_VGND_c_1105_n 0.0286875f $X=4.71 $Y=0.38 $X2=0
+ $Y2=0
cc_525 N_A_776_93#_c_582_n N_VGND_c_1105_n 0.0129575f $X=4.875 $Y=0.74 $X2=0
+ $Y2=0
cc_526 N_A_776_93#_c_580_n N_VGND_c_1106_n 0.00769519f $X=4.71 $Y=0.38 $X2=0
+ $Y2=0
cc_527 N_A_776_93#_c_581_n N_VGND_c_1106_n 0.0208127f $X=5.64 $Y=0.74 $X2=0
+ $Y2=0
cc_528 N_A_776_93#_c_587_n N_VGND_c_1107_n 0.0166185f $X=7.55 $Y=1.395 $X2=0
+ $Y2=0
cc_529 N_A_776_93#_c_588_n N_VGND_c_1107_n 0.001113f $X=7.55 $Y=1.395 $X2=0
+ $Y2=0
cc_530 N_A_776_93#_c_589_n N_VGND_c_1107_n 0.00297085f $X=7.572 $Y=1.23 $X2=0
+ $Y2=0
cc_531 N_A_776_93#_M1007_g N_VGND_c_1108_n 0.00384999f $X=5.86 $Y=0.865 $X2=0
+ $Y2=0
cc_532 N_A_776_93#_c_581_n N_VGND_c_1108_n 0.00210633f $X=5.64 $Y=0.74 $X2=0
+ $Y2=0
cc_533 N_A_776_93#_c_580_n N_VGND_c_1111_n 0.0208026f $X=4.71 $Y=0.38 $X2=0
+ $Y2=0
cc_534 N_A_776_93#_c_581_n N_VGND_c_1111_n 0.00654693f $X=5.64 $Y=0.74 $X2=0
+ $Y2=0
cc_535 N_A_776_93#_c_589_n N_VGND_c_1112_n 0.00521064f $X=7.572 $Y=1.23 $X2=0
+ $Y2=0
cc_536 N_A_776_93#_M1013_s N_VGND_c_1113_n 0.00215158f $X=4.585 $Y=0.235 $X2=0
+ $Y2=0
cc_537 N_A_776_93#_M1019_g N_VGND_c_1113_n 0.00401353f $X=3.955 $Y=0.805 $X2=0
+ $Y2=0
cc_538 N_A_776_93#_M1007_g N_VGND_c_1113_n 0.0046122f $X=5.86 $Y=0.865 $X2=0
+ $Y2=0
cc_539 N_A_776_93#_c_580_n N_VGND_c_1113_n 0.0125108f $X=4.71 $Y=0.38 $X2=0
+ $Y2=0
cc_540 N_A_776_93#_c_581_n N_VGND_c_1113_n 0.0174771f $X=5.64 $Y=0.74 $X2=0
+ $Y2=0
cc_541 N_A_776_93#_c_589_n N_VGND_c_1113_n 0.0105952f $X=7.572 $Y=1.23 $X2=0
+ $Y2=0
cc_542 N_A_776_93#_c_581_n A_1000_47# 0.00321766f $X=5.64 $Y=0.74 $X2=-0.19
+ $Y2=-0.245
cc_543 N_A_626_119#_c_774_n N_RESET_B_M1005_g 0.0383506f $X=4.925 $Y=1.185 $X2=0
+ $Y2=0
cc_544 N_A_626_119#_M1006_g N_RESET_B_M1022_g 0.0407139f $X=4.905 $Y=2.415 $X2=0
+ $Y2=0
cc_545 N_A_626_119#_M1006_g RESET_B 0.0195346f $X=4.905 $Y=2.415 $X2=0 $Y2=0
cc_546 N_A_626_119#_c_777_n RESET_B 0.023254f $X=4.69 $Y=1.35 $X2=0 $Y2=0
cc_547 N_A_626_119#_c_779_n RESET_B 0.0101426f $X=4.905 $Y=1.35 $X2=0 $Y2=0
cc_548 N_A_626_119#_c_779_n N_RESET_B_c_855_n 0.0502175f $X=4.905 $Y=1.35 $X2=0
+ $Y2=0
cc_549 N_A_626_119#_M1006_g N_VPWR_c_957_n 0.00200386f $X=4.905 $Y=2.415 $X2=0
+ $Y2=0
cc_550 N_A_626_119#_M1006_g N_VPWR_c_958_n 4.87449e-19 $X=4.905 $Y=2.415 $X2=0
+ $Y2=0
cc_551 N_A_626_119#_M1006_g N_VPWR_c_964_n 0.0053602f $X=4.905 $Y=2.415 $X2=0
+ $Y2=0
cc_552 N_A_626_119#_M1006_g N_VPWR_c_954_n 0.00595518f $X=4.905 $Y=2.415 $X2=0
+ $Y2=0
cc_553 N_A_626_119#_c_776_n N_VGND_M1019_d 0.00253411f $X=4.525 $Y=1.08 $X2=0
+ $Y2=0
cc_554 N_A_626_119#_c_775_n N_VGND_c_1104_n 0.00707031f $X=3.5 $Y=1.165 $X2=0
+ $Y2=0
cc_555 N_A_626_119#_c_774_n N_VGND_c_1105_n 0.00222253f $X=4.925 $Y=1.185 $X2=0
+ $Y2=0
cc_556 N_A_626_119#_c_775_n N_VGND_c_1105_n 0.00701997f $X=3.5 $Y=1.165 $X2=0
+ $Y2=0
cc_557 N_A_626_119#_c_776_n N_VGND_c_1105_n 0.0219406f $X=4.525 $Y=1.08 $X2=0
+ $Y2=0
cc_558 N_A_626_119#_c_774_n N_VGND_c_1106_n 0.00185786f $X=4.925 $Y=1.185 $X2=0
+ $Y2=0
cc_559 N_A_626_119#_c_774_n N_VGND_c_1111_n 0.00417814f $X=4.925 $Y=1.185 $X2=0
+ $Y2=0
cc_560 N_A_626_119#_c_774_n N_VGND_c_1113_n 0.00701653f $X=4.925 $Y=1.185 $X2=0
+ $Y2=0
cc_561 N_A_626_119#_c_775_n N_VGND_c_1113_n 0.0108586f $X=3.5 $Y=1.165 $X2=0
+ $Y2=0
cc_562 N_A_626_119#_c_776_n A_734_119# 0.00366293f $X=4.525 $Y=1.08 $X2=-0.19
+ $Y2=-0.245
cc_563 RESET_B N_VPWR_M1022_d 0.00306914f $X=4.955 $Y=1.21 $X2=0 $Y2=0
cc_564 N_RESET_B_M1022_g N_VPWR_c_958_n 0.0111078f $X=5.335 $Y=2.415 $X2=0 $Y2=0
cc_565 N_RESET_B_M1022_g N_VPWR_c_964_n 0.00445056f $X=5.335 $Y=2.415 $X2=0
+ $Y2=0
cc_566 N_RESET_B_M1022_g N_VPWR_c_954_n 0.00436961f $X=5.335 $Y=2.415 $X2=0
+ $Y2=0
cc_567 N_RESET_B_M1005_g N_VGND_c_1106_n 0.0102214f $X=5.285 $Y=0.655 $X2=0
+ $Y2=0
cc_568 N_RESET_B_M1005_g N_VGND_c_1111_n 0.00355956f $X=5.285 $Y=0.655 $X2=0
+ $Y2=0
cc_569 N_RESET_B_M1005_g N_VGND_c_1113_n 0.00406467f $X=5.285 $Y=0.655 $X2=0
+ $Y2=0
cc_570 N_A_1187_131#_M1012_g N_VPWR_c_959_n 0.0247987f $X=7.07 $Y=2.465 $X2=0
+ $Y2=0
cc_571 N_A_1187_131#_M1012_g N_VPWR_c_960_n 0.00486043f $X=7.07 $Y=2.465 $X2=0
+ $Y2=0
cc_572 N_A_1187_131#_M1012_g N_VPWR_c_954_n 0.00600853f $X=7.07 $Y=2.465 $X2=0
+ $Y2=0
cc_573 N_A_1187_131#_c_899_n N_Q_N_c_1055_n 0.0158318f $X=6.995 $Y=1.36 $X2=0
+ $Y2=0
cc_574 N_A_1187_131#_M1012_g N_Q_N_c_1055_n 0.0174494f $X=7.07 $Y=2.465 $X2=0
+ $Y2=0
cc_575 N_A_1187_131#_M1002_g N_Q_N_c_1055_n 0.0177324f $X=7.1 $Y=0.7 $X2=0 $Y2=0
cc_576 N_A_1187_131#_c_903_n N_Q_N_c_1055_n 0.00198231f $X=7.085 $Y=1.36 $X2=0
+ $Y2=0
cc_577 N_A_1187_131#_c_904_n N_Q_N_c_1055_n 0.0310377f $X=6.395 $Y=1.25 $X2=0
+ $Y2=0
cc_578 N_A_1187_131#_c_905_n N_Q_N_c_1055_n 0.0170091f $X=6.295 $Y=1.805 $X2=0
+ $Y2=0
cc_579 N_A_1187_131#_c_906_n N_Q_N_c_1055_n 0.0273628f $X=6.485 $Y=0.93 $X2=0
+ $Y2=0
cc_580 N_A_1187_131#_c_907_n N_Q_N_c_1055_n 0.00459253f $X=6.485 $Y=0.93 $X2=0
+ $Y2=0
cc_581 N_A_1187_131#_c_911_n N_Q_N_c_1055_n 0.015605f $X=6.295 $Y=1.97 $X2=0
+ $Y2=0
cc_582 N_A_1187_131#_M1002_g N_VGND_c_1107_n 0.00288831f $X=7.1 $Y=0.7 $X2=0
+ $Y2=0
cc_583 N_A_1187_131#_M1002_g N_VGND_c_1108_n 0.00499957f $X=7.1 $Y=0.7 $X2=0
+ $Y2=0
cc_584 N_A_1187_131#_c_906_n N_VGND_c_1108_n 0.0096914f $X=6.485 $Y=0.93 $X2=0
+ $Y2=0
cc_585 N_A_1187_131#_c_907_n N_VGND_c_1108_n 0.00221029f $X=6.485 $Y=0.93 $X2=0
+ $Y2=0
cc_586 N_A_1187_131#_M1002_g N_VGND_c_1113_n 0.0102696f $X=7.1 $Y=0.7 $X2=0
+ $Y2=0
cc_587 N_A_1187_131#_c_906_n N_VGND_c_1113_n 0.0166993f $X=6.485 $Y=0.93 $X2=0
+ $Y2=0
cc_588 N_A_1187_131#_c_907_n N_VGND_c_1113_n 0.00184885f $X=6.485 $Y=0.93 $X2=0
+ $Y2=0
cc_589 N_VPWR_c_954_n N_Q_N_M1012_s 0.00389753f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_590 N_VPWR_c_954_n N_Q_M1000_d 0.00371702f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_591 N_VPWR_c_965_n N_Q_c_1082_n 0.03179f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_592 N_VPWR_c_954_n N_Q_c_1082_n 0.0176116f $X=7.92 $Y=3.33 $X2=0 $Y2=0
cc_593 N_Q_N_c_1055_n N_VGND_c_1107_n 0.0303961f $X=6.885 $Y=0.425 $X2=0 $Y2=0
cc_594 N_Q_N_c_1055_n N_VGND_c_1108_n 0.0209548f $X=6.885 $Y=0.425 $X2=0 $Y2=0
cc_595 N_Q_N_c_1055_n N_VGND_c_1113_n 0.0116191f $X=6.885 $Y=0.425 $X2=0 $Y2=0
cc_596 N_Q_c_1079_n N_VGND_c_1107_n 0.0323849f $X=7.77 $Y=0.425 $X2=0 $Y2=0
cc_597 N_Q_c_1079_n N_VGND_c_1112_n 0.0324733f $X=7.77 $Y=0.425 $X2=0 $Y2=0
cc_598 N_Q_c_1079_n N_VGND_c_1113_n 0.0180877f $X=7.77 $Y=0.425 $X2=0 $Y2=0
cc_599 N_VGND_c_1113_n A_1000_47# 0.00250288f $X=7.92 $Y=0 $X2=-0.19 $Y2=-0.245
