* File: sky130_fd_sc_lp__ebufn_1.spice
* Created: Wed Sep  2 09:50:38 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__ebufn_1.pex.spice"
.subckt sky130_fd_sc_lp__ebufn_1  VNB VPB TE_B A Z VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Z	Z
* A	A
* TE_B	TE_B
* VPB	VPB
* VNB	VNB
MM1003 A_171_73# N_A_105_263#_M1003_g N_Z_M1003_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1008 AS=0.2394 PD=1.08 PS=2.25 NRD=9.276 NRS=0 M=1 R=5.6 SA=75000.2
+ SB=75000.6 A=0.126 P=1.98 MULT=1
MM1006 N_VGND_M1006_d N_A_219_21#_M1006_g A_171_73# VNB NSHORT L=0.15 W=0.84
+ AD=0.2394 AS=0.1008 PD=2.25 PS=1.08 NRD=0 NRS=9.276 M=1 R=5.6 SA=75000.6
+ SB=75000.2 A=0.126 P=1.98 MULT=1
MM1002 N_VGND_M1002_d N_TE_B_M1002_g N_A_219_21#_M1002_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0882 AS=0.1197 PD=0.84 PS=1.41 NRD=19.992 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1005 N_A_105_263#_M1005_d N_A_M1005_g N_VGND_M1002_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.0882 PD=1.41 PS=0.84 NRD=0 NRS=19.992 M=1 R=2.8 SA=75000.8
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1007 A_165_367# N_A_105_263#_M1007_g N_Z_M1007_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1512 AS=0.3591 PD=1.5 PS=3.09 NRD=10.1455 NRS=0 M=1 R=8.4 SA=75000.2
+ SB=75000.6 A=0.189 P=2.82 MULT=1
MM1000 N_VPWR_M1000_d N_TE_B_M1000_g A_165_367# VPB PHIGHVT L=0.15 W=1.26
+ AD=0.3591 AS=0.1512 PD=3.09 PS=1.5 NRD=0 NRS=10.1455 M=1 R=8.4 SA=75000.6
+ SB=75000.2 A=0.189 P=2.82 MULT=1
MM1001 N_VPWR_M1001_d N_TE_B_M1001_g N_A_219_21#_M1001_s VPB PHIGHVT L=0.15
+ W=0.64 AD=0.2272 AS=0.1824 PD=1.35 PS=1.85 NRD=126.198 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1004 N_A_105_263#_M1004_d N_A_M1004_g N_VPWR_M1001_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.2144 AS=0.2272 PD=1.95 PS=1.35 NRD=15.3857 NRS=6.1464 M=1 R=4.26667
+ SA=75001.1 SB=75000.3 A=0.096 P=1.58 MULT=1
DX8_noxref VNB VPB NWDIODE A=7.8703 P=12.17
*
.include "sky130_fd_sc_lp__ebufn_1.pxi.spice"
*
.ends
*
*
