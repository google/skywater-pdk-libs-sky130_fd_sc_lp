* NGSPICE file created from sky130_fd_sc_lp__o2bb2a_0.ext - technology: sky130A

.subckt sky130_fd_sc_lp__o2bb2a_0 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
M1000 a_512_47# B1 VGND VNB nshort w=420000u l=150000u
+  ad=2.289e+11p pd=2.77e+06u as=2.352e+11p ps=2.8e+06u
M1001 a_512_47# a_229_483# a_80_176# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1002 VGND a_80_176# X VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1003 a_224_70# A1_N VGND VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=0p ps=0u
M1004 a_229_483# A2_N a_224_70# VNB nshort w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1005 VPWR a_80_176# X VPB phighvt w=640000u l=150000u
+  ad=6.463e+11p pd=5.76e+06u as=1.696e+11p ps=1.81e+06u
M1006 VPWR B1 a_598_483# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1007 a_229_483# A1_N VPWR VPB phighvt w=420000u l=150000u
+  ad=1.785e+11p pd=1.69e+06u as=0p ps=0u
M1008 a_598_483# B2 a_80_176# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=1.176e+11p ps=1.4e+06u
M1009 VPWR A2_N a_229_483# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND B2 a_512_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_80_176# a_229_483# VPWR VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

