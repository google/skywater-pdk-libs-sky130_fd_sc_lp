* File: sky130_fd_sc_lp__nor2_lp2.spice
* Created: Wed Sep  2 10:07:51 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__nor2_lp2.pex.spice"
.subckt sky130_fd_sc_lp__nor2_lp2  VNB VPB A B VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1000 A_130_112# N_A_M1000_g N_VGND_M1000_s VNB NSHORT L=0.15 W=0.42 AD=0.0504
+ AS=0.1197 PD=0.66 PS=1.41 NRD=18.564 NRS=0 M=1 R=2.8 SA=75000.2 SB=75001.4
+ A=0.063 P=1.14 MULT=1
MM1002 N_Y_M1002_d N_A_M1002_g A_130_112# VNB NSHORT L=0.15 W=0.42 AD=0.0588
+ AS=0.0504 PD=0.7 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75000.6 SB=75001
+ A=0.063 P=1.14 MULT=1
MM1003 A_294_112# N_B_M1003_g N_Y_M1002_d VNB NSHORT L=0.15 W=0.42 AD=0.0504
+ AS=0.0588 PD=0.66 PS=0.7 NRD=18.564 NRS=0 M=1 R=2.8 SA=75001 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1001 N_VGND_M1001_d N_B_M1001_g A_294_112# VNB NSHORT L=0.15 W=0.42 AD=0.1197
+ AS=0.0504 PD=1.41 PS=0.66 NRD=0 NRS=18.564 M=1 R=2.8 SA=75001.4 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1005 A_134_374# N_A_M1005_g N_VPWR_M1005_s VPB PHIGHVT L=0.25 W=1 AD=0.105
+ AS=0.285 PD=1.21 PS=2.57 NRD=9.8303 NRS=0 M=1 R=4 SA=125000 SB=125001 A=0.25
+ P=2.5 MULT=1
MM1004 N_Y_M1004_d N_B_M1004_g A_134_374# VPB PHIGHVT L=0.25 W=1 AD=0.265
+ AS=0.105 PD=2.53 PS=1.21 NRD=0 NRS=9.8303 M=1 R=4 SA=125001 SB=125000 A=0.25
+ P=2.5 MULT=1
DX6_noxref VNB VPB NWDIODE A=5.1847 P=9.29
c_22 VNB 0 1.59193e-19 $X=0 $Y=0
*
.include "sky130_fd_sc_lp__nor2_lp2.pxi.spice"
*
.ends
*
*
