* NGSPICE file created from sky130_fd_sc_lp__dlxtn_4.ext - technology: sky130A

.subckt sky130_fd_sc_lp__dlxtn_4 D GATE_N VGND VNB VPB VPWR Q
M1000 VGND a_795_423# Q VNB nshort w=840000u l=150000u
+  ad=1.2012e+12p pd=1.197e+07u as=4.704e+11p ps=4.48e+06u
M1001 VPWR a_795_423# Q VPB phighvt w=1.26e+06u l=150000u
+  ad=2.0957e+12p pd=1.745e+07u as=7.056e+11p ps=6.16e+06u
M1002 a_795_423# a_609_485# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=3.339e+11p pd=3.05e+06u as=0p ps=0u
M1003 a_200_481# GATE_N VPWR VPB phighvt w=640000u l=150000u
+  ad=1.696e+11p pd=1.81e+06u as=0p ps=0u
M1004 a_537_485# a_27_481# VPWR VPB phighvt w=640000u l=150000u
+  ad=1.344e+11p pd=1.7e+06u as=0p ps=0u
M1005 a_717_485# a_200_481# a_609_485# VPB phighvt w=420000u l=150000u
+  ad=1.638e+11p pd=1.62e+06u as=2.221e+11p ps=2.06e+06u
M1006 Q a_795_423# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND D a_27_481# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
M1008 a_200_481# GATE_N VGND VNB nshort w=420000u l=150000u
+  ad=1.113e+11p pd=1.37e+06u as=0p ps=0u
M1009 a_574_47# a_27_481# VGND VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1010 VGND a_795_423# Q VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 Q a_795_423# VPWR VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_609_485# a_200_481# a_574_47# VNB nshort w=420000u l=150000u
+  ad=1.638e+11p pd=1.62e+06u as=0p ps=0u
M1013 VPWR a_795_423# a_717_485# VPB phighvt w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VPWR a_200_481# a_310_485# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.824e+11p ps=1.85e+06u
M1015 a_754_47# a_310_485# a_609_485# VNB nshort w=420000u l=150000u
+  ad=1.638e+11p pd=1.62e+06u as=0p ps=0u
M1016 Q a_795_423# VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VPWR D a_27_481# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.824e+11p ps=1.85e+06u
M1018 Q a_795_423# VGND VNB nshort w=840000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VPWR a_795_423# Q VPB phighvt w=1.26e+06u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_609_485# a_310_485# a_537_485# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_795_423# a_609_485# VGND VNB nshort w=840000u l=150000u
+  ad=2.226e+11p pd=2.21e+06u as=0p ps=0u
M1022 VGND a_795_423# a_754_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 VGND a_200_481# a_310_485# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.113e+11p ps=1.37e+06u
.ends

