* NGSPICE file created from sky130_fd_sc_lp__a41oi_lp.ext - technology: sky130A

.subckt sky130_fd_sc_lp__a41oi_lp A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
M1000 Y A1 a_326_47# VNB nshort w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=1.512e+11p ps=1.56e+06u
M1001 a_248_47# A3 a_170_47# VNB nshort w=420000u l=150000u
+  ad=1.008e+11p pd=1.32e+06u as=1.008e+11p ps=1.32e+06u
M1002 VPWR A2 a_27_409# VPB phighvt w=1e+06u l=250000u
+  ad=5.8e+11p pd=5.16e+06u as=8.45e+11p ps=7.69e+06u
M1003 VPWR A4 a_27_409# VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1004 Y B1 a_27_409# VPB phighvt w=1e+06u l=250000u
+  ad=2.85e+11p pd=2.57e+06u as=0p ps=0u
M1005 a_514_47# B1 Y VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1006 VGND B1 a_514_47# VNB nshort w=420000u l=150000u
+  ad=2.394e+11p pd=2.82e+06u as=0p ps=0u
M1007 a_27_409# A3 VPWR VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_27_409# A1 VPWR VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_326_47# A2 a_248_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_170_47# A4 VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

