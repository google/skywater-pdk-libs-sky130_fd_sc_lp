* NGSPICE file created from sky130_fd_sc_lp__a41oi_0.ext - technology: sky130A

.subckt sky130_fd_sc_lp__a41oi_0 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
M1000 VPWR A3 a_176_479# VPB phighvt w=640000u l=150000u
+  ad=3.584e+11p pd=3.68e+06u as=5.28e+11p ps=5.49e+06u
M1001 a_176_479# B1 Y VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=1.696e+11p ps=1.81e+06u
M1002 a_176_479# A4 VPWR VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_434_47# A3 a_320_47# VNB nshort w=420000u l=150000u
+  ad=1.764e+11p pd=1.68e+06u as=1.764e+11p ps=1.68e+06u
M1004 a_176_479# A2 VPWR VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_320_47# A2 a_230_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.26e+11p ps=1.44e+06u
M1006 Y B1 VGND VNB nshort w=420000u l=150000u
+  ad=1.512e+11p pd=1.56e+06u as=2.226e+11p ps=2.74e+06u
M1007 a_230_47# A1 Y VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND A4 a_434_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR A1 a_176_479# VPB phighvt w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

