* File: sky130_fd_sc_lp__mux2i_m.pex.spice
* Created: Fri Aug 28 10:45:41 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__MUX2I_M%S 3 7 9 11 12 14 16 17 24 25 27 28 30 31 32
+ 34 35 36 38 39 40 45
c111 45 0 1.4009e-19 $X=2.975 $Y=1.32
c112 36 0 4.04057e-20 $X=2.465 $Y=2.41
c113 31 0 1.25504e-19 $X=2.295 $Y=2.98
c114 30 0 1.18063e-19 $X=1.42 $Y=2.895
c115 27 0 1.4496e-19 $X=1.335 $Y=2.385
r116 45 46 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.975
+ $Y=1.32 $X2=2.975 $Y2=1.32
r117 39 40 13.5366 $w=3.13e-07 $l=3.7e-07 $layer=LI1_cond $X=3.047 $Y=1.665
+ $X2=3.047 $Y2=2.035
r118 39 46 12.622 $w=3.13e-07 $l=3.45e-07 $layer=LI1_cond $X=3.047 $Y=1.665
+ $X2=3.047 $Y2=1.32
r119 38 46 0.914637 $w=3.13e-07 $l=2.5e-08 $layer=LI1_cond $X=3.047 $Y=1.295
+ $X2=3.047 $Y2=1.32
r120 37 40 10.6098 $w=3.13e-07 $l=2.9e-07 $layer=LI1_cond $X=3.047 $Y=2.325
+ $X2=3.047 $Y2=2.035
r121 35 37 7.64049 $w=1.7e-07 $l=1.94921e-07 $layer=LI1_cond $X=2.89 $Y=2.41
+ $X2=3.047 $Y2=2.325
r122 35 36 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=2.89 $Y=2.41
+ $X2=2.465 $Y2=2.41
r123 33 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.38 $Y=2.495
+ $X2=2.465 $Y2=2.41
r124 33 34 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=2.38 $Y=2.495
+ $X2=2.38 $Y2=2.895
r125 31 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.295 $Y=2.98
+ $X2=2.38 $Y2=2.895
r126 31 32 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=2.295 $Y=2.98
+ $X2=1.505 $Y2=2.98
r127 30 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.42 $Y=2.895
+ $X2=1.505 $Y2=2.98
r128 29 30 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=1.42 $Y=2.47
+ $X2=1.42 $Y2=2.895
r129 27 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.335 $Y=2.385
+ $X2=1.42 $Y2=2.47
r130 27 28 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=1.335 $Y=2.385
+ $X2=0.69 $Y2=2.385
r131 25 49 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.605 $Y=2.16
+ $X2=0.605 $Y2=2.325
r132 25 48 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=0.605 $Y=2.16
+ $X2=0.605 $Y2=1.995
r133 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.605
+ $Y=2.16 $X2=0.605 $Y2=2.16
r134 22 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.605 $Y=2.3
+ $X2=0.69 $Y2=2.385
r135 22 24 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=0.605 $Y=2.3
+ $X2=0.605 $Y2=2.16
r136 21 45 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=2.975 $Y=1.305
+ $X2=2.975 $Y2=1.32
r137 20 45 59.4528 $w=3.3e-07 $l=3.4e-07 $layer=POLY_cond $X=2.975 $Y=1.66
+ $X2=2.975 $Y2=1.32
r138 16 21 32.1775 $w=1.5e-07 $l=1.98997e-07 $layer=POLY_cond $X=2.81 $Y=1.23
+ $X2=2.975 $Y2=1.305
r139 16 17 94.8617 $w=1.5e-07 $l=1.85e-07 $layer=POLY_cond $X=2.81 $Y=1.23
+ $X2=2.625 $Y2=1.23
r140 12 20 80.3333 $w=1.98e-07 $l=4.01298e-07 $layer=POLY_cond $X=2.645 $Y=1.975
+ $X2=2.975 $Y2=1.817
r141 12 14 369.191 $w=1.5e-07 $l=7.2e-07 $layer=POLY_cond $X=2.645 $Y=1.975
+ $X2=2.645 $Y2=2.695
r142 9 17 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.55 $Y=1.155
+ $X2=2.625 $Y2=1.23
r143 9 11 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.55 $Y=1.155
+ $X2=2.55 $Y2=0.835
r144 7 49 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=0.695 $Y=2.695
+ $X2=0.695 $Y2=2.325
r145 3 48 594.809 $w=1.5e-07 $l=1.16e-06 $layer=POLY_cond $X=0.635 $Y=0.835
+ $X2=0.635 $Y2=1.995
.ends

.subckt PM_SKY130_FD_SC_LP__MUX2I_M%A_55_125# 1 2 9 15 17 18 20 22 25 26 28 30
+ 35 37
c64 25 0 1.22432e-19 $X=1.085 $Y=1.59
r65 32 35 7.65801 $w=2.08e-07 $l=1.45e-07 $layer=LI1_cond $X=0.255 $Y=0.9
+ $X2=0.4 $Y2=0.9
r66 28 30 7.39394 $w=2.08e-07 $l=1.4e-07 $layer=LI1_cond $X=0.34 $Y=2.755
+ $X2=0.48 $Y2=2.755
r67 26 40 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.085 $Y=1.59
+ $X2=1.085 $Y2=1.755
r68 26 39 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.085 $Y=1.59
+ $X2=1.085 $Y2=1.425
r69 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.085
+ $Y=1.59 $X2=1.085 $Y2=1.59
r70 23 37 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.34 $Y=1.59
+ $X2=0.255 $Y2=1.59
r71 23 25 26.0173 $w=3.28e-07 $l=7.45e-07 $layer=LI1_cond $X=0.34 $Y=1.59
+ $X2=1.085 $Y2=1.59
r72 22 28 6.91519 $w=2.1e-07 $l=1.41244e-07 $layer=LI1_cond $X=0.255 $Y=2.65
+ $X2=0.34 $Y2=2.755
r73 21 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.255 $Y=1.755
+ $X2=0.255 $Y2=1.59
r74 21 22 58.3904 $w=1.68e-07 $l=8.95e-07 $layer=LI1_cond $X=0.255 $Y=1.755
+ $X2=0.255 $Y2=2.65
r75 20 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.255 $Y=1.425
+ $X2=0.255 $Y2=1.59
r76 19 32 1.9771 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=0.255 $Y=1.005
+ $X2=0.255 $Y2=0.9
r77 19 20 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=0.255 $Y=1.005
+ $X2=0.255 $Y2=1.425
r78 17 18 58.3064 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=1.19 $Y=1.995
+ $X2=1.19 $Y2=2.145
r79 17 40 123.064 $w=1.5e-07 $l=2.4e-07 $layer=POLY_cond $X=1.175 $Y=1.995
+ $X2=1.175 $Y2=1.755
r80 15 18 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=1.205 $Y=2.695
+ $X2=1.205 $Y2=2.145
r81 9 39 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=1.175 $Y=0.835
+ $X2=1.175 $Y2=1.425
r82 2 30 600 $w=1.7e-07 $l=3.26573e-07 $layer=licon1_PDIFF $count=1 $X=0.355
+ $Y=2.485 $X2=0.48 $Y2=2.755
r83 1 35 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=0.275
+ $Y=0.625 $X2=0.4 $Y2=0.9
.ends

.subckt PM_SKY130_FD_SC_LP__MUX2I_M%A1 3 7 10 12 13 15 16 17 22 28 37
c69 28 0 3.23572e-19 $X=1.985 $Y=0.515
c70 22 0 7.26368e-20 $X=1.655 $Y=1.94
r71 22 25 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.655 $Y=1.94
+ $X2=1.655 $Y2=2.105
r72 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.655
+ $Y=1.94 $X2=1.655 $Y2=1.94
r73 17 23 2.67029 $w=4.08e-07 $l=9.5e-08 $layer=LI1_cond $X=1.56 $Y=2.035
+ $X2=1.56 $Y2=1.94
r74 16 23 7.7298 $w=4.08e-07 $l=2.75e-07 $layer=LI1_cond $X=1.56 $Y=1.665
+ $X2=1.56 $Y2=1.94
r75 16 29 7.02709 $w=4.08e-07 $l=2.5e-07 $layer=LI1_cond $X=1.56 $Y=1.665
+ $X2=1.56 $Y2=1.415
r76 15 29 3.373 $w=4.08e-07 $l=1.2e-07 $layer=LI1_cond $X=1.56 $Y=1.295 $X2=1.56
+ $Y2=1.415
r77 15 37 6.44206 $w=4.08e-07 $l=8.5e-08 $layer=LI1_cond $X=1.56 $Y=1.295
+ $X2=1.56 $Y2=1.21
r78 13 28 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=1.985 $Y=0.35
+ $X2=1.985 $Y2=0.515
r79 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.985
+ $Y=0.35 $X2=1.985 $Y2=0.35
r80 10 12 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=1.525 $Y=0.35
+ $X2=1.985 $Y2=0.35
r81 8 10 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.44 $Y=0.435
+ $X2=1.525 $Y2=0.35
r82 8 37 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=1.44 $Y=0.435
+ $X2=1.44 $Y2=1.21
r83 7 28 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.005 $Y=0.835
+ $X2=2.005 $Y2=0.515
r84 3 25 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=1.565 $Y=2.695
+ $X2=1.565 $Y2=2.105
.ends

.subckt PM_SKY130_FD_SC_LP__MUX2I_M%A0 3 5 6 7 9 11
c51 11 0 2.32244e-19 $X=2.16 $Y=1.665
c52 9 0 1.4496e-19 $X=2.185 $Y=2.695
c53 6 0 1.22432e-19 $X=1.64 $Y=1.49
r54 11 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.195
+ $Y=1.71 $X2=2.195 $Y2=1.71
r55 7 15 38.7444 $w=2.79e-07 $l=1.69926e-07 $layer=POLY_cond $X=2.185 $Y=1.875
+ $X2=2.195 $Y2=1.71
r56 7 9 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=2.185 $Y=1.875
+ $X2=2.185 $Y2=2.695
r57 5 15 38.0072 $w=2.79e-07 $l=2.91033e-07 $layer=POLY_cond $X=2.03 $Y=1.49
+ $X2=2.195 $Y2=1.71
r58 5 6 199.979 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=2.03 $Y=1.49 $X2=1.64
+ $Y2=1.49
r59 1 6 25.2915 $w=1.59e-07 $l=1.69558e-07 $layer=POLY_cond $X=1.535 $Y=1.365
+ $X2=1.64 $Y2=1.49
r60 1 3 271.766 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=1.535 $Y=1.365
+ $X2=1.535 $Y2=0.835
.ends

.subckt PM_SKY130_FD_SC_LP__MUX2I_M%VPWR 1 2 9 11 13 16 17 18 24 33
r38 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r39 30 33 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=2.64 $Y=3.33
+ $X2=3.12 $Y2=3.33
r40 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=3.33
+ $X2=2.64 $Y2=3.33
r41 26 29 93.9465 $w=1.68e-07 $l=1.44e-06 $layer=LI1_cond $X=1.2 $Y=3.33
+ $X2=2.64 $Y2=3.33
r42 26 27 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=3.33 $X2=1.2
+ $Y2=3.33
r43 24 32 4.51706 $w=1.7e-07 $l=2.85e-07 $layer=LI1_cond $X=2.79 $Y=3.33
+ $X2=3.075 $Y2=3.33
r44 24 29 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=2.79 $Y=3.33 $X2=2.64
+ $Y2=3.33
r45 22 27 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=3.33
+ $X2=1.2 $Y2=3.33
r46 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r47 18 30 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=2.64 $Y2=3.33
r48 18 27 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=3.33
+ $X2=1.2 $Y2=3.33
r49 16 21 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=0.825 $Y=3.33
+ $X2=0.72 $Y2=3.33
r50 16 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.825 $Y=3.33
+ $X2=0.99 $Y2=3.33
r51 15 26 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=1.155 $Y=3.33
+ $X2=1.2 $Y2=3.33
r52 15 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.155 $Y=3.33
+ $X2=0.99 $Y2=3.33
r53 11 32 3.24911 $w=3.3e-07 $l=1.56844e-07 $layer=LI1_cond $X=2.955 $Y=3.245
+ $X2=3.075 $Y2=3.33
r54 11 13 16.9374 $w=3.28e-07 $l=4.85e-07 $layer=LI1_cond $X=2.955 $Y=3.245
+ $X2=2.955 $Y2=2.76
r55 7 17 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.99 $Y=3.245 $X2=0.99
+ $Y2=3.33
r56 7 9 16.9374 $w=3.28e-07 $l=4.85e-07 $layer=LI1_cond $X=0.99 $Y=3.245
+ $X2=0.99 $Y2=2.76
r57 2 13 600 $w=1.7e-07 $l=3.745e-07 $layer=licon1_PDIFF $count=1 $X=2.72
+ $Y=2.485 $X2=2.955 $Y2=2.76
r58 1 9 600 $w=1.7e-07 $l=3.68951e-07 $layer=licon1_PDIFF $count=1 $X=0.77
+ $Y=2.485 $X2=0.99 $Y2=2.76
.ends

.subckt PM_SKY130_FD_SC_LP__MUX2I_M%Y 1 2 8 9 10 11 14 18 20
c64 11 0 1.63966e-19 $X=2.54 $Y=1.14
r65 20 32 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=2.16 $Y=0.925
+ $X2=2.16 $Y2=1.14
r66 20 25 8.20134 $w=4.98e-07 $l=2.85e-07 $layer=LI1_cond $X=2.075 $Y=0.865
+ $X2=1.79 $Y2=0.865
r67 16 18 9.04785 $w=1.88e-07 $l=1.55e-07 $layer=LI1_cond $X=1.875 $Y=2.62
+ $X2=2.03 $Y2=2.62
r68 13 14 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=2.625 $Y=1.225
+ $X2=2.625 $Y2=1.975
r69 12 32 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.245 $Y=1.14
+ $X2=2.16 $Y2=1.14
r70 11 13 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.54 $Y=1.14
+ $X2=2.625 $Y2=1.225
r71 11 12 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=2.54 $Y=1.14
+ $X2=2.245 $Y2=1.14
r72 9 14 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.54 $Y=2.06
+ $X2=2.625 $Y2=1.975
r73 9 10 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=2.54 $Y=2.06
+ $X2=2.115 $Y2=2.06
r74 8 18 1.386 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.03 $Y=2.525 $X2=2.03
+ $Y2=2.62
r75 7 10 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.03 $Y=2.145
+ $X2=2.115 $Y2=2.06
r76 7 8 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=2.03 $Y=2.145 $X2=2.03
+ $Y2=2.525
r77 2 16 600 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_PDIFF $count=1 $X=1.64
+ $Y=2.485 $X2=1.875 $Y2=2.63
r78 1 25 182 $w=1.7e-07 $l=3.1749e-07 $layer=licon1_NDIFF $count=1 $X=1.61
+ $Y=0.625 $X2=1.79 $Y2=0.865
.ends

.subckt PM_SKY130_FD_SC_LP__MUX2I_M%VGND 1 2 9 13 16 17 18 24 30 31 34
r38 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.64 $Y=0 $X2=2.64
+ $Y2=0
r39 31 35 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.12 $Y=0 $X2=2.64
+ $Y2=0
r40 30 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r41 28 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.93 $Y=0 $X2=2.765
+ $Y2=0
r42 28 30 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=2.93 $Y=0 $X2=3.12
+ $Y2=0
r43 26 27 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r44 24 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.6 $Y=0 $X2=2.765
+ $Y2=0
r45 24 26 91.3369 $w=1.68e-07 $l=1.4e-06 $layer=LI1_cond $X=2.6 $Y=0 $X2=1.2
+ $Y2=0
r46 22 27 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.72 $Y=0 $X2=1.2
+ $Y2=0
r47 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r48 18 35 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=2.64
+ $Y2=0
r49 18 27 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.68 $Y=0 $X2=1.2
+ $Y2=0
r50 16 21 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=0.745 $Y=0 $X2=0.72
+ $Y2=0
r51 16 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.745 $Y=0 $X2=0.91
+ $Y2=0
r52 15 26 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=1.075 $Y=0 $X2=1.2
+ $Y2=0
r53 15 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.075 $Y=0 $X2=0.91
+ $Y2=0
r54 11 34 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.765 $Y=0.085
+ $X2=2.765 $Y2=0
r55 11 13 23.9219 $w=3.28e-07 $l=6.85e-07 $layer=LI1_cond $X=2.765 $Y=0.085
+ $X2=2.765 $Y2=0.77
r56 7 17 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.91 $Y=0.085 $X2=0.91
+ $Y2=0
r57 7 9 23.9219 $w=3.28e-07 $l=6.85e-07 $layer=LI1_cond $X=0.91 $Y=0.085
+ $X2=0.91 $Y2=0.77
r58 2 13 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=2.625
+ $Y=0.625 $X2=2.765 $Y2=0.77
r59 1 9 182 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_NDIFF $count=1 $X=0.71
+ $Y=0.625 $X2=0.91 $Y2=0.77
.ends

