* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_lp__and4b_m A_N B C D VGND VNB VPB VPWR X
X0 a_27_55# A_N VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 VPWR C a_240_73# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X2 a_240_73# a_27_55# a_323_73# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 VPWR a_27_55# a_240_73# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X4 a_395_73# C a_467_73# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 VPWR a_240_73# X VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X6 a_467_73# D VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 a_240_73# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X8 VGND a_240_73# X VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 a_240_73# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X10 a_27_55# A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=150000u
X11 a_323_73# B a_395_73# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
