* File: sky130_fd_sc_lp__a32oi_0.spice
* Created: Fri Aug 28 10:01:30 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__a32oi_0.pex.spice"
.subckt sky130_fd_sc_lp__a32oi_0  VNB VPB B2 B1 A1 A2 A3 Y VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Y	Y
* A3	A3
* A2	A2
* A1	A1
* B1	B1
* B2	B2
* VPB	VPB
* VNB	VNB
MM1005 A_141_47# N_B2_M1005_g N_VGND_M1005_s VNB NSHORT L=0.15 W=0.42 AD=0.0504
+ AS=0.1386 PD=0.66 PS=1.5 NRD=18.564 NRS=18.564 M=1 R=2.8 SA=75000.3 SB=75002.3
+ A=0.063 P=1.14 MULT=1
MM1002 N_Y_M1002_d N_B1_M1002_g A_141_47# VNB NSHORT L=0.15 W=0.42 AD=0.0882
+ AS=0.0504 PD=0.84 PS=0.66 NRD=7.14 NRS=18.564 M=1 R=2.8 SA=75000.6 SB=75001.9
+ A=0.063 P=1.14 MULT=1
MM1009 A_333_47# N_A1_M1009_g N_Y_M1002_d VNB NSHORT L=0.15 W=0.42 AD=0.0882
+ AS=0.0882 PD=0.84 PS=0.84 NRD=44.28 NRS=32.856 M=1 R=2.8 SA=75001.2 SB=75001.3
+ A=0.063 P=1.14 MULT=1
MM1004 A_447_47# N_A2_M1004_g A_333_47# VNB NSHORT L=0.15 W=0.42 AD=0.0819
+ AS=0.0882 PD=0.81 PS=0.84 NRD=39.996 NRS=44.28 M=1 R=2.8 SA=75001.8 SB=75000.7
+ A=0.063 P=1.14 MULT=1
MM1007 N_VGND_M1007_d N_A3_M1007_g A_447_47# VNB NSHORT L=0.15 W=0.42 AD=0.1113
+ AS=0.0819 PD=1.37 PS=0.81 NRD=0 NRS=39.996 M=1 R=2.8 SA=75002.3 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1001 N_Y_M1001_d N_B2_M1001_g N_A_37_397#_M1001_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0896 AS=0.1696 PD=0.92 PS=1.81 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.2
+ SB=75002.2 A=0.096 P=1.58 MULT=1
MM1008 N_A_37_397#_M1008_d N_B1_M1008_g N_Y_M1001_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0896 AS=0.0896 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667 SA=75000.6
+ SB=75001.8 A=0.096 P=1.58 MULT=1
MM1003 N_VPWR_M1003_d N_A1_M1003_g N_A_37_397#_M1008_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1984 AS=0.0896 PD=1.26 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667 SA=75001.1
+ SB=75001.4 A=0.096 P=1.58 MULT=1
MM1006 N_A_37_397#_M1006_d N_A2_M1006_g N_VPWR_M1003_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0896 AS=0.1984 PD=0.92 PS=1.26 NRD=0 NRS=0 M=1 R=4.26667 SA=75001.8
+ SB=75000.6 A=0.096 P=1.58 MULT=1
MM1000 N_VPWR_M1000_d N_A3_M1000_g N_A_37_397#_M1006_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1696 AS=0.0896 PD=1.81 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667 SA=75002.2
+ SB=75000.2 A=0.096 P=1.58 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.9751 P=11.21
*
.include "sky130_fd_sc_lp__a32oi_0.pxi.spice"
*
.ends
*
*
