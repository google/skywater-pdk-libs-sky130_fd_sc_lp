* File: sky130_fd_sc_lp__mux4_2.spice
* Created: Fri Aug 28 10:46:12 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_lp__mux4_2.pex.spice"
.subckt sky130_fd_sc_lp__mux4_2  VNB VPB S1 A3 A2 A1 A0 S0 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* S0	S0
* A0	A0
* A1	A1
* A2	A2
* A3	A3
* S1	S1
* VPB	VPB
* VNB	VNB
MM1013 N_A_110_125#_M1013_d N_S1_M1013_g N_A_27_125#_M1013_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0588 AS=0.1113 PD=0.7 PS=1.37 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1003 N_A_196_125#_M1003_d N_A_80_293#_M1003_g N_A_110_125#_M1013_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.1113 AS=0.0588 PD=1.37 PS=0.7 NRD=0 NRS=0 M=1 R=2.8
+ SA=75000.6 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1023 N_VGND_M1023_d N_S1_M1023_g N_A_80_293#_M1023_s VNB NSHORT L=0.15 W=0.42
+ AD=0.127267 AS=0.1709 PD=0.943333 PS=1.66 NRD=70.86 NRS=32.856 M=1 R=2.8
+ SA=75000.3 SB=75005.1 A=0.063 P=1.14 MULT=1
MM1015 N_X_M1015_d N_A_110_125#_M1015_g N_VGND_M1023_d VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.254533 PD=1.12 PS=1.88667 NRD=0 NRS=12.132 M=1 R=5.6 SA=75000.6
+ SB=75002.9 A=0.126 P=1.98 MULT=1
MM1024 N_X_M1015_d N_A_110_125#_M1024_g N_VGND_M1024_s VNB NSHORT L=0.15 W=0.84
+ AD=0.1176 AS=0.2212 PD=1.12 PS=1.82 NRD=0 NRS=17.496 M=1 R=5.6 SA=75001
+ SB=75002.4 A=0.126 P=1.98 MULT=1
MM1018 A_825_119# N_A3_M1018_g N_VGND_M1024_s VNB NSHORT L=0.15 W=0.42 AD=0.0441
+ AS=0.1106 PD=0.63 PS=0.91 NRD=14.28 NRS=0 M=1 R=2.8 SA=75002 SB=75004 A=0.063
+ P=1.14 MULT=1
MM1009 N_A_27_125#_M1009_d N_S0_M1009_g A_825_119# VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75002.3
+ SB=75003.6 A=0.063 P=1.14 MULT=1
MM1011 A_983_119# N_A_859_351#_M1011_g N_A_27_125#_M1009_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0672 AS=0.0588 PD=0.74 PS=0.7 NRD=30 NRS=0 M=1 R=2.8 SA=75002.8
+ SB=75003.2 A=0.063 P=1.14 MULT=1
MM1020 N_VGND_M1020_d N_A2_M1020_g A_983_119# VNB NSHORT L=0.15 W=0.42 AD=0.1218
+ AS=0.0672 PD=1 PS=0.74 NRD=35.712 NRS=30 M=1 R=2.8 SA=75003.2 SB=75002.7
+ A=0.063 P=1.14 MULT=1
MM1007 A_1223_119# N_A1_M1007_g N_VGND_M1020_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1218 PD=0.63 PS=1 NRD=14.28 NRS=49.992 M=1 R=2.8 SA=75004
+ SB=75002 A=0.063 P=1.14 MULT=1
MM1000 N_A_196_125#_M1000_d N_S0_M1000_g A_1223_119# VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0441 PD=0.7 PS=0.63 NRD=0 NRS=14.28 M=1 R=2.8 SA=75004.3
+ SB=75001.6 A=0.063 P=1.14 MULT=1
MM1001 A_1381_119# N_A_859_351#_M1001_g N_A_196_125#_M1000_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0672 AS=0.0588 PD=0.74 PS=0.7 NRD=30 NRS=0 M=1 R=2.8 SA=75004.7
+ SB=75001.2 A=0.063 P=1.14 MULT=1
MM1004 N_VGND_M1004_d N_A0_M1004_g A_1381_119# VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.0672 PD=0.7 PS=0.74 NRD=0 NRS=30 M=1 R=2.8 SA=75005.2
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1006 N_A_859_351#_M1006_d N_S0_M1006_g N_VGND_M1004_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1617 AS=0.0588 PD=1.61 PS=0.7 NRD=0 NRS=0 M=1 R=2.8 SA=75005.6 SB=75000.3
+ A=0.063 P=1.14 MULT=1
MM1005 N_A_110_125#_M1005_d N_A_80_293#_M1005_g N_A_27_125#_M1005_s VPB PHIGHVT
+ L=0.15 W=0.64 AD=0.0896 AS=0.1696 PD=0.92 PS=1.81 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.2 SB=75000.6 A=0.096 P=1.58 MULT=1
MM1017 N_A_196_125#_M1017_d N_S1_M1017_g N_A_110_125#_M1005_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1696 AS=0.0896 PD=1.81 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75000.6 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1025 N_VPWR_M1025_d N_S1_M1025_g N_A_80_293#_M1025_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.209482 AS=0.2029 PD=1.33053 PS=2 NRD=83.8038 NRS=29.2348 M=1 R=4.26667
+ SA=75000.2 SB=75003.7 A=0.096 P=1.58 MULT=1
MM1002 N_X_M1002_d N_A_110_125#_M1002_g N_VPWR_M1025_d VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.412418 PD=1.54 PS=2.61947 NRD=0 NRS=0 M=1 R=8.4 SA=75000.7
+ SB=75002.9 A=0.189 P=2.82 MULT=1
MM1019 N_X_M1002_d N_A_110_125#_M1019_g N_VPWR_M1019_s VPB PHIGHVT L=0.15 W=1.26
+ AD=0.1764 AS=0.331778 PD=1.54 PS=2.36747 NRD=0 NRS=0 M=1 R=8.4 SA=75001.1
+ SB=75002.5 A=0.189 P=2.82 MULT=1
MM1021 A_817_419# N_A3_M1021_g N_VPWR_M1019_s VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0672 AS=0.168522 PD=0.85 PS=1.20253 NRD=15.3857 NRS=64.1038 M=1 R=4.26667
+ SA=75001.8 SB=75004 A=0.096 P=1.58 MULT=1
MM1026 N_A_27_125#_M1026_d N_A_859_351#_M1026_g A_817_419# VPB PHIGHVT L=0.15
+ W=0.64 AD=0.0896 AS=0.0672 PD=0.92 PS=0.85 NRD=0 NRS=15.3857 M=1 R=4.26667
+ SA=75002.1 SB=75003.7 A=0.096 P=1.58 MULT=1
MM1012 A_975_419# N_S0_M1012_g N_A_27_125#_M1026_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0672 AS=0.0896 PD=0.85 PS=0.92 NRD=15.3857 NRS=0 M=1 R=4.26667 SA=75002.6
+ SB=75003.3 A=0.096 P=1.58 MULT=1
MM1010 N_VPWR_M1010_d N_A2_M1010_g A_975_419# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.2336 AS=0.0672 PD=1.37 PS=0.85 NRD=0 NRS=15.3857 M=1 R=4.26667 SA=75002.9
+ SB=75002.9 A=0.096 P=1.58 MULT=1
MM1022 A_1223_419# N_A1_M1022_g N_VPWR_M1010_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0672 AS=0.2336 PD=0.85 PS=1.37 NRD=15.3857 NRS=138.511 M=1 R=4.26667
+ SA=75003.8 SB=75002 A=0.096 P=1.58 MULT=1
MM1027 N_A_196_125#_M1027_d N_A_859_351#_M1027_g A_1223_419# VPB PHIGHVT L=0.15
+ W=0.64 AD=0.12 AS=0.0672 PD=1.015 PS=0.85 NRD=15.3857 NRS=15.3857 M=1
+ R=4.26667 SA=75004.2 SB=75001.7 A=0.096 P=1.58 MULT=1
MM1014 A_1400_419# N_S0_M1014_g N_A_196_125#_M1027_d VPB PHIGHVT L=0.15 W=0.64
+ AD=0.1152 AS=0.12 PD=1 PS=1.015 NRD=38.4741 NRS=13.8491 M=1 R=4.26667
+ SA=75004.7 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1016 N_VPWR_M1016_d N_A0_M1016_g A_1400_419# VPB PHIGHVT L=0.15 W=0.64
+ AD=0.0896 AS=0.1152 PD=0.92 PS=1 NRD=0 NRS=38.4741 M=1 R=4.26667 SA=75005.2
+ SB=75000.6 A=0.096 P=1.58 MULT=1
MM1008 N_A_859_351#_M1008_d N_S0_M1008_g N_VPWR_M1016_d VPB PHIGHVT L=0.15
+ W=0.64 AD=0.1696 AS=0.0896 PD=1.81 PS=0.92 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75005.6 SB=75000.2 A=0.096 P=1.58 MULT=1
DX28_noxref VNB VPB NWDIODE A=16.9681 P=21.89
c_1241 A_1381_119# 0 6.87706e-20 $X=6.905 $Y=0.595
*
.include "sky130_fd_sc_lp__mux4_2.pxi.spice"
*
.ends
*
*
