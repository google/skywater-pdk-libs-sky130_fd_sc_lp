* File: sky130_fd_sc_lp__decapkapwr_4.pxi.spice
* Created: Fri Aug 28 10:20:36 2020
* 
x_PM_SKY130_FD_SC_LP__DECAPKAPWR_4%VGND N_VGND_M1001_s N_VGND_c_24_n
+ N_VGND_M1000_g N_VGND_c_25_n N_VGND_c_26_n N_VGND_c_27_n N_VGND_c_28_n
+ N_VGND_c_29_n VGND N_VGND_c_30_n N_VGND_c_31_n
+ PM_SKY130_FD_SC_LP__DECAPKAPWR_4%VGND
x_PM_SKY130_FD_SC_LP__DECAPKAPWR_4%KAPWR N_KAPWR_M1000_s N_KAPWR_c_57_n
+ N_KAPWR_c_58_n N_KAPWR_c_67_n N_KAPWR_c_55_n N_KAPWR_c_60_n N_KAPWR_c_61_n
+ KAPWR N_KAPWR_M1001_g N_KAPWR_c_63_n PM_SKY130_FD_SC_LP__DECAPKAPWR_4%KAPWR
x_PM_SKY130_FD_SC_LP__DECAPKAPWR_4%VPWR VPWR N_VPWR_c_93_n VPWR
+ PM_SKY130_FD_SC_LP__DECAPKAPWR_4%VPWR
cc_1 VNB N_VGND_c_24_n 0.0113126f $X=-0.19 $Y=-0.245 $X2=0.91 $Y2=1.935
cc_2 VNB N_VGND_c_25_n 0.012758f $X=-0.19 $Y=-0.245 $X2=0.335 $Y2=0.085
cc_3 VNB N_VGND_c_26_n 0.0607496f $X=-0.19 $Y=-0.245 $X2=0.335 $Y2=0.38
cc_4 VNB N_VGND_c_27_n 0.0118011f $X=-0.19 $Y=-0.245 $X2=1.615 $Y2=0.085
cc_5 VNB N_VGND_c_28_n 0.0365905f $X=-0.19 $Y=-0.245 $X2=1.615 $Y2=0.36
cc_6 VNB N_VGND_c_29_n 0.00314375f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=1.77
cc_7 VNB N_VGND_c_30_n 0.0280737f $X=-0.19 $Y=-0.245 $X2=1.45 $Y2=0
cc_8 VNB N_VGND_c_31_n 0.132299f $X=-0.19 $Y=-0.245 $X2=1.68 $Y2=0
cc_9 VNB N_KAPWR_c_55_n 0.0270854f $X=-0.19 $Y=-0.245 $X2=0.335 $Y2=0.38
cc_10 VNB N_KAPWR_M1001_g 0.123316f $X=-0.19 $Y=-0.245 $X2=0.575 $Y2=1.77
cc_11 VNB VPWR 0.0840719f $X=-0.19 $Y=-0.245 $X2=0.21 $Y2=0.235
cc_12 VPB N_VGND_c_24_n 0.0464251f $X=-0.19 $Y=1.655 $X2=0.91 $Y2=1.935
cc_13 VPB N_VGND_M1000_g 0.0868293f $X=-0.19 $Y=1.655 $X2=0.91 $Y2=2.595
cc_14 VPB N_VGND_c_29_n 0.0173225f $X=-0.19 $Y=1.655 $X2=0.575 $Y2=1.77
cc_15 VPB N_KAPWR_c_57_n 0.00922717f $X=-0.19 $Y=1.655 $X2=0.91 $Y2=1.935
cc_16 VPB N_KAPWR_c_58_n 0.023615f $X=-0.19 $Y=1.655 $X2=0.91 $Y2=2.595
cc_17 VPB N_KAPWR_c_55_n 0.00182185f $X=-0.19 $Y=1.655 $X2=0.335 $Y2=0.38
cc_18 VPB N_KAPWR_c_60_n 0.0105637f $X=-0.19 $Y=1.655 $X2=0.335 $Y2=0.38
cc_19 VPB N_KAPWR_c_61_n 0.0461607f $X=-0.19 $Y=1.655 $X2=0.335 $Y2=1.06
cc_20 VPB N_KAPWR_M1001_g 0.00822137f $X=-0.19 $Y=1.655 $X2=0.575 $Y2=1.77
cc_21 VPB N_KAPWR_c_63_n 0.0254524f $X=-0.19 $Y=1.655 $X2=1.2 $Y2=0
cc_22 VPB VPWR 0.0430995f $X=-0.19 $Y=1.655 $X2=0.21 $Y2=0.235
cc_23 VPB N_VPWR_c_93_n 0.0520213f $X=-0.19 $Y=1.655 $X2=0.91 $Y2=2.595
cc_24 N_VGND_M1000_g N_KAPWR_c_57_n 0.00685959f $X=0.91 $Y=2.595 $X2=0 $Y2=0
cc_25 N_VGND_M1000_g N_KAPWR_c_58_n 0.028057f $X=0.91 $Y=2.595 $X2=0 $Y2=0
cc_26 N_VGND_c_29_n N_KAPWR_c_58_n 0.0192408f $X=0.575 $Y=1.77 $X2=0 $Y2=0
cc_27 N_VGND_M1000_g N_KAPWR_c_67_n 0.056773f $X=0.91 $Y=2.595 $X2=0 $Y2=0
cc_28 N_VGND_c_24_n N_KAPWR_c_55_n 0.00168098f $X=0.91 $Y=1.935 $X2=0 $Y2=0
cc_29 N_VGND_c_28_n N_KAPWR_c_55_n 0.021547f $X=1.615 $Y=0.36 $X2=0 $Y2=0
cc_30 N_VGND_c_29_n N_KAPWR_c_55_n 0.00259429f $X=0.575 $Y=1.77 $X2=0 $Y2=0
cc_31 N_VGND_M1000_g N_KAPWR_c_60_n 0.00746086f $X=0.91 $Y=2.595 $X2=0 $Y2=0
cc_32 N_VGND_c_24_n N_KAPWR_c_61_n 0.00401381f $X=0.91 $Y=1.935 $X2=0 $Y2=0
cc_33 N_VGND_M1000_g N_KAPWR_c_61_n 0.0410524f $X=0.91 $Y=2.595 $X2=0 $Y2=0
cc_34 N_VGND_c_29_n N_KAPWR_c_61_n 0.00767335f $X=0.575 $Y=1.77 $X2=0 $Y2=0
cc_35 N_VGND_c_24_n N_KAPWR_M1001_g 0.0523192f $X=0.91 $Y=1.935 $X2=0 $Y2=0
cc_36 N_VGND_c_26_n N_KAPWR_M1001_g 0.0687615f $X=0.335 $Y=0.38 $X2=0 $Y2=0
cc_37 N_VGND_c_28_n N_KAPWR_M1001_g 0.0510153f $X=1.615 $Y=0.36 $X2=0 $Y2=0
cc_38 N_VGND_c_29_n N_KAPWR_M1001_g 0.00192223f $X=0.575 $Y=1.77 $X2=0 $Y2=0
cc_39 N_VGND_c_30_n N_KAPWR_M1001_g 0.0370388f $X=1.45 $Y=0 $X2=0 $Y2=0
cc_40 N_VGND_c_31_n N_KAPWR_M1001_g 0.0582443f $X=1.68 $Y=0 $X2=0 $Y2=0
cc_41 N_VGND_M1000_g N_KAPWR_c_63_n 0.0476516f $X=0.91 $Y=2.595 $X2=0 $Y2=0
cc_42 N_VGND_M1000_g VPWR 0.0248614f $X=0.91 $Y=2.595 $X2=-0.19 $Y2=-0.245
cc_43 N_VGND_M1000_g N_VPWR_c_93_n 0.0268474f $X=0.91 $Y=2.595 $X2=0 $Y2=0
cc_44 N_KAPWR_M1000_s VPWR 0.00234386f $X=0.135 $Y=2.095 $X2=-0.19 $Y2=-0.245
cc_45 N_KAPWR_c_57_n VPWR 0.00306712f $X=0.26 $Y=2.675 $X2=-0.19 $Y2=-0.245
cc_46 N_KAPWR_c_67_n VPWR 0.00490555f $X=1.385 $Y=2.81 $X2=-0.19 $Y2=-0.245
cc_47 N_KAPWR_c_60_n VPWR 0.00375641f $X=1.587 $Y=2.675 $X2=-0.19 $Y2=-0.245
cc_48 N_KAPWR_c_63_n VPWR 0.187606f $X=1.705 $Y=2.81 $X2=-0.19 $Y2=-0.245
cc_49 N_KAPWR_c_57_n N_VPWR_c_93_n 0.0212079f $X=0.26 $Y=2.675 $X2=0 $Y2=0
cc_50 N_KAPWR_c_67_n N_VPWR_c_93_n 0.0319042f $X=1.385 $Y=2.81 $X2=0 $Y2=0
cc_51 N_KAPWR_c_60_n N_VPWR_c_93_n 0.0265029f $X=1.587 $Y=2.675 $X2=0 $Y2=0
cc_52 N_KAPWR_c_63_n N_VPWR_c_93_n 0.00346901f $X=1.705 $Y=2.81 $X2=0 $Y2=0
