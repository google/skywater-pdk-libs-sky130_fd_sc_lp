* File: sky130_fd_sc_lp__o32ai_1.pxi.spice
* Created: Fri Aug 28 11:18:12 2020
* 
x_PM_SKY130_FD_SC_LP__O32AI_1%B1 N_B1_c_51_n N_B1_M1009_g N_B1_M1004_g B1 B1 B1
+ N_B1_c_54_n N_B1_c_55_n PM_SKY130_FD_SC_LP__O32AI_1%B1
x_PM_SKY130_FD_SC_LP__O32AI_1%B2 N_B2_M1005_g N_B2_M1001_g B2 N_B2_c_86_n
+ N_B2_c_87_n PM_SKY130_FD_SC_LP__O32AI_1%B2
x_PM_SKY130_FD_SC_LP__O32AI_1%A3 N_A3_c_121_n N_A3_M1003_g N_A3_M1006_g A3 A3
+ N_A3_c_124_n PM_SKY130_FD_SC_LP__O32AI_1%A3
x_PM_SKY130_FD_SC_LP__O32AI_1%A2 N_A2_M1008_g N_A2_M1007_g A2 A2 N_A2_c_158_n
+ N_A2_c_159_n PM_SKY130_FD_SC_LP__O32AI_1%A2
x_PM_SKY130_FD_SC_LP__O32AI_1%A1 N_A1_M1000_g N_A1_M1002_g A1 A1 N_A1_c_189_n
+ N_A1_c_190_n PM_SKY130_FD_SC_LP__O32AI_1%A1
x_PM_SKY130_FD_SC_LP__O32AI_1%VPWR N_VPWR_M1004_s N_VPWR_M1000_d N_VPWR_c_212_n
+ N_VPWR_c_213_n N_VPWR_c_214_n N_VPWR_c_215_n N_VPWR_c_216_n VPWR
+ N_VPWR_c_217_n N_VPWR_c_211_n PM_SKY130_FD_SC_LP__O32AI_1%VPWR
x_PM_SKY130_FD_SC_LP__O32AI_1%Y N_Y_M1009_d N_Y_M1005_d N_Y_c_247_n N_Y_c_249_n
+ N_Y_c_250_n Y Y Y N_Y_c_251_n N_Y_c_245_n PM_SKY130_FD_SC_LP__O32AI_1%Y
x_PM_SKY130_FD_SC_LP__O32AI_1%A_76_69# N_A_76_69#_M1009_s N_A_76_69#_M1001_d
+ N_A_76_69#_M1007_d N_A_76_69#_c_277_n N_A_76_69#_c_282_n N_A_76_69#_c_292_n
+ N_A_76_69#_c_288_n N_A_76_69#_c_278_n N_A_76_69#_c_279_n
+ PM_SKY130_FD_SC_LP__O32AI_1%A_76_69#
x_PM_SKY130_FD_SC_LP__O32AI_1%VGND N_VGND_M1003_d N_VGND_M1002_d N_VGND_c_311_n
+ N_VGND_c_312_n VGND N_VGND_c_313_n N_VGND_c_314_n N_VGND_c_315_n
+ N_VGND_c_316_n PM_SKY130_FD_SC_LP__O32AI_1%VGND
cc_1 VNB N_B1_c_51_n 0.0189529f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.295
cc_2 VNB N_B1_M1004_g 0.00137264f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=2.465
cc_3 VNB B1 0.0200157f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_4 VNB N_B1_c_54_n 0.0485687f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.46
cc_5 VNB N_B1_c_55_n 0.0228236f $X=-0.19 $Y=-0.245 $X2=0.345 $Y2=1.195
cc_6 VNB N_B2_M1001_g 0.0200763f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_7 VNB N_B2_c_86_n 0.0266472f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_8 VNB N_B2_c_87_n 0.00386581f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_9 VNB N_A3_c_121_n 0.0188352f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.295
cc_10 VNB N_A3_M1006_g 0.00160058f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=2.465
cc_11 VNB A3 0.00208646f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_12 VNB N_A3_c_124_n 0.041201f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A2_M1008_g 0.00128301f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=0.765
cc_14 VNB A2 0.0105774f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_15 VNB N_A2_c_158_n 0.0285598f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A2_c_159_n 0.0182254f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A1_M1000_g 0.00164097f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=0.765
cc_18 VNB A1 0.0216162f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=0.84
cc_19 VNB N_A1_c_189_n 0.0449371f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A1_c_190_n 0.0203953f $X=-0.19 $Y=-0.245 $X2=0.5 $Y2=1.46
cc_21 VNB N_VPWR_c_211_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_Y_c_245_n 0.00296951f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_76_69#_c_277_n 0.00552299f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.58
cc_24 VNB N_A_76_69#_c_278_n 0.00189378f $X=-0.19 $Y=-0.245 $X2=0.345 $Y2=1.195
cc_25 VNB N_A_76_69#_c_279_n 0.0182282f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_311_n 0.0123161f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_312_n 0.0352805f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_28 VNB N_VGND_c_313_n 0.0444649f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_314_n 0.0146445f $X=-0.19 $Y=-0.245 $X2=0.345 $Y2=1.295
cc_30 VNB N_VGND_c_315_n 0.0173479f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_316_n 0.205322f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VPB N_B1_M1004_g 0.0236801f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=2.465
cc_33 VPB B1 0.0173951f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_34 VPB N_B2_M1005_g 0.0213558f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=0.765
cc_35 VPB N_B2_c_86_n 0.00748735f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_36 VPB N_B2_c_87_n 0.00306913f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_37 VPB N_A3_M1006_g 0.0235463f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=2.465
cc_38 VPB A3 0.00306492f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_39 VPB N_A2_M1008_g 0.0190044f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=0.765
cc_40 VPB A2 0.0247136f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_41 VPB N_A1_M1000_g 0.0249906f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=0.765
cc_42 VPB A1 0.00985898f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=0.84
cc_43 VPB N_VPWR_c_212_n 0.049566f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_44 VPB N_VPWR_c_213_n 0.0124132f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_45 VPB N_VPWR_c_214_n 0.0484529f $X=-0.19 $Y=1.655 $X2=0.5 $Y2=1.46
cc_46 VPB N_VPWR_c_215_n 0.0129628f $X=-0.19 $Y=1.655 $X2=0.345 $Y2=1.195
cc_47 VPB N_VPWR_c_216_n 0.00506799f $X=-0.19 $Y=1.655 $X2=0.345 $Y2=1.295
cc_48 VPB N_VPWR_c_217_n 0.060314f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_49 VPB N_VPWR_c_211_n 0.0567957f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_50 VPB N_Y_c_245_n 0.00132336f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_51 N_B1_M1004_g N_B2_M1005_g 0.059861f $X=0.72 $Y=2.465 $X2=0 $Y2=0
cc_52 N_B1_c_51_n N_B2_M1001_g 0.016585f $X=0.72 $Y=1.295 $X2=0 $Y2=0
cc_53 N_B1_c_54_n N_B2_c_86_n 0.059861f $X=0.72 $Y=1.46 $X2=0 $Y2=0
cc_54 N_B1_c_54_n N_B2_c_87_n 3.21864e-19 $X=0.72 $Y=1.46 $X2=0 $Y2=0
cc_55 N_B1_M1004_g N_VPWR_c_212_n 0.00629315f $X=0.72 $Y=2.465 $X2=0 $Y2=0
cc_56 B1 N_VPWR_c_212_n 0.0235248f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_57 N_B1_c_54_n N_VPWR_c_212_n 0.00149269f $X=0.72 $Y=1.46 $X2=0 $Y2=0
cc_58 N_B1_M1004_g N_VPWR_c_217_n 0.0055654f $X=0.72 $Y=2.465 $X2=0 $Y2=0
cc_59 N_B1_M1004_g N_VPWR_c_211_n 0.0109365f $X=0.72 $Y=2.465 $X2=0 $Y2=0
cc_60 N_B1_c_51_n N_Y_c_247_n 0.00495263f $X=0.72 $Y=1.295 $X2=0 $Y2=0
cc_61 N_B1_c_55_n N_Y_c_247_n 0.0101927f $X=0.345 $Y=1.195 $X2=0 $Y2=0
cc_62 N_B1_c_51_n N_Y_c_249_n 0.0052446f $X=0.72 $Y=1.295 $X2=0 $Y2=0
cc_63 N_B1_c_51_n N_Y_c_250_n 0.00166585f $X=0.72 $Y=1.295 $X2=0 $Y2=0
cc_64 N_B1_M1004_g N_Y_c_251_n 0.0225239f $X=0.72 $Y=2.465 $X2=0 $Y2=0
cc_65 N_B1_c_51_n N_Y_c_245_n 0.0023327f $X=0.72 $Y=1.295 $X2=0 $Y2=0
cc_66 N_B1_M1004_g N_Y_c_245_n 0.0101853f $X=0.72 $Y=2.465 $X2=0 $Y2=0
cc_67 B1 N_Y_c_245_n 0.0422387f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_68 N_B1_c_54_n N_Y_c_245_n 0.00710996f $X=0.72 $Y=1.46 $X2=0 $Y2=0
cc_69 N_B1_c_55_n N_A_76_69#_M1009_s 0.00543656f $X=0.345 $Y=1.195 $X2=-0.19
+ $Y2=-0.245
cc_70 N_B1_c_51_n N_A_76_69#_c_277_n 0.0126331f $X=0.72 $Y=1.295 $X2=0 $Y2=0
cc_71 N_B1_c_51_n N_A_76_69#_c_282_n 3.57705e-19 $X=0.72 $Y=1.295 $X2=0 $Y2=0
cc_72 N_B1_c_51_n N_A_76_69#_c_279_n 8.76125e-19 $X=0.72 $Y=1.295 $X2=0 $Y2=0
cc_73 N_B1_c_54_n N_A_76_69#_c_279_n 7.6976e-19 $X=0.72 $Y=1.46 $X2=0 $Y2=0
cc_74 N_B1_c_55_n N_A_76_69#_c_279_n 0.0210749f $X=0.345 $Y=1.195 $X2=0 $Y2=0
cc_75 N_B1_c_51_n N_VGND_c_313_n 0.0029147f $X=0.72 $Y=1.295 $X2=0 $Y2=0
cc_76 N_B1_c_51_n N_VGND_c_316_n 0.00427198f $X=0.72 $Y=1.295 $X2=0 $Y2=0
cc_77 N_B1_c_55_n N_VGND_c_316_n 0.010607f $X=0.345 $Y=1.195 $X2=0 $Y2=0
cc_78 N_B2_M1001_g N_A3_c_121_n 0.0165842f $X=1.2 $Y=0.765 $X2=-0.19 $Y2=-0.245
cc_79 N_B2_M1005_g N_A3_M1006_g 0.00624545f $X=1.08 $Y=2.465 $X2=0 $Y2=0
cc_80 N_B2_c_86_n N_A3_M1006_g 0.0010262f $X=1.2 $Y=1.51 $X2=0 $Y2=0
cc_81 N_B2_c_87_n N_A3_M1006_g 2.95113e-19 $X=1.2 $Y=1.51 $X2=0 $Y2=0
cc_82 N_B2_M1001_g A3 5.57523e-19 $X=1.2 $Y=0.765 $X2=0 $Y2=0
cc_83 N_B2_c_86_n A3 4.85602e-19 $X=1.2 $Y=1.51 $X2=0 $Y2=0
cc_84 N_B2_c_87_n A3 0.0319362f $X=1.2 $Y=1.51 $X2=0 $Y2=0
cc_85 N_B2_c_86_n N_A3_c_124_n 0.0177979f $X=1.2 $Y=1.51 $X2=0 $Y2=0
cc_86 N_B2_c_87_n N_A3_c_124_n 0.00164345f $X=1.2 $Y=1.51 $X2=0 $Y2=0
cc_87 N_B2_M1005_g N_VPWR_c_217_n 0.00357668f $X=1.08 $Y=2.465 $X2=0 $Y2=0
cc_88 N_B2_M1005_g N_VPWR_c_211_n 0.00591024f $X=1.08 $Y=2.465 $X2=0 $Y2=0
cc_89 N_B2_c_86_n N_Y_c_250_n 0.0037249f $X=1.2 $Y=1.51 $X2=0 $Y2=0
cc_90 N_B2_M1005_g N_Y_c_251_n 0.037261f $X=1.08 $Y=2.465 $X2=0 $Y2=0
cc_91 N_B2_c_86_n N_Y_c_251_n 0.00121006f $X=1.2 $Y=1.51 $X2=0 $Y2=0
cc_92 N_B2_c_87_n N_Y_c_251_n 0.0234644f $X=1.2 $Y=1.51 $X2=0 $Y2=0
cc_93 N_B2_M1001_g N_Y_c_245_n 0.00126081f $X=1.2 $Y=0.765 $X2=0 $Y2=0
cc_94 N_B2_c_86_n N_Y_c_245_n 0.0053805f $X=1.2 $Y=1.51 $X2=0 $Y2=0
cc_95 N_B2_c_87_n N_Y_c_245_n 0.0301772f $X=1.2 $Y=1.51 $X2=0 $Y2=0
cc_96 N_B2_M1001_g N_A_76_69#_c_277_n 0.0127128f $X=1.2 $Y=0.765 $X2=0 $Y2=0
cc_97 N_B2_M1001_g N_A_76_69#_c_282_n 0.00553904f $X=1.2 $Y=0.765 $X2=0 $Y2=0
cc_98 N_B2_M1001_g N_A_76_69#_c_288_n 0.00150521f $X=1.2 $Y=0.765 $X2=0 $Y2=0
cc_99 N_B2_c_86_n N_A_76_69#_c_288_n 4.34637e-19 $X=1.2 $Y=1.51 $X2=0 $Y2=0
cc_100 N_B2_c_87_n N_A_76_69#_c_288_n 0.00623054f $X=1.2 $Y=1.51 $X2=0 $Y2=0
cc_101 N_B2_M1001_g N_VGND_c_313_n 0.00291465f $X=1.2 $Y=0.765 $X2=0 $Y2=0
cc_102 N_B2_M1001_g N_VGND_c_315_n 4.43722e-19 $X=1.2 $Y=0.765 $X2=0 $Y2=0
cc_103 N_B2_M1001_g N_VGND_c_316_n 0.00403581f $X=1.2 $Y=0.765 $X2=0 $Y2=0
cc_104 N_A3_M1006_g N_A2_M1008_g 0.0678238f $X=1.92 $Y=2.465 $X2=0 $Y2=0
cc_105 N_A3_c_121_n A2 2.91721e-19 $X=1.65 $Y=1.295 $X2=0 $Y2=0
cc_106 A3 A2 0.0453016f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_107 N_A3_c_124_n A2 0.00631952f $X=1.92 $Y=1.46 $X2=0 $Y2=0
cc_108 A3 N_A2_c_158_n 2.47184e-19 $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_109 N_A3_c_124_n N_A2_c_158_n 0.0207142f $X=1.92 $Y=1.46 $X2=0 $Y2=0
cc_110 N_A3_c_121_n N_A2_c_159_n 0.0119266f $X=1.65 $Y=1.295 $X2=0 $Y2=0
cc_111 N_A3_M1006_g N_VPWR_c_217_n 0.0054895f $X=1.92 $Y=2.465 $X2=0 $Y2=0
cc_112 N_A3_M1006_g N_VPWR_c_211_n 0.0108264f $X=1.92 $Y=2.465 $X2=0 $Y2=0
cc_113 N_A3_M1006_g N_Y_c_251_n 0.0272279f $X=1.92 $Y=2.465 $X2=0 $Y2=0
cc_114 A3 N_Y_c_251_n 0.022365f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_115 N_A3_c_124_n N_Y_c_251_n 0.00182826f $X=1.92 $Y=1.46 $X2=0 $Y2=0
cc_116 A3 N_Y_c_245_n 0.00320935f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_117 N_A3_c_121_n N_A_76_69#_c_277_n 7.62582e-19 $X=1.65 $Y=1.295 $X2=0 $Y2=0
cc_118 N_A3_c_121_n N_A_76_69#_c_292_n 0.0136505f $X=1.65 $Y=1.295 $X2=0 $Y2=0
cc_119 A3 N_A_76_69#_c_292_n 0.0196414f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_120 N_A3_c_124_n N_A_76_69#_c_292_n 0.0056402f $X=1.92 $Y=1.46 $X2=0 $Y2=0
cc_121 N_A3_c_121_n N_VGND_c_313_n 0.00401871f $X=1.65 $Y=1.295 $X2=0 $Y2=0
cc_122 N_A3_c_121_n N_VGND_c_315_n 0.00941994f $X=1.65 $Y=1.295 $X2=0 $Y2=0
cc_123 N_A3_c_121_n N_VGND_c_316_n 0.00776189f $X=1.65 $Y=1.295 $X2=0 $Y2=0
cc_124 N_A2_M1008_g N_A1_M1000_g 0.0677657f $X=2.37 $Y=2.465 $X2=0 $Y2=0
cc_125 A2 A1 0.0444132f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_126 N_A2_c_158_n A1 2.31618e-19 $X=2.37 $Y=1.46 $X2=0 $Y2=0
cc_127 A2 N_A1_c_189_n 0.00664122f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_128 N_A2_c_158_n N_A1_c_189_n 0.0206643f $X=2.37 $Y=1.46 $X2=0 $Y2=0
cc_129 A2 N_A1_c_190_n 6.9571e-19 $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_130 N_A2_c_159_n N_A1_c_190_n 0.0159226f $X=2.37 $Y=1.295 $X2=0 $Y2=0
cc_131 N_A2_M1008_g N_VPWR_c_214_n 0.00668369f $X=2.37 $Y=2.465 $X2=0 $Y2=0
cc_132 N_A2_M1008_g N_VPWR_c_217_n 0.00585385f $X=2.37 $Y=2.465 $X2=0 $Y2=0
cc_133 N_A2_M1008_g N_VPWR_c_211_n 0.0111381f $X=2.37 $Y=2.465 $X2=0 $Y2=0
cc_134 N_A2_M1008_g N_Y_c_251_n 0.00552505f $X=2.37 $Y=2.465 $X2=0 $Y2=0
cc_135 A2 N_A_76_69#_c_292_n 0.0527067f $X=2.555 $Y=1.21 $X2=0 $Y2=0
cc_136 N_A2_c_158_n N_A_76_69#_c_292_n 6.80933e-19 $X=2.37 $Y=1.46 $X2=0 $Y2=0
cc_137 N_A2_c_159_n N_A_76_69#_c_292_n 0.0133695f $X=2.37 $Y=1.295 $X2=0 $Y2=0
cc_138 N_A2_c_159_n N_VGND_c_312_n 4.8783e-19 $X=2.37 $Y=1.295 $X2=0 $Y2=0
cc_139 N_A2_c_159_n N_VGND_c_314_n 0.00401871f $X=2.37 $Y=1.295 $X2=0 $Y2=0
cc_140 N_A2_c_159_n N_VGND_c_315_n 0.00964305f $X=2.37 $Y=1.295 $X2=0 $Y2=0
cc_141 N_A2_c_159_n N_VGND_c_316_n 0.00775088f $X=2.37 $Y=1.295 $X2=0 $Y2=0
cc_142 N_A1_M1000_g N_VPWR_c_214_n 0.0322194f $X=2.82 $Y=2.465 $X2=0 $Y2=0
cc_143 A1 N_VPWR_c_214_n 0.0244629f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_144 N_A1_c_189_n N_VPWR_c_214_n 0.00133856f $X=2.99 $Y=1.46 $X2=0 $Y2=0
cc_145 N_A1_M1000_g N_VPWR_c_217_n 0.00486043f $X=2.82 $Y=2.465 $X2=0 $Y2=0
cc_146 N_A1_M1000_g N_VPWR_c_211_n 0.00843372f $X=2.82 $Y=2.465 $X2=0 $Y2=0
cc_147 A1 N_VGND_c_312_n 0.026499f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_148 N_A1_c_189_n N_VGND_c_312_n 0.00131759f $X=2.99 $Y=1.46 $X2=0 $Y2=0
cc_149 N_A1_c_190_n N_VGND_c_312_n 0.0141188f $X=2.95 $Y=1.295 $X2=0 $Y2=0
cc_150 N_A1_c_190_n N_VGND_c_314_n 0.00400407f $X=2.95 $Y=1.295 $X2=0 $Y2=0
cc_151 N_A1_c_190_n N_VGND_c_315_n 4.40139e-19 $X=2.95 $Y=1.295 $X2=0 $Y2=0
cc_152 N_A1_c_190_n N_VGND_c_316_n 0.00775088f $X=2.95 $Y=1.295 $X2=0 $Y2=0
cc_153 N_VPWR_c_211_n A_159_367# 0.00168875f $X=3.12 $Y=3.33 $X2=-0.19
+ $Y2=-0.245
cc_154 N_VPWR_c_211_n N_Y_M1005_d 0.00564363f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_155 N_VPWR_c_217_n N_Y_c_251_n 0.0684316f $X=2.87 $Y=3.33 $X2=0 $Y2=0
cc_156 N_VPWR_c_211_n N_Y_c_251_n 0.0414639f $X=3.12 $Y=3.33 $X2=0 $Y2=0
cc_157 N_VPWR_c_211_n A_399_367# 0.0128488f $X=3.12 $Y=3.33 $X2=-0.19 $Y2=-0.245
cc_158 N_VPWR_c_211_n A_489_367# 0.0128488f $X=3.12 $Y=3.33 $X2=-0.19 $Y2=-0.245
cc_159 A_159_367# N_Y_c_251_n 8.99573e-19 $X=0.795 $Y=1.835 $X2=0.72 $Y2=3.33
cc_160 A_159_367# N_Y_c_245_n 3.84994e-19 $X=0.795 $Y=1.835 $X2=0.72 $Y2=3.33
cc_161 N_Y_M1009_d N_A_76_69#_c_277_n 0.00229612f $X=0.795 $Y=0.345 $X2=0 $Y2=0
cc_162 N_Y_c_249_n N_A_76_69#_c_277_n 0.0179996f $X=0.935 $Y=0.72 $X2=0 $Y2=0
cc_163 N_A_76_69#_c_292_n N_VGND_M1003_d 0.0141787f $X=2.54 $Y=0.955 $X2=-0.19
+ $Y2=-0.245
cc_164 N_A_76_69#_c_278_n N_VGND_c_312_n 0.0211767f $X=2.635 $Y=0.49 $X2=0 $Y2=0
cc_165 N_A_76_69#_c_277_n N_VGND_c_313_n 0.0608963f $X=1.27 $Y=0.34 $X2=0 $Y2=0
cc_166 N_A_76_69#_c_279_n N_VGND_c_313_n 0.0178268f $X=0.47 $Y=0.34 $X2=0 $Y2=0
cc_167 N_A_76_69#_c_278_n N_VGND_c_314_n 0.00935612f $X=2.635 $Y=0.49 $X2=0
+ $Y2=0
cc_168 N_A_76_69#_c_277_n N_VGND_c_315_n 0.0112909f $X=1.27 $Y=0.34 $X2=0 $Y2=0
cc_169 N_A_76_69#_c_292_n N_VGND_c_315_n 0.0447396f $X=2.54 $Y=0.955 $X2=0 $Y2=0
cc_170 N_A_76_69#_c_278_n N_VGND_c_315_n 0.0164064f $X=2.635 $Y=0.49 $X2=0 $Y2=0
cc_171 N_A_76_69#_c_277_n N_VGND_c_316_n 0.03393f $X=1.27 $Y=0.34 $X2=0 $Y2=0
cc_172 N_A_76_69#_c_278_n N_VGND_c_316_n 0.00705762f $X=2.635 $Y=0.49 $X2=0
+ $Y2=0
cc_173 N_A_76_69#_c_279_n N_VGND_c_316_n 0.00990565f $X=0.47 $Y=0.34 $X2=0 $Y2=0
