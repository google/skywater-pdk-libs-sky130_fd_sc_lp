* File: sky130_fd_sc_lp__a211oi_lp.pxi.spice
* Created: Wed Sep  2 09:18:22 2020
* 
x_PM_SKY130_FD_SC_LP__A211OI_LP%C1 N_C1_c_62_n N_C1_M1008_g N_C1_c_63_n
+ N_C1_M1004_g N_C1_c_64_n N_C1_c_65_n N_C1_M1005_g N_C1_c_66_n N_C1_c_72_n C1
+ C1 C1 C1 C1 N_C1_c_68_n N_C1_c_69_n PM_SKY130_FD_SC_LP__A211OI_LP%C1
x_PM_SKY130_FD_SC_LP__A211OI_LP%B1 N_B1_M1002_g N_B1_c_111_n N_B1_M1000_g
+ N_B1_c_112_n N_B1_c_113_n N_B1_M1001_g N_B1_c_114_n N_B1_c_115_n N_B1_c_121_n
+ N_B1_c_116_n B1 B1 N_B1_c_118_n PM_SKY130_FD_SC_LP__A211OI_LP%B1
x_PM_SKY130_FD_SC_LP__A211OI_LP%A1 N_A1_M1007_g N_A1_M1003_g A1 A1 N_A1_c_168_n
+ PM_SKY130_FD_SC_LP__A211OI_LP%A1
x_PM_SKY130_FD_SC_LP__A211OI_LP%A2 N_A2_M1009_g N_A2_M1006_g N_A2_c_204_n
+ N_A2_c_205_n A2 A2 N_A2_c_207_n PM_SKY130_FD_SC_LP__A211OI_LP%A2
x_PM_SKY130_FD_SC_LP__A211OI_LP%Y N_Y_M1008_s N_Y_M1001_d N_Y_M1004_s
+ N_Y_c_233_n N_Y_c_234_n Y Y Y Y Y Y Y N_Y_c_236_n
+ PM_SKY130_FD_SC_LP__A211OI_LP%Y
x_PM_SKY130_FD_SC_LP__A211OI_LP%A_279_409# N_A_279_409#_M1002_d
+ N_A_279_409#_M1006_d N_A_279_409#_c_276_n N_A_279_409#_c_277_n
+ N_A_279_409#_c_278_n N_A_279_409#_c_279_n
+ PM_SKY130_FD_SC_LP__A211OI_LP%A_279_409#
x_PM_SKY130_FD_SC_LP__A211OI_LP%VPWR N_VPWR_M1007_d N_VPWR_c_304_n VPWR
+ N_VPWR_c_305_n N_VPWR_c_306_n N_VPWR_c_303_n N_VPWR_c_308_n
+ PM_SKY130_FD_SC_LP__A211OI_LP%VPWR
x_PM_SKY130_FD_SC_LP__A211OI_LP%VGND N_VGND_M1005_d N_VGND_M1009_d
+ N_VGND_c_332_n N_VGND_c_333_n N_VGND_c_334_n N_VGND_c_335_n VGND
+ N_VGND_c_336_n N_VGND_c_337_n N_VGND_c_338_n N_VGND_c_339_n
+ PM_SKY130_FD_SC_LP__A211OI_LP%VGND
cc_1 VNB N_C1_c_62_n 0.0175316f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=0.78
cc_2 VNB N_C1_c_63_n 0.0234643f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.665
cc_3 VNB N_C1_c_64_n 0.015517f $X=-0.19 $Y=-0.245 $X2=0.895 $Y2=0.855
cc_4 VNB N_C1_c_65_n 0.0138901f $X=-0.19 $Y=-0.245 $X2=0.97 $Y2=0.78
cc_5 VNB N_C1_c_66_n 0.00664349f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=0.855
cc_6 VNB C1 0.0014486f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_7 VNB N_C1_c_68_n 0.0176432f $X=-0.19 $Y=-0.245 $X2=0.74 $Y2=1.345
cc_8 VNB N_C1_c_69_n 0.0123438f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.18
cc_9 VNB N_B1_c_111_n 0.0138901f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=1.18
cc_10 VNB N_B1_c_112_n 0.0168137f $X=-0.19 $Y=-0.245 $X2=0.78 $Y2=2.545
cc_11 VNB N_B1_c_113_n 0.0137713f $X=-0.19 $Y=-0.245 $X2=0.895 $Y2=0.855
cc_12 VNB N_B1_c_114_n 0.019498f $X=-0.19 $Y=-0.245 $X2=0.97 $Y2=0.495
cc_13 VNB N_B1_c_115_n 0.0185722f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=0.855
cc_14 VNB N_B1_c_116_n 0.0046532f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_15 VNB B1 0.00548263f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=2.32
cc_16 VNB N_B1_c_118_n 0.0144744f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.345
cc_17 VNB N_A1_M1003_g 0.0370782f $X=-0.19 $Y=-0.245 $X2=0.72 $Y2=1.665
cc_18 VNB A1 0.00291361f $X=-0.19 $Y=-0.245 $X2=0.78 $Y2=2.545
cc_19 VNB N_A1_c_168_n 0.0557381f $X=-0.19 $Y=-0.245 $X2=0.97 $Y2=0.78
cc_20 VNB N_A2_M1009_g 0.0454835f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=0.495
cc_21 VNB N_A2_c_204_n 0.025421f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A2_c_205_n 0.0030084f $X=-0.19 $Y=-0.245 $X2=0.895 $Y2=0.855
cc_23 VNB A2 0.0419629f $X=-0.19 $Y=-0.245 $X2=0.97 $Y2=0.495
cc_24 VNB N_A2_c_207_n 0.0179334f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=2.32
cc_25 VNB N_Y_c_233_n 0.017378f $X=-0.19 $Y=-0.245 $X2=0.78 $Y2=2.545
cc_26 VNB N_Y_c_234_n 0.00207453f $X=-0.19 $Y=-0.245 $X2=0.97 $Y2=0.78
cc_27 VNB Y 0.0493142f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=0.855
cc_28 VNB N_Y_c_236_n 0.0274483f $X=-0.19 $Y=-0.245 $X2=0.74 $Y2=1.295
cc_29 VNB N_VPWR_c_303_n 0.143779f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.95
cc_30 VNB N_VGND_c_332_n 0.00177638f $X=-0.19 $Y=-0.245 $X2=0.78 $Y2=2.545
cc_31 VNB N_VGND_c_333_n 0.0254175f $X=-0.19 $Y=-0.245 $X2=0.685 $Y2=0.855
cc_32 VNB N_VGND_c_334_n 0.0374802f $X=-0.19 $Y=-0.245 $X2=0.97 $Y2=0.495
cc_33 VNB N_VGND_c_335_n 0.00551342f $X=-0.19 $Y=-0.245 $X2=0.61 $Y2=0.855
cc_34 VNB N_VGND_c_336_n 0.0298894f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.58
cc_35 VNB N_VGND_c_337_n 0.0135992f $X=-0.19 $Y=-0.245 $X2=0.74 $Y2=1.295
cc_36 VNB N_VGND_c_338_n 0.221366f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_339_n 0.00500486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_38 VPB N_C1_c_63_n 7.30721e-19 $X=-0.19 $Y=1.655 $X2=0.72 $Y2=1.665
cc_39 VPB N_C1_M1004_g 0.0323872f $X=-0.19 $Y=1.655 $X2=0.78 $Y2=2.545
cc_40 VPB N_C1_c_72_n 0.0195432f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=1.85
cc_41 VPB C1 0.00184745f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_42 VPB N_B1_M1002_g 0.0292636f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=0.495
cc_43 VPB N_B1_c_115_n 0.00110618f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=0.855
cc_44 VPB N_B1_c_121_n 0.0121223f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=1.85
cc_45 VPB B1 0.00589141f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=2.32
cc_46 VPB N_A1_M1007_g 0.0319297f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=0.495
cc_47 VPB A1 0.00313998f $X=-0.19 $Y=1.655 $X2=0.78 $Y2=2.545
cc_48 VPB N_A1_c_168_n 0.0266134f $X=-0.19 $Y=1.655 $X2=0.97 $Y2=0.78
cc_49 VPB N_A2_M1006_g 0.0460636f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=1.665
cc_50 VPB N_A2_c_205_n 0.0115327f $X=-0.19 $Y=1.655 $X2=0.895 $Y2=0.855
cc_51 VPB A2 0.0148479f $X=-0.19 $Y=1.655 $X2=0.97 $Y2=0.495
cc_52 VPB Y 0.0614261f $X=-0.19 $Y=1.655 $X2=0.61 $Y2=0.855
cc_53 VPB N_A_279_409#_c_276_n 0.00252852f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_54 VPB N_A_279_409#_c_277_n 0.0202269f $X=-0.19 $Y=1.655 $X2=0.685 $Y2=0.855
cc_55 VPB N_A_279_409#_c_278_n 0.00302988f $X=-0.19 $Y=1.655 $X2=0.97 $Y2=0.78
cc_56 VPB N_A_279_409#_c_279_n 0.035517f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_57 VPB N_VPWR_c_304_n 0.00426397f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=1.365
cc_58 VPB N_VPWR_c_305_n 0.0555019f $X=-0.19 $Y=1.655 $X2=0.78 $Y2=2.545
cc_59 VPB N_VPWR_c_306_n 0.0338033f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.58
cc_60 VPB N_VPWR_c_303_n 0.0880073f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.95
cc_61 VPB N_VPWR_c_308_n 0.00548753f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_62 N_C1_M1004_g N_B1_M1002_g 0.0269527f $X=0.78 $Y=2.545 $X2=0 $Y2=0
cc_63 N_C1_c_65_n N_B1_c_111_n 0.0100676f $X=0.97 $Y=0.78 $X2=0 $Y2=0
cc_64 N_C1_c_69_n N_B1_c_114_n 0.00165818f $X=0.72 $Y=1.18 $X2=0 $Y2=0
cc_65 N_C1_c_63_n N_B1_c_115_n 0.0269527f $X=0.72 $Y=1.665 $X2=0 $Y2=0
cc_66 N_C1_c_72_n N_B1_c_121_n 0.0269527f $X=0.72 $Y=1.85 $X2=0 $Y2=0
cc_67 C1 N_B1_c_121_n 0.00477186f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_68 N_C1_c_64_n N_B1_c_116_n 0.0100676f $X=0.895 $Y=0.855 $X2=0 $Y2=0
cc_69 C1 B1 0.0533544f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_70 N_C1_c_68_n B1 0.00437424f $X=0.74 $Y=1.345 $X2=0 $Y2=0
cc_71 C1 N_B1_c_118_n 7.42321e-19 $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_72 N_C1_c_68_n N_B1_c_118_n 0.0269527f $X=0.74 $Y=1.345 $X2=0 $Y2=0
cc_73 C1 N_Y_M1004_s 0.0097188f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_74 N_C1_c_64_n N_Y_c_233_n 0.0160347f $X=0.895 $Y=0.855 $X2=0 $Y2=0
cc_75 N_C1_c_66_n N_Y_c_233_n 0.00411533f $X=0.61 $Y=0.855 $X2=0 $Y2=0
cc_76 C1 N_Y_c_233_n 0.0236752f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_77 N_C1_c_68_n N_Y_c_233_n 6.80799e-19 $X=0.74 $Y=1.345 $X2=0 $Y2=0
cc_78 N_C1_c_69_n N_Y_c_233_n 0.00291688f $X=0.72 $Y=1.18 $X2=0 $Y2=0
cc_79 N_C1_M1004_g Y 0.0122402f $X=0.78 $Y=2.545 $X2=0 $Y2=0
cc_80 N_C1_c_66_n Y 0.00263592f $X=0.61 $Y=0.855 $X2=0 $Y2=0
cc_81 C1 Y 0.129279f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_82 N_C1_c_69_n Y 0.0268276f $X=0.72 $Y=1.18 $X2=0 $Y2=0
cc_83 N_C1_c_62_n N_Y_c_236_n 0.0113199f $X=0.61 $Y=0.78 $X2=0 $Y2=0
cc_84 N_C1_c_65_n N_Y_c_236_n 0.00171265f $X=0.97 $Y=0.78 $X2=0 $Y2=0
cc_85 N_C1_c_66_n N_Y_c_236_n 0.00273554f $X=0.61 $Y=0.855 $X2=0 $Y2=0
cc_86 C1 N_A_279_409#_c_278_n 0.00314529f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_87 N_C1_M1004_g N_VPWR_c_305_n 0.00596257f $X=0.78 $Y=2.545 $X2=0 $Y2=0
cc_88 C1 N_VPWR_c_305_n 0.00914393f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_89 N_C1_M1004_g N_VPWR_c_303_n 0.0083872f $X=0.78 $Y=2.545 $X2=0 $Y2=0
cc_90 C1 N_VPWR_c_303_n 0.0101955f $X=0.635 $Y=1.21 $X2=0 $Y2=0
cc_91 N_C1_c_62_n N_VGND_c_332_n 0.00188065f $X=0.61 $Y=0.78 $X2=0 $Y2=0
cc_92 N_C1_c_65_n N_VGND_c_332_n 0.0105659f $X=0.97 $Y=0.78 $X2=0 $Y2=0
cc_93 N_C1_c_62_n N_VGND_c_336_n 0.00502664f $X=0.61 $Y=0.78 $X2=0 $Y2=0
cc_94 N_C1_c_64_n N_VGND_c_336_n 4.57848e-19 $X=0.895 $Y=0.855 $X2=0 $Y2=0
cc_95 N_C1_c_65_n N_VGND_c_336_n 0.00445056f $X=0.97 $Y=0.78 $X2=0 $Y2=0
cc_96 N_C1_c_62_n N_VGND_c_338_n 0.00632776f $X=0.61 $Y=0.78 $X2=0 $Y2=0
cc_97 N_C1_c_64_n N_VGND_c_338_n 6.33118e-19 $X=0.895 $Y=0.855 $X2=0 $Y2=0
cc_98 N_C1_c_65_n N_VGND_c_338_n 0.00418511f $X=0.97 $Y=0.78 $X2=0 $Y2=0
cc_99 N_B1_M1002_g N_A1_M1007_g 0.0151052f $X=1.27 $Y=2.545 $X2=0 $Y2=0
cc_100 N_B1_c_113_n N_A1_M1003_g 0.0179557f $X=1.76 $Y=0.78 $X2=0 $Y2=0
cc_101 N_B1_c_114_n N_A1_M1003_g 0.00494915f $X=1.31 $Y=1.17 $X2=0 $Y2=0
cc_102 B1 A1 0.0510971f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_103 N_B1_c_118_n A1 3.57249e-19 $X=1.31 $Y=1.335 $X2=0 $Y2=0
cc_104 N_B1_c_112_n N_A1_c_168_n 0.00674899f $X=1.685 $Y=0.855 $X2=0 $Y2=0
cc_105 B1 N_A1_c_168_n 0.0235289f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_106 N_B1_c_118_n N_A1_c_168_n 0.0369353f $X=1.31 $Y=1.335 $X2=0 $Y2=0
cc_107 N_B1_c_112_n N_Y_c_233_n 0.0167163f $X=1.685 $Y=0.855 $X2=0 $Y2=0
cc_108 N_B1_c_114_n N_Y_c_233_n 0.00548496f $X=1.31 $Y=1.17 $X2=0 $Y2=0
cc_109 N_B1_c_116_n N_Y_c_233_n 0.00606062f $X=1.4 $Y=0.855 $X2=0 $Y2=0
cc_110 B1 N_Y_c_233_n 0.0548262f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_111 N_B1_c_118_n N_Y_c_233_n 0.00471135f $X=1.31 $Y=1.335 $X2=0 $Y2=0
cc_112 N_B1_c_111_n N_Y_c_234_n 0.00171786f $X=1.4 $Y=0.78 $X2=0 $Y2=0
cc_113 N_B1_c_112_n N_Y_c_234_n 0.00230187f $X=1.685 $Y=0.855 $X2=0 $Y2=0
cc_114 N_B1_c_113_n N_Y_c_234_n 0.0100195f $X=1.76 $Y=0.78 $X2=0 $Y2=0
cc_115 N_B1_M1002_g N_A_279_409#_c_276_n 5.70164e-19 $X=1.27 $Y=2.545 $X2=0
+ $Y2=0
cc_116 B1 N_A_279_409#_c_277_n 0.00394469f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_117 N_B1_M1002_g N_A_279_409#_c_278_n 4.02415e-19 $X=1.27 $Y=2.545 $X2=0
+ $Y2=0
cc_118 N_B1_c_121_n N_A_279_409#_c_278_n 0.00176037f $X=1.31 $Y=1.84 $X2=0 $Y2=0
cc_119 B1 N_A_279_409#_c_278_n 0.0290018f $X=1.595 $Y=1.21 $X2=0 $Y2=0
cc_120 N_B1_M1002_g N_VPWR_c_304_n 7.97642e-19 $X=1.27 $Y=2.545 $X2=0 $Y2=0
cc_121 N_B1_M1002_g N_VPWR_c_305_n 0.00893366f $X=1.27 $Y=2.545 $X2=0 $Y2=0
cc_122 N_B1_M1002_g N_VPWR_c_303_n 0.016682f $X=1.27 $Y=2.545 $X2=0 $Y2=0
cc_123 N_B1_c_111_n N_VGND_c_332_n 0.0105659f $X=1.4 $Y=0.78 $X2=0 $Y2=0
cc_124 N_B1_c_113_n N_VGND_c_332_n 0.00188065f $X=1.76 $Y=0.78 $X2=0 $Y2=0
cc_125 N_B1_c_111_n N_VGND_c_334_n 0.00445056f $X=1.4 $Y=0.78 $X2=0 $Y2=0
cc_126 N_B1_c_112_n N_VGND_c_334_n 4.57848e-19 $X=1.685 $Y=0.855 $X2=0 $Y2=0
cc_127 N_B1_c_113_n N_VGND_c_334_n 0.00502664f $X=1.76 $Y=0.78 $X2=0 $Y2=0
cc_128 N_B1_c_111_n N_VGND_c_338_n 0.00418511f $X=1.4 $Y=0.78 $X2=0 $Y2=0
cc_129 N_B1_c_112_n N_VGND_c_338_n 6.33118e-19 $X=1.685 $Y=0.855 $X2=0 $Y2=0
cc_130 N_B1_c_113_n N_VGND_c_338_n 0.00562693f $X=1.76 $Y=0.78 $X2=0 $Y2=0
cc_131 N_A1_M1003_g N_A2_M1009_g 0.04468f $X=2.19 $Y=0.495 $X2=0 $Y2=0
cc_132 N_A1_M1007_g N_A2_M1006_g 0.0189503f $X=1.84 $Y=2.545 $X2=0 $Y2=0
cc_133 A1 N_A2_c_205_n 4.11727e-19 $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_134 N_A1_M1003_g A2 0.00145529f $X=2.19 $Y=0.495 $X2=0 $Y2=0
cc_135 A1 A2 0.042501f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_136 N_A1_c_168_n A2 0.00432632f $X=2.14 $Y=1.335 $X2=0 $Y2=0
cc_137 A1 N_A2_c_207_n 7.4777e-19 $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_138 N_A1_c_168_n N_A2_c_207_n 0.0374383f $X=2.14 $Y=1.335 $X2=0 $Y2=0
cc_139 N_A1_M1003_g N_Y_c_233_n 0.0062265f $X=2.19 $Y=0.495 $X2=0 $Y2=0
cc_140 A1 N_Y_c_233_n 0.0138709f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_141 N_A1_c_168_n N_Y_c_233_n 0.00933439f $X=2.14 $Y=1.335 $X2=0 $Y2=0
cc_142 N_A1_M1003_g N_Y_c_234_n 0.0118604f $X=2.19 $Y=0.495 $X2=0 $Y2=0
cc_143 N_A1_M1007_g N_A_279_409#_c_276_n 0.0205472f $X=1.84 $Y=2.545 $X2=0 $Y2=0
cc_144 N_A1_M1007_g N_A_279_409#_c_277_n 0.0242264f $X=1.84 $Y=2.545 $X2=0 $Y2=0
cc_145 A1 N_A_279_409#_c_277_n 0.0250673f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_146 N_A1_c_168_n N_A_279_409#_c_277_n 0.00270263f $X=2.14 $Y=1.335 $X2=0
+ $Y2=0
cc_147 N_A1_M1007_g N_A_279_409#_c_278_n 0.00103317f $X=1.84 $Y=2.545 $X2=0
+ $Y2=0
cc_148 N_A1_M1007_g N_VPWR_c_304_n 0.0170232f $X=1.84 $Y=2.545 $X2=0 $Y2=0
cc_149 N_A1_M1007_g N_VPWR_c_305_n 0.00769046f $X=1.84 $Y=2.545 $X2=0 $Y2=0
cc_150 N_A1_M1007_g N_VPWR_c_303_n 0.0135127f $X=1.84 $Y=2.545 $X2=0 $Y2=0
cc_151 N_A1_M1003_g N_VGND_c_333_n 0.00214576f $X=2.19 $Y=0.495 $X2=0 $Y2=0
cc_152 N_A1_M1003_g N_VGND_c_334_n 0.00502664f $X=2.19 $Y=0.495 $X2=0 $Y2=0
cc_153 N_A1_M1003_g N_VGND_c_338_n 0.00957379f $X=2.19 $Y=0.495 $X2=0 $Y2=0
cc_154 N_A2_M1009_g N_Y_c_233_n 8.21499e-19 $X=2.62 $Y=0.495 $X2=0 $Y2=0
cc_155 N_A2_M1009_g N_Y_c_234_n 0.00181469f $X=2.62 $Y=0.495 $X2=0 $Y2=0
cc_156 N_A2_M1006_g N_A_279_409#_c_277_n 0.021661f $X=2.67 $Y=2.545 $X2=0 $Y2=0
cc_157 N_A2_c_205_n N_A_279_409#_c_277_n 0.00205805f $X=2.71 $Y=1.78 $X2=0 $Y2=0
cc_158 A2 N_A_279_409#_c_277_n 0.0377589f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_159 N_A2_M1006_g N_A_279_409#_c_279_n 0.0231404f $X=2.67 $Y=2.545 $X2=0 $Y2=0
cc_160 N_A2_M1006_g N_VPWR_c_304_n 0.00971804f $X=2.67 $Y=2.545 $X2=0 $Y2=0
cc_161 N_A2_M1006_g N_VPWR_c_306_n 0.0086001f $X=2.67 $Y=2.545 $X2=0 $Y2=0
cc_162 N_A2_M1006_g N_VPWR_c_303_n 0.0168995f $X=2.67 $Y=2.545 $X2=0 $Y2=0
cc_163 N_A2_M1009_g N_VGND_c_333_n 0.0149784f $X=2.62 $Y=0.495 $X2=0 $Y2=0
cc_164 A2 N_VGND_c_333_n 0.0162621f $X=3.035 $Y=1.21 $X2=0 $Y2=0
cc_165 N_A2_c_207_n N_VGND_c_333_n 0.00421165f $X=2.71 $Y=1.275 $X2=0 $Y2=0
cc_166 N_A2_M1009_g N_VGND_c_334_n 0.00445056f $X=2.62 $Y=0.495 $X2=0 $Y2=0
cc_167 N_A2_M1009_g N_VGND_c_338_n 0.0081158f $X=2.62 $Y=0.495 $X2=0 $Y2=0
cc_168 Y N_VPWR_c_305_n 0.0180698f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_169 Y N_VPWR_c_303_n 0.0103698f $X=0.155 $Y=0.84 $X2=0 $Y2=0
cc_170 N_Y_c_233_n N_VGND_c_332_n 0.0199879f $X=1.81 $Y=0.905 $X2=0 $Y2=0
cc_171 N_Y_c_234_n N_VGND_c_332_n 0.0125465f $X=1.975 $Y=0.495 $X2=0 $Y2=0
cc_172 N_Y_c_236_n N_VGND_c_332_n 0.0128173f $X=0.395 $Y=0.495 $X2=0 $Y2=0
cc_173 N_Y_c_234_n N_VGND_c_333_n 0.013602f $X=1.975 $Y=0.495 $X2=0 $Y2=0
cc_174 N_Y_c_234_n N_VGND_c_334_n 0.021949f $X=1.975 $Y=0.495 $X2=0 $Y2=0
cc_175 N_Y_c_236_n N_VGND_c_336_n 0.0291117f $X=0.395 $Y=0.495 $X2=0 $Y2=0
cc_176 N_Y_c_233_n N_VGND_c_338_n 0.0284029f $X=1.81 $Y=0.905 $X2=0 $Y2=0
cc_177 N_Y_c_234_n N_VGND_c_338_n 0.0124703f $X=1.975 $Y=0.495 $X2=0 $Y2=0
cc_178 N_Y_c_236_n N_VGND_c_338_n 0.0166436f $X=0.395 $Y=0.495 $X2=0 $Y2=0
cc_179 N_A_279_409#_c_277_n N_VPWR_M1007_d 0.012799f $X=2.77 $Y=2.105 $X2=-0.19
+ $Y2=1.655
cc_180 N_A_279_409#_c_276_n N_VPWR_c_304_n 0.045794f $X=1.575 $Y=2.9 $X2=0 $Y2=0
cc_181 N_A_279_409#_c_277_n N_VPWR_c_304_n 0.0209601f $X=2.77 $Y=2.105 $X2=0
+ $Y2=0
cc_182 N_A_279_409#_c_279_n N_VPWR_c_304_n 0.0233678f $X=2.935 $Y=2.9 $X2=0
+ $Y2=0
cc_183 N_A_279_409#_c_276_n N_VPWR_c_305_n 0.0220321f $X=1.575 $Y=2.9 $X2=0
+ $Y2=0
cc_184 N_A_279_409#_c_279_n N_VPWR_c_306_n 0.0220321f $X=2.935 $Y=2.9 $X2=0
+ $Y2=0
cc_185 N_A_279_409#_c_276_n N_VPWR_c_303_n 0.0125808f $X=1.575 $Y=2.9 $X2=0
+ $Y2=0
cc_186 N_A_279_409#_c_279_n N_VPWR_c_303_n 0.0125808f $X=2.935 $Y=2.9 $X2=0
+ $Y2=0
