* File: sky130_fd_sc_lp__a31o_4.pxi.spice
* Created: Fri Aug 28 09:59:19 2020
* 
x_PM_SKY130_FD_SC_LP__A31O_4%B1 N_B1_M1009_g N_B1_M1011_g N_B1_c_115_n
+ N_B1_M1016_g N_B1_M1022_g N_B1_c_118_n B1 B1 N_B1_c_120_n
+ PM_SKY130_FD_SC_LP__A31O_4%B1
x_PM_SKY130_FD_SC_LP__A31O_4%A_110_47# N_A_110_47#_M1009_d N_A_110_47#_M1002_s
+ N_A_110_47#_M1011_s N_A_110_47#_M1003_g N_A_110_47#_c_159_n
+ N_A_110_47#_c_160_n N_A_110_47#_M1014_g N_A_110_47#_c_170_n
+ N_A_110_47#_M1004_g N_A_110_47#_M1021_g N_A_110_47#_c_171_n
+ N_A_110_47#_M1008_g N_A_110_47#_M1023_g N_A_110_47#_c_172_n
+ N_A_110_47#_M1012_g N_A_110_47#_c_164_n N_A_110_47#_c_165_n
+ N_A_110_47#_c_175_n N_A_110_47#_M1017_g N_A_110_47#_c_295_p
+ N_A_110_47#_c_166_n N_A_110_47#_c_186_n N_A_110_47#_c_167_n
+ N_A_110_47#_c_190_p N_A_110_47#_c_168_n N_A_110_47#_c_212_p
+ N_A_110_47#_c_187_n N_A_110_47#_c_169_n PM_SKY130_FD_SC_LP__A31O_4%A_110_47#
x_PM_SKY130_FD_SC_LP__A31O_4%A3 N_A3_c_325_n N_A3_M1010_g N_A3_c_326_n
+ N_A3_c_327_n N_A3_c_328_n N_A3_M1020_g N_A3_M1006_g N_A3_c_329_n N_A3_M1015_g
+ N_A3_c_330_n N_A3_c_331_n A3 A3 A3 N_A3_c_333_n PM_SKY130_FD_SC_LP__A31O_4%A3
x_PM_SKY130_FD_SC_LP__A31O_4%A2 N_A2_M1000_g N_A2_M1001_g N_A2_M1005_g
+ N_A2_M1013_g A2 A2 N_A2_c_403_n PM_SKY130_FD_SC_LP__A31O_4%A2
x_PM_SKY130_FD_SC_LP__A31O_4%A1 N_A1_M1002_g N_A1_M1007_g N_A1_M1018_g
+ N_A1_M1019_g A1 A1 N_A1_c_452_n PM_SKY130_FD_SC_LP__A31O_4%A1
x_PM_SKY130_FD_SC_LP__A31O_4%A_27_367# N_A_27_367#_M1011_d N_A_27_367#_M1022_d
+ N_A_27_367#_M1006_s N_A_27_367#_M1001_d N_A_27_367#_M1007_d
+ N_A_27_367#_c_490_n N_A_27_367#_c_491_n N_A_27_367#_c_500_n
+ N_A_27_367#_c_564_p N_A_27_367#_c_492_n N_A_27_367#_c_493_n
+ N_A_27_367#_c_508_n N_A_27_367#_c_509_n N_A_27_367#_c_537_p
+ N_A_27_367#_c_515_n N_A_27_367#_c_547_p N_A_27_367#_c_520_n
+ N_A_27_367#_c_525_n N_A_27_367#_c_548_p N_A_27_367#_c_494_n
+ N_A_27_367#_c_517_n N_A_27_367#_c_522_n PM_SKY130_FD_SC_LP__A31O_4%A_27_367#
x_PM_SKY130_FD_SC_LP__A31O_4%VPWR N_VPWR_M1004_d N_VPWR_M1008_d N_VPWR_M1017_d
+ N_VPWR_M1015_d N_VPWR_M1013_s N_VPWR_M1019_s N_VPWR_c_572_n N_VPWR_c_573_n
+ N_VPWR_c_574_n N_VPWR_c_575_n N_VPWR_c_576_n N_VPWR_c_577_n N_VPWR_c_578_n
+ N_VPWR_c_579_n N_VPWR_c_580_n N_VPWR_c_581_n N_VPWR_c_582_n N_VPWR_c_583_n
+ VPWR N_VPWR_c_584_n N_VPWR_c_585_n N_VPWR_c_586_n N_VPWR_c_587_n
+ N_VPWR_c_588_n N_VPWR_c_589_n N_VPWR_c_571_n PM_SKY130_FD_SC_LP__A31O_4%VPWR
x_PM_SKY130_FD_SC_LP__A31O_4%X N_X_M1003_s N_X_M1021_s N_X_M1004_s N_X_M1012_s
+ N_X_c_678_n N_X_c_676_n N_X_c_679_n N_X_c_680_n X X N_X_c_677_n
+ PM_SKY130_FD_SC_LP__A31O_4%X
x_PM_SKY130_FD_SC_LP__A31O_4%VGND N_VGND_M1009_s N_VGND_M1016_s N_VGND_M1014_d
+ N_VGND_M1023_d N_VGND_M1020_s N_VGND_c_734_n N_VGND_c_735_n N_VGND_c_736_n
+ N_VGND_c_737_n N_VGND_c_738_n N_VGND_c_739_n N_VGND_c_740_n N_VGND_c_741_n
+ N_VGND_c_742_n VGND N_VGND_c_743_n N_VGND_c_744_n N_VGND_c_745_n
+ N_VGND_c_746_n N_VGND_c_747_n N_VGND_c_748_n N_VGND_c_749_n
+ PM_SKY130_FD_SC_LP__A31O_4%VGND
x_PM_SKY130_FD_SC_LP__A31O_4%A_726_47# N_A_726_47#_M1010_d N_A_726_47#_M1000_d
+ N_A_726_47#_c_827_n N_A_726_47#_c_829_n N_A_726_47#_c_825_n
+ PM_SKY130_FD_SC_LP__A31O_4%A_726_47#
x_PM_SKY130_FD_SC_LP__A31O_4%A_919_67# N_A_919_67#_M1000_s N_A_919_67#_M1005_s
+ N_A_919_67#_M1018_d N_A_919_67#_c_856_n N_A_919_67#_c_857_n
+ N_A_919_67#_c_858_n N_A_919_67#_c_859_n PM_SKY130_FD_SC_LP__A31O_4%A_919_67#
cc_1 VNB N_B1_M1009_g 0.0231841f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.655
cc_2 VNB N_B1_M1011_g 0.00703468f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.465
cc_3 VNB N_B1_c_115_n 0.0101534f $X=-0.19 $Y=-0.245 $X2=0.83 $Y2=1.465
cc_4 VNB N_B1_M1016_g 0.0255362f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=0.655
cc_5 VNB N_B1_M1022_g 0.00575006f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=2.465
cc_6 VNB N_B1_c_118_n 0.00573352f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=1.465
cc_7 VNB B1 0.0184601f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_8 VNB N_B1_c_120_n 0.0385106f $X=-0.19 $Y=-0.245 $X2=0.34 $Y2=1.375
cc_9 VNB N_A_110_47#_M1003_g 0.0233043f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=0.655
cc_10 VNB N_A_110_47#_c_159_n 0.0297949f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_11 VNB N_A_110_47#_c_160_n 0.00866399f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=1.54
cc_12 VNB N_A_110_47#_M1014_g 0.0244014f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_13 VNB N_A_110_47#_M1021_g 0.0240767f $X=-0.19 $Y=-0.245 $X2=0.34 $Y2=1.375
cc_14 VNB N_A_110_47#_M1023_g 0.0251293f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_15 VNB N_A_110_47#_c_164_n 0.012891f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_16 VNB N_A_110_47#_c_165_n 0.0841486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_17 VNB N_A_110_47#_c_166_n 0.00322617f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_110_47#_c_167_n 0.00177966f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_110_47#_c_168_n 0.0385431f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_110_47#_c_169_n 0.00385932f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A3_c_325_n 0.0160329f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.21
cc_22 VNB N_A3_c_326_n 0.0134225f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A3_c_327_n 0.00805594f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=1.54
cc_24 VNB N_A3_c_328_n 0.019573f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=2.465
cc_25 VNB N_A3_c_329_n 0.0154028f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=0.655
cc_26 VNB N_A3_c_330_n 0.0146228f $X=-0.19 $Y=-0.245 $X2=0.155 $Y2=1.21
cc_27 VNB N_A3_c_331_n 0.00653098f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_28 VNB A3 0.00914451f $X=-0.19 $Y=-0.245 $X2=0.34 $Y2=1.375
cc_29 VNB N_A3_c_333_n 0.016564f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.295
cc_30 VNB N_A2_M1000_g 0.0228894f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.655
cc_31 VNB N_A2_M1005_g 0.019078f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=1.39
cc_32 VNB A2 0.00311942f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_A2_c_403_n 0.0342918f $X=-0.19 $Y=-0.245 $X2=0.34 $Y2=1.375
cc_34 VNB N_A1_M1002_g 0.0190738f $X=-0.19 $Y=-0.245 $X2=0.475 $Y2=0.655
cc_35 VNB N_A1_M1018_g 0.0262521f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=1.39
cc_36 VNB A1 0.0140046f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_37 VNB N_A1_c_452_n 0.0381849f $X=-0.19 $Y=-0.245 $X2=0.34 $Y2=1.375
cc_38 VNB N_VPWR_c_571_n 0.283096f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_39 VNB N_X_c_676_n 0.00689008f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=2.465
cc_40 VNB N_X_c_677_n 0.0075139f $X=-0.19 $Y=-0.245 $X2=0.29 $Y2=1.295
cc_41 VNB N_VGND_c_734_n 0.0103657f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=2.465
cc_42 VNB N_VGND_c_735_n 0.0352483f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_736_n 3.99129e-19 $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_737_n 4.89148e-19 $X=-0.19 $Y=-0.245 $X2=0.34 $Y2=1.375
cc_45 VNB N_VGND_c_738_n 0.0175644f $X=-0.19 $Y=-0.245 $X2=0.362 $Y2=1.465
cc_46 VNB N_VGND_c_739_n 0.002833f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_740_n 0.00487815f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_741_n 0.0183475f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_742_n 0.0038195f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_743_n 0.0121755f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_744_n 0.0186597f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_745_n 0.0594796f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_746_n 0.341179f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_747_n 0.00436154f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_748_n 0.00436154f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_56 VNB N_VGND_c_749_n 0.00510127f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_57 VNB N_A_726_47#_c_825_n 0.00762068f $X=-0.19 $Y=-0.245 $X2=0.905 $Y2=0.655
cc_58 VNB N_A_919_67#_c_856_n 0.0120369f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_59 VNB N_A_919_67#_c_857_n 0.0329098f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_60 VNB N_A_919_67#_c_858_n 0.00780954f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_61 VNB N_A_919_67#_c_859_n 0.00134511f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_62 VPB N_B1_M1011_g 0.0258006f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.465
cc_63 VPB N_B1_M1022_g 0.022786f $X=-0.19 $Y=1.655 $X2=0.905 $Y2=2.465
cc_64 VPB B1 0.00619129f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_65 VPB N_A_110_47#_c_170_n 0.01931f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.21
cc_66 VPB N_A_110_47#_c_171_n 0.0160061f $X=-0.19 $Y=1.655 $X2=0.362 $Y2=1.21
cc_67 VPB N_A_110_47#_c_172_n 0.0160022f $X=-0.19 $Y=1.655 $X2=0.29 $Y2=1.665
cc_68 VPB N_A_110_47#_c_164_n 0.00632517f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_69 VPB N_A_110_47#_c_165_n 0.015268f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_70 VPB N_A_110_47#_c_175_n 0.0159713f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_71 VPB N_A_110_47#_c_166_n 0.00151325f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_72 VPB N_A3_M1006_g 0.0180996f $X=-0.19 $Y=1.655 $X2=0.905 $Y2=1.39
cc_73 VPB N_A3_c_329_n 0.00323474f $X=-0.19 $Y=1.655 $X2=0.905 $Y2=0.655
cc_74 VPB N_A3_M1015_g 0.0185396f $X=-0.19 $Y=1.655 $X2=0.905 $Y2=2.465
cc_75 VPB N_A3_c_331_n 0.00347253f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_76 VPB A3 0.0152608f $X=-0.19 $Y=1.655 $X2=0.34 $Y2=1.375
cc_77 VPB N_A2_M1001_g 0.0188979f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.465
cc_78 VPB N_A2_M1013_g 0.0179997f $X=-0.19 $Y=1.655 $X2=0.905 $Y2=1.54
cc_79 VPB A2 0.00471908f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_80 VPB N_A2_c_403_n 0.00478023f $X=-0.19 $Y=1.655 $X2=0.34 $Y2=1.375
cc_81 VPB N_A1_M1007_g 0.0187774f $X=-0.19 $Y=1.655 $X2=0.475 $Y2=2.465
cc_82 VPB N_A1_M1019_g 0.0233606f $X=-0.19 $Y=1.655 $X2=0.905 $Y2=1.54
cc_83 VPB A1 0.0109779f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_84 VPB N_A1_c_452_n 0.00505343f $X=-0.19 $Y=1.655 $X2=0.34 $Y2=1.375
cc_85 VPB N_A_27_367#_c_490_n 0.00746637f $X=-0.19 $Y=1.655 $X2=0.905 $Y2=2.465
cc_86 VPB N_A_27_367#_c_491_n 0.0392929f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_87 VPB N_A_27_367#_c_492_n 0.0121352f $X=-0.19 $Y=1.655 $X2=0.362 $Y2=1.21
cc_88 VPB N_A_27_367#_c_493_n 0.0238301f $X=-0.19 $Y=1.655 $X2=0.362 $Y2=1.465
cc_89 VPB N_A_27_367#_c_494_n 9.49157e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_90 VPB N_VPWR_c_572_n 0.00910925f $X=-0.19 $Y=1.655 $X2=0.155 $Y2=1.58
cc_91 VPB N_VPWR_c_573_n 3.0911e-19 $X=-0.19 $Y=1.655 $X2=0.34 $Y2=1.375
cc_92 VPB N_VPWR_c_574_n 3.12649e-19 $X=-0.19 $Y=1.655 $X2=0.362 $Y2=1.54
cc_93 VPB N_VPWR_c_575_n 0.0127409f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_94 VPB N_VPWR_c_576_n 3.16188e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_95 VPB N_VPWR_c_577_n 3.12649e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_96 VPB N_VPWR_c_578_n 0.0103398f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_97 VPB N_VPWR_c_579_n 0.0491987f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_98 VPB N_VPWR_c_580_n 0.0127282f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_99 VPB N_VPWR_c_581_n 0.00436638f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_100 VPB N_VPWR_c_582_n 0.0127282f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_101 VPB N_VPWR_c_583_n 0.00436638f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_102 VPB N_VPWR_c_584_n 0.050367f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_103 VPB N_VPWR_c_585_n 0.0133881f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_104 VPB N_VPWR_c_586_n 0.0129398f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_105 VPB N_VPWR_c_587_n 0.00510611f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_106 VPB N_VPWR_c_588_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_107 VPB N_VPWR_c_589_n 0.00436868f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_108 VPB N_VPWR_c_571_n 0.0534145f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_109 VPB N_X_c_678_n 0.00601497f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_110 VPB N_X_c_679_n 0.00852289f $X=-0.19 $Y=1.655 $X2=0.905 $Y2=1.465
cc_111 VPB N_X_c_680_n 0.0100566f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_112 VPB N_X_c_677_n 0.0125685f $X=-0.19 $Y=1.655 $X2=0.29 $Y2=1.295
cc_113 N_B1_M1016_g N_A_110_47#_M1003_g 0.0224594f $X=0.905 $Y=0.655 $X2=0 $Y2=0
cc_114 N_B1_c_118_n N_A_110_47#_c_160_n 0.0224594f $X=0.905 $Y=1.465 $X2=0 $Y2=0
cc_115 N_B1_M1009_g N_A_110_47#_c_166_n 0.00509388f $X=0.475 $Y=0.655 $X2=0
+ $Y2=0
cc_116 N_B1_M1011_g N_A_110_47#_c_166_n 0.00443321f $X=0.475 $Y=2.465 $X2=0
+ $Y2=0
cc_117 N_B1_c_115_n N_A_110_47#_c_166_n 0.0102007f $X=0.83 $Y=1.465 $X2=0 $Y2=0
cc_118 N_B1_M1016_g N_A_110_47#_c_166_n 0.0102699f $X=0.905 $Y=0.655 $X2=0 $Y2=0
cc_119 N_B1_M1022_g N_A_110_47#_c_166_n 0.0192235f $X=0.905 $Y=2.465 $X2=0 $Y2=0
cc_120 N_B1_c_118_n N_A_110_47#_c_166_n 0.00157093f $X=0.905 $Y=1.465 $X2=0
+ $Y2=0
cc_121 B1 N_A_110_47#_c_166_n 0.0414547f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_122 N_B1_M1016_g N_A_110_47#_c_186_n 0.0119928f $X=0.905 $Y=0.655 $X2=0 $Y2=0
cc_123 N_B1_M1016_g N_A_110_47#_c_187_n 0.0012826f $X=0.905 $Y=0.655 $X2=0 $Y2=0
cc_124 N_B1_M1011_g N_A_27_367#_c_490_n 5.81207e-19 $X=0.475 $Y=2.465 $X2=0
+ $Y2=0
cc_125 N_B1_M1011_g N_A_27_367#_c_491_n 0.0123113f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_126 N_B1_M1022_g N_A_27_367#_c_491_n 7.67708e-19 $X=0.905 $Y=2.465 $X2=0
+ $Y2=0
cc_127 B1 N_A_27_367#_c_491_n 0.0214593f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_128 N_B1_c_120_n N_A_27_367#_c_491_n 9.66246e-19 $X=0.34 $Y=1.375 $X2=0 $Y2=0
cc_129 N_B1_M1011_g N_A_27_367#_c_500_n 0.0105205f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_130 N_B1_M1022_g N_A_27_367#_c_500_n 0.0115031f $X=0.905 $Y=2.465 $X2=0 $Y2=0
cc_131 N_B1_M1011_g N_VPWR_c_584_n 0.00357842f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_132 N_B1_M1022_g N_VPWR_c_584_n 0.00357877f $X=0.905 $Y=2.465 $X2=0 $Y2=0
cc_133 N_B1_M1011_g N_VPWR_c_571_n 0.00628379f $X=0.475 $Y=2.465 $X2=0 $Y2=0
cc_134 N_B1_M1022_g N_VPWR_c_571_n 0.00665089f $X=0.905 $Y=2.465 $X2=0 $Y2=0
cc_135 N_B1_M1022_g N_X_c_678_n 0.00254286f $X=0.905 $Y=2.465 $X2=0 $Y2=0
cc_136 N_B1_M1016_g N_X_c_677_n 0.011214f $X=0.905 $Y=0.655 $X2=0 $Y2=0
cc_137 N_B1_M1009_g N_VGND_c_735_n 0.0154209f $X=0.475 $Y=0.655 $X2=0 $Y2=0
cc_138 N_B1_M1016_g N_VGND_c_735_n 6.87633e-19 $X=0.905 $Y=0.655 $X2=0 $Y2=0
cc_139 B1 N_VGND_c_735_n 0.0204697f $X=0.155 $Y=1.21 $X2=0 $Y2=0
cc_140 N_B1_c_120_n N_VGND_c_735_n 0.00160808f $X=0.34 $Y=1.375 $X2=0 $Y2=0
cc_141 N_B1_M1009_g N_VGND_c_736_n 5.09333e-19 $X=0.475 $Y=0.655 $X2=0 $Y2=0
cc_142 N_B1_M1016_g N_VGND_c_736_n 0.00639943f $X=0.905 $Y=0.655 $X2=0 $Y2=0
cc_143 N_B1_M1009_g N_VGND_c_743_n 0.00486043f $X=0.475 $Y=0.655 $X2=0 $Y2=0
cc_144 N_B1_M1016_g N_VGND_c_743_n 0.00353512f $X=0.905 $Y=0.655 $X2=0 $Y2=0
cc_145 N_B1_M1009_g N_VGND_c_746_n 0.00824727f $X=0.475 $Y=0.655 $X2=0 $Y2=0
cc_146 N_B1_M1016_g N_VGND_c_746_n 0.00411673f $X=0.905 $Y=0.655 $X2=0 $Y2=0
cc_147 N_A_110_47#_M1023_g N_A3_c_325_n 0.032573f $X=3.045 $Y=0.655 $X2=-0.19
+ $Y2=-0.245
cc_148 N_A_110_47#_c_186_n N_A3_c_325_n 0.00152893f $X=3.08 $Y=0.72 $X2=-0.19
+ $Y2=-0.245
cc_149 N_A_110_47#_c_190_p N_A3_c_325_n 0.00414508f $X=3.165 $Y=1.075 $X2=-0.19
+ $Y2=-0.245
cc_150 N_A_110_47#_c_168_n N_A3_c_325_n 0.00986262f $X=5.865 $Y=1.16 $X2=-0.19
+ $Y2=-0.245
cc_151 N_A_110_47#_c_168_n N_A3_c_326_n 0.0052475f $X=5.865 $Y=1.16 $X2=0 $Y2=0
cc_152 N_A_110_47#_c_164_n N_A3_c_327_n 0.01241f $X=3.55 $Y=1.65 $X2=0 $Y2=0
cc_153 N_A_110_47#_c_165_n N_A3_c_327_n 0.00113455f $X=3.27 $Y=1.65 $X2=0 $Y2=0
cc_154 N_A_110_47#_c_168_n N_A3_c_327_n 0.00275696f $X=5.865 $Y=1.16 $X2=0 $Y2=0
cc_155 N_A_110_47#_c_169_n N_A3_c_327_n 0.00193085f $X=3.165 $Y=1.16 $X2=0 $Y2=0
cc_156 N_A_110_47#_c_168_n N_A3_c_328_n 0.0074394f $X=5.865 $Y=1.16 $X2=0 $Y2=0
cc_157 N_A_110_47#_c_164_n N_A3_M1006_g 0.0526642f $X=3.55 $Y=1.65 $X2=0 $Y2=0
cc_158 N_A_110_47#_c_168_n N_A3_c_329_n 0.00168779f $X=5.865 $Y=1.16 $X2=0 $Y2=0
cc_159 N_A_110_47#_c_168_n N_A3_c_330_n 0.0105166f $X=5.865 $Y=1.16 $X2=0 $Y2=0
cc_160 N_A_110_47#_c_164_n N_A3_c_331_n 0.00653748f $X=3.55 $Y=1.65 $X2=0 $Y2=0
cc_161 N_A_110_47#_c_172_n A3 6.02336e-19 $X=3.195 $Y=1.725 $X2=0 $Y2=0
cc_162 N_A_110_47#_c_164_n A3 0.0107654f $X=3.55 $Y=1.65 $X2=0 $Y2=0
cc_163 N_A_110_47#_c_165_n A3 8.08604e-19 $X=3.27 $Y=1.65 $X2=0 $Y2=0
cc_164 N_A_110_47#_c_175_n A3 0.0070294f $X=3.625 $Y=1.725 $X2=0 $Y2=0
cc_165 N_A_110_47#_c_168_n A3 0.0855328f $X=5.865 $Y=1.16 $X2=0 $Y2=0
cc_166 N_A_110_47#_c_169_n A3 0.0135766f $X=3.165 $Y=1.16 $X2=0 $Y2=0
cc_167 N_A_110_47#_c_165_n N_A3_c_333_n 0.00275188f $X=3.27 $Y=1.65 $X2=0 $Y2=0
cc_168 N_A_110_47#_c_169_n N_A3_c_333_n 0.00144187f $X=3.165 $Y=1.16 $X2=0 $Y2=0
cc_169 N_A_110_47#_c_168_n N_A2_M1000_g 0.0145762f $X=5.865 $Y=1.16 $X2=0 $Y2=0
cc_170 N_A_110_47#_c_168_n N_A2_M1005_g 0.011897f $X=5.865 $Y=1.16 $X2=0 $Y2=0
cc_171 N_A_110_47#_c_212_p N_A2_M1005_g 0.00173915f $X=6.03 $Y=0.71 $X2=0 $Y2=0
cc_172 N_A_110_47#_c_168_n A2 0.0487804f $X=5.865 $Y=1.16 $X2=0 $Y2=0
cc_173 N_A_110_47#_c_168_n N_A2_c_403_n 0.00243542f $X=5.865 $Y=1.16 $X2=0 $Y2=0
cc_174 N_A_110_47#_c_168_n N_A1_M1002_g 0.0153269f $X=5.865 $Y=1.16 $X2=0 $Y2=0
cc_175 N_A_110_47#_c_212_p N_A1_M1002_g 0.00832686f $X=6.03 $Y=0.71 $X2=0 $Y2=0
cc_176 N_A_110_47#_c_168_n N_A1_M1018_g 0.00481471f $X=5.865 $Y=1.16 $X2=0 $Y2=0
cc_177 N_A_110_47#_c_212_p N_A1_M1018_g 0.0052174f $X=6.03 $Y=0.71 $X2=0 $Y2=0
cc_178 N_A_110_47#_c_168_n A1 0.0234275f $X=5.865 $Y=1.16 $X2=0 $Y2=0
cc_179 N_A_110_47#_c_168_n N_A1_c_452_n 0.00252566f $X=5.865 $Y=1.16 $X2=0 $Y2=0
cc_180 N_A_110_47#_M1011_s N_A_27_367#_c_500_n 0.00332344f $X=0.55 $Y=1.835
+ $X2=0 $Y2=0
cc_181 N_A_110_47#_c_166_n N_A_27_367#_c_500_n 0.0143076f $X=0.69 $Y=0.865 $X2=0
+ $Y2=0
cc_182 N_A_110_47#_c_170_n N_A_27_367#_c_493_n 0.0140162f $X=2.335 $Y=1.725
+ $X2=0 $Y2=0
cc_183 N_A_110_47#_c_171_n N_A_27_367#_c_493_n 0.0119756f $X=2.765 $Y=1.725
+ $X2=0 $Y2=0
cc_184 N_A_110_47#_c_172_n N_A_27_367#_c_493_n 0.0119756f $X=3.195 $Y=1.725
+ $X2=0 $Y2=0
cc_185 N_A_110_47#_c_175_n N_A_27_367#_c_493_n 0.0156956f $X=3.625 $Y=1.725
+ $X2=0 $Y2=0
cc_186 N_A_110_47#_c_175_n N_A_27_367#_c_508_n 5.00333e-19 $X=3.625 $Y=1.725
+ $X2=0 $Y2=0
cc_187 N_A_110_47#_c_175_n N_A_27_367#_c_509_n 0.00134952f $X=3.625 $Y=1.725
+ $X2=0 $Y2=0
cc_188 N_A_110_47#_c_170_n N_VPWR_c_572_n 0.0105259f $X=2.335 $Y=1.725 $X2=0
+ $Y2=0
cc_189 N_A_110_47#_c_171_n N_VPWR_c_572_n 0.00135454f $X=2.765 $Y=1.725 $X2=0
+ $Y2=0
cc_190 N_A_110_47#_c_170_n N_VPWR_c_573_n 0.00135454f $X=2.335 $Y=1.725 $X2=0
+ $Y2=0
cc_191 N_A_110_47#_c_171_n N_VPWR_c_573_n 0.0094624f $X=2.765 $Y=1.725 $X2=0
+ $Y2=0
cc_192 N_A_110_47#_c_172_n N_VPWR_c_573_n 0.0094624f $X=3.195 $Y=1.725 $X2=0
+ $Y2=0
cc_193 N_A_110_47#_c_175_n N_VPWR_c_573_n 0.00135454f $X=3.625 $Y=1.725 $X2=0
+ $Y2=0
cc_194 N_A_110_47#_c_172_n N_VPWR_c_574_n 0.00135454f $X=3.195 $Y=1.725 $X2=0
+ $Y2=0
cc_195 N_A_110_47#_c_175_n N_VPWR_c_574_n 0.00942664f $X=3.625 $Y=1.725 $X2=0
+ $Y2=0
cc_196 N_A_110_47#_c_170_n N_VPWR_c_580_n 0.0036352f $X=2.335 $Y=1.725 $X2=0
+ $Y2=0
cc_197 N_A_110_47#_c_171_n N_VPWR_c_580_n 0.0036352f $X=2.765 $Y=1.725 $X2=0
+ $Y2=0
cc_198 N_A_110_47#_c_172_n N_VPWR_c_582_n 0.0036352f $X=3.195 $Y=1.725 $X2=0
+ $Y2=0
cc_199 N_A_110_47#_c_175_n N_VPWR_c_582_n 0.0036352f $X=3.625 $Y=1.725 $X2=0
+ $Y2=0
cc_200 N_A_110_47#_M1011_s N_VPWR_c_571_n 0.00225186f $X=0.55 $Y=1.835 $X2=0
+ $Y2=0
cc_201 N_A_110_47#_c_170_n N_VPWR_c_571_n 0.00436741f $X=2.335 $Y=1.725 $X2=0
+ $Y2=0
cc_202 N_A_110_47#_c_171_n N_VPWR_c_571_n 0.00436741f $X=2.765 $Y=1.725 $X2=0
+ $Y2=0
cc_203 N_A_110_47#_c_172_n N_VPWR_c_571_n 0.00436741f $X=3.195 $Y=1.725 $X2=0
+ $Y2=0
cc_204 N_A_110_47#_c_175_n N_VPWR_c_571_n 0.00436741f $X=3.625 $Y=1.725 $X2=0
+ $Y2=0
cc_205 N_A_110_47#_c_186_n N_X_M1003_s 0.012114f $X=3.08 $Y=0.72 $X2=-0.19
+ $Y2=-0.245
cc_206 N_A_110_47#_c_186_n N_X_M1021_s 0.0107717f $X=3.08 $Y=0.72 $X2=0 $Y2=0
cc_207 N_A_110_47#_c_170_n N_X_c_678_n 0.00375462f $X=2.335 $Y=1.725 $X2=0 $Y2=0
cc_208 N_A_110_47#_c_166_n N_X_c_678_n 0.00536938f $X=0.69 $Y=0.865 $X2=0 $Y2=0
cc_209 N_A_110_47#_M1003_g N_X_c_676_n 2.33262e-19 $X=1.335 $Y=0.655 $X2=0 $Y2=0
cc_210 N_A_110_47#_c_159_n N_X_c_676_n 0.00513213f $X=1.89 $Y=1.39 $X2=0 $Y2=0
cc_211 N_A_110_47#_M1014_g N_X_c_676_n 0.0123627f $X=1.995 $Y=0.655 $X2=0 $Y2=0
cc_212 N_A_110_47#_M1021_g N_X_c_676_n 0.0127278f $X=2.425 $Y=0.655 $X2=0 $Y2=0
cc_213 N_A_110_47#_M1023_g N_X_c_676_n 0.00213977f $X=3.045 $Y=0.655 $X2=0 $Y2=0
cc_214 N_A_110_47#_c_165_n N_X_c_676_n 0.0103745f $X=3.27 $Y=1.65 $X2=0 $Y2=0
cc_215 N_A_110_47#_c_186_n N_X_c_676_n 0.071003f $X=3.08 $Y=0.72 $X2=0 $Y2=0
cc_216 N_A_110_47#_c_167_n N_X_c_676_n 0.0749102f $X=3.08 $Y=1.5 $X2=0 $Y2=0
cc_217 N_A_110_47#_c_190_p N_X_c_676_n 0.0158673f $X=3.165 $Y=1.075 $X2=0 $Y2=0
cc_218 N_A_110_47#_c_159_n N_X_c_680_n 0.00572674f $X=1.89 $Y=1.39 $X2=0 $Y2=0
cc_219 N_A_110_47#_c_170_n N_X_c_680_n 0.0174413f $X=2.335 $Y=1.725 $X2=0 $Y2=0
cc_220 N_A_110_47#_c_171_n N_X_c_680_n 0.0134574f $X=2.765 $Y=1.725 $X2=0 $Y2=0
cc_221 N_A_110_47#_c_172_n N_X_c_680_n 0.0139551f $X=3.195 $Y=1.725 $X2=0 $Y2=0
cc_222 N_A_110_47#_c_164_n N_X_c_680_n 0.0035723f $X=3.55 $Y=1.65 $X2=0 $Y2=0
cc_223 N_A_110_47#_c_165_n N_X_c_680_n 0.013974f $X=3.27 $Y=1.65 $X2=0 $Y2=0
cc_224 N_A_110_47#_c_175_n N_X_c_680_n 0.0064216f $X=3.625 $Y=1.725 $X2=0 $Y2=0
cc_225 N_A_110_47#_c_167_n N_X_c_680_n 0.0542238f $X=3.08 $Y=1.5 $X2=0 $Y2=0
cc_226 N_A_110_47#_c_169_n N_X_c_680_n 0.00788552f $X=3.165 $Y=1.16 $X2=0 $Y2=0
cc_227 N_A_110_47#_M1003_g N_X_c_677_n 0.014941f $X=1.335 $Y=0.655 $X2=0 $Y2=0
cc_228 N_A_110_47#_c_159_n N_X_c_677_n 0.0184737f $X=1.89 $Y=1.39 $X2=0 $Y2=0
cc_229 N_A_110_47#_c_160_n N_X_c_677_n 0.00653875f $X=1.41 $Y=1.39 $X2=0 $Y2=0
cc_230 N_A_110_47#_M1014_g N_X_c_677_n 0.00383664f $X=1.995 $Y=0.655 $X2=0 $Y2=0
cc_231 N_A_110_47#_c_165_n N_X_c_677_n 0.00511532f $X=3.27 $Y=1.65 $X2=0 $Y2=0
cc_232 N_A_110_47#_c_166_n N_X_c_677_n 0.0599604f $X=0.69 $Y=0.865 $X2=0 $Y2=0
cc_233 N_A_110_47#_c_186_n N_X_c_677_n 0.0429934f $X=3.08 $Y=0.72 $X2=0 $Y2=0
cc_234 N_A_110_47#_c_167_n N_X_c_677_n 0.0220704f $X=3.08 $Y=1.5 $X2=0 $Y2=0
cc_235 N_A_110_47#_c_186_n N_VGND_M1016_s 0.00346066f $X=3.08 $Y=0.72 $X2=0
+ $Y2=0
cc_236 N_A_110_47#_c_186_n N_VGND_M1014_d 0.00334936f $X=3.08 $Y=0.72 $X2=0
+ $Y2=0
cc_237 N_A_110_47#_c_186_n N_VGND_M1023_d 0.00283776f $X=3.08 $Y=0.72 $X2=0
+ $Y2=0
cc_238 N_A_110_47#_c_190_p N_VGND_M1023_d 0.00319681f $X=3.165 $Y=1.075 $X2=0
+ $Y2=0
cc_239 N_A_110_47#_M1003_g N_VGND_c_736_n 0.0100652f $X=1.335 $Y=0.655 $X2=0
+ $Y2=0
cc_240 N_A_110_47#_M1014_g N_VGND_c_736_n 0.00174006f $X=1.995 $Y=0.655 $X2=0
+ $Y2=0
cc_241 N_A_110_47#_c_186_n N_VGND_c_736_n 0.0159984f $X=3.08 $Y=0.72 $X2=0 $Y2=0
cc_242 N_A_110_47#_M1003_g N_VGND_c_737_n 0.00174006f $X=1.335 $Y=0.655 $X2=0
+ $Y2=0
cc_243 N_A_110_47#_M1014_g N_VGND_c_737_n 0.0101009f $X=1.995 $Y=0.655 $X2=0
+ $Y2=0
cc_244 N_A_110_47#_M1021_g N_VGND_c_737_n 0.00996823f $X=2.425 $Y=0.655 $X2=0
+ $Y2=0
cc_245 N_A_110_47#_M1023_g N_VGND_c_737_n 0.0018084f $X=3.045 $Y=0.655 $X2=0
+ $Y2=0
cc_246 N_A_110_47#_c_186_n N_VGND_c_737_n 0.0159984f $X=3.08 $Y=0.72 $X2=0 $Y2=0
cc_247 N_A_110_47#_M1021_g N_VGND_c_738_n 0.00353537f $X=2.425 $Y=0.655 $X2=0
+ $Y2=0
cc_248 N_A_110_47#_M1023_g N_VGND_c_738_n 0.00353523f $X=3.045 $Y=0.655 $X2=0
+ $Y2=0
cc_249 N_A_110_47#_c_186_n N_VGND_c_738_n 0.0114134f $X=3.08 $Y=0.72 $X2=0 $Y2=0
cc_250 N_A_110_47#_M1021_g N_VGND_c_739_n 0.0018084f $X=2.425 $Y=0.655 $X2=0
+ $Y2=0
cc_251 N_A_110_47#_M1023_g N_VGND_c_739_n 0.0100009f $X=3.045 $Y=0.655 $X2=0
+ $Y2=0
cc_252 N_A_110_47#_c_186_n N_VGND_c_739_n 0.00800191f $X=3.08 $Y=0.72 $X2=0
+ $Y2=0
cc_253 N_A_110_47#_c_168_n N_VGND_c_739_n 0.00558016f $X=5.865 $Y=1.16 $X2=0
+ $Y2=0
cc_254 N_A_110_47#_c_295_p N_VGND_c_743_n 0.0124525f $X=0.69 $Y=0.42 $X2=0 $Y2=0
cc_255 N_A_110_47#_c_186_n N_VGND_c_743_n 0.00161675f $X=3.08 $Y=0.72 $X2=0
+ $Y2=0
cc_256 N_A_110_47#_c_187_n N_VGND_c_743_n 8.8957e-19 $X=0.725 $Y=0.72 $X2=0
+ $Y2=0
cc_257 N_A_110_47#_M1003_g N_VGND_c_744_n 0.00353537f $X=1.335 $Y=0.655 $X2=0
+ $Y2=0
cc_258 N_A_110_47#_M1014_g N_VGND_c_744_n 0.00353537f $X=1.995 $Y=0.655 $X2=0
+ $Y2=0
cc_259 N_A_110_47#_c_186_n N_VGND_c_744_n 0.0120947f $X=3.08 $Y=0.72 $X2=0 $Y2=0
cc_260 N_A_110_47#_M1009_d N_VGND_c_746_n 0.00395019f $X=0.55 $Y=0.235 $X2=0
+ $Y2=0
cc_261 N_A_110_47#_M1003_g N_VGND_c_746_n 0.00471497f $X=1.335 $Y=0.655 $X2=0
+ $Y2=0
cc_262 N_A_110_47#_M1014_g N_VGND_c_746_n 0.00471497f $X=1.995 $Y=0.655 $X2=0
+ $Y2=0
cc_263 N_A_110_47#_M1021_g N_VGND_c_746_n 0.00463976f $X=2.425 $Y=0.655 $X2=0
+ $Y2=0
cc_264 N_A_110_47#_M1023_g N_VGND_c_746_n 0.0046395f $X=3.045 $Y=0.655 $X2=0
+ $Y2=0
cc_265 N_A_110_47#_c_295_p N_VGND_c_746_n 0.00730901f $X=0.69 $Y=0.42 $X2=0
+ $Y2=0
cc_266 N_A_110_47#_c_186_n N_VGND_c_746_n 0.0460082f $X=3.08 $Y=0.72 $X2=0 $Y2=0
cc_267 N_A_110_47#_c_187_n N_VGND_c_746_n 0.00195357f $X=0.725 $Y=0.72 $X2=0
+ $Y2=0
cc_268 N_A_110_47#_c_168_n N_A_726_47#_M1000_d 0.00176891f $X=5.865 $Y=1.16
+ $X2=0 $Y2=0
cc_269 N_A_110_47#_M1023_g N_A_726_47#_c_827_n 6.68834e-19 $X=3.045 $Y=0.655
+ $X2=0 $Y2=0
cc_270 N_A_110_47#_c_186_n N_A_726_47#_c_827_n 0.0041981f $X=3.08 $Y=0.72 $X2=0
+ $Y2=0
cc_271 N_A_110_47#_c_186_n N_A_726_47#_c_829_n 0.00395438f $X=3.08 $Y=0.72 $X2=0
+ $Y2=0
cc_272 N_A_110_47#_c_190_p N_A_726_47#_c_829_n 0.00442317f $X=3.165 $Y=1.075
+ $X2=0 $Y2=0
cc_273 N_A_110_47#_c_168_n N_A_726_47#_c_829_n 0.0214931f $X=5.865 $Y=1.16 $X2=0
+ $Y2=0
cc_274 N_A_110_47#_c_168_n N_A_726_47#_c_825_n 0.0870784f $X=5.865 $Y=1.16 $X2=0
+ $Y2=0
cc_275 N_A_110_47#_c_212_p N_A_726_47#_c_825_n 0.00558153f $X=6.03 $Y=0.71 $X2=0
+ $Y2=0
cc_276 N_A_110_47#_c_168_n N_A_919_67#_M1000_s 0.00300496f $X=5.865 $Y=1.16
+ $X2=-0.19 $Y2=-0.245
cc_277 N_A_110_47#_c_168_n N_A_919_67#_M1005_s 0.00276694f $X=5.865 $Y=1.16
+ $X2=0 $Y2=0
cc_278 N_A_110_47#_M1002_s N_A_919_67#_c_856_n 0.00176461f $X=5.89 $Y=0.335
+ $X2=0 $Y2=0
cc_279 N_A_110_47#_c_168_n N_A_919_67#_c_856_n 0.00283067f $X=5.865 $Y=1.16
+ $X2=0 $Y2=0
cc_280 N_A_110_47#_c_212_p N_A_919_67#_c_856_n 0.0159538f $X=6.03 $Y=0.71 $X2=0
+ $Y2=0
cc_281 N_A_110_47#_c_168_n N_A_919_67#_c_857_n 0.00582057f $X=5.865 $Y=1.16
+ $X2=0 $Y2=0
cc_282 N_A_110_47#_c_168_n N_A_919_67#_c_858_n 0.00351715f $X=5.865 $Y=1.16
+ $X2=0 $Y2=0
cc_283 N_A_110_47#_c_168_n N_A_919_67#_c_859_n 0.00645913f $X=5.865 $Y=1.16
+ $X2=0 $Y2=0
cc_284 N_A3_c_330_n N_A2_M1000_g 0.00334472f $X=4.075 $Y=1.26 $X2=0 $Y2=0
cc_285 N_A3_M1015_g N_A2_M1001_g 0.0187538f $X=4.485 $Y=2.465 $X2=0 $Y2=0
cc_286 N_A3_c_329_n A2 2.25164e-19 $X=4.41 $Y=1.6 $X2=0 $Y2=0
cc_287 A3 A2 0.0188276f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_288 N_A3_c_329_n N_A2_c_403_n 0.0187538f $X=4.41 $Y=1.6 $X2=0 $Y2=0
cc_289 A3 N_A2_c_403_n 0.00334573f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_290 N_A3_c_333_n N_A2_c_403_n 0.00334472f $X=4.075 $Y=1.51 $X2=0 $Y2=0
cc_291 N_A3_M1006_g N_A_27_367#_c_493_n 0.0122259f $X=4.055 $Y=2.465 $X2=0 $Y2=0
cc_292 N_A3_M1006_g N_A_27_367#_c_508_n 0.0033152f $X=4.055 $Y=2.465 $X2=0 $Y2=0
cc_293 N_A3_c_331_n N_A_27_367#_c_508_n 6.53457e-19 $X=4.075 $Y=1.6 $X2=0 $Y2=0
cc_294 A3 N_A_27_367#_c_508_n 0.0192671f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_295 N_A3_M1006_g N_A_27_367#_c_509_n 0.00652183f $X=4.055 $Y=2.465 $X2=0
+ $Y2=0
cc_296 N_A3_M1015_g N_A_27_367#_c_515_n 0.013056f $X=4.485 $Y=2.465 $X2=0 $Y2=0
cc_297 A3 N_A_27_367#_c_515_n 0.0155956f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_298 N_A3_M1006_g N_A_27_367#_c_517_n 9.88294e-19 $X=4.055 $Y=2.465 $X2=0
+ $Y2=0
cc_299 N_A3_M1006_g N_VPWR_c_574_n 0.0073068f $X=4.055 $Y=2.465 $X2=0 $Y2=0
cc_300 N_A3_M1015_g N_VPWR_c_574_n 5.41544e-19 $X=4.485 $Y=2.465 $X2=0 $Y2=0
cc_301 N_A3_M1006_g N_VPWR_c_575_n 0.00363497f $X=4.055 $Y=2.465 $X2=0 $Y2=0
cc_302 N_A3_M1015_g N_VPWR_c_575_n 0.00564095f $X=4.485 $Y=2.465 $X2=0 $Y2=0
cc_303 N_A3_M1006_g N_VPWR_c_576_n 6.75329e-19 $X=4.055 $Y=2.465 $X2=0 $Y2=0
cc_304 N_A3_M1015_g N_VPWR_c_576_n 0.0128124f $X=4.485 $Y=2.465 $X2=0 $Y2=0
cc_305 N_A3_M1006_g N_VPWR_c_571_n 0.00429087f $X=4.055 $Y=2.465 $X2=0 $Y2=0
cc_306 N_A3_M1015_g N_VPWR_c_571_n 0.00948291f $X=4.485 $Y=2.465 $X2=0 $Y2=0
cc_307 N_A3_c_327_n N_X_c_680_n 2.36797e-19 $X=3.63 $Y=1.26 $X2=0 $Y2=0
cc_308 N_A3_M1006_g N_X_c_680_n 9.61874e-19 $X=4.055 $Y=2.465 $X2=0 $Y2=0
cc_309 A3 N_X_c_680_n 0.00316116f $X=4.475 $Y=1.58 $X2=0 $Y2=0
cc_310 N_A3_c_325_n N_VGND_c_739_n 0.00422101f $X=3.555 $Y=1.185 $X2=0 $Y2=0
cc_311 N_A3_c_328_n N_VGND_c_740_n 0.00451428f $X=3.985 $Y=1.185 $X2=0 $Y2=0
cc_312 N_A3_c_325_n N_VGND_c_741_n 0.0055185f $X=3.555 $Y=1.185 $X2=0 $Y2=0
cc_313 N_A3_c_328_n N_VGND_c_741_n 0.00428906f $X=3.985 $Y=1.185 $X2=0 $Y2=0
cc_314 N_A3_c_325_n N_VGND_c_746_n 0.0102013f $X=3.555 $Y=1.185 $X2=0 $Y2=0
cc_315 N_A3_c_328_n N_VGND_c_746_n 0.00718404f $X=3.985 $Y=1.185 $X2=0 $Y2=0
cc_316 N_A3_c_325_n N_A_726_47#_c_827_n 0.00613518f $X=3.555 $Y=1.185 $X2=0
+ $Y2=0
cc_317 N_A3_c_328_n N_A_726_47#_c_827_n 0.00998155f $X=3.985 $Y=1.185 $X2=0
+ $Y2=0
cc_318 N_A3_c_325_n N_A_726_47#_c_829_n 0.0029314f $X=3.555 $Y=1.185 $X2=0 $Y2=0
cc_319 N_A3_c_326_n N_A_726_47#_c_829_n 5.96206e-19 $X=3.91 $Y=1.26 $X2=0 $Y2=0
cc_320 N_A3_c_328_n N_A_726_47#_c_829_n 7.37415e-19 $X=3.985 $Y=1.185 $X2=0
+ $Y2=0
cc_321 N_A3_c_328_n N_A_726_47#_c_825_n 0.0112083f $X=3.985 $Y=1.185 $X2=0 $Y2=0
cc_322 N_A3_c_330_n N_A_726_47#_c_825_n 8.49651e-19 $X=4.075 $Y=1.26 $X2=0 $Y2=0
cc_323 N_A2_M1005_g N_A1_M1002_g 0.0301204f $X=5.385 $Y=0.755 $X2=0 $Y2=0
cc_324 N_A2_M1013_g N_A1_M1007_g 0.0301204f $X=5.385 $Y=2.465 $X2=0 $Y2=0
cc_325 A2 A1 0.019724f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_326 N_A2_c_403_n A1 2.09547e-19 $X=5.385 $Y=1.51 $X2=0 $Y2=0
cc_327 A2 N_A1_c_452_n 0.00344199f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_328 N_A2_c_403_n N_A1_c_452_n 0.0301204f $X=5.385 $Y=1.51 $X2=0 $Y2=0
cc_329 N_A2_M1001_g N_A_27_367#_c_515_n 0.0152857f $X=4.955 $Y=2.465 $X2=0 $Y2=0
cc_330 A2 N_A_27_367#_c_515_n 0.00638916f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_331 N_A2_M1013_g N_A_27_367#_c_520_n 0.0122129f $X=5.385 $Y=2.465 $X2=0 $Y2=0
cc_332 A2 N_A_27_367#_c_520_n 0.0218763f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_333 A2 N_A_27_367#_c_522_n 0.0162894f $X=5.435 $Y=1.58 $X2=0 $Y2=0
cc_334 N_A2_c_403_n N_A_27_367#_c_522_n 6.37898e-19 $X=5.385 $Y=1.51 $X2=0 $Y2=0
cc_335 N_A2_M1001_g N_VPWR_c_576_n 0.0128331f $X=4.955 $Y=2.465 $X2=0 $Y2=0
cc_336 N_A2_M1013_g N_VPWR_c_576_n 6.51893e-19 $X=5.385 $Y=2.465 $X2=0 $Y2=0
cc_337 N_A2_M1001_g N_VPWR_c_577_n 6.85826e-19 $X=4.955 $Y=2.465 $X2=0 $Y2=0
cc_338 N_A2_M1013_g N_VPWR_c_577_n 0.0145194f $X=5.385 $Y=2.465 $X2=0 $Y2=0
cc_339 N_A2_M1001_g N_VPWR_c_585_n 0.00564095f $X=4.955 $Y=2.465 $X2=0 $Y2=0
cc_340 N_A2_M1013_g N_VPWR_c_585_n 0.00486043f $X=5.385 $Y=2.465 $X2=0 $Y2=0
cc_341 N_A2_M1001_g N_VPWR_c_571_n 0.00948291f $X=4.955 $Y=2.465 $X2=0 $Y2=0
cc_342 N_A2_M1013_g N_VPWR_c_571_n 0.00824727f $X=5.385 $Y=2.465 $X2=0 $Y2=0
cc_343 N_A2_M1000_g N_VGND_c_740_n 0.001817f $X=4.955 $Y=0.755 $X2=0 $Y2=0
cc_344 N_A2_M1000_g N_VGND_c_745_n 0.00300112f $X=4.955 $Y=0.755 $X2=0 $Y2=0
cc_345 N_A2_M1005_g N_VGND_c_745_n 0.00300112f $X=5.385 $Y=0.755 $X2=0 $Y2=0
cc_346 N_A2_M1000_g N_VGND_c_746_n 0.00457098f $X=4.955 $Y=0.755 $X2=0 $Y2=0
cc_347 N_A2_M1005_g N_VGND_c_746_n 0.00417887f $X=5.385 $Y=0.755 $X2=0 $Y2=0
cc_348 N_A2_M1000_g N_A_726_47#_c_825_n 0.0108615f $X=4.955 $Y=0.755 $X2=0 $Y2=0
cc_349 N_A2_M1005_g N_A_726_47#_c_825_n 0.0037714f $X=5.385 $Y=0.755 $X2=0 $Y2=0
cc_350 N_A2_M1000_g N_A_919_67#_c_858_n 0.0115134f $X=4.955 $Y=0.755 $X2=0 $Y2=0
cc_351 N_A2_M1005_g N_A_919_67#_c_858_n 0.0125232f $X=5.385 $Y=0.755 $X2=0 $Y2=0
cc_352 N_A1_M1007_g N_A_27_367#_c_520_n 0.0167636f $X=5.815 $Y=2.465 $X2=0 $Y2=0
cc_353 A1 N_A_27_367#_c_525_n 0.0154476f $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_354 N_A1_c_452_n N_A_27_367#_c_525_n 6.37898e-19 $X=6.245 $Y=1.51 $X2=0 $Y2=0
cc_355 N_A1_M1007_g N_VPWR_c_577_n 0.014473f $X=5.815 $Y=2.465 $X2=0 $Y2=0
cc_356 N_A1_M1019_g N_VPWR_c_577_n 6.77662e-19 $X=6.245 $Y=2.465 $X2=0 $Y2=0
cc_357 N_A1_M1007_g N_VPWR_c_579_n 7.26038e-19 $X=5.815 $Y=2.465 $X2=0 $Y2=0
cc_358 N_A1_M1019_g N_VPWR_c_579_n 0.0200737f $X=6.245 $Y=2.465 $X2=0 $Y2=0
cc_359 A1 N_VPWR_c_579_n 0.0206299f $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_360 N_A1_M1007_g N_VPWR_c_586_n 0.00486043f $X=5.815 $Y=2.465 $X2=0 $Y2=0
cc_361 N_A1_M1019_g N_VPWR_c_586_n 0.00486043f $X=6.245 $Y=2.465 $X2=0 $Y2=0
cc_362 N_A1_M1007_g N_VPWR_c_571_n 0.00824727f $X=5.815 $Y=2.465 $X2=0 $Y2=0
cc_363 N_A1_M1019_g N_VPWR_c_571_n 0.00824727f $X=6.245 $Y=2.465 $X2=0 $Y2=0
cc_364 N_A1_M1002_g N_VGND_c_745_n 0.00300112f $X=5.815 $Y=0.755 $X2=0 $Y2=0
cc_365 N_A1_M1018_g N_VGND_c_745_n 0.00300112f $X=6.245 $Y=0.755 $X2=0 $Y2=0
cc_366 N_A1_M1002_g N_VGND_c_746_n 0.00417887f $X=5.815 $Y=0.755 $X2=0 $Y2=0
cc_367 N_A1_M1018_g N_VGND_c_746_n 0.00445803f $X=6.245 $Y=0.755 $X2=0 $Y2=0
cc_368 N_A1_M1002_g N_A_726_47#_c_825_n 5.22104e-19 $X=5.815 $Y=0.755 $X2=0
+ $Y2=0
cc_369 N_A1_M1002_g N_A_919_67#_c_856_n 0.00990517f $X=5.815 $Y=0.755 $X2=0
+ $Y2=0
cc_370 N_A1_M1018_g N_A_919_67#_c_856_n 0.0124582f $X=6.245 $Y=0.755 $X2=0 $Y2=0
cc_371 N_A1_M1018_g N_A_919_67#_c_857_n 0.00354524f $X=6.245 $Y=0.755 $X2=0
+ $Y2=0
cc_372 A1 N_A_919_67#_c_857_n 0.0147306f $X=6.395 $Y=1.58 $X2=0 $Y2=0
cc_373 N_A_27_367#_c_493_n N_VPWR_M1004_d 0.00521508f $X=4.105 $Y=2.525
+ $X2=-0.19 $Y2=1.655
cc_374 N_A_27_367#_c_493_n N_VPWR_M1008_d 0.00353123f $X=4.105 $Y=2.525 $X2=0
+ $Y2=0
cc_375 N_A_27_367#_c_493_n N_VPWR_M1017_d 0.00805333f $X=4.105 $Y=2.525 $X2=0
+ $Y2=0
cc_376 N_A_27_367#_c_515_n N_VPWR_M1015_d 0.0092871f $X=5.055 $Y=2.015 $X2=0
+ $Y2=0
cc_377 N_A_27_367#_c_520_n N_VPWR_M1013_s 0.00567848f $X=5.935 $Y=2.015 $X2=0
+ $Y2=0
cc_378 N_A_27_367#_c_492_n N_VPWR_c_572_n 0.00965903f $X=1.155 $Y=2.905 $X2=0
+ $Y2=0
cc_379 N_A_27_367#_c_493_n N_VPWR_c_572_n 0.0211261f $X=4.105 $Y=2.525 $X2=0
+ $Y2=0
cc_380 N_A_27_367#_c_493_n N_VPWR_c_573_n 0.0163958f $X=4.105 $Y=2.525 $X2=0
+ $Y2=0
cc_381 N_A_27_367#_c_493_n N_VPWR_c_574_n 0.0163958f $X=4.105 $Y=2.525 $X2=0
+ $Y2=0
cc_382 N_A_27_367#_c_493_n N_VPWR_c_575_n 0.00133711f $X=4.105 $Y=2.525 $X2=0
+ $Y2=0
cc_383 N_A_27_367#_c_537_p N_VPWR_c_575_n 0.0131621f $X=4.27 $Y=2.91 $X2=0 $Y2=0
cc_384 N_A_27_367#_c_517_n N_VPWR_c_575_n 7.19283e-19 $X=4.245 $Y=2.525 $X2=0
+ $Y2=0
cc_385 N_A_27_367#_c_515_n N_VPWR_c_576_n 0.017285f $X=5.055 $Y=2.015 $X2=0
+ $Y2=0
cc_386 N_A_27_367#_c_520_n N_VPWR_c_577_n 0.0170777f $X=5.935 $Y=2.015 $X2=0
+ $Y2=0
cc_387 N_A_27_367#_c_493_n N_VPWR_c_580_n 0.00667889f $X=4.105 $Y=2.525 $X2=0
+ $Y2=0
cc_388 N_A_27_367#_c_493_n N_VPWR_c_582_n 0.00667889f $X=4.105 $Y=2.525 $X2=0
+ $Y2=0
cc_389 N_A_27_367#_c_490_n N_VPWR_c_584_n 0.0211538f $X=0.26 $Y=2.905 $X2=0
+ $Y2=0
cc_390 N_A_27_367#_c_500_n N_VPWR_c_584_n 0.0329923f $X=1.025 $Y=2.99 $X2=0
+ $Y2=0
cc_391 N_A_27_367#_c_492_n N_VPWR_c_584_n 0.0178999f $X=1.155 $Y=2.905 $X2=0
+ $Y2=0
cc_392 N_A_27_367#_c_493_n N_VPWR_c_584_n 0.0102706f $X=4.105 $Y=2.525 $X2=0
+ $Y2=0
cc_393 N_A_27_367#_c_547_p N_VPWR_c_585_n 0.0131621f $X=5.17 $Y=2.91 $X2=0 $Y2=0
cc_394 N_A_27_367#_c_548_p N_VPWR_c_586_n 0.0124525f $X=6.03 $Y=2.91 $X2=0 $Y2=0
cc_395 N_A_27_367#_M1011_d N_VPWR_c_571_n 0.00215158f $X=0.135 $Y=1.835 $X2=0
+ $Y2=0
cc_396 N_A_27_367#_M1022_d N_VPWR_c_571_n 0.00215161f $X=0.98 $Y=1.835 $X2=0
+ $Y2=0
cc_397 N_A_27_367#_M1006_s N_VPWR_c_571_n 0.00330936f $X=4.13 $Y=1.835 $X2=0
+ $Y2=0
cc_398 N_A_27_367#_M1001_d N_VPWR_c_571_n 0.00467071f $X=5.03 $Y=1.835 $X2=0
+ $Y2=0
cc_399 N_A_27_367#_M1007_d N_VPWR_c_571_n 0.00536646f $X=5.89 $Y=1.835 $X2=0
+ $Y2=0
cc_400 N_A_27_367#_c_490_n N_VPWR_c_571_n 0.0126374f $X=0.26 $Y=2.905 $X2=0
+ $Y2=0
cc_401 N_A_27_367#_c_500_n N_VPWR_c_571_n 0.0212291f $X=1.025 $Y=2.99 $X2=0
+ $Y2=0
cc_402 N_A_27_367#_c_492_n N_VPWR_c_571_n 0.0100994f $X=1.155 $Y=2.905 $X2=0
+ $Y2=0
cc_403 N_A_27_367#_c_493_n N_VPWR_c_571_n 0.0498979f $X=4.105 $Y=2.525 $X2=0
+ $Y2=0
cc_404 N_A_27_367#_c_537_p N_VPWR_c_571_n 0.00808656f $X=4.27 $Y=2.91 $X2=0
+ $Y2=0
cc_405 N_A_27_367#_c_547_p N_VPWR_c_571_n 0.00808656f $X=5.17 $Y=2.91 $X2=0
+ $Y2=0
cc_406 N_A_27_367#_c_548_p N_VPWR_c_571_n 0.00730901f $X=6.03 $Y=2.91 $X2=0
+ $Y2=0
cc_407 N_A_27_367#_c_517_n N_VPWR_c_571_n 0.00181391f $X=4.245 $Y=2.525 $X2=0
+ $Y2=0
cc_408 N_A_27_367#_c_493_n N_X_M1004_s 0.00497864f $X=4.105 $Y=2.525 $X2=0 $Y2=0
cc_409 N_A_27_367#_c_493_n N_X_M1012_s 0.00497864f $X=4.105 $Y=2.525 $X2=0 $Y2=0
cc_410 N_A_27_367#_c_564_p N_X_c_679_n 0.0278195f $X=1.12 $Y=2.095 $X2=0 $Y2=0
cc_411 N_A_27_367#_c_493_n N_X_c_679_n 0.0230702f $X=4.105 $Y=2.525 $X2=0 $Y2=0
cc_412 N_A_27_367#_c_493_n N_X_c_680_n 0.107154f $X=4.105 $Y=2.525 $X2=0 $Y2=0
cc_413 N_A_27_367#_c_508_n N_X_c_680_n 0.00560239f $X=4.245 $Y=2.1 $X2=0 $Y2=0
cc_414 N_A_27_367#_c_509_n N_X_c_680_n 0.00491278f $X=4.245 $Y=2.44 $X2=0 $Y2=0
cc_415 N_A_27_367#_c_564_p N_X_c_677_n 0.0186255f $X=1.12 $Y=2.095 $X2=0 $Y2=0
cc_416 N_A_27_367#_c_494_n N_X_c_677_n 0.00173863f $X=1.155 $Y=2.525 $X2=0 $Y2=0
cc_417 N_VPWR_c_571_n N_X_M1004_s 0.00360572f $X=6.48 $Y=3.33 $X2=0 $Y2=0
cc_418 N_VPWR_c_571_n N_X_M1012_s 0.00360572f $X=6.48 $Y=3.33 $X2=0 $Y2=0
cc_419 N_VPWR_M1004_d N_X_c_680_n 0.00615541f $X=1.995 $Y=1.835 $X2=0 $Y2=0
cc_420 N_VPWR_M1008_d N_X_c_680_n 0.00382577f $X=2.84 $Y=1.835 $X2=0 $Y2=0
cc_421 N_X_c_677_n N_VGND_M1016_s 0.0020581f $X=1.665 $Y=1.06 $X2=0 $Y2=0
cc_422 N_X_c_676_n N_VGND_M1014_d 0.00178048f $X=2.735 $Y=1.06 $X2=0 $Y2=0
cc_423 N_X_M1003_s N_VGND_c_746_n 0.00598115f $X=1.41 $Y=0.235 $X2=0 $Y2=0
cc_424 N_X_M1021_s N_VGND_c_746_n 0.00550255f $X=2.5 $Y=0.235 $X2=0 $Y2=0
cc_425 N_VGND_c_746_n N_A_726_47#_M1010_d 0.00233619f $X=6.48 $Y=0 $X2=-0.19
+ $Y2=-0.245
cc_426 N_VGND_c_741_n N_A_726_47#_c_827_n 0.0118985f $X=4.105 $Y=0 $X2=0 $Y2=0
cc_427 N_VGND_c_746_n N_A_726_47#_c_827_n 0.011818f $X=6.48 $Y=0 $X2=0 $Y2=0
cc_428 N_VGND_M1020_s N_A_726_47#_c_825_n 0.00511797f $X=4.06 $Y=0.235 $X2=0
+ $Y2=0
cc_429 N_VGND_c_740_n N_A_726_47#_c_825_n 0.0139731f $X=4.2 $Y=0.38 $X2=0 $Y2=0
cc_430 N_VGND_c_741_n N_A_726_47#_c_825_n 0.00201199f $X=4.105 $Y=0 $X2=0 $Y2=0
cc_431 N_VGND_c_745_n N_A_726_47#_c_825_n 0.00409988f $X=6.48 $Y=0 $X2=0 $Y2=0
cc_432 N_VGND_c_746_n N_A_726_47#_c_825_n 0.0131334f $X=6.48 $Y=0 $X2=0 $Y2=0
cc_433 N_VGND_c_745_n N_A_919_67#_c_856_n 0.0165439f $X=6.48 $Y=0 $X2=0 $Y2=0
cc_434 N_VGND_c_746_n N_A_919_67#_c_856_n 0.0100107f $X=6.48 $Y=0 $X2=0 $Y2=0
cc_435 N_VGND_c_740_n N_A_919_67#_c_858_n 0.0162237f $X=4.2 $Y=0.38 $X2=0 $Y2=0
cc_436 N_VGND_c_745_n N_A_919_67#_c_858_n 0.103157f $X=6.48 $Y=0 $X2=0 $Y2=0
cc_437 N_VGND_c_746_n N_A_919_67#_c_858_n 0.0642503f $X=6.48 $Y=0 $X2=0 $Y2=0
cc_438 N_A_726_47#_c_825_n N_A_919_67#_M1000_s 0.00584144f $X=5.17 $Y=0.81
+ $X2=-0.19 $Y2=-0.245
cc_439 N_A_726_47#_M1000_d N_A_919_67#_c_858_n 0.00179632f $X=5.03 $Y=0.335
+ $X2=0 $Y2=0
cc_440 N_A_726_47#_c_827_n N_A_919_67#_c_858_n 2.78019e-19 $X=3.77 $Y=0.45 $X2=0
+ $Y2=0
cc_441 N_A_726_47#_c_825_n N_A_919_67#_c_858_n 0.0420985f $X=5.17 $Y=0.81 $X2=0
+ $Y2=0
