* File: sky130_fd_sc_lp__maj3_m.pxi.spice
* Created: Wed Sep  2 09:59:51 2020
* 
x_PM_SKY130_FD_SC_LP__MAJ3_M%A N_A_M1013_g N_A_M1010_g N_A_M1007_g N_A_M1002_g A
+ A N_A_c_72_n PM_SKY130_FD_SC_LP__MAJ3_M%A
x_PM_SKY130_FD_SC_LP__MAJ3_M%B N_B_M1004_g N_B_M1011_g N_B_M1012_g N_B_M1005_g B
+ B N_B_c_109_n PM_SKY130_FD_SC_LP__MAJ3_M%B
x_PM_SKY130_FD_SC_LP__MAJ3_M%C N_C_M1000_g N_C_M1003_g N_C_c_151_n N_C_c_152_n
+ N_C_M1008_g N_C_M1006_g C C N_C_c_155_n PM_SKY130_FD_SC_LP__MAJ3_M%C
x_PM_SKY130_FD_SC_LP__MAJ3_M%A_34_57# N_A_34_57#_M1000_s N_A_34_57#_M1004_d
+ N_A_34_57#_M1003_s N_A_34_57#_M1011_d N_A_34_57#_M1009_g N_A_34_57#_M1001_g
+ N_A_34_57#_c_203_n N_A_34_57#_c_213_n N_A_34_57#_c_204_n N_A_34_57#_c_215_n
+ N_A_34_57#_c_216_n N_A_34_57#_c_217_n N_A_34_57#_c_205_n N_A_34_57#_c_218_n
+ N_A_34_57#_c_206_n N_A_34_57#_c_220_n N_A_34_57#_c_207_n N_A_34_57#_c_208_n
+ N_A_34_57#_c_209_n N_A_34_57#_c_221_n N_A_34_57#_c_210_n N_A_34_57#_c_222_n
+ N_A_34_57#_c_223_n PM_SKY130_FD_SC_LP__MAJ3_M%A_34_57#
x_PM_SKY130_FD_SC_LP__MAJ3_M%VPWR N_VPWR_M1010_d N_VPWR_M1006_d N_VPWR_c_303_n
+ N_VPWR_c_304_n VPWR N_VPWR_c_305_n N_VPWR_c_306_n N_VPWR_c_307_n
+ N_VPWR_c_302_n N_VPWR_c_309_n N_VPWR_c_310_n PM_SKY130_FD_SC_LP__MAJ3_M%VPWR
x_PM_SKY130_FD_SC_LP__MAJ3_M%X N_X_M1009_d N_X_M1001_d X X X X X X X N_X_c_340_n
+ PM_SKY130_FD_SC_LP__MAJ3_M%X
x_PM_SKY130_FD_SC_LP__MAJ3_M%VGND N_VGND_M1013_d N_VGND_M1008_d N_VGND_c_354_n
+ N_VGND_c_355_n N_VGND_c_356_n N_VGND_c_357_n VGND N_VGND_c_358_n
+ N_VGND_c_359_n N_VGND_c_360_n N_VGND_c_361_n PM_SKY130_FD_SC_LP__MAJ3_M%VGND
cc_1 VNB N_A_M1013_g 0.0205579f $X=-0.19 $Y=-0.245 $X2=0.92 $Y2=0.495
cc_2 VNB N_A_M1010_g 0.00402602f $X=-0.19 $Y=-0.245 $X2=0.92 $Y2=2.335
cc_3 VNB N_A_M1007_g 0.0205435f $X=-0.19 $Y=-0.245 $X2=1.35 $Y2=0.495
cc_4 VNB N_A_M1002_g 0.0040279f $X=-0.19 $Y=-0.245 $X2=1.35 $Y2=2.335
cc_5 VNB A 0.0135377f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.21
cc_6 VNB N_A_c_72_n 0.066267f $X=-0.19 $Y=-0.245 $X2=1.16 $Y2=1.07
cc_7 VNB N_B_M1004_g 0.0208051f $X=-0.19 $Y=-0.245 $X2=0.92 $Y2=0.495
cc_8 VNB N_B_M1011_g 0.00402681f $X=-0.19 $Y=-0.245 $X2=0.92 $Y2=2.335
cc_9 VNB N_B_M1012_g 0.0206386f $X=-0.19 $Y=-0.245 $X2=1.35 $Y2=0.495
cc_10 VNB N_B_M1005_g 0.0040147f $X=-0.19 $Y=-0.245 $X2=1.35 $Y2=2.335
cc_11 VNB B 0.0143813f $X=-0.19 $Y=-0.245 $X2=1.115 $Y2=1.21
cc_12 VNB N_B_c_109_n 0.0619356f $X=-0.19 $Y=-0.245 $X2=1.16 $Y2=1.07
cc_13 VNB N_C_M1000_g 0.0634655f $X=-0.19 $Y=-0.245 $X2=0.92 $Y2=0.495
cc_14 VNB N_C_M1008_g 0.0606821f $X=-0.19 $Y=-0.245 $X2=1.35 $Y2=0.495
cc_15 VNB N_A_34_57#_M1009_g 0.0505501f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_16 VNB N_A_34_57#_c_203_n 0.0155738f $X=-0.19 $Y=-0.245 $X2=1.16 $Y2=1.07
cc_17 VNB N_A_34_57#_c_204_n 0.0442541f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_18 VNB N_A_34_57#_c_205_n 0.00643025f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_19 VNB N_A_34_57#_c_206_n 0.00671373f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_20 VNB N_A_34_57#_c_207_n 0.00608294f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_21 VNB N_A_34_57#_c_208_n 0.029231f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_22 VNB N_A_34_57#_c_209_n 0.0251105f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_23 VNB N_A_34_57#_c_210_n 0.004396f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_24 VNB N_VPWR_c_302_n 0.163682f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_25 VNB X 0.0522134f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_26 VNB N_X_c_340_n 0.0244231f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_354_n 0.00412757f $X=-0.19 $Y=-0.245 $X2=1.35 $Y2=0.905
cc_28 VNB N_VGND_c_355_n 0.0138114f $X=-0.19 $Y=-0.245 $X2=1.35 $Y2=1.575
cc_29 VNB N_VGND_c_356_n 0.0414407f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_357_n 0.00634747f $X=-0.19 $Y=-0.245 $X2=0.635 $Y2=1.21
cc_31 VNB N_VGND_c_358_n 0.029267f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_359_n 0.0208137f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_360_n 0.248465f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_361_n 0.00500486f $X=-0.19 $Y=-0.245 $X2=0 $Y2=0
cc_35 VPB N_A_M1010_g 0.0307673f $X=-0.19 $Y=1.655 $X2=0.92 $Y2=2.335
cc_36 VPB N_A_M1002_g 0.0307685f $X=-0.19 $Y=1.655 $X2=1.35 $Y2=2.335
cc_37 VPB N_B_M1011_g 0.0306557f $X=-0.19 $Y=1.655 $X2=0.92 $Y2=2.335
cc_38 VPB N_B_M1005_g 0.0305959f $X=-0.19 $Y=1.655 $X2=1.35 $Y2=2.335
cc_39 VPB N_C_M1000_g 0.0599705f $X=-0.19 $Y=1.655 $X2=0.92 $Y2=0.495
cc_40 VPB N_C_c_151_n 0.13061f $X=-0.19 $Y=1.655 $X2=0.92 $Y2=2.335
cc_41 VPB N_C_c_152_n 0.0146273f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_42 VPB N_C_M1008_g 0.0347356f $X=-0.19 $Y=1.655 $X2=1.35 $Y2=0.495
cc_43 VPB C 0.00751444f $X=-0.19 $Y=1.655 $X2=1.35 $Y2=2.335
cc_44 VPB N_C_c_155_n 0.0435266f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_45 VPB N_A_34_57#_M1001_g 0.0292731f $X=-0.19 $Y=1.655 $X2=1.135 $Y2=1.07
cc_46 VPB N_A_34_57#_c_203_n 0.0106535f $X=-0.19 $Y=1.655 $X2=1.16 $Y2=1.07
cc_47 VPB N_A_34_57#_c_213_n 0.0308162f $X=-0.19 $Y=1.655 $X2=0.72 $Y2=1.24
cc_48 VPB N_A_34_57#_c_204_n 0.00463691f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_49 VPB N_A_34_57#_c_215_n 0.0309058f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_50 VPB N_A_34_57#_c_216_n 0.0294005f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_51 VPB N_A_34_57#_c_217_n 0.00173204f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_52 VPB N_A_34_57#_c_218_n 0.0136101f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_53 VPB N_A_34_57#_c_206_n 9.78186e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_54 VPB N_A_34_57#_c_220_n 0.0194662f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_55 VPB N_A_34_57#_c_221_n 0.0132078f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_56 VPB N_A_34_57#_c_222_n 0.00235119f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_57 VPB N_A_34_57#_c_223_n 3.70622e-19 $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_58 VPB N_VPWR_c_303_n 0.0199564f $X=-0.19 $Y=1.655 $X2=1.35 $Y2=0.905
cc_59 VPB N_VPWR_c_304_n 0.0264246f $X=-0.19 $Y=1.655 $X2=1.35 $Y2=1.575
cc_60 VPB N_VPWR_c_305_n 0.0330106f $X=-0.19 $Y=1.655 $X2=0.635 $Y2=1.21
cc_61 VPB N_VPWR_c_306_n 0.049894f $X=-0.19 $Y=1.655 $X2=1.16 $Y2=1.07
cc_62 VPB N_VPWR_c_307_n 0.0198848f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_63 VPB N_VPWR_c_302_n 0.0958771f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_64 VPB N_VPWR_c_309_n 0.00632158f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_310_n 0.0047828f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_66 VPB X 0.0560779f $X=-0.19 $Y=1.655 $X2=0 $Y2=0
cc_67 N_A_M1007_g N_B_M1004_g 0.0444873f $X=1.35 $Y=0.495 $X2=0 $Y2=0
cc_68 N_A_M1002_g N_B_M1011_g 0.0444873f $X=1.35 $Y=2.335 $X2=0 $Y2=0
cc_69 A B 0.0462624f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_70 N_A_c_72_n B 0.00575432f $X=1.16 $Y=1.07 $X2=0 $Y2=0
cc_71 A N_B_c_109_n 6.10835e-19 $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_72 N_A_c_72_n N_B_c_109_n 0.0444873f $X=1.16 $Y=1.07 $X2=0 $Y2=0
cc_73 N_A_M1013_g N_C_M1000_g 0.132692f $X=0.92 $Y=0.495 $X2=0 $Y2=0
cc_74 A N_C_M1000_g 0.00736802f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_75 N_A_M1010_g N_C_c_151_n 0.00917051f $X=0.92 $Y=2.335 $X2=0 $Y2=0
cc_76 N_A_M1002_g N_C_c_151_n 0.00917051f $X=1.35 $Y=2.335 $X2=0 $Y2=0
cc_77 A N_A_34_57#_c_204_n 0.0363256f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_78 N_A_M1010_g N_A_34_57#_c_215_n 0.00219135f $X=0.92 $Y=2.335 $X2=0 $Y2=0
cc_79 N_A_M1010_g N_A_34_57#_c_216_n 0.0141145f $X=0.92 $Y=2.335 $X2=0 $Y2=0
cc_80 N_A_M1002_g N_A_34_57#_c_216_n 0.0171278f $X=1.35 $Y=2.335 $X2=0 $Y2=0
cc_81 A N_A_34_57#_c_216_n 0.0551295f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_82 N_A_c_72_n N_A_34_57#_c_216_n 0.00257849f $X=1.16 $Y=1.07 $X2=0 $Y2=0
cc_83 N_A_M1002_g N_A_34_57#_c_217_n 0.00219135f $X=1.35 $Y=2.335 $X2=0 $Y2=0
cc_84 N_A_M1013_g N_A_34_57#_c_209_n 0.00130204f $X=0.92 $Y=0.495 $X2=0 $Y2=0
cc_85 N_A_M1007_g N_A_34_57#_c_210_n 0.00130204f $X=1.35 $Y=0.495 $X2=0 $Y2=0
cc_86 N_A_M1010_g N_VPWR_c_303_n 0.012349f $X=0.92 $Y=2.335 $X2=0 $Y2=0
cc_87 N_A_M1002_g N_VPWR_c_303_n 0.012349f $X=1.35 $Y=2.335 $X2=0 $Y2=0
cc_88 N_A_M1013_g N_VGND_c_354_n 0.0128952f $X=0.92 $Y=0.495 $X2=0 $Y2=0
cc_89 N_A_M1007_g N_VGND_c_354_n 0.0128952f $X=1.35 $Y=0.495 $X2=0 $Y2=0
cc_90 A N_VGND_c_354_n 0.027631f $X=1.115 $Y=1.21 $X2=0 $Y2=0
cc_91 N_A_c_72_n N_VGND_c_354_n 0.00266929f $X=1.16 $Y=1.07 $X2=0 $Y2=0
cc_92 N_A_M1007_g N_VGND_c_356_n 0.00445056f $X=1.35 $Y=0.495 $X2=0 $Y2=0
cc_93 N_A_M1013_g N_VGND_c_358_n 0.00445056f $X=0.92 $Y=0.495 $X2=0 $Y2=0
cc_94 N_A_M1013_g N_VGND_c_360_n 0.00804604f $X=0.92 $Y=0.495 $X2=0 $Y2=0
cc_95 N_A_M1007_g N_VGND_c_360_n 0.00804604f $X=1.35 $Y=0.495 $X2=0 $Y2=0
cc_96 N_B_M1011_g N_C_c_151_n 0.00921991f $X=1.74 $Y=2.335 $X2=0 $Y2=0
cc_97 N_B_M1005_g N_C_c_151_n 0.00921991f $X=2.17 $Y=2.335 $X2=0 $Y2=0
cc_98 N_B_M1012_g N_C_M1008_g 0.133103f $X=2.17 $Y=0.495 $X2=0 $Y2=0
cc_99 B N_C_M1008_g 0.0024643f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_100 N_B_M1005_g C 0.00324599f $X=2.17 $Y=2.335 $X2=0 $Y2=0
cc_101 N_B_M1011_g N_A_34_57#_c_216_n 0.0109043f $X=1.74 $Y=2.335 $X2=0 $Y2=0
cc_102 B N_A_34_57#_c_216_n 0.0170733f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_103 N_B_M1011_g N_A_34_57#_c_217_n 0.0139948f $X=1.74 $Y=2.335 $X2=0 $Y2=0
cc_104 N_B_M1005_g N_A_34_57#_c_217_n 0.0134f $X=2.17 $Y=2.335 $X2=0 $Y2=0
cc_105 N_B_M1012_g N_A_34_57#_c_205_n 0.00889116f $X=2.17 $Y=0.495 $X2=0 $Y2=0
cc_106 B N_A_34_57#_c_205_n 0.0114588f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_107 N_B_M1005_g N_A_34_57#_c_218_n 0.0109043f $X=2.17 $Y=2.335 $X2=0 $Y2=0
cc_108 B N_A_34_57#_c_218_n 0.0114265f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_109 N_B_M1012_g N_A_34_57#_c_206_n 0.00347443f $X=2.17 $Y=0.495 $X2=0 $Y2=0
cc_110 B N_A_34_57#_c_206_n 0.0543529f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_111 N_B_c_109_n N_A_34_57#_c_206_n 0.00536393f $X=1.83 $Y=1.07 $X2=0 $Y2=0
cc_112 N_B_M1004_g N_A_34_57#_c_210_n 0.00899751f $X=1.74 $Y=0.495 $X2=0 $Y2=0
cc_113 N_B_M1012_g N_A_34_57#_c_210_n 0.00738837f $X=2.17 $Y=0.495 $X2=0 $Y2=0
cc_114 B N_A_34_57#_c_210_n 0.0268037f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_115 N_B_c_109_n N_A_34_57#_c_210_n 0.00263869f $X=1.83 $Y=1.07 $X2=0 $Y2=0
cc_116 N_B_M1011_g N_A_34_57#_c_222_n 0.00280399f $X=1.74 $Y=2.335 $X2=0 $Y2=0
cc_117 N_B_M1005_g N_A_34_57#_c_222_n 0.00280399f $X=2.17 $Y=2.335 $X2=0 $Y2=0
cc_118 B N_A_34_57#_c_222_n 0.0277917f $X=2.075 $Y=1.21 $X2=0 $Y2=0
cc_119 N_B_c_109_n N_A_34_57#_c_222_n 0.00266929f $X=1.83 $Y=1.07 $X2=0 $Y2=0
cc_120 N_B_M1011_g N_VPWR_c_303_n 0.0018473f $X=1.74 $Y=2.335 $X2=0 $Y2=0
cc_121 N_B_M1004_g N_VGND_c_354_n 0.00213234f $X=1.74 $Y=0.495 $X2=0 $Y2=0
cc_122 N_B_M1004_g N_VGND_c_356_n 0.00502664f $X=1.74 $Y=0.495 $X2=0 $Y2=0
cc_123 N_B_M1012_g N_VGND_c_356_n 0.00367856f $X=2.17 $Y=0.495 $X2=0 $Y2=0
cc_124 N_B_M1004_g N_VGND_c_360_n 0.00948649f $X=1.74 $Y=0.495 $X2=0 $Y2=0
cc_125 N_B_M1012_g N_VGND_c_360_n 0.00515454f $X=2.17 $Y=0.495 $X2=0 $Y2=0
cc_126 N_C_M1008_g N_A_34_57#_M1009_g 0.0195205f $X=2.56 $Y=0.495 $X2=0 $Y2=0
cc_127 N_C_M1008_g N_A_34_57#_M1001_g 0.0103776f $X=2.56 $Y=0.495 $X2=0 $Y2=0
cc_128 N_C_M1000_g N_A_34_57#_c_204_n 0.0235399f $X=0.53 $Y=0.495 $X2=0 $Y2=0
cc_129 N_C_M1000_g N_A_34_57#_c_215_n 0.0164411f $X=0.53 $Y=0.495 $X2=0 $Y2=0
cc_130 N_C_M1000_g N_A_34_57#_c_216_n 0.0146407f $X=0.53 $Y=0.495 $X2=0 $Y2=0
cc_131 N_C_c_151_n N_A_34_57#_c_217_n 0.00974716f $X=2.455 $Y=2.99 $X2=0 $Y2=0
cc_132 N_C_M1008_g N_A_34_57#_c_217_n 0.00208887f $X=2.56 $Y=0.495 $X2=0 $Y2=0
cc_133 C N_A_34_57#_c_217_n 0.00648571f $X=2.555 $Y=2.32 $X2=0 $Y2=0
cc_134 N_C_M1008_g N_A_34_57#_c_205_n 0.00759961f $X=2.56 $Y=0.495 $X2=0 $Y2=0
cc_135 N_C_M1008_g N_A_34_57#_c_206_n 0.0284178f $X=2.56 $Y=0.495 $X2=0 $Y2=0
cc_136 N_C_M1008_g N_A_34_57#_c_220_n 0.00250235f $X=2.56 $Y=0.495 $X2=0 $Y2=0
cc_137 C N_A_34_57#_c_220_n 0.00605635f $X=2.555 $Y=2.32 $X2=0 $Y2=0
cc_138 N_C_M1008_g N_A_34_57#_c_207_n 0.00162504f $X=2.56 $Y=0.495 $X2=0 $Y2=0
cc_139 N_C_M1008_g N_A_34_57#_c_208_n 0.0327321f $X=2.56 $Y=0.495 $X2=0 $Y2=0
cc_140 N_C_M1000_g N_A_34_57#_c_209_n 0.0104256f $X=0.53 $Y=0.495 $X2=0 $Y2=0
cc_141 N_C_M1000_g N_A_34_57#_c_221_n 0.00513266f $X=0.53 $Y=0.495 $X2=0 $Y2=0
cc_142 N_C_M1008_g N_A_34_57#_c_210_n 0.00151852f $X=2.56 $Y=0.495 $X2=0 $Y2=0
cc_143 N_C_M1008_g N_A_34_57#_c_223_n 0.00705928f $X=2.56 $Y=0.495 $X2=0 $Y2=0
cc_144 C N_A_34_57#_c_223_n 0.00718163f $X=2.555 $Y=2.32 $X2=0 $Y2=0
cc_145 C N_VPWR_M1006_d 0.00397893f $X=2.555 $Y=2.32 $X2=0 $Y2=0
cc_146 N_C_M1000_g N_VPWR_c_303_n 0.00907102f $X=0.53 $Y=0.495 $X2=0 $Y2=0
cc_147 N_C_c_151_n N_VPWR_c_303_n 0.0326347f $X=2.455 $Y=2.99 $X2=0 $Y2=0
cc_148 N_C_M1008_g N_VPWR_c_304_n 0.00533619f $X=2.56 $Y=0.495 $X2=0 $Y2=0
cc_149 C N_VPWR_c_304_n 0.0585628f $X=2.555 $Y=2.32 $X2=0 $Y2=0
cc_150 N_C_c_155_n N_VPWR_c_304_n 0.00800542f $X=2.62 $Y=2.9 $X2=0 $Y2=0
cc_151 N_C_c_152_n N_VPWR_c_305_n 0.0165614f $X=0.605 $Y=2.99 $X2=0 $Y2=0
cc_152 N_C_c_151_n N_VPWR_c_306_n 0.0347942f $X=2.455 $Y=2.99 $X2=0 $Y2=0
cc_153 C N_VPWR_c_306_n 0.0209793f $X=2.555 $Y=2.32 $X2=0 $Y2=0
cc_154 N_C_c_155_n N_VPWR_c_306_n 0.00210837f $X=2.62 $Y=2.9 $X2=0 $Y2=0
cc_155 N_C_c_152_n N_VPWR_c_302_n 0.0488942f $X=0.605 $Y=2.99 $X2=0 $Y2=0
cc_156 C N_VPWR_c_302_n 0.0124888f $X=2.555 $Y=2.32 $X2=0 $Y2=0
cc_157 N_C_M1000_g N_VGND_c_354_n 0.00213234f $X=0.53 $Y=0.495 $X2=0 $Y2=0
cc_158 N_C_M1008_g N_VGND_c_355_n 0.0113475f $X=2.56 $Y=0.495 $X2=0 $Y2=0
cc_159 N_C_M1008_g N_VGND_c_356_n 0.00384904f $X=2.56 $Y=0.495 $X2=0 $Y2=0
cc_160 N_C_M1000_g N_VGND_c_358_n 0.00502664f $X=0.53 $Y=0.495 $X2=0 $Y2=0
cc_161 N_C_M1000_g N_VGND_c_360_n 0.0101654f $X=0.53 $Y=0.495 $X2=0 $Y2=0
cc_162 N_C_M1008_g N_VGND_c_360_n 0.00595491f $X=2.56 $Y=0.495 $X2=0 $Y2=0
cc_163 N_A_34_57#_c_215_n N_VPWR_c_303_n 0.0145731f $X=0.315 $Y=2.335 $X2=0
+ $Y2=0
cc_164 N_A_34_57#_c_216_n N_VPWR_c_303_n 0.026201f $X=1.79 $Y=1.84 $X2=0 $Y2=0
cc_165 N_A_34_57#_c_217_n N_VPWR_c_303_n 0.0145731f $X=1.955 $Y=2.335 $X2=0
+ $Y2=0
cc_166 N_A_34_57#_M1001_g N_VPWR_c_304_n 0.00517169f $X=3.345 $Y=2.335 $X2=0
+ $Y2=0
cc_167 N_A_34_57#_c_213_n N_VPWR_c_304_n 0.00192747f $X=3.152 $Y=1.925 $X2=0
+ $Y2=0
cc_168 N_A_34_57#_c_220_n N_VPWR_c_304_n 0.0211474f $X=2.885 $Y=1.84 $X2=0 $Y2=0
cc_169 N_A_34_57#_M1001_g N_VPWR_c_307_n 0.00293455f $X=3.345 $Y=2.335 $X2=0
+ $Y2=0
cc_170 N_A_34_57#_M1001_g N_VPWR_c_302_n 0.00359002f $X=3.345 $Y=2.335 $X2=0
+ $Y2=0
cc_171 N_A_34_57#_c_215_n N_VPWR_c_302_n 0.0137274f $X=0.315 $Y=2.335 $X2=0
+ $Y2=0
cc_172 N_A_34_57#_c_217_n N_VPWR_c_302_n 0.0136322f $X=1.955 $Y=2.335 $X2=0
+ $Y2=0
cc_173 N_A_34_57#_M1009_g X 0.0367994f $X=3.265 $Y=0.495 $X2=0 $Y2=0
cc_174 N_A_34_57#_M1001_g X 0.0217067f $X=3.345 $Y=2.335 $X2=0 $Y2=0
cc_175 N_A_34_57#_c_213_n X 0.00614085f $X=3.152 $Y=1.925 $X2=0 $Y2=0
cc_176 N_A_34_57#_c_220_n X 0.0130008f $X=2.885 $Y=1.84 $X2=0 $Y2=0
cc_177 N_A_34_57#_c_207_n X 0.0378286f $X=3.05 $Y=1.42 $X2=0 $Y2=0
cc_178 N_A_34_57#_M1009_g N_X_c_340_n 0.00779693f $X=3.265 $Y=0.495 $X2=0 $Y2=0
cc_179 N_A_34_57#_c_209_n N_VGND_c_354_n 0.0145731f $X=0.315 $Y=0.495 $X2=0
+ $Y2=0
cc_180 N_A_34_57#_c_210_n N_VGND_c_354_n 0.0145731f $X=1.955 $Y=0.495 $X2=0
+ $Y2=0
cc_181 N_A_34_57#_M1009_g N_VGND_c_355_n 0.00636796f $X=3.265 $Y=0.495 $X2=0
+ $Y2=0
cc_182 N_A_34_57#_c_205_n N_VGND_c_355_n 0.0131309f $X=2.455 $Y=0.64 $X2=0 $Y2=0
cc_183 N_A_34_57#_c_207_n N_VGND_c_355_n 0.0093538f $X=3.05 $Y=1.42 $X2=0 $Y2=0
cc_184 N_A_34_57#_c_208_n N_VGND_c_355_n 0.00162143f $X=3.05 $Y=1.42 $X2=0 $Y2=0
cc_185 N_A_34_57#_c_205_n N_VGND_c_356_n 0.00955596f $X=2.455 $Y=0.64 $X2=0
+ $Y2=0
cc_186 N_A_34_57#_c_210_n N_VGND_c_356_n 0.0213225f $X=1.955 $Y=0.495 $X2=0
+ $Y2=0
cc_187 N_A_34_57#_c_209_n N_VGND_c_358_n 0.0217285f $X=0.315 $Y=0.495 $X2=0
+ $Y2=0
cc_188 N_A_34_57#_M1009_g N_VGND_c_359_n 0.00502664f $X=3.265 $Y=0.495 $X2=0
+ $Y2=0
cc_189 N_A_34_57#_M1009_g N_VGND_c_360_n 0.0105021f $X=3.265 $Y=0.495 $X2=0
+ $Y2=0
cc_190 N_A_34_57#_c_205_n N_VGND_c_360_n 0.014308f $X=2.455 $Y=0.64 $X2=0 $Y2=0
cc_191 N_A_34_57#_c_209_n N_VGND_c_360_n 0.0125175f $X=0.315 $Y=0.495 $X2=0
+ $Y2=0
cc_192 N_A_34_57#_c_210_n N_VGND_c_360_n 0.0123397f $X=1.955 $Y=0.495 $X2=0
+ $Y2=0
cc_193 N_A_34_57#_c_205_n A_449_57# 0.00198548f $X=2.455 $Y=0.64 $X2=-0.19
+ $Y2=-0.245
cc_194 N_VPWR_c_304_n X 0.0429422f $X=3.05 $Y=2.335 $X2=0 $Y2=0
cc_195 N_VPWR_c_307_n X 0.0107254f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_196 N_VPWR_c_302_n X 0.0114362f $X=3.6 $Y=3.33 $X2=0 $Y2=0
cc_197 N_X_c_340_n N_VGND_c_355_n 0.0185622f $X=3.48 $Y=0.495 $X2=0 $Y2=0
cc_198 N_X_c_340_n N_VGND_c_359_n 0.0272774f $X=3.48 $Y=0.495 $X2=0 $Y2=0
cc_199 N_X_c_340_n N_VGND_c_360_n 0.0156449f $X=3.48 $Y=0.495 $X2=0 $Y2=0
