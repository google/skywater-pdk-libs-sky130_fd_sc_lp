* File: sky130_fd_sc_lp__einvp_8.pex.spice
* Created: Wed Sep  2 09:52:42 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_LP__EINVP_8%A_182_367# 1 2 9 10 11 13 14 16 18 19 21 23
+ 24 26 28 29 31 33 34 36 38 39 41 43 44 46 48 50 51 52 53 54 55 56 57 58 59 61
+ 65 71
c162 44 0 5.29075e-20 $X=5.1 $Y=1.65
c163 39 0 4.0679e-20 $X=4.67 $Y=1.65
c164 19 0 4.0679e-20 $X=2.95 $Y=1.65
c165 16 0 9.60268e-20 $X=2.595 $Y=1.725
c166 9 0 3.96626e-20 $X=2.09 $Y=1.685
r167 70 71 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.5
+ $Y=2.095 $X2=1.5 $Y2=2.095
r168 68 70 1.4878 $w=6.15e-07 $l=7.5e-08 $layer=LI1_cond $X=1.28 $Y=2.02
+ $X2=1.28 $Y2=2.095
r169 63 68 6.70087 $w=6.15e-07 $l=2.13014e-07 $layer=LI1_cond $X=1.17 $Y=1.855
+ $X2=1.28 $Y2=2.02
r170 63 65 54.2443 $w=2.88e-07 $l=1.365e-06 $layer=LI1_cond $X=1.17 $Y=1.855
+ $X2=1.17 $Y2=0.49
r171 59 70 3.1996 $w=6.7e-07 $l=1.7e-07 $layer=LI1_cond $X=1.28 $Y=2.265
+ $X2=1.28 $Y2=2.095
r172 59 61 11.5145 $w=6.68e-07 $l=6.45e-07 $layer=LI1_cond $X=1.28 $Y=2.265
+ $X2=1.28 $Y2=2.91
r173 51 71 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=1.5 $Y=2.08 $X2=1.5
+ $Y2=2.095
r174 50 51 43.5886 $w=3.3e-07 $l=1.5e-07 $layer=POLY_cond $X=1.542 $Y=1.93
+ $X2=1.542 $Y2=2.08
r175 46 48 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=5.175 $Y=1.725
+ $X2=5.175 $Y2=2.465
r176 45 58 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.82 $Y=1.65
+ $X2=4.745 $Y2=1.65
r177 44 46 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.1 $Y=1.65
+ $X2=5.175 $Y2=1.725
r178 44 45 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=5.1 $Y=1.65
+ $X2=4.82 $Y2=1.65
r179 41 58 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.745 $Y=1.725
+ $X2=4.745 $Y2=1.65
r180 41 43 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=4.745 $Y=1.725
+ $X2=4.745 $Y2=2.465
r181 40 57 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.39 $Y=1.65
+ $X2=4.315 $Y2=1.65
r182 39 58 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.67 $Y=1.65
+ $X2=4.745 $Y2=1.65
r183 39 40 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=4.67 $Y=1.65
+ $X2=4.39 $Y2=1.65
r184 36 57 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.315 $Y=1.725
+ $X2=4.315 $Y2=1.65
r185 36 38 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=4.315 $Y=1.725
+ $X2=4.315 $Y2=2.465
r186 35 56 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.96 $Y=1.65
+ $X2=3.885 $Y2=1.65
r187 34 57 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.24 $Y=1.65
+ $X2=4.315 $Y2=1.65
r188 34 35 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=4.24 $Y=1.65
+ $X2=3.96 $Y2=1.65
r189 31 56 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.885 $Y=1.725
+ $X2=3.885 $Y2=1.65
r190 31 33 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=3.885 $Y=1.725
+ $X2=3.885 $Y2=2.465
r191 30 55 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.53 $Y=1.65
+ $X2=3.455 $Y2=1.65
r192 29 56 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.81 $Y=1.65
+ $X2=3.885 $Y2=1.65
r193 29 30 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=3.81 $Y=1.65
+ $X2=3.53 $Y2=1.65
r194 26 55 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.455 $Y=1.725
+ $X2=3.455 $Y2=1.65
r195 26 28 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=3.455 $Y=1.725
+ $X2=3.455 $Y2=2.465
r196 25 54 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.1 $Y=1.65
+ $X2=3.025 $Y2=1.65
r197 24 55 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.38 $Y=1.65
+ $X2=3.455 $Y2=1.65
r198 24 25 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=3.38 $Y=1.65
+ $X2=3.1 $Y2=1.65
r199 21 54 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.025 $Y=1.725
+ $X2=3.025 $Y2=1.65
r200 21 23 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=3.025 $Y=1.725
+ $X2=3.025 $Y2=2.465
r201 20 53 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.67 $Y=1.65
+ $X2=2.595 $Y2=1.65
r202 19 54 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.95 $Y=1.65
+ $X2=3.025 $Y2=1.65
r203 19 20 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.95 $Y=1.65
+ $X2=2.67 $Y2=1.65
r204 16 53 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.595 $Y=1.725
+ $X2=2.595 $Y2=1.65
r205 16 18 237.787 $w=1.5e-07 $l=7.4e-07 $layer=POLY_cond $X=2.595 $Y=1.725
+ $X2=2.595 $Y2=2.465
r206 15 52 20.4101 $w=1.5e-07 $l=8.30662e-08 $layer=POLY_cond $X=2.24 $Y=1.65
+ $X2=2.165 $Y2=1.667
r207 14 53 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.52 $Y=1.65
+ $X2=2.595 $Y2=1.65
r208 14 15 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=2.52 $Y=1.65
+ $X2=2.24 $Y2=1.65
r209 11 52 5.30422 $w=1.5e-07 $l=9.3e-08 $layer=POLY_cond $X=2.165 $Y=1.76
+ $X2=2.165 $Y2=1.667
r210 11 13 226.54 $w=1.5e-07 $l=7.05e-07 $layer=POLY_cond $X=2.165 $Y=1.76
+ $X2=2.165 $Y2=2.465
r211 9 52 20.4101 $w=1.5e-07 $l=8.35165e-08 $layer=POLY_cond $X=2.09 $Y=1.685
+ $X2=2.165 $Y2=1.667
r212 9 10 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=2.09 $Y=1.685
+ $X2=1.75 $Y2=1.685
r213 7 10 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.675 $Y=1.76
+ $X2=1.75 $Y2=1.685
r214 7 50 87.1702 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=1.675 $Y=1.76
+ $X2=1.675 $Y2=1.93
r215 2 68 400 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_PDIFF $count=1 $X=0.91
+ $Y=1.835 $X2=1.05 $Y2=2.02
r216 2 61 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=0.91
+ $Y=1.835 $X2=1.05 $Y2=2.91
r217 1 65 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=1.01
+ $Y=0.345 $X2=1.15 $Y2=0.49
.ends

.subckt PM_SKY130_FD_SC_LP__EINVP_8%TE 3 5 7 8 9 10 12 13 14 15 17 18 20 22 23
+ 25 27 28 30 32 33 35 37 38 40 42 43 45 47 48 52 53 54 55 56 57 58 60
c148 43 0 1.72434e-19 $X=5.13 $Y=1.275
r149 67 68 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.64
+ $Y=1.46 $X2=0.64 $Y2=1.46
r150 60 68 1.77197 $w=5.38e-07 $l=8e-08 $layer=LI1_cond $X=0.72 $Y=1.48 $X2=0.64
+ $Y2=1.48
r151 58 68 8.85984 $w=5.38e-07 $l=4e-07 $layer=LI1_cond $X=0.24 $Y=1.48 $X2=0.64
+ $Y2=1.48
r152 49 50 13.7322 $w=3.51e-07 $l=1e-07 $layer=POLY_cond $X=0.835 $Y=1.442
+ $X2=0.935 $Y2=1.442
r153 48 67 20.9834 $w=3.3e-07 $l=1.2e-07 $layer=POLY_cond $X=0.76 $Y=1.46
+ $X2=0.64 $Y2=1.46
r154 48 49 10.5316 $w=3.51e-07 $l=8.35165e-08 $layer=POLY_cond $X=0.76 $Y=1.46
+ $X2=0.835 $Y2=1.442
r155 45 47 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=5.205 $Y=1.185
+ $X2=5.205 $Y2=0.655
r156 44 57 17.4919 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=4.85 $Y=1.275
+ $X2=4.775 $Y2=1.275
r157 43 45 27.2212 $w=1.8e-07 $l=1.21861e-07 $layer=POLY_cond $X=5.13 $Y=1.275
+ $X2=5.205 $Y2=1.185
r158 43 44 108.839 $w=1.8e-07 $l=2.8e-07 $layer=POLY_cond $X=5.13 $Y=1.275
+ $X2=4.85 $Y2=1.275
r159 40 57 7.92773 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=4.775 $Y=1.185
+ $X2=4.775 $Y2=1.275
r160 40 42 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=4.775 $Y=1.185
+ $X2=4.775 $Y2=0.655
r161 39 56 17.4919 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=4.42 $Y=1.275
+ $X2=4.345 $Y2=1.275
r162 38 57 17.4919 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=4.7 $Y=1.275
+ $X2=4.775 $Y2=1.275
r163 38 39 108.839 $w=1.8e-07 $l=2.8e-07 $layer=POLY_cond $X=4.7 $Y=1.275
+ $X2=4.42 $Y2=1.275
r164 35 56 7.92773 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=4.345 $Y=1.185
+ $X2=4.345 $Y2=1.275
r165 35 37 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=4.345 $Y=1.185
+ $X2=4.345 $Y2=0.655
r166 34 55 17.4919 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=3.99 $Y=1.275
+ $X2=3.915 $Y2=1.275
r167 33 56 17.4919 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=4.27 $Y=1.275
+ $X2=4.345 $Y2=1.275
r168 33 34 108.839 $w=1.8e-07 $l=2.8e-07 $layer=POLY_cond $X=4.27 $Y=1.275
+ $X2=3.99 $Y2=1.275
r169 30 55 7.92773 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.915 $Y=1.185
+ $X2=3.915 $Y2=1.275
r170 30 32 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=3.915 $Y=1.185
+ $X2=3.915 $Y2=0.655
r171 29 54 17.4919 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=3.56 $Y=1.275
+ $X2=3.485 $Y2=1.275
r172 28 55 17.4919 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=3.84 $Y=1.275
+ $X2=3.915 $Y2=1.275
r173 28 29 108.839 $w=1.8e-07 $l=2.8e-07 $layer=POLY_cond $X=3.84 $Y=1.275
+ $X2=3.56 $Y2=1.275
r174 25 54 7.92773 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.485 $Y=1.185
+ $X2=3.485 $Y2=1.275
r175 25 27 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=3.485 $Y=1.185
+ $X2=3.485 $Y2=0.655
r176 24 53 17.4919 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=3.13 $Y=1.275
+ $X2=3.055 $Y2=1.275
r177 23 54 17.4919 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=3.41 $Y=1.275
+ $X2=3.485 $Y2=1.275
r178 23 24 108.839 $w=1.8e-07 $l=2.8e-07 $layer=POLY_cond $X=3.41 $Y=1.275
+ $X2=3.13 $Y2=1.275
r179 20 53 7.92773 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.055 $Y=1.185
+ $X2=3.055 $Y2=1.275
r180 20 22 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=3.055 $Y=1.185
+ $X2=3.055 $Y2=0.655
r181 19 52 17.4919 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=2.7 $Y=1.275
+ $X2=2.625 $Y2=1.275
r182 18 53 17.4919 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=2.98 $Y=1.275
+ $X2=3.055 $Y2=1.275
r183 18 19 108.839 $w=1.8e-07 $l=2.8e-07 $layer=POLY_cond $X=2.98 $Y=1.275
+ $X2=2.7 $Y2=1.275
r184 15 52 7.92773 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=2.625 $Y=1.185
+ $X2=2.625 $Y2=1.275
r185 15 17 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.625 $Y=1.185
+ $X2=2.625 $Y2=0.655
r186 14 51 20.0833 $w=1.8e-07 $l=8.52936e-08 $layer=POLY_cond $X=2.27 $Y=1.275
+ $X2=2.195 $Y2=1.297
r187 13 52 17.4919 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=2.55 $Y=1.275
+ $X2=2.625 $Y2=1.275
r188 13 14 108.839 $w=1.8e-07 $l=2.8e-07 $layer=POLY_cond $X=2.55 $Y=1.275
+ $X2=2.27 $Y2=1.275
r189 10 51 7.00825 $w=1.5e-07 $l=1.12e-07 $layer=POLY_cond $X=2.195 $Y=1.185
+ $X2=2.195 $Y2=1.297
r190 10 12 170.307 $w=1.5e-07 $l=5.3e-07 $layer=POLY_cond $X=2.195 $Y=1.185
+ $X2=2.195 $Y2=0.655
r191 9 50 26.4367 $w=3.51e-07 $l=1.39549e-07 $layer=POLY_cond $X=1.01 $Y=1.335
+ $X2=0.935 $Y2=1.442
r192 8 51 228.943 $w=1.79e-07 $l=8.63791e-07 $layer=POLY_cond $X=1.35 $Y=1.335
+ $X2=2.195 $Y2=1.297
r193 8 9 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=1.35 $Y=1.335 $X2=1.01
+ $Y2=1.335
r194 5 50 22.6971 $w=1.5e-07 $l=1.82e-07 $layer=POLY_cond $X=0.935 $Y=1.26
+ $X2=0.935 $Y2=1.442
r195 5 7 159.06 $w=1.5e-07 $l=4.95e-07 $layer=POLY_cond $X=0.935 $Y=1.26
+ $X2=0.935 $Y2=0.765
r196 1 49 22.6971 $w=1.5e-07 $l=1.83e-07 $layer=POLY_cond $X=0.835 $Y=1.625
+ $X2=0.835 $Y2=1.442
r197 1 3 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=0.835 $Y=1.625
+ $X2=0.835 $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__EINVP_8%A 3 7 11 15 19 23 27 31 35 39 43 47 51 55 59
+ 63 67 70 74 75 76 103
c158 39 0 7.73427e-20 $X=7.355 $Y=0.655
c159 15 0 8.34392e-20 $X=6.065 $Y=0.655
r160 102 103 5.24584 $w=3.3e-07 $l=3e-08 $layer=POLY_cond $X=8.615 $Y=1.49
+ $X2=8.645 $Y2=1.49
r161 101 102 69.9445 $w=3.3e-07 $l=4e-07 $layer=POLY_cond $X=8.215 $Y=1.49
+ $X2=8.615 $Y2=1.49
r162 100 101 5.24584 $w=3.3e-07 $l=3e-08 $layer=POLY_cond $X=8.185 $Y=1.49
+ $X2=8.215 $Y2=1.49
r163 97 98 5.24584 $w=3.3e-07 $l=3e-08 $layer=POLY_cond $X=7.755 $Y=1.49
+ $X2=7.785 $Y2=1.49
r164 96 97 69.9445 $w=3.3e-07 $l=4e-07 $layer=POLY_cond $X=7.355 $Y=1.49
+ $X2=7.755 $Y2=1.49
r165 95 96 5.24584 $w=3.3e-07 $l=3e-08 $layer=POLY_cond $X=7.325 $Y=1.49
+ $X2=7.355 $Y2=1.49
r166 92 93 5.24584 $w=3.3e-07 $l=3e-08 $layer=POLY_cond $X=6.895 $Y=1.49
+ $X2=6.925 $Y2=1.49
r167 90 92 16.6118 $w=3.3e-07 $l=9.5e-08 $layer=POLY_cond $X=6.8 $Y=1.49
+ $X2=6.895 $Y2=1.49
r168 90 91 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.8
+ $Y=1.49 $X2=6.8 $Y2=1.49
r169 88 90 53.3327 $w=3.3e-07 $l=3.05e-07 $layer=POLY_cond $X=6.495 $Y=1.49
+ $X2=6.8 $Y2=1.49
r170 87 88 5.24584 $w=3.3e-07 $l=3e-08 $layer=POLY_cond $X=6.465 $Y=1.49
+ $X2=6.495 $Y2=1.49
r171 85 87 0.874306 $w=3.3e-07 $l=5e-09 $layer=POLY_cond $X=6.46 $Y=1.49
+ $X2=6.465 $Y2=1.49
r172 85 86 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.46
+ $Y=1.49 $X2=6.46 $Y2=1.49
r173 83 85 69.0702 $w=3.3e-07 $l=3.95e-07 $layer=POLY_cond $X=6.065 $Y=1.49
+ $X2=6.46 $Y2=1.49
r174 82 83 5.24584 $w=3.3e-07 $l=3e-08 $layer=POLY_cond $X=6.035 $Y=1.49
+ $X2=6.065 $Y2=1.49
r175 81 82 69.9445 $w=3.3e-07 $l=4e-07 $layer=POLY_cond $X=5.635 $Y=1.49
+ $X2=6.035 $Y2=1.49
r176 79 81 5.24584 $w=3.3e-07 $l=3e-08 $layer=POLY_cond $X=5.605 $Y=1.49
+ $X2=5.635 $Y2=1.49
r177 76 91 4.78937 $w=3.83e-07 $l=1.6e-07 $layer=LI1_cond $X=6.96 $Y=1.402
+ $X2=6.8 $Y2=1.402
r178 75 91 9.57875 $w=3.83e-07 $l=3.2e-07 $layer=LI1_cond $X=6.48 $Y=1.402
+ $X2=6.8 $Y2=1.402
r179 75 86 0.598672 $w=3.83e-07 $l=2e-08 $layer=LI1_cond $X=6.48 $Y=1.402
+ $X2=6.46 $Y2=1.402
r180 73 95 32.3493 $w=3.3e-07 $l=1.85e-07 $layer=POLY_cond $X=7.14 $Y=1.49
+ $X2=7.325 $Y2=1.49
r181 73 93 37.5952 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=7.14 $Y=1.49
+ $X2=6.925 $Y2=1.49
r182 72 74 4.55785 $w=3.83e-07 $l=1.05e-07 $layer=LI1_cond $X=7.14 $Y=1.402
+ $X2=7.245 $Y2=1.402
r183 72 73 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.14
+ $Y=1.49 $X2=7.14 $Y2=1.49
r184 70 76 2.78382 $w=3.83e-07 $l=9.3e-08 $layer=LI1_cond $X=7.053 $Y=1.402
+ $X2=6.96 $Y2=1.402
r185 70 72 2.60422 $w=3.83e-07 $l=8.7e-08 $layer=LI1_cond $X=7.053 $Y=1.402
+ $X2=7.14 $Y2=1.402
r186 68 100 63.8244 $w=3.3e-07 $l=3.65e-07 $layer=POLY_cond $X=7.82 $Y=1.49
+ $X2=8.185 $Y2=1.49
r187 68 98 6.12014 $w=3.3e-07 $l=3.5e-08 $layer=POLY_cond $X=7.82 $Y=1.49
+ $X2=7.785 $Y2=1.49
r188 67 74 26.5062 $w=2.48e-07 $l=5.75e-07 $layer=LI1_cond $X=7.82 $Y=1.47
+ $X2=7.245 $Y2=1.47
r189 67 68 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.82
+ $Y=1.49 $X2=7.82 $Y2=1.49
r190 61 103 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.645 $Y=1.325
+ $X2=8.645 $Y2=1.49
r191 61 63 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=8.645 $Y=1.325
+ $X2=8.645 $Y2=0.655
r192 57 102 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.615 $Y=1.655
+ $X2=8.615 $Y2=1.49
r193 57 59 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=8.615 $Y=1.655
+ $X2=8.615 $Y2=2.465
r194 53 101 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.215 $Y=1.325
+ $X2=8.215 $Y2=1.49
r195 53 55 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=8.215 $Y=1.325
+ $X2=8.215 $Y2=0.655
r196 49 100 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=8.185 $Y=1.655
+ $X2=8.185 $Y2=1.49
r197 49 51 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=8.185 $Y=1.655
+ $X2=8.185 $Y2=2.465
r198 45 98 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.785 $Y=1.325
+ $X2=7.785 $Y2=1.49
r199 45 47 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=7.785 $Y=1.325
+ $X2=7.785 $Y2=0.655
r200 41 97 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.755 $Y=1.655
+ $X2=7.755 $Y2=1.49
r201 41 43 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=7.755 $Y=1.655
+ $X2=7.755 $Y2=2.465
r202 37 96 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.355 $Y=1.325
+ $X2=7.355 $Y2=1.49
r203 37 39 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=7.355 $Y=1.325
+ $X2=7.355 $Y2=0.655
r204 33 95 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.325 $Y=1.655
+ $X2=7.325 $Y2=1.49
r205 33 35 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=7.325 $Y=1.655
+ $X2=7.325 $Y2=2.465
r206 29 93 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.925 $Y=1.325
+ $X2=6.925 $Y2=1.49
r207 29 31 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=6.925 $Y=1.325
+ $X2=6.925 $Y2=0.655
r208 25 92 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.895 $Y=1.655
+ $X2=6.895 $Y2=1.49
r209 25 27 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=6.895 $Y=1.655
+ $X2=6.895 $Y2=2.465
r210 21 88 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.495 $Y=1.325
+ $X2=6.495 $Y2=1.49
r211 21 23 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=6.495 $Y=1.325
+ $X2=6.495 $Y2=0.655
r212 17 87 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.465 $Y=1.655
+ $X2=6.465 $Y2=1.49
r213 17 19 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=6.465 $Y=1.655
+ $X2=6.465 $Y2=2.465
r214 13 83 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.065 $Y=1.325
+ $X2=6.065 $Y2=1.49
r215 13 15 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=6.065 $Y=1.325
+ $X2=6.065 $Y2=0.655
r216 9 82 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.035 $Y=1.655
+ $X2=6.035 $Y2=1.49
r217 9 11 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=6.035 $Y=1.655
+ $X2=6.035 $Y2=2.465
r218 5 81 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.635 $Y=1.325
+ $X2=5.635 $Y2=1.49
r219 5 7 343.553 $w=1.5e-07 $l=6.7e-07 $layer=POLY_cond $X=5.635 $Y=1.325
+ $X2=5.635 $Y2=0.655
r220 1 79 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.605 $Y=1.655
+ $X2=5.605 $Y2=1.49
r221 1 3 415.34 $w=1.5e-07 $l=8.1e-07 $layer=POLY_cond $X=5.605 $Y=1.655
+ $X2=5.605 $Y2=2.465
.ends

.subckt PM_SKY130_FD_SC_LP__EINVP_8%VPWR 1 2 3 4 5 18 24 28 32 38 44 48 49 50 52
+ 61 66 73 74 77 80 83 86
r115 86 87 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=5.04 $Y=3.33
+ $X2=5.04 $Y2=3.33
r116 83 84 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=3.33
+ $X2=4.08 $Y2=3.33
r117 80 81 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=3.33
+ $X2=3.12 $Y2=3.33
r118 77 78 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.72 $Y=3.33
+ $X2=0.72 $Y2=3.33
r119 74 87 1.07034 $w=4.9e-07 $l=3.84e-06 $layer=MET1_cond $X=8.88 $Y=3.33
+ $X2=5.04 $Y2=3.33
r120 73 74 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=8.88 $Y=3.33
+ $X2=8.88 $Y2=3.33
r121 71 86 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=5.09 $Y=3.33
+ $X2=4.96 $Y2=3.33
r122 71 73 247.262 $w=1.68e-07 $l=3.79e-06 $layer=LI1_cond $X=5.09 $Y=3.33
+ $X2=8.88 $Y2=3.33
r123 67 83 7.13466 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=4.225 $Y=3.33
+ $X2=4.097 $Y2=3.33
r124 67 69 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=4.225 $Y=3.33
+ $X2=4.56 $Y2=3.33
r125 66 86 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=4.83 $Y=3.33
+ $X2=4.96 $Y2=3.33
r126 66 69 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=4.83 $Y=3.33
+ $X2=4.56 $Y2=3.33
r127 65 84 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=4.08 $Y2=3.33
r128 65 81 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=3.33
+ $X2=3.12 $Y2=3.33
r129 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.33 $X2=3.6
+ $Y2=3.33
r130 62 80 7.34436 $w=1.7e-07 $l=1.33e-07 $layer=LI1_cond $X=3.37 $Y=3.33
+ $X2=3.237 $Y2=3.33
r131 62 64 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=3.37 $Y=3.33
+ $X2=3.6 $Y2=3.33
r132 61 83 7.13466 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=3.97 $Y=3.33
+ $X2=4.097 $Y2=3.33
r133 61 64 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=3.97 $Y=3.33 $X2=3.6
+ $Y2=3.33
r134 60 81 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=3.12 $Y2=3.33
r135 60 78 0.401378 $w=4.9e-07 $l=1.44e-06 $layer=MET1_cond $X=2.16 $Y=3.33
+ $X2=0.72 $Y2=3.33
r136 59 60 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.16 $Y=3.33
+ $X2=2.16 $Y2=3.33
r137 57 77 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=0.725 $Y=3.33
+ $X2=0.59 $Y2=3.33
r138 57 59 93.6203 $w=1.68e-07 $l=1.435e-06 $layer=LI1_cond $X=0.725 $Y=3.33
+ $X2=2.16 $Y2=3.33
r139 55 78 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=3.33
+ $X2=0.72 $Y2=3.33
r140 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=3.33
+ $X2=0.24 $Y2=3.33
r141 52 77 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=0.455 $Y=3.33
+ $X2=0.59 $Y2=3.33
r142 52 54 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=0.455 $Y=3.33
+ $X2=0.24 $Y2=3.33
r143 50 87 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=5.04 $Y2=3.33
r144 50 84 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=3.33
+ $X2=4.08 $Y2=3.33
r145 50 69 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=3.33
+ $X2=4.56 $Y2=3.33
r146 48 59 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=2.245 $Y=3.33
+ $X2=2.16 $Y2=3.33
r147 48 49 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.245 $Y=3.33
+ $X2=2.375 $Y2=3.33
r148 44 47 39.6706 $w=2.58e-07 $l=8.95e-07 $layer=LI1_cond $X=4.96 $Y=2.055
+ $X2=4.96 $Y2=2.95
r149 42 86 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=4.96 $Y=3.245
+ $X2=4.96 $Y2=3.33
r150 42 47 13.0758 $w=2.58e-07 $l=2.95e-07 $layer=LI1_cond $X=4.96 $Y=3.245
+ $X2=4.96 $Y2=2.95
r151 38 41 40.4485 $w=2.53e-07 $l=8.95e-07 $layer=LI1_cond $X=4.097 $Y=2.055
+ $X2=4.097 $Y2=2.95
r152 36 83 0.067832 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=4.097 $Y=3.245
+ $X2=4.097 $Y2=3.33
r153 36 41 13.3322 $w=2.53e-07 $l=2.95e-07 $layer=LI1_cond $X=4.097 $Y=3.245
+ $X2=4.097 $Y2=2.95
r154 32 35 38.9221 $w=2.63e-07 $l=8.95e-07 $layer=LI1_cond $X=3.237 $Y=2.055
+ $X2=3.237 $Y2=2.95
r155 30 80 0.195364 $w=2.65e-07 $l=8.5e-08 $layer=LI1_cond $X=3.237 $Y=3.245
+ $X2=3.237 $Y2=3.33
r156 30 35 12.8291 $w=2.63e-07 $l=2.95e-07 $layer=LI1_cond $X=3.237 $Y=3.245
+ $X2=3.237 $Y2=2.95
r157 29 49 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.505 $Y=3.33
+ $X2=2.375 $Y2=3.33
r158 28 80 7.34436 $w=1.7e-07 $l=1.32e-07 $layer=LI1_cond $X=3.105 $Y=3.33
+ $X2=3.237 $Y2=3.33
r159 28 29 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=3.105 $Y=3.33
+ $X2=2.505 $Y2=3.33
r160 24 27 39.6706 $w=2.58e-07 $l=8.95e-07 $layer=LI1_cond $X=2.375 $Y=2.055
+ $X2=2.375 $Y2=2.95
r161 22 49 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=2.375 $Y=3.245
+ $X2=2.375 $Y2=3.33
r162 22 27 13.0758 $w=2.58e-07 $l=2.95e-07 $layer=LI1_cond $X=2.375 $Y=3.245
+ $X2=2.375 $Y2=2.95
r163 18 21 36.9209 $w=2.68e-07 $l=8.65e-07 $layer=LI1_cond $X=0.59 $Y=2.085
+ $X2=0.59 $Y2=2.95
r164 16 77 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.59 $Y=3.245
+ $X2=0.59 $Y2=3.33
r165 16 21 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.59 $Y=3.245
+ $X2=0.59 $Y2=2.95
r166 5 47 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=4.82
+ $Y=1.835 $X2=4.96 $Y2=2.95
r167 5 44 400 $w=1.7e-07 $l=2.81425e-07 $layer=licon1_PDIFF $count=1 $X=4.82
+ $Y=1.835 $X2=4.96 $Y2=2.055
r168 4 41 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=3.96
+ $Y=1.835 $X2=4.1 $Y2=2.95
r169 4 38 400 $w=1.7e-07 $l=2.81425e-07 $layer=licon1_PDIFF $count=1 $X=3.96
+ $Y=1.835 $X2=4.1 $Y2=2.055
r170 3 35 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=3.1
+ $Y=1.835 $X2=3.24 $Y2=2.95
r171 3 32 400 $w=1.7e-07 $l=2.81425e-07 $layer=licon1_PDIFF $count=1 $X=3.1
+ $Y=1.835 $X2=3.24 $Y2=2.055
r172 2 27 400 $w=1.7e-07 $l=1.18293e-06 $layer=licon1_PDIFF $count=1 $X=2.24
+ $Y=1.835 $X2=2.38 $Y2=2.95
r173 2 24 400 $w=1.7e-07 $l=2.81425e-07 $layer=licon1_PDIFF $count=1 $X=2.24
+ $Y=1.835 $X2=2.38 $Y2=2.055
r174 1 21 400 $w=1.7e-07 $l=1.17584e-06 $layer=licon1_PDIFF $count=1 $X=0.495
+ $Y=1.835 $X2=0.62 $Y2=2.95
r175 1 18 400 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_PDIFF $count=1 $X=0.495
+ $Y=1.835 $X2=0.62 $Y2=2.085
.ends

.subckt PM_SKY130_FD_SC_LP__EINVP_8%A_365_367# 1 2 3 4 5 6 7 8 9 30 34 35 38 42
+ 46 50 54 58 61 63 64 68 72 76 80 84 88 90 92 94 95 96 99 100 101
c162 58 0 1.49947e-19 $X=5.26 $Y=1.635
c163 50 0 4.0679e-20 $X=4.395 $Y=1.635
c164 34 0 4.0679e-20 $X=2.675 $Y=1.635
c165 30 0 9.60268e-20 $X=1.95 $Y=1.98
r166 90 103 2.74877 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=8.85 $Y=2.905
+ $X2=8.85 $Y2=2.99
r167 90 92 36.759 $w=2.88e-07 $l=9.25e-07 $layer=LI1_cond $X=8.85 $Y=2.905
+ $X2=8.85 $Y2=1.98
r168 89 101 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.135 $Y=2.99
+ $X2=7.97 $Y2=2.99
r169 88 103 4.68908 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=8.705 $Y=2.99
+ $X2=8.85 $Y2=2.99
r170 88 89 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=8.705 $Y=2.99
+ $X2=8.135 $Y2=2.99
r171 84 87 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=7.97 $Y=2.19
+ $X2=7.97 $Y2=2.9
r172 82 101 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.97 $Y=2.905
+ $X2=7.97 $Y2=2.99
r173 82 87 0.174613 $w=3.28e-07 $l=5e-09 $layer=LI1_cond $X=7.97 $Y=2.905
+ $X2=7.97 $Y2=2.9
r174 81 100 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.275 $Y=2.99
+ $X2=7.11 $Y2=2.99
r175 80 101 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.805 $Y=2.99
+ $X2=7.97 $Y2=2.99
r176 80 81 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=7.805 $Y=2.99
+ $X2=7.275 $Y2=2.99
r177 76 79 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=7.11 $Y=2.19
+ $X2=7.11 $Y2=2.9
r178 74 100 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.11 $Y=2.905
+ $X2=7.11 $Y2=2.99
r179 74 79 0.174613 $w=3.28e-07 $l=5e-09 $layer=LI1_cond $X=7.11 $Y=2.905
+ $X2=7.11 $Y2=2.9
r180 73 99 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.415 $Y=2.99
+ $X2=6.25 $Y2=2.99
r181 72 100 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.945 $Y=2.99
+ $X2=7.11 $Y2=2.99
r182 72 73 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=6.945 $Y=2.99
+ $X2=6.415 $Y2=2.99
r183 68 71 24.795 $w=3.28e-07 $l=7.1e-07 $layer=LI1_cond $X=6.25 $Y=2.19
+ $X2=6.25 $Y2=2.9
r184 66 99 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.25 $Y=2.905
+ $X2=6.25 $Y2=2.99
r185 66 71 0.174613 $w=3.28e-07 $l=5e-09 $layer=LI1_cond $X=6.25 $Y=2.905
+ $X2=6.25 $Y2=2.9
r186 65 98 4.31308 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=5.515 $Y=2.99
+ $X2=5.387 $Y2=2.99
r187 64 99 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.085 $Y=2.99
+ $X2=6.25 $Y2=2.99
r188 64 65 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=6.085 $Y=2.99
+ $X2=5.515 $Y2=2.99
r189 61 98 2.86415 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=5.387 $Y=2.905
+ $X2=5.387 $Y2=2.99
r190 61 63 41.8043 $w=2.53e-07 $l=9.25e-07 $layer=LI1_cond $X=5.387 $Y=2.905
+ $X2=5.387 $Y2=1.98
r191 60 63 11.7504 $w=2.53e-07 $l=2.6e-07 $layer=LI1_cond $X=5.387 $Y=1.72
+ $X2=5.387 $Y2=1.98
r192 59 96 7.34436 $w=1.7e-07 $l=1.33e-07 $layer=LI1_cond $X=4.66 $Y=1.635
+ $X2=4.527 $Y2=1.635
r193 58 60 7.17723 $w=1.7e-07 $l=1.64085e-07 $layer=LI1_cond $X=5.26 $Y=1.635
+ $X2=5.387 $Y2=1.72
r194 58 59 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=5.26 $Y=1.635
+ $X2=4.66 $Y2=1.635
r195 54 56 40.4442 $w=2.63e-07 $l=9.3e-07 $layer=LI1_cond $X=4.527 $Y=1.98
+ $X2=4.527 $Y2=2.91
r196 52 96 0.195364 $w=2.65e-07 $l=8.5e-08 $layer=LI1_cond $X=4.527 $Y=1.72
+ $X2=4.527 $Y2=1.635
r197 52 54 11.307 $w=2.63e-07 $l=2.6e-07 $layer=LI1_cond $X=4.527 $Y=1.72
+ $X2=4.527 $Y2=1.98
r198 51 95 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.8 $Y=1.635
+ $X2=3.67 $Y2=1.635
r199 50 96 7.34436 $w=1.7e-07 $l=1.32e-07 $layer=LI1_cond $X=4.395 $Y=1.635
+ $X2=4.527 $Y2=1.635
r200 50 51 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=4.395 $Y=1.635
+ $X2=3.8 $Y2=1.635
r201 46 48 41.222 $w=2.58e-07 $l=9.3e-07 $layer=LI1_cond $X=3.67 $Y=1.98
+ $X2=3.67 $Y2=2.91
r202 44 95 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=3.67 $Y=1.72
+ $X2=3.67 $Y2=1.635
r203 44 46 11.5244 $w=2.58e-07 $l=2.6e-07 $layer=LI1_cond $X=3.67 $Y=1.72
+ $X2=3.67 $Y2=1.98
r204 43 94 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.935 $Y=1.635
+ $X2=2.805 $Y2=1.635
r205 42 95 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.54 $Y=1.635
+ $X2=3.67 $Y2=1.635
r206 42 43 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=3.54 $Y=1.635
+ $X2=2.935 $Y2=1.635
r207 38 40 41.222 $w=2.58e-07 $l=9.3e-07 $layer=LI1_cond $X=2.805 $Y=1.98
+ $X2=2.805 $Y2=2.91
r208 36 94 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=2.805 $Y=1.72
+ $X2=2.805 $Y2=1.635
r209 36 38 11.5244 $w=2.58e-07 $l=2.6e-07 $layer=LI1_cond $X=2.805 $Y=1.72
+ $X2=2.805 $Y2=1.98
r210 34 94 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.675 $Y=1.635
+ $X2=2.805 $Y2=1.635
r211 34 35 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=2.675 $Y=1.635
+ $X2=2.075 $Y2=1.635
r212 30 32 36.9577 $w=2.88e-07 $l=9.3e-07 $layer=LI1_cond $X=1.93 $Y=1.98
+ $X2=1.93 $Y2=2.91
r213 28 35 7.43784 $w=1.7e-07 $l=1.8262e-07 $layer=LI1_cond $X=1.93 $Y=1.72
+ $X2=2.075 $Y2=1.635
r214 28 30 10.3322 $w=2.88e-07 $l=2.6e-07 $layer=LI1_cond $X=1.93 $Y=1.72
+ $X2=1.93 $Y2=1.98
r215 9 103 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=8.69
+ $Y=1.835 $X2=8.83 $Y2=2.91
r216 9 92 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=8.69
+ $Y=1.835 $X2=8.83 $Y2=1.98
r217 8 87 400 $w=1.7e-07 $l=1.13284e-06 $layer=licon1_PDIFF $count=1 $X=7.83
+ $Y=1.835 $X2=7.97 $Y2=2.9
r218 8 84 400 $w=1.7e-07 $l=4.19196e-07 $layer=licon1_PDIFF $count=1 $X=7.83
+ $Y=1.835 $X2=7.97 $Y2=2.19
r219 7 79 400 $w=1.7e-07 $l=1.13284e-06 $layer=licon1_PDIFF $count=1 $X=6.97
+ $Y=1.835 $X2=7.11 $Y2=2.9
r220 7 76 400 $w=1.7e-07 $l=4.19196e-07 $layer=licon1_PDIFF $count=1 $X=6.97
+ $Y=1.835 $X2=7.11 $Y2=2.19
r221 6 71 400 $w=1.7e-07 $l=1.13284e-06 $layer=licon1_PDIFF $count=1 $X=6.11
+ $Y=1.835 $X2=6.25 $Y2=2.9
r222 6 68 400 $w=1.7e-07 $l=4.19196e-07 $layer=licon1_PDIFF $count=1 $X=6.11
+ $Y=1.835 $X2=6.25 $Y2=2.19
r223 5 98 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=5.25
+ $Y=1.835 $X2=5.39 $Y2=2.91
r224 5 63 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=5.25
+ $Y=1.835 $X2=5.39 $Y2=1.98
r225 4 56 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=4.39
+ $Y=1.835 $X2=4.53 $Y2=2.91
r226 4 54 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=4.39
+ $Y=1.835 $X2=4.53 $Y2=1.98
r227 3 48 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=3.53
+ $Y=1.835 $X2=3.67 $Y2=2.91
r228 3 46 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=3.53
+ $Y=1.835 $X2=3.67 $Y2=1.98
r229 2 40 400 $w=1.7e-07 $l=1.14286e-06 $layer=licon1_PDIFF $count=1 $X=2.67
+ $Y=1.835 $X2=2.81 $Y2=2.91
r230 2 38 400 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=1 $X=2.67
+ $Y=1.835 $X2=2.81 $Y2=1.98
r231 1 32 400 $w=1.7e-07 $l=1.13578e-06 $layer=licon1_PDIFF $count=1 $X=1.825
+ $Y=1.835 $X2=1.95 $Y2=2.91
r232 1 30 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=1.825
+ $Y=1.835 $X2=1.95 $Y2=1.98
.ends

.subckt PM_SKY130_FD_SC_LP__EINVP_8%Z 1 2 3 4 5 6 7 8 27 29 33 37 39 43 45 47 50
+ 53 57 60 63 64 70 71 72 73 74 78
c111 73 0 2.24865e-20 $X=6 $Y=0.925
c112 60 0 5.29075e-20 $X=5.905 $Y=1.85
c113 47 0 7.73427e-20 $X=8.155 $Y=1.09
r114 73 78 2.96797 $w=3.7e-07 $l=1.35e-07 $layer=LI1_cond $X=5.94 $Y=0.86
+ $X2=5.94 $Y2=0.995
r115 73 74 9.1261 $w=3.68e-07 $l=2.93e-07 $layer=LI1_cond $X=5.94 $Y=1.002
+ $X2=5.94 $Y2=1.295
r116 73 78 0.21803 $w=3.68e-07 $l=7e-09 $layer=LI1_cond $X=5.94 $Y=1.002
+ $X2=5.94 $Y2=0.995
r117 67 68 9.21954 $w=2.48e-07 $l=2e-07 $layer=LI1_cond $X=7.54 $Y=0.89 $X2=7.54
+ $Y2=1.09
r118 64 67 1.38293 $w=2.48e-07 $l=3e-08 $layer=LI1_cond $X=7.54 $Y=0.86 $X2=7.54
+ $Y2=0.89
r119 61 74 7.16384 $w=3.68e-07 $l=2.3e-07 $layer=LI1_cond $X=5.94 $Y=1.525
+ $X2=5.94 $Y2=1.295
r120 60 62 4.83957 $w=4.38e-07 $l=8.5e-08 $layer=LI1_cond $X=5.905 $Y=1.85
+ $X2=5.905 $Y2=1.935
r121 60 61 8.83771 $w=4.38e-07 $l=3.25e-07 $layer=LI1_cond $X=5.905 $Y=1.85
+ $X2=5.905 $Y2=1.525
r122 55 71 3.12539 $w=3.02e-07 $l=1.25499e-07 $layer=LI1_cond $X=8.447 $Y=1.005
+ $X2=8.357 $Y2=1.09
r123 55 57 11.5244 $w=2.23e-07 $l=2.25e-07 $layer=LI1_cond $X=8.447 $Y=1.005
+ $X2=8.447 $Y2=0.78
r124 51 72 3.10218 $w=3.05e-07 $l=1.16619e-07 $layer=LI1_cond $X=8.42 $Y=1.935
+ $X2=8.345 $Y2=1.85
r125 51 53 2.25478 $w=2.28e-07 $l=4.5e-08 $layer=LI1_cond $X=8.42 $Y=1.935
+ $X2=8.42 $Y2=1.98
r126 50 72 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=8.345 $Y=1.765
+ $X2=8.345 $Y2=1.85
r127 49 71 3.12539 $w=3.02e-07 $l=9.0802e-08 $layer=LI1_cond $X=8.345 $Y=1.175
+ $X2=8.357 $Y2=1.09
r128 49 50 17.8932 $w=3.78e-07 $l=5.9e-07 $layer=LI1_cond $X=8.345 $Y=1.175
+ $X2=8.345 $Y2=1.765
r129 48 68 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.665 $Y=1.09
+ $X2=7.54 $Y2=1.09
r130 47 71 3.47949 $w=1.7e-07 $l=2.02e-07 $layer=LI1_cond $X=8.155 $Y=1.09
+ $X2=8.357 $Y2=1.09
r131 47 48 31.9679 $w=1.68e-07 $l=4.9e-07 $layer=LI1_cond $X=8.155 $Y=1.09
+ $X2=7.665 $Y2=1.09
r132 46 70 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=7.635 $Y=1.85
+ $X2=7.54 $Y2=1.85
r133 45 72 3.51065 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=8.155 $Y=1.85
+ $X2=8.345 $Y2=1.85
r134 45 46 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=8.155 $Y=1.85
+ $X2=7.635 $Y2=1.85
r135 41 70 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=7.54 $Y=1.935
+ $X2=7.54 $Y2=1.85
r136 41 43 2.62679 $w=1.88e-07 $l=4.5e-08 $layer=LI1_cond $X=7.54 $Y=1.935
+ $X2=7.54 $Y2=1.98
r137 40 63 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=6.775 $Y=1.85
+ $X2=6.68 $Y2=1.85
r138 39 70 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=7.445 $Y=1.85
+ $X2=7.54 $Y2=1.85
r139 39 40 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=7.445 $Y=1.85
+ $X2=6.775 $Y2=1.85
r140 35 63 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=6.68 $Y=1.935
+ $X2=6.68 $Y2=1.85
r141 35 37 2.62679 $w=1.88e-07 $l=4.5e-08 $layer=LI1_cond $X=6.68 $Y=1.935
+ $X2=6.68 $Y2=1.98
r142 34 60 6.36164 $w=1.7e-07 $l=2.2e-07 $layer=LI1_cond $X=6.125 $Y=1.85
+ $X2=5.905 $Y2=1.85
r143 33 63 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=6.585 $Y=1.85
+ $X2=6.68 $Y2=1.85
r144 33 34 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=6.585 $Y=1.85
+ $X2=6.125 $Y2=1.85
r145 30 73 4.06722 $w=2.7e-07 $l=1.85e-07 $layer=LI1_cond $X=6.125 $Y=0.86
+ $X2=5.94 $Y2=0.86
r146 30 32 24.9696 $w=2.68e-07 $l=5.85e-07 $layer=LI1_cond $X=6.125 $Y=0.86
+ $X2=6.71 $Y2=0.86
r147 29 64 0.241616 $w=2.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.415 $Y=0.86
+ $X2=7.54 $Y2=0.86
r148 29 32 30.0916 $w=2.68e-07 $l=7.05e-07 $layer=LI1_cond $X=7.415 $Y=0.86
+ $X2=6.71 $Y2=0.86
r149 27 62 2.25478 $w=2.28e-07 $l=4.5e-08 $layer=LI1_cond $X=5.8 $Y=1.98 $X2=5.8
+ $Y2=1.935
r150 8 53 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=8.26
+ $Y=1.835 $X2=8.4 $Y2=1.98
r151 7 43 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=7.4
+ $Y=1.835 $X2=7.54 $Y2=1.98
r152 6 37 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=6.54
+ $Y=1.835 $X2=6.68 $Y2=1.98
r153 5 27 300 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_PDIFF $count=2 $X=5.68
+ $Y=1.835 $X2=5.82 $Y2=1.98
r154 4 57 182 $w=1.7e-07 $l=6.11003e-07 $layer=licon1_NDIFF $count=1 $X=8.29
+ $Y=0.235 $X2=8.43 $Y2=0.78
r155 3 67 182 $w=1.7e-07 $l=7.21613e-07 $layer=licon1_NDIFF $count=1 $X=7.43
+ $Y=0.235 $X2=7.57 $Y2=0.89
r156 2 32 182 $w=1.7e-07 $l=6.96491e-07 $layer=licon1_NDIFF $count=1 $X=6.57
+ $Y=0.235 $X2=6.71 $Y2=0.865
r157 1 73 182 $w=1.7e-07 $l=7.21613e-07 $layer=licon1_NDIFF $count=1 $X=5.71
+ $Y=0.235 $X2=5.85 $Y2=0.89
.ends

.subckt PM_SKY130_FD_SC_LP__EINVP_8%VGND 1 2 3 4 5 18 22 24 28 32 36 38 39 40 42
+ 54 59 66 67 70 73 76 79
r109 79 80 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=5.04 $Y=0
+ $X2=5.04 $Y2=0
r110 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.08 $Y=0 $X2=4.08
+ $Y2=0
r111 73 74 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.12 $Y=0 $X2=3.12
+ $Y2=0
r112 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=0 $X2=0.72
+ $Y2=0
r113 67 80 1.07034 $w=4.9e-07 $l=3.84e-06 $layer=MET1_cond $X=8.88 $Y=0 $X2=5.04
+ $Y2=0
r114 66 67 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=8.88 $Y=0
+ $X2=8.88 $Y2=0
r115 64 79 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=5.085 $Y=0 $X2=4.97
+ $Y2=0
r116 64 66 247.588 $w=1.68e-07 $l=3.795e-06 $layer=LI1_cond $X=5.085 $Y=0
+ $X2=8.88 $Y2=0
r117 60 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.295 $Y=0 $X2=4.13
+ $Y2=0
r118 60 62 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=4.295 $Y=0
+ $X2=4.56 $Y2=0
r119 59 79 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=4.855 $Y=0 $X2=4.97
+ $Y2=0
r120 59 62 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=4.855 $Y=0 $X2=4.56
+ $Y2=0
r121 58 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=4.08
+ $Y2=0
r122 58 74 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=3.6 $Y=0 $X2=3.12
+ $Y2=0
r123 57 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=0 $X2=3.6
+ $Y2=0
r124 55 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.435 $Y=0 $X2=3.27
+ $Y2=0
r125 55 57 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=3.435 $Y=0 $X2=3.6
+ $Y2=0
r126 54 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.965 $Y=0 $X2=4.13
+ $Y2=0
r127 54 57 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=3.965 $Y=0 $X2=3.6
+ $Y2=0
r128 53 74 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=2.16 $Y=0 $X2=3.12
+ $Y2=0
r129 52 53 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.16 $Y=0 $X2=2.16
+ $Y2=0
r130 50 53 0.267585 $w=4.9e-07 $l=9.6e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r131 50 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=1.2 $Y=0 $X2=0.72
+ $Y2=0
r132 49 52 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=1.2 $Y=0 $X2=2.16
+ $Y2=0
r133 49 50 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.2 $Y=0 $X2=1.2
+ $Y2=0
r134 47 70 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=0.855 $Y=0 $X2=0.705
+ $Y2=0
r135 47 49 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.855 $Y=0 $X2=1.2
+ $Y2=0
r136 45 71 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=0.24 $Y=0 $X2=0.72
+ $Y2=0
r137 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.24 $Y=0 $X2=0.24
+ $Y2=0
r138 42 70 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=0.555 $Y=0 $X2=0.705
+ $Y2=0
r139 42 44 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.555 $Y=0
+ $X2=0.24 $Y2=0
r140 40 80 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=5.04
+ $Y2=0
r141 40 77 0.133793 $w=4.9e-07 $l=4.8e-07 $layer=MET1_cond $X=4.56 $Y=0 $X2=4.08
+ $Y2=0
r142 40 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.56 $Y=0 $X2=4.56
+ $Y2=0
r143 38 52 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=2.245 $Y=0 $X2=2.16
+ $Y2=0
r144 38 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.245 $Y=0 $X2=2.41
+ $Y2=0
r145 34 79 0.280307 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.97 $Y=0.085
+ $X2=4.97 $Y2=0
r146 34 36 13.7792 $w=2.28e-07 $l=2.75e-07 $layer=LI1_cond $X=4.97 $Y=0.085
+ $X2=4.97 $Y2=0.36
r147 30 76 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.13 $Y=0.085
+ $X2=4.13 $Y2=0
r148 30 32 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=4.13 $Y=0.085
+ $X2=4.13 $Y2=0.38
r149 26 73 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.27 $Y=0.085
+ $X2=3.27 $Y2=0
r150 26 28 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=3.27 $Y=0.085
+ $X2=3.27 $Y2=0.38
r151 25 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.575 $Y=0 $X2=2.41
+ $Y2=0
r152 24 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.105 $Y=0 $X2=3.27
+ $Y2=0
r153 24 25 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=3.105 $Y=0
+ $X2=2.575 $Y2=0
r154 20 39 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.41 $Y=0.085
+ $X2=2.41 $Y2=0
r155 20 22 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.41 $Y=0.085
+ $X2=2.41 $Y2=0.38
r156 16 70 0.597483 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.705 $Y=0.085
+ $X2=0.705 $Y2=0
r157 16 18 15.558 $w=2.98e-07 $l=4.05e-07 $layer=LI1_cond $X=0.705 $Y=0.085
+ $X2=0.705 $Y2=0.49
r158 5 36 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=4.85
+ $Y=0.235 $X2=4.99 $Y2=0.36
r159 4 32 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.99
+ $Y=0.235 $X2=4.13 $Y2=0.38
r160 3 28 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=3.13
+ $Y=0.235 $X2=3.27 $Y2=0.38
r161 2 22 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=2.27
+ $Y=0.235 $X2=2.41 $Y2=0.38
r162 1 18 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=0.575
+ $Y=0.345 $X2=0.72 $Y2=0.49
.ends

.subckt PM_SKY130_FD_SC_LP__EINVP_8%A_371_47# 1 2 3 4 5 6 7 8 9 30 32 33 36 38
+ 42 44 48 50 52 53 54 60 64 65 66 69 76
c139 50 0 8.34392e-20 $X=5.255 $Y=1.295
c140 32 0 3.96626e-20 $X=2.745 $Y=1.295
r141 72 73 1.74613 $w=3.28e-07 $l=5e-08 $layer=LI1_cond $X=8 $Y=0.365 $X2=8
+ $Y2=0.415
r142 69 72 0.174613 $w=3.28e-07 $l=5e-09 $layer=LI1_cond $X=8 $Y=0.36 $X2=8
+ $Y2=0.365
r143 61 69 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.165 $Y=0.36 $X2=8
+ $Y2=0.36
r144 60 76 4.73791 $w=1.7e-07 $l=1.47e-07 $layer=LI1_cond $X=8.73 $Y=0.36
+ $X2=8.877 $Y2=0.36
r145 60 61 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=8.73 $Y=0.36
+ $X2=8.165 $Y2=0.36
r146 57 59 35.3965 $w=2.78e-07 $l=8.6e-07 $layer=LI1_cond $X=6.28 $Y=0.415
+ $X2=7.14 $Y2=0.415
r147 55 68 3.71993 $w=2.8e-07 $l=1.65e-07 $layer=LI1_cond $X=5.585 $Y=0.415
+ $X2=5.42 $Y2=0.415
r148 55 57 28.6053 $w=2.78e-07 $l=6.95e-07 $layer=LI1_cond $X=5.585 $Y=0.415
+ $X2=6.28 $Y2=0.415
r149 54 73 1.70047 $w=2.8e-07 $l=1.65e-07 $layer=LI1_cond $X=7.835 $Y=0.415
+ $X2=8 $Y2=0.415
r150 54 59 28.6053 $w=2.78e-07 $l=6.95e-07 $layer=LI1_cond $X=7.835 $Y=0.415
+ $X2=7.14 $Y2=0.415
r151 52 68 3.1563 $w=3.3e-07 $l=1.4e-07 $layer=LI1_cond $X=5.42 $Y=0.555
+ $X2=5.42 $Y2=0.415
r152 52 53 22.8742 $w=3.28e-07 $l=6.55e-07 $layer=LI1_cond $X=5.42 $Y=0.555
+ $X2=5.42 $Y2=1.21
r153 51 66 6.36606 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=4.685 $Y=1.295
+ $X2=4.575 $Y2=1.295
r154 50 53 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.255 $Y=1.295
+ $X2=5.42 $Y2=1.21
r155 50 51 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=5.255 $Y=1.295
+ $X2=4.685 $Y2=1.295
r156 46 66 0.432806 $w=2.2e-07 $l=8.5e-08 $layer=LI1_cond $X=4.575 $Y=1.21
+ $X2=4.575 $Y2=1.295
r157 46 48 41.3832 $w=2.18e-07 $l=7.9e-07 $layer=LI1_cond $X=4.575 $Y=1.21
+ $X2=4.575 $Y2=0.42
r158 45 65 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=3.795 $Y=1.295
+ $X2=3.7 $Y2=1.295
r159 44 66 6.36606 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=4.465 $Y=1.295
+ $X2=4.575 $Y2=1.295
r160 44 45 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.465 $Y=1.295
+ $X2=3.795 $Y2=1.295
r161 40 65 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=3.7 $Y=1.21 $X2=3.7
+ $Y2=1.295
r162 40 42 46.1148 $w=1.88e-07 $l=7.9e-07 $layer=LI1_cond $X=3.7 $Y=1.21 $X2=3.7
+ $Y2=0.42
r163 39 64 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.935 $Y=1.295
+ $X2=2.84 $Y2=1.295
r164 38 65 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=3.605 $Y=1.295
+ $X2=3.7 $Y2=1.295
r165 38 39 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.605 $Y=1.295
+ $X2=2.935 $Y2=1.295
r166 34 64 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=2.84 $Y=1.21
+ $X2=2.84 $Y2=1.295
r167 34 36 46.1148 $w=1.88e-07 $l=7.9e-07 $layer=LI1_cond $X=2.84 $Y=1.21
+ $X2=2.84 $Y2=0.42
r168 32 64 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.745 $Y=1.295
+ $X2=2.84 $Y2=1.295
r169 32 33 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.745 $Y=1.295
+ $X2=2.075 $Y2=1.295
r170 28 33 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=1.945 $Y=1.21
+ $X2=2.075 $Y2=1.295
r171 28 30 35.0165 $w=2.58e-07 $l=7.9e-07 $layer=LI1_cond $X=1.945 $Y=1.21
+ $X2=1.945 $Y2=0.42
r172 9 76 91 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_NDIFF $count=2 $X=8.72
+ $Y=0.235 $X2=8.86 $Y2=0.44
r173 8 72 91 $w=1.7e-07 $l=1.94422e-07 $layer=licon1_NDIFF $count=2 $X=7.86
+ $Y=0.235 $X2=8 $Y2=0.365
r174 7 59 182 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_NDIFF $count=1 $X=7
+ $Y=0.235 $X2=7.14 $Y2=0.44
r175 6 57 182 $w=1.7e-07 $l=2.65942e-07 $layer=licon1_NDIFF $count=1 $X=6.14
+ $Y=0.235 $X2=6.28 $Y2=0.44
r176 5 68 91 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=2 $X=5.28
+ $Y=0.235 $X2=5.42 $Y2=0.38
r177 4 48 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=4.42
+ $Y=0.235 $X2=4.56 $Y2=0.42
r178 3 42 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=3.56
+ $Y=0.235 $X2=3.7 $Y2=0.42
r179 2 36 91 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=2 $X=2.7
+ $Y=0.235 $X2=2.84 $Y2=0.42
r180 1 30 91 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=2 $X=1.855
+ $Y=0.235 $X2=1.98 $Y2=0.42
.ends

